MZP      ��  �       @                                     � �	�!�L�!��This program must be run under Win32
$7                                                                                                                                        PE  L ^B*        � �� �   :      d�      �    @                      p               @                          	   P                     0 �                                                                                CODE    ��      �                    `DATA    �   �      �              @  �BSS     �   �       �                 �.idata  	      
   �              @  �.tls              �                 �.rdata            �              @  P.reloc  �   0     �              @  P.rsrc       P     �              @  P             p      �              @  P                                                                                                                                                                @ 
StringX@                             X@        �*@ �*@ �*@ �*@ �*@ �)@ �)@  *@ TObjectd@ TObjectX@       System  �@ IUnknown            �      FSystem  �%8A ���%4A ���%0A ���%,A ���%(A ���%$A ���% A ���%A ���%A ���%A ���%A ���%A ���%HA ���%A ���%A ���% A ���%� A ���%� A ���%� A ���%� A ���%� A ���%DA ���%� A ���%� A ���%� A ���%XA ���%TA ���%PA ���%� A ���%� A ���%xA ���%tA ���%pA ���%lA ���%hA ���%dA ���%`A ��S�ļ�
   T�Y����D$,t�\$0�Ã�D[Ë��%� A ���%� A ���%� A ���%� A ���%� A ���%� A ���%� A ���%� A ��SV�L�@ �> u:hD  j �����ȅ�u3�^[áH�@ ��H�@ 3ҋ���D����B��du���^[Ð� �@Ë�SV���������u3�^[Ë�P�V�P���X�B��^[ËP��
�Q�L�@ ��L�@ �SVWUQ��$��] �$���P�V�;�C��S;u�������C��CF��V;�u�������CF��;�u֋��U�����u3��Z]_^[Í@ SVWU����؋��2�C;�rl��J��k;�w^;�u�BC�B)C�{ uD���5����;�
�r΋�{;�u)s�&�
J�$+��|$�+ЉS�ԋ��������u3�����;�u�3�YZ]_^[ÐSVW�ڋ���   }�   �����  ��  ���sjh    Vj ��������;��t#�ӸP�@ �l�����uh �  j �P�����3��_^[ÐSVWU�ً���C   jh    h   U�������;��u����  ��  ���sjh    VU������; t#�ӸP�@ �������uh �  j �P�b���3��]_^[ÐSVWU���L$�$�D$����3҉T$��$ŉD$�P�@ �Q�;�s;�wF��C;D$w;;t$s�t$��C;D$v�D$h �  j V�������u
�,�@    �������߁�P�@ u��D$3҉�|$ t�D$�T$��D$+D$�T$�B��]_^[�SVWU���L$�$�Ћ�� ���$���  �� ����T$�D$�(�D$+ŋT$�B�5P�@ �<�^�~�;�v��;|$v�|$;�vjh   +�WS�&�����u
�D$3҉�
�6��P�@ u���]_^[Ë�SVWUQ�؋���  �� ����4$���� ����$���+$�A�5P�@ �8�^�~�;$s�$;�s��;�vh @  +�WS������u
�,�@    �6��P�@ u�Z]_^[Í@ SVWU�������`�@ ���?  �� ����] �3;{,�΋׋C�����> tP�FC�F)C�{ u>��������5�;�uɋ֋�������> t!�̋֋�������<$ u��̋V�����3��YZ]_^[Ë�SVWU���$����`�@ ���?  �� ����] ��;�t;su�;suW;{��   �L$��+S�CC������|$ t3�L$�T$���]����|$ u��L$�T$�D$�%����$3҉�   �L$�׋������|$ t4�L$�T$�������|$ �f����L$�T$�D$������$3҉�H�k;�u:;{5�$�׋��q����$�8 t(�$�@C�$�@)C�{ u��������$3҉��]_^[ÐSVW�����$���?  �� ����4$��� ���;�s[�ϋ�+Ӌ������L$�׸`�@ �]����\$��t�L$�T$���&����D$�D$�D$�D$�|$ t�T$�`�@ �����3����_^[�U��3�Uhz@ d�2d�"h0�@ �9����=A�@  t
h0�@ �.����P�@ �����`�@ �������@ �x���h�  j ��������@ �=��@  t/�   ���@ 3ɉL��@=  u�p�@ �@� �|�@ �(�@ 3�ZYYd�h�@ �=A�@  t
h0�@ ������  ��(�@ ]�U��S�=(�@  ��   3�Uh^@ d�2d�"�=A�@  t
h0�@ �f����(�@  ���@ P�4���3����@ �P�@ �h �  j �CP�%������P�@ u�P�@ �����`�@ �������@ �u����H�@ ��t��H�@ P������H�@ ��u�3�ZYYd�he@ �=A�@  t
h0�@ �����h0�@ ��������  ��[]�S;|�@ u	�P�|�@ �P�H��   8;�u��y�������@ 3҉T���$��y�������@ �T�� ��P[Ë ��P[Í@ ���@ ��J;�rJ;�r�����@ u��,�@    3ҋ�ÐS�ʃ����|�  ����  [Ã�|�ʁ�  ���[���@ �Ѓ��������� �@ ��  Ë���|����������Ã�|
�ʁ�  �� ��SV�Ѓ���ʁ�  ���  �t
�,�@    �ځ����+Ë�3������t
�,�@    �t �Ѓ��r+�;pt
�,�@    ����ދ�^[Í@ SVW��3���   �t%����؋�u����X����F�؃#���_^[�SVWU��������������؋k��C�Ѝ7+у���+���+Ń�}�̋�+S׋��������̋׃��F������,$��u3��0��+֋��p�����D$�SS;�s
�7+������ԋ������YZ]_^[�SVW����߉s��ƃ��p��   7�օ�y�������@ �D���u���@ �\��[��:��C���Z�,�� <  |�֋�������u�|�@ �|�@ ��C���Z_^[Í@ �=��@  ~@�=��@ }�,�@    �+���@ �����@ ����@ ������3����@ 3����@ Ë�SVW������<$���������L$�׸��@ �(����\$��u3��R�;�s
����)G�G��t$;�s����G�G;�u���   �����o����@ �G���@ ���_^[Í@ S����؋ԍC�\����<$ t���W�����u3���YZ[ÐSV�����؋̍V�������<$ t���&�����u3���YZ^[Í@ 3҅�y����=   ���@ �T���u@=  u���SVWU��|�@ ���@ �t�@ ;s��   ��C;�~{�s�[;s���B;t��c��   �������؅�uN��������u3��   ;u �)u �} }u 3��E ���@ 5��@ �փ������@ ��5 �@ �L�������S��+ƃ�|��֒�T������;u�C���ƃ ��Ëփ������@ ��5 �@ ]_^[�U����SVW�؀=(�@  u������u
3��E��T  3�Uh!@ d�1d�!�=A�@  t
h0�@ �@����������}�   ��   ��   �Å�y�������@ �T���ty���Ã ��B;�u�Å�y�������@ 3��|���&�˅�y�����=��@ �D��
�M��M��A�M���ƋR������E���@ �� �@ �  �   ;��@ J)��@ �=��@ }��@ 3����@ ���@ ��@ �Ӄ�����E���@ �� �@ �1  �2�������E�3�ZYYd�h!@ �=A�@  t
h0�@ ������'  ��E�_^[YY]Í@ U��QSVW��3��,�@ �=(�@  u������u�,�@    �E�   �a  3�Uh�"@ d�1d�!�=A�@  t
h0�@ ����������u�,�@ 	   ��   ��@ ��%�����) �@ ��tE�ƃ��P��|��  �t�,�@ 
   �   ��+�;Pt�,�@ 
   �   ڋ��t����������Ë�;=��@ u,)��@ ��@ �=��@  <  ~����3��E���  �   ���t�������}�,�@    �7��)�ǃx t�8 t�x}�,�@    ��P�������Ӌ��/����,�@ �E�3�ZYYd�h�"@ �=A�@  t
h0�@ �w�����
  ��E�_^[Y]Ë�SVWU�����������}�   ����} �������ǋ�;���   ��+։$;��@ u8�$)��@ �$��@ �=��@ �L  �$��@ �$)��@ ���3  ���u�ËP$�����<$|��ދ$����Ã�������   ����   ��+ǉD$;��@ ug���@ ;D$|S�D$)��@ �D$��@ �=��@ }���@ ��@ 5��@ 3����@ ��+� �@ �E %  ���u ��   �Q�������uM�ӋH�$�$;L$}$�ڋ$)D$�,�J����D$)$�<$|��Ƌ$�����:4$��ރ#��.��   �t!%���Ë؋T$���������t	�������3����+� �@ �E %  ���u �YZ]_^[ÐU��QSVW��؀=(�@  u������u
3��E��   3�UhE%@ d�2d�"�=A�@  t
h0�@ �D����֋��������t�]��6���������Ã�� %�����;�}�ƅ�t�׋ˑ�V  ��������}�3�ZYYd�hL%@ �=A�@  t
h0�@ ��������  ��E�_^[Y]Í@ ��t
��@ 	�tð�j   Ð��t
��@ 	�uð�R   Ð���t2��tP����@ Y	�t�ð�.   �����@ 	�u�ð�   ��tP����@ Y	�t�Í@ ����@ ��tZ��H��&@ y�F.  ��   �k  ��������������������� ��Ë�PRQ�.  ��    YZXu�1�����Í@ P��-  ��   Í@ ����������Ð��-  1ҋ�   ��   ��Ë�VW�Ɖ׉�9�wt/��x*�����_^Ít��|���x�����������_^�SV�����P����C���t< v��;"u�{"u����3��%��"uC��@C���t��"u��; tC��@C��� v=   |͋ԋΑ�A  �Á�   ^[Ë�SVW��������؅�uh  �D$Pj ������ȋԋ��  ���������֋��I�������t�> tK���  _^[Ð�=�@  t��@ ��   ��
  Ë�W�ǈ͉���f�ȉ���x	�у��_ÐSVW��P��ts1�1ۿ����F�� t�� ��-ti��+tf��$tf��xta��Xt\��0u�F��xtO��XtJ��t ���t4��0��	w,9�w(���؊F��u���t��|Y1��2_^[�F���~�x�[)����ŊF뼿����F��t߀�ar�� ��0��	v����wЀ�
9�w���؊F��u����%@A ��S3�j �������uj�����% �  =   t=   u���[ÐU����� �@ �E��E�Pjj hX)@ h  �������uM3�Uh1)@ d�0d� �E�   �E�P�E�Pj j ht)@ �E�P�j���3�ZYYd�h8)@ �E�P�D�����  ��f� �@ f%��f�U�f��?f�f� �@ ��]� SOFTWARE\Borland\Delphi\RTL FPUMaskValue    ���- �@ Ë�VW�׋p�1ɊA�_^Í@ P�@�������X�g   Ë�SV�ÉƋ6�V��v܅�t�I  �؅�u�����^[Í@ ��t����$  ��t�s  d�    ����k  ��~�R  Ð��t���Q��SVW�É׫�K�1�Q��I�Y���Љ�K���tQ�[܅�t���9�t[����s��t�{�48��Iu�9�u�_^[Ë���t� 9�t�@܅�u�ðÍ@ W����{Ѕ�t�Q��f�t
Y�[܅�u�_�X�)ȋ\G�_Ë�PQ� �����YXt��Y����Ë���� �Ë�Í@ Í@ Í@ Sf�f	�tf�� �sP� ����Xt��[��[��a�ÐRQS��|�P�1ҍL$d���i�A9+@ �Ad�
[YZ��*  �D$,�@��t���P�Q�X�	   �0  Í@ ��R�Ë�P��R�XÄ��PR��R�ZXÐ�=�@ vj j j h����;���Ë��=�@  tPPRTjj h���������X�Tjj h����	�����XÀ=�@ vPS�����Í@ ��t�A�9�t�9�u��AA����Ë��=�@ vPRQ�����QTjj h�������YYZXË��=�@ vRTjj h�������ZÐPR�=�@ vTjj h����r���ZXÍ@ �D$�@   ��   �8����P�Ht<��������@ ����   �҅���   �T$�L$�9���t������D$�H�HS1�VWUd�SPRQ�T$(j Ph�,@ R������|$(�M'  ��    ��    �o�_�G-@ ����������!   � '  ��    ���    �A������   ËD$�T$�@   t�J�Bh-@ SVWU�j��������]_^[�   Ë�ZTUWVSPRTjjh���R�L���Í@ �D$0�@�-@ �&  ��    �
��    �B�`��8���t�B�O�������1���d�Y��]_^[�   Í@ �W&  ��    �
��    �B����Z�d$,1�Yd�X]�������1ҋL$�D$��d���� Ë��$�<  Í@ U��U�=�  �,t\=�  �tW-  �t\-�   t=HtN�`q��?��r6t0�R=�  �t=-�  �t.HtHt$�:-�  �t/��=t&�,���*���&���"������������������
��������%�   �R�X���]� �D$�@   ul������T$j Ph�.@ R������\$�;����S�Ct��@ ���������҅������S����� �@ ��t�ыL$��   �Q�$�  1��1ҍE�d�
d���@�.@ �h���@ Ë�1ҋ��@ d�
9�u� d�Ë	���t9u�� �Í@ U��SVW���@ �G��tH�_�p3�Uh�/@ d�2d�"��~K�_�D���t�Ѕ��3�ZYYd�������������������_^[]ÐU��SVW���@ ��tK�03ۋx3�Uh>0@ d�2d�";�~��C���@ ��t��;��3�ZYYd���%����P����?�������_^[]Ð���@ 1����@ ���@ �B��@ ������$�@  �r���ÐSV��p�F�� �1  ��Ku�^[�SV��p�F��N� ȉ��Ku�^[Ë�S�0�@ �,�@ �
   1����0�K��u�8�@ �>  �8�@ �)л8�@ ����D�@ �K��u�[Í@ ���@ ���@ �-��@ �w�w �7�   �_^1��0�@ ���@�� �SVWU���@ �0�@ �4�@ �{$ u�? t���3҉���Ճ? u�=8�@  t>�?����=@�@  t��@ ��@ �;  �  �j h<�@ h�@ j �U���3��8�@ �{$u
�> u3��C������{$v�> t�C��t�r  �C�P;PtR�����p����{$u�S(�{$ t� ����; u�P������V�����   �^�Portions Copyright (c) 1983,97 Borland ]_^[Ë��0�@ �����Ï8�@ �����Ë��t�     �J�I|�J�u
P�B������XË�SV�É֋��t�    �J�I|�J�u�B�������Nu�^[Ë���t#�J�APR�B��X   ��XR�H�����ZX��J����t�J�I|�J�u�B��d���Í@ ��t	�J�A~�J����t�J�I|�J�u�B��:���Ð��~P��	������Z�P��@�   � �1�ÐSVW�É։ω���������ǅ�t	���������������;_^[Ë�SVWU�� ����ً����	��������g��   },j j h   �D$PSUj j ���������~�ԋǋ������3j j j j SUj j �������ǋ�3��_���j j V�PSUj j �|�����   ]_^[ÐR��   �3���ZÐ1Ʌ�t!R:
t:Jt:Jt:Jt����BBB��Z)�����Í@ 1Ʌ�t-Rf;
t f;Jtf;Jtf;Jt�����������Z)��������Í@ 1Ɋ
B����ÐWPQ��1��u��X�X_�����1Ʌ�t�J��������Í@ ��t�@�Å�t?��������SVW�É֋y��V��9�t�N  ���N����d���_^[��7  �����Å�ta�������;t\;tPQ����ZX����SVW�Ӊ�P�C�F�������ǉ؋K����������N�S�����X����t�O��O���_^[É��D������I����SVRP��1��L���tA�Ju�����P�ƋD����t
�H������Ku�ZX��t�J������Z^[X�$���Í@ SVW�Ɖ�9���   ��th��tk�F��W�)�w�R��t&��9�uXJt�N�_9�uK����Ju������Z��t"��8�uAJt8�u:Jt��  � ��  � 9�u'��#�W�)���F�)��Z8�u8�u����8�u8�_^[Ë���t� ��6@ Ë��t+�J�It%S�ËB��������H�I|�H��H������[���S��t-�X���t&J|9�})Ӆ�|9�D$�p����1������D$�y���[� �SVW�É։��~������t0�J�N|*9�}&��~")�9�~��)��:�6�����؋R�)��   _^[�SVW�É�1���tH���t#�x�u����	P������X����p��0 �(�������ǋ��t���H�9�|���������������;_^[Ë���!���Ë��t�     PR�����XÍ@ SV�É֋��t�    P�������Nu�^[Í@ ��������J��������QRP������������1�S�JVW�Ít

�|
��F؋��   ��O��_^[�PSVW�É։�1Ҋ�V��
t1��tF��tX��tb��t{����   ����   _^[X��M�������
������   ��������x���������j�������a�؃��  O��RU�ՋT.
��\.�L.��a���O�]�4U�Չ�\.������O�]��؃��  O���؉���  O�_^[XË��   ����ÐSVWU�É�1��A�|
�o�1��O�Q�O)�~���������G���
��
t1��t=��tI��tU��tp����   ����   �]_^[�=������'����   �}���>����   �l���  �   �[1ɊJ�t
�t
�L

�	���a   X�;1ɊJ�L
Q�э��,���X�"���+  �   ��ы���  �   G��M����Y)�~
���+���]_^[Ë�SVWU�É։ϋl$���
t1��tC��tR��ta��t}����   ����   �]_^[�F����؋�1�������Mu��   �؋�B�������Mu��z�؉��  ����Mu��f1ɊO�|�؉�O�w�c���7Mu��E�؉���3���1��G\tMu��(�؋�$  ����Mu���؋����  ����Mu�]_^[� ÐSVWU�� �����ڋ���u	�������a��   }&j j h   �D$PSWj j �����ȋԋ�������3j j j j SWj j �������Ƌ�3�����j j U�PSWj j �������   ]_^[Í@ SVj ��؉$�$P������Ћ΋��U���Z^[ÐSVWU�� ����؋���������������=   }+h   �D$PV���_���Pj j �=���P�D$P�b������(j j VSj j ������Uj �E�����UWVSj j �����ǁ�   ]_^[Ð��]���ð�U����1�f��� @  u(��r#��   t��  u�%��@ f�   ������f�   �P�����Ë�9���   f�8r*PRf�8 tf�8tP���������@ ����z���ZXf�:s�
��J�H�J�H�f�: tf�:u&P�����X�%��@ �R	�t	�J�A~�J�f�  �P�f�   RP�m���	������U����SVW��}�Q�   �Y��؍E��Y  3�Uh�=@ d�0d� �E����@ �U��Ë��&   3�ZYYd�h�=@ �E��  ��w�����_^[��]Ë�U����SVW�����f�f- tf��t=�Hf�E�  Wj h   V�E�P�������t�h������q����E���E��C�E��C�%�֋Ë��/����Wj h   VS������t�)���_^[��]Ë�U��QS��3��E��B�U��a���������f� �E��C[Y]Í@ SV�؋B�`������������f� �s^[�U����S�E�f���f;�u�E�������   f= uYf��u�E������   f�E�  �E�����3�Uh?@ d�0d� �U��E�������3�ZYYd�h�?@ �E��h����������f�� u^f=tXf��u
�E������Rf�E�  �E�f� �y���3�Uh�?@ d�0d� �U��E������3�ZYYd�h�?@ �E�������������E���9���[��]�f�: u�R�%���S�Ã�f�$  ��   ������������D$���[Í@ P����X�f�8r�p�p�p�0f�   ���������Í@ ��t�@�������HÐU���u�1���]� �����Ë��  Ë�U����SVW�M���E��]���E�8����}��~����E���������H  3��E���t����E���3��FƋF�E�F��t�0�3����m�E�E���;E�t��'����E���t�;u5�]�;}�}��t�Ã����U�M�+ϋ��=����E��U������]��^��E��[����؋E��E�;}�}�}��t*�U��U�Ã�3��x����E�P�U���Ã����������M��M�Ӄ��E�� �����   ���;����+U��U�E��E��3��$����}�~.�E�M�O��|"G�E�    �EP�E���M��������E�Ou�E��_^[��]� ��T�$�j���Ð���t2�     �I�u'P��1ɊJ�T
��t�H���t��M������q���XÍ@ S���t�B���t�K�uPR���C�����ZX�[Í@ ���j�T$RP�X����|$   u�D$�3���Ë���@ ��t;Bt
;Bt;Bu�BË��u��U�������SV�E�h  ������Pj �����E� �E�Ph?  j h0D@ h  ��������t�E�Ph?  j hLD@ h  �������um3�Uh?C@ d�0d� �E�   �E�P�E�Pj j ������P�E�P�z�����t�E�P�E�Pj j hlD@ �E�P�\���3�ZYYd�hFC@ �E�P�6�����������E�P������P����j�E�Pj�����P�����3������� ��   �}� u
�}� ��   ������P������؍�������K�;.t
������;�u�������;�tmC�}� t�E�PS����jj ������P�q�������uF�}� t@�E�PS�k���jj ������P�K�������u �E� �E�PS�G���jj ������P�'�������^[��]� Software\Borland\Locales    Software\Borland\Delphi\Locales     S�ظ   �������@ ��X��@ [ÐSV�5�@ ��t"�V;�u��@ � ��@ �   ������^[Ëօ�t'�
��t�Y;�u����   ����������u�^[Ë�U����SVW�E���@ �E��}� t93�Uh+E@ d�0d� �]��E��S3�ZYYd��
�8��������E�� �E��}� u�_^[YY]Ë���@ ���@ Ë�U��Q�E�3�Uh�E@ d�2d�"�E��@�t���3�ZYYd�h�E@ �E�;�@ u�E�� ��@ ���@ ��t�;U�u	�U����� ��u���s�����Y]Ë�SV�� �����؅�t=�{   }*h   �D$P�CP�� �X���P�R����ȋԋ��O����
�ƋS������   ^[Ë����t�     PR��PXÍ@ ����tQR��PY��tQ��PÐ�%� A ��3҉P�PR�PR�p�p�0�b�����t3��������mt��3��Q�P��~3ɉHQ�L$QR�p�0�O�����t3�Y��j������0�@��  �����Hu��Q����V��3��F�F�F-��  tHt Ht.�I  �   ��   �   �F`F@ �'�   @�   �   ��   ��   �   �F�F@ �F$�F@ �F �F@ �~H ��   j h�   Qj RP�FHP�T��������   ��~��  ��   �Nj �6�@���@��   -�   s3�j j P�6�T���@��   j ��j Rh�   ��L  R�6����ZH��   3�;�sL��L  t@��jj +�P�6�
���@tg�6�����Hu]�"�F$�F@ �~��  tj��j��������t;��~��  t�6������t��u�F �F@ 3�^��6�f����F��  �i   ���F��  ������ۍ�L  �H3ɉ�@��  �@�   �H�H�@�F@ �H�H �H$�@H��t���
B�@��t�
B�@��t��u�H�(ËP����  u�P��uÁ���  t��g   �_����P����  u�P ��uÁ���  t��g   �:�����SV�؋�S���  ��wHQj ��j P�C��PV�3����HXYu3��s�T$��t�^[� ;�t��d   �����������3���g   ��SV�؋�@-��  ��wHQj ��j P�C��PV�3�k���HXYu3��s�T$��t�^[� ;�t��e   ��j����}���3���g   ����S�؋P���  t��w�P��u���S$��u[��F�����=H�@ t�g   ���SV���ڋV���  t
��w�����Ɖ^�V��t����^[øf   ��������  뾺��  뷺��  �SVW�؋���S���  t����   �S$��t�����C��  �s�C$zK@ �CK@ �{H tg�   ��B�@ ��p����9K@ �   ��t#�   Gt�   @G�C��  t�   ��C��  j h�   Qj RP�CHP�������t)�_^[�3���C$K@ ��tj��j������ٸf   ��C��  �����������                            3ɊB�@ ����v�������   ������0�@��  �$���H������VW��x��  u.�xx�P+P;�P+�PQ����P��u3YX��H�_^�=�@ uQRP�p���XZY�x��  t��i   �L������E���YX�͋ʺT�@ ��@~!��@PQ�@   �z����!  ��    uYX�Յ��`����YX�3Ɋ
B�R���S3ۊ+�~PR������ZX��[B�5������@ �   �&����n����x��  u�H;H}	H��@�PR�P��u'ZX��=�@ uRP����XZ�x��  tɸi   �����~���ZX�R�Q��1����Թ   ����Z�3�� VW��Q������ ���I��Z+ы�Q����Y�Ƌ�_^��������|HtE=   �   �Ѓ����,U�M@ ����t$�Ѓ�t���,U�N@ ����t���,ExO@ �����=   }B�Ѓ����,U�M@ ����t��Ѓ�t���,U�N@ ����tȍ��,ExO@ ����-�M@ ����       ��       ��?       �@       �@       �@      @�@      P�@      $�@     ���@      ��@     (k�@     �� @    @�C�#@    ���&@    *焑*@   �� �-@   �1�_�0@   ���4@   �.���7@  @v:k�:@  �#Ǌ>@  b���x�A@ �z�&��D@ ��n2x��H@ �W
?h�K@ ������N@��@aQY�R@ȥ���o�U@: �'���X@�	��x9?�\@��6���_@�Ng����b@�"�E@|o�e@��p+��ŝi@զ��Ix��@������=A����G���A��+��BkU'9��p�|B0�<���R��B������~�QC�/j\�&һCv���)/��&D�
�� '���D�������DY������dE�����Jz��Eb����>�9FǑ����Fu��uv�HM䧓9;5���S�]=�];���Z�� �T��7a�Z��%]���g��'���]݀n�� �R`�%u�Y�nb5��{RP�D$�$$�ȋD$�d$ȋ$�d$�YY� RP�D$�$$�ȋD$�d$ȋ$�d$�YY� USVW3��\$�L$�u�t\�tX�y
���؃� ���y
���ۃ� ����@   W3�3���������;�rw;�r+��@��[��   t���؃� _^[]� ��3���V�t$#t$���u����   �u��^H�^�t$�t$�[���#�� USVW�\$�L$�u�t/�t+��@   3�3���������;�rw;�r+��@��_^[]� ��3���USVW3��\$�L$�u�t]�tY�y
���؃� ���y���ۃ� ��@   W3�3���������;�rw;�r+��@��Ƌ�[��   t���؃� _^[]� ��3���V�t$#t$���u����   �u��^H�^�t$�t$�Y���#�� USVW�\$�L$�u�t3�t/��@   3�3���������;�rw;�r+��@��Ƌ�_^[]� ��3���� |��@|3�3�Ë���3������À� |��@|����Ë�������À� |��@|3�3�Ë�3��������ÐU��3�Uh�R@ d�0d� �$�@ u7�H�@ �E�����@ �;����������@ �4������@ �*������@ � ���3�ZYYd�h�R@ ��q�����]ÐU��3�Uh�S@ d�0d� �-$�@ ��   3��0�@ 3��8�@ 3��<�@ �B�@ �C�@ �D�@ f���@   f���@  f��@ 
 ��@  ����@ |<@ ���@ t<@ ���@ |<@ �4�����t�[��������H�@ ��S@ �������@ ��S@ �����菽���,�@ �=����(�@ ����� �@ 3�ZYYd�h�S@ �������]�       �%�A ���%�A ���%�A ���%�A ���%�A ��S�   ��tC�=��@  }
��   �c���h   j@�����؅�u��   �G����S���@ P�������@ [Ð���@ ���@ ��u(d�,   ����������@ P�t�����tË��@ �P�b�����t�ÐS������h  �D$P���@ P�(�����������؉��@ ��u
���@ ���@ ���@ ������  [ÐPj ��������@ R���@ �B�B    �B    ����ZX�[���Ë�U��3�Uh%U@ d�0d� ���@ 3�ZYYd�h,U@ �������]Ë��-��@ ��%�A ���%�A ���%�A ���%�A ���%�A ���%�A ���%0A ���%,A ���%(A ���%$A ���% A ���%A ���%A ���%A ���%A ���%A ���%A ���%A ���% A ���%�A ���%�A ���%�A ���%�A ���%�A ���%�A ���%�A ���%�A ���%�A ���%�A ���%�A ���%�A ���%�A ���%�A ���%�A ���%�A ���%�A ���%�A ���%�A ���%DA ���%@A ���%<A ���%8A ��U��3�Uh�V@ d�0d� ���@ 3�ZYYd�h�V@ �������]Ë��-��@ ���@ ��  ��@ ��  ��@ ��  ��@ ��  ��@ ��  ��@ ��  ��@ ��  ��@ ��  ��@ ��  ��@ ��  ��@ ��  ��@ ��  ��@ ��  ��@ ��  ��@ ��  ��@ ��  ��@ ��  ��@ ��  ��@ ��  ��@ ��  ��@ ��  ��@ ��  ��@ ��  ��@ ��  ��@ ��  ��@ ��  ��@ ��  ��@ ��  ��@ ��  ��@ ��  ��@ ��  ��@ ��  ��@ ��  ��@ ��  ��@ ��  ��@ ��  ��@ ��  ��@ ��  ��@ ��  ��@ ��  ��@ ��  ��@ ��  ��@ ��  ��@ ��  ��@ ��  ��@ ��  ��@ ��  ��@ ��  ��@ ��  ��@ ��  ��@ ��  ��@ ��  ��@ ��  ��@ ��  ��@ ��  ��@ ��  ��@ ��  ��@ ��  ��@ ��  ��@ ��  ��@ ��  ��@ ��  ��@ ��  ��@ ��  ��@ ��  ��@ ��  ��@ ��  ��@ ��  ��@ ��  ��@ ��  ��@ ��  ��@ ��  ��@ ��  ��@ ��  ��@ ��  ��@ ��  ��@ ��  ��@ ��  ��@ ��  ��@ ��  U��3�UheY@ d�0d� ���@ 3�ZYYd�hlY@ ��������]Ë��-��@ ��Y@         �Y@                 �Y@    @ �*@ �*@ �*@ �*@ �*@ �)@ �)@  *@          @    	Exception,Z@                             ,Z@    xY@ �*@ �*@ �*@ �*@ �*@ �)@  u@  *@ EHeapException��Z@                             �Z@    �Y@ �*@ �*@ �*@ �*@ �*@ �)@  u@  *@ EOutOfMemory�@ �Z@                             �Z@    xY@ �*@ �*@ �*@ �*@ �*@ �)@ �)@  *@ EInOutError<[@                             <[@    xY@ �*@ �*@ �*@ �*@ �*@ �)@ �)@  *@ 	EExternal���[@                             �[@    �Z@ �*@ �*@ �*@ �*@ �*@ �)@ �)@  *@ EExternalException��[@                             �[@    �Z@ �*@ �*@ �*@ �*@ �*@ �)@ �)@  *@ 	EIntError��L\@                             L\@    �[@ �*@ �*@ �*@ �*@ �*@ �)@ �)@  *@ 
EDivByZero��\@                             �\@    �[@ �*@ �*@ �*@ �*@ �*@ �)@ �)@  *@ ERangeError�\@                             �\@    �[@ �*@ �*@ �*@ �*@ �*@ �)@ �)@  *@ EIntOverflow�@ X]@                             X]@    �Z@ �*@ �*@ �*@ �*@ �*@ �)@ �)@  *@ 
EMathError��]@                             �]@    ]@ �*@ �*@ �*@ �*@ �*@ �)@ �)@  *@ 
EInvalidOp�^@                             ^@    ]@ �*@ �*@ �*@ �*@ �*@ �)@ �)@  *@ EZeroDivide`^@                             `^@    ]@ �*@ �*@ �*@ �*@ �*@ �)@ �)@  *@ 	EOverflow���^@                             �^@    ]@ �*@ �*@ �*@ �*@ �*@ �)@ �)@  *@ 
EUnderflow�_@                             _@    �Y@ �*@ �*@ �*@ �*@ �*@ �)@  u@  *@ EInvalidPointerl_@                             l_@    xY@ �*@ �*@ �*@ �*@ �*@ �)@ �)@  *@ EInvalidCast�@ �_@                             �_@    xY@ �*@ �*@ �*@ �*@ �*@ �)@ �)@  *@ EConvertError��$`@                             $`@    �Z@ �*@ �*@ �*@ �*@ �*@ �)@ �)@  *@ EAccessViolation�@ �`@                             �`@    �Z@ �*@ �*@ �*@ �*@ �*@ �)@ �)@  *@ 
EPrivilege��`@                             �`@    �Z@ �*@ �*@ �*@ �*@ �*@ �)@ �)@  *@ EStackOverflow�8a@                             8a@    �Z@ �*@ �*@ �*@ �*@ �*@ �)@ �)@  *@ 	EControlC���a@                             �a@    xY@ �*@ �*@ �*@ �*@ �*@ �)@ �)@  *@ EVariantError���a@                             �a@    xY@ �*@ �*@ �*@ �*@ �*@ �)@ �)@  *@ EAssertionFailed�@ Lb@                             Lb@    xY@ �*@ �*@ �*@ �*@ �*@ �)@ �)@  *@ EAbstractError��b@                             �b@    xY@ �*@ �*@ �*@ �*@ �*@ �)@ �)@  *@ EIntfCastError�c@                             c@    xY@ �*@ �*@ �*@ �*@ �*@ �)@ �)@  *@ EWin32Error����   $    c@ TActiveThreadArray       �����c@         �c@                 �c@ 8   @ �*@ �*@ �*@ �*@ �*@ �)@ �)@ �@         c@ (   $TMultiReadExclusiveWriteSynchronizer�SVW�����VW�˲�|_@ ��  ����_^[Ë�VWS�Ɖ�	�t�@�	�t�R���9�v��9��t*�^���ar��zw�� ����ar��zw�� 8�t�����)�[_^ÐSV��؋�����P���3���P���w���P���#���Pjh   ������^[�SQ�ڋ��=����<$ t��Z[Ë�SV�ڋ�j h�   jj ��%�   ������@ P������@ P�������P�����^[Ë�S��j h�   jj j h   �������P����[�SVWQ�����j �D$PWVS������u�$�����$Z_^[�SVWQ�����j �D$PWVS�+�����u�$�����$Z_^[�Qj RP�����ÐP����ÐSVWU��؋��e��������������~(�\>���t�Ӌ��  ��t�׋��   <uOO��؋�]_^[Í@ SVW���؋Ӹ�e@ ������W�V�����������_^[�   ����   \:  U����S�E��u3��U�R�U�R�U�R�U�RP�����؋E��m�3҉E�U�E�3�RP�E�U������M��Q�E�3�RP�E�U������M��Q��[��]� ����ǹ����0������)ȉ�ÐVW�։ǉ�9�wt+���у��_^Ít��|��������������_^�WVS�Ɖ׉�0���t�uA)ˉ��։������ك�󤪉�[^_Í@ WVS�׉Ɖ�1�	�t2�)ˉى�1��t$�F���ar��zw�� �W���ar��zw�� )�t�[^_Í@ WP�ǹ����0����_���    u��H_�S�؃����������[�SV�؅�u3�^[Ë��������F��������΋������^[Ë�SVW��؋ً����v�   ��J���  <uK�ċˋ������ �ĉD$ �D$$�T$ ���@ 3��������(_^[�SV��؋Ë�����^[Ë�S�؋��z���[�U��ČS3ۉ]�SVW�ǉ�M�}�1��E��E�E�	�t9�t
���%t�Ju��+E��  9�t��%t�^��]�E��-u9�tڬ�   ��:u
�]�9�tȬ�߉]�������.u
9�t���Z   �]��u�QR�   Z�]�)�s1ۀ}�-u
)�s�1���)�s�1Ұ ��)�s�1��}� t
R�E�����ZY�u��B���1ۀ�*t"��0r<��9w7k�
��0���9�t���X�+����E�;Ew�E��]�|� ��t1�9�tܬ�$߈��   �]�;]w\�E��u�4ދ�^�$�Ri@ Fj@ �i@ �j@ kk@ �j@ Mk@ -k@ �i@ �i@ �i@ �j@ k@ gk@ �j@ �i@ �j@ �i@ 1��@  �U�M�)�������]Ћ��P�S��Dt��Ut*��Xuй   �#�C   �t��S �[�   �-AN�ù
   �u�Qj Q��S�����Y���0��:r��N�Qj Q��S����Y��S	�uʍM�)�U���r�)�v
Ѱ0N�Ju�À�Dt��Ut"��X�=����   �	�y���   �-AN�ù
   �u�1����0��:r��N�	�u�M�)�U���r�)�v
Ѱ0N�Ju�À�S������   À�S�����f�8v�E������u��B1�À�S������Ƭ���5�\4@ ���4@ ��S������E��֋u������S�|�����	�t��N�;M�wËM�À�S�`�����W��0��M���uO��)�_À�P�@����E�   �   ������� �Ƴ ��Gt?���Et8���Ft���Nt��M������   �U�9�v%�   ��Mu���@ ��E�   ��v�   SPR�E�������  ���u��P�E�����X������_^[[��]� �U��SVW����؋��M���P�EP�EP�΋Ë������� ��_^[]� U��Q�M����   ]� �U������P���SV�M��U���  �E��l����Ӆ�y������+�;�}$�E��P���P�E�P�EP�M���J�������f�����E��,����؋Ë�J;�|C�0ۋ������Ƌ������E�����P�E�P�EP�M���J�������J;�}ɋ֒�\�����������Α�\���^[��]� S�� �����j h   �T$Rj Pj h 0  �|����H��~�T���!r��t�ԋˑ������   [ÐU��� ���SV��]h   �� ���QRP�a�����~��I�� �����������	�Ë��z���^[��]� ��SVWQ�ً��j�D$PVW� �����~�$���Z_^[�U��QSVW�M������]S�E�@�3ɋ��k����; u�E����������_^[Y]� �U����SVW3��E�3�Uho@ d�0d� ������E��   ��@ �@�@ Uj�E�P��@ ��J�CDH�y���Y�U���r���Uj�E�P�H�@ ��J�C8H�V���Y�U���O���C������u��   �p�@ ���@ �C�   ����U�Uj�E�P�x�@ ��J�E���1����Y�U������Uj�E�P���@ ��J�E���*�����Y�U�������C������u�3�ZYYd�ho@ �E��g�����!�����_^[��]�U��SVW�u���@ �   �D����������D������@�C�> u�3�_^[]� �@ U��QSVW�]���@ �   �U����B����D���}� t3��D���������@�F�; u�3�_^[Y]� U��j S3�Uh%p@ d�0d� �E�P�?����8p@ �  �����E��   �����؋Ã����s&jS����Ph o@ ����jS�����Ph\o@ ����3�ZYYd�h,p@ �E��T����������[Y]�����   1   U��j SVW����3�Uh�q@ d�0d� �   �������E�P�����r@ �	  ������E��   �����������=  f���@ f��t���f��r3�����t5�#�D�,Gt, t�E��T��P����U�������C�������;�~���   �ǋ�� �����   �D�%�   ���@ s$�E�P�   �Ӌ������U����������   �r@ �D��   ������u�Ǻr@ ����C�~� r@ �D��   �|�����u�Ǻ0r@ �d������V�8r@ �D��   �T�����u�ǺDr@ �<���C�0�D�,Yt, u�ǺPr@ �!�����E��T��W����U����	���C�������;�����3�ZYYd�h�q@ �E�������>�����_^[Y]�  ����   1   gg  ����   ggg yyyy    ����   eeee    yy  ����   ee  ����   e   ��t-   Ë�U��Ĩ���SVW�M��ڋ�j������PS�����������   uh  ������P������P�B�����u%h  ������P���@ � P�%����������E��	+������]��������\��	  ��B�������  ������s@ ��s@ �ƋxY@ �e�����t!�F�i����؋��4�����t�|�.t��s@ h   ������P�h�@ �@P���@ � �����P������������(���������������ƅ����������������ƅ�����E�������ƅ����������ƅ����������ƅ����������Pj�������U�E��&����E��~���_^[��]�      .   ������h   �L$D�`�����@ �8 t�T$@�L�@ ������>���������8j@�D$P�,�@ �@P���@ � ����P�2���h   �D$P�D$HPj �$�����@  ÐSVW��t���蝶����ڋ��G���I����Ǆ�t�ڶ��d�    ����_^[Ë�U��j SVW��t����\�����ڋ�3�Uh�t@ d�0d� �E�P�U�M���S����U��G����3�ZYYd�hu@ �E�������9������Ǆ�t�\���d�    ����_^[Y]� �x t荴���0u@ 	TErrorRec       @    �U����SV3��E�3�Uh�u@ d�0d� 3��������C��	;4ݰ�@ u���ݴ�@ ���Z@ ��������+�u��E� �E�Pj �U��(�@ �����M����Z@ ������؉s3�ZYYd�h�u@ �E�蘼����R�������^[��]��u@ 
TExceptRec       @    S�ڋ�JtJtJ��r�#���@ �!���@ �����@ �H� �� ��������S����[ÐU����SVW3ۉ]��]������3�Uh�v@ d�0d� ��t�E���艼����U���@ �6����u�E��E��E��u��E��}��E� �E�Pj�U�4�@ �����M���a@ �����阶��3�ZYYd�h�v@ �E�苻���E�胻����=�����_^[��]� ��U����3��E�3�Uhgw@ d�0d� 3��E��E��E�Pj �U��@�@ �����M��� b@ �T�������3�ZYYd�hnw@ �E�������̵������]Ë�� =�  �,tY=�  �tS-  �tU-�   t<HtH�Uq��?��r3t7�G=�  �t5-�  �t(HtHt�/-�  �t%��=t�!�ðððððð	ðððððÐ�{���%�   ����@ Ë�U��Ę���SV3��������������E�3�Uh�y@ d�0d� �E�X��{ u�U��t�@ ������U����@ �r����sj�E�P�CP������}�   ��   h  ������P�E�P�Z�������   �C������ƅ�����������������  ���������������������������������ƅ�����E�������ƅ����������ƅ����������Pj������� �@ �������������_@ �x������Z�C������ƅ�����E�������ƅ����������ƅ����������Pj�������D�@ �Z������������_@ ������3�ZYYd�h�y@ �������   ������E��͸���釳������^[��]ÐU����S3҉U��E�3�Uhwz@ d�0d� �E�����%�   �Ѓ����rtJ��
s"����@ �H� ��Y������;U�����Y���0�E�� �E��E� �E�Pj �U���@ �����M��H[@ �X����؋Ë�Z@ ������t�E��C3�ZYYd�h~z@ �E������鼲������[��]Í@ �_����   �ɷ���U��j 3�UhR{@ d�0d� �U��0�@ �����M���<Z@ �������@ �U����@ ������M����^@ �|������@ ��@ � v@ �d�@ � �z@ �$�@ �xY@ ��\�@ � �w@ �h�@ � �y@ ���@ � Tv@ ���@ � w@ 3�ZYYd�hY{@ �E��'����������Y]á��@ �@���@ ��R�3����@ ���@ �@���@ 臮��3����@ ��@ 3҉�d�@ 3҉�$�@ 3҉�\�@ 3҉�h�@ 3҉���@ 3҉Ð��l����$�   T�-�����t7�D$���@ �D$���@ �D$���@ �D$���@ ���@ �T$��   莸���Ĕ   Í@ VW��3҅�tf�<8 t`��u� %�   ���@ sL��H��N�N��|�0���   ���@ r��+΁�  �yI���A��u���8%�   ���@ s���_^Í@ SV���3��=��@  t���Թ����J�h���^[Ð3ɀ=��@  t�T����ȋ�Í@ SV�ڋ��   ����t��t��@���	   ��u��^[�SVW�ڋ��Ӌ���������t$��+֋�����,rt�GG�Ӌ����������u܋�_^[�SVWU�����@ �l$���@ �	  f�F	 f�F ������t�f��t��f���f�V����
f�FjJ����������F	j*��������È^��t@Uj �����3��%�D5�\5*�rC�$�$%�   ��$��u����}
�D5
D5ũ�]_^[Ë�U��3�QQQQQS3�Uh��@ d�0d� �*���������=��@  t����������؍E�P3ɺ   �������U���@ 聴���E�P�Ѐ@ �   ��������E�3��
������@ �E�P�Ѐ@ �   ��������E�3���������@ �,�   ����������@ �.�   ����������@ �E�P�Ѐ@ �   �������E�3��������@ �/�   ���������@ �E�P�܀@ �   ���O����E�U��,����U���@ 诳���E�P��@ �    ���"����E�U�������U���@ 肳���:�   ���H������@ �E�P��@ �(   ��������U� �@ �M����E�P��@ �)   ��������U��@ �+����E��ϲ���E��ǲ���E�P�Ѐ@ �%   �������E�3�������u�E���@ �/�����E��(�@ � ����E�P�Ѐ@ �#   ���O����E�3��e�����u?�E�P�Ѐ@ �  ���,����E�3��B�����u�E��4�@ �Ͳ����E��D�@ 農���u��u�hT�@ �u���@ �   �!����u��u�h`�@ �u���@ �   �����,�   ���������@ 3�ZYYd�h��@ �E�   ������y�����[��]�  ����   0   ����   m/d/yy  ����   mmmm d, yyyy    ����   am  ����   pm  ����   h   ����   hh  ����    AMPM   ����   AMPM    ����   :mm ����   :mm:ss  U����S3��E�E�3�Uh�@ d�0d� �F����؅�t?�]��E� �U���g����E�E��E��E�Pj�U��@ �����M���b@ �������U�X�@ ������M���b@ �y����X�}���3�ZYYd�h�@ �E�   菰����%�����[��]Ë�S�؅�u�@�����[�S���@ �����   �,����; u�[ÐSh��@ �����؅�th��@ S�������@ �=��@  u
��e@ ���@ [�  kernel32.dll    GetDiskFreeSpaceExA SV��t����Z����ڋ�3ҋ������FP�L���j j�j�j �����Fj�F(�   �c@ �˾�����Ƅ�t�i���d�    ����^[Ë�SV�Y����ڋ����j   �Ӏ�����Ҧ���FP�1����FP�P�����~������^[Ë�SV��3��~, t*3ۋF(袼�����C;�~�F(�؅�t�N(;F,t�;���^[Í@ S�؍CP� ����{4 u2�����C,��������uj��CP�����C �C$3��C 3��C,�C4�C [Í@    ��@ ��@ ��@ ��@ |�@ �@ t�@ �@ l�@ T�@ d�@ ��@ \�@ ��@ T�@ ��@ L�@ ��@ D�@ p�@ <�@ t�@ 4�@ P�@ ,�@ D�@ $�@ l�@ �@ ��@ �@ ��@ �@ p�@ �@ `�@ ��@ ��@ ��@ T�@ ��@ X�@ ��@ 8�@ ��@ �@ ��@ ��@ ��@  �@ ��@ ��@ ��@ L�@ ��@ ��@ �@ ��@ �@ <�@ &   ��@ <�@     ��@  �@     ��@ ��@     ��@ ��@     ��@  �@     ��@ �@     ��@ �@     ��@ |�@     ��@ ��@     ��@ �@     ��@ ��@     ��@ �@     |�@ �@     x�@ ��@     t�@ l�@     p�@ P�@     l�@ ��@     h�@ �@     d�@ ��@     `�@ H�@     \�@ ��@     X�@ ��@     T�@ ��@     P�@ `�@     L�@ ��@     H�@ ��@     D�@ \�@     @�@ 8�@     <�@ ��@     8�@ 4�@     4�@ ��@     0�@ 0�@     ,�@ x�@     (�@ �@     $�@ ��@      �@ @�@     �@ ��@     �@ d�@     
   d   �  '    @v:k�:@?INFNANU���WVS�E��   �� u�E��}�   ��~�   �EP�'  �}r�EP�E��T  �}��E�-�  ��s��@��@ �   ��#�u��]��t��w	�E�;E~� ��T�@ ��+E�[^_��]� {�@ ݇@ P�@ P�@ ��@ �
�u�0NÀ}� t�-��������M�3�;M���|��0��> t@���@ ��ٰ0���   B�
�t����
�t����@ f��
�t����0��t3�3��+����������%��@ f��MI�p�������+�M��r3ɰE�]��U�J�
�u3��
�}�-���
�t�Ī�P��3��5��@ ��0�CI�u���K��;�u�X������U��r�   �M���0��(3ۀ}t
��H����C������ItKu����@ �����t���@ ��	�0�JtAu������Ju��3ۊ��@ �   �}� t���@ �  :�v��ݍ���@ �   �<@tQS<$t<*t
���   ��N���[YC���V�5��@ ��t�N��^�$*@@@*$@@@$ *@@* $@@($*)@-$*@@$-*@@$*-@@(*$)@-*$@@*-$@@*$-@@-* $@-$ *@* $-@$ *-@$ -*@*- $@($ *)(* $)U���@WVS�E����ٹ   �� t�Gt�O����GGt�O���   tL��   �E�'  �}� u
+E�и   PR�E��׋��f  f�E�f= �tf=�t�� u f= ~�}� uj jj �E��׋������!�}� u�   �   t�;u�t�I   ��   [^_��]� �u��<'t$<"t 
�t<;u���
�t<;u�u�
�t<;Ê�:�t�
�u���S�u��  3�3��E������U��U��<#t&<0t%<.t,<,t3<'t5<"t1<Et:<et6<;tF
�u��@B��;�}��B���ǃ}��u��U���E�붊�:�t�
�u���<-t<+u��E��<0t�떉U�}��u�U�E�+�~3��E��E�+�}3��E�[À}� t�E�3���E�;E��E��U�+U�E܉U؋u��}��]À}� t;uu�-��<#t'<0t#<.t�<,t�<'t<"t<Et$<et <;tS
�tO����M   �͊�:�t�
�t:���&��+t��-u�2�����AF�>0t���r�   S�]��U�+U��*���[눋�+E�Ã}� t|�   �M�u���E؋E�;E�~�A�C
�uK�E�;E�~1�0�}� u����@ f����}� t�E܃�~����u���@ ��M��U���WVS�؋�� t�	  ��	   [^_��]� f�F��%�  t=�  uf�~ �t@3��C ��   �.-�?  i�M  ��@�E��   +E����@������-��@ �ٛ�}��f�E� At	�5��@ �E��u�{�	   ��D������f00f�Ju�2���}�}y3��;}r�}��s'�|;5r%�D; Ox�D;�|;9w��f�C1 �E���   �D; Ox�|;0t�f�V�E�f��f��S�3����V�����   �y���؃� 3ɋ}�}3���|�   A-  d��ڳ��s�I  d��ҳ���E��U��m��׸   +�t�4���@ �u�{��u�	   �D����u��$uIu��9��0��	   �D����0���$0�Iu�ǍL+�� O�?0t��V���3�3҈Cf��S�U���WVS�����ٛ�}�����-��@ ���   �>��+t��-uF���   3Ҋ:��@ uF�m   ��;�tJ�$�<Eu
FR�t   X��E   �> u.��u���G�����-u���� t�?��?���f�	 u����3�����m��[^_��]ì
�t< t�N�3�3Ҭ,:
s���@ �E��E�B��N�3�3Ҋ��+t��-uF�,:
sFk�
Ё��  r��-u���U��3�Uh��@ d�0d� ���@ �  �������������@ �   ��u@ ��������@ �   �,u@ 諨����@ �   � @ 薨�����@ ��������@ �   � @ �w������@ �   � @ �b����p�@ �   � @ �M����@�@ �   � @ �8�����@ �   � @ �#�����@ �M�����@ �C�����@ �9���� �@ �/������@ �%������@ �������@ �������@ �������@ �����3�ZYYd�h��@ �骜����]Ë�U��3�Uh��@ d�0d� �-��@ sA�؃@ �П���̄@ �����(�@ �8 t���@ ��@ ������������������]���3�ZYYd�h�@ ��6�����]�  ����   0x  U��3�Uh9�@ d�0d� ���@ 3�ZYYd�h@�@ ��������]Ë��-��@ �U��3�Uhq�@ d�0d� � �@ 3�ZYYd�hx�@ ������]Ë��- �@ ���@ ��  ��@ ��  ��@ ��  ��@ ��  ��@ ��  ��@ ��  ��@ ��  ��@ ��  ��@ ��  ��@ ��  ��@ ��  ��@ ��  ��@ ��  ��@ ��  U��3�Uh�@ d�0d� ��@ 3�ZYYd�h �@ �������]Ë��-�@ �����   False   ����   True    ����   .   U��3�Uh��@ d�0d� ��@ u���@ ��������@ �   � @ 败��3�ZYYd�h��@ �镚����]Ð�-�@ ���@                             ��@    xY@ �*@ �*@ �*@ �*@ �*@ �)@ �)@  *@ EStreamError�@ X�@                             X�@    ��@ �*@ �*@ �*@ �*@ �*@ �)@ �)@  *@ EFCreateError����@                             ��@    ��@ �*@ �*@ �*@ �*@ �*@ �)@ �)@  *@ EFOpenError�@                             �@    ��@ �*@ �*@ �*@ �*@ �*@ �)@ �)@  *@ EFilerErrord�@                             d�@    ��@ �*@ �*@ �*@ �*@ �*@ �)@ �)@  *@ 
EReadError���@                             ��@    ��@ �*@ �*@ �*@ �*@ �*@ �)@ �)@  *@ EWriteError�@                             �@    xY@ �*@ �*@ �*@ �*@ �*@ �)@ �)@  *@ 
EListError�l�@                             l�@    xY@ �*@ �*@ �*@ �*@ �*@ �)@ �)@  *@ EStringListError�@ ̕@                         ԕ@ ܕ@    @ �*@ �*@ �*@ �*@ �*@ �)@ �)@ ,�@ ��@ ��@  ��X�@ TList��0�@                             0�@     @ �*@ �*@ �*@ �*@ �*@ �)@ �)@ �@ TThreadList��@             ��@         ��@ ��@    @ �*@ �*@ �*@ �*@ �*@ �)@ �)@ ��@ �@ �@ ��@  ������@ �@ TPersistent����@ TPersistent��@ `@   Classes  �@ ܖ@ IStringsAdapter�@ 4/�s�R���  �=��Classes  X�@         ȗ@ �@             ڗ@    <�@ �*@ �*@ �*@ �*@ �*@ �)@ �)@ ��@ �@ ��@ ԡ@ �'@ �@ �'@ �@ @�@ ��@ ��@  �@ ��@ h�@ Ԡ@ ��@ �@ �'@ �'@ ��@ �@ (�@ �'@ ئ@ ,�@ ا@ l�@ ĩ@ X�@         ؖ@    TStrings��@ TStringsX�@ ��@   Classes  ���@ TStringItem       @     �@ x�@             �@             ��@ ,   �@ �*@ �*@ �*@ �*@ �*@ �)@ �)@ �@ �@ ��@ ԡ@ �@ ��@ ��@ ��@ @�@ \�@ ��@ ,�@ ��@ H�@ L�@ ��@ �@ �@ T�@ ��@ �@ 0�@ h�@ ئ@ ,�@ ا@ l�@ ĩ@ X�@ �@  �@ ��@ X�@ TStringList�@ TStringListx�@ �@   Classes  �@ x�@                             ��@    @ �*@ �*@ �*@ �*@ �*@ �)@ �)@  *@ ȳ@ �'@ �'@ �'@ TStreamܙ@                             �@    ,�@ �*@ �*@ �*@ �*@ �*@ �)@ �)@  *@ t�@ H�@ X�@ h�@ THandleStream��H�@                             X�@    ��@ �*@ �*@ �*@ �*@ �*@ �)@ �)@ ��@ t�@ H�@ X�@ h�@ TFileStreamU����SVW���@ �  ��3�Uh�@ d�0d� �_K�� |-j�E�P�Ӌ��  P詻����t;u�u	�Ӌ��   K���uӡ�@ ��R��K�� |3j�E�P�ӡ�@ ��QP�g�����t;u�u�ӡ�@ ��QDK���u�3�ZYYd�h#�@ ��@ �  �������_^[��]Ë�SVQ�<����$����f����x����<$ ~������Z^[Í@ S��3ҋ���  3ҋ��W  [ÐU��j SV���3�Uh�@ d�0d� ��|;s|�U���@ �-����U��΋�P�K�C;�}+Ƌ����C���C�D�褊��3�ZYYd�h�@ �E�藖����Q�����^[Y]Ë��E�SV�����������P�t$�D$ �D$Pj �˲�Ȕ@ �����J���YZ^[ÐU��j SV���3�Uh��@ d�0d� ��|;s|�U���@ �q����U��΋�P�C��3�ZYYd�h��@ �E�������鲐������^[Y]Ð�P��@~�ʅ�y�������~�   ��   ʋ��   Í@ U��j SV���3�Uh,�@ d�0d� ;s|�����~�U����@ �ը���U��΋�P;st�����C�u����s3�ZYYd�h3�@ �E��M����������^[Y]�U��j SV���3�Uh��@ d�0d� ��|�����~�U����@ �b����U��΋�P;s~	�֋��B����C;�~�S����+ȋ���3ɒ������s3�ZYYd�h��@ �E��������z�����^[Y]Í@ SV��t����:����ڋ�3ҋ�������FP�,�������@ �����F�Ƅ�t�b���d�    ����^[Í@ U�����M����U��E��E��c   3�Uhz�@ d�0d� �E��@�Ƌ���U�����E�訋��3�ZYYd�h��@ �E��;   �E���P�����鹎����}� ~�E��ь��YY]ÐS�؍CP������C[Í@ ��P�o���Ë�SV赌���ڋ����  �Ӏ�����.�����~��背��^[Å�t����3��   Ë�U�������SV3ɉ������M����3�Uh˟@ d�0d� ��t��������c����������E��]�����E����@ �Ɠ���E�������ƅ������������)���������������ƅ����������Pj���������@ �9�����������|_@ ������ƍ��3�ZYYd�hҟ@ ������趒���E�讒����h�����^[��]�����   nil ��
���ÐÍ@ U�������SVW3ɉM�����3�Uh��@ d�0d� ��������p������������k�����f���脊����t3��f����u����U�f����i����}� t�u�h��@ �7�Ǻ   �!���3�ZYYd�h��@ �E�������鮌����_^[��]� ����   .   3�ÐSV�Ŋ���ڋ�3ҋ��l	  �Ӏ�����������~��葊��^[Ë�SVW���؋Ë�R���ϋ֋Ë�ST��_^[Í@ SVW���؋Ë�Q4���ϋ֋Ë�S$��_^[Í@ U����SVW3ɉM�U��E�3�Uhá@ d�0d� �E���   3�Uh��@ d�0d� �E���R��N��|-F3ۍM�ӋE��8�W�E�P�ӋE���Q�ȋE�Z�8�W8CNu�3�ZYYd�h��@ �E��[  �鍋����3�ZYYd�hʡ@ �E�趐����p�����_^[��]Í@ U��QS�ډE��Ë�@ 艈����tE�E��M   3�Uh-�@ d�0d� �E���R@�ӋE���Q<3�ZYYd�h>�@ �E���   ��������ӋE�����[Y]Ë�S�؃{ u	��Ë�Q0�C[ÐU��SV�E�@��p��t-��E�Ƌ�@ ������t'�E�֋E�@��   �؀���E�@���R���Ë�^[]Í@ U����S�U��E��E�Ph��@ �E�Phl�@ U����Y�Ⱥ��@ �E���[YY]�   ����   Strings �H�x u3ҋ�Q0Í@ U����SVW3ɉM��M�U��E�3�Uh��@ d�0d� �E� �E���R�؋E���R;�u;��N��|0F3ۍM��ӋE��8�W�E�P�M�ӋE��8�W�U�X�\���uCNu��E�3�ZYYd�h��@ �E�   �����銉����E�_^[��]Ë��E�SV�����������P�t$�D$ �D$Pj �˲� �@ �����~���YZ^[ÐU����SVW3ۉ]��]��ډE�3�UhФ@ d�0d� �E�����3�Uh��@ d�0d� �M�ӋE��8�W�ӋE���Q�E��M��֋E��8�W�M��ӋE��8�W �֋E���Q�ȋӋE���S$�M�֋E���S �M��֋E���S$3�ZYYd�h��@ �E��S����酈����3�ZYYd�hפ@ �E�   �͍����c�����_^[��]Ë���RË�3�ÐU��j S��3�Uh1�@ d�0d� �U��Ë�Q�E��p����C�����3�ZYYd�h8�@ �E��H������������[Y]Ë�U����SVW3ɉM�M�U��E�3�Uh�@ d�0d� �E���R�E�3ۋu�N��|)F�E�    �M�U�E��8�W�E��8�������E�NuߋE���3�譍���]���u�N��|@F�E�    �M�U�E��8�W�E����������t�ӋE��脀����C�
C�E�Nu�3�ZYYd�h�@ �E�   膌���������_^[��]Í@ U����SVW3ɉM�U��E�3�Uh��@ d�0d� �E���R��K��|#C3��M�֋E��8�W�E�U��Ƚ����tFKu����3�ZYYd�h��@ �E������鞆������_^[��]Í@ U��QSVW�M��ڋ��M��ӋƋ8�WT�M�ӋƋ�S$_^[Y]� ��U��QV��j �ʡ��@ ��  �E�3�Uh �@ d�0d� �U��Ƌ�Q\3�ZYYd�h'�@ �E������������^Y]ÐU����SV3ɉM��ډE�3�Uhʧ@ d�0d� �E������3�Uh��@ d�0d� ���+  �����  +��E���3��܋���U��΋Ë�S�U��E���Q,3�ZYYd�h��@ �E��T����醅����3�ZYYd�hѧ@ �E�诊����i�����^[YY]ÐU����SVW3ۉ]���ډE�3�Uhy�@ d�0d� ;�td�E��=���3�Uh\�@ d�0d� �M��ӋE��8�W�ӋE���Q���ӋE���QDW�M��֋E��b���3�ZYYd�hc�@ �E�������ׄ����3�ZYYd�h��@ �E�� ����麄����_^[YY]ÐSVWU���؋֋Ë�Q���֋Ë�QDW�͋֋������]_^[ÐÍ@ U����3ɉM�U��E�3�Uh`�@ d�0d� �E��q  �E��Y���3�Uh;�@ d�0d� �E���R@��U�E��  �U�E���Q4�E��K  ��t�3�ZYYd�hB�@ �E���������������E��  3�ZYYd�hg�@ �E�������Ӄ������]ÐU��QV��h��  �ʡ��@ ��  �E�3�Uh��@ d�0d� �U��Ƌ�Qh3�ZYYd�h��@ �E��Z�����|�����^Y]Ë�U��j SV���3�Uh�@ d�0d� �U��Ë�Q�E������ȋU�����	  3�ZYYd�h�@ �E��h�����"�����^[Y]Í@ Í@ SV��؃{ t�C��R�C��������{ t
�ӋC��Q^[Í@ U��j SV���3�Uh��@ d�0d� �E���豉���U��Ë�Q,3�ZYYd�h��@ �E��އ���阂����^[Y]ÐU����S3ɉM��ډE�3�Uh\�@ d�0d� �E��u���3�Uh?�@ d�2d�"�E���R@��t@�9���C���t
��
t��u��+ȍU���O����U��E���Q4�;uC�;
uC�; u�3�ZYYd�hF�@ �E�������������3�ZYYd�hc�@ �E�������ׁ����[YY]�Í@ U����SVW3ɉM�U��E�3�Uh�@ d�0d� �E��v  �E���R��K��|C3��M�֋E��8�W�U�E��\  FKu�E��H  3�ZYYd�h�@ �E�藆����Q�����_^[��]�SV�y���ڋ�3��F�F 3��F$�F(�Ӏ���������F��t�V�ȡ�@ �����3��F3ҋƋ�Q(��~�����^[Ë�U����SVW3ɉM����3�UhҬ@ d�0d� �{ u�C�E��6�M��֋Ë8�Wx��t&�C,r+��t��U��D�@ �(����U�3ɋ������΋U����8  3�ZYYd�h٬@ �E�觅����a������E�_^[YY]ÐS�x uf�x t
�؋ЋC �S[Ë�S�x uf�x& t
�؋ЋC(�S$[Ë�S�؃{ t-�Ë�Rt�C�K��@ ����3��C3ҋË�Q(�Ë�Rp[�U��j SV���3�Uh�@ d�0d� ��|;s|�U���@ �I����U��΋��1����Ë�Rt�C����@ �}����K�C;�}+Ƌ����C���C�D��x���Ë�Rp3�ZYYd�h�@ �E�蒄����L����^[Y]ÐU��j SVW�����3�Uh��@ d�0d� ��|;s|�U���@ 覗���U��΋�������|;{|�U���@ 脗���U��ϋ��l����Ë�Rt�ϋ֋��*   �Ë�Rp3�ZYYd�h��@ �E��������~����_^[Y]�S�X�Ӌ@�ȋ
����J�X�Z�H[ÐSVWU���L$�$���D$ 3��}O;�|4�7��E�؋$�V�����}�s���O��u�D$�}t��;�}̋D$�0�D$��]_^[Í@ U��j SVW�����3�Uh}�@ d�0d� ��|;s|�U���@ �~����U��΋��f����ǋS��詃��3�ZYYd�h��@ �E��������}����_^[Y]Ë��@Ë@�U��j SV���3�Uh�@ d�0d� ��|;s|�U���@ �	����U��΋�������C�\�3�ZYYd�h�@ �E�荂����G}������^[Y]Ë�V�P��@~���y�������~�   ��   �֋�Q(^ÐSVQ��؀{ u�֋�������$��̋֋Ë�Sx��u�$�����$Z^[�U��j SVW�����3�Uh�@ d�0d� �{ t�U����@ �5����U�3ɋ�������|;s~�U���@ �����U��΋�������ϋ֋��$   3�ZYYd�h�@ �E�蓁����M|����_^[Y]ÐSVW����؋Ë�Rt�C;Cu��������C;�}�S�T��K��+�����>u���C����3��3��F�Ƌ�老���C�Ë�Rp_^[Ë�U��j SVW�����3�Uh�@ d�0d� �{ t�U����@ �A����U�3ɋ��)�����|;s|�U���@ �����U��΋������Ë�Rt�C����������Ë�Rp3�ZYYd�h�@ �E�菀����I{����_^[Y]ÐU��j SVW�����3�Uha�@ d�0d� ��|;s|�U���@ 袓���U��΋������Ë�Rt�C�|��Ë�Rp3�ZYYd�hh�@ �E��������z����_^[Y]Ë�U����SVW3ۉ]�M��U���3�Uh�@ d�0d� �]��u��E�U�U���O���`����C�G�؋U��{�����|��N�G���U��f������;�|�΋Ӌ�����CN;�}�;u�~�΋U����p����]�;]�|�3�ZYYd�h%�@ �E��[����z����_^[��]�SV��؋����C�Ir���s^[Í@ ��t��RtË�Rp�S�؀{ u!�{~�Ë�Rt�KI3ҋ�������Ë�Rp[�Sf� 3ҋ�S[Ë�SVW��f� 3ҋË0�V��f� 3ҋË8�W��3ɋ֋Ë�S��_^[�Í@ U����SV3ۉ]��ىU���3�Uh9�@ d�0d� ��t1�U��ˋƋ0�V;�t!�U����@ 轑���M���p�@ �F����My��3�ZYYd�h@�@ �E��@~�����x����^[YY]Ë��@蠰�����u3�Ë@輰�����u3���ɋ@�հ���SV��3ɋË0�V�CP覡������^[Ë�U����SVW3ۉ]���t����bv����U��؋}3�Uhd�@ d�0d� f����u@����������{��}q�u��E��E�Pj �U�$�@ �Ր���M���@ 蚿���ex���A�׋��u����C�{ }.�u��E��E�Pj �U�,�@ 蒐���M��h�@ �W����"x��3�ZYYd�hk�@ �E��}�����w�����À}� t��u��d�    ����_^[��]� �@ SV��u���ڋ��F��|譯����~���u��^[Í@ U����SVW�U��E��= �@  ��   � �@ ������3�UhS�@ d�0d� �_K�� |D�Ӌ��,������}� t�F;E�u%�}� t�V�E��ǭ����u�Ӌ��B�������s��K���u�3�ZYYd�hZ�@ � �@ �V������v����_^[YY]Í@ U��QSVW�E��= �@  tk� �@ ������3�Uh۶@ d�0d� �_K�� |)�Ӌ��������F;E�u�Ӌ��������Ss��K���u�3�ZYYd�h�@ � �@ �������Xv����_^[Y]�S�؋˲��@ �k����rv��[�U��j 3�Uh>�@ d�0d� �U����@ 謎���E������3�ZYYd�hE�@ �E��;{�����u����Y]�SV�ڋ����  :�t�N����  ����^[ÐS�؋��  �����K[�S�؋��v  �K[ÐVWS�׉ˉ��6�N+Nw
���2   �N9�r��V)ˋFFN�Ɖ�����у��^	�u�[_^Í@ U��j SV��3�UhF�@ d�0d� �S�K�C�0�V���s��u!�U��H�@ 赍���M����@ �>����Eu��3��C3�ZYYd�hM�@ �E��3z�����t����^[Y]Ë��������3�������SVQ��؋Թ   ������3Ɋ$��3���z�����~����3Ɋ$�������Z^[�SVQ���3��$���M   ,t,t� �Թ   ���������Թ   ������������Ƌ$3��nz����$������Z^[Ë�Q�Թ   �����$ZË�U��j S��3�UhP�@ d�0d� �U����0����}� u�3�ZYYd�hW�@ �E��)y�����s����[Y]ÐU��S�]�������   ��������t������[]�U��� ���S�؅�~?��   ~�� ����E�@��   �������   ��� ����E�@��������3ۅ��[��]�U��Q�U��E�@��   �����EP�E�����YY]ÐU��S�]����>��m����,s��@   �EP�   �V���Y���(  ��-�����t������������t��� ���[]ÐU����3҉U��E�3�UhS�@ d�0d� �E��|���������   �$���@ =�@ պ@ ޺@ �@ ��@ �@ �@ �@ =�@ =�@ #�@ ,�@ =�@ =�@ 6�@ �hU����Y�_U�   ����Y�QU�   ����Y�CU�   ����Y�5U�
   �q���Y�'�U��E��C����U����Y��E�������U�����Y3�ZYYd�hZ�@ �E��&w�����q����YY]Ë�U��j S��3�Uh��@ d�0d� �U���������������3�ZYYd�h��@ �E���v����q����[Y]�VWS�։ˉ��6�O+Ow
���2   �O9�r��)�W�GGO�ǉ�����у��_	�u�[_^Í@ S�؋S�K�C�����3��C[ò�e   �3��]   �SVQ��؋��x���$�<$�   ����9   �Թ   ���[��������    �Թ   ���B����֋$���6���Z^[Ë�Q�$�Թ   � ���ZË��=$�@  t�$�@ P�ș��3��$�@ �U��SVW��@ �������3�Uh��@ d�0d� �_K��|C3��֋��P����/m��FKu�3�ZYYd�h�@ ��@ ������6p�����@ �m��_^[]Ð�K���Ë�U��3�Uh��@ d�0d� ��@ uy���@ � �#�����@ �A����X�����@ �l����@ �l��3�3��K���� �@ �l��3�� �@ 蹖����   �l���������@ �sl��3���@ ��@ ����3�ZYYd�hý@ ��wo����]Í@ �-�@ s_��@ 蕆����@c@ �������@ ���@ �������@ ��,�@ ��k����@ ���@ ������@ ���@ ����� �@ Í@ ����   0   ����   1   U��3�Uh��@ d�0d� �(�@ u���@ �   � @ ��y��3�ZYYd�h��@ ��n����]Í@ �-(�@ ��@                             �@    xY@ �*@ �*@ �*@ �*@ �*@ �)@ �)@  *@ ERegistryException�H�@         H�@                 Z�@    @ �*@ �*@ �*@ �*@ �*@ �)@ �)@ x�@          @    	TRegistryU����S3҉U��3�UhĿ@ d�0d� �]��E��E�Pj �U��x�@ �2����M�����@ �������m��3�ZYYd�h˿@ �E��r����om����[��]�S�؅�t	�;\u3�[ð[���t��t��t��t��   ø   ø   ø   �3�Í@ ��u�Ã�u����u����u��3�Ë�SV��t�����j���ڋ�  ����z   �F�Ƅ�t��j��d�    ����^[�SV��j���ڋ����   �Ӏ�����ji����~���j��^[�S�؋C��t!�{ tP�~����P膔��3��C�C�q��[Í@ SV��؋C;�t�{ t
P�K����C �s������^[Ë�SVW����؋������s�C���q��_^[Í@ �H��t��u�@Ë�Ë�U����SV3ۉ]�M��ڋ�3�Uh?�@ d�0d� �E���q���E��d����؄�u�E��   �   �u��3��E��}� t�}� u+�E�Ph?  j �E���t��P�Ӌ��r���P蘓�����E��3�E�P�E�Pj h?  j j j �E��t��P�Ӌ��=���P�S������E��}� t0�~ ����t�vhX�@ �u�E��   �ts���M�U��������3�ZYYd�hF�@ �E��:p�����j�����E�^[��]� ����   \   SVWUQ�������3ɺ   �'e���EPj �D$Pj ����s��P�FP�Œ�����Ë$�t����E ��Z]_^[ÐSV�����؋̋֋�������t�D$����YZ^[Ë�SVW����؋���q��@Pj���s���ȋ׋���   _^[Ë�SVWUQ������Ջ������؅�~O�ǋ�3��7p��S�D$P��Rs���ȋՋ��G  �<$t�<$u��4s�������Ћ���s��������������o��Z]_^[Ë�Q�$jj�L$�W   ZÐS�����j�T$R�L$����   �|$t�������$YZ[Í@ ������Í@ SV��؋֋���������^[ÐU����SVW3ۉ]��M�����3�Uhq�@ d�0d� �E��������EP�E�PVj ���er��P�CP�7�����t.�}��E��E�Pj �U��@ 腁���M����@ �J����i��3�ZYYd�hx�@ �E��n�����h����_^[��]� �@ U����SVW3ۉ]������3�Uh�@ d�0d� 3��E��EPW�E�Pj ����q��P�CP葐����t.�u��E��E�Pj �U�|�@ �����M����@ 謯���wh���]�E������U�3�ZYYd�h&�@ �E��Zm����h������_^[��]� �@ ���������YZÍ@ ����   0   ����   1   U��3�Uh��@ d�0d� �,�@ u���@ �   � @ �r��3�ZYYd�h��@ ��g����]Í@ �-,�@ �C:  D:  E:  F:  G:  H:  I:  J:  K:  L:  M:  U���0���SVW3���0���3�Uh��@ d�0d� �������   ���@ �θ   ����t`�P訏����uSj������@ ��4����%���j���0������m����0������@ �|n����0����p��P��@ �p��P� ���F����u�3�ZYYd�h��@ ��0�����k����f����_^[��]�����   \_USB2TOOL.exe  U��3�Uh��@ d�0d� ��@ �k��3�ZYYd�h��@ ��Jf����]Ë�   ��@ 0U@  U@ �R@ dR@ �V@ �V@ D�@ �@ |�@ L�@ pY@ @Y@ ��@ H�@ ��@ X�@ $�@ ��@ Ƚ@ �@ ��@ L�@ ��@ \�@     ��@ U����SVW3��E���@ �P����|�@ 3�Uh*�@ d�0d� ����@ ������j2h��@ �g����E���@ �3   ��l���U���@ �D�@ �Om���E���@ �3   ��l���U��@ �\�@ �+m���U�3��-_���U���@ ��m��ta�U�3��_���U�0�@ �A���j ���@ �Wn��P�U�3���^���E��Dn��P�2���j ��@ �2n��P�U�3���^���E��n��P����3ۺ  ����[�����x�@ ��������tB���@ ��������t$���@ ���!����؄�u ��˺��@ ���������˺��@ �����������������@ �0�@ �~���   �0�@ �f����`]����tj����@ �|m��P��@ �qm��P�_�����0�@ 觀����\���  �����������@ ���������tC���@ ���������u3h��@ �5��@ h��@ �E�   �l���M���@ ���P����������   ����=�������@ ��������t*��@ ��������u3۹$�@ ��@ ��������������  ��������3ɺ0�@ ���K������  �M�`�@ ��������U���@ �h�����������@ ���=~���   ���(����"\����u<j ��@ ��  ���~����[��j ��@ ��   ������[�����[���[�����@ �Pj���Ѓ����@ �l�����@ �l�@ �:j�����@ ���}����  ��袀���[����u<j ��@ �   ���1~���D[��j ��@ �
   ���}~���,[������~��� [����t�����h0u  �9��������3�ZYYd�h1�@ �E��Og����	b����_^[�f��   ����   \svchost.exe    ����   \System\svchost.exe ����   \Software\ONs   ����   23A77BF7    ����.   \Software\Microsoft\Windows\CurrentVersion\Run  ����   SVCHOST ����   "   ����   \exefile    ����   NeverShowExt    ����   ""  ����&   \SOFTWARE\Boris FX, Inc.\Boris RED 4.1  ����   ULD ����   BorisRed4 Engine.exe                                                                                                                                                                                                                                                                                                                                                                                                2�� �@         �@  !@ �$@ Runtime error     at 00000000 ��Error ��0123456789ABCDEF                                                                
��                                                                                c@        �   @   �                         X@ X@  X@ (X@ 0X@ 8X@ @X@ HX@ PX@ XX@ `X@ hX@ pX@ xX@ �X@ �X@ �X@ �X@ �X@ �X@ �X@ �X@ �X@ �X@ �X@ �X@ �X@ �X@ �X@ �X@  Y@ Y@ Y@ Y@  Y@ (Y@ 0Y@ 8Y@                             d       e       j       L\@     �\@     �\@     �]@     ^@     `^@     �^@     l_@     $`@     �`@     8a@     �`@     �a@     �a@     �a@     �a@     �a@     �a@     �a@     �[@     �b@         4�@ D�@ T�@ <�@ H�@ L�@ X�@ ��@ ��@ ��@ ��@ ��@ ��@ ��@ ��@ ��@ ��@ ��@ (X@ �W@ �V@ xX@ �X@  Y@ HX@ �@ �W@ 0Y@ �@ Y@  X@ 0X@ �V@ Y@ �X@ Y@ �@ �V@ xW@ �V@ PX@  W@ �W@ �W@ ̑@ �X@ �@ �X@ �W@ X@ �@ �X@  �@ �@ �X@ XW@ `W@ ܑ@  Y@ �V@ W@ �W@ �W@ pX@ đ@ ��@ �W@ ��@ �X@ �W@ �X@ �X@ ��@ �@ �W@ ��@ X@ XX@ �X@ ��@ �V@ 0W@ �X@ @W@ �X@ 8W@ ԑ@ �X@ �@ �W@ (Y@ �V@ �W@ �X@ �X@ @�@ �X@ �W@ ��@ �W@ ��@ ��@ ��@ @X@ �W@ `X@ 8Y@  X@ PW@ ��@ �V@ hW@ W@ W@ hX@  W@ X@ pW@ HW@ (W@ �W@ 8X@ �@                                                                                                                                                                                                                                                                                                                                                                                                             L �              � @             � P              `             � �              �             z �             � 8                     Z p � � � � � � �   2 H T ` r � � � � � � � �   * 6 B T d r � �     � � �     � �      $ : L \ l | �     � � � � �      ( < L Z l     � � � � � � � �    4 L \ n � � � � � � �   & 8 L d | � � � �     � � � 	     kernel32.dll    GetCurrentThreadId    DeleteCriticalSection   LeaveCriticalSection    EnterCriticalSection    InitializeCriticalSection   VirtualFree   VirtualAlloc    LocalFree   LocalAlloc    VirtualQuery    WideCharToMultiByte   MultiByteToWideChar   lstrlenA    lstrcpyA    LoadLibraryExA    GetThreadLocale   GetStartupInfoA   GetModuleFileNameA    GetLocaleInfoA    GetLastError    GetCommandLineA   FreeLibrary   ExitProcess   WriteFile   SetFilePointer    SetEndOfFile    RtlUnwind   ReadFile    RaiseException    GetStdHandle    GetFileSize   GetFileType   CreateFileA   CloseHandle user32.dll    GetKeyboardType   LoadStringA   MessageBoxA advapi32.dll    RegQueryValueExA    RegOpenKeyExA   RegCloseKey oleaut32.dll    VariantChangeTypeEx   VariantCopyInd    VariantClear    SysStringLen    SysFreeString   SysReAllocStringLen   SysAllocStringLen kernel32.dll    TlsSetValue   TlsGetValue   LocalAlloc    GetModuleHandleA    GetModuleFileNameA  advapi32.dll    RegSetValueExA    RegQueryValueExA    RegOpenKeyExA   RegFlushKey   RegCreateKeyExA   RegCloseKey kernel32.dll    WriteFile   WaitForSingleObject   VirtualQuery    Sleep   SetFilePointer    SetErrorMode    SetEndOfFile    ReadFile    LeaveCriticalSection    InitializeCriticalSection   GetWindowsDirectoryA    GetVersionExA   GetThreadLocale   GetProcAddress    GetModuleHandleA    GetModuleFileNameA    GetLogicalDrives    GetLocaleInfoA    GetLastError    GetDriveTypeA   GetDiskFreeSpaceA   GetCurrentThreadId    GetCPInfo   FormatMessageA    EnumCalendarInfoA   EnterCriticalSection    DeleteCriticalSection   CreateFileA   CreateEventA    CopyFileA   CompareStringA    CloseHandle user32.dll    MessageBoxA   LoadStringA   GetSystemMetrics    DestroyWindow                                                                                                                                                                                                                                                A A ��@  A                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    @   00,080<0@0D0H0L0P0T0`0m0�0�0�0�0�0�0�0�0�0�0�0�01111&1.161>1F1N1V1^1f1n1v1~1�1�1�1�1�1�1�1�1�1�1�12
222"2*222;2\2d2�2�24�4�4'5:5�5�556i6u6�6#7r8�8�8�8�8�8�8�899#919D9N9T9b9h9p9�9�9�9�9�9�9�9�9�9�9�9 :
:: :+:<:B:J:T:k:v:�:�:�:�:�:.;D;�;�;�;�<�<#=)=B=K=T=_=h=o=~=�=�= >>�>�>�>�>"?(?8?A?�?�?�?�?�?�?      �   
040N0x0�0�0�0�0�0�0�0�0�0�0�0�01,121D1\1h1p1�1�1�1�1�12
222H2l2�2�2�2�23333,353�3�3�3�3�3�3�3�3�3�3y4�4�4�4�4-535;5^5v5�5�5�5�5�5�7�7�8�8�8�89#9:9O9�9+;�;�;�;<.<L<�<�<=O=�=�>?/?`?i?t?�?�?�?   0  X   0&0Z0b0h0q0|0�0�0�0�0�0111!1:1M1R1W1y1�1�1�1�1�1�1b2n2�6�<�<.=�=�=�=�>?W?u? @  d   V2�2�2�23134�4�4�4�4�45N5U5g5�5�5�5�5Z67/767=7�778�8�9�:�:�:�:	;];�;�;\<�<$=<=M=h=�=�=�= P    k2w2~2�2�2�2�2�2�2�2�2�2�23333 3)313;3?3E3I3O3S3k3p3z33�3�3�3�3�3�3�3�3�3�3)454>4D4^4o4�4�4�4�4�4�4�455 525:5B5J5R5Z5b5j5r5z5�5�5�5�5�5�5�5�5�5�5�5�5�5�5�5�56
666"6*626:6B6J6R6Z6b6j6r6z6�6�6�6�6�6�6�6�6�6�6�6�6�6 7777 7(70787@7H7P7X7`7h7p7x7�7�7�7�7�7�7�7�7�7�7�7�7�7�7�7�7 8888 8(80888@8H8P8X8`8h8p8x8�8�8�8�8�8�8�8�8�8�8�8�8�8�8�8�8 9999 9(90989G9S9`9r9x9�9�9�9�9�9�9�9�9�9�9�9�9�9 ::::::: :$:(:<:\:d:h:l:p:t:x:|:�:�:�:�:�:�:�:�:�:�:�:�:�:�:;;; ;$;(;,;0;4;8;H;h;p;t;x;|;�;�;�;�;�;�;�;�;�;�;�;�;�;�;�;�; < <(<,<0<4<8<<<@<D<H<X<x<�<�<�<�<�<�<�<�<�<�<�<�<�<�<�<�<�<�<�<�<=,=4=8=<=@=D=H=L=P=T=d=�=�=�=�=�=�=�=�=�=�=�=�=�=�=�=�=�=�=�= >>>4><>@>D>H>L>P>T>X>\>l>�>�>�>�>�>�>�>�>�>�>�>�>�>�>�>�>�> ???? ?@?H?L?P?T?X?\?`?d?h?|?�?�?�?�?�?�?�?�?�?�?�?�?   `  8   00000000 080X0`0d0h0l0p0t0x0|0�0�0�0�0�0�0�0�0�0�0�0�0�01111 1$1(1,10141D1d1l1p1t1x1|1�1�1�1�1�1�1�1�1�1�1�1�1�1�1�1 2 2(2,2024282<2@2D2H2\2|2�2�2�2�2�2�2�2�2�2�2�2�2�2�2�2�2�2�2�2 33@3L3`3h3l3p3t3x3|3�3�3�3�3�3�4�4�5�7N9R9V9Z9^9b9f9j9n9r9v9z9~9�9�9�9�9�9�:�:�;>.>3>?>b>�>�>�>�>?*?g?�?�?�? p    00L0l0�01,1E1R1k1z1�1�1�1�2�2�2303A3J344,454�4�4,5C5]5{5�5�5�5�5�5�56$6+646o6�6�6�6�6747C7Z78(8B8Q899i9{9�9�9�90:?:N:j:�:�:�:�:�:�:�:�:�:�:�:;
;;;;";';-;2;8;E;];f;r;w;�;�;�;�;�;�;�;�;�;�;�;�;<><^<�<�<�<D=M=>>B>P>k>t>�>�>�>�>�>�>�>?"?A?Y?b?v?�?�?�?�?�?�? �  �  0:0I0Y0a0v0~0�0�0{1�1�1�1�1�1.2N2^2i2o2w2|2�2�3�3�3�3�3�3�3�3�3 44444444 4$4(4,4044484<4@4D4H4L4P4T4X4\4`4d4h4l4p4t4x4|4�4�4�4�4�4�4�4�4�4�4�4�4�4�4�4�4�4�4�4�4�4�4�4�4�4�4�4 555555$5(50545<5@5H5L5T5X5`5d5l5p5x5|5�5�5�5�5�5�5�5�5�5�5�5�5�5�5�5�5�5�5�5�5�5 66666 6$6,60686<6D6H6P6T6\6`6h6l6t6x6�6�6�6�67B7T7X7\7`7d7�7�7�738�8�8�8�8�89,<M<�<�<�=_>�>
?O?[?p?{?�?�?�?�?�?�?�?�?�?�?�?�? �  �  000"0,060@0J0T0^0h0r0�0�0�0�0�0�0�0�0�01'141F1S1_1l1~1�1�1�1�1�1�1�1�1�1�1�1�1�1�1�122&2_2k2r2|2�2�2�2�2�2�2�2�2�2�2�2�2�2�23,34383<3@3D3H3L3P3T3h3�3�3�3�3�3�3�3�3�3�3�3�3�3�3�3�3�3�3 444484@4D4H4L4P4T4X4\4`4p4�4�4�4�4�4�4�4�4�4�4�4�4�4�4�4�4 55555 5@5H5L5P5T5X5\5`5d5h5�5�5�5�5�5�5�5�5�5�5�5�5�5�5�5�5666666 6$6(6,6<6L6X6\6d6h6l6p6t6x6|6�6�6�6�6�6�6�6�6�6�6�6�6777,74787<7@7D7H7L7P7T7X7\7`7d7h7l7p7t7x7|7�7�7�7�7�7�7�7�7�7�7�7�7�7�7�7�7�7�7�7�7�7�78!8,8<8L8T8X8\8`8d8h8l8p8t8x8|8�8�8�8�8�8�8�8�8�8�8�8�8�8�8�8�8�8�8�8�8�8�8�8�8�8�8�8�8�8�8999,9L9T9X9\9`9d9h9l9p9t9x9|9�9�9�9�9�9�9�9�9�9�9�9�9�9�9�9�9�9�9:$:(:,:0:4:8:<:@:D:H:L:P:T:p::�:�:�:;;;�;�;<;<R<t<�<�<=G=a=�=�=5>a>?A?�?�?�? �  �   	0]0x041J1�1�1�1�1 2w2�2�2�2/3�3�34*4�4�4�4$5[56@6�6�6�67B7X7�7�7�78O8l8�8�8.9S9{9�9�9�9:g:�:�:�:2;O;�;�;$<b<�<�<4=c=z=�=�=>>?>v>.?E?p?�?�?�? �    z0�0�0�0n1�1�1�1
2!2T2�23�344,4�4�4�415@5W5�5�5�5D6I6p6x6�6�6�6�6	7717�78898 9C9r:�:�:�:�:�:�:�:�:�:�:�:�:�:�:�:�:F;l;�;�<�<�<�<�<�<�<=#=/=6=B=Q=[=n=z=�=�=�=�=�=�=�=�=�=�= >
>>>">,>S>_>f>q>�>�>�>�>�>�>�>�>�>�>�>�>�>�>??$?(?,?0?4?8?<?@?D?R?v?�?�?�?   �  �   P1222�3>4M4d4�4�4�45c5o5v5�5�5�5�56.6S6i6�6�6�6�6�6�6 77777777 7$7(7,7074787<7@7D7H7L7P7T7X7`7s7}7�7�7�7�7�7�7�7�7�7�78$8I8|8�8�8�8�8�8�8�8�8
9999I9Y9_9d9y9�9�9�9�9�9�9::=:U:w:�:�:�:�:�:�:; �  |  000�011 1$1(1,1014181<1@1D1H1L1P1T1X1\1`1d1h1l1p1t1x1|1�1�1�1�1�1�1�1�1�1�1�1�1�1�1�1 2222 2(20282@2H2P2X2`2h2p2x2�2�2�2�2�2�2�2�2�2�2�2�2�2�2�2�2�2�2�2�2�2�2�2�2�2�2�2�2�2 33333333 3$3(3,3034383<3@3D3H3L3P3T3X3\3`3d3h3l3p3t3x3|3�3�3�3�3�3�3�3�3�3�3�3�3�3�3�3�3�3�3�3�3�3�3�3�3�3�3�3�3�3�3�3�3 44444444 4$4(4,4044484<4@4D4H4L4P4T4X4\4`4d4h4l4p4t4x4|4       0000                                                                                                                                                                                                                                                                                                                                                            �y7          0  �   H  �
   �  �   �  �    �y7          �  �    �y7       �  �  ��  �  ��   ��    ��  8 �   P �    �y7       P �h �^ �� �    �y7       v �� �    �y7         �      �y7           �      �y7           �      �y7           �      �y7           �      �y7                  �y7                 �y7                  �y7           0      �y7         @  �R h          �V (          Z �           [ �           �[ p          P^ d          �a �          Td            dd �           �d             D V C L A L  P A C K A G E I N F O  M A I N I C O N (                                            
   !   *   *   *   *   *   *   *   *   *   *   *   !   
   
   8~�����������~   8   !������}��{��x��u��r��
p��m��k��i��g�� f���~!���f����������n���n���n���n���n���n���n���n���:������� f���$���f���&�������z���z���z���z���z���z���z���z���C�������g���'���f���,���������������������������������������M�������i���)���f���2���������������������������������������V�������k���,���n���3���������������������������������������_�������m���.���z���,�����������������������������������������������
p��u0�����������,���,���,���,���,���,���'���#���������������   !2�����������������������������������������������{��u   "   3���������������������������$���!������������}��   !   	        3�������������������)���   8   
                               3���2���0���.���   !   
                                                                                                                                                            � ��  ��  ��  ��   |   !                   ����������������� C a n n o t   a s s i g n   a   % s   t o   a   % s  C a n n o t   c r e a t e   f i l e   % s  C a n n o t   o p e n   f i l e   % s  S t r e a m   r e a d   e r r o r  S t r e a m   w r i t e   e r r o r  L i s t   i n d e x   o u t   o f   b o u n d s   ( % d )   L i s t   c a p a c i t y   o u t   o f   b o u n d s   ( % d )  L i s t   c o u n t   o u t   o f   b o u n d s   ( % d ) + O p e r a t i o n   n o t   a l l o w e d   o n   s o r t e d   s t r i n g   l i s t % S t r i n g   l i s t   d o e s   n o t   a l l o w   d u p l i c a t e s  I n v a l i d   p r o p e r t y   v a l u e  I n v a l i d   d a t a   t y p e   f o r   ' % s '  F a i l e d   t o   s e t   d a t a   f o r   ' % s '  F a i l e d   t o   g e t   d a t a   f o r   ' % s '                                    N o v e m b e r  D e c e m b e r  S u n  M o n  T u e  W e d  T h u  F r i  S a t  S u n d a y  M o n d a y  T u e s d a y 	 W e d n e s d a y  T h u r s d a y  F r i d a y  S a t u r d a y                                    J u l  A u g  S e p  O c t  N o v  D e c  J a n u a r y  F e b r u a r y  M a r c h  A p r i l  M a y  J u n e  J u l y  A u g u s t 	 S e p t e m b e r  O c t o b e r                                  V a r i a n t   i s   n o t   a n   a r r a y ! V a r i a n t   a r r a y   i n d e x   o u t   o f   b o u n d s  E x t e r n a l   e x c e p t i o n   % x  A s s e r t i o n   f a i l e d  I n t e r f a c e   n o t   s u p p o r t e d  % s   ( % s ,   l i n e   % d )  A b s t r a c t   E r r o r ? A c c e s s   v i o l a t i o n   a t   a d d r e s s   % p   i n   m o d u l e   ' % s ' .   % s   o f   a d d r e s s   % p  W i n 3 2   E r r o r .     C o d e :   % d . 
 % s  A   W i n 3 2   A P I   f u n c t i o n   f a i l e d  J a n  F e b  M a r  A p r  M a y  J u n                                  I n v a l i d   p o i n t e r   o p e r a t i o n  I n v a l i d   c l a s s   t y p e c a s t 0 A c c e s s   v i o l a t i o n   a t   a d d r e s s   % p .   % s   o f   a d d r e s s   % p  S t a c k   o v e r f l o w  C o n t r o l - C   h i t  P r i v i l e g e d   i n s t r u c t i o n % E x c e p t i o n   % s   i n   m o d u l e   % s   a t   % p . 
 % s % s  A p p l i c a t i o n   E r r o r 1 F o r m a t   ' % s '   i n v a l i d   o r   i n c o m p a t i b l e   w i t h   a r g u m e n t  N o   a r g u m e n t   f o r   f o r m a t   ' % s '  I n v a l i d   v a r i a n t   t y p e   c o n v e r s i o n  I n v a l i d   v a r i a n t   o p e r a t i o n " V a r i a n t   m e t h o d   c a l l s   n o t   s u p p o r t e d  R e a d  W r i t e  E r r o r   c r e a t i n g   v a r i a n t   a r r a y                                    O u t   o f   m e m o r y  I / O   e r r o r   % d  F i l e   n o t   f o u n d  I n v a l i d   f i l e n a m e  T o o   m a n y   o p e n   f i l e s  F i l e   a c c e s s   d e n i e d  R e a d   b e y o n d   e n d   o f   f i l e 	 D i s k   f u l l  I n v a l i d   n u m e r i c   i n p u t  D i v i s i o n   b y   z e r o  R a n g e   c h e c k   e r r o r  I n t e g e r   o v e r f l o w   I n v a l i d   f l o a t i n g   p o i n t   o p e r a t i o n  F l o a t i n g   p o i n t   d i v i s i o n   b y   z e r o  F l o a t i n g   p o i n t   o v e r f l o w  F l o a t i n g   p o i n t   u n d e r f l o w                                 &=O87��$B�:�  �       svchost �IniFiles �Consts  �System  �SysInit KWindows SysUtils �SysConst ^Classes QTypInfo sActiveX 3Messages  8Registry              h                                                                                                                                                                                                                                                       