MZ�       ��  �       @                                      � �	�!�L�!This program cannot be run in DOS mode.
$                                                                                                                                       PE  L             � !
 L   >   >  �                                                                        � <                           � �                                                   � $                           .text    P      ,                    @.bss     @   `       0              �  �.rdata   0   �      0              @  @.data       �      B              @  �.rsrc       �      D              @  @.reloc      �      F              @  Bccc            0   R              @  �                                                                                                                                                                                                                                                [�JZ�T��/w��>��Y|Afr�u�A��%�����c�K�����������Ҧ�����������N��,ӽ󫻨�Q�N��k��[�Gc��d܄<�T��lXa���u��[��Ft7���Vc�tD�ӓ	��>V�7����WN��k�~�!ov�J�x^�N�N��`I�<�֒�W���ҵuΈ�P^+�A��z��+��Q*\��vO�����'���kl�^��rI�m�ڋ�t)��$\�Q$�t��'�rL�D�Y�;
$D/��	�6�d��+m}�� �+S��]8/��)'Q�p��2TV/��gBט��}�����6�R�����@{SI:w%A4��;��Xfd���?($�h�}������ֳϡ��N`�3&:eRŒ�d���HƎ�G���}ash�8O��(�����,}O2��m{��AJ�������g&��@��%�����⢽\�����cR9y䕄t_{-��2���rރ���H�����"��/�o� q!�RQp�i�~�>�ȏ��^'"��;Q*�������:��m�;Kj@��Φ~e�1�b��I���H ��}��BO�AE�dޜ�����(;�bk��	b���� Ø��U:��9WZ)HZ�Js(F�[����A�I-	J��˘4���Jӆ���JjZ�P�''��Z�z���Z�����J
o�e��E����6�7"�Z6��R=c�]C� �7�⾑1�ߒ�C�ʹp�z7�]n꣛��V2!�t�9�i�M��A iz�_�^K*n)�Kt�a��~1�}Ǩ���}U��'���L(>�baC�+m�x�0��Q�W��Ǫ�Y������/���������l�ߌ$�btW+W���}���p�L�b?C�OݣI�'mmZؒN�?An�E�>�o�V^�e|:%^�e}&	�� Ҙ�@~/��u��/��|�������q��)c�_�V��E`�n���x�$<���B-�Y�/{Ϧ��b�OB�����3�����x9�2��ډa�&����ΩK��x�В�
�V��1{��+�<�4�
��ܠ���]�'@#�ٸl��v��=�Q��؈81�i��Z����й������%FY���r@L@2��.L��6Q�B�>�H6���:�;���iax\�BV� g!������3& z�Np�.���Ҫ���N��fO4J���-���p�V#��oL���^5�P$�T��SI�]]$&�>��a��*�������D݌�jf����,M8'�.&jα�I�ܑЂ�� �"98���8"5!��I/��$_G�]$*U�lT�zﬔ��ХʸZW#2�/K	#sy�<�s��|��'+���1*�A�81᎗S�8������;FsL�Z�@wЮN�үn�a����{1@}�Ʀ�U�2���F�(!=����o�T&���$�I�".:msE,�b�����0�S���}�m7�@غ�3�a�E�5P:��|�ڸK��$+Nn�a�I��we�r_�D��(�,m1>��:&��k�^v�Jq�p7|2�%��3ߢ	�!��Cߔ�Auztϒ�bQ ݞ��A|pE\�C����YӒ�\w��a�/{Vsf�}�j�lC�N��L-�h�J&��Ի(rY:)V3 �(R��]:`4!�yT�U7�|V-��Zp=��Pĥh���L�ynN���a�Қ�*8����~O
�9����^3hPU�q�'��.���s��̂g'忯\���N��'��#��Ȏ|ǃ@���j���o�/�A#1��8CeӴo�M�wW��fˢT�v�k��
|>�eͭ<uh�q��Kؽ�)�c`-y��zՃ�Y��ew��}\"9�o�6�c~���0o�;���C��i�%�b�6Y�%����0�;4_��t=��`�ř���C�'�s.^��76�3��h裔Pp5�l.������J��a\Q�����L|CT�����ER�*�GG�ua�I�|MN� B /�̳f�Q�L�B�K����5�e�Ύ,v�D@�8�/����;�	����h�}�w��ʷ>^=FIj���QR�$/n�$��NhE_�>���N���Hi^���2}�Kk��G��B�$;��n�0_�+��,*�i��I0��Р��<��`}�2r��Ղ=8Z�(Z�|$+�S{�
6�5]��/䥯���iJ.�Yhuû�SP�r|K��%�̲~��	�{9=���Ro	�&��)���i�H�橈��V���^����P�9TF>kz���ac�!]�|*Z���� �"ѭ��qtA��ҵ���ۺ�w�~D������&0�^Amu;�١|��J�#�(L�)jׯf�Q(8���w��>�D[?��}��a��^>��׵�`|�Xf�4rM����1r|a�$9:�=yi3~�\�e)"�������I��8��<%t�r��B�~{���W�Ԋ�<���i',P�1`�W&���r\uu����G�������|]� xr&6R���T���a��`��"�ұQ�I��p%�ݽ�,D���5;�q̱2�ַ`D�U/��������א���b(�g���H�Ǐ
�rUC�i\�P�f���H�7�\��~�ec�q�������A&�(P�$��ȍϸͧ(^�SE�A�Z��&�>���X��;�FQ���7��\��Y@Eы���.�J��f&�A{X{�ʖ��i�m�a��i2�t�v�{N� O�\�6S��랑 өJ�G>�V��ߛ>L���"�9D�m���T���奐���R�}��i���K���6"�EK�>��ag~:��3{i�w��x����	�^.���n�n�1_AF�-���2k��3��,�Sj1jc\�(�:��D��=k�2>7�	��i�3]���?wwS?hi=8���m���p���ن��g�ԺOMeI7�3�9���\�\O�0m�r��	xk�Rb��]d�б���2w�yU��G�K�g}�tWR��׮�g/S���R2$m���=q��i��YS��2R�{U#��i,l�G������ZʋE@I^)�m��&��8g�D#�� j�յSǼ�/�M�		�5=AE1*�"�-��t��5x��+41v�P}1ˬH���Q���T�U�PC�zVC/�F��
jb��EMX��*�,�x<zw<Z�����y�x3��x[�cV����Gq^T�5�!�օ\y��)Q������4�m�vљL�9��R�C�KF�����I=����B7�ޢ^̶v�bԇ�W?��@S�V<�P�
����Ct�o�d��2��y�@��'q�8vy{ ��^aF�3.��y����hE�����t�`�n�N,zd?$,��?|�0��m1"��Lm�n��ZVػ|1'f)��TG�-Wrr�9�]v��X.l��<Ǻ�H̧�H��(!���kG�������	HX��ܛ�O��;mʂލ��=��̋s��y$�
�J��W����&��.�Yp�8����yꕪ���ϥ�DV�砀�]�F�~�o��g��Д+{��ίԩ��_i�[H%�J[/���}|�ރ9�g�!o�㉛ 764i��Ɉ�ɦ&��Uqw� ��qL��bh���ځ�Y�|2��4�A0�%��ķF&)	Ί�N~QL������U��䢹�ԕ4�i]@�ꕷ���P��
熦�H�n����=�N�Hpפ�p����'h#as�d�ȭE(.�Z)�v��tz�j�>���';���/4��Ҍ�D\@�|� T��@q����[�E���PC�/�;�e#ǻ2��>�d`���>/�'��0h��P���ܟ���5����Y?멌���g2P�!�a���T�K۞f{��J^$\�	.:�[ː0���>��̩�%���o_��+&�{�cU���}�4n��a6�Җ֏[~J�a�藔�I*"^��v,wZĿ�z�ʕj�j+2�,	��]^>�[*�6�c�.2җ�⻹��j�;ﾱ=�J�n1SG�̟ ��3[^� ��0��Kw�� �X�P��
R��'�S��:=�nfz�8(:M� hKۣ=�-Mွ�g��~ހG�b�Spt��p3}�;L�Sl�ˋ ���L{��hr>^��P��"BL��ﶿ�nz/�#&GI_=r��/_e�x��n�+�[�Bc#����c뺡7�ȅ.(r�=�$��L�q�E��������S���Q`ӭD���q��g�W���$�5�����|��hj���-p���� �\m�I���ûDEG�[�,��	ݴ��c?ӟ��W̕U�M1x��5��b.�	ڧ����.�?v	��N��J-I���}ޙOZ�4��{e���t��&�q/B�t�?SX$0X�,����B���x�wX��3���}�n ��4�L���[Ŏ�ƙ�x�]x4M�_4���+�p�6���~cν:S���Sp[E��T�;נY�S�Gj�V��N��s�^�H$W\׻a;�%�6oP%���"�g9'YLٴ�����>�D�jQ�_)�	x�%��$^�ȉ��7����r��¢�B6Mu ���(��Rb�Ӊl�7�D�¢2��Ǎf��"�2�X�
��c�M"{x^���T$�Եd��d$���&�6��f�����E8���/�2|>������W/�;U0��~�Z�@4�*��n�ᰚ��k�.�Ȁ�[���;k��5uM_�Rk�b����HgPg����M�ȟ�x��o��Hr��Y�N@�W.�\��v%2Fd`IӪ̳J���2�z�9�O`�W3�ŽGØ�,���>b*��KD�)I�S[��p�����ej���Y���\���X/
W���b̳����k%A/�`��.x�Uڥ�&c�	>�0½F�&������<��j�r{�S�h�z�0R�Vbi-�- 5�Ze�;��}y%��L�y�����4}JW2-��w�5�1����V�T9���V����Q�z���w�� m�J�#��,#g�uSZx/�4�|�}Dљ#�X�>Fά"yY�GU�h�S2��uT��u���"B��n~��p��T*�U3��f��Nx=��3Ȏ�<z�w�j�f��z"7��2"����×j��7��2����4�n�eK%s��L!Qm�)5��-Kg���&ĎJ�h�������NK�<e{߿cZ�Ĩ�?��2�@S<�?*6��ߌk�8���n�\k�hEi}.�0���c5��N� 雤#�<%Z�1�a{ ���ۯ�8�N*�Q �C�x 7�T��D§�to��B��S����H��v���/�:�8��{��?U�f�ntɎ��(�?�Q�#C��<awt����H�ơh�V0���0�Qh�ُ�N+����|$̚=�dA��F�yj퀺#Ԓ^W�G��4� � ?��b�,���W�R���ؽ�@����H�a��Sy:�B�]3�ԝ�qś�K[��/�<"�B�ǎ�T�^s<����\gU��G���jF,*	!��W]�?��U��fK(��m�h��5@c<YKt=��`�_w�-��TxR��U�sH�+>�6o �~�=�RDd~:��0�K���w�L�4 |�c�5�fZ��z6�YmW��r9`�5Z�Ē����s��懄����Jf�$-rP�|.1�\R�F�����3�
Hɣ�Os�KZHh^5ʢ����d
�!>���]�x�_s1�#�y����*��M[��R)���_X�P�۶�,��O����j���\��p��(�g3�M����G��[Mo8�m�������w#��vz9}$xZ\_p0W��m;T��nH"P,]"Dr��cϸ�T�/�[Y�#/I��f��0�8@$zpa[�@T�_�+T�(��ӄ8�18]ԽJ}[��.l5u�� �x������
Q�}�u�%�H'�;��z0�O�Es�������pV�����1~k2�1ʭ���
J%��<�QLK�]��I���}�
d�sKkZ���?R��ui ��3.m��9J=�z��CXզ8g%Zl$���X&�ܣB	^{;dN��H�^��b[�������Ox�E%����a$�l��{Ivb��>��K3�$�$B�[A(ǥx�O^Ƙ�w��5���Èr@�L1�z�e��>8=�9�ؘv:���#��[����a(%o�Q\o�_��C�
��2n��W�e�Һ�&X����Q&�� M�>q �%��.������O����C���0��4�[������2� �� ��e�Ob_0����R���S��w��Ӭ϶?'�F����?[m1�� ک�.�
�\�1#����w}瀾�,��#��Ru?�-���㡽�\{�7D�F��ۚ)a��M;^pC��G��vO�0��hw\���!�ɫ`��t�����)ߒh�B�~[��ad�}MHî^��>\�s� �ܠ��y��g'�@Gp2^ru��g�j�D�Wc�m��k9H��P&�(��4?2���mo���X[0�Ć�n�P��&27sjU���?S��c������]�ڝ���>o��u�KO7�e�\>6/d��g0_]��NmE���-�ϵ �kaJ���������͜��W��?:{h����m�n�ҹ���T�ƕ��	��C�ǆa�w5� \�a���iz���ؒ�h���k-=���Ur�������"f�\]�ci�ܡ�?T��</9cڷU���8( L��Y��녵�IH����uP�˾Ež]tXNkҡ"���j��8��.F��	�w�O�]$� �T��8����9��'�[��u���������LoZ���,��n�C�f���Q���ңڲ#��Kɻ�2�7�����q�a��B���Ѻ,��0����@�-^#+��,"�3h@W_g�#�{tUI�)�/<�9b�su�:������	T��+�� �v�4\�� f`��	��g����>���Ox��h�Im`��²�&�Sٱ @�ꘒ[��1hc�c�1���izh�Z��c�
�X(��lӘ�:�F�U�`'��}ݚ�S�$�]�]ht����6U��2{�j��w{��H\ ���������X�� �7B`�)�cayƿ�ՠ!�JN(H�����+��Ue=7Bt`M:ʎ�O��x�<���Ǹ��R!��$�t](��6���w�TJ���I�J�a0)��HR5�!p�vB� 8Lg�������o�t���O˖9�ɣ�ک���ta������4��Y���buRZY��v`/�H�H�e��~�NU2Q�l�2{�g܈a�V�t_3[�萳����˟�4P	����[G�,��oc"lN\�H�D~�c)!=���ċ5@,?��K�;_A���WڂI��a�|���6U7)�Gd��)G�ʃX�m��%zSvL��$�
���� �{��xto��>%''��S�ӵ��D�����7�	`�Ϙ�
��s�A�r@
�3yL5΅yӃ�s6��&f�5��Ȍ2It�DM���2��$ b�j6��nc��;���`���*�A�f��'I�U�gkЂ�~�����'>W���EB�u';�ʖ�L��~�G��x����b�Tf��&��xU��O�l��{�C�L,�T���e�Ky�Q5�&a�{Q�.��{��E�.:1�Z:�jw� �I\�n��Ѭ.��/9q$��)4r*r�8��W�o��6{�q��@qx�i�h!�q�y��Y��t����\g�Qcpv{�`��DpZ���q�-��0y�I�$�y�*����A��p�Y�}���gݢ>fr�?	b�)�׈���w�K���^����[^�l�.�3tV�`���D4:!<�.����Y|^�Z�O����ga���"��JL��ɔ�ك�k@���H���b�'0:>R���Cy���t�F�ħ!��ʳ�;�s�͆�T\� ���Vm��U�SS"Ҋ5�J��,�E�:��͝<4��{��'��~�i|���Tn^�t))ƨ>�\툺���,_��n��M7��`}�B'ϟ=��h���Lk�u���"ޟ���aѽ���X����4��+]i��v�Xg���G��`��rV4�H�\�PCV�����o��>���Ml�>��}|>	M��ީ�i2�D�����&�}�F���p��L�_T� �x�`�j�G<�l�����Ą+w�΀�7�2���%:"�Ɲv�;�w7���Ĉ���XHC�(-�3���m����щoͦV���[d��ygT)]�x��8F��П��z��#�iyv�geuR�Ģ-�Y�� �sި�{BD/�r�#+���}苈�[���e
ir��3VH ��Mp��NP�8Z�_u/�R�\����b���ku����Wd�WY���kƌ�8;��P5a�����U�����,�34��I��Vmg���<�0<�H���T�1Q�{���I��3#QG��.W����{Q�-s�걎v�!�z>�qh���'�Ӷ���΀'G\���E�9�d菂+����j��>�\�e����%������T0�$�-_�ħ`ܘ�N���fH�����m� �c1�JՁ�W���g�?l{=m:�q�V<b&�M��P#P��4�}�Z�ET�Ep+`�]ԅ�plACe*�Q�T�an�'�D�W�{�M�Debb�[w3*I��ܴ`�!�քc{r��+U#on�e�S�� �Q�l沕�e#���'��5H�Ϋ���^.}B:��3�d�w�`"����<Z�л��(0z�N�9	N�1�z������`������+� �j�L�#�o�e�z9���7����{T2O�"s�dH���!?� ��z𔁹 ql�����-{L����"32�t���w!��
$"��QӐ���R�E�P�Ξq�4D�"C*�O�.$1�����t<���x܂�e�
;�M����0�u�X袅&�%(!�j\+�� ?d�,B[b��oH���ߓ��d�?�X�o�(4�ʖ�t�ذZ�x_)��!��2TG*Ձxy΢_U�!e��H��a.Z���q�y�ј�`a�]/�v&Ϥ��E�n�q*�
N���{h��!&[�wAA�&����������V�\�~�e�E}��
�#";�=��L��4i
W�~�ed�D"B��$Γnj�+�C�<��ï�s��әY���0���S�y�آ��)⩐d�6p`\�"#&���� ��_���'[A� �jG��Y���W�_��N��Ќ�A�O�Ċl��4�[��k(�P�fa;���(���V�ۃV�>�!!��-b�"�(;C��(4��S5�7�.H��ܰ�M�L���_�W�.�&��G	�-����Ӵ��ٙ�&��BO�4Ո
���Д�8����_� �'��������Hf��a0q�
nC+vP��t�7�oo�ڂ9A��������r��_'h	)W2�����3(�M(A+>=Cԓ��ྠLn	k7@��!r)bG=��aS�-��3�ޯ�/L%����^,��P񹘏1�I�2�7p��8�J��$#8�������&�g�}�栱�
6e
LH�����o��K�/ϻ���	0+y�-mJ�f��G�A�i�����fQ��z`� .l�V׀9)���ufqm�׸�D�l��XgB���ͥ�JQ>�o�������!T�]���)&�d|��)�h���:�oģ�.$��� �&x�c��w�0z��K�`P��Df6=)I*��Κ���̫�e�J� �����!�M6gi�#~hp!+���_j�#B'�̜�~�w�&?J���l���	Ǧ#�K["%�G���0�f��ԃ�)J,����e�G��Z�:��qUv�n}���yh#��䊤/���{o:�Y��[;�T���nf{‎Čg�4q��:Jp�6�&��Z�w�[��X�������@�7��y\��Z쐩�} ��*`�w�g�9�g�>4[�X!,y À2W0�O}Ƿ:H9,QX��ّ%O$ ���Ek%���s �pA��Ե�ѻ�����z`�.�Ҧ43Z�h}�W��7G?1&d�du��SqT�}��`^�W�:7dU�'d�i7x?;/᫨�W�}�P�
�(>?e	I�O�d8�Y��T�k\XD�C�>���2�]fL�Fh0�UK�r�9An�56�|dp����H^�ك���.6H�?��>���V���PG�CH�;mV�,q�6�N�P�j��5��6� ��0�:f��[5�I 	!���/viuݗ��t����ӶYʿl�|�'\�D-��}�`e�v+��x�;��=ԺD��j՗����Ӛ�}�)����+�&�7� ΂����\��Tu�R�[C��h���DOؗ�}�����l���x-E����]�����ɷR|�Z��k!��il���'�D�׼�kg=Z�����ϐu�E)U�G�6'\�e�1�D���m��]-y���j2���Z���´��7})�9LpI��v� N#�V���dw�����ћ����X��VsA����8'FԶi�p!9��߲ϸ�A���7�y,���;��IgW��-y�{|j���*# l}��QN���������H�*�"���s��v�R��y��PQ|r�&��g�A��y`7��0� �*����V�f�͞3<X���8�����.8m�ᤵ��M�]$8MW\cf��3ξٗ�ά�e�V�+������ʞ���i���zY@�g�scUv�r�y�~�P��|2^�&N�g�Aǆl`7i�0�Ә*�X��gf���3<����ìD��.�?��W�����]�MW�f���3��ٗv���%[V�뙫~��Bʞ�巜���V�Y@�Z�s#(v��$�yY�P�6|�&&gw*A�F_`7)f0I��*H�����f�MD3<����֬��.��a
��Qs�]�MW�f�s�3N�ٗ6����-V��L�>�vʞ�Y�\ϲ��Y@bM�s��v��׻y��PX�|��&�Xg7=A�R`7�80	9�*~���L�t�.��Y|�A[���F��K�qa� ��[�R=vI\W��&�g�@Ƚ�!�݉��yFK�O�#�7]�_��y�n(X9�?C��o��BΜ�̅�E��F�Y��v[�����=��y �������nǡ�R�g�����/��xODM 7�%ޯ�p�ug`sn_�߽ ���"R� o�qMN�����0�I� ��+⇳�T�EP���I�`�aDm����h$�r�pAM�q��&��Q800�=��"�Oq��P5�y�v�\)s6(q�=�!�o���&Gq�� 	B�����̰C32�-Z��Z.��tHZ���5蘝0qx��(�LD�����Qf73�X����%�o5z��-=������L�����tJg�CO�K=��0b�BӮV:�Ab�P¸��Z0@��y�;YSwH�u�>�`��֊��/$��f��g:�uX'�kL����
���2}u�Vd�k���2>�Z�����>��Df�"Qe+���J�z�.���2f3�z��䖰ӝ㼓_��/����"�
�f
ւ?}��P�?\ XoE��P�$ȫ��0�P
�S���ԟ�|�S��h�aG}�΄�븎�r����x�������]�
Wo�:1���T��pI����:��,Q�V��z�ۡ�$z �L�/���1`���%��C�)�2���Ǩ�el�N~"���`I�;0=��3>	���̪�7�9��D/EU >�"2�=>9�1�Ƃ�)�c3�(��CF�M�B�L`���p��"��X����H;FM2G����gy>$<w_�?_'�CD�9^��8[|/!�G].��^_�@�x��O�N�W��T��`�8���ES
@|#�Md��*��g&ɤ����t�������n�U��DͰ��#Ue1�r5�d��W3^�RN���H��u�ŗn�Ā�������S7I`։�ԒH�4�n<��,���E��R.|Be���cR�;Kw�.R���eO2�����G����g7�e:�#�����Gl�M
@:��+�<�'J��_�w�O�=I�/��r� D̛y[w$YV*��-�(��M��2��Yқ�{�*���]K�S�m�#<B����^�F��NX�\���K�[�G�&#��8�����<t��Oݫ0"���׏�[�(�w��)�uq٠�9�u���<�*�#�f${ڕ+�_�vQF<~y*1B�ߛ�QI�j��<vb8�܅X�%�$;3+�&��q�˹�ρ���b�TOW��RrD�����/ܔ)��)��9s�p�Nr:R�XХ����ŀ(���hؓR2=� �;�+-�6uA\a����n�E͕fI�o%����Aj�Y�X	t�%T�E"�l%��!���\Z��M2��l�s���I�*�X��LbQB�/ȧ���'�;e�H�Z��b�����zO�b2uY=�1���%��I��m��]��}��T>�=O�-�7�m���9������
c{&xɣq��c�#��,=ے�X��R>˫�(=l�#�6z5�M�W�E���*¬����W�"8�D_�� ��B"�DǦY��uI�]�Y��h�3�����;
G-_s¤��oW�Jm���Z8�1�s�^W$(M�9��mt���2�sZ����V���X�ǘ2�����+Z1�<�e���m�K�w���FN�T�#q�0�#I��Q�K�7:<��~)͢�G�@�`*�<�'kȎ�I�3��ܩV�V������+�`�iy��ͮ��٪�O�@Ț8��c�������������Z�����Negy2�B��$�B������?��h~����抽�Q��Uz��CPDʺ<�mύ�R�E:16��\��̢ (��t-�Bc��7pc[/I�6Y�r[*І�u�]�w�eX(�l��2jdn��ysC<�ɼ�.)$"�α�[�FI+@���,Qg�*��@���/�V+����fI��(ShٹoK2.�G��"�Jb�Bh�2 ]|wmJ�CsBQ�h��t��c�R������ʁ�J�,���
5��S 
X&�	��Oz=�C�Ev$�~·���s9���d(S���Z`gy,�]?"�3�����IDj�Dv���~���Ɗ��`/��K$�}9B�-d�|��{���k��^�E���u>���EbQ�x���*v3D��.-׺����R�H�nտ�fIq,��|�8X/�R�o	��Q��h���=��*E;\sR�yu+��$h�����y8���F[>�4��
�����:��J��ի����T���:�(��?f�����@��b6����-��� �m��#� �q�M��5���C�"r�I����Vį�������^oO]\o�P8c^^v-X4�2
)$�r�f�W��BEK�5�a�v���ڠ��9Xhq��@�=ڕ��� �1�5)qQ�i��
etiG��JE�)��y��w5�����ౣ��4%��|rGX��ئ�VL~�!Ƶ�$���0&N}e�tՕe� �5�w^1�@S�h�J,\bࣴ���H��9��#������]�$��=+!��_���L���T�dyZ�܃��?=;O%��/�ZΖ��^�ۅ6a��K&�#_	��1���9d+����=0�]@���qrJ(D�O�[#ɮ{h	��`
Dz'!g�~X�g"��[+�I�1)���������0�,��'��ͬ|%�|�}�ل,Qw�7$����:��8h��2�O��B;E��*(��\85~<7$j��Ž\�i��9�ڸ�{�q�Z�#���؋}6]ߞ�V��-�:3�RŨ�	R�ήʴ ;�k�FY�Ύ� �2�5�u���q"�;1��`����@����8�>��=,K��"��g5:P�"���V���S�3S5N�M�Bn�<�$���<�|�F������N�����X��
t�;wj���`�k�'���݊�~�$S��~��cL���^Ԑ��u��w/�0P�"���h���s~s��,�f��X$��[����j��6�jx�R�xe�ѹ��c���Ɋ��У��pq�@��0|O�����sG��s�F��p�zd�%64���<����ȏb��p2gш&)�$G	�ظ��:��ݸ��$"0cr��J�}����T\'�U�a�G��_i)#Hz��,)����cᩇ��4gO@_���l��5�)�W1�tKMc.��F'Ӽ�:�vǵ��2�XG5�e!l�~�%�͊��'?�0eo��d�.���'�x��kD���|1�q�Eo��4��Ү�2�>,�Eo��e��+�$s+g�Ň��"�Hգ�X0Bke��|A-Gw����o#d�^F�0������y<���㇆Bn+Ʀ٫e�<�J����4�3B2'��"�-���|`N�^��a�q��V,n�J0�Gˏ�[v��ˤ�`�.�j�&as]a�{��+*H�
4?��3��A�0�)�b��1ؐ>�1����ֲ�)C������=��\m�$���*�^}�D�Q��,}����<�Wv���m�;}�B�~C�����~$��	��E�s��	e��
Zj��$��p=�e�<�^�n�BZ���+�d&Թ�����lV��b��#�ƃLgk{��CaJ�:ۺ��E�s�������}����)�#��v��q�!�9��ҠO���Eo�@�����������o�^3{V� �������j��6�!�Hu�~O1P;0i�X�5
u/�~+��|�<G~����]�1wG��jً��n�h���b	y.r�zv�ϦR˫�$%�����_=0�\�-��a��������
��KڂUΏ�z:b�2-[c����gg�#�y|X�AV ��^�B�/��{��u���Q�'�}������k_�m����N�ħ�]��1G�;�/��"/��l@�uOIR7�}�GTr�J��HK{�[����V\s�O��:K������Ƭ�+0tKV��ۙ��*��n���N����i�-@��[R��e�� �� Y�Ð��jH�yy�i?�R{��)��`4��ÚH�5�� ΆW`�Cr2�AKF	�7��`� @�Ǵ�X
���qV�B#�l��u�aZV0�QD(�.����@-.�b���Ok	�5�6hj�M߿E-]'�����~4�H�y��2R�)$�Y4[J����J	Ȇ��C�ZA�����`	��G]�X����KZVL�O����u�e1Z֘5��L������S2�|)A.듗.��k�~�ն�Ċ��E�U�h
�f����H�ʭ�iЛR{zi)���4��H8"�����Wq�Cr��AK�B�7WY`� ���X
?���BYV�S��l?u.5ZV��QU��b���z1��.�sA����k	G��69S�M�E-����g��O8�E�H���9R��)$��4��Ȁf�J�W���	C��A˟����`��G�wX����K+�VL�D��;�u��lZ�il��]}��
��S�|�.�"�.�k��ն�����E�VL�h�,�7��2_�z좙ů7G=���,<�:����EA�pd>����_�D�����vV������DO]�&ň�[^�SH#��^�L��s�1����
�	��/�/�Ih��k#[�t�1ꋙa >1��4P�Z)t�j�)W�ZU��Pw�u�F�N�f������DTSz$3٪3ՔE֭��ENs��d'�v�� ZgW��/K%S�zV"_�?Z�^2�%V~�,&b�p@�k�۰�{�6"�L���qu��L�S�'�v�h-��~h�� _DL��kc%�ah�z<g�s
0�	Y�!�nb�e��:+&Bq�|����Xj�w�6=+�=�/�+�eŝfn+Du/!�P,P�Y0�F/3��cQ��#m�B�Ȱ��x����`U�t�8Mϫ�R4�+�-knޣo�����)7	��j�UY��%*mx�P��" z�����+��g�T�lz�s�����Ƅ�Y/tX̋������p��=F�����9��iY�<Z���b~�R��#��TE3R�abZ����	��E��X�0h��/�+*�2 F�v��1%'I>g����16��=%�fX*;W\�u*IqV!���-�hh�f��,�8ǵ��;�Z����Ӯ�v��=�\��q<)O�m�&?����w鲜(4��C$�j����B���J#
�f������
v�:����e0�!�aRC��א�2��`b�խ��R���bR��8w#	�a�9��zj��r�,�J��bb�Y�U^��rD�8�����v���+����x����}gy�l[)}�J ����I�/�V��;~�d����,u�al@�gT/Y�c����l�7�U���R���;�^�ի�����Hd)���5X2q�1q�~�A^���-�փ��G���{�&�K�6����*�Rjb�Lz]���-e:�^˶edo��3��f�H�,~�
�&�s2�+u��e{�P��������WQ*zl�;g��(E��`��`<����v �:�rx�v<R�Y&¢\�f����"�P���@�p���k��]v�=�9`�"����@�AF���}��9�ә5�7�y���{���,>|ſP[t�r�V�9Cr�b����̈���g>�Y���;�'!��/���������%K��-�(�pǅ��Ɏ��8완d\�@V>��q�[�KDN(*����-��PE[�6:u��3rlM	E���o&N�ep�E�sP�A܁�E�H(�����P[��k*�TK�V�Â������A��j�S�<9&�$���duME�W��9��~��%mh;�Ɵn`F�7`$�A1���"���Z���������@
�5�W�Z�!�EDu�[�o��}���
6Z�N���|�dB���u�"�sD^�>�X"`�^�#q�	j�њ�M��	b����Fܺ��q��|G�a�h�	����Y�I�鮁��G
��FT/�>��v�Bi�U^A#������@���u\Sn�X̥���6�,H���Eg;<_��?����
��_�k��eP�֔h��I�?�4�~/��hV�6yb��y�G��%��\ބ�w/FwB�j�L�.q�X����fp��S�Gq�%�J�X���X`�˄C�Dzf�SYM�/����)q�_��1�X�N#(�������y�d�0�|௜�a� �>ltP���P�rQ�
���{]�Dɸ"іE���%i�f�-��V`n�+��(���MY�p�`]�m�镘�zwz��bYW@hn�z0Z��KYlQ�������F8�����ߤ=D�Cr���(�.N�ڛV�Dma�5��g�=�to^D�3�i�0�Δ�xH,9�5�ʯ�=#5�|�nm��cdD2^V�jry�t�<kZ�o*R���WJ�{
0��X�u�X�L�����u	��qY>Q>�X�^�ݫP��~i^��"��8q5B���d�����ؔv儙@Y&�9xC?d=��lXmՏ풊w��TEM�$��5�p�<��L�7Tti♦޾���fZJʝ3o�Н��2�rH|����Ƽ<`xy��ar�d�����_��"��Y��(l:�����_��/�yy�D�R�2j1�ϔ�j�*u���7RmK�yAy��6�9�I�w�;ܑ��}�׹Fܚ� 2�,����衡���9/` ݹc�1����O`��YŁ��'%�=8Q���7=]�4�T�����Gۚ�]WZ�s��Jz���a#%�Dt'��i��+�C
me�7����9`�!�򳕾O�ӫ�A1��'�^э���D8c9�����G� B#���?��ͱ)j�JN��Y�W@����0#v��9Fgp�v)qc"�(@V������1����P����v}��9��_��2�a%?�Jo�m7WON)>�U�قX���i�>����z����\Ѱ��T>6�)K�p�2$���Ҩ{j�!��0յ2�q6%���9.�ֈ�x��$L�O����N��p�y����g�����үV|,A<�&�om��bG�*Q�E�R�u��o c�������6��O�!ԟ�/�~������6}����Eö��L��Һ��ycU�J&���w�.��G'�E�4V�����p�$A�t�mL�.����1�	t]�
]4mxT����[�ԭ
��<:.�t�f��k}��_��� ��f�d#C��(��5e��my\��E�Oh��[+�>:�+�	���l.>�]�\�5�b1��9껖*I�{�M�c�c���qz\��2�z�B/�Av����C>eI��"��^�Ͽ���ݗ�\�$�o����f�le�t
���y%J9窭R��A��z9���*���W@ƫg���^l�q��uj��4ܽ�+2���[A�gnX%�7�p9�i���?=yG��8�-�ќ���G��&��}�k��������2��$�9�H%/7���!D5��2CVf�m�f��	]�J�ڔ���p�Z����O�^J�[
���8)p�}�Q<�oV��@����E�K.�4ȹ��*i)g���u�r�	L�0O1M3�T�n�I�Y�Ь�.�~���m���9�ЈT0�DK��O�-��c>��؄��Hz"[�����(�k��cɗD2�r��`J%���h�!'�Ho���l��X�%�(*/5^�׹���G��u��i@���сݘ��h˳A^�2�jE�������X�c����ūZ�f�MEK�أ��s�N��Id
]��ʑ�$,�н�´��/�פ����E�r��C23G#1aT���䪐x���>�ge�fW��"O8����5�r[�b�U�Q�j(�I���!̴�J���agi{;���|�{�es�]4"hs���xL��Ԡ���5~`&Pcź���滿���D�8��F%��M�-Q�sF��ԥ��ɽ��j�,p��bm��A�4w�O"����!���\�J�j���I=FA�~=��[�!s�c�:'�vD����|4�k�e�z�jkI�*�	u�&���MKo��!.������u9�B
����Xƕ~��� wɀC����|��c/����n�G/���e�|0;�]�nuLJ; ��#�3��{����Ԥus��&�t��y\T3_�$���O^��r{��8�	��9P��E�$�&�/f�e`E�	]-���T�P����,��F��I�0e�ګ���bu>nC/�*t�>���Z��F�M6C���`��aV�օv��/��6po����"���	��"�a�_�o�BK���|�Z�Ԇ�dń�Zo�7Q�%�X���{���(\��ѪɴA�ģ�^��!��s��.zܟPi)�-��ғ��Z�Q����.g_�|��� ���L�<�2���B'�3NK��Q�{�
?"��A��|�@jy���!Z���w����wb�?�]���/��Ȗ���D螼X�[�8�r��GɡRP�V��5<٨L0�

���?7`"��,�L�zQ���(��f��o'�t$�P��k8�ǲ������j.2���x_긗�;�4�->��l�ǵ�OU���  35�W��  8 ��  S�  P���g  j�'   ��Y�  ���  ��3����   �  ��B  ��.  ������   9^�~��K
  =��   �� 0  ��   ���  �s   �  �~   �l�   ��3��N  ���'   3��    3��Hx�Ð�����   ��Y�E��)  �Ð�����M��+  �  �1  jh   �=  ��   Pj@�5|�   �p�   1��GG�>  S���D  3����H  �		  �E�U�Q  ���L$�A���P��   ��QQ�X  V��+5��y���V3��  ����Vj�  ��  �����V�o  W�W  ������P�I   ����  5�������~ ��  �F��%����n����3  ��0���4  ����U���@�   �Q�   �} ������  �v  ��@�_  �����A<�  �G<�t8x�  ������D$�@�@�-  ��T$3��
�������5��   S�]V�S   ��U������M�  �5��5�X�  jh   �5����m���S�  +����   ��V��   �E��]� ��  �E�   �u�   �SUV�5������Q�  ���   ����������  W�]���P�   hF/��V��   �b  �|$��  ����   ����<  ��������a  ������  �M  �V�t$�   � �@Ð������?   ��U���Z���V�	  �E��E�E  P�&�����������  �E��4�W�A�-���AN������i   �	������d   �H�x�����Z   �{����c   �E��E�W�_   ����Ð�����E�P�u���t  �����^Ð�����N������^Ð����Y�y  ����  �M���   �]��   �E�P��������Y   �U�쐐���Q����3p����Y�r����y  W�������  3��!u�B��������   ��   ^Ð����Y�/  �E��  ��f�� ��k����U��QS����^�  S�^����t$�4p�*���Y�����������X���������P  �t$�   �L   �J3�B������������8���2��)������   Y�]������Q��A   �Q�����1�|����5��E   �}������3Ɂ}�E  �����F���~�l����  9���  ���^���������`�������E����������U�쐐���Q�e� �E�P�����t$�������2���d��5�����D$�o���VW�}�e ������D> �ǋ^$������~ �[���P�>����U��Q� �����������L$�������E�e� ������E��S����P�������n���XX�=t�k����QÐ������3x�H|�������C����� P��  �G����   �4  �E��E��   �   ��   ���   �   �6�   � �P�   ������{   S�����|   �M�� ����{   h��P�V�=��{   �   � ����c����h�k   ����  ��g   ��Y��  j�����3�_�E��   �����I   PU�����C   ���9  �C   @�8 ������;   �����8   3��B   +��P   ;EY�   �.  ��   �E�P�   _[�=   h���V���8����2   �h�h��-   +��9   P�����O�5   jX^��   h���V���z   �ha�%hj �v   J��y   Y�4p�����u   ��   �E�   �����r����   j@�6�   �E��E;F�I   ���S   W���Z   Ð�����r���h��b��V   ��������t����P   �E���N   �����3���   �d   �l���3��a   j�Y   �v�F���v�Q   V�������N   ���   �   ��+Ί	�   �M�;   ��?   �  �7   �E�7   X_^]�?   PW����S�9   �� ���8   �\����]   �E��]   �M��C����   [Ð����W�����PS�   ��_�   _^[��1   W�P�����$h �  �$   ^[�Ð�����M��   ��  �E��   Ð����j S�   ���   jZ��   ��3��   �F   ��9�   �E���#��"   �#  =��E��   ��J������   @@���   P�%   �M����s   ���   ��   ����   �   j@�   ���   �u���   �6�   ���19�   +ъ�   W���F�,   ���   ��   H�����_^�4   �E�H������   ;��[   �v����
   �.   �   �v�   [�Ð����P�   �U�   W������   �Mj^������{  �   ���������9^��z����3����   ������Y�   �	   jX_�   ���`   �	   ^[���	   �E�P�   3������������P�����Y�z���������u��+M������	��E�H�����������P�����������   H�����H�M���������	��E𐐐�����E�P������������ }  Y�   �����@��   ������   �����@��������   �   @@��������$   �}�������ϐ����+Ί	�������E�H������u����������E𐐐���M� �������E��E𐐐��3��} �6����E������_+�^[������Ð����                0 D P ^ r �     �         " � �         � �                          0 D P ^ r �     } ExitProcess KERNEL32.dll  � GetDesktopWindow  � EndPaint   BeginPaint  � DispatchMessageA  �TranslateMessage  � DialogBoxParamA USER32.dll                                                      ���i���Z7B	       P   ,  uݴn�      `   @                   �   0     "����!      �        �;��3     �        ��鄔3     �        ��^M�2                                                                                                                                                                                                                                                     cyW�ҠZ'�	   Va�i   'B	��Z_aW�a�i��  �   ,4�8�8�8l4r4�7�7�7�7�6�5�6�5j2?4W4�2T8�9Z:�5h8s8�2�9�;=3=�=7#7)7�3�3�3�9�:;�;^<�<�45#5O9.8�3�3:�:�:�:�:;$;�;65<5�4�4�5�2�2d9j9393                                                                                                                                                                                                                                                                                                                                                                                                                                                             V!P~IxCr=l7e0_*Y$VRofbdSL{Fu@o:i3b-\'V$ MWL!P~IxCr=l7e0_*Y$42�U �;�|�N��N�