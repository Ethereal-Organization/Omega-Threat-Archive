MZP      ��  �       @                                     � �	�!�L�!��This program must be run under Win32
$7                                                                                                                                        PE  L ��%G        � ��        � ��
  �  �
   @                                      @                       x�
 l   �
 x                                                  �
                                                    CODE     �                       �  �DATA        �  �                @  �.rsrc       �
  
   �             @  �                                                                                                                                                                                                                                                                                                                                                                                      
�)ۻ�c��
 ��  ,
     j)J�&^r��M��,�M^�����%!�q{����1��S1��Ili��|�,������pB�qc����=���c�^�ͳ������ ���N>�v���e��h�4�ڬ�����u�#��u�d�C�i������+Ҋ,�k�$F?�g�J#5Sa��������mư(1Y�i�hs�ܞ^�����ދz���>�]�I�1.�=�*����N�H�i�!e�:ǐ� �X��̀�!O�δ�C�*,����ug);�_������fb�����ŷ��=F��.����A��w4^���������q>�� k,�=;?c���t��z=�\�m���0�_a�P�:7����گk���8�n�q��3���_#ġ0���1Ui�}&e#j���{�C���:l�mL� �Nڃ���t�(�e�:3�"W�7WZ���A��N�][`� �G���ɏ�.���'��~���`�^Ɏ��[��ZZY��Y�VKk�ĵ�Y�E��V��jF%�&48HP����-^Č*��[�9ѢŹb��E��i.�w��(�l��xu�E��.�g���6�49��$Г+h����B��Lλ��꥽�e�0v ���"m�9�#�[�^�./Պ�1Ѿŵ�?m2��DݗBuC-����7n�!j�eȶ�T��+XZS��V��lR-��`�%�]�?��f��UȲ�.͡�KfGb�|NE�~Sj����������<�g�J�}gLx��p(>:�8�e��s�1�	�K�&1�>��K��x�2N����C�SSDy��GE>"�-�ut����1���|)+�4a�jˁ�ǋaT���;C4<~x-e�ǳ/�6��8���KW����ix7֎%�8�4�G��\iX������y*��'��,Y~�K�潏/㋼C��{́���E��9��-��wŬ�t)_�.͌x��S�p$Ig21�Z���-K�;��3L2�&����u����Lz��I1�/�����@�/.�*
yȠ
~�j����y�~��u�Zw��C����W羭(3���������|�y����r��'��|'٘<���V��>v6�.CՍ詧[֚K��Ȋ�Ά��v��ԡ�-��-� Keٷ��yh`��a����%h�̞���L�܁x������	�+8���P����5����U�t#'�_�*�
д��O��!���@���X��2�D��.���3���:������8�n�6ݗmۄQ5^��q�Q������I��"��wco�9����@�XҜL��q[�Z\�q�CAG
�ucY5��o�
ǅB�3���fS�Ý��U^7��MyQ.k#���iot&!���v�
%��7}��}���$:�!���z*ϛ��m����7d���ed��ò�B;r�GD�{��ȟe�-'zZƃPW<N�1�u���/�nSzڂ���7�\w����7%h٧6w#��[ ��m`h��(SL���?��Wu4�,T���]���G����i��m���!}m�W�r^�����i��d��i|C*kq[�f���B��ٖ���V&%�a�/�����߃H�M�:;D*_�0O��hnZ���!�ձ��G(q��H�9X�����%�Q�Rt�0���S�;���?K)b�[�|o��F�vU\�R�PS����f������������ki�TR��˿���^
ƀlg��g������K���!^e%L��SQ꾾q�^�_��Z��l�(�/��,�I�Îf�f�|�V8��sNw�:�{'h��X��l��ez#b9�{����P���S ��$�������S2�����8��f-��N�����2��̟�P�IQR�� 
�1���T̡黧M���/�mP֏n�������v��FE-�"5���(�֍��#�b���|w8
u��j<����I���b�y�O��v\��}%�Vm����r��?aζ�2qDtl�[�<w��/K\�<i^�o3�U�13gXwQυI�6B���(#��C��Y��B!Rz��K:�gt���~��ݗ�����[+%I�=�?����[T@ÈK=K���x%1 ?u�n:��M<ŉ�7
10�������&�U����/$��pj����P�^��{[�{�P�F��� �;�μR���i"�I���C������)���[���'� ��$��"���u�w�R�!�%(J�^��-��j%�1������!]����[2����&�̀��M�#�^��H�fVf��j�f�.���G��$W~�|V� _N�>"��۝(��K@J��`k�b��R�Q&��P�QW��t2���^u�������\MQے�:cn��&Z��h0z�E�F�#�dY�!��R��;���-�>�o�A$�r�f-�	�^!��rI��|*�)�Ӌak�-w/q� u�����8=�͟��'18�B1��^&��u�;�&b۾��Ĥ�W�#�q@M���F\Ÿ�ʟxU�[��hD�%K��e=�P��� l^������}���?�|�M����U�Ps�����&�?�=�uy���w*�)(��v�U�3z5�"h�l�������O$=����y˷�6�(#^�xҊ���ڐT���\�do�Y���Z��_اS�<(���c�m��X��eh�78�M�K�`�'�A�7������W̠�\~ǹ7����j��I$�Q�Ҥ��jL$k�dC�6R����� ��Bz��Ƒ�|����d34�㡦q�
�ڣ-(J���S��:kem ���>��u�̟�-Y�-��"�'fV6�4�dU�v��I�J|�>m���S����z�۸����A�}�6�~��)gs���|T���0��ɪ��j�#���E�����P(F_���R���=l�o�H���CU��u�n��,�ַ��?f��LV��X���8(��R~љ��ӵ�aUa�|�R�Z�p�=��SB���=��a�Eq�FO�W�ҕ2��V��"
����P�<1VE�-r�q��V�]��(63u �Z�&���ЙTS::Ï8�,ǁK�g@�]_�\[�7,���\��RV����r���5G� �SX���I�d���\���L�OD�IQ��#hn���wY��ޑ�E�z+ �.|q��n�p=&)7��d��v.][��ԏ9#FYQ0Z����fm���KO
g��Q�:Zj�����2�S�HT�7�P̎Im�Ho}��,�q$l���j9>���!�#���=d]6��eb Й~���Um�+��ƹo0z~���ז�
[��-/���K��{�^��,�hB;�B�����X(���536��ލ���h
�O�"��qzF���}���i�`h�M�$v��G�{�#�o�H'j��n�K�^l�׾b�q�+����Mߪk_��S��(VM��ʩ�t�����|�3q�+[�(��qVn���Rd�g�4X�{����KbR��wƹ�b/=.P-���UG]4�;���	����l�y�[�
c����|^���jR�_υ����Ȧ�Ɨ��"�����#>W�	�0;[��k��[��44��fA��Z���i�� hR���n�N1}����#�'�v]l��j����V��l ����N��;�>f ��O"K.��3���?��$�h�M���W����pG���N�5BW�\�2.�R4��t[�ɺ$g&��:!ۻ���_�%�� �+B�H4��P�n��7ɗ�D)�a�\�΋S���A	���
�:
����&�CZ��fӖ��Oi����@��2�͜l��M�N� x\;9����+2�0�ڨ���,f��8����P�4���-�?��R���c�>��D�f�_����gjU��U�r��O	D���2�v�Mv��nv���mx���0U^����׳��t�A3C�A`e�΅Ų'�3Y��	��\07�B�����:6ο�E�n�J�,�<u�W�Ymhe�@Q5AqF�/��DB$l���?�n����^Y���-*:
�Am��/�t��w����ͧ���9O�?�v��*���5<�X���f����*汙��{��R5}�׸�Z����1A�M�*q)Sڊ�p���ޟ�U#G
�˖)��ӣI�sw��d��[?=Чr Q5�^�qc�+�z���h��Q*��uz�%��[8^£��b2n� E�'!BF|�)��5�f�
h�w|�c/x��T��������+3��s��Ÿ�7����R�����C2��Y�ώ����-#^��b�~����E� `��A�l� _y	ufφ=��|sF�K��R�#J�j�j漘:��o%=.��x���}����G��.l_�{t�u6��ݱvX�^r����=�n�V#���\Gl�2��Q���xn#8��%Z�ݞD��M�rYEe�G�t29��:Ԅ���z}�6�Md�Q�Ob�!D�m~%�jB�����M@�h����E�yo�i"���q��X{�mͻs��L]\E#��3����ꟻ�9�v�P�D�Wwg�lb���%!�E#�V�U�3C���,=O�Gc[3_ʇ�,�O|�÷Xnh�g�X�~�5����#�S��?dʊҕ�.Eav��c��Jq\�˷QV�]��hӬ)f���7D$P�%�	���۴@�?ʌQ�M��y|����o�@�0�3��Gu���!�XI����龝B���7�?;�I�K�7���N��29I�d�R�c���~�����nг�����A/G��}+y���<�BFjT�����卒*�D,f��3;!�?����qu'�+Ÿ��Q�s����Wtt� ��~h���/�T�f����?բ苌�'!Gi�1e�e8tg9Oi��Vl�ߵ������kZ���@��=I��r�6tf]��@r�?3�j(����\*��v�{���%�P!��/0������./Gƙ�o�ft�(>���+�c����u��fN9��sl�#�\�e@��S7v����>v/��K\���NyIn��a@B3���̖R�Ѿ��{j�%O�a�i�%�8�<477�[~b��J܃�� 	�2��|ɍ����������Y���:�>M��V4٬�zc�;�{e���x���� X�,�QҕQ�R�|x�l=�H�Q*}[�+�~�zsl�)b�$��p�Zm<*J^s��0k9(��y2��_�9��-�*����3c��/N��Mmj��^���;��'�h���|�3�o���٤�ط�l��Y�;�[�OTU����'ã��U>1����hZY*Z٘'��:e�J6@ҔcUkj����!����������F����݆�)ꆖ�ǃ9��zs
���VÑ�o����<2����SU�8�E�� ��å�yu������L3xv��b�o-���0�[X$o-�=7��f��[L='��mǐ:�F3��jo� �,������p��gbf����H�6����.]L;����LN��XR�֯�{�h��$�I���ֲ�b��Gx��I]f��Ydx&�,wF,}�SlQP£B�^�wuc���
�R� ].�dbMJ��ڛa�3p�f��@��;��|.3�G���}
|�CzOa��Z�;����|ً������D[:aI�-��Gů��%N��om��#�6/x8fw��s*���_���$���p�<�Ф�뽗��l�PBA(� n,��t1��������+���\\}t�����M^-u����g?"�.��J �x.���8�\���T��E/��`�J<HD@X��Ӫ�^�؛�섰:���B��s�:%��sF��V�uk�Ջ���w�b\!S�u��x���g*�)Xr��%�a�2q�X�l�5(1�5ix���0���?4Y;�)mڣ�����qz+���U;�FB�>�̠�����Ax#��F��7�����:[h����ˊ�����KE�kFuz�j�H͐[h�ٍ,u���FB����%i�A`��vT*��B�K��r�[�@fy�C�n�0����N^ˠ�<�M�\]���*�,��N��&�b�XYZ�:/���&1�=��6�5Y�1�8M��Z�+S��\�L�y�d!��}be ����G�F�e�Pڍ�E�@Oޫ򞂭���C�'�.4�������%j-q�lN(O;��zӒW�m5���^���� �dFV}��,{a�Q�����u���o�����T;=�[���~BK���������C=j'G��u_�7��[�0��n�s�đh:tP��:`%5fC oV�P��Ĭe�;�n~�+�(�?��߹�2��"�W������>����HwvT�(�R���u�S���&40�6�5��ZM�,d�V���rz�ΚdS|���#�ߐ3?�ZL��+��M4�g���k�d�� hKo����t�r��FD��/(��U�;JuQ7��e�+�_}�e���nY�8(1��)�;4�A�z̫��~����w���Ԇ���+�W��hs-���tn���\�5�Pۘ��c�?�M��������˃���6���m��K�vn�*�r��F2mR#���΃b��o��[����

��]�rF��f�;I�t�`�]aÂ�q=bz���W��o�bհ���Ƀ,���1/4ur}r\k:��M�����N�-	4�k���<wڍ�7 �����i¸����P�۟:��$7M?Jf��9��p�y	�]t�7�dA��r�w��Ԫ!I�]�:�^汆1���̵o�z��,(��'f�f�	)�Ic��������������Y"��hOG�Hj4��dX�'����U�6�� L��iL�'}��a��@�쾴��gk�0���l��V��D�hh��R����k��Y�&ې'
���/#��\�P�1:��\�W�no/�b�ɏӂ���{�Z�q��W��yM�ˑvy�}�[ !���ʩQ;ߢC������S�[�Z��֠/�/��ZĞ7��o���
�M� ��(C�F�w�����~��>�3\4+�#��Fs>m�[zGA�gz������#+�1IH��
��ͩ���r׺�4wg�1�r�>hB��T�C(F8�d����E��p=l8�?�7����U��l�`fD�zT'���{t�
_`~����vU 甤�i��� ��;���k΅�O�ʄ�R���J5f��,��@�O4-Y4v���y���.����~�on���eP�-5h���ױ֪-��E��B$���O�[Afdz���60Rw��@|��@��t��ǘ�%��ngeE���,�J	4a�I00�U�)�b���T�j&�`Ki`�R�wn�q��}N�) ���3�c<�+U# �X����	��-�c��z�)RZw#>FN9�<��.�3|��'ǀ�fI�#Y��x��6�lY�aףӃH%;_o9Zy�
���K����.1��D�\��޶Q�P�M���y��G�k���4xG�彸��f@�
�S,��_�Ŗ%��؋��+�dX�s'�c�z��$������������%�%��'��C� 9)� /��Rlc�*�|~kό;�c�=�/d����))���q���RC{��t���x��^�O��6ז�d�e�7��������H><�k��&ѳ�:,��|�-��]������=��2�\�QD��6yn3N��T�·�NH�ɯ�3���߻.��}cr'K:�?Hv��ѯ��_㟻��ι�T�M1�S��Зʮ��E�,��̥e�k(�(�����pC�|V��xl:�py�g�����"�@�7�^��Y9���r�{2~���d��5����>b�)������:�7��}Mu5≠-r�*?4@�r?��P~�b6g)x8��U�?�̐AA�U���B�3�Y��Y,���GfA8��.:�>|���1}}4�@T��[����Y��^.�p�x�h˷��Pr���n�X�v��L�>Y��dn0_ ��e1�: ������_��*F��7rH�Z�+���:Ԭ8��i{�"u�F������Yb(���22e���O�პd����Fl�I�3b��;v�3�΅͞f����#H��Ӫ��e�F(FԢ	�B �-�l�^�����$�����18�򁂐�yA���ܴ�@VNSt��u�6R33c~ ����К˽M���j%��{��Yo����*�@��`�:������-�T�ϏN����ɺyHٹ�j%ƣ�6 �_q��A!���1^^��V���Q( �[̧4���K�[ ���2�ޯ�J��K3%�=���� �-:b��r����E!f+Q���³Ͻ�,		�T�����!��|����3
�қ�¼�_�y�x�+t�S�jn[jQv ���_n|��d>=�����E�ew.)�^ڤK����$qxh&xC�p4����v:�0����RXd�6ы��?)^͆���C�	�j��}Ї�}�d�&<� �$X�AߐV?_;@4'�;���������y>=�6h���IƼ@�:�ť2di�.�w�����{���B��Pg�-;Y����:�+0+���
Uut?C�l�x���cHΚ���0�*!�ՠV�����o-�Ƹl+cMF��<��i���_���:�xi��O��O�˹*��~郷$�g�X2�b�1կ�F{�Lks�
er����+���w 5�TE�ğՋ+͐7�R+��T�ݢ��Tن�hD'؇�wy�ߕ������%��G��������d�n����P��54o�������Wu1���H��� `Kj��`�V�p����N��AG���hh��;P��,h1�Ѻ���N��~e�qiCN |� �T�]���~Д�@(�"���al;1��%F,����yT����)�����j3d�	�H��&�"�s�v�L�Ũa�Y,�@#���o��	@�=�J6�
�V:X!;HL���(`ب\1]j�r�
T`�2}«��K�L��M�錧��2QN#�{	dLˤ��t.�m �m�bₙi�aj���U���jC�yAS ���������ךT3<0T��.���b�����zx4�2�����?=�~{�<9 әum�8�'����GO�~�\���RE˗d��ߛ�����%�2]#�E��6�i��/>Q{7�g��-J�z��Ğ���m�QP���h��{ߙ��A�+� -LR�>��N�}q�Lj��MN̄�-�7�&W���\B�,e������s}[Z�*���PJ���w?ng7QG���y�5#݋ǃ�f�Z�W�LL��higX|M��L4���p;����x�D/��=ߴ��W[����P� �h���6���+-���}>o8�E�W}�x����)��ɂ���ԒB���$���-��Y�RY��8ۨ?�5�i^���x�z���V�^v8���4�O��Ϋm�6��ğu��Qf(���n!�o�����b'�7���ı��"3�e'�&�`�M=���hxo�������D}Qx��w�V�ɦ�]-<��.E���C�3� Kt��Ȁ
����r�N��np	��%D�=�>�,�	JlT���%-��h��	��y��ѐxm���'t���?w�+C������	I���}M�A�T�)��z���Ή,�
�\�-��D�:���Rk&��q�ė�[z)���,>:���{�r�+;��Z�l�����_ *F�rBd��s�S�tk/!�E�-9�!{z��UH@�PUz��l�Z�⼅�jL<
Ti��d��0�� D�&#�.j���)�Z�?�`�7̗�u�T>�Řb�]��j�\=$�\�-E!_ӐȺZ�%���G4O�5������wf�1{⼱�T�ҫK���=���f��=�w��0��|tV����-��q�P}ev�_��y�!����t�[>��x��e�ͯj�Z8{��)�5\�L9d.��o��*�������c�\�t��F_�5�*���b��E�f^:�Eő!���nq�i�jHI��M;ިPT�V�̳� ���or�7��W�x�e���4# <!A/�㸴c�^�j�m���>�F�Ӫ>e#������1�䷦uxX	X�5j�X����[Q,�p�T�ބ��3�Rc��ES?�ݖ�>��l+m�k����9oIn��"6����W�t��(sB2%��:�,�<�.�����A�)y��y��W�cfK�]�`i���D��ĥ�6�
��D��uO�J�g�/�io:
���>�{1��{d�9N5����h߱^#jN��r�8�s�^v���j���|"s�O��}�'F<u�[��-�T� �2_d9ʨ+B<���ٝH5=b��[A�<7}��˻V�|����&��sӧ�q�x�Y)5�u6��q�n؆�E���<���Q�M|��9�; 7��Y��1�h�U't����$F�̐��t��<���x�#O�p��j�	��,9HG����A+}�dn]nˋ5��vهA{�;�������U���!D��f����@��nk��v���{���Nٮ��:Cf����Z.�&�J9��_da�?hb���U�`0G��R$N��v2�=ލ1�̖��EUU{ٞSM��L��
��g�������u�Xy4�J�B];v9��Z`����ۆ�FTC�`�S/��(&�;1e�gB%K��+g�'9q�v�[4P*e��-�i�%lȯ S�Q�� ���ܗ��^�GZ!�h��ԡ�5���ꠙee��~��U��W5I����Mԭ��(|�����D��C�v𯖁4�g_ZY^?)��X�f�.�Nbw ��"i���lv�CN.Pq���x[������{�儴z�0�-�3�v}}h�Ho0e#P:���8�Ͳ�}u;���?���*t���*�V����o۷�|/6��&=�����+m+���}:YNлޛID�E�~~Y���O��>/U�,�iE�׏����X�Һ����
SU,앹[�<��>���1=)y]�[ 7�lŪ�|�[V]�K��?̓Sa�`�ה�g�@��qg4���+���-�_U1C�w"8�oE���G]�"��-eB��}M�Z�*�Ȏ�v�9�*��3�^�:��������H�)�P�L:�U��~-�s+#ܥ��%�`.��i�zl0j�1ؚ;�\��4=]�	�cF�b��3B=���JA
JqGn�����*{[����� ��;ǂڊl�*Řk����!d��:���&�k���<�u�e���c�9���ڤ}��0}a���Z���l��F����/C�Y�+4Qj�$��4�J��[@ m�y\����p�)��O<D6����B����\�����I<���V�P����d���A��M@U��-�ã�9揂�L�s1���"���X{������Tp,H��	�<ޏB��Ņ
���C����Y�>#��|d�_X՞�tũn��+m�A�I���6���kf�"r�#���y17r�\r��K�Gg6�/im�wj{\@O����ea^����h�4�<�^C������@�Q#���4^�70�^��O�0#�㟖��$�W����c�0�ޭi���Jp��f�̞�7�;��|a����~�ƯO���^p��&^�Ty?����(��߿��$�z->y�X�p�3��1��!U���D�Ѐ�ꭙ_\�*� 	�
r�'c�'�m�[q��#�/u��߻_}92C��%~	�%Y�n�*�E�ͳd�/:�5�6���q£V�xߎ���"_/_��jc�2��&mF>�vTΓ�Hvx����\+�DI�sɈ*4l�������Ji]P��cա�M�g�-i8UNs������P�\�?ܙ�w�@y�� ��|<s3$�4�*3k������AϮ�g��'�z��h֖�89.�^�H��]���(8&���XtM�&�VwK�������o3b8�)�|����aTLqJ�*�/|�*gB���7����&�,����[���Z�?YS
�S⎑i�r��M����y�	F�*%S/�bU���!�f*���	*�޼N��sUz��@�����)���eA������5���d�^wNο��`���١��5�j,.�9�,����h�俻:#N����Бȼϔ�(�,�W;Y�6�`��_�B�z��$�cNyns)B��F��,���.9��t5۞� ��VT.��Վ<檓��N'��|�5hIU1szU�Ĝrƚ�ZxX-^R�0�ݦ࡫;����|,�eH���7g������{��!�+\x�@Q�Q��x7.�Mo���e��@K���`�*F���G'��3t�>[��3O%������T������	^	�cP_����k	ܝ��`f2��b�\�w����Ex<�V�'u��&!^pϋq �ՆomUﴅRPb%�E�����!h��y���,�-�,��{,��7 �p�0f�9�ȹÙw�c��r�i�<��d��Ҙn����?{h�=������!�Ͷ�+=cq����qz�P{��
��q�7��\��@�`R�,������v�c�/�)Ƅ��=H&�	��1c�EnM\�l�+�z�ik�>A��B�Y٥�X��Fɿ�¾){�z̻#8��������+���ŧi������N�ߦ��S���o�l�Q���U��}�6��?��F�$���a�z.��yP���Ͳ�s�.��	�1ص��[���6�Pz
z%l�/1]*�]�9�ZP[e�$�n.{3f!�,�y��_��?�}���h�Kk��+���%�� V�|�
���e�o?�fvd��RX��Te�u��{nW��uC�lN� �1PY���I�9�vJ"�q��_W\a�ؗ������Yk�8��*�ЅjK��%����0`yI�ȉ'N§�t��<~yb�M)ZV�u�&���ƿ�)�>W��Il<f�A����9{�pAoY;�4������ݤ��(��-;���eg�
��',eπ�@4�������eExU�C���P[�:{6��Sq7�/?4��ﰥ���hq7�h�k�;���QI�z�}����y͡� �X�U�)*(�dz��oӾ��!��_�#��u���� ��d0���l��
$����U�U��k�"<��P�z�����_��a{Qq�w )J�)\E�K�tq�J�U�}Ő;�w���/���`_?��@�24��,n"d��QЄ�K���#Ǜ@�p���u+�D?<�3����a��R١a��R��be6��zd8l(p��%�Rw*z.� Zc�e#lt}ҳ
�U}�H%aDW�@f���.��I�'��bݥW�k2�d����'�e�z�9xV!)�uR}�g����#	W i���4�蚺G7�P���M��P��,onT���+K�TO��	{Y=�o����R�K���8Vm��*�$�^42�`Б�����Y����/�Ƭ�X̊o�Ŷ��kAU�q���M1�<�c5�n��B�}b����*������lJf"+I�N�Y�sf���e��B��A6Z�#����؏�ֶ�Rٗ�fA�Q�\7Ǡ9�W���L�.�q�_Xla�5-��-ٸ��0�>�#y��8�Jb4u�4)U玝 \�d�3uJ�* it,��6o<��7Z�Y�U��3�����\��T�1O%Xt�v�����ٺ�c���\iWF��`�;W��@}�Hh�g�mȑ&}>�6�*��fq~����O�T��y�����8�<֊5tk�z<ET���@k0�e@ OL�&"�w�D��I��w�����o�"�j,�=��g۾ŗ{9�^�Xk�q��.��0
���m��i9�@� ��JP�rAD����V�3u'q����#���Ac��TC�]dc(J����L�_����#��t�����I0�	�.}3	�W���v#���(�A���q�<R�#�}�K{rTt�K���t�0}�SJR�B.p�Eg����Z�A�C�[�7%�y@�UA�&M8\��׾��][��{�I����FT_ђr�J��.����@��U�ؽ?�Ș�._	h �|����^$��L��� ; �B3��ģ��/p��mj&��ba�y'��[���GZN��<�CF�N��t��wC!IJ N��w�O*�6�d?�F�=�l������|��Mn��6�>�D�J흷~Jg��q
��4�w&Ձ!7!�TA�X��LJ�~SkN���2t��:DƷ�\U�5)�d���q�
�s�u����e��"�p�\u���c��^���|ʃ�7�<1˳X�}�k����tzC9���>����xv���l�AN'���]��y�$��E*kU� m��x�\��3�N�:��H��7#ߗ�H�s9|�C%���q�����d~� ֳ�<l�E-���R�C#��Gҍ�,��~jr�bсff��#��l�\�κ����@^.��<0c�vtc�3�_��[T�&�y��3�Q�}��.Ưan���*t��_����o� p���l�}����[�r4͆�u�y�}�c|n0Yo3��B�G�<�wn��uFΟ��m���TX�5c)y���l�)&�ϲ��-�F����V�]�'�N�%����p�,����"`_��С���<�fOH?*T�Oл�Le�a~�`�8���0V�����ᝑ������O�[ӹ
Y�wj�	0��Ծۜ��9���S�Q��O�)_Z�=���Eiʉً�%��A����i�R�"cS�9��|� C;v
l�a�r_���5�Qgu���UV<�Л���yH��'��޽���!�Ƥ���o�91qC6�nx��c�w���ʿ��	��CR�����r����U|�f@>�:��e���* }y߷գB�S��`~�WQF3��o�!��"��ݖSha��g�uX�hQ3��!K�`vWZӗ�ǥ)��}��_���u� �G|��2_�ԗ
^3wf$gjዐ��>q�D�}�L�* +t�U�z�H	��bVVp�,���������8�谆�����_(>��væ��m%di�Ь��c���mY�)�p�3kҒ������x-���.��/SE8Eqe��}�"�A6s���*���7T'�KW����J�-hRYR��d/�4b#�)j[��P�a��=;?9`�Lϭ2�nwhP(-�0�3���?�,x�(6�,�^(>���;�EQ
�-����g�L�Y�h�X��7I�Z��80PL������� �Hn�a���5b�B��.�.�V8�A��[�-"5�H�``��M�	��,3�T)��uͫ�w0"�ӟ<UP��{��|����Ύ"�V��u'k,���ڡ��V������	0`��+�����7��F�&��1���!�.� 꽩6��!u��cgwjLU<D�o��@q�^�e"�R�i6�H���qXtf�>�����i�̈z���!0��g{�����Yz�vr�Q{#ǯ�������seu$��h��V=�mb1��9�dĈLQe�֫��l.�B��޹n���i��y�>�!��Cf�%�6�.jzϯ��yva�j�K��:�YHX�2@?7���X-i]�gRb���*��eAxnJ��Qi�J�^4���3l��a��*)�9�
�ͬ���6���u��E�7r�<s�A�V�=�=�)���H<5l&,��I�\�T���}[\ڱj��"k;q�48r��N%%�j��'��#�e���r�m���ǴP^p��$G���gHF��h{����,Hz"�'�|Մ�lH"l_\] H݋�'6C6 �"��_iTo���]$6��Ǒ��}�XY���F"�u>��x]�
b:��t~yrh�2����z����>���"n��2��/�?�Uv'��l=���ɶZ$�_WD��V
�^]T2|O��C%Eu��@Y����PsZ0#������
�[\�Ֆ�v��!& �P#�'��W�}c� Y�O�!�R�|��e�>�m�
�H�!k�$D(���tV��s�pU�����MS��h
�da`���L"��Q��ϊ�>���R��f�;��	(f=%�5csJ7/��E����<���0��D.T��u�\��i𗩶ET=O|�EL�Eu��/�bwL���#r���
��8y8[E�J��C*1��e�k\�Җ�$՝��٣�=cP ���2rO��|���%��+F��ۋ0KitF1�u�陯0����p(*�MW�.��X���!�'�}�q6�FJ����BЙ��-�A�߷���G����������dP��FW���f�4�b����px)�;W��~[R�8Ҕ\�>J�2.jk�{'���Ul"͊���=
'-�5�f��6ZZdU��n*�� %/��(�����\K~��|��m6ܾ���+�nÿ�LDi[C ������)�4��h[����B�.>�@�o`��y'g�̺6~}0��c�;ZX���hr��+a��o��-Zu��>�g�?E��p�H�jÇ� ӂT���8gJ�Ш�g�/L.�9�S9j�٨��3���@H���tG�
���R�����h��B��@�5�Sځ��Q�B�R��N[��f@&]G/C���:+w��������Uu}鼉�s6jFl��'khvJ���o���G�Ea��@#R�aV���?Ex.��u����Z�:��D�{�zS4�Ώݻe1��S�<5���בâ�l{Q�=�?O���?��b����)��C���W���b����q�f�2w���<e-�ᤅ������\���L�����D�J]����s����Ǆv��9�ܰ�t%��8�Zֵ�Zu�����@Wی��"|ʇ�����𒰙��P�)j1P][�R��Ք�
��� �"P���O�5���幣=]W���Ѩ GP�\5����q��̸� 9lۧ��/2��N&AG2v����ɍNBlБ�ց���{�㖝a��w�ǔ�8<���>�޼I�+����K����+��i���n@��iV�$Q��Xr��^���\Z8|]���{�Nހ�܇zfד�0/�1���)Ks�4F	 &-���3%
!l]�g+���e#N뾚0√o7�q08�Ё��㞟��ɹ ���M�5O�B���w����A"Yݽ�N����San��U|��\K82_R������=��U�%��]ͻ=�;������*{fxm"&�N�p���To���XI	սO �Z��ي���oE��w��8�,�>LC�����ǅ���R���s�:����k�+�}\xgO��"��+ �0�Q�Ļ 		H�㞂�l	S�.<��V�md�F��U��;W/���ȅ��]�U�5�����V"{���غ'�2L����!��:�%��ʘ���nmA�{�5� �g�Tv��T�gPI��M�_iT��D��ϧ E�rxn�JT{����v4�$�(��dJb�T��|�i��6غZ�
ꂑ����TXi ��D����,��<�O�ת�k�a&����h9��q(Ac�xN�����B�*���D���F*<�2��� ���I��U��;J�䏒]j�n+��,���u�M��qрH�xj��u�f|~���͕6�kS�B0㋏~V|C�.ڲ�`�}:��Š]��A[�7P��[bE�"K�3|�����Ƶ@��" l��9��.��kp����9���|%��) L�T  '��96�L�2룑��o�8��=�<h���8����V㇟Ӳ�i���rfY�H���x���g�#���uFu�{I�z��'��ʝ���]:�#����`���!u�}↍l��e��M�m
s�x�AKN�ȟ0m��k�BL|�w����/A���v[� U� V�ڋ�ܢ�LGI�kG�|��ɒr,^X��dC�|}!���Ѧ�]C%�]��'j�L�����q��A/��C�_��>'��f-%��9�� n`{�SN0u:E�B`H!C���OB/��d�8���iF�={��%��+�kܼ��8��9$�>�3M�����&��j���z�7K$�� �*��ĉ|�����8̔�mȈ�l:��;�5_:���"�;9f��H�a�+Ij�������K������@��+!���w�JzP�G�ܪh9���xOX�p�)a���)�R�I硗(���
�����ܩ]�4���`L�6hEv�%jI������i��q�������:h��M����
�g�]ۥ�a�d��d�#��su	)Y���\���PA7�P�h!������'�$c[v����]����G��c�2�k��|����K����А���Ƹ�����\���n37<��ګ�Z��]�aq�XJC|����5��X��U��d��̘��P����
����!��������GJ��3��=×l&��(���B��69���c	R�Q6���8)O�h�ʛ��?yJ�T;t�`�`�u�}E�L<PY�߱�Q��϶?%kɩ&�}`��z$�[�N��h1i[`�KpfɜB���,)���\Qo�]��"U{�BQ���o�?�n4�4W�L\"�����g�ɏ����yS�e�9�J�$^�5����+�eW��u@��*$hL��*gB+���,7e�����ۍ�\�T֛3�n=��ň�湀A��l��{<��&�rL�TNp�ҧ��<���r�` �~�V�%؉ ��F�<l��ei��(�X;!�G	�$���oR�@�o����5r�t}�'�+U�O�V��]��7>xݎP���豘D�W�c=;+w�Y,$��_$c�gB
�xd@A� �>?���!��F���;J5R����<)�,x���N(�1#��:�Х~%gEO�;�||}��(8/�c����A��`:|_4���/�D�h�����h$��T�d`��d]��ZW�a����]{�a�	�%=lE
��F�q^1pKj���o�'���x�T�/��SV;���Y�X�>�W����WB�X:���o̎����!^�� ��݉�3UHh4����J�&x��owjS�g��R"?�<�2��)��R�m�R>���&5F����]�xpCD�OC
 �[�����i�j������.0�N�q�׷ѬZ�Io���^�.�|�sk��Ն�V����c��,T3�����6A���8R�hH��3��s��R��?�7�-D��l��wċC����wW��tXӖX��}d�vw��<�Z���Re�V����1��r8[� �U���:PFy���V���L���da]�@d`�oP��(%ͥ'��ɟ�3�C��MU�S�9��M��O�Y\�s��~ 3�R�A��b�5�L��ns�t_dD`�Ԑ�L�HW��񽥆μ�7��T~�U��鏋��p'�..�6��a�3�m`z��MA���H��#�����9:W���b$QU�S�J�<�O�K_*{30���6q�ot@� � ����F�����$!�+��	1�W��4���G3j��Qv6߻ql�`��c�#��b9�k��x�1z{�r~�;�[H���WHL��'��ڔ�bk�xϜ����M����:x>��7�`K���[�<�˩�� 
zst{�[�O�
�J!�2�Cv�G�x��4j�$�}�2�G��_�ٵc��/���SX��SQ���`3E?hy�d{�mk�E3�hޑ�kH���Yd#��ԯJq����i,�wj�D/h��[F<t"i�Y+�.�|� ���6c��� MO��NM���p�"`k�rC����Q�Et��o��3��gk4g�1Ը�R�Շh�Aq P����q L�M�@�M�?�
ym>�R�6����*[]��r<⚟�Ҋ&(Ş"�͋���؅�8���[9�m������G݋�֯�e$}i897S�����D���w��VM;Xۋ���"g�!��E���f^^OW�Ns8DQ��7}Eވ
�&Y��<)���%Y0V.���,IsK6ܗ4��[��c��f�g8|�F޲>�����|#�r��9g��J�֥��]�I�o�Q���"XF~��b'<DK���7Ǫ�J�`}g%Et�6#f�!��FI*R[AhZJ��@Z����� �j�w�8���0��B��<-k�yƻ�"`�ՅK�������k>��?��y�Z��r�}�K��H�'�4L劣h<�{S����,C:.��ۿ����}l���B���f�V!��>OCYp��M,�����	���
�Z��q�0>���e苼K�1l6��1��g���m2\σP��DxDL�/�tļ��aԶh��%�M��+V�>fx��\���G)�_ %؏��q�CC�s��ʹZlT#O6>t�b(Yս}�/CE���m55�x\��w����w8�C��*�[�o:�/7�,V0��c�g�f�a���H��/䦃����C��餪��W���o���\VC�GI��"�����`��`���Ё�������'w��bU�)��^U�'�7�@���%$�0^�2��{�]�k&m�%��p�	`%�����Z
+�M�H�� �"�1�`q��v��\�2p�c0�8�1����9H�\L��oSff���ľ��\
�����6 b!��7�����"_f�7\:�m|w:VR���0���#j_�8y��\��bXr�3��>��v���@�P3�^��Ӕ���sA���3��oͲ�4�Қgt!vn����^��$��_�A�Y�\RU�Qdx�Ek�4}����$DU��-U�$\ש#둋��ײ_,)?W��	#�7�خ��(�{b!'{��MR���[,8���l꫶0M�|.Z��8�{ƕR%��fKQ\��fmCe�}J6
wh?���ě���&K���<�Ev�G5`ߨ ��@{�M��b�@��s�-�v���>����Y~(�zs~���v��F��h�������Yo���~QOh\�?�eac��B]yxJ�W<�|�����.Xgz�5Hi~��}�*�P����&][����B��f(W��7��4���"� �E�QN��'R!=��F2!�ý2ˎE�N�x%�)��Bb��9Y�	a��[VIA��'S�=M��������@��S���/�xI/Y��J��Éw9ڑ���@U��Z�иha�ɐ!{.���4�5X�g�z���&����^����'Y]��!�~��./"����rw�P�D�����xW@ۇk5D�VX�߲u���Dc�(��������,�7s�W,ۮ��OӼFG�d��u���|}����YO�q�%q���GF�x��Y�#z,��&��k��vI&�-�{��w�}q)L�04X��G+́��F�/D�|��>9\`ʎη^�)�%\�>���#�蘤c�t	&.$M��Fe�Ҿ'T�Xf���L�\������"��cS(����Q�3I#F�4�N� ���^�7dGF�%"�N2q�Le�W���I�|���hP6��>�ٙ� ���B���� ��r��8�~��Ng����������JD����x����(�E�@?��Rǋ���m���x��gQj�1l.E�N�!�����Q�mKT�hr*�>�W�$ai��ZQ�*����:bB�u���������?�Ykf:ᮭ-Q����ߑ@�۱FTN\��%�++��d�oe��v�[A���`�����I�i7?co����ɛ48��*=�OZQ1 *��i�A�#�:�L��*#%x6v������Y�ν\�F-Nآ�bs6RC2,\��
S�")/��\��pF��4*�Z9k�$�񴱽�b����pa���+���*x�(2��e�O½j��k����Nw=��xo�k�1�RM6���^v��6���ύ~�{X�q1 |��ֺޤ�!��lʹ��	��ֿ�A��:��k�em��͙&ͧ��ld8E��*���&9
t(��8�6Ak��zc;,�f־B̯��ffz�?�w�]?k��Ĝݐ�`K�e!�� ���2�P��S�t�R������!��I��r��Ayx:�BZy2 �.o\"���)X��`�MA{��1�F�W@�HQ�F:������A��(A�Z���e�q^|Q��
�ɌT3������{�򓡲����@.�<y� >\�*^m�ًk!q�J7�3�5�䏓+5�{,vSmk�I��1ČC�S���f]؇ZH<
�O�[P��3|0����IK��M��DM3m�[k:%���U�s�]��@D+�����ު��2����zq9R��N�B�����qW�%⟻�N��K!j�bxN-��e`�i�;��?"�`c����\�;���ΑSiw���G��A���~K~J[d�e���j�m�5�;s���x��1���x{�̴�?VSq�@�)ۺ�H�I�Ӳ���M�x����z~�m��,��:���9���i����d���ї0ƅ�9ߒ�iV��Z��KÛ;NPҹun��ȁ��������
.|?�`bY~�Ǣ�q`�xЂ�ܾ9�����1gi���,a�߄�}��w����� �7��h�B��8���ѱ���B�m�T���d'}��p�D8�i�'(��b�0n����GsKRM���5X�/�v��:� 2sG^3RmN��:fb^S����J�ѯB�a��&9�eE"'mx�<���V�+|B��Շt�"�b�҄��������|�[���0���ҵމ��GZ�3-ߘM�[W��D9�e�V�[�_��wѠ���r��-10A7������f6�&}��@ߍ�o|Ѷ��24i%8m�]]�/���'���c/�h���V�N;(�>wl�B�#̾�6&��'C���`F��+!�X�xGj��H6;����\�Wx����/�o���?�2;��փ	��qͼDi�S�{xT�g�M	T�)��ݼ�
��N��_a���c6���R��[���1h2n��%-.��iSaᑬ�{󕞔.X!&"[Iϋ0dݷ��foĈ�"�5�p�̮g��v��}�A>�*O���	�=��]Z�)\�5zT�"8:�_߆�&�w���}�f�,Za=[Ы��ھ�G����J�����m�FR�K�{kf�%�a��	��?7Y�T���R'�{�g�L?z�n�+���t��y��	E�F�g��[�g}��S��G��_���H�|�{5���B6�
�)8o��BMX����3�x����os��6���u��i���j��xE�a}i�K�O�O ���� ~2I� i�G��	�Ρ�#V1DX�#�zy����7I�|��,��F]A��4�X����F(P�i?CV����q/��>3�C$����[��qJ��b4����j����>�<��s)��ś��ؔ�AoP`��⑑�v;4\A���κ�O�ǐ�#�`j��wKCu.��do���)�Ik2�u�r����>�/n����YA��ʪM��ߟ���)�&n���x�ĭ�(����ϑ�����$��~"Y��%�~�k =j?�{��q!�#ۏ���n��[���~�fD�RDw�)5o�8��%�;D9����fx�d���+O�\,�J� /9=	����g&�%�$�|�e���1�mZ��e p �R�6��Qr7Z�Ϸ ��JE������+�"Y�C3�}u}���'o�����m8,�=��F���3	t����k��Bv�g�̨���K�� X���H>�#�_���2�#�6�莃g2�.M��"���d|�g	#�5��~��ݎD����j(�<��W�9��O��ǔG2�e#
�J�[=E��<�R-N��,�쉿��r\R�ZpW��
1��b�.r�����"	v�RV��8��b
�����Z�?�0@0#�^�X��Rh�N���;ɾ�P�2}m�a�]��n����פ�r�G���J�7!Y���R<�����HWY����[�."��,����9�s�%E��pcgASjw��,�-%bo4>����>D���)бܿ��L\X�TX����b3�Q�R�#҄l���H�i��f���@XG�u�(c��� ����1yփB�������3J�����Qh�l^VR���oՂ%E��@�`]Ѽ�;�^�L�䢂������ɗ�&}�
͕�tj��ϻ%��������W[f?Yy8�&��`�{���7�]��x�,��\�����:��� 1��
�p��}[�ܳ�1\r}:���4)FQvt#�8x��5�����T^�k�r68H�o#�6��K�P��h����kU5����^c0Cx+iYg�\���ʞH�߯��B���YGDL-��c;mH���j��(Cƫ$��a�e$PQo��=�{�Z�f�9�Ubu[R��Ul�|�N��j�����ɀ�Y�}8���ͪ���r�ߍxxx���|�(��;��'VEHxt����4$'=���:�{2��/P-x�3̙ߐ��<=�����>�����~�$iy��ۿ�<=x_l��j^w>�$\L�S��$��18́��)1��>�*�^�r�/G�LD�IZ�F
G'D=N���7����y؊81g����8?^��<�sYR1�Չ���&�>(?PC�_,�Xd��Kun��p�O�u�������~�w�z��V���-c�A��O�s�r��1��dX\��,iGq��5]`�|�(���#M���ocm���4��gp�5�@o��/t�N��vF�q��7ɵUz褎#�%�c��Z��Ծ�9[k�'�b�w �
[�����Q�	4�od� g��
�%���o��� l��@�j�v`/d����
{�!�T���9���$j\HC��f:X���>P]��%�l9�o(Q?��w�}���O�PB~�Jp�X

	u�E �|�T��m"�x��w΢�LQ���1���v��_���)�J�9��J�ʊa=�Cw�q����1�{�E�{������\&� Gn��o��׹r�[�&q��@Qh�ͻ�	˥M����0Y�\D!l�ہ���PHI�  ��)�p�.nJ��K� *���D���|�j����qb�ԁ���齡Y��p��!t`�s�̱��b<�_einY�H�fg�� yh���#��'ߖ�V�٘Es��N���&׋&o,.�
�(�V��C�ܷ+��U��V�_�����14譕\:Lb��q��
�;��ۮ��(�I�4_�p�b�t;��(��"�+�#�g�UN��M�x�eA8Ruz�"_S�Q���v'�2�@Oշ嫎~׀�����L���6�|n q�N#A8[�#�	�!/_����	�K�
<�VQ`��w��p(�N?���X�"�o��	V���S�������6���{1���Af��/�$�G�Cm��l�RCm ��g�a�.�#�\��hO;?b�O
����ܮ�w����Z��*����E%����h� �Q�:U���M'}<�2��E��?�2{�}%~�)K���"V�`h8�@�3c>�쩁��)j.�ڙL�=���}E�3�rwVB�oi�v"�.����Sg��a�rK�c ���NԈ��-y�ɥ�D��bɕY81��Ϣ�H�;	{�2�Ƈ�e��<M��'�Xv�.[0����3�j��'4��"3[�pe��Ml�h���\-�>N7M`���?ъ��\�-�%t)B�R�E�6
��O\L�!s�aI�T�H˽Z'ā���U�V���Lk&����O�r}{W�ʸ�V2��>}Em��R�p�$:�E�v�yv��9��w���|�t���*�+p�����w�ҡoP��xC-���cZ���W��ׄJD�z�DġS�iaK����AD�&<��-il2ܜ����;�D���b���}�[ n՜���˗��%5Kd�g�c>�p��c�A��M�+��>�N_}eb.�F��(�_��H}���X}���m�x�ʸ>_�X�3�F�y��	~��F���q���B�s_�u*T��~b���@����91K�h=����g��P�nLϪ�Ȣ�
 �o� ������2�`dF��L��y��졫V�4�(���С왃yϖ29��Du���-(H�Y}q��A�����U�O#i�T)�r�ʚH�	���^c�o�Lu�o$T�&�[���7!]��
,ƕ�"���{oP�*�!���D�U?~67[��Y{f;�ET���w�Յ��3j{G���|H���)�im��<3x�b
������	���ʜ^�3G.��:7��K3��<5�nr���SLRӉ�(�XтZv n6ުN���9�%��)l`�RzU��Cq�p9�ի�U9qG�Uv7/��F������Y���<e�3�~��!��!����'�lK}`S9=_f�kFNq������#t�SC���:Ų֮� yq�ʝg�K�h��n;��׹�g�w!����!�%���1V�}n�Ѽ��G`{�����C��<,�k�!_������Hyw�غj�\+;a�]o��|{�|^����ui�����$��h�[�;�D�8f�>C��+^��������������R�Aآ�(���M��d��FzK��H��y6W��<�3����N#]�ib����*��|����L�����0'�� �Q�G��iR��\dG����m���%�I�{O������Vm~/�rL:��R 3��!�����-D�-�j�S���Q��H�������ߤ����<dڃ��ܠ(���`�b$%����#��S6^Wn�V *W�&K��V"z��QV@0F��>0C�]$x�T���(YC{��WezM⏺p�S��2��V�#>YF���-n���\�ts��tz�$F���F�Q�f��6?ٲ̀�a��P˚R���HDҞ�kіu�^��5� �D��<��t�������X	�R�ݫ�$�n�!�4u�t򖏆L��\�V�-��aS��F�8�B2��=�5�N���d�I
�}𕷵�׺(A��U��[C� ��I@��(���~q�Zhb�U�"�['����C��|,B�ش�u��je�Ғ���a d��~��>0{��a�Uo2Zm����B�i���Н�[�qz�B�ML�E�PW��W�e�7�ʜ\r3�� vX���{�(I���hF�X��0Ge���g;��}>�E�M�K�j� .��٪�+>��AV�r���G��=���X���1M/���`�ރ�SPH�6��8}�[k~_�˜]s\�&��V�އ��q��hiqlh�o�N�:������(g�.���}t�w�2�'d`=�j�3qf�f��T��]��a
�-�e��4d�DI&�5�ߏ��"Z�ƒ6���:fi������e۰N�[�d^����>�r+�� ah��,4�-me���$\��%,X����(����[����z`�?L��8j���/�N j/%*��{�hT�'dOJ(��9��B�9x0�0���04�T1��&[݇8hp$�8*���Ȥ����^��1��[��k�l��2� vFfPD�H��]2��bGA�t��G61(dY��ʎ<�ZD1��&���ǈ�Qd��[����1��PĎ�bQ�&�N��%�U�h��%��, TN���i!*�3��׬[��F7վ��� 4�]�s<�ާJ�<�*�'9���E��K����ou�����N��'S����_�Ĥ\��$��M��$K�2�@��[{����*1���c���j��T�c{+P�d��O[1�����!����տ"���:�E<L�6��9Xw!����{O�:�gӁ��AӚu��x|���=D^0����jm�3�b����%���]4�QiQ8��z��_Z��p����pk#_��K�����iC�ĵ�z/�~��l}N��3��M?���?�����Wx��y5��H�9�^��8�#�k�Y�]�"����|����g)ρ]|� ۭ��Þ,�S\���kZ�mD4H�W�.�q��d�q����4V��q�Z�ZI��&·�9��-v�~����eh���������]HyBaPǤ�@1ǧԨ�B��F�9�^9���@"�LG��l��W����6��Y�H��q�r@qDX.̔?��n��3'�)��5'=a���ի�0,B'�oK-
I;�O��ۗ�[��a�s�vP�a��v��Ά��/OI)���k��")����GR�<�bɵ���2�d�mv��R�2 ֯�O��bjv��?Wa�����~�$��7SZy��v�̺���\�k�Z�j�_w#b���m�ʘ�c�Fߏ�����GJB��b���?�%3�"�H�8�Q��ca�|ņ���´�����g|d�����I:�z���/��^�4L�N���׊M��E*� A�ė�E�y����ݴ�m�ج_�Н ]���9��䬛�'s+�ʢ.�C���^s�(���eU�u�����<[vj	��h�Z�"����H������U��БUɼ�gj)0���>[�y���Ǆ�`�L)B�g󂩗}|M���B��3p�B��|�`w诪�X��Hk��~nN�}c�YR������f�0CX�nn�e���XbP��6mw�3�Rr�sj'}���$%6&Sվ����|7N��E�q�b���1�[.��10BH��93��<��t���`y�2�F����;Ӭ��.7"�*���s؎��EДC�;�l���x���X��q��T6�x�`c�f��L�	Pgn3�Q��Zbf�eRT��	��r�,(���8ěpe�0K��ot$���J�e
S���N6��I�{��R?<H���0b[�5��1��&l�T\2��������^"�O�w9�ep�2�QY��(�z��}�?3Q��f)��te��� Q2�=HQ���'mU�x��|��;DR5d��7�2���u��l#��pL"��ǜ���-RAi�>eNZ7���T���P�����
�s=A��[n���Qq�o��r��_�|ot��Ծ?��jj�c��<t�5< ��b�z�˥s��[����g�_@;��"E��C�XzQ��Uq�)�*3��&�9[�@y�I�򦪘'�=���<-�4�P:
�i!��`�t��9j��呩��;��M��U5�_�e����FfQ!��􉵓)�܅/�D���B�F+Xy�H��;����[�A�� ��pE�z��2��7�*$��]�V2�;E2@n�}���!�i���Q�06Pކ�4
Y��a}�V�jGO	�'�Y캥�x�������2u!�8L�^���T`O�$JMC8@\Sޱ�+aX7�;�
X�E�'d��V(~`<hN`�ZU�R��V4�	P0��p�]�Ja��x��Bn
��TC�*>��S֩xc���w���W������K��5=�eė����C���8M�4��8�/6d�ϥVe�.�E�	r�j#��p�/~�X��	�eهՆ����)���ѴN�~v��Zm�\��~��L/���r73�;$97�%��5���28�*r�(iz����w���dy:���R�*�Q�@��e��p��G���6R�z��t��`3��/���(ϴ��'-�փve��8I��� �5��n�r_�d������M����?[�#�Qx%W{��]Ϳy�ݽ�y�T|�ԋ�_}s�b�����	����7�X��� �n}��k����d7hꓕ3�h���2�3�i� ���18�۸���t��^���� ���f�Wi�hC��}zz��:�{a���K�i�XwT��'MJ����`x?��R0�0߸
#� hW7�Aj[f�<���C�x	�e'b6
d��q�l uN���*�i0#��J�Cx9N�����<���"�?�!���A/��Kߌ+W�@{�j���	&3�ӆ�D��V�p	P��b����]�,x����Q���#�6�]�|�+�c�J�Ȃ֑��tp&9����vf��\G,0羸LSc�����������r��"�$�*o�(̺%�e�LI���υg����HԘ0J^��f��Fw��>�a鯃[9Y��k�|m`S#<X7��\�?\Üt�x���{�*��Ԁ*d��K~���rE��ba�ڙ*j��7�U*��D��C0�Om&vk֐�+�)M.�̏;�& �w��E��I��<@Tf&��44����u�-�8�2�C�n�Z|8�+~���>�a��׍ͳ�U7�G'�.��j
P<C����50�@Rr�'>��W�oK��ZQ�Eh'>�@�� �q����sR�o?�d�g�Il�*�#s���u�!������)��O#N�2���3�R!�涞(��X_n<i<r�]�a'W`?*�2�O�օ[w�{����j���Xa`e��(�i��*�
�㳌Vp!�GQ�����u�m��D��ʞ7곧Zt4�m�����#T]m�k�.�u쎽-��K,���ְ�h�|Í��s�!�0���f&�`�ٔ�C
Q�EUZ���\J�=RH���,Hs�,N��ׇ?�Z������[���9�Q=��f��������99��u�	�x�֊]+���Qѧk�����Y�.�n�%\�JST��sQ@lk�>c����PZh���Q%���`%�}�I�ܒD9 RE��%S��ht��I���s�_��T��Wԝ�on�_n���?�n�<RZAb�G3�O3��+����b���۴k�ɩ8�du�6�ac���C��w�̐��,̔V|�,�(�� ����V�1�I�U_ц�3�x��xT� hUЬq�(0�r�ɜ���ȉ��v��fZ�^-���Y=N��(C�W2鹠9����>�S���h�=	ۺ�Y�R��LG�q�i[O�VټA����V�)�Ӱ��eLiF��(C�r��'j���zU���á��7��sH���rϨ=PؕY[�pV�ԵO՗��e��,7z��� ��<�i[z���UX��z
�	�X�$0���1$�kü��=ϑN@��aW� �*/Ji�b\*�g��]�����ãr�K���|"��E������o��������0 )���k���5�a�dS�������<�n�`߇4!o+���4�w�ԏ�F=��������鱛��?H|���^��:��kӃ
#�*t�3FLW:�ёE�� w\��zlg�&�_�l EYz�x��R��$�]BnO���p�&�h��9�`�U��9L��E��bo�ҽ�+�6�=�?*�%�I��[�[�L	��G�.�5˭��i�"����	y�?���w��|�
LF������U���ڤ�q|��'��Dܬ��R0�����z��CD�@�*.��W����`�Qd8�k׷�n�LW֦�i��Gz��� ��}I�)�)7���ƹP�?�����Ы$% �r�$��)sЌeV o��N�Z)�
��Xˀ��[a�@�a��^%Ŝ|��+���J`7�4E����mFn�%ںy�.�|�.�`�S������)�@��Q
�II#�[�|���M����5�� /lDmt���02j�6������G)� W%��:km6���O��uH� �ld�h�G�>�
]갸�S�X��hʛ��W���}�����4;1:A)n�$~�)�+-�n`Gp��V�-�~�i�o,��о�Jm���,ውJ3&�����c)���(�Ժ��B��/~�bx�K,��:Jhv�6�6�v.����+'S�y�_2ofzaFCf�7���Øt�9�L��Q0�
�.`|�Vr�jz
(�?�	��a��\b�#��:�7��~Su��[��1*��dt������=#ou�V��r�X�)X��[���.��n۔�H�vI��F����9��n�'�C�1_b�ȴU�7h>�-���xP����q_�e4V�	n�G��Xq�w�3P��wA�!�u���{��J4����y����w�e+��$UHv�$Z�J���2`x�e+�L��_��v�ޮ���ܟ�ގ�9�"��H�N�ڍ���X���A9��y��@]o�ɜ���G�b�f��8B)��(Ti�Ņ�.l��xac�1#X܋�ҍ�	�ڣY�Mqz�aK�������+>� ,"��a�K���A�ғ�^j�ࢧr���^��G�ic�鬼�ќ��1$�G>b��G��k�{��{��XC�y�)"m�6�F̧!	�˺�]���n�.RC�'����V*-5�b~��%���[^����$��|�t���4�J`Om������iP����|&�%�#'�� 9u��*y
�?%��{g�,�����:�e��h��}�M��┴W��Z����Nv�=�M�Y��JM^ ���h�҆�밶���RIn3*(�W��A�D��VY�3la���j[�t%#��	��X0���7t辨�2��zi��P��(Q"�镶b͡�H��?��)�p�B�3f��H5�xL��x8�YY�nK��K{��P\��T	��D.ic���x�����;�5�#���E\���m�y��=ES�SϠ���aK��/�Ҟ������R�5ԩ�g��ǁXܷ��6�.ߏ6�s3�)�zHЯ��X�'
��M��	�-��[�-g=���V:,ZDt���Om��ۧ}:���@v#_�CSLi�3�[�ɪp�����;�~lT.Mt�K�|��C�K5��p��DłW��9�d���r�a���Y���FouE�6���Q������l�Y󄈐Y��*vm+_ 6C���|c�[-�߹|�����T�y/�*s4>~��$_9�|���ܥ�{T�E�O,�RR�5�N\*F�a�ڎ�����o���4ދ���o�1����Y}|{�� ��eݢ��E^�(�=�qZ��mֵ��4��{��18j�I���AvfQ��K�t�*��nQNS��D]:�s�|2�r��1F�Q�����q�J�J�pz�>q�{(��e�c荍�0)��-t��_�Ď��ݫ)�����SYoa�\M�֭��
��2���)۳
)[������ �d4�Got����ګ�H�6�;��Q�|-��\�~ =�(8c!-?v'GA��F����(��(�H:h�,6K���M9��-���.�:>��3�,�-l���mAG.�Mҥ��6?oK��>o����KUV����Z��D	�2�+G��ѳr��/�[����ި�?�����`�s�SY��tYw�MX/��5P�F��PKC+ZL�'��r�F����u��_G��k�_�\��ȓ��m�X�G۹�غ�����V�R�]@<�{?�8�fYO���\L���k|�T��V��s�1?��F+��r���풆|�k�:zj8��N����W�d8u�1C�:eZ)����a�osf�'X+�{Zl��q��#��~h��� �_:�X���2&��ŤǮoVp�r�]�[O�l*�(8Q�	i��)ڙm+�D�eÜ� �mV�j;�i =�F�L1�ޫ5�I�c�{�ī�u��#.���?�3�O3v]/vٱ�fnw(�<��t��,�l�����u���	4Sw��ա[����K!n���ƺt�5@,���J�Eۧ}ѵd�u|���T�-)`P	9H��̲,���O���^.2�����h�8���`��6ˤ�!n�h�Ŕ\KQ��8��{�%-ݞ�y�lw���[��ѾZ���|��J/N�;a�cP�`������M�XP"�5J��ǫ|v+��V�RxRM��r�A���WHܳTcx����ҟ�X����v��=k�=�� �\�T��͙���+=����0+?䂭C��2m	�;܃k,��d��������w����4Z�i8�V%X{����[���)���D�%L�w�d�W6��)^��B۰�i�l�+:�Nn�Pq\�xC�AS��M���v����j�7 E܊�sm/��o֘���{�΁�( +xn7۱�_fuUNM��$|��)����m�
FK��o~h]t��Wb�!���S�-�zG��;f�tG�I�6߁�I�?ڬ�%@���l���������u��Z�`�������S���h�!����Jb��/FW���
uRe��:|�\:��+�>W�<Y��gX\�Y5@{��Z��K�6���B�2����%J��+�Y��IM}%�]�e�H��B�����Z%���C�{	�6����$x>j$3CǂR�|__$�鸞��a�@.I��eg�*V��)�.r_�VI�e��u�m��D����UIXD�Z�]�tMӠ}��g��h�kM�3��5��8�m���I^�6�V̓leL^��̵�������9����38�vU@���o�7ۇ����h�窙�H�E��"�����0bQ�Fb�V��1>�{4$ƈi�.�F�v�-wTV�!F�e�ޤC'�\`���R��q�#�m{?	��н>�L��L��q����x�p'����i� �'�U���������ZJ�Q�G���Ct�/:����8{��6��ۄ@���*[\F:{υ�Uqʇi�9=�5��w6���UM��g�N��v�T��4���Ȭ�6�e-�Z!-靳��!;���`�e(�t���_|��g�'&�Ч�I-�M�J�R��V��-PĿ�`�;��ö�R2�X1�꒻�!k�Uzˑ1�����T�J��. �ո�ܺf��m�?]A���Y@��k(���Rj��t� �.���}�H�t�
ʬ$��+ᘊ�`���k����L~5�-W�_�zWW��D�������!�Ԝ��0;�i�m�f�`;�*��P���P�?�$=�CC�)+�|���s�8D��z@l�cv|l|�����(I�X1Bhh����4�=�^Pqȑ����&}��|�i�>�~^�l������N�1X�o�,���h�(ܟ��[�E�bq�	0v�։��"�+�����f�"�wsܐ^δ��/
��?t�����3�F ��ߚd��Z��	�/k��B6O�� O_4̦�i$�j;Bv������T3����96[��Ԥ^��K�r�����Lb,}l{T?�{��o%#�:��H�Imߨ�ٍ�Ԡ�t��^�oZ��A�y�}U:qC��N�֔���P%��vOknQo��q�A`vEr@U�8��=#�,��Ӓm�G�fݤ�rc��A����-�����v�q�'����t�����yS6�����9�d����""��t��Y0�� �t�&�l�6]/\�"��!�\��lə�@�����0���c	A�س�J���I�t������7�"#Q:(�� (��u�|o�ka�����h��i��$���A�Hez��0�1�;�,�٨�$#��x#�sg������Bԧ �3��2| ���ܔ9{�7X�� �����%8e�)ћ���j�ͣ��;[�}�$�ŪG��B�\;�aȘN��oH4�j�咙D�Yu��7|:��Ƶ��XY�
��.9�{�y�L��J�G4t���<�*/dY�\��O\4��=��L���̞kc;{P�g=<����92��U��]��je �g�<�Cizm��Js���ͥ�C,��k���)��Կd���=�}`�Da�G�(��Q�!�ڽ܇�Bۣ1��5kի-�F<"��y�?_o��#� �[��ӗ����k��?I����s�Y�h%��(5�<�E���g��͕��-D������}��l�ׁDR՛���c�n{J��Q�/4�w��~�bP���Q�E�0bwI�+��
�.�I8g��/JmO�W�@���P3�k���x���_҆�v��|��>���L��w������쩱��Јi�m��/��m'�;ųjA�9̔V,ǡ��$�D���0A.lU_�l`�D�Vb�6��Vnk����[���2����3Q�L-���s-w-�G~�
���"�3�j���{N�� ���Avc)����`��8�
��m<��,yb)�9L��o�- \>�y9��	�XZ��fG!������4,0��~"� ��9�\2���Ө"������c  �\��7��?���G$ybDS���W���	_�<}��q�P�
���^E����>�/��@wgT0?3��v�-1*�5�H�-�68���e"E��`��M��6g:�'T���Iv7.��1�����_!�D�V,�>�C|Ҹ��uW������d�e%�K����^��%S���i��!�� b��!���/�8K�\���W>X��6H"���Mbx-��_�Ƴh����r#"��L癘{|���]9��-a]���EF)��|�!��u"�݈1Ȼ��F�!tۅ?�S��Uj |�2�� ީE�h�X,�+HO�nR8o��:�6>�9�Ѫ�+j���l���WA 97[��:�먪�*����Mb
ٞ��YB��|���X�%���k[�q��G����m���	�2�ڏ�b�X+gb	Q���b�6*Os����Q�H0mO��,�H���Q(���K�>�^�jΪ�Tx$���x���[��̾cPa�����1`��L],
)��w��N���^���B9A"��a�"�^���&\u�pց�⎳���-{)������ ����V5f�LV�˶>a�Q� t�ɣ,��/y�Fo]�
n�:v�-1�%�klNz��a�7Y<ݞ�S,{��Be�[�j��x`�_�'
u R[E��M��bK@J\�Z�-[�N�j�E����c��gJ`g���Ī��ρ��_�bs�-���\�T �EDs�HmV�kkf`�>��OA|}w�6����v��w&��vy�o�l���P}�g�D9�����Ej��5�$
:���od�g�
�+a�յgs"�8�j&\p�0�M]p����6H���&�&:_��+}+ܜ࿂P9Y��t6�TU5��k)��A=��X%2ȕ s�C������\�4+�'ja��"r�ASH�6E�S��+�}�=��Z���y�)kCC����ԓ�Ϝ�8��$�ܗ�n�S#���$���~��F��������N�9�S�p��"]u�h����y�3���6��%118��U=a��\D�*��CD�$jO�yދDgKV���Pq���Ez\�w�4N�#?1�+:�С�ޥ�U���ڝY����U�����	ф��'��wU���t���'��'�}��V9����E��/K�r��Z��&c.�� `|-S�FNT}�g�̄��Th8w	<�Ei�,�Uz@]�Ik��u�Gxl��~L�Ք*>�@���t�����v���Y��¬M��L�WW�Ci�F��]E ��1]�zaϊ`�m���<lϩX�<�>�Vg�T������G�����˙3���/�v�n�rW+�{�X?����(�p]�i���d	[�a�8����^�A�o<��oI�C�}UA�N�m��2͕�~�P�U�Hc�D�v��uε��&�{�k@`3g�G*d�=����"�-O%Y�~��PpT�)��+�����%��aP�N�)�BpL� ���[tD���4��c�����:�@;E��+���ի*mh=���;�!3+��{��t��w�zza�ͳ�*�G�����۫����|r�fǦ���G=��S�by�ʁ�.��JNf���oR_�����E+HQ�J�Ń�h�p�	D��b�����<KV�T���;@)�>�{��5�=��Iŉ��i�i~b���h+��c����"Duz��GmȒ�+�-�%�P�ū�R�;�՜�;��*��Ms-_���h`�iܶL�� ��(��U�z�EI�xsB�b/|�Y� �p�xmEA��Nv�0ޡ\_t�:'Wjk��a�MN�!��Pm�%0w�2O�tJĵU� ڎ~�Pb���Õ�)��[t��,/�XѸ����%X�.w��/��k�ڐ1��$q���|��	��Xb�~�Y�$���hΊ��Yq�K��l�m���X�p�vw�3�|�tLI���,kd�9��G�t(f?L�U�n�B8�?��X>F�ڡ��,W��8�.݅��ǿ��6��t�؇"Wmv��(ߐ9�0�ȍL�Go.[v���<L-;5w�t�����-��ˀ"�����?���?F!X�Yjo � b�(�&Y)'��1��f�k��!�1�q�H�D���?�Ɔl�h��׎����r��~��y�� dO�ZHӞ��jG���1
�v��Z�f���Q+|ݧu��,��`�ۓ_��f��7�P9>H�.��a���o����Ǒ@���S��=�r��,�Y�����S�U�t�Wu�
<IݨN=4ŀ=/����KH#K�jr:� ��j�.�t��g�Z�t_���S��}��~��E�S��1}�*�����	��)�����@h�`vM�Ju�<\�wņ��ϗ+�o����K�Ob�T	Xҟ�b���6��/D@w�Ip���c� uZ�ь���9D�8��cL�Hj6�6*Q]2y,$��
pC��t`�o��؀�H睳{�o�DP����X�q���SQ���@���xK�%)��\��9[ R�Dye�i��Jzm��菈ep�$Q��λ�ؘ\|���?��e�X�,[�x���6ed�⥛W�����]zd���W]�����	��۩n�rQ]`i��
�*@q��b�m��)���袯�}���:�Z�AP�OPF�6]����� V�${� ���=o��L���Y�^�Gv�����N=����:��>��Vݵ�����EgTa	�3��p;��K�?��j���`��H��|�˙��04ttp�`���\!8ԁ��HP<>�FF��VхO�x L��M�Ö.C_�D�4���y'���;��桻���<��2��8)"����X�֦/���^�V�G��^i\p5����7��R塪;w���{2K�B�2�6k5��96Y��_0m��F�l�����2	�2	��^Ф�r�)�1Օ�Y/6��T��ކۋ?�p��[/áI��^@ꛗ�����"u����9.��o_�K.?�P�S;�8A{@��#%�ї��A���
;��Ed�8<��2K�k���/y�q6����b����`=�D�M�Wue�,��$ܾ��+��k�5�ٞ�M0c���,�H�F� B[/�ݼNqj-FWq��-̏�����yPю�7{�rY.	na��-Fܻ�ikT��<qOH,''�6�-��v�ki�~%0q-�����_��3�k�� �O%s�z�:�Ug�91��>b�zZ��|? ��h�G�>�_(�AX�J��WZ4Y(�^�757��gT�i�lI�(��_>�b#���[�F�ь�T�$��nV���������0E�O�L.�1�~:��-aG�e_�l�W��=Mr:�����l`q�N}�����~֒�/�t�B�{�&��_����Բ���9P��=����S�ň�}q�\�;����sAAu�Qa��[�R`,JF}q)&n���WxPu-v�B���֖����}d�O����'��%ʱ�P���\[H
n�����{vn�'��� �����0m��?�	N���T�Y

��ߏ��J����wCU5�\{�ĠW|@宎�)R�H��Ff�m�x��'�4��a�f�D������8R�=N��t8	�m�⿻y���|��bZ���{J6#Q����)���ƾ�����=��de�G�������K^}��\�X󘜀����^��y�5f-ڎ(��=,�Z�dƥ��Ps�/Ω7��=�����45���GE�{�A�w}=�l���	�K�ńT7��]_'���W�f�F^J�S�KA&�~�R��ٖ���+��섅L����IfKGAQz����i׮I�DqԬ���U��q�Y!%N9V����<�P����-B��H�?M4l˃\	�ADF��|��ZsGL�g����&�6�d@#0�DػYz���y��i:��5|ʶ�eՂ2E��ֆ �+�!��T���	�<�g�kRT�B�#� LSu�[�����en�5Q�o���cN�(��XߌO#`>>���Cu��)�fXs��h�"w�|��<Nr=�<�)0�a<�uNS�q�o���'�=�j��2�IQ}�� jT	4��s��N�����>r[Ø)���쮙�r�#��[_wk��G^�LX'�P��#]���H�%M�=W�����n�5�����b�|\8�	-)����
�}�(y_r���?_�M��Ydl�~^��I�/��b���'�+���+y�Û�� �Ћ$U1}�գ�����L��V���Ľ��ϋ!/4�|���q��0`/��!lg;⍒���? �-q)���X-a|ԟ.2j'tф��e����Q��I��q|��u�L����ĔlyJNR}�P�%GZ�^]rb�"�����������z큍8"[i5��F��tIJ��)&t�D��<"�q�5�Z\4���e�ݦ��@ڡ�C�\E"�l�qNU�B�K���y7u)2�8���\&Z�G���Y)�k�󧏁�U�=彽���Y=�˧fb/��i����~\�kh@ge�]K�������+я@/�J[�|J{�oTM�>hr�k�k`�be1��Ě#O7�DGE/a��&bҵ��G�4�s�#�>�i[Ӏ�o���c����v%��3Nu8�·e_�k����l�&N�F���XB�q�ZE/��q��X&N� �W9�֎;��%�$��N��pz�7�M�xn����U�۟�G��̛�XyL2}��z���15ڜ��(0�؆=h/��ɝ׵5	?Ь�&є�ن)K�[P\�/��J�=��t�+~9�4�#�ż�^էXj_T�h�����k�8��t�2d¿f��n��L�8��v	b�]r����/Mpa�F.F���,��
��Ơu�í����B�F>%�[�F0�[���23��ƴ�#~�t�1\&~8�Dt�vI$;,�mr�y��x���aԚ	�/�2S���=U_H�2��B���N���x������cqsپ��V?&P��U�'d�ˌ,L���eV���"�E��zfJI�S�	���|�=�/"��a{��V�U��ɵ����39�G�*�JN�LV��������?�SOEkP�VT���j�uCѓk�5"�������a.����J�|k�7^;�X��$�m��H�ݒ���p}
Mr����o+�2���N*��ñU�����8vF
m�Z�(����y=yBһ�V�4a��y)b���I�9.����T'0�c�>�!n\�R+��b��2
�@�>@̛�N�A:gr���<�x�ԙ*S\����F�#��x�K).mYB�?.i�Yet�?ه~Lì>o�s��Fn�H�=�3`�\lS�T�n���O�B ���9�aI�	p&��D&����'���VD����L�H�A��+��&�/L��I�k̀�T�iI1�s¡��6�dYW���z�G3��Z�B{1���n�2�?Y|ĸ�{"�DFФ��w��R6�"ҝ����Z�f|������ӭ��
�r͉��ʡ+5@ZT������>�rq��`X��M��XF=j��(l��K�u��ևM���9F$H�ά�ZL+3�:灃������;�mJϦ< ���DB��_����=�Z����A_�0dC�e��#�ml�
"`X�\�h�"�Y�'x�gu������x���IN �j>S
wt4C�V��+���5x�6��pG��>�4�������:]���`7'��vB
H�	�k���GCZ��Q�
��A�?�U���p�$��+�B|q'#I�urR�"�H���u}���=4���u�M�7�t�f�ͯ;'iА���e��ҫS�Ϯzj ZE1dH�ߴ�R=�+�7�B�0�(���(m����OaLq<�o8�a�;:�HV�7�nG�kXH������7��M׃����s��4��ꎹ_��ҙ#�H�ո1����<�����dAi?�Nj���GNw�u�&Ph�_��'�%���rP��q�q�0�K��i(�\Y��
0�D���Ĥ�4%���y����1J���Xq7���
��Cg>�H:�3a]b"�N <[Ul��~��&b�~��!}�6���V+��^/#C�|FO�v��sH�yr)H���P�:4�|��%�cI�=����wn#^_��&nt��O�cs��\���ο�e=�\iB�08��8��t����at�\y�9��QH"�Qz"rw/Ƕ�-���y��7cg���S��ʯp̢t��5�9���n*!�X_#G-�g�:�[��?w��@.��ҿ
�|P*�}Y��`�(�{){8jg��v�i���E�p���=�'�Nf0���o	KQ�!q�����O�3���gŻh	����<��>�X�ݢٲh���G�Ա���9o�ۥ���/�L�ߖ��7h�&r�q3LͣAcʧ��U���r
�I/0i�R;��@LMX����S���+��n� �j���T�+�W,��"�|����u4G9It���ɘqBX�\7 ��% ,2�S5�"���i��		�Ҽ���z�$�W��c��q��8A,Қ�:�����u�Pz-�}������2��ҽ�\��R��"������	Œ2d�FgѾc���J:�zv�m� W$Tٗ�l���'�T}��a��ωr �pH���� �{�Kn(��<A�H�]��/hBc,����{���`����4>3����v�U-�"L},���]��W"`��t�,)��I���[N�k�S�w�]��ͻ���l+d$��M�-��T���ɦRܹ����v�g�w�[��)��*�J��l���&Ї���+�H�8�^������0�eX�R�cMC$�W~,p�O������AE���dz�`T�ey��x3����;
�N�洘bg;5!�Iۿ!սQ�D��>�˽]�Cy�D��.���ἣ2��/��v�l7��D�c���A��6.�q������F��t���z�-���F�~c69����m ���
7�	.�-xBJ��r>�Ժ.nZ�1�[M���áM�/`Ɛ�g��~�k9p�ćt�瓜+3)YP�|�2��?`\�ǃ���M��νo���UIG�z�!��� �@I�`}ǳ6�^$�ޛ��p>�1b6G�!��AŔ�W�Z��21=�����c����d�C�Z���bbx8�M°�ST��t�ǥ�gs�����[�NcA_��!"17���-?^3 .��c�Aa��QUP+�ru�����Y]�+J�����h�!3a`��Gn1T{]E��D{�ԍ�4��.F7^6��[u���`R��9zk�3�?�1�0c��(��QDrB-��A���+� i�C�<hBo�#f ��b9�U_@I�7�v3�LI��]dj&�J�akY�+����&�]��������.d��	����l�S�invcINx�:|4*]��gSl
#G�p�}��]�cS�-�@:����="�j{�?�e�9-�`vK]������hS�D��)�I��Y���钀�P��%�5�-^G��{����f��������!V��=0����L��?�r�d�����%{?K����Fܬ>��s�����sP4]�`�;�x���#��V�4���o?��������u�F��!�_��q��%�eOņ�j�ʥ"@��i;K�@JJ'���8W�K\�Sc�2ٷ�y��US�7����C�h&�~˞�˗J�2�-���X�V�,S��IpI2HG� !�i��"L��l��<���{��q���V���_�0�@�TZv�������V�L��l*דKV�_8Hh����?���N;�S�E�**Ȑ:�4R3pg-<�!��Ę�e�i}d"�6I*�}3�:ƪ�n�K�D���:�)�l]��cA�����TФZ��g٬�`k�q΢�-5���}z���d;���Q�.���6�1��S9�X[���0%}��1��0�+_�#�����3ц{�K��>�����U^��QO91��=����i��" �f5��׎f4`cTqm'��$b�"Ճ����lQ&`���>^EykC�sn+I].f�j��"�zM�#�J�֊���T�\���dܘ�ç������zg㹲�L13}��n���ٹA��n��3�a]�����b��Qs�0׏�g(�S�`��I��hɊ��Gڱ������X�~"�DT r�(+��P��h�De��c�mU�+�7� G0ˤ����2���:8N�p��]bK=��v�n)�>��wEm�>�8�#��WtQ��V[F�-�yhB�p	���Q�Th纍�9Q[G���c|��~�3�WL%�/�$m��L�?�BT��`4�-
S�yaňVt.�𰜻Pg�7=]�8�'�f�R[Ag���%���qۑ^aGF��h��a�x���[1��!��9�`|8�O��\j0���DB�있�.�QG�S����av��&D5iV��F?l��WP?���h�x��P'O�\{߂���+�c|i���6��L;3T���2i�O�j�6
y�vNM�� �����=ַr�-�ch��f����X����4Ǡh���܅�DA)#��5NhI�����-z�Q/�{�!��&\ڨ"�c�ZA�Q'�w����;��F����Т	G�D�=��q��)t��g%���}�!R���W�dQ� Lw>�-��W^$�)^��5	�����gD@�s��?��N�u���N=�[Zg ���8��s#�3EϤ�J[<��-�8�������G���A��o?0�Oq��
��a�|E���wqr�(�+� �fJ���E�v�Bآ�4�:P�5B%{]�ԟ7t��
	N� PC#�L'�%n�X�S�ڵ���M%����NsG�J�7@s�u�o�6�̞�9lW�~������A�:�%f�깯��6dF�D�*�N�-M��6����8X�GQ��	|4�	���J�nBL��l��}�3����\��d�V������)u�j̐X���S�r9��3�����a$M�c�YN�
.���YR��U�����"�7�a��E2I��V��	�l>D�[!����&8���Tt(|B��W�A��w-F�G�H2x�uKG�=�r����JHq^�?�n�%���mEk���'j~6K��a�P�c&�����t��'-�a5 �ӿ>=x����-BF���Y�hR�v��2
����mad^>0`�/4I�I�%uj�A*�T�4����FoԩJ�����=�U��J�\�xDW�8�����9���X尃��4��`�-�v���&Ժ�2 |[�s�{$:M%x�{�FP�\T�9��	D���F|%޹�5\8c��W��ILwP3��K:ٰ��t��i��	ne�f��&(
n������9�"�:9�Q�[�PLM�4��D��vi���b��G��L�����#�י� $^V�a�^�MD�'�6����v����f���eg?]�5�B�D1��Fvr���f>�t��XS����c�b����@9��!C�դ�d�ҋT�if��q�jγ���z1�X'�����-�d�����m�'9^,c�%����/�ϣrǛgoY��wg�nRj_e��^��@})%z����M��0S��"4��c�CSL��0$YV}J	� �}�J�n�sp.s�h?wu͞���ؽ��S�r*�Ӥ������Ři?g�4�^HWNP;�2�)����n���I�*&��΅ѩdowI`�{�u�2q?(a����6��Zy5u�a߆��R}-_�2����������� :�9m�<1��'�j��"d��y���W�������zdF��Q�N���]u�9q�8�!lc]U�V$�M������!�li����Ad��ݤ�✰�K2������b-�	���L�rt���Gc-�/�f"J,�,�fG�4�� 4���&���
j�GS^�#Rp�x����¥�|�WG�+ƕF��Ve�v=�^�6\׬ce7b�F��[3Q��KV�j��M)�������dJ���.x�^8�ސ#�5'&.�H��>�0.����`QVi��łc��M�x+�+��%�i���w�Z}���3��S�[Y��A��gk{HmԂ��sLi����׭��%*Q�4�T�gȞ����3h��L�^�o�q�!Ly�$�D�"�?\4z'6Yv�(��$ �>U��Uߥ�o�N��(�N�I6<P�K�f���Z����-���pz��)���6 ��w�k2kM�ሀc](I�� 
{֍^|p��s����`�H(X�莅񃄋n,��������U`����	�,v��;�gM�m�z�n�1MJ��<�&�B��PmdU?����3~\��ڍO��	*��|�^Q�����ln�盵�?��t�!P���#\�kx�Q�e/��+i���.y�$���A����I����q��E�H�8�AKL%�cx�?Ț(yY��YO�B9� ��7�1!���+������*D��t8o��~��/��j�Ȓ_b�'�l����&��<� :���^$��m%��
�w��Æ�F~tu���ϥb*��F#ur�I�~M��=�~�~�l:2S����[������^�9��?<h{��j�-c�U���>bCcb2�֫BDH�$�˹���� ������wߨ $g�f���F�E����9I��ܐ��Wo�(�#.2v��;��[��[֚�`���=m��0h��Y!����]��N��b�c�oşݯT4 �k�,-3^��TG�I����"Xz���{лX�J�����
+���C���f������4*�L,"�XC������O��{Y�|׫��w勺�Lm��z@T�(3�<��)�V	���2s7���	�KkGL������1��O��_�s�w��&�"M.���(`�a������#���b�;�(eB�	#.�XX_���F=��de�>(K���[�prj45��Ը��ƈ�VAKx��ΈŦ�&�s�~`%Ua#1tAB�E�FF�C
�,����bK� 1/�ݎ>0�e�$�����=��o��ş?9��u\�2���x �s��X����F�]��Z�/Dť�J�\U �6�`���G_NU}
��^�/��W9�����D
[�����%��%k�QV�����	�'���m�����C�UW	��v*�Vf��߸PS���'س�(u�O�>�s�FKO~�S;�X.�%J��7�tԜ��u�8��û��
�����v��ܟV��x�#k'�h��c�fU<F� �*�uJ�e�`CrR1F�}#/��E�3Lpk{��h=!��E�O�2ϻ-VF����0b��Ov�~;+s�����/A���2�4�!2��=|ӏ����I� ������HS �W�-HO|�ҝ�m�(����'24�u�ѵG�ǔ�?��;��U6F�!�	�v��t28��7D�&�h�J�TOP/,\�B��7#v#����+#���ܦ��΁�ԟd3j��ioӂ� �!��	#�4�=���5�M ���&U<j��e��Ԕ� )�-�9�j\�CM��ǏX:A���Y��y}#آ�Cf0;~$_��֌�c�/�������>��߿��X�<�-� �<���pKA�2�(�>����c�=��cߏ�6~�'��k�\VB?��^�X�6y}|��d��򅋤 �K����R�G%p�_�>|�E��6�!� 3iEvjʟn�;fbPqM4-����>�D35����D�5�+�{7à ���y��Yl�,�J-��HA[�=��1+-@�Eޙ��N�8��k���q�9�Bxk5� qX^�W�����*k��X�$4�:�Ϝx�S�1O�A�n�z�p0�d��|�B�5���gza_�9�, �v��B�T�Ȕ	�M����Մ3���;� ��m����MrH�������Sr����%�Ao�}�+Eҳ�/r���B��6��ew������1
i�D	�H��*��`����[h⽖�,�;ƭsG�y� ͟w��������[P�*�2�̈́��ֵ���5j{ԞF��`?�(�'G�,P���N�k)�R���^��$�����/=���R���:�G���!��>R1��cjm��'�l�$�6$^�g삋�O�w���ji'�)B��j#n,�e�
�]�襤��m��(�~?hv�����%LC�&|�q����s68Q���JX�`��L��2����B3�F��	n�?)��0I��CG;�]9ཏ� M�����÷w�K��0pN���^���'���E*H� ���ߙ��|ׄԼ�kZ���Հ���G�3	����AsQ�SiY�)��(4U�4�o����, ��m�:�Up���-���#'�M�j%�5|HGA�݊*6p��? ���ں�m:���!���h�eζ��Oכ�vx޽լ��0_����{c��l�Z�y��q։v���I?2ǽB�wfMܵE#_�OB���H�h�s�ګd㽆�Y���y���I����:9������*��@�Ҝ<
2)3ھ�P�[%�I(�_dΘ��b�]*`��3��!y`v��e��N�<q���7�%������p�������>���y;{�'xT��P�V�
=,�	~�2agg�t�z�P���%\U�]��>��Q��lf�G��5b�3���W�-h*���Ը+aH�B�;{���Q�>�T�.[ձ��M����E�p�uEl2����ݓ��V�*#+EC!C�S���.��v����W����X�o�J�4��QZW������^�߻0�Q�8wI��-X��&@@t��Yj��7�"���q�������+f��F��<��٦P�,�q�CΩ��.��V�Bnw���A�!��R6�PN� �U����0)ws�|���I��Q�P���^�^��`~Ǎ��ml��/�W�v[�y����FM�n�G����Xg��*���2�gO|�s/k�J�/US����q�ha"����`~��̆�G�۹p����F����4]bJ�T��Qw��W��y�����7�A�/\iigI[�~ٿ^�T{��1=��y� 	DM�L��nB^0��N�շ��J�A0&�t���j�ک�߳򋖮�K���v9+�����v�-�ޔlO����>�/�� ���	�V��9�b���3��~)8��ì:Y��\Y�����T&�S�9�RGh�s^Ӿd�b"�b?@pW����/��C��9����鲒K#Cz������O9:�ˆ����:�ю�V���Y��"c�	����V{ ŭ�r)韮�m�R�t��=�N�Gu�#U�i�D
]��36Z�}�u���,�c&����Ye����ac�	V-�� LP�6��;<�!�����Xh����Y$�
W�L��Q���d�1�قsמ�8�.�`,���[4j��P:�\�=��,�d�Y'�����h#?z��3���L��	EZ'�F��Fo���6���=Ĳ��J�-�7"J���%�t�4i�Ύ>�RT�]Y�ާ�W�|��̙ Ŵh&�d�|����I�������9��-�H��ŀ�2��"�m��i)_2ʙ�������Hd�q% �$6�5����&t��3��%�zǲl���Q	��R��_b������^�i�L��u����y,����:MW1L���)U}ҭY�sZՓ�De	��cB�q~A�#gS�׈�~x�<�B������Vo�%|ο��-�I��U����}����D|[�=aP'�Yo�)0���6��j�I�~1.e��[�\�(�ˠ��B�~������(�| >�����h�1&y%b����y=�7.hAjQ�7�:<�}��(���K���Ŗ�
:��-�e�!�,����� �I3_��3?��K+��e5���zP���7/����QZG��"�#=Ҩ��5Iس7 �Mr~ �v^�!]��i��6�Q��1�(�w{��#���sV�'���J(���~��+�R���FOo�Bg�tK̯�tim�����V�jǺ��ۼ�K�O'>@mF��v}�lv_�nT�eZ)��}XLR/�^@��?QX�U�)/J���z������D��9j�Ds�iƇ8)��aw�˩���G�qda8ը�%m�ac��Y�V����8M����Rc��qth�v+�#��Q����F�G�6l񁫴�2�.���Aĺ*s �������ȓ�fӎk��DP\S�a���E}���{�>.�m��e��H����X��P۝b�*0�+h/�2m�9�����O����2E�(E��y.�;cr��N	u�B���%�`��.��h�g��CĲd�*+)��=x����렸�P�|��
�G�<�l͗� %��$G�j�~ɣ�����>lc�blM��ߑ��9%�fLXI�o�;�
s����x �W�t<Td���F��un3������{b���3~�f=-��֗:%������Q��dқ��L�ė�Eݫ�&�l\ח�,^`p�
��E�3�Ad��~���FD���rX��o�5M*���ݳ����\l`����3�LNX��K�H��%��>y�Y�j�6)ؓ��$=5�������1LA9���b�n���Y�8#K������fq�.wb� +��oJ���C�7�,~i#:#�p������"�yR|:�z������b"�a�rpJp�D��:9e����>�Jz��s#X"�mM����nޡ�1�%���� K:��믈b���D�H �'I �BO�ܚy��iz��4cBYD�7��"�\Y>u'�O븤�f�z{ �P��F�bh�(cB0)?��0�3מ�A?����Tim�}VI܌e5��,��C�s��C��,c�0ztY��G+B�Zw�E|.�}cJ@�nT:�0��w�� XΩɉ�U�__��ײ��]�kdk��l�1��7e��i�.��U�l �G��p?��F�����d>����4b]qS<��r8,5z�
r��-�:�X�Z�\D�MB`J[\$�	�|�Rc0Ga7B���۪���/�c?��Sv�5~�MP���Y(BU�C�Le2��o��Wrb��O Ɓ�l��?������S��>�N��S��U�a�np���F=�߅���C�hDi�$I�<�:'�T�C��/D���
D�պ����>_k[�N(tj�$mr,ާXt�0���w���pL�qnY�_^,�!_�z;o����TN���z�ۮ߼ 2]�ś*����!�H̕�����-�� �o�i��~ ԙ��/4Uy���V�ڠ���#��pA!|���n�FA�$�a�������k��pD�<���R	��W���H�R<��4���&j9N���+��mKN~J6ڌV_`����iQa�Izv!8A�Q��=��@����ME�uWD~
�r�[*BnJ��uM��p�F!���`�<Ļf�|��5�Z��B0Jh�o��&��/�����[�9�}{U'���8�͞�k��S�^��Y��fTOa,���@pJ�uWl^�R���j����)\7� �d�@�����^�pG�}��x����0Y��t�}�|'��.d"���l!U�&���2��БB1� lԬ��� ��j	����@'�Y"���"sv<�(Z$%�-y�,���G��	J3�j	#� ��JM��&�>�]F��]���w���VjH ubI�ҭy����o���%��/Uoą���p1J���������z-e>�����.�Zl�&�=l���=u��T����θoH���
6�]�Ih������a0�mKA�#�	��K:r"��z��,�Zw�Qr����-�ڸ����JԾ���#�9$���&&�ܚ��<䘺gCl�;�|$s��9�l�
�|1�=.�5?�*��/�	�E�'����w�:���܌�.Cpz��>_4	���
o}}K��!G�K�A�l�UG4N�q�.Ef��B�$!�JMA�oXe����&ˠ�E�5��D(G����]�����M��e�`�v	,������1��b���Uc8Lo��ܭ�KAY@}������d=4����ӂBz3$��{������閖mseB�_��_��[��}����8�3�
���J�ʶ�W:�B�c�O�V��[�f��������SWo������|ͅ���z�?A��E��K[=;�n��9��b8�n�s,����X��V� y�A�:>��U�/_7�a��5x�^k���*UqH��?L;c�;I�q� 9@�Y�
T���4��[�|ދ��LT��ǭxԠ�.�9��D�����=�	W�D��hvHo,=�V�i��8�>ˏ���5��dUHb����eK��n�W_yS�h�Q�L����7TZ�!�ʘcUj`9�Ƶ�{B��R�+-F���U�:LT�l���{I��*i�e����\����(d\���3!*��ҕ���Y�T�f�ҁ���M������nA���Dؾ�����H�r4!rVd'2D)����h�V;�����^���6d^�^<�,��2���a�l�����
�^�8׾�}:�ˆyzs\�m������(�P���H�w�(�~���&��#�-5O
���H�o��L'��V��	�����W�`o$DБ������KY�ْ8���q�����"� Vu;��$%�+8�����?^C��xr��>�Ժ%(�4����ρ f��x��x�9��?���|���V61'����pJ�Q��l<�A��K�uD��3���A�k�p.t)Zތ|[��F�`�M�1��M/���9�ƾ����Im�DĴ3�� /7�u�LU�+Z=R肧/�H�{T��!#<n+n�4�1�/������z�-!<X�-��!�^���g6Vд[����'����B{.82��Ȩ�!��.����zO=.jF�wؑ��@��s�J5�k�X���?�@��u����#���btS��a�����08��/y'��/�ҷSqO�����p�y����g��!�g(nS`|�s`P��y���c6��Y���m4xڱ:�Ш����В����-UQ0I�|(`~��Q�z��6��;R`ES���b�k�ɱ���	���f"�<��[����b���&�ww�����}�Ժل��-W��F�8'!7�h���2X��j��TJ�����NG��� ����2�b��oá�C�z����uٯ���͖���-��5�)��.Cx�_|�YP�e�	�{���i�]��¿�(S�d�`'GC�+S�#��.IE>(W�T����Q���� �LB%,�G�X�y�^�zn~�"�U��YN�I�C���H���N  �o�T�|)>8N�C���34/� �]�z�k.��-��e~�)���y��z���	IT~��������oׅ�4�ZWUaS��i�o�hq�Ve>�=n.�UE���'���q����@}�*�'�5" ��خeGbKK�F���2�ol���]���{�GA��f�#���My�0�����o�J��^�Y��z�a��(����g��W�(�~�;Zfp�P��7���d&��$�H'��9���6�Y:'�����C�,��˗�����'W���O8й P|o޾�U�X�������Qp8�c���`�&\P�䵅~���%vp$8�q%���2�noH냗Ή�I��Fh�l#[o��&�:P�����1W`��@-�nR��2����^��lx+����HA�6�h����M=����^-����x�a �u ��Ll�����
$��Y��>שQ�]3��D�i� �L��cd��ʒ��(���*��)r��'|�. �(9���GD��n��z(#�����
�z��!�����҇��9#\YV�/]�}F2u}$�:}������s��u$���������Gh��\��EN��61>�WG�@j�J���5-��	��co���/�p+s�*�6��uGڪ]�:m���%�w�Ŷ���<�R{�nХڿ��DH+�������ӿ�:�{+�T�`�yD.�Xf���"<Tg�f%��f�|���7#�}DI��煔�#������G�tr�7*�k�Q�����q[�w�m}(�� �N��Lá�V�òǸ�N#���YK�$�f��G�1��y��\����׷R�@ �N�}��ՙSD��)<���4h�����6yXYV�K��4"�R|������b��6��&���<�D�M(�e��cd:�v�~K~w�C'���.��)��J�zZ���Ce�6��� ����-����`��+p�r�?�I��qЅ��^�%JqYn����^V9���i��2tL_̴��{0�(�&�8��g9��"�!ԤY3���ǂ�R}�����*��M<��n�S�A����`	<���.ѿV�RJ,��Y�z�Fc�kEJ���Y�$���'!���T��
d�Jq�o��s	�xRi�;��}	�A�hp�b ��ó���8��U|5�,B�B�ȏgf ��l�;�U����%AǕU���9)q{�-.� v�~x!���W�ȣ�qǄ�8J�,�v�X[g1:.M�F�OO%�+d3�a�VG~a�ZN�_Jڳ���aݿ�)��$+W�=yvdR�%rO�__���m��V���=��_�@Č6���8xTR��=��ĳ�2.�^�~X���g�.�PX�M������v�"Io��I�;���B���}[=��V�1Q��"W�xb1�pm ꑑ����@�$|���w�j���W�Ҋ�'�:|"���(%�ͺ1��F�������"g:�A0k�����ݶa��6�U���������tm�w�3�^��W�9N6��Åa�v�N/.��U#�}�r-+T?_}�pe�!�w;؂U'.9�����ـ���		,�ـ<��������&���i�ÄƦ��=^�y���4�kXg���*�V^a��\�1V �&!�����=%5�q <T0��\��%љk�� "fOW�CV�Ip�ϰQ]+7#���o�ԥ��"c�[�k���<�=/f����v�xyޡd^;6ʽ&T�R�L�I��]�x��~�=�`�<4ŲZ���4��س{�����p����ΤQ\������<��ӷ���Y~B)0��/MRX͠^�5����y�l�6tُ ��d-�ԉ�\�̀�����\���)�� �����px���D~nw��T)X�n�[y�j+Q���:0���_���D������Lj�G�ܤ��Naz~��6���6�M]��/�f0��
5��{�\&�CEt"�;FIV0I�)��������� nڅ|+jĕd�Ţ/�8-s��d=}�13Z�kBg����n���9�u6i��eW�M�h��)\���DٱD#�q�;�
Q*t_ܸ(�a���Х���Ql�Mǟ��dw9:$_w�q���L�=���[,�z2���t��m�ϒ��,�-��[ůY ��U0������8enr!��ts���j�{GQ��q�y����&x3\䍤����2V��󛫜�!2�ח���d��P���	�ʻ�T�4H}=��[���+~�C5��ڛI
6��hAmGXܛ_�Y<�5�ȟ����k�6�iq��䤜\��PeY�J��0�rZ��Ϩr���W37m�m���	c��DM5����(���+v���f4D2�����4��b������p�b�]�pM-lN�ӍA���
������xm�n��2
9^mfg>`S09^-�r@%zE�1�����ꞏ� ��u$�i�BVF�;�~���W۽~S��!�R���b1h=�e����f�C�8Zj�'�v@�v���X��|�t�p�Ed����
E܎�:/"}�+�#�B�uZ������Z8k����s��b�H�� ��pN&���I���G1���c���
{�bq�C֢Q��Z�7��8�%%�B ���mWdV�꣱��?�7�:U)��I���C��u��{O���=Y8�^f�-�#�n���*���K'g⿞nk��K�d8���u4L�����&f�,�$�ǣ(�0�-9�X�����*YS�|'�:���a�g������$y�sA��V� :܀	�@ '��.,�z|��27�L<�p�&�,k`2��l>�zY��GC��+낑�f�{]����%&�7v�р��a���S!�:*-4^h�d�2� o����3m2E�7]�.�ͣi��n�w���=�k�r耝�/G��<K�g���V�#�.v��(n�&��Fe Wj[������$B|����]nOglC�J��c���jE	���1�/
r�%9��M��ɞju�ܣ:U�]���[m�'`Yo<��u��=�h(%h!�(�[`�M�<�t9�����/�����1�F��!�Q�&��"*��\�&5�E�Й��cS;9��Iq5��h��u���Z��[VFS@8��^NfQS��FI}d0ֺO��,5qΘ����{#Ʋ# ��cM�~�eUp�ڐ��o]�z�B
dZ:Uu��-�G�E�&��	�ּ���f14���Tx�e����V-8B��+ K�4�:�N3�}��<�!5cDPzտ����|�v���� �Knim��YC�H�����n������ޮ7���`��%����YvG-p�Z(�u�=>s��B���'�<q�f8�u�&�d�&z+�E���S]x�2 c�z:`3Y��d
B��A�*Ǫ��(���bjuJ[�QF�Nҩ�����8�
��N�M&��\�v\X{�d/�|��_�bOD�����	�߇7\Њ/��]��߳[>xat�$��i	�t$�n>��b-�7���)��S�xdN5h��ó�,`��
��*���Ѐ����Q
		��Pr�=�@�\�_p���H���J��!f�`��k~kv�4���c�!�pU+���̃�[$��O�G�b�����P�~V)�Pg�3��]I���J�`�������k�-qS'�j
������K�&w����X�u3��`s��JZ\��8�#��:�7M�15GMQs�,��1����E�d�_��������ԥ�i�b$F�v�bZ^�e<&�6��- �
����̘%zd_��,D�������x����Ke���*���l�n�J!��zFKy�$�~R�0�k:��;Jn\*�MZyͿyb��P���z���|��J�L���~�DN����pe<�KmĒU^�;�\{
П��W�r�o���ߍɄa�`�e���L���#���D���[�
��A�3���F��$��q���8W��[q|�x����yG�WȰ��;�s�)j5��Kĳ�ߑ>�=��V�v~�U�N��MGJ� �m����X�ٙ�^h�\��X��Yj���8��̆( �^w𫚪�f(`4�Ǎ5�5̱���៑�W�X�a�ه�>�M(���-���^�E`�~C�W1�E��L�Vl�%��4�j��e�z�����d���)r�u#1̻��p�UD�ume��|xl�JoK�vJ�JFda��T	fL�*$\�z�Ѫ��t�G߲N�;��fD�ե��Ԉ:E�������/'�gY���Icaa��~�6{嚕�K/��W&iQv�Ul�~�a�c:&/��t +O�Z�s���)*.���Ψ(%�T\;Г��G���̑?J��iؼ����) ��m et�0Ke�����NU�;~�Ô�>��K,X��"��~�� 0۲��v`�n`;��M=פ��"�cUbf��b;f�n���V���)�Z�g����ߦ�Pb�eF���3��������ZOJXVGQ��1���]Շ�-��-�����G��50����\m�Z�ۀ�a؛�"�Z�XkSLa�z[3�8��qcG�\��M*�3�;�T����f3��U��8��Fwh�� 6lX3I�!���� מ�[�,���� ��oMن���O'}r[����p�6:/�r�;	MX�.�9��T����L���zbb�P�t)|A�7H�9,<2Hy��YV��-���_�vl ��33�S9�������U �'��z9��%�Fj/ 'G�i�HCh�����t2�X{tD״ceJ��'�O�L��Ŗ�����	����˕-be�"��RL �ơ�[��`ݾO�?~,�
��qࢃx]h�DJp]�Y�uv��\\�qC.��KbL%+p�c'�犜bvk��\��y�������A�v���w*/��V�dA��+�w�*E���GVLv�k%�+��7�(�p���¼DXҿ�q�-M�(/�"\��#���Qɧq�����_�4@�z��ܟ�D�4U����Aѡ�}ê����6��!���LZí�ezT���<�;N�Ve��:z�jS��}�
`g8��_H���i_���>"��qiEy��99/L3xyY��cIwDC]��z�q�8y��}S�s��rz��P�#��B{I�(�
鼹
��`�A^Z875��%�1tn&�ë����XS��Vޞ�G���Ӡ�����~ֿ�0^do#���Է�R�q�	ͷ-$Y�1	��C�����#.=�"$Ed�E��CwOzOj�}���]:j��rl��w��0��cΎ0u�csx�0i�HH�z��4B��V��fMJy�ף$`��_}�}������Qs3�2�-4X@Z�PH�ذ�Ӳ34:�-�� ����_�V	�Z�lR�F|�M���	�	��G\�_HEv��':)<�&��H@Łb�Ņ�ʘ���ȑ���+Q�m!iu%v�j���3f�F̍��B9O��Ҝ|L�9��I�_=���j��N$L`�#�I1��bn��=��gh�Q��3����.���Sm��\&B�Ҳ�lÁ� �؁�J�)
��<�^���ec�S��ac��	�n��y7��*�Uw/�����j��|R���J�'j>gI<�yK�������@�����l�{�E&��ޤ%��>��2'�U�s����!Y���|�&�X-�I2� ־�V]�����澂�$�$�|L!Am�l%;bٶ5�E�<k����)�M>Q����w1�����`�Q�� ���Y�T|�kN�:��B��xv8U�{��-l�Y�����t{��bDC�	�MM�Y���zP��N��dX.�C��N#D��D�>��3�S/ܡ%󂗮��l��vd怃o�����e���@�4��K�����<���i75J�	�Y�b�*�s��S��zrK�Fg�����������5��_Ad#:������W�i\�����0@���+&;��hU����,�b���	Ѧ�1�XOc/$qab�>���u��b��E�/�قz�}���	rFU�9ȟ<dɔ�Tv�~�U��+�T5�~_�o�wV�`�����k繧��ry[O:7չ���l�A�Q
���!m��V�'yU�X ����(��Mwf�
sORI�kA�����d*��=����h���$�R�2]+FQ'��L~�V��=��Iv9����X^�`EvT��)(���>Uq��.�.+�)��<��Z�w\�g
;��w��O~Z9��BnDt⽸0n%��P.>�xJ��P�g��t��UmA9�TZ�T���/y,}�2�'���1,��@oDy[M�G�}9r��ͅU�I�o����H�Y)rk0�0�/��I̬��vt��7q�����4.��!��g
p�En5�pE���x���7�����|(f�wP{sĐ
�̪�m��Rn_��m�+���0�C�&[�Z+�Rq$P1S	�*�A���#]T�h�J���t�����Cò9pNnHc�`K
�1�=0�x3O��#4<��Z��"��Bua0�R���1����d��*�ds�8��;fö �GҼZS:)K��D��'���i�<��C��K�ݶV�ű���j��NAp����(�9J'�2�k��q͞]x,>����Rվqj�(���'�+�z"/��%�ԤJ�p���ų��|�w�C�26Bf^���=��?�r��G�9V���,1�X�� :���b�qy�3u�u��M���\��Iq��U]�sH��'Y�<�dk�ǫE®��s�̕x7��]7��<��=q�=�>G���Hj隞%lku�86ݚ��n�1�@���8p)r&�O�O^�4�%R㗪q�"0w��z��i):D��%-97�tg)k+Q�^ݍ-��l��}R%:u(�|ƪ�ԧ0�ǡ����$�к��+$R���Kޗ���V$	b��"�Υu-��{Y �)���2 N��1rx������r��	%S.�Sv��p'� W�RK�#o�[X�I� 3������A�5]C_��d��P;��@��U�s�E��3�����+K�|a!�=�0���%�r1z�J{q����k�,�Mׁ��c�CKP������c��5`3ht��ڇ�/���=IZql�d�U�8��Ka�RC.��нl�8��Vb�%w�7���E��C6Ɏi���[�N����1��aH b
��8����+/f	|��ؤ��Tʶ$��������>��w"�'c~���O��ٹ`x;���3M�k�n�j����vQ��xYR�?xݏ@�����+�l������c���r��%�:���E"������"5뱨M�xw�R9J�F�M~Kɬ)�̱��� /���QQu��.��0Ͼ0���HB�h�^,�&)>�5�7%�:_i��8���f7F&�UEy���@���Gg`�zǃD![�H�y~7 ��Y����A��*!���B�^��Ɍ�-��`^�
���������>��zO�/r�CGO(C�����=4�-E�֛T��`� [d�����u�F���_~R
�n8�Y+IU��7����Z���w3>���oh�\��w�9E$��tIJ>Ъ�)����:,mĞ]��W�~��s2�)��#���σF(�͉c�)�5���{&&�P��������@=�B�r�Y@�ҧL�:z�Ow5�V�G�i_����( ��Z�7-߬@S��Չ��[�M�4��nq/��У�lm��������#��� V�����s�b(��cH��ΪfE^ԑ�x]8A�M������+���������ҕ���7e3Oث��+<�K
w-6ϥ`���A��B�0ߕ��[{�C�qy��,j���	-�O��O�s�'&ҺsKUc)�:��i�lh�v.	��E����TAe"Q���NҘ�@���s�j
拭O|��<�9��쳱}ج`��i��'�S�T^V�k����������!H�Lq�1!�#�_Jf�u��;W�����ry�Gd5#�_����Sf���Mp����?�q��28�9a�~>��m��&5�2��������W�6��i���>��K�Ù��oT<vw���*`Ѧ)1	�Y�[�#�s�)��^��ɓ7D]���9O�šxzfǴ���Aq*�`<�����D��c�i��z��T�ٜx4�hº�\w�\�(@H�1X���#�ٞ,��nB���A�v�6�1!?C�@n?��m@(}֪��~��Y��G�����"�-�CW`V�_'ye��� w_@���05���q�[=ty���	W��6x��K�}�S�����lb|��[4�L8�;�C�y�Og*���/����Ki];x�'3�e�t
�y`�"y}ܿŠ��ɝB=(�>7�ףdҹ�p$Lqʥ�Ǯ�h�#����y)�Ll||�(aR���9ը���G�~f+6�k��&�3XHgIn�ib�2B�&P��v�
hz�z��ae�: �څ �8�k�@�vP8]�-� @=#�@i�G�yE�A����L_h��f�
�q�$�z�#v<eF�L�N� �i��N��M��S:���*G��^�w�֚���Ub��wY��O�H7�b�����-l&��ok��Ħ�	�3������#�w�JW����6(K<��]ߕ�x11� ��CE�L&�4}S%X�U�Z��^۽0�YP�=�X|��"V��jプc����]M(9��A�mN�]Iж�ܭQDM���c�ҟ=>�{`�@*h����@H�����1�9�"o�!š%����ǀ��v_����%��l�]2�:��iq;�5k)�6��3yTΆ�=��at����H�b
y0�z�a���KV�oY��6�e�0�p�BB�9f��������>N}���Fv�l��[��.��x���;��%���\�f6*����L�~Gb���տ{�P�vӞ�p�΋�_c����]5��{��X�s���g�h�ۄ38GM���~����'^�5З��3'�:~=X�Bo��IA�"����I�hTopވ�֎"#==qӛ
�ְ~	�)�*,�b���=��v��M���:"��fU�zdT4�o�o�+�,Q��;IP�x�ϧ�a�r�%�qe�2���`�v����e�
?�BR1߾
��c䤝y~bh>�k���*)%���Y�x��z�Y˯�^���h�zCw��-�fuU�M\R��C��" �]PL)�N�ѫ�+�#f�1��ce<<x�2��K��|��XMP)�S2�FT���v������q�g�>�6� �������/��������ɞ�+n|�ƜU:�Y:�8�tN����X�;�_��U 5T���W֣���>yolV3%r�j-�WT����헶����4�@W/F$�����gc�G�	E}�gw��Z���TPbũ����׭"-DH��,��Wb5��.�yR�H���B\���_2���)s-	Q]W;~��;�J!f�Ȼ�V���EQ�%�&�M�2��}�'�LC$��[�wΙ>kɞ�9���t�9��K)��J=0ÆS�N� T �����e��� i�4�g�?J�83�ʘ���HC�X�@�i�.��4E�o}��Y�78}�ڜC.7�F&���Ň���I���E���!^�B��h
��"!j�?22�ӊ���Θ6!����Â�6*T#0�}f��k��*ђw�߫R��ez^�yZ�l?��E0��5u_W2'c�Ga4V8�B��5�l�k�"f����$��\Jq�k��t�c�"����a.�ȋ��W�0;FG(ܢ�6��d]]��6�a���F2ϯ�5x���A�*]uqM��㛼�Z�p�m�o�`����e����e�P��js�Px�C�G�Ҙn�BAz���)�i�JA��(`M)Dq��|x��I+3�|�s���Em�V�#<1Vc"vNC$Q���u)�N�C!�bC����S�tu�3ĭ���i�W#\}(7��y'>�w��}_�h�����SS�����,���#$��SM�8�8-��hiΆ�S���b9��J`(���n��p��A��ҋ=���?�m.U#�2��!���;�a�2B�&X'�R��//��VE�{ o�8��������]�e�����M�"��ko�w�y��>���֦e�]i�b�A�H���:�Lh��M)�����}�0H����E�%�E���4x�hSt>S��G�+���M'c���72��D��Ȩ$���F�^f~�O���]��� ^�K������� �;��Ģ`����A:AYZ;�b>E����qʏ�QǠ�U��BDG�C�he1,ߧ�k.� ��$%�\�?�,м�Jɣwuw@����ͥ����&iQ�Q�˺���w����������5^�j���nvf����}��Ҋ��e	�'�8A�^���,]Q�ɧ;	6�t��b��֖�]Ҧ�y�j*ʺs�q7-X�l��dθW7n���NG���⧿�����$;>b��δgNǱ��
�� �%r�#����V�'!u}U3o�3X�r��M�MNV�т�������o2iw�0�U���D3W�gZ+���}���&0K��(_���#;5�������z�:,�1���]]zp���y�����
u���,D)�J ��} E��nY${K�5��Ѥ��.y�9�x���U��1M�^���W�R壝�2�|L���|�+s:|2���z!�����P2�-<�a���Y�
��\�g���,�uzv�i��Ur�2� �n�y���5uz���$����8ZĊܛs2��k��牕,�r��Z*�_��7"Wҋ�C��b�?��n�PB>:�6�)5��4���~��B�z�>��_�Ϳ^��bԭ�rH
���hj�\��l��9�K�s��Y�9ӋkcՖc��.(��ߓZi�n���6�H�ڱ�K1B�T�q�4�o��)5Q&V�ɓ�Ǧ���$/Q})#X�:6X�P����^7�f3�M���2�z��2��u��y/S���V����)���JM!��2�͇�s����R�'c�B]�p=�n����{�( W�&��ý��u5f��AV�V��-G4S� ��d���*��$�qjMJ��$�,�v�3b�"t���܇��2yi��͡�T���jt.�o*���V�ǭ5�f�f����F���#�.���u|����x��)<P�I�O���#��w_�.b�,��A���O?c��l�U�H�~[F��L�s1ߥ��^�����q&��]Z�4<��m������ ��_ĲHSb^Hn
�0d�/ڱ�/���O�d�<�9ft�Es3�Rd�I�S�#vR��}1R�i���Mq���G ʹ-D	h�ܪ��Ď��o}�LY�c	ѵH��y�R%�p�a�����n��b�=�]���֬��FLԑ���.�Ia %_�g��j]cwg-�C�9G���ޖKS���W��S���d]-��sj"ry������d~�4�TsT�6Y}� ���	��M\��Ȫݑ� L�Q::�����r"��G���v��~��s]vB!���I�S��[��@!J���O�h:���[}@!�3�ǜ��>�HV��V�Ҡ3Zg:�3iΰ��O��<�/��`�Q/p@"�W�,�I�P�8�˻uF�9����.�H�k5���-3[~ ��7����ΉC�R,0�lu��N��|�|����$�VXD�/zo(��*½^]���0�L��"?#]����!��]٩���b�EW�A��D���S�f )2r��&��}	i	{w0yĻ�.������	a]�]��������5:I�`�Ӻ':��6�h�99j0n���;M�y�Z��%ޒ��/�g,&�y�p����ό]L7�k���	Y����t}��gI��	���]�U`�����	C��=��n�(�};%��$�o%ha�_% U+�P�nf�+�|�>ЌUo�^���튊a8���Y�CdH"���>_���]��iA����Np�R�.I���s�
^/h���^n{J8\��z�����5^A��2
C���ϕl�p�s�Ho����-ZQ;�4���$�U2:��K9�(*��.�̬���/���M���y�v>�]|ܬ��3t���e�3��V���P"��ج(��K���
w\)fu>�N�M�6������c���H0"g�S��R�����8?���V �Qc�&H*��|���9�f$Z���t��������oL97��vc����xŐ0k��R�5<�j*��HK����%���M��k�2Ge����C��hR�~��V}<�[�|n�/�ۯ�3�±|��~�_��V��3?S�+��_�(ۻ���c���D@wں�m���&Q�`L�@�fQdl[�z�d���:=���u'�u&>1A�����/�?`��؄��y<��	]����2/sn�Q&���[����;�Q����F�o�-�|82�X9��rP1B���e�i,��F��d�	5��m�q�ߡid(�>_�Ww��>�AB%�=\GP�y���~ڷ���݈�#g���,_�:'����`1]����2WVɵ����[4���Ѯ)�b-����v^�-��.k�VT�������~yM��|T�IΝ�`^���;�	��⾺�:�(Ⱥ���DF�3K�,���@�����V}�[L��L�; �۽�nq �S�~����5=B�2���QO�0b�:��U�q�ĝ�8g�� gd'�,V]����8�V^Y����3뜒�G[��|����@XS��܏�
�t+�����|uV�wZ�վŞ����D���/E�H �#>�yk����M+�̨��VE�ZWW�v
�&�I�G�ַ�\|���d;�Ue��sM�9dᤕ�<N�V8GiG�7p/�h�`e����?d�+���]5�[>ǲw@]6$1[3�u��n�����1���ۗ����GFO��f=�C�ޢ��X����ٻ�4l�x	BW�>7�{��DH�<���"8�yt�j-�/)|pP jR�,�$}�E�@B%E>�83�Le�L�*��fa�8�
X�Y�<������fS�=Ir�[x�Bb[`KcE����Æ�,�7���ٔ%bnPk~��G���Q*�S�0n۪M����&�bP:�?
G��T;�>@��?�����ܓ<-t�u�����f��j&:V�㢀�ឦ�t
�g���F~�"q�����_�X_ �6���J��'Σ+���G�"�ʴ��%��v"���S�$,��@�;��-֥[6|m����O����]<a 1o��`|��5P� ]���!a�z����w:�>pg��-�=��/�F������|��f�����q����1�_�U}
�*��s�*��nV6+@$���ˡ.����cY�g��k�SF���t.���QǛO4�)J�S1�aTX@�ݏ�:xC�U�)Mָ�%�������ג!w:�D�oI���������]�
�W���=�E�Mf�[G���3�F�#�(��M����=��kF[>wv2��:����l7�������tt��e�;������j��o	#o6��+�;E|��yȦE��ѯ�M��i��;X.��;�&]ƪ�Ň�L�v Ǐ��5c3 җMʦ�ɔ𹩄Bwmnl���e!�!d�$�Rw�.!?�jz=��9���u�L�U']�h|���p�%��	�VÏ��ycy��-��*�WK��v8�0�(^������Q&��6�P�KP/!)���� S/���U>����p�3��=��
��+��(f6H��&C�S�?Ĺs9�Bӛ��7���b��g����(2�4z����R���u�7�tԒ�D�TO���=Lߍ���'_�x�`�4/��!Z{N
��I5�
�!�����E|�G�U���F���杆�%7�����Y6�i���t������ͧ�?��`V�7LH�7��,p���!��o��q�,��s�`֔�|��Fۓ������:�<!�w��	�/>?-��bE��_�}�/V�l$�Y�G��iG8���3���V}�K�g�)�EK���z��P��<"o��(�)��������G/��u�j`�+	�<jT~��:Cg;�w�7Y뢏�3�t���$O��:�$�^�'�^�BG�[�Kї�\�U��ZMd�I�R`1~j7_qQa=NO��T�j0��:%i�U]�Y��4�����^S"D��Ъ�*�u���n���X���?A����"8���󀳍^�4g�*����KN�[7-}R��&�Vj�	�A!Ӌ��ڟ>���r6.E*Ur����כ���Jd'�LN�4��D)]�;�َ3���>����7Q�`ԓ�$����&�YW+��IC?��\�b���n��NA���ƫ6�4C��1�ߊ��^��&#$rp�W"�/�/������B�,,DO�u��L�2��Gq��"�R.k1�
���u��aY���& ��q�	��T)\�_!�g�����F��X�۷Vm� �&/�H�G���ϩ�6��ܭl�X���p����:������y!���Ƶ�^�nv?���"`/c�mR�(H�͸�`���+�߲&�L.���[�ob��e$uo#}�Щ�CE��o� �qLG��: �p��+s�BUPk0�[EǶ��H���H�K��������?�`_�
����_ï�����i+�GU��'"i��3?WQ�KP��]%ِqy|Nʪ�Lȸs�����Ђ��;�n�ak���$�ڨ���c<�� GF7�Z�q=����ֻ��������t�M4��B��~o۝[H�r�d���ws쿛�C��Pţ\ �Zt��q��'GmCl�H�=:��aR������_���(� ӇrZ���W�҄>D��� O���E��)?& '�%e��6�fbm�n��XȰJ�T�C�SR�n:��sl23�'F�. `p�0sn6�0�alYuI�[u�(�����@�8�mh�
4���T��jT��i"��E�� ���h�ܤF�׊�b�
F�������j%y1
+�;��Ѕ��o�D��3]���~� ��hYX��K8�
�H  �\0�s��~i_����;d>��V̬Uf��ԃ\��z�Gx�{���m�C6U��\: �&��t�_Ճn����s��pW��<�����{����/|�<�,�3��w�
�c���w��������O����[3���:@4���&:���)H'���|r�?O|�/v-�MK�Tn�!�����|�=�so�U)h��j�F�N��A>�L�v�p�ٛ�N������)�V�L/��]׳��A^H퟾/�ý�
3���_rS ���䕝���)��yC�\1�f�	Znzٍ���S2���
"��j&��3�-&0�<���ɯ=�T�5����m%-�R�魎�R���W⯆���I��E��
&4zs��(=iC-�M�b�������6��@%�,��!��F�5�wf,�Kiu<�P������E�"�e�����P�^*�I q�F1�ֱ~�yrC�Z(��Fp�� ��^����U=é�lR.Θ&8$	I�*��ȗQB�6�f�K;�:z������ʵ����9�
���)�im�HO�	=���y}֜�w�6�$�Bf4�{o�/p>@�o������q��h���4'\	�O��c4�:2��-8��T����#l�w��?c3��0d��Q9����A�u�9�DU-:�^&��!���ìa��h6���4wWknfZ�f�8q��΁�X�&�5��ٮ�-У�G��'�v2c�ʞ8�Vp��(��H��6��J���XPT��x[�[��oǽx��
�G�lOS�כ)��F���p�f�> ��J�P!�A�՝�T��,ݝ�c�F�P �e��m^G޷�M/n#���AٕKy���v���3�V��N�2�]J��n�m��T]��rA�,�����t��x�,l��f�ȿ�
&�^L��	�1P^�N�&\� ���
j��[q������؃���/f�	�q��oD���i������~����O���?�ğ�6T�ƃ+s�G�#�8�"`~�	��r���G��&��k�R.��ä����qE� U�&�,�	z�B�GU���>����[�'�����Z�
�5h	���Ϲ`�ϕ��R��H2ʅ�J�^t�J(
�q��	5��n-�������y[Ƨ��H+��F���p՚�j��(7g�L�b��a��V��M�:��Dq��>࿛Zz������o��TS@z���	gtǷl��CJ�u.���VBK�O=Ͷ_I���K��K���w�}8&��:��k�5��33�\2��\��c�R�R��zݵiyM6�L��N���o�fo?ēG�S�n��Cp׬rn1�>��f#T��s>���؞4&�?���5�lq�p��3��������"��>�{��{�:,K��-i<a���%jP�e(���%�d��1E�_���S�n�.;Y�&D��	��]��XAtV��E�;+��P�}��c���2e4�Gʪ:QiWIap�����~|������Z�����k��9E�)�#���^5��qg$���X��η��]�"=�s�s���q�wc�S�~iu�tW�\�݈�֓�YC'f�g�k�a����B��a��>ֈ�c�p���X�o�� �f��ڠl#�`��¾mra�Lw�b����lr���@Ν���,�iߊ��G
I�]���* d���uł���+�Y��Y���?����314nX�z���VN_��bnk8X�mUL����=�����zNB#M���:Q&��	�������N::
��g�5�iT�3���F��6eqWV�=����C�#T6p?�����P�n���{�*��ڭ8|���������gĚ�Sk�����g����ж_�
\��9^���ۯm�Q��yy�&9��jI��<m�`ǆ�5z
~dג����?&���,Hj�I���q�lĬd	������x%s�J�gԈ)IB�H�ͧ�Z�җ��5h�Ҿ�����y��oi�,��[�5��m��5{�E�I��v���5�a�k�w\��ٞRIl�5l�WKX05�Xl�u��e��s�D��7V*��u�#�Ճf��n����,<7�y����.��8�i�:���Et�
�,�y�tv.���4�g"���hm�B�L�w�u�s�1c�gY���!�+�^�bF�a��)
��@�)08�c�1��D)u��Ӈ���yR� 7�%�T�MXJ�!��1Ais��<���!��{ �,�?�C�a��e<��R���������"j`�RT4�d�8 #�����5�Q#7�5��"�(70d�KAѭ(��[1w���Gn��;�B>򙎔T15c���M��%.��e�h�O��^�~Q;F���CY'�x )<��(����#���1
�e?Ы���\5Z�y�[���	Oy��JZe�0$+�G����j� �X�$��]ö{)a�:�rQ�7{��&��cp��D�Q�Q>d&tY8H�6�rZ?Ҹ��0�3�_-o�b�@W���/"��<�=��8Adt8�H��U�zR�	\�L��Hu�;RVn��-��i� �=��$���9QoG�m���HcC�Zτ�����[~�����THĀ)"KnSS�^��V���>���w����p^ņӼ��)���=߿��e��4���ܚ�v<�����MVz�2��%�dl̈́��&va�)���%g0W��yLj?85��k�~����G݌�S�g2M �I�O�+�V��8U��'��`X��D����w�g�M)F����$�����t���������Rd��Cs@rW�c����a��r(�G���tBeT��t!}8�<���w=�̈�8��es8n��p��9k�=�.�)���g��l˹�a��b�{� T��!��c�D������f0���R���R�OGm}#�̽`�l!b�?��`����K���[�K�=�|�-\Jb�CGg��.בVݔĈ���j�Hh)Qw�V�A��r������k��<��uf���8[����h�WP3	��GQ��X��kL�W"��f[�fA�yD��[rUI�7�1~���UGrf�o^T۷o��b�$k��ǂi��G�w=�է؎{�U2�pA���o��֭g�X>l//G���ړ�%�eX\�s��AQ�ۨ� ��{,�R �v�Z@��r�h��8�B)!R�����RD�K����G�]�H$g_�%��H&�﹔8{���=�r�)����e�w�+1�3���@Tg���F��H\G���d-�9Z�@�����T� ����&[��Q�"Ɏj	�e�mF@�򠗯oh�5�ᳺ�EZ�:gI��_�SC� �i��QQF*0� 8�۴e��ҫ$�u����7s�?�(��E2�xǋd�v��k��ܮ���3�hy����x�?S��
\�&[� j��w�W�������d]˽���S��!(4���rJ�'>���0�2mb˺@<�!�^d�'4��o�9\�s�Wb==�@O1�۹��ݿ�a?ބ��}��spX]y��(99B�*�p"x�n��x���e��Z�\Fc��H�:U�X_~
�{�L|��<��V2h��ۗ�����T�]�E)-	7�D����Dw�giۓ��Ee�{ L3pe���L_��[����օ;><e~u�m.���CH0י}�SPD%JW���TN�J�$ �L�#�%v���SO1����}H�\��6��Bq�0����Z��mp�7��ډ�#,�%��_7����f��y�G��_�3��G/�L.��7y�:?����m۪�rqK���.f\
��g��U{�l6׀G��q�IEbs�a�#*�H'X:ٛZ�S��ߪ��Iq������ׇ�VR�K�K��hv� n��P��L|�k� �b��~�~�ޱ�؄T�z?�]n��įP��|L��[�0�2��i,(4�:xQL�!+�x�̴��|�HY�t'�n�
��}�h���*�ۥܱ%:plA�lMpP��xv��r���-Î(3����.���:c����7�3��Η1��w�v3�"�76��*E��yp�x2`��/Vg%~ �':�y�V۩,�?���h�����9i�����/N��j崹
{�����*`|5]�[�fI1��h`��q�b������Xs�浛P�&0�	�����ʯ���Q�:h��3����p��F�W+�r���`�E���{	�k_�%�dK �C1bn:���x�p�|#��O1ALɔ�ӡ�d�E���auC����4��`ǵD��u��7��L�t��|=����[z���K�p�ة�Y?IF���Qɨi�F�wG@�u=�ޅ�l���>/����R��8��
���Ѧ����^�(��@�շ��.$i	NC���u���@-P�G���I���*�0Y)!����6y���Bƪi�R�N\;S�(���>�Q���W?f�֖+� ���5~
!�K��75��*ݶ?�w��F��	�������p0�8���S�]��)3�zmV��+n󞋉�g����p�9m�� 3i�F$8]*$c���lMV��a|,ZSR���k�W�[�%	����Ͻ��0BCF��"G�b�����f�L�`����P�����-LNk^�t6r����[XYÀ=�0����b�JbZ�[��Y5�Y_�>})�l���֩��M�x�D)��ާ����9�pJ_-!bC-UHt��?Um\�\�J���v���%��FUjW�8#]�]�5��T��]���0i&�I���ՙ����A�% �;e���������C�CE�L3P��joj�+��ؕz�&L6���b�°�ú��2S��%}����+O�e���E�r�,�OP��K��3
"��R~�9��b&��5��_�+���sxl�̂T0l��R�%��T�3��n!�_7 �o��ȧ�~`	� �A�H�`e�x��2�f�v?��|/i�>Wv!#��r���[�d�fs�8=U- �鰼�����ͷ��r�B#1k�i�l�s�H�����`x��a^�)!�E:�^����i�+$������I��Y��&,���+��r��u�::�p\��a���$I�ej���@��l��F{����j5V���p��`#�~�����MM#�B+��a�֝	���ʞ�g��6��/������t�;���G'l�����u���ΔF~�.�N������\����S�ݾv Q��SB/�O�����\���$�H1��Q�[/>��}�WA��6&+�*�.�f���p����2>Vz��vg{��[C$u�Y{��&���9�h6t�P�%����-!b�(
�i�s�7$��I�"'=ɢ+Qv��>��}��!6�[ha�*����5!1�/ۆY�.�H18���A�SJ���;*Yk�cP�t�5�)�%]u�J���"քCz��Z���,��ƒ݃H�x�g��)��05="�|�K+d�PQ�?�7Ed�:"V�4!��%��ٌ:���~�/��qäMh�EΖt�]���nf������o�)U�7`�[/��(���y=��b@�Z����e�C�� �ψ$�c����fTL��J��p�M��,%��H�n=��M��P���w�+q�]���B�E�i�����YH�XLC���<��
m��8{4�g ,�kִ�B�8�i q:4h�L����%�i}w��X2�����N�u&��(�E�Q
W9�?lʅ���E-J�Ω%��Wuyk�#��W���[b6}YL�u��K1,��)%��R��.9�]w���(�̂�������������@�Y�X����޳$�b��WJV�ݲ��I�/|�[��y���JlV7OW��l�6������_<%b����5���Ů&����v%η��~?�q�b��2�X�%PʝL>�|��N��r-�k�'�j��#p`�i�ם��̔t�O��<&�nV�h�s:n��3��7D$��[�o���l��<��\.�z5-Y;(2���~}MGTt �F1�u�������e3}F�#��@C�6d\TI�kQ�9�1�Ο���f����{��bO��hRɼXPN݂X%�����z�#��
>$�q�ѓ#dt��r�w$�ʖ��!ekUt�%�;��I��)��ށ�2ITF��j;(���S����Q�[5�o�&�B ��r�#e
������@7B�����z#��kR#�̐���� �I��}}~����]A`��9CӖ�xڞ�M
��>���A0Fd4�1W����Ę��Ny{:O��V����������%�|�'m9K{U`D�v9a'����	��L�SD׷�ֳ.�'��X��|5��Z�����N��9����1��*��+4Q��r�cߺ�O�����*�6��oFS�h�Õ6��p�k��4P�+����6��h�ߪ�w���u�GRã���np}?�Nck߇߬E��v\���@I۟�~�yLv��!��7�'����o���5CR��FL���Q��ʇZ&��m�����e�] c�|8�	�#�S�l�R3/�HfY.�#N��2;R���i)��݈����_#n�y;
JD�g�|�꒼���"K
3!��5+��C�}���F��^���z��s��\k2�� �oi��)�ܼ��2�SU�f�X�g����dJ�H��z�HF,.k���*W=�2�'^����Ƥg��u��f����v`#����k1�2�Ȇ���k����6\���j��L�S�ݖ� D�����*Z�c���(%���%�Ӌ�o�x�3+Х��$*9�Ѝ+�D[�� �k?������7����>jXw�a��s���%F��?c�ݿ��|X�b����y��y��>q���� )�(R��d�t~��l��M�U`(0@*HS"������1
Wf9���Nr��6g��=!Yb����:C������A��:bX�.�h�0��I����S�엙��]r�#b"ͅ�H$	^]��E��K�I	���Nq,�tbxk�1����C�N�����2|�������������D����T(�)	�َ[�^�)4��u�2dO��Y KA1v�+����됻�%��yr4�|�϶Z ��>$G&㍍f�k�����kY#�y����S
��a(礃�q�=�*��6�ؚ�N]0o*?`T���ؾ0t���������j��d���Id�� �t��ι>�O�t� ���pփ�]�E���Ed̋���⋦�D�[�r��L�?�Z�z=�7���`�Yp�h{"�6*A�� ���%԰?�<��pb].�6��^�Fp�)��{��`�U���U�t!�T�.����Ppm)�Kx%�_	��}������
������ĩ�6������L���l�h>##z2�_�.>�ㇾs�����,�ey9CG��~-`؋�%��L�!̹��w�N���K��*�0�z'�M2,�C� +��}8V��m6'��&A~Hh�J�(GNF�ܪ����6�5�H%·�o]T����'��խIԡE�Dl�?֗�U�}d�H��WoCUHOf�1�������n8M*Q<"o}�Oݚ\��ֽ� Mc|qn�Ⱏ��`a��X]f�Ye�G�#�(^���`:4#+��3�%�S��B9 :T��bEi�=�����;��>uc�Ğ�jD�8����3�Y�-��T�BS��t�����s�
a����M��&]�L��J@�Qk݆�9�ۧHf�������M6}/�.\4rn3`׎޷}8p��tjtC�gY���;�!�`Y�{�Ż`E��m����Q��1Q��@ݮ��#e�Ů�n�U>D��5VgS�L��Z\�i 3�k:?y7>nu��X/�j�����c�������y���5"N?dwA�$��'Z��`�W�6�ܺ�t���#ѓ���5�~���2º��
�mI��U7Ӂ';9D��� �r��%��b!�h����()y`9:K�ܘs�Ê.��"E�L����'���L�H�[�º�<��9�yUz�p/����x�nH�=�U�� ���AZ�U��!�75-[������L5���K2K-�:���)�[4�S���9�`x���������h�ej���lNZ�5������=�_�Ǣ��`���-�M��Z��Icԍ�E(7�sfZ�ٹ��$��v�;N��]/Y�h�0�� �,w�]AN�r�rg���5s�l�N�X�a�s0���)k,�́���L�&�p�,��|��U���7����_�o�s��8Y����s�(��snEJ�
������G�>��8M�j��!auĖ�L��"��Ǌ�	��$OQ4�v�`�+eADko@V��Vf����c���	�=\D�����J���h�P��� ���OW���v���a !�H���a5eWEnh�=d��½���,�{�3Q(�_��g~����*�iV��8Z�9����[F�d��
�K��^���^9�A��f�ߠ�&:��?lvS�]o�C�Z����h��1	C��	��Ѐ��7�'��=}�h�����9� ��GD{C���mEaf�Ok�=0��	�( �Lb��tE~沄f�j�%�.�&�����B�럨�0���u�Xp(�۵>[	j����c&���������O`v1�[{���ڰ��8�t+��P�=����I�����dC���䫗+�ř�m�b�9@�C��X���G�p�� �,~�Y�8.M7OZ��%Z�g#
hx�qt�K%d<�+���p���
K���S��m��ή��Oc�O���⍬�n4?���%m�_~T!���U�m3av&,�n���u�_��ZQ��x���ID_ P7F�<�E���</2� ]	q�z0n�Վ���Y�P�Z�֘m(F���7����p�����4`�Thg8��\ʈ0�}䐺��髒l�X�{��z/�#�z����S���-�Y�i{��"[(��°E'�V�����Jm
VC��|8�*)}U�'��{����T�s��`5��in 
���%�qD[n��s�0��Ce���LFz�l,�`@1J���AB�X�%Ͻw��q�,c�p��I����`N�W�x�lPd|�*4��M{�Tf|������2o`������8O�e��3���ƭ/�o՜���5�ة[��(�^ֱ�޾İ8T�	+�w/�c��bs�6�[t&j�����q�T\A"�)��SR��ON5�C�����7{��=]�����R9�N�8*_�x����NR�՘�DH���_�\���|���F���B0E�q+O��a����W�������|z�	�̺���&�]�����
�Ƞ�=�,�=�~���a��y@+[��]u@�(�@�����'v�ze�n���a� ��L�䕐u��GP��L@.���%�C�ۈ	��7{�VVw͸o�|�yb��Ӗ�zOZ�[���.,�a�J�ay"�$��
�6����	�����x�����ф���3�6Í�5���\��f���5`��#�a�՟�W��l�����N1h�t�Y�$"�SL-�{��{���/�3%�0nU�n���æRW�>FLZ�Ajb��!�>+����8�7�Ȣ�g��n�}m��*DDX�M2���=X�2��U�UO��h���ʮl0�Ak2
I��_�Sc4mY)�]/o�����i`G OM�~��s�M� ����1�~䁁��d	�<���  w�W��ւ��Z��؜U�:)/9"l��Y*sf�Y�x�<����d,mֻC���}}㖆��Գ�n8
��X�}�_ca�����JϩN��0��� �`��[k�z��1�þr�H�kJ�P�}z��G�x��u��l�xe�c��uل`�a"3|�Lt�Y���f�E�N�ꁅfZ�*�.Y��*I���Ê7:<��i�L�]��vPj�c��]m�X�O�.�N'�~	_�E5�S�U3Z�|W�X8ix�	Hw��`q�$�Se�](*��nO�8�R�J�DhΖ���Y�C9��\G_�6���T��.��c/�-��Y���25�b�5�x�� ڂsw��I�R!b����M�6c�V���G�J�-�ߔ��La|$������I��@T�r�q�����^K�{���B��@=A�&�u:��4�}؎y�H��z�s+`��a]���RL���e}���Iq�3ٷ&ӡ��5@�t̮���:��k��3��7�fUD�4��m�D-s��"M;��(��s�	rq|�ns���c��T}M9.;ϑ�����"�l��!v?�p.��RcHfvF��(6�z,U'0��� �Y�C#,��*���,��A��V����h�C6p�����	�J'�6g%^����K�{���(�I=�b���猭��N�z����D�V)���-ړ�t9�����^ݘ|8X���N~��Y�ǘ$��W��qk/��q�K�Y�kRE`��o3�2��b40c�}�%��,h��reD�D#T��:������|wI"Q�*�{w�#���.� �g[�I�̲2-��6���gx�g�i�����M�'�b��g3��� ђ޸_��(�F�k����B/p����u�M۸*'wG��&U@���F�C~��һh\��F���^�5wss�3��Z�	r����(�Mc/:��T_Z>���8i�kЪ�z�� a�%��hѬ��@Z��۝E}�(.�fiJg�z"nL�@��,@�'=�v��ŝG���:�p�7�n~J�@�Nnfco�*jC�^uhR)�	�����t�����a�j����ȋ1"I!���y˵S.��w�-�4��E�z�"+R[�%�DF}vy2kjzW~��(-a�zt����pUm�
�D��GcLj��;Z��i/�6x(����\�a5k��\bv��$�����=n׈n�0��kZ��Ľ,yO�3æW0ᅔ~.JI>	bi���/�i��)�/�N��z�$Q2���Ǫn%h^���X0����y%�2piT�5�tC.5} 4vu�:2:!�?�����s�ɃIr�I��709�����ǰ�@���0\+w�4��_�w��lk�P�bf�EV��k������w��ҽ�>Q����[pЏ��j_�ǚ� �Q�"z"���ϽL�n�#�8v�2��W����f�
A����e���}C-v���(�v�_R���-�wx�g,>��Ɏ���^o���u��ld���y3�����0Z��׾���7'�T#�)�"6���Q�њ*���t	�ѱr��Ej @JQu���%4�%?����u9�.�e%�r�����>�A���O�gc4=�%�)δ�a�ٝ�@{�j�GU��|�Q8���mZ'k��bC"��Y�����i4�����=A`5?m�=�,A6OJ���^���-��׶uO+��oA�(�p�㩀;H��v��Ɵ�=�/��I�ܕZ�P��Nw����Mo�zT��O�CF	�����N�%�E:5���5Ϩ	�މe�7`61�hs�Xy��Բ�n� 2y�EM\�H.�Zh�P���4��X��m#��S����v9E���� ���%'�-�ݏ�l��u$1����ڝ���P�O>>�<�0w�j�c�|Q��7��#��B��`��2����(��ȏ��2D��(|懲��=FK����>\C2#�6�`L�z��<+9i-9��ȹ`�{r���P��տ9:nU,[J뭟Y�o�	�6�LvГg4{xE�1Œ�8U�ї\�z�0�ú~�G��V��X���<�қMu5h�p),�q�u��+�'t��Q�x��d�DS�Y3�[�W��!_A6���d �9�Iw�I������qE�/Y��׭��s)0���������`���\�> ×sg>�xD�M\���&���	*���r%0�[N�!��9��M�PtVs̥/��Z<����7�_ v��<�&�b�����l-��6�O����G�T�m�y]c� �(D����GkZʘ���_��A��P�>���!�m��E�pBG�b�X��kNR�}�����'!W�cJg!c�k�$Z�kgV\��R��1����.~��~��<4S���Шw�H�@$"��Vf�A�.ޮ>MY��C���.���D�d�������p�U 8r~ ��^��@*$Oxh�^�	�|,�i@Ӌ#;�ɵ��hP�u�P�Gz���L	AD}8c7�n�)a�B�@��U}��%��l�1�#M���L(g5��ER��y���n-G� �wQz�C�F_�
^xSL�R
�[�-���[`��P��N��2k��W3=���������c0m�
fN��R�Z4��6�;����bA�h,�o���pۙ�Oqܽ[����YϚ�iӗ�w�-��!�bh��ͨL��O$�?��ǥ�K����E��(��LE�'�JP�!�!��t�l��?��&Cˑe�R
��%�� :�X��3?ilvO?!QS��`3ۚvB��unOt�aӬ�h���u�v}6��,�;Q�����/�]��4l/���|��[�Κy����6�#�X}���O�/������`gV�_�U��Q5em�;���d���K��.����+l�3�>������}�)
Ҧ�f !��(�F�|�Ю y����m�-��gA ���D���m��1�֟:��%�
�fF�l[\ĸ�%���`C�]QP;d:�|Q�^��z���t�:JI�Į�G��q�4��[
��A?�b���
�0���ϴ#%2;�	 42���IP)m�knue^�g��C�o_װbhF@Jd���`qZ�ep	� �`ΦT����ŽWܝ�Q[T�
Uz�p�0T��V��Ե\z�e�͢��>���7�W��a#�'�q�e�0sx�-����ߠ��l(�Cit��4 �/��PoO@�Zw:` ]�E鱵��@'��	�v�VhP�!��c�6R�KM�.�������|u��&��i�q�����\������(&��#�%Q��;o�vNe���]n�^(҄;���4��ڿ��U��,�ۑ[��Q���j#�Vέ�ͮ��q�{��$��t&�ճ�(�m:}7��6G��\�O���V�b�Ƃ�tF��9�-�&�i֊�d7Dx��y���[�'�rq��Qj�.��>k��^�W(�)F.֊WY3�t'�؆�O��?c5��M��%y.6�ާ��}�Q͟}�K[Ua��M��h~�AY+/2�ϧ+���(k4W��"�<Z�pNgP�PB�7�2���_�b<?��:@�����o���[�B�Z���[��\DIwN�j��	u#q�N�a{t=��?o��Q��r�?�����b���~���GF�|t* ���/ms�evT���+\v���D�Y+�6�i���A&��*!Med�V`7(\GH��ʂb#��
�����6\5���i:ۖq�Ƴ��<�ߥ!A�1���%">�{g�川��M���@δ��!��U����X���6Xe\��_�fk���-D�O�
�a6D��i�f�P$�1j�a9�;b���"V�.D���)�����]6� ����4_�݁E���M�d���/o-WIJi��6w(^4s��FI6�/$(/P"N�f,�
�@�^���KUע�V��L@�`���2�m8X�M��s��):��0T�D#ԙݓ��\��^�+Q�V���_"j-�^}�������Rg�Z����1a��B�Z���S���tMC�c��Y�8䆴A	��뭁[HU+*�b���������턬�H{��S,ݕ��N�_t�Q�+/��rp7� �g[tD������*v �&��o�p*�/^�7�mz����oD����,3f�J��m�Y4dQL���d����)���ܻ�/�h��g�PD���S	�C����BFh
��	$�G��f�K�ʣ�ƺ��˹3r�f6�{`��֧��|�. ��r��1a�*4>]ۘW]:I�_'0�Y��+R��MQW�ϛ�@��x	G�`������M��Qp�
�8�8Dj�5���R)H���`|�ʹ/*֞��T��dR�nH?�J��w�f:�`�����]m�s�ĿJX	��Vy�H�aX�}��GR���Գ4M���ΖJhKܬ]���1S�K���ɺ0u�Ó�����g����"{�k�S��S�D]s��]%�<�6���"J��.��"9Œ�*�UB�������ao`h�Y����Dؖ׏v���i�A�������+��֬�`��-�o��8s����/�׃�9�Q���<�W�Gϳi
.��4�ș�u�S��D�� �u�T+Ia��#�$Av�y��[���5��B]wi��e��������-m���zn�Q���b����iBt#-~����&��VvҾ'�C;����q��7�#x˲��vk���+*��fۆ>3S�m%��mÍ��uc��� De:1E�-��Gu�
۳4���I
!r��D�Oq��� Td,�h�ۏw̨Z���/��z�u�M!:���#�6ÂH��؈� ������ʲ�>�4��H�ы{�#�/�&�$�ũ|��c۹g|��`	������N�����2H�Jg�,�Ct:�1Y��C�I�f%��Q� ���^qz<�!Օ�^t/�jY��I׿��f�Ԭ?�z#�
г�~f���UDY��}� p���N��~�\�a�,c %�	t�:���p55���c
P�^���a L�=�eŊH9W�n�7��ǧt̩���*�졄LpA��&57;�٦P��'�� h�!�vh�D»}��[��ax���BiŐW+��Cc�N&k4q(i�~"fq��J������E1�Ac��V�G�͒�֠����gɱ�S�E�L.ZC������n�Z�n!&r>�w�i@�31xxm;�_}�_OR�c�%�{*0|�)V�2�&�<+o�r�۱�`���>�$$�ZmoǴ�Hp�PH�x;���t�]�E<\���8fq�g٪��y}�8 t��-L�����ڐ�����9/�
�%��T��<,	�'t��w��u�ˠo�HEZV3\dݧc�yA��}Zs���Kk+G�J�����Ȟ�OoX� m���<�^�i0���br��F!K#t�_-T�b�Q=�e�<��#���c�V=a�%@i�A �{����.n��K�܈�A3	�?�pN�K���8��=6{��TT�V����\Z�
�X�k+"TV���8x6�C�Z����/ϕ�o���'		�7�v��F	������L)MG�/�W�_i���Į79d��MO9���?Z��Oq�����t���5��nT���4��KZ9:啽�0���5Ġ(W��F�f�8��͂�
X���!�U���j�����\��O>��*��C�0��~�gC7Q�����㣅��lMk��S5QY?;��� ��)V��ڹ\�ӌ��_�\Mv�Lӑ������zt1A�`�1�{�(?)��I���VR���R�p��kl�62V�2���9GCE]�t.��ӵ�Ժ�Ygu�@V��[bE���D����Hb܏��[ �<ҽ�<MA��b���J����Vc���R����Qi�e��0����7�.r֓�7�Zd)�n���gQd  �P���]�H��]�M\&�o��LH"s��',	��u�`��{��I>���}�!�7𑙩"��'Hm�5���I���!\��O��g,ԑ.�!�5�UNe��FsT��ס���J�>������I�q��䒠�N���[��Z�[��6�A��l� ���2�[�W~H�"Z�.`q�A��dXOzã���2׭��>0��l=�D ?�����Ko��W�4���S�l5�[�2��_��f8��SW�,�{uo@!nc��( s���[z�D��J�����W"���Io7ˁ���2��	�q��e� v,��ZGF$�e�#ᯥ0<�RKXM݁;0�O�-&�a�؟����t�,����T��w�e;C��q�U?s�G	�����{�#P�}���V(͎���|��_�P�5gI<.N�4�g����e��iv�-�4��GB�Z$o�/�LǮ�[O���|/��尠�alz>�y�U'��J�z�ՙ�Hn�">.H�	SČ�����NC��fƆ�*��)�-���ż=!n����O���`���
�%������$�.��6N��wM����]l�൅e	���H���?��?T�6�E�k���c->ۘ{O�,RK&�@`����?��~\�+#rإ��o.�⃝~�W�8}�i�lՍFP�S����1�I���JZG��x�d35�y��FZ��0�v{�$��������������E�jj�.��=ִ_��n�k0~{��
[hE�9ٻ�����E�R��Y�ܐo��Iwgs�UmU[����k���u���cz��xDWy�#
땂��w�qӯ�T��� �t<����M$�H-�8���aW�_����@X�٤IO����~�?�H�l&$��v7<b�U_�L�4�uc
r��@�~��BRJ�^�\�O+d"F�l]rY �*�ꥹ��$V��E�̻��KCv�K��6��e]&�F��Â����_��Eݴ��
y7�I~ɒ�� -<�:��m/q+'���=l��n�8*�K?w(ɩu4��b,GC�SH�
��cā7z�P�sH� �74?������C�MU��Ҹ!^��	�i��-
�|���J�ZtD����7?g��wVٵm�VP��5`jY<o�/v��s@��/��5Q�&�����6b���~zDX[eԞ3��B� B���Q���>��4FO�6����'�YV��M{J����t�ד�?l�fl&�ˠ9&��@M�Hj�OvpT^��X9��ڢq�G��d^�׋��ADpSg����.5��J��n��Cq�]y���~�+��(���|Nz�뾐X_�K_[},(����Ѹ����s�5�J�}�փD��Z�Z^�ؗ�F��v���� ���֥�T2�7ѹ  �� �����Z0�_��6��fa�_�@6h�~+�I<��][&��\�U��=�W���(�u�d�KVi��<��D�JЗ�uY5lI;�� ΀���� H�ov�`��o�Qo�_Z���g�٣���Ԩ��Q�,s�����k��-3�O�$�MϬ���(}�\>-OE�t�#OG�ծ�^_Y�.ĝ����:=O�4�<nSe�T��.ѧ�j�����������<܉Z��[��$�슐G���T������$��q, �8�Ύ&0Fr��7�cЖc�
V�R���:��m�}fi�*H��iR������eR#j�i�"W˾�]�Hw�ϟ˥���f�8D�l�h="�P	�I�v��t���@�vz�)�I�~6s���y�\�K�˗<����Q�Դw������%}8�-��y���ȹ/.�ر��"\�i;ѝ'g��\c�������rLU�QGF����8��($7nbN�JҮq�u�6�DA��]�����pI�+���2:s�]�����$9���;[�iME��;A�}	`�@��Ӫ#V����~!����S��7Z[����1or��l��[*�1_�*�:�%�.y`����%��_�v�	Cqޔ�$�"@eh�h���m:'>53W.�y'ѯr�,���]���86��H��nR�i�۱��nM��lڿݘf/Iu�Ow����A����|�S�pZ�xZkd�R_$�a��P����j���,]6�0�6Xt��1��lP���;[��Gz������'J�e�8��^Ot���x|��Г��L,���{����!3m��.R� �Q��,���P�6:2V��x��z]B�4�J���p��Q�cC�@��( o�jV�(M�\E���a�(,H�����AI��7�h�MU�h�'mJS����Ĭژ�e��K����'ơbqJsH��)f�����K�?;����4�vE���87� xo9vv'�y�pC��~�X��� 	�A������.0���shQ������6:��Y7�'!ߩ��+e4U�i�Kf��V�F����1Z1�m*�9�b���W>�H�M��h��0�-�����m{�x1#1��R�^1�����.�W<�g���J�R5��!H�M��5l�M�3Ǟ����*�� .���%�!�����X^G� �F���~b�X�F'�W@]o���x�ȤM;`,���ljDY$��E���H������Zl�Rޮ���D��Y3�D�&@��$���� �t������v&��R�a�]`�˚+d��A����$!v2����6~d�l�#V|����	e��G�R2`�M%��JK� �X (-ؚGfk�ZҩI�������M5a��J��� ��UYe$sF��*L����!�f�&���c�7�i��6��2��	nF�*nL��?�����b>aQ�T��Qȓ�uP��d�K���5��$��X��g��J�k��,��1[2^,Y�R�߼�;�����)1gz�~K̷���b���?��*fn�����ՇK[Jeh��<�BI>��d�Sȯ���7;��G�0�� Ɣ��q�	�|�iȺ#ڪ�}X��!�2s�!jtQLo{8²x�mY������є��~U���i��tR.� (�.}�OJ�ea��x+ƿ\�̎�\�ή�dG*��&ȇ�v����q6^a��X�4�	0��F���ڲ3L>�k���a&��&K�jxMl� ��چ��]�AP2R�g�7���T�&�7dGߏ�y��\�
ea�F�(քZ�%�Y�@E�4�������$�Hj�сՆ0�ʔ\�q�}���3rQ-�b�T�g��y���H�Ϣ.a��C�\~�Խ����w�� 4p��/+��QB����n�q����k$��:`���	��7Lk�
��!rm^\}Y��3H�DGN;����0D�.{0�a��;Kj��M?\�S�1Y���V�S@����!�"�ԏ8���/�9����b��B�#�'��T�W�� 3��A�<-�֠K���4S!6�:���	�\d��Ї�g�M��͵iz����Ы@����.-��6L�:�#�R?�?�A��Q��s�in}��+o)a^p���]܊�� �<�f*����ؽ����,�lԭ���	8o>{�r��T��
�-%��l�]d,ut�'-'�n�%����x����ۄ���m]>�gd�pUt�D��J$֝H�dssӷ*�a��x��z�����U����Haz�s�q��47��Jw�>p6���U�k3�>����E���A*	�gZƝ���(jE@{����O@ӞZ�T�:t���BF0c!H=�ZUP*l��b➳Q�\M����U�?��<<�\�L�>��4h(���슞�lCg����zt1�r(
�7_: �	$˜P�.���[�v�!���=�$�*IIlJ9���{�jnf_��^���`~���<��dd��r{_����Ɋ.�v5�]-X��yY� ��a&��W[
N��yUM�����"6��GJ#�R��l��V�1�)�{�:dIe�8m�V�.�I޿�<��R,�0��{����m�+i}�"�,�`�"}Zdk�c\d�A�rr;�-�Y�f2���G3�#��D�����W��N}���GX�|�XU�0b�|i���>�뵛��{�!�����,Hz����pz�͝��o����S��8	[pT�~k�a����OS�Ē��3"C�	� �gcU�F�[d�9A>��In��!���OV��[()�NW�G!��&�6� S݀�K'308!����×B'){�%u�����2
�E���K?�i����'m��@]c��1z��4�5�����?Ӛ�A_/�;�?���M=f�t�oCת�e��5d9d�[TP�� �����u�
4�B%�׉�-�L��k���%��J]�ϰ2_L�7^��n�l������$��̞�p��?�F�K)2b�Q���y��K�3_ky@�ٺUL^�kˁjݲ�� w�tʸ�wk��[�W ~�ш۞���^��l'歝�N'F"*�RZ
wW�[�)cڹJ�p��';4�:�U�.L�� F?=W?�ag���^y�Kȑ�g��b��]�����О��4���=_Ԉ�V� �Meǧ����=J���ј���<*߷k("Y4�� Q�J;�V7P��+k��±&5E�`%S��2���
��'?u��D��5��!�/&���n�Nٙ�魴��f�ь�7KL�2#W��M[A�E>�4C�\�5)��Vi�sL���B�+����fGW��W��2�ǳ�T��7��͛[݋Gl�y���9�٤¦�͘\:��y�r�UAkJP3���Yg���tq~;Ĵ> J��lн�>d���"O��a��E��g����ц� |� B�y����%��;�6�-��`�2D�ntc��͕F�l9� S���c�C>��Ě��ٻ]��<�F��I��F����+�fne���G~�.��y��MQ:��W�y�L�� P�����:��be� �=��h�s���l����0�M��s������?�O13���q�!4�K ��PZG�W�"~���!~�����V߶���c�SF�CXc>�O~kն��'*��-Ti�A`@��G���m�#
,s�������+��tE���G���� C ��H1'k�ݼ�z������ԣ1y��'�R&�]���!i<�:�J�������b(ߓҬU�2�:H�m{��i�+@��g`�C�}�B��T�Ɍ�4�/��b��c�,-�*F�m�r�JSI&�Ow���������Q¢#�����5�c�*%t�|�9���y��V!� ��w��%t&�k)�¾�a�����eU�	����$�K���{�x�y;G�O�[�b�[>|P��͗���(�ېO�/�X��$��W�.V:T�D���e��n%@g�K]ߵ4�y�6~	�Cٙo�e�i��x�?����0ks�m̛ �@-��`�Z��Fؑ��a�بx��(7tB��iм�,e�8���l>��*��<I�����l�ƸCó�$\B�q���s���T�y��|��;T�~)��c�'�ɱ�D	�h�l6��a�
h��˯e5n~���oP��h@:�:!ؐ���<w�<���������82˼g��.�QT�Z�Ϣ���j��ԭ?�#9O�	�0e��|ۯy��%Z�ae������m�Z��*��څb�И��i��Y��# >���.��@�^w1Ê7�,3�S�|�0�bϺ���C�`�YeB��Ϥ0��Zd�Ta��u�j���"&4G�5���o��'p�R�Ω�#>�a۹[2N��ð,��@ʍM�k#�����m�N��xn�W<��0�Z��<���G��|Y�lp8�!�!N��v�ݶS,ŴQ���5����\f^��$Ӳa�>�C$j������P"Y6:xd�%ω�HfF����~��5ߊ���R��]IuA�F@˾09��M��&B�v��F����%{ۢ%�$��Ju;���2��&��	L�������XSU��J���<����*�
�A�=p��.#�t����Q��Mkx��9#�&hba��0$Q@_�о�%(`�_��G�<5�\���o�KR�1r�%�@\�.d�`��S~��~�*�{Noٕ�s�=^��u�A�h{&f�.녎n�0<D�ٿЂi����ɠ�Os���1��X���)�q�E��h��	�'_"f>�E�84hݰ6�q�C)�Y��	e8�&Pz)Ҳ�5���t�h�&��n�,USKt"�+4[�!U���K�N)!��Qߩڭj���14�Bl3�;x�j�����p@��Z�f%G9�5Ȇmv ���{���p9���{���u�e��*�ѵ��b�NZML���c�//����\�e�7.�.�k^5��$g �e0<���H���$���H|�i5��������_�T�gF�-V�&��V��h8��~YUyJ�V����B˦�YU�_�s���߼x���~m��8�e�S���o�)�P��L�u���U�s���yW]�s-bcL�4<342P�H�@�J��ʬ��O"��O��q�h��.�'�0�l}96�Mn:;�������!O�����N�>��4���r]$��V�����?�~��P���pg��ht��J<�AnoW0'e�h� ����ؑ	xboU���!f��ݫ�`U�YĘ��V�П��d����w���3Rdy�*�Х����+��!�.h�����au�VC�	����G�j3�c�~O����~Յjc��,�R���$0���-��U�����B�\){, ��d������Y�uNN4ۑ��[��(Ё��K�+�U�o�	��rC���w�й;����C�>�3���*�4��/����4}���2�'���Ϟ��B.��J�����v���|\V�"@U�Ӥ�"�4.hqP�2��6��a_i���h��V���A��s����o�]���ό'���Y�rN�j p���8RZDy���%aM  �ܱ���Ǒ�� �[��,�4�:R���ДR�>��_#?$Ky�u��T�|qՏ�V�����P����i��$H�M��1��Zl�q�'�Wl��!����U��2��j�P(����쿁��$LL�h&�*��@�?7
��]`�k�93@5��Y��JPWk�V��d�)o �q��I��|tcE�:�⣀��^�ٔ�w�4�
TV#zt+�D���U�aYd��S�U�d!䏩��m�Rq�����ʄ!����_����e���^:��٬����~�5am�bl� ����@���� �WfB�V�L��������>�-AՔ�1�*���M�/��i��^w�ύ�6 H+��Vi!����e ��l�� =n��?�*�7�,�g;�����Dip��{��qu"pG 5�{��0�vB���T��|�Z�`�� �8[���Dm|7U
kmiC9&�E�R_͌|�jr��,��')~���$���=[ڡ�{���PE�"A�shvV�.Nz :��Ӄ�p�d��Yk����vb�ʞʏ
��jH�`��<���S�[%�:���uI�Y�s�Z�n�[*�dm�Bf��4�m\�L	���la��`W�~���a��ܘ��-ՉA���?��� \���[Z��נ���?�3·v�9`�#�c�L@]?W�(���(�NbM�)z̉-�m�M����	�X&�,�OO�AX��%�Nס�K���*>�U��G��oU�.����/W�Ai�e�z��X�@y<�@��v-�m�$?EK��@�I��0]ׂ�R;����a�'��?��5�e��h���k=jKw�	ϓ(�o�=�E�J�����JKt�<RM���E��ۭ�&��>�x���|t�E'e�k��Z\޼])�iHE(�H���8�Ka��% �>��<�U҈2
(yS_A����=�ѿ��H�C�jڔ��b�쇨��s��cPJ�$t@�q�p�/!Z�H
a�t;����!�9�P�r^ 5"|��Nt�;`-��#�7C���;!�(Q��tNJ2C�fW`Z�ptg�l*ciٺRG+n}�����������8>L��w�΅M�
��d�
9�M>�o"
K�
� �����Ԭ*�2dt`�x��`O�/kD����{g����ڲ�W�D ̻��*O�?/cW�����c#"U@�:"xyN�瘩y��$+��u�53b���S�x`�y>8r���g]��T�5''��1��φ�S� � 9�5m���7�K�`��c�lR��mko]�}Ƣ�7��]��E�"�%e����i��I��
g�� ��L#�DF��>
�������	lwF��'����~�S�6�v�X�!�%���.�Q��ڦ(����L��C�sC�;��5�w��g�8tIW7�\�3��i��7�6� ��+�y�B=%H��`7����X� '=t��m���u��IHqś��d�Xg��D�\�Aa&a�cYIG�w/Y?>�׍����3-ڲx/��/�s�^,UI/"`�Vwi���6T�s
���}�2$���8OL���?D���F�Z�_[��|���9+ei���|���K��#S@����O�(�@������'�?+~�L��qJw���)���kR�*�/���0&.�6q����?*��uɦ�{T�R�	a�TԎ t͋���S��2���˸^ɽ0���A�XJ-{(Gj���/|�N���c�v�)ѧ�ld�
ޥ�#ȓ���.$�jN��&��D����"A�
���7�p Ύ�%`�z�Lz�TYۭ��2�7��F���oiFN��$8 ��>
�U9Z[=r���7�	���ț����mzQ�RY���!9HiG��+W�	dd���廥B<H�Ҋ�TQ�TN
�#���1��m���\�E���o��΢/�Jm�L�ޞ����	��H�<��Bp�O�)?~& 
�C�t����բ^���gn���[�;bb���ɒ��!�m�0���j����!�����h0��R�2~�6����;�|PD�B�w�jo����;��폄��2R��s�����?�����m��� �}�ќ}Yءιb�6�q���>;De�Uz��ڢ���(y�G�*q��4�H\���a��m!�7p�j�LG���ܴ`�j�	:4���x��1����n���3����2z'����p����zoI����iy����L���
�$�����0��Pb�?�7��بX
��F��c
��>}*�~����xW����8 ę��.�\HRr�߭�)�
�i<#Sc�A����w�aU/
xU쒃������+D]�&[nɊB3�V��U]_��O�dm���h�7�����~�R|;��:d��-x�I5;�2��|B�񰳧�t`"q�!��`c"= �v��t��h.!�	�5hЂFd0������ٳ9X���F��K]����ݹ��G�<ۓ�G�i逶�ٌ�~$�1�&�ǿ���$�,��$2�.u���vDX�߬;�e�X3m��jR����{]8Ң�o�n�	w/��(F$�V�Y��t��ν�.]����|�|WHc�����)u�����ױ��m@��h�j&����p�e�����j���u�Ҡ#,�Y뻄&�ꞇٲ�b���nų��Օ|��4�tr��g�����`�Pi�����G'+�HP�X~� �oK>��J�o�M�=Թ*BM�����U��B�K��6^W�}�]Wof"����+�����d����
�W��KH�B#Qu{E��f�(h{v�3)�nS�l/!Ē���k�KF���R��O��$D`�
�6�{�C����ddf6 �(p�[v,E6,F�a��jª�!4�]���U۳����"��������;͕�(�������KC��C�|I;B�B)��3u�Z[�#[���֎���H����N6�� ��cN�mv<}��Qj����a���I����)x�0�'�Y��4�a�$3
f9�)4��E95������n㉽�BC}B��2��q��M��1�n/��g�6�������]��t�c�g�$�L/>
��Gˆg�I�TPy@�7}U��g/�Qc<C�3ks�˝s,`��W�E]�����<�9����
�(w�}h�K���%�Ԅ�]I+EC����ޟ7�'I�=,�6<w�� 5��!tگIMUt����;J�#��&b��/��?���i�����'1�}`ʱ��áGaA�z[��@�F"?�k�����N/�M�ѧT>n7����P���$���v4�J�U�3���Z���x��`;�LHqK*X8�������ʣ��Y���	^�fD�%1���ރ.E.�/ņ�ӵ���XP"-Ѕ��-8.�P��:i���(�/�ծ��,S�������=2��^`l����|D���KDWe��~���U�L\����S�@1u�ua��ܭ��0�)�kY��jR$M(Cz%��ҫ��[Q9��]�:�����iAG�In*N�t�̛#����[��y��cC>{=�7�I��?�q)́��.+䱮h�Gm��)i�Պ�m幽9�K���N�*���u��@rn�pu���̚�c����9�j�{Dw��=�������P��*��lM��6"3�IG��� �jjs� �{H��{#Fi�����&��ƭ��v'F�۾�	@�i=rG�dW3����!~+�ig3.�ҁ�Y�V$-��R_����	'Toxc�a��Cwn�ȳ|��z:�DY�mn�N�0����Z��i��E�3̯�2Q-������zVK��]W��M�I9,fv���d-a�:��Oo��gެ�[-?�+gf��1@'���H��;N�}I�����:����b��׫�F'G	�1b,�hQ;e��*w�T��j��k`"��B�f�LBu �\�al�+]J7�S�5R�Q��0!�(��ڪ�n��,���Ex�#�YVK�� Uc��Е���E�5��@]������j��C!Q&��:1u7�Z��z-�c&���AKφ*A�ɓ)�G��aN߫�մ���N�c�[���}�^��e�i?�겙q�t\������ʾ@d;3�)z`�}k�� ~ '���kcW��H�#�%^( C[�_
�ƞj��Z�xgs��v<m�����у�����Ǯ�0����W	5�Q=B*Z�8qrb�g`��n$�~�a��w�YT�5�gW�n��Ǵ��_p��c1���~dF+U���8��ed�i!hl4C.��=EA=߻Z�$����j�wp�f��1�(�FF����/�q"7C�N)�cC����5Y�zI�{����|�g�UI���Tџ�k�&D}�I�nƶ�D��G�2q#�A�p[�p):����PM�^����a�_ʶ�l��goQr�$%EX#�w�3YfY���]hv
���@j$���
#�̙�,��%��f��KF��քP��|\�[YVc<�3n]5'(���.����]/7Ў-+��j�2x����p����8&�y�gf	7�����#/�v��,��dO���� <����J�Bz(���u�ao�<e8K�w�Bs��f��~Qc煹q߀;�QP���S�k�����s���.��.�{�2�L)-$���>v�dB!��&cN�����M�(�b�#�9�Y�BvvH}�M����Ȗ��l� ���9���"�eq��˔,�;�*��n[G�3���:�}L��l/�*�1`ބ�?#��s�(��a��w\`�����Bv�����ϣvy�0�&�K�M���q�����dK�a[����E�Y��}'���*��,�7w���L��+�{=����U��&��{̂���q䑘���a47R�rq���j��9 wU��ꫀU_Ҥ��������*�q�b:z�QrM"l@�6�Y��^m�����1ZI(�B�U]�Zҟ��g�o��X����������(��)����XI��J��z
���nF�H4K�m�N����$/�%r���ӛ�%aG,T�
,~:v	�3��ϒG��~;�-��ir���n�/h0�y2��F�D��~�wm����o0;�5t6�=V����������V{�^/_k���	�i��#�c�*~D����"�	ؙ���x۶{����C��@���Ϋ�͏8��2"zG���j�ӓr����)��� #%/B��l;a#�8#�c��M�:�=@ �_:�
bP��1�[9����&M���ߌ7���>u?�d�O���O��K���8�C�lvv}�%����Jϲ�3���/��V9!m;��,�t��Us5�5Ov�3\�1v@�\�p.�7Nǫ:�d��,�����%�G@.��,d��s�=mV�Q����%|nvAPn`������<�݂�3?�|v�oWb�*�ӳϏ�~��ul�<Peq��8F�����`(QC]u�Yl�9~�� �!M�<��؟�\�q��?�݆Yx}�}�T��`I
n�-�B}īLV0[����q6>5�8�f����1�>V.B7�O�S��G�dSX,��
>����.��Π���?�(�B�١��z��~c���T����������N�p�Ye;H���d��C�Gۀ�j��IL	�MS���n;4۝�m!d16�����n�Oc��%���"�`�s|Xq*/(��2��7������)��'NQ/�� �;?��I��s��D��Թ�"��l�Nq�WI�-&��}t�mI;f<3x8�ݓ���)|O*�M���J}��n��!�{n/�:Q&<ň�A���|�TI�k[\;��B��7���ρ�ncy8��#�V�h+�H�t�'��=)�����kҢb|�|ˌ���Ÿb,2�f�Î�����S]�O��Sy/�#�~P
4�.����n��ux�It�@S{<�[6ʿ�~�����ڷ�5�]?�зؤGv�����*vH��8q���_k�xJ?C����W�b�e���F��x�eHt*���Y�+�ƻJ��V��	�X��Eg�����Nh��h�|�� b�\_�G|�b�;;��sA����[CL�Bq ��Y�Q�F[UW�c����)��:��rA9�Aqy�=�1�8��.|P�Hf��/S�O�ywà�Ӻs�c�8KJ}�K�w��_+�=� ���G1ἑ]>�� ]�9�8�Zo��Pw8�M�d//�]��|>w�}pV!���n%�)�*����0�/����߲N����S"��?6Ԅ�&�uw�f&q��Mɭi�a������z:=�V���f�~�ۯ̒8`/\��EB��T;�f%�g}�oO�k��?_����,�R�e} gv�*<{Ԅ�݋�s(ZP3���;�5�7����-�~��*��U@c1�+y�u�m;�ބI����"bWR���[�7J�"+�0	��s�蔃9��
mv�ڇ�� �$vM�y�����N�����y#�rDˎE�퉼Ij~�J�:C8E�� �g�Ʉ�b8Czg�8�2������][�O�!��yt���m�k�܃[ɇ��_�N�g�h�H��uG5�RX߾���bZ�ѭW-�"��DR�H��ڏB�ժ<<Ĺh��Aڪf���r�8\�\�y��E�X������C��H5!F��A��Q�Zݳ4WM[|D�]|ϡ��sP�S^i�Dl�t'���;<G]lk�&*(XET�<�7I:*����v��\&yO�v�e��n}u�u˾�����͖��rc Nl<�w�]���<�4h+�bm�b?4U7̳&7�7w�8��R��O5���R�Y�]�3`����!�H�]�N��
�����LZE� ��@���Cpg��7䚗����GmnNo�����-��Fdo�XQA���|C"�m�"5�Ԓ|�r^���F��#U�M(+��f^����c���q�����#��"�#Ga����f�7*p؊]�&_Y2A�&뺃#�S�1sXd��`��J��f�����h�L��'�}G��Q��%'q��(C��4��rz?�gM�@�|%vB�{�#U\��\7��\���Yb�yX0Z8�N�ωA�tB��M[FA�L����Z����HAj �n	��Q������� 5|���\6��Gh&���� �$�S�2f�q��^L~�z5H\�q[Z(��[�x�ʒ>R��{�n�^�G)��톓x��مoq���M37w�X�?�v��K3��~���'�P��쾌���E���`�N����^��P�7�����ؙ��6@�aR�~К�)�C`U��IYƛC��˅���b���N���d��mo9Y�G(�X�Ǜ�����{�1x>�"A&'���)�ؤ�����[�}��,�Ȋ��aI�S-I4D���Pk�z-T��F1=�}(��6Q�mo�;ȁ|ܻu��Jq3�a��G$ꔤ�ي�Ős�L�շȗ���і��O��d�Y^�,�1Ump*@�*�@ǅ,�]ZQ��`&����$��N�k�j��3x�nu�S�����r�A��,��H�y��s�)*.i�[F0ۧ�H��@�\N*.��k u#\uܦ0�����RB�w2�� ii+����w	�C�q��o���!����R�%���pdh�sA)��@���{�Ig���g�(��Y�o,6�*)��W�*lW��ru�1�sZf'�;��'���:��=���e�|��d�<�[�3�@/��K�+=8&i(�J[�[U�#����R6�� ��E~A*�}�/�k�~G�"%�Ϝ%��Z���/W�:��)���*�p��8M+�A��=+�%2��d�g���֚�v��[>�ě�U_e��ضKfv���G���m� o��"1�EU���eW��g]_"�9d��ۺ��RS4UqI��j��j%�l.4�6c,[�T��V=p����� �#����UUv^�Wq|M$�&@Ѵ	�ed��s���Q �����,(���Έڷv�����GB�� ����2�_W�Ţnt|��4o��F��X�"@n��l"B{�z	�d��Co�H�/1�&�9��u��Ŗ���GS�kw�h�>��FL鏁���H5�f���Co�~��q<<�UJ�1�=Ko��-e<}&���*�#����3).�"�J~;��4����z�i�=֛�s/�E���B�}1�9+��q���޻VqI��(�0b�=�����-[]C����t�Wt�$(WP�ȭ�����Jy@M�����?KaH�z�b:���ӝ�)�c }�:��48��v&�o��hFݵ�{��r��QlT�O^�v8_R��fDn$x� 91��r
��;)gZ��>��NWT4fU����Yi'�������#J����tL�/�`: n����]�����G�"��P �?�,bE���<�6�����K<)O��,gڟkN�Fq)�a�Q�/-o�+�jވ�`�fVy�=$l|rl���?G���KqS�5n�M$9e�:=�,B7�F��Lfg._9�4��j�(�F1QB��!I���,�����&q59��V��������DK�,I�D˪�j#����vB٘������s@����Xu���ur��u�c�w�3�d�����Ͱ�C\��k/X��m~�C*p;W��~*jQ�?�.r@�����PD�&rf��.��E�15jx ^��ټ�':�U}�&�]�>ۭ�9&r��o\=�b��� p[J��=�{�]8B��$���p�j�n�/�5�B*{F��7��8�!k9�Q/kh�bș*�RJ��ˌ,�?���]Z@�К�jl�q ��*���F��rk�H>a�[d#�]�͘��I�����~4��っa�V���҇$�n	Iv��(�i#��D�{K�]OV�{�J�ɂ*_p���WiK�t󮵒R�b!��ñMվ������FȞ����q���I�?�Λ�<���Ba�P~+Y�Y�.�����q�CRc��_i7e(-x�D��G�TН�� �(��2-c}��M� �b�S���`���|�A7��Û$`ɒ<h�a27(�* Mr�+1�8�(��D�e�o9�٭�- A8}ecnO����_�6̯p,��ꀎhC?��Y�a�s�N��[���Oh)^k�"�x�؛��=-8��D�&ͥ!�&5����"������w�<
LIVOk�O��е��G��}�29�:Bg��D)N��F�*D5�6Th4Z�no&�h���@Ek��Q��YK�V%J�4]���/z�/j?|�
�<پ~/��A>� �M���
�N��m�ٮP�u�{%�S���P^Vk��m�����#`ƹ��Gl��cy
��9#c3�%M�yb���Z��bq9U��O����&��i�A�zu���a���P�<�`�Oz
���x�U��iE�t���P)���TJ����N�3�%}����r����]��Q��𱽔�5�ˁ�VEKK��`J�7�=���y���a�;Պ奍NXƃEr����h�m��SĽ�����a4s㓍�!��al��i�6������?��s�=�1A�<���	eb<j|�e�Kw��=��6{�#��M�{کjR��h���9�I�^M����je,���Y/沚 �9�`�����cg�q@Ӳ2ɢ���l"H8��ݗ0�I���&���Ϗ(n��(��FkͳI�r2�C!Z7���}�Rqq���+�7#�a�a ^�TV6|=(c���M@5�����$E;ϟ�B�ݬ���Fnp��)�2J��	
�~��4�ĥU��53'��?k�ֳ�d��{f|��u�
�
�4����� �9�:I6T�K�Ы��c������`i��0��8���;�T��K�Hv�G�_�͸h��8���x�}\Ҩ�g���olލ��x�7)?`j�D���~?�.`&TߡJ�Q�hu��l;�PY��P��xx�s���������B��勀ܡ���J2��?@���u���;��vJ�Q�,ln��i0���P��~T�3�����}-Av�.������$��±�|�G�?���8���	+�v�Pa��̭�A�h�U���*۶\�fDME�-u��U�7U�I3�Iz�|��7��X'm�ETIM��J�9KjȓdM`���8��s�v���]p��g�\��^BQ���>��8�9�Rv�+LY*�� �ͺ�NE��D/A��ƹ���r�A��
�0�����V��&���@u�=���2r����Ч)B�V ��T����(���2���Z��!�h��Fsۇ9vWY|Uމ��40�.�;�W`��KX	j׫.B6��@A~�}��A��|����W���'�ͺ��a�����.ЪZE�m�awA�B%ŉ%f��|~��8��Z!�\�-��z�h�oX�.	Q�w�0=G�4���'t��լ���C�Ej!���d��D�y9Dg���~��~��1����!�zF�_�Պ�O���q[��0�篴�(����:� s8>co:�.J*i�0ԫ�{�}�\��'_(�v��-��%W�(3����6�S���T��)�e�Ql�V6tR=�aⰬ���s@x��5�y����@��I��@wUps��%�r�D���WkK�C�$9�i �Υ��SYE�X�}!��϶���r̀ A�;�H�<- O�P���v���ȥ�̏8颗UҤ���z��ZnBA���J����y����~�F���N��F颒�CURP�3;i,��?���B2�Y,���oП���bZHF�'�F�|���+Y)�7�;��x�Ue]�������_8	�w-���,&f�ؚ7���+���GD�:u��N_߷�0bʸLw��DK���c�H -���}c=&h���{q��Dd�I�Kz�n�`T<+ۮ��nn)^�^�$�y��0�bP0�BB�*.I#YV)�
��:9ʼ�/���v��T/<�'�!��@x$C��L	,��Ώ�:M0:y���~t�Q�⯀�bu0Um��8�t(��Z�����3����)T?�~����q��x�oFoz���u���xm�?�� j"��f����h�#rǷ��Qz9�-��k�Y3���-䳡�r�,!�j� t�y�=�6$����Kˮ���Z�'z*~��b���x��u^�0�["8f���S�w��'1�m����g��2�,� ���Fdʃ-�.��޺�n3μ��˱�*�;��$j�l.��LNo`���q��Enr�i/�?��*J�W~��E6eB��A���63�kt�F�ak_���tf����.k%��~]mj��
+�(6��t���e������B���9��ݮw��٧u��)��пk�*J�����M�V)�=li�{��B�[5I�'����,���C,���2�%��Q<�(����>��o�x��4�xZ[��������3�ؖZ��:T��o���^������'���;/Ӯ�S�;�rn	EKVK�k '3��}�2�߈��b��.}�P	x8%��t�ia��̦s7���yz���xN4!�9@ȿ����\]=��,sb3�0ği�P����L�"����W1�-���r�"���Hd��Nn)r��"�MQ��~u7�ÑI`���WU����6�?�;vf|�H�"*/Ć8yi|��U��G��fEܘyzl��j1Ð�iʰ�bl��&���uU-#Tp���ra�f4;wEV��ܾo*�mY���z8Nf*�����g��+�~���ͪ�T��@j�u�O����o��1�O�: J9���#��	��$[E�/?��_)�|[s{n:��En����
M����o$\\�;9����.��� $�ɿ@1���}^��|�V�&�3ۃ1Stkr������#��מ�V���H��>�}��"l��#��'YhTu7�$�]�����;�	�G�ό�Doܹ�aN��X��Ѽ��N���Z�|��2�H�g��w ������b-�s�#���q��oK7��g���v��ڰp���J�y��']�`��tO;D숄�\�x�yH�݈n ��i��s�4P��!���%6ݞ(T��L�~aJF+���3w�I#bk~)�n��kc/��*�	���w��N&Tpm�)��=ӧi1�K��9�.#�ޟe���p���&s;́����B�
����ʆO(Oh�C��AKY�{�tu�*�y��з��^�84� �f4x�B8|�|��֏^C������;F���2d�R(�
&�9l�7��l2��,cq���;��9��K�e?>j����F���-?���_H�%�_�1l�&�.fv�81��ש��K//�]�R.H;�/xx�e�05�ʺ�-�톡{����m�n�1�mU<,��2V�Zֵp�R��5��Y6�T����b;�|u�,�7�?V�Wu���<�X�I����+����nwqF�}�����N�r)�T4��F��p�x��ǎB��؋�W�K~E���/ )nT��59�:����$�מ���Ov��S'��J�DV�BМ,0h���:
��U҆:I��*�+���lr��Q�=�n�w ^���T�v�v��Zy8+A)�B�L�<B��\.�8�p�!!^���wE��)@�.O�������Zy�U)� �S��d�-Ϊ>2�a(��Z
s�z``�VG%�h��E߉�Ҡr�=.�'�g#R;���b= F��z~\F��w>m����b�v����S�E�l�C�h�����k�h�q��w!N������[���ZkN�]63G-�E��y��l����TP������k
�޿���q�����=� �>0\�-�m*�Q����u�[e�7h�T����sʅ��a���ڽԲ}�u���[�8���(�c�����JF�s%��
`  �2YW({3S��#�6\Lw���)Hlk����!��S[]wP�c���;G����=]ʽo�0o�]mօ�bxݐX����s���]3����Wn��-1���g��X���!ȴ��A6��*��ׇޜ�Tڀ��{	�Y���N�c-��Fw�0/h�?d������y�d��/���x�;Wc�3^�2q���4G��5�ɾ������T���Y��3A�ib| ��A��Pp�H��!�n���"%*k��4��Y;�Ղw�q�4U8H�t�{�Ix7M<�q��%#�ۯ\�t`��ej�������ئCb� V�w�q(mi䭚��H����������d�����ü��G�w�LG2剽�e�ƅ;]��-������.E��\T��2-9�&%א�)-��6��-�{L����j���O���2�Y�}��<����$��@�X�R�A�?�bx4��Z��Jq���O�v�R�:���-i�߆����u����Ð��>y��a�6RQ!@�0�\���ķ�i3䃡�>�t�Z�N���PŘqB����;�BK6�D���뮕;Eа�wIW�"��؊Fap���y|�˴�I�X�F��48�&�,��o&P<bnA������Sg���C#�[��Z42�����,��������ts5D�V?}�
�^����|�;��+BW`P��]4[^_:�4��)���j�a
]�>T�I��3�����ૢS�
� X��y(;Jc\��Iq��j�(�f��w�XsB
�'�Fj`B`s��.��&�<>9��7X��zB�o2g�-?���4ȥ<���Yi,@��O���1�V���K��t
�zX̴�ո��K�&�<x�ܘ,�c���w����N3����[��t�k�ЛW��8�iG�7����P�������Ӯ��JFΪ�����mZ,��H�Ó����m:��� 0������j����l`B�������V/D�虒���H�k��f�@�K�a&t9����V2^����rv�G�"�q?F�pL�ݢ+V,m`,r�*Q0���7�5���ݴ���X�$=dK�n�������Li<�Jm�+�-v# ׃����Ô�;��mh���J��	$OR�\�I"����<�l����}��DI�����]E��ő�p:�yԔ�����"5���#E��ʛg���8���/,���x3y-��E˨�K�wf2i�=�s �@�*o��.�Yg��,e���Ӑ�
�~�T�$ /Mꄯ��=\��T|s}��E���ov���q����
L.��W9��ĀԨ �ʧ晆-:Ha�}��3��_���b6E�~?b�T��*fg�H���(�o�;(��2La�ou�]z��Z��o��ۑ¸��x�����f�?w��3{��֯/�p�]ܳ�9E�R]�5�:�#}ѩ��h�dn�k�Q�q��/O�/�����VI�i�1��E��؏yZ��B4� I��/�*�l]� 饗IM�K�f/t� *G`7ԕ���`���ѭ1閂�|B>v���7d�!�e	y����3L{E2 `�Og��j�����-W8�qZ���I����Lq�2X(�s���O�'���B���"b���l�P�ܮ��YA���!O4b6C�u��tƏk�3�4!q>@ݸ�5.����B�N@�gY�"v�_hbܸ7� �N��璩��4o֐��@�e��^g�>X�ا����<s
f� �s �-�l�qe^K��=7�6��ǀ���*��~�4R�.�D��g3b�F��D*�]�B뜁o��ݻ�l2� ��p�H�h������n�w�*���<��'u�O�n��ʘA3��)�^��|N� 6g���|��	�l��I\U��Xܼ}������;-A��HE8�Vov��x'�-Qm��Yܟ󢤿�G����,(�S'���AQNk�.\�x;	��S6*���N�TJj ��/��o��<��X�q�u�2r]v{�������hi|^_Y�q`7��$cd1`2|��}]�[�巢w�<���r��bu9�Bh���&[��y�0�35J<� ����ktA	�����$"Q=�;+b�ĥ�L���"C@J{tǝ{xy�pI�ɷ�JX�S�4^󖓅�-�r��H׻���4�!�\j��u~��E
��iA��*��9dr#��.
h<ȏ����1�Ǫ�{ �_�3k��ś9~�_�e����"E��u�]���n��'5�=`�K���H=_��[@i�R���y��`݊^��*�ӃIg'�|)�0�P]|��~�D�)�?0��q��E;��F$g���R��q�#�?�}��h;���Bܢ��u�Ӣ+��s`~��b�N �1G��B�ɋ���'x��:�2�'h�����xiM4�坳]:�7z�>6�#{�E�Q�U>�r&��+r����|������&������s��)f�mK����GzOY	^�j���_�"���D-�IÊ�:6ãixx�R)������U�_�7Cl0�+����I	��Z�Go %f݁���ڃ䔗�߮܀���=_��0#)�Yƽ�&�1j`�z�lN�t6ng���=�8��E�w����6Ib[���\w�r�e�ɰ&o%6�.`��I��4�>�nȒ�F���$�)C�⃬�a
'�L�ێ�1t���mJ���pef��ppH�2=�g!0WnlJY�1�s�2R�MI!��v���X�����eS8��,w@='��X�ǻ��Xв���Z�[��	$��O6ك��0�I|� x���Ж-V�3�{f{�fPº_�Y�pi۫��"��ܕ��� �O&��8��<�RCs���Ӛ���+���4��g>>>V��8±#nSz����$��-�?�eE绯?mD�iV�)^Ui�hߑx\���䕄��,zc>bhP�>��KB��zkP��_�7�|+��6c)��/D�>P�S!Gʃ� j�3���0ף
����x �"���Bb%�d-��̽d你T�]:K�ʃ�\�@�J=a�#a�`����QNd�ұ���d�i����a9��9[�6v��
��TN�/�9i
������ :���o�m{z��n%Ql2����f�r�r�*�i�M�[$uI��"�=��:"ٌ����Pʤ+��Y��DfM�_�Dμ�z��S�+<��/B/��	�J<2j՗*h���ݹ~S,ć��NZ��+��	2+��  P�8�ٺ\;�v�
,=��_��Ym/;?�+ǫ,׊���\�����Cn��¾-7جE�h�/���7�(:��[K-ܔ3���6���C�׸H���Q���VUW�ހn�Oc����;]z�#,��C��Kci�Z)H���h�Rgע�7��+���{�=�b��j|"}���b�[��3/.8Tt�����E��Z���:؋�GZ4��}���8#d�'�ƤHn���U>,g�'w��x��$�E�*�]h���G�����ŵ�6P"@�҅�nx_k���rh�z�i�jE�-�D1ZFO��%���On�2��YЧ�Z��h�	���H��=a�m�|�0�� ��j�Z������X���禎dk! Vy`ϙg�ԬZHe	�.�V$�&ɋ�
39U؉1h̊�2�2�C���y5)�Äׯ�aҺ=�[#�z�s�S����V�{,Uvw;m|z��mQ9�:;l��	ьZ����a`#%T�ؠE��
BGt�ή\�\����X���֜%O��w�>����b8��?B||^P_]�m�%i��@^g���b	PB��`������,�R�����H��^z;���P��S��-�4b�uǃK�)����.Fʣ$+	����cp�1���\JА��bs� �4�x���y��j�_��u�/Y �:����\�]WG6���a�<����	����m�Dz�_5�j�OX���������ب�X��~P�OP���n�x�M?�OVB����>q�rV>�hqI,[���b��Q�;�	����\��N������G�04��p5�&�~��:8�a�����f�Su?ӇaU�(��P��곣Ǽ^���I���j*&��`��w��.Az��a�vW�f&w�{�\�3">��7P��꼓p?P�9�"Zx:h&���
B���c<�>O�b���:RC� �<�����İ�(L'��W�O"��pA�����/��[N�\��w.������)��xJ@��
0���k���i�`Ü5��h�^�+�x.A�`��t�H��mz�Ey��{�G��g lٳ�2�9���3�8
�~��G��	��#;�R�p���;�ޏ̎��м��YE�GߴT��	T�=xW�����')��v~ٶP,�5je�9w�ܭ��6,;���H�[���L��a�!�?N�)!�`:��e��}��Qצx��¾��k�7t�o����!H�cw�W@u����H�����T��;�}���u}"�a۴�#P�'���G�� ��^BV��P��j�F���[g����)<I��Z٠G'��0�,8xѽ Dn�( �@n"\��A�tM���W��=א����n\��� _� �����<.ӊ�ï�p�y��',h6�P���c7���a�uR��p1���H
4��n�Q�	��o?�Z��/�]s;�e�!���x���ZG�4�sHr���3%'K�s�g�;�϶A|��8�ǟ/��	�j.-<��V}�����w���vɓ/�
��%ֆ�[�yj��`pBSF%��^��["���u�ш���3��zaL�'��X�����@l�骺PJ���uǭq�aE4t��rv��@�~�:v���T�#�5}��^��mF<t�M�+�
�-8�ˊ�@��z>r}����&���h���$�]���]^�	�4�j��)T�=�ӛVW�|\��A_�y]~��%���69��F�!��Ú>�b���Q�`�V,+yr�����;F-�Fu��mX�͝'�s�4�_���rk؇r��З�A�, ��1�q�Vd��0@�f��%5,Ͱ����<xcBc����.�u�hD]b�*�Bo��z�<��P6��[�%�� ��?���:W�Lh��
9���`)[���BcV,��g ?̺�L�K���R^	��3���u,���k��Y��Y8I�8vO�u�d��ٟ��FɄ��Y�/�t���Y�;i�U4m�U�М>ɩ�w���V8O#�����vHӂq�.����BF�p� ��9#���gz�u��uFA�A����g@�b�E�ȷ�/\hG�P��l�C��b���7�*6/i=@�LQ���E֖����E����w�v�L�{.�Qe_n��C�Pc����p�aJMl����:7��Ƭ Vj޸����O4��ac�i3-,��SX�-p�b��윤{С�:D�Z)��0/c��<���}�hb�{$/����I��|B�/:0�u�*5�>��5��Ta�F`�%�� ���{vU��X��	���J����S��
:���������؈�a��UG��n�����}!�� &Y�%R�i-]T���#�h_h,��=���&=b@����e�YE	�"�@�����04&�g�sN���7��bt����|-�A0��R��8d�G�r���'�J{~ �~������������؊���ڳ�G��FuK0��4e��%(�M׍<h��q@�k�}�&/�҄�\����I��d�$��.h�&����1t6o��5?��ɒ�S��n� w���0�,�i�v~#[-*{~�������8���R������{�gP��S*�C�q��Y�UM�T+��T�6�>ۀh�-�Y^uG]�L8����{�=*H���p�ޡnM��l�az�i*P�4��1����q�v��B�"DTJ�0Q̡��������]w�J {� 4���hӎ�I�}c:,˅V��&���LzO������
}�%�*VC���ûIV Ѕ	�C3����о�&U=P�R�h�!Q��.��X�v�m!nX�M�{Y� �#k�*���͡1�H5b��綠��!?��3"YpJ$Qq��b�8�g�o#o�#����~���m] ��_���΄��2���ߵU�-1X�����S9B��5������Q�x�$��K̤��),Z��@��S��TE� ˇK��2Z>��^H�q2v����pG����բ����tp�W�&�FGL^�t�]a"���D�����^���+�j�1T�i@����X�k��u����|�L&�cK���,������4��ǰ�X*�M���*���KV���t�x���b:>�Jz
�8m�_!�!�SO��$Q6�|�y����5�]3͈�����������+��D�i9j�wR��=g������$t�����̙6�m�5�A��8��Z��E�t��'�B\�H/��(�
�A0��<Rn�=LR�*d�	��U= όz��u�ۥ��SgqQu߶P�^1�BD��oۤ�.�d���\*��9�W[j��\�[hjg��L��U�j�j��� /r��B"I�����O�Ay�o%ʩZ��t�ۋ���3��p��#�>5�Pn�Č+�%���+b�T��W�5��Y֙�3�L��K��^8�P��
2�0���_}r	g�#���G *E������O5K6�:�y�_v'���_�Imh��������&�h������?��Ρ�Dz[h�o�+�p�ꨡa��4�T!3�E<�y�f8�N���ȹt�}p��F�5H-���`1se6�}���T�ZS[���N���tQ�ʄ����&���Vۓw9��l+��ޭafք@�>��WϨ����Z�8fm���#]+ ���x�}�s�l筣Y�ߍKBЍ	k���A|-�4�����$�'Ŵ
2�TJe X�1�7��Ia
���Ș���|̡�:Ewl�L����<"��
�~�b��V�最�)���cS��S$VCY�Gt��y^k�f.BȹuYX��k|L���Ǆ�s�/�3��F�_2ߪ�y7�8��i�����@��@��,n�rux=�ؙ�a�m���͌U�B�-E�̈́L
��Nђ0��u�8M�|�8��:��|"�%s��$���I��w�G�����^AbPIN:���<#J��ԥ��B׈�p���
b�&e�.���Q�By�$=B���p�X2X F�TJs���F�[���@�6ш�3cqW�ެ��$WFF��y�a��=8��%����z�-������a�p5$�%⮙zxH"W,G�1T_R��C�d���ywV�C"Q1�������aͫN�;N��`��ce�x��l�Tn9���أ�#nA���$��`s���A��-���4�;�#��E�>�"	*
�p���2���7���d��wH����jiUY�����,� �G��c�B"��:h�{OB��vr�@�Ƙ��9����5�1[j�-F7z��5M�?2Z��r�M��~v��R8<�$�#+]�*���NQ�8<_��.��ߎN��~�O<7k!~�6��m�N,F`u�s)��[��ON���%�Ŝ�$�j���j&9���|:�D��#sWG���ٽ������!�/�ϵ'+��J静ޫiY��?���hd����+0�S�F�"Nz�ђ�w��9�2���t0���\�GE:�$�*D(k��/����Ƴ��L���t��'nQ`�+.ɦ�L���$̘�#�3Ժ������2�<Z����#(�����aS������*�H�����V'���36X�7ˑ%ع�j
�rcke 밟��d���	���b��ͦ.�&��Ŀw��4�o�ݕ�a��c���+�}���:<_������k�a��d�l#R���5�iTxҾ$Jm?\�嗷�B���)�� �,��?�/�shL���s�G躓(��@��JH7���O�Ѝ�>A�q{�7!��CL�n�	UU��N�*�8���ogŧ*C����̄��}&Rx���i�9��i$�Y�b�Q��: Q1�$�S�92��И-&�L�f�Z�Y=��a#�6�VP�n�%�M ��ЬB/!ni��7K�:�s�j�g�� �g.�9�{V�B,+s����;Ĕ!�b_���9%^K���2DDоִN�6`���ÍnO�4�"f�3��5u4Cm�F�)C:�VC0ŶSם������:\h�Y]Tf��H�-KK�R��_c(~+'v��NL��x�oC����ܰ~zb�9��ՙԳ4�����u���׊^0�BCf���
���.#�1"TK�/��[9
��dQf��vV7�]jۅ�l�~��s�,(����_->�1�ge6m�9 [H��4Vdh�N���K�Za���l�衊]��>�Y���w���q/:=S���|��k8t?�c�6���7�ro3�1h�αw{�(�� b�S팸e=�.����sl�>�0�Q���a�M6����JE49�o�S����o��r�I�I���^��RF�c�c�WV~$���S����mZ�"�O�/�6ᬨ����:�.�r=D��'�=W��'�z�&���_��ʜ
�����-[���K�(�s-8&r����i���!��?$敪�*]}~�o�jc>9�ZaX�����'�Z��J[G&L��r��S��b?
_I�l�����N@_�uܩ�
4�K0��*zN���d�.Y:G��ï+~|�/u�%m�J����c�n�^��Ƥ�s�����������=�#�L?��|D����j~�̬dN��6]�sY�3�����m�cw��*'�ͼD.�xΌ!��oh]ZI����m�F�!9��`���UP�b�)S���}��f���g��Dy o'��5��r�Q�v��`�h�:��+arڭ~k�q�ygAR�NH�"sN�2g_��
w���[��c��,�˫����$�G���N����V��?Z_�UHȼ1@iis>�|�i&�:i�V�˰l�#|�'~�
���m�?%��,��CgzX���=�d�'��8�i��������Uh�*���JUʫ�d�?d��2x���T���w\d�y7[�`�ڗ5C"/;3C�4r�P��wg:�j��j�K\�T��X]��yOsJX��T�0��zu��)e+���a���x]"x���
a�e����4f#������˼[_����ɇN�e��B��T������B����C�ri�UnV4�5$��at�`D�f��Φ�o�#ڥ|� P�!Vy'_����_%���x]p$�*}@�*��d�&X:�a%M���fi�tq��h�?+vD��*
J8����8#>�Q+40��<�{JM
�{�3�-b>�&E�_�;��}��XgM��^,I^̟�ӈ~Lgg���Ż/J�<���3�� 𮵒�"��:so���vSV�"o��$�K��%51H��.�����Z��������֍�q%�.��ۃ��cBG_�dYX%�h�:������A��R1�$F�*~�����:Va�t!N�Z�eC:�jػx��1K��J��$��9��=	�٤P�T�̳2�4�����㢤j����gV꧱v���:��o�EP'QiF��#�u=Z�^�3�Ңy]���xx�O]���#����,g��|��{�95`�h���{Ll��*�K���Vo��0��jr�B8�$���F|ߦ���yVb���q��}��-)EJ?�]n,����ǽ3�3���0|q��Eq���͟�g*�ߑ��J��8�Z T�>���DX��x�#��E�b��'r4@����.��6���a��>��Ïť�O���[��3y_3�S��m@���O����[�ǿ�q{� �����ID8��^�ǁ��R6P��8����X��"��N�8`�8��!�gV�:QϮu7�8�g<���n���w������(Ч_�j���T|� &�mk,f�E���I�1��=b],���@�'!7�U�8	�ܗF�"A)蔓�����&,kZ��|�Y-�/�j��	6K��e	���!z6Q�>�m���� �X����~�rC���������8�Q�����I� ?�΃ F��?>!jEx�kI�-dͧ9��!����ofι��); r���ܒ9��6�)s������Ć�a�W�2/�Rw���.�]�o�"�UΨm�lg��Mopƾ;� H�E W�Q����)u9c[Ѿdَ>����1��|X>%���_��UF�a�x�
z�`��
U�?A�<�9�Բ�:ݥ�nT��O!��%�\�W$6*�%4�l�5����9d g3�Ԋ�C��
��[�P�� �f]��]~���4�A�+��GI��V��{hĿ�ՙM�0g�I�{��Q�	$[�G\Dʢ8r�d�Z\\u02At�1����k�yl?�A۠�����:�����{�sk�ë��QZ�Y�o�r�#Y1s�&2����u��t�Q	+J�)ae���tK��0R��PyC������2d��:K$πҾ����ՠ���{�?J��j"glkA������@���"%]Lh�i��j��D��@\��]��N�����0ҁW-�T�6����~�;��Mx�լ�o�\�}K:�Mꖪ6��,���!��`�7Dw�Dπ��I;��J�%��Vؕ���F�MhTXC ��U2�ںՂ��X�u���9��T۬�z����P��V�Y�Cu%e�.�_{[o�d\PVͯ�F+�TE�A���-bW:'B�	}�L����B���R�����ˠ�̟��ç�U7�4 �V�L�U �Y�`?|X��Ӫ�-Ƹ��S�w�q0��ym/I���!�}z;�sH ���w�@,~���� E-�?/��Qhr�.3j��C��e��d�m������= ��fZ�4e#�Lr���I[^�"�	����ۉ=�BM�	0��0)%7�qS�C��p}|&u7���'��A-�F����FV��r�f9�ё�
�@85�G"��^��{s�A7���m�����	��`���@�m���AJyV5��5� ��F�`�|�)~WE�N��ׁp�ƖIg�Q*`Lu,=?-S�Qc��+vT�0&V����EB�L���"�DĖt�_�� ��i��J���i�GR�?CS��? n��F����cT�uc������Qr��D�����N�0���{��[�:D5��	oN5In9K�ۇ΃�LOWOs��j���:�O0��!�� X]�:C�g�.,�mT���=� ����r��q���E'��VC];4��JU#��ta �LE���23�lo��K�B��h� 	�#=�wy�-b'�F����>7]뱶��B���wuǬ�J�����t�jE=9>��&q�R�����	#
b1�b@yfG5h��	���Ľ fNB#��.����n�ji��%�z��{�M��Ձ�0��Cğ�9�=1@����Xj�P�*�?����#(!}2s���["�,?�&�L<0�Q���a�	Z��q��]P%�蠛4(��5Bl��娪J[ԉX�E�N���a�h=1̛�$y��E�k��� ��/�X@�  �9yi�t��;%D����EsE���&SB�LMe���Q�
�M 2`�1:��/	��B���.k��b�@���h��!Q�A�c`�`s��3�Y�R(|t,B���V4]ڕ�}�^+k��i7�? ǉ��,	T�q`xY橯�&A��� �����KW����D3(��3+��l�Ey���u7E@Ι9(�x�vێ�l��G�l���+4�����0��ط��C��}5�Ӻ䔻5��/u�WA�Z�����7�Y�'I�u>�Z��[(��&m��K�U��&��{,(7¼�&�"xu~,�#o�v�>f���z�f����'�k�P�Z^�TG=���MkBd�)�����%�B���t���D�Ӗ�{���0j�:�B�N_�2M��-�������e���B��&����!�H .�!G�H0��.哽,΅�1�V�(}:j���"��Y[A^e0��Q* �20.��͛>H,���^N|���M�2�Ҵ>��ys��z�"q��?.�©PV���@o�^�fw��K���x������~ӥ�i�Q� 1ȣ]�5��r� N*�c���q�7�+�q&�b-��N�~ ���K8�{��;������'����|�f<0��_cQo�(e���-�ׁ6��欕=��՘P��T��>~����l��Ɋ4�D�n�/�|!�����/�Kw���5Mg�a�l�|Ro�D6\ި�+��'�K7'���j{�����g��~��H����/k�w(cr�\��R�ڏ�Hd8Y%߲��?�q�6e�85JKD�X7e'�Hs���� �Z �#˹/�k�%)�]�'�d�έ�?��)�I.�ݵ,�ol��+�������D���t�f� ��ߙ���Q ְƟ���n/�8rG�@��<�� (dԺz�
e��v��]y���+98����D�ݛ�S(%�Z��ڥ�
�_�T	L�:y O�)n,�F�>փ���_WR�jm�Bd-V59��gY'M�`!���a��q���N���d��j��x~��f�P�w#wl�B��E	�ذ9Yw�'v}9�Y8 r��~�)��Tko�os����Ryq�i
 P����nAK�ڧnm;��C�]��!��Z��n^X㖉F(�W-S�b�j�Z�,nu�T�f�
��jL�1cW�>؄�5л�6����?�/���],�T>h#���%'޵q�2�r;�:���RO���e*!�m��^/4����"��9���$4��L��&:�3����%��S0Ƥ��L�`;�ʧ-k��;SR��c<G�
,hC�e"�'{j�A3�Mq܅'q�!�i0�9�;���N�Nci�Gp
�_��01��K:4)�����#�n%A!�(�����	Г��-��?��(ڦ����6 ��Bz��H~Mr.�����*����,}a���lB��.��	N�T���T���S��rϡx�xgn��Bo�2����c��*����m`����t8/['�ۏ�2��ǩ?���%��80��!�g,�5�n,U�
+u��@���.�`���n��Z�9/�¿�]��T��q�����^J0��F9��'Y>i��?�p��6�֢k쿟����>-U�����o_��E!�6WI�=�O�H�+�~��=壾�1�/�Nw$��7,��P�k�l���L�gw��)���n��[��0� �:�0��ؙ)!�P��WH�;Y�\;�,Y>�y�� �c`$��(J!��n�J��F�&U��k��m�����n�̐2�}�w�C�|T@q�
^emS��і�+����H�Ѽ�7�I�=3�U�J�3���W�8�Zѽ���?/���kH��i��_g�jw�ӛۊ� :d#�Ց`��8]x]���&��{A/Mq�ʣ�G�C^�ϭ��o�� ��@��(�%Ҫ~"L�%��Bi���}��{n!���>>��E����7�$� ^1p�lP�I���dt]0b�0g���a���Fh��i�R���4e�)<�ay0��mgg\-��bJ}7�0Aِ������b���~ֈ >�\����<K h��{�$T��Ȇ�B�2���b5gP<3˗��%�h�?^���O�
�fa	�k�Gl�頄\�#N\2r���F����]�g�EZy�q��JѮYd@��
{iB���4NJy��I���!��s�,�.����S6TԆ8L����_�`�ή��&q0p%�xּH�W���_G�~&�^ۥ�Ȯ�o��������R��]�.�n,��=V]#��ɥ���?)�ER�ь{�W�J@�l)�3�2^7��L��5����HY�ݱD�~���<z*c�����4���2��RPd�b�#C��ϭ��ό6���9�P��}=��n@o�l�	��w�pk;��L�.�xܪ	ª͝V&t���p�29Ċ�t��qk�6x����,*�%QCӉ.�4fw��͐6Յ��T�"�:�z:Q_d/j��E[����,���C{���s�#s�ˬt��_}�^�2)4y���3��d��� �i��/�DÑG�0��T�{y����:��Z���Kk<h��ύ�Bt<3�����,\d�	;9�\�xC�J2�ޚ�>p��~�qܭ�������%�sn��|qRB���`�ۊ�K����:QJi���G�dnga��Vd*[ ��
n<�������F��#��,Y�s�~xe!d��%[���^�g�EEmq�r�Ԣ��Lx�7=AEt�`�}��@�+)"�yko�N������-Cn�=D�pe��v��9],������ �?}�K�ӡ�W6�����W9�k�<���j��M���AJ�JV� ������r��9�ؕ�h�G��n½�U�9�e�%�����9A$4���cyV��-�QLZ�0#�>Rk�`�A�"b�Եc`N4�n.��]�L���_F�f�B�:y�1$��X�3+%��,�d�;R�T�(������hb%��4����J/�m,Q&����d�ߤB=G�|?�~�U��!���¶���Y���x�z��N��s֙Dk�͟���/�� "�q%�?+�D¬���T r3�����~Pޗh��ڝ9x����	#t��X��������=�������E�(_}�q\�?*���NΰJe�Y99Nu��!��ۮ�s⛽_��)x����D��g������dK;p����UQ޿��VZ
�5���@M����a �+%C�ٟo�*~bz8dxi4����烯�tH��	����J�]�ˡ��M��<�л�We5ڮ�H��Jn��{��3��$;i���lU���YU�t(ވs����8��>��-��d�"t���^�?���I��v�|����������N��^��y�Wݏ#��ِ��=�&_2�/�1�*��Q��Qkx��/�&��<%�8���I����U�L/�����Sݫ�R����%��P*���G��塏�GYvdl�An�;�g�O� /�#⫖�z������ҳ�Cڬ�t�>O��OF�|7<#�_8?1/w�G�WF^mѴ���]|J�c��D6{�4�_e$�5H��������8�(D�}�C<+H�j�i�mH�#d��a���#e�j�~�^%j�����*�b��^[���M��S����f�h����QL�l�I�J����Y��iOYP��E��*/��8gq�Vh�m���EF�톿ę%��><R'Ma�-W���7�<��&�{oSP����H^��c��M�/����2EOɂU�=)6ND&����ł��_�RAA�"E��: }k�G�T���˂N�ͻ��3�Q:����MZE,:?��-���|��SI�����ͧ���;Vi)ХV?V�SD�(�2���kA�a��'9ٿ���?�u[��&�X�q�O�&�d��+?Z����9^У�*/�Ĩ윏k���/����=�	�+
��l#���*�r��./W7^1n6��w&�������N4	�C1X�����V}���!��@#?/�`Pz㫒i��Qt��=(n�)���,O����ۗ#���e����?��>G��w핥�i|D���f������E�zF��d^�7B1��
�c���[8�<�n)�aW�v�/�H�#�7�.�K0��->�g;�)�}����� ������S~.\�׺�=Q��wx�J�e�jny]&�Y�}�FEn�%��S��O�Xi7��Rv�keA4Z��ux����!r�'v�wY�<Ү� D�$�-�#t��7���1��ɣ�Db���G@�����nDAajNX}���<tYڅϬ�!��@j���˞���+���,�oS��H��P����ɥ��Ğ*�UHL!�x�ycQ��me8���s�b����{(Q��)z�}���A��_͘~����N�~6>�' ������C�;���,i�/�/x��L;�ʁM�d+Fi�����Q�u^̎iS7V��M�/�0���؅]���t�O�2Aw�;\���D��ɥ�_C�)��Q	���=i���4SϦ�Ӣ^3��`��K)�m)����i���~2��4ئ�k~�<��S�C��y�m���B�"$���ZΑ�DOW��|u��cCϰ�s�B��01h7��$Z ���g��z�~�D��:
���}:k`�ʄ���Vp��X?E�
���[��f��Y��|�FDPm�Ab��?��� �kͽH!�`΄]/�&^����3�������ً]�N�ZTڽ��*<�x�z�o�?5~)nv�������ޘ�_�,n�d����Ex*`Ą/L����_�|洎��}牌{!��L��`�[��k&K4����-�_2��i?�e,���4NT�E������"�XS�M�M�Ht��*�����W������;���\zmny@@0�t�@<_ie����E&V�Įk;�Y6�gV</
��������#�A�o�⋔f�X��Wf��u7b�@�(����O�h��AmJ!Π���gM..�j< 	/�G;�:��J\�hR�PgN��s�B�t�D�~i���o{<��0��v.�������U���[uY�e���~�2~��/��;`w)�Ǡ�3�Ɓ%l��,P�坆B���	�納L��Z�V�,/�#�κ����b ����+�M�v#)�-�D]H�ݗn�%N�R�BY��$�����	��C��W�2�FLM��Ì����X8�B���;�$T��k�셜y����')%�Q���5��3�J�S�Q]�S&���u0������M�NJ�V�<IKd�����?������C����iq�����\�C]Jq���� �����ͮfd:_��js峕e�?���i�b��E4��2�DIҏ��9u�4�*N�'��SMF��G�L����n'����$���M~�wα;F��p[}���%X�]T�o�oY tX� �{AMC��m}E4'>/���ě�'͓�bh���wR���(!>zZQ=<�i���%Tr>�E[G�0+%=�^�y����J$�ǽL�`����攌3�	F�U=#g}1��P7�	p��q܅�Tɑ?qQ��Y�u��W���UI-PgM��r9���k�H����%�=��#H����0�HT��5DD�����EXF�v��iN�{ϧv�,T���P��Hld�{����ז|���ɛ�[�f.Dd�~D����)°����͝/f [�a���F7 ���}�3��α�������P%O|J���n�a`q����fR^�cm��\�T�kI�_������-��߄:��`G���cX��R��{���̩Ԁ�`��m�99�0�+��yC���A���ݥ�qz���B��g�wθn�&fE�#��[`�=�?��=�}'��\�X_���b��ʠ���� _��R�>����II����.�tw�L^-:����U��L{ 1Вً��cRWĭ�<�$.���3Xbue��9@��2�7mH�����l�;²�:M�lj�����ܷ�$�YD��i鑳J��Q|�����;R	]{�p�Ůhc����_�1S�r�L�7����J ���-�����~�R� F��L*�=u�)�#������NGz�&ӟ�i��_H�=�N<Th�l[�MS:���pO��,���.����l�*���l��Z$��\��.�D9p�ۥ��/�r�u��e�ކ�L"�x~�5��-���`?����z���/#m���>���pod�w5UI�R����;[���]4����	�������t\�5X�_�J��ga�6�1+Ss�<��d������XC�R�Z!��X��,���������iւ��#ҵ��0�g��X�������/.�:��C�G��_L��<���.Й��Ӏ�{�ӯ�h������U��ym�0,�޻���{�$�:����K*f���bRt}��%%�pD�x�Ve����_7!K�3��V�^`yP���u��A���Yς�I?U#��J�g�i�$9XD��%����S��W�έL�tmes���qS�f�P������zr�]�+��ݒ�'w�?.�Mh܀n���^dQ���E�?�K����ϋ�nT7���	v#Ȏ��е:����y`���w��������1ه��Uv��S�"�����j��.��ڦ�N�*�U"��8X%yq�U�7��x(�o��]bz1{)3����֨�	���!��ޑN��0SUu�w8�)���̲����9$Y7a� ��[}�	��+9���gn]��d�IK8��y�.�Ba��!�#>��n�8rrO����hۙ2�W������U��q�$�u��d�0�q���R���n�0d ���B�\�C@��ݼG���ظ)Yay�w0EA�0�ȼ� y�
q~`�R�����H
�~�����=�r��@	A��vZ��	�N�����v8�NG�b��I֣����A����u��q�F���F���Ġ�Z I�vg<0Z��'H����E��H"�"fO]2�Җ-�	�;��e�p��[�G<$�u���͈���.ǞD�M�y͔�Ut��0<8�,��T�֬t��^�cyM�\�ha�x��JgZ0���
����0b #��:X�*9�ך:����$��B���}��D������Ƥ͍����B���L|/ś-�f-�?��Ũ����oo�~s,J� Ȍ8���򔤺�=��xȢyL6b#
�۝�at ��9�dE��"�+�0˂e;$�҈֑��#�T�*��Ғ�ӑ�0^t�G�4��P���(
I��+I��v�����c����3���5�Z�i��e��˵�A�[�sx��U���s�<�*;Hz2�2)[�cŶ�/H�&ז{�O��΍�:P\�溶��$u`;O��UR�����t��g�ܷ�!\�K^I;��*��,��l�K^�o��n/����\&<m��)�.�+�e��#��#>��o 7�����H�;��3��Tb��x�$S�A���zz00�r۹�TM��a��E�������q(NGqB�0s{��G8�:g�=���¢4�e��6����0��wmʀ�$i�V6iL�ԗ�2q��ل���1�#�IA�Fu9�}���(p �{ �͂�[=���.q�ﭓt���#`�(���n����1l��y�(!	� ɞ�2ֲѡ*�9#�  �"�R�+N��C��F�|�U[=`���1i��t骝WCu���~�rw5ĭʏ��,Ti���W`��e��՟ᘜ��d2��*����2��+�H_6e(Dr[Yl�6��reQLq����ZO:�5~�<�&-�$����%��0�T�TԎ�I�o�&T(C�=F���D�/-�0��GUlX^몊���O��[7h{g\,Q�_�;4>3��FJ_���� �(���Qƭ��G�ּ��2��v�k'��fS9)��=24B�����?�Kfִ��^5�j�c^���_��5i�W�!�E���������щ�hHB �&:���/�/	��a�W���ɸ6��=��@8Q�"L@C�Cӹ���{��i���{}�`���Lp=i- �z}�Û��tK�7~-U˴��j�N�G��Q9��ɻf�1�m��K[:��ܵz�k�y�J�Ks�IT��D�X%Y����bC�z�F_��<�.�Z�m�e\9v"�UkW�t�9���޴��S���,$F^3Vإ�k���b�ǁ����I�߿U���g��~k+������i`ھg�ԢH�k?x��bR[@�&,�Rۢ���2�O�=�u����A/��p�!\���w�m ڡ����U�n#%�o-;���_�������ɓ}�o�..1B���Q�>(4�xὤ�S���҃x	T��egL���~(!2�-
Q���2A�?zz�m�܍�2�"ոr7�b�Ͻ��gKb����"˝��%����aʛ�) � (����1}G(�{���lK�h �����B"�T�7T;&%0A�A�31����_�T,��}�;���Z-Q#��{mt�8W+J���lG�6;h�Ȥ���~���}��;��1������X�n�*����A���r_u�zI�!y������\�N�I;r;��[<��o�Q%�ٔ���A�@�l�%
Ur>��\�WP����l?��,��%��������.���'�ϢQ[+<����lƃh�s�G�dr�Sx��AtF�0��߱M����\n�ѓIRB��w�0u̩���rW,ӄq@V(uk��2����"�#�������~:����6�8'e�X�����6�����֟��RR�;)-R��W��>zn�7�*���bj��^g���HIw�|�p��*��pK��I�:��Oq�l6����о|}�9�.f P$��E5 lt�]�8T,%�I���	���$�L"�p�&��u�V������1t��|wb��)�K{uu�gT(�p	�!�x�vW�̋�Zj���*/11�F��%��G�B�2߯�st��t�^���w�s�]�<1)���'�;�v��!M���E<cE�Nݨ	�)���E�q��SDdo�hn�"8���� .��␽��H��T.�� ��S!�X/M=���cB��:��00��"�+GF�X��o�7M&`���-g��&�?�z�E���<x߾�R���6i0)��/�^��\�ȨRGx5G
�����n۵Ѳ���?.3�LG7r��w!Z��ǰ��d�E8��>�L�<]2�8-�z'�WY�Ь�2��CL���A�.ݔr��O��&
W�
>ed[6Cl�zWf�R�Ӆ�ǔ�c������\�{���^�-ܹ$�G����4�g`,�q[��Q��c�U�;�P�i����襙	.���sOP���j���B�j�Њ����;����tk���u�&<�sp��k
l1h\[OELꢮ��R��1c���9����z�㫌ɜwN���:�W�����!��sUO;M��SE��|��.Qb�Lg�kv\�i=�(���}���`��l  �+��>�Z�P�T��~��)�ӏA�Ye���v��x@AD�H[��`��"�b���	������q�?s[����4��,@Ӕ��w��Y,����^PR&������>����B!?D8
dn0���Q6�>������c_�?�)< �!|�>�0Q�yO��R��֭�u���W�����$��߹I .�x��=o>�W�$2;��J����r݋k�`�W�<���;qQ���l��Hm4�m���{�V{#�Nt&*>R&`ܣIc$�g���Ѧ�h�����|Ĝ�����Ũ�r`]���;�:>+5C�i�1M�=1A�9?�c�@����X|Vd����J��N�~w����g͌w^����B^�@+fv(�`�18=���쁟����Q]�W�u>�p���+��]��4�����ykv�Ux�-Bv�$h�4���d=�D7kb* -����Yk��=A�@WŊ�Wp 9��uT�I7�r�&+v���H6���-�R��^i�.��9�^�K�"��R`1Զ�EX7��7]i��j���������e��������E�0+I�`+�+�\����*�RʈB���Z��E��F�M�p/{��ud�RS���',1�E.mh�ǉ����*��Y�P_`��i�r,Hu�7(
_PA��ͰmSj��L�JFV�=(L�+��E�9�>H$�a��`ݕV�a����*��.a.���D���x�ߑK�#y
���=,�����A<��0H���*N4��^d�CVn�sz	XCN��Tf���=΢��_�"�;���S`�1 ��Cqow��P+��+��>>�ɓ|�~�8�|SQ��Î��L�ߛ	6/�A��lh�,o��R]��U�KX-������;.s�ı&sP�'gO��tl"q�)m�"N�ӞIP|�߂�̋ۧ�J�����nc��č�#鿄5�١v\�Ң{,�;�~L �^�E�1 -�)� �a�IۗW�%B�Y�I�	$@oټ|j����[ ���#<�r�B(���_����]6�C۾[��$)M�(V����)kT�î��[��T���$-�����qd#��VI���������[1�>q� ��z�.� ����*�߽ն�κ���s	�?�m�p����+��26��=��+���d҉&�uK�1�9��!;}���(�k���DQ�qV���]bK�����zQ<^u��
�y�����5X,ި��	%�V�h��p�*���w7�1ܛRE��%�Ts-}�bv��o��o��aj0�/٘W�T�8��W��-/�y.�dq�u�?ߤ��˻Eq�C�#��1p�lYg�p�%��j8�zQ�Ä\C���}�h�RF���� /��|��Ga<d��D9�+@8��u[��/1A�F��l�b�P�0؀V�v�Wi6��j�q�]X�Ŏ������9�U��mp�z�Cl�]�R�B[?���m7Zw�2#5h�5���:#xr!yq�8
����#BH~���~�Z�`�2�T��?BK�FT(#�v�Q;���q`��r�Y�X�W�+�8&���6j����|�1V"cPA� ��� :q�M[f����IM��E\O��b#|�BSxZ6)��e-��##Y4$�O4�ɞ���AB��ܝ5�yt9Ɠ�ܤiCϧ!lnμ���h,���8���j��ӂ���2v�"�1�K~��נԤ��ۢ��vA��s=�"�G�c�\<�金�H��`�,�c�(�4/'��@��}Ůӎ��b�+t���Z��8i��SJ�o�U�Qi���>�`ߒMV{Yaw�����q���-�Od�ː)5R\�7É��}E �+��J�ֱoL&_�9:~�5c^��H](�t|;m��4�4�C�5�JĴ��Ob ���=(M9V5��$!�8g�j/��d�����<�1zOռHƪ�}��0�(:$F:�=�J�8��}gF�������`M��N��6�}����WQ�wp����j�Q3jƵ�7���j�|�<�	c�Ql��M3l�J��9l~���JCsJƊM��z���@)����}8s�6,�/�<�`�7�&|�B	�ˇ%��:�S.��1�4�F��9�%�>!��1n.�Q��T��o�J�31���%o�:.v�i�)9׷)t�ɣ��aʏ�������&9a4@�G��"I�I��\�
ux���<�Vc��LI�nGfB�t|^XKqr o�t�U�������au���d8��$�v3�
�I�����K��8~y^�5:����Q�x�����l��c'�XQ��jgX�lR�sr!�b�ƬS#��͔մ�[`x�60Ͼ�u%ҫ�D��q�}��CkZa�*�'�i����uw9ݬ����c
Znm�1Pp�:���U�{�LӪ$95�u[�d�W@���y�x��\�W
wC�c"�ꍱoA ޡof�����Hr,�DYdY�Z������ڕ2T�˕o�vm͝{�z5қ��7�́8�p��Ls�o}��_����~���s�s"Ib�F<?�!D��Q��e6�lM�bO�̗у����N<͏U�M�տz�e�"��/�	��g�+��g9ܽtmo�ؤ�} %1���c�-!��Sӹ:E�Cw��5���r:��,̾Q�y�|4Fb�M��,��t��[����|���6E ��5�s����+�v�3�ބZ`?�Ἢ�=^c����y���@S�b�'#4�<H�@�MFK�}a B���rRէ�):S��e$���Hr�Ksƒp�����b��)���o�c���*�
y�g��K*yԑ�ը�rƺ�>U�*�x�dE�)�r�ʦl����&��%�s�-&"�'Ŀ+���q��&�~<m?���S*��vZv% o���]袙�e�^���vG�V6�����¸�ɐ���ڙH46>>�F���k��Xs4�/U��1�a��
5��DFi�����\kf�Y���ltYbi�	�C�3�Ի�$°��*�a�|͟\7�<��ŉ� Ѱ'&�&#����r�ofj�/jr�RUg�Hf��-ɣ
Z/|A�7�
�c��u�C�O��<}l��:CB5��gkHC7��ba�J��l��P�I������t̺��N��/�4�V��{����	1jxm�%��;Ɂ���0mB��V���JS��y�*�O�BL���Ӥ�Z�j��Ua���)�����X��Nϊ����:�bX���۵�&n�	'I�ӼoM�R7+��u����+a�L��\�QVV���NE�k�f��E�g+1ѿ�CU���x�9	�;)E'���#ak��Fi��	��n��<�U��M>�}0VH8�e�>\b�Aր���c� .oR��מl9���~���]zIީ���R�}d��A�B��*V����'��Fr����},�i�$�ʝ�q�7�݌X�����T#j{0�sH�J{pu��Mf�d�h��x�PʰY)�Ɵ���e���n�����G��c)ņ��	�����P��=����VDy*��[NE���^O⟑�mO��a	��VvY'��M�ui���p�y*0�^�}qb-Ϧ�˕����ȢvZ���&�oi��4 ���a��@aTд���,����f�l�9R��-������-/���B�U��ʃO�+�
�F*}�u,]�)P͚0�]uH�g$+4�OJh��륡�����*���,�X����5�o�����!69���j����vxkj4�^��J�-�)��C��`̅(���3?��]�f��� �;_q ����Z�!Y�}�����JZ� �
�k�a�z���������=&�?���9�*m�L#��yCW����jC*��ܟ�1+`�ѓ��2�
� `��ث�gB�zJ�|R�k�D�,���l�Cÿ�%j?�4�O:2(C{��NFm��`7�r�J{��t{2fQ���Ts���Q��E\��^	���:���K`K��(��%�ޡǰXYy$���g^���B4���w�5���Ǩ�� c; 2)����ҷk]#"��.3z��PIʹ��P�ݚ�v�{����B�|\�`�y�����G~�?�01��r�{�,ΒE7���?��J^�P�T���b�ܶ�l���K�M�j[�����`��`o+	�:�YΪ�U%9��F���1|~"G��A��Z`%c��R�Ɗ����kW(�
�CxϽ�.:���@ɰ�Ʀf����3'���K)�S^��]v�I\t�洀m7�>-����`&@�<�,�S�� �Si��r���>p �Ib�42AŎ1�n�.� K88�5�A�7��w�o�S�o8�_
����j����{�-��dp�`M`�Ӛ�C�ۥ��j��>A���$^YN��{N�!a2q�w揜��Z;��(�~n��/�O��v���@�E�:�
 y�+�̐�G�Jܒ� C�'s1bx��/w��3���Mx	R$�F�"��?���~�i�'�@EJP��k���P�&V��%\�}H:NP8b�b�����X4̷+�7�h�y�.����ح�`��ڪ69ற�I�w
(���F���;�%t%ߦ�?�����ǫ/��!Cy��y-W����w�cw�g����N��|����h͉���ѱ�̜�&4%�9�|�S���%2*/��k��όz�:��Lȗ�헺��i����NY��5F�qcL��5"�כl�u���'; bG.T����U�o�@��΅"@5B��M)p�������l���m(�{h�i����Yj%�F��q���t$�#G�]DTȒ�����`�db���X���ؽs\?o\�_m���i���P{wN��ΰ���@O(ݧp�L�=�s��qH��h۞׭����#/f�� ����,'��}W�ϒ�|���Dp��m�C����th��|>�V]m��N�9��}1�S����aBFIa�":V"���(d��+�Z�^����/�C��̏ݾ~���2 #� !��|��t@D0�-��?�KSah�
g�͈�y�7m�V�P�&1238���p�?��[Ҙ�}���ߝ�f�
B�ԝ��Ǯof�=/�����v}�S'g��v�����+d�T�0��˞��u/ļ>s�X�|������$Ù���H<��B(��L���!��vwK8o���}�?�-��֔:����/	�y1�7A�!b
�v��L1��dkp�أ�E�f?��8�	{�E0��Gݷɑ`Wp�5M�2yŒ�%�~@�]����^1�J�x���-�Ć�R٠�04&�=j���R,-0k���_8��t�'�1��������TA��	�y��V�	�aM��XS�D_�n#̫���?;�+��>+�Fb�=O�C�T���pqz�ڍX����уy<��D�v�Iq�sѭ�7��(),}�-x������]*r��΀K�J��7E�-��r�t���9��rf�֦4�S3W�a��-�>�>�%��5���ֱ^TZU�G͂��v����p9Pf�=�57*��^���-\(�$�q�(�]}a��5ȸX��8���uK{����-�E2U-h~��X��\xX�	�˄����a���)7����:�����Ǭ��KJH�9�i�u)1=)2w�JH�yi��V�_
��ɹ'U�$�f
��l]/z7q@x��?~˼�����Ie�}���C���ʌpw����b꣡��v���sd���c_j������܎�&�[:Ÿ�p��/������(�y��	�t�8Oǡ_w?���td�\�O)1�����
���mf�{*D	�)˕Ƣ8�;jz��~w�����c;ON�nZЙ�YX�f;��:f�d����,��(���]�s�:���=������H� ��C��	�l�YLk�`��n�칮����Ofڨ7��~�������S�l�c�{��z�������=F��_���7"}
���~�jZ�-��kzҮpt�	�P�(�7C�-=�@��:�e���!�ޫz�+y��#qi)|�8B���p�A�zV`Ͷ�����M��fS�܏���΋|L��I�[g�̘��b+�'FsӘwi�T�%��*D��/����\�vKA禚rф������u�۵g.F���$��%���7����A$6�)�)z+t;�0�c��\�!=�GY���+jP��O,�Х���������r�>-r�7��U���|Ǫ�pC�k����3��&��O�&�3���8�:��0�ʁ��j������Iځ�H��Ip{��}�Lg�.��L�UD3&�������A6���z ������=6Y�m�CTqO�n ����1x����Bm%�����A8��a���jm�)�,������3��*F-�{���;��MmB��/�L�	I�o�<Iy}�#�C��n[�	�I�8e{76�ƻ�|�r{p�W/f� Z��*l+*�|�ҧ�P������1��]��i�͘J`���~�y���!{$eʄ9GV[�
ϥ��DM���C:��I�߻ԗ�a���d%<p�(4��w�g���r���o���v����O����w��m�,'�Iu<�6��w���IM��SO�Է��`���0�_�}DP�$�W���UM�)&�?���0�؎�?n-�*ϥn�8��n@X(�f�Wj8�RL�Ţ�,���q��`�  v��=�ʯ����c�mf'ǼKv�H���{������`��v�x;�>�:9ìW��YW��%\y�z�j�ڿ��X���[�=���:��䫠��o�1�@�~`���E�����Q���R�6x����|��H��n��o���	@fq�g������s<�b�$�8L{B����|�i�Q�/�N6	p=�⊯\��*lAa�I�}��gɅi׻mrj5�c��>�>�!͛�3�op�R��}m������y��+�J�4B��1����^qF���|�q�p\=�k!��L� �H��I����áQ'��nx��F���JV�i<�D�b�D$x��G��x��ƻ	H!�JC~�!�x#�2(ņ�4^wTEhwq�V�H|X���gǄy�l��x�B6���v��I}��c:^Nw����,��ߊ������Ƀ�Ѫ�O[)�\���>^Kb1�K���7Mc]g�����'�|f��(�����UM�����q%��b�m���r�o�6����C(������*�*� L���d�c�,]���4�f�<q���~�C
th��6�dZ}'��
�8��{=!����k�c1�mL���z�X����j�,t�'^���˕�obI���huA%�쉍:z��,�h�1
�����?�Mp}+l&��<-dt��~���؈����QVk�c�`�u	~��@�{@�@�X��h���&ax8�tg�APqI'�	����7!�^�1���=�yt1����^������Cl ڶ[�6:w��(�v��4�����`�.G��KB ź�����f�� �����X~o�t�y��6�:C�G;�uC{V��� �j(ǋ���	W��������feu.qU��O����(Q�öp @֫��vÚ��򃊄�i�v��u�#�ۼ�"��p�V̪{���g-]]�`)S`� k]�K�`n7�?����KP�]v��W7A��'��6�u�O��u����:%��"�e�EC�ˆ����V����|jq���c]���WA�>��B�q�U�O�%SȰ�{Sv�cgS4c�^��JO���^�C��6q�s����$��U|��nR2J!uH�+�����.G$��F(�����H�T/�Sׁ�l���qg�'0v%t0�%��4�(��Nv�!b�l�`T� (i	����&X��R�50�L�UP�������_XW�'5찛�Ǜ�J7��@����vf�w�l'>����7�P	N����{�ܢ��7F�Tɖ�9,D==�Yx�	ts����P���$��Ȏ�M�~ ��&�`j�܋^4����a�i�����(B�G���
�?ꈅ��-W����+�e+-_�>݈���y{k�Đ�,�X��;�A�C�K�j{�9�_�3��6�2)��/w�.��{�������l�S�R��~^�?��'h�����l9�\^��ǵӇ��wR5��� �[%ld��9	����?�ʉ7����\���]���,�&&�����7Ǌ{���c�OG7��L:��+n(?N/;ٔ�"u*򢯸[�x�=MB��c{`�v�@ �,���!�`��R��=O_p�������)�e�;�ҩK�f�T��ZXR��,�K;�L��:O$@B�3JA��d=Py*%Te�a� Wxz�5?�w�>^քhe�o*_�f�cL���x�ϝ�WA��|H�W>�11�*�&P�O���b�r�L!ܼ��o��4�(����rB ��W6���2�;��l4nʷrᇒ\�;sؙ	��s��7aV��_��:��f*z�h�&)��*n����tM@j9㫄���U�?\#D��N�D��{��o�U�+���s�"� �Z�$���rþtQ���êƄ��O�����#�'O�8�sm�zhDJ$�������8'���jy_�����Q��x}*��E���Ç���޷D]�ss#\p����7��ܯ�k����D+zM����>������l������#�s�!�햞����x�kF���*��Z|�L(�B�0.�~=���f@�!Sed��~8��l�2��˂L��_it�Y?O~��t��g4��&�pz��j��	�&�^yN�z$�zzg]���'pq�R@s�\�t.'�>�Y9����M�}��Ԋ�@PqT�\���腵�x�4��zG&�
2.��n˻�C�i��ځ�Z�W������ �\>�.'�?��j���o"�SX�oGʸ������Z7ްG��3�x�J]����Ͽg{�H=��;_��#�np��3~���Kwڋv��H�Z2l� ��N����'wʕm�@�'B�L/����\A#�RP���'ȷ����5���j���o_f�⌟�*�M�@���Fc��,jb�*ƺ�V�M�/����~D�b�=�_�Cm�_M1\fC�AZO�X���:<9��ƜW�d���ݶf�w�u�@��	�k��}�J�#aǪ��
)X��7ٰ+�`���.�:�d;DD�7��S7�}�A
	)O���=\l�ҋ��۴ zw����C�-����*�-T�΁��/*TqgQ��V�-�U	�HT*n,$�}������*E�mT��M?��V��S �+ρ6%�r��I#�^v�a7޲�-�O��X�	����N��c���_g��贵}߮�^��c���z��ZR�=�0��(���[���_�nljK��Ēs��+����
����jja݂ɀS��3�%#�T*ƿ�hɭ���9�G�2��y�`9*��NX���w%C�E*�;K�����٣=#���C�����2I��	�T�,u���S.j; #
�5B_��\t
����� 5F������I�)���$��S��-"G��Ꞻ��-��.W�FO��Ny�9�e]�\[y�3�����U9����Ӹ����K��K���}>n�g�Ee<�	]K�xZN��/N�=�ϛC)�������,\��PF�?ѣџ7�oG	-�_
���s?}����� U0�|��΃D��;4�P�> ���恽;q𳹊~5���v�Kvb*d���Ը+	eO�G�GH��)?t�S�k�^e5��g�QF�T�
g�?Y*�j���n��P4%<,`��0@m�>L�\;�vX.J`�����2?)	��1T�p�L��AAa7�m�����8�Bj�7���X�f�b��S����a�AQ�������}�Z����(�}����m�7�YɨW�pdU�
L2c���|�"�b�}+}O��U�S���JU?8 ��W��@�h�l8�*���Z�/Aۉ�}a.�4�U��!�=�{��"N��iD��&�iM��&�	�/F���Ë��r�]�6�Gss���\�ɍ�&�����2f�S���KKQ�}Y���4��~3|"�(�����[�j�Q���Ja9�^X\�H��H����_֏�'F��8�uOn����_z�B�I�\�����vy��&}�q쁟�@��>�r��R�|pG�5����2������78�i���S�M���	�g�0ɑ{M�P���m�9���G����d��Y������%7a&�\���~�H,�4�$+��afS��lP�Θ`����>�ꥮ`��G"81ͨ%Ao��逛ʘ�X�_X'z�ǖh������2�@1]��aVf���y��V~�-�q�G�:��	���][&2�2�'�o�qjp,X����, ĻJi�j�^�(�b������X���5@W0�R۱�����5KX�Kv8���. �"�p��r9�ʃ����!F���ݐ��� ���C&B������5ߟϿ>��f-��M���e�Z�5���{r���̀��^=r�y��}�?׿t��`9^p��W����p��<��ܯp��B7L37�n����f�T�8�l�H��;"�
�G�~C�Id�J�3W��.~s�,�1��������2�'5��#��@�b�|)����Zr��4��E���\6���۝���~���ౖ�0O�EgF*]Ԋ	�:f�&���pxfyq:X6�W�1��Cq1Rd��U�XiR����Y��y6���]W�PN�����$&$
��KK���
à�1&����x3�n�C�7���M��1Q8�%�#�c\�0ܣ�gs��)O+^�����1�g1�2�s�$�āT|��Zᒷ�	``j�2RY�T5�#-a�@���odI<b(�{!Y����d��&_/�+�hۃ��Hz�(��Q���D71�eLJ���]�c��.+�~KZ{H�/�9Y�j�<��s��R@���6´4�G$� 9.���݌��j�|�[�L������
M�<�LMNJ��b�t�Z�+�=(����غ�#o}+����\��*���C��~{�	p��<�yF����M�0�ܙ�EN-�A���g���<�
"Q�Z�YQ���'ִ)"B���m�E4FB�aQ�tV�E$J�i'Cx���?`���F`0�bj��h�� M��c.JW�R��.�o�9Z�f����q�ы0�S�=W�)4����SGI�����E�?C2��I�2�|���{�r7f��pQ�(���;�Z�����C�'��3dΞ|�Dc{�M�>�N_-���(��d}J6^���E���(ȹ��:(M�H�Fx|c��+���ё�/kl��S�Un���$ �����ytѤ`���2�rTD#��+��TҨ���J���'I)�����A��,(;��b��p�������{�-�M���I��g�������2U>p>�F�����4!����?;e��� �d�Ij�W����I��ʔq�h����qQ���g��kIm�g��/_����RcdK�S�����(3���=�+��L�á�˴�����)�l?����L�W��.�$������ziCJ]8����r��:���a��F�䲛?�� ��,�HqiS��;r+0I y��/��ni�ׁPw˴��0Y�����4�Hxo;��1ϊM}7�Tz��0@%_���X�|������l���5�D�D����d����)_,�-8\�h��7I�C�P^� ���-���G���+t���=��̜��'��!�d<���������ߒl��/��N2Y5��K�X��SV�P����;�F{n�H���7��J2�8Z��3��Z�xu���W��N߫a:�Ѧ�pH�[E���$]h�&��&��m��4�a�¹�,�Ǥ�����P�&��꿑=Z���r�`���~��80g)}���F1��l]��;��R��z(x'�������>��ogT=[9�+'>�}������v��N�5���螅Ꮮ�����A\P�Sw��+~>d/�q,��i"�ׅ'�{�`������N�f�/���J�:5�+^�]�5�$4l.�<�nom�	�;�o�_�$8�a��Ug�z�G)�![��2�:u������b�-��
�$�'������kzFO�3c�:�{+��͚�O�.Q ��[G�.Ǡ�%�B��x ���<�q��;���P�e0<^P�"�kp��ڷ���T���Y���˳���W�,�3�-C��y����K߻�e���@��|� ܈E�!a��5G��-٨;�q2�LFs��$�H9[h�B�v\��ԃ��9�fPэSf��oFP Z�iL����~�	�C��ݝfVFd5f�, ����u2�<@���i�LJA�6�NO���m�?�:&c�Z��t}�F-!���*�z�5N}�svu��OO��Tm�I�Z���{��E��O�A�>}��[�V+�u�څ9�c��?�c��o�%���(�os�l�&v�"��ǳ+)*�du-�QTZ� �A�{�9���P���'Q(�Am�W��eS��u,��>Fxzp�\����fk�~�WX��ny�@|TZ�0>��:j\��(�T�z�,�_�phbI�;�c��!��,lm4�G!ٳo�������J/3�g��L��R9�G�����u��;I]Y	�p3��*�A@�1/DF1�5S���r�<����pO!m8��7��{�dL�{a�U�}:VAə�r<�?q��/&ܯ-�4\�<؉���J5{V���K��&��粧��i>�֭�����@k9/�=����|����z_�@����E$�8��oB�nա �|��@�<��j&����ҵ��M����D���N������"8LS3	�a�HAg�B	4X�A���P�J�~�䐛�z=6��YsQ�����P�x5!����c�%��"+�X#'aQ'7
���|B|�I�	t��ʇ������8:���d�y�����xS�.S)�8�7��8������S���X�	f�g��դؗ��5h��n��֩ۅ�=_D|_L�˥�5�	~l%$�������=H�a�j��}ʉ�����m��a\��}�ۥ��-d[օ&�TO���dkq�3�,\`��e%��ӆ��m(����S�.�@��A�?��&9�
cd�2�b��_���rSk�����]x[�|cA�
���SXj�t3 �:�!p�Zu�(<p1p���36�7�)��A�;Va(Nk���v׾Uf�x�����'h��J��es��/�����=�8ĺ�W�x!� &L�X=�S)�e.��~���^@��?~1R�%v<�� #��Ahڑ��GZ��4��}�����u'�d����
c��[w�أ6h�ʍ�`��q)B�p�Qۭ�.��^���_�c3����}�� P�^��%a�V����	p9�o�%MJ�B��}d5q=B��t��?9���;`7������ L�\3�f!���=��˞�x�A�>E�dm_L��S腹���hM��n��!ǽ�ӡ�P���/t���VH���e#��dk�(au�n.�G��!w�?-�"a����^�J�N1��N�������.aR���R��3�E�D�<���hE�\W��a�ߜ�j���b����*I�5��������@��gؐ�lk�i�����	`Hg�<NY{�q��͘1����EL�⅃��:ڷ����؞�ny��E��F� [d��e��Z����U��ǒ��-������`TP)�쵚`}��R�o�xd������Q�F�ft����U9/�<������)EN� ��G�eZ�?oi���h,��1���2R�;ި��!��B:�[!+\���{8��ä��r%��/ �&���^�g��G�S]ۇf�Y�ҵ��)QG�w)�2�����p~n��+�����П1�~�;��bJv�NL�����"����`� ��&NȼZ���r�xr��B�k��F��MpQ�R�e��CN�1��M��b�R�~[hۚyH4���)aj�R)�����Gf`� m���G�\}�q��M�nԱ_�����B�y{�����G��#���'����z+K��uܮ��a%��J��o&i��b�'�Ȯ&�����_D�9_`���ɛ~�/-ܖ�,����Fw�Ɖ"A,ɿ��Ng��@����������~���'�A�>�
hg1�?��ڎW�cF��=�kA���3���]�\����ȸ��ț���7�^�]4�e�7b7��a#.����!�Վ��ѩ�+�,�����`ꕇ^��y
���0��/|�&m�&����w�e��l��B1��~Fq��(��S[?�X_cOKm�Q���#�w�~� ?C��x�#�;�C�c`QN��c6GD���2�N	�����-�k��۽-8�z<�O�I~�U
�spu�a=�%�^:���� 0���R�P�(?x��P���h����F�[7̐�V~s�Z������.�7�!�]�ͱ��c]��2r�~hiTgSQ0g���x��d�s�K獨*Io�Xץ���ݚ���M�-���E��0_z���������d ^X�9�Ή�!<Ԧ�S��52�'��`�6��h�#�7�����)o@d��g5��٨R(iY��Nc������Ԁp<'��In����9�9���l$[Z!��ʖ^p�@�n�4�ܼ��Y��wwzI�-)������Q��F�x������<F��S�)��_�����,�����O6W?QZ��?��@5��Y����Vh�����ɻ��D�29�UW�e%ֿ�Z�T��8���Z�CՆ$l3P%��. @���i�rc ��F�Z�І$���I����8dNU�⟢m"L)�f/:,<���U���K���[G?T�֒J��az�hܴ����'��#'�
���6���	���;^�����\���<cX�0޳��8�(��x	. ��c72��5���MzՏΧ�wH�f*is*]�A"�H�7Qm���c�M���׳ׁj�p��:�y������@Ws��.��R�?`/C����Mv0��S��!�cPx+�����ɑ��K�d�8�s�c��`e�4���y]��f��z}����^AG�\�L���V1�
uu/�	b�?P��TX{��Y����&��z�zUG�M�"r�)3A'��D������ϴP�6]���4Θ�=�T-��ǳ�b!`.@�֟p��L������-8���󊂛��
hL��S_<O�6�`��x��%t��h���y���:�� `F�X����K`��9��
r�ӳZP��m\2����R WМ��=�ͺd���܄��M�!@O@u�'h �)�JDs�g�_��~�M2`��Ȅ�%%���eL��1�?uߔ�~*v�K���b�� m�}�";��Ց��]��u����k��7���݆c�����#�~]��]�K ��ےY���A��`�M���s�w$ui�������)"��DI67�(<�2#+�����0���c�4XR�Tm�C���Ő�ࣇ�bv�����P?8㊚v�J1?o�I�2$k6��Z}� �ie
#	��P-�e� P�o'�	�W�K�}�������9�G�ֈZ�G��=,���K���	�s2ɝ�9N�5�>-�]~]�S���Wܟ@��/m0�.�ߔ���!͢�T��?m�Ǒ8�iv(Wp��ۊ�f,��/s�z�a�]U�9 ��li%m�=)��A(�@��#)$ڦ�{D+e�L��O!an��;�"]=`��?<�G�a��,�B�.?�{��^4�>�Ts*��M��׭9��Q�Y�`o�l�=k%z���@WV�I,����Q�6�Y5y�9�:z� �4�WO^�M��`��k��'�mȥ���D�gB&g��,�<�-9���ۓ����#u�ku�F�_��֫�I�!sDM�7H�p�B_��}o�}��n$!ќ䍒ON$�Re_e������UVt�{R`�s�<�=���w�o��O����h?.��m�sXkc�ud(��\h(0���
N�8M��<H�"��Ǳ��Z^C'���@��1!�;A2p���]�Ӱ�����4���@x2�S�R
���N!��%�e�~,�����?Y2M$����>JU�Fv��w"���|�����k9�&2��a4c���3��Kyz|��B^���8�����.��	��~|z����w�`�c��v�j)�|���VF���� �X'�VӊV�1�!�l]����,�eGݛ��ʽi��]9��n%�����іYh�D!
wӸ4n$��A���1�N���k�!�'AW���_X�����P���E�8��XX�1ƕ�0I�˘��5�;�����Rb�e�P�a�-���Æf�#g�N���aF����/�ƀ�"�sȟ0�}��6B?�}��h�IEEʆc�s@�m��D���t������Z�pga��yeR!0�T��H�Χ
η� ���,���� F�u]��vWv�.�8�(��{P�f{Dכ�mg���@��8��ཤl�������(FnK�l��M:5��o�ƅ�hQ���SB��������sOj��o���q X$�L��3jh6�.]� �*�6�b.��#��ÞP���D���g�8wY�b��oqȜ����7h�M�Y�A�����#�����G���9R4>��}9���!8K�AD T�CZWC�~�i�"_�rG>����ĝLd-Lkb|w���?��>W2;lX�)^��a[P+���9}�v��D�{A_�I���1 �eQt��)���p�{h�e�d��dC�ښ� �?��^VA��!���2���{��ȏ�O�
�s�K�͗�W��}�=	�M�� ���kr�k�N�\�y�o��~�^��P��&��l`�
�Xǣ��*z��#��M.�/wl����կ����~�QYKW�S��Nr�>^9�W�g䷧w���uĤ� �q]��K���b .��pA�Y�wW��O�)�@�S.49j�O��=����]<�ag�/�HN&B���,dw�8K<'�,'z�\I"aH����*V�$";\��q~�tJ�[��R0�.45��{Y	'��X��*���P�؟���b�az������~*o�]>�0�o���6MtX�٠ُ�����^�!�8B�:ZoW��E��%������0.L|\����R}�a~b��v;a�k4_i�<NK�=�C6��y��*�U�]���9A*�њ��6J] Ҷ
|�ô��Q�kr��+�hb�kV�7���)^ϵ����������I9�_���uEn��r��VB�����

AԦǽS��A�ق���:Nn��i[Q�Z��~�V��.��q Sxp�J�f�h~1�0�+�!���(;�Ji{WM1��M TR:f�QOf���|]��@u7�D4�# D���Ԍ߻ME֟���gU��X�w�A�n�H4h���"���A��o�ђY��M�a%َ�����7��Gղ*uYN��*���P�Ri����	��q3�qZ&���eq:Ʋ�g{_v+�����������Y����y�v��wzW�+�[RL���sk�sE3���.�e$�w�K�N�5eai��#ˏW��y���jbG���D�Kd��ge�Zbw@�N�f�6܊�U"*N��搜�����l�ԁ8x���^�s��t�����v Z�K�>���P;�"�V�-K&�T
S�i�������:P ���=_ܥ�&V;�L�ډæ �I[�.����0M�Ȱ��~U��X��`5��l��]��2{�/L��I��~0���[��eD�G���'[��Z�����碉Aj�n������]��\Eh=[���%R�q��Ҭ�d\�[XK�U�?�$�vT��ǉgjr������<Y��Z/�@ ����^�G����+X����ݕU�im�ǣ���!�����DL7�Y���Lp��_j~˙��&(��
�M���9������_�W?bZ���a�`�PT�"1*�;�p��T�1{J'�������k�ːP'� ��]�P���?v�3�N��N�c + �����n���r��e�0�5.�7�J� fj��+᥾C�yZ��d���Ѽ9gcՅʈV��*�����X��q��6;g�'	{�UG�w�^Љ3b��wy�F��/:v�?�?_�c��x@yʹ��&��xX��Ŧ|��qH�l�����`�Y��d��(�#%rY�;e&Q�v<�;�&�8;�eTl��.K(Dt�T8��ҐT|=������t�j ��	q��|A}�f��<K@,}�@%/e�{�OeCF�
�ʃ=1��K��_8����B�4i������`z�*�
9�P�pm#���c"�z=�!9�şE�r��2�h��Z�T�����y�*�̬��W��U&�EV5�5e��l���D�Y��a������?�$낙�J�B��	���m/�yݠc��~�TS�=m�oĲcR(]5�(��M����Ţ�/��TM����{��sBg���k�:,��ƻHp�i�>�>9��a��5B,�7qU�Ќ��fژ�*R#A>�'�h�i�A|�V�,�z
"`�\�\��Eis�N���{�/����o��䆍�q�a�%*UJ��Z�o�	�v���de[t�.�3?#��=_��S�}.���X��r���'GK.ˉ&�{ʣ,�����-�u���F�4���J�s��̛e[����
��3F��fD2�����++�Out��g�N	�[<Pk�����;�����zG2����~(�z	h8K@�T���Ae������Q~῟�Ű,1ջ�>���CT����#/����u+.���aJ:Eޙ�;v�{�MᳪH�1�?i΢ۤ��0���"O+wZ�H��ϐ=c����Qw�@x`�#�ˡZ�2a� �+�*u�o��w��O���ESC$t�y#���.ϯ��݆��qퟟ �=�����+�<�f��*m�EE�Pg����`�e�3uv��զ�J��,���p�J�������sྃ�["�F�y��y\�ɃC�y�v �+� V�TqsH��]�r�%ߔ��b?.��u0Bq�x��1�/��<����o,e�oÇJm�!�:���@(�UE<�r`�P�%���Gc�B��E;i�DKJ~LXdx|��X~£�\� ������d�S�ڹ'Q�r'qWS<=�2�@ϰ+�y����#73�I�)���jN�YT�z	�%/�B�]l�Q����a�]�=���ȱNO�.J�?t,z��~�V�_I����p�C-Pruf�dW@6Vڬ��Ƌ����{�0�o�Ԓ��0�V���������/��m
\��[¯�EӲÚ� �$ ҩ
[�^����ۮ>�/9��ei�$*,�ɇD8ks=tA�cْW,"��r!�1�r4 v�M�<���C/K�W�	��K�rJ��5pݱ�|S@�s���G}P�8���7<��$����Y��z-+�jK��LB~��A�p��7l�6Mۀ�����`3���)�t7 8���|Cr@؉�/op�$����4y放�j�dNq񍣩��&�18k����Z����D����D���u+�Q����ޚi��֨8����̉�h��u�Z�lүqC���"���jK�Q�J���(3^��'�dC[��4`g{4��ɴa�d录��M8���?�<@��EMa�#0�q���q��3�|_R�
�]]�-��"����笏��t]�; �ҽ$�
���8��b�7����>M���yv��5翹Q�޺C�:q�,�p:����LY`�u����>U�sio��K�3�^{��U'�F�>oג��<��6�S�9sH��HC�{PI���SCZxQ�/6���#������45lϣ�?�+���_���f���k�pZ:؉��C�%46Yyp�be[�[�KZ�wA�i}ه��zD�@|�.��S��+�)1i��a��.Zx����<���ecCTg�/M�J���20���!Ax�C����<Űi����X��1�e�F��5��WCo�bkhU{�̤�x���OHA9^l�I�XNTu�0H	k��_U��fOT�7�Z<����d�@�otzʩV��ʒ�����s�|Dٷp�%9"��QQO��:���CȹE]�c�ܗm�K4������YQfy�1.�°JD�9S��������t��K�[�O~=	x���;�'8ƴ�q�Pp��3�]���&Y��"�ؐlS��i���jߛ�� $@׍��>&�M�Ƀ�������b旐i�ڒ��R҄��Qڝ��o䪉8����'+�wo������a|�?���Կ�ɵ�d�sm��V�m��u��;���p� i��pP��tEz
%�TH�ް������U��XM�ҭ���V��<����Aޱ&�m���l�6I�|��h���[�}��^���#|.�����)/�<QYͷ�B<��`Ya�$d�p��ڄ��ù�]�ܶ�pB�@�['w9����Sg�Ԋ��U�\T�懖;Ë���ڸ�2_J�ԍ'��qL��r�������Ļ���$y�Pe�r��ׁ0�p�D����um��{i��ԭQËM�>���H�o5/������K��J��L�K�b�J��̣��
n��=)�A��X"}m/�8/��o�I�|�_iAU�i�D�A�qjRQ�8�b"���O�D�����F�0���1���q%��`�g8��IĒ�$E0sMz�ɬ.���)�k���_��}� ���U��"���-���?��L$�3E�Ä��L$#�=9�m�X�rA�m�r�,��;�7�h�pW�]�/3��nj�#�āj���t����h�n�X�v�+[��wj�y�WG4_��B���O��C=�[� 3��I&�~��Y�`��U>Z���6�2�w��s�,�2-	S��C�~��̸�f�O���4�:����^���E׽8�_D(����Ӊ5��R�ݥ��=�JKͨ2��#���R*_L�W�2cB+P�\�a��u��L��~b-�N������m}'�� ���\��YZ�{���>(E�׎��
���� ��!Ik3���Z#q0��1l�Pk�G
z8�ɖ:�2c�&��^���ZX���Ӑq.H����B�X���A�2-��I�Կ� 

��@<���r�Z�-�EJ��	�?&!3J~�"�h/Y�q��M�O�IۘDN�~�:m�'7�SA�6[��W�t��t}����0��M.��%�a��RGE�L�ps�>K����e&�r�)RLQ��蟥�h����5��]d3u!A�ߋ���;`Ɛ?��}�y!�}[�i��p�@.�#����4R��#�ՓQ+C���%2�z'�X���d�^�qB��gȤ�d=�J��Q�N��%�ʠ��6��S�*ѕ� ��ւ:���� PN8��Z6��0���� �n\��J(:�|(>��dC���ᒟ�w{[p���#A�NMryo�4猒�!Ɍ&-Nv��W1� e�x��;��z��5��I��[7�D䄪tK��;����Z� �tK��8 �uա��e$Ndoj��*���7��#|�{���Ι��������� �3���gd�<�3kcNؼ��(�b]ݛP��-�`+ƀ�n�FP��l\�>�
at�SPX�(H�mڿx�J�<�J�H�b�'��OO!�/��半r�*�G�ΪR%�`��KBnf���A�{�5�}6-;���CSU��>yv�Y�a���c�W\9���X>����d��xZc�|�/��n��{�K��4��TJw�u��fy�l����i��*q>Hz�L�U���XG�m|~���:Hs�w{@~kʐ��"W�^v�U+ ���>-�'!?�>�	x��.�~���l+.v9_�p�=6�9�72��b8r�Ea]��N�����w2S�0"��2]<�c<�g���lPG���GYE<L�^
-��$�l<�+��k�;i��nЉ~���g �@��x�T"�u-��4�K��Z���Rzw��(�R�?�X{�Cď;pY+��g�2�[̟��V4s����Ͱ�����B`�&K�]z�����Մ���K9�!��/j-J�bq9W}���i���I���5�γ�u��c�
�Ț� h�dQj�T+��{7S���"0��{����M�J���\[��VU8~��9uK����(Q=������QY�H��Y��2�X�_nW�<�˲�}0��-�o����w�~+m�.��D��ʱ��+�(��q90<#�>�h�9�o�g��^�a�,�4��p3�'��$e�]�w�5��a��SK�2ϩ�NZg�_���!�\�V?��w�o��uſ17Jiъ�I�u1X`�gC���c��F����x����q� f�fX��w��)���<7�o�6<�� �˙�N���;�B���H����H��U��� ԰[�U�qBD�u$��yPJ�MP
���TXJ[�"�V��^����L�:�~�WvjV���t�m�*��|�Cx�S���K4+N���Gn߿���;�`��y�|L��!9��
q�EX�Qe�^*��wԜ�\�g�d,|3KP%/Z[� Mkb�&�9IG~Y�t� �}K���7X���M/n��%�P��Δ�,,���]�g�p��l��&�2��	:nI�����ޜ[�\m�a�9��!�!�'�-_�6"rO
٧ʐ�$M�9�f(�-���i(����݀���ƫp0;�v�P�M๚S�b��Po�^y�1��8M,��F�:����^��VR�g�2�,�W��t�������46�!�Zdo����C�F.�����S50*����It��l�T)+�̓iUk0����8Q�%4D}��
y����ƒ>�<_Q3�,���s��:d+��bH� ����GK��C0/Ͼ4�ʤ�� �yrfsK���	�^ڮL�+�#�zo��0�����R��CU����}��I��Noݺ
�{�ܞ6���BJa�*uu���\��9?�A��Jy��r��xʴ�}���HMߎ�f�,�@[�/�q�`��S��j4@TԄ54�v3�͝�s|�;}[A�2*�1aqG��XBdr2�ow�u���w@`,�+ �(���8 ��X�\�4{d��>��X��J���St*TD<a�����X�Q!��������kQ�Q#ù#a��A��4�t����|��qZ|cu�2�;�k �nGy�����!�s��1B�fU0��X�S,Ȇ���[����=&~�g�kNC�5�7dK���5��PEHi�+v�������,܋>bgA���d��Q�w2�ʡ0s���z�1ӽ+�n�s��T�ހ��L#h]���gt���I�����'�"|xx�Ym��TM����=m�]`E>�oЗ��D4t��7`�x�?�P��W߫,���3&<ߴ�evp�{���
?�)���f��"�'�����x�J݁���.���uɀ�πj��<.��d�V���o��j� %%��a�'̔7���[��+�8zu��ghM\�r8/��cr�����m�mA{g�L͂7��X�B���N�]��[胃��\��@��@�����×�B��d��7Y}/_63��57��?ۭo���o�,�l<��-?'Ox@m�g�n�S�
o�� �n-r�@R�/%���\��r�!Z�$�����I�ޑU�/��էu�`�s��H�Ŋ7��zl醁�&���<�ʹ촷	��CZ�~�z\�X�F�F���\t��T�A�����M0�waH��,Xt�c(������8P0M�bnz�>h�8��dQB�����	:�Ȃ$��	�:�:�6�R��6�	V����w4�I͟Go��Ro#������I���1��m5]��W����f��=��q{�� �"46[�[�~!]�O�(��fx���h���]�~d�18�lsC ��d���Z�����\��"mi�c�C��v���7��Bm �:�.p�fJ���`jE��]�S؆1����7�#���Z��1#f��7�Q�'�'XV����,�aT��u��NC�,5[+/��-b���5Ax���+��Y�5Ѱ�ￔ�H�d,f�%��8�Ԉ�6Wi?�"���r9Y|{(Z����(��V�?W)Ux��r�$7�Y�#�9�+� ��Q�f U-
@I�W�BN�J���OK�[�反q��)t��L�v2��(�w��"u�� i��;�z��$4R�Q& �]��n?.PD�ofO����e.����U�D��%I����kAPI�~���`����{��A���u��F/B��ܗ ��_��ip�r��]��vg3I���M	���R�l!B�	3ql�������P�����qs�Џ��E�$(D�1���ƅU��06:/21�@���� ��c3r��SM�n%Qjx���,��,R��ȎҖ�%�n'�`X?⟻ȝw;�©#��atޑR]�;�����I)ƭ	���VGs��A:�#^L>n���V�E��u��CO� *�5xF�0��\ZĒǶ�ɻ����z��4]��3�b�A��WB������p�t� ��8՘!�em�T��Z�s We!��6��Lnu�=�a���z0�4;��!�wp��N�nz���>zҐ�U�_qhJ{[��1�?M�J�݂O�,i���3�0S�(s��H��(��s{�����x���E��rE��!q�� K��rb&�?�8�� �>.�'5��['OJ��Ľ��"������aqF�I�M�7dWx�!�A?�0���A��K�^g���_�,,�qڛ1��Ak�"��4��5�)=�oW�s��C���<�A��A]��z S����XI[�}�
x�y}���`� `���3��
��:<<�e%�|�C ��Y�e?��=)�TK��"r�ę�$d���-ֵۙ���D�ج�
O1}Ca�q����.���v�36�,X<>�C�[o�z�7
�Q���A«|.��JDr��$��]>�ᗨ!�[ScR�PJ��@�?��_��g��)�u�z�����B�g�g�tp���I^�u���1��Tn�֝zS��/��M>%��/t����/E�M���qhF,N�Ǻ�D�J��0�m��|�����y������R� S�z��+��+2�]�ԔvJb��˽��	[�<�ql/��۬"g�\����!~�1������e���Eטa`�+X��I���=H��0��F�|��!�"��q|�J^��T�/D<��P���%Z���6F��u��A�� �d7�r��0XZ�bϓgTy�ժ�f:�w,>X��U��D�nm�Q<m�"�$p�9��TC���z�4*4�dSqtS+�8*�Ar|F��95���{����2Rx��2c�{'U3��f�t.z$�C���Ģ�+9��^�_�|W޼>���X�\X�����'@�6�=浟��r�iH�6�u��O���41�7g��Ik۫}�3��S�JԀ4ʗ�j�����Ȣg��YO��㲳�YQ���%��5��n����`a�z�����V
��B�R"����SN�e'0N<�5��JQQw�F�9��mRyX	�e��*����ܑV;�s�9q�x�p�$Ņl��V�z��M��z��b���W�U��ǰ����2A?t�r�ڡ���͌Mt��x��l�LJ	fI2�iLZЬ���+���4Sb)5LS,�0�k.�S;O	eUr�/P�pZ�kG�[H�~jcEU{"|K���A�1)k�����+v����8ɾ��j�h��7vC��R�o���֒BX��/��y��6iy�S��tV�>:t�j����5�oWs^S���G

_	�-TJ�CWV�UTM_��0�%ҩ���{$b�i���K&b�͂��6me�B �L�s���6��a2�Z??#XԼ�'�@�\7�Ke�E�����ڸ����$;���R5	1:���]p��j��A2A.3�~��,:D�N�J��/�]k{����fŸ�s������y������x�W@����>д���o,��m
�/��a��Uh���wx�!(R��c�
���s/�
��>�������?�@&�᳐>pb�j8��������I�G�]���L�ܤJ���*m�9H�8`�5�Da/]Np5�+1�����m�SUu1�X�|����G]�dP��/�HaMwd���B2�WT��8�ǌysQd\�e���}>���vWoӏP1��A*a�O|�����v[K~�GrG���a	ܩ�[��J]_Y�3������0kU-��)���2�%����ŮX�x���q����8��8��k���Y�@�����w��顲6 e��N�N��$Z�r}:�E��޳i��h�����>�y&��d�i��Tt���M{\1<�՘:`�����x�8��}�k�[���+� �sM_\�ؐ����~�,?-i��/�dɜH.-�{�5S���4��/ZI�·�U�bVu��Vv)�e/`���I$�B7>��|Jh`8Ԑ.ڣ'�$�r�N�wʑ���%��d=:����M�TЛ(��Q��tJ��I ��T6̟�g'ș�S�&��bB�b�8����fy����qY�s6[A�.W��SI���*��4żV�ye)H���Mn|N���\�5��eGLJd�����e;�$zpX�!JuC�,,������M��3�����ʍCO��YU_���B��
��M�ޕǱ��tS�ӊ&�&��l�wy��i",D���fd��=�!$����d�u�e�yɶ\����
� �P|��QW��I��ٍT�R?	2jQ�e1��x��M��ܶ���	K,�]�.�K�Q�jK1q�vv���r \���'�J�rR�N�ի:���2 n����3�.�),O%"�D��P�0�!'�����ErGkw��C�l�Mv��]�YXn�/ݼ�zc1�L@a�����D��a
`��b*e�VEփ�p�����Ё��P�w ���@减�7��HXp�/�Ԗ������OڴC� ߙY�ÿ����҇f}k���&8g"�,��w�I�KSI�XP��	t5�ʉ��w峰Gj#������W�kA���l���ݩ�Ga�4U�#�ֶ���YR|);���V��K�D��E��B�vy!$E:0�a`�K�������fj�b���SөOU�� Ie6�*�3�ǵq\�t&M���X����Ϙ��2i�!G
@�X�[��TS��*&����a�a[�77lF���:�&���*��l:�|<�{�3�z�M��hV��kG�l��I�¹���I:/���oU|%�7���z*���5醴a�j�T
;������;���=��И����\6)$�0{�T��X/gG�Țy��	y`s|�i7�x����Nyߌ��1ͮ�z�s�4��I�@��HiA�������] `|��*��x��(W���\��yY��QJ׀&6��j��4ID�]�G�i-+��t-(�
�E�p�^|��f�0~fB1�g�q�Kn5Kkio�8���,Y֬������2RLǫ��I��)���C��N��k�s��C�37_l�cq��ނ�� ��er�67򾪲��m�ֽ�ٌ���K��b��$U������\����JRUxsZ�j$�5�x�=_�J�U[�t5��0nR��%Ҡ+���2`C�%�
n���7_M��׸��-��\��K"���㖫�#�/cE:`�[���f����J�����RQ�؅���#&����{ԵR��p����]i.\�k-E�OZ���)��]��ЦՑ7��v�����C��x���-:4PC��'��AC��)D�[�4j[�y��psn����m�K���HC���QL�$ ��m������D��=�z?����!>��b�`.6ٻLW%�t_F��b�b���;ן�^<�RT��2�G�8n\hӌ'��8��p�� �%8Ĳק;�7�'�C(�|Ч-�;b|��al��O^���ѳJ�)r^�!;>�$|>L�t*V�]�b��k*!ln�Pp��\z����dI�� �Qy+y�Kψ;�{Ƹ5w$R-nҨ)�nX.7���������Z,�ޒA/=�n떲�2�< 1�:�^�*����ր�!;�2٦�efb0\>S��n������6�h�W��N���o6
b|m�u#�]�QnE��X�A�Y�Ċ�sϬqd�c�kа^��@`�Pن(1�Fܽ�M�W�)��|�gkf��a���g�pT|߆K�L��8$�Y4�iu��`��s�&X<���$M|*�~9�%A �*���y~t�[+H=2�8+�K2:�Ɖ��œ-�K5)b{y�"����umb��M&w��>4 ��!���Wǁ���Շ�����\������R�7���"�8�s�#( V0Ю`�]E3�i�D_Ne�9��
��C����R�a��l���1���fY`{R�oɇS�/ 7�0H�\��q�#?���#ɡ����� K�����ȢʞN�T7޲��77gO�$l��r��Ұ��YA�uﰴ�ţ�!sĀۚ�=e?�qN�dᴳ�	c�S����N�om͏b� Ֆ�';�z�"F^)��_("d���0g�uR8�������7���wFqȊ"{yW����mw�b��0y/Q%��Qʸ)�����P����u��&��� њ�6_�� w�>�Z�8�h�]���i�xm�yQ�I��Χ��^�V�|��l<5^��Y,~|~W�g�����!z��.x�����Р Ӡ��=���<?���M����-/^W@Cj��'�n0��cu�����&�����A`_}i�-�iqȠ���N!J��-�ն�+�8`�����NZD�����10;��B�+�3F�Bj���[��E�ʰ�Nx���A��&�`�g����b�0@xe���W���rAqp{
�ƾ^��ŚJ�hv����r�|Wf1˹ޱX�A�8�s�� �8�ԟ4U3L�Qo��=~
�8�_S{�ly���]��,=��D��J0,��,d��i�����.<��M���J`i��>}���$6~�J��RLf	�#�`0�_VQ,2 (�G���)]��yfi���d��c�O�Ӂ�9�Q�to�m�d���| ���x���:&b;��B&��r{�<!} ���G݂�����Sz>�ǔ�g��9�&r��6Mn���\�{Cok��o#P�FRӞo��cP�'���\�t)l��n~�& �/��E��Z��g�D�z{q�׷_���isH�DM�%��>_���Yn�[B@@���G�&	Ekqs+�
��ZU��b���Q'5;6�L60B�w��X[���2����+1?6�k�y}��9F�'�p5i�8�`T�sUI���������SoZ�q*hw�Y�Th�l�θbm0w?o�B��T����$�A�%ie��Z���ȖD������RF�hwNmu���;U�RɅ�_1V�G q㚫;�wEV�&-��=�ꈥ!�����O�Ы�K&ظC22}�IEe6��L��
Q���f�4�hIU�=v���YZ�d�8�$��65-�?��Z�������D�տ�-�M�\��@�-��v�j��L�O�f7� u�y0'{�q|ڦoeH5N+����[�@��a�~��$^C���Cc�|/U�D�-�E�h������"���K�Q����ۗ[
�P�����JB���*��rA�~;X�}Ku�N���P�+:�t���)yX��٭�y�<���d`!WP5i0�p��?�������뉍~zc^?�u,'A�r}���,�Eí'�݅�j�_̸�K�O+t�
��	��i�s��f�r�M�_z�(�<�m�/��LS��y���9��X9~���SI��F�K��y}�+�Yd�����0P���b�*ұ��t���eQ�a�ٹ�._qu���5�� [���q�^���l߱q*��%�x�o�r�%')r�����"C��]�G!�H�<�k�Ih{�JǲKZF�fm�O	mr�U�+M��!\ʫGp7��ķ( �����5.liL���v�Tזچ?MtC��$η4�5����ư����*���xjv�:w5m�9�/��V���$��ο�Xw��`���gE��	�V+r���
FE1�� r����Yg����>�>T�����DZ�3�c�q�Rw�,U��� �U1ۤ��ibO�Kf~_?Ʀ�J�!{;aD9�K���,ZD+<M�������Ђ�	��[�ﺲ>̍��-e;�����e�&�~�P�kASĚ�gLdL��%&�m�4�F�aS��||w�Cr���7ZY���%��X�h4LE���d�����5VG�e�̃��"`!/�`�L-9��4@��q��IAp��v7����5('��jh��/�-��[��C)�����S���ݢH���=� k���9�3L���J���s���:�o�!o9��<��f�:�J�g��&�<����6ʜK^�4T�:��L/$�G��(��%��$S�W}�M���`��qOy���f�y�h²��8��5�6z�\��jU��|��I>F�7�W���XS��|g��F�c0Ĭ�/&(8r6��F�e�C9:7��' 6j�B<�Fy[�B�YVR���l
��V�֎y
�J�8ι6���x���W�rff��t�ݤ�sI�Ʒ#��r�
w�\P����I���&�5'�㠍�ڪ"��k�����3�2���r��|�����.���T!e66�����&����g�XLFD����%F=��?���*��5:��z>|\m����s\���_�j��hQ�_j��l.��B��������$�xTj�.F_t~�Bt�NDҊ,j2�����i��+cB��-�)/�0]���v�U�ze�~}���d��V��ZOr`�Yn!���0_zk{�����Iw<�b��2Qkl��u/a�5}+(P�jui���/՛�k�%�΢?���ʯ��4�)p⤆n@�����w�)�Ee���G%�cS� ;�6=�G�����������kju�x��3%�^�v��%̵�v�=LK��7f��p�D�D`@-4�/.�M���">�T5��e���X �:#���U�G�i�D0\v!5JQʰ_�����Ugwy�m��	�(�/�ړ}�H��+͉�@� ��B'���=��� ��F$��^�hf��a~
@�z�I8�i��#J��~DF--����O���i5�)�Q���BWĭE�l �f�WarΝ�N�P�Z	��؛U-�f��B�Àz�_�T���_�9N\-����=��X�����㾜�5�0��?����)���J}$$�(0��r�{�y���Ӂ�V�o��&�d�����J�I �z�H����.�ͅ����?�k)�DU�*<�;�%/��5S���G�(�]���4Y�r�� ��y�,�}]�h����e�(����9��p�D�x��P�;al���=c�Q��/	6ž�>4�F�/��7:��~p�X����1���[�v�^�*p�!)�#�P>2*1´�9����b��Uv2}�IrV�4�|���U�4g7�ޘ.����H�\�e@���T\��@ќ��7�ja;3"z�1�H��V+��EV���[7����`e\�\������4��'5CξE�׿P�3�`Q�i��M��	�P'��nr���,���T�@�U��C�c�q��b�d��
ә���bڈ
�f��L�a8�\(O`GB��L�>�UW���.x�\�Ks�|[��p�m� 4mwj!�j�N���d�'լ�p�ݸ��x���๘O�
���(@�1�x���Jm�r���lG���=Rж�.N�☸�Z�v��#�N�&x�����2�0��"N`;n���w�i�^_�z��Լ�A��ToZW��5L��gTԑ�ZMTTm�׹��QִԐ��5�d�5{QK����S���Pٲ͜��q��h���\�_���n��f�x�+���:��7�׫�l���Ki7y�)�^&j"�z��Z�w:x)KF �KX�"�RB1i
�Z8�;>k'���v�-�v���|�Ԃ5��ݳi��~VR9�H5j�x���iV:yA/�-'��$�8�U��^�������B��Re�(YI�������Ń�P���D�Ӌ�c��.�챩��I��� Ps��}����|����wl0�̓�sp�J�g�����}A�����ԫ��X��!G����֑���:ϣ���u5<1wW	�=ܫޫ@ǖ�D,�������{�i`��Z��;	Ce7�9$R���Vb	="U����*(���9�������@I��Ej���:2����9���l3[�tF��VU�a��|~Oޑ�</Z�e<���EygR 3���S���]�e��0v���^�l���k�al�h:�H���]��z"����@�;���O���@�}������~�A�+��K/���M�:��R��ĺ���D��Y�@�{`;��d\!KT3~�As���oqۨm�|:c�6�*W�x�A�n�rc��8��������D�~�&�A l����;�ڳ��ћMkV,���[Vm�������ER���M6�ԣ�!�5T=&������d�u��¤�v*O��ZP���j�睴B}�9��O�FY�'��f!ܼx�'@����K��v"�w����6s����'VEܐ�}i
p��I�I��v���s岐���<��'ި�m��8���M��Ӑ����T���s��ip�`$��O0����#p��'�/��O�C
��o��(��`+��=QO��෾t���.�D�7Mnzi�/�mld+L�tr���Cp0G�]�f�doS�Q���|.��]{��)�%�P��i��Ǌ17��pO[��32�Q8����#ʠx��$L����;�-���"��g����?&��TV�j�{��? "���&5�3¢��oDd����0�@��8ܸ?{�V��as�9�E�I��p����J�I�Ņt���Fc�d&vk�\,֏�	`�q5pJ���k�T�r�������j�+��[����ӫ��2��	&!^�3���p��:�1]�]b0����^����Øs�d�Ҧ�x��=�y6�Ef�ʓ"}�]��/!:��a&�3r�F��~�(-�ȣD N�*��-˴��}ўqL|�����$g*/Pyo*i�N�!���*7��MM�����$�,5�ܥ��7���(��:���6n�2����PK�Z�:+S���	+����a��4(0� ���E��XUc��5�4��ڡLF�@̃Q�eغx�A:���b�n�p��;_,"�ϯrJ� _��I���9 �Mp���OM!;����)�iB%R=鯺�E�/PF�����F8	F�y�2:�O+d����&�����F�5�����`_�3�]N�:�f/���+��BJ��[�T߄k@��mˌ��Uu96v-���7^d��`ԫ��}
����F��9"��������]��TF��	��TA BvfW8k�o���QAa��-�!5c�0}��1�m��O�&�� �DS�r=�a�I�4��6���E�.�W�ͯ���AM/}�Zv��T%��s�[tPL����sid�=�qd���e\�)�e��:�ΐ��}4���,�)j"����S��'}����rE%���'j������Xf5R͏�=��#�WIo��g���Uߴ�U�M�ʳ�f%�l#%Iz(��kT)%T��������>�����K(e�
*��I�AlQ�{�R����X��cpla�i��-�jKT��V��ff<�`H0g�W}�R��X��I������ew���_�/��k�P�]���>J;k��tBδ���2t(��h64P�v����|YX�Th�W?��,s)�/'-CF�ȧ'{ E��@�{�L&�Y*����FG�U~-����y�8]U���E�ǎK����Y2�a΃��}��>uM��l�
��<��P���!O�Q���.�Q#\@�s�^}h�"D���u��C�'z��.�I�^�I�y�l�ر��6M��/z�w{q��B�ͫ�NA
�(���`�{7�Q��֘����A���G��^I�)�˞��,�_��6�${��tLxO�+������w���͸׫c¢�� f`�b5	��z��������v�%��*��'e�Ҧ��@��AZҿ�m�.;�9�n-�y�ɿs�lK��J|���l��2�a'�lF�#{�2�A@�ABd�Է��:��d�b<Y�O���Mg<�MZ9՗g���=��
G���pM��DA��%��G�p�H(�l�:g�����{��-A�!������]��m��哢tn1��
��|So�X��k`Y�n�c�F��	2�SX~b��lm���Yϒ8| ���	=�d!�b[$	�1��,JzY��?�+�3��Af�E�{4'k[ ��'o�"��#&���mqMI�@q�`�¢�v��A@�7��7����ۦ4fo]�B ���Ϙ��`b��K��e��i��l�u]̱����iΉ+hl������4H���m��\	@�[^)R���	�������s��ܫ[�&�'y!�NtN`�RE���c�+?>�sB.�c>(��q��Q���:�8��+Z�� W�r~_\�E��OX�@zDx��Ӥ�&�˥!^5��9*\Ƃ��Ҋ ����̷��?"9�qM�p��0��3
'�F���1K�~��l!�����$x�*j}[�H�lXW� �fB���C����:����q��=�0�Xz�Ao�����%��@����wI�56��;i�_4p���?��V�,Iȃ="��Vf�C;����*k���*�lm�llpRK��d��ﾫ8:g���F��\����D*��<N�)}�ڳ_�bo0N���d�	c* ���r���+�Ǎ���?c O���hǸP��L!�"��ax��'�I֑(U���Q�����B1�ZUQ����j��}���% 9@f�����]M�����#�[E���8G���!Q���#��%�^�)W�}dA�����V��J�<����m�HקDb��Vk��?>r'Ñu���'�*�Ρ��3�b�`�N6ID��:d�ᬄ���nf��R��7�V���.�~���fP	�v�̽b����,�z�I	;_		��Ȗ=��=���&���H������*���|�n9JŞ��YI��\8%���h�>�{�4�H�
P(�U��7�_��\e��v�H���/N0(��j�ΡxR�I0���	Oj����($d����Tb����4�.�w�-��7���=��kr��m���F$�ᤏ�E���FN�^:��iX�+�q�����=O�^i��:#玟��~o\���*B�Rؿ9�U�/д.�*,q��R���>�?7���!e�G�ոo{��`JZe��B>��yFE.r��D4���ѷ+���D��k�c�B	���ѪS��e�a�Փ��̰V��RcC9~�_��i����X��k�0P�ӧ�f8�����k~!Z��uq�n�>j�ud��B&�\ ;��߼��7+����߳��5�����C������N�q*�'9>>ߴg����9�_$� dao��QJu�e�MY
S���@��c}*�n(+�������H^d�`�i�����eMM�EA�	�d�\9���o<��L�?Pբj��g��F�({x7�Σ5���z���p��-��h��i�|ᅩA�=����m�nT��(@[��\�(�i�霜�k��V�����w�H�[,
���*�COc���{	ρ,gz�ԑZ�	���/x�D�SGrٯ�Q%���;�ZɼAh��R�_����H���E tl ��M�\�ݭ!_3�O"
:���Eʉ}�)C1�Wwm>	a�
$��p��p��GT��ן7�X��4SH��ሠ�(�E���w&�A:̸�o�u��/(��M����v�-�*>i�8rH�&��h֨ؿ%�M�v�� �܆hWZ����b䊑�M�v�O���Ж�m�F����AxnX�,�\Q���B���%��o7I7�6>�Α��ms9�n����W�X�n*p[_�8fh{#%������>=J#{����e�/k��������l�u��Ɲ�Cj�H�ks����5���g7;��,}g��O���d��9����j�����H�hLF
-�x�H�!�)����5�d��{?R$O���*@</@@�O6�Z<�Z���q��`�����Q�'|�����
�y��-0R�ibX��P2_��j�������RMb�>��Ϥ^ԵDK	.lE�)f���'9��dm�����e��:��ϴ�q Y�U�Nȱ��/-?FX�-��򑦝n�BO���0�2яܱ"���5t�C��F9�_�s��˺'���TDxL)�V��X�@�@gi���b��}{�~�hn�e!�����F8��BCϵF��+E+��mjO8z,%k+[�#�s��M�#��*k�Z���>����q�ث_�@�w(��x;=�um�����5���9>��[;�#�hF��)AŸr��b�3��,a�c_�%���f0�/2R����!��ʙ���-�F��}xG�U詨�D�[���ţ�b�v�.� ��Cu7�W�L���ik�"|�\qL�z�lm|�bJ��$^~.7I�O�+�	���ٌ�@<�(`Æ��qᦷ��i��`�/�����hۋ٦E+S��1�����o}D�=��UʏNE�l��9�� ����(�5��d�sv��EȠ���\�����#�T��H4������w��k2"����4�RV��T{''���\�Y3�gU�#p�������I&xu�����'��'��WT��!5���f98�x|�Ô�!3я�횵
�-d�����B�jS�`������v��᧯� |Y�F����ia�V֣�/k���Сj~�۲�l����QI����i���D������7;p�����k�🞧�����8�����ULpY�(�f㲝�j�K�ڦrd,��7$�Ur5�O����������9�1�K�Lyp�o嵞h����i��d���3�ܖw�i�Mw��J�hF�]6�5�?��$a��&h���
#;����1�&��	wdc��LAH��MI��]��}�+�~<aH�!��V��]��۪�C��e�EF]#:[�	#1U�	�Qd��kǷJ�M��vB�fz4l{���mC,�9�+?u.�Z$i�6!��O?��HAZ�Վȼ6�v�|J�-��\;LF|�17�`c.���N�����¦h��`�qx2=��+`����!N�ƘZ0�$`��=�G�,c�YHr2�"������z|�İF�H(�ܦ����!j�|Ź
����BޚOk��)�l'���R?�*@�]�y7v�{��e����??��^i,��@�)��r��F���XT�I���DǨ����k��4{�LuY�R��6#5R���VF���+Tn���9�&ot���31�G���ĥ�q:v�:�"Nj4�n�6_?�����R&-�w�ƲhL�RR���!���;�Gpjh2�SK�n�9浐Cp�k%�"d�'����C۬�̦J8;��p��->w�:�)�l O�]*�S��Y�E5`��D')��dU�צ���+��:��(�.��pXdH�JB�	Gb��A��p�m
�&`��yz��	���`�Q���
��0-�@���C��o�,�ĥ2��&��*�nI�V�v��\��sRYV܊��GD�u��x�BY�O_q�����@���/�y=�Y��EMx#�B�S��Q�M���_p�э�J;6����T��� �r��C��5eL,=��9����G�u��-�ك������y�i�K�\���Z�z�01�����������:#���ۭ�����ʣ��Kd�A��/p�i�;�d�':~`�!�g�_TW^=[�����Qd��)8�>���#�"#�3
�s賋7/�	`G��H<\�iiy�V�7��Fr¶Jގ�$SR��&�,O��?Wh�֍T�ڟ��&P��$c�����!/��.�at/`�K�y1�2EG$�;�X�s	�Q偲H�b��nYS%9qYbϺ�ܴ��>�	��;�k0�ʿ�1��u|J.@�]dg�©N������GV/P������Q�:���R�C`];��]�kר�$��;+kB׀cH��3c�f�.<T�3��U��5T�c9��y�O('(��w���:�S`�,���3#��A��$��&�(x=�T��3̡hwh���n-���������.�����a�#��^�g�=�����f@e��N�xe���a$���������ꞁVr��O�I025�Q����WK�J�A*�e�$��^�d�����[Y�m���o���k���?h���/�1��.�H�g��SI�_�2����y��FW�=��=O7QN�m��I7������/�v���]���	�ֹ��:��X
���Ӄ��dB�)�߇*6�w�z4��=����H�T���T�3�P5��!_9�7�uӲ����S�s{l3(�(f�["7�S�-J~Q@� �"p=jD" ��9��5V��2�cMѲxKwN���=3rq�x{&����!�wϥH�'���J �Ŧ��H�������ZCn���y��D�Y�{HQ�*8N8��@X2r��Rڐ���iٜ�����$Klt��}���z{μ�b3�:��j'|��	0Gvp�!tC<ԍZ0�&���.��a��^�|Ⅽ�+�H�=�C��lPٚ�؇P�&Z}j��]�-�����C��lA��ha��?�J,��1jF���0��(|{��m u��sIA��] �T�Q��UΡ�'�_�K^�c���R����=�]��>O%��*J�^ț�e��
?�~E��Dְk�]�S������$���75 "K�2	��{�5e��a>���p�V���	�fF��ϻ��q�DLk?q,X��`��z�GIr�)��эj��(v�eߪ#�ʊ�lZ�4�k��#s�	0z�����T��"Z�u��f���#8����qԿ�`����	D�o�(�v�#�l��}�G���#YA�ʪe/�~��5:���ɳ@��:}H�#;/9�a?���4�b?��K�N!�6:�ʹ�R�}N�a	Ύ���סp,�⠐vj�+��]p�#r]���GC������/h�v�X�������^c6�w`�"I�?��4��$�smG��9%r��n��R
c�D&����ęk����tMp	|�|��w$��kaL~�r�23Z�}s5��?�@��mߦ�$�#^�8�d���έ�t�#�C���N3�)o��C���8!F`ֵ���NU�������H���R�٢r����`�M!}�e���9��/9�]����f��`9�ܠ$���N�@gnV��V�����*��^k
ݑ�s_����LA)*�C���c���r���;��ِ��t��cz�7D(Y)�wM����T\AAYr��+]���DY�~�$��&�gG��"�;E�7$#���M�5^������0��� ��6��tǐ��:�t�:^���x��X�n�ڃ��^�����P'�|�ˋ��T��OB�'�f?̼+{k����՚}���h6������Ħs��?�A��~bqkk4��B�O�V��?y���!�E���@&�{�k�T�z�ol�ErAn�1-9$��.Ax��������}�ꍮC�rŷD�1J<=}(��l�,#^�2j��s������~�O�lȦ�ov]��
Y(��]ن�Z����u�h.�;b���y&���*��	ewвE�����w�&����-N?5s�u��E�1#��J�@�>��A:�x���@��cx!��������W��U]�H'���h):�P�����;��A��D��.}��h�K��6o�JB�T�I���"�\|b{V�Y���sd��} �q�X0�rD��0"��K�S�Q]C1j_c^�܄��3�#i�oK�Q+g�U?�3rڸJ�<�h���S'DuYHH�l9���I�h\M>z�RX�70R�]P�|�ɥV� �
�?ӌ��!"��o����)J
3z"�LM�Wϙ��Ѩ�+8�` ���B�O���=[0��0BZ1}���^,ɿ��O�gLEO�?��>=���\��pN�N ��i���{B�H���mE��Bp�+���R��0���Hr���݊�������;*�����g5	��i�&����1Ƙ�o���Zm4�8�TS�h(�Ȥ9�TH������?����WB�qe�����3z�6��Ӿ�
���	��-���<&)	�Kr'��]`
�{�Ë��@sw���xa���Z��-��;�2���G��>iwd�����g���oS��?��^% �#��m�<�Гa7A[8����h���G������Н�a�X�,Kĺ{bd�Dn������k9��ݡA6�e���M�t8-���>Nd�=:;���w��U���\��r{ۓ�v㑩����Ջ�����gܵ�q��S��fT�NO�㖉�B�|=ic-�Z-#��B1��a�/�D�%r�4�!]��L41�A���� �A�}JjN[�{hd��bZ^�a���'O�?Q���CK�	�)k��a���i�fI�l�i��N$ګV�>�g�ć[�_��huHs�5^:o��0�8z�no������yvq�5�ߖ8l�Te���1=4���K+�;��Rj�	`:��$H�i�5"��m�铍���bedp;z���KyoNl5Fr��ץ�������\�~��EOM��*6��9d]��E	4~�@�+��뺪<M�^3cC1�nȔ�n;�*۬�X{��Űm��h}�+Pw�^j���,L�1��廝5Ѫ[UcAO���p(lڠ�
���ص1&����<I�g�V�)�4ߐz�x��~L?6�PG��*���ۿ��˧I5���O�"A"�B��P�I�)<;���<��2��9h-���ԣM�%س��M^)�Uw�U�F�S�{c��26��w�����N���xx�w]����yQ�
��p�Ra�%����VkX-�y�;��P�c� l����6�:s�1�v���<T�~�,G������J����~{o$@��*�����ͥzE̅ e
|�\%[��kΒVGlN�;�6�f�=
])���=RDf�u>���X��1@��4kdx�7�r6Ei��]�>	�K���Ni�	,.������[��S(�����1k�:�ܘR36����������XL��y�a��R� �)�Nc���9u�s���	��	���1��/[�@�@͕�ʐb1��mF�n<��uH`��ɰ����蚻�2*c��L�g:�O_8Y�XA��t^q�/���2gJx��r�9v���d����q_�\R&�$�[�%�גqc�.ș���+�e�ہ����G��{l�����`���R#S\�:���tc��S �kYv����!�3\�T�-9APVu]��|O�/��8V�����S�̃΢���e_:���zo�M�5�\q��Q�1���敓�sl;�~���J%5G�����l�{�4	�;���@Ryr�9�RI��|q�W?��m{���eY��X%y��5�B�p�j����/(V~���F����o�:��R8�s���<��8�@5���@�d�ް&<�Dv#O�j�]�n����:ܴ;��ͮ޲�TV��85:�ɧ���C�:Zs�%8�AA�bu�\�&���>��كR��s��.�<�I����O@�DI/aB�N���@����>0Fȗ=	]���o�>�FA(�����鲸���jrb�3��y]�]G���ۣ�R$�	���PVIM��p�0vT�;�/q��)�̠CP�n�ar掂�\��rq���l�߁�*�o�>�q!Z,!A޲�Й �
�s+���*� R�х�(�Pg
E�-@���
.����GO��v� �*WZaW�UYC]ɻ�T�<�҈��t<����0������q/��K�V(pIoFɊH�{)�U=E�F�gp� ��j5똗3����yg�}�k}����^���i���9�o�S9Y�ր�{jwI����R�Τ�!����L����{cgB((k��+N��$m�	
�3�3M.�����+�,ٵ���_�V9��ù�$�C�o�?^�(�v$�d	�d��p\ތ��+k�k
N�J�k,bM~�+��a�^Aۼ��y�I��jl�.w`����.Q�37R��KR�7�x��"U,;�ΐ���u�!U�}X�uoߏq��K1�73�5&�`��L�����N���Ϥ̻p��ʢs�,�{����>��;U���BX�	�a'ўo�l�t捷�i�莻�X��p��7$VlE��z���D���b{�|�Q��Mΐӝ��R�.��Z�	�$9F�����
�������>�����0��b���?��bq� e��:�( f�U���һ/]��
;�dH��|��������O�v���#F���UcP��,q�Y�][�b��p��y���<�I@CsՔ�z�v�Q-w���]P���0�A���9��K���~��J[�w�>H�_���jS�ǻNA?j�6:����ɦ�j}�r�X���T�2�T��%n>����ɪF���§��(��mn���T�Y�%��[�u�?�,/�`�q����&���\���܌�_0��<�l�P�����Mm��B�B]>1��)��_��Z��c��U�ց闶?�|�*'Dn�%�6��B��p�:A�������\,	�V��S��b*�|��7W�Vr\J�aU�(6.)��b����р�PVV�V���v֡V�oP&*�Q]w����-�9��[����pRd�;��bo�-�ZB��~����l�1��=+nc2Rc.Jڃ,���-dA�)R���$�T�sh�?d�e�����(�X6�o/�m+lIIML���(�5p��]t`BB����H��pn>�j��f!+#��8�h�w�5QR����>��h�ܘdbb�\���@���Gj�n%X�<��/�G�9H0"�kFp��jX�M����]e�}�����t�?�����sK���=�
�������}h��t�2��N��;�v�.���i����09|�6-WJ+9!
�`E�~#���	,_��9�GV��lD�e|W[;9�w���>"%]�p���]�b��C�|�=O�q~�r|�/U8F�?H)���B�q��,����r�F����V*�MLPhJ�'�!DZ�J{�_=Wa�އM
Y;���D�ޗ���u�CHf83�1s1$J�̂��L��Pi�_n�fgXp+��x�����j�.�����Y� ��+������\���)BQ���f�{.m�U8�S
_��]q����N�nUI�њIpA��S�f��A݉�|��}T�ɿ�}��U���ӝ�)hM���� i�b�s�yK���x������g�8�I��<���x$`Ϫ'j���F�I�-�(�|��B��Pd��~��%�\�<Hx<�#N'�� ��{���T�t	6�,���H�W>:\(,g�"z^,2FoB�F�c���o0����a�0�@r�Ɵ	ʽ�(�/��z��1�a�7`��*��a���C���{��O�3��gՃ�/�CKC�Q��M|����S-�
$�r�mu��pJ���7���S{B%U�й�©p��9�+�bsIQĳ��"B����_�Hp���5�d(��\4i�!:�:�8{���X]=dsL��k��x�6č!�fnK�D=T��$r�f}4�����{+��� ׌��}�u�h��&�E�����u���|�'�+zs�%�_��QL�<4]��K4R���E��2R�U]��L�yt�2@ܩ�`��ljTk����������کN0�@� �J�"��4����OSS�=��
�o�I����Nf���3k*k�=�h��>QI-���	����y���� ����[�ڔ�I��E�_ϊ�����UV):N$�B�!����4��[�����Bo;C96Oþ:4] �"2	S!u�=��y~��=U4e�*vh�E����b0���y���В\R���{�����3�Uk�ԺW�����B#�r��ft����?(����)�jc\�'�xef�A�:Ⱥ �(5�81z��7�=�6e����X>NT�m�YAS-���6ih�#�Ag2k�7�H,�kf���:�-|4A���.�� ��H��i�5/k����B��#d �f'	�9�2���;w4�ԓ���y����X�H@�v���_ҡ�%ɐ_�ƃ-f�3�5�����l��,�!�; �`�I��Y��>d�w3����4 ��yCx�=�9�VS��ޛC#�Nl���+�Q��͖ WhBNZ�\KP����c�.'Gï_t��1ՏQ�̝��byO =�d�e)�tx4"�IΔ<;H���Lo��4$g9V>`��+�*a�'K��Og��~�uR��|!L�9��::���
I"�O!������=_�.��� ��(ј�	��<9�3)�\��#e�����L�9�z�Y]P���p��Jb������dDK-`����z��Fn	9���f_h�n}�}.�hn�;(����\U��I�Дz�r��1�$9%`��&d��I���y��˚��o��sB�7R��u����X�B(o��G��_�V�:2v9�.���y�O6�S�d�h�G�P�K���wع�_�]�{@ѵ�p���4UBV2���'@h�TSJ�/1f��{%$b�y��4��|�������Z��
�P3v(0.-W��Nn�epn�=:��&���6���r�F�b�G�s����*s��ώ ���ii��51�pr�H�Y;&o��E<�,y����H_]�rS�t��Ƿ���X�8f�.&z{OTp8��Oo�g��M�d���؛\��|�ƽZ�#ٸ�u�)D�@4�����g"�z���{�v��S�Ǳ�"}nS��rԊ�*�>�{9�c&�'�&����ˑ7���5�0l,�#y5� %P	Wjw��1}BY�_~��L'�_ݳ!���L1n����0�դ�p؋�"�@)���=���N'�E�ʓRU��@M�1t��y0��79iJ� � �m2h
���{^uȀZ���i��J�6�w�Gl���f���A#^�uH�wq�x(� ���З�w��ĚG�3W"�����3��	�K��-[�+N}3SF�A�<�
7��<r�Vv��C�����|���a�%��m��� ���]	y�*i�MO�'V�k��n�?'����I�1'y��1�u�5[l+��rҥ�ؐ���)Y̭b���5<\r2��;�Oy��B�M�W��LxM+8~�ټmF�����
�OǞc��Y�����g�P�8%�{Cv��.��]e�T\���YB��!=�K�"^4�/�Q��W{��6��������n8��V�o�Gx�_�Oy<Ww��zB~;�Ar�^*n���p�����g�Ԙ�8$�z���:1��;���#Iߋ�#Q�0�x����y��h�<ˋ��<�5�d^�s�������XT3��� fA2V��)� ��[�W#��,&�Xrm�Hq��p\�kKi:�������,L��0uX�0T23l���醕T�1��N��� nm)R�e��{�C�5"�yl��@�-�_w�D��g��9摛�1ӳt����* M[�'���(���`_�e|�q��f�� �9sV�h��$����r�s����gM�	/0�U��^��#����9׃�*l�2�� �Sk�,b�L(#zSw���I�+-��"��%2�w�۹2i!bUV)�Z� ��}����F�T6�?4�5e�V^L]N�S�<�ܿ&iBJgm4"�G���Cb=l԰�>�#Y#hT#�񋍩:���Z	�����_���d�d�1;��K�ָq�f�A�!�{���f�	�[D��i�7ϩvN��L+|�ڬS�15x���g�C���t+�u�u`�ͫm&Q�B�|�v�t�~�S��Ui�w�i����zq��A!R�8	:�Z/F��"v��L'C ��Iq�I�U��=�+)?�P�|r��h���,���h��R�yP'.�x�g��d���4�q�K_�@�2`�m�)3L�hF�⢫��+Tu@��J���Q��!&}}�X��#��<�],�̂B��un��=a��^��^/�F[���~��x8]`lq"	%ћ|�f"����o�Z�r�2d%);~ڈ�e�j��`���o�n�BMvX��/�xk3vZm wH���7]�x�ٖQ�̈́��e���HP+)�xQA�1]�=yꞆ�����m~�������p�E���ч�E��4OٱEQ��.��OrЌ�� 3VR��Gm^�YX��H=��Y��Y;���ЎPC���/5�լ�p.�Tn�����|��~��;��u:�&���T��a�Fa�������M�K���U֜-��o3q��t���;��7��~tp��S�����e�xE�ٵ��Eb�y���b|��
K.��cD)Ƈ��-?.h�ҟ2���m^Ԋ��-�5%�cb<ه,,���o��v������V�z�kd�Ac����ޚ�Gx�G�����#)ũ���,α��v|R�(;�pS?Oe+�68��&̩ȩ˳�VbnX�H�4]{+�bo�̆��f�Ȳ��Ϋ0����r9��ݝ,��PEGr�wԸ.z=e�Y�C�+�}�P���O0�%�5�0|�(yT�Tx�gV�?��Ӊ���L����P)�T1V�'.`���z��3be��.��w��ʤ����]L��K�H��4ą�#�T��ۀZ��D��J�^���:�|����S�Y�_�{+`P���bLY����zѡ�{z�D�F�]g�0vF����f�`u���T^�˚9��+���Ǩ^�Vf�
�)dH��Lz��H��ةΡ���A��Kt6v�q�.W������n�`���B'5��Z&D%����*���&Ya��Ӱ�6�!�Nt{��޹׶�O"C�� ���
��.���眉�C�c�Wk��@��0xsT<�>J��#��u0z���Z�	�y���g�ڞ��|��]������}�J6��1o�̮�o�\���q!��]����"Ƚ��dO�,`e�6�i���/­so��2	�$<>\\��^���ۄ�a��5����'R�n��)�"�P���w�бˉ�DvЍ`�%/C�|�Pv,`�i#����$�̝3��R>��.i{����==;[g��ٯ�5lWG$��O���,^n�f
݈��tŇ�Q��e�T�<�]6k�mپZ�d�Ƃ]�5����y��� ]��$����d��ˑ��_-v��f�zgm�������o^9�ܘ�N���1�	���$9%�i�ۋ�>n����,l�5C1��A̐�]c VH5����ü�Al��N��Tqܡ��ȓ�5}�⎱)9ݧy{��v�:<d�E��E�9
p���M���%3�(ID5��6����fx��L�X���	�H�0q"
�'h+�}`+�}�|�[T�9}�{\ߢ���z�Er=K��A�Iwh��q��ŏ�fқ����T�� �rt���X��^D~�t�n�5:�GLf��"��mX���#��%�W���H�� o�v/��x>LoC�{��b`i5�s�<w�h����4�tݘ_	����Zv� �����d tL�<��sWs�3x�����5�ɱT ���ڙ�-X7zH��՚�z����d��È"*�ך�bL,�F��H�����f*�eCXX+<c�#@�Ox��aà� '��x�5�$����o ���z�ݣ����"�,�Z �A��Dd�,^����~ݹ��t���+@+�K{j�0��:�֩z�>�ӻZ�� �F|�/']�B�N��s~n��A:H���^o�������Y��{�$����,P	ܞ�ݸl��auG.)��YL�,q�f��z"XG��4SJm���.[i��l}��sk�K�2��JT2������ pm+�q������Չۋj�D8������g�:G{�` �)`͖��qr��Z˂$���J~� c�-y_� F��&���~L_٨)%�>W�lB�M���^����L�rt�"P�5[�	q�w$�)ь��6}䊇��5�����0(a(Wz�s0��K�?��$��qT]�-V�G9���J4�E�/�UD�u[���F�y�����D���������?� 9?���]���>o[���Ep�ax�1g�#I��4�d�5,Ks����4���Iv��h�Ɩ�nS�u�B��$װ<�f�j϶�������@��^���f#���=�%�_�As.2����v]G ����+�	;g{��Xy-�0Q��o��d,�4������eo�%��U�cx͕���{|f��\:a6�wp�����PP�ųW,���gu�>ك�!��0���a���h(��i��!-L<�c
4��33��K|�W���ˁ<��L���$���r��+�!���Sg��;չ+Z���n�owlӏV��t!5�T�pƯ_���go����3�};��1��3|��<"��#�}u�lT5�R���K��1�;H�u�/��k�v��R+�e�#ܨ��W%+��@��=��G`*;����Ȭݤ0�w�����kI۳��]{5?d�q�_;�}�Hܪ߿����/X>��|��CN�f��:�����,�����c��wXrzW�9Y�(��첖���(��Y�_�y-�'\�nS>aP�^rU���� ��R̃Ev���	�&ǣhtbM
R��V-��L�t�ǉ����1���u7v#� ��Y�:I/��g�d1�'��`�ى�3�G6z�R_Z��^�G���]m0�kKU�t�u�/ʉ
w��t��&63ۉ"'��S�����-��\���,͇]2*O=�;?��be��E&܌b,V.���=�eQJX�	5�f�!M�4$�N���kH\�jg)uF�m1O)��'���
����iRE��N���"����\,D�G�Zf�}�#���x��HH*��9v�L���LSmp��,��뭡�X��C���e���V��	������J��ԋ�ێb�`�#V1�'N�ɔΉ�{OP7�&�NAt�'o&���h����C�}ĪI!w/wcv�,�X*5�Y�\�l��d�L!͕����mJo."���f��臘:+����\�{�Œ@iJ�	�\���_ɚ���s#S����j�e��b޳BpĢ�,Aă�ݿ�)I����9�Fd�K金-<����C�hw��R�
m��s:�f�L� ǿ=\
��o裀���E��@u������{�����8�K�
���m%�����r��e,#b�w�v�z�e^��I��l��L�:�"�ab'�q��C�Ρ�z6���N�@:�L��z-)iM�8
Q�Ў�jbr���nA�b:����C���G(����+t Td6l��+I�G���G9�^;PU<u�*"����q��[���d�(�18#V%+�O�"���d��.��;`��f��L˒
���ć���'Tɶ��XL�{60�ُVU��?V���*�è�TCFAqx3���� d�B�.Z�����'Z�W /g�k�B|W{���50�)�GΘ$�F�B��n�#�U�Q ���ς��./�u���G��,|Gŭr�})"@���FSd���?��~J�d8�W�����(�ǥ=uW��Mռ�I2 l3Q�M����[}s�E�����뻂A��H �%��2K�ˤ���`���Fqd5�l����]XD��V+v��+ ��������Ց�A��:�Oܷ�n�t���#�q[{��nِG�'T�����PZ,��:�[��Pͺ:��׼C�e�t�7fvI�\���a4+["�(�C����\Z�����<=d��d��Ay^]L	�3,�ۨ�|�3���=�(�B20��s�N���Q4"�4
���%yu�c��ov�s��Q>�#�^GKY�]����Kٌ�<P�蛽gm)2�8�o����Q.��|l����;��ԉ�y��F�M:oGh�����!���}�O]}�R�{���JM��s�a�_=�CCQ�z_s����|{��qNf����ͺjL� �y���;�J�����Y�$�����rw?2� f����?�7P6?S�	���擣��TA����z�ĠP���	:�1ՠ�6E�b� $�br�I��w���l����
�L�����X�)(.d��;ǧ��%R�GxBO�H�t�H�W/�L�:�0l+�;�F���"C���&�EVz)xc�d�œ;�PTR���w��Ї��=Fwa�RX��P���U�~7����z%:"5�kU^r�\����<,$���i�#Ɇ>��>��7����~<�(�7�#�%�Ir\��Ĵ>�%IW�Dl�Z�SuQ5V����o =��҄��gES�Ś{���6َV�}��e�H��g7;Jʒ"tۜ�@���1� !��hV2����F.�,����a��Y�Q�Sm�WB���4(�v��ء���5e:Q���k3g�H�\"!(Ei�3 �38���:�{}���-Lz�GFJ�%M0y�Z��B�qH',Ϻ�����	��K3�o.�ɮu+��D�3��)���sR	���_z*eEm���=D<�Zxgtn�X2愊S���[���`���ŭ��_,��*^�~<a�kJd��;d^k��Ŝ��Hh�=��٫
�J��w�+)��6���TX ��{BK�DH<FFXJIkxjF ��.V�X��N�Z��x�to��_((�737�*�		q�����dm0�S�	��
��2�M��s.�,,���:�|����F�D������m��E"Q�c����� i=i����:��_|{3Ǎ�{�3k��F�e��)�?���@�c`�t��߫M���|q6E�g�xY8�����.Ų����{��zϯ��=+�$�X��c�<��v�>�77&:ja�'�7K��������������	���)��������00��U/����S�Ǭ���?\��=�d�iphKF�\���	��h��:�{�F��b�$!u|W�e�+Jz�����N|��=�2�]�̦{S�z{
�\�!��]�	Ϙ���A��H��:o�|��lk�'��Ԋ�[g�(b+�n���`�}f�巈����$8����+m�S\�!a��r�p�#�&}��������1E�=J��`�/K�ml_�6��0v�������/��#���D��{�u�hj�SU<�L��!�Z�*�>�U��X�7TW�p������]}�QN�&�Sf"�2�t�gC�,ڻ��,�,*]̦���+�[��YW�՘✑i&k�xn����*�7Nk[��B�!
Uy��5�i�vh����)A2�!�R�Ng+�Z��Z��^gw"�"p�	���7�hl��㡻أ ��&��(>�59<��	��uc�Ek�5����_�ۼ��E��9����?%��A��ֆ�1�Iī
��|-�7��$��a���1�Y�:�D�h����.�����>w��H:L���{["#��d1
�Y,{�=C9���'		�L
� ��V�
����ͣeI��PP˯1Q2;�vB�Q��{�t	�2���E>b���Y�L���X7�ȡ�'�.������*B��������P6|��t�'��}���-Ȋ�5�v�l��U���^V��1�w�c�4�L�W��kl�6v��[��G]?8��5D���*k���G�����"��[�/��̟ށ�'ّ'=DV���o������#�L�s#{�#���{�j��ɭ^�p��m��Ѷ�OR�c+l�K]��o�g����Bu��8 }o�7
>�>�6W6��W��?��.�����D�m�������=�Q�@E'�(|'/	���-^}L�}��u{V���r���au�����C-�|D�-}6-����2��y*6;'z�^�����<�)o��)X��2&^��`'�a��tˍf�s��b���!3e1O��-�(R����&M^�wR
1�����"�L �f�:�z+9|S�-DZt���E���<�g�/��ܸW����Y�����ϧ����~��qX����:���ioR�3�j�����R�0d&fAW0����LQ��~p�����*>ȫP��3+��	Rg��z�886����z}(7�eg녅�u�
��p�okkG5y#�c�\]����g��y5])���Xi�_�Y��s��~C�K�-�ֱ��j禘�ȱ�	�gy��~�-|����$߉b��B����]�/B�rQ��+q��B��(y;w�1��ՁX�89H+�6���1cì܌粆"`��?���h�k9�"�"���Ic�0����S�iu~ɬ���0u z�L�~X1ŝ�*�����{�:�3���'�%��ۆȽw�>�/�����fA;qFx|ð�*����'�F���A����:3OH��!��x���/��C��PI+��GT�f�u��5+K��Ih!&6���X�)�/k�u�'V�@  g�X.&�o�aFG��ϸp�@�^��n:@S��p}�����VtV3)���� `����n�1����-
�m,WQM�w���m��k���`~�h薚�ro�|������a;$��ۑB:��;��@`�#j�;'��y��g4������,ē����4볚�u�A6����D-#�K�⒔}qhyցB=Yc�"Tϕ=
��Wd#��B��bz)�=d��8
�S�r�l� -��2�v��q�)Nv#�^'<�/���s3u^��Q��O6�Tym�l�����k`oV��sHgdG;̭�c��o��Y��N�����ct�5�|sp�)��#�E1�i�%v�rݵ>
&~�.���E/�Fu��-�t�+LMۭV	 �}�W�2ß.u8��ۄ��^�΄���xn�M�wjNA�8B��z�x��|���~�/�T��LkFc+�q���l�:=[���[���.ztG�#���a���c��:z�8:}o�i�F��@������L)")|Ǆƪi���ڥ+ɼ��T�k�ۯ  ބ�>��n�U.2�%GD%&�����H<�-�LF�Q���￠D�z8�A1��x���z�zA)�x&IVt���k��WX~;Z�%��x��R:Q	�`w3mmOd�8��c'�O�XFr*%�f�w�n�8�̀��5�>I��$�$t���R�b"�e�OҾ�5�Ax�w���H��`�]A�N~"}�M��ϼ�ۇE�F��]�ҙ��_��sg�;.a�S��;�X�"�h������"+�Ȃ�cs�/����&�d�P���a7���l\�	�m`��ݧO�};�h5�}Q�pF�����f����,&OɀjD�ј��\����+�y�2)o	P�}�^a����-�UBa�a~��Z&��=?�"��!p���?^��5ΪJ ?6h~���s�Q��k�>*�\k�y�n^�q *����'�rr������������q��BR���n�,�(�m<��a�Y�_�����;~T}jEg��	��V1�*B��x��[���x���fUT������a���������!���J/�x� \Ӳ�a6yU?P���،(�}�����[�t�I�Yh��DV3�l���{+=����q�&y�B��s��v6ϫg��l�� ��-7�Z$�����"s���/T����6��D 
�:�A��3�x�A'�hY��s����5��CC!о�12tX�VVnV�%{P���^��hS�q��Yl�w0_o%}���V�&��	�h���*yߋV��ȔF�"O������[��`��ܤ��w��-E����b�Ǣ�)�ݢ�e��Z��h��A%�Ҭ�̇:O=�ю�Gu�����{A�Ǘ��\�E�|�Pr���+�
�CZrd�"ː��J���W�~��;j�y�2x�с�U��Iu�����K��66���'���
��N�v�f�c�3��ֆC�:n7��E�]7��I��6,��eq�y�"兦��`lKTH_��{H���������r��>��Gg�A����Zt�ߩ�@�b���w�q���Ek��ʥ42#�����
�T��7;;��+/.�*uJǻ?��f��Y���e���HκA��1�����w�^�G4a����R�M*���(�f|����`э��{:Nʁ��;�c�<�^�GIZ�F����X��H�/n�
�����gj΄�1�Uϖ*M%ӝ���!�pu��^H� ����<�^u��pc�(�?�X�x�p<�;�J*{B�&�C?����7��j&I��I�o�}L!�	�w5.� �TJ,�E�H�F�2�"�,���������ݩ}��E`f ��e�?9�S'�4tF�E�u+yx�)ge����MuJ5V{��U�z���
�����9����h�����S��l[�KLK�2c���v�_�D�WK�X�
z�I�l�?2w�,bP1��ݨ�Ӡxg�XV��O`nᶌ�|�g� �s18I�_�Hr�q+��H�z��!��`��$�j��+"����q���s�p��(�7�@[�/�m���P\L㖎��s����%%-�m�)O�'��>���=�\��B�8�#��PI�����x��}1;B�y��+6x�m��:��W7��7�⼫����,۳vz%�����ͮy�H8�F�~ɭ�(QZ仃�bl��6s�pvL�pc�4vHE�֜c�O��uM���!�[� � e����օ�ntC|�Wя�)i��P��ZrD�=��� ��%�Sl
ó� ��+��� �F�!ռ�ehO�buI��@��0a�.$p@y@J/����"M�N�V-�]'w��ꂁ����c���@Q��h�l
�2��Si���2�A��M8��A������E��{�87U�R�o!h!@�b���X�4����K:K]\'sa��!z~��D/�rVZ�r���*��7y�-5E-�j�)I��ׅ[�]��a�C����6o"�ޣ�T̞��!��ؕ]C,��NԻ�_%�o\X��\�/�L��3.`��+1��RY�q
d�Q���A�d���L[��3��}��G%�aT�&.�A-Q�j��1$"!���I�C�0V>��F�/�}V�~6��d��'���#5�yȺ4�E$q��K�H
 �q�2̔�s��u����Z�a�!�j_���kE!� ���t�|�S��:��8������X�����xVGK���9#�~`N/���d8��"�P���~;����)rUqo�X�4#�Ss.9e6Gv��	�!т��ȏ����%zD~���5�ʒ���@���ee��ɟ��T˒�P<q����%;���7Dɩ��+O���ر��D�v�QO�z��^�V����=1d9ŅǺ�/A})��G�
3W�Rk��T����.A�y�lg�"C	�|g�Q0c�~H�:�a�\R��!����K��\�A�WDS��is���fƢ�=�MbߙTQt ��w�������bEv]���%|'~��bh1K�""7i�s�����>��C��@}Y����86��a����"đ�V��\��툆��2�-�+8����7��.H�!��.	Z�N�+��3Y�K:AE�:�k)4��2��hN��YP��͠O���Bz� -3�4����aE+"�(�d���b��lќܤ���JK�ڦk�
d���®�i��`��#� ������w���`y1���(�~垹���%����0����[��������s6�&��	�,�uh]��$���kb]y�ٌc�3��״�J�w���V��*�h�x�Z BUR�u]��wH���p�_�`��,gh�䶛�M�l�^�qC�X�`X)�?��I:��C�*��)fww���a>���lD:��fov`Zo���79�Xߌ�/�7�����\��~�����K;����(b dy�x��@�7ռ���Y�YV���X�)��/���� 24hn%�h¾��� J�J�4��P���K.*��!��� ��M'쎟�)�iѾSa��N����V:&�~_�F���,�96Ν۱�KD�䋣�Gƾڎ��F���aWZz ?ٹ ��W�Ps�j��Z��$(�H߼Qx�=-x����iܒp�����l�q�(T��K�ۋ�o�T�G���r������S�,��|D��Ak��ۮ���1	'��Ypǈ�Sɜ�o��� ��OF�W�u]�LV>Y�������9��	K�8�;a��ǝvro��v�->�	G�D�T�vl9��=�1�
X�c;Y[���	kK�S3�Yw��xi�����R�0��*�jQ���������u�G܀��I_�����hʐ�O���+��?� �[+!���� �6[� S�I��F$�"xA�H��m�Ϸ5ii���Dm9/��Z_v��#����`=R꜑yxVS }͏ M3P8K�:r%Av'��
��+�U1U�؉��sQ\��=�H�B�� �ۃ���g�_��on6sX�_�C�μ@�S&u��*�p�0��j�Q�t��i�+��+U;��S��c�Y刎����w�;����]k��kąUe��HlJ�)�B3]	���{�f����N�20���1�F<եo��F$�fc�V�K�!M Ht���&p\? P"M�Bv4�[����w䆏���l��B4}!n��X�a�y�ھ�,A�^�6:��4ým(6ԊG���<�z����j�Ģe�Ԕ�*R�� .�����r����+  ��[ ��eź)���	�/]Á�'��#D��a�&i��?a҄`%�p
@���_����G�<
�U���-F]e�#z�$���T\8��xi�4A���m�U�{�s,k���]�է-��YQ�E����F˳VG���R���Bpl,���L��aV��'�=�>#"C7��5�I���G a���z�#���Y�9�xD����پ��k�js\��xC}ڈ���P�J|�TT�,D�f��;f?�� ��Nky� ����=����՝���������?�g�K�,}R��9[MA��
3T׼������'~�Yֈ�]1zר$�T�i��gEV�N�fp)Ka�6�~�?TR��XR˃�Nm��kc�)�r.&6&�^�+�撳�����w@S�ٌBX�E�qb5�(�s(��B�M��J Q!V?QݍNP$��N�^=�)�ɖ��L���h��j�P�J���F�T���a�?A&���Qo�()J�iz����	�`���=fS~�� ��9�g�nv����'ή<�Â�gs��ˉ0����M1B��~8�=]Z�8��[��x��SXN�M���0��U� �r� jN� {8����|=�*-���sY�R �(8��&������	%:�r�����h�\���1�D����j����/H�Q�3��'�w�ڱ�R����θ`v�?���E\D>h3
��9�h��Zf#TѴ�R{�ojpչ�q�	J�>�iZ�tk�W�O}��j�ai$�x��Uyt��D��p�j;峹Z·���y���%2����6�?գ(k�>'�[�;���#_�-	x���GJ��@J�����\��0��>�ة�m��۲u�q-�S�#��r����wB�uI(b�6�A���c2��ލ��T�pB��z�e��`j@8~nvL�/g�K�e�T�$�u�i�NRb�`�?���f�A�*|r�y}�X2��4%�{8>�Zk�ߑ��z�D����#�=9%�38�<Q���)r�	���/�Z����PL�_��n�+J����E4�=b�)�k�2�tk�V���`F�ݖ�k=n6��@�1��4m)OZrN*��m�%�GQ���3�YAK"y�M��";^��p�^S;��K]<�,+P�2%Qmw%�ù���]�����������0vv�.��9C��eR���Ɛ%x������g;�z�l�mj��'S��އ6C����s!��b�u�eYu�AF �4d�F�;|~��B��9C?&���!e�{�J�sZ�V1��w��+k�T
��>.ԣ�H���~��G_ž�>{Pl�7(W#"���M@0�Ge�5���Lt[���\��Jӝm*�H���HS�w\�i\-M���z�d�G�[��+�KrT�(K��a�P9߷�+�T;�b[�V��|�=��&m��>&�x��5��/"����k���ǫo�����8[)�|�_�d0���8��^�e�A읞�!H��ewJ�H�u|l��=�+�~�2�/�r\�i6o���2NAtz�L�������tq@�,�7Gܮ��D֍� �(����X$ X>V�k�l����u^�ϕ�/�\%�E״�֐iݴ*2£z�YU ��\���R��CW��"��ĝ������x֤��2S�.S�Q�q��M-�Q.ٗd ������--{Kq o �<Fq��qG�k^���z��uj�x�[�]"���gʾ�|ѐy2���m�ʏ;��EF�[���yPI�P�ZG@�I�J��x��-�j�f�.i����
>Cf2��E�}R���c`x.XF\��Z�f Fp�J�<sZ�B7���}�R�A�آ�B�ɾ�g��d�u�ѓ�u�g�!�Z� �(���q9'օ��#���b:��Z92Y
�(po�5��@�W��}�iG�KR_�[�A%���x�C���,7�0�K�L5tZy_97�穇{l&Ņ:$�I��~
�	Kp�c�滐��oJ��q��c��e���q-��[f��J�����}Ɋ�,)�l�.w��F�:�0	�z�����c�_�u��G����%&��||�P4-V��=֙�z��y&j���փ��@��j���z���k(���r���	F��tϑ�Z#
�)
Eli8����j�l��`���vs��,��_e��+B�����J�����!Y�gdW�͖����<m��H�j�>Z�5M2-w�kq% T�R�[�G�֢����%z�v��I�kp���sgl�d�4}���.�)��)Ć�`�`jy���@�y��t��1"'!TmL	��b�����)�l���g��s���g���8��`>�~<�!k3��<�rV��ל��4�{�2cV������u^E"����U�t�����)X��{��E���m� ���8-a�:�{{���SS�@��%��r'Qar>���c@-޲�09F��x$WF�r?����@H]S�B�l*��wy~�	<�F��Ӯ�҃33�#}1�
���G�S���b�4�ŏ�蒽G��,w%o�.Z��FF���9/5o�#y�ø��'AE|	�F�Y�'luK�EQj�&9F ���s���ZF�nwb��~�Z�ͨ`vἵ�Դ�.-��C(��V�Z�"<��Y���,���yƈ���tQY���i�1@��߁	���a(�#U�@c�⨡�X(��;(���S�~��?�W�+
.���w.}q΄���bё*Q"#4����x,&��|*, �`+�2al��;*!�I{������Ж�a�u�:�SU��ï�1#nw3�{��2�17y_����r�P#4/��o�� -$�Z�;s	�4Mߕ�q@�<�!�mF�LY9�ʺF�,�f˻�w��na���*�˂{ � ��I0����3R�U�eY��YB�{�v�E���F�0D8��"zm�=�@62t$�| �/j���,�� ���G�au~����w�'"v�>KfaZ،��IO����0Y�+�>6����2�ך����ZF�PYy{+ۂ@����k`ŭ�[�3mŦZ��m��,]�buN:���^�����`%w�S�hu��Tv�Y(je��m.�{�"��4��	�Y�1�ߦ�k���^��_>�,%
���:0'��X��@��@�5�+C냓��Hndk�� ��S��g��G�{w��9��h�IL��g&�0j1�9�gx,����$N�D��@��*��q� !����x@	X��+��z&�E�jMkSFy���&��*M榹VHu���},k�k⒥T\����B�D���-��7�=:%?P�X����Kk���	��O��U�K�ġ�A� ǟJ���:m����x����`�*���}O�0`�f��"��/$�A�Z��w-�F8���ц&��ԉʭh�=�"K42��'�q�|��g�D�8�]�y�\�\�{پ^�Մ�}�`Nt��߃�<���Ke�S!%�F�Ҋ]����nK�g"�d�����l~�ި�X1�}tw�����]�5x��k�
f7>�m�`����fL]S+aVnb�/(��?}*�Hȿo�e:Χ���=)]7���R�cr�&2=$�3p��v� ��ŧ��$���|ZD�Yewu�(�s{E:��<�!����Z+:�~F��8�a�8��Z$[�.˞Ǜ�����qe?�]Rk��Li%��H?QS�;�؀/D�����z�ұR����s�Ծ�z�YV�9~$3�sy[Z�\((��'�^�b���64�`��^j�@ۉ�}����4k?�KA�I�'�A���P���Pl����u�l�5f0�X	�����(�Xb��{4���=h!b��RXѸ:�?�B&�@w�Zrv:�"{��[�:^I[4~')m<0���/�k}n�J,��ŀI����l��ɸlHm{j�6g�4��g�;%Z3�C��n R��[0O���8huZ�ʷ��'D%���в`�5 ST�{m� ���)k&.Pt���]���GV8��^=��-�-O��_���.A���yD''�h�֊���3 5i>��l�w��fZ;�3�qt�G
����
�G+�!�
�'�R�; dX��p�x��[p�2y��^�S��E��Ϗ4�L���N�8�$�½x�D����nGY6�ړ�M��Y��Ȱ��`�皡@���T���5���${����D�~n���<�����׌u�%�3��SA'����Vc!���řrp���)��� ��*<�K�¢n�H�Q�[���3��Uv����7iQHMlJ:۴�Hu�e���KԼ'H/;��H�,WH5r���l0���y�6J�R�օ�]����kvYz����_ӷ�]UG(>����)�oV_;��Â��r�Ċ|�UQ)���y@hf�oʫ�D���Ϩ��ה�	waf.r$�M�
n,�`q�49S���I���4�ۣ��×�o	Q�L� j��7����k5���0XJ(W�:ޏ��!�H�><@T��C�׮��Xn�����r��OkhSز_�Aw�V�m�ə��a%b�T�o���"$�A��r�?��O�[���\'�QM��w|�F��W7��#A�m�0G�+���"ɜ�4	B_3�ܿ {%�y3�6�G*�p>�V�g:���V�&���T�\^`�,3���MX&:D#��rCV�[)P�ee��7�6Dޯ��-V�K�����_@,8O��ibF�Q�x�A/W-Κ��7h�qi�&���� ���i)�J�=mI;��cd?h-�-G.���fO#ȓ$�6\�j�����NE�e	�:t��1ڥ;�N��0��f~
D�^��Bk���*+�<�9��&N��Pqurl�cD�T�7�[�+�m?����ѫV�����<R�u�L`���W�u��F	���WI(�C�3��������Ӡ�i<o�D���I�F�W^> �gņ���PD�A[�6�5Җ-��۫��}�.0 GZn�*�3Vu�RM��/m����@A[65�����D���mt��[�����H?���F�9���!"yp�c	�0a4�U�G��k�s;y{g$��Z��O�����z2%�������7e��� f7˅��.CI�/٬%��2��x:Mo����N������I�]�`�X�vF/���+~�S�mDܝ��m8�*f��2�0��gK�_���#BW���&S�<�^�ȝ_{�~�ĜR�x-����1r���C3��M�����RG���Ǯ 5E�q�KO{��u������Sv�a�� ��V�s�*J07D�e��qV�N��$�ks4+y���į)�2�#�n5�ʼcv'G�<�͍v#��~���9c��M�.�;ٱM���I�|��4�|qӿ�o�,�J�OeQ(�ȉZQNA;�9���h�H�Q��D�D�0�?a�yS�s��Z��Z������[�<��|��@�=�=@H���?�$� ���a�_�Ei���3��w>VU<������~�\��i;�{X�WZNR��IA@1`�=Nɴ��O��Ӿ�,t���*�nr�b����:�y���y���\��M+�i��Z/����x�֡Hi�4������-[I�\�$QS{�B�W���Y����)�q�)F����C�����	yƛ��4� �&=%��i�(E��_�)�LN���L���"{J	G5h���~��P����Q��VT�S�����ڨv�׭�y�/�J-��R]P�����7��T6`�ۥ�^����3Ά·��~��"J���T?��$�g�t��D������*��4���P�Kփx@�,W�/�$Xy�r+����Ɋڡ/��PWf��pj���Ab�`�l�롮N�a�B���SrƤ)P��y���l�E`]��-�V���w�[���[~$�����ūn`|Ѷ+7O�"�V�V�4��s1�� �jṍ�l�l�|�Y���F���ko�G�l�G&56����y���#b��F�/�}�Ϊ��b�Q�yHI#�׋3�ҩ���*ވC3$�3����͊����&,B$�:�a]�ʵ��F/�B�B��˵�t��偁��+�,�&�/ ;��<��4Z�!	�$Ϡa�E^��sL�\�WI��S5��&h��NYl=Ƿ� ����������z���o`�N��*�y*;/�BH<|m��z���C
���c��<�8�s$&s�A2��>��_��.����ܾߜHi4��f�Ba��	�E­����$LW�њ��í������z���e��
2�o��YXpLH�)+K���,�@��
���U�ܽXc��饋O�LTx�&WW��&�0<8ݠ��'�Q���#�#�7�����:���)�����Ϸ��s���$U�])^�]�<$��m��E�U)����H�(��"$��{2���-�e6�h&uVG�q�6�@�U��~��4eV� �:D�P��r��0ѡUSNâ>���H	�I#�}.98�軻�t
��ՆJ��ӥw^�Ӛ���}��/(E�7�#��o6��d'�&�Z����GJ��/2���Hpr�Ǥ&��U�mg�B1h7;(w�m��`��q�Ux%"n�u��������b0�h/*c��>.�\0H"���R�,�\����}�ZH�So�&$q��m���N�*���\!�L�g��S�R]��yT�^���N.�O�S�i>|�w��Pѱ3� 29�]�e_����Վ	���ak��el�=�x��*/N˯Mv�;2I��G��M���o���n�'?��fB)�ؗk��;���g���a�7 ������AB���XԦw�Ę�����qleJ�ۦA��>.��:��%╦��l��ʎ5YxWֶ��@M*��G�Mh���b��IX�p}�ʗ���˚�,���h�	�.�"��ф�OK�O�W����.N�3a��+-��HJ��'��n4����B�����E�Ȋ���� ��	�j:ō7���(��Z�{�R�}{�DΔ{Ҷ��K��+�4r]��+~�����O���u�2��{��#&Dt�5rg��x�� JPJ������&�0���!����~M������~�z���%ƽ>�Aj�����NkAŹ���"Ώ���I�z3�1��0���f����G�Hx�%�Ow�"-3�����T��m1�#{%;����izW�0}�&�w��g�,�;��>5+�/Y+���IvH��ly#(7h2gIA�X6z~P���qx���&@�/�//�fn`l���T����S}C���k��E��ȒY�_��w���L�]�U[O1}��J�� b�Kˢ�"�6�s��C2����^�e���,�\���~�߳MӵG��0dC;o��`34�?�a�y>,�2ޥ�>V=֒5�ۗg��\�A��4��Ρ���.��\�	x�n[}p�G��L�,Qc'���Yj��Q���AL ��5��;Q��ɑݛ�ή����RR�<-r�<%��������_���LRכL`��?�1p�����KG2�Q�ɍ~�H�Č�$�	�#���mc�`�¤�����UЀ���{u(���=8k,"�qi��.K
t�7�ʁ��P���j��ad��	΍KTD�E���B#dEo*��TUuY��@RmFtɭ�^�K�Т7���FXL�O��|ذ���`�]-$h��d��93���QY��I>��u\��Iht�=��(�ҽ~rM%ϳ��e�F��A�d���PP����8gx��JH9�1�x�� �ׯu�Cʖ���Lb1�K�uZ@m4�.*6�@��"xW�nV�Y��D��Ք���Y)fb4�4���;s��O�D{b<ӈˤLH2'�+�KH���m���.�Z�j�����di?��P�����q�k�W$�����k.{p�g<�����͑X�p���t|��'83�wNǶ[]/#��+���ޣ�r�;�W��v��q��<��ɩH��+Gm��/�$.��q��K��+!���Y��o�3-��\�P�g�?S���go0������u�<��&\p��'2���Ҝ����_$�
|���4)�Z�2՝/Pd�l�'��Y�ȅ3aa�6��|x���\S�O�T ���M�]k@\.�<�5_�Ai`�`�w�:ǧa
���ǈ3aݏ�n���o� ��bE����{���#>��tZ�s�W_��:������K+�j��X���8k���As���P� �D̾"-��k 4��T�F����f�&6d�Kz�rt/���\�>�v��^O�s��7;y�u授��#�#T�u �=
�8���h���ᦾ�� ����I|]�d��,�D�ՠ��*���q�k��Տ�%�����{���a�'}a�^&=ѯ���柳�$�B-�B�~�kW� )�P�L"���0��r��&5-Ӌ1��'��v��<G���;�c&A]�������]ew$��IϮ����2���憜����n���ͳ3ɦ�Y��?!\1�R1�1��}CZ���$�L��}�p ����۾�{0���=�[W���Bd[|�a�]�|�q�� ���+�OPD����/c���Ҹ��o�����/�]vQ�]��*2`���:�
{=��kT��ۊ��VH����o<�/N��x@������������@BHC ��������L8Z��X��sQ�3�3|�{�I�����ސh���Rj���#�?/=���KѦ�|��a��I�r�hݺ���WuRb�y&Q1�\ D믃 jʴ.�6�#�b�� �xLI���~t�hW��)����3>�m%=S�5�@�	����bp �����lwb\���G�B�	�i'�� �=>"a��!Fpsk�:��]�A�+�3-&:'�,���#�
�`ě6Nt"2��jZ��KƳ+�r�E���Ran>� U���q���#�1)�8���ϕ�<pn�����V�3�W�d�`J*�^�-*�	8�Y'f���D��&����n��ͬa�Y(SI��+T�7��i�XPJe�[�J�/�LO�r3�q@j�Y
��ӚQY�H3��%��n{ޢو/���4l��bu�yˏ$�'�+�#��dգy�U�K�21_��j���/a0�X}��|�� w&cu�W	ż�e������we���(#���){%�=�G�ܽH�'��EƇ\P��ʱ|%��(^���������Ryd���N�V�x��$oɿ�F�/i�{�@�KA�9?����W���d�Η�~a�c��
'�WF����E��	Q�o��S����pE|�jYA�-�Ex��k=���n $��'���w+J���_T�-��=u�.�b����;ƛ4p���U]FؤDO��iuQ?Ud^�%�Xs=���Vч}�s�3El�����0s�UV�ì8�W��n	>�P���J��㏤�c�$�[;�S��
uP,ԅ�'Pl�dMJl!`���gC��+����Wq�L�E|w�iy��ӁW_�CqXX������YJ@��RN淅���ݘ�[����؝��xez�����K�lia�҈�*�v��Mt�A6��]�.�W~Y(w�ׁ��>�[�
���Q�*� ��V���h��	��f�N�Dw��<N�׃��r��Zd^X��^�v�̀����G�7�z�AZN�b[����?�
��A��Z�D�X��䟎���=��B��;��	ul��<�h��o�i&{Wj����ow��M�匐�w�e]}�|WiT�����ڪ�l[��I���Q[�Ʉ�
y7�Β4���Z�R},��I�	�����~���	�݈\��">��ɽ�9�Ҙ�E��HkW�B`=��T�`�،�%�3#O��"1�2#����K��� H�'SR�W8����y�A����Gp��? �A*�-&�Ȯ"0���h���N�m �����!��`�YYi��Ȉ�b�u'� �� !X���!�iArR����8����Tt������`�R�F�h-z`D�4��T�GO���z�b^�2���~���=���kh�`�@&�Af��"&*�ׁ�DZ�V&��g�P�Ƌr"���x~�;�8�����,�
��<%M�]w+׷��m/]�r��u��������҅��Y������un-�S�"eF埃�t.C[�?W��ҺBeF`��h��q�Ɏ����6f��)��pܠ੔�e5�þzG]	S%�N!�
��r�cCP���?�u
I�(�$��Ja3g�F�r�������Y�R��N*q4�j���Q���e8)h��J5,ŝ yY5k~�r��d��'�Hm��.�/�;��Zg2�5n+4M���1b�P�����"�Й�^�	��p�<�����o׊=����ۻӔ����Rⷥ�a�1��	�M�\̲�qoH��� c�w���q������� �Ua��wۮA	��ݵ�~�]b�n���:ƅ�db��cJ�+�L�M�:� �����j��H�!�g�f�t���z�e��j�
9��(سיo-4��k�]�wj>�Za'��$��K������摧��2�u�2�����Nu'暚̚����2z�Q�fQr6-���g�%���A��3Ym���&��=����7��G�B�V��",lIp���O�H�}��0g��|�'u�L���$�:�ܪ�].��R-&��'�:���,A�2�|z�"�?ϣ4R����zt�b���ն�"%��/<HKO�ɖ,eKwCJ�K�+�C��QG����,�r��0')��"ǿ:�]NGv�T������3�K܀���->U�h�?5xvwp-�^G���H��������7�=��鷳*Á��J��w��`��F=Hw�!�� ܺ��r�d0���d�bS,ͨ+�& Q�]*�e,��?�2��>�l��V���,=��:6������ϣ=�h&w�#�L��J��r-ӥ�3O������W��=�.�\'��X��sf��G��5��Tx8� ã��Y�n~3D���M��n/˂3� u)��eT4�[�������1o6'Q;��"}}���ͤ���e��;K�L[E���D�><;2�v�{�A�]4ԏ�F�v��*�`���B(�:�5�����@?�Q�5�S�~����R��ϰ�C+��!C���'�{RDo�0���0�����qDJ�_�9+�C�1|�$r�$�����x�dhJq��/���Rm	G�S�7' ��6RM�F�Q�E^���G�tM9��DR�㢽,-1)�{qXw�r���A�^9GM�lpdٵ�ڷp �^�}���;���"� �$X�z� �+;�c�����6b�k��4&D$��
�����������F�5�ڗ׆gFx�"ݗ�Zr����)�X%�>�I�'�X%˂��z'E�$Ѥ����� �HUE���F�A���0��I"��%�����4!?�ke;C��g�[J~��	P�К��������P�5<=�W�y�dˮKc�E�,yFG1���LN�~1wYԸ^is��h#��4ҕ�I���G��D�ǐ����="�,1������	�ه��bN�4�!(�i;-�w���pJ�
�2�"�2�_I*H�l�h�iX�>�č&�������c(�]d�V�_�O]0�.�O�L�b��:_�\\��JSؔ�ƙ{'�!���%�;�L,�>�6��ZW͔.�j��1�-����P�2�Ņ���c�q�H�87I}��������[JK��D�Z�`h�~�>�=sI�o;iN�`6�=�l�_���d6�-"z�r�%.��&�Se�AT�u�h�(G!=K=)�9
�$�	w�xC曉/"���w�;���F9��/%��O��ޢ6�4��qmU)w�8��g�[��`����DQP��i�<1�s���S�
l�'����68�>\�k^�3Q-��$��_j�l�S~����bL�i�<��i� ���d�oDh6���������	����Z}A8per|�;��毶 �g��H�N>��Q욀����Lp�ċ�0c��q�Oc΋pZ�8��|��N��x�X+"}��/�7�yR��j.�r�g^Z�c���ê�3�З\�(in��_��Ԣ?+#�xu�4q{�d�G9m�)�58��[��&��F@9@�)�E�=����R�zq���x��WJ�m/`�W�5�c����xns#��j��6��"8���γm�=�I�b�~<��X����͕_�_�ָ<�(��qi��F^w�v�6�N��+d�����/a�Πklζ_�ءJvmB�K�!X�|r���7>D��"�}�%�b����gi���r�~@	�e���e�C�N�,��ʬsU[��9|^ᓽ�[P�n��]�tk�e��<TjG�܆���C6�kg�����u��WGV6W��/�jR��
"�����I5���O�G%|�ʬ>W��7.4��lR5ȼSc�78q�2[�;�<�����,�lj�b*���^wvІu��]�W�����<hɾ+8�u���;�!����11�#���r�+^�����T����"�`=]"o@�_z�;#�� ��-jF��[���^�G]�������:��>ӽ��@l���N��{���]�����mk���� > ���sG&2�w�Z2xiB6�<|����DrOn�l"��A"�Hy�5�+��ǔ"���-F
�����]$��a�D�^�rZ�1q� B����S�[�|u2�^���2�r���N����OL$F�K��\v"�k�r�+��tk����@ꝈO���G�����NӃ|�R]��k6�U��M�s�$�W�t2�=(����af�f��/H,�fB�[��0E,Vsދ�ڍ���K;K!ւ�j�R]jq?����w�zcw����E�G�TC������BF���E.3�,���|T+�K�<��#�y���������j�@�1�V������e�BJ0b����UI��@�E�����v�J��4��v��t
��,4LBd�q(.phV@k���������?�X�YKf	�H��55Bq�t�ih-~C4Ŝ����@7oP�Z����	y����w�6B���+	>8
X��N���	ln�)�N�Ŕ	��1��y���6Ȳ����/W�>��I�v�Y��Ҩ9yʄ�%�ss��	o�X��{ZlB9��![�Ј��͖�J��4�O��w�S�|6�k[�fE���r��R�	0�b��܊�� ����\�s� ��ץdW"��>�[#WyQ8�t�����r��\ �5�P�
�����DRw:����a�0>�ݔ�����}��@��bT/�
8���2��:���>[��;c�C{�N��P\�2�\_�^����f�J�Y�����g��UMj׆rꦁ�[Y��w������(ꑻ�	��k1��'�;���H�*K[�#ʻ5B���v���d(A�qc�MJK~�KBAUI��"�	&��a�K�PvK�r�.�,���<��:�C�g^&T��B5놚��Cڒ4�6��j4-wyX|�:�&+��~�6/LM�e�M���||V�#�(�T,013׃I1`�-`)�?"���[�$�ǉޝ��M뀎!ٱu{LGa�qs Q��C��nz�4'
�Ϥ#�D{�p�����k�����e�d�����-ͱ����{�h��5�c1r�(��-��$U�o��d���ڛؼ���I^��zMN �n�[ѼߥG�s{l8�2��<���O�D��#'�3M�1
*��+�P���^�I����>����p4r�ߧg�	��_�U��M�Wu��e�|����Z�w�[��C�>>m&���bI�(�ϰ�+��	�dXJ4��|wQ�R8�x=� J�0���/if������jX��tGʩ�[�N����n���S�q8�_6'�Ŕ_��~)75WC6�J���*�s��=�L�]ҧ?Z��=�ؐC�g��=Eê���	� ����i7W���M�]Z� �	Kh��ɭ�I�.Oyc�Μr�E���I$����U��6N7�v')�c���E�����$iՠ׆�˭H�l�_)�ݜt'n)~>���#d6N@"�^2�����.s��DAg?r��������LHJ�c`)ⶀ�@�-���y����ߩ��+�rZ�����α��)�aD�\l�%�*����:ڗ���Ċt��>�O�3�8h� =�����s��*x��خ�l~����z[�r��0e�����e�2�Jn"��lg�j�Rd��A���u-��@�Ek��Y��-�OH������!��Q�gZ�Bвi ��8���.@CǕDo�K�����MV�湝7_<�MxG�����{���!��G��1H�[B�W)6h�A�>@��fx'����0�N��I	�ɲP�D�뚼�jX^>�����iS7$;�q�����広d��L��Z��A>��4��ڳuqR����}C`s�u�����r�nK�a��Wͻ<���U�l<��LC.�2��*v�d�TM��� �tf�Q�pP�)�r��qr3ڄ�녅��PhP#Y�Wa����s��& ?�6%������>.���� �l�a�7�z&r9:��r՝~VP\
6�s���Uq��`�Y`�Y� ��lJ�j�D������=�/Y�Y�r�5�����?��]��zI�}���ZV�H�6�w�	�k��hgxF�Q�	5��5P΀�|�p@njg�h�����q����ӠJS�q�!<;�îz�c-��`�E����Ai�?^�|��ۢ�~��v.v�axDT�rxzj@H�N<�O�H�h����M[�y|g�u|��"���^�����^ ��cZ5�O��>y�V��>;�$b��~�����$�������7l�U�Y��F
pѵ�҈d[S鞈�I+�w��C:	�:J��~\�ڙ}���p�k����ÊҚavm��*�E�B�г�8��40�����)Pg�}�E;�sW�@c� ��v���~�yz\����_&f����v*�Q��j*0B���c+�)(���1�b��R�#$��������9������

z�J�w�	������)5�{�gC[�	Mm��'��c����V �=F&2cK��M#Wf�Y�� U/n3�fq�yk�}��2\k���\�E�v�b��Z�pY��������f&�D��Ƞ���Yr��w�G8M8@��A����f��)�8�u�s��_>�ܽ;�9���������.��.�� d9L0���i[	�(��!)�����V�l�-$ �
��I�\Y������X�zO�s�uD�p)�a��:����k��)�rs��9�sU]�a��@o�y��ۃ��|]2�GK|E��ĵ̂91b#�nN�#�-捥���>\�H� F���N8�*��&R�9��n�x����^_��U(6r�=_�8�N[�7�:���n��o3�,p�=��S�4�񬟈pc�����Zا��Z����|�g4ph}���h��[W��/��Գ�'y/
������ˤQ�e/ ��"�x)l�v�9��k�7�ϰD/��p;({Wh���)+���z��-���%��t�B���Y	%�}Y`�:���(�}�+Ҁ�g��ݔ��3�*���\�\��L[7G8�Mzݱ07T����8bQͣt����HC���=��-�@"';��2~���� ŒD�k�}���ճ���PռF��>|�G۟���P /��}CD��'�!O:���/	�����	ộy��#{ҶڃY��"z��1sþq�*��䌢�wXc�	�ppuI�<7+�[%�/Y_<Y�Zq��U�t/ UA�89��+^��*g�&O˚��_N1ʣĊ����T��&��߃��p2O6����1jh�?7k'�6�\�b7���@!�C�v����r����Y���s��X0o.�'�,F�+Y��%�A�f7f��KQ�NR�W��uxhbn�G 	EW��hh-9������̐@�����@F�6��y!�q��p3r@�M�7r���]�{�����v���q)�ei�z2����m��˺n�;`���4Pq�v��Ug�T�0�ɾ�Js�fgN���MN��H��w+#V +��ĕ��Q�[�ۖらw�CC!>c
O�eo6�㥽�lpö�@���W�څ&I�=<f2c��h��|�=]<��e���Cm��B����Z0��9��D���{gϊ�hp3H?�Ż�L,))/�~���藟��w���+�эlâbK�p���u��	F�sM�f��d �����_�.�WE�1�8�@�N��A���EnOX���p�tNmi#��B,���#�7M��h��fdx^�:���*�i�nm���	O`���v�b�$�����A�3z�ծ��?���H����4��ܫ�(Q��
���ԉ���fo�WXN�Uo��P��"��7:
	�V�Z�xrꒀQÉV��e2a��̋@���˫�šrud�M%�idX�;�N��pP�W�áY�?�o���g�5本��;u[A�V]׆��^�`����̫�{�o�Zb�f�ht���&}x�?m���!������v�K�e F�
\7��,vM�!83�Lg��(Y�G"��%��Q�M�JO�
��Q�S��sU<G[8��@R�+i��Y�8���}���ʁ7NFjT��C@ �{��?����z��<`�D,7�=���"�E\� �%`�:�N\�`���� ���
�tdN�à<��6;��|Ϛ�E�=w��P鏆eg1�]��')��#8&9I�)�{N��YcIn������O]d�L�<�z<|T����/~�'�0�[��
ie�]a ģd� x�Z���k�:Z��o�>zAE�;Zgd6�iMH�u��i뻫/i������댽X���= e����(Q��J*B[���	��ٕ��O�J����"�L�~ݕ�O�U�sL+R{�t��۩���B6���.�s͉{`|۩�Gk�d���?%��p���Dk�{rՓ�<��ɜ�y��ڟ�1>l�)��g�K�v��՟�s@��"L{�����&����ŏ�A���;�"�Xč�<|�4���H�ە�^�Vɪ���$��eE����	�(V�,���v�W���awQ�}7�ʳ��>(���X�Hr�hl��a:=RL��|��C���P7N�Σh��ӭ����yZi���w0��������Ƈ���n[b|Ą�?�񑨹��a�	�J��w�A������5���UP��a������,�w�ʼ�8������,ɐ9�b�?uGn�[�1�� (hT+�����0ju�xEh�av?�Q
������e�[A��T\�	�$�ϰ1���dSY���b9;����<D-r@�2��R�t�7�L�qG��#�BԣW�=
I�CDل�i�P��?��1 �D|��; 1���t��vY�V�-|b�<�[��f�"��5v�"b�ܺ):H�,����:�%��C;� m��́a�Y��F��^�]lsH7���#�����@�J<��LL���m��c"�̅������O�7�<�Z@�L@�sؘ�2�ـ�<�dN+ ���l`p�*u��+��(�"����\����/?/����F����Xi�M92;������̋�ڷ-�����D�Q�=�Ա�������Ä!���K���#��g�6�?��;����M�n^����v2����,�r����V{);�*M�DA߶�0n�Aq`ƒI�}}��< Ȉ���Ak���  hY��d����ˑ�C���W��[a�7�G`h���`�H�m�^��Z�:(cҮ�@�J%X-�CQ�f�����`C޽_��F�{l�}	+8D@��]>K�ޝ�p�o3��H�b�Hs�&v��1cf\W������[z0n�Ǎo��r�/��6^P��|����K����p�u����)��B4F�������~�n@ �	���;���O�>�=�&F���imۿ�����"
"�@t馠-��Ħ9�M��5�&S��~��m��y�[���y���z}���"8 ����A �Z;���2��}$q{`��e��Dm�Xs+�Q��1�!��ݵ�3��YN��yg�-�����n�a��`*��"R?O�#&%�&*{j r�@��2�Cvn�ܽ�(����MV�Y ����`�yK"V[J����1hD8���2���"8%�QzBCJVs�HO��I[�0��ҧ�]6_�P����P�Oͯ�o�m��~c{ǖLL.�NIM���X��ݎ�?��y]��?䐃KJ���sJ(Zd��w�g7���-��h��Q����ع%�tv��?��Փ�وTk���u
��'+o�1��o���y��9bI�k���̇���)�F�Oʕ�c�^T)��ɾ���6�^۔}�n�d����m�I�J�G'w9q�k�V��:^%�C�cbtz�!�iH���K23}mv���O���AUSA�f�^�/�	KR��W_>.޿���H������SQg�r�X�����#�A{,��3N�$�%f�EF��݊��+�~-rj���Td��I(��(���R���gv��;=�`�Q�P��\��0�9Hޜ������w�Fn9��羘	��I^؛c`��{�i�`_����}�5��U'�|tL���������{79�g�7�+�z�k�*�Zk~jʱ��@;�[��H����:'���f$I�c�v��X�4���J� 2U��i��
x`�2ר��t,gYj7Fy\Q�Q�q���[�K@]�G۰3�Z�´X$� �-z�T��`�0�Jڞv[^�pi~� ���M�y_}�_��go;R��i�G)� 9{�-0��xd�8�� ���X�0�����w�|f�/ک_���4��S����n�v���l��!��$�u2��58Y���B�N+f3����� 
�4�`�ʮLyd���atMc'�����[�+�}{�h�ȴ����L�ʭT����.c_x.A#�ianAo,���{pOdd)L$Z0��fי�)�OD�{�7�˾+q�N�l��F��7�:�ϖ�E�=˄K�n�!���8��֕���������i�36}�G�JN)���������F��WJ		�U^#o�b�%c�������|[O,+��T�H�ONq���\�����I�����L��^�Qg�1��׶��� ��(L��W�X��(P����%}p2�,_�ӜE�5��{��W��o"<��#�1�ܾW��e�F��@<�K��ezc4S�f�?���O�_5.9�e
���C�O�J��j�R�fp8��]����X}�t��@��4v���`%�X����|�G�Ø^kY3R06��ƨ���,L�8?T6�R	�)����P���N�)���T#!�i�M~hf�CՕ���Di9^�o.-Q�D�d�B�j�S\�0G������
f�$�3�&(���n�O��$�
x
@�33��_�H��5+:~�%^�A�sE�@��r��v}h�{^�@ojd=�\�+d�ΏA�j>E
a�>�G����ɿ��ߎ��j�&;<� ���C�K:I<M;sVh�;6u+�b��Oo���=����E����q�_���$Yǆ��53Wn��%m@�xپ"�j��H�Yi���Nb�����8�7�,\2��AJ�0W��lK$��j��w_2~���:W}/��ɱ��0�8_����$pI�?m�]�ͬ�ܺ_I/e�+��N�1;J�����Vَ�nt���~�����#pC}���B㑛�?H։�ʸ��M�+C6w�r��_�n扴��Y��~�8�V�-�2�^�X�4H�r/��z� M�[���փᱍ�U��ƃY�Y��0�����i�/ŭœ�Ēm69�(p�����~���������P���r�G��u{Q���VҦ�#���i�H^B�b��\���Y�@�I\I�&�O,r���v+o��،2�i��3����f�p��>�?��	O�:�$��^P�|������YLqp���a
�Ch7zMM1�h���[�f�)Ήs�)<7�H��	udJF@=���9�5�$졎|���N��h� S�K�z�p�Fyq�Ci���3��O��/G����$�j��Z��P4��KL ݼ���V���=6^2Dwֻ���a�`�ʓ�>������.r��΢|��z** �P���x���^#��Ϭ�v	m*�	��Г��KW����<C��]kƨ���|$;kF"	��Z�k���DlVb'���S�����<�!Ⱥ������𫲈7:���I��E��U7L=|��(�[�ɭ����^�2��W�9O!C�L���F�SY[�$|GL�5��N��G�n!a�M��'#nW�=Cv�#,l}'9sK�����y=�N��N��|s&��Xo���~��,FK��Ը�Y� ������޴.��%i�Yܬ���.��8��T��;Q��X���t`�:����M���o��ഡ}-����7��L��+�Q�vz��m	ߛ������EM?���+$K�[�I;�/�����/i4	)ހ$|�.��N��}�-6����q`��.�U��ޑ�� �� ��'�ԏa��;�����<� �d�GM	�I��eK�1����af�<9��ͫ{"ԫ�m�u�Sݷе�֯��dqc��W�~tΌ��2ZE��/���S�4D�?+���Bu�X�B7�6�.�z���'�Lp�4���y��OKj�_+�7�]�Fe�0��R�v�|�lA}Y��7��5��&��n��h����ѝJT+i�&j
�SV�#��ܺ�Km%P��9t��m������'����8�j$@��&��=�e$�ݗJƥ0��[��s�'P�(3��{LE Cq���$ή\[JկS��磔;q�$�F��|�H ͨ����'�V����~���z�G/)"?��6h	��8�z~J^�g��:خg.��?*�йTU�m�5�m=9�S���[�EXv��Kl,�.DĚ��f�>8�^t��Em�/�؝kS��ȧ�-I��Lpw,"�z�ab��?���Nkq���d��V�e��������W`��!j�uB�7a�	#u: "}�@rT���搯P���\Û���ܿe�A/��7C�mj��4�+� ���e�.E��R��/Ͷ�Bm�;Wx�iv�%�2��@��N�h?M�l���+��8��Cy�i���M����( �/ �F���yE�V��[(��9��C,\�8u,1L�c�7�!ULR]��!�d�D�`�D긐�������
 �OHQpR�.��^K�����p�t��
sh�zU���#a�&��6d
�m5�,�r\���Y�  �f�v�.����E{ڿTd��Q��9E�}T�$�	�@��7�}�7Gݟ�xᮤ�#5��b`� ��Yv���vPU�D?���@yz��T(���fA�&�!?�]`�9���P��Tb^9����&�Dq%�\�ĞF���b+%}q��zz<{��V8�!&�g{e�[Y2��+��A��pl�����ҝ7ܢ[1h�{�p�#V�FA	!Ȱ��J7y���'�04������`9UVf?o�u�����x]�����21:P&Ļ�7T�CW ������A5)��zG��{k)%��]�Z2������Dw7�Z��A.�3J$�N�O:�6:�]��So�9���?��[J���@�x��}�sҨ�-#˘�Y�V�p�����O9�t��NH H�4d(�����A��Ϣ.�R1�m����闚���3���M��{�A3����M��^ڒ�~#����u��H�뢾<�H��ƫ7\�Ӂ���50g���Ӱ���z�0G�_ד�xR	!�B**�d��ߴM�yͱ��yf�8v�"�̙�c�q���,�TX􇓣̠��>�b�����?����]�L��tʜ�O@$���Pع���/�)�C�p%�-��3�z�T8��l��9DSdh��%-���r޷��t��}�l��2#������v,�5�ܪ���+���RA�A�@�tp5�E���j-HƧ]�ڀ►v�3w��SeAR{�@��������Ĥ��՘qȸ�Aҡ���)ib�&�;y�+#��s'��5&�����}�Md�~ᅯ�u��;�%��eܲ�, V���$�Bl,ϗ��n@��5�@��%�n8	�"����fV���<�C���8ꆁ����X���[�̛�zK���W�\�Up!qL�M]�'Y�̵�%'Շ��yߪZ����V.��$�&�-n�uh9�MO	����+SU@8��{2J�� ��A���܀��x�g4����U���`��B����z��g�f���8�-�waL���Ue�s:�ցa�!���ѷ ��>7	�o��8��،�V�VEQu�S���Tҝ�,��Wo��8r5�j9��'��mYہv�@%`O9Z�7]lye�\s5�Γ���^��=:7�W��H�A��k�{Q��4*�=���'`Yio�Ћ�J�H�g	I{�T̙"��*BrFh�m����^���*w/�p<\��`|��(b�!{��>^4���n�KD��F��s�ީ�&�;��,���N�l[�
�_��r�w���BHX+c�-��|B$$�����6�A�I`�2�9�S������~bY����9>~/�VFӢ#��rH8��� ftou4-0��%l� �'����m�מ��X2]��K��
��:��!0�ۧ�~�L���d�P?.�:��PV�h�����r�_%��ʓƜ�v���G�_��e�aS�9h���*B�0�`y;�{�ܟD A����f&���l��c��n����ֳ�w9s}���xtCط�>�u���$�59[#���D���98&iۛ�Y�!��f[Ay�<[_G� ,ѯ��\>��@��\S�r���zͳ�B P�ov�1����~��,�&����,��F�8s_�ꔩ��d5�!�Pm��h7���tQ��$YT�T������Rӻ��#ٯ ��f���h��u��.�ї�
R�"�<�]�/!2���������R3n�d��c�M�;��7p�rٳ.�w��	��Pk���wF�*��5ލ/��]���k�:I}��a�dv�c*7W��	S����;���ǭ��l��}*~M���c�)'�C�O�ϟC<�)�:�{��'�)W}�޺jѾ�z���B�����+ɇ_t)��g�~5�{?��>���l0��I�|��_��;�h��pL���Å�⎟P|�?��iJ�^D�S쎬��ׄ�?~8<B��7�*2a	�'��U��u�[��
3�~ل�Ug��Ka��d��ˬ�*�y,
�0�0��pl4�<��F.#0 8��d�`��>綕:;-fw;��0`��δ�3�^�-����zUrm��M尅!qr	]��	3�L,��؛�,g!�f��t*2u����B�֦i�f�B!t�h���j��(�+&_u->�*�RE�>y�3!�KW_$"6�f�BC���a6����$Ⱥ3�}`�F��w���i.,��X=Kc��� ��b� �綞���Qt�Q�ٌ`k
�f��=�:��|L��/�u�1~n#s{f_����jw�>���/ (�����,���AYzr�_�8&Mn�t�B{�|�;k(�V-�s�V�<�b�kG��+�H�d��3� 3'� *S����hr܉3$��1ϝ���t�'��#S�����Pԉ�
�ƧZ�gT�X	dM�pq���]��cO:�a5�[Fm�||�ir��R)UO]�+���:��	�N��"b�cn���}�l8&�U����&�A�9ޅ���D.=/��#s�vZ�o!�W�Ý���%���yA���`&��h���E���*�2�Q���қ�e��[��ͺ%��g�~�FI�;[8���{.��Q6��s���{dF䁋4&]�?��d��T$گ0�Յ�0�H!w9�B�_#	˶M
�$&1,���.����He�.���fhl���u��k��'U��v6y�+���� ;�Aҭ_��V�;��|���
����}��W����c~�s�߅�y+ G����9g��D��P�}=)	�՚r����{v����ش1H� �*�(�;#Q~ߋK�b����V���EHzxf�6�k�36��r@(��qci�ߧ)帻1�C	eĨ�J��b3Y�=�eX��=�Ҋfz���\�N�A̒"QD����T�x�)MEleUك��������-�z�����vV3>�.%���/Rp���~k���� O'oұ�S����l3r�	�,���sqT���'�|I���+bh�җjw�a� Z�[�J��XU�������ӎ��9���xh�V��!H
=�����ۅG\(�6�֦N�7�겈��@��̐�h��O�ߊ&-,���9Rt�ßa∦e��f��t�Ȁ2�E/oe[�)`��bC�9Z�� ��a��Ba�l��\��9��j��M��/�&�V�狠گ(8����������+����`F�G��
-(S���^��t��k���÷���n��8�G�r�Z\&�*Uwc2�)�C����z��W�#գ1L!ܣ�$?����X�\��m���/�����b�v3ȸA��s����M�+�J�Fp��W���8u}5��7+�m�C�Sb�<���D���н+Q㨑)j,=Ĝ��]�1�dD[n�E(C����͢��0�F���0���=i���W�}E	o|�CI��y���K{��� )�� i�Z��lw��
]Q��)�q���j�㈉Nƈ�߳N�f�u��{J�8��MQ6�*ݵ@~�|�Ph������f�"15c_���FG�[�vz�� ��G��PDQ83�	ӗ}�[
��
i{g
���h�%�pE֡��tQ��*������d�v:7RD�<���%�](.��Wac�xKU��=�f���AT�h�)V���sl}K�j���n��\qٱ�CoK�����v�;wt#��Qr~(�ӶV%�9�ti�Xxe�!J���� s�~��X�Atq�,Sf�1�2+��y�X�։�����L1�i��sXzv-��B���(D(�O�0� ھ�$�Yڻ�O4P�v<SjX.B�:վƊE�w,���6���57�5�f�Re	"���������7��Ő��,�iy�,����*Ϯ]]З�6�S�a<�E$9��k�Q��K�I��oS�%x���b);D`�����j��������V Q\�
5��Х�e��?\'1Uz���l�З����ry
j�M�/J������S�H.������_h������P�nWr�����yC^K�� w2��Ҵ�ҫ��� $?�t�����r���WR�g��HL���ڃx%:��{=hZ#�h�3�k���{rR���[�3��'?
�i[����5�~�^���j�"�:�l�,Hl]���ͨ;�}� nt�6�{�9��H���wG\j+P r�����H�ӣy�]7e�#ز�ĂVo�x�"{[��٦%7�t�V�S}�D�`�0o���0;�ߏʗ�v�S&^��]���t0��3^A���*�_�������1�B�ӃP�J��tcѓ@�������c��۷�V۶U�<Fq�CqrA�Z�`9���
���<XmE�{�Y�;t'������
r<�̉Ty�Qi��Uu�#ۀ��v�g���	g/h�#!W�޺�u}D�	p��N-�-���+
!a
u"Y�����a�O==�J���Ev��A�t=��/��Y��&�u�|���;[����rVWk�\��jY_;�P[��'�Q�񆡇�:��[�+>B_X��z3��'�G�yc�w?����*.�&$���08-�Y�{4S����ئ����b�Y��@ l�����ZA[$�s-/�S}�_f18ђ
x����k�P��b]����nl���iG��S:T������
�%�	��F��;����z�!ʉ�L�z�AM0����5'ݡ~��u{��j��S0��H������V��R���,�Go��,T�z�7� ��[���o������/���7��B6�*P�	q,�΁�&���h���l�`6�ge�o�V���]���t6�d�W1=���i���r,NPi)(��<�SWï� jMUZ-p���﷦�`��W
�ڥ ʫ]�ok��g�|��p�zG:ĺ��ȥe���ԗ/�I���>�����?$����g b&��4l�_��s2����z=M�=;�L���B��7dM,/c�՞�Ď���JT�r�Yra0~.ZTY\�^�J�!���L<����7�E�}ОB���"���f!g׎�3�fe�NGpL�i��y�&TN��Ɋ���e�ﱉP��4����Z�=a>�� �Ȼ��͟�"A�Yc�h3D���%$ΒPg���|P�]�~:�1��#��b�L�X�^��DnwXp�at�nY"�<���ҩ��t=���)�8��������6[[�Y�}�o7Q���J�շ��`TrT��n�%�Nn\ܾ�W����$k��Q��^n��KY*~�@\H�Zo�u^3A)$�/�"{���-I0�v���x�ӭ^k�f��2�4��N�bR�C[���Aix�ܥ��u���g�w����S>�4�*�ޒ "(jr���2��:vA�-[o�����4͎s���>�ѷ_�G�t��ǥ������4�qW�Q5�
�Pu�;=!�#pWߧ������Ma6�B-�{d�04˩����Uv),ϸ��Y� �+]���]�r�\�cقL��5����bre�l<�xuz<��[�"�,�ߑ�u�ƶ9��¡�:)����Dg肝9ի�6��F��KN��-ji��v��o�� ���a��!�`��^[U�Ck�����G��,z �L/"Y��6.�W�U�`4���a����~�Q��g��un��f��2J�h;Px�0	uXʎ��T����$��U	��ߺY_.��q���)�-&f
y��I�'~��>���k*����?��mk\��{�┺M��M
h�k�Z�`gWD�g`��� L�z�O��ޤ6�~q"S�Ȣ����Xΐ+�k`u7f��b���d4�S�C�ֱW-��Ĥ/ܘ�v����[���{>��ݸ�2W=5�L=)��ֺ�Z8rlGӪ����x�RΝFҳ�I6����lݭ�@���� ����E|>��mPe��{�_��~?BK���H��D$"���[_�eUڃ����� ^�29��r���C����}����ʞSם��F�ب/1ҖG�L�(@g��YM���$��ޙ�HO��~�,����W����Ҕ3���&<�튊H�I׊�`t6�K��9��
Z=��V������y�o$�-P�f��]�M�W�Vm�A��b���<}���P*��Ⴅ�1sf��r����>�KLf8Y� ��e̵�����oV{��B�BĤ��6=��oy�v���Q��#�[#���Q�@#���T^�ȁ��3�YO��D�^�v��YD�#n$�=���F�{c#��0}�@��tqzd��$+c;m]�݀������v9P9���ɋ�O����Ά�xe�����5sb���~I�iYe]d��ɂ��ڡ.0�`O5��v�%0{#�l�g��Cl�wd*/k=�j6u߅��ac�|v�([��lD8n��7�$f�"T�zڒ2w�>4�?�j&�H�HQ�+�u��S�j����&S*���O_e����ᆉU~!��Ǧ{� �
f�@$��0���Ϸ��%qє���u�
v6�I;qP��
9�
`ټu��, ��e8Ɵ��0�
�����r��m�ݲe����$)b�>R�HM��C���4��"�ɭaV4k�%�J�2���Ќ��� 3�
^fH����U�>׳.�P��t}:�a��`�f�`� ��l��"�ʦE���A.����*�׾��	��1�q� ��39,� �	���$�8]�s�,�Y�m�M*F��G7�b�T����N�����,Uo�>ؠd���C}�}
qK��l�x��C<>���\|V	��}t���Ƀ�H4�'�!�S��g@�?���L��)Ze�
f�=ư�K�}���~���P�Z�\���f߼{F��ؓ'�g�6v�_���'LOܽ�
;�ݛB�]�$�$�<���V���K-����4���v���Yz"�W<�\%�������~͑i�}е��7����8��R�Ó�5՘3K�|A�s����rHd��L��ݦ�a����ލ��)0��*!�|���Ţ�Y�cA��(�(�n�@y�\f#Ig�8n�Rs���5�hmFNB�t��?X�jA� �:F�}�٫Ql������%%��$zI͙��J$�����8�CW<Tq��H����FA�콭��m�	n�mS���&p����h��>���U�h�=��� xº*];�Ta�ϩn~�}����.2w5Z�Գ�s΂��	�?k�4�ͭC����b85��V�V5jdGa��Qrfd��ۦչ
���t�*�m�]�&��y������d����Q���%P�'N�P,d"Z��ZL,7�Y��W���6�)��m����b�∜��s\
fl��o����[֫�\@��r+��<;P3��5��c)��O���ؘ�wJ��:������C�lo�I����(1�`�ވ�H9��~��ިz�}��x��f�k��@���z�m3��,;��6���cä����� H޶���W��H��� �����$.�߮Ύ1GWRB�#�J��K��a��Odz2�:C7ފ��"X|���H��LC�C�Z�
:w�ͻ%�͌lD�VSBmSRK>��v ����PW|��V1o�����F0ʳطN"�l�eԫ:�_U��=HB�fѓJ��L-g��l�?=K�R�n\Ot)�L1���P�P��� �m���3U�y�",'s��N�O���2} �|`` ��.:������q�p/2���յ�I�Z����.���3e��6�K�������s�B50���n��I�,�?:s]C��tʌ~�T�W]v��h��'�^��bX�i�J!��r,�P��X���9��:2����vv>f�k�+�L~0�F
�.����o�*�_���}^6����i ig0'E��h�V[��K)`
ߒ��bm~N�`eZ0�Z��H�B����{4�[ޜ�
��nUT�h3ϓa���.���g=t���u�O�e.�}Ǽ
�y5��$"��1q|�H� S�7;1�q��*���.G��*����*AחY�S�&�R��D�-��<2x�g�L_`�*�`&6�)l��j���k����m	֩C@	��W���R*�~��<T�3c%�����C���Pw����e����6��o)w>��ۭ�!���`�3\�ľ�;e2Y���U��@U����ѥ��ǆX�}�)����I����X7��P�C����!{�U���ȜM��CB���\���zDd�*2LX�<b9FB=�3�Ϥ�f�sMȚ��og`��oI�Ť����P]���@�*�&(K.8�A���_�w:dI�q*{���U�K'�;+�׏�����������y9� �L� 3^�����+ !���\�?Ӂ�j*�C̕&�A�&f>���}VJ2��I@$�I���k躁����}�H�����	����{m��e�����n߫�S�e(���oӊ�B�F�� ���P�0��t��c%��o �?2ī����ʔ�n�`����|km���²��Dp�!�]�Q�t�ޑ��V��EWg�[�v�մ]�� R9y}zFĉOh/�ux�P�pd!���u�S�5��
���A�8|ώ�d~������,t����bk2̖����]^j&{���۝i��yC#�d��o�T�(mO�c�>�$q�=t�D��v�A>z��;�oX`ֈ��FaZ�u|,�R�����)g���܀񻟷m˕%�j|�YB����-b�/����GÕ�,W쥷�"-&q*T�ώ�����l�4z��E��#��롗���w�$7�r=¨��٦���Zww\'d� ^�S,v�#�"V��+"��+a��?�����������#�7}f\7�;ɽA5$�K�;0�K�����H���J�ԴEW��H^I���Jգt�Ƚ�^��ŷ��{�J?�f��1�E���9�a��O��������+�o[���B�t7��U�t�G	`�L����h�[BIS��K �S���Y��
\��?��;�L�ji�暄���'�|}�Qݩ�/?ϛ*�Y���7I�i�bǯ�U����z�g�5�~v�#�Ő�������F{`���i�!�5�g�C������ՠs�B���&$V�Ȯ�c?F��\��o#$(F}�1�Jakq�Z���3{��4��ȴ_YM`�3��O
>L���J�c�~��9�p��w�h�_�PX�C�1H�0��Y�g���HKyu	93��Oe>��s`~�S/Ij
i�g�m�a
�aɽ���x���P^������a�yTt 蜲�uYf�����?5&�4��O��[#u�M�о�#���6&��<o��0��o��Ép� U���ү �<m�C6�M�^ڠi��g��5��ҟ͂0�����O��"��T�E"K!T�$��� ���޳ �?��k�p�YnQ Z�D���:3t��x�$:		!j�~��?}Q����8i�6�R�h܌��	�����c�!�@��:����qL��W�3
I8��s
��x���v��Y����	)JB//��z&�+��5J��.D��:
��8����	�	NDV���B�I4���Γ !�u�	�-���Η�@�J[A��V�M� 2�A�67��c�DF��<�Gi�w��fe��r|�J͑�ԧ�����<�4#`�x���	�a�[�B��֚g��ߌW��~�h�5��s� �o5l�����4w��A�a�B���Y["�/T�.�Ԙ��*�"=O�@�5��n`ܰ�\��yZ!p�d£���ǳ~qFngZ|$��>��h*D���L��Y�(���Dϴȗ�BUS��2;��w��U¤�jD�+�����s��W ]��;!O�	s#Q���#k��=g�ch�|`��� &���6�����)~�SG�󋧿�4�qBe�ƀr�1�r��~�W�97��B�%ڧ�6^�#2]�~/�1�s���ɫaIcȤ�T�c0@*���4��Ȅ%�b=��T'�C�[ZF��!�ωlJֽ����@?�l�n���v��Q��u-\��c���Y��;2[V�B��me7/ͽ[3 {�˦˧v@������{f���mR��K��8��[`��1�6�-���OB�7�]���O\���!+�,�V3h��~H�Ψ��fB�?����{C�ߚ��o�<�LanĜ���%��dUl<i���l-��%)T��CB�&�e�5!�о��_;@V��=՟٢1�R���<��m4�D��8"ݧ� vr�t� ���-n큧�c����W3�E?=�������;���v�=��)m� !Zq[@����A:M��H��P��;�9���M���՞�Em�I���Q\�����@��lb��߷+�B�["��=&�]���h)R��eV4k��q�m|t��h����bwml����X���u�b(�$�-�6Z��pћV�Թ�տ�#���܈��d<�,���l�	�'4�g� <�>�I��E��!<�LWƫYV)��d��y��쉢
��5+���!\A��Q'0���r�N��U<��9��>���{��#9���aV���������ǻZ��X&��,X��ю��W>����^�Z|��NFN�$��X�NHe f-��੡PҸ���<QR"=����1j�� $��D����X�+ԅ��2#�\r��>]63LFX��q5�X����"�c�A�a��a~��}F������9QRG���Ѥ:�^i���l�7��_~U�tQ~;q[Ϙ����_����Zr�d�)�_sƸL�Jc��*gt�L��|��po���� �R���GHw�.~��x}i>��~�E���.�ڹ+p��cbI�i���
Z����6[��w���U=��Wֳ��/��
?��*^P��2ۭ�r��.����f���X�?��}\����ְ�n�obGaX���a�B��U�k�G~�xYI�:_�6���Vv֦�~��G惿m�f���b�frh�Q	`�X�b$vX�"fغʖ��1�˜��s3�˸YAR�cj���\Q��@�P�QN���0�~W�c�q��*�N�7�!��qA��b"2 \g��� ��a"� o;��gw���������b����b7W��gCb00b����z�����#9���Ü5���JER�'��p�(j����QJz�i�2�,�b��Q@]���߿D��ڊ�l,4!4�n>(b3�_���P,Tӕ�6� ��Q�c����*>k{s��A�HT�l�m�^��7S>!���R1�q�gh��������P9i~=s�rv^ρ�y|�iz�*ܵ���bh�bY�[ZC�OU����V��77��g���n�F�?���(ز��'h��U�H�j��<"�O����=�&�#��>�|$ ��d��!/�Q~�vC���ܮ��U�22R���_D�� V*�.\�ڏ�	�Z�ӔS�s/��7�q���4-�=�4�}wU9��Aa�i˪R -ux�<�S��a�yce^�4;�]�x�P����g����-=urn�n������*�ꪉ	<
7h{h��S8��4@6z�z���^S}�e�C���޸�����e8F֡��BB�T�׳"��0���ʡ��i�1q1!�<x���������������:�g���|�ۦ"Jl-#S# �F���e��b�nw�F�x����)#6G۪QיVGH�����YRʄu���I����}�iD��p�IP�\Nӗ��c�F����>���av�0Z��4{	�	,�X�k�wV�~Z��d��z��	�m�������1��)�!��}�g�o�cZ������)K�
/c���Q&������髡θ]F�u��C-둀@��������	����p�>�4��kW�L�j&+�b⋑Al�f��,��A���0�+�#�@�]U�u�����E���fϽ��$IU�2� �YK�L��4���T�Z�����$��ؓ���9��V�a�ç�4�Gf�zW��_ ���8As_�ȑL��8��5h��l�v�#���Q��@�Ȫ����;M���ײ1��g�h�Z��^ʉ�{9{,���ށՉ:d=���mh�X���@.�d���Dj4�D5�
���\�5�׼�����2�#�{A�2����UC��d���ӓv���So�t��5����-��QԠv����z�c��XA��;ǲ�F|^Jo3.mY��{�?��-��e�P�'�˧�z���C���jD��0�l���Wy�%�3�! G��k��m��0s�'AH:�Q����7��kn~�8_F�J�`ү�7�+{AըG�`��F-����Z��B<>����e�<���ϽA��GU��l~��QSD���כ�KU��7�t�KzՑ%������2Ƨ�x�5e�x,��?��<l>�!�;�U�0��h>�$�C�*�W�m!z)ڂ�ǈ���
x�J%4�;-|�-���~���zT�Ĥ� U�@�9��M
됶+K݉�\gE�
N��[�{5\dL#""ˡ��I�]s��n�)��ॸ��м��r�q4^�o��� �UH�`	3����'يQ`��H��S!L�#GON~����My���2��܃�HE
��yUC@�T�SM���������&]�|Ҡj�~���k�8�җ�z�0B� WaC|�~��ff�>��{HF��E�@B�P&1>��l/�S��ǵ����eh����â7� ��z�M�y�74���F���GtO��z}�(֨���%q�0��\��8�	�?>�"<z6����Un���Ha���8����Qҥ8sʷJ
���i���Q���/ƤC�S`kv�ԍ?H��h� ��ӚCl��2ʧ��ҹ��H�n��y�����.)f/����M'H3���{��9�)�1s���(�G`�����0]d��g�OX�E��D
�����4�W�q>r9;IUzI�v�3�3��ǁK&՗�f���2ݜ�����y���vms��`'�B���F�$1*��h7I�gM�Y�ךK�}�:�vq�'e�in!J�GLl�k�&yӛ�$�N��`w;,�����l��ߗrz#�mH��)��ݺ^�T��΅h0Cr;�#8{UR���<gO˴�bUXH➕L�v���-`��!���
H����Q3|���ȥ��RX"=[B%l���Iam؄l�W�	{�L�R�g4�BF�P�J�ү0(Ѳ7�H0Qw��i;�0ʹ����Uֆ*�*��Xz�*ؚ铳 eif2#��  P�jw;�QY��Fuaសi�1�%S2�$�WZ��mG`q��Tt��*���&
m�c+��+��#�h�_����>� �SjX�RS�i��Gnl����t��ꍇ��A�:���H�{b�Q������ήb����`�:X��R3T�]��1��J�i��o /�������_�{Wߊ��Ӊ �����դy��8��1��5 ��	3r�-C[�W�SI?�\r<q���g����0"��GF`(HNKXֻ����u;r1g���zO�p��zxL�Sj�W�K�}�\�/4�&=���t�[��@�燖�K��;�gO�ۑY��u��P���x��x��E���`[���]<Y

&�zR5o�z1Ph退�<wi��g���v�1�+��4!RMx����H���Gu�OG˖"�2�?��j�ҽ��l�58G�,G��f����Z�Y������h�9�Y�]~^�&z�)'�.�/�OۻgD�r�-���c�@&��oEʞ�^YZ�
�uv�Nc;��j����Εý�3���9�}/B_cB|��f���)g�D�0�x=Ho��v���F��d$r���8�����]5�4>P������F���Nb������1,6)X��$�[�/����S�o�)�W1�`�'it�]vwe��E�6���.��8�Ti[��{׍G) �v��E3NNA)��1#��!a���9���87�~V_+N!�]��#VP�p��Qxl��2ɷ[��Ru	y�&#�����t�p#/>���J�Xt%��5<�_&A\���aQ�F��F!O/=��el/�6o�4�$�e.�,�:���!&�c`�`��9j�9`6�>�)�. �Rx�+�R�Ԕ����;���
d�:�Z,���ެ��_�BR�d�:+7�iAi������+_�ZIA���b/�,�rkP��1P�k5F["���Bt�y���be��.�p�s�Y����b]e���$wC�>�1,���Q���!F</���<ݸ0L0��#�		*����!ۙq�Xk��(��0Y�剛@ِ��o* �G�s~ԧ!��a�_���Fq�@m��^�kWѬ���H�� W9pdR�Ʌ�E�>�G�P�l��sihs}��E�_6�0�$�2Ԝz���K�}�J�{!��z���=G.ߩ�Z�2B�+R޼�ʖ���`'����
%�=	�)e��Pὣt��rs�0�B��t�b;�jg�����<SG�+5'�#��cʧRh�g�(���%�L���4��P�_���T���L��ƺ(��J�]EM{��vZ5�t߶�`8x�Z-u\ ��Jԁ�0����y��nh�8���ɓ�>������=�V�5t ����4���깼�syսo^6jX��W�� �r�i>�������^�ryzv28�r�r���������J�o�81Q{�kd@E^�jr2�@�§��pu���1􀕐@HB�F0��b'�v��|:��SD�KY��G��3:�@Z�2 ���Z�X����@LP�@�`��$o(L��kp����bD�"�0��xul7�x~�X�H�\�0�=���VT\�ּͯJU����~i鶼~�m�;��|��6%�v��J��Ո��K���7ħ��#��R A�|v�l�ό�c�P.�&+��m����2�ꉰ����D0l��zI1O�2�T�wmH�ߡR�'�pp�@�YA�P�� 	7}e'[I����`�HF���x�]��|!m4<�uB��X ���~���َ����V �z�Csx��|���.K�^��	qhZGd@g�w�ήq�)��lAD������pʹ}�?�U���J �f�l0*ξ�q�Z�|R�pu��C�Fk`s�I�}��#��^��K�21R���$���~������BD���M�_g�@�~#u97�w�|�PP�>A@�:ߡ�mj��`A�ͳݐ�	NBc?�K��m������<�e�f_���f�R��G ST>��9��j�?Po?;�*�;A*?vV�S	z������Mp- �"�Y��>RUlB�u6*d�ʙ2�mb��%��]�=�s�$�	���y+���̧H?d�f?{Ve-fEN|_�4h�޽�B��/�D������/�����8��#Yڍ�K^�(����T�G���1�L��	�6�w�B��JcZ»=�-H�;�4%dt�T%����P0�<�}N-)}r�ۂԂn.7~���u*N�U��OI����rWh�b�M��!`����{ж]v�5T$JE]�*�LXx$���J������,_nk9f��S_E3:�H���࠽���`��dp���"�A�Mm��6'��n�'��i�SDX�P�w�$�9�D�<^��������xm�%��avk&9 ���[ShyP�;$"tSO�u�Sli���/'ޣ�� V�ONG��Y{{�V��f��*�vOܞ��R45�T&�)6{�l��奃����8����'a:�h�����	��3�U(�44��S����,n�J�H�!I�b�lz�Љ���¬J�1���W򐀶��α'�Ɵ(��X�%�V=�B��Y`�_�2l�
_�I� � � �K�a�\�2��"O�E��槎2���)IRI�-��l)l��?)��9�Ր�����0�}���8����\����M^�Gctݖ�ⅣT��ł{\��H�����WA&J��OQ�IA�����E<�Ġ�L��~ܛˠG��M.�_0X� �wY0��6�V~�-�,�\�b�I7������'�� <�����V�]���6��3��s���'�������ja����%���
q�)�+Ħ8ŷ��$!���>W��k��d,\��m�d'�k"ec<[2�$I��ǣ��d�R,�i6q�I�Y�MEi�ήK��P��x���.w<�x�l% %l�:k��Zܠ4d||j���eAH��0�0y�g4	P�1i�I��#���ɉ�x��;��J�ۥ9�Bi*���i	�+.,*�B����e7��qS׈�� x�-xe�E��L_�w����_�Lٲ.O�X��f���������� ,�� �4�~֗W;ۀ��6����K����=u�&,�k�3OS�"b��x�Z�<���5"�����\s�m֨x��g��&�2�����nD�8��$�R�(��u�=3�B����b�(� ��\d�>���4kO�O(>��$�1��$:��?����O� ��J&�3oS|�@�T��M(؆�o�y���=����n��][�)��6�:B��px�C�]X�-{�~o$�ɺ���I����+eI��F�xv���_���쬂5�|k|�R%B{c|T�4�?�R���V��_�s'*xB�v������������.&s�PcVb,�7^U�|�����!*�L�-fb���»��	�ؼ̬Zx���$��v`�0�"�˝.���Ӡ�;�ꉰT���x\�yK3|2'T"�1�.�����&I�0uӎyC)�yϴ��	~ �E��*$��(�9ġ�f���.��0.�(�W�[��5츾z����be�q�N��ZQ�M�y�B��I*[�Ի\1u��ހ�*���$�M�����|���NL𛋛a�=�$ZQ��^�g{�g�5�ٚVtѫ2�ˣK`��U��Qu\߽�E|�F���S�o~6���c��@m����v؝T�J�G�oB.��1�;�H�����ȥ��.���e����m����Z**X�<�VH3�8�Ӣ̣��z#�g��d�U ?�P�4��Մ<;K�v]`�i��5�b��GB3���6�10`-���s��\�OT/��B�6�B4S
:���K=��ܿl�Ć���/ĭ,�Ʋ�>�#n�V����&	D3
��'bM��l�u��kjq���Q�2���+����yI�0Wd�U�ռ�|��X��t?׬�h��<U���i�Y�&�OΌ����t��-���̎Z�.3 L�� �i���8�@�=Ytō�s� v1=�)����P�g�ɪ����fMI����
F�J�ù�ի�m&g����Qv�Ġ.b�成�9~����(ȧͲtp
�S��+y���I�FЋN+m����bs�e���T�~�����Z4r#.3�/,7K���Q`���?b����'�H�)<��%)$��w�߀� O��WVR����"]t�;lvЄ��E9a�h�=ر��.��i��36܅%����J�aEgto�_�VZߨ<|���GI�[ț�7�o%~8�� 7��T�fs��ti���,)�Ò�����j��*�WA�t`����~K�8x�*v?��D�n;smfE��H�^bgu���;����2���A7M{H�=5��Oj��&-[�3�iF�1%���Ls�Vg�Z����Z�?Xj�2���v �0�.��]�c��J<�W�%�ӠB
i!����yݭ?�����PPoHFk��-�I���t�-+��4ń8���b��K+O����P�kraj�}tRI�D��ݳ���'��N@~�"�?���u�ڼMa����KP��Bn�\jA.�ȟT�@같?-,�2f)pZ�d��ΈO���R/�5Z�ѓ�2����[��xCDN�lG����nQ0v�7Yp��HaQ �_r� f��#�������SAo��Z�`K��uNc��=�<Ώ��8?=��ه<ͿՅ�� !6lڅ)l�_b8�gx�QJ�b�oR*��@[��`!�S�:'&slH��	Y������,�U�$����'w�^5|�r��>Ů�ƋCgT�{pgH�&=]t�#�xi�T��y�u��s��i5�*���@�`��FI�k!�;-���1/*�P�
���	��L7�7�� ���0c������;�&Pf+L��s�@K=m"f�ĕ�"L�<�Q�.U&������ʓ���Y�'R'Q�[)�t8{ߏ�������Ԓ��(��14�G2��y^3��^�FS���Ʒ,C4������Ґ�
�,����l�@o�ERb�~�N!����C��}/P�ԭ�*�@���06g�������� �C��J��q�#pL
�m�cɉ������p���M�a�A6��^�P�j��!�2����ޞ�:+7�<d�yf8�>dTK6�=��wl
�����B�H�ZW�cLo3O.êa�{��sű� ���D��-2��$\��a��T�I�a��l�@���[ě�b��9�w�Ҷ��� �r��t���Ǧ����fn����m���n�����x�Ӡs��P4B���[��bs1Ŝ�#��]X�Սw"x]7b�|��~��A�<`��*����<���j��f�E7������VV(�g�L��bbg���Т=6�#�E1x��w�O�%��Ǹ�8�6ʙrD��k�fߛ�0�~�g*��\u���S��-�w�B�����>�0��S;g��cc�Ӈ���ay��2k���2N�91�[O���X�Py���Dջ�ǘ:�z)\8^�#��bfVKB� &A��s�5D�M�Ia��2�D{/�\_��&�nZ	�e�	�.��}�3*>��Y��g="z}��~bs�+�j.xC<�1 �������Gh���J�%��$�[����|�
A�#�Ǒ��6W9�
crB��n�rý���a�R���1h2�8g�H�趤\��K�� [�1�%l����C9����k���(O�8���ߐ(R_�LqQ�:�%v�a����=f�V��ګb�����0F��>^�#��6J5���u�͌�q�Z�2�L���1�߿?z��A�U�˙\��O�0�gk�G�|�$��P�f��\�����¨4|�c��b�V�xL��}��@4��Oᩱ�BE�6�����? �;(`G7����}���=įݱ��N����W&��'y��4���Z� �����a���_1f%_�e;�gi@��t��(�Z�� �Є�[�uT!A���{XJ�t��Yh���pE���mVA2�;�َO�2#^I�D��U��a������+PTD������?��f�u�9���%��yMGҩ���>|#�y�9�t�4�nh���>'�jL<��1�Wpx_΂��_�?��Ȼ�LDi������E#��<����� ��O4z�sm�e-��t���"��#��E3�����S�n��奆Z{"A=��ڞ�*_˦t��.w���	0m���j{햆�q���%O=�u�Р�;������	�ذ{���Soo��P�C�:9xm�g�10U�51��J�7I`ٻʡˆn�%p�[�G8c��1�.���P|��|������{?�gw�-0��ߕPȋ����Rj���v�r--j���E�L�����i��p��BPhEZw �Iq�mo�5k����lX�L�8���x(�܈�~��Y����}.����
�O�sQ�`4�xx!8|UN��L�L��H8^k��W~�}�Tyh�0 -�����QhcH�FJ�m]6��w�Ƅ������&?�E��n��*#�C���#�U+�pk�_�2ztw�&���]ěX�#c��`�zo���H��tD�[���\2���U�艦��gKr�ye	2��B�Q��pB���1�NE�io�83�L�Ɯ��R��^�:`����������zټP��qD��豲-�?u�^`�ޫ���|�H-�>�P���m��Y��J��7�֨�K�l����(9(���~�|b͒G�~�X6�@-u�B�� �[B�5�Nˠq�`��>GW����-���ٟn��;�\�>V3#+�>���u��%��3�[�������V� Yb�No�9�+)49�>X�9���E��p<��M*4ն�c/h�~�b��o�7��6��L�h"��d{����߿��,uC��p3��/���5��}��v���b�l�h��{�Jӄ��o���=�f����	dھ�?��^�c����K����UE;}��.�L_�F��KA������Ӎ0��¼S��_b�[��	�	��;��uN��fC~�Nl��/���O���8sYr�(��R��h�M<Y�5 �L��dy�IO˚��~2`�~?�� ��N7�U�J�4ě۶��bMr�!�mN)+6M����9Y���H�Պ��:a�#��>*~�b��%4�d$-謈|����H�����K`����jʨ���e3F�֘͸��l��('�e"	�I�Lѩ���Q7П�Rs#a�M)�G�N�	<jg�˯�օ~~*ۏM�2�?���b^��U���os�r�-drL�vױ����:�5���s�2�>ڼ�Ɗ'.����$ ���*�'2��x[�L;,��c�V4Tə��A)ld7�\TӨ ���Q@�s�Pa��|�����\���q�' �e�d�P}@ ��s9�N��u-g������!��XaFô5�S�:�0@��伥e?�5`f="�X�dV�ۆw�8'�L;i;5'BYvӦ���������R�kT������m�|��h'� [B�z-+��b�Ұ��Y�V��êkdD|F%�m-�!Z��|08���O��ylk�fn@��ݨ�����ށ�>Oz�B9;8��j�
��N��R�1���ʽV�i��&�}D�XѪm����*�A���͐���N���Ï�������8�B�!\#zE���H|i-tm�lV��+�KF�E���'0���i(���&��"�D�-��E�Ix���6T\g;׫ ߼��G�Z���OL�*�ȮD_Bs8�.��nC��a��[�I�$d� \1����9hU|�hw�j�G���D5Y~�q��cK�lT�E��Tڏ�N��/=��>K�I�YbG��Z���'qN���\�+�\Rҙ(?כ���?"Y���ǦE��Ds弔����6=��ⷬ���1^���Cf7�;��E�T8	�s��5��Ń��Ā�-�����xԁ�,=��=��ئTר����a���FE��[v½[��;�і�z,ؔ���y�	��$��񮤬%�o�O�a�xҌ��4�t���is�#�>�;�Q��C�d���l��o�:k�
c���b��͢}H�%*ˌڃ�L�珇C�{`cuG[�P��j��>Cl���s����� z�i����[=�&��k��+�G�.�|���+?�7GMF���;]t9։&��g�{N��w1�R�Ꮏؓ������vf���gD�pa� ����&l]yKxR�"�i��odx_��k�8L�h'���y9C���zJ�s:�B�[G�YQ�g�2[}Ӈ����� �2 ɢn�����0�
���-W�c�x�!Q�L�T�F�f���=����,�h����	��T��Rw-��|��Sv�%$ا ��-��B��Q�7n.ú��	��}NK*������E���a:������.����9&��UJ���Q�4�/���Hr�$�S�sh0e�F��b�)�GMDL_�C2�����Lʾdo;w��&V07Cp�{�]�ϯ�F�Yr� �
V��E ��1�Zg��Y,�E'��5/G�i+n��;�ݵw?��pI}*d���	|񉫼Ή�Q�E�u����}!G��
?�X!Y<F�c=��O�Sdմ�3A_�7������O�$�X����3�Sw������\�����c��vM=�H�< Y�q�	��!�᾽ֱ�-�,���=7��'� t#5��[c|��"�e�]�ua�Zn��#�H��6���:?�(�D��kmotc���Rn�u[��UZ�z���X�V��^��bfx��\D��O�9^.,��-̌�,BgK��.GB���.td��.�?����-ܳs(t���V�Z�14*���t�}	%��N�`���6�,!~BFJ�;/:�=�8 m_�>U�HoZ����~yDQV��C&{T��f��2����
�焮䄫^�N��,��
X�rh.��Me���_+���ђd˥��Ěw���+�쐺�r�YP�82�b�WHz�>�}@ e{��H����=���x��`U���	t.ӂ���B�a0�|����t��-��]����^��j.���4�ө��b��&�(����+�����ϔ��
=��@K�x�1#YB�*�y�'r��xC��`��*���k���dJD��,\�k��g��J�=��r�("�đoy�?�K�6�W?�d�e@�"8���uPncۢ�Y��L�b֏&|W�)�V�Td�O���g���_�
��v~qfԀ���h� _���Q�W�4���Y��nN >��:2H�Z���ܭ 2+h:�М8Dߎ~��_=ןo+�/� ���%�U[tz�pVbZ���Ot�[u�(�[�A�FB�$h�M�Nq�G);}�|a����Ey}�q�K�,����
�����q��I�W0����K�[G]?��O ჵPt�3z�$�^��~#���aZvW'�@g�^�'�z����*i����<�B�ŷ���}:�&��@	w�WNT�N��I������	��J0:�ś1��'�!8!�ŗ�YJ�-�e�W*�4��bZ��Mh�}�[^9�7q��-2JK�M�����`0�Iv�p�0@������Kv=!���a4Ȃ�#�p��(��[���o֚~f3I0�czY�ɐ����*��i�;���hV��ʽs����3pZ�_�}����'�5S[����s��(�,b�[��Owk?�b�?��p5H"�x��0n����;���v�ƈ�F�M���E>mcd��g�sI�iV�|��aw[�%��LoG��<�|ΩS�T�gy��x��K�dGI�N����v�@ُ��d_�]���Ťy�x�)x�6��`k|�.D�	?�؞O �>��F��TTs>��7#���8���t�8{��1��ȒCjg�^h�u1��n���`��^�OBM-�b�)i��oy7K�����6,�Q���?��&�9�;�ϡ-k�o7�Z�E}����T؊��V.�3V+���`�%�W�\���V�	|[�Р��~���̭&�i/:�2Ӹ^�?�8�g��̍+�?�c*����$��_,h���h��N`.�;�ǲ׌� �>��˞�\KO9��n�7��)�D�!�O��iE�'6���J�FϮT{^H���5;_m/>�m0�$�V��p�3o��jN0XB�k1�P$�)cQ�zP���y<2�p����W�}�=��{zǤ�o�`�K�9�MW$E��+�~��0�cZ�4�YJ��q�Yr�}��r&�����*B*.Β�ؐ/B�9I���]��p�(qR�o��<��'!G4����`���b��{c��"��g�C��`4�j���6yaq��~&�����J�FM/��k��2
��߯��3wѯ���"�-jjH���S7-���!:�&T�xml�\]�����a��-��8�7B���V�~�Z�͘[v�f7<�c��F}���Z#�)&i��o�7{���1f��XP䆌� �!���[��H�f�}�;��Ty��T�=l��-߬�6�l��-j(n��3�Q	�ɯF.��Q5���� ����m�"n�M�U3�hv\��������o�t�?�y�`�5��wk��V>�����j|��8~�x���R~��vXX9"曡�#�0_E�"X ���2�4��_���5������-�	����}$Gp��<������X��ցڙ��l�������񆳭�f�����$�ա���YNo|բ T0(ue�V~�Z)}Zp֙��9��,e��6����!��B\�}��O.t�[���z��Sd��²_��SŴS�ڃޫԥy/҉��n���o}�6�FH���O�,`��6(�׽����K3��틇:n����0m�N���<�|�PL��"t��!/�zPV�����I��a��c�f�X ��/4�崹�̜��/-C�!{!O�U���EZ�DL��f�`���b+��6����$�Uǉ1������ٔ�
��t�<1`!��z�~2j��Oel'9��Ui�"82�[�J��K@�/��{���FA�ƑC��T�n� ա����]�;��䯕4[�!�q(`����w��C�&u�3�]�d�O@x��^+8�ھ.�N��B-]�F�^k�����5�3~�����K�Ky�T i��a�3周�N:���G�����-��9��d.��ȼ'�Ĉ`k&t�<���_lԂn�l�$�J3��I-�tm�^���،Vf�^��$o�*�3��k:HtF�C7s�;��V��iY
GvvA�g������>G��.�Tz��Kip��̅uriU`u�A�����Ѿ-fϰI`��Y@^c�m�A��p��e��8~�j��Y5��L(�~��FԊ�~*���(��?=N�\����&t/�fNJV��z� tQm5a�bǐ��1ePDೀ�B�ws�!ܭ��}�x�1o���jI��`ڀJq����Se��0h.^������	n9����[�P�W��{�u6��K�_~Wƒ�S���v� N����8I�ť����j���EQ�3�4f���xt_�(j�%ax3����5�>9 ؖ{��<Hc\�M#���eɆ�F18A�"�F��{�~�R@j1dfZ>�y/�8���],���%���-G(� �,��s�`��hv/\���n�0��EqQf��m����]����2��/L;1ɸ�?��T�(�0`��w+�gz���G4,[���r�X1�J"@3����vt���A �#�,%ݝS�f����7l�l�n�C�����oΥ���R��1���h���T�S�0�Vw5;�5�&�*P۲���&ԲR�O�um׫�L�@iQp���G�J��x_�e��q-�:�٢r����/^0�Qq��qu�� �|��pm�G��W(xd�xd}	�g�`������"ɉ�������<囐��Q���$�/"�Ge�q|�{V�-|�f�A�g�>�e�'��Q�$@/�d����I�gX�+b�y�η�S���D���~_CNѧ�s-�Me�r�BW�/�}��|�N-�Q8�2��@1�{E�J.В�[/U��6�q�ƺ��F]<����JkMP9�go����i���\[�.����Lwe�NƊ�
���|�h�x���6��Eclx�V�/�~�niq�IT�2�f�W:x�"�:bb��>�C�6+�	��@i헹�D�{��+ ���Y`*)�S��?�TE�fA^����%��
o�<X!&�<����X�D��`��,���m�5�C����[w�L �<�mK�.LUn�`=$i�t�%5:��Y�z7�/1kX�9]/K��uB�i��\?eSF�"���$Y��N@1���Zp$�������!���^�	���2�H%.���͜��i��[�y�&�=��Z�sأB����[�K>�JJ�β�H�1o-�2�����<
��|-��9qx����F����FU�o�gM�tQ��_#��@}U���=��q8���N
��X�wV�u�G���>��kC{����Z"��~@���d~*Ʋ~{���	ydr����rS��T�q-�G݉�m���މ1e��xx�n�V7*O�X��#���iܷ��y�a��،� гվy�mp�ݮ��.�o>�6�:�'EZ�S!�ݹ��S1멷WF�V�1�u���
���V�P�ͅ.+���d���O=,�D*�A%L.fȖ��mrDJ�ItG�W�� M߉��z�`�ؼ`��ڱ[� �%x�������k�{Qx��J/��Ǘ��U��+w7z9��x��;Tq��e�9[��7&��}�Z]书9-��-�mSI�t��A������oL��B��Pb?���fi�M@ӑI4���^o�,S�D�f]~��Yf�.�C�`� ��+(���}/Crx�(B��vD����ѫrpج�����|�->7�/H��7g�m� �:4����T6q���W[6٧ �"�.�],I-�<9H��z��*������e:w?�7�ELy��Uk���O�s��Z��uJEo�(!���-警�Vȩ�Su��߬>@�lU�ߣ̢y+��l.F+�m����y�W� �g_S���b�M���c���򕕕���E,��`�G19ѽH����(E�b��I��j��mw���Ih��������چ��mdC����1��z���ji'n�Cq��Z� �׫�<�0��tB;��oE�3�нh���ܱDK0���lR�ޢ P��R��g��x80 ��m4��ݫ&�ɇ���่�?��Ƽ�"��;$�M�Pp�V{��67�M6���0�l�&��P)�$���y��DJD2�Xi����'w���(�v�:�BN����*���F��c���6��ۿ�G��a���9ިwl�Q
��XBm����lt;��0�p'�N^H3�����k?��?��b[���د=�nTґ���K��
�ΝO��ڏ:C٫fi�c^ͳ�ۻ�w�?0��N�q�x0v#o�+ZdrSĸ�FV�G�����;(�Ҏ�Aq�L��㜒dv�!_�U4���\��ّ�=���5Ot�(��>x�����0ܢ��w��W]�:�!>l0 Ŝ$���X�\K��w�}��67�_��kw��%9�@��a1�e��ީN�\�Wu�zՈAb��IE�v���哬�a�Uz�*����	����_R����9��bhT�8l�,Re�4��q���-i�--��b�m��%�ێ�b��V�ta%
�Ad��G2b8u0�B���ـ�օiu���VӸ%�i�'H2�H0{�:��*���������|�)�O�$r������pt%X����A����Q`�U_���w�g�ㄣh)ᖍ-e#`Y� �R�!�Y=\�`���%�yU;�7˛0%re����4�r�H�A�7xB���+7e�$�AO�Y�szM�k��#�A)� �p�9J��4N?U�Fڼ����.�Z�+	�]�C�/�9`b<ݢ�9�%�{m��Q�( ��/�k<�ki�?��^��{��}��{�,Z���tӐz����ݣaŸU�Nӷ����&��X�A�P��Eu��`/�%��i��]��ke��Kը����r���H��H��=����bJ���T[��2���v�ES3�X�����/D�����$&�_��S!����u ���Ik����������Ƣ������w�nHxۧ���È�r��Ʊb����3%���g������{��K{>Po��7]}�l`W�����G���v!����A��%��N�1k�aޢ߲����;��x��u43j�� ۭC�g5b��-��C�a��R�;_��j;q�3��]�RF'y�ʭ��X�Ҋ4��r /6�F)�{F�Y���ִ�Ü��n�������FUo��л�2��=݅>�^kcC�{h��ɜDyD���. ���J��&,!Q�w�]�Q�0�k���6�̙+Kƫp��6��N��b%+�}i����/T��ϺZ{�b�
�8�3��h�*P�uˤ=]/jh`և�..�i��*�w~�?�6[�|��h����6_��=ǋ[�+2`��ƒ��ࡇ�'���;Wв`y'8�P���.�X����p�l6y�r������>nq"�P�/���O����� ����q�2Bj@��A9�׆f}�.n=3x%2'O�ֵ"p==�#05�L�!��q��|M,x���|ٓ�r�
��������^͈>���؂�(���]ƃe�ɏ:UL	#V�H�`�k��(��3�
��@��7U|w�L�{�8��Qs
WCaqn��!'�mCaC�p!�]i���E⁲�b�g_-c�����.���^Y��\�b�raĻf��'�5�{tĨ��	믱\�q9�Hf+	l��ҋ�}���
�CM���:+~�/�o�` !=RThi�����ʀ�H07;��+����*j�ղ��J����1%n�?���-�$�D�H2�6
QUY쟁	�dO�_������|i�?�V��c��/���mH�|!���>'�׻���5�j9Mz��[�H���Gα)�� �[�_�>T��T|��횂U R���E��A&�C��#L�M�Wx�;��i깶��i�N�C��!!�g�&$]:��
}D�5��#�֞��?21�ݪ�y��.�����}�e��''<��`Og3ĸ;Y"Zt>Kf'�1�h����ٷ�	:L[����AN{2�x��8�t��x��dƥ�z�iN��H�~5Ti_5��_�:���V�#Z�m9C������ןL��x���W���Y��A�%16I�J+���ʟ��x��_uXP�g��f���8�(��1�2*fe�G�
U��($���(_{4�;1�6�����x)�#���<� ���) 6�7���E*`�p)�����c1,���˸�0�B�Q���y?b��������G`��=�S[eU`/�?�0^���!�����f�¡l��atS�mӽ(AR��xaY��1`�U��_<��\��n��6�Z����tk�ҵ({����D�E�8j�P��{��&C�������JO����Dhn�s��X#1��ᣮ�%\ט$�b�K-}�:@�����d i9.LU*$�9��R5����l!!����|Ģ#[A�eЄ������>cKk����^l�I�\�D��x�ח�໙��z6w>ܢq�?�R�2}d�Q���y���w��T��3�$aޅ�[H��N��`hA��칪��.��� �*M��8�Bv��~����Y��{_
ᇾ`^�����E�����>>sQ�����h�Suimf�m>�|9�k��r�]���7@́��C
1�L��H��-���p�b|��P����Ǆy�A����ϊ,��"nބ�{��4�
4�[p A#�,2P4^h����"���	�_�ꔊ��3���6�p/[ ��il��P���H�G<ø���&�p�ë�z�E����xG����+��K�CG!7􅏩������H5�I0�C�m����D�d���@m���+K����a�/w�w�=����Ѝʫ����⸆�F;�����c������y��Du��'��KJI���̰Ʀ8�9���}�Ūi2a�p
�>��0$Zf�쾀��u�i�9H��0��2K���%Sj�{�B�~�v�>g>��q*����`T͕���㰠?�sv:�{.�ʪ��|���v��J|د݆�m�C^7���	!�)jEq�O_�@�w��^tv�8�9�D���A>������遃�̯��9�X��~T{i��[I�.�7u���\��f+C#7'l���I;@bԽyR��R��at\/���!.�	KC5�`T��� ���L�s���k��[4�1���y�8�D�QF2V���B��H~f������;}�Mb�{��-�Cp�.XYh�Pu	ۀq;���`�,(���^~����&���@<'m$�h���{@���.rI�C�>��p�òv��M$%���\,�l����s5��Op����� �q!��i�Y\��TS5��@7�����o����Ε&ܗ�P�т�I��eڧ���g ���=ʞ��B�,4��ΉQW�5H�-&�tk�7nł�M�f����&��+./������hL����L'߇��6�� ~��MRk�O�s��Lf�ߐ��v)Y�H��i���~dj?�1-�V_����Κ�{7��SToX2 J=����S��`�(�c//	K�<-��<�?2����U��Z��*�ڻy���5�c�$��-J�ӝ\�t`Dh6=�x�{I���?u�[��d֬���TCI�_u�3I������8�M������6յ����W��5���q��7����J0tD����%�Sw��7�[�`ߑ&�8�
�EO����O�1�����<̛=fį�#i�E�����>U/bD
5>+�e
��q���x�{.HD�K��cx�M^_�R�!!�,�,�M���@D$z� �)c�Q �b=-�Z �A��p&,L;�0LӀN4� Tq�!{����}�Ş���T�v�l9�� Z`���=b��Q+���j��I�k�hPj%8x;�?f\梹��� &5s��ᢳ���E�њr�p9��P���8sb����˹�q�Zv(��t��pP<n��G5'Fމ���  �i��(M�&'tU��~)rJ�������/������V}k4M�j�N��<5~�W�9�t�x����D�^�rg�8|�[Q�0�.D��w�̞�TK,~L��ߎ�Ia��_��ֵ�����6������B�����c����7����S��-߭ڔ�>�<�}}_ 󢻁,9���/܏N�V��`̎sԠS�Ҭ�G�����P�H��^��`�k>�f����P�+�ʼ�\Ob�Jo���G���HǇ�n���4KL�o����ǯ�MdH6�z?N�{NU��Y�X;&,��T�턞߷�<��$�q���@H�`G�j��v�!���ݴ��ͩ�"�e�n���WM�����S��1)����:�Ɋm���!�����q��箻=��:�Mx)�I�5n[`����ǐ�;5�}�e�j�qR�{��d	,`�^�4J��b���Q��*IA��p����2�ﾙ����4�	�kS�geB���w=�?πD�{��;V��P��������NbcE���t_�:�8~{�@i}9$�Ņd����e�����̸���r�2�g<���M>�����b���b�*����yFh�T�ޯe Ép�:f������/����8l�v5m��H������]�-ׅ	M�Z�$�c�%3���S��V !�|e��4�E�%�h�k����9��z���O
$kf���K�v�=5?�y'٤_��a���> �z��?ڋ#�;[�H�wq�B�ܡ e��X�a6�k�5��O�W�e��l��ߨ�I�Ǳ���J=�{iXU�J�+lF�%��Q��2 �̪�#g���u9��j�jl�N����\�7��[a�H���>#���n�Q`���{��R�o��.Y��{�^�5���\��_��\�ƢW��b{zD"/�d�^`ki sHC�'�B�p��]XK��U��o�������j/^5�������_�����F�w�~z7��|�
�O����ڿ�W��Ī�q����;�	��VFS��a/�u	�r���ϥ��:=~퐒�G�v)���$�y���8�怩kO������r05R�}B �Q�Nv���h"J���B?�&�/	�_ }]��k�v60w �/J�O��}�����*���>͉�P��&݈}i��N��N��q���IK_��6pB6/yot��*~ �w�[!�z�Z <��wS7TYi�KwJ��o�Z-0Q9H�9-���f�ZB�$OQ	�{�>I��x4���������@m��؟ʄ�r��P�-�q��j$�ߜ���ۚ�1Éni�!��a>0xb�víҵV���w(g��E~��KaC�'�k���;8���g1�1���w���]^� ��\�����%�y��{�9ϑ�� �;��~�"����
ũ��m�C*^��+�E��Ц�A������$C��&����IV¨;��-%Ec�<�"�:��gt���c9�0x����E�{ѸW@eR��6B>C��LM�a�+i�r�H,��f^^�;���*$*U�(�xopƃfͮ���il�ć-�[�.=�tsJ�;0�x��:����v�1�&"�+̑nW� Gl�hIVJ�����ŚxE.�7(�
ЇHY#�ݯ�USZ�������\	����LL°���c������� �Y[u��P§(\����b�||�jF���۱���"J,qk-��q��
e����lV˰>*Oh�J��#XO�!/>JA9����\H��u�?���Z�9�HW��Jh�^�c�.���/H_�?��F��!�H,�)��q�j��T�p�-K���8B���K�P)�ҋБ��[hc*T�E��m�x�j1���8H��Bw�-n��t��.v�\�xҮ���$A"�=�@m�u���Q��L�:�����_0@�������j{=�?��Ҍ�X�BcH�z6XN���HYM����J�¸a� u`��gm��,/��[|�M�y*�}n�NX̻f�ȧ&~0�E�����?�
|:f�(#SnR��x�>�zu�oN�
�9��[&᳍!����� �L��b�L@��Cə�.�lٸ� Ú%��oZ5.~��%����>���x�� ���Q�_��W�ۂ'c��v��\��>��Ws�HQ�<o�E#ݚ�, �!�V�+�����(
�6������F�E����)�/��\�R�nG�P�B�>��1���,2���Q(2��^�py9����O��1P�H͠��/�e�/��kjM���l�Q��Y�~��l�R�`5��H�`ŢPx��Ԝl#�M��Ж�x���1~_)9�5!�q�����nu�qJ�|'��a�
�ѿ�Z ��{zECs��a�g�O+@����M1ѐ�O^���F�۝�UB�����b�o��t���+�KLʳ�����F�?��~L��~'��jC�{�~�C����9}�1�J�J�����Sy	ꀑ[\�Чq��v��	���K�8�BH�Η�.z�07���$��{�� �O�t�EYWY�A�?gF�nr�`. =<��e���5Đ����X����ԋt��	�â���h�Y^�#��,�n��/67�]�]�('�vR�sg*,u��������q������l[m�d�N󦧰V����w�" �������!|1��!	��(�rfA�������G0ӧ�C��&I"�t�T3�*���
���?��2u\����n�}h�Јɺ�7J��)�S{���8����RkI��Q��zchUQ���A���Y�އ�o���v��Q¸=�u�Ky�	�Y��7`2�I!�|B���=S�s-'���ٰF�a2�댃j`v�V��L�΋>��{��e��e���Q)b��v�]�?�'�z`pA"�A��b��i����/,-E��̝1�_�Φݠl�d�Z8�G�K��e-)��C��hq�)ͬ1d�T��I��N=�2�)����8�l���U�Gĳ� ��3	��0�3���w0Yu�Ϧ�	���������j�<��"��|�,����̨��˂J�b��"BPH>'+O�e�����cE�W��=M�MG+�4�*�"��`^>w�G��h� �U��b�wW���+����1��� 4~,A>��hJ|�_�zt�1S?��ǅt�7�^�6���<���W jsiB�z�>k�U�KW��� L��5�Yo��G :HG(��eW$P1!8�(�����)W
�J���XHfeL��c�ҷ�[���[�ފ`��X��bm��r^H���N��r>�.�#r>��F�.)��'��]g��uD��V"4��Xj
������_/�]�����1��[�a!O�����;��7����.C���E�T�БB|N�x]5֧b�ɩ��o���Ж�w��.��Y�Trɼ��B�䕯�tb]#�%���(��q���[���b�
��>�5����?��_fXԅ5X�Ѵ}����=@e���jKx�v;����Ah�fRͭ����O� �q�U�W"��N�M���;v���d�iK���gBQ���}>~*e�;��p�.mC���V�y�o��]Hk�؎�m���hz�ݷ""�\J�}YLD�I#�H�������׷{{�@� j���y� ��\�0g)@M����	��n���^d�=m�� ��Z�_���[�Z�+�(*8B�6�ֽ�f
��*G���Gl���Yu2�����-��en&0�%«�7�05J�����T��_�z�\E�/?�`cP?�Tg����ipUC|D�hF�jS ��Ç�ۑcӣn9~�u�"�L���� ��IU*(���ʘ-���vr�㴊��:˃=_��A�`(��e7A~�s-�v	�����djy�Ռ�+-	���x7p}��O#<��
R�?m1�өHx���I�BL��ܷV1��5��=�C뽜GnB�o�`�>
��l�x(��}��[��B�kp^$]�c^��Fxu;R�X�EY�a�&�xY�1���S/�|�V,�5��*�r�X6E�FS'|p_
�$�u�E�E�V�w�Evd����{��J�҆F<Dn9�4�!I���_ۅu-���$������0%�H wJ�A XY��B�L� �`�k��v�P���R�]�îY���2�N��J��ϋ��^|1�E����R��s�x��s>�#ZB��A�էv���o�bC����L�wA�m�h�{���߁=�C�.P
 ���Nb�U�u�����`T'�����!����ň���I|�ǥx$�g�pg��}퀷�Ţ�,cr���9ݑ^����x���]��S��พ��<�a0�v?]@ʰ��F��� )�z������8�L��G���	�Fֽ�� � �u���4��.�m1���VG����[NOHW��V�[Խ�V�f���dE2e��>7ហp�<���W���A�p��g��c�\5�;��8ٻ���d���^�F,�G�D��� :� �]��V�=���XX)>��K�0K���" �0��B�����/cFzY�4��6�����W�X�ȧ ��P��`n�*�,H��i �%��ZD�D.�a�6�Is�1��g��8̛�<���(E�C`X]��
M�jy(f���S�?.��i�!@����O>��F�g���"��l7if�A�ߤ!�a�� 7
�(��e���ڑ'�]UY�:r|	�\쉎� �`�Hm������.Y����N��u����
�e�q�X�?��ȅ��c�X�{�.�LHn���Dg%��t���d�z?.Iy�k��`�Fv"�����p3��W{���[t0�,�}�n�����뺍9Fߌ��K�Wn7^�J���P)����;��Eݎo|�ռc�r��b�Al:!%�ٮ<��M'H����_�T ���*���c��X��59��r��	�J�`�q!�hg\d�K|�{���+P@�T�uٜj������P���6�X �s������@��˗����jq��?�!s!vҷ,�>F�e�p��`Itg�I�>���s��)����ۀ�.�:�p�ԡ+��=�W��)�+�&����+�r��О�  m}��HNH�+R	�u������j1��-�^]�i�av����Q�#�����˱�i��=������D2l��ԧ��������授W�N�Z��h�7�M�0��v�B��iŲ���]"Y�q ���hf��
��Z�ɜ��5�*hu�4�&P
��Mf��#v"��!#1oe"�JD~j���"��-�9U���|���WbCڮ

v�n
� ��ێ�H���Gþ���9�W��=8`G���q��8*$
c��0}��Q�?x� ܼ�\U���b��=�j�PO������{%P��Y�]�ܲ�g"��K�Ba�'x[@���ߖ�A,�	^���6N60�
.�		J�ʺC��a�D�2�af�g�]��d�J�Z&��^ȭbՑn"/*T���Ib���������EȐ)�Wγ12[15���J�j#s@�E���i��c��ru6�b���V3�`��6knܔ<�Ԫ�m��:������֜��<vL�՘��=��7 T7K���Bl���aU� ���I~)[$�K��2\8Kp:6Qk��w�������bvξ �i���(�9��ˌ<��3]�������.�����"�}�B���a|�v��>���q3�
�X�_yl�ͤ��\�&�$0��zt��ajU�pӝ�9#��|��H��Ä�J��%uD�JGk���R�3=U��]| x_AR�)l��9=�=��M�o ��H%�T�b�'�K���P�4|�L9V{T�Զ��t	����hl:SR�&�Cx�J5�ȥ��̦ɰ7`��q����e�-�O8\G��KJ�Z��yW��ؤ��1�&A���hWB�W6"��78g8�g|i���π���{*�_ (��d7���
��;��S�!rԠ�YM�t��W�g�{�`��0v3S樂�\7JS�B<!���^��������n`�z݈������X�p�,��#�S{�2�ءz�����,��K���Qh)���BS����$�aW�3�💣C"����앑e^L����v@`���t�HW�����PN��/�G��9Ay������Ra��6&����q�ӳX����*7�}��9��U����Ţ��g�@�_7x/���ey�V�P9�䫔��Sy�����iʊ��d��c�)\T��|���g�Y�8�1ӟ��R��M��0�^��?�6qiv:w28�ƫapQ����U�X{z�۝ۀ����޳�)誋 ,:�+�m�4���a�HT�dFLC�L�.���R���n��V���7���Z���`��ho�KsLB)oe�:����o�w����y!�a!�8�+�Y@����b�*R�A1C��e���eu	ڰY�}Y�r)D+�I6�ӣP&�_�0���.:s�FS/���M���p�x ���S�W&Ь%	0`������T]����9҆��@aD��?���=+�ݕ���"P���%�\�Z��n0,��_�8x�� ��~x<���rh6�6�6����˗�&��13�(��}G��!ܢr2�RC��8|q���a&,yԕ��(�|ד�4
�&�"�q�gy��4��E�h�p}a���̨����/�4��jړ��$��f`��� �P�k���P�d�
�wT�W��T�=>���ё�h����>��#�Ҋ�2��rh�/�޲5��x/qFsM��	b͜F�C`�Z��˛�ޑ����H�r�`cX�;�c��5u��3%���J���BP��)w�u�g���h�1j�=��I%�������TE)J�|���F8�ЍCARC�qh�k�}���G��k�wY22����|{����_�m�<h"O��N���(K�&��L���ޜ�!͙��C�/!�]R6X9�0̺���J
O��Ʃ��j�ZwF|��������,����6 ����\���K)�	:�9�`�}�����qKEO%l�3�}���Q��CG�_�c��vG<��n�}�j��Z�`v��"do垪;>8m�ܨ��0�$����9���2�qE��єr��2v�ȓL�8�*�2�*�I�;"�Z}���b�]3�t�/��#K\Iy�X	���4聏��w�Ӗ�zD:�I��bl}�e�іSƣ�.7��d*�>Y,�����d0���Z@�T��C����;�#8��s�����/�v�����qj��s��R�١&�je��<��%�M/���)��ȭ�@1nZ�YWk#����cr˾�C��h���;4M�D
�� h��ȁVg!*�x�*~��N��|Ʋ�%w!':��<o ���9��(i��3?����!��X��_��AD�}[ʰ���-$ ���8���N�&MR���wb*
�d+lwn-y��yм1�����`xءV�M������dT�Ȅ����w����wH�m�8���T�`�Y��+�ݟ �͑4@�;?����5�K86�hE��Y~Nqc-��q[K_s͵A�DMY��Ajp��W�
OZ�} ��P��y����L��ɕ�)��l�(�P;�`ur���zO��zsH���V�wE0Ό����ڏ�e�SH�0ς�&�9:=�w���21eAhVS�L�e6�GC����������z�����N4���ɓ[���̈́]��i�&�yBs��/�2?s��I���L�2�/T�y{c�����E՗�g[�B���W���1i@]Fyݠ{y������,na80�Ӊ��e���װ�|K���-�`�ض�΍ '����k�G��j��͝��Pk�s��Ģb�����:�z�$��H'���@%��'qn���ê�̍�߯v	W�v�̋��þ��{)$:�il��&hG�	�$�5m���Bh�f�<P5HI% ����jb�K�,�R�B���o�I���� �Y�rd<�7�'���^��Z{r���3�!�z\*��T�kLB �8#\���v-u�3]7��cFL¦���c+E�P�{(_]������+��K	z�f�7�axЮo0:	�b�wU��BC2�n1�&j�M;skw�����8㈂29|��'��u���v��D@��9���,�G����cP���{���\�^�EIۧS�N�v�m�[%��C�s֋9䴱Yt�?'��+�AʮQ������3��;Sr�P#˶��$�ݷ�����*>�#h�����=J�<6:�@Љ��Hͫd*�ɒ��^6zA��pUᏅS��q�`�x}e   ����(����P�I�[ur��cg'�#b�o�y<�3���*���NZ0���+x��q6ɾ�zUoy��[-��׿̮�q�EHҾcrH��!��05�+������B�Hfr	L)d��lܖ��{x[д��`�ѿ^�.�[�dT��#�?����$̋�~�;�h�ʗo2A��M��Q��9L���4���~B�8�%EL��h��6W�ƀ���2�J5�sB�I'��G���(�@���iy�uvw^�)N��9^���16xm2��d�#]�����ؿ&��3Ohr'1-��#և��T�;Au'��Ci�o��29�2�;Z���[�t;xe����S�a�X^Qy���l�R��k��	Y..i���|_T�f��廨�E��-$��)"f`/�dg=�AH�%��n�ݸ�A��$�Jc߫��Q�1��@�*�� �ǔ"�T� �c!h�O�u�z���.�t�%^=�����Ə���Tzn��$/1D�I߫u;��C��k��[j�_�����?ï�����!Z��Ӧbͳ绚���=]��&������
��GJ����4����9ݥ1�?6P��8*��J��������#_� ����g���g6N%x?�	g]��
J�U��$�|w$Ƀ�2�1�r���h0�͕�l��n����aO�'P��cHi�iٮ��vfX�z�����Z���s&�H�lH��&��]U,����d�]����\e�{+BK�'�w�f����T�\?��6�o��|��[ af����b��z( ����kJ�}�Ā�A�ʜj
Yi�A�������f�#'���[��xS_�ߐ��M�o��j�����u;��ܪ(h�]x,4#|
��m�wx)I��m0�6�.� �̬EK?ڱJn�J4��}�766!�d��Fd9N��{iG��Z���-8��n�ʿ F��{�,���4ke�z���'4n�� ��7�U Y�W���˚�vqTo�>X�` Y��y;ѥK'�Ρ��
�)��T�v&T�bG���참+Ar~��~d.keI|����>@鬒w/p�L���v�$��	����n�S����rI,�{�jhWk�ͮ�o��Q�%#B�{ء�~��)�-���*P E)��;�|����W4E��j,�u��b *g]�c��k]:\�i�O����Zm
��eY��d�ȝ�nM^Wԥ�	T$R䪠���e��8o�D;z��T��ŉ��I/�L�'2O���W�@����2�,{mS�+n������O� vB���`��V��`�Od�qtIM$u� ����:n$�r2{2<� ?ퟟ�`�f�ty$�H3]`&eWbд�`����7�˸���I�B]7N�]���E��l�FD��g�j��@�g������v �HV���?~�F��u�"�w�%���2�~�ra�Ra��t�vN��df`j�@W�zd���uG�U�6��Z�-�!B��MR7�a���P�`���˙�W:�Č���8��O�u~�m`j���A��❧��¶�^Z�lǈ��2��z��z�8q�f1�c���v�K��y�"RE吻~�,'�xs�<����W�y^�8٫�*X�Z0vָ<�t&�kM"SΦ	�$�D��Z�!Y���%�U���1���"�܈տ I6 �q�uύ�7����@,C/�{�^H��nW�����N|�E�ϱ��o�l���W���~y�b�me�&-W�J��OY���jPxtY*��sS6Yα�9��4�T��x	v�H������I��#��.$l�����P-d����W;z�'���O���E@7L���ދ�U����Um�G�k������`��,OȂ2#�A׍K��*/X@���]ԂQLd�-��[D� 2�7h\IN\PV.۲ȇ"��(��f�ޡE������I��窋'�p��3�q{���W`�.M��:O%$ۏ��8���M+�ʮF��u/C�'aH,�[�o>�e��
l�`�!��Oiu0��V��2����#���U�6i��!�ʙfmT��	;u�3@�P]�v��v��rX5��{w���tn}����ˑ�kd��a���WU�+�C>3]�E3���F���#Zf�3��@_1s32	�����`c�I�����`{�t`w�{�݅�OO� AT.��~�c	��P1c���{o�5�o�6�ˏ2L�@�5h�LP��.]��?</0���%/JhT>d�`:�a97k��8�67�B`?�mŨ�m�;J}�[n��pY@���9���9!�������v	h�)�ѣ�k�b3͒Ο��'�Kgv��eX��b��!u2h�7^�U��2�!{��
UQ�7U�6[�{C�N�֙Y � ��l�� �}I_�M��>�ͱ�gr��<}u�?�`��j<:�Iȑ�V������1vkw��E�ډ��| ]��O���Ѱ����ݝctb���{��|	�������U�dT;f��r1�M`3���Q�Gę�.�S5�Y�� �#�o�	�g���̃��#*&�1�N˚��^�z�b�}1�p�&h�~v+|r�TW`�Xđ��C`���g�HI�>͔>��e�X��+�~<s�n-��U\�
p#�|d�j�wZ�I4�����8Q�sa:&i]Հ[�Y1�������RXeL��9���K����T��,�Tx��{� ���X rܞ	�MC~��|�z�唋\/�䖴��
��Fw�~p��J7�lAl��fBq��h���+0��*��G����ǚ=�N�G[N�de��Vr+�aOHf�zѵ�3�a)�ʁY�����^�À}2�s�2�W�� %�c�v8݃id#Γ���'0ZI����ET�_�a��P<���H̒�}�v��a :6<T�� U\�ꀠ�~zXJ$���M���[��q6^�gh ձ�N���b�s�n��u�P,r4�0�F_(	�����a�!��f-��Ԧ��j*k`�c��0O�\���M!��r�ȶ/��Lq�M�H&@�+ˍF)Be�ĩʼHu�㕀�@��	gf@�utjL��/��8]#����'N��3S�+��n?�썵P�n�s�G�N}��D�@b�/&�3���7�V>r����~q��+�炐�E�0���g�F'��	m�� siBS�WΚ���=70��ͼ��+A��v^�f���8��J_�N�u�v�����@%���~�u���%�\-{��n�}�(G�&���+ե�?���Էa|9�DCLץ3h�5$�l1|����y��=|��D�w)}f��߾�f}.���������u���Z��m�q��&2t����XY���%DK�"�=9��5Eihsg5��sL�����R٭Z
c]��h%�*.���U�;%���]���U�C	��	��ޢmL)������;��t`�B�(V����R�lUIEN�B��JƶyO_�>�B�в!�I����S̮�ce�N�G����cIbi�H�J�v^�{����0�󦪙� �|��=3��1sCB�x����������{�J��cÏbߒ����CI�莬1�J_��tc��Q�\�n�ӎ��n*O��7[�
���f�}�����þ61�sқ��B&��c���K��ߚ^.3�\A�{�� ��S
��-x~�64�	в�-ܵ�������𱩣��Ss� �d��&|��h�7r��/�	�������u.k������U4/?���k�h��k4Ӆ��ۺB	�=���F��7Ʌ�DW��1P�=S�Vg`��!I���o��k�w�V�mh�ٯz�0v������&h�=j�O��Gۊ�L����w�'�t¼*E	����S�E�X�/�����Pg�A�2��s��a.ja";�fe>/��u�����K��}��ā=;�ɗ�0~�>�5ډu��$�{ħ8d(�Z*K��!hA}m���ޫ�g�)��n�쿐�m�(&���D�������3�Ə�ӴHf�vU'����}�� �Z���:
X��R��D�Ŧp(��@���J��m�� ���'u��l%����ח q+}���:��Q)�9�� �_���T����Z@�L�F� �tK���"D� ���V���l<s4�bS���	 U���<n���5Or[C����n����g�G(}B��"_�y��Ƕ����4�vI������T$�$����t���a5�	�W9hIv�(z���G~ȕ���uѿ�!���n�՘����>���R3����O~/�"�C:w�vCud���<5M�,�Xe.��s.�?�Z��L���C<�f�m�g+ow�c4{�[ڛm!�4����G�n��a�6�I�W(f�N�p���a�pIb�ަh�MX��Һ.'/�t0��)���YOH�|���#Xz�[]�v�y������,��	�0ț2|�5,�F��,��%��_�h��j7d�!E�bh�7�!��NS�,&�5�T>g-A$�m9B�y.g�^�ma�����	H�b���\{�JCע"i�u�e�b�|Yٞ��:���-�7ڢQ�2���!ĉ�]����y�
�g��o��=��Wu�G2�2�}}/7 �E�����B��F�/�e�S+w!.���8��qawo�a�	/�h��6��Ko���C5��oB�=Wr"����c{���a�T;������bL2��X_�y���6��S��}����(���
�a/=�k�:�x���8Q=�K<ٝǛ��g�:Ɵ�P�TTv��=�|�=�"��������<Cq�"iJ����@�۷�����!l�x�P9Eb��%��E��7m�\�'�^tt=�t�����H�nU.���^���T��]�S�)��3��1�m����Q�PYRl&l͏w5+WS�q	�*�F6鵼ôNV ˣ�Ԡ��u��!�����@��W�r�~��
������AtJ�s��j�������ܹ�KH����aX�c��(�3��rX{�e=\�s�%T�Nty�4��	�G�� �1�� �:�lc���@�u����oĜk@#.� �����0fm��k~ ���`�ɧ�q�|7ǻZ�� }@ۄ�)���~x�W�	�;0�Fog�ߢ�L&|hr�
Ю�3�J��~^(��P}_Dv��#��!wo92�. ��B��ٻ��]Wk��ъ����˷�@��J��'�)�P���3Qd�O'�=�s��B	�񅭶�h�`�iG��*�G+���1�=�9W�	ˊ�� �5�M����O*-~�NB�%d!c/O��WQ��8B�vƄZs"�/LQ�f��X���6�.z<�χʂ8�N�(7��aaӵ�ͪ�T�K�3���UD���P��,DÝ��U�]�ip�O�j�ĺ���{Cl7����t��Ri�U8������<(l�磧�)
�m��-34'C����{�Ma�8�|�'�^�3o�rr�C�eY+7�80�	W>�g��r2��&��Z��Ev��r>��׎��EK�?D���P��'��$�����FT�!v�Y.u�Ě�o-���=~�O1^����_��IY+����m�O��t��wP|�ۇwW��D�@��Px!&9�m�ڤ��ki������:hC��q8&LV�%N��o�1��A
�K�pD��z�R��'�n��x����Tq�����_����VtT���l5E�ئ[{i�	�
�l�(��h�sC���d�������d�σ&�2���6��A�'@����*��6�;�.}���Z�� `��`��{[�Ctgr���
���9
;i&^�k��j_��6��lj-�k�O�-3x�C���3r�t�&+�0�Jq�;�fa*ζ�j`EJ�$3���*�f�^vݎgt��鈆���B���m;�Қt���ҿ�>��]c+/Jqq�����F2M �!o�^T3E�o��RX��2ΰLD�e��m߸p��ۂ�"�����J�ɋ=󒢟�k��q�ࢤv�+���D&�xf�Ӊ�d`)
'�a�����[��8 5X|��p��b.�M�8��_����ӳ.���h`���+U�m#������M9�T�ػX�  ��F8��}~���I���|�m٫��y.�6��74�8igݎ�MF���en[�@��q��Ҝ-8��\���ڲaRNY�̖���z}�zZͺ�"X��D����ub�V��RX�d�/�G:6q5��3ۭ�o���z��S>�,ks�<��Y��8�Q���[�C8��S���n����\���v�5�&�g8�ˌh�<��� ���.�9D�Q�2k��_v���<�
<cы��B�b2ƍ��ݑ��a���r�Κ�:��I�JQHY_��u��
Iٻx�:���W`�/e���c%�� ��N	LS8x�i��^�^�B�����t�$�z%3 u��ʻlR&�p7r%���)� )�ԟ�%���?K.��\�ݍ�骒�˨��ɲ��{����c�o}�۱Ǖ��R�?!lW"�ZF?�-rv��k�
�v�eO��^�zzZ]W��{��Sq���P	6�V�� �Y�!Y�YmQǣ=���`kr�]H}[Y�α�[FI�j��H7�qz|	��8`�?= �,f�&�^=�����#9b1�>*Z���N�$Mʞ4�D.�h�<F���4]ݴ�\ޝm�(Di�(ԁ)(+8M���.���p��`���9��-P9�,�I�tc�������	b�	��Y1�Q����r���d�k8<�]�-7C����X��I[2��(���NP �؀�w�d@�Eu.\�m�N/��N�#{b ���~���۹h��N@h��e2-[y�$�	˞����p�If�3�;Wp�M�(�>3�ŔW���bk����v�F�\��Cؔ�=-�x8�
�?i;v��s:��_9*5d��ϥ	���M�+�d	$��ڇ(Y�.�>�d*����Qq�"�fs�?�=�x\��G�"�b��bz�N�L<���ϒ� T[4���i���v��<V������b��9(1(s��R^p0�l�ط�w�|��r2Ҋ�ζ���gM���i�x��$�-�P���F��J׀DY�^��;�[�,�GLeO~�cL�D�
[�A�1�ѽ�z���
�9m��y/@!�L�8M$<CߓqLG�G(���ݳ���*��3�kG\�x6��IƵ�|��yyz3�gӘ�Òd5����W߆(���*�T�R�6�h��X�h՟k���WC{	�u0;W��F�lp���tہ���HV��ףPT�Owk<0�����	�r@���) ��C�8�4=`���g��,1�+=��c�]�窵��b^��!܍�bˢӨN�����F�����;�߼��!9���]�s�:%�t�����FZ.3����e��=�u�C��"g��ځ.]�|a>;d���&bc��;�x>����X6w�83���k�J�LQ��!�vE!��Iz�Ɵh�^E=�GV�	�>��@s�D`֮��� 9�#)v9b�)V-SěH�GL�I|�2�)/�<~2v�,GTm0�n� ��
���De�� [�����b�x}N̓ⅈ�_"v��TՀũ}��5�7���@������;�X�j�Ն��vb4���d�F�1cYf��L`J�N�<�E̽�{c�T�f{��8��óuƹf7�7%�&��a;C�7��-���f�r�M�i�/5/5�d����9�h��f+�^ �;8�q&�s�rC�Sz�-���]�$7x-� LT%{�#��h�Æ���7��Sh��씩�`1C�"���ɒ�=��JBi�E����v�+����m�z%_�ሧ(�?B��"i
an���%2_�̅�X�Hꊜu!R�m�hGI�Ua�����Y}QC��U�� 읅A��t-���g��2��5�K����1�^b�o"���3���F]����>�%|$��L�o~_���
���ۣ��PhA�����1<Xv<ŹS\I���~	yv�Ő4�� ;T�"��⿱�����?����Y���N.��#gV%�h�����6���RmZ�Ϙf���|�� 2rQ�J�x6z�����;-*������znAfq�������/JE�nd���cܕ�K>X`��(+��zƂ��8�ӳ���B��g,��8�(2r����F�����Q�gWxL
�-3n�2.��IK�?������X�7J\Nэ(V��o�(�;��2b�E���|��ȹ��-~DJ%�;㓦@)8�ME�a�9�4�ֱo/'�TKt�D�_�נH����(����v�d��Z���
�{*����{&������w/c�ec��8�'��m�@��עU�Qޒ���n��ϥۉ�y� /��l�Iy���Q���(+���_�0(��'�E����q0FX����:�J�F���Or g��D���dP���,BP�6���Z�)�jU�[f���������-�B|h�ʨ'���CX�U<O���l �$��;�vA���Gi^+�=d���o*6GC��E��E:8o<Q�b�Eh�T'�Y���6&����;iU-�G��}�t�vw�_�����)�(�P~��ٟ�ܴ��'v�Aa	�
���tWY�֓ �>��Qܜ�q�W��4�-XcDE��N�6.0�Ze�w;_p���=�y�<jڕ-g�N��k��������"��ԏ!��`+��ݱ�Fb�4��3$�%�䊣F:?�Ȕu���*�V(���'�\q�S����<3��-�� U��8LsB.����H]��S.����ŦAYmmf���w(��;j%�	Im0d?�q�P�{)�.��C6��_����}��f�ᇗt�[���% �EOfρ��R_ns���������j�)pL7Aq��+!RWUӺVS���V&j.�{��F�i��U��KU�h��.�r��wjyT
����.0-[b�DD�A�k���?п�5�^�i�r������"F#�Gr���D���V������g�i����v�i�MX1Ɋڢ2E��Ox�7L��o��� ��|��X�+�k�d�x��"c�@ J^j��湍����ɂۅ�>�x��OO����%�����s�jQjSN#O�z�A����qdc��j�*�{�y݀%~Xc�ҫ�|5�r?�\����U����O���<&�2�^K;�CQ��L�ZO���(��}TYx�cI�3;���Js�eiy�/�1j���᷾\{&�m����c_�@���%���|�ޮ	-�iĞݑ�`o�=�*|V���7�lABL4ڮ�3��/ҩ𯋙\�u�9B��8LG�����wF�k�R] �<�0SP˃9���P�8Bܑ�H�+ǘ%	n�C��F��Yr�I�$ym�IR8ض��z6��Ӯ��-�'ء_�mX<���*��,O�=赲X�ɢƽm] I:�-�jap}���k@���<-49xB�U������-��߼so����jo���D�ܟ��8y1c�(	��g��v�<J���:�E��˙��E�zC�`��;               `� �F ��  ��Ǉ�� ��U|W����卜$����1�P9�u�FFSh��
 W��Sh�� V��SP�  UWVS��|��$�   �D$t    �D$s ��$�   �B�D$x�   �J�����I�L$l�J��H�D$h��$�   �2�E     �D$`    �     �   �t$d�D$\   �D$X   �D$T   �D$P   �J�����6  9L$ts�D$xf�  ������$�   1��D$H�������$�   �T$L1�;\$L�|	  ���BC	ǃ�~狌$�   9L$t�d	  �t$t#t$l�D$`�T$x���t$D��|$H��� �,Bw;\$L�,	  �d$H���C	ǋD$Hf�U ������9���  �D$H�   )ȊL$d���   ��T$sf�E �D$t#D$h�l$x��   +L$d���i�   �|$`��l  �D$��   �D$t+D$\��$�   ��D$@�d$@�L$@�6�l$��   �|$H��� �DM �L$<�,w;\$L�`  �d$H���C	ǋD$Hf��   ������9�s#�D$H�   )������|$< �f��   t"�.)D$H)ǉȍrf��f)��|$< f��   t���   �W����y���   q�6�l$Ձ|$H��� w;\$L��  �d$H���C	ǋD$Hf�M ������9�s�D$H�   )������f�E �)D$H)ǉȍrf��f)�f�M 뇋T$t����$�   �D$s�
B�|$`�T$t�D$`    �  �|$`	
�l$`�
  �l$`�   �L$H)ǋt$`)���f��f)���� f�U �l$x�tu �t$8w;\$L��  �����C	ǋl$8����f���  ����9�sR�Ƹ   )�l$X���L$T��T$8�L$P�L$xf���  �D$\�l$T�D$X1��|$`����d  �@�D$`�t  ��)�)Ɖ�f���L$8f)���� f���  w;\$L�M  �����C	ǋl$8����f���  ����9���   �   ��)��D$4   ������L$8f���  �D$`�L$D��D$x����� �,Hw;\$L��  �����C	�f���  ��������9�s`)L$4�|$4�t$4�D$H�|$t �2f���  ��  1��|$`��$�   �T$t���D 	�D$`�D$t+D$\�D �D$s�*B�T$t�1  )�)ǉ�f��f)�f���  �  ��)�f���l$8f)�)ׁ���� f���  w;\$L�  �����C	ǋL$8����f���  ����9�s#�Ƹ   )ȋl$8���f���  �D$X�   ��)�)���f��f)D$8����� f���  w;\$L��  �����C	ǋt$8����f���  ����9�s �Ƹ   )�l$8���f���  �D$T�&��)�)Ɖ�f��f)D$8f���  �T$T�D$P�T$P�L$X�L$T�l$\�D$\�l$X1��|$`�L$x����h
  �D@�D$`����� w;\$L��  �����C	�f���������9�s/�D$H�   )��d$D���D$,    �f��D$D�L�L$�r)�)ǉ�f��f)���� f�w;\$L��  �����C	�f�Q��������9�s;�D$H�   )��d$D���D$,   ��T$Df�A��  �L$�D$0   �/)�)ǉЉt$Hf���D$,   f)��D$0   f�Q��  �L$�L$0�   �L$(�,�t$�|$H��� w;\$L��  �d$H���C	ǋD$Hf�������9�s�D$H�   )������f��)D$H)ǉ�f��f)�f��U�t$(N�t$(u��L$0�   ��)�T$,�|$`�T$��  �D$`����~�   �t$x���D$$   ��`  �D$�   �, �t$�|$H��� w;\$L�
  �d$H���C	ǋD$Hf�������9�s�D$H�   )����f����)D$H)ǉ�f��f)Ef��l$$M�l$$u��P����$�'  �Љ������H������L$ �l$x��҉4$�Du )�^  �D$�V�P��|$H��� w;\$L�V  �d$H���C	��l$H�;|$Hr+|$H��JuȋD$x���4$D  �D$    �D$�D$   �   �l$��D$Ł|$H��� w;\$L��   �d$H���C	ǋD$Hf�U ������9�s�D$H�   )����f�E �D$�)D$H)ǉ�f��f)D$f�U �T$@	$�L$ �d$I�L$ �p����4$F�t$\tY�L$�l$t��9l$\w_��$�   ��+D$\�$�   �4(�F�D$s�B�D$tIt��$�   9l$tr����$�   9D$t������|$H��� w;\$L�   t)��   � C+�$�   1���$�   �L$t���$�   ���|[^_]s�{�1���$ �����P9�u���1�^�� �
 �	�t<�_��0x�
 �P������
 ��G�t܉�WH�U����
 	�t���������
 ����
 �� ����   PTjSW�Ս�  � �`(XPTPSW��Xa�D$�j 9�u����"��� ,�J <�J � I                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                     *�]7          (  �   h  �
   � �    *�]7       8 �@  �    *�]7           X   xU
 R               *�]7       �  0 ��  X ��  � ��  � ��  � ��  � ��    ��  H ��  p ��  � ��  � ��  � ��   ��  8 ��  ` ��  � ��  � ��  � ��    ��  ( ��  P ��  x �   � �    *�]7Bome       H  �U
                 *�]7Bome       p  �U
                 *�]7Bome       �  V
                 *�]7Bome       �  ,V
                 *�]7Bome       �  LV
                 *�]7Bome         lV
                 *�]7Bome       8  �V
                 *�]7Bome       `  �V
                 *�]7Bome       �  �V
                 *�]7Bome       �  �V
                 *�]7Bome       �  W
                 *�]7Bome          ,W
                 *�]7Bome       (  LW
                 *�]7Bome       P  lW
                 *�]7Bome       x  �W
                 *�]7Bome       �  �W
                 *�]7Bome       �  �W
                 *�]7Bome       �  �W
                 *�]7Bome         X
                 *�]7Bome       @  ,X
                 *�]7Bome       h  LX
                 *�]7Bome       �  lX
                 *�]7Bome       �  �X
                 *�]7       P �� �h � �    *�]7              �X
 4              *�]7           (  �]
 a           D L G T E M P L A T E  P A C K A G E I N F O  T I H O M E               (�
 ��
             5�
 ��
             B�
 ��
             O�
 ��
             \�
 ��
             f�
 ��
             n�
 ��
             z�
 ��
             ��
 ��
             ��
  �
             ��
 �
             ��
 �
             ��
 �
             ��
  �
                     ��
 ��
 ��
 ��
 �
 �
     "�
     0�
     J�
     Z�
     b�
     p�
     ~�
     ��
     ��
     ��
     ��
     ��
     ��
     KERNEL32.DLL advapi32.dll AVICAP32.dll comctl32.dll gdi32.dll mpr.dll MSVFW32.DLL oleaut32.dll shell32.dll URLMON.DLL user32.dll version.dll wininet.dll winmm.dll  LoadLibraryA  GetProcAddress  VirtualProtect  VirtualAlloc  VirtualFree   ExitProcess   RegCloseKey   capCreateCaptureWindowA   ImageList_Add   SaveDC  WNetGetUserA  DrawDibDraw   VariantCopy   ShellExecuteA   URLDownloadToFileA  GetDC   VerQueryValueA  InternetOpenA   mixerOpen                                                                                                                                                                                                                                                                                             