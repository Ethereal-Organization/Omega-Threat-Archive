MZ�       ��  �       @                                   8  � �	�!�L�!This program cannot be run in DOS mode.
$       � �S�N�S�N�S�N�S�O���N����P�N����R�N����R�N���A�V�N������N���.�W�N����R�N�RichS�N�                        0�?'t�Qtt�Qtt�Qtt�PtC�Qt��ts�Qtr�Ztw�Qt��Wtu�QtRicht�Qt                PE  L �lI        �      �     ��     �   @                      �                                      �<    P pv                                                                                                                  �     �                 @  �.text    �   �  �                 @  �.data    P  �  P  
              `  �.rdata   @     8   Z             `  �.rsrc       P     �             @  @.reloc  �J   ` E   �             @  @GetProce                                                                                                                                                                                                                        2�8��Ҝ<�o��.}� ��2�~�t�%[��֛�m̎J��PV�s;�{�bzղ�������֛�x!��^H �0� ����B0ihX ��D�������qµ�����y��>�O	nxB0N�%#��e�K�:ɔ%j���@����D%���@{�;��ƶ��t���41�i���f�����a� �l�O��)[�%���İ@%����^�$��0��;��[������K���G:�yp�"�>+�,6��A����z��cP��A�U����$Lݙ78<�����iH�!������?�D%k����f�22���+��z
Z��o8���Jf�	�������qȊ�r��Sq�A�a3����j��������nb�;�!]���Z�s��p�ݲ�9�K:���ۤ)��y��(���l����������8������c���^�Hac�?������x\����}rt��C�J�VG����Пk�5��|�� q�;v�D���fߘ��*��<����\Ì�����ާp���5K��
���UN�~�5�/���b�tz��i���1�ȉs�tRbv�d��γm��u��c
!�����W�F�L� ��%��׶r�;���d�bYr(⡢!�7���#a4	�B �S�?	����c`'i��$�&aT�7��z���a��=7����%.�y/y�!�W{��`��bq��Cv��Z\��|�ȉ�V�~w4�?)kMzC���+���;�i�K����4sv�3SHP�I`��%}�L�C������5�r�;��8�)�������GM�ܜ�hrE�(��`~{�t���xI��e���4��ᕠo4��Y���0L�A���)��t�k�!tƶ5v��*������/�;�>t	�'E˩���}U��7 Q����:�̫�u:����(��KZ�7�K��Ȍ�d=�QCі C��8���7x�ڐi��m�T(B�1=��q:?t$sٯjK��ԍ��=R�-��@�����;Q|QkW/B�2vHH�qgM��M��X	,��؟��hP����(Wb���w4���,��hn]�s�U�1��2�� �����%~"ٔ���|�s��`�鸕�H�S��!�B���Spk�u�47��򱍤�Aeؽ���#-�E��u+��b�����"��\���ycDO�s�����F�l����d��n*b����\A�~�,8{��K���N��t`0��j�JXK��h�rjN	|�c��64��xԐ�f8���� m$ng������G�c�I���9��y��bʞ��{UU%b0Jq)<�`�=��+���5A�B��&v��謳d-%Y9V�˄�8(p���tM�U�i��t��P\�~�bi���<�Q��-��!�(��t��{b�41�˜�kLS3���&<�̾F�l�t���s܏�K���M=�OS��x�=3?�.�γ����
<ͮ��s�:޳X��jV���j_�Lh��}������[�c�+�N���@V��<`l���+�mWA-�e��`|�,	�FaB0���o�,�ơ�fsl,/��|��]n�D���Yf�n�����]g�{�<��H�8�j�D��D_	5z�������4�y�u��v$}c摾e32�t�	͵SV��h�'���\$����\$��@z ���s3���s3�C��<��[ue g�G�!(�WQ��F���(�6���E��.|Ɨ����t����iE�Bi)d�����w`���슑=(0���x��MZ�1ņ��V���ڒyw�%��ߥu��Zp�ĵ�+�I�V��|;CD�X	�;�<0"K���d9�5��ȹj&�Y�P�A�2������#���y��%,��[�0@ ���@�����KH�_X�������N��F�CgF�R8�� ޷Z��SbQ
a㳳��8ʀ����;Fe��lz	г��3*|�*?�G�B���e4�����f�NP�k>ԣ����fP�#��0�����;�^g���=�m"BzR&DR(���X��Ds��V��At늁���Ua���n1ZF�h+8:$��ڑ�3Ey��i�/���S��h��r�Q8�i�;9��J��x�J����q ��`��ϸ�Д�iÆ�G	P�GN����~�1���+"��#�����*%��:�=xY �Z�� �@�sj��V��������	`����gzz����\�[��t�����z�p�m��/��?�����屽�M�n�L��%���(���&Yf����-�V�f�)y�`�gp����
6���{Q Pb�q0u8�t���5�˪��q�m�L�A�XE���ݽa�D�~�A���#��B���c�x����������+(5MF+�ˌ�a(p�h�2)WZ�o����"����ތ����gD��zJ�|mO���,e�ă���3���K����XG�%�Ó*xV��a%!�4>����r��`����(��ѹ<�!c��Ծ��!)�1�d���M	+���&�8wϚ ��v�/���Y�������'�(Ӛ�C0ü]�b:�̄�h�7D{��/����v�~��1��M��W��;�7ne�=qm\�?kn>k�|���|K�od(ҩ|
�p���1�n܉�d;�P�f@雒�Yv?7sъ�뭶���h��$�?[�&�ش�y8�{n�q�
 �PU�>?��4�%q1�+M���a"2��k�fkT:J:7����(H��͛wЇ��H�|:?�?�d�qD��h����'�3��?�<���������	V*�w�æ���|�ǱB,w=��Dvh	;&<OZ�2C�b>�"AfР���K}���=��8��<+,��]�I�(����-��-�F�0��,�"�"���&2���p��vo^��6����s�W�ʣҮ�Qa�b�MLa�r:�㪝�^!-˷L��r�Ӣc���	)�L/cɑ��	G*�2܂6���9T�7�L���MH';�7�-k��j��R�� ����Lb�s	�n�Boj�R�iLKZn���#)Iop
-k��7Q��*�W&
����:8�b���P&�3K�q�f����_8VۺKh�5�Eqf�LnA��p�J����A6aaAa���R����w�b��,�9���ɾ���S���w��)ځ��W���Q�����Z
�����xq��2sS2�m�F>;0�_����!
��|�oz�DЅ���˫;\}�`q���G�HÑ5����P�"K#�l�@��܆ms\�L�0�)D�"|�I�������#��m�^�n���6Ze T�����B�D�d�3��^���ή3_�yW
��խƶ|��A,��O䱴���|+��
hn�K=Sa�wg�~I���1�E�s����o��b#�̞x[��(4��{fb�;v:�i�X�b�S�U�q��*R�,�9iڻ��H}��%�dп�k��+�h{�jZeD�Y��N+��;BW0MG�ł�r}��v9u�C�nSR��l�=좍�"<�پ��xؔ��>ߝ��o4GHP5����@�{�*-�:�%ڼ�ǴZ�q �Vk{��z��f��M	R�В2~�����D�gC�=TMG��63<���s$.�#1�eT������z#��=���s`.d$�}�e��c���\�����+�ҢO�b��^ֹ������x��K�
�	\��0�׷ e�
��楤���MJ3�E���sW3��G��N^0����8I�fB����	�
����[���+�*��%�pH[�/s��D�*�H��,
����86,���HNlE��;GA�/�VI	ȸ������+AY3j�;�c��C�"��V_+��;
]���Hޑ�c�g#7�U���J����W�[������V�+5�(|�D�r8��U
ܽ���Õ`�z��zW���J<5�jN~�� ~+ 뵞��E�er�O�=��Q9�BQ\��c� 3��`�#	����@@�k���<B��r�N�����d�Ώ�J�����d�7*| cd�\CQsI̾�Abs�tws*�{"<�ʜ��W؜֧$�ڴS���`wʁj�K9��Z�o�����YӸ�`�b����c��Z��=o�p���o�'9�K�h��T�S���C%���@�{���Wھ�R��s�}DX�4��
-Q�m{<VZ�)�VӫIi ]�a=�g;Я��F���:H�,vl�� ��E������
_矲c��p����Z������t����ANo�q�N1��]�vo�B�����(!WY���2��؁�ܔ�lW4��y��E.�q��V�%[��/�Y�{��ꚢJF�_� w���� v�Z�daL�k��jG���O�À�~7X�_qId|d��d`l���rl��vV�FM��$t�h��U�"�Z�Jf �#L"Xw�4�N=�p�>Q?�%R����ӟG�cj�k���{Y�K��k��Al�>Z<^R��H~#j���d���:W����O���N�R?��Gi���aP��\oj<�9wׁ�Mh$��c�QD�C`����[�0��ʋ�O���D)=��ۛ���>u%�!P\?�r����'v'�A7�(Wr��S����/?��rǖ$P���� D�͓�&� ��9#x�X���9 �F$͓��(2a4���Nݻ�|������s[�nl��� �cp��r'�uq�PC���_@%�.c�H�ǧq�Bɲ���$�����0P�*�v<]��Z�@���ӌ%UQ%�s�t)�l���d��.�����kiɶ�@ѷ���uM���1a��m�|�Aև�"��,��T���|(􍅲9��j!K\�6����{�� =6�0!��������΅�!�p��"O�Y�����:�k����^��a��7��w�р>%����S�&��K�m1s����.����c��JET˛���l��ݽ�펏��5�[E��Q��$d�tBT�,�#���U��0�%_�0��9mW�P>�;�D�����K���{��*�����������WO�Q��un�!�x.�+B��O�Mx��{=����Y�}�,p��_�2%�aW�JD�OTXTנT����BT��o*����]{��)�[��h�~,<��_�o2=�|����b����I������1�i�`LQ�8�3�{h�&�D
% ���!}X�JE��j��bz�����X8��V�o'�h-;�ň7]��p5˧����p"#��"|P�qA���#��wxv�4�UVq��:��ˮ��Th���Ġĩ�i�H�g(�#���xɍ��� x?���rV�uS����0+���vA�R���!Sd����0� ���$�j\�/�ZB�%��=��;g��07~�Vb�6�|A��9J==��Ҳ:��X����P9�N8�}^�>�AA�t�hG{�m��/	�`����E��P;��B��.�~C3�?����̴��i�	7�5�X�?��]a@(7h�;-$��huH����.l~�n����,�H�O��C��քe��ҫP�T���ܛdܕ��7�y/�r: ��%Ъ�Q�j7�	n6����*Nϝ�s�	��(ѝ�S.�|H�E90`f3c|°m�Iu��\�>Q��w�K��[E����s����rA`b�*�^6�3��E��=��+6;�t���N�H0&@rk��mI˭�Y:��gy�8RS���^~.����X�cn�	��3UFi�>�ʊf�,�o�4���2���������5���:'�j�fQ�'��v0�x�)�N�<��MS����(Ќ�����b��A;m���� V��	�rl �]S��cRp�����⩝4��g<��֙��K&�l@�~L�6��L0Z
�<�"�2�q>���6�1���)(�`�Ppih�v��r3�rg������w�]��=�����������!����ypqܝ�S|��>���O��OL/���B�Ez8`��MV=��<b1��%����	���ԙc���Ǟ�{U��b�+~�1뗤��<"S��M�uz�d�"t�)�x;|ͮ�t��kh��O��"�S�P�=l���5�/j��  �m$M��hN�l���4��6��#��>�3d-����Z�Kn���w2�}�8�J�ĥ��@�O�^bZ��.��BM� �W��j*�UZ�0�h��ٽ�<0M<''E��m��b��GJ��H	V_�nO���C���/2�K
�����9��?��&�Q���C�_(�#C��HqX4�$�ų$?Y,)��:d+8�z-�(Q3� ����6��Y	�v1-)����&����Y�������ޫ������K��H��zo���Hh>IQ��yp�Rd)MM�f�Bk�:��z4r%^~
�������FV�µ!&���Յ{�P>�;�!��[ .\�!0���@��"!l�%Ɉ���k4��4f���Bq��´��z�J6yH[ʠIQ|��k,���O'���Fe�K�*�M��Uk�=mj�}Iu���RЁ���YQrNN�4����8?���*�8�Q�è�̠�Ĝ�]�т'(M�y�+#�*_�I�@�J 3��3�kä�QK�g	�36���l��ȯ�7sE���|�D������������6H?�@�S�y��q6�@� �UXڧ��l G8�z0MK��������������-+�f���vҏ���c8yN�q�(�3�|F ���@s��m{*F�aUl��\���� �}�L �1��ړ�Qo�c´�����]B�-h�T$6�����$�Yřh���N��3ȕ�Le @cč�O2�*1/��qЇ{���}�47D�1|3���1L�-Dҫ�xe�#�����@���>9�iY1��ų��4��dl�����b�	���+��k=�K�q���^*BY��2s"z0�7�Π�<?tٙå�]���-A!@O��P��m��52���\�Ջ�w��cʬ��.��azSW�ep=\���㽞��ʷ��V��] �	�NPl�	�w�(y���%#
Mܝb�ݓy�bAB�lFj[ ��������3!m�6�c����P�Q��I�1�T>f����U9HB���{�ׁ�c��	�g���OV��n+���)k�#��Td�/���D���P!S,�LF�p��!xߋA��)�K���$����7ʌF�j#��ga��Xa�ŖU�xQ=���Y�#��ĵ.��<�C��8�֪�O�5�$�m�������l\�@�Y^��0��0Py�7�w�k�\@����g�j����$(�NV�&������� J��B{�б�,Ε�U��|,�O�ɑ^�]9?O��S��D�l�)P���AU2����}-������x����M��F��U��D���0r�ﰣ:ඈzT�������?{���^��*c4}��*~^d�/�M�ǰ8dk�W��u��<v̝@��#�����7B��u 	���K�ΐ�4q�=H�k7�C�,�"�E�9����m�u�>}��uǤ��k�{�g�ڲ�j��o��OaB��v��)�^Ľ�O�K�u�}�M� �" ��&:2��hdzR����cM���mKwݯ�����>o��o#��f\�=�[���ᷪ1pz ��.�X�Su�|5�N@�Lp�r�8ND0����
F^�	��7��kW�#��~?�Jc�pm&�sv��J� �?�3��#x v��=F���J�u�e��E޺�D��}����UX��úHyJ��a�� D�3�	�6���4?��1�l�e���&/�|{5��/�C:�i"tq�[�8��ֱ&5&I�ǥ�	n�坌E��o8��y%~�Y9j�t�m|�ϲ��8��`�@l�a>�VV5[-����+�o1����7��b{3a���%EK
���F��P:*"�*H�u� |����@���#�لf����!��5�4A�n[�3������D�����{��irz�'��ӂT�T(dD����(gBn-���בI��]�&z܎4#�R��+m$+ Pp�P0�+z�/��[���F�b�t�]z�U��j����M�iD��JCN���b��/�b0��5u�7 ҆a�Ft}*�5J�7�Ǔې��=Y�����$w�9�I������Iԍ�gڣ̭c;��o�Uf�3�F���1&" ���|�x���Ĳ�n=����!��Zi����!�>�QhV��9h����6��Q��B��<�rjzd�bw�?_@f5�7\X�s��-j2��-_�����$|�>k%������uP�g�����S	��^c@�������q��g^��ϲu���ڊG.�S����P�U��r��[��4�)b�e�����%H�lLJ�5���0���}�~-�H���t�J{���i\��z�>��$��
�.;pre��ԑ.+-��qI۬��4�۽�OU̢��[�m]�D��2�UAE���9��)b�t�����D�R���}���
(A�3�'��]UX8�Й`�c ���{�eT���ؽ�e���S;,��m���=���,X9���_h����[9�]��ξR��K��@Lp=�r)U��&��;��Q��D��go(ْ���Fnw_/%�Z�=2�¡=�:&�:�k��+p%��/#ѪoI)���"��灞�_��B� ���#��c�gf��W�, �0�H�͇5h�����d�6�K�:��oB^q�5FN����HbV�5<D
���=inh>>�;��u~�w��L29([��X�����d2K�C�M�GB�]�]d��bW��%�Fy�LV�}���Y���qr��i�r1�燾XK�Nb�%}�ݵȬ�:!����j˕�	�W"l�s��Q'=`z�\�5a ��L`�w*\-yy��D��4��ci�)s�\�Y�ov��+��u�3�E�����I`u]��pFm����ˇ�B&��d��Frc��$�O�P�Ao.&���'�r���r��Ym���G~􄕲��tsXt���-��3|saQ?v�&�&�?Q�#��+�~��?���8!�A���75�VoYL�Q�k 8�U>N+<�G��{�~z
�~���{gN�dL��|x�!V�CƠ�9�������^��ֳ�Z+n���^x�Ow�+=Z���̩#��0�@�d�4akD�+B{�q�̫�%�
�}p����lz쾍�,t`pT�l��D�yS�l�,l>�i�Ny���{����B�	-@T��3��|K�W7��ת+=�>�̦ۗ��
�:=�|K�R� ��K��}39�̫��1+o��\��~��=k>���2�o9�nVY�����A&�G5x�����~�|K�4z�9p�Nة�?��𩡪|K��L}�.z��|3ͩ|K��*(k`��A��4KJG��(D��;n��E��3̩|K?�ԛ��O��|�A�ϞC&�S;n��|��ܥ�8�ͥ��n=A�#]�	d���|��i�g)xU��7���[˽�K##��-	l�"�n���.���x��ֆVt#�O�JU����z)���ɿ��14Oϣ�h��|�����fv�ķ6�Efi2aC,�E �(���Z��lǋy{X��D��4�o�R�rȅ>�?V��׌J]
=��B�ǻ��H�P��"�q�wr�֯��4T�f�'S�$|V��Ql�P쪵W����V�;Y-��^���uJ??��:w����x��n�4+C`��b{Ar�{T�����>�"0K]����|޸�L{uL���愠eZ���U��xg$W�XP�h��a��0��Mj�8Oz�%�M�5|��`��z�Q�NbS�O�����#82���~aOO��)D9P̧��:��>��
YBiR}	=Z�ٲ��SM丵7j�g�$q�hg ��*��d#����z�<�a�m����7;��Y8�����)@>g��qɥ'����-�9��~A�SJI�ډ�������Y�N%�&8fNޖ��Z4?`�t�/?����3�\*륡�������ӹ�O�Hr%\;��&:�d���:�c�b�GXݜ]�9x��5�P�&�y'� �zDH�W��u[D/�he�y)���]-
��^3��m���YP;�g��s�A�njN��O��9�OmcCO�g�ݏ2Q�RJO�Q��a��"��"U�{�-0?{���`��&E�R��IJ��`�G�uz�3"7�T��_���GV��t��%r*YU���X�c���R����cOsˢ��.9�$�n�0̦�ܸ=،gKE��<�Щ���\p�����{�\��5�採7��^G�R�
�����'c�1tH��@���LZ.��ې���mL��$��U��ؑ������b�!�Jo�A���+��1
J̐��!���n�"!��M$W�`_�i=�D��Fe�8}j6ƞYkmp��F����8����^���:Q��T�f��/�+��HHeq�$��/J���,���h��W�w�YX�C@���E5���S'+k��E�&��������Hn̔�b�=wn�R������rF�Cy��vz�$�0��PE����DVf7������zM2��E�8y�~ȭV�X�J�ůy{
mD1��u���8H�xXs �1��`�Zѧ�مќ6kK�kp����^��*��_�z/���q5���pj�r\k�8����'��RS(G�8�Yɐ�~Y{��r:J�I��h'/��� ��{�^F����2� ʗ7��Ǽ8bX?� �.y"]�	�{��Y*�Qź�H+K$���x��k�=_��$Ì��'&s��Z8�=��X����^�^$�(�[���sU��:�0�� �*��Q]P��Br�ݷ���;<�#w��ND�P���e-��a�兔<K����7/b|�(�W��G�ʆ�x�=	1�x�d��)�bD���J���3�ukf?����@�ͬ�d�5r=h��͜�=^�?���6�njeԟ�:0|"x��Q8qh�l�q��6�i��#:�g�n��C!B3t�Hq5���<wd�o~���/�֏�6
C��>�`Wq����g,؅�9���?�])s4¹��(Jڟ��i�jA Z�u׿��%\�D����<C�V�wj�]� "��ׇ~��EFS�x��/����j�P"��G�Oqz���F����"��IlLC|"�Ӱ�d�}�H�J�H~����l6�#z���VL�E�H�w���v�n�(N%B��ۧI����Isj��P�>��n��%
���o<���RK;]���~�ol 'ҞS�7/�����KP�i�"��pUq4�'�����!�e�$M�BW1Ӌ��c�q���(b�%��Y�-��M�5�����^V's��[**w������N[()��]�&I�s���*�i��W�+���^P#���ƽ�;�tT�-,�\`�픙�}�P��Q�.��.bv��,�O������Mp0R� d	���~!�v��-JB2��f�c�R{��	� �F4x��g/5��w�Ϝ�G$�p�k;a�\��.�/ .ԇ���=�ťHk�فq<+ԙY}�X�
q���*��m�W��@+{�L�l�ո��a�Q��.�vGs?=w�dS?i�����:��J\�n{�&1 ��@���vr���.)]�Y
�Dʺ��(~�m[U������v�i�]��h��p��S"#g j�d��k)��Y�6�	JF�DŦ2}��$l��8*�3j���1�0�@���G��?�~��)����t>@�W��C{�WX �Z�]J�zX�y�#$�=�����Aa7Z�d��r�uf�a;mG�J]�%��vo;�SS�њD�|c�g��k�
���Gz�~���A���u���H/�0�� �x��&��K��Y��n�m���W%zx�@�<�7���M�J��i�C	�	���G�S��}(6�����l���'nR~�n��(����h_*"� �Y���j��"K�W�%�^�����x�Z��=g�4�����~i�V�x��3d\��^����JI��y�ӵ}H�%�T"����'����@Z��9X��gQSS�0ַ�H�e��v���Q7��2���z��%%��M	ESX�a���+r�̚d�.�T�'��2Ҡ`?Z����\~�a�=���?^�7�Ч��ZM���ҿ��}h�<]h�*��l�X�˄�y�ҍ�ͳ�:1PE1�x3?��1��>^�k�ժw@8��d � �,jR�2u}*ӭ�J��S=�(��k�d�-K����M�C9)��vAz	�\�S=�(K^][�Mks��2���S,l�pʛ~�޹ݙ7C�-�T
}��Ϫ�����f9����"�D�l�����%�N[��������_RtݩU�GB����kv�U.m��u���Q�Qy<�Ig�g�T�ǫ;#PP�����{��b��ʷ��Ŋ�Ny����O���b�fV*�D�X��s*���>��zx ���1ಀ(IS��և���AF���ݼ�Z���aC��,��VtWd��s�hX�OR���#xD*u�t/����gp��._��&��ʛ�k8?�qA�2��|��RO��(���S���@��n��_;c�Lx��2���"R�t���tR�Q)C�^ؘtz˾s��V��:��Q��<k���b�e����3쩁�h+TR�=?�l�D��J��
����	{��?�@��v��Ak��$�ZI~xS��h^�#��,�A�Á	Fh�yՙ�����^@A��L�p�p��  ��'ɉT/��g]%������3�-�Sh�\�8@��<�|�7�H�Jj��������jaS9D]�M�J�	��uX?=��$b��G��[ �?}n���Ȑ�D�/a�._��⑷� d@$�ڗWj��h��S����V8`�짩�5�LKY&�̞�O��EiE`�1��-�� y�(:��F����FE��>~��#��<���|Ϧ2,��5 ���'ŹIoQ�0��V��qլ��갩�\�kx�3
(���_f��w���I[.E�D�~m"B��b�`Y�%p�=����K��׍iMG����k�~h��[�������&txn|��\��ی�w�RTM¡E�پ��֐����@㨄�U�X�Ӛ^;j$��n����'�h;e�i�\��Cz��O�m��~S�l/���x�R�/*�(��&:{sK~L�T�4cR�A��ݼmJa-8��Y����?��>u����jv�}1��Qp��UT4�e-i$oC^�I�G�	�dG�Qm��G&�f����-��h-R�
,EV���>A�^��Z�k�Aej��� �[]�h���8|,�Y����S���d�#ԭBM7|��1˼�g�?2�󃥀<Ds3�۳�JE�\o�����@>%��XV�2����1�-�V�=B�6�DJ�W�wÝ/��d�� �S/�&ddи�� &w4fv��7��K�a�v�I���ר��́�Bx�ǡNJ�|���:ǡJ����"�š�IH��ʭ���@FT]#�l�[�#p�Y0�����G{w̺�!��;ͥ�L|��J�ʻ���uh��P5ja���SƵ��B'X6=�d"�l������G�Yc�w�~�����\�����X��r����C�_<Q�5�X�V��1�JG��K����"��N<�D�mek��M0�I-�J~AX���y'�`5�G���ص'���9�5��<H�OirO��ƕ��gU�Ҩ�X�24���7���Z�����-��sڛ�����s��+ȱ6ĵ<�c��H������1P�Y���&���w��*�ʄ�T!$��y�:<�T�̫mz�/�cR�1>H�xPB7@p����@u�G�[#B�0�w9��������m�Ks\��_F�.����Bt]�&XqT\�["�R)b�I��J���#m"�'�R�\ޡ\�uO���w5��8��̶�ˮf�f���z]_\Q �b�]O�ʷo��[1FIӣ}��[�/=��F����:OH�)�=鼓�Ve`�) �qa�/Ц��`�����V,�-�w&o�����O��Tz]'n�q �	;����t8����=`Z�4�%=����G��M��o/�vb�������B�u��Q��?#�3�s=��пG���8��-k���N������򀂐^ot��)^J7t��N5�ېfB�$v/�>=u�������~��O�
*��jy�L�Z�߽�L^o`�l@�R�R$�n��)bX��/�ʖ�*�����nVZe���,�F�����)��V%�멌n��3����.��
�J?H��%sBң!(�Q�$��B�&�?�ʴ��ǩ�����;���|�T����n��ݯz��fl�?�E�[J]S�\���O]��2��4L��L�Ӿh��:[�pIX�۝�Y[���\ z~
g������z��+�*�����jj;O��S7�"~�#:@�� ������ছ	1Er2�Q����kcC�b^�����0�#P��ɥ>2ޚ��#�V�昶A*F���K�'���(�z2k�}�4L-M�ͤh��"d>sx�/�u^ �����Y�ʱ\G"Fh���rK��q@/A߅65�PH�3�mA)�(���hW�h���b��|o��U��E�H9UM$X,�$���z�k4�4~�c��/���_i�ց����V-Ķ?.�]����9�q�� >�����	�(y��7\�ĚmSb�G\�tNp]�D��tk�C7�n��I����w��ֱ�h.�7
�,��(J$2=��C��l�P�c�����Y7q�Et����sՇ�㖫@Y_���^��Γ��x�(���G�>��z�N�up��g�S��'�J��%՛Q�9	R��b2ў@��qL��Ew��
Ty����`F%B
@��]ɮS��������Z ,G�<{w2���2fX 5)�35��y�����q��y�6�q@�k�.K��8�Z�O�o������.i�'G#
fO�4ǈ�ka��l��U�^Q����5�-��e��G��`a��7�uvF���%�c�q��Z����[�8��l�S�M�"85�l6	�F�/[�.�#�Q6������w `W�- �Z1��#)�V�� ���%��e��h�Zip������f� h���gy6�wpQ��Z�2'EѶ@XSǴ��7=�J�R�V�e~g�,
�7Т�bӆ���c�f�K!9��o��r��EmǗ$s9�|����C���Q��B��VP* oC���+�!S�<��Kd�y\�48*=�-\�k�TW��Z�}ʧSC�m���_��
Pkl�Py�'��ƕ(�n4���k��,?���/C����`�b��Iv�8B�Z"� ]��&��Z�����C��H<,B{#B ������������Z�&mY*���Z�s�hq�f�$ڤ$�]�$G��חX�s,g�m��H3�>��Ҝr~��z}�l�I���{ٞw�a��a�V1�e�U��Ja[0��su���N��~
����pz.�|�A�{6�\���������H�s����R�*�A݁�_�(��g�j,w�$Ӊ�!��V�ud��6���q�VNr��%Ed�GI��bc�	\y���Q��vTR����Apl��c��o�ܳ �mҀz�?C/��l\C�~w�i`�	E���A���P��ʻf�6��������������;��_m�'�TT�����
�޼��a��7Kȷ�$���[B���NA`ӀX�q�xw�`����_���H���l-�J�o�͜��^���X�ɨ���y������%A{�����BD����49ó-�i�D>3�s�p0cRۨ�&�~]{\���4��׵U �~f_-Fs���
D��Mh�Z�8��zB�=�/qw��쟔.#�%G����_\�5"����F�
��J�O�B;vG\��p0����@Z��br{�iTvQ��p�ַ���4:ή�ADqdN9��,ġ=�F|�JF!�p�"�0���օz�r>^N:owf��G^{�H��vF���O�s�k�nY����6�X��w���gR}�����=�@�(�����H>�I���*�N�'��Z&}�BoR�)�:2��hE��I�R��g�f���M�J?�h��F�f�m�G��KG,���wI<j������Za'�wP8s����åuT��8�
�u���]��r���ہ#Y�Z~c��,�	�S�7�^B�Z�54�z3X����+�`X*�I�&�ez�V9�<Mj@� Zhb����T�czC��R}�K��Z>���U�K��@�y��U7x,}�Γ
i��t
}h�Wk�~P!��r�8���_*��e)S�����cY��{.�9�A���2ׁ!K�0; ���*�,���w�{9 �L\*��N�"Q}�u\8,��X&��VB ;�E8g�b�n�F��$�ų޲NeOG��Y���[:{%�����	�l��w(�������D�ne9��9V�� ��y$���x��TD����}g��IU�UJױ�)A��O�ޝ*��8�ϼZ��oG���_|�'5&��x���� IQCI���/�R���v�M`�y�|̳�P�Z����u�[s@��@�����H"O7�D����8=M��3�S��H��=Z�2G�2�z���t��>œ�VQ��T���VR���E����pMԕD��n�A��r�7Mqe饑�}K?9�4� �A�%F�>����J�'�a߄騝�k3�j{S����+˿
r<2�O��|X�?��>/4���_`�&�� )9?#W��z����{�g��v ���* $��ed�ʣ�)�u�a#��%ʖ`�\E��1%G}.f��y�G�b�(��mk�G�`|&�"�����i)��jʣ%8��C�Q�~�����/uo��\\;h��� A���
�Q���5f���K�B�?n35|������IY��cT���\�1XJ˂15q�t#/-_��H�,��XdGI�ʶ��!��q���"�/�7�n�-@�d�N$��;<���P�_O���¸P�ZY��~�дL��Bnګ��,�Y0 Ia�b�/�$���s���I\�4����v�X|��:O��
�&md&w������7�S�B<��a���Ώ���߂o�&Z9Z)�uV�Cܠ��\;�Q�]X��<�0�+��VD��B��j/WV�c���:�}o�T�z����E<�r�����������)Һ>�l)K߇���<ͯP�E��C�O�<)������L���X�d�L�x��::&W��j5�������0�1F������{B��4\9�)~˨jG�$ؑ�sT�2��:�zAc������,5uD��f����X[&'���2a�m��ٻU��d�QC\�
lI��r5m$p�-D.�u/Ĕ*�|�_}�u
����#Z�����P��?/H�������
%=T�{��m��&�K���Pw�7�X�{f!!
D�T��c�$<�X��-�ޛuj�1���'�U�?�H����Ih�s���c>=�lL-9�lu�v2.'2/+�h��}r�Lr��� �f>F�<�[eWA��ӿ���n�PG�jgiY�sB$�t��(NbFXuOӇ�3������� �鐹���ެ+z0p����9Ax�Y'R.��9�Z�'��݁��T�B:�W����Ă^�F�V��g�dG�,=Z�u��ad������ZJL���M���品	�)1v����@'�e�� ��9���ЦG�W�1�ŭ���rR�V}�Mm� �Pk�rKk�r�Z�1Zu�!qД��lt�Z��^͆�+\��گ���M�Tt����"�B�[�h8�cA�\�D	���wnz�%��7�#h�7���\��Nj���S�Ka:��}�8�,�Нr�����tv�ӂp�Yy����w���g|�
�Δ�������}�3�:�ږ�	x?���^�S�)~�r4^�uvf_0D!�ڃl@ԏ��@ts���I̊�MJʙB�g.��4|���O�25��g��5V$��}��s/���%�n묱����Ak���[t��0�����*�pl�
>�:��諐?��޷[��`�T�|
�ŵ[ϒBx�����.�f�� �"�o	�Z����c�z>�Q�'�+� {?�f7��~N�����P$��QG�g�	2s
����	���!�ן�:�ƞ��>�F��M�3���ʋ��yؼ�I���������.�O�_8yБ�|�\[: �xșx!j�Ż��4{9h��	ɧ�.��q�з��EO��9�O���i���b��CkҶ9�`�����ѭ�$*����n�y�|4i��i����%5�Y���66i�,��K� ���I4>�ޣjX���,��&o__��Ý��L���5G4�#��q\i��p�i��*��)�T���}1J4�C�	,�� ^�����a�)J�xQ"DP��}M����{��gn� �1&�9*���/y^��(�_�2#�'̲�P�K���i9������!MUW
����w���ݤNY��j�a�]'��HKg���Ny}ΉM9?a�te��*Z���+����N�]�@�q2"2�x��1"AFbݝ��\�kZ&O�ύ��R/��ɓ��#�Mr�!ݬb�B��b�Y�:��O�p��X�+�6o'ђ�QjM�;IX����䣩'N�F{�#�n�(��wt�<NV�M�C�xu���.�zk!W�<����{��p�O?��B�� ���ٕ#<,eը�5Y��X�
:�Va�˦�o�+V[��%J��%g�.�O��~5�~�<8��O������x�,�E.&��#�u��8��ҹQ^�J�<����� f�,��Ƃ7��P��R�-�L���>7w�8F��C���SNl�B�g�O�5nn�5l �>v�pn,���޳�y�j#�0tJ���t��mߚ� �}p�K��0s��t���`��zIB�{�	ƨ�h�$<���h�B��tZ���S����`��o��SN�pK\�����!�E�ԣ���Bu,<�M��`k[~�{�b�0W?*ɐ�+��f���廯��,�A��ȶ�z;K��(���7�kvT�|�F���ʎܫӆtm^�[���gtδ|'N�IS�@Ĥ�w<����:��i%{����L1d�XwR/Dis���<�smB؅���u�b��Ym���,F\x�,Bу:������/���+��C�/��6�1]J�v򡷪oa��%(�Н�S�J�~�Y�kc�@���V�|%2���2o�:�Lȯ�W��bf�/�g5�����)��9_8���(:4��/5iN���&���<LK�%Ňi2��l�R(�S����w��|y� !eM�eӧBˬw,�䚄ռ�&x|	��T�K��H��*��[/�������C��͒p	�dvK�4	Ţ����ү���ofIRX}mHiLG�=1`�{�l��r̔�bK-�@)�^*�
b�2����	�fh�<��q�>#Tmk��UXZ��|O?����X������AU�7Om���� |f)���ذ�o_c�4@F>�'�:@��MHDh"/I���J��7u������H��Rs㐚����~��4�<�q��wY�����/�3u�z��"����W��;Ki�%V��?���8pς����4��Օ�oal�c��<�#�QD��.�`�h�<���ͤĬP�eq�a�;c�1+����x@Q��Ni���L�/���O�3��1�x��sg�����1�(a$i,L�R�ho���$�`D�M�����Vn??VJ�m��z?�������+ym�R�1�f�!M��3��W��:��Z���!3��۩V{Ct�f���Wґ4��gN�(�/����o�'��׍�?�Co���f�����l5�G��x^�
�m��gѹN���RZp��{*�!字�Ы�C!�T�x��}Zt|�hZ�;,���y���hN+����GW_%�#͟��K�_	�ڦ�*�W�S;��B�&����� ĳS�
��V;j���;�|F{��F,W��TWIAl��	��d����s�<��X��y��t��є�k��	�~�fЅ{y7�}����M�VX��T-�ݟ���zK_����2ѧ��� �v��,��@a�D�F���Q4�^~�H�6���>^埳~�O� ������
@��i�L����vW�b�u↺�	�}�#�
�5��C�
�'�X������BK�ҍJ�n�m_8�?�6-DjW	�O2un��x���6/��q_�b�/>"�}�r]�����m��uS�P���e!U�>f�U.���̱�G�C�F����m�޶q�i3�)���?�6��6��H�S?��8Ic(�'��	*�l����G�����С����M�P�%Α��W]�h�#�&=���@�煇C���	#[2	�fae_S#�H��&��X��D{E�W ��x���Q��_�ް$*,�A_�܈{o�Z�t|+�s7!� NF8���&�#�҂-/�.Ă��{E)��d�~~C�VБ�w�a9�2(��c�|�9��5��_�$� �rc�/����}���/�̠�;���-n�9:�ّ�Ҥ4�D���0QT���@�[��D鑧H᦮6��'�\���$� �o.�8�5�
b,I���2���l�2�z�(�0'�}c7Q��?��l�V�3@#$I���8O�J�}����=L����*x��@�H񊺋~5��z�I�RCZ6�M���Q����w߾)2��1`���s�b�W_I�*���R���f��s}����^_��y>��d��r�w?ޙ���RA�/�b�s�A����}�^���G󰜁���E?�"9�B�_�V;�3+������-%�t~�@N���Y�����u&��w-�G��AA{(`tZwǱ��#���*�$��Y�Cq#|���9�D�r=s��h�,�'<������؟��k0)=q������%.RTa8�G�ΣB7�p���|�UG��$�F"�^r��'��D<��
�z��q�NE	�~չGb�� �,{��Z�pTF5W/ ��;~�����Ц����t����}�^a������*����x���Ľ�FI��R�	o[)x�It�{��Z�@v|[�tC7>b|��]`�G��nh��
Ξ��.;h�K��l;cn�6��$�{��CcOb_��z��O�kD� k�کS��V�GO�a�ꚴjKtp�����V&�	j�0��,�R�s�f�)��� G�UU kJ�ϩUX��>����
D?P^�[.&�Jw�;8φ��+G��"�8L�����N���/>*��|P�fۊ�5�/�Bvsw��1�$M�P��y��u�y���%�`J���aź�����Ҫ�vɦ����ʬ�`"��*+�x��?��� % rϋ�&�wc�řޚB��`_�Y���k��s�gڛ��z���r$�H-�~Fʭ�� ���è4�Zcc���)VN�`�L���������L��dG��I|Lx�e�,�����j�(ֻ]:Z� �mm��{����qR�gC8;�����K���kG�D�?�E/�C��Py"(��J����hB5���,d΂A���^���z?~-c6�r��� �ˁ���+�J`�RH=J�:��l}��x��8�Ț�B6����75po��Q}�|�������#~��Z 3��"F�1������\<Â���|�Y��q@��r�^�]x���ZU��䥠��1`{�b���i��~�y:��I�ZU�����Y��!n>�(�thE�6H����܎���S]����']���׾ӭW�x���Z!=�ZL~�,U���J����t:�K��~%�+�qm6����v�{4��s�VP< �o�]���<��ӫ�h�|gAm9���;@0/����[��v�u�]R�hN� �Ѹfq~K%f�V]h��q%���і�������]����m�+�L��)�t�H�k������;���n>�T��$?�\��MF�Ĉ�oa�R���;��i\��uTMj�kk�J��J���(@�#�\�i�ya��z���}�u�6C a���{UDܟF�p��	��`�HG� vG����`�Z����J��q�@��֘@�������Kf��u_�������J�&ZY�h��Jȉ֖P�:
w`�Xp��
)�5O��w,5+��(�Hr�9ѱ��h�*�7[bG��	�|���1�٭d�UWKL���k�����o�$�偡2�.+.���@�#�fb�;S%����n��y�x�wbx�'qꌃ��D���J?;t�V���ɽ��V
�#���ڴ��q��3|��^��
��z� �yOȉ5.���޲�ȓBQM���2?_W��t\�')?���t}��J gw��:,�D�lg�������Ku��%\�����?��	�����_����^��^�׫�.�I�.�,�3��_l��۠�)n��g����OwR�ŵp1��� ҿ�$S�i���n:�j�.�e@Yӧ��^��2�T���s�ՠ�i�} j�F�[V⋡��JK:����d%�h(��Vy�+6�48N�?�XB'�ű��)SuNA�o�����<N��X��DLU���#z�'�A���44�؏q7{�m���t	.�@3_r��ph���WC���[I���	[�rC=���e<����˕�b�}�v�pt�~�6�*y�}���wF�V�n��{f�7U��##r�S�Ky_�*]c�h�`A����Y�N͒�7��m�ɫ^rt+ '��;��iN#ë���=�j�G�ok�r�B9���$���0P^���VQ�˻��!r:�R�쒅�R#�^���D ̓�T��d�:O����"`��U�6��Kǽ��W�;�$�|xW���`H���)���&�yJY=�ڍ�Dk�����a�'v[�۬��A=�=����^)�r�]c�~�>�У���	0+?o�_��P��:��c�q�-�k�`��"�?7����C���/ehdb����3�ɉ��@��0�d6d��Ƙe0W������w2�afBǘ��,)ͯ��g�I4^�h��j��)��B����6�Z��W�<�'��Ջ]���8DW~�
���!��h�/ �:�SPӝ���4q�����;jP"����C֎��
F�c=�L�q����jb����5��J�sG�V>��ڴzw�{�A#F�n�(�����{RKЫez~6v�l����{���u�)���f4DY��ϊ�[N�w�}K��.zC0���m� �i� s+����
O_���瑇|0r��6�%~�h�β��	��a���s�`Ͻh���_�U��w���!����Hh���v�L_��7QO�*(ς���(�H��[���i_$�����"MX��P�;� �ߨ�\�N��?�Do��1� i��Jm�. ����B�V!*)�L��� �t��+N! ���Y�B�P���b�J�'v��Z-��{����4�QG�)	�U\��vxv�-���C�*��'^S��	uH�����w@i,/��`����q�Sת�
=;.¢�by\�/n����|��90U��c.��j��r�N�y�sw,of��^AЏ�̢R�53q:m��a2��N�b���`�M�ZL���b�1��@���x
�wsd�K�xWY�Yt�)b���,1���OFlz�-�M���\p���O�SM͇�cD�#� $�_�osisx��}��y�ca��,y��YZJR�6,�2[b�B �X8F���K Ѫ���ȕ"RԀ�,��l���G����!��^����DE�1UT������һ�D] i�;�] �������:ێ�H�w�?A_����ԙe�@[�}_:y�(#]�����\�v�צ�beE��m
�L�J���� ��BUA���uWզ�i4�*�̋)t2����������)[�䤲���O��:J7G�H6d�1匰J
،��<����*|�\n�!3�{�&i�$�3���ڃ��E�K���82�($�i�Zr�NQO�9���-�3��c^��y'gI�b�0��z�+��:fo�]�kv!&��~�|U0GZ���@�x�2��S�����]�0A��x`��*3d���Q���m�DW���:b*A�n������3+D����[)-�|L������"r��b�I���r��g�uCO��u��|QtLmQ+�C%��|%ejk�E#]�b �Q�F�0`�U�N�������Oq�6t7E4ⴁ�z">C�K�_��ѳB�=dD�v��q��౻��Eu��Q�*4�I`(��&K���M/���@[�%�[����b�����;'���N� Ѭ�1L�1"h��1Y����x%���äB��)�Z�o���4�z��.b_��W#ՉI���G��$e�3�w�?�g���!��⛚F�q�n�o�^M�־�G�������`���<�x��Ze���AG�A����s�H3ǃ5�MO���N�6���ԏy5�H�������!���<����3�C�����2(n�~����Y\_ýM�Тc`{� �	t|��I݅h%��jbWY�F׊�fs�,ut��!����2�9�_:A��B*���Y+[�v��*��j�cI�akw��ƈ&�H(f0������� ��4�g����օ�1�1�؇߭>���@A7�Y,����\S��3�e�6�5]u�
X�j*��f�g�G
J��C��O��Ss��aOE�}�,~l� #)Z�#�B@�'q�b�&�s�y��1Ĭ�@��ع(�9hp�<%zP�O%�P�R9�8������T���3����.��#P���6���5��/ �[���c�S�O�� ���;�BD�w��N!�}��s�	�1H�(>	H[ͫ��Ե�3,�B��'텔�߮6�=�-ꭑ���)+Y�S/���E��:��d�ϣ�w�`C�9�
���.����F=��>�˾�^%~�lO�N����k�Ciǭ(�������Z�ѱ�%�~w?,n�rm�`(/������g�|�!}��}ls)�}���q`��p�\w��i���~;�X^,^7�T����� ��s�G��Ax���r���(w�/���3_�}���Z!�IkӨrE� ���`TT�b@:onl�e��|��~�}�\}q�)�����4y�_����[R����w␖�e���LS7����A���ɍ/E��+w_�ys�� ^�"���2���@��bǞ�_����0CHB�r�hL�TB;U2�Z^�r�4j;_�( pз��;\��d�8	Z��M�3k�tJ�ς�ky��yV��Y	&>`�#��x=:*�C���?,������2�_lT����8q7��R��ȅ�~s�5�Աj���e�۸Q�.�83yF2���r��X��[���?�;g�>.H�t���5E]�%�TM`���c���M����!0�����X����߈"+��~�X��p皞�f`$���*?늡��H�Tґa����3�I܍��s��ёR6��t�����:O�:G��}��4��D���KA�X�~�Qy�H��Ū�)��BhTH��{�x�-��H����~qQM}��`x_$x#U61�{��D�q�]we079#b&V���A<TN�D�cہ�
�;m*)��&�n�fw�*�dw|N��H�*h�Δ�X�7��t�c�s� �@aȅ�p�6!�!�>$�sƙx�I�o�X�FT��%�;.����{�fv$/��t����-���-b#�_�R�S��$�	�p5���״I�&+�iR��1x���=I��ߩ�	OU���'i[ۯ���cAhh���pa�����!����G|n8�%k��Џ���N�v[&g�ܡق�'I�qz�OK)��Sbb��#y���@���So���G7.
EFOڎ�����XQݯ�S�`��~�Z�p/Ԡ������{Oz�@ͦ�����B��|K9k��K��<�=��ps�|K�*n�L��z�1�;�a�����Z���i�3<���M�|K�|۵f����y�e����i4:�v��>��|K�q��9|�
γ�*�V��x�{K�<Ϳ��@4ߪ|KǺD�L@i����T%�`���"ap�p���]�K��Ak9}J�� �.%�1��$�$V�bз���Y�8��n�%�/����̣	&,!�J�c������~~� ף�D�S ��Q\����6���+-��H��)g��i�+���e���K�!}���uf���z=��v��	���[O;���P�W� �:`���h͒�|R�Ș��9le�v�_�[O%�
IA�k�R���!5A�Ѕ�~�hE�*���j���3/�4_ Fx,p����R?��$�c���`��]Ҟ�N�@!�|K���o;n��� �w�;K��C��|���,΀�|�?E2������g3<4|B��3ѯ�o��y"ޫ��41ܬA���<j�ָ*<6H�w�x����*<P��|�vƿP�*j��_׆eL��|Z���S뜯>��|K�x��|��ܥ���*f^��|�z�քq}P��|�A����̀�|���|�՞�o����4@�x�L+�o��|K+_X��������|K���N3�gu����d���|�ӆY<�������q��}���;^��m�*U��� ����fy�@�V "6 �,BB��D����4��̠�̃�Ҁo����|KA���3�6�4�o;n������l�lY�QW����h ��Y�$��TYY`Q��z�83$YQ3�Y3���  T��ϗ�ޱ�Gd����i�1������"�C�ܺ��ұVv1fzcOg�7�׏C�Co�� hh�.�	�̜u�f3��O/�
}�P�d���B��p��Z^PE�=���Qu��tB��O&E �(\���`H�~��^�(E	"��R8P��2r�c�*��-Bzо
��a���㠆�em���4��ٷ& �0O�g���3ȍ�¥�2��;��z
O
��+��!,S'�, �K}��Zu�����q �3l�w�����Ot���\J��hD�.e��QE�dӮ �4z���d�Ј#���$P�:�N����`յ5��+��3C���ƔȆC��G% ���S� ���~���]��^�^!�ʖ�6p]m��<�ľ ��~��T��6U��I-J#&��e����ʖ�4_��CzН�3���u��d%��?S�t$��VV���$Q�$VLI [Shֳ��[$[S3�[+���\$�VV^[S�$W�$Y	�YP�T`: ��I	�+�X��E��Eً̋	���ü`�T��`��$Q�4$��hu�^�4$�����h    ^�����WW�t$��AIQP��X����+�W��_��S[YS[�   ���2   P��XV� (��c���4$^h58�b+4$��R�����Z������V�|$��h@[/O^�P�@H��A ?0�XVWh�À�_+�_�>^SV^V3�^�  wi1{��h�kZ�G�PY�k�z�W�����[6���<,��7�u��6��lp��Q9&:o%`v�m?Ȧ�K��!pPz�o�%JfX�6�k)I�7H�o�Q��� �#��f����.�Vu�5��i"���<�W%HB8����r(}��<����ԥ)6~g@���T��Y�8�"jr;k@��&0���Nߍu�M]|�Π�/b�l��⋵~��D�Kk�ͽ#���)�<��qu5�X��襁�2�^���V�zHʦ������3"�M=6�4����iK=�F��f|_��צ;���G�V> �w.�b���C���xC�3�$L%D�Q�`�UB��~�:`Idt��œ^�p�����3�ŔY둱�('����S$� -ؑ����R h��R h�$��Q�@ 
 ��7���+�Y���$��aWQ�YV��_Q�4$�4$��WV+�^���?��V�`�$��S�D	+�^W�8���2��<$_��W�D 2���#�+�_�Ƭ�}Ӂ�T8�,��F�5�V�<$�ϋ��?���"<d"`3��x�7�N���  lSt2P��s�$6�Iĭ�"��l��a4��c;���T}gz�Uޞ��60ܱ�5N2;�m�L�ͭ� ^�ҡ���sf��y[���������c��Ǫ�#44yMC�_I-ʛm�9�[�.����r��(�FB���4x:���fi�nbwA_J�C�H�~���+,�I6�������4f�K4��ӓ=Zl,N2ڨh�^4��]�u��n��@:�.7��O����x���!�Fе7'k<$t`�RE�G��(Zt�V���Q�b�k%���|��b:�Z��"�N�E{J�P�B�qr�rZ�c^�bb�f_o��F}ў28 *�38���Xf*�1V�Z'�T���rh|2��!�`�҆����&P��s̭u��O�o��&��0�
"�/�F��3�=�A�1=w�qq��~�z���6��?UL_�B���^@ܑ���+�5�V�g3ǁ��A� ���h�Z�C[��C#�ٺ    ��1�k����B���;�"��$nn-�9Fn!�8[RV�����  3�3�13�*w+�H�Ƹ   +���%-oQTt�    `3��a�Vh�.l^^������-�->{�}  �6�?��A]m��W�����
��4$1iT�;�*�0)�p�L�|�I�aw+��V��Eh��	��췡B�ٯ��W�lshL�5a�aI���{Nzlb0� ��z��m\�z��� �){�
��r�����e�C���ZO���bUxu���=�C�w��9�V1��t`��Ы�+�h��? ���gl�y�!�(c�<����42Z�)��
����1���}�C�4l�d���<|�e��;r�['�yא�*fM����p��}���4Ђ�Fq4��
��I��,��v�����B��{�XN#����|<0iy	7��Q�Ӷp�&�z<ds����4+�3"�ۼV��R�~��vEgշ�*�Y<���*p�4T�^wB�ߐ�PW_V�$��P�$   X�W�B8�(���]�+�_����T$�� �$��ÆI�|ΆocK�����^!K}}��P1�	�,{��v��+����/%��#ҝ>���>��"�V{j��4ٺ�:�P�}N,���j�_C;l�$��N=�O"OVVX�dO( ����V�2�ƙp`k��^�����Ӂ� ,��p`k��   �/wz�R-�ѕ3F-���K=V���Kp��zFo�q��I�Eѿ�X6݂�S�|)O�0�������z�6)J)�� 2$p��B�)[q"E)�;?�j(e������e�h��3�_JK���ғ�z�=�c(����A4B��R˝z��2��ύop�M!h���s@Ԟ��~ִ,E�^-*<�`ZmZ��ؙ�ql����$S��קht��8�yC-s!��IyEʓ��z�]73_쏒���#t�4^����n�p���n�p�t$�VS�<$��WV_��   ��_�>W�,$�  _�>V��_� �4$���+)tm��Q~�+��O�+�lN�HA��޾�s���y:��r�)O��jC��0^5�H�/zz*3<6�{c�����}0l�L*�y
#N�v�}uD��]r^�/�G���c��:���k�
53�`#��    3�#���@� =�u�7�jG`�ȁ�`�f_��3ҁ�;"0���C"0�E�h�G&^���ȷ��V��    `���   +��_cY�   ��Y���+�Xt�þ�  �Ƌ���8   �D�n�   考�x�	AZN�������n���b,�_�9ŌǵRWQ�a,�b�5�Q&�>Y�QYGQ���YJ����   YQ4�Y_Q��YZ�E�a,�bQ�YGa��wbJ���   �j:�C�&�r+���s0M�);pk���-�w$ܲ�)v�l��P`������	W�&+R�>ׄ9_|C6|��i���P2����)����&�)T�.�ݗ5��A�`^����ߒ2��@��޽��<;�K_ZyWR$�P�~g�W�I0z�@	�$N�Xb��Q�WW��јaC��Nʩɾ�ݒ�47w�� ݗTZ	L��c?�k��,���;�T��;`i�:��7Y�f�>s����.c�+^09��f�,��Y��?Ob�zy�м"j�K�P7OI�OH?`9$W�f���LP���6K�[�h�P�Ǡ�>�'��Oh����%�����E #.*��yjėr�x��8�@�NA9����l�q��[z�&<��Z��8��.��rj?`�}�=���-�@m:S�Tjb���$���i@y�k���-��z+a���d@�t���&���Φ�{L��$f(*����w9]{����3��)�F@����q��l�>�#x��V���*yIiW6-��1�D��z��]���!Ih�����wE_����ˊ6M�:��:0N�:��>�?�Y�Q8����1ܼ(u��>�詿��\=7�)��?{��tg�����D�^k(�f%/\�L�
�̍�X:�s,ܞ&x�K��Yo�k&|N}g�@aCG�N�x�X�p�CY�)@�0����0��<e�Z�1�9E(�&���ѶZ�z?�a߹�塺�Pt�ɣϯ����*�p@����C���@j����Y�����(�_��L)_���+��LSV¼�V
��K�f0Z��;�2���Qm��=�\���fL*E)���@TVƪ�9�ܝ@��ӳ���z۰Q�� ]j���$cL�yĠC*׼��������p��y_��ԟ��dl�Y)L�����1�0[ Ǝ�<�t����!�����ٺ,�h��X���]����`�Hc�M������˲��,������j"6��_���vrx
��_��M��k��I�b����Q�k�0�ѻ�Aqh���h\�S
��`��!�K_u����C��?�F�,����_� Ә��V�h�f��R�_뎜��(%;�"�
��:M�s&<�7uߊ��b?D7�1���w��/�!�l��:)P�j���0Z���o�RFB�O��nTh���j���%цsj�J��ʦ(�vX��a�\�r��[�����'��nX"%���1���������2�����''-�; '�>\8�л��%沭fTS�׎��?U1�p'� ���:S��RX�G$9�$��G�*#�m3�/���kle��<v�$E`��s�m�!�#W�o�Pw� ��P��uԜmt�y�`pq a>����,{���&,�oqV��

�pO��⚣�)5����=ț�;�Pu]�)}��Kadޟw��C-�\�/S��?�ב�������a�c� ��2+Uht۱e&V�0�4r�7�������t��W�E:���l�\��WX�
@�C��no���r�G���a=7a��H�lV���O��L�c�.���ŧ�������L{<iT���y\�H�"l ����?5Qe�ꝥ���/��ʛ�g]���{��C�FX2���k�ՕE7z+0lG���L�#�X�¼KQh[�`J�����>ɏ��?��ޥ>.\闑Ͱ#wF�+Kc,���/;y�Ȧ��h>���d����$����ˊmF�b�I߾�͉����bx|d6��nzTM���K!�����2�
�"�]`d�����6��̐Fu�B���!��8�)�������8o�+��[]'��\�\P�\���BeH�aUA����`��z����N���'��zƙܛ�t��(�y���\��
�w�ӻ�dP �(��C�X���e�t3�e�b�\���3K\�-�B.z�s�Q�ǅ�Wi��Ğ뮚B��N��{�2ҷ�bNʓ(0���j���k�>�xF�t������ɸz]�'N��}j�.6^�pF{,ς�Bi���ԸwFma���(�iK࿚�p�����[Bim��?���+3UP�;�T�o��K�7Eܪ�
;>���a�wp�b��\����!��jgG�k�%@r�<ʕ9J���o��]��w�����ʑ<�{�yK�.

\Az�2��h��܍F��j �<6��4�*�e�F1k�#MG2��,4w@��p=\���	QN�/`yP�-��:q��#��=�=��0W��xR1��S��3�7�և2�ek���HI�q�#S�8/�£��&P%p@�����p�6���,�{�0rG~G�� ��3�uВZ�^b���A����Ts�
V;V]�C����eQ�T~�;E9�\O�c�z�+��ٌ��n�a�_F���fޥW<��6,���j-0H�#cD�u�[Q=Ƕ69�ݕ��.N4!n°a�=�%G����a��`����܆{�V���WB'�SW�Y��"1�1��q���"�<3%�e�&!�x 5;*�L&�$&@뀆������f5�?�b�y-I���>�Ĩ��4���W�r��ǸL�����Ȣp���# !�y�88���R��qH[�� `�G`�8A�N k���y��ͯ��I��H��_��Z�� ��f;���uy�	V��By�e���*���(�����Ewa*z�ǳ����B��mz�i�l������9��Z�HB�H7�!�r	�����1Y:*Z���fS��w�9�L�i	�nBw��I"%��;�n��*�hrT�m��W��ݗ4D}��8��]B��	<����Ѯh�ŕ�P�=��w����\��>���S��٣��j:��`�	#�U�;�V�����:7���,/^�u�E_�$.U ���Af�����1�^�D#�O���'�Ȣ�c�q�"�3����dӬ�9�A���YW�H��D���{i`Gۻ��'l��A]e�A@��w�$��T���y�6�Û�I#Ĝ��x��+ 6�n�h�mj��[�;?h0�5;�'_"o��/{��<�\��Y&��lTMё��4�8���c��ͧE��g��7�o/��=��2Ҟ��,�@|u���8[<Ԁ�Ѣ�� �-Ɔ���NMWH�(��x���h���<�L�.��A\�!�7��15홙f��'s9ujb��x^e0�-�fY |��;#Z�R��?��e�%w�V����#r�5/��6�E��"i�}�{,s���r�#�K�D�x��E(p�i�|q�nL����b	��༽C H���`�'g	;:z�}X]7J��y�� �����X��UQ���l�\�G@9�ʸۍ+Wh�K5��1����(��	�d�c"Y ����(d(�u�t���"���b�}<a��?�.���~���# `��9�%V�h���C"�V�$@'։M=m�c�.L]*���q����!g�/EAS`&����)��+*3v��j�g�{geCݢ���!�<�t#Ţ��{{:t�oh�-|ď��S����4h�weft�Y������puR���A�k����i/�
�t��S}��5��k�JY��d�M4��N��۴��h�!q:Sh���^��D����c�|�A�@�g���[��#��\�~�Wb��Io9.&8�/��r���p�o���^�_��J�r֩�%!�:w������K���jϖ06����[u��~��xN�kD�`��?[���V�;9�1�M�����sT��͵r�+O��d�������9�=V#���U}�l�&p^.�*��=��pn���u��X��Q� $;�p��y�d��
=6޲'�.[`#�Z��=�"OC�~ �9�́��Π�ݜ�`65%��wB+�۠�ǋ�*�M����T�4�y�4���jݨ��o��Y&���FtMUQޘ�]Q;
!#{,D)L��r�a�E@c�}�K� �o�2��e��)v��
�=,�'����F���
~�"z	�a,��N@`]
�V������e��WhC@�{0�,�e[?܅��q����9-v� �&���:�Ś�ky�(v�3�hv�+[Y2��ج��T�F ��/C@�B7�kB�&��3���̿�;����c�N��Y�*�`��m<sH���(a�!�8��ԃ����yV����/���l�;��量�T<�آu�tp@R8Zd���Rd��9�1��B�9�)`���G�5����J������9;�G�퍻�����!4���Q���D�n k��Y�����"���5�	��a�i���2��Qǂ�ȟj�����l n[vFs��٥�E#/�_Uؠ��[?[�X[
��;�p�T����������|��d�0�
��$�DnK>-{�fo����[���}�+��^^�s��uj�$��tw�}[�h��X}laߦL����\�b$/�pB���r�6���HH����'��U�{�B�dSy���ְ.�1;8a-F��Ҋ�]���h̫KKJ�l2�pe�!j�0�a����6:��?π٥�<0盎�H>|򵨻��W�ƛ(v���g�B���Gu�T�8U�l�/�WK��JND��t�KG�w���ߍ�LH�^�4��Gȸ�hi���h\r�K1E�9�Xq4@ᨆ�� ��?��������=��4e����D���j�+�rڷc���=(�m �C�b����~�l�����b]����dm�p��������(v��%yJh٠a���ǵ�+8b�)�l���&�.	��T�rw�ǻ�yxp�U�f�s�K5(&��G|��4���,�?n)^��0���� HX ���Z��&!����:��e8 ��7�TbOvF�l/;^	�p��R"�K
����|�#N����]&��"���z?�?�c��Ωt�0!8�����D�i��O{�m��Cx���w#�Ľ6�(���24�,��\w�AN¬�A�>MUhnٟ\K�D��D�U�`�L�KL��`_�B�̀�:p�93�x����޻lu�J������?��g7~��1�����R[ [sT� _TL��|�j����J5b�U�	�R��۟~�_����X]
$����'��%R	�h��.tQ��x[Y[����A;����y���=�	}J�8�:�$x��G����(/��I��`��_�pzFn�{��һ��S��/l��'����F�3LYVP�����6P�b|}5���R��J0H�Ax�0�����`V�s��l׼��Zg��i�������=�$��Z�'?���|���^�y�"z�B�C���J)��q8S�����K�DgA&a7,|�����>�,Ԇ�ܱy��d��a�8��>�|��r�L̍%�i�9���p�R���v�k�(�R��;;Qvcy9��l�&����RiwK���U�Kl|.yX�L_�/:*�����ֳ�m(wסL+�G�R.��O�X?՘&����
��Rp�H9I����� �*�Β���<�L��gH��Bw�?�"��
�J�8i�7�\�<�F�x�m��t�s�����Ġ3�)[����EG;�R��9pZ�Ε����½��3_�G;w��<l�!��:�a�"���<n���f׽~+�+J/&b5@M�YB��ۭܞ�^��A�p�V[<��c3�1H�S|W.>(\&��蕱ƀxG�������'��)�&�)���E�� ��,�TIA�7���SǗ5�t�d��\�R�f�c������$�p��#ȥ�i≕G{E;Ν�(��r����{���r���|1]z��9���w��)�tB«�{;�F �D�֑�c
r � ��I���֙������)��]il|B(��`W����v��P�z� �K}fE!�y�qm� �AT��� �#���J?�����G��Q�4��G�8���d����U]�+�uǊy~m^�J փ��Gan��
8��0s&���6�$�3U&%�ɩ0|�JDt;T���<���	6�)�X>��"T ��ՋS���Ρ~J�UX8jy��~�n�OefO�=��Ij`��E��/�IcJ�s�K-<"���>W�������2�m��Tٛ�9I[��W�u
� ���V�BL,Ѓ�0�9�1��+��M}�Kȱ��u�
�$�>(\O9Q�-��M��>خE���*y��D���C��|:,���ס��=��lA��8��d�o{�p�.�n�`�3������� b'��A��5���6�v��l�$�O��n�`����x/Ҽ/���{K�aZNA!�Y��5�sq�-ss��HVuQ�w�����L;�^��䰑�߯�{�(�?\ɯ���%20:����|�6�
r`��A�Q��Hl|M��r���)L-#e��&y����Bv��)�iw��l�'BP�K�K�B�ȥ�޾�w�_O��s�.ƙ��#,�8`2d`��/���рؽ-x�h\X���p� �޷���F�7��R�5�>9QM��,�X)�=�sR{��<�@��W�f;w#q��}��}	����^6
Θ�[E��L�� �f:���g~��+�x�L*Q�Y:�Ybf)JSW���XVK�sr��P4�1fe��2F�m�3z����H)�黟�Vl/��~�޸n��ׁ==(ז�����k���G ��jȿ1&C㑲�h�������r���~�Sk�޼���¹�c�.@�#���@��/�G>�RQ���S��� S��r�I	�e�A+ۭ�nb��Л�P��:%���"���d^i|�J��ц=���r�iM�eO���N%>K1�aMp���R�p��iJ���uO���k��V���A�|0�8#%LFIv3�C�d�����w·h\ŧw�%�� -�"����?��$���L,�"a���j����
�*��c7�ܩ %lhͥ#%��o;r��/mfB�L�����JxT��X���G4M�J�p(��v]���2cS\ң(6�>P�r?�m3'�±�=�,F �N�t�}JHG�W�#Ť%��@f�'�T��%|]�]/r��m����>6Y���b�v�:� ���-���R�:<��9�̳l?ݺ��<������;RzZ�:R�@-RA)�I��X�\M?��ԝ��%�ީ�YI�4}׾�\\i���Ϩ��A�'�ox3�Y�N�>�y�y�v1%ý�FX��ކH��I{�m^���
�_�1�VIq�8��dn��M���Α�*o~�N.�'_�l�H�O%�X<k{��Nv�C!�؋"{	b�������8gJ�lW���8���t�[��p��	B��LD[��Cp�[*�2�<z�� k<>�a���P�bМ�������������BE�M�?�����`��/�e�"��'��p5yK��J�v?��q-��� �ec�6Q�(
�
�
%����p"���[���+������1�ڲ|$��V8@N���,g8�Þ��|�d�/]���pJx���M�o��D�T^'y't��
����������iGj����g��n�E�9��N��ˑ{��Y>2����l�9i��2a:�9v[!��!@GŦ�����+�:�+�{Q���5�ӯ�ۺ�����w���ۘz�7li(�6���)h�!�*�eD�Q��:���wJ'd��BȤX�X8M����ϲ����b�j�|N?c'�����t�_�1�Ő�[M����ޮ���/yP�kj��f��\[���	��lo�[��i"���)'ϟbQ�X�>D��W����#���S����V�"<�.����'��O޼5�;���ޣ�ٓ��(�/����>B�*<,���@{�+�Id���q��3�<\�ZO�;���}��.sZ@짡�*��do�v ���顷t����1*إA�_�z�W!�H�c���@�A�3�� �E�p��>K����vz������3d�禆���`��R��N�����K�SD�1���m>�t��wO�}W��[�=�I[����߀Q9U6<|-����.9�ђܣ���zBN1���'�UzwD4��M@Q�?�L�g&f���F��l��Eu8s��j�U=O�-�q����ix�k��>����k@��B�
Xi��HgƆ�m䰊w�cߊ���R����Pr���UHΛuZ��g}��/f�2aq����!������BK���fԥ��M�����E�I�7<o� �&�Wß����M��6�*���h���E��7S���Z���9,}W^<�>�le��Mf��avkJe��f]y�&*��0?��Â���P�V�$�x�/�T{��#�'O`L)��A��3r�^8f}�.<R��M"
j(�� ��n�	.FN
�3~�k���~^!���"����!Arr�2�����+�T�֚��D��	E��\�������T[H%���G��.d�_�';��v8����e[�X�� #k�/$-��~��e�E.
IѢ"/�럽��<h���K3�}|�3R(+Dtp]�����<&_�x[�����ѿ�r���(R�i~ۀ���	1ԟ"z���f0�6+���YV�>Z�i�(0�{sa�������P�p�2��������l~!� op�E��Z~c�2� q3O7�L��T�L�̻��U�]���AC:iKҝ��CT���V�T�����Y�Xw;hk�:ӟ0�H7O�Fg�������H�fyL?�w��r��ߢK�}�����W�X��V0+� ��~ч�^=[��y����?�b�Yq�o�M\Hٵ����5��������Ct6�����Y���r��
�2��q�Vc��N��0��єI���R%�U�*;����*�o6X������-�ds��kEwz?#��m|wk���%1��r�8$�/O�x i�t��G;SP�/S<��X�RV�������F}���J�I��z�o��NJ&8�ӷ��<F%h?�,�&I;���8֍;��/�Via��"
��0w[� 	>��H(=欲ф��q�a�4�h��Ru��0Շ:��yq��������[����h��#�*�b&8r��e�1��6pO9*E=C��S���;*��&��g���
P���"��b/�� �TK��0ř���i�&��_�?,�S��(:)�����������0�e�Z���;�p����.��\�>}t����o�-qo���c�BG��1��#��mԑ_�[&9���ju�H9j�xpkz�'����"�9�╝�P.�����đ�1�*�y�F�be/l# 4�D�H�N�K�2�,A�k�LY@(��6:�1���}R��ך(��6X�K ��S�Ӈo哛����h��O\�k���6�y (�u�Ev��S�	ؒV^Q�3k\��lF{��xz�h(�7*��+$ނUhz��y/9��%A�'�������P �l�e{�ټ������?	����K%���鳨h�*YJw�\�Ν��ʭ���14�ԚP����#S����!n4N]�ș���;[�|�dR�������h�,��8���,]N�[�����]��^S��@�vE�g��L蝝��$P���y��R���Ҥ¾���Lb0�f;0�
�h?��+tf�|��dB�^^���)���[^�^��*��(��B�kR�Y}�N���i��H�t&48}�_�FN;���F�"�����&��6B�B >gs'��rK[�c�tw!�����A0w:��mKC�5��|�����p�H�94��]K����P�� ~>���f�˦t�M�v�o�<fl����T8�o�T2�݊㢼�L(C@�j��+D��͵��f�*2����]����X[��Mad�S��՟߈L7�j��DS��'���ؿWkݑ��kQ�:��]\���>�k\{� 5ԫr�$���H�f���ښ	0�&���Ah�q��Z�HPď�����'�<ScU�Է��%����d�������E9Ҵ?����qH=s�<55OF�?��q�����
���.�+�OHE���3̕���Ծ�������;ݓΒ`VڜƘ��}<�ͷ��Pylf&�aH(�b�[&r���8'���_���Tԉ�ͬ���%�*�{���e}�(T�C�rӍ�[!�{�xm��n� �a�Y2�-&ȗY����w�9e�D��o�1�}qz4=J���������0���dd�G&'%�����O���	�R~��WM�M�ՓFF�6um%��,#�t�#���=�$7�됬�mM�]K����3=��a�|1�'��l\����#ir��0 ����)<'��K��ř��H���Q�|l�:-��.���M�$$/&�ݝ���J�2X�e\ӯ�:�7|��wH�����o-�蟌�u�U&i�NV��:�d"�0���B6{�(;�M����3�����)=0k{`�q��4/��ϥa4���L�n�_�y'��'җw�>g��1��p��`��%�ѼƼCڿsC����,��C�t�
>�C�,,�2-��<&C�2����'���)+��쫹��Ѐ�Ėk�З�i�9��2���Y=:�����a#͒���"��������S�����}�(�y���N
ʅ-�M8SJ���R�ۯ�X$̉�Ĺw�������qO��r;�o��YP����x�"�t�rjp4]S�>9t1��K�+/���эn�p@:(�f�+�RǢ9�m��s�cM��� 	$��x���Eٹ�*y���6���2����r�mσe(�V�y�Y}�Ho1�A?u�z4x6|Kī�`䖼������(v2��f��7e%;		�����B=R����݁���g(=αA?��'�)T���zZXp@�����W��D���4��lSÝ�+)���R�/����{M�_o���!~����h#
�T�)A�A�����#{����U�͇N���P��d�O�jaF��ҟ΀�t6m*�f*��p��Nc_8�jk�|ƌO3esY\M�����?Eݯ� �����g� ��3� T����lO�E�1�P�Zc�	K�����Mb��j#[<��8`w����H�Srt)���]c7s�Q��17)S2|�(�Ѭ��dtW¡y(X�#�&�T����T������4q��D,���To$�m��/)R��) ����:�i��+*�ً*U�B�x����p������hMiJz�|�=����� ��9�[�?޵.�$�����{�N�KhY{���H촏�- ��|��Б��[ܱ�ϳ�'����Z����
tF�B��w�421�ԧ�wdB��?&��cw�l��r����5�J�����z���2q�7�v���4�`�H�_�4�H���	Ht�R�W�Sj+I��5>(���፾����~t�s=ݸ%
�=�b&��������wߕH2�q�w��>�!�fnc�a�L�Y�2n��@�`|ܱ7R:����o���Gf�n|����d��ܵ�����.P�)Ax$�k�(f�4�q5;r�)e�&*rD<b~��7"E�=fh�`Xo�킵Cg�� �(��vM��d��ƹ3k�.|ROP>���Ao���31K��	��N쁚��r$��^?]��g��U�+cZ�,�9�1��2��u\ŦV���ky{�dY��
�'
f�u�df��W�W|��2��gU9�o�CV��p/�t)QS�� �g8|�?�30��9342H���χ�Il��5</yB͐���Z��I�u�����l���h����$�0G�j;����܇��HZd�V��@7ǒ�}qJ�
�q�&������j�b�gl( ?y���s�n�p�M�0�%���՛�	iR������ϣ����i����kp�el:�8�����Ų��C��ŀ#ݙ^2�0��<	zU�?��	4�H���Y>�ig��"p钑/�,���1�����l�]����P�]у�0+�&�	o��*���de�|Rڇ�x�בP����q��V�a�*���?��kD���̈́�J��6�� b�~a����o���+�ԃb��>�I����.X�KI8��B�����f�%9`��G�L�ws�a��w8�r
�x6g�C�i	���_ȟ�����zb	�YQ�í�����w���`�H�x�pg�2f�ƥK;��Y�3|�Q�(�LU�1Y����Z%2 ��Ƥ%��{�
���`<;�ܓa�^����V#�q#Y÷V��n �kx���1@���ĶO~�eM�@VO���#T�x%�!`�Aosɯr�'l��^W�B�묤�eUp��!Ȍ�Pn�1�w���L�����Fa�z^��%+E�o��z����{A���ݰK�ξ�B�����ot��:t9t$ #���7�Еv��h�E�?�)���F5G%��X�^��9^}��o���-�1h`�j�i6&�w��y�o��yo��tT��n^UBi9�K��Og�7��p�9�Q�F6��3�Ow�Q��c��5C��\����aq���Qv��mS!^%�p�C��-�����1�8�F\�6U6�e5n��]7�����jr�d㈎�4�9j��ߪ�b킵7D@���˱�ZWy&8u�G^ݏ�QA󖎩�h�ڞsNP��%�p\�́Ozp\�?�������2<e��^�:dw��^�tI:tuGj~gWJ�pOW�@�R~c7^5��c�׈�<L�^��ލP)�`57h�U�5qJ��iDC�^J�@ ��5�AĲ������3���y�Й'e\�EZ�{�[�ט�m����Ы� 
�\��1��͹ީ�� ��/��՞o��+)P�����{��^C�wB�x=�$$���2ܶZ@�i�\��L�ٿ|�!�9�_Y<��N�3N��1�tґr�䑻�(��
�kaE}�%d�:����j�P `�v��+�|��o50d�>³7��꯫%3�*�[���7={L.�4�ݽ�;��#UZ����~�~*��
��FkВ��7��+b�*yͣS�>@�x�r�~}�����d�r��q��z�4�h�&�y&�2(��Q�ݾ�T!4�|�^��3��'p����Ht(��)�<;aW+�<8�y�l�{�;;���~9�N_eF��K�5�{Z�e)���
����ʯ���3D��
/,0ڌ�.�B��>��[1 ��bG�N�a�JD��+c�k�F��vq<^}Dh���u���w����X���:9/��x�7�u�~�%
")�Ug�w�ꗡ|�W������c!̰;=HA�0�����;v���g�)��w�|r�)p��-������~ɜT-�ܯ��l��n`wI<9�۴����o �!:�ĥ.M!�z%��ѳm�1�v\�������6�@yZ�E�¤>�2%E:G���y����#?��)<��>/�����cxn����֠��h�@�k��x|�[�R�Ɔv�Z��qyg��}Z��E|1�9a�g-��C[6BNk�&����G�����
aJU�A�k��B�������O@b��!yT�tB*��c�L`��� ѯP+��Y~P�ӹ6�}��}+����6����,�p<���-���� q�=e\j��F������qj�hP8��x�(����w�'ˑ��VIͤC��Ɯ�r'��aF�<��
tGл�����5S�%x�|��%5��i�PP
��g�Ut�����A�2B@�DP���&��eL&b�Ѭ�ᄉ
P/	2�|(aG_��E��K�M�-��X� O6J����/�[���1���缀	l���=�	fl��x�5� F��G0�{^�=ED46��c0#E��5�aԎ%�/�z_J�X����#���y�
\�6��3d���}ľ"��J\i��bq��q�

v��gn�f3q1�y��������dI�`q	���b"�\����L�=JzxT�u���03�4�ڤ���^1�׃?	������@�;q��~ v�(&���s�	[τ����b	FEsu���Nx�������q�f��_� �CiPn |
���͙�U|�/��a�"_�d���kgK�rYֺ�G�vp�߫�� ~���9>j҇C�e	�8x����T��g��XI�����g��\��x��T�J�����������k�#�u�`�_����i��� ��P^5�>��%)�����������핪�0�I�3���$.�A<�?��)8↘|��DƯ�.�"����1�U}��������j��f7�k%E�.���Ri��"|�k��
�L�fi��W�u��G�7�-`��Ώ{�b�V1TY~y�����5����^ϩ�' �	<��uW��^ݷ�	���JV���7������.���9�݂���*�	d5���G�%����kIn���'��de@����h#���㾴�ȚVg_<�� ��D���.:�������x]+�>��wƉ%�Ϛ6|�,F&<���jEd��
��6��mü)֔��,��?M�K��2ͤ?�q�35�q,T?ξc���J�&�8�l=�������ŉ���3�9~�L�A�u���3? s:��{tEW9G�H�r�4K^_|�l�P����~\��T8c' �`0a�N�VFR���6`�f�t�����H��/sh"�$�����r$GhC�(��'%1���:�^�E#;��/CP~�I�	n�,h�T�T�X�wI/ p�h�d�ǠV�9�rzx���짂�=���	5s�o����z��� v��t��b�oB��ۨ��_��r��R�C��\�-�8e����>%
�.�y����!�!/"��Zmүu0�B���$48�wN%(���
��گ����jI��Gpq+��>F�����v�k�S:U\��u.�`�ʻɩ�*.�8�� q��]ܙ���([��|������u��޻o����1��3�(�P�r����'�/��ǧ�tk�W)i?�	7�`�0��I+Z�,����?���,��]�[|��O��Zߗ�=�[�/�w�Y���c����A}K�o}��_r�y��}�/�a6����sV|l[V��򢢡�3��Lho���;p`d�O8���(��wv��g�f��A�$�V�:���s�2����I�'���;�\Sf5L�F�9D��D�h:d�2�0���������D�J���}E�*N},�a��e*U��Ȉ�����&�I!P�E��ذtv�� �9������ěL$�*�ˢ�����35z��Jsi��/'a|�Jn(�![��K��7�{g��E���ư�5"���|��/_tr�xC���C�C6o�:hn�^�Ee\X�:J�K�O(f��L��R��+��
�(5�f��g�V�J'ٷ��Lg��s�z6<]��2�<�bO�����d�!7B�Xp�l�_�P��/H�?+j]�Ug;�Wvl~?�Sx3��l��-��*��'����4�rw��,�<�<�����=�5<(���V���$6��~C�t�X�`I�!�_���:��_��I��̠��Z��#�w	����D��ы���!f�n������0Gx1�s[�f�,N�P���֝��֛�2��D��̟���6�]r��s���C^?=,�)~��z�J=��B�X��!s,wl6���d�M i���/g�ò��l� �&`y�����t���<2[��Ӈ�.�����u�Wqhs��e��9p����G����Bc����
����YC�ml2Y#��x²tN����e�߬����Jrh�����)���}�-�%�%t���Qj���
���l|:�-Cu�5If8��Q��Ϟ�3�'
�:��bߴ,,��)N&���"'��?ߒ+�)�$-���瀹ֶ|�vñY��ۻ������-Jk�6څoӌS�"h��'�ϓ����������|B���γ�񽵻��7ݴl�{�9��y�*���YvV�QTNța����wc�=`4)�0a�^�
�-reS�	_}��pue�S�[0���B��{�{E?���2�g�Ͳp��Y������c���Z*\=)Y�q|��E�yt@}҅ү�1�Nz"��8�^2��ڋ�"ӏx����b5��ZCDV�,�¿���ӫ(:y��Llͯl*�K��Ӄ����%�����]9���g�*Ґ�U�0q�<e\�]I\D<F�v^Bl�]'aXbS�#Xj��Qq{���Fx7��DRe)�RLHw{+Z���jpK�;���s�d��r�����!�)�'��7���ɱ�7Ig+}� tK�fc�*�>zy��g]ĵ�],�6C�)����Pa��,<'�p�l,�ρ]h`���]%� GQa�?
�����Nr2�}��]�Qȴ�:�d����$;Zt���:O���W��	 �P'�L�p<�k2hZ��w��+v!���3�""��w(�e�|�yܹ���T��`�T�x���n�q����j �Z����[|lK����������M~���j�{�agf�ج��5m�#�pxt�����b�n@u�ɠjJ��3Xj�I�i�z��~�t����fI�������������tx����]y�N_k��[Oq�{ߵmk(�4o�;}��,-����	a0��@�3/�^��8_M�+�F�nT��(���\���c`�!{�
��~q_C��^�H�}|9#:�Ew݃��MKW�jG7ez��n��G��p�䀰x������e��	��J�kCb��3��K�q`F�q�-�9��;�G���6�:���t�H��HI;k��c���:���gB���E�T��=$d���7_��5PczQ�1���R�"�:	c58�����ݍ���&��0��C{UU5[���p��P���r�i��uLFŹ(|�P"�xs�q�I/'��.}x�pq��3*s�&d�����(~iG;5�ZGw���J�0>_䓺�S�(��k�A
�4�5��$�az �N�t��J�d�~(A:��(Uj���^0�e��m5!��k5��/�rSU�}�Кgǩ��c�x�Zxb�^ﳷf�vk���Լ�YJ�:�g5s��!�c�61�2�M�_:kk��l{x���b�9-�x
�����������@םS1�p�x��O:eǑ}�qf�>a������!CD�Z���p��@���_�:���~"��"�ĩ�"�%�@Z.����Z�tZ��T�@,�����G۸��J���yz�
���	��ĥ�%R��F�K����;�{u�����a�{҈yα�S�����+,&gޜ8���2�aFs���_CE�צ�Gxu���?0�!�J�c�Lk6��������ա�պvKC��%�6|�^r�	��
z{R�,�ؼu.P��­�fb�6��T�Ȗ׶���ش���kġ"�&{d{6/|�ʷ#i��F��0�8�~�+;�y����/y��l�� �d��`�]��)��T�u��J��(���+o<pC�PP�W���M��k�
l�j8I*Ue&t���L6�
�O;����n�ʃ�?r�/g�N�"В�2�7_UZ��Bo(saANC��2cC�ף!��,�V�2��:6?��c\�ߊ����+}8Q�qY�2�|��?ț�'jF��;����h��&�O��F�����1'�a%c'�X�Ÿ��cۛm�v]�yvdK@��A"O�al�n����R�h��=�"�W@�L��j��[���ޱ�\��fbX���\g�5�v�e�A�/���'aQ:���@��~:mR�/����ɑ�@a�^gj9�pIۛ�O�sw?/0��}�P�a����1����fi~%�f�e��?0�ɬ���M�$�g�!��+�˥��k�D��{�d�)�A$�+�m�v�,E����m��`m�(l����_�5�W��c#Ȍ�ook1�:����֎!��A5�p[�-l��Zf��םR"V�#�ް�Ev�@w��)I���/�;w��߱|L)G���@�q�w�z@��_������4^J����)4V�1S&ɶ�ڂ���n9�N�eP�a�g��"��c5a�_�b1�wi����tn�.&<N �X�시c��	���ɿ��{��ö�F_�:_y`���5�N�p��6���#r=�0�격;�"����L�i �[��x�>oV����Q�"��稳s�^/�ل��Y��O�s�G>�V4\�>y@q��[����~�@pi�W���j�������o��̞\��(���n!��uZAo�2���r|/s��e`C��G��`�!�N�8���H��0.a2��Z�8A�fJ��h� �����h��^�#�ԆxF�j<#�ftC��:-�x81A���e�՚��J<����I��E:�v���I]v��H�\���am����������a1
]��Y^�<k'��ZmmE�����NvPƼ���U�A�G�>^��w1�%h4��b���,��@HɎnt1�?�����#�I�錮^�.o,�`ck��Z~�.�ա�����<Qָyߍ�s��%����dMfF���F�W��� ���OP`��݃rDw�u<)��X���r#-�7���9�:��F*h��> �ݲ�`�#��?uv�l�c�T2�s�ʣ�G\r��g`�P�F+r�b�A��ؤ�n�6��V^ �����0�a2V܀QV��oA.���4������_�;���&+F�ѽC��W�=�`��ʴw��V�}V���s\��z*^x����a�B���o����\[I��jfFp�@�*���w}Q'yz���1����ĒO|��/���M̓`K
�=�(�@��M�ξ�·c�q��B����f4.��q�7V��O�sO1�j�ӧ(yq y����y��e�!��-"!8k3j��m&Q����,�̢S��ځ�c�	?�g�z�K"E$�$�
2x�[�H��Z���������, �"�n�R]犁<�a��ŉ�P��89�/#_Br��P��|֠��hQ<��t|<���5M\�_�EðQ[����e�g��4�lx�W�U�@:P\�8��bWO|:�f����b)�8��*q��䪔�K����Y) ��n[L��c;^���1d�����m3�ZLw��(lj�����S/ �/�����m�"����c�<B�<1 �������p9}O�~�v��O��]��;ڜA�z��#�RH�v���,V_lxa3]_l�}$�0���7��`��6k�7��ұҺ���6��rtC�S2��Q������fḱJ4��ڒ@�SD���	�!�k�Q�x�1`	~۫8��.6uf�������oޮ��ť�x�	3�0�E8���?�"dX)}�d��
����
A��T�&����Q��̾e�b A��^�1�#I~�E���y6������jZPM9o4e��׋ݓ��+�V���"A���fO��ԥ���hmS��+<G�$��A�[�D�*3����Z�pXg�~���;�#��QY� �{�=��񦤍����Ք���
���ꏱ,���@v2�ݬ�������҅m�P��A;z��˵�f��LA�$�Ղ�%�T���,_u�(��\=ƈ �a�I#x
�;��zU~ӎQj�Zo/���B�#�)B�l�(E���3=<1�,m�^LL`|�C(蝩 �(����f���l]ݗ�u��bx$�K"�"�wkFp�0�XD�s"y�i�y]9��<�q\iE?�I�{�-��]5�P� ��������W{��Mb��|U|U�_Q&@r��̉F��X�cG�����9��d%ܭk	���v��4��&����4��/{@�n�1���8�N�JL��t�V��ٷ���#$��������<��_2��g��Bʜl�A���Pr<0�y��x���m�j*/���d/��tS��5�l" (E�����X� �[�:��IjJ_�ƻ�_�`�� q��X�Ka�D@3O�����=g<��*�{R�|�F��F]�o�d��m�Ƞ��Ʃ�u�T>Y�/^�I�f�O�d�v��[tc	�&^�O��-�~�;��|ԫ�����'�հ��Ӣ��Tr�@�"�G�NY"w����G�6a�|�v)F�(���ja�k�-���R��̲L��`�0k��p�vq\���腭_����p�ᨹ�S��:�a���Q���V8,��KTg#�P���IB�۳�kg�,s�֓��jĤ�Ij�;�����n�6a
Qs<u˖q}�&�L4�VeL�=J1�z�ݽF ��$�xM�D���kTF�4p�:~#B#��U��yJ[�rQ��0�6��~���,@եi�q�*8�d����e	�yJ�I���I<�����3LW�un^*Eh��RX\�{�0�oj�	V@˄�2�����|
W���VĢ?�H�����V�!RØ@��D�ή�>3g��˱��Hɕj
Ê����L���hs!��i(/FO�v�����������u`��)ּ���B��b���DWsC��'2;.�%��2����~�~�.�#��Aa��Cf6�G���ԭ�P��5H�m"f����q$��KK�L����6Ԛߦb�E��1 �KR��(�z�=��6�`%_(�ά�s(�	��ڏ�T2��҅�S�.� ��o�Z�iش=>�,��Y!��L$z�c��X%��U �i�ȅ�R
t\�ц�r��YU�YQ�EVV}R��@�<K�ţ����]�m�;t�9��jKoW�AOc�dP<�$�O���'�MI�L�ylP��4¯���`�Y��h���^�O������ �X�u��X��I��Y�⎿e���@��)�'��,3����E��B��3��	�d�d���]�7�
̩?��152�<�?]�ҋ�ӿu����"�)e&�hV��:��9Lu>�*)�+���e�1cܺ��݊���q��m�U����rΤ�>��P������7�tm--	%���9?5��H��I���
�B9b�U{�9��#��è�7�v~¯�����8n�ا��*K�5F_�>FϏ�@���V�o,b�x`Vb�iګz��l�n˼ C_�715!�/9A�&���^-�
����-�v���__����a!~א��y�F��Fgd\&�s #��r�VpV�	�Bpw0�b�\�p��̿8.��ʇ����H�֖֘3��8�=x�v�/E���l�c0{������Zk���H�Ġ�I*� �|0��Ǣb�v��`��Z�W�.�P(L{��bK���LH�_Eŧ�<Ϛi{3���Mg�rdȔ���.U��,})ghԠ���㑵���qK)��1����T��|-���#��,Y�/Ȧ��~4:���%Q�o��g��<Zj@�d��ч����Hh���^'������Ⱦ�[�U�d6-���O�-�N��A��X.�0�ǍvڳaV�m�5㦺��me݁E�]�oc_ֲ�d���(��:x�ś�4UuP��fѣ��6�����D��B�RbD8����T���y��B �{��ůeN\��E�3��'Ѡ�Ё'�n:�?:�X�uO���L1�d��!�t�5�MoU��t�2��󽥘w�֧l����z,NIv�^J=,��D	N)?�Iw��Y�)�#춄U$�s�4�h�e*���H�Ru�K��O}l��BvH�8;����]>:�����g<�c|h0�>���(�$�J�d]���@_���B1�igV�C�)������Z=�]���#�N�_�ȟ^�L	ɐ�d�P��V�a`;[J���̂�\o��g���m(�d��dͫ��0%6��)]�4�"</��	�
P�\���̪����R EM[:�E��!���x)z[����O�j���F^̚�&Y���cC��z�Sc���k�"~}m#��i��z�(�e�O�$�`%"�G�;ۏ�a7R����?)�E=��S��v��Kl�B�10��u�E�+Vj��R�5�daظ�h���K�nq��C�5��$N��,E}�1D36������L�:n[�!,���-���V�紼�e] y"����N��C�v���Kf�X��]��4M'�ʧXl��v:v:6bͮɎr9���\!ί� o��:a�7͞Ĕ�Ҕ�l_�=|.>Z\W[�� B'�a�3VЉ�Ϣ�21/pm�m��f�� 5��M��B^cD�T�/��f����2�0�}��ĘX�jӯ�ܳ�-]~4CN�px��
(����=�x��}�Q�����T�(�B����؝�O��Lh��c�[[?���m���#�����\�:�|�P���; :�>� ���M��~�T=�?�)V͝|��b�
o~�-�S�i�V�>�#��j�8��,�3}3���8��P�$�����"��c�2����ݹ��/�rG#�i�"E�а{_���َ����^-�=&��,h�콡���,P�O�|�4�͘2�8���*�Ԩ)2F�4�B�����(.�d��.�|�װ��J_:�E.2�G� ��Ǌ��*h���\�b<��;���;m�m���%�@��a���Q��M�/c�uL���H�2N��KB"R��@�����k��Gz��7��fO��\
\jp�/'j� =�{�36����Ӣ��8���wK�6��h�R�9���O�N�6�
�n׹[.[��cCU�L��5�E���i�\c	�.טp�E�0���YD�br�3op6˪+g��mjJh[ۥ���SbԠ^�vi/PˊE�����qB��{�,��0�xZc8?��;M�(gS���+�*W��~T�v׭c���"{�K3�7:U)N�fG�A��9���&�U����hO��2-�j��9�kv{�ͤ�O+�)ґ~�]�/y��J�˵��Eh2ص������L�et^<ɢ��a�u�U�h/�B�G�Y�n�`�8���W�_�G�k-�M����E���5�T��>vB�赟F���a�2�e��0�q^'�>�K>E����&��򎤓�ڵ��8vN+1���_:���b��j�cE�h1��E��1�E��V��������(�������yx|W>�t��E)9TT	פ��q�����Ц���xs�������>�֙�uVBi�`�30��a�>}�#w��įb�ܳ�� �~�9L�]A���
���ǒܲ�'_�5��ʬ��O�4���Y���P)e�ջo�8 ��f�>=�zS]�m�|��M�k��6���Y��e�����W,��E��yT�r�?��2	}�s�&=�����yZ���� Ä�]|��GNEe8w噵�):���=.i��Y��&Uҷ�W���IkNB��Iy�~KWx��%��(u$�^�o	�Vq�5�Ɯ���M�>������>g~lx�n5�2sE��g�����/|�f�,���l�L��Ϣ�U,[#�J��i���㯺���*��4JL�=ʒ��=�̒M֗?A�=�z+B�S��ЯX�](r}h�Bά^(�O~zj�iы���˞/И:o8�T���װ܉�����{�8_}���6�$z�L-[?��^{YYM� ���C<6���̶'���HoT�#h��&+{f�P�w_�	�[,�Š+�b�� ����	�ʗ�Y�`�η��$��Nw�	K���)�w�Sh� �m�u# v�DfDV��C$��x E��tō�ქ��ԑ�%R����.��U(�#Y窺�If�H�,��~���&��4�wy��`{'G���n�B�d�Ԥ� �sE�rGF��4�������ܿr�`���?�%�O�x46���_},���3�`܏y��_\��5���8B?@����;4<F�՘����P�i'1�#��V�2����^�/Ԫ���C���������ȇ�G��,�w)\q��?�@E����yeR��u����E�4���*G�R�}���-�Y8V�Q�0���9�U�]�/4y6��5p����n����hQ�'�����pE��*n�z~Y��c`�������
��l��>�����4�_�Xm�����y�Ao$}���)��t
�+ޠ�.' ���"�Z����O�uf�ތJWD#��"s��\�6���~�����-��{
�[�U!��Y5�\�V5�ϥ�����_�H0
�<��h��%�C��d%�S��.�I�R�=�b?�������Z�_a��2`f���P�k���+ ��~N���yl������KL�\D�I;3�����ַ�F�0��į�\J��җ�p��~��X����HJ0(=��p5+6���F א��/*N���=M��-�����'���}��� HƸ܎��B�C�_{X��#��OGj���������M��q�:���gNY��%�k~nY��ɓ�S������y[?�{�׺����QmeW'p* �Z[�����T�'�=�3\��{�DR���>ׅ��2��V�U�q'G�ֲeP��.8S$m��
�C��jk�4�> I$`Ԓ�wo�=�K%�VC��
+���Y���]��W��C����YT�߸ F�C�=�����-=u���R�r�$ ���s�sD�̶�Z�w�����4�׺xl��K�N���"�{Yu8u/�c����"N4%$���XF�+�u��YY�9!�V���r9��\N'�T�ߐ��qY9y�������gӴ̝�/�!�0���S�ɫ�	e�p���3rXNN��3P����=ذ�����~���02g�2X!ևP�2�d�ѣ�;x�3�K���@�U��+x��;����o����K�����У�L�q����Xþ[L �~�@K
g)�9It9��6q��u�Oğ���E���Ch���1=�@������yl1m�H3Z1�+��f�����Ļ�6����)������t-2��s'���h�г�"l�/>[܆
~�Q���\?r��C�)xJ�#�g�o.�!	��x���
��l[��?�K�u{�:���
_2��p:��B�iR�W���_�V���XP^��ږ�Ġ�4Ƹ݆{A}���SI��)��x?���d�ӭ2�zV�ҭ|ٜ*;�Ij��Se�*
�}�)7��?�;�+�ۉۥ"�*��;C� � ��ݤ�k{��]fƑB���n���O��d�տGt�c�KA��]�(�iz�v��P�d=�*����=�}��f-M>��r������-�Z�8p)P��H�-�Xp(M3S��;��3t��3q�t�g��:t>�&��\҉�Hy`��9\Ai��5
����h}:��/[�΃O����!cՄJ;��8�c8=�Ĕa��v�Ph�M��q]o�F�
xEhk6�=-9Hu�,��y�77+���\�m�~h$��5N��\��b�����;k��yd���0D�U$ge\0����`#��&<]r5�}��N�UMb�KZ�!�����3���\�Zקt}�4u�G���W��4��F���P`
�5�Õ�KѐkMU��mL��:�^,�FR��0$`Џ���"�r�ڀ`u�_����I	ӫ�5껡o��@O7d��EPh_�1!�ٛe� ]Z*�&< �������I���k���8c�D�\]M������j����ST��Y�~��E��3t�v��8��TjH�=�-ǚ��t�dv����By�k����S&֝+�
p-��^��Ҷ<	��9�60e�}�LoTu1&e��{�O����0c��!F:T��RZ�#kI�`�I��	��G0V��iضЦ�J�Owy��+���܌Ѡ�n�n��9����ť�O$�'-
i�w��rv�1���Y�B;Ew�{���~5��x���\K̡�x��N�~l��m��#ד�:�8繲�u*�]����5����5_�BٙUì�Ў�޼������1���G]��?D�z�:��N:ac?7��e���%��M�N=Di��L�{kő�������I\N�0seϚ�yнJ�u�i��zKE#�4�oInɫ��=�QH߯Y�f��n�x�~���}�MӿV@#
1�(/�K��ܤ���*Y�Q��V���p����W����>7p��i�u���n)�@m2"1H1_���9v=D]M����[��s펱��H[ћ���N ��Q���{� �TǶ��iz4��nWF���S!���n
����R��Nv�`�p�r�t��s	�����,�|�]�?|�����C�f�H_�2u�9����'j�I��6�@ln���o���G5�7�[�D�� ��<zk����̮<(��n���8�t�r�B�>�8`�_�21�w��	�n;�-�E貍=�$H�B����8pM��
�N���:^N0�"할�?�(u�.Z�H��oJ�4�������_&�����=�8�N�^��M���%^W &C赪��>�=R��xAl0��=���(?��|o�'�u��QZ`iDPB׻�_4��5��ˈ�ߙw7`�!],袱�_�E� ҥ�MU3R�i�˶���~�A�h%�oE��f6�-�lDN0%��cc!Y�r�J�m�&��$mY~�l�䍝J`���E@K-u�FA�|˄��wf=��*����������FbvK��96&�J��N��n��������3o��^�O/� E�j���g�&��	-n�9�m�����է���I-��wȴ���_��J��ͧS����˝msp=�%IytН��ɐ�2�4V��d2��n�ʔ���\��w:�c��l/ԦV�W�#ߕ���T���7���9"�7��Cc�J�\��6^n�0>�s�)ZS�����~��>Ra�؊pg�
�oi�����S�����dr��kH��D���;����YIc1=h��v�긅-M]��	�Lyg���= �b��o	lpf���U5Ο�Rr!GGJ��KV��*���(�%@>�Z��������toǋ�/P\����.���Ð�~O3,L��!}P z�'�����2���>R����R�\^��/�]�������K.@�=� ��oСޥ7O�v;���Z��_KN8�'�ݼu_�X	E�y�>:|S��f=���.�������m��]����Kd�N�5�ɺ����l.��v���i�߻B	�#����#m/a�lp��G�D(�ܕC������p�� �X�,���X�~��w��c<�$���?E���-�c!7��j�;��=����}t���� Ѓ	�&��#d����~=oL��6��	1�1=��sSY���N�o���=�*�vl��b��#������[���-��2a�3 ��e��¾����1��!������Qe�ds/-��΋�YJxc[u��W[�g(�oT!"{���i�&O,��kYmm:͹|F]�pn������E�Ȋ���g��A��z���>,��lW��t*��֛��a�����,Yi̢�	!޷Q����
�e���O'#H��yy��O��U��7-���5�G�Ρ�8�2��Vg�(j�Q�Z�d���k���˭����5d:�?����h�U�T�>�{�8@B��O�E���U�l��� q�����\!7�da.����Ս������H v�Q(Ъ�Ar�����q����Қ1��Q�X
Z�_xf
߶�o}�ѥ���&�t`��!����9ݗ�[��R%w#KJ{'���&d>nl��]�c����چ�n�V�mbTg�к���'*��Ķ8!���s��2yG� $,���yp:}�����ޯ���� �ņm����ـ�%?1�h�RY���7�����LP�U��QA�{G�n�v����v��C3�;}�a�q���������sVN�9�2��#��+�H��A��r��z���Bzgs��
QY1�l�1������(��:ED.p�s�^���n���㳧ֈ&�Y�{��c
5\Z���-�uAΉ��z� V����]�K����l�y���[M�2]��|0�
����4����mu�5��Tf���*�[ۈ �e���I�gٰbS�na�m���E��''�9Ct�Y^������G����c:۸�1N�k���\7�Էҷ�QP������4r�S?�nz�?a��P��&��������ۺ�C�*��3m[�Ih%J
:�`Q f��*��d��Z�X'XS#8ŕ�� ��� ݱ[ԥ�B�0���E0�3�r�"I���+9[�s�hV�Qr	���	���{i��ي�b���b��r��g��+��kǔl$�����,�&޶�ĳi骶�Ϳf�QE��3{�S��c��|�YѲ���ae�'l^Ȼa����s�'��{|8���.��1�[��u��t4�M�n�pXa]Q�ݹ�1���R|�Pi��Z5��"E"
�'�c����%z�s��iK4q1��|��4�n�itMߚ~�brX�m�:��s�čx1�qH��l,k��#�u"��Stj����MS6�^q{Y�ߜ>8�V�-'�Eԅ�#�& O'(]�u��S|���W�#7-�p �_	��k�&�Un�ۍ��y⎋�Qy�ܟ�o�����<#�7�?e�����FO=^�"<T��`�d=��7̀��N/*�f?k�Pq�Ԏ
Mh�Jp ﳼ�R���{��xh���/��:��bu1{�NDu]o�6�\r�W�V���F1a1�%M=t%��G�'�,����Zb��FX@Q��	�����1xE������qn-�a��Ui�D�	�X~�@H,����%(<��܏܎Wk��gK���s="r�M���<�/*(�b��FZ�L�S?$�!���wiБ��� UJ&y������MXWi/��m�^�qr�R��@Ԑ�n��1[�+O��lӎU�@m`�t6�Yq��q���Q�Ǩ��_jxKĚ���ŋ4������N�5�)�p�bt��Z�B4�ϬL�iq�u�;z#RĞ�Q"D�΅a����0Z���k���d�oJ�ncpmC��������z@�C�[�d�)��|����p���K{�h����F���P�{�l����l:��WC�Ql_)��$��@���0��^^7��T�zW��=H#["��c̩�i-Z*|�`E'����-;��ey��gI:��B�)L�DJ�)ٲ�n�@����C�,M+1��V�@��f�Ϧ5DW�dy<�T��Rc!��c�I�gS�p1�-�����$��vT�$�v6(>ݙ�2�n���-$��zGkD�t|�금Uq���|��"�O=�oK!��:sl��54��L܅��p�"
�t�M�N6���0�)ь-����-R��jQ������p���!�YS#�	���x���9�b\{�H�+��������O%�r9c��7mU)��Ԇ�r�:��~�L $ꫬ6�A�~?̪b�p���(���2���}~MyT����Zm]�Y����SV��~~�m��a�j��|E)WF����3rZ}�@4�d8�����ܮ�3�� }	
��?-@�+�IB����JY�	���D��9"f4��B͵Q8�p�(W�g�ܶ\K8����$(-*p.�߼l�j#܊8�Y��'a֟)#�@�Zcraȥ3A��͋��nl�׸��@+1��ɃD�n�[s3��oR�Yu�A���^�ޝ��^`֟u�>���z� ���%�b����#V�@��Ľ�Mu�?
#�+-����@�C��2VBq8��'�>�4�b$�0	۔읩nZ��[�0?��&h�ݯ�H��=$>�_��5�)�W=�lF#�;����K�� ���z|	��$<9Kb:��pp<̫y�N�<{փDT���D���2k���e���ŮR�"�oV�|�VXt1�#�P)�Wx���Qs4a�f*adG�Z�hTXe=jQ߮&iI�F#9��)���|0��=�7pg��7ݦ�N�Tb�|�1���"�����$t�������?����	{8�}8�>�{�~��_���)x��|J ���e\8x�C�V�%�6���U�$��K,R)��@Kr�bt��u�M��A�ej'�DD{=�Ж�#�n���4HV�&w��T���]Q��L�����p���k�T��c�msO��~zM�_�Jƍ�v�G�%�~t��<{~�}G)u9�'?s�0QQ.�Yi�rj ���C;��kr(�~X�"�� E2'7�M-��ɅRMo�&Хߢ�� Z��W�����i7��6�2�z�'7>ʠN1/֣�P�<�p��Ɵ��V�Y�kt���C��� �4[0jty�ϴ�	�^ܰ)eQCYf}"��B/,ts*$��������#?�7����}�G����4�w:�.�r�T��{V??g���Yr,P4�c�ff-���k���so���&�Q�7�B�>����� FI���S�)k2땰�O�������{���?j�p\i7��n�M4��U,/�)�O�9?���A�j�o�puMڊՉ�AR�ss�(�5��������E�:ΨJ���"	0��m���iDyՏ%c�� ̻%s�y�$9V�����3T!.W�����v8�aɵ�U@�P{6�e+�)��X�����o��a��V$�f�������u�9�=���$�����2�&|{��Q,n˂AĄ{A�
/�Z�|�u��"$d��j'Fn�/ �h�C�F�ew�o��{_Eм&��_XU���)��z�/#X�!�I�m�-k�����.i�l"�ɴK~��z��M��PpZ}�gG~�B�y���5���\�-��iYB�ׂ�+���kQ,�1�1��Տ<��W�-�uVMC�� Q�,����~�ip����A�T����W�y��3����?���&�M'Q�Qp4�.ߔ�W&;��sa���1{��֑֏�C! ������Kx�R�jc �٢���y�>p�m��Ǳ���l��ٛS� 9�r��BE��#��:�*>P{e@�0��lX�kl�;��)�е�۹��vh,�����<�WK�2����eоU�����f�֌#���U͈^4�\dP�B2p��+�j0qN޳?Ք^�o��b������&d��a�1��r�ăC7��zm��ԩ�Q,9l����f�kxhjS�2�HD����k�|�g�� ��RY'WFv0���[2lŽE��b��'���_qq���E�7�%���d"���Q�p`LQ�e�w$�Z�g$�C��~A�a�ISe���<�RV�zUk�a(��3o��J���V�yb��ٖ�59䳐�E�.��y�0q�����(�W���`/�]�@N���D9E:�GT��v�8��$Ϛ���o  �w�i��(g#F��F��ņI,5޷4�|gFTQv|�L���vr���ղ�d� �W\��?BG��иi����6
�b(�R������I`�WQ�2C���d@N��FBr#(��<�+�� ��'  `�=�W���@8[��]2�~� �;!Θ���^��D�g=^��v��B�vƷ�	ȳ���]*ۻ�e���C�ϟ��V��h�y�Z5������V'�<F����
�~��W�#R�*5�B���٥�����b��͒cUu��gC�9����LL@fYP��!�¡Q�3�Z)T2����������ԱPm.��yF��;Y'/GT*��s�>��8e_&�������)l� ��KU2	�Y���;�b�f-O��J��N����P��~�	�Pn�i.��R$]<5����m��nB����=��������J��ƹ����#��88}�e}h����ct��>M�O�Z��6bȿ�l�R���eB:4�@5��K��+�\|���.+T��o�	i��rNRqA��4�˴�����������⬨>S3I�UK�!���`�a��	66OS;�+HOa���\�=��y��D�	
o�AF�����yM"V�˄!c<���q�:.��g7��uu̍��f����g�Qy-r�%��VM,��h[<Zi6��y���
�X΅h7���@n2�#�J���R�nY�c���MHA�L���~o��>����{�Ff&��*hS	�]���a�ݣ�c_cje+y�Qh*��jL��z>,����r��S޺�b�B�*����"ZL2�ʁ��ŋ�Z��jJ���V���4f@�և��*M�{_3AH���6s�"̽?h\H�ܞkjԓ�0��vV��Qf!��xȓ	q��k�\ *�@f7^Ⱥ"!u���&���A��1���xGY��0h��U���p�L�M�j�'H�{��6�j�&T�	��t���˟t���!�,	������W>�W�1�����K][{�o�N!6҈�sT'��Q.U��b�1޶�׉�t	��n�E�TE�td���ݐ�*�~��I��#�`H�ڍNT��GN�Hoj�~��F3	K|�E��ň�1R2s���~_���v1�C��'!�7��#B�xh�a\�E�˙�w�^�0���J1	I����ʦ���O����7(dR���o��$h��R�\w�x���O�'�8;�Iy��Z�[q�����a��v��0o�pb.q���{9ۅY�ř�s�zB���a(\�S��|*�E�Q(Ŋ�%���%c|�֕�e ����"�:}���=�Q�@
��(������5iwm��b��Z��}�J���c�����SB+��iע�j2*;Q���������iHo�KĲ�x^��?3}I��Z�K�:�S�>0��k�Q�����SH�F�m�8����mN���S荣Bu��B��Π���-�^0zfB�(tP�q�rdS#6�lU�I>ׁ\���kw��`rge�0�i�sN:a�D�^>��;j��C��\
�e\�=���=���.:��C�`RV��6���wl�0� �d9,�>�����T*5��p��������,�v
�������R/,���=�6����c+���p�ns���*��t��n9گ�[�{�C�I.T �@��3��̌�lvG�����a�tY9&��D�)���rp�k5�٫ĥ��0C���TC����e�;"I�|��i�b�RKR������[���W'9Ȼ�r�$T!6�Co�R�:��S����,�=U�ۜ�;�fUlχM��iK0�ˮ�^L���ŗ`��T ���G��(f�ȿ�'��;�e6�Y�l�N�~_%�a!�9�+|�JXA~��4��-����'۠%wc��o�B����R����rq^m�m+�~�HZ�'*��^���e�1:^L�>1$a��	���4�� ���|�W˔�9����o��|�I�=��>����K]��r}��T�Kh �xNuo�$�yx��ጋ8�G.�(Z�;���W�B�G�����y+m
��%h	z�f=/��h�G���/��S��S8��Y�>���3i��Jam����{}���ґ��tkg�%MJ��Y������� ���d��Q�{C�����B4��c�	λ����>���<��Y=�}�EA:H�gmޯ
���¢�I���#s��3��K�ⷙ\��IZQ���]�H�f���L5fE:�	V��+�q�ð�3E�j��XѬ=�A)~i'|,ԺZ=��ǩ�Z-�+�����QB9�|&��D���4*��Nr%�Ц*@`�o{H�<ّtް j�i'g�_���0�]l��Մ�w*�)��?��s;Ϊ����R�]%�:��Gj��ю�x�V^d��\��J|�g�|=d ir�����x�)���.���S���k�4�mOq�>��P��ٗ@D���PHf��~xX��|�M�؂���)�F���D�I��X���tE�E��&(�;�r)O�H���:)l�IC�?��O��ۍ�u1�b��Y�h��ᐭ,Vܦ�C���]S���6��쫙v�!��GH����������w���]yl�㮝�Z8U���ܚ�5?�Xx�]ڡz���KI�C�O �e�q�q�iɈ��&Y>w=P���<UŹ�i8ы=�OSϕ���4����1�=Ė5lng�
��'���u?٨v�.�#������eS1Ny�wi�[O̙���c'.��߃��B��*�����8�Fx��J�G5h�n�ꕇ�Ze��ă}��İwl]�EJR�f��\]�q	ڠ���~}p�+Bw����w'e����zٰP��Kݗv�63���L�Hצ���+˻v����1������)M�w��ݍZ�iQ]��*�4��p�]	�YIm,օ(÷����f�@cƸ���8 #�\6ONNZ�L��4&#Y���+f��x���jrl�v�+��jgl������.�W��2�o|�p�@*�1&�y��z{
�F.��\kB�s%+�Fi�M^��s�`�����Őte{:q0��F<��7:�_����R�E��Y-ʁN/��M:�4�np����C� ��"	xmg.�#�/ӱ����T�����|a�-ur6��/(�����8J�jo��4a��ހJ(&kB���Uu�f���Bg����bτ�R�f�NڞEV�It>����㵙<�%Z��X��>;*5����I������,#~�D�$�J��4��m��4�C���|W���i_`2�i6 V��3>3��z���5��LB��}�G.�g{iW�WO��T�KAE�~+��v/)gY�M�z)�#Z��͝�=e�d
q�cÁ�W'������8��jg�.T�0��U�~Bo�@U��w��k�? q#�		ȼ��$/�ק��m9��)�o�ID%��H6�CJ���`>���M�b��>fU��d��:��po�0P���M*�(�&��'��^w�_S%�� C�Q7����.(| g��I�;�4Ϋ	?,�<���	p�yѣ��.E���������m��Q%jPF��1�&]��aۭ��y�!-r�����C�蘀��!���a�ۘ���E�����6+�����Ͱ������.z���`�Ny9�x�.q^|�W����e%23ޞƻ_�t-��~ .�q��'�3(`$S��G��4�I��{Լ��cY��Q�ZM�^G�)|�AH�{Rn��@[k�j�H]]����Ǜ��5�B���=!�S���!_��`����?^-e;t���0����Ǯ�H��g��^_T�[.o��L4#d�w�l���� &,�0�B�ŧ�W�Lǎ��-�����'W��p\����{�����|o���3�
�`�V^<�ϗ8c���3���k�B4��0$39���[n��<#Ӹ�k	�bEaR�N~���A�ϷQ�r��9��D]P�b(Q��,��*12�E�Ǿ� l"�*x�Z���+��H�t����|ZFvϜ�������P�m	�L�9�J�%��G2� ���7��e�X����A:$u��Cy�G���N�i{x��+���M,�W�T=q�9u/6�̛�������m���x��i��s����v�}Mc����	���pn�f=G�l��t�uE��gs�D��>�SI�M�>s��_� ���cb�`;��s˻��Zu[i�=��sfHu���~<ɘb$�WO�Z�i@�5�{{�s+���#�z����=���!�a���!ۥ�e�J�;������1vϝ�4�|c'\v��h��϶n�u�ʚ�X�O�!�л���G���ł���l �C�XA�"��O9h�8e��߄�V�r\���&ߜ��h�~�< X�b���rć����v���ߑ�=�%�����?����7�t=�m�*���O��Q��񞿠/��}��1�<�P@@��1�Z�jN�|���	Uþ�\�n���w#l��ތ�dY�dSr�ۂ�=J�$5K���;#���HeM��'��j�������R�J��8����0ܱ2�@hFD�� >���2}�0������Y����!/��_���?���0�Ò��ʛ^թ���bQySGG6{�'���=�mnU��zF���'��L�l%�/]ʞKq��U���so�`�*����0ԏc��H�j����V�:��Jb��u$-Aho���/���֠9�D���q+|�Z��`�g[|*�m��^�Q��*�±n�Ѫ�� �d_��k���wmS�u�QÐ�AX9Jp{��s�����ꚡ�x
+&���X���u`ǒO�yS�88��61��"�'�2��)�Wx�^���[�v!*C*l3�#)�����NN!����fc���-�_ъ�T
4)�c-D��.2��=1�ϧ.�HZ�xLE��l
�07�K�:`��Wd�~9"ۜ6���LY�<��h�C�n��xC�z�w���T�� l�BSr\CV2f��8�qN~�SH�B��9"�+H�# <6;�D�������tɰ������d���bx?�͎�nj�����j���^���$�������'jiNϙ{�t���GYS~�}5ͲEq�8]�ľ��If<#��d��߱U�o�1Q��֡��1���n������0���OQ�ٲ��U�|M"�IdaѶ�yo4���n�s�z���>f!��?��~�y�Ԯ���~�i=G���J#���ɿĄhqEas��j��:6YFy�92'�"�J�O�@E�����NU���|л���-���:e�\�S���suF2��ipI���3�����:�H����:�b�����u[_���t�������*T�٬���/ j�[��k�+!���* �V�t�'
�������l���gZf����$I��m̓%����Q�����D;ҕkv�1����3�q_� �LX���1^N�	Tnّ4c3]��a-�񿭡t�L�=#�{F��M� I70�7���By��RRW�J`�D�o����<���?_M�s�߅^L��5�f/�
��B���hM�AҖr��'�1�x@�x ��]gu\�[�1X�U�?2�p��4�@���>�cH��#��c��У��|���g��cչ7�D� �F�͋����ì6~'���>���k����F��F���űІc�aV����	:Q�$�6���+�Y��ԋ�'V�3㋧4(^�m��"`�c����@h���	�1�["�?/���elxg�����B������,��X$�^�B4I�M��;���cH�&i�����N!�3��y�e�PS��@���Wd�CM����%�����:�A*[�N{��U�ͳ=ٳ�:,�x�����dKٍ�w�֖�����7���1��צ{D,p���ݶ�zL��d��$��+���0�	6�iC��Jr��HJyd|N~�x��}+�1i���!@NƧ��ۿ�Vގ@o,.H�s�w	Ų����֐�PBA|�4�e4.�������:͆Ow䐍
���J�N�G99�s�)s�ܧ($/\20�8�t};�Q=yf�}?2c�����(�Xe���_B�4�N��XK:C�e$:�f7ח+o?��qx������W���� �E[��D�-ݹ�c]��Rџbx�;�ܱH�M�pm��O��v�&�|H5ʞ������@7:��e��aCo������J�s%��Ŏ7��p8�$:��+�4cJ
��-kh�tG����'9b����\���������
�rZ݅�9�.�l�7��4��B��$-D��gj�4iょ+<7�9�A&�w��A�Vd��X5 l�/ʟI�_�y^�[��`�FP����:�_�C&ۙ��4{
[����&P����K;Q��ȵE�6�|Ja��ܠG�}Q N?�����m$� �imr&�݃ZpL�o�� �n��~O�"� WKJ��jD�Ȟʍ�����H�7L� �e�߽<��v�����m�F�~���!�݄�H��\�	CɅyzY�ŐHI�B;�Α��^{�6�X��JL;��FX@4]҆gPȜ/J"VQcbТ�ưw�'~\���t�e�B�����SV6����W��}m�ݤ+�]�x��M̨�lm^2hcIgY���L�>��?��?�΁�ފr��	=�N;��	�-�˜�c����u��96|�Z g�؍Ij9ʌ���29�I�0Ñ������3}K��w�h��f4�^����Yx#6��9T�c�4�����T�0�����b�p�O}0�',�]a��$��?����&���d� ��W��,5Ww9��}�$�X��\E��0�Y�6~���#7���a�$�g`e%Q�z�_A����. ���n}��va�!�T��]+��a�7�O8��0��������סYV�P�$OQy�Hq?(��"g���#M�������#��ma|��G�VR�K�쐖����kخ�28���SE�6o��3�.�q"����Q J���N�J�
�W <V�O�}���SIfD��o��_�B��t��q2�ś������N��)R�ZX˟��io��7�������6-ʎ���#�	�:�`�L��z�Ċ���]�M�D�3k����2H�:�z��&~���6^r�^a����`ä�ܑ�W���x�d����s�Q�y�9�L��z�zJ��i�K�6��O��Y	&�7
�p�"��Do.�c�,��ȻG�@ҏ$�N��v�2���l����)�\��:�O�l�n�=ј�(8��\���>X��?�0cQ��َ�)�׺�i��5J�|"���ei7T7<Ùk�Io����
��H�	���k!h�|�L���#�?r8���#�\�Gi=0xat�	��Yl'��^�1�2�*&Ѳ��a�"$+q�h��L�v����H��8޷+�˶��{g�]J�����o�Dt_�?ɂ���䋒6��;_�9 ~t!`I�mR����9P��X�O
&]Gn�~�	l�{�M�H�31�ފ�7�q���ߵB����ƙQ'?���(�v�����V �P�"��uQ�,Y�WivFM,e )���&6@��[ h6|�&U� �49d�7x�^�[�r���Y��A<s��G��,CC��k�Bb�E�{��*�W����.��8���}�f�B?���K�Z�"�^���*uR,�Tv��ń���zLO��m�K��!X��3�����%�A������?�S��^*��>��H6�� iV�0+�:�T>�b�]��&�n�shyx��z��o����<�Vᒘ-a������&EH�ޏv�bŖ�Pj�����Y�v�vl@.�0,�MF�=��oG&!,<���Te�;�����a�LĜϪ�M6p��R
NѐRڟ���%��e�S<&5!X������r-����k��q�!�aJJJ����.:�[rb�Y g����N��=�� K�Y�ۍL+}9��d���;uO����pꔫi;�v�o<�՗��r5�2�c�t�$�v��9!뀋�#V^CC�j�g�TA��`8�G����ñ���p�w;��,�,M�Q�H�,�Ʌ�'�N0+�)������������q���wN��rk�S��#܊�]$�?E��EA�i�aF�I��+-6��+D�M2+d^�wP�/��RKM��µrבը_���TE#���@������{;S�A�/x�;����z��� �����!K�ܾ�2<���e`����d�l�2�x�L�c���P�ݶ��)��Z{˜We��)p�X~!��������;��<���#�\CH��g4��M��?��ZW�8�$������,ܤMs�wԝA��eֻ��8��489��߷��І�I��L�eP��� ����:�ZHo��A�Z��-�Ca�C��\����W�ӡ����Ɏ��̌�(zO�Z?�?Iv��ͫ�XMź!d�d�Ƭ�{~3�4a�Mf6�Y���F���c֏[M���\�I�J_ۜ�a�A�į�RA�<�"�ֆM���ς�Y�iW���E�$Kt���P����A�rt��^��+�"�q�%���>�2�$|[+i������d�-m������I�p���?mn0<������{ds<��VeOd{8b�#��y��*>�B��7�C���?0�Iz~�~F`"�i;W��9#�u�'�R��]8�� �^6Q�V�%dp[X��;����)�~��c-�}�n:棂� �e�_�>�NN�L�60褐)D~y�8u�2@Z�>�:���ׯ>��D6��m���?cP:/���;��1Q/y��v�#�hk�����>�J΃7:�薎�a�����_�E�M�[����^��.Q�ˈ&+���A�ע��'&n�΍���*�#y����ŏes�ς�t��a_D�X�CwPo��t���ĝv�x=�MXC�\�U�E���C#��Q�Id�������N��˴�+d�<wN���a���9"S�m��$u��sZI�R�/�����E����8��-�r�x&	�f����]��*�߂�@�܏�WL���H�5}�c������w��@��-�/ ]�uHajF�TF���(��>0��4�1x~uCl#x���y�H���w�W&	w�u��|gn��% ��HhyY���Ι)p,{��`(8�^Ў:�xX��p��!�g�؉��aN\���	�'RG�~*]RA'\�h�DD@�<�۠yw�r[r�Yj_����B?g��j ���A�,��	F����s���]�؇�"�&@�o&FF\V�D`�P���J�����<�~b�l�S�E�������
����S�0e\ψ|�!Cؿ<J2�bL��^d��Iy�c�tB.�2>n�>�t˿ߖ��f�������>B��V�&@�<^�Y��9Y7�6��,��@��U�l�K��M�Nӷ���!IsCF�� �!@�Q�Q�No]���{�Ɯ������]� )�kI~ı[H��ѡkW��1:�3��+�|�iC�/��m vF�r��� ���f=g��n��ih`kw0H,-�8�s[��B�����TCڛ�C06vX�(���%�"G�@���2��d�w���¸�L���j�a���i�R�!;2��X�*f#at���|���"�)�w�_���)^i�EqU�*��V�Y���
�m��3
��K�p^�b��TXV�u�x�)e��}y����1��!o�t����T�k��ǘ��ɋOe�p �p���v3�a����!v�x���|ܪG9
2�"�j�O��m+�e����̰1�&�+�Ա�ck�}F�����mm���~
�#UE��#{�(nI�oH�������d�g �H���U1��!�0t�]��@���u�Fq��{;��dݓ�d	.kbk�$ǘ�@"����k������}��f8N����S��j�h��̈́�$%�jf����2`X8�+�e����u�=�"�y�#	s���f�f��j&�ZP�W"wjC� ��8��foe+e�����"�+l;w��֯��ك�����y�2��J4��A�Q�d�=Vâ56�f	���$])�r��i4
k4}��~�~O���g��(��c�w!�^��x�Eq��aR/�P�J�دC9�����-���vּ+��#��@zmy7�����_�����Qd�~�>;-M�S�nDPs�m����)�Jk��������m���X��ݡ/��f����/!MhgP��
���ރ��?��+�zH����&s}-�����P���x�W�L���Z� LZ��+����I����x�y��k�[�Ic�<=�Y�+/�d�L�^�3J	���^z�*Ͼ[��$ޅ!�y�H�+\:e�C��U�y�o��i���g���O5�0���Sx��h�Zq݄���X�n�A���:9����t}$&Y�0"�Hj�:�Y���~4�*�{
i��/Oc��4�D�"�D(�c�oX��zd��-�q8:D��Gٻ��*���UDjs�E"��]�����a�z�i�����7��؝�v�ēE2�r�x��M'��j�1�W���u`ӯ����H����3�]6�{+���W���7@]��x#[��+�k���@LA,����l6���J��=(����6PO��=̄k6��~�VX 
����0A���iP
c1�jl�*J)������o7��o���E���up��Ez���祲�Ȑ�2s��&�P���!��^4��� ��sގd�[���F��&�d�Z����J.F�U�Ӏm��֤���B�DWJ����끎%��ڸ�;$8]6���]��ϩ/�>*�5j3�ܘ��:�ZԞ�ȀS�a�
m82,;��;&����h,�Ɯ;����#T�����S0{zw�8��j��f
=��q �P|&�5�x�ү�KwǸ*>�{�GV��
���qVp�?��5�-�Qh���XK�{�r�'k� djm}�-!1������#߷�0�r�[��zrx�f@�9U���Rl-���j�)�����U���������2!P��/l��q��;(�H�E�/Od��
��OFT�i�qM�NE �zު�΄��pG��n�X��R9�F\�9n�"Ǻ@]*&L�SS`��P%ir����r���~n��-]�B 4�0��	~T$߽��m�Dg���;�h���88%R@`k��:b-JK����C[x��ƾqdT�5�����|M�7�D�����	|�Ty�Jgr,�2Pp]<���u���E�����Fj౧��z���7�W����-;��r[4q�3�M�[�^,=x6�i��ӹ-��x�:�y?�B��ڳ�<ȏ���]��?���#W(>�N�i�/Ŋ��Ή˼����7����24vo�Z���^��ض��QfI�ĳE,[�̴8O��F{����oAf1XS�G��������{���F�O蒟�&��W]��i]�@J�X;�G_���Ь���*V��c����R���v%FvX!����ΜQ����d�;se�Տ&3�VZ�aɉ���DS�fM��c-S���}������UϵB���	R_�䪾���KUft�C�����Ҥ��J�ܪ�̼w9��D�ڐu>�AE�C;5̘j�pK�!�ϭq�f�U�4q��kۗ��xK��w�
�_jkΚ|0�Oj^�*�v�7��q��+�Nb�����W�0{��U��=7�M�kw hL4����ׁ��Z��`nn0�g�K~=V�d^`GY�ג�Jw�ʯk0��傌��4�PF�-n�����&=������x��;R�#��8�2^����%� <iq�>
b�ٌ[��ߍ��[So��*��$�"�>�8��b[_�K�T�02W�D `Q)5&2�Dw������G��z��<Έ�l�rZ"ݢ���Ozۣ�}� �����L��ɁC� S"���
��τOi�bZ��y��&�Ө�gS��D���h3�b�"6Nˋ�L��8b�O$��{a�Lͮ��Og�1�V��E��w���"T����WA3���e�h��R5�PE��T@���o30���{���\��݄�K`{�Q��>8ѳ�v�H���*=[Xܕ��GIĸc|Z����z�x%s
a�Pd�:�b|�/����Q��µ�i� M� �q��:6��<;�ASŦdƽ�|:j�P/q�K�!��F�\����X4[���`������oV�<Ԉ �a~o��Gī�_��ʲ3��p��杲��L@z�$��ؔ�jz�Ř�fu���zy�C��F�v8�x�L���>;��*�r�VE+�·N�����.[��R0�'���f�u+��#�

7�A�,jkG<��W} ���;Ӽ��C�u
���s�vӎjx�^��J����z��2�����A��	� �"��>�6����`��ḷ����5	]J=�2�2b��P`_�'�{,_{� %�?�����+f���$���TK2Y��]JQ/:���| #��n�snJ K�s����p�}'��T�m^.�T?�6���Y U�/��.K"崁�{������}�8�0WM���#9��r�V��C���5�f��/���zj�Õc`��8���m���8��d�E�/�t�*������=���:C&y���SD���\�$�$�������
��㜦�R��·�VHrQ���\W02 x�&Dc��2�8�mu�5,~�6�j|k����zި���l�z������O]l����rqV�N~KY���2�-�Q��$]��2b�i)K���RTl0I�zTA4(�(k�n���mX��9���������k�� �&d�^ �e��g�"�M�����SO�:;��E߬*��ô_��=��������<<�@����(3�"��=�o�SĎ��E�,�V��;�@�=��er7p��ΰ��^M���|峡gyN�^,y��|���yd	���;.�^��d᧪N�}:�;pp�_��}Y��a�R���՟ٚLn�s��.&�n�,���q|�
M6�Y5xR��U�@��4o=UU��jWv[c��a#�}����P��Z&nTK0bC�N��v�SVS�a��L��r��yo��J����p�1�Q-�9W��9\/T�[�x�!ҾN r���䷼Q���mU�yud�u�E4堛}6�v�|ꥮF������y�#y+ֿ�����ض�,p߼�!QM,	��8K���ǒ�sh�Q<$�W>2׶�&����1�� _ŋvG����b���j:��5��RNQT�MCӭ�Ur�Dښy��������t�o�Be�� H"�˞���%��4ő �ɖ4���i��:h��H�&�	���)��{��S̞����?�����lݑ��5��R|��v�ǻ���;��4*o�r?8W�� �"	D�~W-X������5�Gv&�J��9e�>1W�lYn/��x�G��U����l�w�h&�a��%�Z���(���6�sݼP$$ۘ��^K���=&�q�iJD�uZ�o�#䪻VՌ�r�ƴF
2�L�T�F�ڏ�eVϨ�nڌ���s���C�����9<i�Y��" ���l 
��Y�WIl�%B��Li5p�n�@��Cx�.����o�@s�_#�{�Va�my����{�M���6 Lʆ��Ye�`��0�H]Ǝ+HHP��K���GS��Y�s�ܝ�Pjf�Q$�o��F����*<��<f(���Y  �J��<ac}b
ݻ�kC`��4ġ�^��\ ~+�&a�NmՍܨ�?�	L�IC�D�cO}����P�1`�E\���p�
K5�C�����RB"-Wګa2KL$�^�2�𦼄�y�RN E
�9���X�" bB������K����Ud�_�q�}�ND"�{�¶�����p���S=Y�{m�����8�����;P[�Ƭ�S���1<~��(����4i��������╔�`,�5���k�
��rHQSDKQZD�L=L�|�;0� ���r��[�y%B��a�3Qd$U߱��s2�*���4z��fF�z9b�.�T-K;�Q.��U_ -`�^'�����]�A���`��f��;-�u2}< �ёTj}3~/����튿+����R��6S�I#+��r��ua�omge8M}1��G��l�ӻ�� |��V�b��D.���X�e�蒐���-Mi�k�'�{�؈	�D�c̏"	r��"�:�Gf��>K�
�	{t�2���,�=���E��0�-�J�c}��t�_?�4o{���q�9����rw����[�On�c�O���5��j�!�����}Y�A��M[Z�T��L�}��G�x*�� �8D&�C���Z�����*����a���>=2�]�m�O-��Xiڥ���,}|�0B&����ˇO���N���1̓O����h���`v"��U�S4�p��
#BBg$8<�ەӄAg��I�1P�O��a��h�r�=/zH�(�:EG��.���KB�M��;�O����V^;��\l�d3�������)�غ^�J��~�/r���K�6�4�R�u��<�i䵌P��̒� �U��o�A��0$����Y55jU� b$��v; ��1��K,��(!gV�K�JL0.z9��Kh�f�i;����XR{�hlv�m�#����zy�(ܞ?Om�]7��g�M�OJ�SG#j����إ�`|7�������s9N���x�����a��E�C�,̡,��r-H�رH�#J#ⓔ{cbΧ��8S$I�s��\o�k��6��I�e�e�'y�s��a�,�>_�JB���egR?3��X�b�2��l�
�[m�t���i�_�?�G�d��W��]�NYhrH&^/�(W��Ž�����L�r�_�\�	��Y�;��f���wm�'o�'ww�k��XSi4"��e��(���Uđ��豆 |�Q�/�'_y��+�hN|.l�!n��e��"��s3��ʥ�|&���
VW���w�K��5(8�2Z4<���(�u'���o�w���"�3f;`�eU��G�ɫ��Y۳�'�����粠`0&h��n"E�0V0�_,S��e��,M�����	�Mx�J�<|�f�W�i4�1H:��1��>sX��	���:
��[��y{��o.�����x�e����S���ƺ�n���c.�o_�g���9dì�.v�E$Lͩ;"q�); ��z,��2��`;�������Ne�Ƥ��oƓ`]��x�A�٨�	N+(.Y|�����A��$�V?R�}�q[�j�{� t��kx�B�n���*P ӫֆn\�"N.lɡm �yd�p&�����.���r��F����BF�_�%{KQ�UF5��k�Q�_G�n�ɉk�� F!�$�=Q�C (�D�p�}��^�ѽB��̡�ڔ��aAh �	_k�)8[��f
�����D�+��LiOK��tF�)W3"5��/���M����=�7Њ��e`��1_&٥:���_�o��*I��z�B�9l#�1��Yk����+І�݈��j��eo���\Q6�)���ɛ-�gv�\�S$��(�@9}ү(������˻���x0���@��|Ћ�F]N��l�M5d�����K�Mh��;�u�ys�sx���H��3.z���$P��;N��ҏXFw�"�#Dr}px�ߦ�䉎H6�r��8��e��h�#�P�F¢ᜇ0*�RI�%����1X��J"�$
6���!�>o_�.<���td�&���'� .�l��	F���7��o 5$�V.�Dw�xA��d��N�LNK2��,�_�- ]���V/�A��;"(w�*oQe�8�m<�M�Ef�	�`��ʼ��Bd.���Y��Ҡ�A��ks
�'���i7�dl�?��u���i�3L˃��Ʌ7�a�:M�A�c�����^�I�'��v2�ɝOc�����
-����#�pd�#jM�C��(&�7�M[���C���PѼGT�����M���6�ߓ~7Ss��S�	��IU?荱M	U�z5��%P8�����6�
�X;�jYة��cx�6(�ok��I	Jg����s�(0;-���&����pty0���L	�#ĺ�#�c*�r� �����2V�&Bg�R��]9�{��)g����Ã�'XJ�G�I>�D~�V¬�>V�@-�)e�hV/�	���tR�AVsT`��P��g�όcE�v����4���EI|�[H����߳4��I��LqF5�i����=wUP<qސ���.�:L��كzld��S�a-##�㭞\��8��J�'V�E�ؿ���#�H'�m���!+
̸z���"��$^x��4Ei�[KT,���g�O1y�$N+A��.Lԟ2Z�:z@W����4H� ���PV�;~A @��q�{�T�{�]���.���p_�.��'E��I���zj��;z���Jt�1��g�s��5���3=��$Mb��!]
�RόPb��V��<&�j^�G½�R{�I�#+��F�7Z��T&s�ܝb�{��2ыRܯ-��͌�=��z��	aeqtEIΫ?��^���/�ÚVV,Km���ӀT�z����3\x-�j�ݜ�J�OR1U���w�H�"��]Q�	�/�D���m���8�&@m���Ŭe�ɲs�i������8�׌�0n��y� {��7!5ٜʂ]����D��Cf�k)�>}�٥���d��{����4�(w��JU`�m�T��G�w�3�?y��)ن<���%�S�ra_č��2ǁ���:<041��fH��V���˕!��Ҽ�GO���{�g:�"�HLq��΢!�l�(��I�H."=��I�~��]���+TT��9\fA-�P�ݴ��=Ƶ^����0w����y�=c���7|��h�V=�;?qw2�PͰUi�����xePX���N��l_�*�;���c������������F[ޚ/�e�C��
J��b!��Tf,^�i��-ex.f᤻�jF���X�jC�4'�c�cV��:@��u�e|�}Sz������#���5�^zH۸
�+[m���?Z`�Y�z����+%�����#�%�I��V��Зr�
W�0sfo$O,�Ytd묘?&�����΃%6����I.�.>�%��j �-pMfA�����`}�TVR-�I@���2��A]���&n�Jp���p� ��**���sl�G�i9A`�w�WU��[�Y��r<u�
�,jVh���_���'��g�}X�@�-	ϹO�f:�26-+)�?\��"uj�A��@2�����2�e�30��U�r�")i�ӁV��'�a�5�$_������Zb�k�r�gz�ˣ>�:*2��Ǆ+��W*��w��:��=�`a^�݁�k��ɗ��YGx]�6��ʯ���.�,)f��j���ѬCXs��ܽmj��ٕ�T@������vJ��LW�E6mӒy����J[��o�p�+~�(�\��.C>�K������1`��
�U�5�Q���P7�~�v����9�N:���a)��,inN:�3�U:C�X�m�R�� T��5����£]C�Z:����d����[tj����J�P=M��˺W��!�1�p��m�;fe�@�=���@릓�LN�\z���]E���wN��,\	��[�r����ChuZ�p>*~�z��,B�4ßc����~��F+f>`���^w�a���L����$�o��.7���"q`a�&`��;y�p�M ��2)��bCIz}B��0@�i�W��S�s?��0n�x����[� a���C����/`�����$���w1X!E�d�)�w��Lb2'Z������H�����SS�`��k�����r �$�����,���t�V����2}��{��`����{/DVtYK�L5o,i�1����oL/�-2����d:�=U �$�j�h��it��7k������3��~OZ~�H��$ؾ�U�#�u�oCN)+�F �_��%��3O�,^�ۗ�$|>ݺ�{C}�T�?��2��ؖ��o��(
�6���q�ʞ~���³x|F 2�t��os6�$�>.��vz�G�������Cی1��Ǽ͋�������c4�+Em�%����F)�{Cu_��͎"n���rƧ�S�&*�vؠ�6�D����%Ҭ��~.0���y����}۵I)и��`�j�NM�X-�Z�w�lpр���/��A��)>"oA<j5�a�n1}�۬=�+���vG:�Y�(��������Y�ju_��(x��o��4t��?]�t|�yH��N�N6�j�_�!�)����R��{��Y�T��eE|Ԅ�#P�*�&���~Fp��2�J���R9�uu��o�Z�(К��n_R*>�r0B��[
G%촏Q�[����_�ÄWi��|�o���j0:�%*�,�RgX
X_
l9:����X�Z�N����&~��If'���NK��O
 r%Tb�{<b��<7t:�~�_��o�v	j�,W�����U-h=(Hl���"k�c��U����SI����Q�]� �Q�[ƹ
��࢈(�b=�M�~���xE�)|�g��!4��د��NlvqH�{��~i^Yt�מ�)�~�A��!��P@'�~������(Y)����*�'x���;�
)�<P �]�{RA�R���	�#jdܖL����3�1ƪ�-�:������ap}&ۓ��h�$��F�u�d;*��m�p���s��}�8�c��迋R�ȯ������.�2u#�	&F]S�чHC�������A�1�$-'VEnz�R�Y�Y���o��uN��Frw{�Qu
k>Q�[EM��+U`�nŝ	�iD�V	 (\��4�ǹ��_�F ����dy�d�c��:i�U�Jg��v�1��F�v�D��sCJ챵�sH�h���U�:+2h$��A�^k�AԌ3ߡ�1�� =Pj&�מ���y~F�0^c:����pL��9u ���A2~�о��}���ef"ł{gs�/58,]�sB:�иή%�&�!FX��YC9��O����N,�P�`�O鏉M��Ή��)QB�N*����W�_�}J)֓�;NV�:D��-��T�+��n"񁃉�髭 Δ�?�N�`�)�é�' 6"k ��SaȰ[�����j�`(X���nu���"�(�E���0�A�ҏ]}��%�TZd�g
�	+�"뉱�֝^=��/�E�X�ѹ�ljaOF��i	U�\�Ķ)ۑ�� .�=U���r����΂:M���n�2^\4���K:�|XZ�Ц��x����CVl&*h��}ovi[���qꟖ�]�k}��]��2j����U�f*B�ͫ��[��6��=� sx��l����6���d��klD�z���$�ə�7z�h����C,���^����@"����%����w�ê��(RI�D<�L�s.T��V)��>l0	=Ew�Aq�{��X���*�Y ���$pi�y3@��arj��F͵&,7;��-��"LG1���m��%�L������'���|��}m͛b.��f�< [� �s�m��,�PLAK��L�������M�վR�p�J����Ѻ�mo~���g����[Q}o�b��[f��v���zc��6�ª�ں:���5����F��0���3U��I.��,�M8�}��Ҵ��1��,�TO*	C����ӊ�A~����s��E5ɴ�oӜpx$�[��������s�Hu�Rn�a�IY�<`!g$���*0���x"�Ī%����Z���0ܶR�B�Ҙ*��}�0�L�� ;���.^/=��I��%��E'5��l�e֪!&���I����&�&�����ٜ�M%Tjm$˰`�[�
n��,^k�*�d��	M���*ԫ#��k��P��l�G�P�������a��"��K8��B0C���4����w�X�/�`�x8�ib*}G�#G
�z����Y�5�T|��߅ݯ�y��5Αj%q;����e��S'��N��z~FLi1�eD�ɻz�j
I��4�:�{LtcDeG��}F8{��]��߬dC�[��Ӑ\��������rߓ���/��M>�Ψf��8-H8f'�Y5;�����JXF��A��y����=R�$u}c/�{�����4k��p��]���Ѷ~H���7��"�'Dq1]Ê](7z��e��6<���;�0��lc�i��){�VP�8�Od�Y�<�!�8RU�4.j?y��B��@L�g�2��O���\P�������nk��4z;�������=����3��WmCJ���h���(3Tϫ�������Xݰ���P�<��:!n�?�R9�N��{�8�<�����U7g<����E�X������]zg;8�sD�a����8��̸��t��ol�3�3�҅�}Yۺ��4���tX�����.�e���N?��k���GXr�0w��QP��V՘;�PǝG���!P����I(���~�ٿ�C������ۣ�{�ޤ�B�h��뮫g�Ε������gx�.�@A</�_4&ɿTK�W��Sx��
p!EB65$A��U�ӗ���k0�^����	�����Są̂��������XS�P��Q����dy�I���:�$�3���[��g��߿����1�XS`�|��t�Mn5�q�2O��{�5�8c�V( \�t�+��j�R���!;����uo�������I��y�!g֨i�}��C ��g���d�����\���$��l�5,?��& }�U�`�}��Τ��'���v)�pj'�Ug�݁X��&�I�w�8EȾ_^�<��3��>��r��Я"\��W�À�mX ���i*Z��j�5�R�J�� m��J8��}�>�$�9�6�9Sƕ8�=NbB
���閿��_��nU��n�R��-^Iv�uA#ʎC~~cf^E�%�U��Ui����n�K͸
�Ndgc��<{}�ڮ�(|������A���՛��۠iq9`�<���H�3'X��ȼ����큵wn�Pע=dߖ���#_����Tg���!T�Jʰ��c�p�h����檹$<9���#��pr�<֜b�]3(}�K�t�/1̖-I���I�.J�PPIlM�4�L͆��e.�wcr䧟C��R�G��>�o$Ck��h�5n*Օ-�."�2�ES�ԶT�J��k5'�c��o2��t&L���g ��{�
�ܟ��N�VE�$Gf��\`v1 ���������L���P%8��)�������y��w��[��G������{O��	�ȥko�y�����'� �7bm�ի8�Ik5����>�]:�9��C��gW���3�&� �^�.�LqRH�s�?��7�%�e\�$�"�+�Wfj��s��Ʌ��1>O�D��/c�U,I���c	���F�5�*�l��Iv9�v�ǌ�ﯩ�r�9����M*�,I�p�͜!��L�_�|��:�P�"4��u��`P�D�'f�?�a�	�l�b���t��o����QI|�b-���GA��e��x��h�t*�x��_u�N���w���1;�흯��7j��Q�-�FrݥԲn��"�)`yۡ��7y��4U��꯫��Q5��~������Y7�KΑ��1#�>sy# �c��`k�A�0��Td����k��l��^���M�u<=��\3>���#l�_j̙�e�V(AM����S<�7@��Ŀ\��#`mB|���!7�[-{��9,����Hiĵn+�8���鲩ǹ���G����e�D>(���A�$����P1칠U�'9�NQ�dX��ëd��&U\^���? 9��	�L@�xI��-��+�o��`�ڤ��P��������Z�o�TG����r��^���T	�a�.V�B�G��(�*�G���@F>�$�F�7�`�u.2O�Y��ZP"����@`�e��?CLj�[����<�B<Z�p�V����q�B,8��ۊ���c�e�F���FגȰ���>
���������{Ёֱ���x�
JE9z��N~�g��A� r�ZB΄��p
n�GM�ґ-HV��qϸc��Ĥ���OV�S7Z�
JuĮz�c1�����ÑD�'&^ B�C X�}fm���5�Jᝁ��
̮�sR:n/���&O�*�S^f�r��N��;3֖P�u�$�F�ЪiR���6"�p�N�Y���s#Y����hPR���O�n�k��k �5������9��E�eC(��ɱ�=p�r	���������AP�7���1�ռg�<�a��(~��fR�+��B�<!��!����v�Jl���Ե�P��G�\W�<�*���i��d�ˑ6�Vi}�k*'��{�~�AG�?UxZK_��s��v�q+b�؇�~�����:c�1s8����}�|���V��SqaO�t��Il^���ڥ�c�1�⎲�U	4��>�j;�x��s�n}��k�16I��x�;TP��w��Ʌ)��xһ�Y��݅E�s�P	x��&����ػC����i6���o��>V���2��v��!/�2|&�<�� ���_Y
8Yd:�9��.�F�&�F
ck�������n-w�c3Qݮ^�'ѵ����Fc@�y U:���V~? e��0����/�P����6b=��3�n��Q!��jЯ��VK�I�����c Ǘ�@	��t���K5i&�l/������,>_}0ʊI ���w�͊y��$|,3�Xg��t8�a4P�r�R{�4d�X���N��	���>��8��=7����0Yw����Ṅ&b��N�ȥ���Oh�EaVf��0���Z�_�ٷϔ2鸹��E������Y��b瘳%��c���5H+
��eF=�c6YnO�
�$���2���sH�ݲAZ'jZ��d�p5�}���I?�T�-�{�s��K>�H1_��K-	X&T���V�����o�e@x����W9��yp���p�MH����6��h,no�NtC#��E�e��HJsz�	�Pr�|J�|�Ǿ3����GvH֖����4��iۖb2�-e����ԃ���T�90� �A`K�����v��d��BS[5�{;1[�xF<�~�� ���f���~��\�AȂ�����[d�d4</�jV�jCD��P쒰�@�_�u�&�_V���b���˓Ў{�|�?r�G��}��J:����צ��a�%=��-ѻ�Glq�Y�28�[N�j+�ɦQWK�"
Q��OMl���
��h�b�~�5��D$�Մ9��a����g晡��wp�H|ÿڥ�����ݹ�JF�[�	��b�Ų��a�݂)�C��^���e��3�������_M����"	W�d�_(H�<4�����G�yl�+��hz
�9J�����X\y20����@tQ�# 0���<��NǪ�ӊt)
�K�=u�Ć��NU1;to����b"���cV���4R�\D�Oe�~��Bi�m���D���+�C���~˝H�f��HӬ�ǅ���<kگ6�L}>�[Y�ƒ�3�(]#�3B����F�zL�d~��I5\�I؛��Z��]]���~��Y�y9z֫��I�Lw�ό���i��3�2�L<�U�M�Ũ��(�E���Η$��)�N�q��a�a1��2�[��N"EC�B}P���y��{͏�R<��,]�F���P��_�՗.���G��+8�E1О�IHS�u����)!�S;R?���")�N�Y\���
�zF�T3�O�3$x̩�A�?�S��"2�Ŋ�k�G�윘E��J�5A������U맇���L�ᾫm�b��>��o)l�e,��=G����~s&�5�[�$l���.v�|ذ4X䴳Z���� m�*Պ�9���׬8��h�d#<
X��X��99*)�Ծ�V\���Z�~�a{]X/�Got1�%E�2B��Ů᥾_/������غ(j�w��T-�줇y�� $=�C%�r��~��F��`��1�[��/�8�c�D 9�l�+��7�B�+h��y�� B�x���E'����٧���Z{ֶ>��W���7��4�E9�8X�*���@��
]�Y���~�-�����cM������ڰ�*PTb9������LHQ�[2\.�<�U�jYV�81T�N�<[��sw���:�s/]�Kʻ·��<ç�oo���*������C��۝;��l���L�}^0��R��j�k`	q?L�0��hR��Z"�)pbA�J�8���
���>/t��%x�g����dq?v�6D��뼹�T3�<#8�)#c%ևv�6M__ٖs�����]�j��}*����1���Cﰺ.i���GT���>���q��'Ֆ�y��3/D�:���纗�IZZ�΢q�'%��<2Oi��BX�����y ���θ���;G�:� �M���W^џc!ȗ�S���-��E�l���� ���C~�(�}4�C�hv�L�l�b|��u[)Q�;����}�M�x{v�ij\L \��nͽ[�9IWa���j��c���j5������r�@�|��t�~�8G��D�e�����5�m���tՠd����2�����Y��dƼ���k��8&��{/�(۩�@�� ʦg��h�:�������S�JgRK2�޴H	��H�;ϳ��b~��2i���)�h7�U���1��it]�Lޠh�h��2G�j�I<��]%��|�a�>�M�<,#�/�l�������a��q��Q �Vh�LE�r"�^$9,�F����I� ���$|L/�0�*}y�0�@F���JY��!��;����>��/��.����z�-�.A��6��?|�}�]8�d�P�Ѡ�&�T4ě#�p�̝�=A~�+�.�7��3�MT$�6&?s��rc�
�9]�:�F ���&;Nw�fl��Y�#�:��5R�?����]}�����>r�,}~l_oȱ� g[�]���ԟ�Y��N�C��YZ|��r'6�q�)a�w�>A74�5��K�X��,�X���(Q�;�7
�y

y�;�"��7��~.K�K?�P����և���>`(��aCNL׸`�y`F0e��!��;g��V��&	چ�7P!��"F*�!�[v�z�ik�e�ʕ�ۄё%���z^�J�F��j!*E�W�����^lE���)8��!�E� b:�G�7}l�<Ǳ���v���+�*&�Y���8�
��C[��k=�!+:��~��]A�(�$�R��v��).yO�DL9���`�6kG��P�~��i�Xk�rYT�ˍk��7q.� �Jlz�f�K3C5 ��3��4`�-i��D#�T+��¤���W	F�U��C�_�q��?����v[���Ԗf@c!5<&je��mI+g�$�=�<�L���+0HM�,�Pdgq��k����*�C5ّ_���a�p��/�z�'���q��Q����ݏt�(`�c{̀ "`4+}0���?���'� ��J�	!B=�`D���9=�Q������mw�_7:8�Z�ĜRv�����g� � ��T��B�h'¥s�FrM�l��=X�y��Ԧ�rl���ƵT�`y�P��[э���y��0�"ϫ��n�u�봿�<RK8�A��W�;�)�T	�pU.Gz���%�b'�5oMM46��B��6Yu's������ju�:���T�<�|��� ]~�
�_�d���{Q��&�"y�h��V�,D���o�q�D�����0��6/���z�'�,����Ci�Ӣ���bgIM�ا'�ˢ������7 ��0�7�-�!�BoĈ��˿:��`+�Xr�O��X�2�#�`�L�-�#�)�V�6#�`����G����87g&\��*��>��){n,ؼ;�
>n�p �!����"�\����Sy�+��<�1z��G���D�ݡ�-4��|�8�w�Ŵ��TK6nLGl�Ϙ���YYpqb�-�0�}Z�P°Y�?(�YY,�h�1Nm�)#F�B2�h��Y�J�ڤ|p���
�,�X'?�i�	䚖*!����aʾ{���f<:c�}tЄ�}��-l��X�
��*�:<��E�M��'��dN0\���gł��wl]j��Yo�3 �$K{�*q:G���Ri����*㰭�ţ����e�w�S��V 9y������}� �,���W�	U�#��n�Ia���V-#�Fy�ӈ:�+�"����`V����g�9H�-A1�2�6���1bO_�w��P~z��u�һSQ%n\�S}�U!�:3��*���87}��G|9Q@н쿹��Juĉ=��cr<�35aB�_���j��y�G���/��m��wWr��z������@|�������|e�L��17#����̷��7�7�d�N��˒�L�^�j�ILM�����:��	�6|�Ӵ�(W��4�	�M��/�@'z�<r������#���ſ�g4�z�#�z�.�-;�uwM�(�����(�<��Pw�b���AM&�5q
�Ab�I��?zdD!�#���u�4���ɔ�o ��-��FOŪ���@����l`W{�':91��!���|]��St&P�����Vt�"���#__�R����$�w�[|q�0%�ڬ�KO[�2%���y��m�M;@8l�O�f�F�Oނq\ց[M��T��/�z�#$�Jb++g@*�-�͸���3�J�^2;���Nm��k�f��ظP�����E�7+�7ϣ\.y��,��R���ߐ=���m���K�x�)�g�Jǹ1BGYl�M��r�M��B.ذ*޳oӺ�P)�`�ga�9[^M"iq;�?���y�-u���&F�Լ�����c���;�+�d=pQ��#�?��E�$�2H��=�q����Q:u8�q;�'�K��P������W���o-N���lc~���������9�aJֶ�.�7��ʄ/�Y�	�?/���2���ƥ��w�E}w��CƵ 	�
�y<��YRF���Q�cK�"�˞����O�W~t��*��&���������b���.���Ż�3�i9�Ġ;���S_�z�"K���h�$�-�DBFt00�dŁ[��7�N��jb��Ȝ�H'ijL���m
7Ti�[E��pȽ�"�Z���.���*�c���~+"DN�g�,�Y%���U�V��3�ޥ���'W�v��+�cQ�0��R6K�إ� 	�����.	|ʊ[
��rrTӻ	�~��7��fk�!�b�q����8+F�\���lݤp��c�w���{s_3&����w�l9�9��/QbNn�nc�嚌�.���n�)��c�fW��1P�YW51v���sfύ��wL-����"K�"T�7j�>,��4="��at2���h$�V�(����|��JOR��u�X�C1�%�)��'9���㋈�>dC�_�X/+���(������1Ԭ�1;����`���e�㕯՘�S�4W�
�;Ƶa�gt�ᗼ�gɜ(b�J}�-�BX��V]=��ɉ�m�t\聃ʚ�R�^�<�~!jV���Q", �)�;d:)�*KՠZmƏ���/LmjtymŘT�p5�9Uדs�&�v<� (�����	�l5�Y��%�mY�h5i��$P�V��E�(c�T.�+��qo(��R��R�	,*?�}�
YK��H�{
~~q��J�Vj� .�D��{��c_X�Z��i^륳!�����g7M�">5���� ��@J��df��Cee�}��eqD��*�h� �$��&g�	�Nh��P�l�c����T���I��f��
�0S]�^e�_?�y�>�yϚ���-����3�V�K��_P,8Jr��e�#T?��"��ɤ�-����'&C�����d>Vh���Nԛ�rJ: �l�ܭ�a�&���8�,+����N���G����O~�a�bi��/z�k�"ż�:k"���K6��V㒑�~���S����XB��l����=��Ω���90�����ल��4kBױfO�q(��J�:yh1�$F�W
%��/�ue��n)��m�:�6��t�!�����mA��d����V���)�H��.�U�<>�P�"_�nd��ZI��v�m��g+�z�f����V��pb�5� ��JR�^w\��[�E�;�����1�1���h�H`�7D9o/H�h�IR�W6�?�P5�f2������4ht� +!t�4�˛9)[�����
��o�qs��x��~R*���P:M�G�O��(��7��i_����'۽���&~Ki���`�?�B���=�b��|H��./rn�)�
=�f�x�����ؖ-Y1Rm��qD�)�Y������)��=��b�>i�Wo�-&^a�O�g�`Y��q�$����h��G����b��?�)�P�=����]0h��
"MU������f��k���-V�,���#���Ҝ;	�6�V�=�Pm��5��RVe�k��&�1����X��u�҄S��hHkAy�;����++MiEqQ�;|�hK���������{��v���dQ,���0A�?jo���)���7S<M��_���kʴE�����.?�Hǆ�������TM��Q|���rȹH�
�YHT��� ^�����,�g��eOW�C!oN�oƉ���9_���T�~A�+Q���)�37@huv'T���q�2������r^��iG|�.[�����c1�����<BGI�*pu��``+h�~�#�i�ۇ仗&�.z�,��� ��$*aZ�����lӘSp���"Λ'��T=J ������J!�;x�~ߓ�%�cOs�?GiNlL�� �<�Rt�P���_e��(^����}�Z���Q���Vv�4�m��Ո�U>����T6���ġ�Ԃ�<B5���=sc�KGs��r��}��w���2���N�L%�:Dׇ#�:l:wDN!�O�.]@k���ucH������Hd�
G��<����%��E���h��b���{� N�W,�3GT�|�}��O�ZO�&,�9�,�+�ځ���M�K�B^@����ܹ��'zYuX̴�2Cdt�e�V��`����'f�f9��aU<d��@��0������XQB�Wjqh�{e�\���@��a�)x���p���\ҝe#�7r뮢��2j?&�
�>6����C��H�U�ϊ��>��#�j���W�s��Zl9���%�Ů�r��ъ�����A$����\FJL��O��9�$�W��!�-���$v �=qe��<�)�����3��Ϗ�%�Y����Ou����C߱�V��/�U+{�F%bЕXc��}�?�!ټ�t��B0�i���r��W9���6P]����ۼ����on��QAe����iN���GbU��C���$=����(�X'��F�G���u��^�[n����O�(U[�v��f��|�:�g����;�(
�Ok�w��uM��`�~*MG�20�R՗����m8q���ܟ��B�=��q��`x��Z�^�(�"� �>R�E��31^�'��|^��ك�vl:��Y�1ǦuS`z�r� �m��^�6Is"�^�}x)��z��7�,Z��lY��/����y ����\9��<�U������pފ�Y�Νe���t���1� �C���3�w_�Lm��-$/��#��j���}��ʢ�)��9`Y]ڙE�?�D�L����U���%��p�Oǐ�e!���Aΐ�,V"�dZڐ��z�Y`D=�y/3i���W���z)]���EN隁���߬��$��B�
��4T���㸞rcJ���������Q����0'൙��jf��Z&u��Y���px�2�5�_Y��/��ٺO"��\���_���}�GӦ�7����?�^yV����P
|O�=�2 ��c���3Tx�`����j�G%�ðQ�dj����Q[�o�|���|�}�eTX�9[jC����;Ϻ�Dh�w����z�46$<�� )��+袲��ֱuЋW���(�6ɔ}�t���{�.���Qx�n1r3]��y��od�H�!�������[.�I�$���n����,��ޏ̐;���c�ǐ�}�9DӮZvZ��NK>�r�/n�� ^?�#U\����-��I�A�Qc�{��������7�R	�38�
��}�v1k�4�x�~+����!W�xGׂ�FY���Y�y����7)���� �11s:��%l6[B���?���R(��*�r]��;X�a����c�1s��֑���{���h#9��r�bΝ|�cg��F��_�lr���T�&z��Wb����������|i�n{C�ٯ��7�0� -�HƠ�W�!��������梺R/�� �b�5���'�o,��3����I��5o�^�k6��L~���$N�S�(l�X�xJ1�ce^�#�15�^�=X�[��+j܁f.�o�^���FA��Q���\NN �\�+P;+��r�ifJŘ���S�op7 �;�8�hA?)�_�~��J@2���*4�W��Ce �`Zɵ��ɼx�H^�ɷ"�f��Ķw����<cy�=����=1��=[�p�ǥ�ט��E���i���)��bj�6��L��G�V�-xl��C�a�|�E�`��y�Tm�]��m?��n8e�Wh����f4
���� �Y�û��@^G�C�Z���my:oR?�4�Dֺ�󈗶���r���N�`���Zh�Q��)�;�)ǂ{����'��@��an;+���2��W؏X�أ�N%���^==��D���2"�@>��D	qG����on�ڥ,t+��i������M��F����<_�'9X���t��r���O?��4@�Y�-Ⱥ�����;�/�yױEk�2SD�;��:�F��4,�]�qF��gSz�{r9~��iK<������ �<��bJ�I�o=Ňf�����HZ��>���	I��LT��6�ld�� �>/���'m=ESd(�G�2d�HFܳչ{*E��\�K�b�M4e�x�����/�ӗ�$��I{ļ.���wL���]����q��̐G�]����,�<o�R�qa��'��̇~@�"����N3h�Ԅ�{�ӂs���vs!�*��'D�g kV|��k��7�$O��n���v�mX@Rɐ�pt�G�~ǅg���/��(�_�C�"���|���3BR9���Vc��`{�U��jm����@a(��&�J�{��K�� �&�z�.�Љ��"@|�<"905x=.	G,a�x�]똨=5�
o�{� - �0J�"ErC�X�b�b5v<D8�O����	~���#�5�bf]c�� � Π�	~g��S�,��U7��J8Z5�n���ҲOE�oWF��'q��ĞE�D�8Qb�Ӝ���������Ʉ|雍�e��h��i�ڔ���'�!��l�@z�4�]ǜ�C���PqflL�#��{�\�b52���
<�rm� �-ŵ��(5$5V�_��A�$T��z���]GJ7QwU�L�;��
�ȋ$)JS��k���-ƋS���@xö[-�ʻy=턈�4����Av#�-b	s�1gV�dT���ѩ�~�ZY�-e����A��&��x]B�22է���{�����Mސ�s��o�v�{��%|�����91�,�w�6M|�F��&r���3�|р}�Ө�¡�kz��4Y	-JJ����x6D����'Cz	v�8s�t�3�J�\���Y^i=|���Ĩj�/L����KgrT��ϩ(���g?y{!㩅��+�K$���9�c�g.=��Y�J�Y�n��՜����2��۩�-c�|̩Ί��M�g�܋@8��5.�Ǔ����^���|�y�v�wob����(���)_4u����P������4�OtL�(*��(�q����0�D_>�� \*�j��2Յ�(zI?.~Cq��C���Ei;JW=كQ�M#`�h ��E)�B���C'1iɏИ.���.|#'��N�DF�"�PŻ�9���g�(���؏3����e���ކ$1����<$�}�i*���6�Y�Rp^M�����kSȁ���.��o��fzE��A[Iأ��$�o��*��'@��tò`�D�z��'�R�
��E���5�S�d�}KD]�����nu� ӻ!hһ~b�`����sʙ�B���?G���\��Q#�����;Y�G�-j�"Ъ�,>Ԭ��:߁�$��Mx����� ���=2��^�p�x�)?4���ќs2���Ѿm8c�������W���R1
��h�O=7`gf6��]�}��$�e�����`e/sdP����j���|h�>m�5}2�=���>ﮦ���k'
^a�Zja�ͫ�zdn� �=a��l�U!ܠ��8_�������U�W(&є\N�*�g�m����Mp	º"Đ��eϕ�Bk��O��9I f�ާ#�7��<��`�d�G�1y>~����o�5�̠��%L�-����R+����#N�fF[���y]*y����ϲm����!�%=3�:O?K�x�`���1>�9m���O�7G��*�L�1�.��t� �׉�&�������u� ����c���ؿ2��b穻�ݎ͖f�=a=���]9�N᮪q|�vf�u�=U���Lv8�M!ݨ_tٻ�7M��q�Prtq_sN�GIfH�UO�a�3"���*Ky��j����Ic�ӫO'aԝq�rJ�߉v����F~�΅H|���!���% f���e��
�	=�q�(M�}L����*�9'â{Գ���:����@�	��|�R����)~�r��j(s0*yM��ore���*��p�wU�(�iZ�\K���9�W �YQ_l�:���n��o?Q:�Y�_�,#��EpL�>�;�UB�����	��<K�G�1��:���i�v��_7��skh\_t�k�|l �x{�*�d��E��$����C_(�
�|.���w���ZmY���vP1-������4��8cW�s7t�+m3��&���ChU4�7��:i��P��H���F�/�z�1���H�a=�PN*�C�͚��7�ky��{iŶ	^`=u(��ф�CVy��aH����]��b
��t��˼a���A͘��A ��*����}K���
��3������>�K@��fX=MQM�	%�(76��cy^�����I�5$�cf��dz��5dٮ?� �H��?�*��<��|��y`����^�۝]�ܙ�9�k5<D��8Fa�v'T!̏`�]��2��9r��=`7�7G�6c�_`xS�N��y��U��/���r��I��0<�,�~@B|�H�y(�D�.D(�Q��3vR#/=�n�e���%GnG�����k�T��D]ѭ�����\����BS���3���g<IqN�r�	#��:��3�P�|Y|��WWC�x��D�J�I�LQH�S�1߶SDb�G��/��S&B���ZN��h��W��z����#�L8q?�7Nh.�}	�Ȣ�u��6��yI��v/1�{����l��BqٷT���fO��䮝`�1�#5���ܱ{u���?�Y�-�'2Z7��4�\�S�R�������of�p_:�����~ù��`
-�TI13�"�W0�
Z�J�o\
�y�H���+�1J)V�|�&��j��1-it�QF�����Gt˧�׃V|;�E�|�̙I!�Q���A(����>�����.�����g\���*�`tl�s9=�X`�`��F� 3��\O��"V1!l����s�gcM[�y�K����aK�A"�8����SQ'Lw������|j�0�T�ri��#�D�F7�zA��7B���J���REfߜ�*��1�®���<8ꙝ�١u�����:����x��}�xU�7��0|.J�Y���	%|�����+ Ba�>.����o�2�7�m#�C�_�$nf��}aU�?�}��k>'ӈd4���g]Z=�Ӥ��n������V��.���LS�(9���l�1ϰ�8���o�AEӞ�ӍC�	&�?o�K�0h~ʁ'�RY�
��n�$3�1����r^I��1" ���+�GQ��������X\ i�_���M�;E?l��݄�|;�~��c,�JK
>��4�7+�(Mg�R���9U_GL�}/�W��o~��so*:G����7"�B���62��h!�<��n$�����9e�Փ*�?���J��Mڼ|H^2�7�"3�&!��iar���m_籆��OJ����#uk�|mX�6�ա�R	Zz��G��rA�4m&���S8��V#Ԫث]��5(�������.];/��Z�-{�	�4��u�6&���k�:�
"�-����R'��T��2���7�   h��H��b��c̾h��c��s��r����r��c��s��c��rE��c��6c��j��e����p��@��t��&n��b̾h�� r�� c��&i��c��1i��4o��3��q)�Yq-�U3�W�S��Hu�   tLi_�T���0�i����\�-�ze}�NSW�s��ò��k%�
O����|6/ �����#ǃȍ����US�����=�-[����(3w[=�v�q��^��3ċ�3���	V���F�F�`����ya^`��Hm5-��-gla,t3���S\���   ��3�3�[m5�@��  �; ��   ���T�S��j}!�?*ō��1�J��]4"rLxtX3� +�=�?";�7�:P��_�^&���3���n�� t=�b�%J�<X����X�3�X�#�Ã� u��N���[��t�=sa3��+�3�5�#O4C+�����Gf]�   -�0q��5_Ń�L���u ©M�0�  ��ǁ/|K���#�K�������rY���t��������%�(
L���[�3�_ g��߃
} ���A!=X��$�-{E �>M#����}	��N[+��^~�xѯ_LQ9k�q�=~}�=7x�W�S�   3�%"e�i_3��ȓ�2#n����W3��3�#�[~t�XW��3��G�1�#ƁǢ��43�#ā��   ��O-�)�7�Ö   �������������X�^�W�vW�lw���@9IS3ċ��ޑ15&Ed	�a��g��āÙ=�=:0���
k8I�_�Q)�|�W��   ����W���V   �J�:V#�+Ë��]��s�F�QAY^`+�3�a,�t��[-g�C_Ƌ��3�+Ƌ��^q_�[�<X�f&_�/<�5!P��-3���PZ�&P3��3�X�'���<<t#3�������z�>�ĸ�e��%�N�M�	,sDS3CSraoC coirtaeAeeC8Fpte            3= �<                     �= |= �> �> -> @= �= �= �= �> �= �= i= \> �> > �> n> G> > X=     KERNEL32.DLL   GetVolumeInformationW   GetProcessHeap   EnumDateFormatsA   GetCurrentProcessId   GetStartupInfoW   ExitVDM   GetLocaleInfoW   EnumLanguageGroupLocalesA   GetLogicalDriveStringsA   GetLocaleInfoA   EnumSystemCodePagesA   GetVersionExA   FreeEnvironmentStringsA   GetFileAttributesA   FindResourceExW   GetPrivateProfileIntA   LoadLibraryA   GetCurrentConsoleFont   GetTapeStatus   GetExitCodeProcess   GetCurrentProcessId                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              