MZP      ��  �       @                                     � �	�!�L�!��This program must be run under Win32
$7                                                                                                                                        PE  L ^B*        � �� �  J     �/     �   @                      00               @                       ��/ �   p  $                 T�/                            <�/                                                   .text    �     �                @  �.itext       �     �             @  �.data    p   �  &   �             @  �.bss     `          	             @  �.idata   @   �     	             @  �.tls        �      .	             @  �.rdata      �     .	             @  �.reloc   �  �      0	             @  �.rsrc    0  p    0	             @  �.PEPack  �   �/  x   8             @  �.xpr01       0      �             @  �                                                                                (K����4O�����$C��X,���\��!�!=CՋ$`"�2AA	��xx�e}k�]�)}��T�52L	��R=�����!���m�+�w���^��w��m�p�d�@j�Z܀�/@my�� 6��my[y޼���wy#v� ����{�7�x[��������{��>������y��g����$���g��Y�l� ���l�V�pX���>�h+-,�ZB7�9�a�/�H*�c�q�������C���gj�-$
�sP���j坩�t9����K,��9C�N�v�N}�H�S�����m�W��
*՜�e��X=
Bb�ML�n��ؤ"��jC^"=N�+�6fu�����f&^ѕ����I�+�6���F@��Z^͈�I:�Ճ�S���f
�dg��Z���~C*��Q��9�h)���;SC/������V���C|�	��ck�2���yc�J ����W�֓A��SFe�@�r�|�G�t�4�����_�Q�#�m�=�f��֐��$�9�&��csn�=vS��9f��c��F)�Ŝ���]�������G,�����6�G`Ze��,|S8�t�/�D�'��p��竧�.���\<�x��\�G䩞��P<��)<�,�i�G�>JY��~H����~��?��OdO@�ƞ�rǹ3��g����'��`�>��=��C��x�����fG���0�!�}5@S1yj�gG�?U��=�e�j�����b�Ib��ee�3�3X�X��b_���MOΜ%�<���3���v�Ӏ?���mq��e$�me�5�v�{-���3يA�zfWXP�HpI��PDX�=�q$a0=8<���?i�s	(9,�Iĸl5/�fD�\]%�a�ľЉ�����BH�r�s��r��:Z	P8�r75fz�*g�iSQ����58�&p��,yPp�<��Aู�<f�2-Z繥Fz�OY���U��"����F]$i��?Dze�b���I�B�O���)�/N��t];�VT7 c{�����%�AtU8�V�: ^�(���'���Y�>��xKЁ��DW�(�E�k �a��Gp$	�_ 5bY�C�\3�8Q�i�B�*V��=�����l!l����4iJ���밽�j�?���i���gzrɟ5t�5�_P*�0@Z@#�i@�����+�M��`Y���^�dW���=�'�/��L>�oױ<p��]�:�{�����׌���K�7+V	ILR�h��>��Ӛ��|�� |D�C�+"Gy�V�(}���)��H���%�����A��A_\�(��w�Dm(�ps���7;�ޜ�qy-�T�2DS6���2h���hYiԉ�	4k��u�H�%<K`*F�ߊm0��u��+'˦W��u�-��j[ވt^�� �.�y����U�U�EX
�	(�S�)A`x�<�ڬ�)J[��$�fA:�ю��#�l�7�g�{җ(1����St����z9Ox�_Is!�h���A��"o��j��*��`��E!.RYM���y@d�t�H�2��&蕠�F�^�y�{����z.?�/Q�v������Π��+A��"]���tb-����ȶB�7¤H]��&L���CNɗ��!g�7�P0ɳKh��~j���l���_��Ǥ�4K�vU;H�i ����hb<!�F?]�#�u�8���nf�����"�Y�Q1ܡ(�-��?i��D��-�r�#_du�KP��kD.�.^m)�<�?N�r� ʜ��H�-�Ԕ�*f�ʃ{�^|�$��ڦ�z�۬ N���˕>�`�r�wSV����R���n(y�����N_�9�j��iϻLIm?Ŕ%v�0�����%[��{���5MQ�1�*Gd�dӺ��b�z��j!�?
T���VwW,��]y��2�D+Q0dU�X'daW���ѝ����heYC�,�Q>8e��"�)Dh�q(8Z�"2$�0��"���-�Υ�g�Γ�Q���b¢���Y㚽�[�ըա�҆nMz���21�M/�;��m��S��D8'dBT���`[߄�1�V���
3f�W���A�&s�[��2�M�$��u��bWԡ�����ͤ��GI�2�[%���s�;vr��}��Gt���B�7����"*,�w���q�#LP���x��K���S+��.�T���0M�d��Y����8��ɛ7�jr	�~K�:�h[6M��R��O.��nBK�P>���A����`�vθ+i���8�㘽]�pL��Ὓ��F}bKٻ6�	�������<cBm3��eV���'*Xdo� �za!n��O�*t�AX<�Kd��鵥D��+���=]t5R���_��pu0�� �AN���Z�EQ׽V>��{�7�h����
�hL�Kص�bQ�Qý$Rj��$$�x� ��uD����Bl�ַ�R�N��������ƫ��V\�g/���S��o�l�0�%��*ud-��?���ER�-�;�;����1x�)l��Q[[��HH��+�<����m9�<	���x�`t���
�N;6΃M��ü�j���#�
_�%�BK��D�2`!%��HϽs�"�1�L����R�&��[��Wa<�ֵ�����@%�^��� q��݉�B��[)K^E�6���k�� ��H����(&�� Wc����f=��vgV_/]6*L�+�t�����d`߰X�"L�3!ZP�#bT	�[���,�U�u�Wa^��8>�cMoP�Jڃ�^ڈ��yW��`�`��Q J#\=]g�%�!_fQ3UV�V@�Y�P��
�Q�H{
B�7~}�$V�(� �Y�!�˪���$%���%��&Tj���I�F;�ʃ�0�a��6�4�A׹E��cg��Hth�P��Db�2#	p�Db�m�����T5!�m'��Le����E��}S���;�0����p��oA��Ԃ�-U�Q�`/�W����֓dL���Ů�tI�.�Me_撞6��@�1±�~	�R�QkNGrD�g�"p�E'ݿ��`iЪ�Rgn�2h"�g-c�ƺ�v!����H+?�h(�nSe�\��A�1k�Ł*P%�����A�I�9�4��~>+��6	*�˂��Gf",5n���%/�U�L;+���C!�z޻wI�Y:�e��$��ϝ��%ga+����f��C~��*�n�*��	1.xЧ
�)��宒�"�U(X�s)�T*O��D`>ϓi$2�T�Ĥ��ԁla� �
/��,��-]_�p�J?/�; ��6^��.��r�y�
y: [�o�� 0��%�&/q)R*�O��;���l�}��O�G�ˠ���sk�?��`�Rȇ��O�qǝ֢B�Ll�gj�n�j�@R�]�X�^E�ų}>0��n<�E�-�d�����Dq�>��0�pZI�ÀW��L�Ʃwi��V��(@<� ����n�����H�()���(HeI�D�Z�,�1��˕R�'.�R���0'W
�iZ+����]�_1I��6�J������b`e�o!$ۻ�kތZk��㎠��,�S��x�l�B�\AV(��'L;.�)G,���d���xx������t}�Ij̆�<��4`''�P���4v��}���K
�3�5 (�����;B>5)9v����du`��F��[��j{��TZ���~�U�B�Yw`E��~Q���t1���K��W�"�Äg��Q�;Ysc��Z��BZ�w ��	6�/ajM������@�&�����#��� ��:��u����cuY�x	����a�`��N�k9�BȺ�	���>�J1Ss��?Z/Ӯ�;�~��(cS_�����j����K�h�4��K��X�M�]�nZ��Q �D_BK�`��ԏ�է,��փ��jX	E�Np"��|��I!���������g��Z;���衬���/Zp6ԳSxp����eJc��"��^U��׶�7������Z5C�H��ʔ�ǲ=]��8t��򽘑[3=��8	�ىqL�U���%8���M,�d��?�@���v�,��{^�]�ᬨ��R8f�]Bv��8�Z�0ٸ�5����E�!��|c<�5�q�Cf��␮͠�a�3���9�K����SX�s���LU�#
PW]�r�/���A Wz!s�:��}��*�6N�\wJ`�R�׊�� ������WI�K�4Ǡ5P
��`�I�Yň�	ۏ��`^q�S��F�1��&?����t-h����6���p�͇�|�ϛ|ĸ��.�y�B"hC8Y����"� �ꅝt�-����Bj�k�N�sܩKfc���ٍ��zR|��Z ��%�H��"L~��d��7,�n�MR�ͳ���&��]}��� 7`�%rj��������d[�-v�wCŵj|-��0ҹ��r�z�����\��.$��/�׾Rz���`�T�,J ��n��.��gP����j˯�ʸS�S�l��V�T�<���0�|�v=ʇt�y�ڃ�I�/7��/u�⬂`SnC��iJw6<�7 e�d�	F��{��-'�Z�����er��r��S�p|(��#���cG�V��(�b߅��x�ҡ�z������3�� �\�8�pn��.f��ȁ�_b��(yg8{]�Ao�׭�݄JRL^ߕ�3�1��U�5`�h� ^�J����g~$�`N� ݔKmH!���e�"s�@}UA����)�(�kk�a�a��+�FQ1��������%W.:E^% {�q����(�ꔩ���D�)PKW�S[�����z��S~p|�%�;[h��d��i*��ԑ�;�
�C���}d��Qz5�����5���?����6o^1���|�A�W\q5�i4eC7v���Au�8mу�`֢^s�'��;�HB��`@�N��V��3 ��~�]�9c��Y�S:B�`UĔA�=�Gy�1�Q좈y"M�����M.����i*��OgLF؊p��*I��5���%�7my�g\��y������Z^��	/A������?`�m}z�ffm����m�:�I��<Ț��e�<D"u��-d}{�)T��R"K�MD��o&7<8��j�MB�:�s�c�}��H�(~�������h)4
�%u�e�٩&�q����2$D��X�.�D��K�"�ၢ?@��~29�\6�Z6�|��d�nB�����P����Ad�6����e�r���������!�
�CQ���HN�)�O؏�k�$����4�W��e3�Q���8rlo��2� 5E�E���L�m�<�1@��ud��{������eN�6����z�s��t2����ДF��X�0x��ƨ��"�x�ѩ䌹4\Sc#�'L��ՐE6�������F�{���)�Eer��g)�o/]d�-��|�4o.�Z�-FCe�0��<�	=5��ed��U�Vwtܹ0
t�}��J� H���$�"��VB͒N������d�p�QT]�͵�D��f%�$���nY�M���Ũ����%��ǲl)zl��.���l�hxY�sT�h�j��7��e���2-�ʙ�`w(��B]�� �F�����m\_�6x[L�R'!�V���p�,�6�M'�Smp�η[  �ρ����v+�5mt������c͠������ܰ$ƻA��((�;ow@��&3A���v��&"�d���q�׭?�����~V�*��yd\CNh���{k�[�4]�L�>�6�9���`hE��V�J����\�Q���m'Y_?�(���l����U�4�|v�<�J*}�y�A�N/l�����Q��I��~�1w�h?e:X������ڰ���)��Dߐ\<�"�O���D�M���uQO�&Ŕ�`�����M���_\c�,��;�\�~���5�Z@H�B�� ֱ����"��
�f�5I#+}����jW5�#�Z��*�d�v��¿���������F��'$�Jr篃G{Uv*�+�R�ٙ��k��&�G���a�pn��)�qj�L�^��I�V3��0�5GU+
R�6V��IZMe?E�-��,vb>JK��_iف��O&��b�^@@�G?>�"7U�J
c��Y	Z���mNh�GQ��98ME�p���l1J$�b&�Ų����yJQ�1L�
&-��t�/���mS�7�����}��3���D����A���i�n�HW�~��o讇P�����3�]��L�����T.[��=���[u�Ɣ��<���*�U(�-dl@�xn��1�bM"�IqH,��GL��*
�2o���V�M�pi��hCJdS��*}�Q�]M��?���%����B��ԫ'W2C)ͬ-���v�0�:�A ��d��ʩ�Ed��ʩ���,>G4�N^�����[���@%Z6��`Cʛ�ȭR���w�_k�5�ٝ��&Iǥ��4g!�����dp�aF��#�x�i�O���Ǹ>��2J���p����bT]q��6'*�K���j�X����چu,� �I���'g�G�H:�`�'��~_����)[=$���/l��q/�/�L$K���������c�[��l���+�y}i�r���L�h��%L�t�G
p�o�(~���%QE�x[����S{�B�2�/ToS�v�k:�K�����l�VbD�P��T�͎�Z�-x�ѣk)�G���_�4�w�U�9�$5�o<6XcL�wmj�?r�nV~g�]��*&�'pZQ˺d'+��gh��&��,��w�v���U��"��-0����,Ga�%WJ0�P+?��\�Y���8S�(v��HF��-�}�ɤ���J#�3�`4��i��V��+��SU<��4�s}ن�iL22�B�^#�'Q4��#k�q���=:������j0Bp?m������'�_]-�Ж�N�[�k���qK��2'=��٩mS��7�0SV�6��@����T�5�K����f�%���\R��_6�Ӷ��[�Ϙw\p�%����n�A�N�J��ø���9���W�>��%��� ��o�V��ʽ�9ސ���	�����\I��T��*҃����l��%����ޏZ�	9��"���hӈ���_�ph{�z��8� Pt�8L�%ek4BpƗ��t��V�|�56#|�2f_嚞a_�ʖ��`���?�6B�ٜ!�di3�(�|�G���.� y7#>�7r��,K��(Yj_�L�d�����n�xr>��S�َ�S��t9�"K��>?2��X�`n�TOqM�������I�T8���u�@h�����MZ~���2�s��_V�9s�n��[�tĎ����.e��Dv�VI�-�$�W���d�}�	��������@�,�+���k����8KJ�Z�O��])�nB�b'��� ��]s�O��T�������Ch߹��y��?��/��kJ������9rǫ+���窝ג���2ۿ\(�c�a�*��a�k
UQ�V�o�=�%��CV�myg��,��-%��ي�u��yjJ��C���}���<�'�#���2kL|Ü71o뙪]6B�"��r���yDl�訶��g��s4,U�n�<�n8�c��c�y%E^	ӟ�������/��Y>������Ed��`$��Bd)Wz�`�7Y�tJ�6���)`X�5����_�j2n������-}�B]ҌU2�3?n����v˭6�3nC&\G/eydH\�7*h�(I�j9�����ZF�}���H������mA�BO,�3;�J��BG4��e�fM��i�lh,�J�x���)۪ ��z4Rm��0��xF�ӷ�w7ZQ~���\W�ԫ��Ɋ��=���c���*�-���Z��&[)_��Oخ_׃v}�`��Kp
�`E�t�/V�⿬�~�h��+�P�q��3�k�RX˗�4b)�d��L��������Zо��$�����Gn�93>h6��&�pj�pd�����Rx=�K�&-`6�=X��Czw9^����gT]����M�\5�4)�g�=��7!����鏢v�C�A�bU#s���/���_8-Y�D���a��q�<@�6#ؘ���7/F/^��;�h5�*t�7��̟df.�QmI"SQ��ʡX�W�`h���N������!I��ٌ�5-���)�5�{��V�bw�����%���w�=�Sk�@��ڄ��I�K �h�0��la����?�Qc��E/�	�f���݃����M�TU�d.�	�	z�/��U>7�a%/j]��S�O��a�W�X�%*��M 7C����
��T5jV�	R10G*�����94�?5L������h,�^�e��Sa�=v��g���T�uR�Rx-Q����?��ʹʚ'����m	H\�/�7�h��z�0R�L�FNy�N�(iuxYVl����1�M���Fb��lH	T^�Z�7
��*�����(��9k&����^����TdW|\HAN��oa�ye���~)�}T1m�TĨ���wo������e��W�����\n��@���Qx��v+WT���������څ)�y{V!���30r���LIu�6"��K�`��I֢��K.QE�W���d5D�FCO�SK��Ed���my}���8��EE�]4�0�1(BX�xW��6�ǳ�^cd�W�S�)�j�9)�.|���wi_��
�B�7[�3�F�&�$ai������bF������x���m�W9�(篒m��ѓ}����J���*\�\cd���Æ����iI3V?w����l��Ӌ�U
T�����:鶹}�
||��#.��GR���� 
�MC�0����TA��9xm�{ ���ںb"6?ꂧվ��1$�=��D���\�ۘ�&
.��O敲�xX�u/�(��i9��;¯#�'��nՔ��b(ꎊ��<Z��T������5N� ��x؝�ⶒ/��Boہ����=jU�h�M(�t�����%.�À�k˾�dR��#f/i���-~L��T�����au��JK��[Y��c~���΂�o0pq����V���^�k*���s��g�9v�Qv����s��]g�
Q����e�˯-�	��.�p_�~��1����^EE�Y-��K�!7�`���Z}+A�N�Z�߯��rk��8�Qm��X�W���V*cu�|qȶ��˥s{��&y�[�v�=��]&�����_��bi�b)N�W����f��L��*PO���o�3�������mD�G(�,y�u�H�M�޴�G��Γ\���+@�e���&��4K�������J~xX�S?@2�����H�n��)�u��k�K�TB4����[7H�)�"PxC�2}�<��XX
a��Nϙ=R/��tݮ�]�R,bτ����_����&���v�9��yęQ|����H�4��pGz{�Xb��nFl��S�Wս�wJ)\�">���yUe�\*'��F�o�Z��Vչ]Ob�3������i����Bx�R�i=������j��Қ��ƨ�Cs���9�MO��MO��Ix#H�w��!��?ٱ۩��k8L��:�{"��s���;�\[�.
c.~����G���VR�o^����5q}9~;= I�[x���RMv�~������s�y(��6ޙRȳ
�'T@�3������9��Ҹg�rdl*<�/�F�Q��(�½y�9�t�W.}�VE޺l��'�̢2��p~�%U��L0.R/�������$��	 տ��vϪ�ׅSR~����.�8�W)l��7��՝[�j�6����<"l�B���Q� ���u7������O�����F�Ѡ���u<�<e�5�!j3_�KhZ �ѝF���J�Wa�W���PR��sGv ��hr�BCA#�WI�����k�x 7/ӽ�#���I��Bs����h\b�Q��.䘃��A7s_�� �n�t���S�W��M7��hF	��u�Ib��M��fd���?�X���WuTw�؈� kEEL������L��d�Y,B�F���Wֈ��d��kF����M&��cER�L�Tʖ�5F2Հ�q��c_m�=|�s���π��A�y����D�d�*���&3���h]�����w�]�s��q�s�7���������{�<��>������;��~|��5){���	�m�5��nY-�89!���P�8�um!�7IU�*9��g��n�N����J��'HpQ�$/6��,�e�(�샐�
C�N��w�+1�7����Uڔ2(���")��)�P��X��n�t����ܚ�.��ꯙx2�<{�q��[jx)���C5#��A��T.!d};����a��#!�p����(��=�E$�:_�;<.g4�NFG*�>֫ʞ��;��� �Ͳ�s�c�v�(J3�"r����A��4�q�]�D�����������z��>&�P��F��M�MD��^�?�byN%����L�#��O<���� �
�,��j<�����xX�?uCE\	,�bU�`���)j�����f�ME���ʷQ�f���u-�i�?6Gb'�N�Ѹ�2�^�1�?�Z���ѣl~ڍA0�K/��A�	����K�չb��ײO�D���TÊ9��l�uUڎC�8�$�+.n�ƴ�~}F���:B��~�0�X)���y�AU<Q��q�U�EV�տ��vS���J��ޭ��@�b�[��ƌ���0��QLԛ��ѴY9`�0� ׇ6��k+�?�RT����_���܁�)\%� ȽC�]�Y	�H�_�v����~ײ�y�ѿE�w�+lVM�soG-7�VŦ��-2�[f^��W�)���Y޹A<\��Bt�|8!d���B�3x����)�����[��Ѳ̏�[վ����~��L5/����K~�T]�z`�O��4�]��Ѵ����WQڤ�V���@�MTI6���Nh��|w~��}�����S
�58�͏̲�%�)D[�
VL�''U
cT$Y'M��(љZ6�8�\�$p��G��v�Ry����"�Ӧ�j�t�Yg����X-=!up��jʗ'�H!xѨ�Գ2@��9��Ɨ>���ޡi7��O�����n�F�L2K4�:�G�&{���~ �34m0�剆<v'Q�����[��ޢ��V%	߾����6]���K�Z���eXOE0�󌆩�����Л|
R��K�6��t�N��9�uC2��H���N�R���j��TA�s���;�pSЏO�Et�J/	�_�%`~�YV�6�Ew�y�\����r�Þ��im[-
�״N�N�Ю����:Зச)[���n�L�����2n��,i*�;EX��Nj�h\c_���N'\���x����	7�J�F+��W���0hL�U�MW;Y�{��q��+�(�cn�¾�r�a�<� 6�2#r^����{��_��7���A4C(�셌��v\Ա�_�r�r-J��r�0}�}�R�䇼���ݤ�2I�R�^�N���1�N4����T^>4���M/jN&Tq�kQЙS���^0.gQ�wF�CN?Z�D)ܓ�s ��L$B�w�w�g�FzR��e���A�r<6�W�@OJ�Tj��s�����j|�x�%�>/��7���O�6���k#�8��]4�6cd����R7��h�B���gX��fr���E�!Ao�kh\�k��iuPҖ�g�ߵ騯�T����n�����/�+�GPv�ļ9����ȑ�yRŝ��O|��kT�{�Fj" �;w�#��zЊڴ�c�/t\��5���I�^�g�ʝ>��*�k�ͩg*'�E��ǒE0��s����v�%�� .{�SC񦳊��v�+�6q���R}�X���������$!?�tqOל��M@�����`��r�����wß�TX���8g�(�@`�|n�5<S�A�yܖ���r]q	�7c���1*� ���b�=�e�>{���̾�Z�ïg6��׌���>�Jd�"�T<S:;����C�H����oy]�6y,��v�P�҅��1��kU��QOE ���l���v��=6�{f�zS8F���$��{t���R����0���^�LTtk!��)!�%ECG���y���[��K�^�L��˖~U�}Ⱥ+�j�*_��1�Jd:��AƠ��#qf� ���xf��&ѝ���ݲl�Rgg�Bn�}�r
�����nKb���1�C�^�U�� ]��F"��yQ�%�[!WpƬ��b�=���0L+�~���{ pRU��?B�n-4G�h�4W1êk�[])ڎ��>�n���;��c��QU��U �ΪL�z�̴�U$�5U(�J�в=�V_4Q�up\�ƌ�AŜ�I&���ϗ��^����E�z@e�� �\� ��D�^=�.{���ݭ���/��tpt�Bﴔ����E7�t����ދ�b�!H=+���&ݬ�:�u��l���U�@�f���'��U}�vS��Qĝ|܋��k�衇��Q�>&Kᚗi�h���$i��2��<M\����t��@�0e#MC����cB��X\�LP�>�	���!$�6�=���8��P��Kp'NU�\Ǿ���)"x֭���_��)@RP�-J93,�q$�d�S6ð<SFӶ��T2Z����,�-%��`�݂��N�T��~͖��ȃ-E�F�v[�eS"1��^>c�J��}o�[�M����H��*jU�,�èD؎�i��o��~U����)]��]�q�������ǧMu��ۣct���u\�p���v�s���ҏ�X����t"�5<������;A
�s��[�_�\jH�,jd��A�tfsս+R�w(u�:������x .L	�æ�OԌ���_~�H-��%F���5��<gW�X5��l�)�+���f�җP��N����b��OVk�X5�	��)�f'KTӾ\.ѿJ_S��r�i�*y1�X���P�9���c@��*_j�˛���s�͎��n	�԰
W��c��I4�2�J�}�oxh�Q�L����B!#��[�*���]����+�`0�{����&������A��Ӡ��O���<�B�!a�O��%��5y8�CIgS���#[�TQ�Ū6�}��^L]G�G����t�݌]�}����t�̼=<[�.O:.ґ\�ȴ̧\��˫r~�W�o����x�O����Hu���G����<�vX>{|�OͻG>ð�x���*H'��'-`���=7%�X��
���j���|=`��U@���<�ۑ(�?j��Y7�R�Zk�{��;�O�qk��Gy�;JH���#IA=����`��c�Q2��	�L�a�"�tl:HsM$��{*I����bQ��Fv�]���KJ�9�% �"'͗��x��;��X�ݥC�~!,��s��-xlo�G[�_n�GS[f3~�R�bD��7��GV��h�;;n��)�W���'5vA~�M��S;�i2�|�uv�`Kl�?#�R��f�%Y�v�����Z���Gy,��W���O���Q��R1��i��ṛ�.KDL�7^�T3�vQ�`"�FR�'��.+!��F��$rQ�'vG���(�܇HKPa���>�.I�E���Z@��a�H
��"g�$��d��dv���h=x�W�j�e��?	B�� ���Z�ң[�^�J�c:G�c\Ҹ4/�s�����@�q�a�e�Ƣ܍�B��}�|�z􄷦�"�aU����*~Z���P��
ɢ$׫>;/p�~��������G�Q;���] �UN�5�A}�-p,;��}j�k4>�=0�HCt�R���88��;^"t=�Kp�����3�ϔ���.aS<}��N�<L�g�E˚��/�uo0[��v���l��{�
�k�',3s[�|�ꭊϚm��~o.�S�Tv����sT�נ�݋�k�;%z��eJ�����q ��%�I�M �	аgV�^�}ݟb�}���I?:�����k~��z#o���r�a>ڶ����g���v}9/A��k<׉{@�#��a?�ۇ�t�E��[i���y�&<�ǽ���J�=>Q�&c�Uˣ��jb$�\�6�k;^��)H�D�U��|�s�/&\\z&�?��q@���y�]`ֻɍ�(~��W�x�k�rsX�I�&��/�|Ur�a�;�w�D6̭��A9R�"h�$�L�.�)�#����1!w������%�<��l��}� �^�3�@JH���_t�����έ���=���Evfs��++�"	�v	X��(�zn���/�-#*�Sbd?͊p�S�*��?����سD���2��:�H���N�D����P��7+��{�N��'>��%�ԋ��3*U��
L\V*���������GW�}�M��vV�ȝ�FN��"��u__u���DcpťE��C:«u�� �E�k�q������j�4%䆝��kFy��z���;I�Zh�n�Y3S�7j�{h�\��\�_�b�"o]V9c�.�m��k�j�+@G���V�zq�pz-�Nw�M^αn�7e�<�Q���|�3��G�4V�IᏱs��/X��׬�d��g�^�S����L$�C�):��t��$:�#�g1_���-�� q��P�c]�G_���(��83�O�^L��6*OK#�
�%�>A	��:��i��~�IϯB�\1
�1��汋����e�gS2�z��ǽ���ο�~?vl�Q��*l��j|�w�k�I?M�ܟ��uK�����*<�+�
�'�?C�/T<Z�I{L|�S��,��a�p今v�$fx5�4��?�:>���֚ �rX�M�t�O`��&[p1��8�=?�Z0cIa�6�'�J2��
��T�+���_C@�%6wbV���#���/kՓЬ$y}R��qǻ*L��.O ��c�,�vR�囑}��7z9B>%lo�~h�rA�*K��:^ �}��1+�iq��z�<��nC�>J������㗖��n�S�ʢ�9M�訵'L`BI�M"��&s��'�gqf4��8_ؤ��H54��_i[��]s��M2p �6n:�����㾯�,�kl'7+�q��Ѥ���S��ؙ���ԼU��]�)Y�Es3�n��z}PJ�
��d�]���\DmKQ��X/���[Rn܈�T_���]\��l�ޛSTq*#g)D?͍�j#�98#�8��@é)ІA�q��8�w$y�=M%Z�JԳN��br��"��3�sنX̘��[G��G�>74���s���e�����%.�R���ySg��v���e���u��(��\)9�#�rl,̨\�Q��41�Q��Ӽ���ul�[0�V/jw#V��& +{�$���7����(}W��ꨩtS(�?��ѕ�WZFT�����?��@�+9v�/ �_�˛ai�.Pa~�Ӌl_6!�l/�c�Ɍ�G�)��+��Z&o���Ίh3��� ��G(��Ѫ���?ѓ��z7�½��@ɦӾ�����9��I��@��&��L�w��M2K�l��:jO?� M����>��k���ߞ�B ��U�.�5Gt�c�n�|�K�6<]����[��QĞ�1@��K���L���H(�!�C 9���(:��� ���y2��A����T�m��k3F!�+�h��v�Ix"5��+�(��Ӯ���ݼ�J:���q�D����Bޡ��S{_6��s4}<̜6�6^x�VQ�n�`�%����1������Ix�d3]���٭�֮���l	Z��r]U�H8+s�����u�z37	&nJ��<�y��t��<a�I����\buWG[�fo�LG�|���(��I"��"� ?��T,=����s�0;����<��Z�c�BU��A���z<k��7[?�۲�����j����;��]�]� &*�L%�SC8�<U�"x�3���7@���R�9S�\>0h�/~��EP���ӡ��a+�kH8�J	$�t��g	����ߺK���>V�$�%��������&��$@���-�Ê�֚�H��8zȘi<V����H�"HE|�O�]�IIB���Ș�#td?	��x��!3�S������KX1�}7��Wj���c�A4���@��0g�OJ��#Wf@��㔆��z��T��g-�����Umћҫ�UV��1��E����g�2�\ˑ �@�A�2�|���'.V��ҴQ�+����j�+Er���"R�>�X�(�,�������+� Y�,�	`P	� ���4s��
�k&?eqV�P�邕c�� ��L>t����Aǃ�\A�-�lX8���8 ���7��Po�B����,�g`e�����-�Q�XAL( ����x'h&X`H������|�=��������[���q �PpAi@o�f�,���6���+�X+ ���`���!G`U0��N�r	��	��	`P	� �@k�}���^�8�y�;��-�k��8@����`߂��hXA��������b�>�s0a�*]
�Q�XAL( ����x'h&X�I� ����B��z���q��wp[�!���xo@��YB���������������0���Y
8+�)� Bv�O�M�K�L	 �8�G@k�}���^�8�y�;��-�k��8@����`߂��hXA����������0���Y
8+�)� Bv�O�M�r��� � w�f~n��>���Aǃ�\A�-�lX8���8 ���7��Po�B�{-���,�g`e�����-�Q�XAL(�����x'h&X`H���t���ax����. ���C� ��ZB��Y�~(7���J�鷹re�#�gLQ�to�[���+7xn>9<} �(��\L R$~�-C��>E��y�C�e�.��� o�T~��Z|O�:�u0�i���g>:��$ ulv��ۦO|u<O��̭j㡷�;ɞ�߃�%M��i�fN��.��e��9��Xt�H3)��
��W���������2&��3�<��(�I�8�%
�x:�p���:���b*k&�Tg�'i����eaahv.�G��\�����=ij
�⅚�MWʕ��/T�{�U��-R�����Y8��r��X����?IG�j���/^�z-X�IH,ɺSW֗�U%�Q?6����x8�.8�J%J+Ti�U�E��y1��mx�E�����.L$��ު2n��������TS���4d��O��I=�1ٌ�$ά0���S���6�o�D�b@L�"���c�jT��\��R�#��,�0D���w�U`�<��>yuv��vn{��^��T&��R�m�U?a�"C��E`�KC>j��g��.��
p�a޼ufE���5��k���aه6m\u}����3�C�'��l���}F���0!mލW+R������aM	��"oQ�]������o�'d(7���D��I�ѳ� Y�@�K6���+�X+ ����1�/PZ����)���o���.`/a|���̅��/��惛`��ra��=�{������@�^���\��-�p�q�r�<��.�v<9 �B� �`��� ��lhqAŅ�=�q�ƅ�=�{0����
08�=�q���É�,�� ���=hzഇ�Cׇ{ �!��xoa��,��C};Y��t$e�EX䙀ol�	(�˵FF��4������&|h���{��7�j	��;�	�ު���x��.���mFX��ꕝ��	7����u]�ބ�U_?���$�=~%h\m��{�"�Ҵ4�%����G^/����%g����p�����u�����_0���	����cR)U���-(z��y=iab�1�Y�r�⣾tM@>����5<;C���p7���Gf]&4'��o[(����z�n���U�Z��5 謤,.2V7J�kM�����}���ߜy����.C;�ig*:�6I�����VXf��-6C��U��#=Y��Yo�u�������\yT~�v?�������p�@0�Q���Wm���ue+��U���FK}蚀wVr���U�+^x���G2��3X��b��c�3��}�9�f�֫Lf�vM
]��?��h K(�Zc������get����N��z����OZFX���q�g{�3q �r��|�l3��z�;Z��]�JC$W&]b��-�J���$���q � s�_(���Pk}���s�}�y���!򞻖�(�P��Y�Z�VY*�I+�\�?�rhF{A�	�QR�K~QƁ��L�f���.��&>%YG���Vh��yy�?�e��
��0[q���N��;�F���ਏ���\@�Ƀۃ���D �F��\��N���
���,{5�j�w��6�C��pd��p�I��o�Y���H�&l�z�6H�U�"b�&�^� ۃMX�Qww�TٚZ+ui�vX��7.T�VU��$����f�t�������7��ãm�d#���H�൴RϹ�TP]��lF�؇y�dG�C>yZS.�y9��O�k�>s�k��_9�b����+~��yS��l�»K��1!e��-�_\��T���L�nffhc�!����C���ź��>|�R��ha�a�����r��aEs�oT�����\.��1�5+`�����������&����wq��/k����9^^�g1��a#�V��,JU���7	�i� ��8�1�F��$e���ɣ�f��[�c�cߤgWJ�����c�Tc�]v����b�
�k���+�m�1��-�q�U��Ä"�ђ�V]���.�O�we�: ]\������$�E�������:�<��/#���ye�hv"���<�\S�'| �r�#R*��W��H�f
%��S�O%��
oŧ!���.��"�\�����U˲��⳦�W��&~T��'+�ޣ3�P����X���3ωU�;�At�`�їFE�'J΁o��ă�|nTcC]�S|�{b�q,sѰ�2Ǖ]9���6�{!Qʚ�-��au^T��1wp�rY��v�Mo�fg���
���մN���-h��״7����3�P��ce)#�����Cu2)w;��ƴp�a������V�&�5�!'�N�"�cwd>���%X����/��m����G)"V��>�!y���
"���ѳ�����҃����G�ʙ�C�ׅ��4<�P��V_c\�;���4A�p;� ���Y��6���8��	��ey�{��7��OPԮ�y���Yz�|��*�����sW�0c]�Z��m��b�V"ح�L>v�YvD������lyHn�|u&bˑW��wk�h7M�vL�j�{��)��������q�pN��ۖ/Y����#��.�}��1z�.)�"wŴ7����k���ǌ���#�,Γ G�����2�9�H4���Ӈ�I�?���P�|��DM|[ɔ\��+]��c�aL��A?ַ��c���7b�ĵy8���3��rSc��y�f�����'���@9��qN�+�� ���r��Mo�!��OZ���i�m�)��;~ʚg��,j�H��㌪�d���rw���C�[P�8�����wI��	�J�:�<�ӛQ5��\`R���:Z����������|�+Pb�s�*�P{ũFur2E�I���?0��^�)[W���\-퇶�.�d�]�9n_U����Ӄu����}MO1+WPc�	P��H7<�Qa!$5CA6LDZ�`&�1)�)ˢ��	�6ف�2��P����-ݝ<��<��.Q�!15A!)ʝt5w��~�`�Uv��"��A���������l"�!9NAϐr�j�������Ǹ}��N8T�v��ޟ���/�f[[ ��~��w%9��I��q�|%�\��q_Fy�%�P�1	U>c�q:��$7ES��Lع�j��q���*����)YF ��^kEF��*����1}9w (]���x��˫^ \��Δ&yh��p%�w���}�,>rUK��J,NG[�J&q��_O��γH��	�O��)P����:��pŒ�[���;������#8v?\~h��t��4�x�����|����?��k������uX6;�ҫF~-o���B�",lt��k�J���"��Q7ٻ��0F�����2�G�:	�_8���]j֍u��n_|�uÃѲF��m���f��U�g�R�I4��7���j_q����T2�2u#���g�Y�"r��A����Q�������C�L�}V�2����6Ř��\�S;V-��1{��T��Yc{:k��L��0�y�l�r�5��ɾi5���r}淝W#��㓖�KvE`o�g���&��V<�2����-������O�a��Ő�������a^��~=<�=��<"ϭ��e�s�U�P�����;����}Z��n�%�����w2\)s�Pp[V�k��Za?4�p~�����L�&�x��z���wv��'s��w�/��ƽ�Ks���r��T@�-bZ�/�0���h����j�\("��!x�(�JD �3$F"�T�_� $H
��P�.Svmӻ;�"ݻM�mB`�8�����J�5m�*Z�{y��$���t�v���.ǁ�{[f qE�l�ap��z����_�.�8B�mǥ�}��U�I����{�{{�����j8]��_��~������)�k����F����T\�����L���~=�{l5��ۃ��4�R/�r��I�E���i�� ��/����W��-�+�%��{����^YPKү��!n�Z����6�N^vqe�pgM�ؐ���g>Ya�\��i�,\�L�y�zP�gD\�kHqd����Y���
H%�����PY����u�cΦ=]�g i��H'�qP�iꘚE�M�@�M�r�}��F�&����y��"z4G�:�l��W�~�{�_ȝq���_7�@	�I��fR"���<e�=a�Vl]�Y�+�����P\�Z>u9�/��u
Ɋ,Qs9�/�����^����t��h��v_��*��M��� 05�r�{�PyW�"K/V�l桡|��Ä����Za�Z���S�2�p4i�{c�ww�e�i(����� �^|Ҷ�pb���mH+�������̧�.�:��*��ay�*A��U�Lξ%����Bnt�g�	�B�yL����dU��2��{Y�o�]�e��]����_�2�Q撑��'�mg$�%�_<�OKS��ƅ� xi�T0k�ȟ�2��^���S��׼�t��i�5��#>ڃ��`C�}ڈ��J,E��'{����	KnGO	'�X(�Ys�=���bl��.Q���,���2�Km�'����������1� vY���d�q����^0�$;4.�ĸҍ �y�i@���д��H)�EUB��G��@b�:l����v:��+3�d��h�8��o�E��2T-*9Ɖe���~x\�y7�`},ٴ�X귉J����h�M��X^E�_%��/S��fh]�:ﾆ��9ԕw�z�S'��(Մh��ߛ�K�#i�R�~�)�9��ycR
'�,L���}�q�Pd�K^-v-c����k��4��,;�����9���ǲy��^�[:��=��¡�A^2S䫥N��&
Q���:+�h4d�HaM͸z�CRv"����(�Up{sپ���-�I��5�"3IO`x@������z^���w���k��쁻�����	��Ӧe���-;n.��&��{z\��N��n!�D����d&�&����d"|C�U��[�n�	�=��(Z�m%�Q�&���\����&4Z�����d�l����w .ڿ�w��+q{�	��n���~�*���Ϸ��'�yC�~>S��q���*�%�]%e�w+x��и�Y�l@$v��|w�/�x���� l�p�-�-1��,��|{���Y�I;� Q�w��͛>$7���������c�R̷��t�wڌ�I\G�.+3_�Rچ��G���-Q;a'��Ɲ,�'Q����x`0�bܳ��K7
�T, �UQ�@N�FpL�νT�m-y��t��7U���Ab�(+�n�C�Ik�����sr��%���XN�]������t����5	�F�_Y7�J�t��N��/bm�:M\�UgN٩6�gF�����(b�#��[v�w��5D�-$��zJ��v@�M�~����R�o;��ˠ?0P�̷��'�˦o��1<s{OD�_��d�;؛���R]�j��.�}��%g����*bn�%�B��ڗT�Y)ƛ�����+ۦD����҇���u���Ҩ�U�c��\i ���w1;331-��߸6.�T��Ǯ���Ո�V^2�H��Ko��p
m+���1��P�b���KgzF��o��qF|!k�a�M���{����:���X~����ٽ��
]sGU�sA��-�q�[2�y�k����pD�tMA�;&]��@�4`Cx�j��|О�ViQ'/�fM&�89�<_f�Ӝ�V������e�>¶6�`1H�*�q"�BIFж�fIՕ�HIқ˟�-s8��n�.���O�E��+}�6�����a��0W�sP��O���U7��7[~)���H��f�����w-`<�����(6O��b���{��u5�Sؓ.q�9���	g���Ҏ�����bnγMey��	&��8IWе"@=e$�K��.g����	
d�ا�����V:Um�p��u���p��̲�璻�L�/�hP��aVC��n�`��[I�X����2���J��������	��pE����U8uOf�f��'�X��\'�U����r�@GU�27�t���ḾE��j7�( S\x>��+B�_�L��!g��D�$�HE��%���$��}ZiLF������+�^kk��ˌq=�Փe)Y)�����xN�HE%Zq�ӽ��8�����P�����l���n��:�m��[��Ph�LgB+2U8^WV��M���ױ�����+������%n��&<��^958V��S�o;��غT�ײ����ʟ2��Q��Gj�M�D8��:|0��
t���g���������×U��6��y�]��ӨBU�K��h�����1��h�Kn�1�:�� Rg�c��j�)U�]n����Rd�����q���T�(LN��`nC*v�W/�#1)wËlR�u���d�d��6.u�C×�X� �P���-U�wN��NE�N��	�>"Ѫah!�z4i�*`n�fн<�+י��Ӆ�W�$���&L���V�.�$7��L���Kv8ל�.�o.@��U�6�?.䦣i�/2Y&I|_w�kzϠ�;��p����9��h�ĵ*��݅�,��g蒞�V�3C?�#ZTY(�L�g����]�}A&�P>�)��긑74VْϨ>���B���S�&R�egy�������P��]j|�ubM���Ӆ�F�Q�g�[Er��:e&��9�!���Z��J�Lؠ[*�L�Ϡ"�(ӽs�`&�{Ql�.�Fؕ�)��5a_�@��(�ɾ�ԋ�R=X-�xÄ�Z�A�>��9Q;��3�����{�X�^<M��'�$����e[E�޸��ǒ ���*�K���q��h}�c)sL�U��z5�j��me�-��!��Z���(���W�����vª�]��Q^��R^�qIŭ0�Iԣ[2�p|����nx3�'�Y�gk����� ����wg_�v�H�B�,(�*<%�s�b���.���ꅕY��U
��qb����^�\���fRPd� �~��A����!3����f���������7��o��q"WyW���i�������-���L}�hm�h?�Ux�XZI}��0���Df�<�G�%��N�ꒉ��j1+2;ʶ[if�v���GS�*�w\�<�9	����aF�L�O2��v�}��ȧ(d�*��^\~�B�� Ң�����n_`�k��@�ⅷ����$<Hw��
�}ذ��&F��jA%�P��)4�̇}~���l� ���Cs%�EP8dp����}}�����t��Z�iQ q8w���w�(зj�SP��Q
}�� Z4Zb?4yg^Q�Qv�U�=F��9��4�;�sX�-h�-�N�ú�w(Z�]ml�~���O0l����V��^2��@��I���{����w#��tߌ�\��4p�X���)���-.��4�
������]?:<��*��V�,���,��8��nn��1���wW%l��q�ۯ��PW��I7X#`J6k4�7 �����B��gJ/��c8��qQIh,�O���A�"�Uf���z�*�R["�n�E�o�E;�m���:M�m�W}�[W̆J��󆉊�K��n�5����ݚ7[� �)�U9.���G\��	�>z�9��כ4ˏt S(�*�֛�g%�_�f�����jL�5�L�ϴ�E���)���.��7c��ii���`���̭-�ݭ�t�MW�dF��	ᦪ�E�L��S�RctÆ�q�Lt�ϟU������J�uOa�y����FU/7dø]���UG0�2n�$��b�$R�x^f+np*���7����Vr��Z���pЪ[��i��,a�s��O
ը�V�hff1i�(����~vgnN�S�V�8�q`n=�&�}Qf�����ٵ����s��g6���fv��w�G��dz��c�x1�ڷ���v5ǭ2ʃƍA��I�V����O��7�Vt��xef��V#{�}��� ���j�d3����q(���s��Z�U���,�N�wJt1�Z��m�)�4�7�Vj� �S�@�:vmǪNJ�ڻQF6p`�h�Ƃ~$W����x'r����Y]W��i��� )&��2��7�첥q�6LK�g����}�c����+3Ȃ�!�X�O)6�+���&�o�9f�@��3W�`k�*|5��ʹ�7��� ����3�����h`eF�X�j������;�����a�K�:g��d��um�ƭG�R�@>�~���nĠ��Y��'.�{�h�vz���)Ap%��OB\gDh�� ��֗�yM�ˇ4Μ���`9�pk��r�i��kcq����&�-E�L%d�C\�>v1���y�6b��o�	\3��qY.���pP���#\�~�	�w:Scr��TSb���:	��;�ʄw*/\��2t+�����������갖T�^�0a����:�\$����F�Y���]\���2�ظ �Na��.&
~ɍ�6Bb�:dHFF�k�ن�F�,��n$=1���+����^�E}kB?�sr�չ�-Ys��3�o.U�^K{�P���^�]��ze6�|`�����#?1� EpP���N� �`b1'q�I�I��"mx6!�0�>�9��D�����������-�=�<p�G26�����)rw�TP�7e��U��R�*���E�F_��ea����,/�ؚ}�b�gɕJ#��ǂ���L�r�T�>�(<�6�`��q�~��}R'5�h�R��}m��r�ǅq=X���Y�������j)W���f#���R�"���
���Ǽ���&jڙ��!Ve*\l��*��	���=�=x�d-��ꉢ6Q	�AN�Վ���ory^Β�A#�/&[�7��f8���e��omC�����38�2z��[�+9wDs�I}:9�AU��" D[�>�BQ/R�Ghs�m���|��u;6#?~hQE�`]�� ����\otie[E��e�=�)�;���&EW���8
l� ��f%p�Sۆ��3#L�X,��h�e*_zTJ���(q�L�e}��@���"�`q���e�i�[�e�g��]5w�@(�|X��	��NU�һ�8���EW��M������ϰ�g@`�27�.
E�S�dx��!�|��/?�� m�"����\���I�����ك�e,f$�!�۫�,O,�KTj��o�)���F��~o=̀K��fi���"�:+)�}e"�BTZ�b���������Y�eZ��T�T:�y�� ��0��p]�<e5��悱;�i��^QC}F��IH`�ξ%JZ��c�Q*"�*��G�k��R���A(���.dJ�3�������HA^�E&L�i �6%&��д�'������\�W�e�,>z�ak�SM����Jn�˧�/�$��`�3��#¶Y���dk^�v�"�Pϼ7��
}m�I�1vxXI"X"��v�E��꿊(��IHz��!��L(<�$RAd�a���&Ȇ���閩DȞ��\&�(�휠�40�*�Bׯh��	%ǂ��;�LԪ�|Zw��k|��o|3ڨ�u�IG��+y�2��&�����aR�&#-�L���ێ�t��<�$���"��F"��,0t/�M�nl�I)0+x����)C�4k�<;����:��޶��x��A����,�R�7�����c�3�e��� ���L:�z����󋞖��,.�>�o�y���tq˰,�-�;�W��%�5�D^��PcJt�uf!bJ�/���9t?~����'��)�����������p��n�u^���ղ���`U-u�_Ĺ�.&e�k>�ff��͝�P2�@���բ��s�m���Oo�Y�e�)~���3#L|FA9�Ec0U[(��Ǉ�%��`��ukh�E��z�y���k�;���W�ʣ��J��9�i��W�6�(!l�}:ê��(�����FG�d�l���3
�U\�U.��IHO�C����l���{��䯁�Q�(j��2�e-�ПQy�ʍ��M��w��h�K����sCLQX~G�)�>��g�3�ʎ�`�­���L��a�lw�hi99�ǆ�O	m�u��.�?���PZf�������p(�����H�I�Y��S�e �D�Rl���̡V��L����7>ψ��@|�-T�U��?��jF�<a�uɼ�/G�
�fP�u=HV�?6@$fu�ə�;"�Y?�>��U�<s>�#H�E;P��ƌn92LFS3�� �d��	���F[�O��8�Ą�o8�i��i�D�
�����!	1q]09x�)� ����~#���2\%�k%JƷ[팉����g�9��`Ώ�f,�F�3���-�V7�W�U+��e �c`6r'�#� �>�h�Z��@�^�$����X��iTQQ�գ{L��c��-9G��/S9�kf���b6��)���%�;��� F9'�@yu{~�E�6Qɱ��^�^^�f�޺�i�΀C��ɹ��
̜ԓ����Uk(�E�@}�?;��6�(ct�Lmu��A�2��5T����0H|��+��E^�+u�G��E�ͪ�=?���s.c�:�� �3M=�������{�P�M�Vj�S�8�YP�).��4����V@�r�# ,*X�w�r��<�PGB�D���60ҫ-/��U�_Y>�x7bTeɚر����yѭ&`�u-{lG�����3�D'#:�����r>�A�T�֨��1v���&*](0�!quj����� �N�<y����º�u��<�[�)���$۲�a 있q����4��Us�+����1��9)В�#���1�6����e�G4|أ-wյ1r
�^\�tQ{�%���}؟�2JV���-*f1�;��DS)����%��� ?Ф\�:���QR���D^Q4'�%��v��M��% t�u�&'8��UK���S~���bK�a��n]�5Q2hۧ��N���C���Av+L_Zq�ϋD����``ˏM�y�zk*�8-�o|�nd���l��s�c�)�n�'q,fa��	{����$��c�϶Wp�m����}���?�>����a���F����RDJ�����cn�=����~�L�3����}��RA�QZ�Jzm���Z�S`���Te�h+�ƿ�vp�d�_��x��ꕰ���M���$'����e<
���y��-�X��yh�Y���Gd ��v��R�$���b��i�����Ѳg�v�~�~��~�T���7j�5q��cii�����|����ωɘs�3�3�Y�
����H�'�v8��x�Q��5�_��W���z� �w�����o}�F�TL�l�;'�5�77����SS����<Y���%"�O�/OCO�s�H��U�|�X�'�	��2u��[)YTdY���П�h���,��@X7�>�	�(�ִ�]�o��`�|�D�&�5�v|Y}�s���w�~ۃ_~���#�;i���˨�vf�|�����Qr>Hx�]�����$І+��,����O�t�]<��ew�Z�-]HC]E��:���ޗA�(�!��Se����l)ro�H�T����#�!--�-Y�N�Q�r>u���k-���"Q_mJ��t�}��&F�H�+��T���8�H�Ԗ"$��wu)E�[>K��|� �P�nԧ��	��޵����C���5���l@��
��QO{���ڵ�}E�0X���5fPٞ+[^�m�����7��p���:��ހ�y���$?�?�'��ܱ˳���J��䯠��z�꽶n��+��@����\�Q�85 ����Vi��3T��:�հ�����G/UGިA��� �C�D4p�!�u�|k�*�p��j{A��~v��MTO&�l�S�����@%�/k���L���F�P��ĠEO�A�3Tڳ����g�?"�� D��n�rW�3CK@�8�Vw�0j���1ڞ����� ���DH��a�\i���+�'b��4>�Λ�΢�ތK-��a?��C����7� �'�O�´��[�H������E�bZMn�������Vs1�^���A�C'�kp2����Uw�+o ~HfƤj7��5p�zj�i�,�Oo���(���C 6J����%��
��q��Q��V�G"N�aE�ĢO��ϺE�-�}gb�_�"��O��=8�CN念��Q͂���:�Q��ۄOs.i,�Q�}�͉���\4�&��r�V��M��^�Ε��×_;���+��K,^��{;��'�$:��s��_���u3�A�S�I���zf����?5�b�T�!�m|�ԙZ�T��uG�Hn�v��3�0�[�H�^���*�f5����j!���̊M�b-�O��+�zng�w4v6�b�����-E���0� V������J���OqB�6��@�4��8�����C�,9���E���T}�ݹt맒���V�ɤ���O�l�,���ի�>ȓ�ir��*m�5����p��6�IHp�eM���G1EVO�S9�����)�Z�D�^x��$�>_�i+�u�~��N�&KHf���h��t���A��?߿\�W����!�K�i!����dѭX��
\�H@�AS}�. �� ��^O�6��&�IL���*QIyԭfq�� ��WݢĲƴ�(�B~xC���^�M�2�DpF�c��o2��DȤ�ٱ�ֵ�/��sZ���i�����7��jR���N��a�s�}�֓�~�Ұ�?*����q/{��K����W�9l"B�:x�]VG�����5/u��&�}3E��%5~�n������y�e�x�������%��2�|v�=�P��(F_�)D��3�G�Df��U�WR�'i=��A�F�ߨ,j#o�������T��Jb���O�G%�D��c�T�u��Ԏ����n�m��͟��jf����j���t��_d�F���r��X�����p�{�6�p*}D��ʗ�^��~'���Ą�O���?j��eA�C+�ߋ�s�&��/dG2+3,�U.��m�9ec�}�?Ε1|-d��A`���.b�sLG��Vj�����A�����.I<��e����bw/�8�cj^ Z���#��P*��-@�C݄�ݝn�[aw��Ѫ��(�4ہ=�]Y֚/�f�ũ/�,ژ�ѸL�R>R{���s�1��u�N�fB��i~�AA�k��ݶ�'_)2O_M�(�X03��R��M��s/�C�!xX��L�(Sp����:���_�5D��q��F�4�	�d�i���V)h�� -+G`cۢ�ϡ�a\�ٟˑ$�4]uAaE���nS�ihm�+��^�U�qFl"����Kf19
��CE��P:$���0���%X����
��So-<�b�2y�U�O�^?�c�Oq���ߎQ��Y���K�4q���[.�\�Eq`ܡɺ`�,n$]�>�^��~/����le��?5)w�wξ����P�]�
����Q�׽�f�,0��P����J��D0W�'hD�]��q�+C���!�z���&�q8�B�/�ʇ�F[�Ʒ2�bYm]2����cd[��q�<�\1#2����[�Դ��JX���K2���+
�xWG��F\����!��_ZKƢra����a95��Wk�)>m\�:�L���v�T��.���
��=Xv,�����P�IZ�5�-1�s�̷$@o��Vz�ھ��Pa�����~d,�̼{"e����?��\[H3����2C��PvL�:"޺��/?ٳ��Q>r��q�
7��5!���2M�/Hú`��n��Q��~��Hfi0�r!B�N�wk����0^����ԸY��B�g �p'E�u��<�c~���
?���>��fAÅD��{G�K�:h.�j�z�"z��ޢ��>�#�)��#�C
�/�.�����~	�5��ׁ�w-Յ�����P��/w1m�>�B�a8�Df��/�Fgj���R�Tj�(\��?|&��R�Q���o����U���k���_���Or���)o��a7iM���'�wQ4m��9H#�}�(N��+�n�*)�c�X�HNԠ=�������f�˪���3�Zz����VR�Q���~�yh+� ��Gflt8tdm�߳��*�$oVD�8��?������E��뾦M^�9"��>��?�w�)�ޘa�ۺ jC��`;nxh{i��3c����3����}J�[}���"0������*�,���Y��@M���`K�e���mbw�t�o�?
D=D�s�T�x}T�&��m�wN��|fIxz�{3���� 5Z΄�6�38�\Z��U�ed�b.%��fcy�C�(c ��5�A�k����)�H#b��->#��W���Ϥ���bԦ�YvE����M-[>P����w�{�r89����$�v��1��� ��fYjv&��<Ӏ�B�7)�Qu)����?�����}͈��!e�gv��w=�u�C�UGy����}d%[��.�~�R^��=����C=����J������34:�H���wr�.�R�J�sU��w�������JD�{��ϳ�Vs��CMwN&��TK��7�m��s����M��i��c��>�O� 򌦲���n!�_y2��=Y$-ȱ�`Q!�bqW0�̃̀Jp�"ת�7�"<��Cǜ�ɬx�[s򽎻ʁIÜ��1���F��Y@�<U��/��?B�BU��fWe}����e�/zfp���i��O��rc�DP���� �t�-���#�n�Y�A��	6�B�������w;G�K�8�������+��FR�{m�;�n�2IB���V��̚����#Ь���!c�`lF�RX.��~�y�Tŕ.� Z��w��Nj���t�T�p2"�_g��K��H4˃,��	#J�n.�����3��!�C�$�� +�Y�r�@���x�tn�'a�Do��E�	��܎јI�Dl�y�#��M�&OՒl���F; �%��c�x��r		c$�-ʄQg'�bW=��#au�R锲	��*�]��\�]�Q{G�t�{��\��R�>�A�D��� ���sC%�!G*�6���*��$�u��+f*'SV��H\$i�?C�MȤl����`�D��&<�o���ɎGE��7hˎz�d��47��ɟ'��a��kو�}-f�W$/��c�'P?���
B�^7��p,��o�Ɣ�m�+.Y��I�&f�YM�e`xcf(cp���&��m�6�����n�[�:g�вM�-f^�PI�Ņt)��Q"1��G�=U��Lkr���w��ۿ�����ϧ��_'��4m�۾p���&��tKzl��1?o�"�8F���#7�(�)WP�@鸀`��q��翟>��١�7��Ͽo�?���?zv��ϱ�c��ۭ�2H2%� �Fz����*D�	uΘ*ƍ/�"t>F�P-�ʆ2�Qq^�hu�V�JG�	U�UB�s�\U8	,��%]��
��[`�����!��^&4���̓w�7ԙ�2�+�c��"߿�$�ԃ�I�DE/!^�H/6%i�^U�F�!��'/��P"�A$�d�x�*e�Կ�(
QȀ_C.J�5��'�%���ę{=TbF蕔	dK쑞Yx�R�$�Թh�[4��^�	Q��W�,����u�ͺ�W��
��r���h	ܵ`�P,/R���P#���h)ċ��VL@�$kC�̇��-ʖ��3w�XE���S��^ �+[]�h"��sb>�7.��=���B@BHBPD\"2X�d����Vl�J,��Cu���s��T�8�ңa0����/R��uv_\3H�x{��{
: в�r�����9d�|��<p�Q;� �J�LX�\_������n�y�w���=�Θ�R'��c�f�FDb�rE��$��Nt�ni(6��}0"t���d�\����K�e�Dӂw��%Q�a�����0�|0?J0��K7��|�>rz�oaC���,�Us��)�'�L8��q���|ȕi��S� �� h�]摋7�=��>���g�g�_���D"�q����3��Jp�Z�t�B<�%�]������jb�m�	�MqL��;��i_[�����P8���D�I:����N�V�VULT�TF��Fq���R�gV��p2��e�Mڤxw��Y����L6E� �@�_W*���Zo#f2�Ⱦ ��*��1��PLm��Z\	���f�2��J`IP� M&PH	��)�;�L���Z�1b����X��AR	�1S�o�3v"P�W�gLT"ˁ3�%��P���	�b��(Bb�!(&�W���iH��1��6u��u~�E�\�NG}+d*�"��ؓԶ&(	o���u��/h~�]9{"�� �)��@bM�O�Ǥ��|�V�9YkV�1����R�g �?y���/hm����m��|�L����0�
&��ؕ���p�ȃ�Ry��=���6�d�[@+���Ѱ#GDh}���҅� jT��T���;t��M��:H�SROh5~:��Vޒ�dJ߇[���*	]�}�a)R��,�h W聧��"�P��&�?l�[��W�&��=�L��%+��$JҦ'L�WS������{不�[ � ���
� �5������Ƚ�ƍV��"ƈ"�1w��<�l��;�DH�������z�J�lTQ>]�m�y8�fmݓ&#����D�����p���\�|̃T9�(q��p�H��(��-�o����姡�=�A�WH����K��{ݜ��>�x�x���pV����]L��� �+*� �T��
p��7���'_69�yN��P�"I�O��ߴj�yW����BX�ǡ���F�b}:��	�c�#S�3������VsTYzDp�%�)Og����>�� g)32�?�&/L���d�x����&^^�3��^��.x�^���'�G�d\�ˢV���m���>m�<>�׬hܞ$\�S4㚻��Z�"t�n�$�����B�P�F�
C��mgH���M����it4/R(�Ɛ�ҙݍ�.$dE}]q�U��(>�'�6C����ƹJ�1ff�ƻ�t�>4F��u�A]��(@m��e ���gw �벭��hnL_~��ي�ْ�Fsw)�k�3�~�0S�HA��Z}U"��p�~�PG_��l�O(���86]���]�k�&���;B�s
���oN�r�N�6P�뵹-y	W^Xek㛫|���5��ʯV��XhEhS׋ͯD�V��������i:�0��P����Q�h���o�e���ե�������>q�F��=���CC��~h��,
L��I&�fB;���;�J `X�F��8>����c����Ÿ�I���P���C��tDǨ���4X:��C�6�˷��7��]�A�aAG���z�p�!*����ea�Q��	��M�����k]��]7�]
��7z��4�"֫��]g%��:!��}�u���k�g-0ʹ�݉�A0zNL3��ߧ���ꃼy�'��1"t�3(w�������u#L��u�� �P����R�W�{���
$�6:­���kmyt�� �V��N���$Vlï��8�dj�:���N!#璪$��T;ܸDSn���|��UAT��^�s~>_��%��0h��o�u�ezPp9�L�G�o��
�J�����,�K��Sk�|	��?(R���p��]E��po&�g���<d	����>,}G���I�&��o+�&� �t9�Q �qZP���ۉ8�S�Q�6����Q�ɏh���f*��Q
L8[0��[�U��Cꇯ=AaD�,��hc?�.��;�-�e��w/a���3:U��/�ټ}�>v[�o��8�2$��Ug�^?����eк�a�.B�r}�۱�����$�}�&ƿ�Td���0e���?�
l��y���L��NгiTa)A��'����Gay����^D`
��f�is�#������GiŤCW �VH�$C�p���]�<�W��pO�ǜ�������7��$�<��~�J,ʟ߷��{	\��\�\S(HXg��Q$a�Q��n��i�bv3��gG*y�q��E�u��n�cc�	m���y���VDb�n^��3Y���E	�s���Kn�kjC"��&�"��j>	0& ����vE���>ݓ���� �;�ȓ��|NQ�,��j��p��#E���1��̋<��5���-\9�y�Gk��@�
�᪈�<�็����m��0ߌ��:����:�hg��}�9��%�A���\isE�,\�t�ph]+��0��Li�.��}��l-�Ņ܄�zb���<ɳ"?fD"Ϣ�\u=�^�F#�h$[��Y�*y턃������	`���v�M�腓��G+ �F�X���1��:+�L�E��aw������j�g:��mzgQC	�S6)xM$�"Po~��KL�I��M-M���}F�6�'N�c�=�:�5�:��P�QBa0��c>���G�lX���I��� lg
�iu�F.��ީ9���IR2kԳ�DPz?��bbşXk��8�WARB������j��Qi{�/�	\���urI�H��'a��^��ë����q�Kb��|� ��%X� q�#����LŢ��{�U�o�[��m!OWN�tH⨑�
�8p��'w:d3����v������<&S�	a�"v�z��q�F8�5��I	x��'M�[٥,y�wÎ�c?lݝ�|Q'����;�c=_gp�0ƚ	�if�a4
s�X{قI:ම{3������h�X�������}�aE���]�F��?�f�Wp�d����(]�g�	��>b����{��:���fN��>��?  ,�0eJ�Vľ���E�L�'�����b�0��5)��]��o����^��{��l��a�c�1�'a��N=���T�m��,�^����/3r�m��'��:� 9_'%ފ��^�t_����7��l*;vIU �:�B�Hޜ��3Q�ⴇ���Ӂ.�ilNI�vp.
44d�8HA𚂶� ��v
6�eIˊ�qA�����=������S�"#S�Ό4����Q/{����8�5���<
Y����C�_�MT��r��=�L1Ts�Ԛ�8��9\O�UG'\P��LJ��<���UT�+t�oeƯ���I���4WB0��I�{��Fڣ3ԣT�+��;��]
�#K���O� )�ڃ�L�e�d�U�ߓ�Z9�l�w��׮�u�w^5C5h�ϊ����������b��*�.��������ާ�M�~d�W���r��T����L�![L�ɿ��˨mmB����Z��ō���F�.�@��8^y�k��U��hٛ�/�H�s�(щ�ٻ+��$D1b�W��r����),�c��kڐj��Z�ENX�Q���G_}{e��nG����A��F8�?��,v�!t�Dm�ք�I��ד�7sٖ�e�nt[y��nP-/����&��h.ztx�m���m�G�p��'����7[�7�.����_��Z�]�~*~�:�C������OkڰU����ʹ�#�6�����$���8^vZ�	�ݪ`g\4%��}̢1�d@t���Ys��p�T�F�E����@N��ԣ�m���63�1h|/�S�[jP���x+��c"���@��!I˩�X�2c	Q�c﷭�}����&�"�p��W�׽�-��(��a�="""-5��]G�J�+sx5����$F�ɏ����~�+���'f�	t%7S.�]2С��������+�X��>~����ʋ�gxY'!�m��}��UX9���G��6p�' �`�A��U|X6� ې96z��jD�P�k�u��T���a�8�I��}���R��I�]���~��\t����Ja�V1v=��1�r�Q�����'h�#�8sӖ K>͙,�q�lT-�Z[�mI/fv�Cխ�f�4� R����c���
<�̡�"@� �<�w�����i��h7�lLF�8u�'+��֭W�1�aB��g�j1<�'��C�;Ӱ��x�.���OmZF \r�&4�F,4�wjL;���L]������a�*&�ղ��ZBb��6dM�E0��!�%��s�!"����2s�\_!o��� �
K���!
k5�chx��m	���M��'���CU������Rf�Y"�g�1�I��WS��ᢗ������pG �	X=�(`ہ��kF�Rg��iV��߸\0�� ��Jz�-j/m�B	����Dq:[Ai���Jk2&&����xsǳ����909��~��˕ƉR!�Z�V�뽂���o�EJr�����C�����z�z#��γm,3�f�� [�P֨	`�k웱�9�(`��o�`&|��3M�5I��u�L��l�=]����J_��+�R��>��g|��%����ђ��{o�%"���at�r�X��]V�����H�3��n�yC|�1�b_07_}����ǐ#}�|���L�)����X��j|��>�V�Ü�*G�������%[��B���������"-?���0nNC�ԉ����Џ���~`�"{y&�]e�(̏�j�����f���P'��NWY�U�j߸�H�6MLɥ��T�M�����$�5�4�D��u�*� �ee	}h��c�(�74��]"���b���Cz�oT�iļ�_Y'���8�q��D-A�F�6ԖBl��=���,<�p�^��1��#$�G&��c�����AZil��'�,˭��X��XBطx�Qiv�u)��9Ɯ��n.�u��{�c�h�SOU 9ޮE�/�sluݚ�wL�H��y�Y	�L8��ع9���7�)_���I"l� �E�P(Q�`X���l�o��6�h�% ����Sw�O����h������n��DqYl\��o$l�����` �=�}�/_S_�O���x67H��y&�%I���l���qa-��4 X�41��X���@�t�c�����K��ߙ;���H)p��zC#߲�����[/� ��y9e�����Cxs�aAN��ef�c@줺5��2D����y���U� �[?;wȔ�/�k��d ��e����cރ}�(+�lo�����mi�� �	�6�>*T�C�m� ���廚�A8{�� 0П"�p%�S7f�h�M��u7�\�yQ�mQ��ʊ;���V��%�(-�n�H��e#J%V���O�QB����m�����o�f��"kKy\�
��o�6w�wk,f��3�m8��'z�;��w�w0c	 1�Cn��hI=��T�=H��MGc�W��!����3��^VI�ߝ��<�[�M�?���d���\.Owɴ�Hu���7�~ڮ_uqt��[�I �aD m��'���k iV��߷�\PJڣI�omj?��ie]-nܢ���i�F�=�'���Z�2���^��X�Ͷ��@��\��'��j.p�U�����G9��oE��SC�)z�p�t��!���ɉ�6�i�4�j�QY�߂���@:[�ijZ�9߭���w���
]�ٿ�þ�<{�o���pX�WM9�X��`�`��ݓ��^J��Q?7:v�}I�j�q^t���no�Sbad ϛE,���4�7���>��zf!�QM^����
��w�M�,���Dl�����R4[�8|k+��m5e2}��<���Bއ
%�Ѯ/*���9g���`;�N��"a�ز:�]�/��d��FV��>�W�@J�A]�����=.�W��P-�I���N�(��u��i����4Ƞ��W���V�����0E�Y��;�O�4�{M�q]wھ($��߄߲�Ɉ�et��A�tC"Cv+��X�gt���xQ%ff_cS<bگ�[(*EA��l
8=�7�S&|@-��XU��o��j@�c��N���a�� iM.���Z���N�0�0���Ƭ\�2mc�[��oa0�,'��5����f	.^G�'�2�XF��Yt-����޴�>2�~�ռK���6E��)��,Ӝf���ܪ�b�i��q>}� ���KÝ�t^��ޯ���)���ɭu�8�%�̗��>N(L$���7���G����3�������A��p-��п�����\�k@Q�)�����'v���kN�2��'E��kÎ� �b�rUh&�b�����j=�D���{F-�+�P�DY��}ݫ�Ph���=�-�-�~~E����m&���٬SS:s!��ʞP]b�jWj��t��-���rLOH�nm�Y�ߝ5Ιȁ���3��Јw`a�vit!�|�ڨ^1�<���9"�܈�%���x/=Ȳ�4|���={!�\��w�4\m�l{i�x�L'C��!��6c52�g��.�5u/_0�N�˅��F���K.=���|���_&D�d?a�����>e�?^O��(��⃅���W�{`4�R"�M�
 ��gyc�k��!"86Su�v�Sv�Cz�oV3y�:��r���u�.>(��{.&_�mNbcU0���*��7��������1o�c�+�)�z3ٽE��%��N�}�3T������)����?g��n���6�WB�k �����
X7`p �h�(�bej�զō�`�`�V7���F�H�I�6�&*'X�C=������f���-&*���ِڵ�i�o�#i�fz�ڪZ7�E������-�JLR��6*[	jU\��i�s��WƐ�M��e����'t��V�6 ��E�8�x��x��]_��h3g2�kb|ؖ�{��d���FD+)�
����%u�v(���%'F��6�.8�LY\�/a���Ha]̰�����q��A|�],{4��� ��%~�s��X����|����ID�	��Ƈ&8�#3>
���T�,��o���r�St�� �G�@�j�[Ę�"�U��!%�-�EU S����]���g��!��AA#�7��gj?E�k�/Y.-���m8y"��r7b���D�/�}Y�!у��V۞�t�����@2�d,���vУ�4���5����@��͚�@��Y(E�mk:9���ՙo6���)�:����<�xk�5���zx�8o��N}%��aIɿ}!�~��xӇCs�Z��2$�����S����. �r�^J�
mNC��d��+aGK�?ö�����H'TK���Q��^p�Z_T]=z��-�X���c���6R�z6^]	�l5c��3����%2��>�eiE
�6�Ϩ
yF�[�m(�DGo��0&Ŕ�:PȪN�gUhNhT��v�&k��S�/�;�m��sao�ɏ��?�c
��2�x!�	"�v�t���Ým��̌�هͦx#�]�`�t�z��rϪ�i�E�����a�nҭ�`5��� ��_+n�S�%���s@زϲ?.�8�����|y���ܰ3(=��)�C��>��9�
H����W*����kl�{W�aOO���(�>��U>%�I���D66��������f�皎��w6�0���D����W��#ڀY��%���L�
TG2^*4NWB�<J�8i}ݭ!�����;��b��� ���Џ<���� ��y%$��t-s��ƈ�BفE�+�!Zmk�G�'�df��c�Ӭ��N^G���C��M(-�/��0����B�x��C�p�q7�+m����LK[�A�`����qY5�a�s'��i�d��Q�e�U���O>:z�4�����	=�=�X��%a�>X8�φ�A����H>@?/��?��P�|����fg���?�L����\�{+�6���50ƌ�eD�ڸ=�av�DF4����2H|͋���M��A%�.q��҄��vd2���e�� ��8�T��攓T� �4ͳE;�7N����T���G����v�a��ڬe^+��� ���t QYG k#��A��Q.�Km�F�Y{0+/�2�Z ���4^�OL��U	����	!��sÏ:	��z�+��3�<\q����B�Q�j�p/dk��Sd	B�f�{��®���5���iA�ǣ�F�����v<k��������5��K|0}����Z��V~+�����5iZ��~��� ���E'u7�_AQr}�)�ěn�O\�K=W���v|7�<x�n�.�s�M�x��s�=3ހ*uH�/ճr�t�M�a������rw��E��ɥ�L%�7'O��q,=Q��p���t��w�Da#��͆r[��+y�-���z�ϧ�hf ��s�=lPS ���ҏ��S����"��3��!��o-,n8"}�&X����+�ư���?ZB�$�{�`�*z�ܙ��:���`ۓM�Ƙ��E�!Տh���3�M��@�F�}n4��oJR2%��J;�?>�=AJ\N��煛��rV�W�7Kd!�CA$2.˜�G}�%�BGҝ�2��~��[��ý����=VY�xx@�uk�xӛ������#C� ��۞��q'�_HNbi��&�p�>*�
M�^Z?��r�;֔�U��CxP@II�N�)���zzD+�z�~�G�L+�f��,�Nbp?$g�����V]���_@�dM�I ��*nԐ?��\f���.��9�����)�ы��[]m��h�^D�1GW~�Р�$� �a��pj�����E�E��_����21���A��N��6`����H(�l��b��g����l�Kw�{)TO]}��(��'$���9�x��N'�c�D�&�]<�ud������������Bm.���/W!���r>��u$;tz����<��*�ܖs����Φ�gRD<T+wn`t����ƳuJ�N���ǕFT�Q��~~�[$��'�k4�K�=H�^vӚ`Իȝo�F�vRO�FI2���}�)R��+��D���C��������I��Ÿ�	1#�
O�&dJ��^�s���0���2�։v�~��	�-�G	�2�L�Թ@��:���V��s6����g	p^���p�=n��gc��q���g�&Z��S3�^Zpb���$�.AFk�)�"C��k��w�K��;Cf���*��E��Dm���j�&o�8�ѫW��JҼ�X������8��%D*������>,�{3:���9��*Y�)EtnN�a ��j`E��|2�f�'�QUח<l�G!q�y*�ۍ��w��)�{�5�$���k~��V��Ic�Nx��}�J�oa� �m����@����A�}�`�a�˟��{��8��֩��m[��$?����,fB�1,��J�����,A���\6�!ŕ[�]9�	�c#EvAO(���J�����}(G�a�ja�2F�]6�بN�=��f}5>[ �S���^�`i"��G�i@��H������{�Frx%�e�U��G�d�W~�����n�Ї��D}tIA�ܷ:E{W�ĪM�4OG�嫩�����+~�,��{/�5� ��=���G���ǳ9�x�����u�P��J�qo9-t�����%'���"L/7
[�cK��l��X����,���h���oI`}�&	(��:���P$�r�
�߷��ޅ�c�� zJ�z��:���>#����_z�j�*0�F��B.��0�ڲ��S�7&|#)GD�����aR�Φ�d�����`{Z~�v��i׸h�kS`<G�t{!b
�=����ƿ\!La�4����h��c(C�$)�`ѱN=`I�
��P�}	˄�1cĢ��C�%(�x�ٮx'��_k�d�"=�Wg����'��w�u��L����\�a8lt�d>��>ҳ�AJ\�����ƴv��*�g�TS�	t��w�%�elj`�n|=��Q�_����,���s&�Mƻu��\��.�{ϧҐ'c��*�
S~������:A�e�̨��F�����Kb��(�Ih��uN�P�@���TF:��4b�$��&_�����z7_���͔{GG�.}vx��<̡�Y3�'YG6�4��&�{o����
�b�b��uoȘV�;��	kK�/��� �+��}�:{�nY�ӷ�|��ہ��<���f{��߰��C`z"�\���I)�j�|�a^?D왥�?9]���q����3����{
آn��Zp�j*�z�[|w'�*�wiV=�Q)<��N �����T�\�D�)D��q�yiT�lc�`+[��!��q��������,��"���EƱ+'����?��#L�1�{�bg چWc��DhS����_y��#Z�;wv6s�`��i�`�v1��>���n�%o�OF3B.APe*E���R�{�|0VA��0�-DL���xB�6)�R�Iu���!vc���S��:�l&q-��ah+25	g3!ߖ/��5"w��]:�3�vNnQ��.�uȀ��Wz]�[���?�X�U1�|V���}�2,T���y[F>׸��L{Ҽ��'bn�pٍ�R.�`���+F[�CU�n8[�!�Ȓ/8�s��[��ⶹ��l�W���}N�!����,�U,è�Bĳ�&6�*}��0�.�	���չ>��@����`�1��C#v�2�߫�(�h����ܴ&k7L������=�$TR��b�8��%"6���Iz� +�;����
�V�P�bA���,�%�}�cÈv�=vQE�^��vy'���!]��B�~��C����Yه��\.�����q�?�,��
��(5�@��"1|sE� ����Yv�ڐ�^+�`���q�IW���g�<�%ї��[�y头O5�k�a>u�O�9aV IsF��W���
L�z�HF/v���.���g��j� �
M� Z�`ٛp�8��l�[�,�ٜ��a��-4x3~$��FՎ�Z���s��(�M'S�3�uQt�fm�m�>������3~�������v�A�'6e���&NR�%���ᵸ��B@�냷`<�ȀL`�� ����^������������_��"�f�)��_�����*̱��a�χ4|��#��\{cEF!�Z��BM���V���)*g�
��#6j��V�T۫�O�n����8Ȋ"�PO�+L��㼷.��5�ff<�Z8�RK�|�m�e/�-�-�C�J��4���u�bPq
�8"��6�x&����x��*�ԌF�	�]�"�_[�Y{����������� �T7�`MU��=��1/���e5�
l�'���a@/7n�U�K����K+F�O���`�mZ�1�g���rǛ�0�ڝ�8gnr{z�C��}��}��5����h*g��o<�5�
�v1�yfi���M���'U�*�b0v>�}��*Ѥ*�֌���Y�aLY����=�=J�h+�ኔ��j�d;!	<�9��m�L�fy�<j���LY4c��TȮ�M&��\�G�I�ݒA:/b[ycRlJ�ޅr�m'�Ԛ�1���%��2w�O&�@���jܫ�K^YI�'��K�t�K���DEK���L2l4�u���W	/paq�Eu^x�ȃ.�ת�ȓT��?�]�3,6��D4=��OI3���W�j��W����Y0��2�'�q��[�L�S�X���H������L@�A���
]/�o��Nt�"��W��Mu��-���^,��^���w/BI�wQX�1����t5 �9��d�R�U���`U�Ms9NX�P���T�.igX^����\�������҇L�S�	2�`Z?�R?�:�G X�A�b�f#��}�Ll�r�>R��YYl��e����	}1GY_�P�8�ĳ�y7G�7�����D����E��h:yX~Z(|Pd�*�-N�_�����Q��h)m�ZZ!J.�b��ij�$fWMG�\1�9�AV �(:O(-7�����'`N��4*DE�c��Iu�A]ɱH�R��L���3��9~���׉�^�c�����k��p����xgAd�eq�>�߫��ϰ��vt��:�P�R�L��l^��uPU�lr�	N���U�H�t����~��aP��Yɡ3a���s&����~{"����0���@rH���k�HDE�m7d�89'D�p�u�!S�C��M)3f��#����x{X�vc�@S�߭��,̂�G�4�2�V�z>�%�~hg���	�4ǈ�pB�
��v=�o	�m� ��*@WU$��L[U���aa�{hT�DD���x��|����`� pA��`�^�
�b�I]�������R���u�"�2�B�]���YZ1P��ʦ�ev"����Y�T��ʐ+���
�J�euº�Y�Y�ZZ	Y�]P7쀂=d��H@H������������h����&"��Ď@o���� ��lϳ���&l��Yg�!�$ma�֪��#���&lfC�Pnik�)A�;�>�giz^|V�|�K_��?ʃ������W��w�}�Р�'<WBX�\�=Han��6��M��߽-�e����pYX�+W�=)�[ �Q�)�,x�vϑ�;�a�0���«����J�8ǋbىi7��(�wE��V��t�}��h�����(hU%r9rG�vd��	����7�3wЮȿ�(���$%ZIp��O�G�1���f�e�I�-E���`��S�ʒ���B�� ����%���o������+���_l��O�-�����6��ᆉ	�*g�*��<�����-�yQ���>���1Qc�����N"�z0_��Ex:K��ˈ��0CO	#��%5��YOӥ�P*��4�{H�Y�ْObD�z[Iس��;#��Y�ѵ��'��X�,�]6��u���hƎ|�S���Xձ�=^�/p�k�;N< g��3��'�vt��;���!�����=D==��h!ϐ>���1��k�z��Aؖ\`ܢ6�����V1��A�6�tR�CՐ%�oF���DO�p�H�Y�{�!�ʴ��4��]js	�>�KD�d��^�9��կ"T�i���Ώ}V�L��JA��2A�Au��sm���x�� �&��俷�Hv�=�c��$�@$U�s�b(��w-���ĔQ���Xb��F�o�C������1d6G�h���X��,w����l���]�旂�|_NN�~,��N��cD��Y��M�~�5-�A�j�j gֺIci��&�����'j���!S��,�u�YT�(_	5X����z���G�=�5��~a���f��2|uÜ�Fa���G-i�$�8�K�HW���'m;kVR*�'���h̹y����/ɫY�������#�=����-dΗwg��q��Ӻ6I�mz|>�_&!'���u5�r�\#��F8�˺��/�m�)^���n0�:��ܳ�f}�J�4G�а�!
����4&����V|m��jm9���'`G^��`��S'G��]Fr�*�'^HrWΗ'��1���ndυ�����|���a�F˺`��O�?!�
6�)�P��E>�B	gЉ�Dd}$W�'@�k�����&�]���[6��݂�}��d��<x;3`�q�B0���a��w؅u����ܜ�m9V��.��M����KۺA7�Lr�ϢА������P��D�.��7��m��V�b��DI��PhWϮ�lP��i�@��� �9�C���%�1n�%~U��B0E�1�L���+�6A�O�l��0i�g��H��3m�.��L�˜���v-ƍ*n��9P$g��=#3����� ѥqJ��?>�Z�����,!|!m~61oƭ�\R�h����d�5��=��(��4��VqP��JGw6�X�ΈZ�S�B�D�p���t��xy��-O)VO�^��EP�q5���7QiZa��ne�5R?7h@��+�OJ���GB�^أ
J����K��ٿ6��;,�Y�����;%}8Je�r^��V5�o݅�3�Ax�1-P�r��, n��<�A<�O�pց�'&�� ��QF,%�W\�
��艷,��� (��F��zG���;���1�`�%�l�n�xi�4��X��Iɶ����0��N�"�)Т娀�p-K�*fH�G� w���� ��eA0[a���&��g�����M��DPYL#<�킮�ݫe5ʀ��ށVnɈ��2�z+�����5�5���p��8x6������f��k~���l�v`P��!����K�CȨ-��lJ=xp�T�c8'H5��&��^F d��o�>r�E�Tp��l=��{��R�e�3q���HG�T.`J6懽��V��Z��,�~X�����O��.7�����D�a����K��0TY��ѹW�tM�+9> �f�hz�
�l^pS����L�Q�1�k��_���@?�i�s��F�CWo�> �+]�q�ړ����' �K���7�E��^�S�n������6 ��=۽u��J��d��|'dc��t#�A+QK�aF��H�!K�j Ī�p���e#�"l��R��׸��� �\�*�ނ�(o�G�'f�UN�e��E�M�UɮS��h�`�`��ܽ���Z��%ۙ1����FF�<�q��7�Yk ��	 �-Aȗg� i���#t����]��)g1	�-��);�ұ�!�f�V�����:���I�f��#�	�Z�;
��M*�y�g�L�	�b��([8�
뽍g]�1�f0آ�EZJ"�=�o���=\=�(t�z����X5v��x�v؍-[C^	��K�0�¤�8ۺ(a!S�Ň�q?�xr��d-�_��p�C��5�,��Ɖ<r*��Etp���.H�z���<�#Ls���q�]�^K4��޲�K���ܩ��bW��֣��(G\�H�j�3��j/�k�cH�7��{3~i�KV&�A�iwYلӷ�=���';?��n*ʏ6 �O!��g�E��k�E�.MX������s�N�����j�3mi������0p�5�v~��P��.��x~�-��!�U�g?+����h���?rh<'O��#2���4�!��G�P�Qr������=+�c*XV�ɼ�@� q��OV��S��T����b0#�*���k���V�������gm9��ڼ 8��πk�Q���k���|�6n`�����EЭw�:@
'���h'�n`�&��5K�캘s��c������kǫ�qZ��`������J��`����E����]�,���
ޱ��ܩ ex��20JA�h����"�^����фbE�'͆὏���|���Tōck�t��隴)��Ί��JD sX���YR�C�����9����`�-p<nSZSI��m��OH�1�`0�w��8[;�gc<J5B� �|6�ˣ'�,��k-���ِ�BڸsU��l20��h�{��������,�Kc�g#w�,Z��w?��T�aKQ�K�0kg���F��?cW��+5�B��-��.H7H8@����vU��}B�\,�^j�U~Ϩ�?��?�kν�\)dW�]������vK�Q�|8������L�R��:��	7�����G78(+�z޳�|���(�9m8}B�XG������?�$��q��k/X�dL�uw�E��˸�8ǂ˺�`�92�<�hp�$L�G}ܦR�ݬ�#\�5����w��)��U��S���.���@h�}����X?ĩ���F(�2��D�<���?9�.˺y��T�Je�fվ&�at�͋I6��N�$3������ݻۑ���JR���~����o5�Ϙ��&�t�D�sI�Ԋq�BbIMT��-�����9#!n��HE����9)���8=����$��JF����-.%S���<Ú/��r�fq��s	:�o�="\h�,!���Ee3��϶�N�~ʋ9���s ���9X�ӼaJ� �0��+-�M�ዓAǜ�!���q��\��Jf�9��h���f�-݃9<H�K�v�)���С�Б^$S��'�Ŋϣ�M�1g
\��/�������O4��x+�nuo���f�p@dD�Bzm�c[�S��L��\�d��2١��~�5�)���0?��d/3�Ø�iS��}j�՗��l���I1#I�[`Jbd�U�	��3*0���v�|�K_��s�����mj�L���,x�;�RbdL�F�'S�'m��}�LY	���!�w|��c*P�#�'n&��%�%MLj�̄��֖M�L����O�ܒQ7��5e�`�DY�����Ș��ŉb8D�����!N���! ^Χ:˪���V^��(��$"����>rBw����Տ��Ǩt)K�4��Q��"m�T�3ڨ�$:m|=��l�)-���F�)����]�,!�f�![�#��V:d#>��H�n�G}CTڡiKo_�B���Ĕ���<8��\`f���
SX@�9�Fm�ے+]��:��n)[_{Eù1��d7)c��tW�#A��v~�©�w�$�� �Z��t.i�n]��Wp���JkeN��L����g��{�T0�q�����aNk닌M�|��2U�-I~��u�^y�݉	~:�Ǉ[FA>%�]*��k9�D�s85���MΪ�	:�㮃E�2��Ҡ"�-�9z�������A/ۭˏ�؃��A�KQ��	)lj6�,.6@ �����,w6#� [#���M��K5F��Pd�x�o|�$`B+�	��UP��b��s3rW��
;�	�x�:/i������^�!�ꓧ(;�h����I*rʬ;k�&�����/�Ѓ5S[����ko�V\�y��O�XG���x�jH�⦁����ؒ�R�`{��u8hq�lZPZtr��N�[�cEQ��Fȿ�^]�
�0iv�p�j`��2#r����1#�M�Dui���	I�Ա]�5��!\����ک֘TpG�:��pt�^S����۝KeW������1�I9vD�#<!m���G���,|�@=~��ַ,x�c�2�bv�6�~Q]":���̓��FOy��Oy�;YGC܋���ڍ D�E��#MG�du�8�<�ݶ��jh:������Ȑu5���Yh��B4%>�4	9=��<�-RJ�ܩ�c� ��sw���g�\��� E�-|�Ie&欱}	b!�ͧԷ��
�ۏ������wf�Ye�A��(���6��sn�A���ԃCZ'������SYip4G#��":��<dF�E�W�*_,�k9���z-�`�り�n h9P1���(����4�dlM����qGe$^ʧ�TV�%�-���Q���GD �'���_C��(��T\���~�-J��|��h���G�1��MX��ek�ա��[:/-��R����in���d"aC�,Xh��(�h^�5$`� ���i����}��t���G�t��EzZ��a���*:V5v�-���-n�V_AF��cp�QU�,��|e��&�����Ԏw��ͧ3;�R�nNT��R'��mcR�o�:�m��3��l_1x�+�$x��4��?���خ4}�sIߋ!���-ky�5��;p��-�s�j�b�9Ft��Qwr���V+�J���b�Жɀ� ������2�����OQ�l\�+��>���X�dQ�G����� -�>��ɫ���㰡`�_�bt4Ux�JS'��H������/�ڹ��:��e5�	i��͞��� ��;}>P�&P�NH�"S�(�R�S��\qBE(�"M[l�܁^,�S@�풢��7e�Y��`�����t��қ����@oָQօd�}�.�B�:��?T*�u\�#T՜1'o�x�W� ;�]XW��; s�J>�ã���rB.���U�l�o���"Tč�ҕ~M,���*��%d�SY�U��մx0G�C �G�e�ivɺ�V��@8$7�F���|�����0��	޷3�cQ�y���j�u��W����)���,��?�N�3�[9�"�G�~��e=���U��Tؘ��O7bؿ�c��W�<��=g��<5i4�rBtt~�Վ���i�<g|�IM	n(<8+�Y�F����D)��_���)�����7^�|Q����$�ܳo�u��G���[�xW�4bVE��`I��Q��7�\\}���υV� �=~��vLX�.sf�(d7��hg������E?&ijR���D���z�ȏ�F�4�����o�1��p�i(8A�Y�).�
���0n��������&�%4N2}��!VXu�10�/~�li)<�RC�b��	��J�����FZ�pjQ��Gl�F���t�
^0�"�&��g����{"�FId�>y�����L|gm*h*:��!*"[9�W{��s/@j��5dϱ����t��G�E�?���'㻢�'ė��*���	l�,d�f���c���%�B�t�1S)Ts9ѐ�aH��T�:Kv�a�8Uvw��k&�)�����+�Z��q�;���i��}CrӞ�#�6���j��7I;�tn^�tQ:Mŉ��O�y`����|e���=ڬ�*�"$��·C'�_97C���k��1��I�����`-��
�]�ӂ�
�bڣ%*����t����� �)']2-�ĉQ�_Qݻ3���a�b�%��w/��n�Z̤��}Ȯ�R��If�8ێ�	4��F�u���n�r��=`J�ۀ��%��|����݋����<���٭��
�L3`��"B�l��0e`����Q/)~�&*M�n�:�+7�D�Ѡ��Q�J��8e�L���>�s�#&)fͼ~����(z�!������VCi����*��:��������B�ʹ���iAB4�]
JT�&z'&�'^�B��\���M�:�y�8S�c�ʡ+�Yt&ѩ¯��,F�p�n+Q�$"���?B-`��8�TR���z09v���s�_�$Ѿ�N�u�OFdC�ۀZ�ܔ���!)R�:�ț�=d����0ٴQt��8v�=�T��K9��疰	.��e����e-"���=��X�	��n��1j�S�
>�J�B]*f�UF��0 n����C�I�����_<�{�y>��t�"ų���S~3���Nd����lv�4"� Fr7�[��j"\ɟ�$EӦ�|�KPE�*w�D���N��!��4�y���R��!l*8��n���5��
�%����O̽�\"���^�f�:�PA���+u��iY��GCmј��~Kбʙ�NQ�C�*�\+8��$ͷ������B�5y{U�d�3���Z�2�ATj��2�6όB�ޖ��)|>��C�
x�s煡u�NF[��������zIr��ۈ��֢��nb��X�砨(]?f�p�_>o➀��g
�$>�9Uԃ�m����׳�p%3�
���,��m�����H�=��yƫn,��?�n>�W�0N�pO\�����]J����8�X\6��>�:�Y٦�y�l�CX�6G�H�0LH��'F���%��~������0m7�o/a�6�^n�����}�т�Y��o�����{�=��JƸ?N�X���F4G����!?�KQ)Z��6sv�`��١;����6��r.�����e6�ug���KN�w�c�-\lSV��	ҝA�^�iYῠĸ��KCxc9ƕe3~Y;�,V|}w���h�МZ/��w�d���d��f�0��Jb��������� �������k��k}T畇-n���l��t�%�pP�@�ϖԷ��	:՗�蓲���X&<�EI3�ȉ��.���O��qG��h�_��o-1�LF�1�� Qڋ��Wq��0)�l�M%A����ݫזq�mB�����^b)K�����9��#���j�휓��p�0�?�~A��Ё��,g/·P�0*�Zp��w�%�W�(�c����w�O�C,9EIZV{z����Aں��Ю7qY�t�	�hڐ��{����cH�'�
�t�����j�\�]�j������^���^ A��a�����dZ��xC)q�R׌���,Ga[C}h$0�u�[�p����Q7��c����h��ˮ.�_�LG17�Bt�+�~3����8a��g!�a��rAK(�<�ﾎ�E�Oqe�=����65�F�יhx������2�_��WOwڟ}����5���)��.�&ʦ R��#���m����������'pB���构�,
]�H��eaV�L����e�W�`��w�2��ݯ�	)Nk�_���d��>�K:�\�W�~.�qx$q���h�o�M� ��q�;�7#`�([Ϯ	�  �Q�ծ�m���R4a���C@���h�P*w��re�44^<�آE,_�E��g?#/��8�:맇Uc7�$o��k�Ri�D�4�}�4��^yX��[�iuI�
2�n�d��r҈�{B��#=2��16�l�ӈh:��^��'������u�C����Ù�-Rjg��~�>�o+u���S�"��V�O�@�-t
���c:��&gr�JR����V�}+���e2b,��|w=^�>jC#���!:��B�U�<��0�M<c����=�f���E�>�𖁶%�I��O��٥��v�X�1IoM��N}�;��[����X!�r���T����Ջ=���^�R�>��H'��^i�Z�(�������Xa��EǬO��(��8��y)H>�Z����VM�P��yC?"cąW�:�#=�r#O�W�h(Y��)f$ w�oC��D4B�{� ��2�[p���X�6��=��*��w��")*BC"�����<��Q<6��^o����'��q/�1r�����x�cD�Ea��g�2gB���L�5�������K��_�q�Ep7ٿ*߀Nm�ʭ��/�����Qu,_%�`�6�Pޒ��W�r5�+>*�9��#7�=�/�� ��p�����X2U~��[f��2T�.(x� 6����!����|U�Q�^��3����:���Á'�>��m���ך/g�b+=h���K툉�I�DU�W��0y_���(z��!�2`4��&�N�xEC���g��H��жtKx��h��p����W:�@�H��H|h�_��٧�5,z�r�u_�w�Z�k�Ǒ����4�
Iȑ�7�� yvx5$_���Ť��k��G�?�G'��҅�:OEJ}<��[���$�<-���Gi�����u
��⬄����*���G#������+�P)c㶁 ��m�
?)�O|���B�;}�T�&��S�����:|���>D�E�prR�c7���!S��=[�7��i�&)���n���p��fnS�+2��1g	�?����_[j�Va��=M\���(��cN�a���8��GB�rxƲB�J�pfo86�?3i�$_O�O�Y/�Kk��w��z��#��^���ȱ���,��ƛ�l��d�Ҿ��ի'������u��4Q?|��y6�C��%��{ٴ�
�q玡���Ì�$���0<��K/!�q����r���jx�}�
#�Y��$|��p�{�Yl0��:(�#�k�U��8���A�e�'Mx������KK�5I_��6u+ey������9氠���:,s��x�[N�F�(MK��y>�'B�}~�p�E����
c�:���~�ݨ�:�c�Ӛ���}���� �|'�k<7����@� dB�R�I�F W��%�����<���1LҖN��_	���VS��4t����?bn�nM��.n�|P�W�R���	�	]�m.��]|U��]��z��wVg�{Z��5y�d�P��y��2�}�g��P����bU�[����4�\��ds��~�?
#�_���}��Y��h���5�i>u�ͳ�*��v{�K,b�W�����\�0�Rm�l\H�����:�y���]>���-�)�*� ���Sy
���<~�q�
��&R]��*,��QۺV���Q

�H�P�J���7-�X� �	
�!�d��k��+�v��~{s��y^�[�>&!U�Q����12���7�'����797���Q;�5�ˑ7�������]�FO�Mg�3������.�l~]j%m���,C�{*1���7��H=;|��[�;H X��he�ƽ;�Yj$0<#Jf&m���rl �!G� �:!��
 lˎzJ�T�����.�]�H�d*n ��l;:B��6����s����ޕ˰�4����/����h�㰳ǁ�!��j\�Z�9�xQp� �ɿa���w{��q�'���R�EV�v����Խ`���D�~�0L��7�����i�m�U����ZO��nGK��|�?�6��"�g>{��Â�v�S�5�GL;��{�P_r����K�?�\�S�J�@<�x���,ψ����e��O0Pb]�f?�����#��Jr��o��7w���/�W(LBO��s}�F�����Q�m�y�m���>�d{YsB�p��9*�Z,���7+�	>Ip!�η��#�h]�Poc��0�P���gcꯇ���4�xft�.nƏ���6��&$��}�
�ލ<���"##������lC:��oo����{�?H�jͮ��6#Z�pU�GsӲ(��0��@�o���%�_����LT�s},�3Jά&:��v^R�������΢�����s�v���P	zZ��,�ǒI"�{�3Q�Os�=�±^�c��u��H�_g4�����4rD�º�	Cb�<�+�H�M�$;KH��$��g��,<�_P"\�_�����WR}���f3RU071���18���[S�*��ݰL]���>/��s�\5Aa��2���UU�B�Y5�}�0�t:Mʬ���o.�G(+(��vE{7�f�:
������J�W;on���r���������P�7�X����&��pA1�����wM�e��u>��>��
�?�� �d�e ]�2�;�G2S�Q[K)!*]l��5RzW^���1A�v�Zd�͜tƅ:*e"rs#þg
�aA����=H�5J�o��{)R�[�_ގ
�O鐅TGU��Nx*���nt�jk�;eИ���S�[#(�\��_�g�7��lT
�S7s��G�,Z�{Tr�x�uG�TB��'�\-���J�;ᙽ�JA����\��M�D�xճ�'�¢��U;Y���'S+�C�Fh���*�p;��jW�>��B��T�y<Col+{��͑A�d6!P�z��._jЧ5ˌ
Ɓ�3��:e���x��t��1���.y�C5�_�/C����1!��x�[�&�O�t#ְs��^)g�d�2�1|LϏ��7��]��kh'�X�Aj����B��r�,���_mQ��� w�D���v�b�s��2���s2���q�O�	Py`̸Wi~S�t�Qk��W����Wb4{�47�4#��%h�	��u6�: ��w��ۦ6�|g�H���������	<��j�\Nh�q���]I;�=Ts�px��O�s�	�U)5����y��?�?��_���!�Q�:M��P��
f�ka1�ۦf��w�ww1��l�؏Ll3����������Fc���/�����G|���ë=`
Ր�>W��w)5ְ�|��X�����{�[b�	�6D��M�k\����䫾����M���5W7���6[^������Q�KI��Kw	�(n}م1�w�#�?���ʎ�ʈ0�>��|S��	�
�V$��"�B�M7�,�w9M"��C C�V��.���݆͛�p8�f���L��c>oC�~r^<>�o,6]�����d���`z�H?��⳸�D�;(Oض�qݵ��N�3���gO����7z� l���P���b6�� ��v���M CӦ���	h�Q����]H��<m	��h��:�OF��9�>n��/�M
 ��f���i�
Xd��˟�O�fCSe��yO��J(~��p]�8���I�,Y6�@?��v<b��L����ZX�-"��𢜷������x�C����z��=���
W���r�4�#��6-��%O�+�]�86��,[���3@XY*~vl;<�	|2���U�v��u��98y�g�tŚyu�Q"$�X��fu��Vs4�x�2']��3�<j� ����#�]�~�����'(�g�u��Z������G�w��`(84"�.]{��\sB°���6_����%�ÇU�-Cҥ�޶L4���$�-[;J�,q-�:�� � �U��c	��Y�#_�O��G�<&۶���*�U�蘒bA:5��&`]nH�����:�ł���!������5F9����bWZܩx:s�è¥�m��A��v�1w��M�C�) 2'��yN?��X�NXχ�h���얺����,y��?�&ɱ���w�T���6�2�L!H>>��mw��n[��n[@ ���L�˛�b�L�_r�-�cg�9�,:��@��HC��ܿ[WH��~BG�B�0�4k6��ګ�D�}U�fH����k�4ސ$���d`�X��/?���Թ�+$���;Z������4u5�@�Ɯ��'
�!��հ�=O������q��X�Ǖ����K�Rmۅb�a�&���>��F��&�?dX��� ������=2p
.��
H��!���z�ufh��&�#ܜ��t=�|�Йx���7�}uq�ć�������A ,�魟%�/2r"XтRP�/�`�zX<·Y�I�B�s��ݹ�q���Dw��V�nl�d����N���Sp�!J��kE�c���C��\�ĆL��f�"����,�ˈ�����&�����y6�C�����Gg��@����!�jM_���S�ȍ�sIn��3BR�$D�P�v���)7�)}��XY�����"zTU��_'��������q��ךr�n�h|�$���<���v �jT>�o^N�_�\�U /$���|�"�s�!m�w�%�!��ͩV����-ǞzK�s�]I�I��
S�>7�&墂�#C��L�$:���ہq):E�*���:~��rBIe�魭&J����m��*~��+�FfhQ,��i�'ٷLsn�M
���zĊ�]l�ڗ��R��	��M�{�FBu�bhu�F}��ȧCӨ�"�P�k�؝����\�/끭��m~�����L��<��{2jA'V�e�E�M�UK���@��+b\���ЛdIf��p�U�����E�~�����i�4��K��� H������1�q���f Z"WP��[��o��~�wMV��Qω�+�����+/7������n��e�C+3��bw��Y ����ۑ��AX"��L� ���l�q\$�q@���:W�<`��A�F��� ��0�����W��aS�
?eQ o�[q��>�"ā]sMDW$��Qb�Zy�����R�@t*��pϽچ5D�*CD�w�(
����4���R���ܚ�E3�����h�CÀ��a���pU.j?Ur9\��`Lʢ��2�z	s�%�e�$;���C��T�0�R2|�;��-�&}����g�]��׉�$�e��t�"umd�A������{���|ꦅ��t���r
�Ѕ�zQ�:�RQ��C��{ �\86p{��x�D#�0�vyH��|���o�6'�c"d�B�f�E�g�����G'�}Ml6C;劥�ߓk�t)[����C���P;�"$���[0�O�ªBdP"�RXi�-AR����1E;뱟�2�N*��� �0��=����B�r���~���M���'T!�eT��3�+�����)��WH�H�ӑ���x��e��rQ�F�m�`���c篥��#˙* i}�~�^cT���N� �c_����yPk��H�-̄�(����)Ρ��t���E���؊�o�>��K�A�+B:�d��+xH��9�رDT�CF,:P:X�9'U\�QA�.���1����g��~}`��Zγ|?t9�؟�u�0��9�|�q��i8�~��ՔKν"|�c;����ԓ�FP̨��[��Xo�/�_��� �U����R=���οW��Vsn��r�?q]3~:�w�[7�3V��n�~��f��N����3��V\���"hegX;w�ܐ3sgk�O�t�5P;�h�$̟��y$�Y�N�w,r@Ξl�g��5��h�v>6d��w�.wZ(NTb�cE��:R#��,7h,.*^�|�;�yR�>k����)b[�����6bZI�iX���ZƮ���~CF���?5�DfdJv����M L��|)=���h��U- �
�i%$����hA��,H��}��lZOAMӷa���Ϻ������펕�j��{&��!}���H���U�[Z�r�{��Fޮ+�C������L�8f�[U)^o|w�GLw����8rO��&�er�x혥���ዻ(S/lj������AB@GU�!q��:����'��������x�)x<�\�p(��`9��b����wN�G��T��&L85I��'�	�X$;�!�WdR�قʭ|u-��wF��Ι_d�T�>��F�uFzS��[���3Y�U�J�)M�PX��u]ެY�����Qh��^��QXT�vE0�ij��7s��� �0w5(�q���GxϗeN����������̞�+�4x�����?'#s��X��M%$5���Yp?���#�Y���=����o�YOjA<���J-8�v��"��qlʟ4�`9__�	��k3)A����b٢(����٘���&�$���leI���p��I4��L<2�6[�����4`x��|H�V�~�F�i);i�S��~j!�\��}���A��|>r ���q��~�NF*E�`�1�ݦ8�Y�6{�n/h$:��{|ְؼ�mr�G��1 ��N� 0	Mz�d20$���.^	��_�u�2�W���r3�:&m�+�ENb2�E�I�=�p� �}'�"j���K�A��հ�X��r|�E�؂�KJxԢ-���8�0J[�<#���a$�$+��^R�33��d�د�Zs�A�����=�5�S�ę1XV`RO��`�|F	&M�ٱ��,�H#���V����||��=:VM�=�Iw�urwꐸ��4���R9�NT�ԉ;%��	���U��k����h����ˠv<H�9��[��qC�*	����l�*��3?�\��q&(�.��a�Al Z%t6-+<ݵp�S\���Ď�,B�8�%]cO�+Po�'�MKA{��5g��% Ѥ�;����!�lx8bd\3]`d`rg4���>����N��<��m{6��b��b�>��k쪂�3��N-�E��G�p�`7k�ӻ{�� �?3�P�����𰔾A��]t����y����S�fi�b�t{�΄;cc|���jk�5�X����W^j�|�C9��J��W�r�U(�<|����i�pZf>7޼M��7<�`Dx���k*k�X:�fX:�"�ea;�e�U+[��Vז��� r���"���"x+v nZ����U��?WO[q�+��z�6��ϐĺY`|����'��6c .m��*��-F��7��e�+�=���I�I�b1Խ��z䟘2Y��9���Oo2�׼���_�K���5�>��E%�ߞr��t;��t����]�Js�������-k�i��=V�k����q�@C؟��(	����_ �^��`<���2���Z���}��T�����Tk��:t�oj�+(��� p�����
��"ta��)ɴ%l��޸�����#H�vR�)�׋Z���@~�]�5W�	n�ѣ�F�ml(�9���g��Z$�,��Za_�h�-�U�@�o5\�����.ez���j&�U���o��|���T89`��n-$�.�V�8�-��Z���I*�!�]vs7�9�"�b+�\7iF�Z(��
8\ED�bH���a=���近Z�:�Sl��B�u��+�fW����ն��Q�͞�`�x�S�O-ƨ��ϐv����3�T$l_�:�2��#��l�-���J�z���
w~�E6�"����f�����E��n�q�(��á������j�6jJa��/iJ���^�ѷ�����誳�6��ڣV��#IR@�Ւu~՚E�[[p|��T�{n�4	�;�Q�V2�%Ci�2߃Rz�����F�M�ں�}_�\6� ��y� Zj�׏�}1�s�\n�dh�3Ƅ����aQ�	���8Є=g�$^מL �>���V�����3)�`����p�/+4�ao)�i,O� V���c�ܶ��o������ Vg�^)E��,K���P��r�FFEn�ṹ.��a�T�p�0� S���)PK�:���خ�I�\�4S�����$h��mP>�O��}�"��=��&�q��7�Zh{� &2-G����P�2��̃��RnA>�����^�.Y����s
YApÔ.��b^$�7��<{e�s�%�� �byo���CT�n�k
�[���]�)�\��Y��$������!&ڛ� YԁA�<�:څ�Ea�Ϻ��dzMv��]Z��ǀ�wTz��]EI��Ug�xq��_��u��s��bY�HB�ŅńӢ�� �O:N�#�g"shCB���j��>�՜��?:<۾V|�$�RR�Í��4&��&������o�4 1���AKŞ"Ǟ��>�ӎ�Mg��'��?ڪ�Pi�E�+ys���}ߖ���<��Ҙ@���	<��Ror��Z���~ 7�p�n�N�l����uz���A�~�-����q�e<L4�T�����8�(�/`�&I~G���d�GF;2G�U\�×�u.a����4����^xMz|��fD����;i���q�%�Pط8K��1�⪅�Q�F�z�MAS�ז���+85P��;�ᜑ(�ܝ��-Rv�7q�;�肑�9��OV.�O����{el]���;�E�2���#��j,cYo���7���U�D'��a�r���)z����TK������)�I�^]�@U����|?/S7����zq�<��m�ۨ3A�\�2�S�v��w�_��z����	3Rg���4%���Qw��i�~N�6
�#�qV�Z���� �N؂%�g�	-5��[�&�e�����:W��Q��^�д��2����Sq�
|�)��9h[�m0&��_�S��ީ���':LW��-W���S)�x�����(�ӗ#�Si0�z�T���;���0ⱦTz�<�e��.*ӡڏJ\I�GkmxbX7XBT�?��%g	Ν�_+2�ELj�� _H��l-]A탭�b�J��+�{p�(�kk8�k���6�".V�_s��s�Xf�8���`b=��ͺa����M����1f���oYN�����@X6�q|����|@������i����}�(v���v.�:��$E;���ѿ�����h�?�+T+�Y�nI�G��?�c����U	�H:��o�v0����_�ުY��ե��HgE�?!&�z�d�/F��N���>3���]OV���,��l�߸<�w�<ֲ�>l���&5au�zI�@}��j�6I�>K+�@̞+B��uhv�n�C�9B�\sh����\�h&���u��я,�
B;)35�`�����kH����"�^G�j�:{6Ӧ�ZEN�$U
ޜ
x5G�N�7�R:��4���R{��*�'�A��"c��� �w�~+��Vw	��|�SICe�|��z���O�l-w,ATV^�#(��\�5e��~i���e�r��>mX���ʳ��V�����jZ�,G��|'�q�N������	�Xӎ������qH�?����nF�y��K���Q��'���?�@�$v��P��v��z�z;�MH���Č+5�,,�4W�泑l;�ܑ4�?�0^���������M��+�j�;}�D�:k�Cꚰ�O�i|("`\��\��{2�w�������`��f�R��R-A�����7�B^s�r7	�'+s�s=ss�����g�X.�:���M!Sz�Yc9S%Z�����1��{��8���0��8/�7}��ȋ�Z.���抎,�Ӥu(���8����8��kȱ�KFn�������ӎ}!��L$B,��j����Pd�^MN��'u#^�m��D�o��p¢�Y �g#��y%h�@B!�I��l����}�q�-�[��D�]�3ĭ�[Va��^�Y��T��f�M12p�^�B�����m줭6�28���kg�)9#QSk!��ݘ�� �����v8$�"�h���<�4�2k��3y�P��H��,g�s�����R�O`Dc���Ҡ� T"�Ͳ��Q%<�I��2�>�!\Zb��V����c��-�-�*H[�_� �D⤀�zω�EdM?n���!�"���L�6���j_�q*����!���!�Z�&T�]4Pt��`5%��\��&��R��]?�P��9XyY[EY�I�m�����A�>�	�ٕ%_R̝��@r�� zC6�[���4�s��k��3. �[dnUa>�c��jq��5��C�s{� '��Xux#����ezN�F�S:Fmv�}����j1�����K�k�;Ȗ{`\6���F+r� ��zl
at��.ז�KT�r��lY~���!��"��Hq`c�o��c᧝J��[h�s0~1���V�b~t1��:��T�ѓm��W4_�,�5�6"qSf�Q tgzՂ�jlCD�9���<��¯���s	����ؐZK��
�r�%r��P��B� �\,M|��H�/�Z�-⊧-,o�u�xk-+ae�k�U"/�c�y���mN6��yq0����>��N�\¹�oM̿�#�Qe��u�Q)̯�D��	@5-a~٧O#�Cŧ��5y��-��kG�A�/�i�v�O�{T�W6��2y"�����Nc�{f2����FHS���l+����W���mA��B�����RU�'�:<�#�
�~�5�{w�'ӏ8AX�8_���9����۸&�]1鞐���#d�O�4����7�_%<꧒��TCݸ]�d�o�%�2\��p��2i�4�2�gȒ�4m���TCR��i7+�Kw�CF&�,��l��Z.��g����)��+��[�6I��	�a�7�/$�^#�g����⠱�g�|�5*7+R��-rt�4��Һ��T��$q�fU�p�KA���~�ʏ�y��v��@c�hR!:�n/��fQiz.�r���l�av/(�����r�,\�Q�E����D����k�е�B]s���i�1�e@�s�6�*�=�(�F� ���2#��&���+�rt�k�n/�VX�zL��ϳ�� Ȅ��5�fg�B�T��_���ѯp��~>W~�U��G}�n�"���;f���T}��l��K�VݠnJ��Ȏ���v���`C �ac�O���v�_���_pvl�Vb����/I4�D��3�hg�;\���G_ǚ=�cT�.q n8�T�*�Cf�yiϔ��R�u��?ї�_��bĬ����1A��:au����k	�b�IO� �MO� W��s�T����[�C�@�׋=����e�?d�P��d�B͖g�]�4�ߘϚ�W�k�c7�DD� ?. ��$�d6�,t�|HWѓݦa��S�.�t��so��7Q���=#J�[����J>#��S��L�c�k���LT�R�W��x% ��?@y�͜%k�1"� �V9^��y Z���"�
�i�4�8�dV �9�����h
��LhS*x��\����,U�[�Ջ?��tY»��9e?�]g<�;���&�C+��i�?����,[܀CUf���V3N���� ��$m���+�i+P���#��тY.���{~�mɸNX�	�V&|V�TT֦j�*&A����D��G�o�����Sp������WHm)8���	L������\y����ߍ��h�x�%v2��
�������p1� �֒��j��z�z���V��z�y%M��S�V�n��RPGF�}K�</���ޙj#��cߒ�cȔ
%>�����L��kt���'�;jc�3����L�y���"�e�Q7I��ć"CCb��A��}�^�B��兦
�[1	!���Ȃ�	])~���V��Rk-�Ү"C�F�v��S�3l9��ѱ~%|ǒ�(%�L�gxJ�l�V�kA�#A���_(���{!���	_�i>sFb�a�8-49�D����P��L&E;�LaϦ��+�����x[s�m�!1��m`G;�,E���U�_��q�n���9<vx�/�m�Ԡ�4�E67H^�I���ڏ�L����+���*!7Ɛ��x�c,��GSѫ�y�]����,���S\��x׎�"����3����Ym'_�g�0���W$�Hl��t���%4oa����9���B#�Y�lA������>A{"8U��/_s4{2<�֠i��	B�
7p}Y�t󺄼1%�4�b�����셞��p���Z�]�dk>�#�k/�Y�xM�rج}���S�.��5���k����QEH;L�]~�5YJ��N�ON��c���)Nŝ�(��+�l9.$�q��')-}���^��� ͷ��9�[�;�I��-#,�SX2��cdk�ҭzj���YN���A2��9Nlʮj���י���P��Ou��"���;v���%�拓#cw����t��4�kv)����sS��'�r��[{�oVͻ�/�I[y�4�+�޴	�t��)E�̺�B�\}|Q+ jK��eB*�M[~����/A5�#H�w�d0_��s�A�����X�(�*R�*qb�B�R)�Jj�!�yy�����uj�Z���n����+��+=O�W�C���K@cP��,���G������ 4�oOR�订k=�
S	6-��r��B�K���<T:^�m������T�h��?>�őQ1$c��4՚~(�����
�[},VB���i�͌Gy#�P���,(?�%���i0/�9!g�.�����aq����Pxa� �1K�������=7����7<
��_-�V��_�ַ4���*g,���
}���-'#~�OR
8�N8Y=��U)r�2ffiF��A�q&QxXϜ��);��lS��Hkq�!�N��f[~|�����9uM?��s��#8-�3q���A/�B���5�XN��=Z�bkm�|=�>->acP( ��v@�i�V������<����Л�X�k� B�<���O7�ʗrh�R4Ҟb���,adU�������/�����V��N��o޿����+'}I�ڠR���������b��q�jn��_�գ�ৣ A��<	>� \������6�J��p� [CWn�w5foIS�[���� Y�y��{o5��YX�ܔ���p�M֣�/|��Ul�nQOUG?�p{�o�T��(����"V�����#{��X?���`$q�����4���M��A���}�;�ARҍ�Qh'mZO�,�>d����k9��L��g<*�碡  �V�鞿��-!h~N
�]x���j�O��[�����=0��
���8wr��ڛ�c?H��ũ�N,ﺉ�L����8@K��S"2���d����p�83vE	w�v�.[�w"��rQ�Js�79��yT�(�j�S�+6�ND��M�F�3����Rxi%v��~��^��3N���-Z�ڨ��ӱ
-����A�\t�:��فG_���QF��`�����@�>t������7z!-��/z�:���x�7�鹃6gⓕ;w��HWW�0���l�T\����w���d���6�Uq�T�Xۋ��'-���I�9zˠ$'����D:�/!�-�N�£��F�V/jD�pB��"��(��Uh��K��������&~ੋ(�7UX��(��Zr?�|���CT=�^�k�Ц�P�/��U�~W#ַ4 "J��K|�CY�ي�"	
dT٘Qз��(�R͌!�r=O���f�����A��N����Ϩ��P�+c�o���Lx0�e�;1���,ߢj��uNY�Ki�>}�����@SP� Mn�QL�e��f�z�ZS�� ��I�w
  "���\�����f�,OM%�г{�>�+����pY�@t�nl���ua�*�j��S�9��o�6��C��v��g �W�������ɑ�I0U���@��<���񧰓����Oܤ��3��x���>$}?? �h�c)� �Wru�)N��픴q�e@/�Q�"���b���eM�=ES�C؟��l��WF"m����.��
���J���&./Gè��~wN%h��-j9#��2#�kf(IT�� ��Q&�8E�k�ʷ�$��?��8h >'�Ӽ�MA�]�]6�5�e)���K��o
�n����i�����Ɂ�¶���w���H� 8���t����
��Pл�&)+�N�1��*�;\0���ňK�t�QE����1xd*�w��l?!	� L^�qww��==T���lx�'�׹����9�0hQ�>=|�ӛ�2��Ț�ns��X4�o��Q��Cg�:��i�D�����!��}����C���Iq�V
ν�����P*��������X���y%qǀ��=؄`cV�.�K�w�*R#�|n4���zv���{!Z��:KP�2A~�-(tWOȽyPoD �:�?�S6W���eZ��X�~솇��̧/J.��������Zz�ۺ�?xm~pg�ǰ�U`Fz�{H~4Y� �
���K�΍N��OI�R������z(u���W�ѳK|�'"N�����M�;/�̝��yʞ�['�̯�g��2Z�F�"t��r�BT��o�x�l�ƑI�6�]�<���;��d�a���c��g�z@�9x�=��	�?e�Z:�� ��~�M�=�8�ߌK� @��ߥi--�\��\y�PKCm��p����j�&���2K��|�bb:�8{�<��+�`��#'o�ȍU���<sv�M�p̈́��цf[��g�����~o\�]l��f��_qy0
:���R �7��e3�$���\�t&�����O`&"m
��_�MD�O"�~<��ҕ�MF&�O݅xKE��������h��禥P�J�q���XX���ے��)���&\,L�ڀ�͂[_�]h��lk7)s�I���;��l$��V&'��\;膯�*s�Rz����ܴc�*(�v�ah�wo��t��rDX_���&��|KNt��L�ɉ�Q�F}�	��\i-d2q��r88�w�?ڀ-^�.Th��Z���fVr{�ߠ�Y?�pk�!��o��|�$h�L=z�<�G�=j��X"�G��q3���3z(���*�J>~���*"lҵnS|v���K��`ec?�W��i+
wMf�bG쁈�Ν ��p�qD11-������k�5��c4:���6��0�{0���7h%���1]|'O�x ��1]�����q)�~���$�ʳ�Z��דF��
��[��,�Y�V�Åܻ-�|�#�Xa��L�.}8x.KF@~]y���`��V�<��@:�RT���(���l{k ������y���y���AVq����;엶��ǟ+�\w>w%��^=���Qp��.g�eE>wƛ2�z�ˇ	���s.g�Ќ�LFG6�u?�2��r�Qye�]��R��v�jԍ9�xA_�R2/`��o�Y�ws¦Z�{�7Ȣn�'�r��^�<ägs���U�>�|5ߧBo�B����{� �'����y��9,B z���>ϰe�S�S$<�ن�x|*'���{������W�_�ܶ=p	��
�K_�v|�C�֚�F!;��j7Xh �-q=��6V)`F�F�y�vY,?6	=.��K�2 �x��h�X��>�^DRm&�FU�M)i�Cz�#z�MpyJ(�q�g��,��2ز�q�EW����t�f��y�tio��[��s�t���ޔ4Nm��
�=R��_��k{v��d��	����݈ƹ��(�zR~��I�Ӈ�̖̽q�ܵ�Zg�Q5۹�r	|Ͳv�sԧYb�ֈǖ�T�77s桊�^������r�Y�0S9�·��;�\6�#)�"�ؖ��Ҟ��[դ)�e=�O��R�� d�s"��uWB�CH4�"U��J�U���b_9��M=V ,�q�ӌ)h|~�<�V�zHJ��lJ�Y�s)�D�e�܄�����5��B6\��l�yN8*��AN()0g�t�ș����J'��g?��|§SWA��t-� h&",�|��A�A'���v��a#�n����nIc�s4�'߃����OK��w2hh��t�:ƦFBJ�vq��z��-�j	���-͙���w������`P ;1iJ���b�~$�U�������{���uu	Oe5i�BL��T�d�����wi�=-�[ϧ��V���9J�'�O0��v^ʿ�3�wG�I.�NE�Zs��Պ��୹��hl%�D7`�r--�UT�!�1���n]�n�k��(���\|����#w>~�/*z6�S��qmʴ�:���>�N)��e��j�qݭҴL.�|%9}��>��1��"��F1Y>5&}�X�Wc����!r,�X|�6�0x�x�6�1 ��4�E�.�������a���\8X9e���3(B�̪��Pk'BY�&�����Z$c�T��ěC���ĕ�"b%ݘ�d�͊J�r�Ҝ�W-|U��GZc�3B��m;��m�:Ɩޙ�����������,X���-v�|�[f����`D�['s�3~ׯY��^��o/���]}u�_��Zd�s�8ٻ��豊lq��A�<Ͱ��w�l�W����)����8/8U�>�^x �HVa!�&�u׿���1T����o����������sq ~
����~^!u��h�-���1���В���v��zq�](�~֬����11?��T��ǳ��
��[�R_�ˇ{�FCVHuc��U6�w�-����y6�_jP�J8�]YA���M���`��z�|�W�q#��'jH�[�J�v~���K	d�>��sZ���{!	,��+U�SR�*1�NS�5�����dQ��1�c���ǁ�ޑ/�ݭS���A�ǆC�>u����\�L����%lt�;��(������m$=�]��׺ �=	Ehf�If8d.��{��23aa�d s��D-{H�O���F�`�gC��9�ߞ��"u�E&�r©��oGM�?��E��!�U7�S�
���4>�������myȔ�U���u���R����y�ȬX�-��+C�p��0P�Kv�d&��s���\wW��C��#4|(��r8���L7IQ��k#y���+QQ/T��N?�R+�.�twf��	�lέWk@څX4_F@Qƶ1�J���_07���5}�o��溡���D�t������8nt�G{$r��/���Z_1g��+o�O�j"'S���v�0[�(�T�P�,&�6M��`�#a:��zT����h�IIĕ�E�\v<��##���y�^�A��� �p��	�'m�Qk�ꋇ�/�����/vF[a\�����ɘ�E{Z�7��vyF�!i��	�
��lU�W����E�<����Xf�Z�M4V@�g�/4PBߥBaCa��x7��@/oq�o�x@����p�=�z1��ze��ɨ��8����BM�,cz��p�¿��A��+��ra1"�j�)�L�W���-�u*?�e"�"�%�?d�eJ���º�M?w�
(#��u�T�������54W�ɾ��[p���rzs���ҔB����,��J���/G\@o�?R�Ѳ����}`3ę��՚��)nҁ����iyP��(a;16|`^�Y�
�q-�������"����HԀ�+*r��Y��n��^xxW���oyD5m����o��\<2�KS(�`��Ac�/i��2��KwW&�-������fA*�d�t��mF�u���eGo�ۡ�:3d���V2��m���tdH1��h�XV�oU2��
(�AU�Ϫb�d�ŧ��Z�`?+ӁJ�:٘�V��ahQf��Uqc�A�5F���P�l�}0�'�'�˰$�뭽:(\�Z+L��ӳ8���᭼~j(4��ϗ�-�|yg���]�%��E��{�]���`zY�����ް�������N���/%"�����L�ŀp'�� ��Z��X4)�c'Q�vDN�����
E�g����+�㪗,�llW4U�h�_�����+�	�7`=�h���P���t��7��B��(�UG�Շ���Ө�1<u@�P���y�T��ȐTU+5��-������Z���COH��2J����2������A�19kf[�Ĩ9�k�iL���(F܆e�iKC2��n��'Ϙ�R�&!�U���n��E���.��8NwAlE&Ey�`�M�e3�i�$�J�b\�c�P4�h�@�����v��2���G�JwK�8㶺.]c��`��m��_��-k�נ��[�z������)�!@���	\�rX�����d��y-y��6�kChC;h6�Uy����뿘B�o�R���W����83a�4W���y��nb�&=1u��q���ʗp�[�]p� k,?� Myg��a3�o,6��v�W�HU�Q�/�?[���vj8���yV��(���'�
�����Y�G� g�Dj
V��	����{�<�P����͔<�0LEH2n�� �8��G��e�L�]�}�4n}��& �ʚb�y�A(Wp���4Q?��)�����X��6��}����`	h^��� ��n1��'J]�T��*E�L�9��T�v� yr.�:MԞyt�Y���'m�M�O��<[Ӭ�?�h"�A�P&B�t�`��������!�]��g���#��gOc�zt��H	*�R��h����M}_�ߘ{��8�w*ya�w���>*X������3��g��ǲ$~�?Z_̪����g[��lL~�?��?��?����/�C���RžM�u��`>����r����a��/����E�8�VA~?�1%�j}�K��	z<p�_l��]%1!L�4����P>i�!�^���Lڴ�ŭ2���6YƂ���Ze�p�7�n=�.�h�S�C-�@.�k�i{]ާ$S�^�lؑC�\ᜨv>���mՌ7Th�_8��gX�(-��$q�snҮ�h��`��ܒJ�+�af�p`�%8�T�PT{��!}�8��n7�E���f�H�]���:�PZ�}�cX���R�c�y6�A�{t�'Uh��� �b s>TcB��2+45'g/h���XV2lj�>!�r��e\뵉�����LckG�4r%�����V�<(�J���w�7�Xt���*5�Q�oP(E_�L6�$�#��ܸ*��m��e��KT�8C�UZ�*�NF�E�"���vd]zÞI�p�Ӱ'�3Uܝri�@��ڒ;r4��AB�/O��|TnaE��Oi�}��@�w%[YzH`s����ߣ��R,�I�Tj����d|ҜE�g��D��@��Nx����n=��* #���-�j�+�nXnJ��i	wA�J�V�c��Un��vX4Ƀ���"�\�
V~9jh��E q��a���}�Q�d�H������/��+���a�Wr魼kOH�\N��Kp�Z��#*6!V$U�@�������E�.D+J���P���ɸ3L���]�&\u2E�U�B��_|k��*���.�w��U�Zi�=(�W�NIB�]e���ۻ{�M��`�,!�&KF�C�2�L�����/p�<��7Pzۦp��T�c*�W�Co��(�:I8<E���������
�a��+4lxRw��Tg��b1Z������	�	h!�8��Vr�>g�F���?�)���T+yE\�>��(M��Q&iUڳ~?�J�g�b5��-/QWj�S	D�|]�
3qu�NN�_��ڎ?���4j%A@��菌b$"7�� u��W0�����e����G���%�������j�V��;�-i�E���<keo}CyP%��l_+�$����,��ّ��<��<�7"�C���-|�X�?���rз2�q�8)���r厡݋O�%
��Ҵ�&�����=7ߩ�+4�9st�h�w@?���E'9Q�V3���z+p� �fPjm�qd�;�7G��]�k~=�����13k}����B�3�I�_(���@����޼;��'��T�k�-��3^�[���$�eњ�#�u,�ݨ9���VXs��#�b��|&��s�+����!����6�!�g�
/|�ؑ�'(��{�}g�n�EN&G����9�XWb)�p��>�v]浑Y��*Ьs�}0���Y*�h뎶��J�$���e�:�(A- y^Z �$AD	du�	s3�g;� C���}I'g�
UU����L��m3y�\�oI�8K�4F�5�J�iT:ې7�z��>�����(Wp͇Jbq�|���$ZSq0|(���ń���\f��ۉ�d��B�W?���@~q^�3�]q���=�,4:�'4%8�h^:���a�'�������.\*6LFjb%9ӊ�c�<��[$έ��;���Z�Y����0Ӟ dX
�D��7a6Ơz��7�5;ܥ�R;�Gf,<7�����@�O
uŨ9�@�Z�w��K�eć3��(9�3��xŇ3��|�Ø��$rP�e�ذg��ݳ*ǿ+���0�X
W�h0Qug}�Ξm��_a�m�'�ҜiКz����x��w�1��k�a(�\<N��S&��L�wp=K�<�#XG��3��qxQ��4���D��֞ԏ�E1wVK'U'�_p�6��h��-A땦RΥ���b���<!3.����$?�o��7�Nvy·�|2�]p�T��r48��3QR�h�-��X�uh!��_�������Yk�]u@�z�u��؁��	�L�'��kV��q� ��"��^ $����L�X�$����>���ø������R�L«�=��2�KS��(���v�����=e4	��ۃ|�9@T�e��C�jdu�*�]�҇r/*{�Vb<����G�j$�@τ��q�����/:�*Ш�^~*2uY_�	�G6���n3�z��Y<�{_e�c�D� FU�j�����2���сr2�O����\�sn�{#���Wmw����j����������%��&i\��{Γ[�\���e�0��I�w*�.q*��arEq��A�q�'��`���_��WV���=n}�aD���5x�-
��	�e�׺&C r� pz��	q�<�<�~���#�������U����x�F4	5e1�8g(���t7�}��7��=��>zO���2lZ��x���5����ݭO
�����"�/�WTL��cxl�̏��W�+�a�@@�`�;��/���eܖiJ��t�IO}j??��ɉ"���a��E���;@(��d��� Ĕ�?Q�'��=�k�h��<㞯�c{��`���SRK��V]���I%�'�����a{�)����}��Z��Xէ?J��F�ͯ.yS�=ۙ �����}bI��
d�%��+�����̻AĩS��v�����H沿�Ї?N�@��`ᄇ��|��a*El��E�|��5m¡�Ew!��HYa���7�9���9��^���G��J�% ��"��-y�q��0��W|W�K�gn,��2/��[�O��ؕS����P�+H��b㊅��.QAYŖ񧟅��6�*�L�@ldy���{���a���k���A{�_?`��4{���WvB�FTF *{���[��Ch����	z]�Ri�i�����a��r���5u �&���';��5I
P�Ϳ�0�w��^Ғyr�H�7����8��-�Y�M�8�\�Sy���ه �"X?F�̶2Bq�qW����<i/I)h�z]������^� �A����e}�)7�T�����Nj�.!~aged�P�x�'�X��xQ�����p����w_����R^�P�ul����O��F���"sP:����#��W�X�%��Rޤ������V3�$d�B�d�9�6���APqc��8_�qs�a��Lr�7?܃ί��"��&=d��
��͌Pb,��r��S4ӈ`K�Ux?D03���Q���U��(�-BߗXy�іv����^��OS��eocU��)v2|?��_Q��ń����e��H�ڲ�:���A3�yB�`cb�|�{xbx�w=����Z� �����/~_Ne����t��m��p^s�R�a[x���G�\8�8�۝��4,k�c�{��9��E	bn"6��Z���ن*�g�
txa���">%�B�*<JchɃh�Ȏg�̂5�)�Y>6�����w��q��=Wj�6~,�]�Z�(��w�e�yi �w�Z0vFY�I��wq��-� ��&�=<���D���������"Y�C n<��$O�^<�!<�^���ho�O����u�y�k�2V�F$���D���p��,�	���k1�ѯ�ܪ��{vj@�P�i4�
0pF���;�s��Jg�B�ym�Y�����Σ"�7Ǐ��N�I���3��䱝�6�)v�J,� �i1>H�����_�8q_d QC�3>�鹌L@10Eڄ�.=ҭ�Vy*����ը �+~b��[ ����&˷b��G`�A�JP�4{1a�bF�.���C�P�)�S����>M�֭<�Z[
�QX�@��$\s��!��C�4���w����c��4[ϒ� �0>;K�qE4��:d��G�Z���Y�5�wm�,D��@e�& V�/~�h� c#^��=YC lc?9M3y�‧��iē�{y����R}x����������x(6�P+����pI@��-�<
@���`|v!��ddw�b����Z^�<�5�_����ӭ�x�O�5l����$f�{�%q,�4�0u��P��A=P[@;��?4�C"�"� i�� �f��s�42�0�X�mȳ����|Ƽ<�5�E�`+���#Kת��ϬjH�76YSx��K�M�qM;#9j��n�ε���@��T	v��x6�E��~��������(�n����(O����0��ج-��A����+�Bb|����l��l,l�i�9�_�;�(m�.H�"K����fD��9 �2�)�p e#����?#f'�G��1X��ܮ��b_~
R�4�r����K��E��/f�W^�C�KPk��(��  ��lH�
gjFwLpϰ"�ߺ%�PƜ�	 ��8���V���eP��<K�1�M׹�e���~Gφaao�����1�q��3M�`e3�m�� � Xb�$�(C>ϖ#��L���+������F3�*H�-��}w��D-.U&�0���X��mc:ʻe8{NQ[�q�
rr�ZEҏ�y�c�9gZU�]u��C�UL=��h5	�����3zo+>r%N5r@ ��W2�GDtӹM�pi��P��ʊ�Iۯ4 �&!��ԋʜW�I-mKL�Q��ۦ�<�mI�.PxwnXT��sU%���H��R�� 4����t�9i�Y��]R�*FcmA �(��ro=��8P�t$[|���u�"�'���/E���͸/'��J�W�r����N�T]؇>7}�	��J�Pˍ���l�A�;�]��y��m��єA�,���o�*����#G!0_>��UCw�A���Np�wUy�������")�߿�&.�>X~y����=��VG�
��r�L����v�1%��L\��4�2ֵ���Bqs���~���5j�cL�sDK�C=�e�4Nj�L�K����>�1��8���_�u��2?�â�%5=���K����0����d?h�F1��-�f���\�ynͰԿ6��� ʛ�W��@�#�4����wR���s2�GcF�!�b��#87*ᵛ��j�٥%���u�A>��ε�NBZ���j����`/-�&� I%{(T\B�%J����|��8X�QN[u��F���E�HZ�Z�+��N��n�&{3^���C[-�`��1��Ty�L�-�:����ϸjW(=�	�0mޚ!;�DJN�"׬�#9_�yE�ީ�`��䈜����Q]/H�Ż��^�
�XN�q��nLt��L�����> ~���WX=�=~Q��Q>(~���O�R�7SWȴ��qpR1��ۄ?p�+�_��u��.D�꿄����փKA���@s�>L�M8���J���+�S�h��)���Y_/�"X�]�dEю�	����"��=}��w�����`�A����p
U�,��5!$��F��a�H�b��Vj�M�ʃ����w�F�mf�>�"�)�_���@VZuE����\��c�s�E�vBD�����7[qdvP�l�v�l���#��KΒq�
��K��8%/�ĺ&d��s�%Z`j�����(�P����E�i�.�S�3��ֱShd�%�&umN�8�����ե�
L'O���q&��)���E�)v�}��qd?���s�#���z�8a(�d��Li�.��Yo`�JW������&�������<�ג���U�e	5ʣΊ.�Gv����]�^�����k��8̕�!�n:�iy1�誠.��ʙ�f�P�IFfKmvq1��_��n��;�2jP���Y�+�J$��~b���&�1��g�T�9��R�M����s~����P��*h�d�x/\)���d���f���^��~:�hpg`'n?�9�$g����"�/-"��X�5���w�95g����M�9��k �۟ �Xȋ��0t�HTc�r܊t�"�1�N��dl�F�@����nO��� )R����=9�� ��R���F���ub�b'M1�r)tAx�*���k��>t̿�A��'[)����VI��t�y�	x2��ϯ����:��]��A�����8���w���8��<ɝ���������p�'��d��2��C���^��g�e͏��!����m��:�Z�|ܑ���M�Vq��VC�,<:���<�8��1W���.�5G�1��x���.�
�
�0v����?h����5c4���8�W�v*�b�g���D��ϕl��+��qCs���Z����� d=R�Q�6�/�"�*���=!(C=�.�*�L���M�]h-\�2O塟���C2@�B��9�����ܛ�*��n&w�V��c��#K㌷���R�����N,���NH'���{:���\Tj�h�q�FI�U�/�j���[}��9�+� e�<�Iqw?%b�tg|�:�|�ꫠrI����zŃ��	�q�W�.$���.���YI��)�vĹ�3��*:����^����u�y��A#��WW�f���E�%��08�� ){���פDX|�l4�d�$�E��-���\mK��[����ص�$�Ү>%���5'[������Cdt������6-��=�k��~��$7	J#�?��gHC�QM�qb���-���g�[L��9p�zZeh��@oL�Q&��Hj6����!��"�9�ڶW�J��QZFe��oOe�(d\$c�5�,ET3?'.�55`� �FK�e?�{1d8���h���>�$u�/�H���Ot��Nyq#��~��W�;��1�G�+EY(ɿ�Ǆ��d�D]h#���*!�Zŀ�qt�^$cY�{�W��h������وN�"h�Ѧ��H��G��2����ŞX"0�vD#�Eռ����/�D]-$<���^�^��ɼ��9=��(�[�Wa��fcd���kG�"'OF&��P)�.��_�pQ��t%��8��,5�my[^�:��1��Qh�`)�a�c��^ϛ����=W2���8�!�8�eQ����0)JQ�\)pp��R�Nߑ�㦪��S�̄'s�|�����9��!Ew�/�!�pw�y�|���w�s�nz�|1%����z�2.&*�D���F���x�>OT�Az)�=p�c:�aj2��j�7H�2n���2�G�=^>%��F�.��,�Nk�N��?�?��n�&k��[py3�˹5XY����~k����:h�Q�˄c��v�H4�J�j&�Mtc^�X�MNxou�-�C�7�+��/0ϗ
b�Y��Q��F�|���$k,$!Er٢r���fMB��Ж�����rה���Xk��j���f�g�����%=e*B�m����ȭz�r =������+�g��T�!�2�d_�ng��WBz	4ًi�ra�p&��"[��6���_g#Y�꿗��0w�vB㘌g�R�"/we𝕬�R��l!����!���u���/v�QG=(C�c��ϗb�����$���z�Jûlk�G���^��"n`�V�X�7�;�2���1��s�o�y�F����oG�~7DW��#Ty��X�����*�
)
��Tm:)�y@��rgN�hƞ��%K�L-[5�П�IsЏ�?�d�̖_nN5%��9p���깚����tt���V0r�, �l��%���$>�hL���3�������Zq���4?_��I����	��� �x:���u���(T^4�i�\@��d�_Tu��:5<��<r2�C�{��`{6$�7W��F���kS雄�H|����(|���>!�s��]�Cf\3Wo�1��>����gƐ���!g�>*���h�P�x�d4<U��PUw[,���B+l~Sm��d;�y�I|��W��Kk	��XHF����&L��E7�y'���9 �������\��&�ח�ʟMZD���抷%e�YrO�|Qy(�Y]:X����ʹ��b��j�s=_��lc�5|:���uL��|����^~r�!wN���*���/
ZL�]����6�3`���i�]ֲ��-���0[�n����0�e\4��&4X����K��y�w菱8��������������f�?��~�|�����W��QE�_3��I�A�_�	�gg�Y����d��P3{a�� ��~�.��EIBS�>�<
z���-�-�-�)�[8[@[HJMB�7
p�Z�Z�S������Ak�k�zp��K	0$Г�������)�^�)�S@�p�����j!KBԂ�!z ��jaj�$�/х���"����E΅�����/<8R���Zx_�Ф�I��--$ �`�p�����B҂�p���r���;�!a�|�C�%	 %ߗ]���P�x��z�X���#XC����FE��хb����x�H��c�K᠞�.5&����B����[3=�QЊ�1��NY��H��g,��9"~�9�RXl�6¢H)�DȀ=H�2ȭR�ڇ��x�j����o9D�.�:a�z6��?L��68����ݒ�֏D�v�g��5<C�
��p�p����knq���#4B�,������1�j�2Ɨ̌�����W���X�>*�-_@	��:q ��2��h�T�'!3�h��ě2��l�o���]�
hL,����G��00�<n=���&�����0OC����~R!Ӱ���>�@cvw%y*ݡ����Z'���sD_�
P2(� �_���*>y�F,UG��nSf�;ㄙ�x��$�tc�F�ռ��T�<NyO?Xα��?���LO<��l���Z�Gh�l mH��gҍ���H�
Tu�������/"��	�]q��rP�"6N�H�G>cxh��[���@�T�����]F�鼙1L&���Ŵ�O6Ԅ(n������77gb�$eQ�jvޯ)����)J��$��7F�Ui��6L�.hH*ͬ�b�h#�L���t&v,���1�4��
i����V��h@�,���Nن#�E)��������k;ؔ�6��^3�2�N����~�K�OZ�d�����n΋�.	V�?��Rk[b��n���ht/�$y@*ݤ��y:q���L���@��"���$�A�1�v�&����w���(ȶ�Z�a����:[�Yr���KE �Pvt��M��֛��Ιu}���3�ZoR{b�$�	�_ls���	�MO���$������>�*ĝ�˥�s�o���y4f�(��i��S��i'`���=v81�O*�l���g��>j���K��l��جRez�T�IH���`t�/x��,��������;�\�#^l"iM��8�73J��#�'��Ts�dٷ^����/�va�F��H����{*���}}w�S�~�Jt��T#/N�
((�B�������F�	��s�"2��6î�NܣϪ��Q��kW�N�`R�w�G���|9x��N�%��� m���_l>vтpv�=7Sb��ZCo���c�����,�`F�p�PvI�ʤ��u2�C�<s�嵭 ���v�7�m�P�;K�j}��<*�e�׼;/�.�{Ԋr�5B�@/�kd�,[�/BE4�\�ĭ��+��vζuzH����;�_������iV��?U�j�nX�1s���̪�?�-pG��4�ɩ92~��$Uk\�>���A!�X�2ǘ�`f@8������
�?E�������lmT�:�9�:W��C��\�L�7�wp���)jN>i����u�W��A��A�!��<�D(_I�Zn����g��PW�'�Eu�kǠ����g/-X�r���y=����a�k�>m������� ���6��X�x����Mm���v��ty�7,��ӣ`2�{6��
�j����A�'6:�M�L$�h�������:�?�~��Pj�&v��<qN��9b$�yK9�.���RB���@�����y��:f٦�$ʜ,i�-��p�I#�[��V�t&��J�O��3�K��ݴ^�sD����7 �[�<�}5kWe[e�Tc�&�{�
P��R�F���G����'4B�+uU)ף�"w&��7s�fb�p��?R�@��S�<X%���|g ������,�I6��5��\�Jj�fg�m�:�JXcU�e����Ӡki��� D�\`�%�n�k̈́Y$�c�e���P���,����A����t�Z��&$y�)�;<���ǖN8�jG�;�s��M�����_�����C'x {<�����I���&��#Lt��k���d�虷�Zx��Y�:��H|�{�:_�������e�Sy���`L�Y����'/��O�z�j^�O3��/k�>g���<��]��Z$�� {tCW��yd����'��tƙ�%6MJ�Ԁn�V���5)�č({zbj^cTj^����j�x	�J�sq.�P���Q@܇�H���n}��gte_f'm����7vj�XM0���evb��x]ZE�i�����F��݊�S��p&l����w�����k�x�ɉ�5-d�Le0J��q/e]�4T�gg���naC�&�Q����S��0g�� �W�Z|	��"
��>��I�<2-�I�2v�	'{9%����9n���IZ&@a�NUԕ#a�e�F]��bM���.��k�?|Ňv�n��:�\�×�!���������ӷ�rf�p6^~fkKk%���~ZRyjg��L��_ȯ<|��[���&
0�����#O(2���"�D`f��j��l����n��92I��6� ͳ3�����������~�'/^��?q���U) �Z�GGb���6��4FZ�o�B�1j���}-��J��'�,�S��R�Գ7���U�JͦSaܾ����	{A鄰��0���W�B1��*�0^�*�_詎 ?<8�����jJ.6)����cu��@3�:;��)
���Q�n�:iӂ����Q[��J~�-�&�Z�
n�z�0LJ ��4%(k�ِ71�ɇ&�(��Wd�@G:���W�I�(3�1�_���B�=�V�Ev>��rJ�O��>fvl�t*�r���W���މ����z�0"�.�荐��y(v˙:xЃ�j[ؘԋص�+b��A�q��`&ޜ8�pM;-y�ʫU�fB���4#o`_06Of3��Ǯ��G�
��]��m!Z���&L���D�(z��V@��<����r��o�_H��gF��7ga���=rlP@��3��������b����!�C��}���-j�6��^n�����+���)A����ƈ�ȭ��yV���-�����cE%�'a���$:�oM/wD�;��E�s�V���X�m)_�y�r[F��&��a���)�>��7=�"���C�R
ڍ�G	9+�iǨxvڷ4� �B��u$�:}A�Q1݇,�P�,���g'oy�w4_w!з��,�xYz�7V���?����Zh�5�.R�L�B�<��9$��\��<ai,52���(��ڦd6��Sz�}|��U��ޙH��W�4W�H�����	/���K�dy�9&�O���j��Q�u��^�jB]c�`Pl�k��_���BI_d�|��D�rt������/�veB4�qYP7�C�����"�n,e��l֥�R�R�&����	y��F��Y3�а��!m3!��Z �'����G��\�2(�����.+юB�cJ�<��?Δ��V��J���Y��
��&�l�u�_��]xC[�Ї6��LgHsD@Y��9��̮'ڭK�j�̶���*��b-r8J��g�!�dHL����m�iXs+�lKSY��Y��P��.[i2�Mq~ΚΦ�I�I��$�u7�!�`l�T��78�y`�X.�u2��	��m1��^�=�H��&(h�I��i4g���i9	#Ȫa�@U�*�p8��1�eYId#LW�[/�z����MU�8f�����`i!��@Y�� ��w@��Y���×&&��8LUf�cT�uKf9���EQ�Ҥ�o��Xň5!V�"h�,}�LD6	��c��FM�{j��rpPL�%���vT���.�O4[���\ތ�|�b/>:C�=�9�z�!��9$�GE�g���ᭁw�b�d��idW�%�Mߗ�����_�G�
��e'�dP.�I �!̚J���� ��+ǛF�oݑR��u�♾9@��$��I�	z�LS����#�,y�jLX�5�E��;!.�qS��w3��6\�ڥKfVS�V0y��e�0~���v��Z�@5 x�%)�t�dX������莥���R�(��E�����q��c�5ֵk��E���F�X[N�Z#��B�l�#lҹ��-�9.?<U�b`j:IM�;
ʴBÿ�s
� -�,BVY�Umg��$waW�R�󑢏K�:u%ש�7����'���u�����֢i߆_�xe*�V-�Z\j8�`���	�6$N��(�y�e�Ev�!���@[��t�e`���M"T
�b ��@B��M�GՃ[���E���C� ��_l����[���>�����h��<(��<\�q*�j�����;#iʳ
t�%��?.Qv�K��\�D~��`Ϸ¢ӻa`��W�[$�.�z���Pu�ĩg~I���	��p�2�Ď��,�X�T#,��#%-҆���=��K�^�-*-\}[=�*���6�!�0�FaT�����UB�f4�@e�����S��һ��$pf�~ރ�h2{����;�!����Τo��S[-��J�ż��1h������'�!DQ(.왹��vs�ϣb�R����.�~�, b5�cs`��6���q�f���o�jX�M�w��/%Q����S��,��	W�=m`�Ṇ���$��CF���b#���3��	�Ш�_�5�96�|\�������9�z�^�`�h*Ÿ�S��9�ƾ�
��-�FO�j����S���;�c��GY,�KE��S�x3�퀸j�>��ٺ�S~��B_�ϥ��^�kF���(��7)��J	k|���zT���&PJ���1~����
�X�(�	��.�~Q��CS��'�\�rG�P�(�(��m�𿥵2����!��H��I?�2��,�m�W�`�2��Eݫ5�9<$��9�)�ru<�BI��&��P�9�Y��Z��`���3M �6���,o�A��!!�v�=:"�a��zR�CU�q����z`
,F�tk�����R���il��1��z{)V��>����Vq@���&��
$_�Jrb]2��!.� ��d���1�����mNN��6z@P��fչ��>�M���ɽ���p�f���(0a����T�q�Tr �o���?\����gD�e�Rncg��I��<*�^rN`�J�,Y	���=�u	!D�2��L�+��w�V�/�*�s��Y^�c�E4�#�����ѤA��-�r�҈����?e ���Tūݞ ����/",CF5���7���A������!�4� ���G��;}c��-KPn�q`�hB.p-p2��E�����F����Z������X���;�V�/�݋0���9 -R��k�H_���� MWd�u(69�����X�~����a�^�{u��sK�}�7���:Q+��U�|w;�;&���B&��q���pY^T�D�!^��X�UeM)���L%��"�h
(P$�h��˂��K�>1�4�?�x�����Q)�d��ܧ�aw�&�5�3��4(�g���ͩ�%�E1�05��q���@@5���V+0"��ԫ�{��{�oC�`�� ���Z ���h�;�R�X�D�RX�h�Z�d�:����42S��ql�N�?�~� �Ѯ�n� pY.�l�Xז���(�I�jj��|MmFC�����{���P�2���a�_�Bf����b�t<B��=�e����, �]�E��L���V�s��3 �Ӿ�Q�,�����䄳*����/���e��ͷМ��`�I��_��1�u���{�{V��'������|0-�ac�O^\XAJn�j��7�n�/�弪�J=�;[����cN�*5�\8G��Auj�l(_pS�v2 z).0E�و�6]p���z���<���Sg���2*l�9���V���s#�G����kg��0�%��uq�q���2�ЧJ�2U��Os�l���@[��x��]>�*}���C1��f0������Y�g
��!�����ïk�~�������qbS�|�B��r��r9�B���rʜ��j��~��9�;��j�W8ۧ Ĺ��L�%ehTT���1g�ҭ��g�;l�u�P���H�"g� �Oyc����QWM��B�ܺ�y]0�1[PӲ�p�!����j��a��\���:u��0����]@��h�٦j-g�������	x7����n��5Em����\�x����%��L���m�;v�1h���2G:�w"���z���N�+����軱�����a���.��7;�[�.k������^$m�]4l��>ر4���M��}�|�uqg'g��Sz�th�9��4��;��G.
*�S��Q�VC���[�@S0�D�v�F�XMՀã��^{b��oٳy�� |�/�|�B*ض*���=����u�^.����f�4��ʥ�q����߈��0Uݳ�!��>��|�L�vAd�:�������7��)HFo ���Yn�E����>gG9'��ZE%S� ]�m�m�����h����E��훉"��t�=qI�w�����膍%b8�<�0�	�z�&}:3��)ȱm�a���`�!/Q�Pk&����=��L�i@���]����r���?%�A�3�{`���fBr��P�ͨ��#Y�dT:��)5H�����`�ծqs}�ڟ<6VMA5=O2�z��3�;���U}yM���t�
�ʹ��t漧�+Jza��ג�'��dJ�U��Jy��i_.b�\���v���WFt��cE�7��P?��t(��8��
g#��S�p�&ԍ�1��J�{C�P|�:Z�6�~iT��Jͧ���5�'��a��t�Ź�vd���sh	��z4[��D���T�?^B���@ø�sh����P�C�дm�#4�J�N#/��f�C+�Gdj���N.d�)�����.&9�6@S7�u��(�Q����.�H��x��Z� ����U����2��pC4�fs��:%l��i���Pt��.b���y��i;%,&1��+��E�&LҬ=*0���d�@.��'��vv˃�E���7~��#!�f*�#�hG*�y:�fXԺ(�	��8}[(��D�t���щ7��GH���l8��1����ȏ� -<g������=��L�i���H���l��yn��DkҀ(���1���P�����&Y��$�b׸�w��y�'�n~�����g<fiÐ�h��7���5'�7&��?�2�6oqQ�[P��~n��w|���bũN����h0�c��(�gߙ��f�S�fS�xpɷ��a5 ��n��A6>_��Xn�/W(}*�i�0��5R��,<3-���pOj���[F�@^���:"{�f�&�2�Ki����}��9o�W����:���_=?��)��+pA��������}7�S#���Υ���hh�&�;�δh�ð���;��R���+ɞ�@a�I��j"k۔qZw�8(u5D�#��$��J*�x'�T�ߺ�����d�<+�@?w�yӃSqL{��1y�L��j�^]�V�u�h-Ҭ��L�N�C�`�L��S/�&�L>�l�L�ê�"��A��b�04�%��������FvG������1�w������Ö�࣡)t�aw��M�'D�幄륈Z�tl���3���zz�iX\�N�jΰ}�*ݝw��n.h�e��x�-��s����x@
�xa�_����E)8x��9dd>�\M���:������J��3g*�2۩AE.�t�I �O�����HD^�b\8��Bfd��*D��
xCYT!E�t�	I��Y���:�ˏ�~��\#��_ε;DGDf���\���l�J��@��UD�	�]�F?�C�o�mhM4�u#6�d8!�'�9BU
�֧�*4���f0���A	G=.ᜆ��!�F7�$�H���KX�lEϝ���?��f��j��g��u���2s�r2��a9n��P��$ x�� DN0øH���s�O��BS,(q�Z��)�
�	 ���W �A�qpR���d��BV:1���l������V볩D)]������|����r��.���8]��cJ�H$�(|j�j���u�%}�<�� tw�o}�a����zl��q�q�?���4���!S���v��6�6�8	 5i��=�aX��[%�����ik��P�W�{�H*gm�F��n��x���Iafb����.0]b�kd�&\��J��@�S��ow�N�Z�7K���jh�r �^>�n<u�.��`j|�VC�����l��d'½��8���I_j��T�މb�P��mw�h염�Յc���,�*���ˣM�����U�%��Oe��*قO�Q�a�����J��y95e ��!�a#�D���4��W��ގԹ�GTG},�Ԏ�tNb���%���/�ʆ}bf2y��T'"ԃ��kO[��Y��X�fM��?���%�vB}*��U(Z�:�?).�vP �����f��&�*��O�6o�����h��lԩ�S^=k�m�d�kJ��*��i�R�XGbb"�ٖ����~��:�}l'HvؖƸ�h85�Ab S�}{ב�K(ƭ��K]�K�ʜR�^�6@��%-�ƶ1����>��p�d������h��h�=�h��$10�W�T�^Y�P���&�ս�؃�`!%�Z?�M7���6V	kɃ�U\�C��]6N�rT��� P���%
�`(��BP�kU%Q8(�dd��5 ���|#�O�:+��m��m9�l���C�[�{�M�Ϩ�-ʆ���Paa�X�DRr&
�A85/�_҂�A�̎~A�Wߍ>��=6J���y:O�Ƥ'@(<ʇ	eaM2��o��o}��N�&F�Ao��%Ÿ�-x���ʆL�^C�%P9v9ШP'��皚(Ut	��^d{%2+���]m��p�7��7%�+]�o�W�X[��|��@5��bC�b���h�[	�N�E����|fkF+S��Hq�1\a!�v�30>�8���)=}�4U�1��쑯/��i,ū�h�Y!���wӃ]��ݗ��|�PB�a<0��,��-^�8DP �x �p�1A���EH:�'ӥB�������%l��4�kA9p-�p]��z��k"�.F�,"��E�dɌ٠��l�}ZyA�����^�a��xJ��I�Qt9M�?��c]4��aw!�[w� �Ǩ^�U/o:�
Z�_SAw�%�x�̩��z;��ĘE$�$�MN�l�}���rw"
��S{#6�.]�	f�WhC�:X�̃X�?a�Bc����FRa�9a�P�[A���'��*�H���]�$~�a�߆\��=�4�y�h�[�u��҇჻ik2�`R��;|����a�Z_�!�b�S�����"���C��_�}�S��rdps�Q�{�(���J��3±�J��̵��h��q!u�p!���$�~Ώ[�k�6D�dw��O��80���a�~�����b#����\>\��%BJ�܎�s7��tv����Okai(��I�KK���${c��VULA2 �g<R��K�̱�B�/�K��̀�]{�9�����5�œkGr��N&�}ǜ���pk�R��ߥ�ざ`T���[&8�\�{X��lұ��(̭.Ȗ=��ssF
��[PŰ�#j������<7%`6Qp	".�'���6H�+w���;D!!��b�߸�a�1|4�0d���Q�ty�
2�UB�>��O��|��c�0��*G��^�%�x٭�0�,�ލ��(dd{�'�k}���+�;�����M�w}�.'3�j֯��e��ƋK�Nrc�អB1n��7WQ��	&(ZGGݗԲ:(4-�!�Þ-h�c�v��o�r|���d~�	:��Bڀ!���ܕ��U���S	����?j��w|7̝1T�I����|&7CЏ�ja�al0-�����/Ж��.7����?����A��]��x5c@�M!�z��V����$� ^Yr�C4	q����{T����6�\�u�T��Q�F{����ɯT�즲>��:Ggjʬ�x�r8�` ��{���� VPO�m�hעn���} �w�M�(�$�$KK�7�~���B��^��@�Ihb����,���^"h�~�:�+��9�lܳ;(�1��i��N����Q��rj�^�4dCE6�&S?��F��fE�=<]�b�^I�����p!D��Ӌqm	��F8`%��	Wz�A����pI��2��N!A ���)~@*g�%����M���F�"������'���h^pـ�պ�B��s�pwdT 	�S�� �\��-B�V�.����/k%V8 �ju�@킨�lq�!�iU=!,DG��VCJ���r�P�.�=�<��Ǚ��qn@+��c�����r��j���Y�ϕL�Fgꀾ��g�>�)�S}+K&Q���'�eUϻOҷ�~qC��r��&����?�#��a)�p *�6����f��Q-�+�#���sj>�t�6w��\8&�u��\L��o������iht&�I��y�?���C^-���G9@Žye��8Fi铽�2=cI+�|�UOf�����|������T(r]�Y8��~�:�s�O���ߍ!�q�E��J���N6�� ��N��U��x�D��# p}�&�r�rخ0�'���H�g�E�exN����������V!�.#��eBU@��?F����~�d�F/�:����q/�o�U9��U4��±[�	�[
�~���#��J��Zo���Q��/M�(���T�v�4:���0F�����y����6�n����`MS-�G)GU2`<ͧu�O0�v|�q���3��<�Ii����ӊ$���(75��e�����P�����UA�����îd��8�c��`�}s�W��{�#���H!%m�e�,�m�6 �|�a��a��0�k硫'���5v1��-$?=s���=�}l�ת���D���lWc�fD����?�m����O�G zCfc�tI����E�v�
�Vm�ag�U���b�����DߌgA��	e��Ϗ�
�����)BQD
hAmB
���-�Q+�O�z�f�~Ec�YsV�p
zI�wE�M��P`��~9�a�e�Uht{�L�?�8sZ\�"�TR$2c�'�i�c��*�IAh��ǀ�s��'����^:<�0t�{V(�5b����[�+v�K?4�䭰��Y�bL�=�#>]�z�b(�F���eIq�b���絷���d�������LV{iCk/�*6}���Ea�� �� X�-2U&��6i�#��A�|���H�ҧ��\A�l��z���q��<��IA��9�ً�Q��Y��x��R�������+�@��݊�A0�� �E�j�p]����vp���~<8���2��d ���e���� ]�=�/s?ۻH4P?w��V�A�|��H�DK慨�;ҡ��1ޟ����78;��ڡgvp�R��7��dCsd�&D7VfZݪ�����<>�����U��i!��{|�<6����{���Y���d�_�5V��.��𳾰�����I�-����	��E�q�D���^�p*7'�����e�	;4�%{0�|�8�L���Gf"�s���XܾP�	?�)��Ae!4�R�>t*�\�|q����M�E� Ǖ��F�h�h��u�d��a��b�I���j��_�ix�C-�q�-��l��ٮC>��6I*e�ٷK�j�+����PR��R�� fH�S�z�?�5 �s��À�[\P0;�@�-���pt��ϑs���=��}!�}�q�I2=��g��n�b��z�4\	n�{�0W󇊳 �gU%�M�D�ɐ�m%	��R��/*�¯|Z:�+U�?�:�LAH����|���_-;���n�X��AJ��%��0�����̟�(��Oc���Y��̧C߇�SL�B{n�E�V����}�l�Ǵ���$�q�Q�^X1%5��l`��7����I�z��|W.�(�$�?iC��)2��$t�5ahH�Ufv����	:�=$"�-}S�Sp���Sh��ebHCun<h��M���N��L�UD�H9�fyڕ�֠ڪ3(9Hs���̙�<�G1�w8OB͋�u��w�� B��y���g��e#��-)����Ϲ�'_N�X�trK��&�MR?���1P�� F�"M$��2�^{�^� �ֱY�A���R璕f~t���?1���,x�#6���{�Z'�H���LՍ�Oޅ{_�E+N�7k���&43���Y�,��s�d%u����'���VP4��ެCu���ЏH�#�$r��mꕆN^6	d/� Sm@l�GMjFǗ����ז�O.�������iª�S���������s��6/N�2dl�}:��Xt���/�SGl��ww��V�����I.���:�f�_��0	�+X��g+Z��)tCo	�g[�r=��;h��#�V�A6�����G�z�/=$�w<ɔ���9X`�dn�ȼ���7{z?�ms_K7��'��Z�t�$t˵~N�+��\��<�
�� {Aܛs(�g���y� �� �A�W�)��~�3���m����J�N���vo������Y��d�f��,ah��Cb_E-2�~+��oXX�e�e�ҴV�?Xċ�72-l渓���d�'�Sp��/F���7�ZS5�� �m�'��E�,���7P��1$?C5�夽v��<�>��I��?ޢV`g��`�^Y��	���?��,�1��P�����./i,�)c%��*	��_��o��e�xZ-���RԬ;���t��&_q��pӶ�K����;��B��opy��Ԫ���{�����A��$����`�V-H��h�����,���5<�:�z��F��-��/xz���}���N������v�~�J��3��?V�Kdyo]��,M���z(����ҲuM6k�&p��Q�X��P
�,2�}�I��&W
8��G�>OR�e�|��?��Wxq�­�rw�Pk����}KR�؈?�a�'�`_^�g�zP���%Q[��ir�'k�sl�GDRY=�e���2��&xv���H�).���g[V!�q���A��p}�p�键����ը;����(m#i�^��3��p(���Q����	\��j�7(�>��5�M��{�h���[�P�G��n�*�o�{z6K��h�U_��
�^�0�u���� ����i���V�N,$/����~:����R��i�a�/�n����%�e��7��|h����l�hຍ�������m�Tq	�$Ӌ����y\˧�!	�"��ch`���JƔ>��"�lAj몎�S��[K�u�_��}��(��vW�]߸%�_���V\�����v����#0�������
}9�Hbw�'���dЦ�}�>�����_������%�ꛆI��3��nz��և��G��Dˏ����sLF��z����9'�nj�c�V#Ɖ*���e���ykrO���/���$ft���v�D?�
�+�t>��䨏X���Nz\'���ë�w7��?��+;^�	!�"A�?Y0|�Ij�NߊΥz�DQ৯�n?K��ǁ���̵5U����9>nF;ڝ-6 9E��7t|�S�6�
�0�t�����"i@ǯ��"�c���_�,Ȋl+�`,/rJ�����A��28ۆ�|.������iT�;�ޟ�-�:����Ϸ`��SF28��M���r��[1�&j���e�8�Y	v�'�i��yQ����Ő�G|��7!�� �\7{Ө('�G�;��<��:!��܃8��}��;ߦ����$P;a�yܼp
�^p~iq���!��s�&�xl���~`��#%]��-�19a��k�GF߇]��|]��/d��Љ)��G!�>�̙:��ƒ��S���k�k��T|�m�SDǃX,����_l�($��ܼ� ���%˭��z�����7��p]
�ch��~F:>��3�\)�-������|d����Mцi�玈��r�B��]�AZ��L�B��.�]���qf�>Y�f߫��
D_�䭽�U6�9��N��k���h�6?$L%� 
Ud\����Ms����m2U�g��"��j�$t��lGEƁ�/�����s�ϗ������=֤t���}6�nGk��]�_�L�[ɬ�A�v*�ʙ	��g��۱�F����\z1�=�Vf��W�T�@u"�rl8���"sϛ�$@��Ӫ�}#JbCj��,6e$�`e� �Ǭ��`�u�0K��x�O1���	���أ�D�M��}��b�R�"���y���^�y&�o�J��93�E븾_�d�%�@M�焑 ���=3z;����N��#$��Yp��2��U]���$=z���8䄰�ʙ�7h�x-ǵ�Y@`R�2��=�+*U~�FO�2%�e��=N�u�(U�s2�@�U� y":;[O��UTDp�؍�����{U.�p!+�'�h���bb�۫�偆��V~!��]ЄB�V"p���ib��`f|.�ӻ�/�>`�5�IB�W�#N��l��B���"��E���>K�ٔ��8Z�����^#�|O�!�E���q�H�J�Y��k�֎_�՗���/��J�E;(�%��,Y��wyQ�r9� P�[��G���X=/H��6� �]�җtC*HP�b:�{C[g�����F=+��=���ڛ���}�-o{��YyS��J-��!|�r�:����H������`v�6�вv��K���F�?�c���5�����SiI�O`%���r�C������4k������wX?��c6�0�-��f�Y)co���Q�Y�p1�:G�����m${�s�
��Z��ג��̓
v�p�{�:��ڻX-��7g�����d6���;����Ѐ�,�<gv�}����^x�_-�1�}ߴ�1۾��JNϭ{�$�{���,31��Y���׬�i}"������Kv� ����j�2�޸J�������'�r��"w^�'o��[����
�ص,��J��C#��Qm������!�L�=�F*�W(f|�#yJ�4��/��9�u*��{��O��(B�e����~97p� 2����յ��g�V� ��ת
Y#�}�ȇ�,���Th��T��	�T�B��^ɻ�R4�EԸ�֕C�d�J�D��+|5VĐ�����|�)s����(^@�9�+.`	V_�>)���&º(�z��w:3��:����8���5;?i>��䠅!ʼ�%zT�1I�����d9=�"F���B��]���� �j��H��#	cQò�*[ �j�����c2nz�B���#�,�d��qI�2�4���8��@g#�\3��VKg�Cn���yJyؕ ��O�)T�b� I�{�pS4,@�x��tђ4��i¾R\O$��+ޖHa\<P�h�횞S!�Z_톔vM���T�#��dWV��
Ƚlժ�;�: ��l-r�_J\��;���>:��O��@��~���G-��,��i\L��{���d��f�K�;����*�����&��Q�l#�@X�����@�4��d\������*&8�'+�nc6E�������u����fr�T9����gH#�g�3�8!��V��>�m!��I��o�x�$�Xd;�F�R3�/E�����`=����\�2�j��Z;^'�V^�O7�}y�������-�\7[��I^fBa�Nbq5�0�3c[�{�7�fwh���Q��Ԅ�=If�8�6�7�v�{����~��n�m��;m�&�in�n�6�g���iշsk��cf^�Q�瞼������7w��a�����������\��1����%���$��b���'"�z�rr��6r䡤(ͳ<���ʓZy���{�=��
ܾ�y���>�%xo�,�R�xb��T��ϰ2�h$�iΟ��]��� �CW>JN&OP�M7�����.�߰�,Yh:nzj��S�*tW�W�f�����UJ1�j�⢋4J�b�7kD��wj���*:��O����~��a��727�+�d\��ӕ�̜$�V�E�}9<��Q�;&��8z�CK,����wm��M�-:�4ध�$jlٔ�7'=�cA���.���6?���~P��їX磊�a�����w��hdO8���J|�C���s�*vP|`<Ǩ�m�=�7��wB����.��nAxN��1%
������dOoϢl���G��@ml�܊�Ikc W���$��|�_��?�#"	�d����L�̧�z�04��)N�9�G|�k�eH[��[?e���r1�{5��D\;=�Ƭ7+<�}��Պ?l��v85Ꟊ��⧥�.��ϯa�����)�a��OwP!����QE'�H.�s1\P�H�d�LIf8i �ge��0���m��z'TOu|% T*q�A����1]�1�#3C	�l�F��G,�B�V��˺q'Ѱ�H�d����������x��U������'���Sj6ۊ�m�����璛3 ߺ���|)ޤ;K0���n�F'���^Y�8������~=�~����!��C��F�<5�ْX�&��b��}�)��5��V���LĀamڇ(���Uf��;^��/���	T�Q�\"h��?��zgر\,�O{'��ٔ���xfBI�P݊�6RԿ���Y,7�scGQ!r$F�33Y���v���B��m�{E5�hU��S�î�˝���ԙ2� �<���`_-��i�s�ꅒMk�ǎ��~{ewv�砤J�na�~�+�2t:(�e�j�8����+��gh���+����͡�(������ ��Xѐq�B��s���X���z���$�ஜ4a����3�V��k��5���#�l	l{�Wѻ	
�7��G0m����>i���e�E�Wx����&�hɞ&4;-��ETx��߱)��O�m.r7�D�Sd��w�E��?sBާ�ã�Hv(���W����e�/��~�+��ަ�V@�9\��>d�g��?\pE�OP�s6z�~p�7�{��^�۵Ob�-��^7y��o.�!8��ģ�#|�`4�
}f���?,/$�(�,��}�|���u�k���)e����������l^6�Q����@I�%�%��Er<��LYPꙝ��A�e�V����Ī��;�8�d�Vt�=(�,���zaZ�;�Y��{�vUY �+,hzd=�= V�	�"�x� �sM�#5�f�?�D��R�py� ��ɸӦ��ʰH�vf�R���Q=���#f�Ϸ Ӻf#�sɡ3ݷ���D&P9$�Z��%���Jf��fKK�_�	����,:�����L��Q4}^�S�4��ӡ�������e"t/�FHo���M�޺�}NM�L��ͤȩ��M���7�O7���ߜ�'���x�|�gnC����yL���"S��:��ߖ[+�u��������ɳ
�$�|M��B
9�e]��s�H5�`dǐ��MV�u5�|W��X �>���T��O��qZN�B,kv6�`:
�3Cj�F��]�^��}��V,���a�Z�q	o��,�Ϩ�Y�1�S��^3[���e/���f���zdIݦ`�_��/�k%����Od�,�33�n�(�E�z���y�|Ood�@�����\�]EF���E*��3MD�/^(��AqRz����z�X1��Y�ӻ�X�޼��M���0�Z�	����\���N�o�t��A��28y
��� l�4��8tK��:e�|�I�%럮��=3i��l���U�G�8�������;�����Ÿ�V�/��M}��C	4�E�:df�a	jx�V����n|�����z`u[����O��5��(C���r9�l�z7���2O�=��nh4=8��w�|l����kN!nF�>��Cc�SBhD�I�>&zL��3�g$ƓLY1D��m�I�_'gc� M�9~7��G�5��������d
ɒƻ�3|^�5���f��v4K�'��Y�񻂚ї5��i!,o�"|x�%���������x�Q�d��WI! �x�Kx��@�6 ����rJW�?@�_���)���d�y�#3���y�B%�.�o[e�Ø�;���ioI�>�sȂ�C���������	� hf���jF�XS�д`�v4d�d"���DlW�����/��k�sLK�� ��_3�Ώ��f�GM��
�� q���Jm�k.��@��F�n^1�ɎwФ�l��˱��@��)'tJ���8�xّ�rkǧ(ԑ�������/e���Pi\�G�)j1(0<r"X�S��-�KE�p(s%Gl2�<���Azhfi�%��1�g|��%&��(�C筹�
���%(���㪞�Kd�	G*�$��i~�O��%�Ȣ#Œ@�k�_��E�����=X=d9�z�s��A���W��ƫ����X8c��p�y�[`|���-�#���OI�c�t��3f@'���γsuwj��r��Ki�_-�uI����8���E���uH-$�$�$�$�/ �.� �R1�\��)7��X���vn![#�������|�[��u��m�\�Z/o91�d۟Lx��@8�L�uOG�@ӽ:�S���[�d@yg�a�I8�O�-�Hl
�6�.S?�q��s�#�8`�1Zg���\����1�軾����+���������� �T�u��]\�'S���l�ꨞ�wE����+�p� `�Hm���?�r���ι��4��i���ǐ�5 uir�=������7�~:����u���z:�m���I�>���`������J�H+{s�/J5X
,e7C���C|�����y�ݯ��4x���T����켮��I5�ۭ/�I(Wd�Գ��d�һ]������:�\��j�^c_��_D)��SC)-�cD��Ͻ�^�F3�N���W�`>�B�u���[<Q�$n�oU���F�ҷ�̞�FAh#��n�8o_�QW=T�
_\�)����4�Sр��Q�#}pk�$�GS�;��B���V���6����O�ާKw�3MY���I�\ßot D�5�@	R����cb�7�K_	p��r���m���Ly����;�Y�x��h���(���<�C���x����4���咿���s�}��g�7�������B$�Rp�.�	�&��[�� �0��BH��˔6��E�S�&Y�+t�0y�_��"��� �͓�B���x��ǯ���=��@�R�ff^�zn��|ɔ��`'߶���u��� �'t�sO��ֽ�=���D��n�z�͘��:u�-8
���U?V'�%_VK��ʚ��ت��Ǒ�ӌ�d���m~͓��Я���KIqâ�&��k@��l�D�J�K?M�N��Tφ��D�
��*,�M��͵/�E�Z�,��m�H��Z�n3�O|��_Y�7g�"n*���a[ŁIԏ�L`OK�&��G��������r�&��bn�}�ֲ�����'�o�쒰��؁ �R�p�>��D��Г�a�/h�� ���a���}a�H�Qa��.?ku�R}�W���F�1�t]+����z1m���H�A�Z63�"��R|�ç�p殶6+��~F_�p��<��ǵ�]9GتaH��!�N�5��.UD��ڬe���oE��Xl��Y4��K������6���� -O��,&.K�,\x���Q@4Mm����D�9�F;�c��]�s������}>,�=����}��J,��J�i+��a�J�?�7�N|�H�c�?u��Hlz5��EY���i'Np�I1��fԑd#\���{��r�P��N�
��#/��U14�^���g�8W�݊Oq:
Mu������x��x��c���i`��&C&�a�T���.#)Tju���ߐp�%�\�`��!c��������jZ;>�*����r�_�ۂ=��R_������^*q+�Ю8�&���:n¦GIP=�2���#�\؝�L�̀�o���S������wk���-�Kb�j����N�"�`>��9�0Fy��H��Fw�7s?��l�ɣ	yb�Ⱥ^����vc��\:FaʐDtH�c�������A�?��S�T����_�U6{�L�V��p�u���Ds���iq�)�ɑER�4 P��#QpP�6 �*��)��3�d(���i�O[�1�2%r�e���������L��yzY;{�R�:*���~��%ʙ�rp���O��w+�n�������%=��$�T�@���z;�̸?��S��=y	��I�.X�S�Z�0*�}�`Zzf��jr���{K�rg׊������[.��0[[6�	��e��R2�������ݕx��D<�[|_A��E2d;���i��Y�#���k	�t���z9���z��������a�e9KJI��o��:&{��C"hI�?څ��v>�v�ɰ���D&���ށ�����s�9um�DqRW+�AjT�o�L�3�n�s
O�G��vtc��_��Q*���.jP�����gӉ��#ag)������\���_��˭��^����Ā
l���\����%�p�����`����6h�����>p*}R��!jHv#C��p�� 4�܊k\�B��4��C=\� h{���ނ�Βѵ��\��[����)�t[����XN3zh��U��`��3��K�n���^��P�5�W��_/7�T�����$��q`z�m�x�>K9Ȗ��R�x�AH��Q�������aD���<�ș{�^�XY4(k8DBV\o��Y�xQ�͚����N���&����9��I8�y%J$�����S%M%N%�U%P%Q%R%T%V%W%X$�J�J�J�I\������%�KD��.]%e%f%g$�I��	+A!B�(�C	$r���X�D}u�_��^��]�v�T����-�6�(BrC5a�iq3�y�:����ӟH�>�֥ �q��O"v�H��"�I"�J#IS#P���S�׀��+ J�W@�E�*$N��DO���f�Ub) Ur)�U�)�J�i@U�;ph�H
�|��W�V+@V26P%�, K$F��D�	l���K����j*��&���F���xU0�0�W�\a`�0
"3ڂ�<Ei��R������}�c}T�|*�#��{5,qq"���Af�^EP��P���D9o�k:��9&o����bm7�������K}"��>�_��r��few��H�m�&���l���:>�H؊NT��y٪��S'rY�-��^�ChLpIE�;J���\�
�eL�W��ˌ��Ʀ5]��������*���֋�7t6��1��+�6Q�/E<�j,�t��J�2�/6 �ȧ��@��
T����y��.�_3k�쪾V0ܨ��`���H�;��#S���@�<�#�Mz{G�:T�
Cd�)u���v�<��h�n��{�w��NQs�0�=���
���E��L�E����7`~y��~�
;;�o��W�I���=�0�N�!'��}8|O$���.��$��]��O��~D�M(�I4�j$�	��NcC߲ǣ-�ó���5^����s��z잠����J<�$��)g�9_wx� ^�s-1Pj�[w���9&Cg����2�^m����G�ȡCC�إU�=d�t��n	gbwOi������zɊ�)��dJh��L�@���xRv�� ��˻2�(�?��_e��B�O���\�����[�sYfP.�y�yW
�X�V
�#
��0&2@��Q~�2�f���%� �����3���@��%ڠB�$�9�
p"�Wh���lγ5E��A(yІ�]	+Շcj�;s
�^u���+GU���ʚR��$5 ���@f�2�ꢽ�1�ק~�P���ח��ǧD�Ϡ~`����}�]!t�8��#)�'�̭g��iE��ɸ��*,�6M8���caE���͢�4�*��p�$3wM��L�� �K�����|[z8�(������ҬM5��\����!�D������4j<\=�A�t�c���_��>R�rɔt�X�He��󊲙N�@����z�^�eK��Wx"��k`�݄k��1b
TzB׵m�o9$�]��-I.�l4�ET���$�\��~���:e�X�d;'������u+m7�#�����4_"p9*��A�6T粫�*�#�v3��@tr�[;nO�O�w���YU$lK�nn�n��G�+RP�]=qu� &��5�?�6�wtD��t���5��Q��'J���Q��i��xvwJV^b�� _�X��!;ǹ(mT���-�KfA�Գ(�ƥ�,{���ymfZ�E��Dzį�9����o;��"#���~�!�|���G�PϽ�ؐCAʄG	��k�s��������M��e��8�3-�+n�E��yi�gM��`��C�%jK�	l@L´����pr����3-Ԁǅ~⦜V`���k$N$��I����2��a.�e���#!g�T�����̷R	;˯��ᯂ����6FS ���D`:Mz��;Kzof7ӦB#a>LX��#�E-=���o!`s�
X캃v#��13�&b�����0��v���T@�w��Az�x�5l����-c�� 3|�!������9Ҋ���2�S[�3�`O��\ټ��;ٸ��&aZC,)���dϦ}�Ě�G!I�˭��z���8X�$��ғ(�	9T��@�1C:2@�ϸτ
�� t59��Nۻ�lm���ri��Y�mw�rÈq�����9����:H]��2�=hn�
XSDf6d�p����d�{�O��!�?(��ڳ��W�B�K��&\8FX���� �� �d�&�x��w+f���F�,[��U�JUÚ:̂\��T��CP��_�����{٧�cLD/U��O�vU��Sp_�#	���^��_��<�<&�L=+"JxT�7S���"�K|Ư~8ɎY=Pt�~�"�k8c��`��w��L~��nX���:7��Ư�Hw�9�E��Q3��3����k���N�^������+pU��r/��F�+�3�A�>0�Y�T\V�YUq�,����ua]ǫ��Wz����v����Me�TYH�}X�����P|r�>XcUl�@������z%���H �0�:����n�&`�\b���f��ۥ����+"�0�]�;y@��ΔTh9$�>�Kj�����P6��X��}�1H��g���A�y0a��p #U
�X}�W�SA����t�}O@,N��Tg��
B
����H��iV��`Ħ�q\�j<v$��g�A�^k�1r�6�p%���0��Bs���V��͂��>��Ŵ�����X���^?�[�=%H�Sc�rf8���a[�j4��YXo��hps�=/V'�'rdp8�kZ}��d�*w�m~��'�Fq�.sF��:@qf�Q7���6�jyz���?��
eQ\Q*]��|����cX��k���&<Bzo*��g��C��=g�����Rp{�Hߵ�r yH��왍f� %d�͆ǀd��9�3	A���b#i�԰pXڞ���;���s����JJ:�?{�o<�ǿ9<(���S�L�:���C�l�����vV�_���M���d��ϟ�I�X8K ��t|_ӣ0��7ڢ ���JQ&����c\nZ���|..$��$�a�qI{�gR1����R�+ ]l�� �=@3���A�ƹ�3=TՀ��� ��T�Cd�-:,�2���Q�n�.����k}��l�t�8ח��:�"X�J&5���M߸L��(��8��pp�b�|P�&hBU1���u?��Q�P�}� 琗���=�AIK�'��YJ0�Z���Ҧ��f���wXD+�Wri7jz!��[��R9֙N��F�pY��~�j֫�~:D7��p����B�jfa-���i�f��f^?�cI_1��di�0�p"�\4 Ƽ����q��w8� 1�N����5 yH��v� �(<d��xI�"L�TJU�읤�4I�Gb��v�@z��)	P8��yzXa�<��� ]kSpVK[B0)�l�ۛ.�ƺl��6r�9;^B����e$v��Itfa��`u:K�/�c��a�?�c���?~�d<��FW�P��kۺSd̦f|�A�W1�u����L���l]���e������j rVy�8|:PT���z5�x9rg:�p�o��Lv-�w�h��熢�cD|Χ��gh�g���\,��E�+�u�_�/yGr/k2�t��4�L�g������Ph��+a&���7���8�k����8F���0���8�"k�imזһN��T�{�,Ah�vMJ|��zQ E��R\|���P�_�������n4�a�"�����	Y�ױn�^��vb���ߔKB<g�� �4!�ˡ����c0K�=��ծ��ÿ�;�S�7E�o��{�x�T�^�⏎�k���$a/�H^/n�VMzCR
��W�Yf[&Ү�e/���{�=���jŕ�v�J�Dywd����#��V�,���h�Q<��d��>�ER��4��6�vX����N���#_+�N������:Юk��S��b�Y�Z�eI�Y��.}�[۳Č�[o�8H�*�K�T(ͬ�+��P�p�Q50�>tIZ��7=��L�1��&oD/1X��\h�;b�D�<��z�VR��\yQ\Q�R����<�V��`���Q�%��H�B�lDc�?-���
����Su�z'�B�c:�P���Ug���IZ��ü�@�������*���y-Y����L�z.D ��(*�P}�{H���uC�>HrW�u�0x�ل���>h1ɏ�ڛ��f��ut� |�>�`t�?� -��d��p���f@��L��U�:�mD~������mBاX}���ȼx,/� �|�.�Vl��S�-Ԥ���թ�?�zINz�����(8�.QS��E�]�J�0Ӷ �K��n\�5���[o�_#��R&ƇRM��C�Ms_�����e3Dx\��z�5]�����ئ��8M$i顫&��Ұcj^6�����+Lj�G@���{,���r�c�9���N�׻� yHr|
��<� >D��Ӱ2H���rPs�d�q�8I��L��@qg^��[Mj���f5Ґ7&о�a�+%��~���:\K��y� �22�����%A$u����+��l7�p�A�lѥ)�B{����W���C_#�q�(٨�N���B����7���Ԧ��\q�5��s�~��!\��P���ͳ{B��#�=��^�FcW�~(e��>�q���H󡆇�(�?���i��>��}���iy�A��S	�ƧG��)H)c3
�ÿx�e��{h �)�`5se$��8-�Á�����C{<w�?��X��wg�U��\(�$�� ��8I��$N3Ƥ��љG8��^23���>�Z�w���z�l�T��KҨ�*�:	ы7��˭���E�ʠj�g�4 ��v�Զ���ku�҃O�2� ����Wl:B�BX3ꃘ��>i� ���c� ��T��u�bhjyR�O&�iM�_Q[fQ�j�\5pC>4A�T:��)F���8&���Ȕ� ||�e�,R<��u�?�_91 ۖsuF�
��5.l�e'�KӰp��Jɀ��6N ܔΖ
8�`'��Ӹ_��NiA'�XP�����-ly~��߬��PT;o�X�]�x\��YPAʾ����Z�V��R��.<�?�&ڇ���ݍ������@	h.9x!01[F-�X�[,��f�#_uy& -��
SS�_��ItzC*s�,���鮊L�H\���>�L��.�TՁҞ,.��X�`>06H�ţ�X�`�*�l����e���`�����l����&P�Tq���K�Щ�*r�nr 75�y��À�`g��@ꀴ|���5�u�А�q� 㭃�H���	�_@�gM!��tC1���;�	>N�s]��?���lIbjy�_��Sj�S��c[
�PAe�6+�f[�*۩�ÍZ��y?�J�Z������Y��~Pʻ!��t��m����Jn�m�5kZAE�7�����sQkC�`���+1��s��N5k��{�q	�dꟳ5��Jh�/����'TtֹD�6�go��z�b���7`���L|�d�5A5ʳ��3^�V����ϔ�)�_ X�_ֳ\w�$�S�p��Ze��*J�v�A[��yP�j��m�x�����I�A*4�*��g�	�P�F�~�X��G5j�?&͵��B�/y�+lF��:��;4$Ė�UQ&�
�����{��~�3��x���9x�}L�uB�Ѹ$��g\���W�����6��#��ڍ_j��J�>Y�;��O ħ?�J#	�;�����oң��W�a#o	Nt�r��:�|iuD����ԃ33#Pd��X�J��W
����r|�{4F���+=6m1�/QRn��"mo���{���.H����g�bmO��U�S;_���!��/	o*'ҥ��2�5��=�f���/UZ�;�ն㮐�R=[����0Sfnv�Qw?�{�A={ȉ�7�/!�6yO �O�}�|S�,AHQ�`'a�R\��e��\}Q�񼌣vVwv��^��o:Z�G��� J7��}/((�1��z�O��qu�N1-�⼆���Z���V��آ��d��t!�Ϡ�L��G�c�>M���4�T�/Tkb����6�3Xb�����2��,���X�΍a�7Oy���z��@ny�=7�rs|=�m�:Q��̯�̛� l>��^Ǚ\�Ru�UN��Ĭ��r��jgD�[�o{ȟ�=
�SGL�x�G��R'�0���zZ������Ju�Zڜ�D�*RB@�����) v�}��ck���n����E����dM�nA�lK�����l���������粦7x� �;{�����SN|��d3�S8�:�ގR��4��pk���&Ax��Ca�dr�������ש�F�m+��M�(p�>k�Wz�B���6V�gw�*]�����O{^�	d�k��u�z���E-Ϣg�����;�l=�9"sM������3��8Ap�U6wbl�J�_F��w����t��哆��^@�z������vn+�疟���s��B2Op�[�6���QX�|�MG%��h 
i�5z�-ͅ�^<�Q��E��On�8���4e�>S7�F�Rc6	d&�ħ]�zr݆y���W�k7��o�^�Һ�n!�����
�EI?ѯ�xj���JG�W^]g�Zߜ��a� �L�f�j�vE"ͽ��h�{�d/�������.����=�����1p�׾"
���1��/g��ꮈ���F����,bi�e�Z����q(��-ls�q`|�ʸ��M}5���Ӹ�V�7"2��zo���Uy>ANg���%:�_�v�Q4��PGm���Aj�L��ϑ�+qd'�!C�GU`�b��mȳk���b�;LO{�Mĝ�+���l���۝#�3�,]�-� b�Lݍ�H��{>�q����&�c��޶M��p�a�3�����]���I��s��=��])T��^�P6qϴ�^i�qk�q�N�� ֫^7���q���0(��my\�1�ѩ ��l���5�!�I1~D�69������`P4>b�)�}S*�(�n�db+E�D~�s�X�y�|-�$5Ut�,r��Oug�?KMv��Q�ә�b�;�x*\w]���|��ӧ��Ja��+��M�����&����H�@����r&�����}��H�F��_��J�܂�$�8;�Ka�1�x��5BJO�9��B�;*���:K,�q9��:�RH�\+��V���g,`�3u��_�����6������J�w�䮝p�e��K~U�
/��_����YN� d�?�7۰yY��9j�c?��U	>^7��#������˾!t�}��גp���!�X��y;�K���^���c n�`�(1}�� �:��f.�b�.�pZ5���i�xxD3�����g�:��;umٶ�õ
׶ۀ�D�>$��4^q����I��~���;����ˎ�X���꠳���G�i��O�R'zT��F���>��ﾓ��K�ڷ��j� 1�O1C�������nm��0`Fo�o���1 ;���]T�Y:�'M��n�Dڜ�M�&e�mgw7�ns��pZ�10�3\�o>�����_��-�{�j羀����M���v�w/p� �S#��Ykف��� �6�&��B��P!�B����������`ʘ`s��< Ԙ��Z),�3���n_]p����ۇ�y�Y�oU��ē����
������feC��)��	N�z.��~D(���$�貱!����q�����a�;�8�1(���7S���F�+��w��ޞ$�킴��tA���>�Iz��T�s��u'6Nu�8�!\���@�k�M�#E��(t�~�������k�v�O�J�K?	��Z��nٛN��<��.��ə����
E7���(�QD���~<�GC�5̘ �hQ'�!����)�UѾ���:!�0��GĪ�.�#MiK����FJ~�2������L�s�l�!A�Og�����2�*Ba
�*P1��<]�d1�P�`6����Ɏ5hg7�1AQ�xPR�mU�MM����=�j�jF��u�_aK�N�R��A�0 ��z������V'�.����mVHz������'K���N�]	�E��<8賅)�%e҉����8=u�Z�����N�1qqG���
X&���b:���QvS��âc�.9C����[�y�G��u���K�h��`M����=�bQK���!�ࢗZ~{��p�Φ�o� l�r�@�^���Ÿ����6 ��1��搔r�UQ*L��U��J��v?|vvN�����OU�)�����p��fQ^�օk�hDZ��k��dƔ�`��Tͽ�S�[���:�~'��*g�o���1�nM�=��r��0�DM]Z�R�N�`�;����sd�f���n�ǖ����n��6F	������3��w
�΍���IJ5�]�����v��1o���)3[�y>\B�γ�D-v�Y�߼O�<ƛ��h�P���׽y�=��R��q8E��c�*��>�MzQt/L�)�Gq3��_I~�1�d�݂0I9;͓�R]������f�#��&��7����#1�H��<|��s]
�d���e̪�e�B+�	��vf����~����u�5���v�&����	�7�����h˾���>yzm���<	�Lѿ�h��������`�J.�ܟ�k�=Zfc�O�Y23�b��
���o�����X�9@w�xYԪ' N(��#[�#�����B�9
0i�0�˻��ǭ���NmQ:z���O���� &%dL�g�.I���,f�f��Xo��=�L�T֪��g��	�Bܡ�o�l�t�dSD�:Q��s8����F�T]���'LhUin"1��a���� �u�2��XXr��U�=*�W�O�3�ԧ���E)\��_rω���nJ����z���C�
�H�0�擱l��B��snڹ&�|� ��2%�jZ�oh�^�p�]�;ї�r�x��")�#�h*��;�p�g��h[\��f)��4�/ {֓	S�~P����<�<�1ҾfM>���5�P�:��KWd���;���og��;-��dǭ�w�:y�	t&��W��$��مoLN��f��eZ�L����gDQ�o8P"�@z��3��|�5w$����%Q�|�S���BI-�@��%jz�o�o_&���XE�gmo���oY��#`��YP
��^��w�6%�c�����k5����~D(D)E�J�P]����|�'vU[�������w�L�����K ���E?��~��C��O�?�.�~�O�+���I�ɳ�ks��Yg�g��{�5(ylU��ȷ�J%�P���`�U��6����Y�,�g0w��ou���L��lC�6��Yٶ;j��R���;f�}4���B�Ƨ�,�S�-3�#�1�K���~^�1���UF�enY���+3�;���2���H<΁��&�ѻ&�6��_ADA��Y�.�K��B��V��t�<��+)����w2f�	Y�U���W�ކ��8�}�~���d�Ǆ(i�����\D��ؼ��6��Wa����{-�G�ۣ���~�V��>0� .(N�1T�S�f�,��{�=�2�vK�.��}`	�E҄K��</���p�n�uK���KS��=����i��;b6W�OG�FnJ@�&k���-<jKp�����z�-�j��РL�����oR|������1ܸ��s�$�-���Z�,�K~ƍ{X���P���v����n�A��'C��V�#G�W1����`��t�#>����[� ��N��g�>��C8��tV�/8����l hM��!�=Y>�ſ=a��H'�	�JrW�eI�ă6�?�%�B���U�Vzܡ2�u������#=��E��6z��x�P-x��������,,��O�����3�,x8J�ҝ��Uh�rQ��Giߊ�.����ﲑ���}.l7.����[Ԑ'��tܸ���j���r=Ž�z��m�I*�X@f�I�ȏ�,���?do��WX5�Y�|���?ݨ�j��1�b���@3�{'^Oo:L��(�'�s�cg&�@fdV�����JW=��EM�X������\�$��c�2���İBf��K��e�,R���t~�i����:��F^�̺�5�)J?�T�O��;vm�ѣ�i�h�����Վ�$������ET=��U6����i�����4�=��5Væx)/;���֢�P\2m>�O��ݎ]���e�cEel�zl>�`�NRy>�XG��Dx<tm۲Y�$�?b�䇟=��M�
�R~��N��E(�0܀=���?��8kK��U%u��u�l���K�h�ӓv\|��wZ���7=$�ͻ���
�#͎�E�Ũ8��Ҝ������[}��D��t�C�+z/�HUΦ6�d�/��*}c�s��	n:��7V�4C��ov�� ����z6L��c��<�?��Ƌ��;�B��_N�"���z��.
��?��Bug�Y%*�fM��n��]Y���_Nyp�=�s;��퍹 D-G�3��*=��a0I��#�g�Q.3��Ó�X���fr$Ʉ������/�`�yV����IH��oM�Vo������<S���ȁ��QU�Z�~���̶��������z��F@�W�	���ڝ�G�&�2�^�f�RA�^2�|�p|A���f��-�������ʴ�L!w��5��l�4�B>�iw������me_b_��52'����^+�aYS�#?v����,�?��u��w�|b��ǁ�3�1e�nq�\�xe��1OR�Z�E��t�
[Y*�W��}�~Te�� �����S���E{���5����VԄ�&2�_tv��:y����u����� ��v�R:�~4��`�Nt�C�A:��&O+��Z]"�������s[E������ز�o�z9�������M/�K�����sޤ��k����~7T����/M�<<s��̠�9���Ikd��De�k��d)���$��;İ��&q���Z�,Ew�W��& ���c���2z�Q��;�A� C�ӑ��ԵP�����&4/��e5Ɗ��6�0���n7#�wBx^Q�E�㩕��]<�ɯ�i|��I��e;��i��mt�����;P҇�z֨g�5½� �Vd#K���\���H�1���7<�R$���7L�.��O�����6KHZ��>5�f)�O~���#�������^�S�%� w�6d C7�ox��Ca;Џ��u���}�c��E��/&0Y#�w�^�E�5�>r&�0p�&��g��#��h5��N'/�*�dH��0�,?��Y������D�;���S�d?�O��S�H R#���@2,/�,�6#���:u)	��<�ҳ2*a���>�T���������hr��]N�e������C���ErZ�wѲ]|��uZ{d��v?����ۑ[�5u�q�ᶇe��B��3����������}�UG�w3��n�isU\��[l�G���=�j����n�SE*��c�-m>j��%�[�&MA�%j��_QBxvѯ��.N^�ǭ�ۂ�Q���� $:��\oE��Y|�ޏ�1|�[�n�*ۋ��6�bW��Y�������N܊޵Y�U�����G�N���7�#�m���i^2A�o�p���W�]D��N:�� W�;��p�_�����/����YC��fmR7��l���������1�?���g�[^ƭ晒���@��X�2���ߔ=���:T���~b�D�P�SP��@�Be�Hi>:��fU#gꌧ��YH^(X�!��c�ڱ��$�a<lK�D�斑��9�ˁ1ރ�����ƚy�X�����c�^߲S�M��Eޫ_�n��=���46�@k�_[�1�?Bo:	�]���j�����&l���B�F$�C{#��i10�|��Zw�!P}O	/�~��ʺ:IOj{��1�C���;F�Oޠ���tj��k`���=:Tʩ@�q��p�]%���v[��
��j���<�e����۽��Z�ꂆ��ܼ	������\ q*�K��+�c�_�C'_��1���i�T��L�!��8�D�7x�wP�`|��^N!R�?D����,�;�Ch��M����ݜ/�=�q�k��O�y�A��2�<j��z.��D���{��#����Q����4�=��HpS*�?��E����B6�eU�Ƀ��������͢���9#���e�iج{����b��P���h�$�� �>��Z:�i��������m��qx}H}݈�.�������;�X^vׂ��$iS��5���~ �e�0���� a�r
�"�k����7�#�A1`���K2�G��e��f2|�i��멳T�cF���T�v��o�&"�IՅga"��ڛ%?�Q"�9�ET�j��%l�JU���pyB5l":r�w�3�S �&ouׄY= 3����9�Z?I�������V��%�p:~�{�KR01���R�8�=�:�4�;%�9��µjB�zbLɰs������5� ��:p9��,�g@�m�U^L�X$�?�;�V.t�/m�1f�|�8xm:�s��{P�FVgD�G��O߂F��f�\#-��:,O��\I擘ޝ��{T�)�#�-�>`_��D�辌��I�e�{��b��"������<�u#�Q"Y��u�As�GB՘�R��?�ؒ0��k��[x��QV"�53�qcM�t%��q�e��|�f�n_�]�{���i���q�emM�%ԊU�жQy������nRJ������f8�ET�J�
;˄�t*gI�����-G)ե��4�dS
� ��q���`� ��X�y=�' Ç-p2C���5x��6B��&�|+�m���ez�Rm��"���射��p���o�x���S�Uޢ��W�&a�S�5��b5�Y��Ch�D�G��!~.�����`��o}C+փ�5Ԁ�FJ����1;k��+X���xE]���4����eS���G�8��7wS��8|Df�˶�K ���d�����w�,X^����Uހ`	6lO�:m�Y��7D1�|�q�wi�ä":U�ʰ֒�+.QL�A���dL1�<�A,]@������:�2sE+
����{|_H1]�y�#T���+�#�+���~�u�B���G�Q����ޟd$c(e��t��g��W<E�o/�*Y��?�3�Y-�z��AQa���3-��mIz�-���V���uP��7'ض��q;��H��QR�T�5�6ᯕ�]��� )�BY)|�?	�*�+յ3.Q0�W�~�>�9U��?ֺ�E��g���T����l:�|א�Q�J�İ60#�C��A�uk��C�A���m�6$; *
M5p��	�&��8� ��O�YAD��t�O�Xç�����F�Z"�(��{��%��*�?��ST�\+�
GЛh�F<��L)K��ɶ �hQF]^��`�)Dv��j����i�ةT�}�×cQ5퉲�����G��v/�Nʫ�xm���^���j�?&�c�ה�k9��BuӪhY+3�H츸��db��t 9�"��pP�걎��:#��=ƿ�i��/|4Ær��zs��ٽz�sV��h���R_��#M�Y�I(5~t�5m;��5�����F�r!
e!���me��D>�z.�ŏ�ݶ��eu�_-��<=��^4�����`�L/fh\�1X;��H�yjE)vr�sWYd�y�����k��s���>�s@�������7����3�W�EÓ0a��Ϣ�~wO�/��,�3��Fġ2���oLa����6�L鳵k1eHvP�d�b��`��<��>�2{qe���(����.e�G��G�F�q��򤕄�4�	���s�V����5�T���/��mt��n�k�x)9���N}��8!_��z�_��~]V�b̠��<�����Y#l�o9��-�������"��s���R������ɼ��r���c�2ȸ�{g�v|�1)|Ԭ����7�����ܓ.����or���f����I��Y��W=�� ������E)A�3R̹�rtH{-��T4�J��:1 Q�.6��_n��-Q��bQ�S��'n�eʻ�J�FO���B�<�n�A��#�;�U�M�U)@��v�*R�)J�:��zg�y��A�x^@{N�Y�Y��]��kһC��Q��K���M� !!��y��1�#���G�-��]h��~��x;�ו�0�4�$^�h� 8cwݿ]���P��S�ޢ������[r�l�x�Æ�F�O�}v����C��ɼ�s�?��f����ϖ�! �QHIC>+�IO�jo~W��k���|'(P8��k���s��HQ3:���L���>�,z�)�xoCD;
͛�|�M�k¢����6�̩��}��`�KN�Ɣ���=�z9�� �ˮ/FCaG�	��.Pj��*��.;W���,5�͊�Ռ Ę�p}2ǒ=�#��î�0а�K��m�xR[6�w��=������K�T�R3���m3)nYE��ViA79�6�PM���>I����#Y�[�0{q.�a)���P	
g�2RoJ'+�[�B>؃�鄡�H��M͍f�~8�ٝ
��F{�+��C?l�Ʋ{M
B�0j�w�?����eg�>b��҇��� ������=���ʶ;zR��;<��"@t��C��x��}����[4$���i�
!�~{1���ĕ_t�5n�a�t�>���أA�3�Þ2�:@`n<b��46@�/��H��;�(��*D�.<������0;�FٽM��y�)�_�x��N:���c,�n�Ep��_t!� s���.������?�Q�μ7j���P��}Z�{��\��Z�����i�*�	4�1<�6�S&��~Sak��;�q*n�1�pts�bƿ��5�A����#!(�H�d}; ��$�#0�� �
�M{S��/"�e�	���t	:��[y�L���}�}�fᝄ��_%+��ƀ�k��,���;2�G�!���(V�o�����k�gd�,:��dx+��o������o�(m�d����nA�G|�t�����zXd�R;�0���������e�h8iZ�0�=���M��C��6��u��#���z|s��e`�kӐ��"�Rd�����-j��s��0�f�0[m���@D��c1dgZ�ܭ�F#�S{M� �YȠ�k��?t�Ύ�����qâXD�5��,�NN�7fW��Z�CW�o`��n9S�;��=f���B���,�J�J��w�m �Pq�M�;�'@������q�~��3�at���I�T�yD���6a�������f:5�r�o��Y��۝o�}�o�\tg�9�t���1�5��v�<��:�^{G��jDf�ݨL/��S�'�:�n�� p��-R�
��t D:N�}��Ӭ8[���h���4r�8�ְ�����"��ʚq��'8��\� pCu޹��+8�#zL2W��=�a��2��CfR$`�D�?2�)'pA���h9J#f̥�МQ}M�Y8�������!W0����&o,����#N�.�H�J�ey�
���o�rP���g?����Y��T��E�/�fXwu�$�������J�&��i��D�3�b�!v%��7\rq=Q�ً~�������D�̚ޒ�'����JN���o��C�mM	���k���ђ�L�\��;tR���xpH��P��B ����)�A/[��v@�������W3_-NI��6l��<͸��n���&��i�R��H{��!��Z|�I86Jסm�Ǚ�8�%V��?�&�p����Z�wm�6��	����̳6��l���Y�:���t��F G��CmF]�.������*X�_���_�煆�(�c��������MVR�=�����!���"�������OYc+�$?��˖v��Obc�I�G���$IVK;9�Mڗ2d.~�� V���h����I�@�z���ev�^�<�m�;I�n.�(H�T&�љ%�u�)����U<�6�<��u�I�#�浫��wW��e^�Õag�������Z�|ۗV̝��%3w�f��g/�EW�@�!ɡ�QX�ӡ����mr����G2��	U�![��!��m�!#�R�w�8����ׅ1�_�NUmr�Y��3.����Z���6�c�-]��d=\2�썪cg�r�D���"�-�m� �gm���$�`��*�fķ+(�9V�r�`Y��\�����H��Q��� [YD�?��0?񾝡6��((�v�X��x���~8s*)v��$�3u����Sk�)�,�p�o�H��|���9��!���9Q�N��$�英����Z���m~}su�:x�3b��.��#���5�@:u����/���f]�X1UYV���u._��u7���뫚 ���)`E��s -��O���(c�ĵ�7���VsK��Z{�r��7�Z�K�#샧���ϓ��!N�5Z$����(����0')�j��YHl7�q�l��5��m|]t̄�|���u"��c)讋�ׅ��D�"�r���>�ex����]	uo@��ri�&�td��!d�<C�z�3����-䴶������k���$��h�l섗���І�ޟEX�*\c�j%��!g�t�`�e}��NmuC�V9Oy9�y���е��F��m�"�����7��Q����5�"�Ĵl�n�m�t���Z}��F�JS���rSn��p����&7�aVt�X٨��٨�ݏ=��9����[M9��c]]q�]����zW}T0p�������'_�#�������l��(1V�GK�������"<��1"����B�$;RH|�q{���Vm����VQa}W�����C7ZT�2���2j UmŰo����v��eCSs�����5:K�N7�|���B^����5���m���f4~���$,`vj�!��ton�w>����S~��EJ��Z�,�^1��6ڡ����O.;<�J���8���:���Z�C��+֮���a���Ljk\���![�鼝/��!VHZq�A�*�q�[3�^�j'lr��
U
�4y����}����`��=)�>ٜpM��*	�$�Ӭρ�5�J9��V,$�`��[��7�k	L%2��-T�s��$��?���z˩hH^�������+��*gC#���&�䩘T�N�ͮI��%w�nU�@����1yZ~����p��x���w�}h(������ڵ�?��X�o�l�ĕ^���[Z�?��b��o�^�g�2�?�Y���8+�����+vw��i�!S�e=	
$o,Ū��}
��It��Hv�Hvk0]T�ik�[~��Tq�ǹUX��Z��m�,�-c�6�Rh\��b��) ���O�mT�⸆�!uƻ�q����t���)����������L�����4;�ஐ[+�ɇ.�?�a���S�U���[�lNW�D��+�U��9�:�_�}�ڴ$_��V��oI���Q'�r�\�/�n	Q�ֱ��d�#��0�8�ޯhk$�ۃY�?������5+�E�9E�U�}��<�Ey��3�q���h���� _�� |�[d*X�6(8F�r�(N�]c��}Y�j�qE�Y*�i�rƙYmy悴��7Rh��F�u� ��R�`�Y9P-��GT6h�	��}s�J*E'�+7�������ү�C��$���b�qd����$���bb@8W�|���~�\:�(�z�M+��NdX��}���o����>3̟o4/�~[a�Xo�ݒH3o1Bw�*�4Q�i� 	�j)xm=�v���m�`��qw�JN]�5����J*1�K�*��U�=��Ǖq�^G���ӂ��{�CL�0����Ț3��5�Zq����V/⧠���ā|L��@��{Ԋ�/����@�E�|`�%�RD/��4PY������0/:��]~�--��������x#�=R:XT�7�y�Ѽ�D��9�`1�����8"��� (Kv�a%���L`���0��X$j�)�)�\bQ�^���9t��]��V����>�u�&�M�7�E�����2��~b�p�i�m��:D�|P��ب�6���w$�OV��ec�<��)9�on��4����|5�b��-�%��+t���q<%�Iږ�o�A4�fQ��J�|S�%�7 ��q��H�n�ph���㠾<�p^v��]�����>�P:�`��>a�n���S�@9G���w�h�=%�.Y��i����>��O���!k��|�@"!#8	8#rX+�!d�f�̊AX��������PeVVVJ�_f�eC�:�J�;H- �m�Lt�Q��M� ~�'H㩖���#�:���P ��M��`���`��vدĶ,.��/-�?�ij�;,P���m����d�"+��8e�=\a�����3��QW��!8�Q���7��GJi��wBq&����L���m��Q����AH�h��]e\'�_��v��bTP�~�3��_rm��2X5n�l$W��>���
���J��Q��=()��:�!�e=[O���:�4W,$��k$��'��!_��U
v��K�e{B��Y7���>*R�o��ih��$ey�(�?�K���Wd|����٤���=-d#��@���j��+�_]��	�@oS�lZ���$<�`�5�r�_z�RI�=������Ei~lɭ��{�-w!�5��aa�>z2�ഈ���OZ�l$]��0<�q���b����Gn�΁ltǀ-I7nbq���_?���)샾�,�p�u�^g8�(H?o�$��b{'	�ai��|/�Y�P:i`���w�]��q{ra�߭�D�>�9l������%������O�ǳQp�8��Ĳ��*}��V�����2TB��q�`M���;o�H@߸B���|���͍;�a�]����q�,��y�"L���I8:������OW���Ȅ��h;o����?t��R�K�^���Z�ؾ4������9���:�n��L^]-FE��lf�%��73-xx�D�o>���+ۇh�r�7�3_Ae�(~9�=��^�"ת�9E������>T�omAblw�H�͠��u]I��0�w����l��0EF��=݀rpե:ʟ��l�e�I��i��	�C����E����+�u9�@��䯐bؕ�B}�#dࡾ���;`�$�7C�o Ū`Ӕ ��j��
�ag~���P�c�%*ad�+x5�
�ڋ�ӔS:o4��u��IF�6��|�G���5.ŝ(�tԽ�wâm���PD�5I��yf��N��Y,F~Ī�X���O1r9��D��[�z���˅-���[ �4�Z�|�$ϟ$[�Q�������a	��4ϙl5��Pʣ8�d:���$q�)�>� ���qk
l+�u���B%�s��b�o�dk�k���#y+��#T�U~4E��u�>aO�Hr�ˮ<�G�!���*��ŉ�̲9 ��ї��.�΀�{-5�XI .�G{��_�_A<9Q�K���х��cұ�Y�����n
h$�#�6�J�Ž��x�K���
����
w�V� �aC�<9-�j�3 hi*�1���"�nI,����"^O0�!Of���^`�^��ΚP��=�8�Ե�Sa�v��Ȋ%]3��y�^�2m���vmrռ7A\?��=��_?�}��Ta&�6��P%N�Ž�8&���(��J�>L5<���.E���+�EgD6��c3�]����}m�r�Az��{�o{jS�V0O�Mb�n������O�΅����"Z��E�Yn��2ycn��D.��  ���,�߶Ǎ���x��)���f�Jc<~d�t||�`K?�yMC��O�%�O�TV��;�Ű�W�aF��xĵ��ܷ��D�HO�Ȍ����e�@x��R-P��b4����ߓ�&��#����NZ��Bo���X.ԩ��F�}��e��#�N�hn`v#�1����+G������������㐎q}Ō��¡��`e��W��B��tIA���%?��*�ѧ��3��o>XǶb�IS�C�
n�f�#�I�y-@�Rb���f���� b��/������|�a���$��k�X߸�V)� {P�[�E�1n񏯔o��� T����#���^.�tsc%��l�j��O�Y6�3N���P��0�'��?��#ˆ�`@��h/���R�������{�>�&��{ވ~��5�zn"lI�.��䳜��$��-ހ���1�5F��{5�|W�Tq�{y"�(��t��Oױd.�s�c?���L��w_��կ�H�H��F��8�m�}�C��.�����짃��UjX�Ī���E��^�Б�I>�W锟����}�	�պV0����;|�r��T��[}#ƛ���`��^�5g�`}$y�T�� q�<~ͤ�3�,�3�Dr3�
YkJSB�ӫ������.[�o)���}hz2�W����*>���@W��3N(���m���N��Y3\��$�!C��Ds4��" �S���]<��� Q3���.�Ow���� �'���KT��KP����'3Iw��T���he�Ka,[}���s��ʉKC�N$���(��L�O7I)�hD�/5�����b�&e؞%  �P��fKI��WW�vp�ɵ�>k���ݢ�|X�n�9ͱTm�}m�85��+�3�7����[Uy�'�>�I1���;o�������^� W�FaUe����c1�� 6�sfl0�v�G��!�����l�8�NG�U>¼��n���BA���_o���s��n������۸�v�%�N�m�]#Y�t�v}�VQ�&J�Y ʏa�';�Ӈy�`��gL}����y{��) s���C��y�>O��\��z��}�b'�n��mtG�~6�s�~���rp/���}N�,��-���Vs�fzk8����'��V���+Z�@�]/r���&��}����!*���w�b�p�WP~K͍�ii~dɦ�`���r�o���X%��Y�:]~�yd��nk���t�+���^k�Z����!+Kܴ@��K�]��m����mC)6�9>�1-�+�`yٛ��9��̶y0��w��3����o�I��R8������NQLZ�N�"�7�L�.��u��'kv[����*�$�f�|�6�j�G�$L��3�F�`���}
E�IN�=d1m�M��m-�'����"��'�H�dum�	���W��w&����ဉA���J���CuGS@d����"! ,��5�HE�)�W�%��ĳz���uR��+�V��/��L�j�p��6���f�ΏVLBbp��½'��Yd[��k 5e `Z����1S�Jރ���7�o����.E��*�C�
�j@��� �%2CẗY���}2=�u����}�s.sƭ�\	��=|;�j�|^�1�X�j<ũU�P��D���t�d�����U*_c2���P��x`
����=�|XԼ4S��E�Ѭ�t��t�(�KG��S��kA�`}���<$o�$|1�D>��!?����lB�6Th�F�T��*�e��/��&�{���·ݖ�O	E�C&p�ټL�\�'܅�X�X�1�i
V�03�����%"ߤ<"�jX?g��:9�Z�'J�.�(lL2�D�ʤq�L�iJ�|��3��{�����ڈ0�A�hLW�+��u���/� ��(�{�踕@0��P���	���o'�˥��W�%��Oy	C�`��a�s��N33F���d^I� zEF�`�U붹�y`�VоC��_�	��9A�%���� �M,)&dI��^Ǳ�>�"0�)[�@X$��x�a,�dL&�{���Fn˵;����Y�4>ţ��E�ׂ�g�D������ZP2��6�=I Cߢf]������7�� � � 5��L�)[ɽ
�.��<�lp�0�>{d_Tb�z�l��,϶# =oW�O���k���7����E�e�((i���U���[���/��*t����Ek@��?�0�����b"�@쩐}��ˀJ�b�Ng�H�_����)\����&�Yl�b�(�.K���,��榐��>Eb�Z�G}A'NJ�D�d�#����"�Y#^�|�Z
%Ul#W�0��p��E�����/I����ϴ�)l���.g�:A�����,��C��x5��>a��G���SWF�	|����Д�)Ibm�Bn�X&	�̫�&��;(*�63��ݕj`�ԋ��52k.�`��ҟ�*�7�"������_:sҎVkͤ|��8.�h����v�R���|��pp����_��{�>䎥�&K|�-��.�3��Hk�_�̅^���P�>5c����[I_��E�{p7p({480� ޢ(RX�!Āɼҗ���].��$	�|Y��� 36`��?o^z��wT��o�\N=�C����imf*]E�ܜC�ɘy�=�f�V�����#��<SM�H�gLD�ë�P�'ޠl��B@��Q=�$���p�Ձ��3���!8|7�Ø�Y�L��5��_K�JG���-\�&f��F�7Z9kMGp�\q��H����!���-�!.pFͦ_t�������)J������D5�*0t,{��H4n��J�N�jN��Ha�/�5�t�ߘ��ͽx��U^�_s�=���/8��/��^AꜫD
�4�W�*6(qZ�M��D�j
�v��Q�ߦ������9�E7}kJ�ܚ�H�Jхt������-i g��h��5�dֹ\�~G��җ�1�P�X߃�!�|��V�EuS,Nצ(Phn��ٻ�VpO1��ށ#�`�Ly�ǽ(?�[h���7V#�$�yEc�%��tz����]�e��绁�#w��{�Yb6���5\iHTuϷ�ph@�y���j���b9�K��׺maZ+ov�� ��&ZJ��U�#`DY��=����iLt4
aTa�q[�ҙ�zDZ D�p�g׋q>�Io�KNr�f��,�.�A�c(�m���p/������S���2��c ��w�%�/����E�n�=�eM�D���7�$O�o޳o����^R+=�!XC�F0���I-���B�VW�)��{�2t��X�:�|�m�y�N!�p�T�%���޽k'���F��b�J�s܊�����qw�lA��<W��	�خ'�;;_G|g�^�	�i�]�^�����������ll�)�P%���r3}�b��O�D==A?nsd��"+%*<�$�g?
n�hY(��� �{�iAtn��Ly�8���q�Mn���� ?��@w:aΊ����Ɇ,�����F3�ee�� �р��6*��c+y7�Ap�M������Oir��J%���4f�Է�R�eE�5+O�?��&9"Ӱ�oʐ�zk:'=�x�P�y��n��o/�A|s׏/��VOy�t�$���c�$�k�Y��񁴑��Qe���0r{h�%� ��4	JR�jF��	5)6�"����S�޺����D��?�7+�p�qW�x���'��Y� 
7�&F���p�W�g�{���~�{��N������Y��w{ƚ����k�������쪐�����\V�j'�	V^��R*���B����zՈ�p2!�Rg��Pd3<c�Q�ؖ��Xz�Z
���8�*����C;�0�"sh[1���HGw鿚u�Y_u�Mj��oȉ�(� �Su�����&����ʪ�o��P{K�pV�~�-�);��>ϙ�ҺT��ՂAf:(.�Dά-/A'�{z�Xl_�G�9 ���ա6E	�)(ty���~��I������=�P����Vm|QY9ooqG0���GZ'q�/�\�JF������trr��%i���V#��g�j�/ +%�jX�eK·]��Z������Џ~�V�U
��Ģ����=��U
{$/�9QuH�������[=q�t� @A��	P$��� �>9����\q��͇��ά�죓��VJ��-����B�nS*�@��ӌ|���<$�+)O x�;f��/g���ڤڮ}3��a�p[��GNu�`(x�D����n�z���J�n\=ڽ��ʫ�3o�3"$�G����$G��ltT�z3����fڢ�r�� ��y��'ߌ4���Q!rgGD�-�j�ū�y��"�ǜ4�h2�l�icم��bjB���k��~�`܀��a��y�[q2{m���+��QWE�"J�N��g�H	� ����>�D�ޑP���=�7.{��Z!z�ܰ����4��UD���<�`���ݐG��Vջ/^�Zs�d�is'O��ML��j���:�|U\��Q.)�e�0K)�(H��1��oK����Z(�HDօ�����փv�Fso˵K���Hk���]!�A�v�l��
Eʠ����Ĥ&��ѡ$a_0r;�P$<��Ϧ\^sqAU�.C*�UU� ����)e,Q[�$��<�4�!IW�����Q ǆh��9��5��A��f�h)��I�~@N�y�
�y��ׁڴ���X�E�����ɞ�����PK˺�P^���Pݗe $�-t;C��j�1���л���0�ن�̣m99O��u�`'Q�����Σ-�림Qљi����1'A���S���j�	yt����z���ﵢ��}I?�|�ý�C@[��ըP��*4��_�]�8V���q��A�aYyVb�����z�/�F���^��oj�}��Pϑ3��MLt�IUhVik��j��,v��z��nk�ZKP�l�Fz��1�RQIO4DI0�$xM����RX�-
�7����k�+$r�X�D�n_@WAV,L��?�$_��p{l���"��h����&_��!͠b(�d��rN����1N&���	X�G�N/���g܄��UZs�^�fz�~4�jp�ۇ5<:���3~Vn2!PT���zr������ �G�;j\�Cj�T����f(:��o++Q_�݄&dS��$:�M��wQ��?����= �~�U|��^G=O��Z*c��z�[V�/k&]�L�������	~��@��Mi�zH�,�:��}j�0�����=��E�)^�<	�Jsm�����f��ވ�ݔ�J�9h�m�oBܨռu^���QC����ҏӠ'<^V4T�����k�n���ݪ������O%+��Z� �q	\�U r��'yT\bSQ��I��	%�% Ӣ}�����?F��=�\��ӷ�rͬ��D݃��J=�n�}U*��jT���<�@�w�������N8,):�sY�1�(���;�p(�Ҳ�����s�����n"UT��)y�u���".�����h�������`�z�[}��9��g�s9��m�Xۈd�Ў℣I����':.0��/��4�Yƪ�[~k���Jr��d_��V�o����1�q��q�O+��$6G���$c���+�'�E��4�İ��$�{OG��A�>��f�}��ak�!!���abUO�a18(h�%#���)�oȣ�����>�6<�
�Bϋ��,BQE�$�!p;�♺c�]
 X��Q&B*���@���?��'��>�uRG�f_&�Y/�>[�S��j߻�THl�(?��qq`F��Dn���K;�⁤�)h�Bk�aO��*�`���H$�����c�}�4Btsr�z�T�$��=�w��~�ҘY��L�K(�����M�D��2� B��B�"�4������܃A8�e��;F�p��)^f��T�Q��"ӊԹ�N�ϗj��c̉&�ٍ;W�]�g������|�+1}P�B��}��,	���z�>��O��yd��9�_�V�&u�ٰ�o�&Ω�H�κ�gn;��~��R���s1[^�4���W��>X��<{�9k}�I���pD΢���gnv�	4�
�̲X��e<.O�|H̎bRP�	��lU���.¸R��QY����Ԩ����A��BJ��Own�o��z�:'�ԅk��(����膄Vyv�s�N��s��t�b�Y}!),]�y��&�;%c��o�w�����J*'�� ]�Uv�l7'k���F�F��-�g�����߅w�D�V%U�ӫ���6�v���(^uiB�
Ǎ��?���K�S~��
�8j��z�Ym��	� �HCxʊ@�΁�O�kHD�(9ٟ�]iUFF�SgB��(�4�i��*�0,�twn���u��^��8�p�3]'4��o��ri���ł��T����0�qpr�@2�خ5�5J(����!�ځp�C���t���vg$͎�y=�^�������.���t���˖��/�K�ب͚GX�u�&�p�rsX��������!0���G�6hd����C:�}U�F/���b�r7@�6��.��1\��۬r�Y�ěG=˧y�!}hY8�!���l9����C���-'��H��㸖���F�����<j��c1�9n��p�	B�l�y9a�l�P|�5`ke�~,���-;6�;o�\�����A�馥���?޽
�%D)��;A��)Da�* 3���O� Q����،�K�9n~���H�V��bp�J�S���>6�G�Κ��"jWrH�.��XP�V�� �V��b��:�%�v=O�������J���Zw��
�_L+T �U�����pN�E�%�N󖔢Sn�пׄM9��$7O[n�I���R�����X��@�B/$�T汓A#���]�4����1j�'�O��`'����6�:�'*�ge3S�����Ո��r �UqV̓����G<\��F���9��5��cpǘ.]�r��m�*�ƭ���o��(���a]��c W�rd�>�>0O�+>�⯟G���p��)����Dh�	���^�S��)�T
�L$I�ǚl���[j�)�,��D��_z�t��[c��_])�B���b Zcs�-������M�-B{6�c�]��">^�v�_*Y
�,���|�N������Qz��
����u������!���?g�¼�!�0yuë��m��51f񈋖��ZJ���{���{��e�t�� �I����L�dK����� {/Ӿ����-1`��mC;3�#0���շnǀSIn��Z���΀܌�,$�R�M0Y��/���9����f�N$h��e��5�-}�'���Ԡ���vDL@��va j�hɝ����в�,�n�P%�:��r:W؛h�-I���K��0�6�h~��aE�.+��U�#���FqR��J ��_���NBֲ��:�����S��p�"��<�llȗ��B��h����P�/x��F�/)g�8_b~��Q0crD���Y� �BP��˨�oQoɣ�?�Xn�)C+t��y���i%g���
�t@���J�%t�Xe�}�|�l�^k��������c_Td�8E�kZN�f�;����UA�����>)qt�9���e�2�|1�=�b+�h��h������޶0�J��;hW=h���0�2'a�Nųrq���i�?�����z�$�"yf�P����k�6�F��o�{t�T�.k�>�O��Po}j 8ß}d��;�(R�Gg����i�e'�u�D�ps��ۿ�3-k}������R��\W��Znp@�<�?�Ar�Ȉ����|V�#�%#�dS�&bN1�
څ�mm2":
q;��0�K��J3;�ՆBu)C�m��X#؊�k�P��b�Jᗼq���[��3L�JM���C��164d�EZp=�S��ɥ<�����58�;P���[f3�e�x-Ǳ%m�{��A��s��A���A�Qa9ۺH�#~ԡ=���n-[N� ����s���.�*�/4kgl�ἧ$`=2��WJ�Y�$qf6r,�&0�~^v�.O!v�bp���U�;m��9��7��6(NY��,���b?I��"����lb��E��RyIZ��5���&φ��N�`t��Z<����7-���HTiI>�1Wk��]h�I5�>���mA&�?6�{m~8u���o��Ђ�����e��ַX�\��v�o̡~uU��>�vJ�?��(�n˫�w���n�W$ �<�Ml�j/,�����yY�?�ۨ�T��I�Q[�.��Rq2�5 ��ȃ��������mjI^&��rng9ff:m�!�7��?Rt��q�
���W���Gs�����u����1Z��b<A�+�v?S�Β�e�ÜmTq�#x���#�9?$�v��6�x&T"`͛F��A��g��He<�À��ٓ��sv��x�A��J��f��� �sGs��-���gri2�Lq�?<-�ǶL�M��Z0��|��s4�/1�2x�)�s&N�v$�.~Z�[l���dr:&�q�+���������r}g�;I0��s����ɼ�i5"�������;w{��$���V�aAA5ը@<B�)�V��3R-~���D�z� �wD�Nz�*�Z$���׏.R�������v��+�8�n�P��=�C��I\�mN)ޖ�A�4�� ����c'M���H�I��-���z�3_
I��j��l���^S���^{�&�וc)!��Ը���S��:v �(�2��Jk�꺄�����v��Qw�]�˻�a��j�C��LTWt�w�x���ېz�!� d;��T5ĝ;�����ܝtV�G o�A�s®�ڢ�t
�_���Y���u���N���ۖ֓�p]x�o�.���_W��܈��,�gh�9�7q����ٻ#6r��������m��7bN�վ p����G<�9�Bmz���L�/6�ڏQ��"�`�ʃ���x���6�+'��kKב�K��������u��CU&3xv��Q���W]�!�-��b7wt��wp�4��l�D���=%c�\�ad�����:���V��8�{i�	����C���,W05zA�& O����Ɗ\���#�X���t��0�1�B������D_W�2��K̗���'4y&!M��$�z��6���I�>C$�O&�bƠ'���CC}� tWګ���Sإ���/�K$��v(����c�"5*M�Qܐ�9��|̣�tۓ!�l��9��sB�B�T��e���w�_��o�)q�W���ڕ$C�RYH�M�>�X��Qj�:њ�$a�cM��V+ݟY�V�h��wd��q~��;��� ���Ğ]<4�����͖�F]7t�vxk� 
�b`��wTq=��f�Z���KǜrmI��!gG�����6���`������I�f6*IQ����MA�%��OᒓK�S���)&q�q]K XY�����	?V+X2v"6�ɽ�U$3�+1�9�&��+��jU�3ݦ���n�:D!7�/Ҥ���Ixc
�F�m�	�TN@��G�s�F"k���Ģ�{�.�F٧���z��pr(��'0����:7��wWf����� |������B���z0�\�kH�By�����O��8[ܕ�ǔ�i�ܯ�S��F�E�p���v7��a�E�`����!~;�ɽӜ�ecJO��E�Y�D�!}K���}<��^�� �F��U�[�y?c>߆��4> {dH�*��/<�����O ͡g1�=<��������!9t�I.kp��O����0�I�X@p��/t�^E��%�p2�Q��F�'�C�p�sg�2���'��o�l��y �%�oX_ւ(��x�	�7'RS���<����pF�D�����0Py�:�:�ӥ;9ɀ]�/�@Q�[�>De����#��b�`|�֦TR�@����/�7o�x�Hgk5�y�}�A�z��\"�ĥE��!�|4�vu�S$��c �	-=7y��S�,/�>�I:W��W:��*�¸}+��ȡ	�e4�G�ce�y�qZ�Z�w��L�:�lo*B�$����,K�����(��־NUN����`L9�Z�J��
\��8�A��`9g�q�,�*��?���l���VSqWHR��(#��~����͋�}'r�V�ω��U~�g3�8�?"�Y�`5����$e'-W-�O���NZ�G�r��d�r�*��T_��j�����}�{tiL���NI�C%UrK"�w�pl���mt6��f<1#H�E_���:fO�e\��j�m�����X^�*�N����#	dφ�s
���7cǙ��j��2p���2/?��	%V�:sbB[ػ%(���ML.]eࠃ�pj�ݙ`#�^�G&��D!� B�	7�i�L<�!�"++�!�e�~E�#�Yo"ot:�O���5�q��s	�ۅ�TD����^��5��ri��9�P���)x9�q������|N��t�P���8�ю#YVT�����`>(�I����L�"'2��Ip@hb�װ�p��"��A�])<��u=/S�r�Cq��A��3^C<7N�;5Y�&G��ͤÉz�ȹB��뽀�U�z����:�gh�LG�m����-@f�%��b�}D�ޤE���pd�.���j��G����:h�/_ƹDuNP^�7�����&�m 7e�R�7��{v+`��պC��r���� T�A%�48�̋$�~$�M9�ӿr�
vm �nmA�Iz��P��s����;�aFc�m�Rg4d�r�9]�js������p�V[:�Q�ɣ�0��tƞ�F^�+5:Ҥ�j���.g�?KT�a	�zDN��'S!�e	C�摃���?��������/���~�RJоW+ρΔ�c8ks`?��5��s(�͐�/+@�Ǭ.}p���ضY�wߊ
k5�C9�&͸�7�
�ͼԧͯ�ǫJ5o&�㧵���Q�����OQ���$w�a4h�d�d���4��r��/�5d��:S��6*4�O֘bZ��b�?>�z�������+��^0 �7�j�������SpMc������Ĭw�9����a��/<��Q!����*A�� �1*D��p��ۇ/o��@5_�Q��|��H�7��F?���y2��r�ƙT�6=8j=��0�|>�)c*���v�*'���5��B��8���-�ǰ�I��٢���]B�cJn�x��<ZWs��p[��f��)��s%G���BrV���c���z����D�;R�6��=��B�x�zdgzP��P�:�����y���*��������,y��Eh&14cN�d��{�f�O�g�ȕ���;��@[��:�=�z�*'ma��s�T��ci�bp�!'��B*�uB���9��,�_�G6���/�2@q�~t��$H�1�gT貓�F�Mm�2�!�=\ެ��Ȋ���نǆ�B	��ݤɑ ���\3��:����ݩ(y���Bpu�ɽ���o��Yq�l��~W/9��K'�wG���e\�Ӛ@;g��2�k���z�BYdⲑ����TF�N�:�K����&��w�����0�k�T����藛"�Q�M���=P������M:Zo�o�a���SKq�$�4��o�U�^�;�Qs��̈�l�l`�,Nv�/�zӓ�yF�ZdM�k�6���R�xv����	4'�/4�K�v
,N���j��e��c��5P��z��cA�T�uj�n��1*�a���4��w��xw.�Ӷ���J|�	�����aޡ�{y�0e�ĹŮ��w�����>a�-��~�R0?���a0�c':�XP__)��$�<�?I���h�z������~T880���x\�>����xZ�H�M��k0�#kP�tAf��,���r��;v���%<mv7T.�E՘�:���{�L���M���$��-)�T��<*��Z��l���OsՁM�4�KSoxcKv�⛛c���ŏ��`4�9(߅���4o��]?M��%T���p����,ﮟ��8)?��fU+�ҨzuiESWI�P���I�4�P5G�)F��R�T�ʘUʠUf���v�G
�6�v� �t��V����7,`Z�A���Х�#�I���M�����(�*��u5`��:�������Ǚ*k���d�8��`q����2]���֡f
R��f�۟�1f�fA�"�m>=1�L��4���)K��VeL�2�	��!�Y�X�������n����e�׌�=73��c7}��ph�kS��L��<��V+吥=��?���(��<�"��6��0r#<�l��l���Wʖ������6(�R�Jn�M�cae�A�[i�qSV�77�e��k�͕��R�pl@�Zn�-��I����{��y0�$׋4����x'5YB��(3[1U��b��1ll�(6��g1\�9ѧ	M�
^�n�&�8���m6�T��Y���k��L��M��JK@�U���H��%����na���%������F�"J�Z���M-���5c��]����f&F�J:s���~R�땧GY/d�jj���2�).�,�O���W��1U���[`��?BVT9�{s(��~%��&mMP@�Y�g�W�7��觟3��������}�k��#j�-������9&�+vz]�f�}��Z�˒����N����|��#)�f�vy���}L��gp<��a���ciθ`?��\+GO=��y~�r4D�4=Q�q l� �ߣ�����~Wq��1ψ'���L��\<��������x�$l�R)+a� ��3�\�U9D�;� ���Jyr��!�j���(�"~	�Q����d���߅_͍��Y(���A$d�Z��H��(��m��;�B�lӦYZ�#I��=)����X' ���I�{*�݂(���Р�XtvC��x��&}�Q��b��vDb�Q�\�.�q'AhPø��_����^R�Y�����Ab��4����EJ�f�L�"k�J���=������`��0���N�2�:s�8���%���$_��s�c�DC���á�	�'������P��*
1`b��#>IR�F�㛗��{�(x�
�?����ڃ��`����AKZ��?�򃻂��܂)�G�Q�h�렧��������H��C<{�c�t2a�˻���44$��R���AcPТ��FCP���P��G�GCG�G�Q ���R�H$P��R@��H� ���a%���&�� ���,E��'����[�ΰ!0`ԂP`�1`��2`Cb`��K񪙦+$SN��
�J�<�	��K2���W���a�3DŭEbS��F��r���#��4��\��lJ��̡.�~�Wk�A\f�� �Ep����1��ޱ��ӡ�k8���c��
(���_�vB}mUn1����[b䜞���MO���O��I�h��
{^���x���{�k�9�G��wR�͆Ż
�$A���k�k�����N���Q�q������uEn�7X.�����D�� ""� ,�oAN5C"�.Lkl��{�Xn��k�i�gGp+Bm���g��g\ݭ#r�*u�I�O�9�ܴ��Ǟ�7D�����ϊ���?��~�mUT"�+��G��;P60�6�C �t	��\�����m��r�B�������'	��������z���A��zh,I�Mt �����ۋ=K�o���3al�ц�D4O�9��Z&�sl����*�-�Z5�t��n�Bk7I���Q�Qy�E��9
���N�@����eT8Rr���
�2{�(�t��&���}�#!�n��n��E6qˇ���Y��F�сh��Wo����~�����V(F�~���dh��[s`ٱyQc~Ǔ�>�йJ�&\��0n���8h�Fz��cE��V�[8�w�x��H(J6�(� +1TX�ǌr��N`v�^��J1�Q�9/`+1�v�X����㢴��@����)��tFb��L��_�-��j�@`m`W����PF��ߺ�L٘	i�*|ʧ�*O@��z���@&}ۻ|ٷ��=�F��sXpOAC��L^K܀��c6b[��;��ٿ�����^8�`�U��	}nGRq��0@(Jt;i9�����ϸ�m�o�����*�]��U����G�$&~�r�sr�L����_H�}��f�f�Mf�P�S����Y��` 5ؠB��eI>G��?�o=�X5��%)C'�HcR�#5�$��N������-���Q$�Ӏj�@����C!(��Ug(�޿7sE��;��N;}Xwr``)���-#��ӢF�ˆz�*΀��Ȧ��E��OߜP�m\|�4��O��N�
QEC'�(]�_uP(�O#^��eqݒ��UZi|wd�}�1w�>w�B�iF57���a���S1\h& �_y	�w|u\	����_�S݀��j�]Ul�?)�|_Ԣ���pU���|H��.3�{�7�������޾�k�ߣ����Vfj��͟�>��ץ�|h>����f.�(� ��(4�͟�6��������xXW�
�W��15j|'��¢�?/�U�f�h�	w1?qb�W��y���f��I���P��<��pR�:�����(����ME�gp��q�7���$��y�0��ee-�w��b��$Ͻ�G� ��)������-�6����)��?��,ʙ�⺨�y��x���e�å�^V6Q�#hL�y��Q;��o��5�֍���Ҙ)�g.jקڠ�W��{�UlDw�j���6hn7]��k��:gl$˲�=�S�f&b��������e��9/��P�=�=�3�~]�g޳9�.E��MW�%�~�ݧ��&J��X]:�c���F�7�����
]��MN+�I�T�<m���Jح*�?7���u��4��F���`E0���������ߣ���rF}���x�H{'�!!�D���2��W��W���[.��l�2�MX'Æ3��� �s����MR�༆��bB�=�:�!�3���6+~w�ޕC��������!���iQ�#�f�C1�+C0ZN/"��x����4f��xRt<3�Кp��S�f�!�.�	t-��<���M1s�X6��ɍoF�#�O5��5�HJ`�� o�XY)��*(q?��C��!-='�j�q ��(���#{���xP# o����lud�?w�^/���L�UH��9���&�f�Q��i�8!K��l��n�îm��`d'�ǹ��l�&����ɗ&MB$W3�y�G��@��L�K���:{�N%� Ѽ�3��_��y䓪u�%�F-�B�庒��k^�����z��r��<�^���gg�,.����[��4�N|��H:nd��ޟ��4yE�uf�iH�O���K�Eʒ�tٵ�5�fVDS9h���U�����n�������5JVΏ	{��LN�5�����7KkNj���oo�J�f�(���0]C��t���X��L!����O.D����hk<}��yY$*R��q�Kv��?�sص�*�Z�_�+⺑F�AI�/0����M�:N.��r���K[ӟ�&�K��y7}�y,�gq���5g\�S�Z��B�+"3�nH��Ԉ'޷I���Gxs���T��:�.��C��*�ڈ��,���M"	a�BK$��F�s�q��Ҁ�pAV{���A$��RVq��\��K�qw�4N��x�HL�x׭T���0��PۖvI@�{���mҋ���VN���|q�×+�N���0o��D4o��"X�Yoį��F��w%��r�ES�#�Hsak�t�G$�3�˖H��[b�b��p�&��J���r2�^E6Z�i�֨=��P%��閣�1ɽQ��f�����ma�6�Ƃc&��{���p��M���`ی�	�[n�	����9��Z�eu��p��Z��\�lWzs:0+����h���Ը�dL��Z"�Q�G����Q��g�Ϧ�@�%mB���<x	 Q)ۖ��A2o	-�l~	�)�iB�+ĂNf�ƨ-��}��?����(��d�죕
�[C���S]���B��$��1�&r��=ڮ��3N\=�� �f���X��A��ʃ���yGm'�h�|}	Q�J�':�ȉ����qGo������O��c6��:����R��,30�,�Cǁ�L&�f�:h�#�����h�����R��J�Q�u���X�1��\��B>�>X{�b%�o=�0���gے�w�j��I��&�4T��X'H�)w,���2�7��Z羚��pd���j������O�����P���.M�2`r���)&��cs|Œ��<��M>v��
v����>���s�b�?�d!�`y� ϒ�k��yݍؑMb�Ez��6>鹣��	���z�د$N���$hg<�%U����Q�./�\�X~䟻������4����#7K�ԉ��i[��rǣ�
�H�+�5Z���55�EN�Uh�� 8�Ͱ�ˏ����bs.��f(��5�GY�.{~�xCiٝu��(ǵ�|�C��q�[���lBWt NY?�$%����g���b��i�yc�&���*K��	(A�g�T�W4dn��9|��P��gHh2� !�Ɵ����k�����Y���D&��3��*c��l�v:�
$e�$��6����vA%��>e��n�N��gD�\�*�t�~+/����W�n�F�� 2>�4xw�D9��۵̇0�w� ui�4g�Zkz|�w1����i�@%�:��4n>����'�,G��S痏irR���p�^(�ZW�o��'Č��ln��r�����I��W*8�=��?<���}��%H�NuzA�a�S�8�Vi��l�(��u���^�럣��[���<��ġ�le�!����F�q؋<�dhT�M� ���q`�Q��Cv,�Al���"�*f4"����[�Z����V:@R����s�Ō!�̙'� 6���lB{�"�P1���Rݜ2%7ː"Ǐęt���(2 �R����¯�w1L��"���5�`�>e�sN��_��S�/��#S4:Lo-�� Ғ@����m!,ͷt9�5�d��2���Y�]��6����EK6^�A࿑��˷�:|�9p�5o��n�E�E�/�d�=VT��-~��twe8�.�=-�L&���%33q�)����*\�U�/�Q�����k��rx��T�ׂ���	Q��Z�1�˜����ZD�+\qr˽�Ə��T ꭧr9|P�NҴ�F
����b����(F�GH����|��r���-��TWOi�}����,B~�[*��%c%�u_�#g�0%<��w���P�57vSx2@TM��I;��W��Z3�-�K�^g����C�s�FƜ=D@���ƖQd���J���+_��b%�kJ�'��V�G-<��rԡ��I��}��$�x>WY�ɖ�T�l��~�խ�Y��lXB�r�C����+��aD8�8�Զ����Ƽ�+��nG���'����+���rëL�Ƣ��9S��_���H�������&O�CB�����Ē�'���;��?�l^�>��;�ZދYs�!����蓴_��>�CS�BA(�=��fj7"ZX'��Hx����s��m������5��%����Q�k�4��_�FFp��vUm)�Tդ�����2�B/�|1�T9���ML�]i����+�V���u�V>��H
��Q��>;�c�+D�?p���b�]���SV��(��V��pS�,rmh�@����lU�w�lq�����e�G���.C:u�ڭ�z`"�}�D���Ld���{+76ߣ���̌.2UB�/3���b]d_(�i|��R��ҝ#��v���.m��C)�7D����)�.�l�~��Q6<ы��h�6[՞U~ٵ�C���Ŷd����wR�1m���P�<�put���ST@ڶQ65I�=��eV����I�a�$?X<w�!�-����p�ܯ����m���7`%�Y\�j����!7r���60�I����蕱��e�S�x��pD�+�t�K���<}��WEZX*,�p�,�1{qٶ����=zf�p�[���anC\V^"�.�aOM۔���̊������R�W� �������V.�Z�F���G�斫׍��ݥk�>��U�V��c�ȿ�4i�_V����;���GW5EǏ�^v��s�)�Q�U���L������U^2c�]��`�3��p�4XfEU&����|^�X��<B!^S�h�T�}��b����w�6��M�^{�6q_�V��+S�lC�ڋ��\���T�y�iH�㧆�1�ƞ���N>jT!�D�Sθ��������'�'W5L�=S�ظ|�>ڀw��b�]�]G"�\J;o��?���Bz�`�ظ��p��q���$�ْq#I?rM�g�	#�SI�]|�bB,B��j��P��a</�]���S��YF��>�sˁ@"�x
��L'\^l�����nCk���{��⃹�X�*�ו���ɇ�lD���7mWg6j`��I�w��˦]� ��D�ř��c�I�b`�MV���P�Z�M#:|l��D#6ǜ��/�W)ƶY�V��C�B2e��9PP&Ck(5�T�e�N���-�e��q�w�ФFa�l������\�^{��T���r-Q���z��� �i{X/��m��'�;�Nsn�|n*z��� ���^_B �� 	�4dw\����KDO�=Q0�9�8g����m9�~��y���IM.<��>�ڕ��BSH�䷭�V��~Nɒ��?*��N)@<��މ�R�M%�I��ޅ�p�:��'���$g�8���<���@�&��h�b|��5��v�%�T����p�5m��A�@$����t D��>��|�n�R��t/��X�x� >�/�_��8I���qQb	�:Mu�ū�H�~NX���-�@3HGC�]ޘ� �=ʴ"��M�#7y 9�q�U4@2��0�FKUIGl��5֕ȨL�h�r*K���;O�&0�KЀ7WI0���U�2��2mTD�'򷡘�Uz��OJ��:�͓�M&�w!e�8��L��o
�>O��7���g7֟�;f�-If2Q�Q�.&�䮠�oG�ۧ�&�����_y�1T�>����
�C�T�д~�c��I�&�me�m�Ծ�.��w�ܺG�d�nz�q(V|���	��-M::f�x,��Ϸ	�;h}u6���(�C��m)4/�|���H1��T?˫^�WF`��;��O|���=gdb+8�d9�ĉ+ۭ��%��]p8�M��y h.��j�4��c����F��AiF>]t2�-����wv���謫Z������OP�\���
bvDH��Qku�BC�?z;������7�0�j�T��2I��9E�h��7}��fCy.�H1x�M�1[/���Y'���ևl!��n��Z���e�6I'��,�K�����	TTC�K��I�،�M���q�$����w������ZЀo<���9���x`�z,Vz+��2�N9��L�b	l�^��QU���&m��w[��*��.�0P�dqh�b���Z������m��;�l�gQ�j' *�8\�dɅ}&�����J,2#��	`^�	t�gu��Lې��u׀�SQx�G���(�sU6c����kr:{�5��?��u-�Z��YA��;���kTծ�\5��#P-+�� on��k�ʘ���w�-CtdVXdURcB2���Ŷrɯ��V���J��|�:����� ��H�"?0�򈈐�4�3b�s��Z���W,߭��B��^B�g���hD������ vt��n���h��1��	��e	��:������V#1�l�GV�R<VHa����t�-��n=r[��-{�Y�ݖ��y�)~Ȍ�6ѱ�$^Y�6\2�;&zOqR2k}��J2Y��uL$F�ŻgĢ��t?dS�~l��Ho�c뱪k�4�{i�'��%l� 7(�S��������E�&7�{2iZ.��Rm�$�wA��Ru� ��˛��|ך]�6�V�%=7,�<( �=��j��L�&�%o��]۷�&#G�"�J��Z,�_�ba\K2�dvrX�i7�9a*��5�̓�|�S���"z���#d}�U���2���L�[i:�K%>�F�6%E�ʗlYt��u,��Ƹ�D�6BK���Dz`""��lh�h�P�ҐQ+Q�h�ƈ�3�Ȓ~Ũ�2���Ҏ�k�B�����5	��	���U���(1�s�L2���̍��Q���E�'�����	b����8�<܄�!�go[�Gw�ڸQ��.�:�[��`��N�T*��8c��5=�ȴpcޟ ��-�`yVêX'
�1l�"]�:�QU
��R�h�/�B�H���lsv�0��&�C[h���U�h���T��]�';�����H��'j:�E��*�O�I)�J=�U�����Đ�g�T�x�z9­N���]a�/��}/�� ��!m���&�X�����^�׋Za���Ă�2*L��QBZ����XpT���L��^�V�D���I2�S8M��u���>���ы�BC{�Y�u�	$�e���JU�q�L<�b"�Pl�����[�U\� ܅}x�_c>�/��+Op�dD����U���nu�\"U;��2`EPMTv��{��x'�~�ElT� R�[���PG�A��� !WRK�ܨ��ψL`�K��xU\�R�S���-�0���e��"/�}\�O�Ę�gX��]�>���	bc����;�`��*��~��Z���	��Ktü1�0�S�/i�mj��RQ�P����q<���#���m��dW�#��c{f�<(����J�_���m����֐��h��a!f�(M��0��&��䌨M�$c��G᭶��k&��xs7N�7�U<o8V��j䵇*����0��~��v��Zo�&r�S�F}�l��y��t�b������IG ��`�p�Oz�耗�!�{Dz�����|�'%�$�����'T��J .��4H!=�-:o컽������	Ơq�n4_��?�a��iK�t�hkg;��d�x�pG�_�� ` ��S��LN��"5$&Q�h�:;Y�D���j�!���)wv�L�
˅�b��U�&�%em�-��UhQ��|�Q���6��sB�eb�������9��c��~Y�;�|c��#-Cf@	!]�,z����FQ�_u�`�_��0Ș�de��^(�%p�z;�Tz��\;�uاD����Éuh�g�������l�  U�9�oW�g٭�|�!zjp�N�У�	�����()�"̹�����e|���A3��sP�2#,\~q���}�$k�놔�EC8��Ȍ� T��ky�2��1y@��=p��.U3s��khǿ1p��A���ܩ�Yg��0�@H���Ņ�����o՛��z��R�
�v�?��|!Wz?F����#$5���́�5i�G�+�Q4ĵ�6s`Vț�L���&�S`���y�՚�W����6�{�[h�	J֍X�+*,�z3ϒnUC� B�G��3x%�x��d�-��D��<-�A|����\�`�%�>}�.W�����P�s0噄FgŒx��g3���g�*��ضĖS�1�9��T����g����26A����zl�  �6:��VC�O�Ь~�Ss���#�٥*��g��')ksc�h��+D$1��*�Lea>jx>�'6C��#�\�j������; �z���;�KOpP�'���'gӨ={�2!1�7�Ɂ	�U����Oe�zl�fV^�!���b�a�E=5�n xc��=LI1M"�X)�Z���� [/s���iɒO��{���zʞ�fҝrP��Ӣ6ʊ�2�?rys|0,����� 30*-��}�m�K�g ::�6�YO8�BR!@4g�c��>�#�������^���Img�0k�}	1Ë�]E!-����e��1D�#-�`4�-,���z�b��-tVi�̱���Ș��'>�jFN,0t�1@����������-9�,�Wܔ"� ��v�Y*��p�M���(�6�tO�&�VaƁ��0�2��[Y|z�K,�[��_��_D��%�	��?��;�x��.�;�z��Q�;{W8�|Ķ�f\B�l*�U�u;L#X��<�Q/{�
���s�OL4`��">���-�Z����� �*�&+��H)���*
���>�p��\�|��Z[��N�M����p ���b�$��y��*E���rӪh?.z��|M�̑�$�9@��7�` �@�Oq��W�	:���؅&[�����݄�,��;(Y�Sʧ;���n쟪��7��#}$�� E.D��!�%r㧮�M�]�(a`ǅ�#n�~�m�8R�_7��z^���)޺�G��ƁE���__��~���(�P"�tgD��{y��E[C"��Lyql�c�ve�c�	�:�'WA{�/b�=`.�b����6XA�m��$7���~�X�k�9��Z'6���"�s|�g2���t��%����,^q���h땁���˂�K����J��Tޞ�S��:p���*]�܍�`�����]����*��z�ۜ6b�Qp�n�mKd���/�de������Y�z?o����q/��k�Ԇ>~#���«-��|�3�����#d���y�Wp���X�Nwu3�X��H�c��<כ�[��ˑp���|�� �NGt�%Ukvke�
SL�+�ODlF��5���-�qNv$��/�J)���q�h^h֠�Q�AC�ň��&����*�Y���@��S?�{!�Br�"�����[�7�X�RQM��RQ��� b���x�r��8p���4�Y��ұl�mR1O�%�c�H��
�ԈeHqg�z<X��*7A.�i8,g?y��ϭV���F^X�tv�������nƻR1'�w�j}�\��@`'&� �"�V��&1���ե�B���t�~���"8�k�0i�Ґ6-Àݧ��Ϗ�!Pv���!W�f>��q�%\��!%�Y�b�L�K���,��c�(�l)H���cs��D<�/B���G�����]���τ��z������9E!a��)2 ��Q��c?����~DcP��ʣ{8T����qU��ww�1�=S��M7�:����S	b��*dj8��߀��%��UrC���noo��B����}违���k�X><�nU�'��a 2-`f���'Z�1��0�u�C�L~b��/��2�p�Z����w^��wr�)�cZ���]�r}�?�[�+XB��dr<ŌmM �}9�+�ͻ[5��
�s��0�3gp'0����; �7`�A�Ҫr`���N���A�@�N�K�zA.*��#��vS�0��y_���1<U(B-f'E����Q�c� �IÊ7Ț�
'���=��W�C*k�$��M�N+���"�'���M�J�?~�HP���&ڢ�[��
d���
����DMo]HN,(��d�qs���`K(IP�z>z�6�VԳ�x'gH�U�}��U���.����G�XB�Q�U5�r�����["�?�<(�?ѷ�ˌϫX��'���ذR��²V/��'������.�*��z�Z�)Ҭ�aQ��ZG�,���DEi�O��������YA��
����z:2�H���,&��-��x�����g��4AX��.����`z+����;�_�&08z2�19 �ntȱswQB7�%R��:"+��2Or)���=��ɓ�:{�֧���@H��h�o��fQ����?���H�r!�=kݪE�ސIo!V�~x��ی�HV�D<�
�Q����p���G��T!�Uʯ�]�&���3J�x��8(��-Ie�8hG�E�P�lF���|�eW���0��`�ԍL�b�1_ǵ2�<��F�*m!��H��av�fX�a��ɽ9�����#�6n��l��a�G�s=Z���5#�,�r!���T��D5%�2/z�f���hk�Us�Ե�;cK[k��� �^d^�����pz�t�4&�%�oe`��t�`�7f!��LY@�f1*R�%�D�9���G��Zg�O�-`h���P�<Ɯ�y��Ѫa�s���}��u����p��1	EBQ�5c0���>�X�=$�����=WQ��X���\/����� 2�{���R�iDӓq�nqA~��:Ff��{��n�G���?ޘ���Cﴯ�C��BS�	��!�olMnA�&���Y&d�d�$���R)Y�'�剆$n��ιu)lq������B��xS3�T�%���Ǧ��:uv|r�1�J8WMx�EM��r�x��j,m
���vZ-�Fk��-�q}=vǯ����m��sn֣r�F,�q�-F�%�E�P5� h�1�U��K`4�if�)C6��� �-���Vm��
�]Q�<b���ZI����(�)�T0OW�����U[��A!��n�0G��AF\���x�ͳ�E�����JdyԜ�A�l�����՚8����l]tL"���D���T9������ֳ> sFp̜PLF(I�����Bnό�FK��+t�<Ϗ�)�?��J�P�_�
�]S9'{uد벉�@EO����R����J���?��t4��4�z�/~�S9 5&�x��z��nE2�	1�K9
�������_Bx���95w?ƌs3����7��t	�_�n­�/�^���M.��[r�`XTa�W��h�OA�83
�R����8ƪ�x�?(G�3F�GJ����x�F����AWsO�Μh�_B��O˩��oYV �>�Y���g>DӖW5{RyKkL[�A>J]eGQ�&b�t�y%��2Ѯ4h^�O��fs�ڮ���W��7 ����3-Qkd�z����I���΃��*�F��L�~oE:�J��U]�"���҄<`�s�gf�]g+��&!�9� l��+V�q����w&&�kܗr������K	��|�/��� A�=Ì�|�-<ܠ�m��ٰ��-����
��K&ʵj/4Ų�kD��!��?����у�-/	<��
Q�L�H��*�8e!�g�i,@_�������f�r�Q); Ӫ��:t|f��z�댍�q@�NKg�����\�ï|ق�������L%�˨�H�`�N�z�\�!RP4�Dk�U
`�''b�6?�9?����p�`�#��ڀ������Kp�����x��!��������.PF����fsͅ��F���� t$[0 >p.z�J���\�s��� .H!p��߰�&�0/	8^2��P��C
�M,1��h�/J�L�E)(����s_]�}���1�H��*�q�B��UxLYқD�;dY��n>�x���hQ�6C�J�1�Ho��\�fXx�_�=[[
�L���j.�q��qQ1����f�9����G��}UH��S�}[�଀�hLhb����4� ����{لR���|l��)��xuK���i{gy	[D� ��&������힖7�z�rOH�qF�a[Q��/lZ���(�9��=hF�s��LR��V�9�5�[�ك�1�Hn�g�[+�ȼ�؝����i2S��7�6�>>�ϥ�O�a�>���R(D����jy��4侈E؛�����Z?��-���g����4C$��O��-J.�Z�p�5���߅���kv��ҹ��w�ؗ�W��.�
��U(��]�+�ܐZ���,Ÿ(>t���,9[�HZ���sX���I�3�O�T�7� \�:H�-��<�W����y�z�6���^L��i
#���q�߱�k(�e�o'�;�y�����]���&Q��2s�$݋��=��ځ���S�վ�:G����ထS�����0�L%CW]E��8M] �X[�ֆ�P�U,�d줈DZA�������#B��dE�R�@��a�RC�W��۪�rTE��r���rQ��"��Z��5}T��@�j @^����������T�1��n-H2'%Vq[��1�r�E�Fb�W�o��
� +������z�m�4R�C��Ճ�gUr�;0�X�	fF�\�'��&R�RAR�%H� �A��Җ��R����-}HR�*��_�G����[���?��Ѯg�,�u���E��>�f�����"̋�6k���@�1SpS|����
F���pE� �
�ŷ5��
/���N�	�� 	QJ��z��&9_bm��S[QM@ߗ���e���Pi@̐JT�
:�$pdB��1T�R��l�\�ҥm�E�2eI�.{�
X'�ܒ��k�`�R�J2��� �T�d�҆�S��⅞��֎�S�C�ٕ���8�p��N��;#���|��A�8&bB�]R��z>��R��@�m���ඉG���.��,��J�-&0zI�W0��+ ��7�"?�i>��Il>g{R[v�H.Ѷ4H7\Ѥ�Ҷ�G��m�ښ�G�B��1�8_0^�����L.�k8s�c�������'n��[{UM��1����,{�x8�;3p$������]jTj�%�;�1��7�q��0]ԁN�2�~������MH8U�7G��|���P8@O�ę� ���<��؀��60L�u�G�Z�9^����
ʩ�A��T�]\mz�6��XF{�T�m�6�����a�p�v�X�1Y	׮����~����j|G66l�6`@bMx  �&�q��m���16�F�3��$m�`m�*@���w���Y�1uo��_��������.��ӷ�j%j��8U�m�\P��E�ޠ�.�|YKVx�hiOGQD\��v��y���W�`/\�/]  ߹ף�ԛ+t�>�;=S=47������-��jUmq;~�搿Kw��'Q�ӷ��;~h�
u5)t�M��$�9*܊�0��{Y@�Q���'���J�%A�f�]��O5Q��X�qb���Ƌ���Q9�|=��>���7*@G7��B8b�F��f���1��E��+[�C�g�����.{$��X�:�ۅd|�ԕ��=C:Ϋ���S���}��6��	�?������l]&�jŭ�ʭE��}�Dj��M<������ʗw����?LT�;�����Z�XMGu�3M�����^�eAK��2ƌ��y�|�e��J-ҷI���}~�4�Л³�҄���+�3�c�6�)�W����^�/߃-?�)p�p��%����4b��(?�O�.j癶X-��h�_�O�@"�@0�Z�M�ܯ5��:k�w��QR
��Y`�v��fdc,�A*�����Ԃ�����K�������o���B�ט��%�6����g�L
H��c4�t��$j[�F�)r��Jch�֚�����]K���B�[ZR�^����d�p/���ׂ�0�W��.	�7�ؼ�_R1����:1��V�ܖZ�@,��8>��u��7�=�D��k�K�5o��V��Rjn��p�Q/�M/����hy/�K�|&_��o��s���o\��UtU!r5�4��������Y�ء�:�+��5@8kLh��Kޘe���I����o���@�J@�VC�9��+�v+��c����j����-F��he��j��,��MOf�v����-)Շ�|���T����.����/���W��c�̈3�ݖ���++1%Mk�5��`�W�57.�]������Ui�D�Æ�"�h��Ȣ��x�D`Km��(Ru PC�9Cq�X�����KN�6�L�uM[�5kw0��?��m[�9y����v��>�x��:����Plb���t� ���%G��LƄ`�۾�y�fJ�G�:Wy�=l_�y)J2�\�]jFm�J���?F����!������M�O
�D�nv>� gk��5y�?�X�S�R
������xXq��H%���f�+��H�/r���2���۽Ih4,��a-�+k��VUC����I6�n!{�\d����$
��(�����n���"�M;P�h%=|�,h��e��{B�AeY��TF��5Vh��Dhx�XR���A�4�
����)��ݹ�����H�[�P����<�f�<	�v�4�q
n����W/��E�9n@ΛK��J�F@���.��\t_�Sf~Nu�	3��I��[~<nx?I�)ǋ���G�����j4���Fx��I�%��0sM)+8�Ź �經�)��c!~W'MĀ!��($��dP�b�H�� w�re�:?���o��y�w$z�t�Cظ���ʟ($iC ��C`�:��3H�!X��N��
�1���?B}!+;�����h���_$��q�%���/��)��HAA�xϯ�VfF�C�k��B<R��S�r��X���QO�t�~�{��v �~c-�7�"�_9c���(���O������`}p��<|Vc��}C�%G�fn�[w�<�OmYGF��]=�WجU4�IM(Фb���x�@�Lƣ����NG?�΂;#ˮ��!�D����	�~H�m�r$����CeVw��E��;���Rg�T�C3s랼)S�A�[4�Q0���ߣ�(���8 T��A?ש!��t��MN�Z4�����Kt����1&M[C��ي�vE)	H(�Z��8Є�.P ���?������/Q/�l�˝�4M�,�3���'a�����Kz&χ8�t�G��X/F���C��hI��{���Ao�jD@9 �gN'O��Q%�w�aWX� 9J��1�+tƙX�,�2��{*S5�tv�����,W��T���߿��^Bw2�9����_'9q�>u�7�C��0�9=Ũr;���^0���!�V<�/�����,��\�+��%z�4����ԋb�<���<�^�L�/YU�Bi�id
,I�8���ƻ���q���B XY����8�3|��G�R����IA`�-f�.��>\bB��0ևO�ظ���Dܼ�����гL�g�L�'�����DN��d�,�,XtP��N3�>ͱ.?rנ��zڠ�4��5tb��8#��=�}���9C�첿��'�}�ń���m������W���@�<,~y�篠��j����VD9�	��@J*����ޞ9��\
��:���KS}�<փ3">,OF'�N��RT��+��~����;DT9O_ȃͿ��<`4 O>`;0=S�v�N�,WUǄx�ϕ�VT�`�{���!����I���6�s�( R[�	j��C��W�l�EG����>���кʦ����v:C�H�݇X§0Qj�6bDY�R�M������4Q\�&y�0>�F�?хd�?�8�|0�0 g���|�Y�Ѧ	?�X��ѹ�)�h^s�	c�!o��a8',�ȑ4]@�k�L^��s�i���ڌ�M���J�4��@[��w�#���*Q��e��E�HW�"����ZΓD5�P��<���B��X=s�kH�C�@�4GL��kJ�Rצ�'6̚��;�5\�e7��,��7&�C���f=e΢�yh���6%�����Ѫ���4���P���T�*o��d�)���,����˂�6��[�\��B��-�[��A����D��WԴ�^UC'�S��/��\�f��Q����8��<��U�T����vQ��2�^r��.��@�<e>0Q0J�R��$|�^AT4�z��BKy�{�]pD6<����ίb�̳���1v��>
3�̴L������s�e+Â�����6�9����]{%O砓¥���4�K���F5:� /D~җs'[7)��� �z�?K/��F	� 1�Xy6{2����W���;�:��<`���bC�'E�'��aWƇy���r�Efֈη�a4�H*/'`2�Qx�c��N<�^Q#-�Nj�W����.�h�����M��ǃ��5�M;�G�Ǆ6�����8E��k<�
�@U0a$��=�T+��\x[�y��?pBH/�򒲃Ӹ���<nq�-���aT�GX�:��@�O�n���#��cE��8d�5:���i"�C�G��g���P���k/6��;��o���=g^�|��zy���P�;�����Z�KTU(�EX����&p�?�k��5�18���rXr��)�o��[�;SП��A���,�;=��?:5�wDc�U�����įc����Ruvl`��6J��K�����j�l`�K��t|$\��n��h2��ګ�Gp^�Ѓ����(�%߃�l�Y�i�~Q�D�^D
�	�I��R�3
����Y�����A؎|j�G�q�[�N�z�vM3(<��fT�E�y�g�}�2j��F�&����j�]$@�CU���{��s�w�	N�$�/�:[�Z�.��c3Wdh�虣�5�d���y���edcB��'�p��S�:�/*ngc_% �����\�&_5!_~$��~�И������$m#W\�M@���i���>Vґ�o�ȁ$@����lf[���j��M�����-�0a�1n"(�&��I1������	�RV	p�����b�W��	�ky5�ز��W-�L���ܜ0N(_��s2�8 9tg&?�C�x
�GָA=��Umvqe��kq�ƕ[v�n���l�����/�9�CH^�0�U"�!��<���ݗ�/���([��rZ+��$P�ڹ��?ԊN��du��H�cݜ6���q���&��pG�}vyX۽��p��s�ػ$˔���|��%�)O��P����'�0�����a@=x�}2=̀�`V���a@�ׂ�1Ʈ��/���Q1��k�P���4 �=EO������W-Oݥ@[��G�ʝ]/5M�*Н`��`�}G�7_�z7u�}@��f�h�����.Hh&Yڼ*���=��F���'��F�^HI�9��������_���^3o�#(���dZ�r �W�f&���W@" �I�S��ı�ٵ�-PB����g� m\i����C�b��_��D2e3a��	G�k���s�����m���C2Hc��g�x�뭕f�lUL�Z0����!S�.M��q� " E�`d���A�O���?�Z�ʀҿ�_oʨ�gY���@]�������Hk�\G��4��x!�M��Q�`�L��yZ�ʜA��ob|�]F _�O�3<�_�&r�~�.�q�ؾ�>텻(�����6��w�b�2OD�i���4-EJ��ᛔ�{e�`7Hk�1�Dw�/�L��/�6Apa���d�m�"��,z
m���,�l{(:��ap��4K�#��v�%O�@��.�ӁW�SOŋ�w������Vr��vOz	r���찁dw�3@�.'0�����g�H��F׾v6�|M�S�:+-��F�X���MkH7w�=D��u�i��E~օE�3җ��3 ��U�ݓ��~���_�����S�w����~�>1RH��>B��C���%=��T�n�6�8Sx��{$�2珡�Y2+9'㩱aܾ�_~w4�Rke��0�6�2��ə�і���]^�G*TRI�4�8���b$|Q�MGJe�����X5#B��+�·���W����AZ�f�z��3���pk�u�������4UԶgڬY���fʹ�}-�����γ�C���kI����1��w����������̍�h�.=W��+�Oh�b[�>��r�Рo���i�6��
w�hk�\:�h�ļ]ԥM�!���\`v~�JH���TkMQ�U���U�g>�3w`8pV�R'�1j���G�vS�]8��d��'��@�9���s#�]%ju��.���F�sQ���� TF}&ү�[U9�G�����8��-)�tdv4Ws$��p�^�~~���}��|]dqggL����"�s1G1��+ ���� ��F��vy1�C;z�mj�M�5�˪����]��g.�U���������u��)�Mc�qx�4r�8�"s�C�,a���MQ!�F�	�*�e��u��z��i�\�^��+�!�&/X��!����KB4���z�ϻ����v����+�rt��{���8�U��C
8-��
V���:�"����5 �N�����&����3� ���f�Im����L��|q��6���%�J�N'���7{j�<�7�ܓ��n���܌%%Sۯn���ޝ�Z���9��w>�k(v,�zw���� hU��^C]rY�\!�H��mt|F�U�Fc>6���T5����"v7����s�^v�̰Mi4��k������'�����5�F�@�����~Ͳ6%G�t����M4�nI��	�O�C�i�]N��̣�m��|^²xc4�	
�оx��a�#W\��|{�e>�9�rJ�(R�/ݏ{� !(S�����zO	�Py�d��?�31��h��m��`�Ln)�E�{���`fI��t�֥/t)\	!a����#�������v���a9��lMY�p䌉�)��>X��th�Q]���m3��rky�*�J�33
�އqW�o���2�+Bb�Bॶ���b��^t`L�*��3���� ]��Y�@��Ko//�1���;b$�}B䰩p�/��:��:�;C�5@���@�;�åZ��.l�IdȠm����䡣�rorƆP{m0���&U���Y����>��'��|�/
�bZـ�"s7��r���,D���z��Ԝ�y��jDx���#�7!�;{���������������h��"�J�^Գ"�R�*(c^�3�êT�X}
n~O�BO�I�狏����<.��	�S*����{�$��b~��M�.����_~����k��
�����}k�����4�o`�F�D��4QnH`BD��؛���c�&���{����.!-	h��x(p��r|%��F��kEP��4-ia&�3\Q��}2����4�/�ρ����u����w1��i���V���,�g�-��lZ�VaT������4�驮�'$��~�F��r��&���l�#@�UU�������;R<�r�����ru2��U��3v%h��7[�?]���.2Uf)r�����/]C!��$Ҍ2�ʨ��b�xp,�ζu�UI=i?iq�����)��`c���;J�;㝌U����ʩ	_�e�������W�Q�s4uZ��`q�"��Me7x�MQC��x��f�v� ��1��[�-��+���8X�1����$��j�x�D�o�I5T`�#�~~^��E��@��,�C��?���_��V�siv��ſx9��oNhl1�^��Q�,<���@�	Od�YK���ͥs_��s����$�I�KqQ���(�t4�|������a�͘%�W��tA���A�zї�1�^d!-:<���e��H�`Գ������ߨH�S����la�F������PY��.��?N��wZ���sf2z���Z+�l/�����,�̀�i3�6�|z���&��7g9���Dg�#9S�r ���H��Uy�A�I؇�dOZg ^zNVkz9�J%<8!�Ƃ7�s9��{�p�C|#>��@Y�TŤ�C]�XVIB���Q7��c��s���t=b�D���u\�Y�l�A͑�����"^S+�bWk��E��O�Z�Ww�jNp	�g�Z\D����l�/�y�"��'N����
#�����K��>���Ɖ-ϰG��9����}�<����H߷�v�[\�ϲ>H�"��%�$��6x��Ǎ�1�9_��LWO�Ef�:��4�)�ui��|u6��}KH���Z�%@��w�0M
��6Z��Sy����g�=�-��4�i%�a3rm&,�����sQt����!��r2�4̜w/���L���>jɻ���վ�������������i�H�T�FF��\�Q؛�I���}*
U8�(�\�#',���"Ԭ1pz�-���U˘�xI�YA���;i�����	�3���C��S ���6��%}�ѭH�%ur=��[N����TH�\��i~nO�[f\����s}��H��<�Ō� Gk���Te;�&��а!��e�"O�R7 �~���u�����.xo���0&F����>�k���]���&ק����>�L�~�1��<��� r�M��l~�U�8?�3nzl���P�D>�$bؿYD�#�\B;�ť:���y��%����^%�����d^�wOb�*D��ZD!�y���!�!���+�ހD=��&��a�� �e����C[U�Of�e��to�T
SU���'��z̬�߱���qrL�RېU��)��R679��3�J�.(98o�B���HC�0�[�ϫGxT���}7���K#�?���R>~��;�$B�Ӡ�*�\��i��ƿ�����z,�OJ��Wĉf�J�(��|q����z�#��^�m�]=9d�����*\N��\)���[rmB���=,I3��>�r��`Dɫ潶���а7o���Z��,֝��Ȍ�d�jR:�S�v�2�l�B���Fl��UI�����SW1!AYZ���o�.�j�{uSp��G��lId���$��ݦ�n�M�/ C\>>@7��KM�ƌ�<�����0�ÍB���P���Zܡ�d6��4�m���dlK	͊RѨF�<�� �Na�MD��_+.��Q������1X�y�Ȃ��l-�e#j7�ʭ��%�j�/�d�0�gt1{��
RN"n�"���8g��P@�PJ��k#B+V{���ʽ��H �$�)�/�Գ)�:�2˨��ԭ�c�T�����U2d��aK�M���Ru�g�����E��G#��L;�0�łI��$�|��wj���L���b�_*�8�9&!-R�R�=�4�j�,,҃1���/�B�`1` Q[�]7w����`*�=�*���ǜ����#���`�p�T�9 K�Y��ZJ�����NE���Y�uu�� lb��e�s��c������G�B�����ÎӒ*��}*��O̏�z�*���I� k02mZQ� ��KF%�ŒF�����Wb!y�0�d�|D��P�f�`�I1$6�xA��D���}eǀ��7W9�W�<l����ك�B���4��A4����f�L-�Y{�)|�/@;��Cd�\�&#�̌}��oy�w�ǻ�u��@W_S)���us��9�G�J�(� �@ʞ�Q��܆AU͏��.��j��6�74¾�O����B�y�Y������Ϗ���i ���8����H�o�g��h�/#9g憦��A���������o�4�v��X5�E-~�AzLe��@�P7����\�Ê����{E��f�x�-�]���@�� ��h6�j>#���5.L͜M���* �S�Q,�>� [ȅ���ҿ0�������,����G����C!	+�5,/�ҫuo�[d%�,'?{+�!
�T�]���<3\}�m`G������R�|*]P��ބ�Wɗ����#G���@P3�3|�ʌ2)�]�ò��AKЏ�b��]d�u��c�����g�Jݏ�������=�U�a��]
i8Ak��C{���DJ��س����YH{Oۻ�����3�[�jC-`>�Ce�&�2W��[�I�s�9��O2��"6x�Mix��SY�y�;|&����0I����|�Xˆ@}�9!�r�Yn#s�������8l�-8uf;��S�#��_��7�w3Q��n�Mr,CH#%����+�%��5Xp��z�O��3�%֎�+G�)_"�Z�6ʼ����V��龼�}B�WS��bFn�X�!	��T�jck1�	dC\5�0t����8'h��R��7:'��g��G6����Y񛆀��Pn^��NBGH�LCE���@P�s�}J0f���$�
d����""�%����:�E��m���O[QV�A����b�q|��*�R��a-�Hǵ(y	�ȑ�)���� n` O�t
2�u~���ޤS�&b��#+I���u��.�������J���zD����_�Z�,[����8�.�<ȼ���'ʦ+�%�/�s[#�oP��OC��qnT�)�Z�c0x�gǽ���nU������jd�n�Dt<����Z�> {�+s��E{r ��2W���נQ=+!w��s�% ӻ���V2��>�i����rK���ƾl;T��2��=�x�Ha��Ahۛ�r��ԍ0Q�)����y-	q���$�[	�m��Z��Д8tx�M��c	Ǐ�������N�o��W��G���*���gv�
���SLf9d�S,�K���+�*F'������ޒ��irA�ӭ�R���B���{eIO]��)��y�<F%�:(obԳN�o?�фGmt&�8�j�	8uj-����:l�*R��S�6��X苣3����@��]���B@���w����䳈�s��$PӰ�Gb���z��m�γx�s����W/'�pW�.!-�l<_]���h4�{hH�4�q|9���T� �T���?��+lPy͂��'�l�M4h�Y~_�&��t�
,[#����ښْ!�;�k�����O"�_�?��,Z��xF�}�YE�_��꩝�V���G���V+@1��摏	�R�]��>�M�x����8fm�D��H�W�qe23��M�t�S��A����֔�Zq70���^�S���3{����.i�$�������%ps#����V���"�7��`D�>s�B_����)�c��7�*�?Y�äl����Z˱��7���/�]��T�#��`ܖB�0��h �W�
#��$o�uU� �9 �]���j��}��A��f��i��M�,IK��m��LT�OYhZ��e�m�(c)��5�A|�=iG�;�z���O���K8�fs�6�Ei���D���z�1�������̂A�9��r�,���xF|R{};�d $$A0�����I�q�]b�64�����^�:J����Ŏ4�^a�|�Vr'���b��aZ.���UK�)�8�9��7~w}�<�xoI�0�75�F�8@�i���[�U�ſNr�)�$�CJA�-��Y]���INM���)�8b3���D�PSZp�sJ꿏4ݦ�ݽd�ۚ�{ֆ�b�Q�=��_���Q*#��2ڞ�z2��^���u>����ң{��/�kKyR��'<��œ	��4w����U����L�2�qAD�%N(aE� GM�40����+�������l[��۴���-Lp8@���o��ӵfԔ�� ��jOy7��l�}�g�x��l�E:	�\�� J6��2v+0���Ӯ<$��CW��O��zD�ae*m�Oğ��'j:cV`8Р��Y�䧸�^�~C"�~�5o��Sb�t�D�2�����$\��r�7����M#9s̝�+W�5V���#d���y���Dr�z�@������ '�P-���4^��q�{��H�5�O�b���~e���P@�l�j0X`K�!�oA�������xU�~XX���`�dr���g"���t~^d��ǭ����o��� `)�|Z�c\�=^G!z�=�X#p�\�I�������x6N��<>Df��/�ﱝ�햤���;�!x����I:�����:��c��>h�}�W�h����Ɛ�;��#�199��i���H��h�u���\pn!(�z�N�,K8�����)6����J��|XY �P�r��ը�N�����;�w��CL�s��I��s+��S�0;u�俵r�3���9�S�K�6�k�@!���K�@�<s�ЊYM�����y�h�Zi�����9ld�7��X�ڷWPz�,���a@�9��P2;����^KA^lL�y�
Όu�_ ?xW�7�Uf;����C�B���P�����<���Lf��Ȗz�g Hg���[>N��o�#�a����#���j�g���T�|M/���q��4ڂ��m�,��e?h�!��@l�����\ ��6��l�ښ�g�y��[�A����@���`Y[���@����3_6��b�[x�.NsRי��ؙ����(v���S�.�M��(z�C  �{���72Z�6�}xe'�/����#��J� 0-Ȧ�M!	CZ>�O6D���U<��u3�B���t&qqo��*�7=��E�~�_7)Y�k�~Ԩ��PM��c�84�F5�$� ����g�%�:-�"#��#���z��M��8`�;���΁��”@��
�]>#��)�*�BK+���5f�(�;�|���~��@�s,t4��(�Ϲ�	��E�'ws)�� ����-h����~��<H�l��+,���/�?�*b=9�U�t�����S�/�mg�F�����������N�x��G{,6�'|�Tg����C��:\�=d��D"WII�kg�@�wDn��OƼS�x]3���f�~]X����Ѝ�f@Ch[��k�˧x{r%��Ҙ�EЗf�0� ^���O 41E�bAg�.�)К��(*�2�<���#��8�P����<��>�c����ƣ��?�M��<(�V�{��:^ٿ�!��o�G�r�S�98< B�R&���'g�����z�0w#�C_s���c#Z��ɲ�\k
	yh��5B0?7��sxw��c���p3 ���bSv8���r�.@�BG�_�C��4'����nA("[\��Q�����y��?�\`�*�a'���^���D3-+��B�H���4�i�oR8n��cޢÂ���S	ɤ��4|��y+�rrH@Tn|�H-��a QS��泚,��.z��b��a{���!u�Ux��Ă��w��fG��들m�HU��d��a��-�\���f�c`8
͜F�e��o�fgn�Z����Ʃ �I���4�E���M(U͚����B�Y�'f43>��Y�L���������dl	�DX��Y��-��p�����{Cz�Mz��6�Y廽��d,�i�-���e�1^3pf.]�d�J�Ny�[�_k���wa��(���m���f
�i���.��/��}��W{���1��&�W�[|�^�W��!V�&,����o��%w1>�`v��v��,Fq�5`z��	� �!9"PT\��ʉ�ao[+���9S�"�Ҡ����]rYZG�R� x��Z#]�!�/x�o8$}���-���BEsy�+�΃�?|E�~+�(�W����`N"�h~�Ȫ��9�:����O�z@4y���'��d��лq�XC����)�ܡ�V6��Fj�W�D�{�"�tiv��R��O�d��Qco1��UȂ���fj�Ȑ�0����b�J�I6�����q\�u~f:D��&*�[�7˸���r%'�3���7i�����͈��C�KW�a�ª�R��8�1�]c��*^��Z�=�k"yu\?�m���J�ִ����C0���Hjb��K�P�6s	�}1-�?�D��k�Zw������U����8��t�=��������bs̉i��Uπ�<Hi���"sb/�
$p�}7���	�X��˲�fK�,��57ѿ�wZg���6������1*�d�Xt5���`�a���ȼ��L�|��O�K�$�!L�<� dS�.�����U���͢�gq��e#=��֘�k�bo�?����4;�E�D7�����8�����,�T��i�l�+=)�����yb�S6vā`@�1�3X�!���ځg<���A8Hѡ�`D����䲧اh�����K�&���{��Oox~�R��� �E1?�I��n����®�T�Ze��,T_��v����W�,�E��_|����[[��#��w�#�J�Û%.�}\�!1ސ/V�If��a*�n2mg��?�' X7�%�:����� ��{�ƑS�H�1�xk�K~T;��.m�}��6���%#.a�C � 'f���v����'��D���ւ�H)Z�mڬ?�@���54�FNT�S�������-#��X�tYۂu��ș�T����+`J�uM�L��y��G��͔�M
� C��(um�L9�fٰ1���c	������0�C�]D_��{!d��/��'�M�P\i"hPh5#�H���/���CJ�����2E�v�W;�(d]켒G����izfj�
�"@�eo��5�{'\MտjBfG��_e�>?�u���3�I&=,������6OؙY�l~o��<��}L�H�G�}i~���S����R<����0'�z�������o����K�=E�U�$y���3����L�b�ݘ�e�[��,iH(ҦZH����%����^F�Ԫ�+mm� e��N���� �{�l��:��<��ל�=�.��3n�m��0�cՄp����m� c:�@�7[� `j�l�� ٰB)O=_�7���g�a
�~s����~����sEb`k�H��@��#��t�4��QV�ǉc	M�l
������/�D�6��j���U���"���"045��9�M��lb��4��(
d���z�w�%%��l�s�>|=��F�_��/f>�a�Z}��%@Ƞ�7�fb%�voKR�W�t�xG�Z��z�lv���_�ۿp�3�T�ﴇ՛�{'�8ԋ�&�1�uݜdKʺ��\{�
Q�\�$LO��X_:�Q~ȋ3h��o=��p����.b&۸T+��r�}��#�[7YǴ5q~��P�CG�/����0����xnU��μ[ ��u���c,�	'�T��_��y�sp�sT�҄�-��]��USV���l�CF��c\���u�����N��9�o2e/���:P��K��fz�-���bڰ/���(�'��՚ֿC{� ?|U��jb�����Ɔ-N��:�A3���j��dڙ]�$̺դx�Ʋ�/zU���z?~T�ϦO��M \����=ԩ�~�i�g��]3��str_��B��i�+��z�h�^����}h���԰*����z����Tk���B�Ӗcr�*S}�vO<<��1�V��#����tߝ��+*�i;����E;�U����ҔK��T�^_\ 	����n]�t4�(AH��)G*-�Ѥ��ū8�����m&䭪NҞ�O^�8��X[�����;��X<����f���I )n�!i�R��0�c��W"Y�B@3��
�ʑҒ:�!j�HY�DQ�3?uD�i�q�#��J���a�U)��`���h(��j�$���f����ӒD�}C��d&���a��	"z�^�`�K�!(�<���q5���$��CmtJW�Z?L��2�炾Շp�|h�V��Te>�����*%�{�}�YIM�(�J,�:ny��z��1�j2(o
z>'YF��T>��8�J�<NC~�1��C��T3�DM�߄V��f���h/}j������rOp)���˚���~�����)*�.�v�h����pk�w�gl��$W@q���ڋ��b��'-1��x-��x3����!���w
�)�wC��,wڪ���A�� ��C���n�����0rI�����nߖ����Y_�����}��h.'��8���&ʓ��u�n�ڑ�Y��;��'IE�aR4>n��a��z(�4�/���<�ǫ&�����m��Y�;N��3?|������f��v��K����C1���sH�wt#�0�^�C-4C��$5��h1�j�.MY'M]�c��4>�+���Dļ"�i6�'9@�vH�zubfK�-n��I�ㆻ}=&<�py}iD�9F����?.��gb�C	G=�k���������#�`�w�Uq�KQ�9�S��&s;fl�\~6c*���Nፁ���$}/��]��p�>�Ѡ�d�aځ]3B�o�sP�ԼJ�Q^J�n�����m��̑>@���l���2�LlJ���d�K����5�>j�����	:��俈���7����"0��s�����yc��.X�7�P�b���͂��2~bQ-��=�&9�Ѽ;(Wj�3Sl�=���^^�]����C�ҥA&�Ud�o�+8��|�R�7#,�H��>��q�x���4�uub����N��$3WZ����* Z-����0��N�9!M@���H�-���K�A��X',���NT�W��B<N=�7EЏ��}݁��Ui ���:~�xu�a�:-އ��fvo�"ӣ���7=����T�j��auD8�]4��F$5�#(F��]`��9!�̷�?��ѿq��F�a(�xDhs)���d���d@<d0ݗ�I��[�)�J�E��e�@0�O��c�h��[ ���a�3B��F��3�A墈D��i��;�j�,D��;�HT�)!wE�r��4���"�'TtW��!Vl1ݵ��>�3����̓�Z�0+�,&tG/�k�_>%%�󅀑4�@	�% l{�`��KEh��������"�M����wi���'��4��йy�\U���bf�X��z����h���J�>�Ւ��d�H�I���l#�p8Sq{�32(F�h��i��%�8`D_"��ׅ�H��d�������33%!�&!�m����߱L4֥�6��IpOU�8�Γ���j�4+����&�%��=�kn���D��K?�I�	���Z���'4D�[���֗��\$��?�-����=7�ńt�|W�1e��߳{�O��'LD��Y���/�����Ö�s��f���B�.N*�Q;��o�+o$͜�#S!(ҙ�f��er�\����o���*0Z��o�+����0xA��X� `�B:�����Gk�rc"�f���4�R-Ze;ty�u�L%.��0�i- c}%�4����&�5P�^=���¥�����A�züw���2iuhy'-j
�s�W�Ai�wB��`�E# v@�)����`d
��A��$������+Y7��W���W��v]��BeQ��#��-D�䊻a$E(�$@K=��}��M�U���7����X�7z@��o�I-W$z��k��jb�k����k>�1%�\��;`7�(
�^��� �Z�yA�]�	ٌ1xO��cs@(G�O�*�-Ԝ�d�p'�(�[���;�鲫0�R�����������>��n�q��T�g��Yr�Aw�o~ͨ�����:O<W��-RP�Y)<F�o�Vi��-�~3� ��|�m̎����?�2��BX�v��L���cB�"�����I©�@�T��&�}�����ɀI��kdQ=��1#��X�U�p���Z?�H�C�^D��@{�CS�"�Ƽ�4���5�e�fT��\&��ZS�Z�ɲ�&��8{�޾.�Q�Ϯ{@ěg�]�o��:uu�TL�M�"�%���K�_�F�C��ذ�~�5��m�O�6�r�S�+{�H��҆�$�����_"Y�Ft	jt�xw�,[A�P�b�!Mh����p�,?���T_ґ�>=M��e�}�NۦѾ�6�F�S3ɂ�EE��v�eY�2�9���k�z��T �w��ns-[���{�/z�33h������Ƿ�hN�Q��g��o��_^4�"���M:���|ժ��j�w�M��8S���u2��Ք'�/䦑۽շo���e{{H��E ���q������R�GB�Q~��k�9��U�P��w ����پ�b����:C�) :�T������FHW�;#DXטT��fN��h��ǜ��
$�SS�/���g�����~�r�`ɮ��O M��9p����W��L�S�۾U.l��j��8�L��-�{ܴF�ÁPp��㔥�ߠ�o�Up������ȊE����68$nF�z�8��� ;V��\�<�3�����Bx���=�i���2)�6)�)�c@�f�8��MK8�/Q�c�(j\�jmR�0��%�RQ9b�0>���h}���~������F�|<��c8mFr"�b�u9%�o�5z����c����č���Rwm���~��-����m[;��,c��DW&<�L,jNJ��6�0�'=I����ߢ�s�8��.�*����'m��Og�㮉�s���2+�w�2�&X'Z�R8ê�LC�u�K^�KE�g~C���`��-t.�T<pe�Hr2�P��1���X�3���q�}-�ً�.Au�rO��:Q9�/,�A~/Ԝu _[����m��LmQ�s�<�+cv�E�Bb���t�W��zw�c�U�k�iuH�'��z���r�  �:~���!��j�DĒ�m�*�h�e܉���#�c_S�.f=i3/3�V�Q�
������N1vCΉ脬<t^�0��{FLΔ�z� ����4�k�n���_�)^٢f7�ே�L���C����kX���#_Z\J��F@ ���d���|ה��i�x|��IB�q�;�d�%~�P>�;����t�	��rw�'�& a��x��@ΓF���*JplP�k�v��D�T�ں�d�ˆ��Wz͕����*��1�w�j�:��U|��s(,���)�V�Gy���+��񻬦Z������~�ϼ㡓��:b,�wPq�u��_x
�w�&gA���CW3�U�;fwu���}���7-��ժiJfv0��l�S�9{1��[�9�9l��3�F	�a��x�8�M�[�ǿ��.L�9H��� ����N�����n� �s-�ߔ��$��S[�!�Ԟ���2e�ɨ�Hژ-O^V%����\�V�Y�`�+O��=�zpQ��ρ�:G�<N�U�x~ZP��1��Hy�o���M��SQ����㼉D�;W�Q�����Z�D�g���E������MzU�*����-��ju���h���:#a�	y׏%�KԶ���a��Ɔ�xBUͧ��		�S&gq�P�o�3��F��@���sK�R�e5�ѿ��L@ϙ����b0[El)~�+��f9��E�ŰlOm����lA[�K�1p9j��&�v�N�9�1]`v��bD���p��J�+m�"4Z1� F1���?v%�t-��,���p��0��K����<R�50���OU��-c���F�6�aLd+h�H0gȈ@K�o���:�o+b���4N��C���mu0�_���ٷb��G�^^��+���:��n�A$�h�w�l�K�FĤ��K�,\�W0�|"P� �l���q�D����(�/uh6��`n�O�vȧ��<�`�L��z ��|�A�k�6�����W�ɎC/���dAM��3Y�H�x���d\�+��t,7�F���m��0�nOn�{�;�y�5��0H���֟���;h�y�KB�jc{����q��x
�w߹��6gX���OkTk\�4��g��'�H�XO��*�#�_~���R����!.�$iA�$\��1�	j@���o}�NB��v�Y��r&��G���|�7���7��5���Ã���Fr)�%�#�H.�y\�BV0�n;N�^|Xzu�y�����'W��������µ���i�:�#潧���ya�	u���\y��y#1"�J>�c���$�t�U�Dy�l\{��򭝆m��p��@�U>���j�Whô������#��)��z�65#I�R�C�C� Z{�����s;m�?�Qz�1��̵_0%� ��UA��Iʾ��@z
��$:f���ã�^KL�1ﭿ9Q�Ģ̥����R��[1����@�ݰ1�2�:�����X�5Ƚu�=w�	&npu�;����|h�g������U�=���p�m5���dͼe���H2��e�E_�5�A�z���,�\��~��E���Uug���I����l�4-o��C��M���?IWt<ɔ��f�)\���?�@�!��{`ETK���C���z}I���B����4ďNkۛ��~��*G����s1jI�wY����5��-��y˳����V ��d���k	_9tW��t'��I�wm~�k�'N�MMӹ}W�|�n���"����vf�k=̌hf�f�u�>O�TR�5�5��"q�ޓN6���[N��ɄB�|�u
�w�<�&�\�{��,�*X�ޔH"�=K>�S�1��i���4CK���A�����B�L�A��+>d��A�Tt�tz�7���Y=�uC_]���ЋF��ἲ�P�G�nG"��,�!�WĽ޳�\0���kz�g}�oZƀ&应;1��'��7,����[�w�x'
�f��}���.��\�Q��N�����xR��-�/�R�J���9��Ż��Q��"��5���Ё�Oxd��s�03��nA��2Oc��(�Cl��Q��]�������*�~u��F'z�	�=/ٽO���6L?oA���"A��g���;�㻖�0EtA�W|���D�\g*���fA3������5��(?��4�<_��6Y�1y�e
�<I�?�g���(��	
�WL�&b��k���+\��jR$*�)}�C�� �n���~H;���U�M(�CR<�K۬��+e��Y
�9���kwc�m�{����|֐���<%YV9c,b�q���}�	F'V�s��&&���o#�ӖZ��Xtdئ�z�w�	�k�;`�g��Sm���655p�	����V�阻L��Ԉ���.$)߲�:�����%��ޓW���ix�c�H�JIW�_]�TE��z(�P=/k�����C�vf����S���j��?˗/�EU�J�h��J�&NE��W`I��l��P��� �z<����nB#��7PP�Ǔ.~���c�L0��;���F����] 1��ޜ����dr)[��ILqJ��E�/mֺ��y�P�.�^Y�l�`JQH^�8M��%_�����h���x�A�[��k!/��s�t�<K�6d��Yx��Q��<��W?Z
-�����~0�x���m���ӄ����O��2���HD�I`XE��U��8����n<|���(f`���=����\�T��`J9�9w�>h����X�x����Qh�ľ�X3G����>�Hj&Ix�t�6{$��+��-�9����V�<��|�R��1s�B������w��Z��DzJ�ǲ�ݨHS�3|͐��M�GhM���ف�F����[��!j�.�P��w�D��� �H�8eSy�\O�W���������TSaB6ܒW)4�ͭQ���a'r��9��P���d�A��m�T*ٹ^�f7�1��?.~�{��YC��BF�8f0��W|ű�D�LeA�=�}#&F$UJ&�ݎc��/��:���?�żxD�B\)ʦύ0	-0V���|(���9�A���7���Vۧ�>���Đ��;y��#"Y�B=�2�����0�C$�ݲ �����1b1�a˻lw�E~�cq��	C��#�Ƕ�7=�l8�9ĝɂo�8i���Z�LL��ƲY�8���J'Ѻ���#�@��`��5����s��(�G���w����r4.�.ˢ��	.ʄ[bp.zH|��{zX�'+�R^B�nڀ�3�if������b5�f�'���	�j"�E���dC5��:Z���i>���|���b����1I\[-���
�Ở5�	��"lC�jTG���-���Ni R��6�+�"JYCі����w�[4�-�.�j�/$mr'ɓ�]�<��`�b;7��3YY�3J �5V재�������uhJ��-���� pG��-ZM�e�7y����R�ݣL�l��Y�kYzO�Qr�/�_��@&�hl�����4��yn��UE����?��u�����V3�q��ֽX@E���Q�/�x���8�r��DޞB�oJ�@tn���-��:eaG��
����SUM��Bd$:��gz��ʭ����+���*÷�uu�����sڞu� �0S$z���T�
��sGȇOo�:��5���o��u��	�p��|��=��8̒�b����R�d��l�1�6u�.����-i.��P�GRX��Ɗ�cmWm��{��e(�[&$&�8��:�%<x��JJ#U�ƭ<�Щ5��R�@j�+�LP$�%jh�YE�k-z,A\��d��:@�n��k%�;�F�H>6�*��#~��0�:�M:u�ԕl�0���{f�&�e_߹�Mj���R��WG$��Or�9k8~G�݇v]��lB�sc����`�ɲbj��.����'�
}Pi'��y7���q��]5kJ���X%x���=A6����O%i�#����ZIV9Ҧ�y&�MPn}R�Df�&����	<P�	4��� ^@���N�8 ������{�6nB���c�r���]��)f�{*�����"��㔒c����s�d�U(���:O;2�2�ĕ��<VO�*�4o�/q�jg�٫�_<#����/��~��o�k�U�s��72�e�q/nG����@l?g�K�o
]s&�H��<�%$���ME�I@�[��#}��䖻�<G⍺�~Qt@8@�h����_��QBh��"��l(�aS�I_`��G9���n���%9b�#�|Q���N����E�����6�8�0�z�d��W�yw)V�cT�~��*cO��5g̴��B��-��y��&7�T�EV��o�+�߶�'?$YG�L���a.��2�f��%��� *��*m���׿*ORt�$��Q�G�ה�Jx����\�\!��B�<��|'�1�A������N���Z�3�˟��a*�b��O�ၪ��H�ʼ��*5jМ�5"���S�cyV%V����D�{,P��?�$NRB��Dxe��u{|�"��
�� ��m�u=9�E�XI*x&�֘cp��^�ξd�h����|�33�k�mxA�X�����{���B��A\BĐ�A*�{�j�/�)x�l.���M��X��������u�
���J/���e5��כt�ݦ�փnrn9N�g���)��n���<�uuz�$(=�Ũ�aJ���^����=5�E�9������k��<�K��p�`������8����6C�o���s��f"��)'���g8n<cOb���o �������	}Ud������0��9ߑ���9]�kͦY������YeW���V��G8�W�6�M��of�fDjU�������|u��8�A��5��o9�L4t����]�3�y!8'sz}�I���'����@�p'��'&��"UZ�>��6��َH���1cJk�q��"���ˣ��"�/��GUi���J�s��2/P~(W��OO,F��R��"� �ТȆ�����Ѐ�7�X��$[�9-3�_R$筀~g�i�'aCgM�N\w$�w}���0\d8��h0�b�n���kF7y��y���2s�m6��΂�zgg��mic&Ʈ��7^��F|K�%ꂿ98�;I�7��P5��m��J.<��Ӫp\���E\����|N!;�B�Q��+E$Ҟ��X��VJ��?��Cظ��J�:��c�{��º0j͹���p|��W��(tC߻>C�DNcqf�è6-9~�����9pҸ�OH�M����5�$+[%6`;��ܶw���a�GI��}��n��B��
�z�,�2�J:I;�=�o��V��u�{��3n�^ #r�^8�s��F�?�i�j��v���n¬=���oxP�+1��oiR�<�޴��S
o��> �E���q��lyyr�3�'S5��uy)�Ea�����S�����?ϝ7��'��m����s>��"��(�y��-����)[�f7V�	ï�L����d����lx(�?��W~�Q+�=���H�����u���(�U!��Kq���D8'�P��5����K&��$�{����h�P=�*�=��QtSm���9_�3�f%�/6�>�(�
��b�X�L)�9G����1���*xP�I��^�QZ8q`��+���7��ia��h5�!���c�84bTeu0V��վ6$��쉱bt��n?��5���.���14⎃3ma��j���Q��X�y�	��Z�4��z��h-��@'(�Q�}Y> �	!��Y���|"�]{���!��G��vL�cK[������� /Z%����PY��,�1�����>�8e�����H$j�o��%�<dr9�!F�:�y�ȸڷho̜����S�H�0#���,;��^Ә|��ّ�hB���ODI�w~.N�IPs�����^�P,�A�ec��U�)y�0�h�=F<�����.ML�@���5[t]�|����b�3H�}o�ݓ�Q�6P��90Í�yya/�~��	��\wY1���H�K�3�XE��R�Rbr�S����(~�If�W��M�%Ω�ÑmW��mR�7���~�<%�6�^]Ś��<�Zy���/�Gp>�6�` ��aVl03�Uz]oOL!<[�P�؜�2F:!�P��+�w��F�@������S�����[�1�a�V�1��mҧT�	�?�����YOL��
���P�υ»br����Qc��1ͦ�����l��6�J�O��Cy�����h
_�O	1�үAu�V�y��%n�I�]��l��W=�OS��Z��O<�e!��E�X�H_�%�'�%�I)�۪GETܟ�l�o|�����]����"�7�8����'^�M�٨�(�ǈ���F'��H@���)}�M�ꮨ�)�aL�s���tD4~"`�a��7�7�_b�q�t�>A��q�ɹ�G�Ze����H>esF�븁=i�X曦8�R$��R4��s�b�z{V�s!����bG�g//=�bp��͢l	�C/)Lp$�ה=����H�Ei+%{Y����K�F��|N�:{8B�GB��=����RO6�99e�āZ�����s�o^��Rg� �ClQTT	���8��-ek_Kw'�}j��Q.|��rs�k��uaQ��G�<�gQ��N!e� ���VM]-4!����Z�)���Uz�[��ۮ��Ħ�v{'xeՐmb!AO�ia��m}f�H_�
�놡/�,�1	F7�R�z~������]u��U��m�>��c����N�"b�����#��=Ki��!g]���9Ĭ#�Y�X�nx�³ �:oA�!�qLm����AG��گ�ƨ�����&����{9��9�ڮ�u��l�����ё6�?�[ު!C�%�r�A��3|P�6X]�Lf�r�����lsn��	�n[B�c�9���Ѕ��G�ѫ��'�~],�ks�D��53��� �H�r��\E�q9Z�{�Q��W�P3�xI���e_�O�w�)}�$��o�jz��Lp�F���>�Ҥf�?��2��!���	���b�TEZ���p��_�לr��h��DV
@;P3�|{�n�M⩁���=�M)⃗tF���ԅ(ysv1����6���/0
�^dDO9/,s����{0��=)���V
�L�K�G{�*�1x2�����܋{R/����OD��<$���' �&Qa�C{���f/�0�q:�Z�0]���ʡPۯD�:�\<�)X�Y���|�K��a��溗M6�3Qov3vx���1������O%��fA-H+����tg�%0�0�E3t
!^dE�ה�D��mS�3�� ���I8�U��~�5�`y6{�]���{B�'�\rl����|0bN,�m�׷�	���Xf�k��$�B��J3��ډ�@����#��l�F)�k�4y1;zmQ]�*3@��Mx,��B=��P(�����O��-���Jۓ�����'�=��n0a��-�yx=��I���a��A΁��������e�u������I���F�`^� ��C�Sl�D��R��~�4u�� `b?��	�ȗ�L�ו�k�����+!}��!t�2�@��V^k���0�T���S���_D|����;�^��5�7cj85�>R�v{UN��r������[P/nR^�#��I��v�_9
2T�j�Nf.�]ꡞ �s�5'k��֗���������9;�W�isY�{k�U]
��G9�e��4�w��B��>�jT�HR�S���99H�QB�ё�U%�v�4 ���l���1������n �5�=�m����t�y��� UD�;:t�;�d�!8����1�r8��Y�{�v&ٌ$Y��N�+&߹{��%�c��~�h������@&���5���z<l˭�+���ɻx��L3zuօw�_�%1X;y�ɫ��x��;~��	��h��U�qd˦���$o��i*� �+rU̯��+j�( �k}$��
��������v�(s�>F�܎"�����JטQ�j� ��K��r"0�ꄌ��Յ�7W�ż<���dՀ�n��q�a\��_C��_��Z;�D�g{o���w�@ԛ=�2r,97��i|�4��|h�(�tg���$7S��+�=�}rޕV����4# ��]ܔe�kb��%}���3_�~���hB��B,[䤍�L
��BF�n;9R��r5����r������K}Y�F���X�F��>̻���2�#Y�?q�(�F���b��V��e↎��k����� ��D��`�j�4:٥E��S���10o�]ޜQ��;qZ��О�?L�ؠRK�n��0ڗ�tQ�� �D��\�q�����[�'P�Dx:U{�&^F<{���~�0��]B�_Y���TsՔ�aU�g�����c��K�o;�]B�����՞%��>{}�g���!t<����WV[�5o� �����$'v����L�����]y��<v�n&���r%A��U�6�0�$
�ݻ-�t���km���]3�z`Q}埶d"d~	�x��PRqJ
�9=Z�A>�v=���]vFk�{Ɍ�X�WQ��*U6�~�5��Ӛ�0G�ҔxJPF2�p����S���y�T��I�W�eʹ�L���)�W#Ȫ�p��6q�r��+85@vN����84`M��v�q�4J����AEi>�U[司�M�E7�i�T�����_�?t��+t���\>9�HB�']P���\�~4���ku�JΧiZ��|g����J��~ѳ�ם�8+! 7��Q��NУ��7b]!t}��^�[�B��!+�::�Z���M��r^����ލ�K�4,�8�۱7����r�E�[�Կ�K��l��4ZС`;�#_@w�)y��*��!�"_+1 UM3 G�R� ��H[�0�ԎP}���*S���JХ]�k�2
6��H���J]uv�}o@~���4&�^}Enz*#9(�!���vQ+?���!,�~����`�����Y�q�T$Pǰ�C�K)���І�� �Nw�}�f*d���5S�6�\�vw2?�\������6P��~����H?h�_[�hT��!�Ӊ	�d��F��7�M���Ux�k�v q�KS6��*��4����L�Ɓ*�qЯ������##4�|a8	R6���E
��H��q��
e�t�S�-�MW�DS���FL����e��M�F�ô�^��UD�$H=6��#\ld�U#����z�6Y���E%-Ҙ��毐� �M�<E.�c5��J� ��&���k�U7�
�| �]}8��A� ۧ�ch�:�Iw0d2#�^[}c�{'S���}�t6Q*D��B�ښ�+C¨`Û�UШ����3�B7j�9�~.�J��%�|�� � f31u ���*�Խ�MK4�X�� ��W:�8��[c�����`(����0ʢj�)�3��W1�O����#�Ym��)�.������G<\q@e�D��Ojj�Օ��vu�iF���3�e�U�T�P�+ o��T�ڒ����7�mLtw�W¬��*yY�2��}����Ǡ��=�v�\���xÄ>���9��R������tF��ES�U�؋�V�� ��XMh:j�ٙ
��I���C��# U�K"��� �ۍ���`V*���4�}���4��8�(�t�yxRLW$tр)�T�Zq7�����M�S:�T�t�,��&�
�}m�������Bf�ϐ��hQ����9�	H�qޗ��΋�v�х�&�
��/���Rc���	w͉�J���)oa��
�Ċ�Kȩ<�/�}��SE,R%�`��'a�L�	0�/��20a����@C�ʛD�f���e��L;naa�m�n�-��[���i�����9���q�Ӝ�\�Q?�f�ơ�60ӽn�	��ߏ0}{��������z���m���&��p2��\��*�W	�U�{��f��eu�s���j�˖0fl��f� ��=o������^<~r�~�{����/��d[��{�md�fF���~�YCY�,ʖeo�o�u�؆��J�/|K�	{��6^��Kݒ�c��߉{�[�-���܈���ݧ�aFr�����$[�ۘ3���ܝ%�q%L%K$���a�<�[�/*1[(5PT4�%r�(�� N�m�/l`�imL��
�2�"�0���2*�ޡ΁`L�؁�F�7g۩f��(��� p� Rd�mqIM],P��v�i��X�@Ya��@7�Q�t�|5�Zΐ��0U�J@����"�sO�s�FA��)�0)%�i�~�rL6����[�T�@&���r�z���X�Y�7^.�!,��8%��{$�������"j�_|�͒:u�Х����pFv4r�XF���,��K
ɖR�/�ޤ<u|\�W��}�0VP���'@�0!�q0`W�*��d������.����ֵ��9�ᡍQ�T^����W�^��!��z���$�So�,�Vd�h��������F��6�o�[cA�(B�"�U��Y���;y�c]<V��[?gmlHÜ�UuO0i���%��GU��~�8�mkjD���������|�v��Y~KYOݹ��\k*��_�Q�g1�I�t&|��{v�ϗ�:���|U6|�u�%x3X��Y[�6��`e6�'j���J�IY~"o����j��i�s޿R��3�+��3����t� ��Ӣ܋-���t�C.3e�!�Ȍ�2u�g�ϵ�wp��)�0vy�K�&�T�o�J1�рD��^�(�#�
P�����KnW��~����/yzɌ�P�$WA���j�3� _,��*¯��`��%�]�㝟�|��O�y����Qf�����a�Q�ȷ`SN�a��5�ߟ�6_�[�~�7�W���h\���Du}EE0:��gŤ>�+��Cp6���=��<����a�!�Z�ߗkV~u?:�wb}� ��è��e�l���֎�u�.�	ǔ� �$�1x.���Z�%���u��8%�΂��,�r+��c�1�EL����Ve2��!�>���qO*d���)$��^ԕ���Dr���q�H��-��rm��$�Y.dKؒڲ�^���pI6�y��e`X04pj �+�%4��� �
 Ё��}�U^��SW��c����^Zv�%�d��@T^��`UXdO�g��f`,�Ѐ�Qh=��m�	Z��f@��:���`v�g`������JZ���ZS"���?R �z��B�ɶ�T��i6��0*l�����^��-��a�`�/��-�7=�� 6�X���]�r`G�+U/Q�Fh;TṦR���ʿ���Jv�v&�t��:�ym��S����PO�Zr�f+f����L��״I
?����W�u �n�(b��O�O?`��ªU+��`lA��#�;�ڨ׿��M��������		{�eB�n�S�8��u�<u���T��hoӨx���h����ͪ����6�f-��±Ҳ�:� 断׵��E��ʛ)T�5ہ`)��(�}�p�p_՝m�~M�jH/j�H �2j�'�sTeg=M����Z)��(��-P���]�ޗ���O�ū�k,TPUAÂ����J=�XB��vۧ�бФ%�~�j��;��π�L�P1����4�����u]�>��g���Ḩ�W��
@wgi���BV�=�҆Kp����X�Nxh&���	n�����V��F�xAx�JL��鿩i2��m�kH^��}���N��U��/]� �_��@����X����?E�a�P��1@����½��E�礡j*(��:m��ɀ���=����n�}��F�t �`NH��!4bD���U�Z�AX�Jا�������T����@l���]Qp�idi��wZg�؏$$�G����	���0i;�&D2����@"o�HY4���-�L}���@Sw@*5 >ѥVp���;y#~��[W	gЎ�\�m��o�khm��.���X�y���B�\�&���f'7ҫ��6�W�B���
�ꬶ�`�����?���#�l	��;�CQ�\�Z{_���=Dc�?=ٜt��͝�V�X�ءV�6�;�`M�Y�b���}'���p�ѫ�vA����j�CzJ�a�T>e���DR�5^�����J��E�8�BqOW=��x��Z�,�@*8�<lU�ig����,t&������f�����G�$y34�W]O���Q�k��sI��WI��A	E��?���)�h��G�z1���b� �N������5�t]�(��Y�5G��s��%�XO�
h�##�!1ߴ6iD�<h;�)�	֫{XBk��'��R��_ZL�5��X��?�����S)��KO��.�)q;Y[L�Z���/��.w��2�q�[����_>�·�o(���}��nv�R|�5KO-|I�>n���"g���V��r������g���5VWԣ~Λ����y/���p�U��|��*� ʁ(8͓[S&���P���_�-��A>u�aAҒF��e�n	��<��R3�z,�c�]�������b��,��2d#l;ɢ'�F!����%y;^E��y�<W�؏�;�gz �2U8F��=�*TG�KQ��J�en,�C/_�C���=�!�aⱞ�����Ro4�:*RGJ=��G��'�hApV���D������� �V:�꣺�ö���������A��Y.�ic�֩!���R��`��w����57;=�������w�Z�R�7s�~���
��9�30(-0zd�HJH� ᝗�� �-l�/ݫ�,��4<X-�����˳깖����ݝT���.��A` �C@#�G���%L�`��(�:�ql�)��$,�d,@/�{³��v�[Yz�	��4�vڿ�@�YpN��A��0�Y���5M�� �|g2�0w���x�p@ӛ|����S�r���k-<EkD����40���:�o[��y��e���� }җ|�3�X��z%U�O����I�zy����`T`�}��-
S��9��GC'��]�Byq7�c@p�໾79��q��8"_���Xԣ�FssK��=�Ȱ�v��5��!��5�	
�\�|a�$ZoW�v�DGy�T�X@p��S���]*��`1rn�r�%���κ�H�о�1�Ɉ־��CA�1^.������g������h'��������kJi�)�'���~(Kr���-.��o�-����RdG��S-�?d=q��~�Ul9�Ʃ����c��Qa�&�Ә��r�D)	�j&Ă�(�+p�V��o�2�^��݈�zEc:Q�c�_�T�n��B)$O�T�<.M>C}#�VEkN�l�:�Dfɗ���FJ�z;��̂�(Um�G<7f2=��[�n�|2�mXv��r�؄G@� ���+�e2֐����5ѥC�S�b
�-a��dFİ�^�1�}TS�u:T�1�<�y��h47��B����I��8���8'���@����0�ǹ%�+�)�$)>	������ٜc�qbNN�I��H�
Ђ@�A���KR���֢GD�[���
��C�z��+h�ڴ;��	�0K|m�����O�Žv���~�X�3�:M�uG_�m�w\�U:[�x���D��
��QD���蛕gЃ ��m7r,�&��*e�~�C_�r�8�	f
)GV�t0o�rUң�֝D�����?��N�Hw|�)��9����GK��r1��������>��l���)������^v�R�b�v�h�h�q��n�V��r|\�}W$����ռ^���-S�p=���ԺY +�#���2"3�=�h1��89.���k6I�hFBȤ�l��D��RS��R ?Z4>Aa�,*F"�~����*��}--�Qsw�:l���	��R���'�f�J���	�N���V�W7��S��)ӭ�
�t�D8������T{]�$!*�TB�@�o��5��U�z�at� �v�N]y��(�L�^?���l�;'���4ż�"�pW�L��?x�׼w�U�i�4�^o�h��gH���Q� "�᪊�7��٧�0�G.ͪ�XO�E�y_6ǹ�F-qWn7O���N��?g[�K��
I��}��� ������-�h���D<E(�8�kpP΄<G����c��.����
�t�"��7��/[Ϩ���xʼ^���-Tmp��e��c�����>z��X�[�G�z.�t��#=�4;�D��E����R�y��W��:ؿ�d<�;���L�:^�|H�1�c�S���l`�r1}_"ƫ�g�������5yc[O�`�w��S�E9A�4fl�~U�<k��whݲD Ak�>�}�4���}�UUJ�޾��J�u'��Z�Ӳ@��Q��s~k�=��yݬL_oޠ1�=+Yy��A�_��G-�'}N��';w��뮚�f��V�kJ�w�I�^4)gNZ����X��K�h3��k(@g���
9���ES���=�O����k�nY|�(��b�0j�ܟd�	�m�'ZrĶ:�r#�\bq{g�����
!�j�g9��i?Ҋ�}��ʢw���c�� ��I9�t9y�B���	�c�����C��d�!N*��ə�7B.��b�H�D��P�x^jSGEn[�����?���d/�5��F?_Y ř��B������']o�#�r�"W�Dǁ�!@�#�]�K/;���[��Rq+�R�31b'�L�!P�Y�/�o��I���g�n"3��w���N.��ܬ����l�>��η��=Е]ȟ�BN���w�S�x�&���9:o�6�瑅�H�i�:Mɠ�C�!��GS�A�'/P��cʑJ�/(��uA�ԀJM������P)2d=i!YvZ�AVd:3=�_�w��(��vƿ����z���&��;c���ePC�0hu��P��Qγ� 
;����S���������׌�#�wY���R ��BK\����䖎҆��p�Po��z�á���ӑ�+z�?�˩���+t$�ߘ�tO��3cJc]u_L�EH��ͨE��/��y�SC��ɮ���U���YD@�l2���I.0��l�P@���EdT4F^׊GO�(^1�P�MJ��&�$?��_�$B(ALU�OԒVދ�gK�*A~��[Gv<��Q�\�g�w%.�t/�\T��q�
���>B����7"4�D���Z�{8,��`rY��]�����@����Wˊ򄥌W57n尋�)�4x~M����~���.A������z���:^z�E1X*��0>K�v۵��k�S�Y}Wj������;V������������4��e~���VX �� ���	�ܵ���J�������`؊�?���M\D9 ����p�|o,��@+xUi���8��X(���ƕ�L��Q$�����T���2���8-Q�FZ�g͓�� 3�A����)&��"�X�*�
���w\,��b%��
:׏�Q���ӣ�m[�~*�g������dF���"=���P��W>]���!5q��;{��us�Os�� ��PƩ�h_q����@*�x&U.��-X6k���D�x%�MVkBs�2���o�ˤMF֊o��g�6��S̞��W�ƀ��1�/o�^2|�TT	����';�/m;�@�T*(N5ʉ�9
(eD0�/��z_~[�s�R<�&�����Ў��0;���̅Wd,S�k[*�1�c� �t2ha$!�;P�ϫ�G��!C��Uqak���j�V�@v�5G?���u��V��ĵ�8��[��Q��Ҷ�����|�I�I�v�<��{��gQ�2��3�Ns�N�dʽ[ʠ(��?։I��'T]��XI���UXf��\�ߓ�����j�-i��R+Q�����~�%6��]��k��#{͕�,�9�����s�����Mہ����A�Υl�3�\��[sZ�lN���0/�,.�5]�*��Ѫ��Io�_��Av�C\�oZ��}��"��%�G�QpOzQ�T��Ϛ��3/��\C���-�5��c�jȈ��i)i����+��@<� ���%Z�Ȱ�_ѺHԢܑO���w/D���X�@^mZ� .6"��q>��W�J�xT��.�Q��ج6"vjӯ��rn	��\�ud�=��K�F�x&�#�� ��+��[�=�J*-��KH��<@HRס�T��y&%M��g[�S�* ��\d$�/	��M?�6F��Ap�؏�R�k���M0�+8�(R��Fe�/����>"2ۥ�{	G3O�O%������
ӥɻy��yQ߬���|�)�:�]�o[_���<�;{�|�N�?e{a�z�<���ꉽ-�`2����8-Tu�% �1Gǻa���!�+;R%ˊ��U؇8�����aVk���T�><����}y� \�9���C��ӾZ[��c�:P���@(�?<X�`� (EGh<�_�/������l�z��B}�IѠq�<v�뺀�N�v^7�X�@���p��ְ�q"Ӓ��ʏ�\�4��ʒ4��&���#�B��(����&?�D�
��-�B��+j
���&06@�����j7��Y0��������ۚ���}�v-�i~���곢l��+�f��e�Fт���R�︿��}������#��Mk�&sd,�	��"b�Yǆ�	j�ÚAPESV�DM��K�	c��{<,K�dO��~0?'�Ы�+�Br�#@�z^ǀ��W�7sb͂U�F䛉}&=�ѳ�9,Ds���0:�A���T(��|.�%��Hk�-��Jz�vdH�-�r][�f���_ߌ�?iK�c����������Y�Êe�+�+&��y�� c�R���*�YU�,j�3?�{�NIf�O�َ�t��v�r�1Q��l�LO^�(*�ٻ���t�M4������H��b����h+
�Ѥ��Z���d�M���{S��M����Zz�"����%��-n�^jr�N6L�N7�PZp	U�&W$�����`���Z���8U��n`l='��۹�����xlB��A�N��3|��\�����/I{J�MD/��6Bi�����?D�+3mɩS�Y��R@�-��;�=�D<]L[��I�nl)u4
��O�}jA�.���RY��Iy+���3c�܂L�J��y��o��!��y'κ���5 �"Z�0����ޞA���s�~S|�	��:��KKtV������swȠ��|��72ie]���1��mQ)���'p;���Z ��	q�<~��L&P��+���^�n�?�f.�0�R��~���;��3��<e3�P׊������'VC10�)���@��.d�t_o1�6�~��2[���V뼑%�6Y9�������8m���~~b~tl�ԅ4�}9���0Y�&C�����f�x\�A�o�#C]��HvMӶ2����J6g\��Bsanaƴf���� =�M���=�J� 	x�PE2CС�~��	�i�TC�~��qa@�4 ��LP1���c����k�$U�P��?|��e/wպp�te{�-X��f�@2��)�EBK�pX����Ǽn(>�ҷj�@C2�¨�:6<��l ������Zz.���+�/}w�bƑ�hNU�^?2����ͥ!�iF@)D�CT�P�X�P���\d5��e�o�T0�?6|�t:Rg�_m�_*+�K!��[q��	�gc��������M\��t��ׅ��M|��0���(T���y����D�#٭��oiv��y�]��X�&M�嬄k���G~�^���:�ک�AN(��j�
a�S��m�?`;�j:2����l��y���h�k�X��w�~���f�[2^b�q��s�v�ۉ?��@]��^I����֯��h���0��]��yH>~��	�ЅsvxQD1W~rx�o�ڨ����/�q��<��*"-~f$�"#�̄�S)«2Z�M��.��'��j�i��(7c~�	2d:0�ʘֆ��������"6f+$Zkb�A1�&�~&	����Fm]b�fz�^���vC<��>^���x���bS�!Ig�E����F�=f�Z�=�ɒ��H��3�Ooo��+U�oܴ�l�tmZ��S�}�]�¶-|7�@(��Ό1{ʭ$��,���r�7.���:�>�J��\H����:�������)� Y+L�G����ꇛ�@'���e����r�5��"i�ސ��
�وH�_�OF����A]s4Zo����Z���$5L�q_#��*��ѐg����2�,�� ")��~4j�%����W�ѡ����;��	��3ۮj�d`G�U�OA8K3p�m���[��(���Uq���
2�j>l'�ݡ�n�6�^�l`�q뜺0C�-N���m�n�Αx���읢�?:`��l��?1�(��Z��U��!���m�3�.��MF�� p7Oh�/q}��
R��a0��Icc�e��'�6
�T�,G9�����ZZ�qV��5�_���p-i��<f$_-�����<z�
x��T���ZL�+�u|?=�0�D�@$ˎp�JŎ�Ǿ�b�*��2�\���<�J�O�:z]hY�2���F�7��7�勈=� o�eI?
��%`5K��5p���в��_�*�B�SA��� ����ݸ��$.�C��oI|��"����π�Xץ��P��+tŞ�5����~���g�$�6�z�,�!cm���up�)a��1���w*ŵ%�������f<Ɍ!L��Ɋv[�ީη1`@���_\-o�O>�8TQ��pͥ Y����5�M��A���zl��3��n�� ����)ǅఈ@�X�D�4��ݗXF�� �����O%��+�jQ�R�ˉ�F>�Y!�����AE/���*X_;����Wnv�M׺i�>����.A���	��M��Cg�G�?�����ʯ���Q�<U(C�q�C]�}��$�5��8�ċ[z`g�誛�=`�k;f��&t�<���G�:Mg"f�{�M�h��?S�?p>��FI^{�;����B���#��v�m��=Y7�@��j�3��NE�ߞi^|(>�x�������3��;��VH��������\�hl�9���*ס	z��W�p|��Z����'������N��9�+u��N��s������(�=��&1CΠ�ԅ�;�� �dE�\	����ֻYx7�J����S�Ċ�s���I?P0)���a�V�	ŕ
��}���7���O�J����]y~]E��V�򖇥հq������ؑ������J���c��ꪁC�d����d<^�Ͼ���@8`�t�

wrc�l��?I��P�㓑t���ດ
�&!f{>���|;���4�4�
���d	������������L�j�\�-u)1�?�C�L�^ ��� >��JE�3}n�����9h�^ ��^�,��m/��*�LD���t[�E̎]Q�ȥ��'%_�v������t�� y��RzM;z�̭w�nekb�k��֝���l3�^=�WvZg�����>)��W^5�>���<硉y����p��T-�&��-�U�!l�����rͿ-�xz+�dtf���A�:�b���6�l�s[|�!��⬞,?�b�gj0���Y����X�W��5�;CԎ���9���b����M��4�ڌ+m^ z��c�!~r�YR.����,U�IL�����LuM�؄k �Ȣq���������2f�n�7)F驯S؂�� �t[\'r�_hGK]�-�j��՟����[���݆�P��H�S_A�6J���C�6Ԣ����vl��=E�^�Z�9@M�Ԯ�ׅ�W;�7�C�t@w�1��ݠ���H�Q��q��	|�W$0��='��N�aPo������4�0��~���Chz�הD��-�c�R&ȶ��w���'*����?�fb������j*W��1�>��	���_a�ی��[��E���J��gI�/woU�x��m�M��ͯ�H��ml3l�3����JQA��zOr����J��;����|�V���
0����<;x�4�zM�b� ���Z>
ߜ�ᣈb�˻j��H��E?_�@���p�2v��.
()pZ�`�BN���à���s�"���ǘEp�c/�υ�o�sފ2�,�{�����b�����C�l@'�a{��Y=I�l�u��"&
�����Q�CвȬ�C�?k��C=����b�r��R��E���ș�܁̿�y�.ȡ�!K���$�� /d�ÉD�� �V@� �Z���48�,U%��Ɇ������}�7ɜ������zw�$xA�y^!�>4��8-�W7��;'����%��I��d�da�Ia��� -�U���\��G�z�~�weCӫ`F-�����Χ{���\��}~�>6}r��~�V�P�*�&�N��iJ �X��==��-[��r�d���� !k��xO(�|��b׾ߥ	y+��aS�1����#N��:����Ұ�-�,*^r'�����">��ea��h6�����PzGn#��I��4 '3���b3��C��9�UxXnw�0h�y ���b���:	�d��\��+1�=�ܷ�_fl��z6�����1n<Vo!1���>-�'?�2dE��{��&=�z!A��B�D��o���5�I���Q�&g�3&����Ƭ�[+c]M�VhAD�Zks����s'���ѐӀ̊䬑�3G;�_$�ߜ�c�,��2͈^�2�Kt����.q�'���0U�6 7�!�|�y�ф��n�v-�B9�#�>>1z+��_H� ��z>D{$�`��\Lx�M��ѝ*��� y_���(* _	0\�$��ՂJ��y�-��I�E����4 �/��nP��J	(W`�� '���~�m�eN���6uI�����`�u��^GSJK)`T��ed�����P^xÍy��A %wlf�)\�)�C�Q	rK2	����(5r��T���*�P���|��g�6����^6(r,�(b����^o��JL�S;�=��岻/^]�X��A�_,����v�͙�{�xI2|`4�;��Zw�r=�o�۪I�:;	�^���S�\�����&<�@|WM'>�NR��v�'0�c��~�<i����/��
�?i듎�E���8,�I�B��!N�,7H��B(q����
d� ֍!;���z��f�z%r��]R���;Li�7�۸4`9NVv�w�	f������'&��Y��\�},��A���h�z�����э`�}� ?����nnX�m|xd�HX��GV�6=&�����g�sԐ��Qp��Q�*��:��0��S>��/���F���rȦ��,"yuI�4�u�¿�:(�1��T���y����FA�L=ՍL4��(�jz݂��
n���$]o#>��v[´r�+�U0$
ʃL��om��C��l�$޸� �ߔO�z��	m�{	�V��r�/ә�vtk��Ǣ��<�.�*�{R-�@��V+[Hvq��!�z�=(M�#oբ���r�-���Cm��� �*��v�my���K^I�����Z(��ǱZ����,y g�
A$��!4�h��-�����v:K���d�}��ʹVPa�{������TA˵�PE�3�ɽxl��oT�����}4	�TB�X{�W�y�Oxf9IRW�p��]�#^Q���ɷ�:���ݤOq���������b^�q1��{�������/��<�y��DiE��l�bƊq$/�X����\��I���
����[ǘ?&Dm�]���#�{��}tS0�!]�X
�̧2J "
yh ��Q����hԚuW"}º5��ܜBIR��b���f�!��:��c�>.ꥱ1���h�N�k����b�Bi��z��Ԃ��9�
Q���`vmi�`��1h��͙*�FJ�lp5�$�4 Ԗ���u�@������(s,a��{�CgC��'�+"���T.��@0L��*ej���(���8���e�Nx78�tă|o�'�d��g�3�#�Q)�3�y)�
4j�;�'�>�
��W�W)v\E7��㒨q��R�bx?�Р:AA��p�g��_B*.�I����U|qsef���4��O�绔��=z��ze'T�����!�(A��-�Ӓ�����S���E������x�F��m8)(]Ґ����I�PP��%�gX�U��0�s.ȯ�OK]5'`���;�&� �|�=��	��a��X���������ٵ��N�@�$���r�o��|ͭvߒ�6����4�J��ק��I���N�'�me$J=S\<��u�����1A��h�+vFpC���l�*����_����\t%�3���z<�I(P�d�X�W������Oy��� ��o��j"�Ӷ���+���.���e��}�f�օ]���S�X�=G��D�J�0�d�/B���,!49��E�C&��Azf%�P.f��7�a4[�C�eՆ�cR��V����H%��җ�0(�k�)��"��G�Pf���7�Ɍ����@�`
�l�h���#lK�ԛ��䌰oq#+��3�������V;�֒U������RG�ϯ��\�w�J��H��)�j����J�č�DJ����d�5�T`�]߂%TZ��v:�V�ϭa��7O4�1�^�{4�c�����%��* 0s�O��a����(3h �1癥E��9��£��Ix9����fr
U����X�(���e�0`����.��p�jI^�Q0b��P����"�#�B
*���S��W'7<��T�Z*[*�p
OD���\���W���	9�mk��d�ʹ�if�]��Yi>uM��̆�!�7����9�)�@jT�܆����-��(!ܬ����h487�w����o�$Arh3d�����7�{UnmZ�1�M��vUؾ��?�ߞ��j�-۾�� �{�]���������Ng��b3`����v
�m��[�so|����d�h;HlsT�3�%�����U��k#�ں@Ѓ�X�iL�x&!*������Ҵ~��}�v���|8jPM�1p����U���E�F궲��U�꽚%������i���f��27�N�g_��I�غ=���D4�e��?�N��Tx�9��)��oa�)Gh�g�`s���#�2^6���mJr�#���W�����}n�P��8�:r�`˦�c0������0���a���<�*�!�w��	�P�^��;�b�V�U�ic��I��ݭ��Of�j(�X	�C�V�0=��o�>�2�U���"���!T�6�Fa_��r����+f��$F2�E�~��"�WFnd�:�=��d��(t��;�0��;�����L����UHɹ�����Ym&�BU0�U�!�2�L	S��3Wk��0�j�o��՞d"f!ؙ�f�҂��6	�4�09f��o�6��0�����i�8ZL1���s��{��l�9��Tղ� �����8� ���u��׿��:���7���)� *�h_��c�rQ �\AT��ؠ��$�ʻ�	��`L�0Ȍ�]���x#���`�c�����,���/�P��0�X��n�]1L����������kZt�7�s�Ս�![�J�	�/��
en��vݺ����K�**��*� ��ۗ���#��e��}w	3A"?WVx�?�ґ4x�'`XO&�{Z$`���>�|���Ȼ=J~ ��Z]ZSr����>ȩ��؞�{�����N 8�%��i�} ���Z��0�C0��=�"�u���#�x,�6�:�q��h�>�Z�7��?Ø��������G�Q0�N�r?3�Ǣ�p0��s�� �̗�qOZO�S���	��Z\�vp8�yG�)�����3�[��kU�X\^jG�T)ǿ�	�qD��%PJy���\�9�c."����A��ll��k12�@s�͡�D��Q��)��y�x��JoIV�65��I��,�T�`����XI�F%��'���Rm�q�{� ��݌{�����c�-�/[ăX~M'�}�*�K�7��?_��F7����5�N���D��AB��v_�s���E�5O�_L%�{�f[9��Y�Zϡ�)�����b⢭&���Y�?8���2�3�%A����2����|iLH�?5�7|<�
�5�zG�N`#v�����w�^�]��H��1=��G4�|�Sɜw���g��hD�V��QH �oƓ��;�Y���)��h��0�!�R�D��$�:��P9S�����IO����ѕ!��I9I��SEOQ�l�tN�h��vƺm�B�Ƀ�%�,*ٶ���P`<3,��*�ׁ�^�U��I	�"r=��8)�n�����=gAsd��ڵ\���4�A;�~��´�V�*�s#�m�j~���'�+i��b
�Z��|�n.xJ��)왚mHa�[�H ׷�0|��]g���I(������#�%�s1+��#8 �;<�㨞u`l�N��t�9��p�u�۠�礝���!V�R'Z/Ɠ-�I��+�l���8ò��� ��l0�,rx�9�ENK�@t�'�I �(]*��B$b&�L�$%���2���uX���.W�3ư�u�"R����SE����Y�7�<W V>:�(�
���-��l�gJ��t�m1?.>�S%�K~#5��� ��K�������+�>��w�&G<U��#�����B'���r-z8�o�h%�1�Agwvj��N�n�g-7�kg�6%,���ܢL>��1�h�ى}�j�����'��7jT.��\1�~��'Qܥdm�߫{�Ү&�*�4����ed~u���w�$�̐%X5�֍B�:��=)�h�4&2�}�=YS4d-W���ۤ^m�Z*8v��&�u&���ƐM�帙`i 4�Έ�A�-��W������{U��	_���-�~�<[�F%ZFK��ˍLg�S	b^�N�S��h�?�s��4/���"<�Cu�|��E����0C(�xUtE�OS��J�`�7"�(I�;�J@<���g�8b	�nI�������ApJk&:'H�%���;#�)���+���T=��	4t�_C{B�OD������kT�3��}�m��6�M��i t�!E��	��,<��M�~h@z�ӹ�=`���9ݻ��N+��+i�=}�����Ɗ�������F��C���@�;S[l[�F���z�-(]-�0G7΢��q������)�k���7%�u���_���2�%���[�~T����Y�6�J\����j�2�;���A �8]��EԹ��R��sa�0������ ��_�W��@b�o/�ŏ��E2�0c�M	˝�?��4 �����Y�;+�D�g`�6�@l�ټl�O��)�ց�����}DT7M���߼Z�,,qfC����.���D=�|����.�h�����,��j��	�G�ej��Q)�����s `�����6�@�wf�E���+<v4�]f8��qev�!�:�L��ү��џ)��ھ P���>w�b�u��@��L/U�iE\'	C��P|���c�s�����_�j�_�lU����7�/+��P�˱}��4mT��_c)�Qd�c�#�Qz��Q�H��J��>?��������G��fy_���N�)�Ϸ44��&M�sw}u����Ȩ���D���(x�����|�m"O�	Z�=BU��Y2�M[IT��ټ�����U��}����P.�.Z]��v����G4sƭVu6���$��rhOSY8b�(ҹ�slC� ��-�s�M������&���)N^)��=�iXA��Q��;e<<p�H`��{{���pl�[x|�[�]��W#Si;Rх��rA�S�w���������Dg$�_���'i�lN��Η�{:Cӽ�c���#*Gl N���a��5<���s��(�$�
w�b���	0��b]D좚�E����/W�G�ӱ�|�S.�0�X��\?�>�g2�|�ӫ_��5դ�\�e����2nc
���`��<ˁ�`r��-����ߪ��.t�[���l�6�G0U��n��@ ��[x:����^3�AEn�L�+�8>�I���F�sW� ��7�fjΘ�ϛv�8a���<GeP<�	Q�{����d���m��~�~�0Z��˾MR�^˴�y�(N��Zv*Y�V�q�rM����x�5�UsfK��-��%S��j&�z&�xZ�+�ܶt�����B<�<Fa��Z�N�rƥ���ߐ^��C�0�+�[��3.��z��w/������`:N���3y�C�h�c19����Z�q����o����f���4{]D��87���'�15�ZR�r�����\��P�cƗɱ�2]u$2��t�J�"'���b����L���1�����Yb{Ά�bJb��A��� ;�<x]�
�d���t"��37'����� %����Pv�1��-�^z{u���mђV��E��?��h)��!��8?|i�st��$��F�"��.)Z)e�T��\c���9Sa:�7+�0�F��0VH�sC���ޤRύ�.������jn\F[�[��!/�h��h%lÉ������C�@�]+��6�&� Q�=�W�b_<AQ�a��a�t�7|�$��-�� ��g(�Kr�}��)h$��P"�թ
{�����؝p�F�#s|�vqqV�qy��,�s\F�U���;���3���yp����ញ����z��{a����>V�x��V\�,8u Xff  7�S����u�T7ڔȏbӞҲ��%V���Ua���}>#g���ߩ#�Յ��of��d���W�1B�zE�&1]`��ϺeH�Wc�4��T�?U��B<��c��QN7�H����4�����Ǽ��_�̎K������a�<��m��pM�0�x�`�m�0:.�f̋i��]i[���^�+��[�kTm���{$S�7���oD�r��`|[c�8�.�lۃf�C�;��+��{�,��*ܛ���%�����|qè#�<��$h�+���.BW4���Ι��
���;'%H��Ÿ���$pկܾ�Y#��繍x(�gL��K� �!�eO����<3�Q��g�9��,�2�Ӹ�Oȋ#�j���!�W��*������BZ�3Ϙ���6�f:�y~���/����,����O��Iec �+Nc*z�؎��|�;�b/qT�;������J�#z2�^�S�щ�-X��N�]�x�F;N�<Õ`��ߔ� YR�_X!Q ~* vw#��u��C=�h�D7�<����thZ�}i��j��Q�������+b��<�)HiҾ
�����	ia(��q}5�Mx�<x9n:@K_h�IڛC2�k�t\={<��js%ijѿ3��y��D�*�;P�؞��:��<���2��r�E�n7�8�-@*:�j#�bo%�@;>�ld>9]1�P`��	J��g��KCS`[P�HE@`��3��.U���a�;�` ����ޣVDm�Kd#fƾ]�o^��AE�k �F0̘�<X�uږ?��A��"���FC�d�۠�u�w�}��A��5�L��*h�z#S�e���pdD}i�
�C��Y<ֱ�a`nZ6���m�npկ���Uy�Z>����p���K�GQ���l�Ȫ�@C��k��ܓ�,�����,G#�{ƈ�e9]�؋v�CI����_�@�)��o:�u>XP3�E��C�0}��Lv󼲓�u���1=�"f$�8A�0��Q��O�S�6��[�ӠB̯���
ֻ��uq�QR4�E���Gs��{�-���ѭ�L��0�:�o���#]�[܄1`����1?w�l��}��~eL�'�L�k��|��w�m��1D�]ڙ�MD5p_VD�r����j	̀,����$��8�t�D��i�a��%�}Ȃ��0��h^�90��%��}}�7l���\Y!��ϙ(�C�P|�n�i�;U��%�p��)vV��>��D����/�	a�Z|���]�"j{�����q�5a��1���x�AU�OD��uK�`81J���'�;�U���/���׊e�4%st6� �J)�bʃ����6Ł}��/e$G1"�'�
�y�����} ��9�=d�ɥ�E�Fr��=���{VD�5�}�F{u��0�p-o���,��A]��yzJ_L��Gy|�.� ��>�)���ਏ�����JǦ���w}1���v��Q"p����A	�ćl��Q������Äd�xt����Z��I�6�~�Ef�����;���&�� ���yM���Y&�L�OO��Z#�͝.ly}�e��z�533j0��NV�t���c��?��;�8yHM�p���L�s�����u�{���R�����0�z����d�'Z84���{��b��a��:��Ka�uF�����'��m�	pD�L���߉�q��yɓ@V�Y��ǳ<��Z��;x�-�E�B�p��L�L�e1\�g��A�9f}��,M@�̧�&"�[{SpbpL'#�?K��^���J�+a:�e�*B��2+�#X��d�2�*ܷUm�4�g��)|C����+�ЇNŜڶ�M�|����?���˄�7&�9��IHh�W	�.�}O4�1�%���l�c�CѢ.=�ӚgWm;$��{K�Gt������(��7���e��<hlܞ�+c���3`e�4���U���L!�_�2%M^1Q�5�b�.t��e��l���pT|p@
|q8Äϸ��.r}20H��M�|.q�mT�}���]�f�k{�͏��҂������}�(۲�����GL������Ӻc֠�ӛ�C�y�s�8�W#�9��<yޮ�i�)Z�+��b��cjr��f]�x���$f]��&��Z^�q��N�0��ds��_����Zw��f��\"l�����$T���;q���H�P��K�]c]�2�$V���gT�,.1���Y�fy��������r�7t5Ds�IKl��y���V	!f�(�>�Ѐ(Ћ�>�Õ�Y�6W����c�W2/a7�o&ܰ�#�+Q��g�<��aDA����Y��S蔘�2O�|�i��"��6��T�àV�����^�G~`�ă��[�u��gO����Z/��\4�F_}�������utX-�I�R��cG��,P)E���pc�����ҭ}p��zQ�b˅&v�g�
�% �����N2�Ś�),�N]IVvE�
��g�%qV�����]���̛�t[�n v�o���$8��si|EM7tH��G��wP�X��l^@|Ül��e�����9���0� �H�P��O��^�Ϩ6=��U��T��L|zǉD��c������4W��#��?�Í�0qʹ�Y/KfZ2	���ЃF��M'M��%��TA$��0T�!P���[؂Пp(��f��L�ol5�Et�e�$��נvY;a��N �*[b�%��́�?G��7����/5���N��Z�E�E@t�zO֤��GԆ1����Á-Ŵ��и�6\콵�K��E����T` ��>�j���0�Fw#��� =xs����#Ȫ��68�"JT%%	\A\,8
�p,��T�_G��v9�b�q�D?�.o� ��;Y�}����8�݇o>*���Y�y�FJ���Xh{�V��(�ݹe���r�A���5�~/<�#���`QQ�6���
�%~�Ɩݬ2/�`��{P�N���.wfP�-����_���=���1�4�v+�@U��	m?	%$��Ki�X(::��1�e�H��N=���^�D*�珈 ����1"��0I50� �G����ù�"]���ӌ�	�a�_@$�#%K�]L��cK��+#�����C
�����bj���v�8��*��%qIL�T��/aH��T����b�2�ԛ��T�(���a�c���=�L<0-��&�ШE�6]�*8�E:A�<�_|���4�ؓ��R�Z�^�1�/���/�N���{t�õU��KP��H�D������Tg�9�v���z��S�:Kv"3�{���c�U汇u ��ꭻ�t6\;�8�ފ�F��k��`�;���gTɪ*Y<`��Hi#�1�8`#��gP�ٿZ�C3 ������6���!a�)_Y�K�(:�H���>8���uv����1�ц~�t�i�ɘ���(��1�Y� чfȈ��F�&湉���k�A
d+?Θg�^�����
��.;��<�ok`���J�L3���`���S�Ɓ�X��g!(0|���K�g�5�`˾��P��R�`�[X��$��$ya�SC/C�}�7�QQA� ��1�0��!�ƛ奔!�{�^-*����$`�����g/l]���qUw��f��n DG�>�����Q������ډS\����)8��ZW�	����a���7�#���㟮+��z��tL��gT/ʿD�z�Ϩ⇯, �F����	0�4N]���_�>1�֞�����k��Ap�kq���>�eZ/jM�3�q��]HĖzN��ڸ1�	�q���6P���A�|�}��.w��l+7~�IɁ��'y���*�z��?+vJ7"R���P�qvj�>$�����1�H���V^vM)���;p���)��`t|�Ҹu��F̫N�-�W�n|7�5�A4��SٳN��l�0�����m�[]-ݺ�uM3g>�:��f��4q.v8e�7�_ʍV�ْgi�J�ix���d͒;�=�L�#(���g��mm��XVd�ڗ��ʰZE���a��n��Ҙ�Cn*f�(�^]�}I�����t0�#tr����D��ٱ����|b��cڕ4�A!v��7�UT��T{O?���t�y�|�(S�{��n��35��'���␼s6�Ba��ϝg�M��*&Ґ!J�?
ViG�X����
� d�0'��X�$��t�W�d�A�!�F�ta}��k��Lq,�y.��w����c�V�g='jV�y��j�����.y�؈jb�ߞ��j�K�����yW�T;7@\�^%�χE%m�!?�i�	9��<T���?I��-y��o�[Y��|bH��]�Q��s�-LΪZf�I7l� ����������)��uxpZ�F����6dy�p�e T��[�n�4�/f�c� �,����#(������D�0 ���Z�㚭~w'~�Dz�rk�䰳�o�K�a�L�8b��ò��ݡ�t���+͖��ma~�#�+�C��A�f��1P\~�͉:�E�~j�/2]ä�+��cg��n��WPbJZ�ԡ�<[��z��W�H�z�B��Z�?����Zc{�/� >���%��Y��b0�1�������/������	sO������V�1x�Il-�C��H�
���`��\�S��u�B�#�[>�ӂGdχ'S�.OķY�v2f���� ������4���k,q���.��>7�@���8�	�盪�{k�H�'��Du�J:`��E�fSE���Q�s�����(��� �t����{y�q��1Vށ ��8�`;����(��ȱ�qڡ�f�J�M@��Lx�#$EA:�S�cK�z9����c���B���e��A;K�$��7b����1]�	��cR�rB�O���:c�-ofjA� ���?,��`#��Aa�U�zm=�6��m�tΊP�&�F����>}	� �I?��aqJ�B�]���G�S'*��2ߚ1L`�B�ŁJKſ!��L*!���B4D�FA<g�=�^��I(�)e1�~�n��,�HJ7��^�y������՜�P'��3�A^+��v� �.:[�(ӑ+f�rL� �՗TH8�<�|�05 �����eFFƣg�ZA6Q�9r�c���U�a�)l�k�VxNӔ��'�o�l0��55�J�⬣~D�-#4�D_X�� �[�;�!$_�L�Z^�}pi2^˷��iGI���Sƚ���Er*0��%<&�JxI@	�5h������M8Y-���7�9�7�����B4ȸuE&���x8�"���)Y�é�P��t�u��u���G]t Wc��ju���P@PR�?��LZ�j\�4�Hj����@P@P@Qewe)�xOtN*5��&�B�5u@+�e@��+ZW1�3�Gj8����n7����]#�L @�9]q��}��h�$��R�.��rS�
M�sk�2.��Kx�Q�k>hP�o2�=��B�&�j���f�9�2˹dkU��ͪX�k����^��_ >�|>�UUu���6�M���� �P�h�^E$�Y��FLPO�-����X��Ԟ2:�0��I�c�d�(�-��"(�����!sL�J�N���E=��;d�	c�P����(����ºa(V�#y:��}֚��q;�(��J���w�䆁���Գ�ǀ�-��qbS��¿Ĺ�������)+g,:Kx�W���m�΍?o���������9t��&w���YT������7u�Hr���Q���q��8z�py���d�y����&�SQ�yu�w��o����>��
����c6�*��
��5�w��v@�P\^$3�M6�7�o�i�ۇ���ˬ�I-,����Q�D�A��˒T�#C?+e~|����D_�"��������.�ݭ;��>R�rS�u�=�2�'��D�x�.nI8 p ��p��T�꘶�hN��&3�w���>5Jx�U�g֞y1�xX%}~�fqf��hc�-��}��p�����*P�����C�]�_�Z����k;��K�A���	���>Ր1&#�ڗ�Lpƨ�x'ߪ�\�Ҽf���@�H�FH�aͯ�9ͻ�;�#�d��(�؟�n�16/��6�`��Q�(;~�
ȍ��Ws]�������:�Դߒ��m�Ɍ�AR-8�?Z��+�V���b�;j�x,�r�%8B�1L�5�	�ca�L�U�i/\ZWҰĶ�rd���K��ے�����c����9�#*����\{���I	e���)s�&�ܝ��F�"]v�ε�p(W+V�bsB^\0�M���u����Z�0�1�'gQ�kr�)p��75y������=}g���X:l� ��7<C(鿯��.2�(
��j��~��ì�W'�iX��������rRB�!52
����Akk��y���[Ӕ�� ��[J��K���q����Ѕ����%�c�Г�1�9��Ƥ4΄��#/3#~����@�'Q�9@�
N�5>ʄ��3ؼ�!Fz��,8a#�!!AV�78�0}�t ���K�M��7����|�	Fύ���M�DޥQ2W@�y�����fA)+q�c����a;!v��1��K��.q�l3��'��?E4�&�3��x4��x$����������?,E/��4�@�N�T�~�*Q4S�z�,��5�D�F�l��We,!KRbh]��xk���d*Ni�0�	��B��A)$����R���IG����"�� $�X�^���݇���d��P��?a�i%�:S� T�F��ls��(��M}H�7��Zg��룎W�Ƚ�ƒ�-gΰ:j�I1��q���ݝ� s��l%��QE;\8�*w�����U� �*ET޽�*��TĘw;VG$J�=��ۍgm�����ً�V"?^?��4�trf��e��u��'w���Wp� 1C��? �춴�U�w<]��	�7 *�@���캆y��u��^�(Q�تd��Hz���S�4g�4V��li�������7�{'���g1�*���B��
�-�?�t#�Z8�9I�Q-Y�D3C�S��:�N��6�Q[6>#1:�q�>mAKP��7&� �l����PƯ����a�̇�bB����h�p����rw87����yv�;�sK?Yԥ�$
��Os&YJ�u;���a�x�N�Xua��V��Wf�3oA���*@i� ��3BQ�d����p���Jb$���1�fA��{�(P�	�i�pܵ)�����Oӡ�JRH���;WY�y�?P�أD|�����"��ߐ���o\aծ�1�M�i��%E�>�5s��d:D���x��t���#^���+h"��@�W�W<r	�*�#^s�'�B�Dbw�.��J���������s?�`*�>H�k)���J�T�F�P_��Q�B���G#�:��f���֟?B]V�5��hm��-3?�t`�?���AC��NL ��������*(O�����B�%� �7o	N	�a���S�g('k.Bdb������m{
vF���ɥ��A�'��%���Z&� d��=A��U���	��ސ�~��$yon҄�Lc,3�$���:Cn���d�����4Me�\�Pjܮ<-X��N�Ш���Քn<gn�GIu���x����诎��s�V��r�Ld�Ȑ�I(;���,b ��g��������q-�*E�@����#�cju����A����`�fW0&dUTȄ-�n���W�tC����П�xP����F^�g�N�����2��y�eK ��-�<�acoM=��$�cˠ�h`�)����R��#&�z�p?�� ���/�k��!0���Wψu�ҥ�u��K>�4�����i���ӸE8�����Sk*A@�I��M�ק����n�à:�i��g����"E;'�(�x�{T��z���c�d�u	I3����u�c�;PM/�'h��#��
���ҋ,N��Pk��}�!z�
�L���ѝhE�ݗ�����&�l9I�󁠩"��ha���,ί1�	�?�w���Y����#�t*ɵv*�����=z��u��5uoQ���']�-3�D��q�o0�z(ɐ�nK|?9�KF���b���3���� q�Y�C��ߙ��uZJ�=t;0��Ay%(}��9}Uf��Y�zf�d����ۑ�d��q/R�!̐�#�~w���}�I�+������w.6�r��z4���MH�N�m����/*�}�.bM���4���C>h�0�e�Ff�`c��I�m_=���URK��x*jI�D�w�C�VP�8aN՞�P��;�=�S�&)i�t�<f��E��3�pw� ���:����u�x0�}�RQgb&C	�,��na�)� S����Gu<�`[�D�5I���L;*�������)]�5��N��������lw�n�rw
�����:���rF�Ĕ��"�h=ɬ����9��ڐ�ʖ�G��
�	<���C��Sh��|�YY�ȥp� bj^jN��2MQD�=S�!�ew^��
5[(+W�5�1C iux�� �n�l!���֖���|�?5A�3�	tXr3O.�
�L��\���w%�A�;�����D�m�	����s�����aFm���ͺN�����C��iq�ޥ[�-qO�=�2�=�a��T�<�E�&�^����ٳ!cE䔓q�r`����d���!��o)gK���P�P{�Ψ�y�(�mH*�oK��SѰ̙X���>K��RÇ-�4�2Oi��nM��0K���
A7�b��"��32OmS��x�����2�h�0�jk�!m K5ܺ�)��d���IT*���8ћݒ��i]�{r��3��ߐ~��������&�r�1]�b�dө��oDɸJ�l� �b��k;�y�uKxL���s<�:�fo�j02��ѳIE��#��NRV��O�#[L���Lp݄e�)���)���E� ��#�;�
������B�	� P���H�m񇪰2b��-��Q�*��-LҼ��*L�1��rFd�z[S�c���=B�������;Z�*=�ms$u_�Z��o����-��
�
�K\���2��4Ԃb�"��R�o"��p�^Ƭ�!�?������рk.��q�w�fx��Ƃ�P��Zo��xA���}`�A���-�2��ng�-b����ɒ��ck<`�) �W-1kB�Z�d1���,l!�b�\�9q+^�\f:�:���(�n��\&+\�?�x@Y~А���X�?0J�?�R�* {��GTD��t�͡���#A#��${��|�t��	F���,^��l8��v��Lȣ�z�:_�`�4 �NN�+u(�P5���hZD8��"���.mT�C�Q�`�օ���8����e���９�}���u����͓m����a��w���P��X��������Vo��,�,ݓ£���9X�� �z�A��$�{�/<��~	�V�,ϰ�����	|�`7#Y>��a6K�x�����A��~��z�Tߺam�+���ӫ�/����b#.-e�<�N�ě,��2�����Db��he�]A˩�tC��������P����u�˻'�[à��KR�G�o��]u�:�Ro�$|A�g��6}S#�ީ���6���QG8.}��k���=!d���ïO�`���1� �w�P�$~g�?#=-u�}؁�I$�����ߊ�n��Y��t˽ʡ{Z[�� Ov)���x)�Qר��͙y��_'�pc�<���7.a��U$T��`𾫬(��HJY�2�s��dǨ�n�9��n��ʍXEP��z�+%����t�ŚA8p��E� �����Ѕ9���%�/v�qO�R��R�o�~J5�&`��hy�P���L�Bt�"��H��,�(R�k棷�,�f�@/�&��(}��)i���4����|䬒�%XmTY�x�v��ڤ^����к >�ǁ��s=���h��KGO5<�%����V�O��h+^�tGjuQ9fzD�o�&|�z���Оop�$EncL���΅ ����L��MV��wϫ�4CB�	�R2���R�j\N�V����u5I1V�l����Dd���uC���.�`�vw3���çI{�~*�$���l�B���]�؂+_a�l�G]����洺d�ݸ�T09	¢
F�����ʏ�B����>`�l��PX$����n�g�[l�1c`�2�a�d�i��k}7�#)F��c7v�mlKPK/�rn�����r��~*��`b���ą�d5D{�n'\Յ+�T4M���4֊B�O�C%���9.@�s��?Sw3/���	a���Ř%����C�x�ܐ �!�pT1��-|M`޽Z���4jM�ʃ7�7���I�272Kh�'���Ty3#�d��[�,�S�_��)���~`>y����Gq}�;��ۧ��]LL���0޲��'�0�/��0-�*B'N��� /Zd����������Xz��
?�K�<�\� �W����׋�<t6�6��֩��P������պ�-@�17x�����Ҡk	�d��)�7 �.'ݲ|B��7��]�H��<{P�1�q��%�T�E؏T� <?�e��q_[�x�
���
���Plۢ7���{`��g�2��#��?膧u�ޝ��D���-����i|ͱ��J�L	�O޷x�A=R��m8;����6#?@;��<W�1�>���"�k6ᗙA��2����,�8Y�����֑�!�QmF�b�7/&�KΥz�?��r��������C��&�ۡ���c�c�M,c�em���2��C��?� \�fU�`�kլ��h�#��Q��e1+z�A��T���r@�y�~������"����*�Yބe�}C���ٞu��ݥ��T]�!�K���U�j��m����I�!�M����l�cFMV�6�ent�M��[,�3z�ٲ��$���Vٹ�ͳ~�m��Yu`�ӥT:�s��=�L���m�9����~=��v�������WW�~|c�҂>�@�Y�kyg��5�
�nl��8O��P��1.�KĊ�]s�ERAU� !�#k���?����� 9�7���߯�^�}�kKi!v;]<v�*��Ff��)u��Q��l�֠q�<�w57c	�����ӑ�2�¥���A�d�)1��`��K?�A�,���s�/'k0��
IS�b�u��Æ�d��W�3���lZQ>�!���Oc�ڇN$��=�����c?�'cNӤXl�X�jW��c
O�jX��X�V�qחJ�������g%pYN*zB�/Ys�Ő��c��2Qcs}z�G���QS,w���-��7MXp���s"�v�/�n�~�x��'=�]�^���1��aSz�D��-.�9�<�C�
ο�
�_4tZzx�!UfJ9KP����۵MT�t�~0�_�wMހ��ؚ��L#�L!��-]j�Οi�̂#(P��[3����Zp��5��y>�Km���D�z����c_����{�h��s}�Fs��I->�|���������!i?-��B}ˮ���f�@�`?������
�y����8�x�r��
B�e7��y�z�sʰO$��[�u��0����0N9r�K
�b+��Ϋ��t���/!���k�9��#N�R���@�P���|"�\�+�^6N ַw1���+bR)���j2��LtyV)	k��_�(��_Th���iwO��W�/,��{3�5Q���H�boh�/�׹$*�ʙ�W�W���^��z�ݳ�ɝF;��q���G���01��da�u�W��D)���I?4�Gy���O,u�bn:���7���n /�n׸e���	d�"<�LQ��� U�X�(�R��Z�J�;��2�� �<`�2�%+P�W��$��Ɂ"���6D0����2	w�QH���=˅�]]�R�a��}�|���ǵ"e�|�	�a����=U�iL�.���<�G�p Eo�!����-)��I�J���,�#�ಓ6�=r��[��{w\)�\?c�FZ�1<*&%�+�;G!{�
��Yī�H�e�S�ٯ�K/7��69�����~$�og��L�J\�)���g���t�f,'o7`��J���Z���8z�Z�E<6+�� ��Ӽ�����6J'�W��V6x2 cv�\|����[�o�v0yZ*uEI�_�|B�fн/��������A']���v�g����ժn%%{�}��,�uq�<��D�r[dk�VG����99-�:f�R���Wԭ^�Iv��v`;m�����y�R;��ΔQ�������)]��8T���Jfe�bC����j�4.��Z�!���:@��� �0�����oa�*s?Wd��w������͚�y�y)Y��)َ�Ʊ7�ʝ �m�DT�b���p�bޫ}�D��}��p����!P5�����$����X)�o���@8=A�8����B.>���A��Ht�*�ܚ��S�\.Йo�&��Y���Y������(�:}Y�t�^�w�j<5�G��c�Ls�W����*�`�t�/��;^��-;d���0���ޞ!���~W�к�֛���P���j��e����/��rEmOq/�le9_�&�z��k�߷��������蒏����\_��cz\�ދ���iC��fd(�]jC�v�5a��m�ɒ�B�Ux�޶�hn̞a/��g�c�4K �T�Y,���̦�Z
bt$��g��[�&7�sH%�_1���j)���{�Ɩ�j|�PP��Z1��5gZ��GV�a|��je?���,��M�;h��UY��N�s9���D �̱!�b�3j��~�d�|J�Y*αѕ)���eH�>{=H�S�%��E;�a��6lr��dRיRuK����
:D^�~i����O7�ஶ��v�0 	���=��G�m� +��jQ���mQ�ʥ�-��G�H轅)���ݩ�$3���K(v���5ƿPg�t5��n��0�T��rJ)�Ae|�!@Q� \7�Y5��X�|��V�dp��
3��nEu��F)�
�G��L���Q��[-��x@��F�c�)�SA���3����+���@���~����R$�|�����`���1�ؔ��ܠ_����������A�3�;3B��6	�@t�ķ���	��GE��v:��4�����k�fW�F|l���8�(�-)�]O������G<j@��\��#��D>kN��d��k��B��B���L9LDf��Lh�M��*3E��R�Ȼ�J�.$�i�O�'2�O܏gYY7�����/�̿����,-���R�gnކ����]Y�mf?y6̽�z���=V^��'ds:i�0߼�����Wz���Ms=����t��]��i<��������>��c1��E�ٯ)#���M�_��z�X���ȓ_^F�$��)|��O[i^8D-�"�#��J�NH"�<��	(��	,B��
��U���+�-9"e�):v���؛[ɮ��TzK5%�sD��ʓk-s�iZ��m�����)F_�$�m}8�Z����0�,��r�Iٟ�Z�r{W�S��2���!�G�/�v@��O�(���v����?���ǋ�q/K�@/�j�B�� ;���$Kx�jS��Q&�B�J�<���ʀ���t��ρ�6�G������@��jsJ�pƯ���=�*�;w���<$��8���gw��N7�0v��y~l�/4X�V;=S��?�w�=������|Ak�,3��p/�8��l�$�w�k���O�S�G����:8y�������B�F�9P\����cxס}�4��6^�~1��5�B�kN$U���d6[�@Wv`���3]�젒��j>�M�`o>� �Tv�]� ��54�m��dF�(�y+B"���d+�%�IL���w2۱�z�%Ί3CQ�=���_�(Ƶkf� '������0 �&������>9��^R���r��[�9Ye� >��8]�{�C�D�����l���|M����Yt���ԝ,'������㈾E�ٸy�z*ΖGH�,�F�,֋���sv�>=�B��]wXQ�i���g��q�\Ȟ��7,;0Ղ�)���-/����}(�P���G{8�83��<7��Oc�E�ß�Ƨ�x:�<��y-o��1o��V����d����^z�d�|����wO*�}��D݄]?�'��"�;�[g���5m�EG	��������H� �0ė��ؽ�g�謻��x��?\5���m,ܽF�Y7�	5Z2�6�M��	Y�֝��a�s�<�+'U��2���iI��58E�	Z+]E=O��?�5c�Ftn1C:2��jLm���kt���
/R·�����7P�%9{���V�|�A'9�c���H�w~���z��)�5�&?m0��a��MJ����x)�����Y�
m+^�}\&Z�tC3H�Q	Ɏ�ߺRv�����-��"�J�U�L`>��whz���L3����D��.�w�z�YL���J�XD�	`2zq<�`�	�ev��$�vQJ��+W.��/p5��l� <�Ǯ"Y��]���8V/���䴭�Os�Ϣ����m������ʗW������!*z��]��/?֩*i���������<��0��[��ql���\ޗ�t����"���/���!���Q�{�������>��6��Q�����O}v�D���&~�Q���D�w��}���'�K�Uy�>�G����~���U�-��R��Zb����}Id�-��w �3h�٨U�!l��u�:_���,�{Hü~(+��O�B��ZO�L���e�i�SrW|+}b"�E7i�#��l_B�0���M���q��ѭ4#a�>9�5�����#�QoWQ��C~!����UC������oF�<Tl,���o��"O�A�ʟ�X�$���;w����F�9��r+���[�q~Tk���P\��KM�}i�>�T0M`��&�劶[���y���ʜZ����!�<�Czj����پ\&�����F��#�/O\�d	�toR[,ƕ.A/ ���������I����;��s�4�U���C��@:��(4Ay���og�=���TPߠq�[���o�ݨ�&�8�ɸ����e-aQ�WV؀!�x�	�:�G".eNVSK-0��ɻ�Nl`Y�\5���hdD��m����w
m&���l����{�ɤ��tN[��߆�9˰E��tOÍEm�h��>��:�
����U�EL���m�6�9�MV��6�k  �8)����nܑ��Ѡ�)��9HA5�����7��ڹ������Ѝ-�R����W��5\�*3,;����C���ή[�'�Z�C���Yl�Z�~�s��<���k~#P���ؘ~<���4�����)�}�gX�e��os#ݳ��K�\��2��1[�7�H�Y6��٫+~r��믘�wU��Y/~u�9��O/�U8RNG�A��I�6	M7g�!;�b'Л6sͱo63Y�ڰ�G��;ͷ1e�ݰB�R|��2 /0~���F�<l���z�jfy��ꅅ�y	�c�̪M�SǛ��?+JG���M�u�awu&�X�Z�.5k�{����r�-�-���qvޖ:��탞
�&ùQY�Ԕ���8]�Q����5�`�>o+����΍��5��M���}�|�����/�|�E�`��=�A=`p{�-�O��8F�<�}=|J�Z��+z]���bY�7���o�v�'��Mq�04�&��t���9�7#A��л5�� ���3����O�WH�O�]��Q�S�Ĭ�e�S��E�t:�[��k[��~��V%��s �8l_����Za��ÙiA�����\\���d�`Z�'����yz;z>H�b!��g��,�� 
qBB���HǓ���p�XI욽z˩D�S,xn7�2���&�����j��\y�P|6�g{���O�{�_�7��G���u�}!+xkP ��Y����)�����	O�d!�5�$��L���wp�>�.3Î�G���x6Z#�[`Ѐ��`��}J����Ǐ��9��l*�q�ĎD�&75�ZF��4Q'�9"Pq)��7� ]��Ii"��������c3M"B�8��d}(Q�c׺Ml�g���8�
u{w�[Ue�_>���M�-#�˛����ž0|f���~`��+�{vp��X)��݉.�.'3�Z���i$!�p�%�)Tn�������F��0dMD�������=EV�p���E/T��$닐=2ܢ	t��ȩ�@it���ǡ65U��ۀn���C�%�R�� ��P�k}��s+����0��g ��̦�mu���Ë���rÒ��>{�9S^5h`��c��7B���T�&�L��RPE-��K�ˮ�������ʻ<��K��<�k"���*�ܞ�=2A�P
ӎ��[O��,L���6RkQTC���+��D�:�@}�EgZr8���.���w�岔d{��Mͫ�A�Ul/WIv8�_a�V�33iI<JY���px=h#�Զ��K���'MZ��V��r���[>Ck�n,�Rv>���50�t���3l���lCaP0��Ys�������1hk�p�g��]ݢ�Qf��I�1�U<�SD���~�M}���:�u����79�N�l��\�Ғ���#ѧ/��5ʋ���\��m2"NO�G�9�bЇ���G9�lf�:���\�1G����W$-8ȫ�?B  Hy��sU��*�^�����D�L0l%�W���ξ�o��٧��N�T� S7
ݘn����9u� &�"_'��K�Vg�b��:�1�ʓn���͛8�O{C����O�# �h�s��c6{S����\G��J��?�RL�c�Cέ�#�"���ߠ�t3���2�AK��R�I� %p�#|�.>����^���_i�}��|+�U��乇��5pU����BWw�;ȏeF��������ly��&�~��5�3�,P���ӄ�?
���f!����������c6��7w�S뇗�-��H�M�Eu�t�)�+�D�?4J%��^�oؕr��w;�?~߂�����8=��}l�/!a�s)�6<<�9���!A�8s��r�%�C K�R�dd��BZ��=�lIK����Mﳠ"]�"�!Es'z$
�ϞH
�;�� �4>������桠���:�ix�͑��X5����"�����ڊ��Y��p�!9��7x[��횱�#��BK+n�'��F����;3K%XNB3�%ߏ��q`x;����8l��4|�4 ֗���B�����zJ��~�-k�����{9f[��?��䄷hA�}�0�,:2;�����^���	[!`�8���b���	z8�@�u OL��/�0##	V�a�B?�z�@�����{�ZD�э/�����F7~�RvjWb��?i;a;ķ���E#~��i����lm�X��#X�8���y�U� �q� �#�]���Z޵���)�b�����!R+��2�'X	@��*]�R����	_�5Gƣ��'�!ߩ�����ᣨ�� q��d��r�-�c5/�so�	r�,ٿ���r<���2��֭g���9�С~,r�9�o����;~Дb˿����X~��[���.&c\�{����N�:!0Aw{"�hb��y:۶E�|���^��a���?��ҧ�L5S�����}Z�?X��Ț����2�����'�����:l��t�H���\o����#�8�	���sM�U>�l}-�^|��鹥��_�ަybb,���~ 8�r����{�٩�6_*��V8��n�%���=�D���Bb��&3��������g9i�4yo��u�A����s�l;a��E}��^1kO� ���|�/��-��^�F��.<�='� �S��+.Β�\����X�z���m>�i�
��^V>h�#	�ͨ;�;V�0�;&O�3:��_K�7���h+�×�t��z�a�L��To8,͸b�[����u�#��4�u#��U��34��.r��_�7aS-Ț��8St�w:O?:¤7�!���e{�_�/��5�|�)��n��6��nL���q��P�{�r ��DrDI+RМ�Q���n���Wj���B��Ep}� 0X*H���ά�6�鎫����
���M4�l��R����(�5�g,�r����l�)���4�Ƚ�Kű�PK��~WӁ*L�t��Y�:���Sg�5��^>��5Oc�z�o�Ab���A�����N��x��+�S޸P7���hm �����	nMZ�aѽ�C?U1<�w}h�\�v�MS����Uܡ�K��Z�^	�A�G?��m��=��9F��ST�W�IǘB�f���N-6<h��37��_��qȼ8�rϦ��[���d�A���G�a�^��$T����O�2F-�"N�3IT]3<	�k�p�:�܆��Of곬��مSD匤?�����H�,$��k-�9
�qh��@W���w.��P������
V��>�anل��缙}�,L�Ά�V���L��{�EJ�޺S����}r���k�c'�c��t6�Z:O��ކ���z�+SG��=�Tڣ�&&85�X"^J^t���K�H@��@�"xS��6� ��A���Q����$\���ܳ��oH^0���H~�k�=����a�Uw�Q��%B�u����f�/t����<��*�{��Cf�!�S6q����|�NS��H����D�W�E�i�3�n����n��A�W-y���y�4�D�DEU|�bV۸a&�iA%l�w@mr��O�,��D�i.��a��q��U�}:`.��P���x�Ή��3<���G|���DU�i��F�)�P�2�a�y�q0����d�!�F��^�0t�Au�����j��|O��;�_.p��<�-�!̩��d;�h�Ⱦ�YH�y�LL�.q��1�?R�� ~�<C���/�Y�bK‾*h �7 Ƚl��X��Qo�iP�@�s����Ė�֩1��+�F5sCB��60� &5�D��0Y�0��/g9ȹ@���i��S&
,���9�E����ZE�LH�@
�1�
�I:B<��@	��O������z<?j_�� н(q�H�>f1X#�.Ʀ��Í=;������Ũ�(�섭�5��t_�K��@���l��C��&�$�F�ɣ�ޖ("�:�bi����"��B�F��٠�=-�O*!������x�R����HŲQ0^8���)q�_*8b�E�����2޸d��� nO�T�4v�Nb����a79��r�B����{/�M����2q�-a�X0�JM�kZ�+|7XZK�X�����|��0k��E����?:�W8�PSA�6{�}#��`@�.�ۜ�t�܎?���2"�;묍{��Nl��x��{�]E�h�i�4�%�Y�;s�B�S��(D\[ѣ�ǋ�X��G�>�I��9$ �&/�A��v�P\ł���?�Ưlz!��Yc��E�3R��^xd�/�1�ߤx�)��p���t�p�^.U<��dE$@��� �E4Ӯ��f=�X�}���kX�5��W�(�öw_k��L�`�Eώ<4��V��mG�r�������=B���k��%�Og�Nڞ2�	�+{E���e$�KS��}w��� uU{%N\�Mdog1U#Oc�I��
����H����O���ޕw&j��,� �ܷ�͚u��eP֐[�ɓh�����]iJ��)�Q�Q�[q���>�ٗ���kK�w�ƀK����,�����yB3������R+�ò��}�l�(�&u��R�=����c1}����>a���-���Ϫ,����S�K܃�xmV�ۨ���0�<��v��Y����&��Ⲙ(799êȊ�#/Ut�R|�D7$�VP�ٺ�z����UT�0��L�­�1�gE��x��z�8�`j���)+񼤫O��.~)N>�gvXY���f$���y!n���)\��Z��(2�;�ک�1�*�Zp�/7m;N�0 ��4XL�[3�2Z?Ƌ�M�O�9v�Td	��A��i�Rn˿��[�Ό�>	��Y|�K!H���<y�v�cwK;I�o��{܏�j`�RT��6y��L��j����z��xu��w��^�9��~Ȑ��_���c� �/²�G>-��ġ@P��%4���iƛ��j�(�`�-?z���\�?qt\�����2'���i��7�\�o$��VBo����׻)L��yXD�	M[:��yJ��%���u�ȶbyR�j
l������k�P|�4�*�lIj���=yW}��s��F�i�n�X;�B��<��.  r���t�Wpc�tI�ur~Q�?����/���``R^��~�.�6�(� �f@�ub�|�mt�.Z�Ň�=k������ k�f�d�&����W(��u��0�M�����lnԞ=_�YЖ�Zu�0c�5�vJ�TQ�K�h7 ��YG|����+i
B�yrJ��jvR�$��(�$�-7ſ� $�3�4�~�Y�Y�1�A���$�:i[N�4�.���ڔ@�B�ڪ��M�x�zz���ė��AӇ4(�VE��3�l����(��ʥ�,6����ա�&J������t�^�5R��A��(�z��n�׽Li��jr�yVC1�r���cR�l����g�%{�^��j����,���o���BrJ�p�=�]Gk��DeJ-��ZMo.� ���p�%��$��ъ�Cg�9���l2r�&M�BK
��7]u:�,Ƀ��zꠉ38�v�z�'��9�$�[F=��S"�'�f�(oc)�5W��IL�k?�(�ε����;;��|5�:%�M������ �`|�m�sꋞ���tf�:{ba�L5��n5�(8"�))g�����5K�m���q�T�V�iv�g�"Iv��BծNS#�:BD�.��vvJ��+"Up�Ϻ����X��.����Ͷa�c?pO+���"���=�*�A����+<�.��Q+X-^��%�Z�R�;�@aA8��B��,��Y�Iޜj����)ޮ��!;G��94��"�z���!��1pW�g�;�[:�O:��d~�Wb "�fU�`P�?k���:V��Z�?̚�S9�e�|��\�§��-��&)6�Hf�g*�n��T���F8��+��	�)z���u��U��l��G����r��(��kN����R��ԏ��U�R���	8Mb�����7��r?qzrSh��������?���>er����n�ں��5b��A�zv�w%r�@Wkm��g�D����z	<m�:�0�J�iZ�������:p�r�]e��NeF/�4�E����0������tE��R>K�[Ӊ���b�$�P�>P�ꘃ��S�Hwk��n1�9A<���=J֦�y)��<�68U%_V]a>F�<��?��IV�ۣ�F0��οD���kB:֔\7�	��m]���[6�L9sj��ŝf����!�F:�\݌�V�э<�/��+݇-!��/�gj����~�T[;�Uf�@�_q����̒�[�����l��<iR�"y��f��J�%Z�8�ͷ:ʂ|��N(z��P8�k>�v���\7'ȋ���.��H��{.�p�Z���/2��X7���g<��7�O	�μ�N������+���\�Vpvұ�>�����s�K#��t��~�N�Z�Sf�737�Q���� �6��$���g�ޅX�p�H����dP���x��˝|`pq����u����B4�|���R�g��S�.0��$�ᜁ]�~h�J���B�t;�(qf����W�$�-�P�UZ��
���S����KY㘝�vp6����@-��BԜu��'�ߦO��(2�`���y@���qm.K�I �H��JH=(�H:)m|N�v���"GI$i �ƙ���1�N���i�,�Þ3��դIC�F�&�:%>��"��]1b�MS�p�!�e_*�Lb��4E�����65n�n��^�G����?J*��m��)I��d���ƹ�3jA7�y/o�&2���쉰�n!�PfA�v7���:c!8EdⅬ���#�R{��y��"�l)�Vw���t5��@9Z���H�p{ѥ��γ����?lI^?e���1���>}��"_u�l�ZT�&��&�7V�u���=�]/�&��wZ�~O���@_4(K;�����E��~[Xf~�f #��ʒ�,��H���(���h��ȟ�n\'� �����7eI^�y��}�1�U*T�$�4b{��5���#�1��l�m�i4�	Z84��}�^�U5�͑:k�?VU�A&��^U�ib�R�b� "�l�4��hji7��=��_��*�w�/p:��H�u��e)�6g[�X��v���$��{�H�W�6Z8�ZY3�{F5�C���j-&��8p��9����$.�l��ڋ�&f�1�e��ʄA���_eX�`$u}ت�	1H
0hs���2��]�22g�w|h7*�6
�rw������-*7����S���Ɖ�VS�[@Q�yk�������	M�+ە]ϥ�j�Bcp1ڴ�ȡ��h�&��s��0֘��`��p�t�G-#�U?i�NnrLŭDg��Kį�]�Yxod����?A��o�;��*�RN����i��^�w�A����%�Ěg���Y�љ�
v)���}M�4$1>29=�oF�,-����A���dG��m�j��j����7?�S�������:���V�Ҹ�@�����%VBo��
�V?�8��\ɬ9�Z�/��1)1pH��-!h�'��l՗E�9��d�-�T�$$[E���z��/�Q�:�2v!4Bx���mLR���yBWǁT��
��4�������&���M��Jl#�<���s�,msB��M��U�=��g�|
b%r��·���N��S�=����빚�@��#6�u�����ql�"n� ʟ��sZ���5���Tv��
lL?*6��:I W�U
W���z&@(M;c��qg��~W�H/�S�F.�6��,��
l�ƣ��|I���=�4c;�	�2w��"��?
�0g29���:��&�Q_!�ޤ3;d�R�R��/�^
��^<�:�cp4��?���V����ŲU���/��p���z���sEi.B$����:��'{�@i(w*�7�S�c��&.D`��
� ��P6��zh�.���U���
A8��9UIBxVl����#Kp �)��p�KV*a4$�S����>��t9�#S;��+��4������Y��� ۑ+V�
���S�j{bw?~�p�[_7 b�rJG�j�S�)�b�6��hּ/����9m&�)�n6F�E�Gʰ���Sy�1Zȹ��\��;��M{�x��J읫�N�������L+��o�����gMh\�B�ù�I�)�PyN_��gU���z�Ь'�hK��g �Ga<@ KS�俰�ܙ�^}r�u�g�����I-�;R=6���:;o
�v�`Y�3I����Qm�e��� �,�f���d�7�w�,	�)"�M��s;ʺ���{���gFSՋ���z����l�Z��AQ��s��)�ʚ�/fZ�k���$�����=����̨ '�J�1S�idހ��-ߔ~2Zt�v�)�s#<fbE#Dlp����(R����]po��+V�9�ׅau���o6�m��θ��+#k��N��1l�x˚G3��x�lGV^4���/�w^T8:U����D+��d�9qfN
b}�I+�JPJp��H�'�V��=sa���<kU���n-����C��lo|d���¨̂�=~8��X���'
��jx���/�n���/�Ql�.ɔ�����.�o��i|=�H�B8"b�ak�sK$�i���w@ �9?�Ga�P�ч��������O�6
^	���E����JA�efD_��|9�Z?>遞[�g���W�Y�U'ᣮ�^¸_�Uz=�����,&veA��Ei���4x�l{�>�$����� Mj��4�i���^$����Z�5W�a���s+g=��m]���U��E ?�*z���"�$�
�l�:g!70*!s�)� 5� ÷��6;�q�7X���]��g�����cp��h̵��B���hӞe�l�h�%x�R�}5,�4� ��\sΏ@����;�˃Y�7b5ǩ���9��
�D�^��[��?�[w�,�������7M�#���h���W9���浘����|n���5�B� rH���'Eo�q�v%; Tr)�#]���A���A�oB|�F���=��`�+;�Ĝ=;��D�����?t0�5��<ҕ�t�cUxB�(P�ФV���?;����n��&uuu!�jԬ[g�X߄�L�V��k�qr�(�0���K�T��x�9�q^%������b��ZJ7���@�T�����[|���>l{	MKA3XI����Ģ�RU~o�`�����[;����!2��F�u�(@���^cE��z��׶�$N\&+�&Z ��S�_���LH<<˱4B����6ΘFL�����co,�ͳ����\nl�f��kU����L����s�n�w���J���⚱+"61��g��׾��}z~Ns|�!u��ch����2������X��tlP�!ځ�
XҦ�3h
�T�wFcF7%��
��@��N��~��A�0��z~'��U���Ϭt�1�-ֵ
�!&\�P���PxDuNve�JFxJ�t�y3͟2��"�  �@����W���1d�F�5��?�C�;cĨ(;aؗ�L?4��}
q>¿�Y����،9��@p����k����Rh�d�n�5;[���:b\hN�9d����D8��ʒVP����3�L�Fר5���j�Q�DOQ���E���C�Ms:E-+��6^ǫ !ǽ����y����Ƞ�s�{ ��!�����L�G�e��=�V�`�8"�1"i�#���:N��M��\xb��T����Ǽ�Q�0O*���F<M$?�T9WtUEG���=i7{��0�c���/W��/>�
i�"�$	�e$i�%��T���)���O�l���!!<�Fy6�{0<Z����t�#��2}��
�as�����*џ���j.�t��m�G��G��	�o���	iN�e�Ҙ�� m�)W��QfI���/H��ϭ�^ �Z�R�I�Y˒;��i��e�/x�mʇf�	�������j?O�S ����=ʢ�|���&KF"^t��|�=#=�U��T��s��k����󜷷�pwr��C�-7[z����38x[��(��<h,|7��x�qW{,��aL�:���@Z���&��Z��'�hZ^a���:[�\u�L�2aZ.i/
f�~d��`x<��ok*o�z9ьR���W���//���Q�y�$=C��`sX@]�ƒ����Di���]u�,�<��#��8r���l�q���S]���D,v���|p�\��6�n�ȋ6ٔ��b�ꋋ��*�D� ���`m_h��������Wr� )�Dl���������4Pvf��Lɐ���#��j8|�ũ{&2퉗��7'�V�Fn�I��k�B&���" *����B˓�h�iɓܭ,(�� (r���~��Է��7�[S#�&���l�K DqԷz��HMg��1���*ӣA��Y��\���c�k>d�߇�ԉ��{ 0bP��������E@m��lCL��ʩ��Ǉ;!��\��m��p�q�[4��[D[n� �
��*�"���p��WNΈkd���*iv�mx���^�p��]��-oJ�k�iـS�����2��m�f�$�-���D�sI+�؏�\����Ne��#��DTBi���0�j�]|a�,M�iLe�r�2!>']�4J�|^��X�*5z� j��,;��)��hMA31����Īoyqj��b��n��ɇ��v�>�ʫ������������;�������	N��p��vL(�740f�
�>��8� ���a�@��'�4�D4�:3Z����t�����b��wgiy��S.�h�d���i9#t�1V��0�<��\�I#�v�2���NK�$�8�L|-���(T�X\_P�O,H�0eu� )Ϙ�:�2:���@w�8H}9�+u`�,�� U`�b�����-y��1�A(��jl��:Յ�c�ǵi/��]Bܢ�����wkDX��بõg�rZ�#@*U7��(,}�i�yrE�G4eHK�{��˄��v�j�׿����ki�"H{-6��/������l[�_JX���gR���1��,2 a��³��mĢ1��V��Z�x��s-%��8;z���Dh�����:��`�}O,@j����*qϽ��D�d�/��L �f.9ˮ2�A啑9s;E� r�t �|cz��0<z�K�R�W=
ߌ�p��̭/4����p�O��v�H<,�9��91�"�r��m�d��M�оt�������;��u{*�p.�.�pO����R�|ʞDj��"c�"ۮ��TP{�K�g���SM�{�Ͳ�
���T��
���Pi��'�����P�s�Zd����q�'a1=���f���!Y-���l3:�Oꛓ��C��?�?�h3y�T�wN�%��%�?���H[o�
����R_9(;K#���m�M7C�"h����r�<z�Vv�@1H�G������	5y��)�|x��M�(�F�b
.���d?{t
Kpʒ؅�����
�R�����ꐧZ�9ڻ�|a�T&9$���?P�S��݂S
�:n��磅�X��!D��GK�n��b7��p���3��Ic����{9,�j�}���so%��z���
g��8���S�I:x`O;Y�:�H��4���t�-k83VY]�n���]ݚ *5I�6�s�K�����H����c&s���w8���Ł�&F�I���.����^�kPF�|g6J� Q�5�����v�,��8�n N�HB����H1�?����J��]0����1^�൶R�P�\���h08��NP�&������t�*�K!�,%�4��sؗ�4�Q�5E���'�i*�b�u���:��׬��̜�ʽ��9*�x�P�y�8�����~��w��*r-��@&;]�e�����4�@��j�7�/k#��Q�9b����9'�v���5sO�c�q�.��m�'uw�ǻ㩟?Ϫ� �A:t;M���G!B6ɭ_I�=��î�i���|x�ʛ��f��~�9���	
��tt��<�tW�6�{kSU.�'Z��a��R]�ژ
&�LY8A4` 2X����0��1�Z_F��������W_��| g��L�q ����t0E0#�#�A&0������g�sqN|�w��aiiV��?FCF>5�t�r�G�H��#��r��J�%v'�'�9/�Ճ�_�������$�@頒@&�	��Hj<�#�&�V�Iík���
���]h`�%��зn��t��%����`��>��n��4ԇ�����}	F��̤W`��Z�\�l�9�`Ή��۪�_��i1ʒڪP=�j~������zfҰ�ܦ�S�mi��@Su[��T� ?�O!�� ��s���ݝ]��cF�(�p��l�-|Ӥt�"�+l���D<|^��^W�}<s77Z1}YU�O7GJ�4��5?�%Ǆ�H$bؒ��?��h�g+���R�i[pː3� �j�( ��g7�ꌉ�,ꄗ�m����$��?�V;��U���{�[�L?>^�
1��nFA����*9i<�C���}���s)���&�R��u�f �)��$r%	���˖l{ [v[�O����3�e>\��^�R*S��tL8��8�V��py~N����fwf3_S%�:A6[l��D�&='[p����p�-���k��A���w���m��OA�s����� �z��o��MW��A/V>���GB�z2�&�s&�8N�V��`Y��I���`�����mjI畒�#h[(�Ol��k����Nk'�P������A�#}�ҡ��U%����b���������cb��y�������1J��
v��@x�tY�;��¼�Y�;���=�b��b��*��e ;*޾�ZY=�j�A+��G!-��L�9j�K�P�n�-J/�$�!/��l����kq$��ة�h�8�E��>�:���L7��x��t*{X����)6^m����8`�[Ǽ��w+;N�,~d����Q��V���W�{���]�:L�!&��(ej����I����t��t�+E]���[���%�D˧�m�?H����§c��v[h�я[@(�K�̟���\:B���p/h���}C��C��FD�ZC-��T�0�u$��)�b����~���{C����4~��m]������ї_�O�i}.��-H�b��IQ�4*U���@�&:��E�&��Ύe�����#��J��|�j8)Qa��k1�����\�s���V��h�I���J�fXU:��.�φ=�=h�;��u"iu��p�]?E���Sg��`D��>���e�U���>�f���SK����NR]��1WA)dс�J�SV��
ml+s%M�
酪\���\����˒�]��%30�v��gdi�I�a��S\#�ߟ�$�%W��؂�����B��H�1F��Uw�5�m�G�e��OB \��{а�A:L���a@�*�3��7i6�Fj��}�*"��4ͅVx?Oo�5-�IsA��<-f}c���3�������G��,�u�}�BYd^�\	z^�hKX���u��)�Ċ�Ȟ~Oc&�N9��@'��u��2$��$>ek��zv���]*�v�� ��ߗ!�FΌ=f���q��)L��t!�)4�d-��_H��B~�;B��DC,��F'H@N��&�z��%ə$�^YJ��^�EEcr��V�%�{����n��x��Mlᚒ���������\~�={ްd-5-7q�)�O=�#�$�Ă�>R����y럃N�)�0�m,�����(�����ۦ���u�&s}�hl��˯y�$�%����s��c
mKW�K1̮��J蕘H}-7�'���#h�ɠ� ��, ������\������9���ɤb���*�&}6�5s�=���ZܚL\<U���<²{��R��Kbp���O��m���>eQ�+$��b\T��Ec=k�˭hxڀ|�(�q��E�3�&�\�n;uNV`�B�~�3wDA�x��E��+[%�n |�^��'��y��ނ��`�`C�5��{��57���i�>\Uj>��*�����+��o�y�����sΗM�$o�!���t[�r���i�S��gU)�શ��Ʌ�J��#1��$�%�����5�7������$�G��,���Nrg���D�ҸB_h�0_�BuEFD+=G��HgK�WfCQ=#��7f��c��g����J4T�����o�A}Ԯ��������D���h��%$�2�����B�E%
�� �>T�G��S��}�u���%��l`��<.���xf"uKœÕ�lES���N�����L�OHY;�κ�%��������,In�b��5D��P�pE����J����GBBj��<4Z��D�^_�xn��]���ч� ~E���K�~���J��%Z~+K���w�Qvɐᖈ_�ʻ�e`y�����J�C�K�>|N�e�z�C9AZ�^F=Nsl��ž�[c�~�s?Gf�Q�݉�(W�%�@F'?��b��`L���.�f���#ի.�b&ҋ$�ju�¢n ~�T2+ӿ�T ��aD�O����h�^D�=��27m�?����϶m4z�P��<"�s��r����ѻ���ޕ<U46���N(���6�*TA��7���賡�Y155�gC���D���}p�v�S(¼W"%�~�� >@9��	��o�[q��(x�>j��$��_��l?��>wR!3OǬ��Wb�N�EA ��PX{㡅>��-���c<7����A��_#�D����!m��AF2h�
ios@;潅�>��T2q0��o�I�ao���HO������G�U��ڮ�:�i|>��a�x�
�s���4+��:ͨ͡�Yhᖢ��(j�Ve)�x�Ⱦ�q�ɪ��hkm�NRZ������	)j�_��:�C6̦�qT)A=�Ĥ�jGj^��h$�DT��$��y�����/�ی{���|���,b�'�hmoи��1nj�o���)E�&lɓ���8O��f#B'���ջP��ɇL[��ަ���x*G���� ���;��2��ܟe��vYy	(��~�U:�5�fs��Bu1K�u�]%U��ܘ$:�I_A3	����.�t����멭�5��j�r�����K�@�	XD�A�&䉚��<)�|4Yn�P��>��:s;}	7���@����>H���Q��MS6d��d�2v���OS&p%4M1M��!��2����F��7���a�'1�oVG���%���v����§F�[��B�̢V��Wst$��{��a�dt+ۗ�n�Vbķ)y��E��i5'�\-wz
K����Ks�M���x#Ud	����:����3D�$����NBk;?�]����<�(�]��J}W�X^XJ �e��.��JO#����^,f����f�8=���/�)>�b)�6�>���2")2q
ϡ{��ɔ�_|�c����YMy��]`}wVVU"�MO�:���D���GQ<��$"?�su��b~�~/s�Ǟ����+�m���y��������z�z���.,[t�6��.P7R� ul=R�#�Uo#�6G1�^�v�\hW9ߓ�N��T��6
��RL8���"�����a��;My^#�F���<_Ƽ4��T��.�$?S�ш�4:�؊���`�9�x�G؈��#��^�M��P"L��Ɩ"�ӷ�P��o֓y^z��GIޙk����p�}R�(�̹����}���]��;�M�ЍA~����7�"��C(�_:�e��/T�=����Y�]@*?�XZ��UÎ��Ck#j*r�~%^�j�2�&k���<���}GMkɪ7"zM0'�����ݨ����U-���$�\���<@�|N�+Z��=�>[Ǔ8xy,����� Î�	�g�5��U�v	�n�X�Q�F�Dƣ�)��{2b�Ȍ	�5�2� (n����)gѪ.%K�w�d�5�~������jppd	�v����j���R���n���ƛV����6���T(bV:�U�
QŔ�$Ӡ�P�ܩ.6>����j�TΫ�$�c�Kw�se"0PذJ���A�ut�r��C ���>�h`3-wD�fOk)�9�t���*��V큄�]j��}i/[����'�~W�@�o�e�4I���6�I��SS�b� .�/��Z`GW��P��7O�vc�{m%�,���΄���.��GMp�(i��S|�=u8��v=�j
Cw�@68kb�����B�	$�Z�;�]��[g ��<ާ�V`���^�$�����K�O��V�W��f� ��Aӡ:�����k�H*D�L[�^�xP��KJ����.>��Gp�dN	g����ĵ�,�?I� �1jY�@��
pN	��j5BԀ2�?�@�&���V��Kޜ����o�]߾��EEv������4�D�P�r
�eEh���� �bñD�t�ӌձ:: �/�}vP
���2��1��p �1Q��N,�c�M�JDx/1�����O���-'!p��W"�ڤ���Ӻ�:jXd�0P.�����O�8��A�H;h���m7%e����b̊��Af�P�XV�����0XX7�i�Z���;:�Owtr�����`��g�Rk�&�3�t�J��>*s�ic����$K3��@�h"P�̱a�"�ZR��b���*(�3�B���B3���lD�O,���U+��X��׳�F4c�=A��_�V���_b�m�����,�
I�s�@���(Ër����Ш����$�>W����!(�&��1�������3߳�7t"zL��N���\��.-��k��R�N��1r��c���`4{:�aOS=�*�r�78>�Mѻ���˿m�l�"����_e���<�BF,��gv�:Q";��:��2]~rY���}N��S���c���8�����y�?R��Dm�-ص7��2�3|˜�L�A��CV�V#��5y�ֱ$�n���Լ+^V�͙�|@�?O+i+6��Y\���ꀝ�Xc`�p���B������Ŷ%�W�mu(�İ_-�t3Bu��
�Bd]�����o��HT_qN�j��[fk�8�9�hKw��.lޫA�/�`E���@�`_��M���19�3�v�!�~��+�������Jl��͓{����9:"
)BȄ�y�,s	1���^z�A�SB�gЊ�����17h����D8~-@-Vd���a�/R����_3.��r�\˔I�Z�Z�����E} b���U��w$�B���Ƨ����$�#����Hz�gL�a����>/�n��Y)2n�)�`wF:��:yz`��M�G[���h��WPϠ�t�H��c��rM(K:��F����khW�=u�#�k�+!	�ȧ,f�XR��	L-B�#m�-B�ؓ��7�$�ګ?]��P�0 ��8�B8����3\2v����x���û!��*����c�5lx��`�_�f���-����F'��b�^�y�6���� X�k��fW��9��`d������6��x�V�IJ���JrA0�Y`!4n�;qZ��=8ܥ%^�S)#M�yY�{߸n�8(jm�YW����/?�	�p�p#J �
�	����4N+�ꖀ��\*ϊE�O��TT�M\- *�F���HW���%f�N:( W
ϊ�?k� �2R0o�&*�i�g6����\�->���<6���
�z/��k�	qX�Tk�U�,'��
(�t;�,\W��G>5�S�SyQI���h��$��!�Tn�i��x��k]��%{��o�?^RE�i�񫭺=X`�C�0" 9RZ̻p_���Q�2�f|�-S̉���jI[I���+3%'
 � �{UTf;�T��zjL���'�J��-������S ��'Q1PT}*��~��6�⸤�HG�F�^�MV=�~Wn�˶��)�2�ҷ5��1�o��~�a�v<!�~"W������Ǜ��	�+ڈWﱻ�Z,���4�N�m��]��N���������%���� 㞌��"-��� Tl6�P��7��)Q		���ٵ���/�g��Q7�[��h Ё᱕IUG*�}<�󌙘���S,��ĝv_KꈵRX�+�W���� ��
`�Dm��Jp{�X��d�|���d1'����"��M�w�旸b�D�u�0煝��p�ݿz������!o���0�҃�lZLq��}>(	��a�{���Q�P�+od����R���Q����'])�z��Â���a����p��+�n`��r��vH�U�$�s����9��k)Gjc���5E����z�.���%P��6�mFIY���
��P0E�7�V��:[ �$K���]8!ܚ�V���~��UJ�,�sS1�;��d\s�bc��k��uyH@���t��2EC�B�i�*��)�IH�Q�����_��@��ͧE8$��T���E_	�x�?�\�̛A��N�mJ�V�-ͬk �< 5��>�R���4��0VsMtda��]K-�Z�$������r�#OP�
�Yj�/EV���U��;���Sl�&	Jq�G� y+�fX	�$jk+���EPPk�Gy�}����¤�\kޙns����Ѵ�|ɥ�*�� 7�9��G2�:�}e�К$Ĝ��V�F�
?⬙��=m 	�|T��$9�G�As჎�^����eA\�_�H�uQ�����D����Zq�5��)Wr��s難a�H���葂rE�ȟ���r���S
O�a��|����J����`���Y���ϥ6&%xo���C'Ԅ`�,�E.�O������u�(�Mt�2+�Wxd �pK(� ���G�n��u�7��o�h�E�J�_�ak��_"�-���-�Z�$p�|3�%��s���q��N�6���9l�i7�#���F�V>�R]��6����V��m`��zJ����W+��]�B6�&�$�)�/�y���͠ȄP��Fl>l5�CS��PK�uG��-=Z��H���وW40t��ԭC��ہqM��ȡ�9'��-q�K$�������T���w����]T��=��z��
��L�C����n��I�J�Sh�8@hU&�/�U��[%��E0�tXcU�y�/L�6<軮O��O��f�Tw���ߕ�k0Q-��G�f���A�m��+���@�qFX��0fiw-)ȱ�32�����E�ַ
$�� %�OAb�c���Ķ=���T| 3�@�)�
����:6��J�~,O�c�2�q	)v��?mq¿���3#�3
���S^(��b���bq�D����Rǘ�MCV��V�q���Z8vM���m;lELK���s�!+����+͔�j�pj�C���H3�i2��k�X���͹�Sɾ,��z��gS0�U����y�lR��������(���ڮ�/�5P�mA|�^�Xv�R�߸X�4�fb{���/�9��� �:��7~���xv�uՂ(�Jl>�5h+��\�з+=c�QӍ[��q�[5���4jl�ψ,)\s�Ź �H�Y	���=q��!{�Y#I���v��(�C&ծ��6үw[�u��AWZ`p$�|�G��y�b�qS�D63ſN�q w�hQ	>3b�|�28�� 8[⎭�|�{G�n��q�0�W����c�['9�s�� ������ϭ0��C�d�����%�]Mi�g$W�A,��3\ߤU6 ����a��S�K�>���k<=����dnn�O,m\�tD�L����BI�Pr-\�=Eo	�̌2��g�qc"59,G���*Y��qʚ��1,[�0z�ؚ�2R�cprǳ���$Zh�CF5xΚ7N$K���� ��՝�&�a�R�-0X#`��(1��؄ݨ��O�m�_l��'��Ϙ�G��;	2Q�`�n�RG`��hN��X&����-q��������xu�Z���fJk������$�z�)�BB~�4#,ݧ��c�lT�8B�*�-��斩B)�!I�)5c��D��q�|�+�6�	H�+Y��S�/%� �T�H��UBb	��^��E)X��|4�!�t�4O�pɃ0��8\�օd)yV��t���9i}��}r��Ӓ"bRt0����dH��`�Y��ȧғ��%=BS����ҡd���;55�Ν+w�d��=���}�����m�nqBIV!�*s�)��C�����뒔�yq�v:|^�Hk��\|�����~ի���	�T�D�P��l>2�@nn��i�� ��P�z-u�fQMF�K.�aH�N��݇�Q]2?İ����2� as��4�zBlc[�++b�PŖ�Y����z�XVzc����q�_�&#c?�k�W�%J�6
�O�R(l��EEP��UY���>��� hJ��q�@�����ɱ����R}�v�L��҉_���{���o��@JLjU�PG�< Q[h�H*9h\�=ͽ��=)�Ep�!��� �8{T�E	� d�	ڲ��UI�u),�J�yW$��{>U��y/J;Q��TZLx��"�O\_�3��,5�2!�t�,�bޑ��f��%_��K;�	w��m[���iۘw:����J����.��U��j�`���#	��W]gB~���y8�>>	Kh�A����d�,?�#e}z���@��8e�%�}��[ƭ����n�8F��g�p=�Ṉ	 �k81e�T�2^�Wz](��zA��'XB:5N=:�i��vg[���τ@���+/ݢ�/�|��7�#�.���R3�}�ঊ�؋�\�V�Em���.&����
�� �̟9t�o`��uW�\B��R?�|��o�����68�m_����̙?��b}��''"rˮ�A�#1�C){|wɪ݋���ڵsa�qJ��mD1�<��D�0�O�q�5�5R��F�>5ܞM��n����z�2o�j"�ۅt#�h��e��;�w�L��R���ǛV}�� �T�O�H��I���������l��6��̅Hf�`;>6�!���Q�G�m��3��@�Y����@4��#܋i
�C�q�RR����6	����X'����n�v%u��0��dץ,�/t�Ky��FS�\ٱQgW"��xoͭ�Zw��F�4���h.Rƛ5��e�-B������~K+ޚ����7�Y����2D ]����<ʹ�{�����	NHTj��6�XW� �(9;�I�F��pC�NX/eD24[DJ��"7*�������7f�ȑi���'�QP�B����[����;g鏣+�,�x�Vl��o�;N`�a��$ �rp�[zĤ��hv�`�,�ſ٥�떣'�͆8���q�IQ��6��OI�y,�@��$����O*�nz)U� �w�7�)���.�߿��~I�n��v�9�ռA�ʩ��nW#�X�x\�#_ǈ��S|�g���O����!��=��v�ܝ���cIY�h:(0P،|� K�\y5}Jİcl	�P:�*��b+x_iyC��s!=�:E���&I��g!��� p�����Sf`�]�ڑ�<c��Z��=�l��©X����p"^�`�n�W9ߙS6�0������0�%��ЄWRʔج��YtՁ26�Y��%+B6����[��UD�1��Y�K�"��F|�Z9����0�U?6�c\o�sL�c���vN]GBn���忖e����?荮�Hw���㹹(����o�^� 9�S#�s��&p*c�&E碧Opp�T��-D��|�b7��| ��Vr#��� �m�Yt��j+Ӹa��^�kG��~��ͻH��$��,8g���Yo�\�2A��U�u�����{>`���4�}4Bo���m����"�ǑA���H��W�Ś�ƞ��G�|��/�e�+���3�`�q���c֘�hgP��]ܫ�>����o\�SEU���� |��	��1@p9lb[S(Ileh��-���^�Dx,��X���U�5Ukۃdԉ-�D�CDӵ��Kϲ��o����Rsr�]�/��ј��e����9�Ѝe2�ފ#i�/���Pc��ys	Ӂ[��.GhE�����fg*���UK�M���9��V _�"y�)�Y�WF��#2n�'B[�E���3�t��n���+.�8��:�ZDf�����+,m)�� :���F��}��������V~�^K�Xh���FyiM|����$\�hҴ�	i9�M��P�b��4�52�󉅿��l�>���"�K��c׶�r���1gd�S�L����*�����9�P�>�9���Q�6,��G�ҌWt5;��ڳY�#~�s��HUcj�E��JN�JQ���b��?s'������Wx�Hk���kt�Dh��n�K��x�Ɠ"�q��ǰ����X�=�ݿ�����ѝ:�����;�I�>��x-�ገ��P*o�t�a�cTu� ;V�]�É+�����K�m����cPx����J����\�A߰B��C��ٓ�L��V&�t3/�1	��>ˣ&�_�ej��g�<A��::-q�����ʐ��8�ƒ$'_��O�<���tL���J����`��~��[�jg�#��n��j�n��p;ME�Сەb�KR	Ҝ��J������;0�BXLH�J\kh/fZS�����lO���"Q����K�&5?7�9�!B%��p�U���Vr�6�����)����#���F�PS�?"���>]�ۛx5M�؊4���h	��|(6�W������
t��^�5�왊)f�id�WB��{��r�)O��볰e����I_��-{r�I���&s�k�gU��ϤYf$r?*7'{�!r'M��wGP%�I����p1R|��̪��;Ϗ�ӓֺ��eڵ�\�"s�=_s�R3a�t�5�&WzZm)՟x�X�n�2�J-��F���k��W�rm�1%�C9;�,��T�
�)��\�pR���W{��ϩ�D�2���zE3�>�W�����8�2�S����Ȼ[I��Fb����^�����Ԇ0͉�.idy3�®֏~�Y=��#��k�[����Cϼ�=��N`�U������x�
�Z	t���e��?��<�Lx��?h��%��J�n�k��%�͇��˛/����A���ن��a��C�����7�0g��o*P����mL�<Ҍ1Wa:��܀RX�����f�8Z����5Z%���N�|�������8	o)輨�� �	���?�Ҝ ;�����o�~~*r���������ڄ�L@'�Sq�=K�?'��mJ��r	YG�?�r6�˙�\�ن9C�Ba����oT��f������ ��e��ל����0k>���Š�_畂z��
r\!T�^r,�l�|5Q$�]W�. gH����$m�L�G&���qk��+⁘�W����%�l��+�F�3)v��F(�d�E���ܕM�h�`	r�Z|S	��.q��c#h/���V�$�O���Ne�75e�gy�aK���5a\�6N5^ߠ�ͨ�g5
�#vj	��8Yʎo��x�xS���{L_��K�Eҙ�-�ET�17狑.c��6�&u��677�ҋ���kS�^���4E)��R��:�o���yP{��M�	C�Ix�0���S�� ��k�9�D��cUUτ�1�ƽ��V�6����DϛxA"A�2 �-�G'}רW��VH��$�-!!��ᕓQD�d��c[`�3`��ʹfby��S9�E�YL6�8*��9X��`,�wc ��Ƥ�'{+����g�x���|#��ٵ��E��2I�� ?�d��d?��`��TZ�
�4ca@����y��2�W*r��>��7���`A�����S5w�������p�����J����*���U�XY��`U���k���z���i��Χ0����j�½{I+L��/_��ز�1na@mP�x~�6~���
k$S������ςi��g!>j����qY�q� �����|�Co���8B�8ސ��j�:����DB��.g�-{{(f��&��P�aR6]���MEk!�ʳ�]=��t>�q��ў@�2��m����x��>��W�Ň��\�(�i�iƛbU�$ͥc�M�-b�:�c���Q�n@��G$&����d/�d��v������|i05��BJP0�V)�yύ%Jt7�$v#���&�]�$m��*�78�܎�z�>�h|0�	��%�̥��D�U����~�IX��������AΑ�"i�D��P\���fAk\j܅ݭ���Z����Ƞ���jW�%-^�&�ۥ������,M�.���)���'�z��aL����<X�b�; �v�~�`�z�O��3�`�D�^��$��C��8�\MHؚ`�ϛ</</</<P��~�O�W)�[e6'��z3L��7�����>��d8���]�B>�{��MU����pڧ<�@�}��[�
qY�T"ѧ8���(��+U[}H�ΰ�Y�(�[�4y�^zU�A���6�� �^�2���8ŗ 絨6gD�[�����;B�m*�m�$���%o���� NɌ�q��ầu�a��݃]�5�J@#-7S�	)����ώ�b�u:����=��?mQ������y^>5�Ox/~FvYF�+�1ޏ�
K�IdC��$�rFP�w`6��M��x�2���v�8�l���wp��\.k]'7�T�q�r:��JR�OZ3�l �&�����F7���c��"a�|S��s1[���~e��!�?!T�S�6/Sf!5����Dn���䄭"р���D�~�S�����
x� ����4�βW���f,9E��^0I��й�)	�̓��le��8��$g�:I��£�3��Y���Ihc"�܀9��z�:#!���=��m�~�
��_�K���O�26Űon�c�]{��қ;g��m��U9r��Gݦ�]'�]�.�S�An��Ճ�̌�5@nB(Z�X���]Uǩ�j��^ �4Ng,���/���#h�Fdg��d�?�S�!��N�T�v`[h��$�d,�cHjmd�kͥɪ��M|D����	d~@?iY5����Yb�y=�*���n�����&�u3}n�;0<�E�l2Y�6M,;��Og�1�LT,���)k�U��Ad)n��@������z��bDz�^QC+��*��J�Ga~p��Ѝ�p�z�=(�І�<ӊ%W��+N���kk�R��s��KD�r��D^�}�I�i��ѫ�CVh�멏��bXM���q��8�^���.G�I�i*J��Edu�$�>&A����d���H=����Y��RR���� ��-`�'���+�+���$�s����V��J6R��1�t�H�1�3�B)��F���Y��7�A��Z"$;v�B�[�}�vJp���SC�-w2d˻Ě�.������3�_̚����>q�g�-6�m�����H��뢜$H>0zSk(M%���H���i lt�<x%��w,�=��Ν��@&��Z�-x>���d	&�����/p5���+dN?>0quYN��5}��t��0��Y�XL;R�	��VPG���n��X�P-�3�6x�~����L�#�N��k0�wn������Y��Q��B��[SF5M��=���ލ��{�F9� �ݍN���9ۼ�0�G�x{�F��Jt����!\8�K�G���7h����l[�T���N�� ��١[�-ϋ�'I���셲������d|�DT�E�>�=�W�s<yZW=I��ftqc���	h}`o6�?��������虦R*��:%�"T|K�n�0��������͈����Qt䓦1,>~b��f�߰�v��=�?��Wp�ۑ�p n��'�e���ŕ������������[u�@���z�����xޓ���=x������ŕ���v��߈�`T��20�{�k��
|�KѼoR��'��[�]�F�*������W{�J6
�E.7��E�TOɏJ�J���QU��l��68]��z03
�W��x�t"�:Z�@CT�8vFC����z�] iB��y�e�$���	�1��+�FHh���tNRJ?�7b��+�T��T�#��i.u���ڴ��14���X�0B�ҧ� )���x�X���yVeOyk~�D/ �߷�l��y�@\>�g";P��v�sR�Sª�Ӏ
є�4 uS�;w��};b���GP�^����:�y~�T��h�����=eʪ�BZ����吂WQK�KD��������D�x5���1S���k� !�ku(���j��yd~�0�]Z��q�p>!Rj���y�(� ��n`%��~
(�����l�j�GezKW%� h�N�a�����*\9�]�{EXg%�y|�I�M:W���}W��F�\��/��	�K� L�S~<�^���#bp�<͗�i�4���1]��#b>�V�^fY���?O��1ߢ��F�x�P����7�6}�v7�(^���Y�}�m�ga;����V����z�,nZ�%F8����5�E�8EQ�_\� h�Ĭ,<gPy��W�v��Gd3 `-��cΡ� GA�%w#�2O#S��W˚�����s]�(%VӻS �z���)
j:�o��v���VYP%�AO5NE+�\���:\r}�ST�у�5�@A��7���m^�RH-Ý�7�6����Z���#�E�M*�Y�6|��ڎ����,�)�9)w����MpΦ;�1#�:�q�/���T��7���[x��R.��J��� JZe�~	�VF3xi"��M61�_�M��u��H��J��8P�t���4�>���a�ރ�+< vp�6���N��D�~a�U?#%������?z�@���g�i-t���B��V������&��a_wT:[i�З?T큞T���� ��S�ᦨ�����c��+�(��UT�{?t �߸s���.�MC�D���-W�tW� �#���7�6i:��K�V����i��gE�.dX�|f��6��v�������M�+�j�%jm�6�lR)U���T�j�i�]�k���iq��-%C]+��I�1ez���СM��Vɰ�:�5�8��4�~���qf�v�~����[�Eۤ	�ݷBx���g�A-�S4����v��Ch�B��H��)���ىD��\{��nl�~Y�.�*�����)��4g%�B�J�Aڮ�(���9��t�+�����PU�խ�,�oԪF���N~x�݁;DP�T̯N�533[��Λ�3�ck��k��^)��h�1nf'Ʉ�W�㝣*�� ���i�]9�'9�G��i�K�A�GUo%�#�������O�.L;��q�p�P�G�#��*냻Џ揮��;�������;��Ji�g=`���u�{ʏĢ뭑v%�p��j3	�ˠh��|�:a��2��m��!�.fp&4�7\:n��gFWg�>�W�,�I���_��9@�43��(�D%�w��U��6�<��h=d�o�fMVh����A�Y�`0� x��)T2����^��*��<��U�=)���:��n.Z���ԋt<��i��篓N܂�"�3���&�e9��V����!�Pw�Q�B��$(Q/_�_����m��r�N���/;t�S��_*�G9�o���U��.��qL�Y�sY]
��|(�@��FS7;�2:WYH�o�D\qF�2�)a�Q�7��Wܢ �77,��l��rf���v�Mp��Uא66������b���������e2M�0�Ng YE/����q�f�_����@�a3w:1vnA3E���=F�c�}�<P������)��&[o�"���(��b�S7�d�륳�
����<
�P�5�9O�c�>-=-/�|�@�����R����n�_^��*r�f�+UL�\��1	㴂�P�u}��q�'�G	�P�Z1ߠ�NI^R+{�[�����8���\�o���5P��,��^Q�����n�y>, �XQ�Y���m0��F!���Ef�J�Y��)f�Q����E9�b,hV��ɤ
ͺ�o���h�@�dt����p5���8?�GEr�[�Ĕ�ځ�c� 0 �[A��X�Ɋ�ĭG��6��J����v�0�H�����xH�b��o\��=:E��'jЬ'�O\��ja,V����=�~$/���-E?f��"�H}w7m�ߪ�y��:9zU���He����r�>L���.2��|��ה�:L��E*X��(:��1\Z�rK��{[bJ��8C�	�)qv���gw�J���<aj�3���ۅ &cT�vuo_�K���:�E��Z��5D0*(�G�d���=N�T�XDGׅ��V@ƿ��R��*i�S�:�i�������D�>U�׌4��$k5/�`��L��IqU-=Re��H���[dPȪ �D7�<��r)>�C���y�1��)i�Fm������Nη�D����u��-�'��˥k�e��r)v��琌׵��"vO/�-��N�6yɡ��z6���֦ �Eyh$]��:��iJ�*p�K^;p�I����Z��bT`���G@�U0�"*�].�����TH��L�ak� ��x����>���E�<o��R��_ ��cL��#��.�3�8�\Wۧ���W���&��-��;��X�Y~¾�̰f�ύC�_�4���
�;.4�����mh[��S?]v��.�o��׳8��d�Y���@Z�����'���T��(�zW�\G�ITPuxQϧG�٪��=���%`���g���vi/4����.G����� �*a�8~���˚����t��)D*}���9
Y��i)9p��ɧ����N�L�M/ 0���9�� `��ޭ�Cuݬ}���!\���Ѩ��v�h�(wkr��u#��:_���"�;?���S)�vX�5{)S����?1�k��цkx�xq��}�KX�\?pv�c���Fe�4���kq�;N���� ^J4��*{���+��X�M��a��冄$cbr㒚��Wv�������;�S>	�������4x��-0���)�0_��uϦRPp�<��.7�sl�c%M;����#����4TG�����7��9�w�J�����	�d�p��M"���gM���H�O+�S���+fS㭩Q[X�=�A+i��b%�,̮tm��;3KV?n��[�ʇ"��Hׯzi�[�&@��Q%�$��	�t��u{q��$�}�#6��r7 ����T��Ou��S�
D�VG:*�ˤ���B%^�.r�����˙�:k���:��c'�iIo�3��f������+ޱVut3�?�^��Sc�V���P5������-'�i��߱Y�"A�t�����ڞp7��B�D��xE{RE��`��:�<�ư��0y�*� ���{.����|?�C0������)֐�R]�Uڿ4��~isB ����6	1�hЯ����hB�R/�4a���$|�t��[��OҘY|��5_�,l"T�B�C_N[8˗�&e�5BkyM�Nh����կd-6���hR�K���t�q�>��E2|����lM�\�P��E���l4�JbZ�7l�\8(o3T�'�e�L�H����0X����|"*4�$�I)�範H�ֳ6'�y|�P̡�
����>-��<,�-�f|!�_x�[�Le9*�\\�u{��A"��Gt�-P��SHZơ���eL�<�C�d���c6����h��v�϶�A��aD�=!<��=��YL� �:�0�I�E[L�/w����;�>��h8n��v7~��L?��z����(��Q���݇ܙ����D&P<�����a�:�'�'�#�09���pZ�&uڄȕVnY6��7C�L�/cY�І�B׫�Y��d��ǟ{si�����`N`$q�N�ǲ׫I0������a5�����~#4���B�!\�)�nô�56��"�@��25w��v���Rv�,kUS������%�"�͗ڍ�`�;���q<<,(�W1W�M���Ҟ�"
=a��T����� Xkүe�V/� ��f�T��m����&�S����)}h���T*t�6���9�o",;qծ���rn��BQ��6�}���]��e[*�}C�ͷE��6�dEy�p�=���n� �H�$3�.��F����r���E;l����R>�v���S� ���|tt��S����"�,��/�w��i�}T�՟����Ň�v&f��h�s�*�^$�7-�u���ef��������f) 4 e�a�ًM�'.��ǣo'h+K�����w�	�1�F��D��?�I��"*�a�� ǈ5�3�_��^�iq��[S�uCTx�ʌ�Q�R��L&np���E���
*��+h����>��<�	(ee��k 멠u��2j��a�&�vl�Q�s8oh�d�J�;�r��g��%mP��h3��'CN�p}����;�ji���B����uf�sH�>�i-�6�[���?�k���0����^B��൜�A:�U�"*�ݤA ڭ�������2@�oEr�+�C菋�fgOX��2څ���&V�O�ģ�U�#ԛ��5mo��1I�FRF���%-� R|�U��+�)�4�_�D�%���Q�s;�d3��l(�j�8G���g�9�%h�W����IN��o$_!b�����z��iq�ԃF,���S�aAd�H�nڄ+�d�]n����Y��A���(����76�V����pĹu����_�˜�d��}���~^W�j<
Hy�#�0��A_6ɭ�@�j
,r�R$�Pv�_КK�!�*�ށ�R~�'�3�x�C �qsT3hV
C�mA�/*Fw#�$�"8-��$�1zS�y��{];���1 C����a=���՘�X����XZ�e:�2cOq�Pi��|�I熭��e��|����1,~�L�Y�;8-����)�$m$��얳�����u�d�8�א�y84��y8 ��~	\��"	�X#��X��c�� ���1����4���3o?���a�V�M:��'�Di�Ca��Cآ��M��JBZ( ��*׮�ڮ�v��9������3���*�!�R?�+ i{ T�W��$h4!��ʎ�cŏ���^�Y<����!�"�E�՚%�W���d+�<�r�_2*%���� �N�t��"X3
-�/*��E�,>���&�1�k�='Ǳi�-�Sg>�I`����H�@��)+������dZ�7�Ӡs}{���2�K��0��%y4��U���<��Y�,v�W_m}��.�XR���A���H1jU�c�lL�����n]k��e)��;�/�NQJ���;���h��DS���� �!�&;��Y=� K� ��2����7�e�x�eժ�l3#Zu&�^�"
?nr`q�.��ǭR�Q������~�e��%M�7����O�^b��j���yR Т��@�K6B���*#35H�eG8��@�z���ٹ�B��<�X-�H$�+��?�ښK�R����_�"j��t�D��$%��C9{���L��8��BL~d*b���^ &Qb�	�pX�䙓=W�_�lD򽑶A��ނ�C�� s{f�
��p�C*u��t��Aw�RŁ���˛9�C?P~P`:=j�A��k���핇���P�vj2D�]�vd�k��tn��X��d�̯�.���>Jij-�H�m���D� �@���.L�S=��~�#��}��e1������T�F�w�P��e���{�q8y�K�͊�-���eK���6,�L����r�r�x��`*������W��o�$;���)�����ϲ�L�<�p�]�I�l4�P
����Yy���V��]��̻��>R%�a'���]����0W4"����8%xζiL��6���5oD:�P�9���3�4�k#эE�#X���f6)I���c
�Q�����:c�ŕ��[���$Q e}�^�:�s�{�A����A�ŵ/�k�\c"�� ��u�]c[��$š�'/H/1/JZ"��<�cH2��^�>�1�g�)�˗5D��/c0��2�s��k��͵<.������E��4\o����$��r�UgK��kʈ�d�����U]<��!�������NS�l{����n��|b�9x��Ú���9�/�xp�i�� �RI��|�?$j����ii
/@��^���0=�K�,���[�8�"piԌ�Х5��YzR\�}= �J8�r!vdֿ�5�6��<��%�>��:����JP�D��t���<^z�c������y��
+��o���#>4"r�{��3�����d�4�
.��y��sR�--�;	�Xc�el��}t~�.$�{����T���z�H�L;
��I�5v�l1�1F��#�*<�����m��R����]��^Y>����Uf��Q�G��&L*�* ��ur�lz�Gē.�w~(�d����E���s��1b.H��~!9��c������R�Rc�i��^Ћl��gt���v�g9�1��)iT��B�1��oaڌx_��&�
DV�F^Vg܎ܧu��%���p�2�#���餇�ӛ'C�n��Ѹ��<��5\�R��r,�%���,I&�A���t���RM�U�?�$�S�/���nN� ۮ��$�BV#���6�5����g��t����3�٢(����{٩C��R���$g��B)����.��ݎڡ]g��0��o
��O�Ԫ��ᾭ��ݯ���6^�#�Er��v�3 ���6�	?��Q/1Q������NCx�����#}��D�m G�~#��^EA�Y׮���aj��@�b���i,�6���NU�}��^��i���E����=��#��C1����b35�B��(~�NE+�� þ�g0	*���$s��q>�c����� �5-��Q3�>��i�m�Z�׌�|DJ��|_�� ���g����3�LT&*+:d�20��v����<,��ُ��a���@�T:�rfO\-�V3u�Ui�&���s��y���I6:�iN����^��Z��ٰ�>��~�W�G����p" ew�lշ�IC�kɞ Qz��{�%�%��l�+�|gl���|C���d�,���lo�o>8		�-����ܡ���hk]�X��|-x��!��k~N�v�6A��u~��-.��o녻�5�L,�_���>�܏�c�$N���w�|N_��:+�{Ua�1��g�N��J=���+@:U<�3�s��x�����5;:G�:I��b���������w<�c��n���PtZ��Ɓ��֐ٱ��>@9��i��p�vf��E�.�����l'v�`�W��Ly��Ĥ�k{�Q�f2~*�/�V�oB<XC˞XI&��vH�����[�rَ���3@6��C������� ���y�ث�C��%%���0�xbO��ʖ�}���8�!�Ǣ#�5Ʃ�#J���U��'�G�Hw?\9�Sx�̛��LK�Yqd�I��<\��� ����-�|5�gB�C��:��}���Ǔ"���1H�)������6��gN����Q�@�K�oǚK�=m�➸MPMdOD&�&B��7P��m�������#��7��N8��)����#�=&����,���ڿQ��#�w�}Q�{����p���V���k�(Hxק'�X*�^y��-+eДGBeP�D1'B$G6�0=>e6��dKu���jR�I�T���0� �f`4p5��]�e�KJu�3����)���K4H(`�Ė�3�]�{��ˊ
O{�ƥ�.�9��*+_r&�����G]�Io��3��FTݞl�&����b&\Џ/��R2��kK�����b�hD��I�5�qS���I���S���C�U_w�#�k#ކ���k�?3F�kYm�Y��ˎeXe>���������}���عN�\ҩ�@zs�۰~o�g9T��l5��ϡ{�VK�Ȩ�c��n����vx��WJ0�ḟ����j��6��EY���raR�$O��C���ZL�qIy- �t� [��媍f)*�r�DY�����}�����3<���6}A�y��5t�vd>z(��F�]_�P��j���CiRհ��i�8O۸,�?�D��GK ��c��7*k7qTg�3�ۂ�I@n�3�D�	�A�dk�>��Ô>�D�G ����k���lY؀_�0.�,#�]P37Q�	@MH��ҋ�T*9���*�@����r�D��˂u�K��Y�L����~+@�s�оa�DD^#}�����jSk��'���B.�j�}%�{,�x��� ������V+-�8ݓ�f�F?����Թ?VtD]+���P�$��3�������c��l,��ͤ{d��z�1%; Y ��F_���g�ؿ�8!\�9.����6࿄(x��:9���u�|�4�c�F��V�M�[����q�s���-�V�6����`������Uv�ξ}��~	i��|�1%���W��1EWT����w��2�=����6�D*�	;���sq����5�����.y^�zOc�5qȏuixЅ�s��\ڷ�w^��F$�lEH;P\-�U�b��ȟ�
`Bd(�7	������m3�=���߈&����H�ňԾP��g�>�4��㊎.<���J�.vT��S�KH��Vw^��)ȚX�_&U�Z�g���w�����z�~A"R}���p�5pc���^�_4�y�����\�����\*�jo��t����,�|�/����s>��tĻ ���/<p�2MPN�rao�~:i̙�i+�M�f@0�ޭ���s0$�׋��d�o�[�Bd�.�iڼ_��$F�=Mi0�QP4�F*3�G��d����}#1pR�Ƞ	�Ѿ��n~tN��ݙ~iO�\����J�c�Y�P�<ϡ>�yD���S$��t��/M����͞�[M�6�;=���.Yy�B3 �2����YnL�������0���Щ��QgsP�.��{�<Q��Z�m�h��=�e:�����h6Ң�m����6�ݞ����s���wpˑ�oO9a9%"�%$����x6a��;h�v���Mn�V̝� w���^פ�:/�3�`^z
C ���3�'n�\ƚKQP���=�qR�x�E��4��U�J�'��U��^���yS|�~q��~�b�������͖����l��CP�5-���I�@�Pl �b$��GcrĖ�5�\�)!�F��3��q�|���n��<�@���j�;g�LF�l٨ݬ|3���ۥd&�`�o���0�g[,7e����=������a �	�J2{���4Hc�y{D0)��"�k灑;0���6p)��f��{����)�:�O-x����n�G:��6��P'��	��;-�Fo�U*z�j�o����F�	7��k\�S��G�pp�b�+z�R�A߲M�E��9lϛ+T�g�U�6�%����CZ'��1��6-�:p)L(��#|���*]iX���J΅s�fR�\�P��;2Y���d��LٚT�Y
�SQJ$� O��3�Y��Ko��7�\	�9r��j��1,<�5�q�.�5�Ƌ�7��_��تڤN-�8�R % ���r?��ɼ�n��K����������4�'gc=P��P��yB��yJ�)���I���^���:���.�[6�n~����v�% ��R@1U�48��b�H8z`���$$=*���_A��!e�P�]�]��Ec�h�@�~��E`���3<c$&���"b�����5���>�:d�f������� ߸ɇ!��6��&�T�2�������+�,L�ڸ�3�3$/y����B�╁�������?f'��+d��[�}]B[ހ[��������bD�Q�&8���W�'��}(���x����ᇻbY#��?f?��^'_`D�]���&]���O���LX`�f�vjM�=�j�&��rVT�� ���줥}a�ܘt��-�%6K�)�A7,����5W������z]w�cp�"{��섩"����jo��Q��ODk=�!#�0(q� � ���/��)-3m
��8�jw:j����# Q���[ȡ�y�V��&�Z�t���򞏝Մ�EQK��D��:�QB�a:�X�W�DD:����b=��i��xb*3�۠�FC�v��C��/g���)[O�r ޡ�'fo�)���ٓD�]Q.;�ٺ_ 0t5=x91�Ov?)���j���}�fG�WL��09p���I��bh!y�����-�EW�c=:_�������k4;�`�m��A�aEe�z�!��	ϊ�]%��\5F�QQ��ta�M+�[@x���)X����m۱���aaU'�����0n����(����]�a/��4�"kM�lW�06B㟂N�H'M#�q��Մ!���fG1�
2��;| ��N-K�J��֧hH|��G��}3�|G�L�\�Fk�����`p�mڇ��x�A�Q�̥U��.�g��˿mt�?����8�}2���m��5<% �R�VjS܁�"��;I�[�gw1=j�D	�����O	��;��|-)>�	������Q�����6�0�ѷ����|�ۆ��q��u`�� pe3הk�&_�!]ޒ��s�-�q}�0w�j�!j�d{AJ�\r_�52�P)�a�&Ή�UN$3"O��@)>�EqE�S߭h��+|�Tl8~�I�a���2�.���,O���vZ��<Ꝅ�6�h���QџJ57���3�KOG��T�b?��O��X ���,N�(��������7R]��A�Q,8'��Y3˂��d����r�s|.	�{�4{��x���?��G�����C8����R���b8�`nt���F���W���v�׏H��[��_�������oa���X!S�ڒ�Xς��.N�����2%!��KKo8i��rFZ���k����	����z}/0$p���N�\�!̊��{��G)uk{��3�O�I��eF��e�F:�[� �Uujj%�N�~0]L�����z���3��{�R��C[Y��
���g"\������ǉ�1���
�F������f��:^O�Y9�=�l�\0811������a�f�6���a?xO����l�~
�p_�蓐�(����<�P<��Q����=�͊��:i0U����/=���#͟T�z��]!�󛅲i��{~����h�Z#�LM���t��:�M��s���I���yq	�mX������%+Ӑ� 4�.hew:��}E��J��M�B��� 㲮Wt��w���cM,!&þ�G�C~��h�?,|��"A�XH��cɯ�������x׺�⫸@�f�I�B+�M���pIDdBh�i���:��]���}������.7��t�ynC����\�<���j������ES��C�O޸�¿p0Jɯ���Lv���͟X�N�O�:�O�jo�f�Hآ�f�c�b]ӻu�ѩ��}I�.,���g[�����Ԍ}e.��o)��OVE�z*���}� A�
�Uo����VM�
s���v�}���wm���ֿɷC�)�1RM�bV&\y���K[ʹ���cEP���Z�Mځ���B�Z�����{���� ��b�ԓS �bipw���a�R9�Pl��
��ek*�Y����wPs��G�h����z�h�"9娇K��@�i�g�lg�-���#�E��"� <C<!3� 0#Aab���p	�|��P���	N@����PDY��`��0q��DBh�[�ސh�Ɋ�����
U��Hξ/}�>���� � fg��8����+�E�Ft�h��B!l��������lC���ip�J�M�0؈(���������D3�Oz΁\�����#�G��k,���  d@��{�?>������S�3��k�;�"m�X���o���`�\1�i�*Ijy����皿�~)�̰�W�Է��ϗ3ǲIM,���ǌ�f}^]7W���x΢zKps��R?��c�Y2Z��!�������/����������Qo��\{�	e�b�q��c��*L�b�F\w�@�VU��J$]<{f������h���,FL�X��`��A�iv �I�H,Q��4g��߸9����*
m�.K�Dh�&0t���ijj_U/.e_LZ�O%���fb^Ly��������iO-�L�wU�䅤�`e�+/!/�ݽ�L��v��Dy��y��&ҳ5��xG$�^E���J	0[,˔��	�y�(�6�~��>��$��ٟ\�|4$��!����C,��=ݠP�����̒Pzvh��qo7�*�R*rx��C��}#�n��+C���b����h*K$ޙ/;���� +�8��j>��zpʇ?�xt�(���J�H�5��/�$��3�W�|��Z�e���7�/�tZ��n݊˕��u)��CT`m� �t�f���@E�CO
��yfb�`��l�Y�|gT�Hnۑlk�Gan�o%Ҷ]����w���?L������+��V�d[���	}��t/�e��%lS�����ݖ�Z�m���?j��hZ �®�Y���X����[
��|өH���(���Z!w ������$��1�����hS'o�uf���؋�8'9P�R ��*����i=�y��H*;j.V"��������X��}����_�U��d��nb�gE�w{4
��	���0���|I5�\�t�='JXC,����2_�34��w�����K:Nu�*f�}�u��tP\;x��ܾ<%n ��c��?8H`��L��+,�)�:o�s-���%'��K6�S\�L4�?�� ��ўi�)���p�elA��/�D�G���r��H�V�=�YFXl�h�8�1�G�CŇp�v����!��摯_Ym�82����[�C[�ôw���C�
�����$
9kC�@�l���T�݈�ؽ1���|G��h�6����6�޵�t�~��;�8F۲/`3w���]�NXe�|G��`E��Y�bFb�j�.(��?�;'�kEr�(J����Li�������
KT<�+�V�������ʙ`Ɩ���01���w敒�Y�{��8{��0
��l�}%8η+�6��`h%�B3X�����n{^��#��,f@ա�BG�������G��� Vt;�#;U���s+���16�d~5�z:+:��9Z��܉Z4%fߠd�b67�}�R��6Y�ՕY篣���f���n�X�H7c���9�|�ڸ^�X�u���M�	�翰�w{�����1�ؓ��*�f/5��z*IL��n2@�4`U��M�����L{����)��b����4hrWma�V��u'1O���r���Wk�5�5��qB���'�\�l6�.}.{�����7g�2��T��<U�'��y=ۦI�C�Q��#Ƭt	�U`�N<��uK����7�9��G���p�	P�<�Ģ��(8�Svydڶ�M�s4��S�$�B?�.�)�b�H����)��:���af��0AbAr�z��f3��LSzi��Y�A��h��tf��~]��������B���;׆0Eo��ir7��'ցzʼ,��g���z��Ԥ|x/�À""�l$���:�t�v���)z&r���ia�bJ����9Jm��=�ҳ���8�ot�������qH�N�����(4���H4آ[��~�?���֝CyH���/�+�񄘪P��`�I�٬�e�7�0�F9f�l{�ی������_U��^C����@��t-�s���J:�RS��`�X)���M
��B��i~�ZI�M��Q�̣����6�ܹ�))�<�9�@���\�~�]��]
�	M�VU%[P�:_эНe���:�($��S|�r��y�0;��f�e��P�P���2׸=D3��+?�,3e�ϗ�" �ɘ�:+�Ǧu��:��Z�U���	�`��y��'������V���|�-C��;=VD��?Z=^����QL��LU���REe*u������Hi�l��;J�%�NG�
#4�yO�����.�~�Er�0cD~c�#n�[ &|��0���g���I�rH�1���S\��mQ�r�gjK93C��&�.h�(���RՑ��ˠ��8v׼�a>r${�&B�O�AיZ�pr�)Bz�I�q�*��=\��8��zD�0�3#j�!$��S1�K.�[�sL�-�!1�U��=�����8�dp*�軴���*�TK:���s������/^,_��y�տ5K�;z�C���_�a��b:i�C�7����%�3+�V�T�yu�4dW>`�A%Y��H�4�)�.���p����-|��r���7 g�ui����	q��Z:d+���X}gM���Z%�i>/*�\�s�I�Z�E#�fA�g�ۥ+�3K���b3'g¦m>�8g�SiK<0���M���L�/2p~����Qo!ԨYb����������gte����6�0���E����� ��2��X"J�0�<�R�m����1���Z4��d��Z�aT���Q"��#s(v�K�T��qmMi,��{M��4JD	3 ��Ƌ���XQsm|�r"�u᪰��6��4�|�E�fX��.k�;��Z��e9����g��e<��.��ƣS9 ?d�۝p�v�=���}��k���2㨲£T�����*��z�Ǘ��e�k�brm5E�g٥>@�OG�^@��ϲ���!?$���'k�Ph$�4bÐj�eq飡�)j�B��3�=��E�Dr��CŹ^��� �(��l�xYz7�Q�a�;YS6��������5�Tj�.��f��A�Yt�����;���������Ў�7c��[P�kL6����2h�W���Ʋal�#�FZm���	�&c��6m�vJUh�j`�-��(�poR���A���Ms�O�h�ӻ�r7��||�>��	�+�	i�mO�ͦC7�����k!:Ҁ�6�ݞc�*/�pHfi�R�b�xX��gtE|�y����T�5���ZS"탨��<3��|v�Pm����Zc�C��n���n���H�!&X1�85�4�:���d4�N/�Y	�}k�K ��P�'߭	����h��*/���O���ﱍ\�=4U�h4����>��f��ۅK�&*�DE͉�H�1B�S�����;�������N.u�(�c�}�Q���y�&uW��<�9 ��H�Qi��3P"s�f����igQ�s����ĵ���+0��s�B�/�2G�U=0k��?r/kl�~
����%E�(㜎�S�+|�zD�Q�;�&(Q�c�Y�P����n�bIN�(�����PM�1��u����c��^	^̛�
���Bĸ��(D�LS�?$�����1ays�lcT嘋�~<@�z���n𫣵���A��D���G��Q�:�?�l��y�j�K���H�L��'1!W/O��բnA�=���I*/��+.s���cx�f����� ��I��/�-��x�x)�=��|mҨ��+d����7�fS�#٥���ݰ��uA5�����VW�.��X��q�1H�4�<iO����
U������,�W�-b�b�k�@
s�\:`|�tQ����:��%:��(���J'�$���*h>��!�o�i8�$�E�p=�ͧ��v�����w�V�#=���,�y����.��?yc����l�S��r뜁�Yd���(�.� �	��9����r[P��X	:$��{`�;�-���y�����(pt茈�@�Z��ݥC�!V�<m;?^Z �;�>���#���Z'���ˑ���w7��lY�S8k�;��X�]����� +H���8f4�I��7�G���Z,S���.�Ũ��=S��&4�/B�B��kHx/,m��S/&}ٍLm챓�z���W�P��,	[�'��m�5�Oyc�ˉ'p��Z΋u���`6�՟W:8�	��yg+|�:w�!$�O��WTb�ѲuK�#Ev��i�wt�Ԕ�q߮�E���:vA�дD"_:��aL��QD�ph�뼏��|�̟�^V���,���'ͨ�����12m�hH�6�����1H��h�Z��`�L��o�թ�`����Y0�r��{�b��t1A�N���'gLgL�$�ґM;���0!�~��̥!���?u�Z���li�I�n����Ï䪜NBhWU���t2C��N��ۙO��?4��ଉ�}�W�;�!#�Hֳ���JN��G�3�H��r��.�a��=�4@�*2�	
|�Ř:dH�΅�	kֺ�x�­r�E}J�Evn��2:T����E�`���q{�GG�1([��)U�[`E����r0�U����T%����*U�hύ����i`)�oA�B�^�W�"cikҜ�83v����;Dg�y�V�q����%��4[�
Q�h��Mp��u�!N_���Z)@`��R�O9$>���;I�p�P�Xm|�tQg�i����KK
. ޭ�k�'��]Y`��h�7��w^9�R1��b������s�A[���u=%x��a?Cq�8�|��@�"��?Q�Ɖ�,������N#Q/����7�7��c�����Nz\dl�d;�m}��cz���S� d&i�2�5�:V���r�B�+�r�C�mu���h����g��$�	(AO1������
��oD>[������[ܜ��1ӆ)��;Rq�f�=V����iSk��5�@�5,�	�KݑFz1�S�G����\,θ��;-�\�ъk�$l�aVz��g�	2��"|��2!���o��w���>$vL�B:LT23Α0lD2�FQ�+戻���M��ꡩ�)�X�O�zD�O�G-������ͽ���S�s�Г��â�����W�	�ޖd����ϩ(M s#�V�Ӄ�J�v4Kzz>�:GF������6n�c?����iCez`��z<��3��S�ޒ�⊎V+����\?��s�kB+1��Љ@ܸ�M�A�l����AoH:u/�F/��C��z:c�\Y�V�O`�̊Ot��Tҵ���h;��˽��Nz�����w_����Ճ�������s�F��0�0�=�#K�NU�ǮVl��� �;����ufZ�YT�g7<��uG4K�{�_՗X���X�?#�7-'�B��z��0�$Տ��O��Z�}=�֬�dt���}S#Y&��:���dK�g����C{H}hR�Qe��>F�;.IG��k�c�`���3��g�����/�-/D����2p���v��;��紦A���\Z��{�7����>�KO�RX8��ҩ�;����:�Z�u0j�5.!�LN4���SR+�����f t����FP����և�ϣ�JDKϗ��( nG6+����������q�f��l�1#�;aP:H����s&�����ˡ&:N�e*?ly�oY^vi��r0[2* uj���Tl��#��{��D)��p�w��;�wZ�DL
70��\ `��>��Y�5h|�'[@��q��x�<rʿpU�Kt�"b�!��4^G��YB$}��|�[�%�o�����8����Vi��`V���ͬo����8$�g'���Ocj����zT�	t;M��ésKh�櫾tGx-_saB�I�E|������̗ε�z3�S��u��+�72Ք'|H���̀�]�8R�z:�}���g����YW�˵��D��H��%J��x��}̫̲{ٓ9�q�����`N�	E�Z����Zb��������%kWm�@*��Ki���^��J�J&�кv��J��;Y��N"��3�١�>(�5$!hYh�����D��y����B�gSmu�z���y	>y�7�?��,��z�����m8����s?�%>O�P;%���*Z#v�dH��qop��,�>͞~��:�q-0�,���Jj�n�o����K@(��.��o�ٴ�H�џ��3���L&����>���i��.N�uL0�_I�Ljl�#�ֺF��I���5p��+��b^��<�%XJȮ$�2�ĻTS�a�+���nQrT��M�i���Y��E���C�"&���1���rb���´Qb�~�
������1���@�V"��;ThCD��<�$�ia�y���s;%��'xf�%��W�*n �&A)�<�������$Q)~�̜�Z`Ս1^Q
�{e�acC���-�5ڧ���:���(���� o�n�웣,�7��\���:��*�+��|�������-X(ͳ��N��)�L�֒)��6���tb��h����{�߄ۏ!�0�q�W�4h!A�Vʐ��:t�n*Lg.;G+q#*�c�ђ�艣�֬�lW]l�`�cw����T�]��l�
��2�hP�MU��JU�pJ�%��@���tN��V"�+
{r\l�޼�Ǟ�䗙�Qr�L-ް)�gԧ3Ŝeq��KJ4A��/���k�rb�v��5��ؕ�8+R-�񿣞��F�3��!�C�� ]N�����I�G�t����k�$��K�U��^?E4����E�N�j���$hW�al��P��I�ɬ>�cJ��5����3Q�x���k�0G�g�Q&]�yV|h�!��!���0~�V訦�
~�Ǿt�1�6��g��^�k��$c{�!bM|�| ����oTm�!H���r(�V���/��C-�9z������]$b�M�W˖*�q���e�m0����T�-0umA�P,�Z|�7sL7�$Td|M�l��O���8���Ƌ�)0�?b��#j7��+Rz��O��� �� �0�+fB�=S�z�սz�&��Ԫ���@�k�}53��O���p!? ����P%��M$� ����sZ�Q�D��$ܬ^�*��K���������	�P�?U<]f�^�C�M�f;�Q@'���8åYye�\��Q�8�X��7��L(��:^��N��3;��e�	w�ԑ8�1��鵓�+��\3�`@���CH,=��㲒���)��9�~���O�G^>����'_&&����h"p뢄��ǚ��l���@��m�mt1����5�s����B�(����c3fdL?�>�ޭ�U�&.3�� aa��Z�|v��$j�f,ar���1vw�A�+��T�_!*!h؀��"�,HE�
u�1���yZ����Y�Y�|g�xb�&��q6>^�FI/�J\�(�檏��]�sA,HY|���ɯ��WA4Ϲp�E�^38�P!ƊG@@TJ��c��O֘p���J_c��q�وt~��Z��7�P?f�H�!-h���y[d�k<�Bv\��E����n,x��9�V��O�w���Y$���>�b&ލO6��*��6Kv0GP��C۝�ė�,��B���uF��%g ����*�
��L���LoV-hg�!����Cr\�3������fe/�!>�<�g�ts�>��)nv&��%��W:>V�')�H`�F�!Ҍu��h&OEt,
��M1veʏi��G��������2|��v����Bp��l���;�����N.���ɴ�,b"G�#�}�8A�w�S ���B��H%�n���\2��C�L�,���.�r��Pe��,;���l� X��W:���'oѡ��m2QAǧ�_�E�S.�0�U{��7\�AS�a
��-L�#�2@R�y��2��e�r�yӮ�b�ZihF��,��f8�򼼾ʾ"N���r�e�Hd،vQ �Z��Ԡ�:ﻧ�7a����Y�-�~���q���l|.�qwo	��T�������.(����5���b�Ϫ<Y����^��[rK���H\E}�- ��A�q	8�q����-Vn|�M� k�n@O� f(p~��ť��fC���M�`�c��t�ܶ%�ı,DN�D��0@H"&��%�1���
"�`fUt���?ӵ�����\����4S���h��\��a����:3#Z}�+Y#4}g�w�cۄ�r�ӁiL���Z
�Ҙ����i!
����N��k���U� ��^�ʾh�Fl�绺�Y�2بl�1���Su>�Do�}:?r�?a8ǆ�"`wn��޺�-�W�%jAhr��32�J�I_IG2k���A��?Ͳ2Ԫ^�"��<ר��:C�j7&�����C�ʼ6��.EWK�&�W7) �97/#�~EcIW$�ѳη�m[ba�3��f�S��`�W�j�P�g���Zai�9�?�Ӎ`*s�������M�g�A8-D��#�݁}���V��YX'�����z ��h'�/��@k��F�J���`�I�|[���s}v�ӽ�m�g�Gf�į#G�S����!���Z�#�c*�[�}���mQ���7��0�Y%����;&ձ���'��3��z%B���|��}ٍ���ݜ":�e1�k�Ai,f� �gm�9Wli$�"V[[A\G�Z҉�R*K;�x0�pt��Gg�hH���9�JP6I|A��:�M�R���'5�(-@pg�O��e6ۄ���I
� 릦�Y-����	���,�)�/"��D}�V�9-K�MТRb������F�ky��n��Ş}�A���a�*���V'H��*�>/>��/1�;	���uDv�	6I���	��|��"�k)��{^��q�Z�WY����7�G�۷�&�E���p�JĠ�Y�\����:��H����\ZC\�טE;�	Dn�ψ���
��e|�ug���)\����*�4�kkM|;i���yz\��N��Σ��؏B�������(j���V�D~����J�����~�d ���h�5ލ��<2����}y�x|��?>k�7�3�B�ͱ[�\vi	�a�|����Y��\h�u�,���F<T���j0'{�K��瀚�����HF!�i����8,�q8���s�Qp�����|ĩ'Hz��6~��*��v�����X$����i��p;ԈS\@���a�#!W�>Op�%�A�c�����A��mxVz�5��ת�6�E1�	�v����䟅F��e�����u0�e�[r`�u'���c	��4Tu@��w�	�]�:�\d��Xmʤ��F�0-}��%��s6��	G7Mo$ɢ�T�rf�	�y#u~+5�,�Z������&��	�G�玥}A��K�#���
��)7�Ԛ��6�Y��#�o�����]�TTOhX����zO�M��۳'�e��~s���Y�C�]�@t�?��;�`];U��5���X����(
f�ӳ�L���48��k�?\��IiCe�'�I9t��}�伙�Gu�a���CLbd�.y�q�^C���q�	�"�q���L�j)�S�&Z�	�T<4���-��r�?�:Ҋ�����x,-�d����( �G��uּC�{�\5O�D�x�w��ޗ��#	wx��aȾ��j"Ə|����NTe�){L���^:;�izI��_d0F�qd�R�:��s̊~HN<��0�]�����ߩ��v7w��T�&�[��e���N�N�ߡșD�DaG�@�ǭf��B��!��+��3R���Kp�øk�y�ڈw$�˺!S�Ә����S�\W_�z�rX�����Ӧ�U!�\4�u�U�)�?yPHI�N|e4-�����p�}lQrk�5lK>�E��>�>2�w��Pu�cH�'*��kZ�$Ց�v�P$�GHp#�k�Kupc��¥E���F�ʌ9�+�a�L5�u�Х�jW�F�a�l�2�	��a�%��v�~�]y�O���@�mzy���S�9-�,ü�z��tl�v�e"q�a�'�[�[�W�$�"��*�5ޡQ�F���w�Ț=�8.��¥��b�ytc���z������A�����{�|i�$4���x+�&�`��^��UD\dz�w�F;>�\v#A^��\�˖[�*6�RkN��h�%��u�9�d̦I��w^i^�U���㦙kx��&E@2�02���P�4�����h��7��b�Cf��{B�U�3�� ͇ѫ�X��2;A6��^X��� n�fUr3}`�������p%oYC:�E#�`�=x��eQh)L�d���7�0Dr�qW����Z��u��Q�>�Dn��[@�	!Z%��v�Ҽ{B�>���=w;y��a�l� _;p��)����R��v]����S���rn��Y!�9(�3@����e���j�5/e�2G�~j=�)d>��!�T".�f3�߮���/Oֻ�FAؒ��	�fcL�9��uL�ZG��L9�2��>��W���h���pËL�U\xP��7gJ�����v蕟�-ܻ��.&iI������M�*�����n��]k:~�֭D���F�f��PHn����ԙ���.Ǎ�o���,^ S����:vO��j��td�\;�c�k�jh9�-c����'
����<���H�1�*̀Y� ��z�.?�0�7�<���A�286
�[h����d"Y�V�5F�
q4]�L�58|�2>�F�~�o
�m�\�t�"A�8&o�T�C�O}瓁>�y��,u]�>���D3�=�3�}RM>��A1�Sz����W^��ڀ+w�������v���"m�$3�V-��>>&�=�C������#��?d�l
�̺	[����<n�(=��C���,j��_���2���&����	252`���?D�*l�[�䝄��h\N��4��S�'Ck�KЙ�\�~��xnb�C �%!����e$!��!�S�(��ҩ�m_�c2/��˪��]���a�T����YNtӔ�6 �^3���Ҕ�e�{����3R]�(��I���d'���q���o�pѾd	�᳿�f��#(�7;_2�׻�����s�
��!��� 6H�z�Ks�g7K���)�s_JeGe��������	���|ؾ��Q�����H�U��/3T�������Zr*��\�䗣�	C�9�u�H���&@�k3���f1�/}���M�G��&!&���24���ְ@"��ĸ� 5()��6�#/h��A�3������4b�kJy�����<�����u��\RP[M�X�Ȯ<'-"�cX�M#a!�Q}񢿸��H�t�;-BKC9��������/?��W�>�=��0�*1]��o�!{-؈��������V�� 廬
�Q����u�j��w�����!Hօ�b���=�ϲ�I=�a1�Dd�f>�r���S�Rm�T�� ��o�P��J���;��_���R�}c��K>>f��_?f��~��/�c�H�q����tU��䐲h�Bq��$M��J�k�V���%�!B��#g��h�fN{q�����RػKE`27�X���$G�&z�b���E���/_�N|K�o,g�����F��ߜ�<ϿV+$�$�5�%�smS8�X��3��_}��oY���/�-�Z�*�Ӵ� [�B��W�������o�o��@8��K�]�������� �H�����������<bl%�ȑL����F���4�ƴ�G��9P`��ڌjzIv4�RU����Y�|H�R+[T�+Lbt҂�E=���|-%5��_��bه�L����B���[j�9�V,r<CK	yT���D�p�RŒ��xƸ5�v��N�}w������+�s̰��p6>W�LK���5�1"_�I1�v̤�
�wlg�{��K	C��¥l�hS�*���B�z�/��g���ѕ;y=+�7���/�0_�<�0/qt�d������0tA��||AZ�� �EG�p�>���@�N�Y���"x�A��W;�:�$��A���hR��7�V�[{�띑���6O7��U:���Y�sܦu
��q[R�����V0�UM}^T
����C��)��� ��G㙰��4����5��� ̳흉���;�wv�X�߁d�W�w�4� '�6�ZYS����h��"�OW#Vx
�!|����)��}i��\�W����$g�A�v�MS|%��h"�4g�>M�^L+!���	�A�fہ�l��2��m����d�lJ�KQK�R����r�D �`աJ��H&d���M����]B8��~�<0[��|C�]�I vb�L�X�/O4f�j��	mB\�%	:
�rđg�2�O8�mC�p��E�5��@T3ܯ?��<4:ևQO�d���,H�2aj����n��S�_�b�Y(y�6���,3�W�@���րJe�P�ˬ^�^Ƚ'"�ڋǢ�Q�,��m�R�_*0��=���vM=\�<�M	�+p�o沾Y�td¤Q�tA�ix���L�/&g�?���xN�/�,�mK��s �ܧ�Ŵ��� Y[��Ͻ6%�t*K�AJu&,���þ���|C�E*P͍pi���*�W��N4�*ӁôSt�v.Yhm�{2v��A��Ѫ��F��q�8���/�5o����|/�,7���~{vచ-�8�p����1�����e�[3*��Vx7yԨ��� �n��:�;(x�C�	}<6vc�hh���Rb��fF�'�D��d"a�ԝ���0;%��fk��ZL����Z�N� �������F�>���nrCq�ۛs1�Y��sT�3����I��<�9����������U���Ȑr�A��
� "3`��zЏ��f���d]*��/W���du�r9����6�0���g6�������������l�v}����7�E��
���nB��"��ɩ��c3|XoV}Q�)�zfN0�#�N�N���̃��5��[p��涻L��� ����� ��������,*q�ȹ�58ח�f:QK���t�*WJ]��\�-�jZ�;+>�"�I�%sJ���KwoP�u9����t1־���:�M�K>���a��d�4�j�.ԺTt�FA\��@�j|9���ȳM�`��z<���v��1Fl8��B��x�y���u.׿�荛!Î�@�m��,��OG���؞��+��+��젏�ye����
2��x�8�P�A�\@.�D��q���	z�C}F���+��?�n/G��H�1ƛ��]}0��8�G� g)�.�HgJ�Y��n|���غ<(9��o6���]�6�h1��e\mW����Pʫ�
E K�K�j]N3�0v��UIa��p�9��H0����V��.�K0��;d����8/��}R2-�4bwF�^8���o�9��RV�11�� �´q��׀�;q��b��G�Q�����}\�\��y�w�@~4ꄸ�М��2�`�z�'px��qLY�})��l�6#�!������vO�H{��p�%	~��騑�5=z�9z�Dar��^���6��HĞk�\IsU���L_�����[c�P�'����d�eH��*S����*U�e���8sy��"?=fȆ2�d�Xk�J^�}�Vڻ���f�Q�g,�"�]�ڋg�@2 k�/J���6z���ER&�e+�r��D�b��ܶ6�J��Dƪj�|h�M=�I��&��Ѥ�o�؎Ì���H��H�¬��6v/��(BrT�`N���Y�kӓ��z���L��&�ʨ	o��r�߹=7�k��O�V���:���*���|�!Uf��_ɖ�Y�A��i����"�5�"���q�� ���Qrp�M'�\a):�/���5aͻ�]���íRv�k�
����Q<z��3"�˦R������ȶ wJ�S!(K�J����,HL!��%X���.?� �х��T������l�����J;�n��qв�R�P]�^'i�&�z7c�c�
@n�I��/���k����~˝���M��2�P��}�@�A�C3��S2�S����ņ�~W��Q�G�iwi�6���}T�TWcZ���T;\�F�C]G����Bl�A>K�H~V��b�&��n��tC�G��{n
���Y.��Hk E_�%Uo�Y�[��	�x�
(��VO������H*o)-ʫ�d#T�
<�+q�f֝6��y�1Fǔ����nV�G����h_��m@�#��P�7;y~��
�s�H"(�ݳ�Q���X�Bhi}m/��+�D�]�˗� �����N��zZ�	�j|�i�<U��mp��'��?	#T��eLƺN��%,S󷱕E�,��13�h-�JA�@��NJ����4*&8�,�%���9�-H����ѧDV���.�&��ɔ��$8?��T%:7`��s*��7pM��<w�>s�WG@��cМ������������V��[c�Z�R^ˤ����nɼ]�Ț�+FHnn�xC}���8\!��w��\@�#��[icq���*ۭ�t\9�ofP\hwŲ��z%�%��Lb=�}�'�e�3 �F�C���g#B�Bp��u3�����A��t�@+���(^4�����m�&����5���^ȯ�w:�5�F�1-�!6�[9�����H�q�@�S7��%�s�'��oḳ�Lf�cH@�dv*R[o5��ڲ(�;��ղ�Hj^��%�w4���h����K��)S��e�-&��Zj��$FU��&���ݚ�����V�4�M��̞~܇V[�c����R�̤?q�'TjOV�XqA�#�V�g��%�H��>q����­��VpD��+�F̓a��jZ�O;�T�ЫG�@!ӭӴ^�/������6@1�����#)�霷��*:���Sck^E��a�c�,@.���a@(��] b!'�H+��$�2E"~e����a?y��j5�eD�d
\,�
Z��Է[�m��wT�We�?�����=�����ޙ�>��L̼7�'��*�8 }�k#����:�<+��������R��j������uS?��}����^#�Z�����o��yD��Z�[7�n@X��bK�c��7�# >o�fD,\`�"M�$%~c�(.�uUN
X�%�CA���[_���GO���o�MC,E=�~g��Æh�m|=�v��<2
r��rix:vT�8���=�������"�:ID�����d�x��Guo�����z��VU��ƶ��S���XɌ��̡������O���		�����Ǒ�����$�L��WBx"*fU9w�L�����::ڭ�[u�>��Mv�3�R��30"U�x^X<�ʛ|L1x�/��}��_)����N�Ѩv�K06�2y�e��_[	����O�}��Q�э}�K�O�w�7��n����K�a|qMo�VO�OCQ�NN����8,P��?<A���g�|6���:��Cy�����*��h[/���2�?	�p�`8����	�σ4N�����G}6����I�_��"@��_#Ѐ�(�Vˈ�$��z�5ſR��W�(б ��z��K�p?T?�Bb��=y�?_���4���izID($��L0���e��o/���Ku=ю��Ԝ�6��j_�ԙ��IS�qkysb�Y)�r%摖~'��,��}���g��Ň1q�����$�Ob/܏;�{��4>�j�ױtu	fh�#�=fg%��-��0���Ƈ��H��y-^�H�3����Pl2+Q�w�nߥ����{�i�{��ɛ��[�?�i�R�����]�&bF%w!�{�n���$������i$M�C~|]>?m)^�F�OY�:Sd$"�m���z6��9���9��ꃕ��񾻷�)�U�>b]��ϒ�ӛ9/j����x��e-|�+�Q�D�)y�O��jD!�#�������!�v���{i�D(!l�S*z��U&�̃�	rʌww!⾍~����i�����F�^�:��S��q�\����y]�ӯ,/'!W���w��m�W���eF;��DB���� (=&�A�T,&�P�O�/�B��YQ��ܼ�)xz��OwI���K�fY@�
p=PhpCU^ [� �ʏ!��eGk�U^����M�PR��'~�	͹O��P����j��<�UB�`�Qpb^"�ƅ�..��y�0p� �ܵ�Ay8���~�s��
a�iF+iS�Y������Q���MM���n��P�1^����c��K5/R��KF�wn]�<�$̈́��H`���"��ҝ-�Szh�(I:[�Sj�=����M>����%�\mG)�K=�I���1kԇ_|�Ib�k�v�Q�K�tB�9u��_�L.d�%�wO� Q��L�x�����e��wZ��S9{�E�M�@-}�T��iVM�g����``9܇݉	b�����k.��"P�E� ���F2S�LXdS�V�#�yP�����3��n�i������a��i�<����@,D- !�E��H�@jZU���E�n!)���ǲ4'&nG֬E���U�B�ա�?^�ؖ<��s��Q��)�Dj]�`��Zi��kzW'<����[`s}twg�x��E	�D��>���M�䌰շ�ƕ��z�(kӈM<TxRyv�A��������]��~}@��h��P�q��T����2 ^��F�S�ӈQ�/	NT]$�O%o`{`�hM�X-�����N>����i�%1}gD�d�Jh�5��P��~�hM#��}Ι�K�x��s  ��\����<L�O�o�a��{��cY���f8��:�j���L�'��I�krlAEJ�"M)�JH�xWN�R
<,�V�}pO���o�#+{��+�9� QO��c�H|�V�����j��.I���^Gt�Ǯ�Db2���҂�n���4��x�����y?�����P���2�b7\��11������@X���V�Ǆ�m��[PR~�
)sn>�b$��t0𓭛,٨l��U� X!"m��%��>�DY%6/M�6�e3B|HI���-::2���T����0F)�F}se��v�S�Z�2�*�:a�I���u����I&C��4�Ǌ+Ղ�?ZU �ʂB�Mw��3,
X�~�>��x4�����1`��9��V+�!��v.R�dW���7�Δa��� ���P�<��)��N��e�L{$)K�G�k��Ep|X&�X�� �n�R��v�>r�M����X[�e`Ne��c0��7����n��+�Nihΰ�o��e#�Z�GJ��P��qG����^�aٳ�Rggvl��k�4���bN�W�Wj	��F����v��4�f�*t���UY)}E�^:�pH;g���y�'�l�V�%/N�F�jS��/��O���2���;`�E�{AXt�W���t9�����s��9o�@u.N�S�A����'U�i�f�Ƚ퓀�4^\��E��uIa���&+��4���	xŪ,�Q(l��q fͯ.����F0����{d�b芋��fQ��C$��V�-����2��ԧ_��**���
��_&,S�]#K�c����ñ0v�c`{7o����-��q�^ �h]��d��U_Y��=�:�X�F��F�2�͇����M�V	�	y���]{3��^�����u�V�*x+k�z _�����L9=?��������V�L:s�bg�~��S�"�/����l-����Mkf�]�K���
���Ʀ!��j��ۙ�H�L�^�q"��^ڀ���MѾ:m`���x
�W0�� � �cS��:N�`M�aݍc�G�P�5G�3�x6
�T�)�*9W���p5��c2wk>�N��~��@b��jl��\ޭ�\���2cYai ��dh��äN(d$!��>|~��W͟c@}{ċ
�BO�)��'Ƴ������O��	H��;�&�O��]��	�����`IG��	ҽ23�O�d�����.���;a�p?�~D�D"�.d/��|t�n89z8V;e��K��C�C[���l�k�z4Z2����k��������xi4�T�\hh&����)c�\A�2��JwK�"��7t��u���S����"^�ٟ7�Ԫ^��=�ud�G�~*���7+���ǥgى�&��A������u<3�u�$P�����C��-8$����p;9�L3Z��q_J@����%A����,V
poC�X��憛���g�=@[����"���>��LB��\�juu����^���ª��R��W�����J��aSZ-w��Z�l*[p��K�|{m��/�B���ĵ=�N
�Z�Դ�����v*HU�!����!�u5����{�������L=�{�=�on';�jI��*����]���i����V���]
�_��#rf5�
�<Ǣ��5�
-wo׏�K.Qd�U�ìL\�@%�n��ސ��tw��n� f���@Qߋ/�����1�9򻘄y�P@�G�]���E�f!*�I��ܽL�q�^�GnkE]��BP��c֝r�d�%>���qtǹ����F�{��#��.�i�4�I��lo$���F�v�4:���Mŋ�z���Qԩ`��J:���]���W6������I�����?����(�}}��|���YXkH���XZ�s�A���� 6�9�X� V�LI�Z�����)jpo�O���S��Z��d����I��,���I�fs�)h�·Q��0�! i�2a0AS[Bd��f��Ձ�U������K���	Eз��G�L9$ ��ǃj�퐛%�~q��H15t�g�[M6]5�S���a��>6���!��oE�aJ��6��Mx�n�?VY�и:��:��!~�2� (����)�&� ��.��f�"�h�S�f����d ���*�h	ː+�S�-�� ��Ą���S��Ӯ�Yd ��|��zB��#���E���7�*���� S~π����)T%����}=H����D/�H(�..�{g]y�$(���i(��� �G�D�~���H!�մSw���`n&��8���-l
��W��*��Z`<K ,�@K�5mo8%u��S���1�U=ž��h?�	Z�M��Jm�+$UͰ*4�6��|�雁L�$��D=��th�����x.K��g4|4�#���E��������oދ�~��N9�D��M�4.�ZiSg���`538�"��]PC<�XZ@s��X^����?�#�Wĸ@��B���{�0߇�Q�$�����^B���j�j%x��l抹<���2��o���O�X�z՟rdju��08Ƅa���j9���&�8	�iݼn�4��Ĳ�q�ɓ�.�� ���p[�}��"YM�k���i}�S���^�����M�3�U:c3�y���Q�-Ac�J���ȇo��5��/l,��g��q!����FNzl�{E��BI@GEU���]7�4*h~l;��5}l*�NG�z�mH���w��iE�`q�B@p�;]�x/ӕ�F��i`��� /���$�>���sYފ�Y5���O�vf��π��<�a�m&AK$��$�!�TB���a]��ݪɍY�S���-Y/��� &�F^֝��W����uf����w��r���Ҁ�N��i�,=E���,A�r�\r{7��os�_�~����8���m����!ߓ�%��U�XKE��f�NרU�z�Iaha��?c@�����ˉ��� 	��7�`~��Փ��*l�o��Mx�����R�s
ч����|Y�i൩��#����2 N��
��x �ă�#�d��ޚ�˦�P��?��?�����8�c��Ov�u�X��	}*�Ǽ�z.n�9��[�F��VQ@���Me�-��S�8����;�.q� �q��C!҅ѫ���r���۱"�>�����K�b���F�A�Ѱ��pC��l��@�@���������fpԸ�xH�vy���ʐ�o��<Up�{"E��=*\;��'4x�<��1H��eC�Et5��~&G�9�~\�aPC�����m?�����L����c��� �Ah]6�oxUd�����(*<*�Tr�j�?73Z������2F��N�c��Pc�N�>���mU�G$���9֢
3���$��HKj�0��z� es>�����RN����d�B��2�q�U��q���^;)lqp�G�>��`�r�fp�����ب�U�r��Nq�&m[�̋���	��M���9�ڸ��N,�ŉ���nj51qY��n�ɕ�n�uݙ����K3c�M��v�9}����]pJ,��#���#��u�ʿtV�h����Þ?�P�[0�� �ߥA�>c�u �]y����r <HD���ؚ�Ǒ���GT���E��q9�&��N�$���"��0v>	�:�/�s��:c�;g"x0`U��؈g%�9��i��1�����S�If�7`�C��ۄV~�E�<�p����Ib�w!s���p/*�����њ��,�(!vK1���t�E���?���<�s�n7�j���-�콰O=�Nbzfv����nx�BUêT�Kc�$-�b�P�5�|,���=�|�'氺Ri�"��kCx���rO�+���>7����kגʚ�]�iD +�8<c�����08Q�GU�PsLq���Ry�V�O���K��2MM�#Ix�����b3gp}�GW��
s3�T�D��wf�#�s?�V��f�n&SAs?`z�b��ar��h�DK J�<�?�ߝ�X=˰y��̰h��7T쀱�Ө��,F�T�3���q�'p�lb��r��P�W��G��y�R�.�Z8�1͠�<�.����T��X����C�Oêw)g�#wW��F���<�E��on=z0��I>@J�1{�岏+�3�bS���뵬>R��?q�����WӢr�Z�U��'�;T
�bE�}���}��ʢ�����0y;ٻ�a��Ă�

���Q��$��?�	ϖE�$��F�Ai����C�Z��(�,����ˮ��r'����<���__ؔpb�u�Wof�f��L+m����s���D.n��o�<>G��&v��@]٦Qڨn;��;ٝ�:Iشc7v��\,��y$��3�
�����C���c�"\"]���@��m92��Z���9�F�V�eQnx��
�����~�%硦��	0�-GH�1̩���8vZ"��vz���g�-[y�Õ���yl�|W����o.8�d�E�����7���x�E�m8Oa�������S���1T�����r�LE��U�d#d%e�5@�� ͑������dk�����ӲL��	���o�����Vڣ|���1�(�$�Γ�[R��(�϶f����/g�5(h��aC��m!�l!��8�+�V݊��C��,�?���m��:��?|�݃��YoZ�PWG5,��ې:�WZ#RʥE�g`��ko�9�>0TTN7�e�����dS��S-��9��*I�D�?�$Z]�����,�*���5P������a�4��7_
y�T� �*��N�o����"�wh名��8��a}RU�Gbo�3'�uh��yc2����|)�`<�[1az⊑��>�D�^J|�`�'��>1"aU
�Z�m��]\�P�H2i�c�&��E]���;3 |����2$y����\��ؘG�0K�2�:n�7������<xt�԰�8:/���5���b������ldFq�=n�sy�g�?]!jw�?��Ҿ��7�K��n!�p��T���z�ɋ�C��a�MSO�T�VV�,
9��9% >FW�۶'��=ϫ+a-dU�@)�m�hK��C�˕=7ӫZ�7�+}�g�4�ǜ�i��k ]�]r��>��X*B�R籭)���n��6֤no���������+���K1��!C����6v�l���r��^��aq�Y�UY!ܹ�q��NᓜUuKHU�3��ba�� +ة�l7�������}����*?�sxo�ߤ~^��)���!���23Q�q��O�t-����/������\��)9��WSJ�Z ,�6�&ۗ��I_�<X��[�ʌ�i��"����:}�G �i��n����cȻ����#뵁��< DJi?�BvJs���ԧ�*�v���1�@�c�8���)u&u�&	�+L�/��Z����a�s�0�b���W�Xp���ID�蓿a@�s��4X=[]��0�!6���6*��7���7Hɗ��	*�/��$yG����+:���pE��(�l�%B�qF�kEU��c?�����wa&����"����F����`������0'�9>����>�%L��Ѝ=�I�o�;�&����vs�9P�	�α��n��c����5�"kGɛ��m���v�t���E�b`7����w�^ΏW�ׂ��Ac�9�{w*�9ׇ�̚�S0���<x�H�6b4*?��G��ѿ�TdC]֫#<-��=%�o^����g�ZRpM��Jʂ�n�~�h�G���J�)�����C+�@+�ʛ� ��lC=��~���I�-�@�t��(�C����~Ud	m"�^U����8�h��B,ظ�٥!ޟ'�ʕ��$�R-�A;�.ƅJʌ�����i{��a]��-X�&l�'-��aK-�Q2�YPD��A�`h*���������I��lwE�'��Kğ��\w�� ��`�.Y��v:���0�0� ��Jz�
ܬ��ȷ+�ue�+G��_�P�a��E����iҒ�6��Zty���w"�D3:e|�g;��;�LwH���Z�w���4��(5!�� 9�A <�üV>��ۀyҮ��tU(��yxB	tI�	'�M.qA�G�Ο8�20��c��Ek} /({QD���Ԡ���x�5��lwc��O�*�����OW��ʑ�{���)�zn���s�YꝔ�#Wh����m���Ԉ]_`d�z��t#o���(�"� ��Ar�QZj4�v�2��F������S�?p.�oU��"q*g����D���YV8����:�y���9_2���8��Dm�������+L��,�O$v��#�J4�0N�>���O��٣�qbD1����%���a.m.0�6J�7������?ƗN�=���vat
HF-Z�B�`�)d��:�W�����Px�8�T�x|c��� N��Ҙߥ��U΀��yq�c���[��S�CR}�����)�I�nq��θ�%'�]��~1++4��~���3�/��� .��K�=����x�iDE	/c��<=d��-��؉4LE�oW���d@@�z�mE����	Dze�4��y�Z#DgHY8pɿ���Y���;Gͼ>^}�-[�q�Xoa��̱3 ��gw�Y�[�(ĵC1)W��ɧֿ\P;�S���Cp��!G>4�1N�*ě�$��4�>d��t�-z%U��۷�Іd%>ȭ'��nNY*�YP��B��G��1~P��ER���������}]��k����\-LƳ� .��m��IǍ[ی�̧,�ȶ��:�����R*�B�F@�T��`J�^�z����ތ�>��K���῁�]��z0������.�Ic�+�[�ãw9��ph|g�_a��#a�	_La/����
���� �gz]*��j����r�F���L+2`����0p�}�i��Wn�]��]�2ẹ$�W�ό=�����" �Ff��b�:�m�b���+���'���aT��n�	�=�*	o�T ���D��xU����V��ZԮa������R�K���q�j�$V\3����RX��~�?V=�>�#
���?��~��O)����1)\�x&�!�#;���8�*�?8՜���=��bQ�:�&�l�C�F�ص� ��y��L�xGE}�ܖE�tpO��崛N�1ͪ���9a���H[��L^#j�Ui,�Nv��݀,��	���J��G�ǖ���q�<������~Y��<ܰ�]��G�tZ��'�t��-�	�����	��������_��0ur����q*�v���f{\�MѨba�
i>Qf�?��;6'"�TL}�D����2$CeR�_X�����h�.pT[Z=)���(�IB����(.zL?P��1����e��o��1��]Qtas�C+:��G�C��^;G3�"m�XN�A��x�]��2^n�P��H�Ǘ��&3��Z���=>�t��9��'(n���	a^��(��Y5��\ta$c����D�A�����<4��_�8"T��H�T���"7��$�{�m��v���$����"��<ƃ�׆��.Uw����y��/�N$�#�pxh+~ԃϮܶ�XF���̑�ub��:����;^�|��
i�ea|s�nSa����=j�V򁎸�>�E_~Jo����E[p�'��-@������C��88����Цx��k��x7���*�v5�x�^�дD�	�fJ{�=t��'b�N��JZ�	���d�|�<��`Ⱦ��e��h���o�fTN��U?�[�ͽU@׬��!�Ue*,,B� ��w��NP%3PL��]����a5!�#��9���-��x	`u]�rl8V�o����~T�#���������8�4�J_k����$�����7Ђjx+�����5̀�5�5��!ߚdaM��;]PO����_ya>0�&r!dt�M��1p+���"]2H�=W0soakn���O�ˋ��G���g[߽7�<J�}�o����:�K����2�P�B��V��)H�3_ �#4^Pr ��GZ��v��\�����֓�T�ʁZ\�t��U뒞��k�S�B=��P��+ꕊ?�>~݀.<����z��`RM���!�Q�NM��W��Z��*u/�C�x�B���o�}=\>{,�|�O����� ~�@�$\�W;Y��l���~6]�~B"sx8�?b\���W.��5VE���Z��x;�5��F�u��CcQ���7w�_JF�7�$r>'g*ȪE}�ރ��]���-��q�/��Q�C-�Q�gۋ���{�M�~��N�|���;��2�H�a��$.,LdE���mn`?h]���ϐ~#�֥;�*�G������'}8JU݈
�8L� B?�z�ߑ�ǅªՃX��~L�Wd�/ķ��q
C\�G~\v���铌2��$XL�Z�Hv�OqP}w������)�Y�i�#�������hL�-c�,e���u�tL�DMU ��I�יB$>\ Ԟ�SF?��S�G�X;���I��J����qW��&w� wye7yĠƈ���Ym��1���ЌBI��V��F�n��сn9m������5��7O�����l3�q��C��r�sa{���������^<��o�}������WRO�Sl(#�(7.���V�,��:)UBP%�m��s����2�!8}*"77{�����Y\�}.��^����q����nR���p���{��~%\�(���.�n�s������[,JM�{??�[��?��}�V>���}��e}��8��ش�U�����c�q˜��S
T�����4C��W2O��|J�r��?��<��;2bct��m��D���4�M^��7>�$xpn(p���ϱ��%�]��üD8� ����Щ��L���=��!P!]�R�v��.�|#=��X��9K��|.�k^n������;��gUhA�w5��9�������z��{����h��Tt�p,9d��|��/���w�rȾ���<􋘖���j
�"F#m���k�Z��'�����q�׹XJ�pz�N��_m3�N~c�HQ�X�:ɘ|�%l��8Jk�A���r{����g�P�7��@�/Z=͘���+���i������6�H�Ӱ�,��¡���j������YhLx���^�˪�W]H�A�f����ƾ���Fl�s,,V����$�T	#����4R^l�`F�+���S��ϋg6LL>؇d�.�hN��� ���W�-gJn��@6�ۻ��CZ��1ѝ:0� ڈ����f�{ڷ�F�����C
�	��-pa�_�����@8��Ѕ? �U�O
{��+�M��{���� ���ہ4��=��-gkIl�V9C�n/�ĭ;�Hs/D3C}� ��m �2�q�^ehc��F�L�ʫ/ Hȁ�Ú�3� L��)��}c���D�pM���׭�ZH^�L7�~f���&uf��{2!����9�P���6�>O��>
��f��wɧ�Y졛<b�������L ���O���=�b���{U�Ғ��|I_5deD�?n�����D�g��8��`)�Z0ɩ�ٶ�X��f�/�-�"�Z̗`��@/�G_����b�	��,�U���X���K��B\�)Wq��G�d�n�V�J�m�kFrͤ0΢õ�Kn
�ս[@�J! �X�HD�g���l�i��&F���*�PP�}�qנ�"Јl���~]Lb�#��!��9 y���e���[Q��<�����T+�΄�?�ť����_�n7��%*v�@wk"�� em�w��٩�_�!_����e������?�y��Ԁ]_�p)��?����	�~A�_�AG��� �Yl�Bb�&�y�cm�B@�
Dv��X���s"o����-��u'5-��M�5��=f�����j+d�/,��v`�j�T�L�4�RH�����Cj�!,�aŕ0����!n�lH�I��}Q1��:]�S����/�J�`�L�3k�88[Ujm�"Z������.���ZV�,�OS���d�^lz1>�72q�w��}��ԋ��l�^QDB��Y��ծEYwͅ�e?���pc�Y��J@�3}QIU$��W܈ӵo�?�c�/�'(��z��U~I�un~����E�I3k�G��in��D��6z��.D0����C�4�N!���Ȍ%A���K`x&}�S	�`�6ozS_M����K7yD�印ۣP�\�y�p![fB!����8֧��D�Yނ1���05mz�W��&&���$��p�j�8ھ�u����E$\5���d�W6#p���&��9����睰������o b�^1��%�1���ni�'��"!khYe�Tt�Z��\�0=�#�.h$x3E��_}���ԢǮ�a!�,cE��%���U3lF<�g�?�����<ԥ2q��uդ-�w��Eo������9Dc��NJ���|s1A�oQ���C8�DG��AP2��)�]:H�h:�#��jn	s����#��@��:^dY�^�d�H$�v$\���� oIy*���B�}X��ն��x�IP��όrˑDFX��zT��(�Υ���Tq0�E�6�am�����5o��V����(t@�*p#��������(�YΞ��xa�O���l���eb�SϹ<uO�.k<�V+�?�q�C�j>qcL`L��H�sa�폑�x�P�N����3�u�ҡ���?_���aq��ʏj{Ր�@���6���r�3Ig�S��2e�^���S=B(��'Jq�*��٤k��d���h�8�q_����]���f9$`���j*���P:�聁B���>Өi�ֹˉ0Ŗ�/�7h���iʠ-zff�q�`!�D]4�l�[(_�O�|�W]��)�װ���VP�r{���;�a��v %�k�'�a�hvL�'ȉy(���J�zQ��I�	w?�3�枱���oDr�.p�1 �Ho���TyB�m�Tm�9�	i
�>��6Ьrԗ��t8��/`=˷P����G�����_s�w�ٺZ6"�� �k02F=�.�EQ�se�r[9a<��=@mq��-�J��KP;-�Ο7�s&vx��2K�np1�k$���w�4�0]�)P��������U��OθAg��*2�����E{��|@=l!@�H�D�$���xr�1x).�����48B��3���-T�?0¾��>/D��߁�Mh^��K��K}��4T�V䱰k��8l�7��(�k��K0X��ns�}}�k�I/�	�����;/kA��,���6���jv�9R�k�Tߓ�|i<�s���4tU=�2)�.�:�1oa��v\���K[���U*�B1�uϳ�+���R� �&���VJw�9a�a�x���6�	��`#�@bo��kbIIK�cht��˸M��D@՟��������ύ�����Y�J"/�55CJI�k𽏀�O8�|H���H�lnc��漤I�/���k��^L�.L���3�s'�>}�N	�3~<~�Q�.���E�pd�	Z��e��-�Vw���I$��%l�8�k�8`w,�.υLE,���Z_>b���7�����VS�o�*A{M�	�jf	$B0B��tV��'�_�K)�һ]P����VR��x��i�c,oܪDVa_�{���0`��+S��M"+���``<
8PUGJ�Vr�9=���
������l�PIh]�7�9s�����P����o�H X�l/��T���ٔ�#��!pN_��	�|x���NAc�j�[�CxƯ<a�]���:v�I<��D*vIT!P�#��#��`+��[]u�=��������E�ʭ�����v�7�G1K].+2�$��,Ĝ��o�{eMߖ?~H��w�F����>S��������O���`Q�L0�y���jdW=O �_þ}����}r>49�Ш�����.�=v�LX`r'�y��������� �#���$0����T?�WC��y�_}I��5)���0�6�F
�gI���B�E�g�������|���S%����dŐ��`e@�3�tLF5����/7��S^�K ��@"����!�D���r�AfֺR.խM-k?G�o� �	��I��>Ab���Z��wj�j%4�	��u��L�t!0��㠬�,��������\�E�'$�lY�]f�Vu�z�
�"k��� �4���($!m(�fi54T��:6ZēD!GԪ/�Z_B�o�B����{�4�����=���w˺v�	�W�x%��G��p�V�f��6����<���k��xN��P�')�,�s����g�?_�r8�\g:�s���`��mƯ�E���קB2�^[����&����9e�$צU����Z�˶��ɂ����*�cD��O�8��!*I�cڼ���C��p���p����v7�S�].#f)Mb�ϡ)9�2��.Z39<�q�̳z<1'o�Zs{Ͼou���R�M�2-�v��6�RO{H-�K��6�[b-�8�}�}>�ʓ=�iȥ��
`7R��phK�\�lj����S�^Y֕ ��Yגu�k����ڇBU�A7,�=[zdߖ!�D�=��tH�oV�4�N����ޖ#k�Yl�j:�ULo..@�h�(Y<�u<ں�����7��M��%��T�iY�oJ0�y��b�0��F9;w6n���d�*�K�D	�pTMz���@H�6��lb\�ǩ�)C��lGK0ؽLQȏ��^DhVWa!�/�&�������1 ����T���J�"#e5�0�U`މ
�����*σ �g8�>�I�,!��"?�wa������L��_J��Z	^��`��͠���^��������o�C��1�m���r:���ˎ.�܊m�W�t���MP�z�-;ߩ�.A��f�]/.�D���Ư���Kc�.���e8-v��![�bf�����s���L��)���P`Y/�l'�_pv�Mm�&acN��~I#�H�(�s��E:5c�d����.CSg���˪+�j�ےc�r�=-�U�S�ڣE�]Y�sqǰ9�eA��T�h��Jh�%<���oR�I����̡bc}�cwt����Z����Q:��Ӛm馅��0	ᨺ�7B�缻yv*�p��	�Z�Ì�WVO����Hq��T}�VT�w�w]ũ	9gv��Zӣ�S�0��3&&��������n(5ę�������]��7���5
�h�e�A��5:�γF�1xA� 
NB����.WU#<����^y������unK[���}��~9�v�:B<���ϟ�7��kU��1T]7|t�]<����Q�\���ϋF������.Wξ��ؿ���<oG�v<�Dcs?�% �\�*����/�gr�2%%��\�R��f��1�,�LƷs��:�#/���&�:�g���w_�^8J�]�|���k��P��}2��X�V2��ӼL_E�����գv��P1ğ�"��d�͢���6�Wh&y�L�?L�9
�h ����K=q��,|�E����x8}lz��I����B%�|��h�1��4%A��Ŕ	Ew��mf�ҷ��sˀh϶����Ft�#]�t�:�>np��y&�"67���F��O���pa�3W�g�Q�cNdW
��ڰj㒠���b3��1�X�N�Fl����[�ZԤ~�%2�*ӡ��+p�O��A����K_ӑ�[����9m;_�H����t{����5�P���g����u�4Ɯ8@��P��_�u���T-�W���yl$�O;^�g��h"�ʜ�d�Ҙ�;>/t���cW���"YD���ٕ�J����P'���;\�0T�6�ӄ;�(�m�#�� y�K��Y�x)�?���
?�|j��R�b� �	Gb���̫]_u}c:Dʭ�b74�=0�]��C!���F��~S���
'k9�]�6���eޅ�h���z���L�b�h%۽�V	`� ���٫��7��Z���B�K'�ª����Er��"bfU��`�aS5�u����Y��#��ǖ8U��~��y���Jb�`�Ԣ���!���IW�o��nDB�%�l�xI��s�B)I��r{.�[3�A�
\��De���I�*�)�Ir#,��o.�Y)�kz�%�&�M���(GB����0^2�
�@����`���k��?��J�T���!'ye��������'q����9��C{7^�J��B�8N9����in�;�f�}<e��9#bOŵ�ּO��p*���d���D�N�w/�n��LGb��B�3��=q�4{��Ȃրb��e&2�'ú��eܹl�[M��s,�NIW���d^�	)��[{VAB���4Z�����i<�t������)�
�ʩ�ꔽJK�ˀꎽGTU�(:�W��v��MR�g��o�l�8β3zj5#c%nt_`q���S{�r���,�@Ţ��N�'�@�Oj��[��J�	��m4O`���y�oN�Bϙ�_d����쾮�J�y��-�&a
��%�=�����3fE<� �����+��>x2C�<�"�됲��z<\��YP
�J-mH�ã3����j�r��1	���Y�g���c<Kr� �DS��^B��
�>�E?i��":�Xug������ۂ������s�.�	�L_N�\t�\���բ�!� p�l]����0�cCP�4��+�u�� B
��Leg>��7�I:{�e-�Gn3X��ss�](��}g��dDQ�Oa/�!,"^~���-0Dﱿ�(FBo����F>�6-�U84�ޚ��<,�K{�;v��]ߍe�xzn��?v=�~n���omT-܆W��J%'�ZE,���>$62"�1��KR3�o�z��΅�&��'_ֵͬ�W�3��]�ۛ��������D�F5�7/#\��	��_�$]{:$�S �4��7�'*�jhM���4�{=E0ݰkЖ�P1mq��T�k�{���RZ$�m�x'�2��";�bt)�4�nJ��Fy0�bI��1�o�S<�u�-��o����ԦAA96�,�k��f�wf����u��\h����BG�{�[j��aX�Ob�^��a���L$-RX#D��9�Ҹ��BP�)7�T�{}'�r��O��^qB�X�4ON'g����ǜy�u�j�!�ߌ�Y3[Ce��#��&��N�JK���%Ks��֪Q���!�N�䘫�_t���j��G�K��Z�C������n8�����4�������MNZ�'C��S;?K������K��h�� жK�~��a/�R�/۟|ښ��(zz�+��`��p��ג����lt����mI��`CSq��b"u
_,�d*B���l%�in��h��4��4�w5�a��^���Q�����I�j�|���1��0���R�?����G���9���k_����)hږ����9$0��(��W	QO
�oK�ib%���"����5��nL�n,�*�T������˛~����X�;?��e�m�s8��4�1��6Jl��M�:�W욟ݵ0ۮk%?����%�"���O ����뚮a�#4&��f�*JS�.�L�p��ѧ�j��T�_���T%b��f<&O���+X�d�	��>LVgvJiI#���C-���C�}TE�s�/��H���WܙY�}�u �w��"u�v(������Z2��K�nY�Y�Y�j�r�_h:n�>M1�sM�5z�b�[�k�V\�����e�]C��
�7[��&��WU�-�E�mh��K�9�TH�>n���G�&��(�AB���xz^/�zR���A�!��t�T��U���ꦹ�ߠ(��ã�x!�XUZ��^vKؤ�ݖ	��hR��%���L����4��¤`�dS��y���:ץ}�}���v�����>a�X�S��
����G��[	�*�#��]*Gz��e���S�Z. %$��ж�� ����z�����	���?l}K� �W������T/p ��oK��_~��#�E"���\�[o{��4�[�T/��,Um�Ynlշ����j��?���<�-Q[x��Sq;��5�~��Ca��ڻ,X�!CU?��ݏC���<��>���a�c��y^�}�PD��L��H�K{l.�W����5	t�q(��[�9��.U�O��� �r��3�	<؛i�m���gjA�ʐ��0|�"ӓ�@�PI9�s��|YzL�êX>w5�
�[v3�%�Sd��ݒ����켚��Ϙ�	nwk5ʿ 6�/x�`�x�������!�h�J�����@S�},!�`_�J�M|����������ơS7���P�IL�TT&dwf\ �.�Q���x��Eק�4L`C����3E�(�
�]Y���Q՘}�H���^I�C"�b�˴�H�$az*2E~�aPEFc���N9�5B+�*f����!TS4�P���@���-�Χ�'�~z�BeS�UK�����/�J�,_��`_�m��G^��߬�MM�l����׭���԰
����]�Kq�/�!��7���/ݨ�"P`�z,��ˢ��F�U(�
���ѝ��F��&�E�@?X�OW�������q����?�����4� ��F{|�Ӌ9U����&�#��{��V��kR������u��nn�+�X8�r]��p����Ao�w��N��^'���en�ŭ��N��A��������Z���Qj&�ns���Q��&zu/�$s�
x_x'O��*��al������ �Q"�3\XtF����٥���?d��!m�T'�u��!L�]���<k����=z����ф���ϒR+q��_i��E�K�WB�Q���,4 y�^_4�y�[e�Œ.���-����;��e�\�����f!��je�= ����
O��p�&����"/2%��Z�m�>U%��� t%�8���\t�m����Ԣy��`�ț���푶J�Od��L����B`"jP,R���i/����φ1��I�3g�|yL�V�/-6lb�i=�y�9R��=�wo�S����s��j�E��$��#Kr�AC,MX9ŀȑN�%�Э��'��w�pWih/������K<�Y�p�=')Ɲ�o�=9�����dʹ����4E��ϖ��`[7]�D����;SZ0R�Oa���-� �y FD��/]�$�줜������d�
�/��蔗���;��җ����5�Z��D��{��o4ֵi�'W,�*d�@?��-p{�[���/�)Ǒ�^ �K�����ԓ��~r�<�SD[{畩�Q��K����F����6�A%�h�l
�_��r���x�z���-��E��;M�D�;<B/Ї"���j��<�����cw��U�`�+�~c�~�A2�j K��-W�Ov|W��f{|���U�"��FO����D��WT`�8�l@�5��z��i��Zт��g�d���x;?9��}��y��6H��ꇁ� ��M���1.�
&d��D���X皱�=,Ă�3�\P�y���&��7��I7xDq���z�[|+�~��aε���Sn�w�t5`w<s���O��K+���5o��Q�S���E뼷b�_���P�^�W��c>w#AM�S�I֤k�R�3�f+�-<�ܣ8�js�:�'�a)/.Lӑ����A	��S֢T�@d��88 
���w1�4#�<>}K���x����(��,��[5�=O��[D3�~+Cډx(��ڹ�������}�׮�HŌ�="8j��@U0��O�~�񵸓W���{���־<-���)�l�4vZ��M��6Qcv[�p�(�WB�Z��N���1�d�!�YD5��5��$#һ�7�)y��$a2o�D䍢�Uhز�=��f���fӓ���j80Ҍ�SDOÑ��<]f�J�I_`}4�� �T�:j�+/b�p�Q�s�O{�����-��+�G̕�M���eo��9C�:�>��R��8^k�Q߁Q�"'��?�^�!��/�j=y�l�:�K�P|�_*]WiR�BmD4􀶉�j��m'�PM�j`��J��}��x�0Q��ni��^�䎖�&�K���H�B�q<lO�
�7!`�CqO�e�+�Ӣ~�V��!�5��6vř �~4&��*b��qVe�4�_�T<���Z�BV��Y0�(���;)%�Q�L�m%cFT��{ʶ�ܿ4]���fX����B'~�M�cdaP��:��8���4?�(���ۥR[��a���y٬}SGb�������t�:ca���xv��=;N�%�p.����`�X�dt(��aEk����_�Í%�r�@b��_~��a��`=~1�ёcB�
�,lX��Q���J<*X����M@*p�Ső#H,�\�Ud���QHY@��teB�"�P��+a���	�(� (l
8F��	���is;Vg.�!k|�;�#����2�l���oۓ��|��xh�!�SQ�Q�Q�HƳ�ew�76�m�l�p�t�1�3�B�0000"�{~��;{����5�Ʉ�Q��E}��I�p����C�%��u� �)���/}T�ਢ��r|��i��J�ኜn��/ߦ��i��䬊�W)���|� }io�߿D������
���,�*��",	�4ˊ�Ԯyq�q&����_ȋξ~:�V�^�}`���A �ԭ��s�4�?�A�'Xb�������6����P�M�P��vf;��+kw�M��U�)ة9B����'���n��k�J�}�9R�"�6MC��ٚ)�[����b���Q���Cs!��BV�>����@\���!���\������(`�>_;�t�>1\�UXp���E�=.��`����U /?��Q�PG�B>�d_�?Q0��tBvЋ��Z_�?��"��:��FU�wݗ~����-DE��G#�����"P$x,0>�	 N��'�H�$`�@I(&~�	&��(�)J% � $�AНe���k���� D �68:vl��'��$�5�x�It�t���[��4^���4��ȼ-DE��G#����ݥ���2	DE��G#��������# ��D@K}Zw!�F�*�JwΙ�}�D&���0������r��i�NG�����ՓO��1�?.� 
fU�F�q�f]��k����VC�D������ykl�E�
��,n�κ#2���*��Ю�$/�ܹΏ�Ѻ6f���K��L�+���4L���p�q������:4�lQ�e�#d������n�_.��J�3W�#��y��&<El��&��m)p�a!\��V��3����v_%�`H=�<��y��Ѿ��dx~7b���G��x�����U�Cq%���Q�eyO٧�����M3m���8F]�Nn�D;�ҙXD��@>��􄯏�U�H�ML�ҥj��z�-����Oc)�$����I!|&f<����Fث�o3���-d*�`&����gk�=y�i%�d/���Sb#�[��]��X%�$?6�@ܰ��,o1���ҐK�]U��W�r��<O��(Y�F�L̢��{ ����p�ĺh�= ��]P�N �8p��#�=so~�#��6��qп�1[l��
�g�'U�9������������:9��?��4G��eɍF�i���S�!�(Rq�Ve�^d��⳶�>H5-��R1Wj��^��-^Uθ�?�����,�:�̍��{���'�%���N��{�5�+�@2�4������X��ݳ.���ʟ�O�{�>�ɇ�LU?��܉9B�-�D�UEPr�s�ĺ`�zDm��+~�
ٻq���� ^8J>�)V�c��`>Q!q���C�n1%/9H�l{|�L?�i�̱ù'�O,.Z�WNv&��؁������1��/�V'�7m1F�(���'�U�����?��A�Ŝ�*�nS9Z~'e�ʳ�_��[G�8>Q@.y�����g&�DGJ�O�zr��T�m��-V/I忨ɂ����O�x����_�2W����R/�p�10�+$��9��� Z�8����?qt��������8ZQܪ�<����Ч-ە9��B���TJVU��eA\q��ٛ��j���)o ��U\��D-�U�	k���~�xݹS�-X3@]CJ	�1T|����mh.h���Ay,�1��
7�G��\�pG΁��t�9Q���$��kAUh����T�=��u�s���۬� �D-�XJJR<=�1�?j7��U5�;f��M\y�%�Z
���[��yI��
��;�r�_1N��]*n�x�@Pj7�U$'��(}�����Cz#�n����ޯ�t����������������������������������������������������������������������������U��k�k�k���� ���j6�-���p���&,���ܲ���iEU[�5��]C+a_wX�uRO�8��5����o�9ʣ����Q �ϥ+נK�a2�S��Ք���^*q��]v��w��U�!	�x�/�=b�ʉ,q���T���dë�? < ���@C� LDH �2�0@@e�<��`��fh5� B�@ �$ɀ�"�3�TX\r� ΀F F@F�" E �;� G �ˀ�@g�@% � K �>4�p	� 0@P� `p
 �J J@h %@40VC� � %�4P0�	h	p ��� Ҁi`4�h8�R��y�U������m'%����Q��b����I:Ut��m"��Ke������i�K�Zm�^
T�����i����K�ѧ�L�__-���-����.�|�x9R�JU��UQ�X���z����(�G3^�_F��W�p��(g���b(#��u�WL/E��Ig����گc����BU[R H�Y�rS`���M��(�>Nc��J����ע��m?��R�͕�-��Ǧw�#��a����)Wv�+�=�U�U��^����!��,�52B���S����
��îbW��ٳ�������O��ET�\�h��P?Gֻ�����.�x�%W0���+ˀCé���b�cd��[���32�5(�eI���|6�f�f�&�VR[�msw��{syZ�&�չGe�?�x��t�|�/s�/���ؼz��}���翧��������\�������� 3`�����b8Ǌh�4���2L��U��!�m�cn�:��W)^8�W<}Ǒ��p��zm�ޛn�����o~���~��`�m�F�����,�R�6����@FJ�%L%��?�5ɤۙY\z!���b2N��W���C���)�����}�؆�X�kp]���D�~em�'�ɧ�5ǹ�dy�X�w�M$eK0`�L}cjf�)��.�ⓦ����x�!'M_�gO�bWf;5��ɔ�u�rTom��;�ʁI2��ѩv����􅓂U����6�H��|�|5ٓ���:��y����sVβ[�M�J�����v^�&o�� HI��'����39�F�m�D�ʺ	���f�Ѳ�'��S�d����y}�����#���y��+Ұ�.�R<��T��JÒa�K���lL
�r���c|�&�@������9��(�C���_���?|G�/�-�{�U������d��-�ڻ��I1ğ�"���G�?
�4H>���TUh��Qdn^��Pj":�=9K�2HF)�'sY��ƓƐ�WЫ�YۿŹrD{�v	�M�Ɣ�Bo9����
��}!ܾ�}���� 8��h�!��c�
8�A_E��7S�8��3�$<�ڜ��L45[�r�~t;ᑥ�-�y�~�P֫<V��­B��W.�>�P�;&��Ej��)�藄ao�[e�	:�<6m�‗�D[�H��0��<m�i�=Qg����o���po��ƐG��Ws��G��ʒ��enR9v�o��T �6ܭ��ɒ���+#9� b�#�?�K��ĆL��m怔�%*���[�sPݺ��\B0G$fm����,�?�h����ɚ��}7�rO���O/��ц��:E����Q�ܽ�g���b���:,&��� �����a�4�
C&E����4wR�j��Ga�p�՗G��]ES��H��D�t������1Dp 73o�և ��M�����'���	|�v��~�9Hs �CQ�������P��ˢ�EC҃��C^b��~�=�?�P=�:x~�5`�g!���p�z=�#�Bؙ�P�A� Ɓ���g�BT7b�g�@��@3�t�YE6J7NP%��0��hE�,VjN8����@� hf�H'Z~5�V�&*����5o]8b�gf�z���AG���EÏ�P"�fc@e�Gp�%���ą�G-d�Ac���G�I���G�^�$x"�'d_F������Vs��XR�#��X��+�,�A;����`v!@@�M�l8����-�'e1�A���E�.��}L���-��>�1���� �9�Ձ�ǵ�7el���#�bmj��%����>�
��0e��sZRΩ�[��8l%3L]�^U�	��&�ph^�autPX]0�ں���S���^P��od��h�?�%أp��̪sT�8�-ڃ����al tB�l���L�
u\��r�o3¯J��fH�Jj��˚��u��:�Ђ�©�����nz�56=A��=��NF�NHZB!�ـo�4ȁ�pyC���8�w��u�q�\s�VNB\�#VF����N��a�
>@�Ch���8�
s��s�	H��=~9�	�q��bC��D����J۩%�		`�g�����{3�亘�����;x:t�m�C��^:��9
���<�?N�^;��(�E��?*ƺLJ�VxO��n�9���� 6�o��P��+=i�%KK\S;a�Yو�h�G�[n!�h˫���
5'J�U���1�)���#��@TH�T��J5�ƚ�д�<�XH�4�������떗�>f˥y�B����i8�n����>�/˲�s]�7��o��0obsCe�`��j8
����H�h��J�x�{�$���#�T�M�'�a�����g�L��ncl5���qYl�*���?*�U��A��I�6���r�����A7�'��X��9�n�D�J��v�r3.����;��NŒFƐ��I��Q�ϖ�,4��>����94��񙖋_��݃Bf����y�E#ge)I��g�s�~/����=��u�
[��PG��e�j��:��Z{Յ_�T4j�ԐD��6횰�̈́>}n�ΐ��;�y�<Co���#`o�;/� �A1Ǫ�����~Y=�g�Ȃ(���\0��X�:���@�f������cF�)�5�F�������9K�V�Z�ٟYҚ媼܍���|�c�e�i��]߽N�G�I�����?W��Ѹ��^�� J�/yɮ�S��'�CT�����^�8�N���Ȥ�3��/;��~͖�A�g��M|������銽uټC�e��*I�d��],�U�����	��$�&�0�_�lI��ͽ�Ѱ���k���sD����[�W=�ƍd��e����s�)�1����V����a�+j��p-�����LB�qa�Tď�s�W|����C�pe��Q���o:^0��1����!x�<<\&j(�]��p҈�A���v �R��8[�LnwKJ[�!Ք-4c�3���!V�zs�3��� C~a�֐��#Q�נ
BSD�	,h&[��>�Ξ�AA�qM-�T�����IGtܽ�K[,�E�e�jNU��� .@g1��F��Q���}h�~�!���u=�=�<��|EēCR·���U�IE�����!P�0�3�>��t��y?Do����:�:��q`!b���"��`�:��\z���F k=����*�q:�q�udF7:@��&^�g���U�;�f����h^%��`��i�xg�g	�l�!��'��%�s�X�Ͽ���ە`a����%�p�|x� ����l\̶���B�r8�7�l��Ì �M[�G�!V�(�xd�����q�v��`�a�NS��ArJ�ϧ[�����<���4V�.ݚs�?du�l�ŭ�s�Y��<���� /v�K>u"S�C�9��4���F4�(���ʟ�۴%_�K\��6�,����lGP$G=�I��i�r0�,���-�I�6K�6Z�(�o�Bk��n����~J2��
�]|�Ⱥ�+��r;Y�����l��zC�2b�.�f� Բ�|ml}#O�����e�[l#�5�?�P�Ya��1z.��`��3��&�H4H���HUǝ5�^��^=(L����
:d�U0����Ak3 �K��$�梈���vHHR�����Iy$p�~�ɑ��"O���|ɽ_a��p��������^��?4; *��re�`9L�b�$Ь`l��M��hEx����m'�!�
`�b�����F��y�h����Ǟ��8�Vji �2>G�:0H��$�.fM[A�D��Ő� ��j��kWӪ�r�n����h���;�8%<���F�����X�_�ⲕ������f7�4Qp�h�8����úξξ1r4�v��0���Ӽ��]�8W%���Vc ��plBH�8RCx�C��u��gP ݷ9k�4z�,vtt~ w�v�O�Ǖ�2]�+�G�|�*�� vk=�\����5.��̯��~zx�p���)Ǚ\!��&��c������Tx����mً��.)��+�|��OX���܉f�Oy����*��Y�J�taݿ�����gŽ¡ *o��I�HZT��8�#�/��N���=�����l����Cs��͏���p�}?e��Z����!�X�8����i���)k��LOcx���9���a���O��e������C��Tou��V���9�2.��&�?��<�h8�A�6�T�����>�웚�(r$q���MA���I�qw)͈jk����1���d]}/��b�g��Jxb$�g�^�&}�Y{�yH��
@YJ�m�}Ψ%����T[U�x�:������_�m�3�
 y�V�E���1y'���ی~��DV�O�@|��#�}vv.=i��,�jH6p�X}P��q�#�"`��l��[B�z�~8���.�U�vaQs)��S-$c`m��V�6��3a�%�oV��:b]��L�TV��$���{>\��������K�|iԞ�����V�����K��]�W^�a��F	���\�k���\��<L<c̽��$B&��W�0WV�������.�����)��\�13�{�K(>��t��`ﲯQ�����V�<ҝ�1�����E�S�y�ܾ"���������o����Q���ؒ q�I��m�M>5%���O�-*�\0�a��.Q�#���:!���V�.�كG�\c�T����(��ź���2�`���lAa&o{�����1`	y�}�>3AG3ϥ̆�As����m,0]F��8. ���h[� (j�
6pC�>B����1:�����-�EV9-��YN���Z���-Pc"{7�op�y�BS8CJq��r��t��x�9#�I!��y���"�.��X���Y:��7��}A��ST���e��8��g��\	6O�Hw��Ou`{j�9P��C� Ha�Gu��r��n�ۺb]�C�yt��c��`����߰h�c�W`�Id+H�Q +���q�պ����:Ӄ2H������1�O�o�c)&3� ~�d'�����m(\Ţ�w�86��&������{�H�WK:z�t�摧
��2��u���q�Bq�9*#���e>�O�.6O��R�;�����O�i���1���k�2� �ho<�XA��_h��1�Oҹ�ui���d��|%��s��5��Z4+�������`9Yv"Ct��^�_��b,�F�w�H6�mE�P�9/$�"�ɫ���b�D�7n�?�Z|FzEL5P灣9�P]�
v��I���z�  �QR0O�ʋ�@pb�8Gad��M�0�C9�ۺ�UP�O5�ʛI����z����ZI'�0��W[��N>�f��l�u�!��~B%˄Џ\��cb��i��/A���$�(a�J������A&r��,��ɣn�#��lɉ�3��p7%0T$�?8�{�����p� �4��GCa�eW[I��ϬuH�,8���3d�7w���qo������XS1�ރ����<�����Y�n:�$���L�!U�c;n�=cs(�zI�8���Q[z���J��׋�Зn@�L�[�c���/#�����Q�w�#�H��ӄȷ�SAښV �K1�bí!�M"-?��i�f�/�M��;�Jߍ/>����}�w;�(�^8��w(�B]b�X�tT\:�ߟ�'H:���M�{%���|�٠tg�+ߡ�H���ƬY[��6�p�=��3�,�=�a51l�A�$���ZZ>��_�g:����kQk�2���O~�-�I�hC��tg{�k��������,DZ'�}��y|2~����� �7��%ఇ���ͪ��PR���%�Պ6�����)���/���mBAQR�gûb�B:�'bFו��s&��pGm$(L.�٘g�R��ػ�d�]�vB�I��V�P�T>�����+]3���)ԉ֚[1���,}��;/��`����;��D�c�J����bD8�^�@ivf�<	������0jl�㽾�����Eg+~\�r2.tG��z��7pi{c�����i��'��z	D+4�,��H�I|Y�^��r����eO���p�U��:q�4B�%o��ȷ�YY���w`l`���Ao�ld4�ŅJNm�O��ä�:#
3�~���u��0�&�Q�L��K�x�
1�q�l��>�p�߾�:+�[���]�=�홗��*���ḕ_oO0�?�G�9�4\m���ϣ�?�zC��LF�i�qρ9�5���egEל��I�2OA������Z2������201�:���.���ض�k�GGD��\�_� "��WT�G�5��VD}�E&�S5�|�/�*?a���w�Pϩ6��@,prqY�Ɋ�*��6��m.h�����lh�J�g!�����)������]�l���9(�zd���%!$�Q��#�^�3�fNm�ΰ���Z��ʖ��|b�XO�oWIxu��O��(��~��E¾�d|��o�7���(�Sx��m3h'6��}Q�dQ�Dsc�-P�CVXBHP��)H�G�]�K�PIK#В�dil-4$ՖrN	8�E:�����<HDH.��r��[�Z&UBt�_j�(�,�V{����+���i��FKϺ��1x¾�3���|�;+����/g��W뾪�jV?�X�Ko��Ay�k����=)M �'zJ��qo�,Y��Z����F����A�c�8�t^>��uF�gkR{�*���͕�x�L�{z���2iѹ�G�[#��1	q�G$�TV��d�D6v[�,
PZ��S�)�@)�C}�&49b�NZM@�Nd)wh�nq"�e+��b������F�ӗ0�q�ɲ��S���=õ�?�AS���g����*�#^g��Bؕ]}�\1,(��S�_7�)iL������ ̓���dx.�����*r�KT�/J�ۣo]��& +���QYg�q���E�,{���*��nB��'+6��}�%�q���]M�iR�X��[x�T};��#U�J�@NS�xr�rp}�~N�P���Ә;t�����f��A�Ό��0^w��b��K�Ub$��#�;H���݆nEe�o��?++�N���:7t�W�!I|��qv�V�P/�F�D	LHGo���6Z�n�^CA
��֓�_��]
K�Sz�����C�X�:�hx�k7ದ�]C5 ��
��#��b��`Ť�V��Oa9Q�5���@)+Rj�)GX���Q֨����Q�����w�v��=��O�l��,UN (�F^��@�Q���?�?����a��O�J���V+S��K�۸����#[��د��N������Ȉ��Qҋ�5�pp=R\<�9<��@�e���f�k�&��I��~��՘�XL?��ǲ�K]x"�3_���+�Je~�F�"�c�,�3'�����>��1!m����/[�A��K���z���~fҍ��z�3r௃c ��(�؀_����<D�g��9l�y�5����ݼx{��.��QP.�(�V��!w�\�/�t��9�JG�T��ڮ����9:ܳ`+��D>B�Y��=I�3M^m��7���kA� �ӷR<�xW�v�������AS��L�~��f�0��Y_UR{(v \���,[�/:^UH��Sc�.{\z�u0�E1f�	�O��'7��*�F��6�c�vq=��^�Gò��	ā�,�|���k;�#!�?
��]�V8�7�D��4��g+����/u�����ʹ�*�@ն��f�:zя����'RF�ws*�M����BC'Z��nZǄ�r �"܎�����_2�ȯe�����NF�>rZh�!۽F�8���Ƅ!���G�1ď��8���oAF졽�,!�Yv-\��H܏�7��:���-�߿ZZ}�I�\�m�1��c����Ҹcuk�g:�\����ӥ���Z<�+P� �e��;㮊ɦ���d��	��˰�Eu@ ����9i�(�	<{|���m����l$F�o܆U�p�e�l�zEÓ��J巙��`>��|# w(>�3G�u���a!���������#az�9U�$81�i�������2��"����l����3d���ɋrL0��7�����"W�4P3�=�Ee�?�Ɩ�	����(��w��$y�Z��@���������}��\���.2Q�b�a�$D&���Z��C��}[�iFl|Y�r~��>�!�"�G��{��nb�д,�Qm'��Ȩ�ޒ�)�a�����[�g�A8?�5����foVAȗ�� ��l�dU�x�e�ݴ;�_����~��D_-�/JӴI�b�ޅ�^��\:�|P�c�}�	㈱i��&r��O��$?�K����x��<�vi��+s(æ��1��O�+Dvp*`�C������RT�LY4$b�NH]��S0��BHgd	��p�6eͅ3��:3�a.�Xfɣ��y������1<��^��
I$̓�����>��ݫ�ᔨ����=��H'���r����w���y�����-W��p��8����&�TU)Y���	>,���/�U	����l���\�~I͢���X��V�Y��q/��u��T5.н���NV���gkt�{��s(z���7X+�b�����'�׉�r2�[,�2d��<�I6[p��/m�/I�͔h��CY�WoO��%��V%�X���g���h�u�l�oË�>��>�x���!��P��S�[����8�
W�X�����]�" ����L�Oh=uZe1G7Fקf�󜪂s,GE�:��o�/pr�!|8���3���m�������X�s���H��=ŭ�S=<��xDt ܙk�׵V,x�PjgX�����z���s���ޝɳJ���H���$�o�'�eՍt�؁b~��w��t^K���!?�w]�J�z=���l�PXA��ւs`�o���H����>�Ē?hK��'���X����jD�#�)�RDK~�����S�3_L��5��{����nent�-O�%^�\�'^^* :�~X����t��a[�_Uٰ������b@�x.8�)L��p�C�)���?Ǭ��&`��e�3��1ϹSj���r�T���������<��涴K9�I�E�΢�u&]~Z0ɛ6�9��v���Ju����o,WX�^X��C,��H�>3 f�2��`U'	�5�^���O���:�z��D;����TN����p1��'^,��hN�RN�����5��^���M;��b��G����uP��/�u�/���k̘{i*�yqk�NE�m��a����lRZ�Wp��CL���#p������Mg�i:o�(/�?�9��d��5m����E�)2�eg�z�5/��q�<|�|���O/O�ӝp�jH�����2�� ����q����������]�ͫ�R.a� ���_}�	��3�u%Ȩ�@�pT�91�F��* ��X[�t]*��ʠ���Oϱ����#�����
��!�ڱ����/��8m�]N�����$C
����O�H�V���B���oD�@����D�L�nJR��'Gi�S��m?�i@d�N���)/,��o��|j	U�$'�y��C��(��d;{+�hX�,��O,�I�Q���@��4!j���jE�������W�NIA��g�w/`GV|�o��3j�]	�&��� ]k�bvk�L}�d�P��_k���֧�л75���F�ػ�YT�p��\���a�k�o7��`)��������	�M5�U���+�$�ߙ���I$�A�"��a8����$	��Է����͸Bf�!�?����WHL*�$e�^O�_S��}ĉLVR�,�aW�F�#�w�C��#����5��a�:Z���Ӄ�P.HJc�.�L[��B�ޮ�����m�����VM�9 ��0�����̄�k��h��?L��)�ɲ7W2_�����FϹ Q ^�C�>A���V��c�����yuˊ(�� b~��5ţ�x�[
���؞�g5w(ќJ�6��FId/M��כ�B��<�^'��`G�l@��푅A��b��V��HN�7��1�מx�TB�Ni(�GWJ�K+�]ɾZ���p�oN�
86m���2��2!
g��e-�S��}X'���Kj#&�&��Ɇ�	�<	����/���
߯�\���̶8O�.W8b�u�+�!0�7c4!l�>�l8V>���=l����=�ê�&5������c�qTd��_����#%�vߺok�e��¼�ПNCMxS� ���t_��-�c+fdmZ�g�Z�}A������8�G�	�I�E�,g�Ĥ�ú�d�.����O��èlO���*��7��m�����ϡ�����2��t?�R�X���.�c��B�)�����łx|&��}r�r�mt�Y��T5x�!*L}��h9�5;�>�ky��uv]�EAV�z��`���.J4nu�ϳ��5x���!�)_3�s����^�ʛ�:6��4���O"[i���R
�̦�Z�7�X��+�U�m_>5KW.���n��х�u��*V��-��������@6�\��? ݘp�vĳE�1)s#�6n���G`$�9��y�e�즎-7Bu�
�C�e#ȵ�ӝ�Xz���`�3^� ��!��/`�"���Ṳؙ̃�V���2�T���T_���+���~
�r\�;d#m��\rр���8�%�6W�!=}3 ��T�L� � �.y��7�2M�����=�{Y�ΠJ'pr�'g}%�`r��+� �uQ�A���k�;�5����+�a�eL%�%�� �l�W�5 ��mbq���'�
\�߱�����|Ql�c_����x}sL�u�WE�l@B�ʿؓ}}�9r���!��#��`��B����[oY���;o�,��=	�l`�A��Pd�����R�(��"��=��������1Y���;��v��xQ�=���z���		M;w�3�\#E��tQ6�e�p�tA�+
p�V���r �F}�6 �w�%L������R/�8���)�N�v	_���W�1Cj����,�����>J�gPf�h��6��	f��m�m��6�E\�G���&���{΍3�C�̚�>!��,��{��e.Gn;4-���r���Xz�T\ZG�6�����^ݑ�=�(�"��5���y.ʢJvY8&�S9()��N:���sN`�<�q�ۚ3s/�%��w.;�Kp�Ӆ�Q>��5c��0y�?���D��
�ﲀ���Hv�nȑ���w�w�A.r�F�]�V�«h������=���:��o�!����L�HwDWp7�Օ��rr{�W�9З�M��~��8/���de;���M��͝'�ﵠ@��Dr�6���冞4X��q�d�RE8�����]��Z��NRg�� Q��o�}ԗ��GӰ��d)1@�[(+̈́qY�W�m��Q�V����uw�O��ت�E
���..��}�&���Oo%�˦P�!������$I�LZL�!�^��=g����X�ܶ	Ǣ�	����ow�
��љ��f���������^�mI�$
da��;1e}_�c�wn: ���'S��Ln{OW�� Z����Kf/�o�N��$m��|#}�Ϯ4�;|��2�9;1gV�V��Nn�\��	�tc���A<;��ZDbP�f��.�B������F��р`�|Ɠ�n(�NN�\[�*�VY�,~BO�<�D�!�a؂��zc6&�d���z��MK l�� �+�jT�ץ0F�[|t<�%%x(�{�O��-^�����#����p��6�������3�LU>�u�U|W�Q�˞�k�b�.쨵6�Я|q�i�G�$������
���m�Q)��\>j/_!�D�xgo������_� �ZU���!<_�\��rodÇ�Ǣ�b8���ä��*�\��lK ����e���ؙx{��np����ax �q��G=�PX��l+y��b���p���K{y�[�Xx?Y*�c��J
���W���@����{�s���d�d~el�	�節M�&7o���o�j�&
R_߹���R5�Dg\�6M�k�L��G�����SY݇���`h�K�S��������s�5T��ǡY��"��>4�/���v�e�É�Y@�R��s�ӱ5i7����Q[�._�6�WxE��������$���N���	.�C�kn�u�uW���}â-����N�����^��,��>���.{��ޠPU�^�Tz0H#����W}��0s�2{og(���w^p�yO�����d��_��:���}=����D���$`�g�Gj����mBn~�k�3���#��g����CbǓǆ|��QD~N�������q��k��������L}-sPk\�B�J�L� ��,Q..̼j(��':��
Z�X<���oau��z��
l2��,,�J��"�Ny�=O7��Y�Ƃi*#��^��i�W2����t�d֘|�,��"{U�w�R ���m������'�����$�Һ������}��c�wNp�d�����٣�����I�Dmf�%�7�p�`�?�觍��2:[��s,�0ʨŷ:D	�6��������0��M�����ͦ�3I����f*[6ws�b=���d���X�[#�^4+�!cJN� ��r��Y4��8~����96;����?��_	���̪@uK����]1[��e�+��Z�M^]����׍��ŧ)�u���˞�e��N�/=����9���Ͷ��u�S��������H^���8�r2��Sh���l���,��/��t�6�6���^�-�ҍ���*�Z�����`�_�����ӟV
á7.��#��L�8���Q�o|�U_��`g�x��bHi!����ؔZ�	�؍z�r�����uʊ�=��v\��3lq��D،�j~����q��� ��;�l����=i�Df�9nwV��.~/h�su�믡���>r��tY�)~Qh�G�?�G��z��"C���S���� �G��|��A�3V�3#
�̂z� 4�5~w�OV�ڙ)�Q��nS��1���Ntnhv(#Wcm�|p�8=�;�U�~AB�`�*�+Wc����7i75�^�5b��0��c"�'7��%*���v�	�-^r�$��{� ����|���>+A��v	��}{�O@���6�ۿ��(f���@�^&N@��f�KONP�pJ�R*�h�8���������M���K��FJ5 �����Q�|�{d��Wro����|]z���PV?�]��M�{n�K>����J��(�,�:��S+���q�9���2��Uc��Q�zd�R6O��-��AV��񋶀�x/��������{��Q1��}~�q�-z��}�V�:�n���v��B?WF<�O���i��.&�<ѭ��v|��]���*4ρ"u蜟f#�g���:L�	��"�Yu+z�*�������_.�_7c�����x�]B̓|�|Y!�wF���y܎�>_�7S�.����M�!�1��p�	��W8(WgD���j�7`.����9x���M�
Yi�^(J^������h7��1�d���4���_�Oۜ��-i� ,~�
��j�� ��%!�X��ۚ龨n��.��\n"�܃8ѐ����Z~�������R��>-A�:�ɾ�`�2 ���A7u���ú.T�!خ"���^�`�2�q�z�l����p�$�	N���B��Gzy^�#�sfb����b�!�g@fƘ���G���L;T�P�ʤ�ǧ��Njs��`>�D[�<�>HI��I�������Í�4��Iئ�¸.�S�~Kٻ�|N��?r[�79D�(�Z��`�ϊ:?�ѡp��d�_�Ua�{��{���,M�_�����8u�}6Sk��%t0j?�˝ޭ�
�n��Ä�"�Q�O��-��ջ����в�����d�o96ʎm���栺��Ϫ̝� ��ǉW��bG������kH�l�VR㡪iT����'�X��������k�<��/�q������k��/v�.+�Y�
D�z���4�ƽT�Iu�M��4_V�� EQ�N��Ì�(d��ֺ���
�A�p����<��I
)�@]Ttt2Sɨ ��F�+�l'%�oa\����J��>�j�w��M�6R�Vy�H�@1����}iY�����&� ��/J�0b�TUCm��f�ƣg6��P��q��[pq�oGR�[Lm�]"�ݮ�ġP�:����]��]|��EIU<x�06)��|���k�g<����&��>��C�[�-�]*F �H �3�&�h�`Ͱb�?��;����Ҍ��v�N���3�F�ns��= �k�-T�E��틶Od��1>�ٳ��vD��v�`�z����-�*���Ш��ASh�jܤ��#uy&s���cBq�#�-s���츬+�����}H�z]{|a�l�v;��^�w!i쁡4l|S���|�O�����E�Q;U'V���~��!�3F�~�y�Z����Y�𑥬�u��J�'��xn�_���
gۘna	��+'�C�|@����'ퟤ��1�*<E��\���/�b}��*�NG������4���<�)�?µā2�"}��F ����4�V��m�g��Bq��0B���9H�I�����T�ګ����dq8b�z]�W*�� ��O�?�����Gw4�ܩ�E�B�0��vb���{=��!�7��O�O����!j��
�P�:�x(�����`
�(mBe�{�?�]Q�#s>M�>
)��0��h�^G�j�SI�Ց��I����B�oh5nK��"[4K,�:����v��Hg}kŶ�'I����cnhrW�\��F��� ʀe�; RC�H�>���o-$�	��/����b�L^CPn�s�R�"c�����L�*�e�p�%I�r�Fy0�V�n_#�
1%�0��&�7ma J��f���<r��k�ʠ��K�����R��ʋ��WW��}�묢:-�����m�Ukg�0~�C�>�v$H �W���b��p�+�J��&����6���I�����8/ں��O���G�Zz�(���Ob߼V&���������\s$A�΄@����c^M�e*V�?w<�A0v���X��mj i#+�/���E�B�ɷ���?����Q���=	�u�z�W%�E
�]�C ����Ea�rN�%N�V�����y�z�%K�qا��yt���Z�n�Bџ���ﾧM����_ �^q�J��+���|+�O����:��X��Z�<���;,���h��Nt�J� ��1���,�%������t�tE��Ȳp՛��-ܐűg!y/`�I��m����Rw;��w֏RekR��u�7�q%�+�O�$9�F�﷯�)�P;�齔Q�~�_ۑ=�kkYE�z�&�0�[�t��(���UKY0��JЃ�mm��_��wN�[�i]x���^ {���{.�L}��SA�l3R�u`K�NP��o�����e�죓Nb'�b/.� ׋JC��,RK�3�?�e ����r�x�"5���%�t��<�J����س��O�������@*��ii6�'�mz�E)-�,\e�B)I��f�tQ�tA'I�'��r'N��|����ˁ��8���l��J>X�"a{[��)��M^�4�=�m N�c�:��*�"]|B.���^�|�$�l���W#��F�W�"R���o��R�=��K7X�[W�4$}��Y�u6
�l�E�4`�K��8���=���wY#aq�=��HQ��;�U�mZ��6)�A��"\�������h�"V��_͠�V�HB��UWw���c���IAEg�{,TمZk؇Qt��_q{Q�{Y��	�-�C hz����`��}ε?:B'�u��U=M���<�[,��o{����]fA�7\#P�8��iu�8�{�L��e���Q����f�k��9q�
�y��S� LJXU����
L�Cl��@µ �ʹ��c���R�O��b�
J��}�[�a�_W���Ӧ�����b�&7C[�7	2,?��v��N�0����a5��"bT�"Di�ď蟬 �ZL sM�/��t�������_]ӂMT7:�U�_��_1�f)���>��>���yճl���ߐy���aXՓ�Fb���)����*�����V�?�����
�D=/g�G��qVW#0�^�����=��s��:3dm��_B�M!E�m)�����Q����`��,��2'+�^�L|�����L�����P���'i8���Y�ۂ�Z:�G�C����x��e�޹ԃ�~Y��8���G���"�qg娍�z��i�G�I}�z�<aZ���%�0Pr�}��R�ݢ����n�S '���i�R�k&�t��0��֕��_=s>N��>�����n�Ƅ��V3D�s�|��H��T��N��Tu�J� :���Zf�Dqb�!����N�U��6�,X�ԘP�:2s1�%J�w���
\NP���rוB�W%�� LՀZ.�.̯8�;��h68ڂ��R80� �J�bu�h��kB^(~{�����?ʺ���,�M��"o�Q<��<u���r:��KV5� �/��s��0�L(g#�3o�J�gA
o!�Kq& Gĭ���W�wͩM8���P��9���f��Y�}�9�}�����()��$X�����f��j��B�;�:�*�Cś�����֏��� mhE��ކ��@�=Qb�^�P<YN�?�T�g� Sx��"Ϛ��1v�6qE�'�Ȏ��R���\�b`n�y1���0x��o;9�� X]K�rw	o��{�}渷�dE�d�� ��_�c"]W�L1�	S-�&��#ϊr�v�P�,��-�RW�:]��g�."Κ����j�b%4;O��"��@@cj��^�,$���_?��c��4	SԄ�F��v�~kYl}=���r��p��l+���)�lOjt �{8i;bk)��ې��=A�&D<䟢a1_X�%.n\b�I�g6?���a��Kǃ6b-@�CWC
�5$E��`�^�� ����C�L-�Q�.u�|�_Q��1�0�#�S��<"���j�	�d��R{�Q��G:�2h����+��r�����
0��E�&�0�f\S�b�O�evfS]���"�>^}���ɓ��W�zx}�Q �Í��Y�6�"����UƲ�x�5������l���ǰ;}�#TX�K]����<����q4��>k̽�h�S�(�G(=,S"	
��oD���.����-py�'����ǢTʏ�(���O�>͂s�6�	��D'A�b�o�63��_���J���%a�h�!�;-fS�~[̺\��J��¿�٪W��jʔ��4�e\m�kv���E>Qb�Lh�4<�'=���cK,�q �?�w8��&����'���;�R�OfDV��'��1��Y=�apJc�`9�;���M�l�ˌ�~��t��fb��+��C�������{P���:p~y�D�3q����z+a��|L��_5��h���]Xɐ�Ũ��itPl�c�R-[$pĘ���6(���@v���Ӱ~�|��-ѽIM!Љ9j��|��b:��sލa\յ���܄C�mfC�=�W��mm]2��x�xw�Ec2v����:�*��-���ۊ�TtR�d��:��;�Eʥl��⃴�5=�	��T$<����M$��.��uMJ�vvE�D*|�n ݺ��N�����I�4�f���K�{6Ⱥ�f�	�]���T�~�"z�<�O/�DD���xpЄ�"��)�UX���g:o�w��,��AX�>��i�=�jYי�A�sϟZ{^T��{~O���_�=1�0K >EI�W�k��s]���$��p�Gʷc
g�W���e�݄����NFz�!�F���x�D��!q��RtA�����e��H=��lY��w�\V�{�~a�C��"q?/�L2yL'g�=�x�Ƈ4�y�lM=Lcݴ��:b٧`~pz�ҋ��E�5�#�W;{v	G�
a9�?�g~��$�P���j$'�n��n$�O��,{ƫѝN��yq�Z}P1���L�i�ۏj�C�ds��--U�H�,�t9JC�*Z�lZ�h�U?.���/z�.uti�u}���&��d�>]����Ā����jh���5VD�X��ԩ��S��N�Z��:��Qd�?�ڢ0�=:s,Q5[�)
M,l�ZM*!)��%Rif\B\�Z���n��n.`jxm��8��	���������ʴ��O����rUgU{J��R��X��E��b�Zj��WM��EH�;AO�)�Yp����P��i��}E@lfV�%��|m��[R:LCh�q�*�|���P۟��>�]��(�(�(�)��p�tE��'3�'��BJ�<��CMp�y��9 !��#�Cd^Z����A� ���\��ZӀ���94(��oނ�l�|r���10?�{��5${��E�j�Wzp�~[a���T�ހ��ya����73��4�^(�z��[c���������\���?+`��S��B�|�R���O���,\�j���n�w�*�O��-��^q�J�ɠp���������v�U��綖l���3�*"�r[g��v�_��X0'8R�������Q�-�h�*.�l)�A��k�k=�C�0OiJ�cu6�꠬»]�M���;鵿t ����t:R���*�:�s����Ԁ+��H�*j�G��O�����\)�����PR�R4u�����G\|_;5-~il���i><�_h�x��a	-�A��Kx��)�EmQ��Y.��H%���[�.2a?	�%=9~���M�cNs�񵢱�.E9wX���v��`�?t.�_�D)���H��1�yMNzU�`��̆<t�`]7_��=���/*��蜻�rɌ�8����yl%��l�q���ӓ�m�K&ծ|��:gɩ@�4�)F�\uA/�Ԛ8�9�k���R먗إ-�Cqt�(����P�9U�њYa��<�q�C�!O��:`hq�A��q�_�;j�9q:�Win��Nt����Wv%8�6����m���wOA��<N���U$v�سJ}�r��u6�}D�7d"kaݨ""����"E,�T� 3E9h
b�`�M8r�@�E�	㼤T�Y���E(�y)�<�� '��)�kiyS�kR���^�O��c�9�G��/�FZ�%�'F'۹I���E�GHo+@��|������rx4t��j/�CC���>2������{�/(S��{m?�MEo�����S0"��r���=,oK�`��d�-j�`H�V�+��Ʀ\�|�ܣ��p)�$���g�u�Uִ��V��3{���Z\��֪���!'V���:J�ܠ.r`�=H��S~�䒋����q�������g���QAG�V!5/`�R��d*�6���9�X�h|]a[�FT��y���?S�<�[�G�H����`R�r�aE0�?R��$~���8B��\���h<���Z�[����ϫ$��:��������!&�f��4ʟ�����i�C��`�d�ko��j�i"1*���L���v����(cBM��I
�I�EH�k���=�����ΕԼvf�~E1r3.Y&��s\���>გ�w��8�~#�yPy>N�ѩ$��
UUr�=�W�8�iF
3	�¾�<+5��M���q�Hqn𰺃~+���p�h�뫾�В��z:F!�I�#���CGw%&�?� C�ʈv�VCS����(Sg�Rۦ�ܪ��7޴�]�U�j+�V=�59���J��$�K����9����w��J�v*F�j�5S� m�)��<�0T �c?nrz�o�͹�����1̈�1����CC�?QC?y�`tGK��\�+���}�#ZQ#[<ѝ&m��ӰjJ%��|��@>������;Ol�S�ɉ��mU���f7F��`���|;%[Ysk����:t+0k6ÙKh^P�Q�37B�~�*�6an�u$��S�*���JhP�y0^��]e2�*ğ��iNA����%��/-�
�s\%�'�l'�䊊�qD�U��P<>��؛�ޫ� �m�x���]|�'�������B�]��Y��Ik�/;ܒ�֗��%��X���>KIw-HG�DE��M=&m6��o�68�L�H�F\�Ӓ�`���F�H��1*>��ĭI=�����W��9ʒ6�CAG��RO����*U����F5���sF��V�"��o.�g�{F�LRG;�V�"'>������,�,j:v�2�W�J,*�O3���1�iS�㕉K<K@4X�N�W�<B-��8m�/[����"A����T=E�6���n�U	~�#;�(qQ�nd�m��
A��'��	�f�I�Z�F�	Q�4��!�{����=D�di�n�ۄ���4W�����l]m��죯]>#�b �D��hF����l
`zSY9���;���*+<ޫ{B MD+74��l= �L��4�9�a\vw�Ĉ�a�w�3(�)�����o`r�
�|U�^���x엲�2��$<b���2�	ׅ���e
	��+n�|�~x+�6��6�ujE���y�cE43զ�F��P��$�a�F����K� ��)|W��E�w���XɷFXL�w��
�[|��$��ЭH��������bЭH�iĳ�m�x��>j�ճel�Z +9\oe���t��՝~�B}:K�/���B�ݷ����Ak�xÏ�_�����+7�I� �ɸEl*5$��.y?�[�e�4��eg�p �@������K�h�~���4���TE�9�s��҅��}j����H8*1�U��R���g�U�2O����{�ω{ ,�/8"�I��<��c�	�C��-�(4�¡Q�eq*Y��Jz�2�2�N[�+��Tc������(�;_��O6Ф�c�]��fa��ټW���H�<���tiŕ�X�(E���z�8��z��x�r�#ɖ��>�����`��AҬ�|SϷ�3����
ͅk�Iv}�!���p��Z����$|[�%^�'l0Wz����Tq>�|#��VU_��
E�cN9T���e���F�L�g�GVl����
L4�>j[��9?B�Oy��z~���ΆE!�S���ƟU|�vIc�x�C&g�������#��T�k��aPep�8 �JA�����xJp�P��Iŕ����	+�n�݅}��x�Va���=��8�0ki�����C\١�(��	l����7M�Ca�nǅ/wU���_}Rh�T��T@=TH[��SZ�d�`�8��ƪ�D��w�<z.��k�}9���Z�����/u���os�� ^J���1�����O�0�%gk{���,�)i�بW�S�kF������O�gųy|�	�!ЕZL�cg%�#ɾ��9�:�˚�F�D2��J�N���;�m���]x��{L���+2��/�_'�~�i"�I���. ��v>���D�T����!uGRJ
��}P-/�	�;&�5�*�6'd������˾�\�99� }-��ҕ����џUa�M	4)s���b��H�r�*|��y�JLj2�u�8�kk~^@x ��/O��{���	��{�wp���s$��Js�̬����\�r5]c5�[d�� uqɑ�&�:����5m�"���LQk���w�yiT>�/�h��M���$�C2����+6��/��
�"��QwDa{�[�[��y��|;x1
�ō�S��(��-�|Y[b�"�K�C)(�NnF���}YPhl����G'���=���\���۬�k,_����c>(QC7kԛj��ob�肻�-N5��A~��QUd�9��Ongǚd����=憋18񉟨W�r�[$u���H)@pԤ��l`ۖÏ?_#VO[�~�^�S�mt��,��3�������}����:�1@�R�f�i*�-�u�H	RI�fj�7K�^��C-�)��N]�d
��TC�����ph@.��5{ǹ3:�A������:)iE��"]�ZC;;t���gD�ᅻeU���!�kc��
ĭ֭A!�q�#�Cz|���qg�w��hI^����JXN}~D�bhy(�Gp�_��|r�L�H%gHU�ܑ�3Ue��ظ]8Fu|���&!*߾O
��{�K�}u�O��z*����2�/��qS�08����.)>�t�@� �4��t�;|�� ?r���h���t��h�
B\�x:`�\*�:e9\gdb�l�,j�#J��>�Z;)�V�I�`�v2Q}SFV}��F?�Qz:�N�:��smy�_c��*���'o�ޓ��ɔqG�<�.u�X��6���ޚX��m
-_�s5o�X��ѯ�1*��o���y�,H_��-��k䳏��� s��
i��*tJee�~}W�f*��w�~*ڤ���辏 ��1�+ڑ�7������j�Vz�'���߀���x�U0�cj��4�=�aHX>����ÀD�u���Ɂ����������a=�$-!�Uka��?D9eSZ���Q����<a�Np����\��}���J!����(=(��Ȃp@�u�0��ic]p�#��z:b@� z8zPfF�L�/�T�U.�CY�k���>`~h	ƃ{pEw���r�Jw	/~j��Y��
���\��A\1O���Q��� yF}*����XN����y<�UC����@��Akp�	Y]�B�W:��5�� �X0�B� ͙��<~J�DUഴp����A���qP8��Ձ�D)Tuy �R��l�'!�`W*����fJ�h�Z!Y�����Uʲ�� �0@,�<U��������P�r�L"]V�?L��aą3�ۊ���E�� o�������D

j�qĤ����������&[+N��|����C�?GM���?�bZeH(�q��ucjlsI����=�=�:i����� ��@}�v�G�N����D>ܟ���/�� �!��5|9���G`��0U�o���$-w�g��B3}EU�AA6 ��#�p�9 uV���C�Һ';�}��&#U#k�����j��SI��6� �	�4�����(�T�5[F��bdh7O,�I�CA�|n4-��o3`h�mC�,G#��d��"�W�V�������=���9��$P���h*���@��Nn�����r�I~o/�R��(�(kS���aM�C=4
�E�29£��]�>6^m��̬����w�4��_m	8Q|7_�r/W�^��D{��r�o����b��&�s]ݛ�Y1�bބ�{}�4�I�7�¶a<�xgB�S�)�w`�wsf�e���_*�}n���_Q�л�k.kE�3�[�ߖ��W�"��������j�߃��6�����O��K+���NC:(H��}�c��������塞����r���x�T��J�.8�iG�EN��܉T�~�����#xؖ������n�bI��1#���S��s�;'�����Ј���� Q	@�U"��� V�dK-�>������m��{�!=@RS�g�⎔1OS
Bi�>Tf�:@���k��tp���5�ؓ��K���7��ϲowW�CdB�W��$�Yi���T:�u��a����9���~���������B���I�B��s�+�x���l�g��N~����_��� ��r���BG�K.�a)�#���k`_�<0Ʃ&"����2�A��x��'T���Ye
�e�A[���xPXK�>�َ7uM�ƀ��Q6��aw�r��hB~r��u�9ܑ�F_����2+oR�0U������KY����hj���lM
���:H��?���\�.� ��$7`ahum�s�*lh�f3���h��sE8H���=9�Z�"*�Z�H�	��mS9x���{�3�蒈����{�I>���w����KCV�Q�E��O�AY<�>����F0�$:'"0d�A�j�MZlrQz�)�_:�gJ\t,ioB�ԝ�Lv�`/x6���K���P	�o��opK���-z��<-��4���9���K�b�-�|���9ci��>v���,�p�������Q�)8��#�ߪ���L o������}�c=��g�@u�i�m	@�`ɓ�2>��%���C�x,��$�zSW�a,3��Tz����ݱ����'�"W`�����6��+ -���0�Ŭ��
Oʌ�}e�4ˮ����ݸ��2�	(��7]G���6ͽI�q��]���E�^ϱ��8o�1��¨Fb݋�Y�K�[��(���gX���ȳ��[�2@�sW!c���@��
`Q�Y.sy<O�؎|S��6��P�,&Z��G�@gu��K��?f.<L�v�>R��4|���*p_��l%Q'J�c˧lM����g.5J���+nd��i������
hg=�u�u�$vP�o%���x�HV��p|T�I���ʊ�C�I�9�L\�4�=�.:B��	�p��Q�_��J*�ay��K�Ɂ��N��SD���^���Cy�;-������c��3�fs��
?�Q�L�M(~p�%�!ޡآv;BC�o���u����I�����:1���5�lX�
�{9�d/��k��u��Bs눔�������%ߑ�+H��K��ղ�۟_�!���yH��T����� #H}��;85�<�>\���L��<%��ϲ��n�
_����|�d�e	�z�ѻ��w���{��>�����Em��U�#k/&���ɦK��P�{����@A�y�V�Ť���Bm,�㵫�1�d}��,/=�����{��7aokdr\|g�5�����cy4�蠚@���5�&n/F�@Qq/NK���~&Ds�Tvť���ȁi��.�����e���gr��64�9�Ƣ��V(�x�d�� d���kaw�F_���RG�g�V/r�V��������0���C�	�zkA-@Eƺ�"Е�~��9������������+���V��φh��#ھ�� y��eEX�$|m�#���l��ӏ�j�Ѯ˛��
g�OhgFJ�/�=/�>����P��������[:��/l��m�I��wZŴ/@Z�=�&�]O�9$�q���c?4U�`�l����=W��D�ҼK���B`�H9lZ����1�q);���� ����;������l�a�\m��0Qgt�#�|}^�4<[=����7�޸������҈	=nt���$���BQ�EL2dފQ%����<�!�&��K��9��P�������B��R=�28��޳^-�p����� �qK�څG31ӟ =AB�fOׁX�����Yw��iU�����ӗ��B�4nyS[x&��J!ms%eDZ�����k���=�r���������>=��.ۏ�r�2�>������@�/��*���K����r5Q��w|��m��N�7���ՏZ��Us7�O � R���
��x>0�D����]��v���ֻ�����.��[�p�}[��`�qe�>#�7.S��_Y�$���"y�T'�2��f��[F��F#m�9��Y�SWx�3u�1eWo�W]x�����8��G}�Go(�}�]3,ڝ�S�O�-�4[�aSntj��^	���Lf��p��ȼ��(��ixQ��'�UDj6_I� ��
�p��[/Lw٦���'����l.�r��GX0�Ƣ��<���g��>=O��������g��`�Oa�
�'�����]i%�z��V�<��ģ��hN;�Mn��ϳ D�tي���N�������}��cl�����q�6,���q�d&�����<HS������s&���q�a[m-��}*�me/�0=�9�(>d�A<���<$�g�CQ�xr`%����4��&���kh���g3��j%��� ��ЏGM�=F/�&*�����#�幮x�m�� �ٸ��Yn�c�h���}Q�rTi�u�!&a59��]�򌗁rc�x���a�iw�<׍uF�6{��&tQ�Z��eE���g���I�k)�9��U�!����|W�%I���{Z��S�'�q(قg��gg<TIsT)U��{�_#�փ ���瑩I{;�`��s�����W��4�l�HG��rr�)�1AsE`�;������ꉹ� �m�r'�"��"�7j2���'�5��"`��m�8�ll��4��V�0��]���v���xf������lt��,W8-~y�w�������o����"���:hh�"!��c��o�ni_� ���#�r�wb*��j����;�7��)x'n���_��)�)�ä�J�aN���)��%
�誢@���W�SY���g�{w8(�'`�߄�iݾ|�
�t������lZ0����vq@I�?C�7�p���(���5�0=�L�e=���Z��>��y�דn�����:�w�&�fp���
��~������=��Cx�o�����Df*Ѽh�z��G2����|�L�<��6'����5
��JR���G��"*kꑰ$5M}U �	�O�:�����}tb<�V�7��D�@.�lj�c\b2�rm{�0�ϣ��/���]du��*���w�'S5.���	��B6g�x��٨
�1ܙ���A7*��3��ݓnh�A���M.�l�+�[ż�i���٘�8v➿m����a�XT��VS��0���Wn�Nc�]p���.х���i40��S�A�.ۇq��6S�7�q:�^�����M7��0���&0$E195[$�+���nm�W�b�q��@'	8��n~�6-31���q�E���x�f{���:� ��˽ݑݚ��]C�>��Q ��Gٗ�>���ǒ3G?�ԕ%�lSf�H�fl�JV�X+�_�����PA��"g"��Lg�K^����?�/d4�|G���ݍS���`�^O�DV��M3ݢ�*]�`�H?�������	�,�1Z�Wt�o�z���h�ylm�t�췽ӧF�w
��� ��Ut����/y�E�}Vg���{,��+��ò%Q�"ޚ���]��-�U]"�u�[���x�%����Ș}_��2���HL湾�pq��PJ���`N)�K���:�K�7��g�Ά���M�"�[g����,C�!Ն�y�\k���E��9��s0~�nգKDY�7!Y����`_D�S2��uB���H[5���[���qN�ğq��Y�@n�;;��X	2����pOt �X^0WJW0U���-d�N(p��ǿ��ӱu��,l�Y&��;Y��F^P������&Eͮ���??����8H�ёĚ!��������y���]�p��TS��T�LH��Ë�Ηu �8 f!�lM2V����ǋ����w7	1@Qr�T��xVاm�a���&<��Dv��ߢ�VEX� ������}���yIYl�ϝ�v��p�Gf��#�ru�g����� 0�Bh"����4�-�]�u�Ks�0��B����FK�vlf�K�5��:�>���q&���nsև
��/��x��l��[�K�g*��?U�15hv7���6Z�\ܓ���,	W_U���&��`��=�Z�;7G��˯�7	ن���l��b�	�Z�O �zD�(�*��_�>�[���t�j�-��-y���Xw����#��]I@-��"�Ջ^�uIbB�
���b��:��捡bh�e�,�*���*�)�ujXE"�v��?EF�:���ĝw?	Nܩ�	�Wob�t&�t�/��=BT��6���(Yu@{F6�����5�~�!�h��|�h� ��ue#�Ą0,*�[��׍{B�G�����\�P�U$阂���Q���U>��k��*цW�s׸�^�/�� /[����ʪl�~�\��t�
G[��ʐ�ag�|x�~�fa���j��[@��0��3A�5Hu%� e���)-YPQ`���Ͷj�j��@ڔ���(�%��y�GAG���<�)�~Y�[#��Q"(�52q���S5�[b"�
�0b�맙(&n,�4�n�uu��z�����fyf� L/�h�}���\�i���K>���A|]�������Ͼ`��A������s��^�����;�@�S�����v�WJ���N��R�W�S�*z�����I�Z������w�Rk�����B@�u�G����@�����f�T���^b�=-)��\���D��̻�<J@�`Y�̬���,���b:��a����Q'^���>�R��79��3�mX�~y���3-��0m��,��F��z�s��o��^����V�{��D4���ؓ# l�� �R��쉶�����[bl��m͑��ю��6���g<g�p��9�ǃ2f����{����ؾ5��{�}���� �`M��p�v֫R}S�1=?R��Z$��\KkOʹ��-V}</���Ģ� q7~V�.��HlY��r�ؠ_
��^��l82�oc��� ng���^��M��'���^�9?[Uن���,��o\�߼���̔$b����
q�f5�`hP���-��x�U��9c$�6V[�C��k��=!� �3C��|�tc*�o��WqwS�0�&�f!sUK���(�Ƶ��W���5�^x�lP"�s���	L����&8�.�`��	[���w4���^�XZ6~�؃����vY[��({�e�
�ng����e�Q��Oz;BB:�_��3T8Jm �d� o@����ĳ�"�~�z1/-���0��S��b���\J��cR`b�M$�]�n�(8�M��h9�n�Uݍ�c�`��:-jhI�S�P�Nz��^�b3,=aT]�'T��"�q�n
��"���܍�ߚQY���!Jj>�.��Kf���R36,��[��!8�����r�b��G���A_;����.�th��Q����r�^�xI�PLU��}ݼ��:tJk��%;��>YV��U�� 5����г���9��z��>�F?
�������V����@��W��b?!]\QjV���
;�p������;�F��0x��v��O0���C�1��4s/�k�O�e� ��.���	9�����W�$P(p%5�}&��mC���� �ؠ9�l�8��/���cvx[t������S�Q��oL������.��dTe�9�zCR=Y��� ���E>��7HM�!��}�}�� 8wi�l?�8��	hE���k3�Q�p~Y��.������u$^��ܴp���TрΥr�l�����\;�c�'f8�b�V���]g⸬�YtO��:��D"k�J�����ܹ�3�"�jͷ�L��;^=qqؐ�*�?���V�*6�:q�k.�O*���^�(��h��(���:�\.�L
�;bb�#��	w�,��@�ҝ�ޥO�Y�3�8� 4�vD�AC`L�֣�D�CLb��N`��VG�� 5��e�-�E������`��ˀ�I[�����1�պ$h��G��٩��h`v}ҽqi|������~�V�h�0x��c��啄�񓫿�x��	l5�EQ���$�x����63��-� �.F|1��3��i�6�)���r1Ac�U�nI�Ȼ�Ӽ�jV�
[�.�#}|��E�tՁ�V�"����A����e���8��>Y�a���#���3��g�U#6��X�b����z-t��q��D��h]��3z��K������;��m���(-�xM���g"R�*X$�j����^/���l!�BC��ZG�O�*�S���I��Vm�Y3����
����~��c%q�w֙��1�"oTz���q��*=���'��V�'0�I��8]q�����9ўH>��݁�@S��a�b��E�]	�����_;ٍ��͉���7��Ըj�b�?˱qq`��ƾ�>��������J, �K���G��u!�We@x��#0�Gb2Pz�9�76߯�M����}h� hG�:���g�WG9cl��>n�e4��9^�P���ߗ�&M0�1�$t�q�}��k��Űn��¤��.e�G��1�ږ��M�QN���Y�7���k&j�+���7 �g�r#L<�o�֪���'�0L�Ȩ�iG����{���0#�;�E����E�6A�N����&>�O˥�g����k�-�ɷ{��~��˭�*�_P?���V�	K��'J'��2�mؖ���_���Km�>r��ë\� ��;��BQ`XI�������S���U=yqÑD�mX�k�{"N���r�i�͒�j�Lq� �y�$a�GZF7��p��q����r�| =��}k�<�ec@�%3�7�R��v�W��_�ם*U�����'�6Z��I�Uhҹ�����xo���p� �`T2}w�F�J|_�lI��<b�k�6�.�¢WBT���j��H����huYɔ�2r�+I�d+�9O����h�/�lW�9��p<M�c�T'�o=2�gs��ϳ�ʓ�B�І�W��nu���B�8(�c�d.b����O�����V�����#��Q���3'ݭ���t�����D#!��@Ó<@�d2�ЪD�,3a=����b^�F�c��xU��ߌ�y5h��|�V��#��vpwR����Wou��� �9%���u���-��rw��F�-�ʓ`hW �@L����_���;�ŃѠ�ϦDY��;&u�ED���k���-4�jҧ�`s�L�|S���4~�8�.h����Uz��;�K�|�)7�`q�{�U���Ƿ&`.+\���솏4����{� W��/.��/�֙ciX���)H0�v�?��y1�g,/�x�>D��Pc�zI����TM	�Nm�tP9J?{����_�w��IY
[+��m��7�ﮀW�C���uc쒨��id <�Ի+rԚ`3���H^�� ��aX��rǵ��5��k�ՑE���3�wx^blx)�}�hbw��թ8��mF���KYi��rS�e�s�e�7} v�J|Ұ� ٚC룔��,��up�d���?����,���aS��Ǯ<�t�P|�$キH[�Ի9�'����*j�C6�v��|��0�P���r��S;�q ��S�t���w)+�"���V(m�0BFV�1vgQ��RC$V<���w�4�)�W�-��h�״�wa����Tz�j"���դl4��͎�k<���~ c�=�
ɤFZNp��b��s&��ik��m��;��O 5xj�G3b#YՆ��/��|%ޫ�ʜ'�d��p7�����I���Q��h�]�U��pP%/#*�P�?_�7��X	���#\[�Y!`�YW��5U )���ft�}S!h��1eغ��#O� f��m���G1�V-+�iv@C#7o�n��e�m( �n�}b`bN��+#�0�i���a9�랡z]|V�k�Z�5�R�H��6�o�A=#�A��$��Ԍj���z"r��
ĵf�E{�Ɉ�eT�I�j�}Yg�eB��_#>�#o���g�
�Wq���曑3*^��&�b�w��A��}2�����2>L��i���>�v��颐�)�H�7c2j��(�8^@7j���cJ��L�@��,/e`ϭQE�M"ز
G�b5�����g�}u#� ����[C�/�;v�Z�NW�cۑ�#b'̍H'���v��WE�*�^4��VS�Ȼ۬��($d0�Y Q90^�4�HQ�4-�=�4�!h��1����3���G�g�g�! `<Lz����G�0�/�?�� ��Ǹ�6�e#�k��x��]Ҟ�_�K��t�b�EjY}��/[v��i�h �	�Γ�*b�Ğ#��aw��,�ɪ,�xf�o~\ k����o!*�E�:����[;i��E��*�б �6>qC�i�F��w��|��e��:U���Yf)Y�4����WdV�f}����z���x���u�8Q
�4Tr;�lc�F��^���j��X�!�<�F��k�|��(b�@4�pHٌW�g�g���&�nU��,j��m��*z3��:eYW8T8T��6Z_xqh�{�Xα
a|b8�fN7K�j�]p��q�yP��tp�����4,�3z�t.����O�Σ#�E�}�/a�ڭFҳ:a�������z_z��G t�]Fw�q���W��cE�i�U �t�ł��e|[���;��%�����n����5gJF����I���ؐ�R��+�b��l���J�κ1��Wν/w����x�6v���2��w\g�R�@�P�?��ʛ}�6pL��e�2��/&�B��]k,���k���)�J磑s������n?Y���f�P�|uN��kt`�7j�l��h���9Kg�m�m#T��Z�U�ظ��"�rx֥�+����!���2�e���g.P�Rz u O���g�lN�nE1��KW����,���᰿A����9��G���kqјv����Ҟ��,��n��QK������
�%��iϭG�>��ͽ���0�D|�C�O��*�3sc6nId!9�E#g]i��c��\G��9s���*��5�db5۹A�r$��%1q��$zǊBu�����%�(wj�����Q����q�}dTl*�?Q;�&`���&a�`$�����`u+վ�'6>�1G�l=�ZZ�7�OL z��3]2l��4P�M'�����B�Ўzg�<;�����L���q���aږ���K}aϚ��W7B�U�p��]4�~�*r!:�s�Y����5T�4�vYm��Z��(���S
�Al��T�T)��vW�$21���ʧ�K~���E�)�\�����r�o7E��5�#�	��kۉ��%'p�l�ۓ
���gJ�5���('�+���a{��vC�cQ�Wt�bխ���7��J�0���P�BٷJr�HI�kooX¥Y���#��GN��j��f�����(�g_�I��;����3Tߘ����`ꁿ�;+�S�>��q�� ���P~�#6��S	�Ύ�&��<�{���]X]�XΡw ���P���8�?��_�nh��%�i@
��qB��?� ��!��4��6]W���Ȅn����e~��z6RN\Z�:��*�DwO(�&�z�����d{�q�b��o��*T�D��]L��.���Z���&�����ʀ��o���^[U��]y3I�ԭ�k8�6}_m����lT�\W���kt�<��.[/fB�|.�C?�="��ס��6��[_`l�E���a[�z�)�n��ƃ��W**p,������=<�c��l�Z��M�b���Q%YA�b��(Tz������OJ��E����م#�1u �8�1�\�xz�oG���� �*�AG�)t�}Qk��P���!7�cˮ�=M �a2B��=Y�|�Å�yL��A��_����ő��7j�3r��V��Q�J٤�c�z�l馘*�̳�����RU
��&/wy}k	$-�`=�X,Ȩ�uԞ
���T&>QuǕ�0z�M�RKl���W-����2U�ͧt�*k~�>~A>��F���n��&��y�дLz�,7
����V��*�Bh7I4���f��]%QN(u[���-$�P�w���EAk$�nD�g��d�1����X��-���8'�G��x�������aa����C��ٍ�|���HҦ�s����˩0����l�93���6��ðj���Ӧ���^.���� �t}���Ll�~��Iᩏ������0��c�`����1�bTO�� b�����l�	6bx-&4�E���Rh�����QQ��#���F�d�4yV��R�1�3G��=�t]%)w8��U�(�N쿴���ɀ뀃�=����ϭ�=+�W֡얢lHYO����=������+��3&�3�G��F����_�Dn���z�,y`j@`�����_������^�+B�؅����^`-�e��B@d}�"��5}�9��}`��?��G��&���Y:���o��@?ijl�b����9Ńork�t�(�G�?�19�zT��УT.��ȑ��(A
`��MV%��mx	�\L7�P�}g�? A�����w]}�Y�hҞ����)Ea�ec,�_V��鐉DL�5y{�~BO ��GZ4e��Ў>`%������X���Nabs��B0"R��?F���d3?Pc�� �A�0���$��uM�C�$j��m��3κ�R��ܧPFy?�߰?r;��]K�_S|.֓��~�9��"j״B��cǔ~1?Q^bY,��.�dkg��)A�����8����"y�ۘ��Z�s�	�"��*u��:���9�>7��.V�}_7��3�̿L���#xr;��,3!xJS��'��
��v�36�+ޠ�f���Ek�x�4N������r�6= ݩ��R��9I���ڒ?�%���xm�g<}GD��Y)��wU�M�Dg^ڵ�T�=��L��J�f/��c�j �:���/��'���2i=ä5�GqkL>�%�/�e��rw�u[�;ڞi}��������v.�	��p(=j�[�Wku��dϟ{�x]/U �"���Q!N#'n_Kf�j{E����S��N"��qP����o'Y��D��q-�YR�v	Z	��!|P�,A3�P��	�}��pK�2���U��D���2��P\�i���cl4T7�{*����ƺ�55.EFK���k�s�eK���F$,������50�	Z��Q���Zn����t�}�'����I�tb��&�K`�n_�ME
S�Z��"��L��5�L	[55�u�sA��|b����d�`��9W�<��?�=(�ۻ�[S/�;i���X��pk�.H�ɖ�¥��}�t�S�ۧ���<��n�\n������n��7w��:Q�?��3(H��F
�T����e�x��Z�I#l���	C��� f���k��>]S��_�I�.�U���`�k�������/��}!po���M�,�����%����NV�m�br������S/�]���Q�H~�x�g��RU��H�X�~��s�x�ܻ^���!u��6t(�q7�m�����cmP�t �Y)���`��wpAp�5�-�ȥUyu��5l��Q�	%~�h�)ʴ{P��?"2�B�Xn��Z���h��Ǆ�j%�XӃӧ	<�i���%���֥l�LIX�`�*��mt�Pn�l=��kZ:X���Y^���J�x6CIM�T��1�t�1 o8�Nl4�X$q�P���؏2U��=��4�9��k
�5T0�V��**�vQ�^��
x��VLq�\��K��g�z.8��=
�j|�p	�6d�����}�,x��j�.;�T�.�F1p�Ǧ�F�d_?rMui���e���}��|/2Kf�Q�kZ���~�WjxO��J"�13w��H�TYi��]'EKf��]pjfu���+)�
�����f����nZ=0�1t���i~�#��0������h�y~8h'�#�#�Li
U!��?���O�4f���J����g�ιCy��k+��}�3w�����+�γZb�iy;������r��g_O��(
��-��G%ٲ�}]3xx�{b't�§�����{rW��d���B݅m�������~<Ԯ5��U���~�
X�N��cIk���X��I*9�\D6�?1/T�k�j8�ASM`�@�K-&�qۈ���+<�q,0��ހ��=+�c�04�Q)T�B�u�n�1�<�s�c�X��'�'ae0T���dj!��� l)(z�7|�XCFU��9TWW;T�x�q/}�	$�6�-���ags�O࿧:KCc�Ws▼�2���8����Lmr��D��ZD�1�+��s�oO�e�|v��OW��Ty���3.C\��pǣD������2�<�[M�����c�&�:N�߶���˳���������@�L�KHН�%�J�c,�P�\�Cv�'iRwf�
�lWv%oF��_�ƑU,�md��������oM_l�[�kKS\�U����������h��u�;KX,&vh�]E�P%�y�K1re��B��҇�V�����Lk����)��c��u$-1�yt�]R��%Ж���H��F�C}���qI[9C����H����6�R������
H�Sx���<Y�ӻF��9�85cdY4���;�6{���͉5ѯ�줅O��J�$w��@�3����L�ak�K�e*��۹�ƃ�ҕ��b�"�)���*����5�>u�5�Uу홟P1�4��sȘ ���t��I�{B��E�K�	j�|AyRs�^�����;Jp	D\ICk��ַֽ�#6QL���h�r`n�vV����V�]E�LR'7��s��/���/N��`�s�?�� ��G������Z5x�V�U�k��g# ��OaA�ﰅ\�9��0�,>�$ӻ�d�p��v��3��=�^|QK��`$��Xӌ�;D׌Vt���:�D-���㈕k*����u�D�\������&��Z�x4>����)��{���O��1����>r���ݻ����,�����s�l#�e��$�/�~#��ܓ��}��V��$�j�s�@6a�^U��)S��M�M��͝N���2�fsir#�3�z��lc:p�\'���o�����O��	�q��L*��3��r���Qg�Z���."��9qjO�4x��Ey�O�6˫,�0Unū�!�I::�N%N�4���l�˨�q%��J�d��?��3��Ij�%��UaSc�I�8�gb�$T1H6S4Vn<���Y���/E����ڕ���c�_�(!��!��8��}���֜�N}�H5U0(V�)��y�f�6l���
w~p6��=K� ���M��M~�E2��`������]�Y$.\�x�Ќ��<v�Up��Q��`�����?��ﵴ�-�G��ؘZ����i� ����Cl�_���v讖�U��L��i�|4�Gq�	�u��t�/���M,�(
�bCUIgx�D��+��w��������L���� �H�ePjr��y�k�l�05|�������o@��E��7�F��9,�WN#��n�{�������G^�4�h�k���b53ő�}��� a���(A�I��c֎�*�*�<�)v�[&�X�m���Ie�ǩ�e��0F}d<��J�C�;��*���hP[Kk�[E�/��� ne��aD/�6
�c�k�*=��E�_����隈^���nh�T�pu�����F�u#y�C7a�T����v�diI?9�*�+�_�fD�.� ��{d*�xDm���w�.s��Y�
���|�ٯ䱡'��zu��)��[�O���5��W@͓y�9'��`���d3�Q7���l!��>���d��T��Rl�1^�3ߨ�����;�D�˵�he]|f+ iV~݉��y�D��MEUET���4ezF9�F++�&�ڙs_��-���5T?¦2�n$<�Q7����3�� .��-�9��"�@h����O���[���2M����ǌ���mS!�qG{�!2n�~d@
2  ~�7f��T*O9��T3�J{L�y_�
q'���·��S|���C�D�z��������	J>!F�����u��ދQ��`>��ɳ�Uy��Ŏo8gA
����R���<H��`3����*�T�4Ә���I��������u�H%t�9>h�k�FJ�2��oK����kW�Wf�/��T�f��Fn�iV���<
���p����$i�+�R a��'La��$�C	��J��N�l�&�	��*&MG΅�O��k��	���{��ώ���,h�k�B<�8������\3�D���u9Fѫ��D�lRR���5h�ª>M����P{��]��Pm��Ofդ�e�cd6:ڝ~$�<�ƒ�h���@�4�d�xH��W���`�;��B�e���	OUj"]�m��vKk:Wz[�F�g���hY��k�(I��]�f�&�4�b�C6���mM�:9�dx�9o��>��� e�0]f�(��X9���L+��
���y�"HNdVɱGpWw�E���h�R����"Q`�P���5Q���R��x�1�x�Ћl5�q�8�؏>K/�.|8j;7&��iM㓁
]��IzSO��p�W�>����\�B��8ɂ��P~_m����g3�U�/�%n��rM6���{�Bצ�9���5�5��=7��T�*��)��Y��`?ˋO�� |��9��_D�Jɱ�e��/G�.p�����S�8�Ì����=�����a�x�œ��X��OA���qյ;���;P�*�]7bV��p�)'�����q����C��d���RZ%��n?9��{v�����Y�3�(���R=�_���}����A��'��������f�F5>%4��A�4)�T����Y�� �ۯ5(K]'��)X#��yF��M�Ȯ�iX �a����t��k�M �� J!B8��N�����q�vʮn���/�N���9�y�`�ջⷈ~RC��� 肛e�TB?s+��s��)I��鵟��D��r!�
j��H+*���p�{���^9*w�v�X����n�QH��E"�E�)R(�QH��E"�E�)R(�QH��E"�E=��JJ�K
KJyr�⚱M\��Q����)��C)���������
J
JJi�4�yM@��RTSR(~SH)(�R8R:R<R>Q9N�~ЕXI��ّ��^�)6����p.���3n���[푴�
�H��鹦N#<s1)S��8�xAAu{E��ѣO))���v����m�
�˸���Z�FI�f�n�_�$�Jե�we0E��"��Yg���9�Rj�o
g[��r5�3�+M��r�����^�ܯ;lR�y���=�xH�̽���t�������N&K���o����D���a����h�D$����֬��!tHl�E���ĪQ�z�(�g�z�K|D�)o�����yfahӒORl�!�)Sf1��,1�b�)|
�_���a͠���Yd����8����M3)	����<�nJzq�cZB"�<2��bD���� ����s�%D^�F�P_+�LRd�('���|'���͠2�A\�v����}y.���EP��q7ia;��C��,F�֝�ŀ(n|?t�ۢ/#��Si�!����nl���(H%�1���0��hԱ]7j}��]y�������b��%�%'���@.�� ���]9J�Y��K����suA��
䅇��j������u&�#�="&j4M�;Dk�	wI^5�]��+2z�Fa��,#�&H˵=?.�%sΠ=M�?�mA��X�<���u�D���1K�ii"�W0���_�s��p����c�t��c*h��91��s0ֱA�y�X�2����+c]!�8��$;G���zki6�/�õ3or�Ѩr饕��A�6��XP�	eMPa��i�����[SR�H��]�S�p52�e��fT��㇒��ט���V`{R�M�ԔN�_��!G
��Em��'5h�����H�t�@	W���*w����j�`^�4TX-��C�K����;�0����'�8����	��RR0��0���"��_st��re��J.^(��x��i���E��,tX�c��4h~���tK^-�Ȃ���Y��g�����	��*�6�4��y�v�׆�h�E��Q>�EF��A"�F�Ig@6��*p�Z��+l%hB�J=(�E
�P��w�ROdt��^��na	��浨F�?�B0���A�<*j�F��괻���A�c�/�]����v��8V���t�-�g�k�we�b���W��C>߹�H t3��tP��ۛ�3#��_��im�V67�]s�P�H��<��:7�Ā.�.I&���|�:'U�yxm�b��a����-���3X屒ǲ�e�HI�D�I_6Q@%�b,�犬�Q
������ߌ���z�S	w��>k����b���� ������F�A�8����������4�H��Dǌ"�V�����a��<��Z��H�I?�ż�╨���B�մ��J��I�Qc��A�u����!�I4��7���j��~��̣�K����,&`&ڠUG>UQN�T	�,/�U������,������N��
b6�%�T0�Knz��lc���QE+�C�e��R�Ͷ���+:so�_I��Ec�����3�?NX�N�"��xC�fh��	V�i��{^{_VI��:� ��/kv*?N�QV�)kҪ�~�eh5\�OF�@&����w���-PD3F�e��������h�uE�^�d=��L�dꋘS<'~���x ����(ͭ}p��PX4�\c=���c�Y@�T�-��7ߓ֚+�Nq�x}�~���F��.�'6.�:1U�Y?�Zm�vz
B����Ћ����1ר�N6/(O�?�p����>qO�5�q)@�W��q1��������d(4L����\*�YOB� Dn~���!�pc���|L˃ИD��R)p}�sJ~L��抋w�%��d).�X�������BfĘ=������#]�x{���#��̏Y�U�࿷ �C ΰ�����Q?6)T�Ak9ϧ����߫� ���+�u�M$�B���c�N� �A�)t15�s�H���1Z����K���A7��C<��� �a�1ޖW�
</�i<e�2޸��EFl�jQ,t�ϑ�A���n�W��n�Y���*5I�1�A��b���)[:�y�>$5��=��_jNx3�W�e�[<�m��B΃�6��)�����b�t�C�ƈ�[�Ƥ]��;�'�U��d�A}����?F�=������bnp�^z��Ph�oɓSX��-Ŭ�#��Q��d�=�W�3��E����҆�$6�ʓ'�k�f&7X�Ʒ�:�=��Z�t��g��4�4��cL��`b���h���'��u�/����M��B2�H�%����ό|���!��V�^�
.��}�<CP��j����x��;=�ihL�YR<S83�#b���3A�cD�l(Ҹծ�XK�@�Z��Տ?%L�E	�;p��0/��9N�Cb�� E��Nʷ����Qf��g����g��x�hQ�����S��23�1	g�9�����<�;�ôXT؅��7�9�jpZB���Y勵`��g�!Oܓ���灞�A&��p�e�>��������{ڮ�0���޹�6�.�:}�(vXB,����$��q&�y���:���`�ǔ��3�y����Oy�9�͒�Q�]�~���{MÛ���������� C�:�D��倴n����f;��.&+6fmչ3+��1��3��|�G:����{���Ϝ��=�Ʉ�end�G�#��Zs9��k�vcv}|z�}{��_}���n�h�|?'#�U5Qk�*N$�V����!I�/Ө�e�of=w����]yW��W<��r�{\U	��[9G��ːF8�r�޽Ru��S��q�7����c����׮��{����9o�� v��h��ޑ�1��E��� <i�_b]�a��h�X�b; �~k�Rt����u�V�j��	��=�) 1�cj6Ӆ�Z��Yܠ {§���3�/Y/y���%��&�M����[��]� ?8��ė\�Ԉ�hW'�d���i�D/����Zb�A�X�;k{�ĆA`ŻR����
ʱ<<��:�5n���OR��@�,c����v�6�b�����M;A;B�l->�#7��qqZ+�؋L�-F�\�wB\��E�K����F��S����?�"`+�""u	�h�v�A��62;��[��q�<�3)�'�{̅�(�S�ݹْi��ib�|ʓ�^q�R~�U��a�Ĉ�5R����a1Z�b��y�x��p�t��5.��QhB�&��OԱ�N�'����@�2:� �U �Z�_z+���"7#α�u�]s�Oظ��UU��$~mԽ�c�K^&C>M�� ��b�~���� ���B
�n%�1515ZF�ٯ6�������$ㄫq�ܱ� [��mQ�|�kN�fHn�Gua6�^Ӷģ�b�\fs�)���U쭖!�
�^�ao�����ϻ�ɛp\���=z�&��:�R"�kEn�X�q�/~v�	Q����k!9�-��M��V/|9�#3<)�r���8���7�\�����_<�����B�M�q�x^�� ӻ$7=YEk_Q��s�ub��}��g"����O�Y�͞�W�=��D��XL�#��.Vh�*�@�Θ��nA��B��q1��m����6+���%��/�/�3��ּm���N��&���=\�qD��?M<��<[�!����^`���C���H�))�؉���ԇ������l�}�ֹ���\�;��YZ�~[~�����-}��Wֵ��d��Ql�l^ў���v2���M�{�A�.PĆk��V�Z���7v�]�w[+��>2�{�lj$��Bw޺:�d$�yu+:�,���v���w���qql��N��YBB�w�&��;�E���d;�2��Bqc8��^�A���[�R������ҊR��I�h��"��J�_�v���ĸ�.â��Z�Ep�P����\hfQ�AֲǔR�����/���X�/+�jr�J�;%��O��C���i�`3(a�H�)��?a��bL���m���\�<��od�����F+uX�R�;�0����R˶����c�26��ֹ��iG�탿�;x�`{���Gr9O2��\���c0)dr�4.�&ӫ������˝SD
�Bg[�Q��7�[�b�z&�O�w��+�t�����F:�FC:���JWZu�\A�|��CYo*��!W�$�ϲ�h��T�{�18?�s:� τ��߲��3��5�@j&Dѷ2K��`Ǔ��ZW3��X��ևB�1��4�un}f��ؑӕ����F�Ğ�K�[z~r���R�<@VJ�v�-��5�Z �e���R/�)�O�E��I���P	9e�p܅s*[	�W�x��-��V�,�����'��"P�R���T����$=!}/�*O�YY�	s�J�����GU�f�)y�(��΢�k�g�nW�T�%�=L6 �o�s�\xj���E�b��7�4�T��xT�����"��"~��{��퀹aZ,��FpX�E.�:��;2ʌ�mt�/~W�A��G�@<��O�!ˠ�� ����C\���T!�"	�g$�o?������V02xE�����ѣ����EԱ�#a,;�ɪ�	~u�Q!Q~f�����<�]<>/RSR��^�FV)��K3M�V�emM���D�z��>�ћ�]4�b.���@~y�3A>{m��x����0��K0���2;��8���P��C��l9R�.lۈ��o���0��	Tq�e���e�u��P�(b�A��߰�"sUT~�C�G��`�\�⼔K��Q���z"עT|	�iZ+��@� S��u\wz?��c;���.%Tԡt��;�@Z!s�^����i���_y?����V]��9�m�^b>B˧?�:Y֏b?���y�A�w+G,�u������ړ���Y�>)���SU�T��S����P*v�"�,J�j�H��}J��Ƙw&�,)�R|��!x%������W��7�d��)��Vs�m�t\J��Jr���0�ׇ%�.��-�#����1��4�BQ�"��d.��~$���u�U.��D%ѿ5yu�:�k$m�1r>���s�G�%�4��&r���-��q�K�"�/�:����+It��fi�*e:�]DZ'�	��M���W|H�Ax�ܳ7�9�*��)�-]H|1��I*�1<Z�v:ױ�1�])�!�F.���.�'I����(
�	��$�;�)(9�i1�����!Q6D 6"����31�Xp"ӣq�7֩;x�:&�$��F;�v��F������ RNh�M9ʀ��9T_+p�4�4�
�%��Z���澍�Rs��U�B>z�5���|�V��w�k��K�1*c��9oq�İ%.5� �I�O:�2od(�鰣����#� 3˯v��̺w���Fg��ܺ��sT��I
��~iԟ6j;Hz4�L!F��[������rI�p�USj�v�v�.��i��J���b�8���^���%N7mOA�����bD�b����ť�l�`2�k�;ګ
�-i���O�=/T�5�ͩ�9y� ��F�ࡡ8`��XtHQ�=	�w�\�4+�p"�D0��hy�A<PP f��{��q���Q��Q�R�	}0�5;΄�g���58D�r�q��UݬƮ~Ta�]6VV���1���킉�oS<�V)�)4����ڦ�zF�����cb��y��2�.�%U�P�,��E�;!��s%;ո�T���P;�-v^��o4Oa���ݔ�8��l��ciT"s�|�2�ԯ�*�#�Ԩ	M��/uM�V�U�lj����Iϙ7&�>�a��6��%��_�-m�no��`{��;�.�(I ��$��<,4j�,Z!�Qт`��q�̊�ט��W�F�r�%c���c+��fh���|�r�pKf�i{K��!�����<��a��L��@f��^��t��m�W����ֻ�sx5�@�kg8�
n�B?A�$��R@�3D���K�σ�j���:g�D��I@� LM���BJ �s���:'M�eA�<:h�
t���ў�A?$���⧀��C�o|>�}8�",���X)�\A^k�;C��
���sÿ��>���1"����d�z�W��,z�#!�(�̠�5T��B �>�崙5p�Q�p>
�����a��V��ر-li�Κ��f�����#:���}��0��h@��0��U�b��R��r�"�c�"���� �"ʟ���	G��&wfB����Os�f�9�ZpΆ�*��x4�5+0-��'� �E�t`���^@JA���%*Y x�*��e:ŝG��_-�+����#�hދ�3=���q���;y;2;c����b�z7G������w�`�Z�+G_L'ue �����>w��wZ7�HZ��R!���k�Y��'?��]�f��	n4�1��no���!Ѱ��Ґ[R�m��t�ñV�rag��� }�q�����O�%��{��L /6G�����n� L
=�#i�i8A��Q�%���ܗ)���$8����*/��V��tݔ6Չ���F����i~08�|[^fy~I_�#��Yh���VvQK|p���[�a>y}�2�e�mg�F�A��ֈY (�+4?G���0<4��ѧ^`�EXZ�	K�C+��r�m̉���枎O��� _�m��hC�bbU��M�cdS �z��d}�[�*���U�����Y���j�����ಔ"���0(�)΢�XY�h��B���	
F�ꯨq������$ؒ��͵�b�d�M����N�� ��GbA
��T��;1E�� ��ƴ����a9�I�l�#�dh�9�y�������6u� ��`�L��ӡ�J��߳�_�M2��*@��9 %����񧀸�!R A��;���n����R��`|�	$g��vpVoް��b�cE��AAy�y����5�^�����J��o�ص��WO�%���ȧ���t�]ϳq,g�k�W����HA.~5nE������G��I�%t0s'�bBJ��1�L�=l�v_����׽�J6.��r��s�⺑odg��s+9t8�l�!D�%?\��P�h�CU�n� �����c"g����m�׳���|K��*C�A�EhS�O�b%�����a=k�������LV�2�Blo"�0L��HB�oQ�4���B$T�^�{~
*7�b
>��4�Q������ �I�K����C����ȀH�5�ÒW����t�C��`��r���s�A�D|_G���W������i`�d*r&����=�ߨFU�?�y>�� 5Fm�t�uͺ ��_<G��9=�*x���pՌ�B��0޾�[ 
����� �HAr�����
9�}rND<�E요]�U�bR�X3���w����@v����ǅd������:T���������Ar�`A�G_����AN��};�pm��$��4���܀���C����!H���$#g�d��3�4�:gኲ-b,"�]�Q�0+W6jĊJ���X�z+1�A�&�X�ՒDM�_��#GO�"�~Y��X�Q�ع�G\��u��9aښ�w��P�C3$��u�&���0��/(�'�Ի.%\����=<`{���z�}�I��,ۭԥ{n7Z���s��0�!�!W�0�L�L+Ad΄��i��w����ԅ#��3��-���W����Ƞ��b�F�l��GQ�a�W��r�]W�`��$;i�������	�+B��2�]]��%���R����IȨ�!K(4�n��
�?�W,~"c�!�,΅,~41&S���ߗ�=/���;09|R�y׳<�R��\K 1��k����������8
0�	QC��I9��B֋2b,[j��!�5@�q���(T�4��
����*��Q�1h1�'��2��-��+m����dR͆�KX;�+��*�{35ۭ���F�C�gh,6!�>�yj"�%f�eOc����b�aP�׊�����Q��P��{;zP�l�k�h�x�5v6Ƞ�.�ڎ�R��%E�n��]4l!t��*27u���[c��I  z��VτO��$ I5m˿ t7�4ɗ)+�/uū0�{\�H���Y�(�	Y�!�����f
�i�jP`z��<��9T�n�_�H�_�'$�
x�~�qz
���1��q��ǘ��pݴ`�*����{G;J'���"��:(I`/�=�,�ɱ�&����$�j�Sp�R�DMT��
�lAM(����M��u9��U�N���|$��/��/(�|ͨy�*�^l��s�#�[-�Oh,����x+�&<
9N���
���w��F�Xj�f��\j�e#��S%��,TH��$�A�2(*��I:J�IP>��ϲԾB��}���iMs(���_P\/�V��1��6�kޠ±��bCh	�7K�Ü��i$N����A���<���Hx�a��O���A�O=.���� C�"�"�\��u��k�]D�7�3х��Cf	�{&��ВOȘ�Z4B�^�&�h$/?�	ƛ�ޅ664��E���#�����X�C�k�����KX���9��7��/�����S�x=���7*2���U�ዝ#b�hZ�!N�{K"��πT|�6���N�c1��@S���s�����!����+��"�L��e��^7�/�;�:��6>} |:t;�Gf��>N��!��8S1�̻7]awp��c�L����-�$�Zf�s��i]yޫqh3˨RE���)��/�7�!T��4�����'��4޸�������mt��U(4tAf��gv������[�]LQ���M@���36�
� ��v�l��Jt�D�j5��w8��J��x$) J����b��Еh?˶������Xw;OE�X�]fN`�ぼ]V��iX9�x]��g{�-�Jj���-��l:����t�`�]W	�^�[x3���]$/i@E&��0��,83A�jy�Ӆ�tj��CQd��4|�,�M����U<�o��[?���i�i�bV� �3�0���A66���Gyܫ�"du�?%��!s~+�5���+9�I���~�ߎP���U8��e��Lg�Y,�v��r*ǃ�eD8Q��R5%U�*�%IP砹b���
P՚�t�A�������d��ēnTJ*���a�wG���׽'�TR�X��iJ��j��㼳7�Hx�k�Y�wȑ7��U볔g�΄��Ո�D&1]�_k	ZSC5��S��*Hid�d$�o"�K��l~r%dB�BUK�F��� �ĺ��JR�Mc.�/��3��As�U����;�:��0�EU3y�[�Xϛ�#��\���h�|�
����Ve;�nA�H=V�ۋ���+_j��!^2�3�St�7wHT����*р��dr_��u�����B:�;9�҆��j?VR��5�`q��K�q'���B�k��+I�ƺnVs9w���L�9��W+=���!J�tsu�wⅨ��p:B�� ����T�j��2CM�����úf���@� w� �:�szi����˿�N��%\Tջ����0��F����A����}��g�����Z_�=WeL�Y���+���e ���@���Q���ߝ#�:x蠘�����#\���4txB�*��&Toְ*q���=RpoPW���F��cz�} m�3�z�9Y�xC��ڡ�A���t�Pޠ�X1堈�ޠ�א����	~�����P��%�oP	��I�.W7Nu�.����0�҃
ک�~�!��U7�6S4����1�2qJ�&#����K��P5Frk_�W1X#�����v}\ֽ�Å{�i_XQ�ғ�8:$8��z��>H*Ӭ�g�,��i]s6�O!��$JD�ڜ:U��U�5v�i�m8��&��.h��@j�/��4qh�5[�3'��٬�7Y�D��I�<��d�=�a���c�X7t��� ����0F�MTy�;�@'�i�i��RՃ����M�U:�0Wu2�e�=pӔNpp,NU	j�IXTb����$�5���E���*��Cx=)X>��.}��8��d�$��k�D��b��`�����f�8e	��R��9���lƊ���F��Nz��?jN�t	������Q^��#B0��?Y�0�I�����F�A㙪)�weY������N�"=i5��T�H�C�j�܈{�X��Q�I�I���)X'�=�un�<�c�5���~��#JQ�p7S���.&�V�9s�N� tøl�� t���e�Z�1�I1�N]�q%4���] �w����{蓁�6�!���D�@�����{,���y�n������5FL��/���uo$���I�eep0r~_W���c ��rNg.�*�A����+�6X��y����i��Z����'Z*r�5L.3YA&� x��_	��ex�z8_��"VP�jh!�0���b���ҍ�u\�zh"�}��&
�D%0�c�&���%�2�ŵ(Qxȳy���唼q�O&��&=iP6U|,����i��U^bp���n5-� }Tg���r��MK:����0�
���Q :k���Cz��!Ng�7:`.L�/�|����P�3���M��=�q�6|Ƥ�R��� �i*ay{���T�O2}�z!h<���|]mP�]k��A�A(�ƴmް^�Ϭ��G �o/�Wu<�N>���i�x�~:�j
��]��sc�������B)�S�➩XfB���n�ҤHtw��%}x<��a�i1��t}��đk��"�_�˔G�@;��A�� L7)���ɽh�Z��D�E^`7�I�X�)1���Ϫ5�I5�s����|�o�8M(�г
4K����sMj<{�qQ�`��{���2��F
����X����Y���3��Vq�E�|�p�#���X+�,�(� �������޳��etČ�
|1Ȋ\������myxeT4~ba%��x�#ol7 �r	��Z^h��XfS���Cg�xhR�?���]ϛ�;I0�N�����i����#���o��J~㪫��͓��׏����P��g�T5M�S^e�o�1�2�x��?��܊�p����d��n�z��f���|i�QZK��<�+���F��B#�q�-���\�My�#�K��'T��B��鰑CW#���2H!�h�7>�(�kNQD�O�W�C
�d����P�T�!-Ԓ�"u4�fSD�F]�u'�2 D�r�>��j3I�~�e���?��-)!%DiG$ئ��h7�fJ����"9�R�99���?	[oSԯEn]�}�4�D�ZR���i�J�ML��blb�*v�sK0�����S#"��A��j}σ��9z��	G"��+=�`d˯:�O��Dެ��E��V�|���=��.�?y!z��eO��R�MQ��J��Y�	
ߌR���{��T�{�W�$Q{�1@�)���[%f�Ú�,D�"�n��,X���NZ��в�#�G�IA��q�mq�8�r+Y=��d�K�2��ş4��6|Wx^��侖��;��hS(@��7`fD�|˷�<�w4'��7�z��h5�w�.�*'ӌ���(�8��"C�K!��>i�r�
3U�\B�إ���T�H�]��PN�����ʋ��_᧒%b��G�f��*lɳ�:iFgu��r�ܽtg+U�,T�"�d5Q^����7��rܲK��h�S�1��~y����x�Ȳ1�28��hW�7惌����,��	��rJ�;��C{+S��GV�\X`�C�?LE̥P�/�Q�����bM����N�V��E8�cР8�ό~6k��	"����wY��N��2�(6 ߧ'2V��x�f�e��ܕ�į�2XD��M�虊eR�N�ݙ���Ъ�.ߩK0U��#��?���,�����!5K��vV�8�kx���N��+G㧌��YH��.XmI��(Ɠ��|N�{'|K�BMN��w݇$�!��v��2:��Sؖ��`���0-��(94�-�M�Ų���+M\��8BV��=�}���V�ihV� ��d)�hH���9M�*q���q�xW�-��(@���L\��?�Lz��M�}kIZ�eƒ�U���M3񷓹Z8�ޮ����K,"B&9�A����nmzAs��!%�V��~y���3_�k��$�6�RAD]?!gO�i��wHO�
�¡P�V�.��o,R>��Tb���w � �����R��|ԏp.�ٽ��lLc\�7
3�-���y�W�:�y˷�'n*;Zi5�-k?z���lN%�L����m��T=���`��raR8hO�Hm����w&s*����զ�ݩ\�<M���K���ݣ���ص�^�0d�7kj���N�Y\��"ؾ���2'��
h-��JO�Brȅ�k� �y2�A�<�$�n�n�Ba��~/�s��4еE�u�����K�����M�l�I&�zR�UF݃�FP៶je�5��_��� 6]�׍h�"W���	�+�2�]��W�+��c�G栶s^��O�go�����J��E�_�]�5h�2�9	��#N�ݎ��&l�i�KT6��I�wk�
QA��h�Ad��%"w�����P_�Ŗ���'�1��F�=�{cPl�.���ze�C�u����[>~0�&������;"��:es~W>��*���8��Ĭ�"uR?���3�m|�_����3�GH"�����`9�=��/؋�o��yd	%���M3�Ħm�O���%[}g�/�k�ڽW��=�dC�`����v`�|��������=����7ͻ�g����m�>�ԂyB�K���V	�\�_SAIO�W<�>i���̠4���<<�V]��6gB�8�;��ݢ��wm`}������16=�{1YS�Hn��ԞI-��0k��$��	~�za5�k�����Z3G�o�s��z��0kb�my��O��!a��x�[��>MW�$NM��|���S���qp!T1���w�sN<?��=��4%e��z�Eԉ@(�Ȕ��|t���ȓ,�8O��r�-�hy�?:��w�%�����$�J��F�R5�wx"�M�pL��<&�ٳ��s٘�BȪ(d����,���	.��x�{�gj����A�G�̯�x����M��9 3d`ӊ��h��8 ������}5ۍAG(��.)�,��{�n����\ U�%]�$�������|������_]b�� �}b*��Q����:���%'�S��A��|�_��O���"3�X��D�t�G~m�5�>���+�z;�U3��F�������=���ptG��d�@ї�5%Y�ҟT�wP{��0h�K�$ɶ���B�x�QZYV���v���B��l=�����cR�V�&8��K��ʟ���g�ձ6r���ˇ���s��|���9^,�n�/�]����ܹ��r�u����/L8��F1.*(������	�ڒD�V��6F��6f��6v�@�I�8G��>�J��?"�Z��}e�Zx�
I��9�t���ಙ��sg��s�F7��Z8�x�J7cM6L��9 ���gxI3��8�ex	vVՁ�%OhX��1v��R��"�(v�c�H�<y������(4�w�?�������y�(�3��c������{���ڠB�*Hj�q�OϚT��5ی̍D�6��o�����Z�M���"���3E����J�[�8S+��7��-��m�m�Z���O��3K�л����=)t�S����:Z+�`���y�)��`������T�W@i���L����tQOk���~�ʚG�gÉ⁰]\���!Oj�QZ=��V��*���е�hQ�7~�����6��'t˩!��iu�P��֊��@v���Vz�Fٔլ��@��3��W��������9�N/|"Ms�S�J��"Yq�ۗ�$rx�i=���Č&BSr�7�~�ӯ�[��W&�3_�����_�5�GsA-A���?&ۗ~�FMv� �>�^�[���}�:������8}�����	4o����5�ȹ
�~df��X'i���������L�,!��#6�0B����9��G����.2�F"9�Z���?z�<�]^|�d���%,K�}ג�bwQ�ّ̐�Y�O��g ��O����̌��z�Ko�q���	x��sd�ѧY�!/1���yW��uAV�8g�P�v!?��7�@ju�e6Շz7�YJ5�>�.8��ϓ�j��'�pyn13?��)8y%lQ)��E<�h�.��Í����6�R�unT;K]�7+Q��6,��F;����I���K(�[�H
9���惕�S�9x�s�7��6�S��x����;��rq�<����w���zz��T���`@�ϥm1�����<���^��ЫY�{���p�+���ʥ���4��)�>������~W7%":8�G�6e ���NM�6DkF���3Z��i�d�����<��Ϡ�����\�n>mv�@�Qx�g��L���1nN�ִ-�}ܙ�j�~j��+��]�W��y�rV�4�wWR�qL~qΩ8L��e�d�}����s�Ulh���t��k�\÷w�i�h2o��A�n��
#�K�A���7�p��]�RpOzG�۵�I	�(]uM���^���jn>Pn��A�;�^�2�)4l/�pO",0��@&��'K��D������EO�x�c-����!���D�=.HU2p���j2��(e���;si�_��M�Cq��{�l��,xml�j��j� liEQ��#&���,"f;6{M��:����0G�#��w����)>����?E�3'9ೡp�6��+o��%�>�p]�c��kїq�������4�GX�S� k��+\�=�d~�JuT,gI'�&^E��e{�u}�T�����k�UT_��4-�uP�Ė��~T�S�g��A<�8�T���)2��ݯ*�V��.��!b�)q9f&s,��n8�W9�;�!��S�+�)Mai0»yO���������[�����N�����K(gK�,��)]s����m�M�4�h�zX�����W�)�}�N�`����8ñ�|��I��?��Hp�ަMHf*�r�0��go�ӆ:�A/�3s �eIԬ�����oc�����i�W,!zD�$7�S>�_]�ȴ-t����@ ҬRn"�Z��"�RȔz%D�"ط��*��j�t%�I�D���R1���^ʆ_�w"�� F�s�e�7;��m��ND`���򘾻U�=���
��A��	��j�L��f&�����.�>�˩��c�-~_к_�>o���:��Le�] ���H�:wVҎ^�v��o8K�{�7)
}�� 7��5����ʎq|]\=&��w����r ����2�R�� e��J�Z�4D���J��ϲ/�y�J��8Lh|4`�%�ͱ�ӌ��)�Yt��跈�d�\)6��%o}֖LV�����%{�D��!������Xt�.�I�f�N�����zUA���^�������/S%�ӽS����F�ǲ��'���U������/�	�'G���N�QK{��w�gU}�!*�|��d�¸<yZ̹��)�R9vQ���X�oݎe3[��S8��nh���~�9Bz�a@�x��^sXB���hPy��;�O�y�h����h,��p��d����xr���-��m/L��/�)�5F[,��
�Lg��:����`jg�5hKځ����׽�/����5�<����^�m֮&�Sbj'�.��q�d�?]��O���Y�ô�ÍT_�/��S��2�},Vm�ͳ��V��ӆ�.��F�,����ֿ�9d%�?��n�u�[M��Ŷ-�}6�(a+ �bi4�H_٠*{�]�3���2�33s�
����W�(Qf>Ԍa�j�0���_Bz!����+�G+ ��}���P������CUyW�<�}��9�J�k�5���~� ���o7�٥R�����("єQ=��^�Q�/���펌['�H^o$���gi�6XF��֏�zYAv�(=�@_B�sjWH��!|��j�33.�
O�Z� ��&s���+o���05�6g*��h.g�q�s���e8����ge@Vf:À��9�M#����l㍹�=���~[�s�?����C��_)�2]����avnR6gfٰ�F�PU�Pd�v��]�;w�߹]����{۽2�z��l���Q�m��8�"z������G�)�����|�'�P�1r�G@��#g����O3$L:ոg�mV�����ɴ����|��>�������ҙQ���ژ{ /�w �P\w�	$�=`O�e+��0�B��V��ϰ�e�r5\�-fw���7+Δ�U�"�����Y.$*�o\K�d��6wj�-a����%�Q�i����ۊ5i�zz���~�i�ʚ1�u���CS����-wM��Ff=0�@�̓���k{�*��`�b����J{{-���~]_���|+�у��]�F6��i�4����@����k��`|_��7���;K"�@��F��͠#�O	��$	���L��'�*�� ��� �&u���ڄ���H���f�}�v'�l�+��o ��'��&>;o8��ϊl;6��WÎ킔�Ռ�4C�XP��s���A
��JP���O�	�6L��i���IJ�����C|�������c�`1Ǭ��<_��1�A���6�l07& ����*�D��tL�c]�8yo�^�g{�FM�rQ�5��[�W+�D����8�������섑���
n:;�$����U�b��	-B�T���W��OYANΟ0�D��$xa$�P�H�*�î���N]����\\�nK��B�a?_X���������o8S���ɼ 1�ɶ=��)�2�9�:����R�K+:�;��geI��r�(Y8�m��)1�9�+όVn"7�=�H�����D�y�8��YU2�����4ch!��;�$ch\ȝ��֝��u�W����zk�[���K\������"�g�M��̣A��}�D$v_�n��/���X^��9�	��
 ��|Ǯ4����Й�x�Ǟb��46/��	Q=�a��C.@/�v�B�y�z_:d�(�_��%km�������̩y��>��BZ: ����	'��2���x9v)���!&&�?A!�3/iHv
��U.�� �I�w\�%~�n��&�[������;��/b�o�koRX���	��j�6��C��tCU��c.�j���0�m�4`�#��,d$�-�2�����Mxi���Xm�9���G2�]��b�_޶�� T7�f�p\LI/��:��L���s����V�m�����p	�(7?#o�&zq��-����C�s'������^wb~�-� ������g���<�m)٤9��
Y!��7��}"��_��r\�/$h��_�r9|b���o�7�3cV�։+��Vx%hz���}���KY3Tk">�:��1)D{,'�`S����d|ژQ���8'Ta���3��f1Е�O>3�KIP�,�����j:��R���B���0�)����+�C�d7�����װ�]�"�a�R�����2�2��ˁ�Ps=�Q�����#�,�wGp��C-�H��Ӄ�I�T�:�6��;�/�~Y'�(�K���J���ӊ૤�#���Ǹ,��SY�*bwQS�Ke�ǝs�E��gG�<_�%����Q\!�=�(�X"-|9�Bц�ޅ�#��slC)wv׭ȋ�z���$0�B�!�-�����C{b<�sUy j��[7/mt��xߙ�0�<��GR��@�{� ���]�)� ^�{W�5f���a�4��P����^/��"�-O� OmK������ȣѢ�t�\�Je�5bVp��C��Ì�7��(j�V��v��=e[�m���`oզ������Xl�htKv.>ث#m�z�ߴG}j��p��]ʬ�*r�U���rL�5Gs5�s�!-EGKh�`v0!V�W����`ZP�F�Oy.�J�%d�"Xo���`m�
R��yU]a����H�����@ā�mҶ�N���L�k��k�`��u\.��5�%�nq	<��kwh��%��PJ�*f�Q[ᢉ1���e�{} �yc�-���2l,#�A��(BwX�t��	�dִ�����y)�
"��LJ�@Cd۾�����U]��у�"
�V���=�'F���C]q����Q��ZӓZ�����u�9�Q��%���_�z������97��RM]}k͌-Tr�^֛� ^�/,Y��Ylz�4c��t`��?<2��ݳY�!�rx*V���O������ݍ�YB]����Y?��ю��sb��'n69�hc,��p���kţHM�G1M�a���$��A-@B D��w�z���VZb�ȧ��L���d��;�@d܌]��9��u�~6]��(�ϱc��B�����E�o��f]���O����/�y/�='uDR|����|�*���_�$C�͹'�G*s�SB�\*�Zi��O���F�u� ���X@q������:�����Q��4 �NTT��=�M�<T�Z=�
��Td3�jC�4ȔcH�uG�0h�9��K�Ftw��:׊�Eb2���gşy�U�J�Na�tF[�$}UU)Q��H[���w~�/�_Dq��ꃼ�f!V��x��f���+�n�e�����y�P�-���@*�����w,�q�h����� w��74=�o��Mb��.dʍ�צ47�J@7A[₟.�{���}�kU�V�S�+з�~�l��6J#����'d���n��|[Ag�_C����$��o7^�l&�}u,۔�����D����X0�ŉ�߸�J.�k��	�e�T�ѯc�����l���Nlx��Fu�	&���^)��'�c��+?�UQ�y
�i03�V������4�\��O�9^i �m~�A�cpfvc=܉��#���D&z)4�����[��)�UέD�����g`�j��=_U��a6"3a&��M��Pbu-�B"���A�$`�UJ�
5v/���a5�Y��<�eM`cu�n�ђr ��:��7#��ݓ�&� [X����S��H�"2gi�F�bx�E��;J݋��x+�H�9 �	.��,p.z6�L|�e���t�h%;�8�w��+±
��-�;������1������r���ȟ���:_!g�w�4N�bw��ͥ����?���A�TG�a7���)fq`����� Ru$�.R"�[Q'1>)s��!Ѵ)c�9�p��c�
X�4q�=� <�)��@�M����Ѓ���������N�$�l�loޠa4�C��W�Q=H����lG�/l�9�T��j.N0Y�js�"�Hڵ٣��cH�}�WU��Q[�i�}�.�Y�6�O0�1y"��*]ܫ�[�v��a�B3Ը�P��ʖ>��o�`��K��A�{�+l�M�i��=o2�m�{�a��|³���aUB1J��n����jJ�&� V�x��C���1����9���g�*�S����W�مu�^�`:H���v)dn-��Ze����`�B��~�du֏�������*��m�^����֬Ǖ��v(d��h5m�������~�jR`nsC���.�_��n��Q�V�A�%9�ɤ*;����o�	J2��Lha����YK��A"
ˌ�俛�6��^Ki�
�W������"�e�4�ϩ�K�ً4̮�Nu�6�N��˼r�	����0#*��6ﰔ�9r�q��]��EWs�zw����ʺۣt�bC�a�v�{d�ymȷ���8�\�K,���z�����l��V7x������F�@w�<��9���Hc�cU�D��$��b9����UG�A��;�%���e@{A�zm�gH$���Mg%��(�B_����L�Ȟ�u��Z5~u�L3R��c�E{�QS�I{nt�5�>a�.ܡ��'��R�:8�������YxX�a>~�1�:�y����ZO(��uRU��v��LS�Û�Ga�9:�R$���V�*�͙MԂC�$�K���Wx��2�G��n���7ݼ��?�\G�nc.Ďq��d��Q;n)�ݦ��ZE3L��+���w<���<�7ZG&i�C��h�R0b(@dpnwPy���%J�Q��9��:L�5g�է�
|��I,���z𫶉,P��{���+ȤL�nLW���ڊZ�,kZ�%��	��Sk�ˎH��t�5�y�9��>��՘o� �k���<s�ŝ���{x?�jn�W�h�#OoC)g��}�`���s-ؖyΠ|vg���C����r�j���J[���GB�8�WQDuIPʆ�^]�< �؅�ڌ�Q'dŒK�U�"��uhZ�m:�42G�D|I�V^��Ca9�K��QOq��6���O�ȨwO��:c)�nX�)�t-�<4���϶�"�4���祣���0,�9pَ��>�e����O9]�O|��B~�6(�Z��O����-�
Ӈ�	uy:k
6Üb��:�(����-^�?i�p�^�����AV�hz0�����ڞ�? ��V�oP�x�fy�x�"�� �?9n���s�����c�	�:Mq�t�ϵ���~�ψeÝ<4���i�?��35�lubm�%�0=�0Lx�H$��\~���p�8��1�@������C"ٗ�.e���%�Ҕ$>�e��G������|��WF0T��N=��N� �Rn�*�"�B�:|^��D���Y���%aT�r�\ϥ�w�uq�fB�6�$�|:&�S�1X��C+Ӆr���H�/��"y\��Յ�@g%\��a�-s�C���UH�IA�;�m>Q�p��h�4������e^e�9�.����r\Q[��5�(U�W�j�5���~"�"s�S�f����.�Cm�
y���d�g��"����e�� w�i�!�B��9��� �m@Xz0T��2��V�#� ��ǲ<��t��͕����!����?Yo9!}�c4���lCÉ�"qZn�wK���A�j��J�-|�2��T�$j����7Z�Lξ�_�<͑���8��o�J.��k���ڋ������ ��t�#��S���j<������j����ǀY0<,��i[kOHT�i�lE�;6�rp��ta�ӫ{� ��X���f��NX�;��0t��@�8�+0��j+]�m-����J;a�5�;���=�Mך�S_-gn���Ǆ�Mo'u�v� x	���}��ht�v�]�����5?���A�Yg�Xj8�6ᘉ�:��RUg)�_d'7�Z�=��"�p�v*��V��L��9���L��ML�FVMʮ\�O<L��~_F�D�0`2��%��lIn����a���q���2f���SOY��J%�+�+��.�Y�eYjk�40�U�7!�<�{K�e��.�	aH�	���6Ŋ+B0i!b"{``��G�=>{G$��Y�'û��;��n�yF1J�Ήܠ�������X�m�uM�,��*C?�\��3 ;h��:����E��� ��jS���(u=�n����;W�2*���>	̸5������*:�����*}m����z��F4U��d?��	)�̸��Uӑ��r*����	���n�+�a�Q�M���,u���L�u=f8]x�p�p�,~.%�YQ��''�k�=��ٴYb%GY5�6�R�\�hUW��(b�*��3�w�PkUH�[v.�NQ.��%f��F��瘙�1�G�]g��֯�wE�ZU��}ڽ����<��󒂿O裑�����qJ,����H�z�d@��H�E�G_�}��E�i�94ueb����H �����(d �!����au|I
6x�Q����hhᏕ4+[�<.|a�k��鰄��^&v+��a��Cx��p�߽�B�Ɋ�}0ʴK_�~헬��Sz�{.x�t	
�l���ׯK������5�^�f1mŀ�$S���m��Ʃ)���[�!Z�RH�a-�m �� I��Q�
!� ��lіE�wh�I����8�h�{�Y*�|�e�|"��ɹ��
�o@�8���;��9 �N1�*n�	��
�S#ZbU�}�Ɨ�����3c�VloS�ٌZ�^��¶M��d°�$�Q���>�w�S�-�K��NL����Y}�E%N� imz��s�FA� ���<gHA�ѫoi`@�۝�ӕ�r�Y�����b�~���C(��	�=i�?��9��W\��t'b��K�_�ו����/ڕm3�^��<�S~�ʖ+���-@��m�aGq�L���:��x(eEn��R�ݎ��G������xNDWC����Uܒ���ٹqaGTCE������w����x-��`��1]r���8��:�����#|ǜ��{:�1Pz�,J�p+ <\����Gǃ�3��nV�^o�&�'L�P��c��[��WChJ�����&�y~�ܩl Ϸ���3y�K+x6v�6�g�'}�Ub�1{y3,��ԲV��K&;H��	������EPS}���'����t���B�Z������e��k38�4�BqS�xl�H��Q��v,���ϜOʤh���B\�$;>�
zk��p%�=,�-9,w#ƃ�3�v�E�հ�a^�l��A,�"{�.�����f��Jާ���*����PKd1Œ
%d�F;�0fE@lb-9��A
�^9�M{@ڀ#��ܱ��]�#\|���Ή��5�2f��/�����	��I'��g��MѮ�eS�N�iS�[�0�1>k�W�	�����3CJ�"Sv�Q�]��z�D]��k�
EraPWr���ASP��6%jH�.&��GV��� ν�XH�,$\�wK2���i���	?�T=(�*��$�\��B�)e�+�c��j�
J��)�d�a8N�F��j6��,���@�ti�X���&���J�da|��+����{�^���hG�Zܔj���������~wg�y<8�O˩66�WB���x�3�dKW�ߌ>{o(��u}� �[R��e��b���͌4�|�Q\m��8��%!�x�g��H��i3�1i�u"��z�_0P���򛂷YI0�;H����N�M:�q@t�s�hiP�������^�|ʯ����Ll��}���=����;!l��M�%�1�0��s�'uc�@��P9�`�zڲ��t��g�ߙ�o�?\���H@�j�8�#�\yf���!9�0�P�?���/�~-�UI�4���Φ{/�O��C�4�d��{V�zg@���q�I���S�T����L�]��@��uYk:��d:
N�^�i�_�M���֎kkV,�hs�^��L&�L�9�-E`��ţ� �ρ���`.��&@��F?bG��G�p�
X�	��Q�Qp�����#Bc=�~����Ū�����@7r�	`>;3�mv�~&���A	�dn��!��yh_+j�Q�pa����%��@򠏀Hk����6��+�[�_�:_W�݌1�F�v��x�蛹�9�J��}q��Bk����j)�Õ�{�Ī@�d֦C9k��Z�hp8`�McNU�4�#���CC�C�a���R.$X?���X������M�r�L=���
"V؝`������V�o���־�T��ɞ��m�7�d ����L��)m��9�t���?��p�d���Z!m�F��d��*�1�@��p�9���7я,>��D@SQ�1�K~�g���w�r�2��� �1��0R+��22��D�Mg�ޘ�zL�cs7SU�[b�̅���m�k�z^>?�R��Ч�y9\�E�c!i/n�"�9����B@����rCDz��s�&ւf ��u=٪f�=?��3��Y��1�y%[��=���rN�Nۧ[0o��wW�p��F���zX�����U2����$^����Rᤎ�j�E@I�E���2��)�܎C�C�׼}�n-�6ru2v�V����:��>���d�xb��KQ���&S�ȹ�8�B7�͞2�I5g�����LV��Y$At�i�Q#l�{g����g��A&�L"��pvF�14�[�V4�����n_]ޜ������eqP-��s�ai��{I&`Q�7���d�i^8��V��-q^�̤����� )���z��(@T!(���g�{�E�Ё2�d
�I3�'��g �qh>��tS��ڵ�B�D��Rƣ��Z$��ݨ@]�x��*>)X �Cm�����s�[t�[�-��*�w���O'D�be���m|�����_�R���K�y�-��2��>�~qJb�xDA�qLAir6�Z�r��9�Qq�'#b�-��M'rE}�(d�P�lOp�	�)�m�ÿ��?���i�����e���Vn�H�J_V\���;G��r�z�W/��O�[:|[|�)1~}jZqz�7�������6̭��j��*��٧�����#r��i%�90W�l�@��Z��jk����ꃴ��3u�u����-t i�\�3���e*�k"�����C�y�w�>W{f�&�	������L�$8��>�F@����h9>0�>`=]�<X'_��1�6�o�w[��P��5���_�L�~��y�i�G�r6�wDg6�!�=z�=c�v�K:m�,�So]�X,�l�v`r���3�)3z�p#�ka����K��)�R����Aj����o& l���#TU�y�~���AH�k_�}Rp��M?�#���Z2���R4�0
a���s�%��^�<U���)�;�B..&��E��W-6���+&8�e�/��!f8�S'd�lD�%�bi�Tk�V�P�w��� ��O��D��x@����S���l:�΂�39��f���fN�F�k�ɂ��	Y_ �k�Wia�(h9����+���f�z�9�){tq��r2z���R�cICA�����m߼/ w�ꨦc�G�|e�X�_'ȭ���]'���<��Ea/}�ų��L��k�##�naӡ��%�g\Po��+���N��{�V<�y�c��e����~�ۢ�GYKa;��D!�Ӿ���(K�̂~5�n��	�إYo6k������ۊ�NE�U���iJH����d~�!�`�~�����&4n2"�\$v��̀'�!�R+ ��|^�7���nEY\��x���h<����S��Aa��;����`�������"�%TTN�X5}^4Ǵ3���I3��xh��C�F"66X�pb���C��$��(�BTK�D+�9O*����<\�|I׼�����BcTW�ЗQ�3%�W���u��mFB�X�Q��(���Tj#��D2�<�l��n��̛����я�EfҶj,�p��!�(�)�<��R[�������*�����}Y}xj��-��5Y���RE�4$�� C��X�0Nx�f����e���_���%������y���B�^*t����.����'>����I��n�q遱��)睙2z@�\됦4Ǫ�tU��ֻi�_��k�J`�!S�/���HcY�Pi+[X�]�J7|Pk��+(�q�Q�(���k����6���s4 J���p��ܰ�Q-� Y�ǻ�c��2�Md����dc[���VN�:$ew��}���{�ڠ�t����z2��Ο�D��n$�~>2�lB�A*�I 1"R1$��b�ha�W���	�qSb!xsp�[H�e��T�!c�U�R'f�A��DBx.�������ƕ��P����[T:��l�����#�w�2�O��D8�&"��/ W��y;p�6p���FF��d�D��0��מP$�IP�k��#�:�چ/����Z,�슒ɻɸ>x��=}�!���[Qѱ��u�\0$�Y3փ۫����	Z��aϧ�:y1�n����vG��V�+<�a�Ҏeٯ$�␚S��ښ/i�/�EN	^.8/+�Vc��N�(�텷�Q�N��U�ڀ����r9��#���׬A� �����=a��Yo	{*`#��ͼP��l������o�����5�[<"�Q�O��5O<|@�B�*A�3���XVL/���Ⲕ��HR�m�6��
"��8;�Q��l��%&�l�:�C3�p����TH���ʪ�2��Ud���WE�u:ߠ+��MvZ*(����q�ѫTU��a�h���t�&z�:�9�~�Sڲ�͙��i�s�D���E&��Fyo�2��'�J0{-5�A�T=Oǻ���	_�<��XVJ\L�Ⰽ��˳>ԋ�m��-��Q��J��MP��rKeB�6D ,��#�y�zI~RK�D�=|��=)���%QxSh��9��q'��$����^k�2���@{9��CQBO�\�x'�%@A!�F�WB��t5ҭ�A".��+p����ob���Or��D�͍��e�T*��a_'�:qj�J3�Xay��h�r������5C�|B��^&ޭ
�p���k�>�eޖNf��������p�)ƵO3\3�c6fF�R��.rj�c�,��Nd��$e�����n�nĩ�AN�Dy(�==ò{��1��D$Y���z���t`B(7\Yb�VgcUh��z[���H=��^�Gms�|�5/�a#��9�a�0�˪��yz���R�2j4��q]��g���B,�e���a.FY��	����o�5L5�;n�#�5	ZI�?9C�2�h�E}�<�i�y�y��-{�-��$�ꔢ��AϢ��$�W!�)���c��'0�Ed����ݚ �zձ���h�A�B�}m�g��оG���N��I5�P�h�ܛ'�ȬVr�G���U�_���B���	���e�bќ�G��������ߙm�qǑ�*��`~��6���(C.t��G���K\���#Eev|K.��b�s���6ɧY{%�Q�3zF}u\���B�>���}KZ���.����t�+��h�A%K�A(A�´P�T���B��]We������ZK���p=�p܂��X����$��xP�>�iD�~����oB��:�"z�1�7�Q������]:z�MBj�nЬݩ-���Џ��Y"ѐ�ޕi�}t�K.6Bplo��-�5
�ŏ���5�+4jܒ�� Q�"�ŉ�<�u��W6^?#�mk2)��h���O�G@iw���(9M��7���7���r{6�g��������&�P��_k�ADE؟{]Y9A��Kcn^���nN��Y�Xn:-�����~��
)x�uVl��q?O�Ŭ�|S�]�v,�W4T�F�9r1 �ɎZJ�~{�1��T$6���M`
`&��s��W��3Ra�GORv'�a'�����G�z���#$�_k추�2����R���˪m$슐u�QD�1,�� I�V�xʤA'`(�H2yz�E�r��ߤ1W��m��rao��6����v�Hv�j����+D�s*�py�0���!e��s�F������6uN���5�z|��t8�F�|�G�x��;�1 0��r2�*mm誡b��_W p:�<yF5����z����Т���ِ~ɽ�܂�5SC?�#�R��}���\��gɳ��Y�:�Ϊ���,���q�$O���nA�Y��R���+�k�����VY�����u�����1������P�
�ʸ�B&�tl;��;h�`�3�z�t�����9d�黛o�P*�}<���s-O�kj
k44}��۠�46! �����Kҁ�iSс�K�*���[F x�a;�.��ް�8-Q(���#GB�����\g���\D��N`�z#x�z����^�3�l8D�Yv2d �g\l�t�0���ނr�����F������y�i훢��|��A�S��񮽮�I{=��UK��x$�X6)�?����-;��\�ѩ�ĮS�K�ts�������K�jݽ���"z��&O�S����I�P����Q{2��t۶�7�������`���������<\�R���6�!>͌���|\�bi� )i���nt���?��^�7�M���q�{T�žr�,�q�;� �x�	K�j`��� �'T�@���o�C��jTj�r��?|1�GtF�[�/=�<��m�9���^��P���{�J`��B��Cw<���KtN�`H�}��G�;
���/~:�aDj�:�h=���Q��>oi����%���06~zH��T<b�?)� ;5�|P}S�:�8��U�����W�Q���[�a}|K?���$Ҏ��Q}������>I���C
T���i�R���|&�Pf����~]��V/4�B���\�$�@�9�l#	gL8Hx:*���x�B|
������/nM�n��C�K��iA�����Q�"�/CCjv��~�dH��t���v����4�onչd8EFo;�R�i8Y<r�*o�7�Z�K�e�T�u�-~�w}�V�����H��i�-�f�T��N�k���te���+�MS>+�{8��M:cB��~���	A*���v|���5^����1�
�m���e��}v���4��� �o�ko�������-���&�߃�ނ�4��	��o��{�Lk/
�/��b(�Y��~��mmE�n�"_Z{OC��2��Px�m�dN����m3JcI�m)Y{�h^0�A��+334��(E���)O'�-ÖR��/�I<�9v�_WI�4��t�rܠ�"'Q����?p�����>^����O�J�+]J��C���/g��XV+��zX���>qհ��L��ćDH�����^��·�Ϟ����ff�B\�P�SE#��Qݐ<�������\+<��5��><�P�깞�Ս�bj"��>r5��Q�,�ӄX��<
`���¡���z��p_N�׳�{Qx=�;L t>^-�+x"�_`��?��^]�����lvQ��G��m�������>3�!N���I`ڭ�a]�!���Di:��S�U:���|�&Joջ
E��W�N��BJ	����%�S���#�'�p��H�4gk:�8��A�Z��d�n�~�K�@uơ:
����|�*����>�F"�m�c�UjE�@�&	����ֶ���YծW����O3�r��tq~f)��ѶcT:����#�����u.�8kn��OG?n#9>E'���0��"���K�1Iy�Za�F � ]�����;:H��$���	�j�x��,�&z�� �e�gpN��]�B?�5ί�Y����f�;�߂u�^�(^v`�k;�@�1�
�S��YYk�k	��<���SVrjx���j�[�gmg������<ZE(��p~�dS�x�>{��%)]=eN�8Q��K� �����d"��md1>x�N�y��\!��O��aQ�I'��!���Kt ��H��ߖ����:�jA0٤�A�+@��5��n����-�S�OiJbE����:�� �n�

���G�O�[szؽ�&���Z~���I��6.�C�i(bÎ�	DQHy�-5�!S� �BP�X��c���b؁u����N����](�Ԯ&5����n6�zQ��QCi���nt*�H4M�(��6Mɿ6�tm#���E	5�,���� ��ӄ�+�K]���h��6%���ld�GցL)����(�����=w�_��*���d���]6A=��_I��6io7�v�ݣC��E�X�$��[Cix'�ک&(M$��7�VZ4\*T��&���I�5Ģ�_�����y�c���ۋ?#<Wv����b��@��)���w���VT���Y�;�mγfO8���0�m�ZJ�'���H���	R��f�|-#�脏���E���o���*�Ǜ|W�no���i��|�Bc�x��Po�ɾ �E�$V�#h�蠧<o��g��K���9��WW��X^��k��܋�!	���:<'IH֥�q�>�,���%���J�ry>:a�� ��b=&|M�42h�wf�"����PC:��"+X��:{
�d(���L�y��_-�7L�b�=����;�Jt��&0Om��^�GN��~cd�
��&�6�fM���E 6����oF$��/0�q����W�	 �vcg��9�J�C�er
��4�o
�Z`��Ճl�C�~�cp�ts?3�ӝ{߸�78zkMOX����j�-׶ջ���6�o��06�Y�m�������菨Z���C�M�-������lO�� ��"�<#�S
��T��U=R�J�M��nͻ��r���\���H�5�S���l:|�|{���x���?��o��V����a�d�B6R`＞�������5�x��B��]���f�}AF�*o�����-d���՟����M�+���ﻝ.�Pp�}��e��J�97�z+#���孾ꙫR��W�M������'��հ!�FI7�|�h�r�#�px���f�i $"`ϰ$�
^\�-5WN�T�ݹdLDp+�.��,a�2�`I`���~����K��u�7��FW�o�44Y~oN�0�ѾSU`�\��VU_K����@4]��C~�ڨ��ܥE}w+Ѡ�W�'�q��^����ޫ�����zn#���]3�$��~���N<���'ӊ��sW>@�b�*`�3��Ҟd�JX���?��,XⰜ9�Q�m Tc?�m���|����#�/�|��W�_���H7SO�Og���t�@|�-��9u_u��l]��ƙ�&;�ˋ�\���u#gjaˇ)ɢգ��d�g�������Etn���$1���R��L�6P���%�8�bl�0�_2ܿ��-�E+����&�P��b�,~�)PGז�n"�������Ot��bj^�����$����&ΠM,�[)��#�[�%��a�w+:Y2��7\\�m:%�s�7�g��"�bW���
R��~SԹ�����qy��΍�;YU�� Ф��
~q:?�u��Ƽ��r�_0�2y����,�犋?�����S�>W��G("H�3�A����(U����:{:�OZ�OjASq�^�TPU?���Xś�sXfЦ⭰M\/04����C>���� ^ ����F�Ks��*���Τa�ܠ*s}N���Y6A���v�-n� J�x�.���Y��uS����_K4�!������_]�&F�a��a<R
��L��&F�2K�1kx�s���=�!�UD��{��g3j��ͬY6�ֱ0�mp龱��BAJb�K6�r�zA#O;��I�\�n蝛��{3�?�Qv���4V�T�lΊ`	�Le��2�[H�WH���]��<��7e�:c��u���U�s9r��i|)�[t���M����yjڳO��$/��v_�W�?@�q��>W-n&�b~��N|��GC�i�zkH����H�x��:i��s��t�J}T�������J�_%#�Ȝ�y3���}�Je*}�)�K�]���us�T�H����H��s�J�^G�� �B+�Q��5R�C�_��T�8MʱX���-�'z���_��L�+� ��<�U<���$r�HM�ń�#����B
`�q�oIz��`|�!�~/\�&�Zt�LT[F���,�p�Tl\oKf��E�I����Z3L�aV�0�s�����)fC=�ZoP���W�
Z�
_���(uO�p��p��K���*������Ʈ�j��m��|��
�{��m���
�[
�'���H9��,�q2���XIΆ��^E�o�% �Z	�r�7�E��G���b:>q�/����I�c�JJv���_�N�AmdMY��5��qq�#��S�y�KCwlo��^�#!L~jq��Z�1�*���ޒ�q�\��5�/���O�W�����Kku"1M�P�69������F����z,+�6}a����<�~+F���9}�~R���A��-��!�ĭO��E&^����e��|��";~�%�|kt�5�_S����o%��
�*^~
_�9���
���b,�㞬�¹�Y(���Ŭk��?�;�EH�}s�j�0d\�{�v%�`�[x�l��MT'�kaԑ�0����$�CB������F���|[�_��̋Pn	L���%�]�_�r�e	]���')y�Ѫ�Bռ��|It��%�W�H��$A��$:�sU�#l�g[� Y�>Ӹ���k�l�L>K >�_"��v#�*�t w��A�9n�¸���sA$��	��Sj�b�S<Aơ�#�G&jL�<���3I�Dɚ��5&n0L8M���0M��4�:N&m���$L�3v0e�(��Q�R&l���X�%��5�0�z:�i\�C�1�Y�-� ��W���:T
ɬIR�s���������-Q�P��d|9�������Àl��#�L��q�f۪�4�ީO|�7/�ɇ,�|�D~��\��x��	vV>����
���9�Ms:�k�
��e��c%�E#��-�(48�5L8�F�
��!��D���)�M���;�gi�z�U�t�n/��,�g��J�T�V-;�d.Ė�'����O��#�3<]O���RX*z]�l��Gٚj{�;�1m�Ŷ	���^\�z�V�R(U��T����g����zI���� �r�T�����"��E���R��H�Ĕo�3����RH��za����w��&�83$5bVK�o���!&��M�G��x��gr�n�Xq���5���K��XfKj"ot���hג�#�,?l�'D��/���I�KUFoM�ZxOP�����[=rmٷBXZ?4ʋi�YV$�� |J�#J&1��e�U1t�+Y��5�z����l�;>5��m�+0�Ȗ����n-��|xvhbN����oT�`��5/;��͟ㅗ1�X�Ѿg�if�����S�5�_lb�k5-�N�k�乨F���z�Osl���h<'�k�(���
@R���6��BM[��ŧӊy��,���EM3gVyC����Lk����Q�RV3<��?^�7���^������o�2C�OY.ƫ2-ȼ��(�6������U���c�w;�����E5N��bG��_PRd�� ���5�k
1W�7Q�nCA�lB���:���a��c�%	F����#�(��-R[��/�i��CX7������l8�1;��B)7�s��M�h�S��LG�~~b�}���"�K����wȫN�3w`�TS�LW��El���䭽�<I,j���&�W�`Q���r���.�H\:��(�2��t�1=g	�FeWc�.�ؗT+����r�D"ң�Y�BK���O^�ĝM���ſ�<�����;5{��Q��V0���n����Ls�_�@�$;�]���J�䯪y���J�L��FŨx�=�i��UR�^�*LP���k�+N7I�E�EZ�Ԥcl���tY8�̠�g��1ߪ8-�����U Z Ex�1ϋ�����M�M���W�>5ų��
9�O�_ʹ>�h|.F�\ݴT��?�WW��r�-�8xcr����P=��1%�OjE�,�8�5R�4�Jǅ��U)��:T� ߺ��9��,p��XYcAk��n�� ��'��� M����Gɘ����P��y��� ��b��D̜Py��"�v�Kʪ0@y�M�DS(o_`^�f_�?iл���J��ѩ�)��O��8`�-D��� �Q�_m�\1��Vw��~)����R���� �H2voԶ\�
+\��W	BZ�ԗ:J)y�'k֌����������<���!�X���@k	��6��׬o�V�,����Ώ(U�iaܓ�pϧ��b�(��iF ��C�6JΡ��;��sUs�n����-�\�ȩھYl<������*<Exlq)(�W�#�,M�C����:�����!��(E�n�o(�����a�b|����%>.�s��U�ȍ&ǍƁ���,�:�`�����&���Af#}��І9î9�8"�l�?*!�A9bڼ]|; �]Q'*��ZA!.����r@.�A���H��:Q��d��Q�m��Q6f�-W��뀙qʹ�;�Rf,ά��n��@���QrX�XUye��]�ਬ���*#�ˎ��O4�?T�� I�\�x]���j7-yn����t���L���ƶ'|���G�\�M����{;�HԘ��:F��k�d�H��}B�N��l�jFS�5�k`���`��Dc4#P�P��Gd�����v|��3���I
Qv���~�W�ͩ���{Ӟtws�E]T}ܮ\�c��I�ˇ>��œ[����{۟
��//6`�e��dncg�;�e��}���I���`��99��ns�c�P��8����"n���FU&3 g
^��U������� ���	L���v[��M�y�:21՟d���U��j9�,���i�4��8��.��lH��Đ5ht������ s����O�A72�b���/��[yDǈp�Jh��_!g|wO��)�un�6���?j�X�ȱ���~?&_��O����
I����m��+�>MD���ڥ���j��8g&�g����Av(��s�#�m�p��jo%������^7�V��V/9I���HūĚ�w�{��<�!L�t�D��d醿���rL���jf;��&��z6<��8e����M��Q����T�W�B�M(��f�W��е�j�~mR�?��羻:�v9�� ���������5,r�D#�A�8�9s�%|��A]&DOgHqp�]Wcaݴ�^%���s�{��Zz�A�^]��r��]aQ� xp�r��B��-�%�p|)/���Ǘ�ƞ\�X#*4�U�jb�u,�psQ!���,ᭊW�-�f�m�IYV������4/YfW� �4MJ�&|>���X���Lh�#�g��f&�/:��[pS��G�IyU;�1���3����[h�oN6�DD
$�: b��Q ��;�'���7
�ǥE��
/)Q�d�,z� 8����%���W�e[��#�����Z� ��P]�+Q�*�����8��$H�t��������q bT��@�zp4��9��*%��?��M4 6`&�(2.F����Hu	�l!��� 5(>�l<��;��@��ddG��vo ��z��4��5����w�(�'SB�FԊ�J�������}c�׺T;�iE1��{��
R�N�|1J��<4�߿X�:�Sݢ������� }�BGC߆���QA�I�l-^0�����7n 6�Q���J8RA���Z{Bh|lD�Cz�]�4|�䤣�A�֐������0l��� I��A�2�-��� e�P�5c���7��9[�v{�p5{C��_+��&��h�u�N�&�AR�̶v2D�_���I���NyiQ@�~���t�n�t�%���0EfR%é͒�9qQ��X9Xs��:>���F�#�UW�T�Wˤ��@#�� ��n�<��nZQA��;��BC���j��L�S�'Nr�:��LӻIn^3��N�M��4�:��5K/������!��o����4��T�0���jM$4�jP+,�"}IsL"�Z����B��q�=�\����ٙ�/��˞�e t��S΢���,��6�l8���*KH�N"m>�٥����$<<V{	�/��;�t�^��,(ƒ@¼�B� C���*R��;���3/J?�Q2 콦-�NBE1ߝ܀��sba��*!6(�+������ͩ+�p�Ma�P�U<y�wY��K"l��#0��D'UJ��Fcc�,z�r�T�:b�M�����3L`vg@v�_����0L�t�i�D�l��g����9��E�BRg�Z���~j�*BX�4\Ӎ|���2�M��-�X6��v�>��~���M���#h*�JA�y�(���X��S��ŏ,lx8:�Z�.\���>�b��o��8mW�_��Z���Ö��p����O&�|���v)b���;�=4w�W֑�F�#z�g�4;w�s�P���	(*LyW��P6q�X��u�p�B���J��C���){t��PLT��a�=�;�|I#��/vA�W�`֡�;�X�UKZn��·7V^������xKb�kl̹*�.��m�U�3K?{�TPd(ȩ����B�C�%z�@����27q7 �������W���F���k�Aj���r޸R�K�A�>��{q2-j�$��̒n	��[V�Xd�C}�tzv�wTM(��)J��0�l8���lb��W�>
��f�*|�?/����(�f�"�� �Kb���ת�Kd/@�lE��֝��������s:����ȴ؉�
YL����$M*|=0I�� �f�MN(��㞑PȠ�O7���kG��|@뮑��pwY��0 Bz\4��"��Z�H�tDy�h:�Dm�ʩʢ<�[G�n�P=Z��~�}��TC+$=w�������ظA=� ��fA�#$Gَ�#�b��}�
�*���m����������Bժ@z��w���k�����	��|��
>���Dr��{��?�o���|Oy��O�5�j1�/�1h	��t�s�=X�E�!Jya���O��;����"�����*�+q������*I:��*���?r�1����|W|I8)9�m�%�W��R�o-_'�ז�����H�LvO���A��(j��e�E�vh�'���Ky����Q$r�������5�4Z�cA=���7S��e+�Aפ��6���gMk�u�t_v�n�ŭ,0z=L����GN޽j�'W~u��;�I��JY� >�Y!���>�A�u�h7nj�LM{�p���t���Ih�H ��iTT�3X<h�z���ҋCX$C�y��R�H��^��z�c�ɾ!�2��������1i�M��ʺ'\����䃈�I��C-�<�Fm.���!�[��u�E���
#��8\�%أm�J]p��`
ΐ�rۧ�	�f��tkٿ����#=ӯ�Z�A���-�9'L�_:�i3zSnw
+�Eɟ�k�F�<'N�P:|�j=���3st�l'"����2ϯ��;�.#,�+��:��	Ƽ��З���Nzr�+�R�:96�f:�B�)�ُ�B*��rＩjX������ċiO�y��-'*~�>�ƀ�/h�d�W����bӶ��>��r����Pz�+��;�<>��{gܰN��.y���y�迮�TB�* T+�M��g�lX��sP�ꌧ���"�j0��'��h��ꄟٳ�d�/�"��%"&n�0/�ҋ�څ܄9��2���u�KS�K#����:=��s��C�^_��.y@�$x�R�2 g/TMՔ�����b���<F��w�)��K�e��D�ʔcp�k|�����u�ڨ�TU:��F'�i\�k�l�2��e���>�je3�:�������������#s��Yf�.�p .C��s�sw"�s���iw]� �wAz����v�P��-c~�އ�<�VY�w�;`���\��Mɼw|��Y����hf?�g}B�?�ۊf3����F?��{��~��>��R^���F*R�x�#�FGj?_k'�,)�I�-E�������=p����ǳ�/n $���y�|$�h:tw��/$8C�t/�Ϡ
-�CU���e����aPN�L#�z�D�����?H�2��9�:��;`L�X�(�D�J�;&ڮ�͑��|N���9\�ڮ�ӈ��(rã������/L���[΀H$4J����U����O(�̏74�	F��2�X8��RA�u�z��q����%��S�m҆�P�m$���$'�)�4����.��y�c�v-���j��	������Y��K�1G��0����B7C~O9�u�JO�)j!�^$�F���V�XXT�Q�#K ������B�Ş9�Hs��;I�k��������/���&`o�x�C��r	��Qm_������z�����s�Q_[�-�`;�����>���S�Ó�n���)ܖxX���Җ��$�|��E��澫��'�7��>�h��8"k��G�Ѐq��~� �xʄAqH��H�����c� qT����/�\����ݞ����F"�M������������]���Þ��"�-�s�U�S�aT���W`? �r|�6���jR:�`�5�x2�A3t�c��@4T"�D)="oH��*�Df�BSb���c���rG[?���`�{*9u�Gv�l��"C#�W7`���_�k������-?�#�B�B���0�˗h>���3 �`0����f �� cV2�@	��(۲uW�S�d �S 3��z�g�.X�����NLsx�f�i���q�Jd�'�y����6_��5���R%�j�8]p�!�Y}�?���,�W���]6\9��b���<3���ڂm��H����X����w�6���T!��YlǤ�a�X��N�#a��� ���j��ٍX�mKVC������=��-}�;��*5W�c�@5�CM���F���|mZ���e�c��aj�A��Λ���\l2 ^�l�<H�2������(��Œ}�W(Ux�	tYMy1{�	�
�!�r$l��PN�Bsq�#AƋJ�k0�ި8}j�?҉�$R�����o@��7�ݣ�����L?
&
28p��eD�D±#ylġ��&���cΫ�<�;4 �'�ǘ�%�OD6W���;���Eh�5Y�A"CY#���ǢPwp6�i����Х�6��H/�k%}�3MA���@*���I+�Ԋj&���Ӑ8FU�?�'�|i~|���n?Ɩ/<�钐"��V`���u��уXR���H��j>�e��Ž^?�@� �ZC�0h=EK�I��O�e%��������1}h0�GS?k�����Ө�iA���`+#@�r�#gP]��/��E�`����O���v2�;��Uz'���B�c'�;�A�6�	`�o�N$@�	쭁`\�O�>��ftڛ�̵7di��D���LM`'����m<�6QO��^�Z8YS
��=��#kaI�� �#. ���%AEa���v���J0����E���b#E� f7GPѤ'��!1�� �cJJ�d#Jgc&��K@�BS���1�Be�LAi�MGEF����;�� ��a���H�3c:!V�I=b��L����ڲ�uit�#�8�N��ӆ�~�s۷����R1�%zGA��U�'
�-+����eS��s��4�mP�rZW
i��^������W������ yU?J6Z���vˇ�J�gw՜?���0� _kb��=������M���Z0�S
�b�M�O__ƌgc+��K���<A.��[��'SG$G�r��ج��x�8~�u�	��r�i���\t�ΦZ��<��ӭ>��r�g*����7yE�@�k��G>�Qle.
F��@{e�uGࡿ�Rt墧�1���v9����P���^w�DDZ��{/o�|0�*!��t 梹��1"Ń^�3<�\,���������_8)(�q8��;�R��s{��4@��q�x�!?t�3?�40{�>��f *E��Jd1�pŲsH`���r�o&$��q����>\�'�:xi�뵀�ټ~��`�=fns_1���NO����7����?ɟerч�p'�VN��Ĩ�1-������vm��~T��-��%�\��Ws��6S.w�'|*x�LyRJN�m��l;�K�@��f��ַ~�h�O�����i�;h��u8<�jU�&��!������~���^XX����BFg$�\��@�V�I���E[��2�q��[�A�),#K5)�P�c��;p�(�ti_��D��YnAi�-����Tbf�F��
�nr�u`�h�҅��C���N�F��ӛ�,��-�F�@���q����\��=@�ؿM���ǀM�/��� 	���Hn:�W����Ou�\� �R"��i�a��u񲰠o	�ic�N�c3< @O5�[��}�Li��.�9<�'uO�Z	���E�v��+.z�r���h�Q+Ds㛤�m�Z};m/l",��M3�Q�<*������W���AG��f��)��<�<�ۛ�L��������.����d�	���|Q�6AZ�:&�fT9�ӡ�@�ʡh���+ܒ�~�UAa9re�QB�*�%-v8�D���cR��,��Q��8Xc�c���Dt�^~���Z´+�py�L��ێ���	�GMN؛?�V��u-���%5;D��>d��m7>�v"d�>�@����y�&����r�%Yc��:�Rű�v�u�NR��
鞛B������	�����X7�
^�wO��@/�1B�s�H>6������>��������}}�������k>9M�ai�ɮ�n����2\d3�2=��Q/�v���#V��9�v�
�?2QW���1�qڛ��4��W�EG� HB��m�ƞ�A/{���.�I����b��m��k� �`g���K�y:8F׏'е�z��%����'�O �2xbw����X��J�U��YP�iY���&������S�[���]�t�Q�P�}���4���%s�)5XA���F�����0��(
}�6�S#���v/��8�[v#���C���OϊZ��8.l���(��_^i��|��\������\�gLh�=&�?��=�ʦ#侍ͯ�8�fa��3.G3���5��?�|7?���SS�ǤS��V���R᤹Ȁ\�4M�Y���W��ї���
v�vF�5ɝX��<jb\`���0FFj��bm�7�:���z�z">yJ"L".L1�F��Й�1�A��\�ƕ���r�@<c��)'3�\W\�l�1p��>�sx�?�&�5/?Ƀ;o`6���C� ��O��C���?�q�c��TB&�	&H�)#Hč#�5$nH*HRHbc�=��	b0�d�LOh�L3|��{�L���LK��	&��Voτ+T�J�����Qe[�Qi��ł���]�h�e�+��~_���&�4Un聍3����ï"�89�85��S2t�' �NE
ϡbj��Gj�;�5�%�R�L��j4�
�tR5��(6P�Ь�nm�Ǯ=��Ӳ�M�d4�3�`M��:�9�iD�Tq���E��Z�勺J�$I�ݘ�u�b����=���E�ozn��	V��\n�6cCqˤ�C��M���7w��ŋ�Z��0_��y/VP?{���?��OXP>�a��+��Ln�,=8U��W83�J��z��@Tn�8���<� :�	�ۿ��P���s͌��X�+� BxOTdI�4�pY��a>�))��ŝ
�/��By�x|������mB(�J�Q�30��q���ɒŘ����y'.����{1b�
OU��k?�9JB�x�O�Ҫ��ϕb���F�Ī��^�{/��U��~[��yq(j#����_����'d�['�$=�%��22!?H�%���C��C����)[ugkU�{T�'�,/	l*O�fmL�D�k��7�V�>�T1��bt��~�$�ݐ��Qf61�JnSLECƾ��Q:�aI���E��7H�އ�ŞD��@���~���+�����\����ģ3M��!4�G�"a1�sZ��S`��4M�B��%7Ì���r���Ҋ���}��UW{�~��d�=�uc���o�������[�b�O�S�3�R�eU~HR;�цc�d�Ea�|��<\�{�M�6�����ʀq��.�x|y� ��.>inPF��kQ���2b��3+�V��=zO}�d
Xm�ǖ��w6m�SZ{�SzUb�q����  @���3������D�#�7H1m�LV���٠Ƕ)���	�X��n�����W�w���0���k�B�����1nӺ���tS4lT�7'~�*Q��#P�~��~S�M���=.7Hx�{��c�ѻ�0�l"��UM�e����]���?X~��Y~-�f��~~��d i��J^����@6jeu��sGV[н"R�'�μ%��ȺS,7�ڜh��k���XA��>\Ϸn~���>��UT�w�/[��B�� ]�8m��X5�oh��z_{���Sk)r�Y�WdK�8��Cf]�6�{�߲e��1آ�H>e�.�ʚQ2��r��9bk��Oc�l*��t������#(��or2T[[����_�l[��ZǷ���+-�w����BL26#%Nt�@�W�X���6b�����ۏ����^��WG�D���l���/��z�����pc)��
�V?p���Bz'Iw�9�*���n�*P/��������g��ح����n� Zleї���/>��krn��]��Q�i���]�:���\	P!�nbP�*5�#�D]��W\3��Q�}W�EY}l� k`�!B-4�q����X_�d�-��i���O��ԠN�o�eZGГ}ڮ����^���%qm�DUOʙy�w��:����hc�_* {C�*А�Du�w�@� }�6o��Ѷ��z���mHW㝳q{+V�Y���dd5��\K�O�X굤L��:���7Z4���#!7�wC*���ܱ��Y3����JdW�_�i��V�~��(������0S��\�ҍ�A����1��»"3C���ĥ8�n2�A��p'd�f5�E�� V"�F�@�(HU�$��$�U����ɋX�%ծ:8tb	��J�Ս��e�ቸ���2�|�yq�"�H�LR�8�Ԋ)�Xo�se���44U�t���ѨF��Fj�1�p�"�+Pb�k�Us^N.n�n��Ys+�n�,���=��þ��4^����Ł!Z����&_��jD����w�7>ܮyv��������"��-oE����<�-b�UYT�x?`-V������e�����fz�7�-;a+k^�|�i�o�&_��	�;Ȯ�t$;�4{S���R"���َ�R��M��x�k� ���r�y�$�2����Ė��)T�V����jk�x[\��+���Ti�K�W 7�]�j#���{qqu|��wj��������C9j��Շ�'���r�f]=2M����-���³ѽ��B�Յ�k�jt�.3W'�4��d�~e�↕���s��D�����\�)��V�\��!�s5r9訡�*H����m����%{<oMw��m�)k#�ͳmJ5s�0,�ad0Y3rЃ$�N�g����r�;<k<¶��? �|���%�T+�ܲ �ʈcY~�.<:��>^�\���۠Ԧٟ�7>Y~�t�K�m��}��\��v���Y�2�d�	�g�2�b[�7�~��ղ7P�T�*Qx*�������卑#�����
#��岎 ��!�j�[�H��9���oK&���;�Mo1M̜I�e�� Yq=��k/�G���ø���K��Sh^���՝�ق���bl�*Sb�}�]���Q�ׅl��k6�hN	g����@�w�B�-�Ց�A�b�ʢ}e�	����oY�Y���1�uHd�_H��xc�7<�z3��\�[)���J�����p��� [�Z�%k9�8&���s�ӹ�tM�'���~Z����##�\�b��ڈ�q�	����/U�s�a�rw�Z����/�˫�3Zm�;��9����� �K�<KE��H�n�����ھ��_d��ԝ�&[ses��Q^-�����"��r˧g���ɿO���V������sw6񱶢9�ci�6׽�~8����>��o�p~�����m��.��m���
m�o��2�fl�GK[���:�ً9e��6m����9뙜��ŕH�p�Th穮�������������}>>����W�hw/7�k������a��5�fZ�=q39<F`�@���YC��\�b�
q)�K�u�_��rn���%���Q�"�af���/4�Z=&��L���׻��l�k�w�~���Fԫw�t6@�dcX�{{�����1��럌y#��3�#�3�N��ƀs�?7��3Y����5]fC����f��4-o�f�U�%�s��q*^kk�͇Q�'c�a��C�3�|��p�% ƶgͅW��(]c�`
��e����±$��
���@#�	�h���\��&9���bZTr�R�����o�IU�q��������|.��<�G�Yhj�(�GB$T�gc��Y��0Q�Gz�<�BhU=�"��)/��&���p{��EC��j�8��\�l��aճ�x�fAd%"_����Z�L��/�Y���5}߆A!&���΢��� �y��u�t�~�P��)^��Qc����βӉi�T�N�M�ҹ|�� q�ԗ4A}����S�w���R�,�38,
MtU�RR�D�b��G�  *��cc֥�F̍�����&��O�}��˾O��!�ޱ�Y�Ojl0�1ߞ�/c�����4~�l����j$�L�������x7�m(㢜(m�(��ƈDN,��b����q�p+���]��W���Qt��<���1	�9��>�#:Xo-?��x��T-�k����)|�̟�'��y�Oly�e�Q�_��a��-�4�9Z1�u��`�>�Y��A>���t|���x�Y�Q�Du݀�zΌ;��1!t�#�G�������vc5,�s%>�W>R�	\9J�QY�S��=�����t�:�����'�$Æ+5G�ˎ�l-��/��i~��ۢ�g(���u�*� �?��#����%3<��Z�#T�9oOU,i;��ldzLŷ��s�0��� [�at�T!����s��1�����*����e˘����`	t+<o�B#���MJ����}~k�*+e�<.V73���
6=���e�Éa-����5��`�iҋ�A��n)�^5�F ��v��f	�@)���٦@]Adݥ���oF�����?uɐ�+̕4{ؔd�{$=a�&�§�0�C*炓��um$A.j��3�G��Ņ�ͮ�\dJ���M�Sr��\pD�����"h�}$'�fƙ�����lc_٩�Y�GNtX�3���KmK
�~�S'��n�nٕt�����"_W�#ck�Hk���&�$ey�p>�n�����ٛ�i���Q�Ǳ�U&�WY�v��s$�l�i���Ơ�K�q��p��Q�.91su�A��	�]��Sw�P4�D�gL߄,��2ny9�;e�9z�&t/{f�+i����|�����m�m�s�8��[v���+S�q����*�؎ǽ8�����"�g��j��$���r1�+%UK��6/!^��m�J	�795Q�9��I�ٽQ�|��Sy4/&�W3��9��[dc��2|S��og4b�iƭ	���u������0Ug�&3�酣�5�'�HU�q�ճ���v�ӀܓDt]��{��!G9"��՛Ư�f���v�5��c��y��vC!���K��#���9ؤ5|�R���:�" ]�2��3�ș|I�~8t�[[�`�����DdGp fG���mB
%V$Ab<�*��M�����*<�'��j��=g�%�[�2�r��q�̩��S~��S��]'�f�%ivӼڬ2���2)G����f�m����7��6�:vK�i,`Ƕ�~aԝ���vm;v��������*G8�9�=`��_]�Qb���S�Hvsͻك�|*�-�/X�6���y��[���S��o�r"*�n+wMsĄf|d���M��8T;������(O�lp�0�H�ij��D��27�RGb�Y����>O��p�������3���d��Z�]��e-��_��?u���ؒ�+��o���U0���f�0UmS��\F��%}N�yͷ{�t���s|7�g��OI�Z�##���x�%#N�y,��C"��N�b�K�Y�<r��n�73p�O���ZսSlaN�,��<!���;��k�MJ�������-g%&��'K�$��_L��B��2����A
��haP���p}�j9<�D`*%\�Jx�/#���c�;^����Yz�!NP��ĥ�a��C�̰!Qo�;��d�	��7"����kk�ؑ��i��Yj*����I#��.%�Jk�Т�@\+��+��˿rʉs�-ʙ�:�n��DA��<��taw� gp]s���{��.?���-w��R��t��8^*��C��B�0OQ��,p�嵯�+ҥ|?��dgD Z�p�N�PXsQR���� ���;�&�hwT��34ib�xZ�<��ݓØ <?Y�ڇ��>�K��8���1٣\Jh z h��N���~��K�ܰaj���a�2�W�}i&��N�S�
T�i�r �cn
�9F�P��u��{�����W�5�����NTbmZ���BZ{��5Q��s��du�m�VJ	�V��9���!�:�Т�8o��O��mAؾ.N^���
�޳�X���r�pTB���ξ�S�. V��P�h0���<�+��V���V��S@|��p�^������?P�T��H��/Q����w!�qE�:)�I�"�x�l�ϡ��S�M �i(�T�B�zsM(���H2p9�Xv⣌�;��w\R{����&uM�\��f��-��6=��x̹1��Z�n��{{���$���<>\��OF��B�����P�t�bT�k��Zi�W�,fv���f�"�\�3GMN�$� ����JLfm�����fEW���5����M-&]/N�ُ��%뫧�FgLֱӉulW֜y_�� T����,���Q�a^�8��V��pM�hzƚ�,Jq�
�G�^�������)�s�-���G�GQ�5m]�q��N��n��휴�K�O�y�x�6�{�\�Z�η��Z��z\L�Ra���Oj�Q����4�g\��-�������-�L���|����y���L 5B��Ag����(�G�ً��f��v���8Y�M.S�ǱO�e6'��E�/L�`���d��+Ԥ>ȳ�[m5�G=���B��f*��[�,9�*z���A��+�S��L�x#p�#rd�М�1bR��bR�'�?��R���."�b
J�ORy�L2a�/�#�ՃL�Ju���00�[
��Ksb!���oI�k὾��ܱ�E�Z�R$��_��Ɓ�����V��m�d��i���q�a\�z[�V��	]�#3�?^+�c���G�F�BnL^�C����o�C��`����ue+�؝�:�"Ƣ<��_��a��˦���N��E�'��r8Lq�X��H4��LzV�L��aZJ	9���$?$^>Dp�謘6��N	����zX�>�zYnvҕ[xB�����K����k�"�Ƴl��+_�����x_�(���ܗ],�]]���#Qc�<�)��լ[���؜D/Y��W�_8�J*��O-���{��';U�� ���)xC�h��SP�%g�	2�)"�HyO/Yz��d>/���@�6f��u����s"-n̿�y]���|�aC�(8Rh���=����v���{���"��q�-�ףw&�2i�9�Z��JL�C��V�����9ZdȂRy��Ҵ:"�4.�<�D­�G�]�f�z/.��l�Z���a��^�v2c�eiYp����8�unX���_��(!��S1����F�riLy�q�����DbjG���)&��$V�
<�M��v�k޾�ٓ�Pm"���H�/�������8�X����CU������V�G�fxa/��Sk��N׎+�0zX%��M���� +/��EJ�~rdg�_�9�$���A8�ĥ��������7,��'���J�h�2��,�s)9��&ꋏ�x8R����P��e�Z��u�6�k[�E��6�R���i�Z.��C�D�]@b[d�/�te_��ڢ��V��K�ν��^�C#<��ٯ�쐭v������c5���,�,hp��:i��F�Ei'���
� �*�1����J�:5943������U�[Zx�����S��-z2ҀV��?;��m����Խ��U6�L�v�}.�\��ՎxZֹQ|+�(z��m�s	�����L$����/��d���z�VCd�%�cs�܄���g���$�j�L��~�~�L�:�>D����^�e�G>�N�m�$ɯW�qx:����Q� ���Vх��6��+	��="�~QG�$�e�*�Ϲ�-A�UoQ��E͑ς7 �/}g #���LYT�D�z	���^����!>�r~@���}�)#��P�Uv(J�:oD���1T���@E���=2�N�E4Kx/H��d�1ph<_��B�9�2��N�>P�����MkbK+�]xf��������Ib�0*�qw7���>u;������=�@�d�r]��0(��k��n�e���k�L!���A��N� ���2��mE��������$�w����ކ�����^�h��45(�42(�q`ji/�|)��P��y5F�2�ɵ�)A>S�%h>�Lwr�Mi���}�UY�շ�r���E��Ջ>������(�P.����+�����1��nߝ��z{ap�۲n�m[{��x���.j7P�3F�Q����g�S�.�4��7�6�V�1�b�I\β4孷nR���'��RefDA �f�6G@b�"��̐l�^^�{���Jn,�M�ͺ�`R�:�6Cv�hM��~��{	J�xt��~7� ����;n�W�>��-���q_�����E��NqYt��9� �#|D!*Rw���fw2����U��塤W�p2c�V2k�埯�]���L9�f��u�'-	�j
`�?�,�nE_-����;χ���ڴ।�\���q���FI� wM��!�[z=�Go�|O�o���h
ؒ���d�HB����լ1+�4��'���3[	�����S���q�w
��b�r�pΑ0S���͹�TB�x,J�Q;1I�Y�-Q�ˆz�����|&X�U�"�>u? ����>)̝Vn���Z�RIr�*��*90��ky�`5����569����e%Ɍ���L=n��eM���l���T<PZ�ִp��2oQ�!����B9�M�zƫ��Db�|��Zo�r���ڒMl}�R��ޒF�����឴g���YxdC��\M�ܲ7�Qn���J�h�ا�.��6-t�6��N���������m�x�L�j��!ҧ4ޛ4��8�����2IS���&�ӏ�3Cu�����*��7�u;k[F�Za��˙�<TY��+`�m(����D�+e��*Q��d욾��_�� ���b���h�Ӑi�uY�����tjQ~�T�&^�Y����)�d�Uoy%�$-�P~��S�Nױ~4�+x��>�E∹~�f��"t�Y�V���5ÿN�(aɿ;�l�b�h2�3Q�_�b���^�&m�z�Q�?�0�˝ �L7��wW�(u�6��? ~2c8-��3�p���c+j���+������R���2'��V��DU�s?iN��5&��/����%|�1��Kgů:�:!���9]$��dx��Lb%츻���Ȓ���~��<���N��o�:�K�/\w:�a<��8I�o��
���DC�sNE+�B�o��C{��@�+�a�<��K7��!T�L���m��ٱ{�`����%�If��p��
��ԞKM���d)��'��%��Ϳ >��^���zNPYJ���GI���^d��W�Oi4�s�; ?9Dh�C�6S�w��9�g&��ue4�S��t��q;�,���f�~T縚a���A��P}z��+���ʻ9������o1�5�5��CҍS����?;e`��[���n%��m�b��s��u�lgO�����/-���E�+�]�;$B�frHjJ�ً�n��T��~)$'>�{|�%�D�ZJ
Y�J��~���M>�4�����gW����#�P��P���$������I�$���ɬh�%���fn�	��H���2	h_�Җ�"�Z��ڇ��I�����/JjW�n�G�/�/�����1�ސJ�P�|��I(�r	H>�x
��<���a�~��u�a���c���~c��g���gBѤ ��~�Ʊ�ˉ��z�@�hZ:!$�qK�u��(��J�
%�U�	�OdI6$b��QdY�8)��D��� =A��ڀ��Q������Wz�7��U�`�*�'QrO��*z��4����Q/�ti�D���m��Ĕ|���\��t
�:c�Yp�6���3QA�G�%<l.�K�T�NV���i�Μ�N���7��f�������ۗqeڙ;��8N�[�F!/�zz�{yj�oJ%RG��B�>�s��27V�"H�?V=� �����R�f�;^��΅/�dߑˎ��q���S��$��{{�#4��J��v�cB,�����|��T�v�^��uݚ49bE°��!����VrMv�U����l�	���kr០l#�jx϶й���j[z�w��j���t�݀���.<��^����A^���x��j�虾3��t���<��s�v76�oOlb�c�:8VKy6���/����X�}_� ����@7�e���?E�TgZ�}��N���4��nb����tϕ�V�j�{Q����P���x��4��Z�`���08��_��3����%���M��w������S4b�W#�JD�B��&x�Qm]��~y=赽��Xgq[��p�w=h�'q�Q�{���^.:���������c7��kmdc��y.�ɸ\@׹7P�	.�ϫ�>���
�Ie'rnN[Ј2c������-��>��)�S�FJ�M܃��>�!kGX8��9�%��U:��dó���)���s��~J2c���Lw����]ÌZ؉�
N>���j�ށKu�`�W��0��g�P��.�{�Z�¶��C��|�O���$Z/��
�vǷZm>x���+�=�����*'8�e[9RMK�
��Ґ��i��)RO��K��Rk��'|#Јw�9��]>�k�H���E��f�+�W���E�Ȫ|�?��I�ёA�{���̇�V�.�ק��|�=�JZ�'�1�(ɏ��Up)���Hf#�c:�B��=��P}��y(��0���1Z{؉$��%�����n����S�qtf�ɝ�~_��xn�(�
��/�˴q��kv��8����S�Oa<m�z�O�h���Y3{_���Y��(!�[�	xB�#7s�����q�h����G �JG
X��Kf�Px����c]��2��ɴ�	v�©��~]@��9CQ�[ï��h���:�z���:��u"O���N��E��/?��V�R�׾)���ɲc�f�j��9P��{U��m�����H:�_�oC;Z�Ri�[�3���礆T1�`�`vD:(�9��=0 �}��'9�B�	{L����%�*q����~���U=-M*�VC��q�㠒���@=pY�e��^��E�>y|>�ح4�5��:�`�]�JO�WyVl�������:|DFn�㼗��㭖<�<�|�le6^�I�P��|,����)��a�Ў�Z"�-��]+R�Z�u��H�,~5~���VJ�6��㺚}��g)lp�sQ�[?f N�F`:gP;��k��GMo����R+&Rτn8������=ok���U������t�~���IJ>�}3�Rh~�1?Z�����Rꒈ���U_���\U�Y6���2�FiD�X�����%���\�O��剴�_&�I�Z���4�8eҋ�
���rvS��>����5$t��7�w/��0�D��ԷS��F��_�&h��-�,ߚ{lP���n���ء���F/#K���B�h�v�:�9���g#W�L���3嘵+iNx�G}�<Fv�6ֽ��_�����g�"Ґ��$�&l�R�����c%[����S��,~�:=���Eks�|���2��VyPr� u�$gO��ӑ��X[������;�0��� �]5�߳��9���͡&���[=>�����W�y)ڇl�������/K�@���r� �_��6��(贻���)8=)ոp�O ��5���=G�0�����d�~��߶�H�P���	ǯ�y+!�:X(�a��� �9�u;�7TW�|3���RԽOvУ��n��V�;�^S�5���R�Ĳ
��voWu#�q������`K�<`����q������oC���:����Z��� t�T3��I�<}��㉱�;��Xn�}dO}�?�K\`��O*O9��ӱɃ�<��{��^�k�vmn�p��a��?Ƿgm�S%�D����X����J6 i��nD�Z�,��x�Y���QFW�����v}�O�E�q));��q��}SjrӨ:���G?�M#�4۾O��#P��y"DU����_/z}8���:Rt������ˈyK<;,�|5�X̫A�q�k��8��T*ک)����R\��7&8%
��b82GGTp~
05T&����aִ8�S_���a1��ЎJ���xQ�샠u���l /��m6 Z|�ο�px�u,`�-��fJ,��𭫞�[��켎.�KX��:��O���5^x�� ���3oe8�:.�?��q��uv�`Ժ�@�M����O\� ��������w?Ij9�o7�p:��)��2�}5u�OQ�����U�D�ؠ��݁AP)/(�[���?Y8(�I��H���6��wK9���z%�����M�-�'�Saf��4�hl�Kt!2۪����H��hR���RZ	M�H(8=�:8l��i�@5{(U�����y���7k�� ���SC�<��z��+����o���uC��бE�P�Sx)L� ob { �:S�B]g.�X���ػ	9�y��6��A�I�vPW�c~����ӁE�`?UN��-�$��xK��8G���mY�dC�����X��i��-~�pL��!����Tp�6ܔ��V���zDt�ԦT���զ[�p���F�6v}x�l�<�]%� �4P���٨>|^����	@6�|O�˃t��I�g�U�AH.�N5�7�"���XG���bbBU0�9E
� �d����ED��E��'�L���l�H�Z�>�L�h"�O"�S6/?��	�5�>+j-�+/�Xl�8��aʝ��d�����
�oTTF���WCDԶ���0���MKq��L�N΀DԲ�<'Ŝ�����u�����@3�9�OW-�$j�"Xa��7]��Az9ȁ�F@^�y��}�Z[jg�P�1ܓ	�)� ;h���q��3
�3 ����w��b�П��l	�e;1[��~�%@��v�bfW�W�P��`�U/�y���1z�HgH7q�pv�@r\��fWm/�A�j>�"�ҷ4�>� |b<%QLg!����y��G �F�|G�[ϕ�Ȑ�����cS�S��]�I��=���B=����S}�uo6����&���?����:_a��T9����,=@��kw4jHe$ͤ�P���I��GVベ�o�/[�������e�'޴�U�0ȣ��Tm ���ㄺWu�i	R\�:�%[I]`�����-�T|2�X�2���j*�&-pD���Qh[e���8+B~�a������[����a���B|�I���T��3�n ���ف���B�q90_�0�jmeG��Vp���CAJ���ٴ�a_QM8��CA��F�4U<��9ALԗF�s:pt�Ɔ�@4#��X�r݄��!"O�J���6���Υ�N���CQ�3	�������߻��!�[�W�`5�vA����X0�K�Ci�cI	0� ��A���ǅ~|>�σ������᫂ר��n6�u�ȶ��m��b��]�XN�c�tLk琑��3F
�k?���E���z5�m\�{-�����&�4�,��|0���Y���0�LO�4�Urqx�VځJ@j�+�WU�I�2-�W̭j�g#F-N�W׫�ܕ�I�T6w��mb������jR�4\B�������"��J�^�6��t����9��4iPi" �vXr
R�6�3�A�é#�=`:hja������2u�D6c���" ƘM4+���4��N��ER�O�agP�>���u���6t��o�G�<Vr�]�H�^|��iN��Kz
��=o��n�qn�>�b�T�be��k�Z�:��A���6����W������ � �!��o�`߿�d��i�q����$�2��5�x:�Bұ�����1��Z��YB��Ȋ�� 4��G�f@�il�4|ފZ<#���t$E�3�:�"]���[,��P��7j]m��� ͞a�G8L��H�31q�B��Y�F�������d�V$��Ę��ԌV��;��bmJi�_#��>$P�R�Za�a;�	�)��/�4Ts��ޡ��j���Crݲ���_-9#�ێ**@�!�L��mu�|	C�IԌ��=���F��{�٬��iBq�hٻ]�f&��:�^�N�N렽�A|���l�"���h���(�Y�F ؟�5��F�}bkO���Lֹ��J�5�e�j�&�W��yAzP/K逿H�]����Y,|����h8iB\�%��k�|�%��0Z�0��.V��T&�'zi�L��l���U(��,9��0��	i��'��'Ku�8��m��F��3`F�Ym�q�efd枽��6��:�w�y�K{K̍JAj.
�6b�J���`nE�9IIx&h�< A;ll�U"�'	�|�S��/����.5�yP�ԇ�"cm�W�T�̃�A�d~,"]h���;nR��?k)
�"�ݧ	��ҷ���诱_��߾ʐE}٩�uh����"z~Aeđ�^=Ÿ�z�H�(T��
q�Me{��]�?N
Jt��2�]�OC�ƕ���R���i��*���A'�?\�#��,ѩR�n��d��3(���r�L��������ŋ�܎��D���4��P����C���͡���&�*��S0��歨��1
��.�1�t	�y�u�÷���ɏņ'd��o˧���N�í+���v-ݟ�ݯ�u�:=��IÓ�c0��"��Z^4V�x����H�P�$�Q4�����h�19{�h4v<g^���9X;��:���CN��ٟ{��NK��ń���ȽBI�R����y':�4���IǪ��3�W�ٝ{���ۤ���6-6���U~T�����s:���a�Z��T=���F@or���0x��,�~�d�*/IUv�+�+�,a����%�77Ϸ��Ai�-B�:��>���ܢC1�<��`�iYUg]����aWC'yr� �g�K��T�L�6�I����/�czў|��z�\x"�B/u�W�Qn�K�d�Pb��&��+���3�x������s�� �������u����''y��]̰���j�W{�e�_���������~�6����������*�h��K*�L����)	�d��
YSJĪ�'�d/>�"�����ǫ�td�ŇB�܄���V����f�n^=)4�Xz��Q��	D5{0�Dq;��!H��7k�pJ�g@�DNS���@�d��'��*�&A�n�>��AHq���0�� ��H��C-+L����ZB8�&��������9�w�㟕ȅ ��s�p��e��)x��[C7Qe˹�3j��Ă���{�7zx���U͟��Mez����w-!�@� �v yS��+��	R���6؂+��k����A���Z��f7B��?a��h,U�쿅�(��F�b�v~���Vv��2�Q{΄=�M�#��j�0H���#���炊�3$��_B�:��^h�ć���d�i�^�q`
��Կ7�/�1���A����F8U�#]U�ۜ�կ�6���6�)tN1�{�p�εP������q	���'���X����A�Y��~zrKw�Z_�n�
Nn��H�T"�-km�p�y
pt=Ɖ��'�k����^y��B4:�	��� k	ȟ-�y,��_�a9+�1[�\�4 w�`�J���N�pEҐp� ���.��<��$�
}�8$� ����8ʣ "��� �N�Э+.����)(�]-����@�rI�Xp=�F``J��$�}3�&��� �n�Y��o�y��f��`�a���G��@�6��!�|�`b�#l��P	�3�=�����[�p��kC�A�H�)��,���]~ ���}*Cá�{�C��ԍ���2@Gj���՛�4�oY��le9D���n���	ו���,$AU*:�lV<��a|������:�S�:����R�`KOZ :@�;2���0g<3�e��TCO �$�5E;HF��FDsvp#^�@B}P��yA%5�o M���И6`����>�kV�v�]�̌qci@�U�q�sR)��At��%��Q��~0t�ֵ~-��*,C��|�+"a�B6Ȋ������;�N�.�l׊�b���jى�EU'�#�9p���htk�P�Gps"�~���Ơs<?�@�wUi�.-����Q\�Y��a�k}�5O��wwM˯y���h��^q-j">��Ar~�A:�E�q����ےF���O�s�Z]z&�+�$�\b� ��Q���&ѣ _~����{�[6�3Y`r���zk�!�5�c��,�Q�`�Q!��8�ȐN]B����g�M��vT�o����l�Nig����`rDT�IfD&�>{�v��¢%��$LH&�Ȑ �I ����!�Ƹә�X�?9ƈ5h�X��8�)Oi19��7	�Pdb[Ք/���H����Z�^R���� ���5��}�y 0�p�־�s�}���v�w}8_^�&�
�Z9��
��&�uF�I�������c g�Z�U�^��@}��`�{��ep�c`0:��3��8���a"��-ѥ��w�Q��ӵs7\�b��a �nT�L���*��Go�l�	|1����c�O�K��cJX$�%-��Nm^�_��P-�8h�#΀��h�h�aǐ�_U��w��1wO�Uݐ�V�Ł���*t``TMA��h��#Ł�Ł����X_��G  �,��Qu��tH%T2�><+E�*�-���^`� �̀y����{q���|��@�`?��t-�]�8�h�:�8O=�1�x\y�zJ!�� �mX�|;�+h���R�����|y��7ѧj��r,�$��b���A��>�S�#5\��}�#k@�q���$>�K�p��3`�M�f㬆G����3��K����虛��$��330����&��E"T�+���"xY4�*/�-����m�R���/��{+�������r�S�c�v2��ld����}~�s������ϒxl�6�f/��&b��ph����l���%�z��\05��a��"���mݛw����sԚ�A�bg�u=J���g�Pxxs�s���y�k��2~��0��D��&3'�\�ODl�� �j8';�\9�,����*4>�]����JX�o���+�z8��{ ��V���d|	n�d��u)�z���-q��5�?W`=3<�(����N� �����a���������L��7Yۻ|����[��	��V�mc>��U�����Nn�eFb�?��O4q�U��G����֊WV+"+�f��2�r�h ڄ�>��ni��_tx�ڼN�o>>&�pБ�<�����x�OB��{�5�о��ltV�~Ǚ���W��sB���𚬑A"}AN�#e��si�sO[��N΂a ]�E����}�3nQ<��B�Lbb?�e�й��i[��,�%�JD�oI�5f�6��y�[P	(��������j�Vܪ{Y~*;פ�ސ0ۮ�e�w�{�m΢(c����p�s�b����AK]�/���^`�rg0��KV�m�7��v�V.�UvS��T����rg�2��n�=�w7ex3>Uj��p*�OeG��T����/u��ԩ��j�Ge�� ����\��<���A3�un��[Z�i� �^����|]�i��p%�%��� X���2��s�9զ��Scy����<�ыQ�iR���($Kf�eilfM4#���#ߩ���2Z]�̴�.��Zj�L�s)��R��SM����%T�>�wg��q�V���{ȴ{C�>#.X95~���[�vvA���_w?)����<�D �H˰�����ag>:VD������9e<�s���HVR��'�'<n5R7�B6�07�{��9��mt+���h����3�|Q�Ef.)P�'9#m���Mθt;I��M�2^�8���O-�N:�˽�:�z;s2Ը��oZz�w��Al��#��D:����^��	��5��h��d�*�#���&W+ǠĢ_f���p2v�6�p�	�Q5gV"�p�1���w5M�5b� v[1�ô�Lp�f�#?OV������>UyL#,����_\"z�K����b~�'G����F/�V��\_|j�?��V�T3o"�Om
�n��el�GsN:[�M4p�G����AI�%�
w��҇�S���<�1H1}�g�Ն���ʵ��}�kg���j���[�ao|u����&������L��G�+�V�U�l�Q9���mn������$���}���A�b�w�`��(pg-�
���R��b�n*�1B���Ӑ~;;n�xٛ��)eQ
z����,�� �c���Y`�e~���,%6������ (m�E�F�=��~=�<��J��sw���;;�j�@��!^C�"X�a��P+=��*q ���V�c���xE��ғ�1w[Yyc��q/W���Yx{6�����a��ʈ��6�K!�6"n�6�pZ�JjM�J>��Н%b;��Iq��#n���!7*���J�e�; Z}9��N�=6u˶���IW4�Ipc弁<V��QJ��ް��1+_��{c��H����Q��P�`���j�� ᱋��`T6�IP�A�u�S���~`�5��7or�T��4GP�*x�5~ɵ�����(o}�K�3-r�{Є>��x�����"J���h�ƘD����eA�t26V�"Ih~�H�����\:�
��5�a"������К���'@(�(�������r�;X��k��N�uα�9��?
�x�R��ؽS�<�H�]�����e�ڥ����5�Q��� �AK�}���.I^�)ցA�-��h�Q:`�\�n�r��Xu=lH�&�Z�3O래��kV�g\���+��b�;Dh[Y�Gx����/��T�6��Gv+nBn�͵�kfzi�K��M��O�l�T�?<^PtD����_4��w��M�\|Qi,�X<��ñ�6qd�N:�|7N!|�;�?��ٌ TKm�\�+.��G�/CM�S��x��'ӷ>���&����#�I�Z��)�)781��(Y��C;H�~r�q�j�PT!�5�L|L�nvS�C+N͹L,�a��M�3��e��r�g�ӏ�����2Gy��n���M)�����/ADnz�A����v״&M������!�г�i��b��pϔԚ�d���_ȳ�.�	$��Q���1d�Eeeok�n�x�L_���5���jH>�����@��^�.'i2�rD'��UT��a�
j��2]a��36�DL��wY);����dB�$4TT"�9��0�$����z�1YOmĽ����JB@ə2��߸[���k��C���.�"d1n��� ��sM;zaqu'�k�Ҕ_u5��32�`��26�B$hUi7�(� y��.�:�z�.�N�:�l#�ζ��De����Bse\�N�»?���%t�Ɩ��G'���&��G��Fpp��@WO^[bz��L�-o�O����F�\��*��P�͒������Fd�zbz>�l�� vq|鞊��~ٲm�8Gr�aaP�i0�%OE�$�e�	���� R	F�׀x�Z)yg��2�t�޻Y:�@�%�k%x��2J�u����qU���Q�fv(�㹫.m���M�r�p��u\��UGgV?<ם�]��f(���&u�[��>�Xy@E��N�;��%}sdJ�fy����!�*�������P��Ɣ�����_���?�z��k��;=��=��s���l���F�8��p/��9>ϩ<�Ւ���{1~T����^��7�@��,�p��K�j@�i��|��Q��Ԋ�dm��ƚ��1R���j����_��?O��b��_��Sq}z��� ߨ�ŝuf�3x�7��>K����ܴDZց����dz����(l��Ǐ��pz�~Wp�ɜt��6��b��yY4*z�*C��6ǆ���k[�)���� 	�Վ���
3�3��Ŋ�4�NJ��pn��+i�cɣ3�T��#�K��ƥ�	�w|��E~�X�g����l�N>����=�<��Kg�вh`�6)d�´3���d�ǵL u,C��1rL��^�<�_�q���������C� ؁^R�C���x��s}O�Y�=	�+U���>�MY~x��ʂ
k�� ����ꡋ��>�*Bo�ӣ�|��!��?����#�k+�(N�=�<�]ْ��u�`�����_�]��xs�x��¼���ƙb�Π��< � '.5=fN��44o��"���Smex�<�s���ho� �A�l�/�pA�*�����s���2�5�S&��)�
�����!w�	Z�2y��Ŗ��{R���K�A����[��o�W��W��v�������{_w��ϡ4�XI���W ����RL�b���I�=B�bGk�� �v�`��2l��8�h��?!�Gڟ������]�az�H�G*`4��~�7B��6����j�m�H����Ӿ���o�)�[��@?↔��7_*�yY�i�F{&$�?�sƋ���:F��/�����M�H_!�aL��yvN\] ���B�S_��V��Sj�Օ��,MF������Ϧ�n����_"�da����j&&��Y���wt��o�)�ж�p��
��3�Qd7��.g$QA�����^�r0}��U��M���u +��Y(���N<Ĺ��$%�LMt_���g�<ם��q��ha"���h���W'Q�MX��Qv��h�"[B���s!bT�4iy�^��E���9�%gq�N��ɸ��F�#c�U�a�?����DBl���f�8y�����S$;�E��ߋ�{��/�k�H:�s�Z�|��^�߾��V����h#'���x��\�ap���S�Tۃ���1�C��>�]ǊV$c���v~��-�W�&�4J���4�N����=6w�>-��&DcO�&?[����P�8;	T���I�R�OX<%�wr=��R{�����Z9������h���xq'�d��MU����66j��|����#����b�r6�a6�TM]S�l��m����3������p��w�8��+>���F*���B��э�6��KQ����P٠��X�W�=���w�l�7���:p�������-�o�1>~C湑��O�����!�j� *cd�A��2��$��%�������o�����x���9���K��yh��3��)<���4�l���ď��{�eۄ��%�A�RE�Ε��s��(*xp;�:�*�J�,~�uk�6ZYfM%��T��ßRrypD�pҼ�!*%����������xhΏ�B_�����S�W���[H�{�|����dEQ)��?xUA�`j��љr�	�GS㭰"�L>����h�
C���1�˞|As��_>����f[�:�S�.�V	*�z�"9:nT�P�_%+E��D�q<M4O�n�QΣ�ON����*4Pg#�g�p3��ao��r:����KUf�!�уA����A-7�Ql��^�
���df�µ�u������T��:�@��«
��*�0��«���Q:Q}�� Y�/FcуƨTH������(��ADM�x7��V������W�F��_�W:X��Z�i�
Q *�C}�KH]`\���d�&��W巏�.��_��˚�!��&,��tc�Cf;�<��f>O;e��>����~Dp���~[0���A4�
R	�`R�R��I(R�ccR�`���q�R�����Q��A��������R�Ɩ=,����xWP��<DR�JX*9�V��A��<d����u~r{���c��!�g�~ȰJ*�>�.���0L��<w/-��x������?�x���f�.rA�� ��"�ǚ}�I��h�&�����~��q��L�� a�gl��]���x��WxpEG��ʹ���0����C� �@�H��jA��F�{�#FH����H��u���p7�nbR���?j���l��9Ql�=]��O;�Kf�� l����	��
���v�)�,T�7��[����N� gf���&DUe\q�W;9N�e�}�_��\fYc%⫭�w�{�F{�̫_u��-���F�s��w-��LT�X=I�#��_i!��H�RV	��Q�>U��M:2O����I'��{T������l״�Џ�қ���|�R-�RI��
�UU``
��5q��M��1裀Q�O� V�phwf��5�uJ,�0O�偀�B��[<ºm$`���I]�L80s�ym���S8I���:���a�,⾇k;��oK���l����uo�̦�&�z6�����&�[w�@A2R8[�xQh��4��3Y_~Ή@g���Svڮ�`��H���Q����}�ȧ���0�3��U�k
��v��@����d��>ǽ��rz]�3�W��!�����}L�dfI[� �h'ήM�	�"�aA�ZNи0��;�U1���a{)UByzͱ�`�_�vع(*4q��
G��������"�S�C��\�m,��<W#R�7^:�}���9�������U/z��c`��+���QK"�د�*1}l%�*����+�`
�`)��!�{��v
�K��8��xS3����+/(Xh�xz�V�ZJ
f������M�U��~&6��4����I\�	
��O��Mg
�=�� ��<8)c�� ����}3Ĭ��E6��;>b�e���e\���it;[,O=�Wv?}�o�+��{��g��cF�t/�Z)���k<�<3��E=��?���G&���8r��p2Kx����*&�a��`�C�I���YR�ƛ�:l^���ӓFEK�%Ѿؖ��>��HL�3�����=�J��>�Q���-_N�h�dW"靀�rq�&% OAf���aHo9!/�'k�慂qn85D^\U��ė��`�#�?�l'Φ�I�e�úM[�	����YdnGS�ŷ\Ih����:�/Η�����u�re@��7ˣ�;�6���Ӳh!M9��S�O��$��8y	��b�kx��kǜ�F�!"W1��C���1����VA p��kN������ė�:���'���V��Ͽw��Ž���,�X�XJp����f�z<��\p�B�p�tb�%y��;H2�C�g7�����7����Wp�ل�fOE8'KBfJq-���O��t��"��Ӿ9I#@�la��Y%�����f���1����������^��5� ]X�%fe����X�9x���a��3�����̈�/�#|+�kj������@�w��=μv*�9�y��h|N���x�d�K���̲��>+x<Ô����i�.����qO�����Y�>�޲[�D2J������{/�c��d�u�d&1o8"/�X�`s�"�I+I�ց�BJ[�:�g��wJF ����i+P�E�R��x�[t$Ŝ3��}ίi98�`����&�U"Γ���8���27���%������
v'��ͦH��>m+ �����/�ZZ⎷�ʷ��^?�,\� �Yu(kE���<傺�D%(���C::�M�!蜎,k}*g��R���%oW�Z-J�����&Ķ"pN�0�?��KB"[]��jD�	��'R2 ��!���e>���O�4@f�x~C����+~|8�ׯ�J�������:�z��~`�j��
��e���A⩯��
ڦ$����t��K@�S���'x���]�K`�3<��Kzᠷ�wI�s)�Fd��Sj��n�p'.kIڦ)#��x�ʜF��d�����CcJ���T*�W�sF���Y<q=M��BmD�.ub��j��Mgs.�R�0Hx�%/Ax���<\�0x�t�����cp��"0A7�r8$8���	�����ДP2}�*7�z�HUA�B�ܫv.*��5@� ��.�v��@��[v������Q�C�]<�&���P�$;��J�Qٰ�BP�DP ���ޡ�N�a���H-fӷ�e)�������y�Op�ٍ;4�sݵ����uR��ذ͑���b�ŽC��l������-����a� &�+�:�)��f��ލ�3=M�t�O{~R��0�k�)kB���{x���$i_Z!p܏��'&�Q�H��A�m�ε�&�G	u<��h)oQ�*��(�À/�O��0gs������g�r��_�R���Ⱥ��j��	�g����Ho�ڪ4�g�`��TChr-��U#l9��{�=kq$.p#/���E�Yΐ�%���h3@���Y�c��1Y�k��߰�e��?��V�y�3U���QSg�J�?��gT\�`V�$�ad#N�6(�ޅ��w@�1wR���$���)�U^Y5��n��(�F+h���@ˬ6&l䃖�����f�⣁��a��H�~�|��@��µd�Z�YEI��꣙��O��\��vl��:7���:0��t�ɱB�!-��ϕ�84��r@+aIA�岶jd�f.�D����`��7ױ����n����L�G��E�>u+`�`�qB��po��WD �\NK1J"���M���C�
���i>IK���>�v������T�������^�C��M��6٧r��㌢�
��I��8��z'�3�o���U��{����Z��旋���`�[k|-���+�J����'�^M�
`S$ �9��zk�$e���P��5]$�;ׇ dPq�6R���UQ*�]��s��lU`T��eP
����K�1�-�[	]�C��*&uʳ�U�w�����6����X&�N0�g����~�]���^��|��,;�e8vؗ�K;d�������6�d�h��qdفŇy����H[�M��Gv��o�4�DR�I��]�`f�NWj�˰������k����n޿��]�s����%ʋ�����bKb}�~�F+�%�H��s� ����!t��G{��/��A���n1;�f�b�uy�q�^y��������1m�r�1 �hJ����u_��&�f���s������8$W���z2�G�����5hTX�
�勞�r�O'�P39�(xL�;!�o	>��+8�����\��$[�yNr��59iv2)Vm��pB(�҈��/�����'�:Y�aW�	���b��F�IX�L@48�C��>��n����Y�"�:!z�`��GR ��� ����H�2uj�	���	�/Cgl�4��!����ԗ��{����Q���%c��1���'��]�,������^/9a�1�S ��3�/̊.�Y��P��ަB0o�O�󭫡&��*ý87^Qd	?c������m/[mF��?�0�i��%S��8~T�M��<�f�מ�K�S"�䊔),�뽆5I-��҄{a���f��r�x�Ҩ�+9�(��-ɾ5Q����Ʃ��6Y���U�P�8�Ժa���A\g�}�WTISh�n���v@U���˘7� �z{����/uv�ϕ�2uon�qh2-�-a���UY�/ 	���Tċ���Q��LL�нb�IX�v���S��H���ӳ�FF��U"A��Y%����h�7�.4�opP��*q��4�]l�R����+���+�nF�3�<19�4�@��m�:tp�������r����f�n�����yW	*��������b�Xw��\�fQb���S\�gm�l`��Wc>
���lj�~`��\�ZC�W\��!e��ɿ��N!p/�z�W�����\�fą�V�^��n�}�J��`.�,��l��՜=s�d\��u��<!1��� ����{@J�+�"�x�Ɍ��%���~|йJ�ۻ����>8ߠR��Pd��gWB�F�D�>��uĀ�ث��� �Y<J /ί��i����/9���Χ�h @]Ҥ��_L����Ä�l����g�6�}�GH ���T��A(�FX��k���@�O�t?3���{_7����g�ނ�k�܋��+BI~�N¼���l�e�r|U@��J��p/V�o��ec/�����i�>M)\7*5��=��L.'����d��PU���y!)@`t;�i�����u���R@���O�Qt&Ɯ�^�x��:oF"�
�}��ӯ�5�W�le�K�n�����B�at'�'0KA���{h��n����.{	6k�@���%֓�C�E?[��1d-����0o1��oE�H� ��Ta͠8��Ik�o�e�1Ip��Uh��nvp�]z�4/���j�<u�õ2_W��bl/ѡt�[�2��g][i�r��W���Ub����>�ǽ�[OP�h<�UMP	P��eB�;�"�ML+����S���<�YA�x���X�?�>���HZ��Ui	4�& ��)p^��'�N����/��x0�Xp��j]!��Eh��G�Z�8A�4��Ñ���/���E4�Ǫ���cA��e�Ќ.��ڍ�K*/.��8Gq���&'����FW^�gu���-�=T�ɉ@)@d���T*!f0o��BtZ˥_������X�W&0U�K�c!g��Z��@��$|w�O��Q��r���''���	���a����;��K,��{�Fw�h�GywMc,
�y�bJ�(���$�;J�Ѣ�&������O��3����o v�R
�u�c������5�g�ݓ���Ap�}]R<KJ�^l]7�G,w���2�r�z4�e�{%p�%��fD�����7�}Ra�8�����?��Sw2F�����} �J����+����Y n^�R~XVm��y��u�8�d�Ej�s7�fu��0�r	��o�92V��'4C�:H H�=݂x��7>��h�i�d��{�Ы�����=G�j����~?���&�}�|#ҹB�����N:�avD���5
~�{���k<��~e��?l����s〓A���'�3��Ir4q%�R��%c��Y_��'p�hS��;2���>R�Z�t��G6aD��E�4��:�k�#��2�P%�6aD��%�)V�-�ClZ��6��θ�Q�)�[S*�h>0tX����j'�$8�0�ʦ�$��沘��j������bi�j`3!5R�*�
d��@~(��ƨ�h�|�����<���[��pO{�Ay�`_��+�n$�����	X�8��^�F�=O�i	4�
&3=ذ���=�'�"�g=I�;�PK�e^pGz:h!}9^�h�ЉX?�.�w�?Cq�N��S�@�!��d����$���`�S��2��x
,�,H����^g09%�l�~	$�EJ���l^ē/\�'a��`':Vy��8��1�O��M��<5� �*��n>'����h�kiҔ��>i51�/0*F�$�)�����.���	y&�t�<\���r�P�hr�n�أf��H	Μ����]�#�����ߘ�'oߔ�J�WCd�L�p����S��}rN�W����b}.K�ʴ����#��A4��L|��ԌQ�4���<�;Z���R������4�o�d���k����S)����-j���2`F�!��^�f�r���h�j�@��+�ލ%����� t�"fn�"	l�nÍ�Z���L���7F�?G��J[���ʒ]�6zYI��Yv�*�x_�N�]XB@%���KC�$���ԔA�kI���Q��B�
��W�k���le*�OH��ҬNQ�CG_у~��\�	�h2lU����������}�U1%E7�<V��G4�|���x�]�(��E�Qs�{C!1���l%���I��#�+MD��lFUX�!����R��QQ�"<%L��La7M>���_��Q�u��T�1�3����{c_�i�P3��j_o9� xT��[e�|Ϲ*�ƚ�b�rE�Nd��,�����w���	�'Z�qué���������D	T>�=�{���T�Er��X8D�����Yf���kN�;�'�j8?��81��<���a�hة��i�� IZg�K�М|�E��:l����H@�N@.k��"���/��0tIv,�+ �m娂A����T̡�qu��y� �������*>3z�%��On���nA��v���J_�'p.��1����#�΁H<�u�p�������`���K�鮵���e�	eJK�[�����1�$!��XA)�eb�}x���=��V�L��'n^Dҋ������?����wu0g�hbՔ�!G�3�G�awX=ar�|H�Ζ�lk����i�ƁB�}��jf���I^���~�f�K<�2��-T�aK,>"���5H��4�*���CE!uI�$��w�,��2���� ��)�����H�*?��Hu��LHJW_�:�D�ɻ����]q+v���,���c��m��uv��y�bS���Ҟ _c>�w�S��D�MΙQH�d��.7i��N��l�ҙK��E�Ce�s��v�s`�xk[�����s���b��e^�W�Z�DJ�rڶp�2�7	(O���-cw��k$�@�]��D��i�]s�R����2�T�L��A	)a{�R��؞*�)\���^y\�17� QIفL��;"WG�r��z	Z1X��F���`c��T��2n�"������>R}gC\��-�]����5��̜l��*'K�I^�A񁀊W�{�pi!Wyk^���qh��nT�u��,����\�E�7���m�_�>#Q"R\���<XHQ���7&��{�?���Շ��cȝ�9�[���		��w ����X�;M����w�,������W�`қM���H����۶����#�9+/7e�A$��O�o��u�s�:�Ð���m�3[����#��k�X�\2����2r�զ�Y|�n#�:��pQn=���4@Fz�ɾ�5 p);cȵ����}��J�~)��ڴ(�a�U���uЍi��ĐC"�Y�i������rلH4�jQ��)b�9^V
5M�<2L�=�t����ֿ�8,"�6;�)�n!}R���ޝ����.㩲:��! �|
��PɸRJ�s�T���}�N�@+�#RϹ��)viM�/�!_������N��@��'��'���4���1���%rxv�6	y�]xH�픀;E�q����6�M�S�̚�@^y��镎~�*S��9t{vmy��%���N�U#�~>:�q��Ƣހ�#�W�j	��K��;�e�%�7�la�=���F�C
�V13��&9yY��B��5��R_�=)�4�Rzi	U	64� ʔ�]\S������5�-#%l(�neچ���g��\k�u���q8�h!�	:n�^�~YX�o4~	�q���P,	��΁�)?��x��?sȉ�Q�p��2�����hi3�ڔ���{���:�]�8_��ʩ﨩32)��;��tKn�������ik.�A12R��H���hㅓ#t|�y�	�l�s�Sl���.�_j[8��������!g��ٸ;�Ě�hM{�`I'���jj��7ӂ�6�y�oNm[�i!�� f�:!�W�ӋZ�,~�RS��R�G��)���\�j��S��鸹��4��N!/�A�ٝ�F_��V�'7�*�Ҿ��Т9L�e���^
�:ɝU���q������|d&�Rw���B�A7H�c&�Q'z$2r����<��$����5ۙ�7�%c��N3s\��ن����£�o?q��`�}lKi��m"�CzfY.�4�K��6��د:����p����ӎ�ԭ�*Ļ��ϭPؖ��Ȟg��@�x�u]�,70&�_�s��qG�|u�|����boW8���>���K���RNP���3�'�z�*��$�_��xc�=�aُL�z3�Ɲ�EF:���t�sװM�SJ��*��f+� J��1����ę��d�ì�����̀0���}B��d�l����*rK�g��-؉h���2T#R�2��� �Cp߾P8ea4�Ӆ)�G�{ތ
dgՌƹ(d���yaV=ǚ�끑�ےAVPa��i9S0'HJ�t\�s88��ݶ}X�QW�2͡=%��%燼/o��x�Qx�?�o��cu���)z��c���F���8V>��������r/��{RqϹ�-���9��
],�C�y��@WI���i4��'���0~�!��<8�E�l��Jw%�Rʭ2���%����@�30m"��C��ʉ%�]�B�-6;��{�R��dE_F()oA6k�L4��I~�5c����Y�OOr�ʛ?!`�0��s�r�L���%��l5�� W�
����%�M�~A],��3�55�4�<��CR��*�'4�����c�=o���tG�h��7��@m2�])�[��2Ad��/-G˵�K�H�n ���b��	1�#��^\.(�������7����[�\�1�k, �OJ#��*��u9i:�6�8ꖥi;�"�\�/w��v�>�����2x}�P��i��n��B�]��Nu���fwE}y��!Y��d�FpsDS����>p�Qx��B�Z�|�D�H���R����_/��p(�v�44
^$��޶���^��3 �g��9i?6��Je�8�aN��Zpgn1�쁶�"�R��� �D��?����,W6���iMHFH9�� �jC�u�d�-
������BX�Z���̫3��6��)�XSgN
)��d'[�C�s��EP�H��@����>���p�95ԁ�U�j��@�$yI�xb��x��K��ŧY9%��-�v}i�����Kbq�X�!�]�[��XF�!~���9�(��/M�KB9f�o#~lO��ӐΙ����K���D?��U���F�#:ys����[�Ç��E����y�p���&�*l�X#Q�#Xp�,����o'*���&�`0Z̎�9}8�M�	Ȇ�����Sl�Cq#�J��r��S+'����D�H;��4A�n78c:m�-u����3@��,6г�x�*T��eD����j������;�yݻ+����,띕T�����X��@-���7:�_9�~��|�9}�&޺!� 6����_��hG!1����T�	���l˭����?EK�m�s��"��D��`0��=eS��u�x���<��j�ҠJ�r��to�;XFF#���MR���`s�[�䥤wݧ����"ٻ�����«��DWb�#Y��D?.��].�]�b�uC;�꾹��}�+'�y�h�qc���G��5u�1WD�)�W�B�515��L�p�4�M��\����	����<Sc��2A$0�5>0r�A���M2HT�`<o{d�a��ܷa���0��%�/�~��\8x=�a�\��E{-ƛ���t� a����˼�K�Q.�D;����;��,�����>�N�a0�����9-r�����bщy���i��C)��@���^��Nl#1��ni���,���9Wr��J{�i��t	ˤ �w�F���ū}�6�''��Q�3{���)�� �T�[D�����M�B��B�C�]j�}?��e��@e����-���p�jۙ���|e��c��;�?Jɓ���4����D�L�ن�t}c"�4��,��˥� K���LL\b�-����b�jȨ���wp�R��-n�}psN+��r�}��L溯]���x�'�5ZY�ۼ}��ZoƬ��SЍj����ڀyS�ͅ��GN�g2�nC���~����-����q���b��k��ن�ͨ��-��s+n0'�L�wt�V�=���/�wa�__$�]��tw�R��U��IXL@|�4�GR�w~�v{���3��KS�l����#*cy�jt��`{�F��qs!���{g��:��P�ɐ*PF:���hTB��dP~#!����8[6�bkx�'Zmէe���ɘFa|Z=��m7cp�nN�l̃²���Y���&A��&���d�X+|k>��\=7��r��Y�Mzv�{�M�1��r�'O�I��_��BY�C<�"���B�R��T6�C�T*T0T8�4�^�\:��˄iz@y
���[A�`.�$7v@�|dB�V@���wK0��r���଎x����\���o�a(��z_���4$!ܥ�/7�:�ֹb���c[u3;�Ѹ5ӧ�!~��A�\��s�܁��0"���gk�-���%}�%UF��QU	i�(� *"���h�G�v�R~��̛�7�&}v^���	hZC�P=ZYg�@Z��� ��̍ο��3�=�а5���;A��]��>�Ƥ-�+�K$' �V�� 9�G��p�6�mW$ȳ�8!m�ꥻQ�q������x�`e\�ԁ �E�qm�-�������2��	]���%b.�I�}4�h�6ʉƏ�%����2m�^�E�޿���D������h� k�$�z��	���=e�n�¾�G�Ԡ^/T��n�!���|
'�tɯ�,w!	e�4�wD�l�wM����&��#eč�޷|���cиg�i�I<�+�ʩWر[͋Ľ ������Loip����>�e�.[J���F� 7߹��J�-��XZ�9ъ2��<gJ�׌:B&��GE��v�<*��B��H�i<	YZ]���,�Xe��F/u�b�!u4���?��9�C#�̺��4�{o�I�W, ���!M3[hz)5���H��o�|��A��K��
7�rgԵ	�V��h�?���@W4Ӥٸ�{����E����Li�q��CI�:&:Ϙ������Aƕ�m��ɚ����;ɛ��� �`��)�m��G<�3Q�D���V�$�p��mh{	�������L>r3�~���p���o��L�~��h�(�W!�hH�y�@�����3�_��Ի����W:ݾy�ǙU�R�%�p��wa:�z�lE�J��W�򆇜[���α�K&]�a����@F[�&��f`��^"�@�!�����u$@�ћѧ�M���<�S�oM#T��rjyː�H��**#���8$�᥇�<2_ �4Q_�]�`��c:�~�����
�*c�����%}�F).�C,��@�&���[��b�uʾ1)K-A*HRAA�c�����'9)h�Uߢ1���Uߵ���Ԏ�On���.}���˒5�����H�wh�q�v��J���2.�(����������H�0[��S7_���ĳqnQlK����	pC��B���׎���3:-0.�]��'�o/?���o���-[��k���U����`ݻo6���_�����ʣ4z�Ay�
�����MM$��<�~�ٻ������n����Δ��L�jDN���_���J�K��cw�8ș+GĚ{�`/��1M��F�^�TL��#w+.�p��WwL�%5d�T�^��۫�l��a��2YG�h���#���D�O-+�!�w(i���\��+%����1���j���4_1����LBg�dmB
��"�����V��]�c��S�)s/T�^8E��p�.N��R�a�~5%H}0�QrZ��}6R�vA�6(��G�)(~�y�Y$ >��D}K�v���[~XM`'��7vsU�|+}����BT����!�y##�����d�3�=<��bz����H��N���2=y)����%,�z�*t�c_�p��6I��1gI��h��i�(�ڡ��f>�X���.�^h��m��d��w&�iI?nc��*Z���k=}�LD`�]��^���|��9�)T­��9��&A�
��q���e�š�3Ԙ�hf��Cq}�׀�pU��㡹m{���NQ\��%rj?�+7�N�j65��]��[S]��(���C�?O���3����;��f�]�2��1|ll����D��7�D���6�јq�	�B�(я�A��(};�+Fǘ��_��۷���@ځ���'�����Ī�!G͒�b��Х>m*���ʸ�l�;���
uk��]���Rj$`<��ӆ˃���A�=��/3�
rČ7���һG��D;��%�W�\]���}��l!�?vl�U�e%�m�Y���t)��������ڵ�?�[�X+��h���HQ�y�+}�Ύ�:�z^`0�C�=(gW��pl�/��G�$fӞN<��S"\<���;�Q�e �;Wh�44"��ɞ:��=[+��O��]I����Qq����f�ۮ�ű���Q.�ѹE�$�Q������%��!�)1�T�'�%×#��+�K�AY�0ˬp�C��?^0s�����~���k�^[��f8s։}C/Gb'^~MCN#�u�E���P嵄E�b���^�[��!%�KO�$�Ö���+��O��k��^R9��ԌV�nS��6��\Aת� �p�A���u�z�ys�xӍb�O��t!j�[��	?v"Ȋ�l&U�[s���O݈qY��؁���9�˃��|���K��z�B�Y�&��m�׺��9c璆J4 ���<76\��	$��Y��Ӏ�D|�G��J�_Ms»W�uU*��F�9��	d����m�c��"�"���p5�}���]��� ȫ��8��D_�3�d�)ӈ����T�L�XL��.ܷ�D�2��]@d2�yj�F��-�D�d�t�'����Bf}����c���N���j�߼t [�Z;sE���4�uhYl�����lY6�^Z�����������g�G��r�~Mt�!l���W�Xz�ʱ}��>-L},tʚ���C}w_�V�@����:B%#�����H:�w����͢Ej*�%j�a|N������+�+�ɕT��Z��5��If����˪���=����4�a[�6�袴��$3L��3ZJTo_ݾl�ff�D�U�xs[MҷmG��!s���o�Β3*xx������a��j����J�b�#R5�y����T��k2!�-��_I����=̲]�~��-�٠gu0����=p�V�6��2�Tm�
�tҍQ1!Ҍ�P���[y�������6����f�r_-�:3��N<���0�h�/]<}���u����fgn���0Z�uK�Ǝ�e���|��䱌>ˤ_���Y�����x����Ґ��3J~���(�	.�`�ɪ�E�^��Fw7��\�����M��8򫿀kF_i�S�z��|�<N"�P.:�s���\����-��|g`1G�4�T���G�Ɖr���*� ��a��"�z��w�������4��'��=��%L�g7W[k}+�\Q��-&�ƚ� K���.c���8��	��T�n7��d?��2�.��	�J^=�\��9&nꔻ�5����+�z&�������`!�ZlKt+���L���C[$��S�p�x^���
:���U��٘�����:�۽��Sy�X��#�F��$|\����y��6Yp��F�[h�l����o~��c��D�(�+ L��IH����KՓF��z��Ђ3`�XBd��EF'?���p?�?����<�6����j��h`H��ł�c��ԛ%"\����V���b�?�U�aU�t��"�e����c�j��Z��*9�c���{2��sE�gO�������Y|�@e4X�Ya��"��U.[b���uF�W̻h6a�q���s2��
t�u^a�b�[_��.���eۇ|��@�Oϳ��PE�}�|�\B��6��-��e�Q�CN���-vW@$*(\�.�eؠ�Q�s(������~M��H�	���5Z1�^v�kz���T�cV��Kb���b�,�ƌ�.����e����	=f��6���Y@��S �n���}L��'X 2�� Gp�����
�c���>������%�&I����~�c䪪}�/��'�/��ȪK��6�,�ߩ��e�: ����@*ۍ��6���(ꅡ��jA0�Ӟ�|��G4a�Pd��YG�R�� �GL�)p��]�����HB��l�u�i�MW��J�}�2��#B4݆̈�H1?�`�m�]�S�z��`D�Tct����-}��9P��C�+�O�u�WV��� G�tX���uC�j�5D~xPt`f��ZqSq��'[�`ĺ��#K�F�{�/���2`���]��Z�_i��x=s�U��Z DX-�/�ۙ��?Y���Z�|7+qz�;�k��J�.�V�0"��H����V�P7� P7.� �g�el~��\�ePߌ�kDbMaz��]Nׅ��D鹲.-��������]�k3?r�!�D���ʬl��D��t�����Jڜeԅ���D~�OWn�AV�{�A��vk�^�����I&�����@͢dB�a��5��|�1���B�"�RC�/�ub]��P!�
�9|bI����L"
�7�G�`Њ�?�c�#r��O>�J��z_�o� ���������p�_l�^���p����u{�y�.p�����
��W`Ŏ�:�V��r�Ѫ��g��ߧ���>��֕�ŏ@�_*T�ra|?����S�4>y�	�����Qj��^�wJو6�$P[����xtʴI�䷤�l�g�5�7f�=�p���Pt�cH�1m�T��&~bMe��y���hX��	����'�N��RDKj��\�S[њk���BЎ��>�V�@2�X�� ��0�1�k,B0��g �F`�`0Y@2�f���B�J@��2�q�Q�wRM�����.M�d�+��W�.*�!���n�V�H���z��mi���)��4�i�ʣN���a��c�N�ǘ���+���"ɧW��Y��zsXq��x2�і��HD�+#N�ɯ=і� �Ѡ��V��}����ڧ��n�v�;����+�am5^�����&_�
ܫWy(�%-�6*^.�v�Bk��\s}Y2�J1���w�|��Rgڽ�ω��q�Q�<�C0A���v��i�X RrNe1�V�̈́�_�grM�X��Iw i���]�?T렣�@�z�K8���,��(��n�]M�RZw�?���	Q�m��+2<�rV�쒇1����EJ/�+ű�-$����2n+v���K��
"�%���W<M��&fT���2�<��w�hW�P��+CCL&��>�6Y���\��z��4�������i'yol�ңV�q���"O��#D�ڎ���S��G+�,�v�d�<�װ%�(�W�ؐ�-��WdP�	<�NR�/Q�f��z4�ɤ+��\��Tןλ�`M��|��^B��g��S�3OD>�{s�^�?�"����V7�`@�L���z��֤a鮕�b)��[�o�LZ#>H�H0�}�2��X#�
A�s$�z�9�N5�N�h��$M�n���N��\,��p�=���ۜ��)���+c�yX�ZqG��[a,K�7��w�~����i���5�2Ü	�
��qÔ��>4]���։�������IP���NQ��<�i� �B��Bk5�e���G9�)��Ѭ,��D-�uM*X_��N,�/�T�x:�{p��6��Dh�N�{eZ�s�65p����A��b9�y1��C��*c��e�<�d7��A��.t:�1Ր�ȃ����8K���ͤ'
�"�Z��E,�4���>��"��BM�5 =vwp�<8R��S��1����8�����8_41G�ǐ&$��|B<D�c<'X�0���B�$�n����j�d!���Z�l3.U�I�Pt<B>��mY?�S��-T���&<R|5	X`pWx�����v�׭f��Ϥɵt��߁M7|p��g���Gb����YB��L1(�����1px�c
=�\�Yiw+�f2\L��x�iK{^[Zp�=�V�!��QOsޛo�͕֓Cn-(���gG��.ܒCU
�C?Y�s��L����q��Y��J�����u�;�l�+"c}��[{ч��;ȿqL;��]���7�OR\�[���4a�j/P��(�F0��r�����|�hW�}�0M�/�f�l���7SK=�mZG�����а���T�t�?xQ^�-<2-��L2�G̞�XRB'ijh��B��(�*r{3�5u�|)�Ts��l�&2L��v^c n�,3-�9U,�m�K<��@�c��5��I���1�y���	A�㓸Gb&�[9���ZÈp޿�iw@L-���93KG�*k��u�2�ޚ¢�3B�����3|�PV;0���xB�+�#P1�s|ߥ�eJI=f�ji�� j�՞�
5T�^#+$��n�Z�\�Hz����	>x���ǀ0ZW��_�f��9'�;`�_Y�@��r�qm���Đ�w�r���YD�vE;��t9k.7Ͻ�7Ŀ�'�"���_5�/����&���̝��y�ߏ<2'��G9�"v/W����4��1���yӐ}�+����u_�'���˔�����1לpY)W%��K�跊�]��mN]��.?Rv��ٵ�z|Dx��fp/��:�jd�p�/�t����q@��D~ج'w�C��?m���92.;����'ќ�쳝��(�_��o�h����S�Ħ�eT�j�0l"��J$!F�Ĕ�)Kk?"��/}	��!�ĞLV�c����,X�:�2b��E�8���>��l��J�R�{�	�.	�������9��;��X������S��qu/D�o�D����mԠ~�R�����1@������V}��[K�(i��r��n
(Wa$��U���mN�lb�%�R~m�5�.h�l��	W�	x�2���a�	x.�[
� b T!�6��Clt1��% �g��Z)`-��-i�f�
j	XL�i�f�����CF�����9��k�rj��g/ ʰ�E�6�� �0�0��u����9C��`Mՠ�7�0��M։�k��V0�̤��eމ�o�B���e�s�p��a��2�2�R^4�Di��hK4��u}/N��������eB7cp�2 "�Pڊ�34m����1�UM-��\�#���k�������`������<y5���|i�@����B������^q�fݤ��q�-̞0C�q���rc`��ϡ�v���n�w�l2�-i�)�{P���Sb��u���L�K�{&�2��3�5��nᨉ��=��1_��.c���N6��~��2pb����>��S�c��8��Q0�.�B?KL��[�L��:z;;����5Atu����� Xz�h��Y	����!��?L0K�I��.�����m1�^3�q���l^(��[6P�Jj�0��\�[ֽbz@�yM �l$s��u�C�3sO@�i�7��`N��h�3�*c�z�vB�<�ݽo�?M�ez�?J��M��ǳ_\t�tg|n�C��N��I(��ER1��6j��"	Z�U���#6d��5�v:,�X�t�ұ�� m��(؍)��#<�EB�ʱ��XW�E��lVَ�&�KM�@�<[=��bzB���17����y�@���] 2�����`�:�B��X�me��Rp�
o�x.�C�0���%$�,�N�?d�l;�-L$��!߲��4�D�%kad�Q�~�����zx�5�GW$4\0�W�e���zk�^��%k����L�Q A鲴����񻮅���k���4�������0KS�.l�"=��6'�L�Rw�uiAl|�u��[t����JÝ]�����霶}ʼ����[v�tq��Jܼ��!ӪPK�T�w�.��v]j=��/��~a���p��3 |L�;v�(�3 hǂDH=�jR-�k�S�^֕=H��-��Z�٥��Ƅ�4��{�c�V�{�w7�+�U@�Q�4��#�}��UNՕ��P��F1�T*��EUШ�Y.��OT��{�c��T��,���8>���ߺ��)?'Mî_F�RLsX��[�4�Kĺ��9�D�)�)�EJ!	�R<"�T}�Ʋi,���뒓����T.[�@���w��� �"�i��fu����\6�|±��~�!��$�,'(ù &x"&Y1����;�zIQ�(�0$�����9�}��~Zm�����?��0��ZU�+�ۮjͪ����l��;[:п?hv�{@~�q,�ӓ������KZ�j��f5�� ��n��KC��;���%�w)�����٣��$��-k5I��	�c՘+a�rl��e9Z���`?�NE朖yf[	�R謩��v�����������n%�Р�X,��������QPd1��ce��d�ūG�Pv���b�ө'����oл��ݔ�6%��D��e�Ŷ�Q��������,[���K �y��͖�����z�:��Zė�����=�-�6���
n��3ښc����Z���Ѝ�O�p��,{6���v�(g�)�f;ݞSǘ��Ud���k-�&h�2�K "�%�P�Q=�:����P���
?���Idb�z7�c���;�D�c��5
B�VN2�-/h��m�l�����Y_>$J����r���E��M[A�$I�O?|x�[�֝X�z������������w�Xh~�H=���t[��˟�o/�b±t��e���*a�z�l桀fJ�!rLR�
k� �s�&Xd2�e|B�W�\2H��ֲJd0��o�����dR�x�νp�ʹ�����+h��Hc�Nv�@�0@:�v�r�_d���R�P3�7�8R�*e:�� ��;�yFU����C9�h&�Å��e�t������^�w'4�j!!5HӪgPÖ|9K�<#��w=���D�����?��z�g�B�#B΍#���\�tPa�3����ǀޥ�P���E\����X�^��e����
R���ڞ�eZ���lg��m|5�$L��2�Z���l?P�����[tYH�F7����q��i�FD`�IA�a��9��(�K�a���2H�A�ϻqYNdxx4��.=��R0��*�ҵ��!Q��#F�Y��Q��n��S�"D�E)4����[n�]��h��m�m���E6݊z2$�L!TO����_e⟚.�ښ��Ú%��N	�A��c���yJV�=���0��x������v26\	���K��\�cn$̳�9��zCV�"̴2q�:i>�K��*��R߁xkG���D��{]>zZ;"pn�7y�aShr�����!�{J[�=�2.I
�,d�,��n1�Y�L�T��g���Sֳ�u�A��4�h��/��n/�d�.N�����Ro�������k�+�tE���.]h{�)�h?ՄN\"R\jU��'V����DbpU޷���r5ݷ-6$�T��q����TZH�@�X�_�>�U^�2�W���
�`�+i�����)�^a��i���P����ldڱ'�a��Y|3e�%Nb�N��|k����I��Q�������:�����+��j���
��xB���8�leʎ�S؝�:q�3��B���H0����`�� �B0J�C�%Ot � X���C��a���Z�'HE�*g�VMtÜ9����gG��b!d Ø��,P,��OA�W
�5�jy
ɤ��`��ri 2V3_����1�:�HP2�A,�D�B�VR������/i�alA��3�M�}�+�5����7��7-��"h܌��wj�8c�ڋ;�������r�[����օ�����ݯ/��� ��.oH�U!�4z�`��KJ��(7�1��C?< >�	�O����a��b)	�|��׵[��]I��x��m,p�Ů��w$���P�Z��X��PӺ7p�Ma�j�+?��h���"'�|<�����6�4�2xwH�^?��Â�5������,���r����n�gw�U�C�Cv_5��F�j1')�Y&�`�)��������!qV�d��u�-������3��l��ũ�k��:��śpS̀�n)�Qs*Ar� nep��Y�����<rSDq����oZ�2£2Yv�TcU��d�ɔ<�i�C��Z��hO!��{IZ@oJ��k��H-T���_\����>q�;A��ځ,���_G�3fj�]1!���H�U��9姱(��Z'���%6�K������Ģlљ����w�Q�� �6�	ɷ$�rjI�>����tC��Kݽ�f�/_"� ��#+�=c=��1	���69�M'�?mSJ8��%������My6q3���ŧ��>��3_�1�=*S�T`�$mj��n����x�&��+��."�!Ʈ�j-��p#�Ze s���֡N�����ꢞ�L��"N<�E1�oN�q:}��2t9�Y�D���B1��"�B1������R]�%YgYQ����h��݅1�C��X�C�W�U��y)��M20���L�~�mʸm��{u s�ҋ�|K%dV75���u�{�~c�|`ͥ�T<N���^J�0����=�bo���q���:�.��Lj�P�:�ά��9k�%�	�=�ќr/�e$o�§Tt'<rw%�\��G���6�!f�@©֨��I�y�

R�V��T�JReS�p��ԅ+iRE��F�a�F�TA��A���*KB-�T�PNv��&��ͥ�y+?�I� ��4�?�M����m%	�tuanV�ײ�JB�����[5eY���<^5R��FѤ�f�Ė��d��O ��W���9�ö����#���M;w.���<��޻9�Pf�e��e�?7��v�󾯙��2��~��],ot��Չ����4qN{Zsbw��p\��Ӫ\2I�`�p��u-�uC6u)˺��_�'վ�p���)�Q��&G1L����5O�1ՃB�v����bp���bmH�^��G�ɡ�}�)��Ѧ�<FEg�NM^3�X�N����-����L���~.�7-z�g�N����Ŭ��?������S�_;���ˈ�7��+N=q�]?�3��yJYx��40������j�W���A��Z������3������Y��,t��u�k�ŞO_�����֖�\�Ú���:k����5�*�L�\*G06HĆ��q�$[[2� ��)&R�ǌ��&�"#��RSk�d�}-&F6=���_F3� �P t�s:0o��,�N���%��h��xä�gͺy�E}o9��'�@��T����&������W�@���4���s_o=o�iw��(e )�����4����y!�$��7�@ɴ��Չ����Bm;�w�&��q�nN{ZoS���ӪFʀvh�Q]m�߆D��@3N���d}�I��ɮDO"�dA,C�+��dC�?E�YȾ�9'�p:`.f-�>��04���u"��L���-���8ˤ�l�Ξ>�n���0�����K�]��֢�SԮ�t�z�A�1��n�Ow׽oi9҆�8;'L�� ��f���G>d��˰ܜ��MMBҘ�A��*���@@>^@&�U�piq�AC���
S��Q��/�����q�X�l��6P-9�>\����[|Pd�N�-�w${aLXҁsp�DnH"�et�C,�>g���pfb�$���Q'����i#�p�V�'R�%������8����v��^v�k���#$a��ϾE�>��śPg��?ѻ7�
��.tr���3�y����te�ŝ�j𠨼�j�)�R��.<����|�@a�Z���N�~p)�r�D�}}l��bq°���Q�����ܹ�f�ܯ�>���@j�Q@��*#+hڕ�j�"�NA"�QCiPe����v��w�=���̬����&�ޭ{�S��3�=������sy���$s}�p�;�g�q��(ŊƘfa�����R}.���'m��lv' 8g�����77�Q�:�S�<�T0t�'΂}k����q�ʦP~c�饓�����8킯��i��94D�%ܵ��]J
9r�YE�c�w� 4��7
��&H���X�7�.�Y�h�;�LV��k~�5K�t�l��x�NRLu�؆�����r���OXh�#��vu�09Ȝ��3�:�s���pZk�p�=2PU�j?����k���A�� e>u~��RF�~�T�"ل��s��eXNK��d��	��7�&����+�"Co9��<�w��|�5�`��.�!b�#0�%h#̊2��r^L�S���v�8cV����cV0��k�����J[/��6�*ڸՆ��X_���}��4�U��м@��F��gA��sm�3��=�fbz&��ȱ��AI�s<x����19u�t�9>hT*�Bn���E���d�;8�D���`��������MF̟����r��%{���O���ßoY����/L�]/��b���z"�����;.x���"x�����ys<��1qƤ�|žՙ���N5(.
.�.c��J�u!�Ɏ��RF4�"���0r������N3�?��$��b�:b�}|������/<�C&k3t��N��*=���i#F���,8>jI?�C!l"��"��B�k'�:�j��R{Q!pvW�n8ln�٤��I�TO�S�����`�����ۗ�q�V�K�I�c�;
��?^|�iqM�z�9;�� �
G{ �v�mo�L���ޅ;9��m��A;L)�,�5��s_��ɱ�9!s`�T�	�k��_X�9�8H�2W�Qz�A�F0d�	&X�cm�4Ѕz��{�n�+]s���tL.��Cva��B�!�$ʻ�:�	��w������8���Qw������Ia��Z���7���A#��X,�m}��ϋ�C2�3 �3��|�M�t��V6��QEe=����SɭYk�R����ëJ�Iư��%}+��u��y��=�Y���ܴ��3�+�J�Kb.�CfJ�����wҗ+ػ���v��j��c��'��M�Yb��u����@�u��Ы�P��
x�W��֬��U��fiSJ�4cS0��U9V�Yvڭ�k�친��6�jH�^~]œ gf���=a��	oͼ`_`
�s��ZtS<���YIʃ2���vsߍP	ad��,���V�ȍ]�b"��P@P4��݋�I��g����m���!�	�T]ۧ�]����V�߬��,T�%ڈ��.�������St��H�`��@��9a���� ������������߃�����jL{��s�	�QSl~�`0M�@�8��{zd0
`�P�-
ހ�B��[�}b�`A�6s�8��������v3� ��O��?�G��iu��u$f���_�\|���!묰m-�e@��x��$I�X��C��P(�6��nq^?Q���s��t Lu���s�՛ %�N����)�!Zs�=9Q�<�'�߹y����U�	v_)+��5�9Г!�6�^m �J�j��س�^��Bfߣw/D���o�3������5��:�L�g|*s����}�Љ�I����<ߡ"��4�V�h{�(f�ր�	�S�nstI�&��V�x����`4�n���3`�9�m�q�ɣ%�k�jiG���"kBL��������QV������y��evR��x���g��Z�B ��:o�z��Q�2�U�^*��:ٷ���v|Ĩ�hS��uP��k��~�~��ݜ��C?>�sg9w[�\������E�~�T�fY��X����O���6��Z�w{�/�fp^]�5���������np��>���vj��Axm7�	�2�E��1��_;Yh �I�?,D� 4˽I�5�����M�A��\C��b��8��������_X�	�n%����{��x|!�E�����SV2ݲ��lc��Y �u�0�����B�M�+�����˻�CF�[�h`���Ľ�zi�ȫhZ�dט+��m��u���d�'b�BcT$7cF�p�7�U�0Hb��� �wc8�@ =>q�/q�t���<����*�A�!�e�5��C"�@�orO�8 l��B�cu�;Y��� -�Oܰ�̚yNa�
��n͢h�ŗa�X��۪�ըqK�+��B�E�<d��I��'P"R�i�4i~`ߌ����B�e��!�  �t��1��E�,����"��~�%��p��$Fldg��D�O�t�̝��_לd�j{������s�c����@'��P��7?���p� ��;yh��\����C�+���u������;�����s�B���a�C�^b��s���E�Fl#d�H׸��)}�� �p#{�;)mk$x���{FgF�N/��CF�DF�7��<�([���:0�=����c�1y0?I-�DK�δu\*$�"<%
��#3Uj��4r�]�0��R��)oYQ� ��(@~DɅ{�$�|�îYC�A����A�s (7x봑��]�J'�#��H�M�s2�s��Sx6�ve����H�y�-Bq������Cw�����[���@@�ԗ
=ӃR�4n�f��h�-��������^������Ñ�?M̨F���&%?rE�lnmc��GW졫$�ᣲ�ՀT�o� ��5���'�H������a�R��y�ȯ�Nd�B��Y�$-m.�r�;o�O�HIT;�'���cn%�n�
fa��s�yò��]��8�P�fN�DfrB�8���ߎb)<Dbtݰ�1���C�â�u�7��t�Qß)�'��~<DBtݞfC�d�� Å i��2��a�|m �������Ih6R�t+-VŲ��,sjM	��-�F�Ȓ�AFp�{����j�:��a�,���ͼ���map��}O/������K�����͓D5�
�;w�(u0_{�}u��d'AKe�+����rD%���f�8+�O�`g	SxZq/	�|�߿�-j��Mg\��\&I��[��|�%�b�_������Y��7��L�G5nU�^~5�$CV��P��X���Ҡ<e��o�\fC(^��B��&��4,�YP�����<8s���1=J�UY5?%�-�j�G�~J�)�1�R���g��8�;k�A������ٴO�'7f�s"��@���p��p��p�������
h[6�d��2K��a�E�͑�d�Y,�%]��7b�['a��~e��0o���%O ع�H��'7��X�ݥ�vT����t����`@�#6�� ic�qq[��ٍm:^��C����ڦF�<�K@g�����-_O1�	8��SJ^���0��Nڎ���6���2����Z8�w��:���#��;h.�Z�p6��5��G;�3���m����ӻ9��0=��q�?�MnG���-�Ү���y��W�N��ق���
<���4<"��b.f�^����>��z��Љt'L&�N�K�It��{�UtA/:�B@�m_@���mʁ�5q�9�+�+2>,�C�Ua���=��k�gQG�a�b�'�K�pS䰧�QT���#�m�LL��hi��9�O����2�fKM�O ����WoG����fh4�L�{i�p� ��J��ov��K~�{N�z�����9�5D-`{"��¾+˫jwo������AC�_�i����m��]�����2�V	���7��el7�p9��t��Q��i]5<��C-�*	{ݓ7Į��&��ϺZ\��L��rd5��!�\���H���!�4��܆󲛆7�0��Wfh{u��$2�!EUn)i���]o���f$�u��T�c����m:~�|�bN���\&թZ���/�8��ٽE���4�}�~�����Ul,�;i�c���޹���Q�W�H��������1,8�����u�����*��}�}�����Y���]M���~�� �P������_C�	�9��7߶���@՚a�*sD�HF������O���۽��R���N��$5^'��&�b�9��0k3���c�h�18��M���x�����0�0�0�0�0�г#���!/�{�s�d2�dM�������J1��� J�ŵ���l�=�읽�'ƴ�B�?���x��j��n:7�l��>�ݿ!���b���]��O�eF�"��,���rί��kE�c����s+�!�t�K������+|��'��1�A\_1M�\1du���l�X������Sِ$ùϿn76�t�˚m0�_� ��}�0��I�.L���F �.a��\n֗pqȰ*�HS�IaO/�}�*#8�Ѝb��7�3�sDm� �]?lԀ�t�pۖ�$"A��Hy�����v� C�*����kvPL�Ws���Z�[FH�mJ�k�N��$�e��ru2���I�$5�Wf�V��3}�}M�"�'9�Z�bB����f%k��M%x�ីj��p"�¾��(�9��l-p��񂁈ǆq+��է�Sa���K}
H3��x����lU_kLJ�Po����׀NO ���=�^(轶��%���	>
�TX�@� +�6�����u~T�"�j�,|L�FB�R�}
S��.(�>�.0���e�ƕ�R8��[��R Kt ��O��SP�9 �S��= �T
BCwx��sWx�������F����N���r�¶����)�ՍO���q����C�xP��/��!a5�;��pT��Ό���5=(���N�ib�&y�c;ʻڔc�N��YTgdP���fڨ�j�C�j�OB!�'C4Umc�@j�|���)�\[f��(�؋`�:�
��h�n�-�즯=�G����2pz:��w�'��[��HG��S��=�e*��u`-��@��]eՁ���ƤȱB�BG
4I;�ge��-�_�G�JI&���鶶*<�z���4�?�V�=E�]�\���^\g��k�t���(�01c���7%�^<���z�)��h�x^Rq��ra+��
W��������XOh<�����SG���
|�X#�m�b��*<	"�E=�"�e�X���0d�L��n���o���+��*��aW��U�� 3�a�X�X�f�L�z��R�Lim�g�c�������:k���~M+L]`<ಐ�!��%��N��]��cA�����A���) �A�yWwfi�Ȑ��.<��;�j�U�ق�!k
܅�+�$�(�:�'qw��nF
���CQ�|���D���K�^~Gtφ�b�';G:�7��R�q$����W�j���sQ�7��¸":��*�l����m^��T����Vog�@1O/���ʜ{�v�lӋ�lK��0���
��9'0��)@��E��7Vr$
����ƃd�����7�����O���OM ~��bi��\�~���h9t��aV�h�gM�����n�����8��&�|U����0���Y�q�q�E��j蜨����\�[�~*�j��7v�h!�'z����M�qs���$<
�Q8}')g�?�J��+��ջYᬏ�Y��k �-�Ymá��0�n�n�n�5��Ҷ�FA�>�i}��>3c}ʾ��}��z���֐�kC�GZ�ց�����cX=h|��
[�����J�c� u��36\#u�/n��	�gfɌ�q�D*d1E/!�šYʩfb�5�<��+�5�II,�E{z��V��p)�<xF����� �h�s/p��ߋ'���d!��׷�%Aw���g�>"4�'�O ߑ?�c򋽍��D�@�{d^8p�y�IxR0�r�ʞ8���$w�+��DO�������:%`���+�D�/�	�x�����*�藞�b%#5�F@o���1�jV��\{E�Յ뙈#�h[�"�ﾱ���W��c
\cQ~٪��4��b�=g��_�|/JHw�T�q��jҴ�݇|iN�~��K��0й�^���=��i�_��!�q�AHN���.���3ܩ/.<��܃m{�'�lJ0�N@?lL���=Y��_�Xl'=-ؓ�k���.|\����7�IO���l��y�S%��R���֔dAN D�ho(�93U}�Q�E_?�n�G��3�k�ݯ4��G�>��<��!ke�}ƺ9�r��}ynl���;�F��́ar�N���s�>�tE�b�v*D!�R���e�0w1oD�e��c��`����%��¾���x,?�w�dA��" DPH$ ���� ��-�gy��"���k�/w�kk� �:$��bt�.k��|�Y�8�~~Q[�g�1*�����t���O���ҕf���H�=� #��5o�$|�%�cp���_�vi�>]� �����:��%��-�@� ���{�GH�|�D	u�uЈ��"��!��
�.kD�`�L ����nL|�Q�#�G{��ҏO�_���B� T`�Y�(����#c�$��䦛���!N˅~0�_߈�+�Q���ܝ�ʝ6�Y�߱3t���t�6�	���M4��^��#���+�	��br�!XM}o�+�OK3���0�!�m��p�-���<[����߼���Ow
ml._�Z?�DQ�A;����R�ώގ��Y�γ���w���7��fze2'���eƙG�I����kK�����#Ǯ�M���IX=y�s����|��W�#�}H�B����E��u�v�Xm�����@,&�.���w�J[6�d��8LL�N��:X#�X`�+�5�D�E�U�$@��X�!�l��7]�(���4��1k�i����+O���B^�F$�\{dRv9�"[�8A��,���r����W"��)���Q�ދe@T0�G���WxY�?~���gK�Y�i�P�У>y�¬�,�	_���-㡪ޅ��:�����-��������[�d}�w�[�{|���A�x��R�V���W�C$0&�`M���!�;Cy��
,\0Y(`�He�cC�|+�#�Â�����7���M1� q��7u*�|��c����M(foش3��Ŏv�� �K��'ޔ$ڮ�a��n(�^B��\�����������k����l� �^{��VlW�/�}��a� �b�D����w����b'���� x���tN�n\`S�S�w��+I.;����4O��<<�-И���)�w>ka]�1qf5^�6lJn-���Bv!n�I�Y���eN�>b��)}~���ˇ�aXս����xm�r�%�td��t][R��B���*@;��L�<PXP�!b�������Eƚ3�k/���mJ$��ԛk"��lb�W���( ���|4F�Q�S�@���P����h�z��<+�X�J�a�S���G�"�qy.g]D�c�Rߞ�	�ƙћΗ��,��Rh��w�6�ӣ���+!4�~߂�%
T�E0܅���M�����ѭj�\�b��<�)\�[����	��.�D��069(�R���E_~`|�F�E��.�/��b&�Er�Q���]Yx���k� ��՝;'��S�Xꄋ�k-\�
¦N����M'���o=�z�����&��Y���
�F㵔��W���X?�VTȔ�[�#�h|�����L+��F;��bg3Oe<y:��U�������׻4ڪ�]�s��f�:!�vZ[�Mc�.�O����h��i�9m��4�5��G:�Z�l�m9���4�$�*�LF)���;��x��X���:�J�c�����2��o�gى�3n*]��c�E?0��������h���Qix��8�g�C&D5D�vzPӌ���:��:m�h��˴�֝����d;~к��0�W����Fx�`?TW l���̌�g�i��G�R1Ng�+�5�hb��>I�;|���ߘ���ʨn�,�|���}��[��>4�h�Z�tK�T��#ä5$y+�M�Lzu�I��_e4@|)�6>|���J�/�G
����?6R�bb۴�f�b�;H�+��S�J˯���ڎ,{A���G��ˮՇ^��Gͩc�ϻQ9h>�^!��f��Pr����k��c���:�6�gI}H��=�	��|p�,=�θǪ��tL��)�<������E
v	)�$���¢B_ �R��g��S`F�N��hQ��EB�z��<1g~_� Wðxpk�xpK�5�eX����oqV�O�¼�+sr[-`g�.^������'RKױ�u����P���F�Wy�A�L�K��&�4bgTV��ω���x�/��'��dJ�Ҋ�*1�Cf�4���X굎�X���V��jܨ0� �d�"N@[���ZT�$�w%C���cu�e�h�H��������l;fE@�l
�v��m�`v��S`�R *��L�[�M½�Z�����;���ৣ�E�$�E���j>�|R�G[I���r#���=#F��$؝�K�b�;��eh���2}˰�'�+���(�ɡ�q`>F���ŧ�>C��4R����۱s%�m� ����Wcr��%^�@��������;F�i�qؖ�Ç}Qm]��{h�z�G{�dX1P�"�{O���jZ��S�>���J���/б�Im��9��@ M�G��U�L�'����O|��y�gӚ���Z2Q,�ڞ#���N+�w�4�ΰ߅������m�qnz+�����Kd�뽃��6�ֶ�dۀv!�nt�䜹��挰�=��J2(�QT֜�FX�.�){o���L{x�!�e5m�BU�q*���u��{�[���������0��`�~gw��#G���do&�;�$�����k=O����T����v�:$������P}-g��m �.�����Z��5����n؉���2#�x \��,(I��0$�q& Q�@q��H
p	(��Qm��Ba�g_�������D���Y��i�(��y$	[�$(�+���k3땮����j��cN؛1��O��0�T���T �1��7Ѱ/1$x��K��ۈ&����
Κ���Zq�R�{U�ztq� [}@�!!���ۈYM�*��
ȔdAM`F��G@�)�:;�P�G��T`}�Fb�1W�J��dw�b��ҍԻ'϶���ӻdj��u+���_%D��,s�u@�*G5����f/@L���@[����!�(��<��8�y�!���nC�o
��s	�����Dv�1'���n`�e��Kn��,_Y�2?�P�;���&�K>
X\�az�?���?�
����Tb�-Id'�nk~8�M�i��ެ
�|F�!+*��0�i����A<y���>�[NQN=[��;�A���r�a&Ke��� �ۢ9�FǺg�iKY�g�p��t�>�'?�Q�Y�n�_�Jt�����>�^�#ε �_˕qZ+���*8F�j��\ps��Y���E������+�=�ᅵC�ﶚ�0q�ȟS�,p,rdK y@�eC��S���R^<>���� W��`��+N���K����I�m�C����M�������;���y䝊��`������k�V��%Y`!���C����
�t�Q��Zz�����	)���"6���^�	��r�cʿ�F��/M��-L|]���w����w������[)��Lu3X�fa'���=�x��.;�[�1�j���0@�	��L`&2dA2.	���EM[Y��Kٴ��}�3W8��4l�[2<�깪q���k��q!䲡�@�j�G3��p>�&?HR�aQ}-_e���c�`L �՜��B�U=�L)He)�L���h꜉�n�����	���Ux�Y�S��I��l�(��x��K����1'�LՌ7�
�0�DHVY�b#³�4{�ץ�N����h�y�����6�)ct;zEc1�;�eb�8�d;�E���9�����.j���Er��/��ۣ��,����%J�����N��V�S=J�L�4��N	=T0���a���L� ���~��Q��$��g�.��-#���2�Cz'��Ǎ�X���M�������$2H�!�*ٺ`��X��92������^��Ķ�H�M�
�S!R�YJf(�l#9^j[�8~JoI���/Ͱ��r�0�����i8�ӉF1�Ľ&-p�~������I���8�ǂ�e�� ���}��?a��s�cJ����cw������J�U29Ŕ\��̽�!��l��ͨ�MƦ��ԍ�;v2:N�����2��g�����{�h� ҷd#��Io	�H��nI�.�����;*KN���\��e���3?9n'��=�l��!�-O~Cd2p~F�]�����T�O� fvI��ޛS!]Hϻ=���ʜ�O�"������<(cÿSZR��{�cϹK���;�.��촥<o���<J9�������y��L��^`����'~I�7�rRr>_&�C]3N���}��u���;qQ���t�H"��e�Y=[��f��S4������犾���Y�.�3]S���h�]Y�W���dC�����#����5u`�]R[êÆ�ӡ7v,;*+���������
�mYkk�	�$�@ݍ���/�Yj<1�W�$Ӹ����T"g�<U{4�	c�)��e
İ���l��Y�r�g[�T�Q�o����hzd� X���Ȣ����u��)^ Q����+�A�_S��)���S�H>)p��v�.�<�ߝK�ݘ�UU.y���Bv8�]g�%�R:�c�2_p�n`��ㆫ�%��Ō}]e�}������-��[���{z�n��ߧ3O�zw��QK�7DEV�v�f�?�i� ˳������f�~�%�Ҕ|���H���ywau�tԸ��� _�/T��ǂ�Ƴ��s��'������!a��;/ͮş���V�3���5���{g�[8��9@��Wi�Wҹ��7�Tc(��e�f��q��Hm�⪷�ӛ��ٵ|�0�Cmj`�knm0��6��>���1��$2'�W�2,��m��D�"��Ԉ����kď�a-��#.���:�\���V*T#�A��w��#���>�ʴAճ�2�q�ޟ4:��y��m���5e�,X�޻��ܡ<sJ�~~!�4�}ᬺ�8W�ɸ�Y�V��b3���9gEWGk�|:|�~]�������ob��B�,eȾ�d��6�_��.DZ��aDcNc�l�Ej�D�F�CldJ^����y��d�h�m�r�5`�X�X�CL�D;�2��>���F_�iR�1(���E@O���z���(��ęf.��cf��Y�ct���ӭȽ��w؎���xZ;�\�}����|
��Ԉd4QY�­���:M(���Ȟb��De��j8��Q<��Ǳ�<Q��Q<�?�hS�i�MN��a�h��$ �b���$�1O�%�N�g@�jQIh��yIR#;8,ctmg��9H~rgB��0���8�D�<�]���q�ft.��sY ����^c��n���T���j���{)U|�JG<L� ��[���k+��}53����>@� N�_!b���q��n�N��u�q���vj�B����q�I�3¿�D���Ԫ��/�����O$�mJ�;;q�O/�����ߘ��ȅl>OQR��}��s�Og��0Aw/f���夠�%	m$���r%��ڢ���b?S2�D���~���]aϣ�7|u�x����g^P��i�<!w�n>��.�]�D���ֹ���6L6}k�W&��q��5�I����	����6�\7\�<������u�1��W�+߇��9�/ƟN��|oH����'z��������ʮ�^�����q�t�"kl�O�q�*8�`�m-��|��ϫf�B�7�a�r1�`w���n��WW	�%����yGa7 o�Â\w|m�<�������+�l�3��np��a_�O��FB�&�F�V9���x��o��^j��Uq�g�)����U�S��ʶ��٘��[	��#��kC�ﭢ{#�����}s셹V f{1c�_ݺ��a�?�o[���F��z��<���ؿ�pF̿}���	�����S�&Vc�u�.�����$w�S|<3���O����o�,q9��y���}D-�?"|�P�+�מ��<��j�z���&X��6����~�u�ϒ���?�z�B��FA�}��F�#:2�Dh�0���k9B�NlAz:�7���pkѐn��ሧ2&{�z?7f�!���"=��K� azȂ�|i1����}��#�$,h,=�i(1/�"ɩ���d�v0��2��xh�1-� �zHѰa�v�G9 ���q��s�S��z�+e����a�������ay����H1��ă�j�H��i0��u��w7LL�6?$U�U����0���B��>9{���A�̩��� ��`u�u#�~_:唙<ׅns�6~9�NX�j��'�q���;�<���12;XcM4P
���H�SIGX�kf�$W�J]qMt�y�Y��E[V�4*��ʠ�w<�Cڥ[�-�4P
��}AZzE�bd���Z��((����V|�*�ǉ�Jd���tף]�8f�?��%y�gxS(��C$ ��ݷΛu6{���=������G���DX��OI�P``Ey���$"&TȏP��$#H)!߉�	�./�$y�
 ��x ?�~�|���~
���Ы�S�ĀV��F����EE���`$-j���O�D&֤���|C�Х �Dp���O�W�'9�p��Q�n��V۰w�����{�AZ����l��@
�<o�|=��h�N$�+0���T��q~L�O[���/�`���㞌|_A{~8�#�C��
�X	J7 ɓ�,T�����x��(�?n��tP4�]F�7E�̂�!Ou> ��r*�_
	�4��KccֈQt�x-�J� ��x��<5��^SI��:P2I������3�w�D�A�:|�a�U��U3�*6����y'@N�z�}s��A���qQ���������;-�>�RY�LM�保��`�o}8�(dLNA� "�D��C�8��{����	�ܝ��c�"h,�Ī�����h �nB��[���M�����L�9��G��&3� ��?�^y�3�A���g؂=�y]�t_��JlQY�y�|p�ԑպL�i
��M[ۑ���Z|���KH�d?m�mW���t,٧2ܸr�PV�U���UJ���ez�h*�Qz���_�T�/P����J���'��\����:09�بխ�b\]��i��N�Im���ƛlF��$�V�r:QwǾ����Z��쵺|���.�y�E�mPm�"nq��>�ŕQ7�R����}���0�d��t��L��%:߁�%�!��%�۫��3s�}f��w� �K�4�o)�n3 yj�7p'���6w�%��	�+����#v�[�!_1NN�Y��ce�ڡu%j�j�o��ʹ�hk�'�\���fe�-�l�����~V(���oEW�'���(P����?�RW�� �$s�>�`G�u��X1Oz��2��~��<�s~.
�mU�V:���(���=3 F`=o��F�TЦ@�4#@&�����SU!?�;�`	T	|*H4���+ݝ��5/++n�SW����:�1}�ZBU�����=h\
z	\	LL���4��ў��3�b�}_��eOR�O��RX��z����6l�/�L\z�3��[�?E�*\Ap����Faձ�����h:t(��\�ɼ��Zߛnco1ߺ3���rn:7~�R���d\]�9���40b/�O�rχ1��(�W]��n���rh�"x!�L���SE�,oX�5������v!dˡ���nA׼���q��~� HN�0C�ڹ��zfGdKЌK6��B:fO��/sV7�|�+�@kX�u�Cl��Eg�f"����$CdC� ;"��ɵ˃Ϳ��C��*�|r�~��$�}ń�062BI��P�B#A`�2BH��R�� �%]	M.��LK�X�)8�H{�)�]W��
��~�`�o�UF�J���3�K�W��Z7��h��xS����8�n X!�$'S�~as?u���1�����di�R�8�ta�Y�^-gq��utW6s���P���69"nh�@����yQ�U��~t]:��J%�y8���RfS4�Y��c"`#[���
X9�
�Vi��A,����n����L}�����U��Q$Ed�i��d��ύ�%��,�2��2�,\��}���uFC�U�_�S�f�r[ڑ���}#�Q�P�.a�&�NB�ْ�e����E�+�"�6[���2jH&��p���o�'�Dw�������d���z^��`t��]
�CV��F�G�Ҝ���uܛ��wD�xqJ�]�j��+�~wBu�>PC�2�t2P^�x���ZPC �(���W��^��]�Y~���o������y�c7]6�
�-�(�f�� @�����R"��%x��~Z2�~o���Dsg�!芳F5�H!l�k"0�Q�2VF�JJ����|r�M���NI�,�uWQI�\;���d :t���{�-��{�J�6n��2�����}5~�	#�d�yG�V��=� ��B��#@���@� ��K�L T�#I�	�P��
�Ia.J6:KU�-02�J� #��@��T�!^h�X�
��M1Ҁe@H I�K T@%�&#)�
`�
���]�@M���� ����0	��h�
��N2������� ��TP%�&P#I�	�X��d��M@M@�@��S�*���z4S�Q���FZ`�xp�	��,�
hz�`5�"`mN<;G��G(�y?>���;JMd�@28�vW%��s����+�ndNw=�n-�*����[�6N>0oˍ+�n�r��BO���l��^��ޙ����D���/f����&��X4>
�d�'d���;�X�h��}1���ȩ".��7��W�آN�9I�d�|s��8�����obM�� �IN�9G��W��vsg�+��pR���8�ͱ�Z�5�ȉ9p�Y��� �O1̵����Q�����G�������a*d��������F���;�#�v^c�S����!e�:d�`(H�闘���E��_S���Ћ'�#&c�J�C�϶q�o�O����V�1��ds�P�oh�H;�ٽ�E	���n����J@*���'�6�\m72�h7%�7
��C���5�IG��Jp�i����7�bP�}0?FC=>_8|�����S��<��9��W�/��}��6���R<A����7�/�� 7�~���S�]��ٍ�Y�N�|��CUNg4g��^�&�_s2v�ԃ�ҋx#8�#˲���ǆ��2u�� ��q�?'����R/ۖ��wZuDq�ָp�9�z|1	�w1������F�S�?λx��r���8I��W"���8�#V��0o{���w|�֥�)S��h��	�r%{{���̆y]K�Rn�����!�Gyˢ�E���G����T���iδKxj�$��"��C9yǴ ��Ol�:���ii|o[~��Fa�����;C�wf��z;ڨrQ^����^,=�>�#A>B@Asե��@�^#����I��ɶ�]뙴��R5W�H�r=A#���m��{.��?�|��_rp�����m��+�"$���������)���}	�����e��f��ɶ�s2O9�1�a���9{�M�:��n^��MR��{�����]Y9Ept�l?']_�^���r��0��\a�c%?�mѴCFF�px��5�oJ�q�����xķ�8����!\^�3�%�]o\�ִ�v�˸'�X�~8��h�g�f��6#~#�.�r-�ǝ�7�Vn՗g�_�}x�&B2;y�B�W�	w~����mV$H�ޤ�Ǥ��<b��H@&6B��aă������q[�n#:���JO�8nK��o\��������<��(������WL��S;'!��ޓ<l�C)	�}�'��\v�k��U�xl�����!���m��=���ݕ4ٺm�=��#"��?�< �q˞ofv �dV����kN	q4�qf ]O�B�z�����Zf�3���ya>�'�R�k�͑�G\vwX�����ۣ�93 �$T����l����Sz���G�S�D��ayk�Z}��no��4������3�9u�î�!�7�G�W��=��:�Z]��a��̡���7 �5|t�5�8�Rw��'��VԨj}�D�@��?�X�F�(}�������*1���o�uQ2k§o���⦲q����&�%�]07=�}�a7_grJ�/B��� �����i�^Qv����Z��}V�5GY!�k�f뱝oU��to[��U~3J�>�y1ǎ�z	�w=
��6�Pc2n9;�CPj��� �7�R[���z��j�6M��hQ�����������/iÁ�D���}	�M)!Og��y�e�f�V�TMK���-t�]�=���ǋ[�~��6� U��%h����FzG/�I�W��6�F	��͞��\����k�@B��
ח�0��e���4��v(�F���[:��5�L|��EN���i�uy���5٤%�0Cp�|��gӟAt
a�^��a���^��e����V��qu�/d@��dV�n����9&��r������:R0��C�X���&���/0�� ������
�YWT���Y���� <�v�c�:��CDI"�߲�#�Y
p�߶�1h��"���e_��4����/�0��(n6+WH����Q�[+���������\G�z�ݾ֖$J�`�f�o�6��Hx��D�Ym�v�w0��Q,�;���r�Up����7�u��"SK_r|�E��S2P�!~17q�;�Zw�2	B�����7KVH4���K}je[S� o�KP�Ԙr�D�PD���a�)*	�~Y�(���8E6J����r��-3vY���`9>r.��K�F/��H�M5n�;v<L]6r|��kf^Ux��/���3Y���خ�1Y�0T�ݓ�b�,��<<���,��NY1: �zо�b�@��}�Eu�+&N$
�<���I70T�!���� l6a,,����`���dr	Hm�X�ݩ\k吘��VKX7�E��h���Č�ŉ�b Z�{���3(}'��W��Um�	"�c8|Fz|*�����Q8~�A�+��Ȝ>ɦ�#ԤWBz�ǡuF�h$d�a�R��oR �k �Πl��r��-	Z�:t����>���*��O�=[[q1�е���#���*P�Es ��J�)\��*r8:`0T0�<�~�8P���l�o����W]�ח�4@�+\������9��د��:����A�5�r9yw�ŎW���H��oj��̨̪�4!a��0�Yka3�޼T�����I��������(��g_"���x��@b�|?B�@BLj�d�ꨢ3ű����^a��
d���&�&�s�D�/{B�)N�eZSx��Mx�uר=|{������@��9%����Y��}��
3��ޖ��+�:0�/�<�Q4jv&�ه���`���=�'��^q2��\$���2( ��O6��Q�(�~P���Cz�����D����[8=Ŭ2���O�-H��^ȟ8�¾�����,-'9#���%bdSK����]�~*.5���F�c�?�֞FC.|���چ��fP�n����C�$��Wnޝ-��K��C�]�����<g(��n �O�N�K�� ���V^q�|!�:���B�X�I�?�HP�c��DJ��� vyY��ʷ�+�%��x��3���%���
Ɉ]�x�c�Ƹ��\*+��#�U���8���5o�?_�%�����e������|��$���a�q��BΧ�ꉁS��V08�����̥O��?�s��3�xa�̎��q~�vh��+�y�rc�� ZT�������~+r#g8n�e 0t����<����ָ���B�mÆ�q�3�
�@��~*��R����,	�:����NfC�<5�Ӿ��K�S�c�_���dP�I�٦n�0�/�2�t��m��n�}�O�%���m�̣�A�"�X}M2�P��;�Py�|�o� 	��x0��$�8�8�C�EgI���o�²��x�V˒�V����K��触2�����%�ơċf��)�Fv8ӻ���u���G��V���a��2Vh���:3ҋ}��(��)T1�0�3k%�#�T
	�5��9�����rm��xO\ 9߈'	闘	��T?˒P�p��&x	�ԟ���Z�2<yd�p>%�y��LC\��������k�B=�8Q��T��* K�2��o
���\& Ʃ����;�J6�*�0��acxC���+7��,׌E���� ��UY
��I}e�Y�������X�X 6�}���WT�V���2���5�C��tM��>���D���Ҡή��6�+�m邞�T5Д�����'���q��x�Va%�2	줼���^A���a*���.�TL��x���>'����C/�3�tZ���A�&���8��ZFƚ�b�k5�x �Ö�.��jz@;)������H�-�=�����(F��UQS1�s8�m]�]�l��.G��m����j��U�Q��$[aeA�+�,q�b[���ڳ�O�o�!E��}����9p�L���_>�t�`:�22<Kd�htbn��n2^cp��3A1����S�<X�N�]*6)�ܢM����N;IЛ�5g)�]pM�M�/��EIn4�n;sr�k��L�U�Z�[�.�!�V��讠�!�P�ʽ�Ӿ�= ��?��-x���&��<4�ܹ���+l�=9 �e��K��� �f�l�E��4aI[ZȾ�RѪV��Al�jEs�bN��}
r�y���v�q�3T�&��ϓ�~yM=��J�dʑ��_8TGIfiK�L�t�P��P���[vS
�j�����?B���-�J�oi�����v����A�g�q�R"a���ϕͅ�`�V��sL�����Ĥ~;dQ���8x��	��ut0c��r���,�.S�F��+ Ye���$�d��X�
g�۝�)��$��<l��ڮ�@�9hI�̚}�-<X�����m���#%9d�:���R�݂�K}rzR!Q�h:kMK�߯��hI�]0=��ϔ�3%q�L�;H|o<�>+���	=�č�
s�h����o:o��T�O���>e�A��Mp��C�Gɞ�ikaC�k+)�0�u8���s�<��_��O�[�X�GD]�?��H~&bw�
!�|m��O�k&�i/x�-�Ҡ��������]�o�{��{�RO�����&��񞢎�ں�a����B�P�wx��v��;�87���8?���3X��P���hh�����*FI�y�Vܘw�FKx��*��(��ݵb����_+JqԂ.Y���Qѝ�r���.8x�3�= ����2�o�R ��M��p�Ɓ�$�J6i:�W{P�������E��~�]z�k ~�^牫e�B���l�B�B����E@U�hXU@����t"�p^Xs�Z_%�M�0�rcbIhg��㈚Z�Xs{�T������ޕ��я�TvF��9flm���� �w٭����e�wH_[ĵ+��p��h�����L3O��b�n�X��1���]!$?�����;�q;��e���*H�O��U�h���Ai�ۧ�%��8l����l�XT��\�IE��P�*q.��Tt�ȈR�Rf��� �[���ʔ��D�g�K^������3�`��M�Qv�����C�8���d4��+�CO�!q �^[����/���ʍ;%��(���@���D%ʱ�����H�,�s}뽴����[N���ѡ[�?�s|��Lm!����O�ꩼm#��'�"X�i�B���|�w��|Ϻ>�&o۳�qr`q����z&�x����&����>�P��s����ǎ�>b��s�%�8m:�R|Gy��,���� k�QC��f|)(�w���������
�������9� sЁ���0r��Eh����J~UA0HN' �� ����.�K��n�G��I�b�A�h�cL|N\g�9(��W���~�L��}\���?Nl]����zuӨv���M:|nNF0��n�]c�N(�
�I�MTN?6�n.�lwvd�#�f7�;���#)��Z�p�k	�F|Yq��燗�E�t�,mX�,��$�ȸx�)�]>O�I����r&�U�ۍ��
�N�)���E�a%.�WO���v'(}��3��
�S|\��~,�	-lE�ӥa��ᖸ�0�I�]�h�Z7������њ��WW|] Ш�u��'��r���������lnWK�n2�G?[O��=폡�ā�u�V��
P;�0�a(���	C� ���ƛ���0��:��Ad�iA)^�83 �	�4��DB��	��z��t��i*
��n���׏���rc��O�$y)�8�ႍ�Ԯ�Z��xᝥd��(�����]��F`p��Yz*��ӎ9���y@K��S��Rl�-p�]��bH�b�A)�7�e���aL�G�Ù�y ��0��w��bߟ��Ù����}�#8g�+wxJ�8���~ax�;����ǻ�`�gP��x	���	Uj�(H$�?��&)8p�Z�	�$k+y�a�h�b�
�S����8W����U]�C���#�!�īo�������d|�1=��R�up�yX�9^
�L�C&7t2��F�`���zD�M,!0����]�v��=�&�5�ϝ(R��3�:�RQP�aO~���\#�8XuG��#��V_&���|�7�����AW[U���O����rOJ8����:/S���q���9��r.��w�~��[�z=rVٍ3�`b��]�>��ͮ��?���k~w��&��Yjc%���]��{/,�_C��C�!�jt.�������nY�w�-��E�j�Z?�8���q���`ֽ����Q�V�{���_p�d�;٬<YXc������Ҡ֝��
ݖePF�om��Y²��ƹ��`�Ƈ(I�I��d8�,v0�ȹ�?�6Kl"�3k������Y1�&�E��eȳD˾S�[|S���a\�&�#��2:&�SJC��7��|!�q=��F�]c��
c��[!X�og���������<�HNX�w�TYV��qϑFN5��`����?�ķ�fwv��dy�w��-�����@
�/��\Qnjp�z�j�u�=-��M�gzH��cx�
>ީ)?�{�^VTd}{N�/���	@8^x��#�8S�P.��q�2sb ��8�m�؍�wfY���;9CH<RSCT���@�Bt��<�F5e\��+ [���s�"}���[��Z�p���x?�c�~��������;It1|r��k$"���A�ΞS�/����Q�9f�f��[n�e�~�f-��ӵ�%nvǺ%v�ۡ���JPQw���k�)���!��'�2���toV�L:���ã=�uS���ʶ����ڣ��V���Ы������$�i�l�*x���w1<=��A��������~W�^��MI)_VԷG�g\��W]DS��L�DOoq�~&��TՓ��]�B�T�3�V�H�b� &R���:-?I�x����y�Y�5��Ϳ���w��a$'_�3��Y�e�_i��1���p�ߡl+>�"p[�������_n������E�ґO&2����N��\� �Q�H�n��Jt��f4�y[�5�Rw�m�=�Mc�K���#���.�k��/H�Ծ��_#��p�~���	�>�x+���U��9��� N�K�h��"�����Y�-g�!C"W���r{ٿH_���ԃ�
�K}�aI,������ƿ? ��+L\�}���ު�E�������������E����O��:������>�}��RͿ\�)���j��>���L�g�������S�H ��AWT9�� J)��-̘�|�;�l�q�m��dldUP�������,}�נ�9�&� �5��H6��׳�J�����_F��`F4�}V�C6�����E�p��u�P�Fq�ת��?r�E
v���]�-��IX��4�׾cDg�EY�*����Bp�R4P<?A2Ŧ�]�(H����1@�VT�t`�U;�.��E��(�^���oNw����mY��.Q��Zf�lG�4�@�����A?K��xhy��Q!'"�^�3לyq�ͣGa��,�f����O�gr�I?��oߜf�dG�F�E��Fm�W�V�O�t�ּ�^%oOwV.⬝gQ���l��^ '�����v$x]�xqz���[�3V+d�*.�y5�U��p�y,מN��t{�t�N���E��@�SWmv�B�j.�(=]��x�$Eq��eZ�_�Z��$?�3^�{lQә���e�����M��,oE�x�;U�li=O�w���8H�k3_�t�_pG��1{�Bw�3M��k5W��C���~�?n���MH�p�S�ֿ�M,G���
��=J��)8���j~c�yҹh:���l���?�>�A���^�^�ǝ��i��G��]�O���a
6��L�l;�-|���z�����H.�j�i[��X�
G+�s��(e���\����a��l�r̛����J�ģ�di�#_���y7V�1;�/nґ�p��������%�~��rq����b`��"}%d?����	L$����6U���?��Ƚ	6rXY*k��̧{�4��<�i��s���qucu�O�u���s���J/ֳ�OȮX�WC����"˭�������}t�<��B����0숀��S_�i��J,����K)�a�I���U5L�UdN�!v�Z^I���� ؀�g_D�5�������T0��ӊD~/�H�R +[9H��?NR 5k�8�:)�0�c�Ի2K�ٝu@�6!�?U#�9w�������Z1o����{f��ޥ �GQ�ZgdEJ�.�u�5��~%��S�0U�oúYa�G�!Lq��- mm<�x�e�{H(g��i�Y���V)n:�,�_�����zH�C�1�0���FC[�ey6���>�'h:��iQ����ןX>����1�Z;lc�={���q��m�5�zzc���V�#i]��R�K$c��\�+a.�F)���ӪU?(�lÙ�`��N�B]��!͜��C�$D���C
W�4��rI-�?�cߧlv�o[۬n[	p�s�)��}��;֐�T{�а��������l����'��ЯI���z�1��)!`2�G��x�43��� ՙE��n]8(#�z���頭���L�����ME�G"���!�?`��4�����M�Q�l��6��A�Qa2���q�zW�)�
�
�qJUW�5�u��!�B�'ݚ_@�Đ�o�{�;���熐��{���-������Z9}�v]�z��%��W�a�Ђ�m��Qˊ�+��;�^'�*��~J�*v
:;f�3�p'��|3�]�������)�9��]"������P���UiP1����e������</�l7K���Z����������k�l��M	������C
ԕi��c)�<#�3C��U��ħs�*�)�2p{V0�'f���J1~������:�=�_��g���@}s���by(�r�V�=����r�Ks��+�X��{�	p�p�o�������*pw��LX���GS��jW��V�qd�n���(��V^C(X��]t�UI��W��8�/��5����-Ӳs��w�gYD�/��Z����B�A�{��m���q?�.�;�U�H�C�p����"(c��>2�/���ͩ�p�d�}�?�&M�v)ꛭ�������y�Lߧ�x�O�\yԻ���ά\p97l�����q�ѻl4��5U냧� ��'H75�-�x�]�7j��B2B2B2B2B6�Hi�YZ|*��Z��@�n�-�B�(�]�m��A���`��Dc����BS��/=Lд-�[T���k^T)^�mt����[����qm�^������ �����ߩF>oiH�6�L=<>����1+���7 ���	M��؆���0�K3`��;w�m��Xn;�Pw��+�w_�9p��Xw-�nl�t��ګ͇�C\k�R���廙n�q��1�im�{�i���d��� �g�O6.&�����2�p��,/N��Ǘ���Ԝޑ@�:7=��SLl���~���Ն*�%�X��A5��7��@@�U���uЂ�	-lFP�\��`F�Q�@��������J�t`.�K���5��у%�r���h|5T��<4	Wgg���Jz(�ʉdX6r�>�b�4�ʋ�u�yhnr��t	��MB4�h4lu�,"I�����F�y�?�ҙ�:F� 4Z����tw�"�r���3��Oy�G��q��:�����Ԇ�`�:�`!��zp�5 ���%�M�������&�4���q+�U�7��pVT#�Ȅ��HVEJV�� ����ډ�����b[��]E����Q[ٯQ��b��6�0`�h�
���~��jR�>�b@���~���/���|����?/FH4� yr-�}�c�_��\>|�u��$�U�0
N�ޓ͠OW��pVNj���+��>I��/��@�+�����>��Σ�3�h0'���ok_{�?��I��ރ�h�����2���fL#��~����[X~�2�г�� Ђ$j�^�C�d�V{s���5��c^>�gBi���D���f%�~�"{|}x�[�[�:^-[�+��<
ۡq�9�FJb^�+[��0Pϊ(���b�wC� �Ye�T�%���?B1؆�}U]����h^�
�Ґɜ� ��o@嶕��zes�w
�� d��4lM�ZL����|�={��7m�``޽F_��K�Z֯��Vu��ٶ�hT2�="�<���?w�2��&�]��w��2�J�~��Dz��U�g_ͳ����<KC9�u��	�X1����-���.��8�E��p{;{��昚��lz��E��[I�y҇��Gy�{+?�j�/�Dy��=�`ɠK��aO�-0*Ш?Q�(B�Z�\��$��������L��\��\�Gi����a������[(����t�g��y���2;�G����4]��πf���Q��I��]�UVJ���<�W9\��V��x�%g*���:,�T�󭤭�0L�f@��E��E�m�񲱔�N!Z��LQ�t�����o7�Ag�ݯ��$��P�ʘ� n����v���M@:��-x�i,����p�n���`��<�:������d��zT����]�4i�9b|X������\j�Y�[��K�0`9��v@�)�.;m��Op=�d��Ͻ�ˬ��S�'���dKN�$��۳d83}��A6o���v]U�_(�*0Ɗ�ћ)m h^�pk�Yr,���\_l{�[z��KA�/�6T���~oqH$��.�����Y����v������J��T�ك�I��6ƞ����*SSܕJ����[@V�+������d<�"l���ҭk�GP��~�t2_*�����4��d_\���vlC����4LI/�cu�H�ԛütc�j��.s&'����'J��ж����k�-%����ʒ�UпM-���^�Z�X̴1���SN���2BPn"�����0�5�#��M�G}�o��J@=Q��zS~�'���6"��X�|�g`M��!�����֖ETZ��b���Eh�=�_�$/|0[L��=>�d=��4��>g������w�ʰ=���I,� X�ˮ9p_����i0?k��w.f�v,�u����ǉ�=��WV,N9�dR�b�l]�$b��m�����cob���ܶt@� ������ "%Ԛ#(�!�x���f;ʶ^q�͜���9���ln6�3qfV]j�
����f3nG�M���w�d��kp۳����Կ�*�q�����ǿ����m�=�oD�>�E�4&�Q[��JzF��X1��|fØ��H ���_�{�w��}Co��s׮�삤 5+����:��@1&�7������P8��V90�y�������-UL�Ay:�qk�
'1{P� =EN��Ę%H������/�7���sn��}�
:�2(��
	W�pm�)�yBꉦ�J��S���Bw����V7��EcyY*}Pf~I9��:<I�}S�Δ�Jw��=ٍn>�HL�3�oB��$�����M�x��B~�B1���[�),#���q]�=�U]��5a�t�711����6>+�bU�j|]���} 1�W/Λ-s#ݯA>���n�����zB��BZe"UW�\K}�O�a,��%�BZެ,������%'|�x�Y��HO��	U$a���"���^�]����NDG�؄��Q�p'���n�]��<?��k[#;`���7��%g\{3�N8t�Z�[4@P��H��F��.Qe�D�����D�Q�`����Ѻ�Q��Mhȗ�k ����sAz_���W��|*_X���E�9��j����)�D6��5����L�5��Rξr>�{qw� /Va�".�Ρy6���cVDw�~�J��޷�����-+��nǸJh��b<�,]�~VB�Ql�ٚ�*m-���DV��	yd�حb�;�-�����E�0#z+?!�J��R��:M�������l�mu�d�|/��kpT+fM������JE�+P��<��k��A&Dneã���&o��~�E��1N�P����������W��?�b�\��QU�J3���#U��R��.�gk��gWe|�h�1����>�k��J<�}�⼩N�*����k)�r<����r{�e�eX�
d�B";�DH��sc;�Q��D��hY�	��qK
��")`�L�+�E�X����ܸ�h--��>yFfF��#X�I�ܨi��&M&��
嬜)�n� ��a��n ���MOb#M�0)����)H9��f'�nn-=K5��˒���%W35�:+�G(�]lo8f5�i�	�N�EG�d���nT�1-a%_Tu!���ˡ�[�&�up.�zl_�a���G���8�]X�bPs�K�+��(���Z~B���8ЊB�+W,ǿ����`?ҟ7≎�cqC����V)�#7�>PUXѯ�!jj�6PU_2ɰ�j`P֍�4��h��������;����|�LV��(�������yߖ��v�I=i(������"¬���o���L����ً���>l����M����� �=�?N��`x>�9ى�"��/���&�@$���Aw~�����.���ϱ�[�.��'�REk��F�7*鱔t�V�6eI+0b�ٮ ��4c'���%�҃��(��'1��?U��G�I�� #�\���U2���o��`�Ø�'���Js8����l,ETj[V��Es �x���s�I��̾m��V�L\�N���oNɡy��qE��e״y�L�'�E��ͦ݇m�@����"U��d��y�h$�C�a%�i��(��:�M��c�wbo�"(��%�lǊ��;֋A�J�^ʭ��o���	��>����ͱ���޲�r���*H������=&P1
�iwq�����2	�ر,7��1	o��zXڒǸ�:��(��W�M%������a�:���"��sڷGnqΏS�&�P�!n�|Mc��t>��s���;���7AdrO}��0�����Mr߳K�i���1+��ujɽG�`�ԍ���$)rR�b麒���Da�����v��&+�m���L���o�ûQh˦W[���Xn]������A��k��JF��+��o*�������o
?�a��/s�`7�`S�t���n�-�a�q#�7F�C.�aT�',ۨ�"�;)�xg������^���R�=E.�`$=�ϳ�b\A�]L��M]Z]�J$�-�~H��v�K��dR����i�*/��.����ԄZ��GJY��j �1˗s?�$p�aM���cS��OYq�M�V�������U$$oWE��%I��g��aH����sq��<�HyG�LZ �oKr��e���]yȘ��)�ro��C�u�}N���rK�X{荘#A��U��v��Ƿ>�{�2���|��f
]���ܱ)��S7z.N���a�Ԏ���8Wg��u�]�	�^�qO�D����Dԕ�'�1�6�y�H�T�:��)³JX���3��	^R@貆]�X���('֯?mdJڋ�>l#��!;�XV�˼ֳ*&!�׿=d(�I&9����9�ob���b����)��Yɸٮ^���|����D2U 7c@�T��f��D4�7'���%�=��ޥ���G?�?�b1�l�Q`W ;l�o�1a_�d�&�U4��3���=[S��.>�b7d�om����ķTV��[���]���U%�9X���X}$n��nk�X�.�ԏD�����P)1M��G	,z�8�8V�7v�#4�]�H����{��N�$Wvh_���T� ����돿y��̶�}߀Zp��&����3z�X����6�1`>�ǋ8�魟�:�����Qro�P�o�P�h�I�ěi�bhm�:f���;���m���O�u�\JM���}�#����A�`ǧ�Ac����͍�������U��c�
��s� 0ZW��\ ���I'�6/N7<ǁ�C�]Fy�&D�\�'%��،�8��A�,Y�[��ɩ����/�c��4��3�1��dS-����!�u���K�Ci��̐ F��}�Z�oz%=��^�����/��e��&�}5��"Ǟ��R�yK�ʷW�$����teؚ �����6R�I��'^U�G6%��o��6�=�C0��"/��ڶ���]��tHx�2.�
�E�n��A~�[��^/W�0$���e�͡UP���;���6�Ig�L�I$�lI.\Ę?pk�&�E�r��&R)����c�����͚gY0��Q����J���6DnwRx��I�����1'k﫬�J�P��ë��1���1���v����f�2��U��i�H��mp�%r��J3{����]X�p��1r�ʅ�(ڃ~�=��Saq�g�K����uT����5*���zB ���VP����(�gf�]�9B�$�*�
�r����UNq�}%�ZB���qC�ܡsNg��$$�guC��."�Mhz�1f0� ���g�:���q�m�\m�����.���<�=�5N����|�[3n�u��ј�"C7#8zF�6+2z˄9��XL3LPc�R6�N�h.���� �Ծ9af_��� m�]����k%.�RA����=D�.b�z�f�Q��5ȵ�e�S+;8Q�%�
=��|I~v�oIy��n��1��X�Ӏ���o�`�!�$�U�`ѷ���PbC��׻B9���1�A�'� |B+|��̎?�BĢ���f6���2�Ms��̲������-a�H�Yc}�T�� \��I��e��a�H��fDg��&��qfYv��
�hX:5���㙐(_�M�܍�d�0T�)�SSf����I91Q��
�����6����ټ�;H^Nd��q��^]Ixϋ�౪r���5ZygK�5a�m(_���1���9m���<��)���
��wMM�ML��ib$2Ӟ��^��`�zo�7���������T#o�>�5W��W�R%D���j�KO����fȉH��a���tRUKI5ku{��RN����M�H��{07N* ������Ԙ>G�,�i��U�'٦���Xgu�x�'��wN4�������@=���"AmYOp�_��M�A+=9t��I,�N��[��f%j�g�_W���tB�-!���i��M4I?�F�Z��x4�߲n����
n�	��*�[�ʅ���8p0	@&e�oR}���=�t�`���N�Y�VX76p�v��?�̹�]�_���N꧳�(���Y���� ��MgW�?� ��n�u�:��~f=D��e��1�{�52S6#@�AD�jY�LHF���;���-:[݅Ic>d��Sɱ7T��=��� ��H��uhL���(H�#�Dچ-��"x�$��[�����h�T��<Elm�s���ퟤ�'�ކ)�k�yx��e8<�Kd��+ډC{�1����ԅ� �Z���T��Xy���,�0`Eh	�DxcQ�u���+Sk�ɴ�C4��-� md�W�Ox�7�� �(-�8�'4*�� ��bhǘA�Dԝ�(m.��0��4���L��~����$����dτl�&��bK�1�ؕ�F�Vg:*�ER^�N��+F{*[�%�nl�g[׺��=vI~LM2���aI�f�j�G`-�8X{��$��Ae��Ond �Ύ�]��ϲ�_]�7cH�%�:�;��׋v7f����_L���8ʉ�u��Lk�o���b���JM�{�������J�Y��^�=������D��D��yr�� ld���]���J>?�/���d��y�a*�-Br�p�:�p��Fq/��:�/�� c�� �J���DP��I�����\�Y�a�5wc��nl�)��ݖ�����E?\�L��$�	����Ք��]���+�B�����E�U��"�@�w����C��Es={{�������x��7����n�����?����bT~e�W�Ф4U��>/��ǂ��=T��̫[�j�����/�|����2]m2��G�����{�m�,L��"���*n	��ׯߙD�T_n��O����G�r�_���������HG�FXp�H�A�'g��RTv"�ljF^�2^�ہ���{]n��A�Ņ�W>���,C�j��{�%�[������ƺha��?,��eh��|�����^d14| ׃zÕ���7�K@|.����Ft�ፀ^Kۦ��C�-.%Zz�={��@I|\�K.?�W��,�l�^I�����e����l�ՁDg��C\�]ǆ��J���5B��}�*j\���X]��r3Z���A��j#J�I�~?Y̸�l�C�8�&��X��c�66e���yl�/+��o5�?N;2���M��.�fc�M�{��3t��2�k��({H@�}����M�<I_[�CY�~�N��vaol�d���Q@��~�N�N�Jm���)a��e�b��z,`¡j��%���9m��z�5��"¥�m�d�}�K��6��o)�ۮ%�c,l�i廫��d�M_��a[�;�4�e��d&{!��$�e6��jX�a5ZK Tu0^P̆�GOZG�Y��S���}	��6��(���F�j	!?�tN����(Ur��	KE�ݧN�S{�Q��f=�^$x���WF[��Uv��T���Ǟ�)G1t�Fe��6��2Le>Hɧ� ����3�R�8v#�7�-r9Fw
9ߕ�R���۳ȓ�_+���O�s��.?�50ס��A��=4ii����(�'�R�:��F=5�8U��9+#njP��=�mT�$��6��r�B	%#��:,xm1�������^����uN�˝7�R�e[�_�0~[��F���sv����#1�DqNDh�Sp@24bNAL@�]Z���1
3�7�� h.��,Ib�J�k��
q� y樸��1u'��`	F"Q�-���RÄ4���m0+�}�K��h��ͼ�Ui,��3� ��h�&G���흍���ٰ֘���ʩ�W��q�5�L�|�����
p�v�f�P<�x@��Giblx�2�i�=Ż|�YQ6��Co�1�,�ރc��A��-�Th���&���׮�w!kEu�8O��+��X^��x�g�Ӗ4�I��C��h��3�)W�\�h(zS:���ED�ܫ#�*�2M�C
�b���?�m��?f��3.��s0N|5���LP�*E�:�L1����"y�Ȍ�sn�[2x����4�9��}6n/��kF;@W��Hq���=&��TL��͕�Z�����/��b�[���&��m�X�Џ4K�f!ߊ� �!&'&O45p�Zac�Y�q���1\�&��o����0��H]�:�1�3�mZ:(� ���2s9,ʭ��0�B�p����;��o���p���� ���+n.���#��-�Y\!����p�S2�0�.L��<5�_�X�9�^M�n�#a��Eܻa2__��h2N�y>�i8��f�|��w_}I�B�U&ԧ0-crbU>(��G�4����K����{���G�m=[�zA�c�C�k�0�U����� ��w��\��Zk�ބd�j���^?� z�ɧ���^[ր�������{��r�E�O@���TϽ����Vݕ���+ئ��Ƥ�h	�7#Q}w��c���[�k?�,�����Xӗd�~�����e��v�!����q�ބ�c�[�l�<٫1'�(��,GW�B�E}H�+M�ߓU�չ��ze�K� �k��TuPV#sj��k�����Z�˃�<�lC5媓��?Ml�c�P[��D���!vɿ��_<�᧤MC��xԨ�u`NN��Bd#CB-"S�$�_�p�-�e�t����������-t�Z�r ,���訝�6m�	K��Q�JJ��#��!(!�Y�3&����O��I�v��ҟ�)|��J�������\�FĴI�;�7`gU@_�+d'*Q_���E��N���Q�80G��H����º��\ы��e�q�ո;�Y`���[2��g�����p$Sg���<���5��Bʚ!��r�KZRZ��O��O"r7�����ߎ_��z!t�wl���+U������pz�+0��mm��zV��>$;�[��nJ�~]z����c{߲i�-���O��8�̅=�^ɢ�^��cp�K-$��}�H�N�%�K�F��ǁ	�tj
��H��ɪ(0v������&?t��{�5�4��bIM.�w�@ãp�m�%�~��r�F.�J��Dv�"�c�V߉p@��I���)��o�iո4�n�P��+�Tx��]�;����*4����t�f_�5����m=���
>�A�3�܂���BOG��"6]ؗ��
.���'�hlz����H�K�X��])�R᪖���pT�b��Ѭ������UGB��l`18=E;��}�2��a�e���Ch<bP`�N4;��ߠ���kL�T7��ۧE���M�O_D35[����%f�m�!{�/wT"w�@�r.@���"���@l��6QX-��B"�8F��
~��{h���E�y
ާC��A��?D��:�� �-�X�ыc���b6b���]r�3q}�6����_�_���_�R�s`��ask�U��|���{�1)e1ɨ�/J'�i��J`�q(؝�_�oNɾ����\H�كE��N�Qf�W_\�0p�Qa�y	���]�����hY���"�跳�E�.9�!�4��M�C>�F��P��8�vu��B���KC;T(<fp��Ү:��B����}[,,,����,<v�Y_���<,=l^��[ɔ0=sh`~�mP�'U'���Ĵ3�CC�q�wa�j�����O!�,8?�y��j�뼜oP�O�ç�%���xx�C��]�bv�������뮯�T<,�H��Җ�N�u/ʺbzW|W�*�o�D�Cr^� J�S��pҾb{B�*)ϽY�zx���i�yVR	%� B~p
ќgG2���n�k5#����ZL�߈{�^��P�`�\��AZ�=.T��js�"�3zt�+J��
'ҡ�0�4��n��@�ܵ}�û����~3�n��)��J�N���]���%l2�j��*�UJU��:��ʝ��Y7`���n��v�v)��ԗ��s8޻3������ۭ}�9�{l�
6?��&��\n�����Ǻ�#�y"'��v�]��{�)�����Z:UA/�i���1a=FE�E�J�"V-c�Vq�B�N�>��ߋ��xm {�TS�Vl9ѡW�F�>��1��z����E���4
�*̕�dW\}�����j���9.�l���D���*r�2�&��d�y	<t9��z��S��>\����m{>~+��R�����:l2ǗJH��{%��Cўo	Z���J�jp&v-��'�gY܉ɣ���i�|<r��$&�O'P>���L瘾4Ca�*	�$;�9l'
G(�}SՎ�X���J��[���[/Y�s�p�wi��R���/.S�o�sg�*ğ�%|�M�����Y��􋝪4x�49��\�<a�ȩID����Tg$x��&���?�I"��������l0V��O��D`��^�HIk�+#r-��9&�C8��̛Ќ��Vf_�ի�h֙\3:�/����I�k"�A&H>'$�/�
_�\ct6B%�����G!) ����1?[p�^���q�d�~2.AL��c��RW�f�|Jr�o��g%q��4zʭ���D�kkϢ�S�PzFֵ#��i�kOF���d���r���oa�3����i�S<5�M�5��Dk�g�S�QM������Ou!"B��ȝ���T���J�5�>b5���;i�P��;
��#T�e�y^�!��h�u��M�����)�����`_;Hm_�� �2�qPE��<�Y�*�R��ϓG��1 "+W���&5c�-lgu�: �R�վpƷF2��d��熶��>�#�|)�`�E3됑��޿��	��%���;���1S*\������VѦy�������TR/�:~�zn1ӟ	y��#'vK�oo�}��"LRl�\gU�폯,J�I�%0ne
BG�-\���&@�o���p�'�P�6��P~�RU����;����hz1��o�)^OC!��1�.�#�#�*z��9�]M�O��F��4�#�q���0�q׃9O&�-K�KF�!�ng
��e`�̸$�^|456�]W �e����P�����m��ło̎4��g���2���������E�b��?�;8�BG���T]�}(ȟ�Yg6���������� gғ��A�E��#�s@P�H���,�Z�������`�Ĕ�}A�F��c���n�z0�O
I�T�r�m$l�u#%X�HJ�EJ��`b +�6�w�ٵ')�-Un�2�fa��P@�2��x��!�X"?�k�Tr,!R��r�q�X��ו�C��5�Y����=��|��M�m~���hYP��P�0���\��$�^`硍9���8!���a��,4��}O4��}�@�e_�v{f�ຘ��D���@����������1^�
�LǓ���0�7P>�������.���ޱYg���TJ��9$l�mh�b�-�[�(�TF	u(�J���8�<v����;"����h8?��2:D���s'�X6�*���H�y�-�z�r���ob�����;�׽w}~q��'g�H�R���8�Lr&Z�N�Qo�/T�`E��rw,��i�-�����y�鹨<P5Ff��$Q�ã"�B�S��JirR�H�o�=$����F����@=I�0����iŧ�?|4W�tH����v�L8w݇
�E�A��4_B�����5�M �4/D%D� G ���� ���@&�(A��"�ʀ�Q�d�p�aON0�xI��Σ�;m.�p��/�82�N�S��Og�}S�DЮ���HI����˫�PlQ*�� ��|+��T�����p��5!'��O������g�O<������^���o��V#��爰E%b��[=q-�J�E�/qk`���i{\���Μ	��1���#��p��1Fh�z���#^�u�J$��"��)BX�}yy�_��-�d�0xn5���AQ���ݪ�*ҤǊr:�odz�Oa~" XMAah,��8Z�1Dȸߧ�����w�30��A^����6�	��;��r`|M���f8��1u8Ri"�vsd�R��5L�+�;���r�Nɝ��,�W���
�W�	���5����/���AÞ?w��maogn�굁p�����?�@*2�>/�<y�P]�I�%����������-��,�%(q=�XI\6�*k$	n�<�S{��|�L�:�B-!V(�8wx+��+�����5�Γ��J��W!	6Ɯ��d���*���'vwGIc[ԥ�:�&��\��Z\�5��#
������d������̬����Hj
�*��
?��)W:���܀���*8"N�iP�K�(:��J���O�z��3��1(bL��4�+��e?l��3�F�t�m���&�DdR�/��b�0�Ng���]u���Q4e���ek�6��Y��烱@�R�Q/q� ��s7�F_���E�'��32Y��BDj�l^7~
qඛ֔o�{�+B��8!VF�T'0ag���͊��?�����'y�k��V��:�`�פ���j�D5=Π�e�?������ �H�������)��E�+�2�УI�r������U�r�q�"���@P?䏠����"��{R~]r~�ۨ�x�@�h���w"G�2[v���s����*;�Jz$`ȕQ?�A�y�¿�:�.q^��YO����<�'kˍ�&��ƍ�c�n$t��{x����;n���Ȼ���ל�#u\���%T<p4~X��X��k'^EB�0+O0y���a��A���J��d]����6G�Hpf� ���Ϡ6�#��n\m��Ȃ�R�Z��Y\%��=���K����RI򞐎����bE������_���w�]Ye��2�e�D�L�"��A.g͉�v����WVƅ�to�!�o#��U�_���7\>��f=��Q�އ|�_�+�f*���!ԲW��j���u�	�*��c{+Cp(z�9�V{c�q�"yO��to�L���A��30��9�DЌG�9�A��"��#���ll�yؤC�B�"L>��T�(�5�]���Q�O��s?�Ά��"D.��	�x��u	٨&��-�����[�ꑄ���T�N�����Đ]u=g���[.=�o%P0��+H�E���bA��r1��˸��?�pGg�k<��fE:� on���=ݿ�]��l��S}8���}�x'�u?�sN�c�}F�6�M^W�`�9����[ۼ�s�m�\U��H��B��0���Uj�֋���Џ�tݣ2���� ����l�� ��cC����!C������0UÀ�-��`sOy��!_f.ZȾ�mo��aJl�C���`]\c2�H�tRw�|}4gP�b�XR�'v�ANh�����F�$�h�7�{�Dh(�&2�F��6�y��]�/�ĸ�8{�q���>�U�a�ɡ��E�<,T�UZ��Ӫ�h9�s�K���5�[O��Z����[u�7���"���"�����������E�<Ur�[Ov�5�lCP��Z�)	}et��#���ҽ28%���Z>�N�c��F<�l��w����!�z��ㆲ�lu�n�g���Y��9�G�W};6�0U��]�A�����x��;)<Y�kx��NΞ$F%��"��� r�ڥ����ҳm�֝��H���,@%�C��v��!j^H�`䠠�>H>ga�t
I�!����4�$�g�N�L�W[H�VK�OK9d� �{_���� ��I �3`����y�咴���1���
�M���"�O�]`�F�6��@.��C#�4m���2��B����:m����!� ~S2�C��Z�%���AQ�Y�v��,q���1��d S����G��xoz�d��Uta�Oɹ����CK� ),!�_ۂ!K[����D�أ�
�k�VŖ�. �Z���Z�$�&�H���r���<����0�h��}������H#��>PKY��9��Kŧ�/4�. �ke�7p��Z��T�BId������U̓��!(+������Rt,
Wb��	"��ٸ�R��7d�Ƙ��aQ�_�Y��z+�m1���SC��͘�ھ�%5�;Fq��!V�h�̻��~[�J�ȫ5~�!��h�|��$����>����t�D�{5�p��������>q}s<�_��5_J�:-0� )�� ��`��"�=z��I<��B�Ɓ�d�)�������9��6V�`[&1ǹ�[��ɖ�]����%���*]���F���!$Ҽ�
 �I���_�B��qReyQ9�n�%�fr'V�<��⩰�n�8;���2����$�؅q*ʏB��� .})d�vZ�k���\ͨ��(�IiL�硬�?����jJ���c�Ù��h��_�f5����_�T:�H�e�<ǥϧ!��/5r��Q-l�:�����QU�k�'0)U:�G�J���2E�+��Ǻ�A��#��ר,��0�ҏ���ZYCp��(��>��M�l3�'K�e�I�/�W/���(��g��
C[,�}�,���u�hMg�z�����}�:_�m-IXUϮP��vu��<�_|���9ç�7���,�ܜ�� ��R�RK�usa�N;<��l�{�N������W Z��-�N��L+'>/4ȶ�L����^6�b������Z����Ǔ���h�8QT��f: �ʰɶN9k��g'ʪM��(I�t_Z��Ѝ�_2��9���V 4� I� �&�I����8��������G�80�
���䘑�{؊9�J�%14���X��x�{���N�`�4Ö�(1B���ÊD�ѪS���ڏ�("�����@�EůVW�U;�Ƃ���S�e7���葃�L��ۨ�K��j��87)�۲oy�E��!�:�l��W��-�U��N�&�I6!���u�+T5X3���P�rf�������^{��'��	�1�W4�[�=�'�����j�~F?lZ��'����' U�"�=.`>�\���<�>z�<�z�W�ʐu�X�H��vgr�#�NȞ�@ ���6H~;y����Ⳛ�B�6R�G�����(�F'�L�����Cf��hC�ϫ�^J�������b��CL�kM�ڸ���q�	��S�<�q�l'P��.#zr������=
��Le8�ǯ�:��{ȣz7V�*�<�W��jz��ݵlzQ�[:�������z���X��(>��=B���x��V�*�� �Iw�Y�"���FѦ�D�;�5�vs�L�����<��˱	JE#ֱ�.Q?d+�/ͽ�w�I���	A�A�DaU���ħ�O��	OD݁f�GR�.��O�+3�c��%6�����~�%>
}݂qR�L�_M�0�'��5�qV	4o�^..�4�ɑH��X�<iz��(�h�x�D�ߥ�=��Y������C�@;P/�\�x�Z��bv3�!�B��1���s���MO���b[���Ro���H�x�Ӎ�h��xv�CՍ5��N�]v��ո�'�Ba1�����>?*�}&ujL=J[�+�Ȩ��$t�����}8]>�d��<�Q�Q�|��<�i�MD[m��3�1�J���;�{T�=�F�#���Vs�L�//�Ӗ;i���jl�n1���۱�B>t��P����+���&�e�a��!a�aR��M����u������S����e8��=�L�ٶ�C���±�K:�$+Ա��a���|eBB8�.Z�w!�%��ǝ�������jY�̈́s�{��n�o0s�:뷧KW��٭�Q�=m3(vY��,Ĳ����,4!�㮶Hh�J�_��	��6��FB��G��������&p���fr�:D[�ᑴLj��*=Q֟��J�=�m�n�����0G�$y�zG�_�j�0�����8��	b��(���!��⽾��f^�1�:��àE4\ʇ�n���|�R��bH�e`椡�?0��pK���f�:�E' ����~<2�v,x�W���;���ބ?V��P����bGE�r��N2G>�{�C�	B��bq�3�R�*bk�'���s����q��R���f=B3�~pP��s*� A�l�a����<ܟ��S͔�Y��Z�>�I�d5\�@�L��M�(ϻ��#�D ءO�{�#]�����Q�������ąLD��M
�T-�r��l(2��&��m��OM�j�6�6�fg�G
�9v|�Ƅ4�g[�(����]R<�<싽�N�w��]a��m~�<����������Ο�0yWm��m-��Cm��8솧�"؞�fl�m���8�[|6�����M��8��s�0������2ʊ*�˴��s�f,�*�Z�e1�ץ��^���-�w��'���=��S��B���Pࡹ��Hx���`�'~�Vur��\g;���
��P蜻����y�g�<��;���b\F���y�вu.ptO˒�AT5�b�<��a�/���+�6� ))��(�T�ĥoj�(n ۻ&��o�� ԝ�O���ۅެO$%.W����_Zk�+h]R�_��U�*o
���
��t.���`��ew ����5�T�,P��H���r?"�|@(X�xP�������_�s�/5ۘ���C:�k��`��Jc5�b� ��<�|��R�f���w��`Je+���:��d����I�/]s��u �
�&?�WI΁�!��ӣQ��ۓD[	�8�/6*�̴3V�ڐ��D�p�VK��le�X����X���?P��*����t#�O���w�p�y%KIq�▜g!�?&�7:����
�"ǮG���_�'�wb��l�'LZ>h��H��w��� �=�A���4�9]$�9�0�Xk$.��'h�`]�w��&%&˝�U|���z������E���*CR�_�|{~�l�?�L>G�eM^�n8��Ug-�+�v3��'�6�@ˀ~e�o��>HՔ� R\�{f^�'�v@�շ�AN�_�eD4m��Nˋ;��q���>k�����dҩFz��L�`u�!��,��9��'�.L�̀�#o���$�*�AM�e��W#x�p-�e�"Є�^56�?y�A!�2N��[���nHf�b��c�u�V�4OBL�պbCS&c�2je/��w.�,eެ%q/�O�O2[�.\���k�oo�*��DV�uE�K�|Ǟ�k�;՜�ĎzpU4�g��K��ih��TV������zV�n+��!��5҂�9`�b���Ś�>~	"w� 	��q-�ue�����4�st�D4߇4dy$	8W<�5ߑ���q�
g��y�O�K�Ie/�&������'gS�Um�FH�7f�9�6�� ��m�&�N�ݨi̜���� ��E��:$���pO�#���2z-����5��yA-��>g�����������;�ׯ������0�����۞�|U�ZI�2��lU��k�"q2!d�d��x���.��������.�e��R]�i���}�(�}�2w�D9pӜĘ+<7l����V�1k���{�mCo��+�uzkG��˞lT���cj9��������t+�Ħ�RlB��:&�o�>_"\��4����\,��!e�R�8AoM�ԗ"ߞ�����9��[K�x��4�ɐh���
'��q���{_�z�Me3¡��H[s727�W��V߷\�6��M�q�&��r
}�����܂��s�1�����{g�۸Iq�SNw�E�l�s���C$q���w�F��U��#ٷÖ'�����i��� H�W�����L�,O�&y�dZB�U�;�쓋F�{NY	gx3k���w�V�l�Rw+*#s��0�%��>��d�oy���D=����A�w��&K�Z�4'�0@�~8
��J��)~�fO�a�U���<�᱆+C����>D$�R2�k�%�� �T<�?�9��=����F�c�h�>XS�]͙(bUй�"�g�YO �A��
L�v���_�~�իx2bܰ���5�B�o9s���`������15�D��߭�����W���\{9�0RΊX�ͬ�������Եd����T��QiRs�#�k���33tf��h8��:�D�+|?��� ��:G��cZ���:�"q�Ɩ_rl���ؼؤ������e����D�6�S-4>Y���h�լVB���#/Ԃt�a�u>�����h^��V}����`\k �����2�V W�-Z�8�_hO����=a4r.ȿ���0Y9u��hrM�v�}oU�ҞE+�ġ'M���r/�$��9b������ޞ��;3.��� f%(|���;��n�w{Z)�8��ŵ�T�1|�0/`IEeŶr�"��̹z%m�r9�RڙMH�|��eN�\���Ci�.��r��pw<�?������"�ϩ]u��fظ�y#n����l�I��8�	=�<tl�p�����%m{��y����,K��F�����嫻_�=?�0����]o�
�/楇�m^�}�L�p��
�����������ѱ�{����G&5��A=R5�R)9U*�Ud��T0�I�nI�u�3Ҫ%T
�et_x��5�v�2p��	q��nf������d��hd����g����o�M�5"�!}­q(��=4jk�]���9�E�G�OAЅ����(�$ƀ�Nc{k!7ihP%V�>���n�������hv4���W�D��:�5ԺI��%|gD��-o�ӄ��rқE�uP��E�#-�x�����37F+��i;#a���M�.�[��]��<�A;�����5��P��`��Ǡ��J
%}݆wV.�ׄ����\R��I-���YKC�XL}N`�)�:�]Ba���R�s�`��?{���h������M��-��WJ�{���8w��&��"�r1Zə'�c����a_��-@�l`�C���a�dH����`t�'�qC<���PIP��h^�ƤD�:�dr�։M7$*�iK�"X��S�W��x$��O��)E�]D���A&�<���>՗U�)���Q����3��3su��<K�ք��d��o�і������x���c���fG۫PӤ��Dd� ��!*Ӏ
��pǬfq�iN� ��8�ΌÀI�v���e��vW�&��8:gv���7�z��KV���7H*�2����a�B�HA�:t�"9cWs�0wJ�������а2�õ��ycYv2*%�1��lg-��;�P�ЇH�ُ�f���+n~W�V�F��;鬏��H�='����(������}��7����WniT��b^���| ���L��Eܞ��K��Q���Ԥ�����	RNs_��ŧ�^�{`����+�j��>��8=yxK�����dx}��1�}hɈH��$�7���/B���AM]�P�&Ϳ��9ru�?��j
b�)�	E�sm��
d�M5���Z�q=�<�ʸ�B�[��uɧ����+��(Ɨvf�k]M	�cJ�v忮�B������Gg���p��+� ���B*Gɵ[����ʯΆ�a�'S�������_�^*�K\P)� �Tqu2�V�r��2��R�eB�\� � �:�I�z�a��W�<�sԱ"Z��@��{M�5�Ay)�C%9� \�@��qE�����0�%�$�\�/��A���)��L�u���cyd��ިa*v�2�ک-�s�B+k���6nX�Nl�k���(�hg�$k�q�SIɜ��P��ݚ��[TR�<~f�m��,0ԉL�1�_�Ū�����h��-�7Y�c�!���؎E�ma�N֡��gMP�
�R܎>�o�5|ַ�Փ�w�@���y&���d���U��i:	e[^keX/gs�0�w{V�SR몕���t��	뎙Oc���|�d�<�K@:��ܡ����^l'��c�%WG�r^-_:+J��@ ��0a�\��Ɠ�܋�z�h�}�����T����wN�̋º���P�^K7	;�	�Ct�/���<���2��{s^NI��Y�C}��z�wor6{�:Q�Z�|-��gY��L\JpS�<]CY�����R��RHY�n�n�i#>EZO���]�p䱏���a��N�3~�'�K�M}�k�C���qa���s���*��2G��`���VN^��s��#�z+��_�(G��}.G2k��09��t�k]��H�~��I:�A�Bx?d�N���׷�����;I�٭T��Cc�ا�����Fo�Y�Q����,�$�[�}��/���)���z ���]z�֥6��3w��c�tM cĖѳ���m������Qp��5�_��b��G5��{7��<�F�`x��w��7��&�/弑���S�;�=���eK�N�5�j��3�
%́M��Eګϖ�����j�eBəLq��H��/{v ҙ���r���2�q2�ɑ^����B���f��������̤N�/�T��J)g$�,��[��gw��QSn퍙��j�d�a]k�Z������-ʕa6�0ʹB?�L@����@�<�ɾ���c���P��
���Q}T���U�MO��pI5�k ����/�������kWYɍF�������{���;��5�J���QȓB�n�H;̸�YC�J�Z�����n�;0���:e{S�=#�bg��*������2B�^S&�����kQ�D�b�+�����Wվ�KxϹC%v�MYIw�-l>�F�Fo�k�mڠ�P\�$
:�мiP`t�H���U��Z�Ե�#��.3�sPJ�[Ie�M$���(@));	�4�z�ϋx����E��q (�H�.��M���vU�Ņ��e��A�aA�+k)�J�[��RU2ٚ�.���/9�/)�A�o:ݪ�L���ֲ���4���/Q�<���/��_̹�ɪ�c#�JV2�u>�ʸ�9M�0���4Q����ض7��!ϴ����Q�h.�
ysg����a�OW|�ͷj�`�c_B��kxϳ�}xAb����8�v$��{���Le�ϧ}�f�'=õ�|V\�^�H��b��毶-�٤ ����=޽�!=>��E͉2��{B���3��=����5z{�&�.�:|c�'�����������t���<��r�݊�eH4�׺FJ���#���8��Q���q�L'e��2/8�#�D��-�dS]O ͏���نL<uQ�=Y��hί�dP�UTp���	ٯ�$��@	��X,�2�6�@�P.X��������}��(��r��.@L��E5d���/ăؽ�{'r�z\��O�?p�JTCbfzJ��WiL�)�{"�/���Ӻ��T�fP8>y�[TnO;��ut�������t�!����KJ�è"��Ji�]�7��*�^���C/��S6����Q(� e
�[ ��E�j3�ܴ����^RI������y�&�s�Lmi�������ş�8�ȏ����H�q�$�!�`]��8����c���
O��GLEJV-�Rp^��)�ӫ~�FjI�.M��<mQ���~](3w��
A���x�cq��a�<%�{B�OC��=HOv�Fq�S5byA�����􏳞	gae�G��O�<뼬���ǩ�ry-�<����aSm�C���X�zI<����if*�@�-�X���ZA��M^�
4�ۧ��ݭ��f�y�w�[	�lJ����9FQg
���f�~�ɖ/z���g50J�T�8u��>[ݹ��H��;O������lj<�ץRz��u��դuV�i�pV���>����qIJ�����d�|�FF��Y�U[�,	��Gp��=�QJ��e֘V��6�8.��%W�N	3V_),�Ӎۤ�I͝J�(*��@uS���(���V�4�E~�b(�~��M�r�:K���Sby�XM�.ٙ���+x����f|J��Q�� bw�>��������P�f�)3��U,jJ�QX�rJ�	� �]/gP����ԧ8`�39�����^�u�a�6�	֡H�柺���9LS�w#��B���P���h��qT�tDh�4Z8:1@� G"�$�e�rCG��	E���������,*;QA�j�3');W��Bf�F<?ci��GCA��U;&!���W��Fצ2��� ��Yb�h���ŚƉ�����H�CfZ���$E����x�ݑ��:�`1�$v��c����Q���f�����~��������\vO���@����E���
,��º�I��b�,j�h1t4�d����!F9^��*�C���8B@������M�fњ�����,����b�2n�p�m�rCYP��q�TcHhn,�"��6o`*�z�-k0;?�u���D1���Hȍ�rj�,�.�,C#�A?AkC���Ȭa	����3���������,��B�81��)a���d��q�<����ep�����)�������#b9R+����9���2:`�f�ř��Wx�8W�TGE��N�5����4G#��I^o�
1f��D�[dC�!���ž2�R����������'+�0����F��P�" ���M���d�8,�A�������x�B2^�X���i
8�%�Ē��U��b��B�R���%�m�0��=�P�OWN� �X#�]P����s�"��+%��PR�Qy@
�R���p�@*��@*�K U�� iK@i�*�U.<���^^F
`F/0��4��� �����@h!' �K� ���h�D)��QP_��F��B� ��N�g�h 3� @,�AC?-�_�t��'��I��}f��'�|5��)囷�P) � K %��%� 	�r ���N '@��;.d�{n���
��F��g;�p~}�#�w-ʚ�B�������H��Ln �'��#��w�����8�]p3�ЅVY���?����	O{�F�,M�lo�!�}��Sպ"'��ή������ͻ�j���HZ�*��>/E�	�r����a
&��n�J�s��Rw��LLu31¡�������C��{���5h�u��y�;(ꌸ�X���y`ܧ0ؓ��V(t��M��3]��1�A�W#�231X]��;���1�X]aܑa���HO��TЎD>0D2C~8��9�z^�����oO(�y�J)9�WCb�u��;�+�1�
ђ,�_�6n\c�e�d�ҿ{ۨ�J�E>������ǟ{r�3�[�[���}����{��I��K*���"4{��?�`��򵌮�߽H!?�:�I^���?Y!��v~�ʈ��_+)xK�3��d��YjQ(P��pl�ַ��b�<���������t�+���>�gx���+&�;�_�d9�^�f�a�䊺dy�wY+�J	��n�0v�@i2��j��y�\ d��v9>���{�<�}8 ���:�w��-=Ws���к�pJ�6�Z��z�~f�%r�/��8���;n�d���Pގ��;����Q^i��Ӭ,���Ze4LOL�	E��'��T�4h�6-�Wϣu_[Ғ8�[�C��/S��-k$�˦Ja�5���%j���y��h�Q�������3\��t����u"�;'!��4F��&����o!�Ew"*�_j�+e�(�<=/����o�[�C�D�rfR��!N��s%R�f�2F�W�W̔GCa8�X��9���j��^cã�׳�m� P�ٮ�m3��L#�Y+��!�8��[��,���������,IZ\v5bP#���~8S��3엂t ��N�|2����
�2Թ�̘�����ZJȎT����O(db���k�fE�3��JvȻ���mY*3@~�(���K��ds���Y��d�?	�L�G/�uRV�
X����9#���~[�ZZ��ԯ¦��	J�6Yj��2#�Qg��Ծ��h��G������^LP&o���E�nmZ����Y~|�/���	���F�-3$��Q�����Z�w�o�ۃ���@��U��~P���L~2�K�G��&��VaToN��'>�`7�k�#����0Pq�U�%�^K�Y�t�6i\-���Z<GJ���Q"�ġx@�	ŀ#���	�ڣ?���F(1�H-/�.U��o+�	�@���ht}2�CPz�s׏P'ϏF�I��ZJ�V�.��"Ȟ#��e�<	�_�gӫ�v�f�ӷ���.�]&�w�Jwf��gj�\<�IS���gx���3�M���1m�y^�!�0>n�7�ϛ�)�82����\��ߘz�r(�D�<J���׿�߰:�_����~��hŬ'�/�Ì4R/�MIf��/9���u�D���������w2X��O����0���׭|Q��S���w�O:T��v��h֜��)w�=�+�!�3ٮ�1,6wd4�6�e���q*����T�j���r���~A"5�m�?AL��Ӆ�T������+XC5A|�КV�h6��]9zN��s� U��I�; �-�l�e5&tKe'�X����~��vl �]`v�(5�X�V�����# ��1>߆��I�h�Uv0`1�6�`����i��@mZK�	����k��5M��#���vaM���Mi��:�&�v+��4bt��<���Z����P��"'���|�!�i��X���ҦYc�"Ů��J�R���v;_էR�j�j����Hc�� Gi�D�ŵ��H�ct��3,��3��r��W��<����۷�6��=��f������a[��-����߯/�tgѰj� [:P7&���g���q�,+pb}��2�.�y�^Д�)ԍ��g��D!,�]�	�~uj��{g��6�e�r0��<^T��e��ʶ8��?��*R��b�V��{WR�P'���w���T�[
���F��~�ҚI-�[!@z	DQ ����$��@j�����Tpm�����%�5/�=����,j ww
�S��L���J/�Z��%:&Ii�^?R��%N���qIJ+7��
�L��;�!3;r
�Ў��nx��o0׊ ؝�MI�ݚ���C���f@�5��WF����5��{d���A����$ϙ�s�|�vR�+�9��5��N\CV#�'���+ȃ
�J�៓�O�{��Bg����k1��k�. ��R��0Ӝ/fDOs+^�[魸��o�˶?٨S�K3v��s�(��å-���6�QӀsL����'�ǈ�%����X�%�In�$�EM�Y�������Q/[K�%�t<Sa��q��+��VWT�>܊4}���Q� ��3��wx�{bt	�֘_pᢍ����s���g���+i�F�r��2��c�Eo�]L����0��¿�<�q'(�C,��hUTy[���T��GbL��%i䷆�G����V_(��gyH��,�,���׼�w���Z&�A8Ax<T��q��S�R��a��6$�w3��������3��p�,m�r���o��tL���#3���9���nl#<V����k�u+L���m�22PI��Zϰc?0��p��D}uPp��$	������שW���d*ɔ4zLL��$�[S��I��k0�)ϠԧS`�Sة�(�츪;p�� ��p6QnYQI��E))�3]M�����_��)�8����z
�o�t<,��Ԣظ�:t:[e��K�.�K\���GC����Jí�Q�2��F,�ꩠ�tV(�*+�m,�)+��TҪ�~�V��	'k`ЗN^���'��Z�CߍaS���9n]��)�+˱����4ˁ�c��{g!ʧ]��pi�8V���ީAP0�HWd���5%z�i��\H�$)��-�mz���s.�m��⻬M3�ʜ��N�2 ��&���v�y�զ�JY�t�2!�}z;5h[�{��1>�x�8凎A�ǂҲ����d�WV���I����\#%		�חx�#=���O{���V!ў�%���r���l���e�����9�4��w{wM9�ѥj,o�%��&3�V!*Q<����fGY��Qᴪř����]��t�ῢ_�]�)L9-��@ $������G
�B�l��y��mT�j�V���SU5eN`�T����fQU9Y+9��j,��c��Iv���.�(B[*��_N���01�v�(� ��+������~^�9[<j�~�A�� �L��:�/�/�����4?gL�*"���l氽|�)�X�ԭ����}w)�4�=���T[����Lx�������ʸ�g�8�,���PJ���n���k!��`����n�E�x�GIr���p�_������m?/=����:�C��<���O��B�.��F�J��ƽs�z���6*zH9Ab@�"l���ڄ�Г�*����P���4�v��Ȥϊ��l<`�����7F�覞W��I���%��-����<�!�UpdB7H��/N!��w]�Q��}��_ '�@���PK!�l=��w�������bhA�!�!�W�BRZ��l��|�~M�n«۸�W:&�ۼL��yޖ�ȁG��I����F�l#Tܞ�Senǡ%iL�h�O�V�	��q�$�5�Xz_@Nb�)��Ǫ�*�ρ��]��N
��u�`�k�g�rծ�bT�
��(���*G�����Zy��f�p��cx;�8�o}���[7��`b���C#�F�ϕ3�Q����:��g�+�䳹Y�F�wۙ[��[W�FQd<.�&�H����tcG�xj�
n�&�0��ъj&�K�W�$E���b��0��M�{���Fn:ka[{W*�qǝ��/�ݽ��=(�j
���3v��;�-yACj��s��2�!�;��6^*ow����z��iC���(���2j�{��S(�춁�0E�*���{��pyG[�Z����.tf���<��T9 �a����~<���w�f�@Vx�
���=1&#|�;M1x�f���es8se��N�xN���ӫ΂������m$c������؈1�+ �3�>��;:��_����"������A������U�>|�/ݬ�h	6�n����cOۦ�q�1��Jd�Mu�	�L^A�F8��H��a� X-/��+rB��awa���$W�c��ل�j�sW��y��	����]�4(sa O!���&�sREY�!.�n2;%7��V _����<*��ň4�`�bg����&��+8�8�|]�Jū��	�`�"��I���^�L=�26R=ھh�.ɮ�	�4��H��`-��	Kk]D�������ǵ~n��%�?��-m'�����vl2�ڳM<_:h$� 0�u�w��,?��t��b{�[_���f�1�'h�^���N� YB�	򵟂_�f�Ow��87u�s/�+�a�j~�2x2d(�OwVr�3�[��dzv)�dm�J�b�F���b-eԚ`i�!,��6<��l�y��K/`�&�ρF�ԸՎI�[h�b��{��������O�./��ɾڸ55�Vk����H&��<W/}��Ch���hZ��h�O��>)?*�M�u?��+�~���؆6g��y���A�S-r)��ݗ!�θ �N��>Q��2Ж�4l�Dt�!V���d���kt2}0�3��s��3�%�-납5�2���e���H����i��I�}T=�P��6��1��$]�RKUD�P�6c���G>Ew�d�EI�^��Һh<� �������/8 ���d��SQ��s�����*0�>E�D4[��:TD�;-��1ny�nG�+��^�Q6b'�a�;Zl`�,�h.��O��吓����]teF���n1��!�i�w�l�������̑�h����"�;����KJX����f鳴���P��lc݊��6Қm�z����c~4�)�:eR��΃l�Z(�I�`���l#�F�;�.��i��< �T�v�s�j&�EC��c����{-�5��qt���z�@�r���{�4��,'���g�8R�t-0�3>%>�����q��'�5?-ބw��0;q�7�'��#���H��I��h� �FYh��	|�w��h���<��B%8P��������lJ��kl�����DO5�OB9!/d�(�����F��60�����zst�D��.U{"$)t�|�)F�wԙ���
�e2��w��$d�ֽ��G�p�EѨ��%܄U`�&$�����4H�����i��v��ؐ1C5�L���8>�?ڎ�|Ә����ޅ<�y�������Xk4��,gZdmO�5_��ג9�jf���(�?�[_��MZ|_�&�Q�*>�e�}��Kyg}��~�ჾ��n��T��bk<�K�4�>R����1�����`����T�����:�@�{����Y|���͌���=�6 Cg�L�
������\�}[�,*���溝�i�c�f�*�$��ak���V�$)��u�e�����kS�d��^]���w��-7k��@�������1��(��?�Y;�����B�ͱ�Ӵ������P�ܥ�q701g��@MA���Ts/髜��w	�o��-{�.װ��is�VStJ���$���øQ(�o��؍��b�L�����'O�����;t�+�_���Ċ.2R�$�y�8���#ͦB���	�R9M�UU?�C���ߍ�^Z�/��m�7�������bH%�TI3{"�������M)�������n�o,AK�;ٲj�sq1{��Gyf�p�7ψ�a�G���2�q��<��)O�r����jk�sP�bf�Nx�iB��ԛ	�!<� 0��nK	���*_�*vFZ�P�P�*��a�=��#�^ǫ�iছ3�� �$���T���Zx��vx�W�]@�kCɝ�ǵN���}C�sT̑�����������ǬĆP?�|�2���r��wy��F���$�I�b����s��
����$z[��3��_��s���W8�eobҭ��Ac`t(w! �j�Ȗz?`=]�
a�Jr"�B�*6��kd'_�dH�s���2���l����Y �/�8�R�A���u�E��>1^ೈy-��CIL�4�K�g[����T��fo���q�{����1��$��K��3��H�5�T�[X�ͦT��c�`�YA���4����Q����o$��t�m���{�h�����'�i��ޱT����-Lx�9K���"����]v]�@�+8�	H1�g����F�N�w�-�N�pA,j�(>��u������:
�&F�]3&�R��FBI�%�^R����Z���u���IY	o���),���Ѩ�T��_���k�}��2�� !<A@^���B��ca�H0r��*h�������m��b��v������5��ԯ�r�jAeR�r�b�wcR)$�GPѳ��G*V!��Q�P�G r��Z**�r\G�0�4�%/�IsIO�y7�Iqa{nco��m���h�0�lP`��k��, e����>Ќ/���٭�"7�AK���e��]W��R�@%G�$��*�.g7�l6m#�8��#�ͨ]�5?�b	��_V�u�����3�Rnߵ|�$��^��h�4:��hڵ�Ĕ���X<�P�	�A�'iAT�1�����T�F�ݙ�X(�Ì0.���b5�O�J�孂�d|A�����{
T��.Ka0��hC��#{Q�2\^�ͻ�m�AkjF�2:����k3v-��s1�n�D. _E��E��G\ˀ����3��q���V�	���Rx���NRݽ��1\3nm����cj��G5>4���4�\����TӴ�Il�b�g��̑��[L��ͳ6��s3<g�n�����<���yg�_�73��������M�hlq�{3�M�DK$Re^�I9�և��������3Ɣ�Ži�
c�n��M���i�4x*xbn�o�Q��u�>�?��S�\@���j�����ޗ?;�BY٧�".a|�vwV�ZU~�=4�=M��ä�_��V�%�_Z��+f��9
ŏ�]2�����n�H���t��n��FR�zY!���G;c�EuJ9v�)>]�;0P�,|ykɹh��q�WЯ}�Z�~M�NTX� �L�m�!��Q��_������M��&A�;��(���x���1գgǦ��ܜ1sN}*��C��hĳ&f���\��C��l2��F���z�܂������E���I��Hͅ�(JF!dx'�E�������X?������)�t56 -��?4��T�I%�pcQ;�tl�����#�e��0'�.��9�~�vr�.�+�I�ȲB��R%a�BIR" 'u���x�y's�Ό$��E�_"��"4wJ/�?TՉ?�i��Iu�d��d�(ӸVb�J�HZ�*��.~�G��/]j��:��H�ˍ+EH��'�8:�#�H��4TZ�E>�R�(P"b���S�#���Z,�mN�tri�C�r��8\���xS�,���'�F)�)F@Z.��@��F%��u)h�bC��o<�X9���J��e#��"�Z.S� 4]/Q)�W}'�����?z >�?�c	��]�j�]�NezC��&�c<�b�e!c����tp��o'7vY����&�<RO�uf�e�in�!��4X���|�]���h�'��y�	0SyC44(${�oy�"��M��$�������oʸ�o�# <K��f���)k�'�y��rh�3K6��>X���r��&_J֩�4�ھ�����XK������";���G+�ѫѿ+����K��U�O�4��0���5�Q�!�k��b�,mE�e�L؈�i����l1��maR@�խǊM���N?g���|���!�t��3������������Z`�()���� s{բ$�
S���^2h�e��˄�`l�2|�b�/d
Z�g H}:��1��_i�?T>�i��m*fH��+�AT�x��ŉ�'�~�����!n{8uD3�P�^�}�k;al���,�h��-��̓���f�cr�:��`t�h;-���
f������:<�k����b���p�c�����H��W �9.�k��76���˛�������M���/�3����ab�����vgY���k���B�^��	�Ĳ3� q���te�w_��n 6��MѨ�,׳�Z�����'GG�qa��Ai?���f��^���)��iYBO�x�x/Ʌ �u���>��P%��Ha��U��}��)����x�*r>���n#"���N5�2FUV����&�K�F���~��
&��T!\ә2W�͑�>�� � ��S��X��4"��(����a>q�z��\s���ðK��}?���]�����m%s(�gѝ�Kj��`�;nв�^�;��S\���%F����m�Nx�vp,�%I̓�fY��(Zkm٧�B���Y|^?�ē"��TYi�.X5A���t��@_=ǆ�Bϒ�ۄ�@s}-D*��CE`U�����+vp�b赜�X�&��\d�U���������,9��8�9���Z���k39,� <�2=�f/櫽����-�~�Q����2���k�GȺ�o�k��M�C�g	4[0�й@�HM)aR�
�d��ӑ�b�5~�����б�髡VL��>�б�be��7l�ͧ�Ksߞ��3�����8w�y���4_�h��G�f{t�1��[�+�������l��n��=I��V烒@�k��.+V��2�騗ڛEҀa������]�R%<�Up�vx��VpmE���x��H� tX��H���%�����q.�Ȗs��V�b}9�Ug�ù}'_q�0��}�p)S'4�
(t<l����RQp:-TM��%4!L'���A���ւ���	�!�q�)Gq\�9�O�
�:L��C*��QH�C3�
��':�-AsdÓ�Žj��.q�Q�*��MQ��U�c��)�7��R�b��-tn�?�է�MV���N�r��'8l�r�� .s�Q񸫖��`|�S]=�����J�ا�^�k�7�&N�EY������u�^��B�.JL�qq�>L��z���v�Z�]Y�j�Rk��c���O}
���H΂&˗
,iNL�6��8��;�<��Y���z����C�*�⩩�ee�{Q���W�"f]6j��Xzq����\8[��{�"y��1���iL���Ĉ��
J[��������Y��1�G&̻��X�������XfM�%�m��s)g{��w����&��־�>%����^qr�O�w��n>c6��&�m���P;�8{�@����w��@�\c#�;兟#y�,�|E8����$��C��}?�R{6�X~��EI�%h��E.8^�8��{��8����9/4I��賕��!�k�I�MHOG���A���<��ۃ5@n;�5��"�h99��z��T8�Z�����U׋>������Ɓ�a���:�p�m��շ|aʢ`�Gn��4��x�_���!�_V�D�c���([��]J����ZE�D�RB����Φ٪#^�k�ᵽ*g��u�Bf|���$5�7�|�?&�,0+|6��r;�	�3�$-�� �C �01�|��*:�m!�pHd��V�]��e��$]y�aa�n\#1�e=@����4�^M_!N��S"���Gg�Cs?d)Xv���ug���p;:NX�B�k���T`O'���FM �U%=!{��Mx9���g���<�U��}\A G�Kѷ�8��3���xd�U�b��W�t�6"�[����Jƒ�#敊��!�h�n"���j�ϡ�������Dl2	TM'�Cg��\��ྥ��?3|��!�Ѭ虸R.Q��y�g�4K���8�@�n��|\d1��f���Yg(�G��L��Ǌg�yzs� �c�bAZ�����qA�6�#��<��Sڿr�o���1W�ϗ�<\��NQ���>��1Ϡ#�~�K�;V&k�^J�AB!&d�����y��`��oɗ��X��~'iӯ{�l`�E��� ���!xG�}�XK�%�����XxJ�o^�e�3e����c��j�?�28�� �M�1n��+q��O]��+��Ի殲�DWW���(�>��4�z�fn��lm���*���ɲhv#�R;�=t�*�͠?�c:V�b���"h����~���8�7�]Ŀ"���M~���[#��D)Q�������[+��.n63�t�X�}Y�+U�����%�F��*���+�!�>'�X&�}���A��$nJm(����[ y�NQ����S%>��a_�SN+�2XyR��;B��5�v��7��B�����4�W��č�3�^�h��5~�yiY�}��]�D��Ul�p�/ww�yy��X�V�j��IՆ�5^ȥ�>4�_^T�"�2aATX�Y��O/�H�e��Nm�SWFt>��~ww��T��ƅW½$���}���]�W�?F�_��o�l[����
��h������өl^ob���%+1_.�q�i��p��hZƒ���Ũϕ(/n_x���7�G��Ι��ӥi9��,#��kb�&����PhLd_���L9��ǃ0"E��e�����Qĉdm�^�UR��|������X�Y|jbͽ�$��X����҅y8Z�'�<5�WTW�*��_T�!��$�Fq ��#��_��?��m0'd�h��d�&�y.3�V����V�ֶL5HU�->@�9���Jv'j�pf���u&���Q4ƴ�#*����+��x=�Zޔ���z\/P�!����6i#��D��gω+QJ��]�����ΰ�0�☥mK�B�E���,Bu������\�Kd�UI>�L�9�Q�Ss>�%�T��u�E��eP�t�7��,=r���h5���A���=u2K���À�H�f�h�l�og���l_������%@��G�D:H��?��vU�䙃����tv��ʋ>f�h��K�ҟ���R�/� ҃JpP� �s�\x/���;~�JB1)��ݩ�n�BH�m���n!:EX��
�	�?vO3����C���V`�Ým5	�dQ,�V�Nd�㖛W��4ɴ��}�*h�9�a{ L���,��>G>A���K���)�g��y|.�d�B?�$p)��l�L�&g� ���	���+�TE$QMf`Р9N�.,���c�(`	F�_屘 fBy5/�>4뻊�D�7}1��q�F���πH�.S;{Ӊ~E�΁�>zg�I�UaG(�3� ��C;���`���7�� ��1pIK��/2=)�f��62@���z���&����\�[ \��
�Z;�:�O�w��QH��ʗ�Rk��(�7!X9�E�]	N��*W��)A~8Ц2�),�X"9�+����������5csS�;l���h�?Х%��� Y�nlj�沋uh4�E6|#�
4iYm�C�u(�R��<�l{�A�К����(����<��q�I!~�VU+C_b8���Ɂ��l�s�´6Y����(�5mŌ
^a��)yS9�3:���xP5��ώjs%�֕��S5�Ź�����1��/)��Xm�J4~�j�5;��,�Z�x֚��,�]-�'][Sr��I
.�	��� �:)Ī"�]���9#0.��]��f�	���W'�H�8��uH ;A@.LԐ1��,+螆���^da5^����i����r�.SY�B��-wo��YK̂|�2��
)y��b)y�,, ��3�M�%��1K�{30c��^[���8�Od45��́�n@��I�����\H� f�	�@�d������(��b��,��@�;���;)��?<Z�}qpbx@
^eo5ށ��,�� y�D�xπ�//+� ��v�O"�Sz�_�ꔠ�reW@fⴔ�KV���`��,Z��1_f�ծ���L���+�%����}���;G!#j�5���'�v��2P�B���2��u�O&m�* ��@U�(� �x� ܖ +J����(
4aJre�]����Jf=#���*@kw���ds�p��݆��큳[ɿ�g�i5YT ���!�����@��-���'#e����&��3U�$�����2��	��F2���� :�dLJ�5B.G�s�zO"�Sָ�E[U�7%x�F%2��^.#H1?Gt[�ڱ�M38Ȓ)������x��ـU�8U� ����4R?�́�1��3q���h�P9;�~!�ݚ��{�2���8C��a�� �9q����� �΁Ѝץ�J�S�겥!�����ϕ;U3|�9Y-�����
��G��풱��1��@߳�J�a�ҿ�Li]��[k�Ҟ���<'�kǍ"���C�Ӿ��oߒ`[$Y&6[�,v0�t
���7�A��|�*���h�+�TlA��jpZ4�x��:[���~JE��5ур��J�d�ɀ����v���"I+�۞�f�N.Xmm���*�C**��d�/i�-���)i��i4p�p5?��+0��;MBg;��b��Y��aR2C$��`�q�yb3rF��nK2f6YE5	��R���|�K�V�CFIjW�e4�q����ŏ�r�>ie��e�|6U�&F�5,,�@LU����.|�(uv��\�r6���ωEDГ�7M��Y�mW"Z<ujA�@O�m/^�y/��V�q�AF	��~3���v���Q4%�U]``r�M*B��ʀc��p������Κ'D~��VB��	~��$I[P���[�<�g�$�vj����'�mp4�`c��%'O�\6`�ϊ�
���IX�[U�
 3�4[G�3h�� h�l��ӻ F�5vJD��j6��[���*4>6>8�T	�K�؞]Ϫ��7c1P�H8z�d��'��$�{��+d������2F,(�;yn�w�cJBW�n�b���7K?+�c�2�*X�t����嘰Y�̈́�fi��
�&{X"OɭV����?��KS��t�t���U�~(���TA�\$O8�>γ �ݕ���|����Գ7_�"�8Qy�]�x�\˿� ��X�����\�U�>�#�G��F�6�YE"�w�[��"7�]f
���Qd}��Q	�n���
�q���Y94ja	^�,��^M��fd�Vg�i2�h�:~z,��9_e�XW�D!{�ՙ�X?Z��>����E��͡�/ij�nMڰ����^i�VF���]>�͗���D�!�Of�r"uEhSNuP�ص`���|�F�C����[o�vE]��n	�ݠ��w�T�x�d̝��p���a $��7I<� ��6�h�?'�\�`��{n�Z�Վ�t�\.O*��[f�,{�R%[�x�4�ۓ'X�^�O�2��E�%AvJP��d8@$@� H�"�� ���ʛ��˯�/M��)�	��<���NU�BS����/� )5b%��)��D@B��K��Ǡ��Ȱ�x�4�d;�����e�
^˪Gv���{?D ���g�_�%���1Fn�|�!�t0>�ɑ���]/��^�AҬ)�"%2/�U��[���Л)wT=o,.˽� EB_n�]� �K^r2�K��l�2�<9���8�%L劤���ꖃ8�݈�"*	ZH����e/4�� �ϐ���F��j���Or@�hz5P���3�G9��u��

���ɜ�(��v�hK��T�+��;B�F��3�P���\/�_5���V����a�3||	ʵ��hKk�׾>)F7��fRy��},��C�����v�ZvY1!�N� ���Ee�@�(e�L���j�!#?�u��pփ�'�x�ʌ�hA3�9�=jyt�nT%�e�xe�qX?��Ji�aĢZy����S]Დ���d8����#*UzL交��'|K��"dC�R��b�i�eY�6��P1yvM����w��]��1	����+������Jv���o6��o_����&��X� 'r�Q�����a��t��*c�uW������������Ŭ.g[�|ސ�U�a��v�x�^%�l�a�
���,�v����Pz?I֭b<ɜ�B��`��	�˽�Q���+���wF\Kܼ�\Ip����ퟫ��ˑ2��WHS�+��KYA1Y9�h��+h��`��(h���T
�̃��x��ܨgU;��wIWL�P�l��Cged%v;�Ϻ���{G�p�z�W��{Z����xn��/���}I����H��T���*�e���І���!oF��my�qm���KX��C���_ ��y�'�]Tx?��|��F�!�RS�Е���H
�YJ1z%*F���9S��U�Ep��Zj0?|Vf@���h�u��ݙ.|����IozY2b�����>�0������w}8+z|O�����r.��ka^�Ftcu i]K��R#e!:�51�ȣ��\7U?'@k$��!�m�	w��J���?Z���j�Ex=u��j�qX�۳�ڨ����*��G�==M�
�G��uQf����[��9/=a�ȅ�$����I�wM��z��w���w�O�U� �B�_Wͯ�3/_��^�Lh��R�u=��P�$ �/U���|K8ԙ����e�� �A�,)E��V�*�	~��K�8� �v���0>��}��8H���ʂ� �:����&��9�@rK�[�X��HhG�a�z�|[z�	���(�75{?�d����xVh��ML��vM�8?�]!{�<��\+����a :���
���"��M�GQ n<F�.Ǹ�Lk��s�OYh
��Ҏ����᧍xCM�Њᛣ*=Z7y��V�e�D��}/�W�0̥hYקbz��h�haX���ׯ�Cw%�N�f���q'MiE��˼����;�Ur�r-��l��;��	N�]aW��d3�9}}ߤ��X��GpOJ�l�Ж��
���%}���N��#{�T�_�г���o�S;��!ۦ8�Rs�����BS��eH�jn7��a���	ҷ��iG�l �r{�͞Q�;�gz�r?��O�=8m$=���cwN���Ry���y,H�����2hB4�o�|�ӱ��;�C5�����z�P`3A���^�|�. #P������\ZO��;�Ց��S_+�Z���kY4w��d4��U����X!�"�c���@���Fs�]�j0UT%��&��׫`[����|
������1 ��d[UW'���5�@Z�=	�O^�+МfZ��R	���0�v��c�E-G� �T*�:m��#���h�d�۟�������!�m��񵗃�%D�����B��A��#�W*omH*��ٟt}s�tL��:�g�T�������C�FO�r�)�R��ֿg-l��Y��V fj)�9����k�QR*�i�2��ғK�1f�,,'�K��o�Gm�	 �Y�}����2p莴B�+�׌�K�zV��s�i��H��E�`�C��Ǚ��W����r	X�j�/�U��Bj� ��������F"�~�ؕ���-O	Z����0lyi�������й�9��p�i#Ϗ�\Z�5!na/80C�Oj��$d��j����������7w	*6�84�b��u�/�*/
鳆b\cX3��m`�Ce<�t�]!|����	
jިYhze�j�og��Fϻ�YddB�f��걉����ĉ'Q����}D^t�B�:�O�+?+���@t�9h�6�8���#���YhG�p�]�˲pri*�$d��+�F}�y�7�6�)��%#���!DP�H���/���dd�$�
�����A��2�ФG�L�����u��e�YZ�M���Ҥ�zV����Ԓ���,$_6kg��O��(�3Ȕ�Â�τ:#�L���\�	�0;?T���� ���}����#�צ������!p/��K#|nU�ډ�I�*s���F��������]aD�ٲ�!�o�:w��G|�g�N�]�9��$�9��D��l������Џ�K���5�������E�)��;����*������Dp6�HC��G2+� R���D�_x��v^u���"0L���Wv�m��Q�$4!����aN��G�C���Ǵ�S�׾��f�����ژ"̚���E�XVD�u6�6$�c2�	\s��wBG�L�l~��0�U>~��a�y�AR���M1�!c��_��]/#���{6�;�ݾ��E��}��9�;���V�.,� Qe��,i��9��0�I���䫧�n��I�mUS^�}�rY���55(�FrqgA�T�}�L����'1;�u��ad+"z��M�u_[G���KS���%ڍ�B �� x^0#��d!Or�	J���Aնp9�� ����<i�xPR{R�M����B���?Xc�Q9�z����.�(��G?���~����'|e�\�*����]�_Ž��g��)���mzy]�dlZ?�TДdF �OsxG��D�H���L�X}�=o�]Y2dt�Ti��)����$*}7_���z�3�r��J�s��^������|885-�/��tJ��J�[}'�,�2���ҋ��/�9Ei���(y�X��JI^���P�.��3.J�-����QXtl��гU�'�ozr��%��\1��Y`ދy��Ҕ0^9_^�SS��4a�k�ǥl���?��lBR�Lj�fhP�얘�0���_���d�/X8��Q�szk�:qު���� ��\�U���t�UI;_���g�Uj�p�I�҆U+�߾�e�� `�~ު�<TZf�R��5vHLu���K6 jX7����2��lgQ��H힊�0`[A�P�t��@/�=y�4��d��&��hR����%�R��dƢa�g�U`SϠ�c��F�6�9�w7�®E:�E���{����i�Ea��E^6�	/�W]!�ԋ�NS�[�}�ll���"f���n�m<}9G�ɍ7ꁪn�ڣ�S�|�H�c�Q3(��z�A]��q�6�S��D9Q���������mI�5��ւ�ȱXBHNlLwu.y� �>6g��ڇ{�$S��{��(��H0J�Zh0�wi���n0��������!ԯy諊V譔���$s#�=o��J��:Fa�_	��?������a#����Nd��S��`�Z�;*�-�6Q.72����.�c�~���k�OKC�e�f��k��D�K{AdN�I��X�5���-�k���:ϑ9<q��)Y��X`��C����q���ݯL�µ�1J�7�.ONV������F}e��������Ġ����µ�z�g����s��?Y녗�����1�)�X��ć�mN��i���A��y1�[I�/���	���H��ۀ��^�C|g��3�-�B��a�t@����ϰ�ɦ�G!
�6�;Qֺ��U&v��5:�oZ����Z61c�|5���7L)應� �)���V��%V2pɌ2��j"$�.a/nY�'��g�'A��~����][�� �wL���#Q<nG��_�uBb��=r�b��P���3�g��ԍ��=����v�¥2��q�+(}W9�¼ȷ�#=���dB�
��f���[��vXs� �iC E��v�o���'�䂗`r�ϐj:j,��S�B�Nj���N�l��;8D�
×���R�޻��'�`�Ֆ�b
���k���΋6~A�*�p��䮒"��L��U��.oq���]}�I>�^��$�*8r�B¥.�~�鎷�	Q�B\�9����O�s�u�~������+�wr�1��֧��������G�?̷B�yg1
#Knɝ�.�k�O� �����S�*�_M��iIU"��&�g݌z���z�hφ�̌�l�jn�6�`y���5��<�p]^z��֕��b'#�᳣2"�\	ٙ
e5!�2��}=݄�؝�w�� ��`�����8i������txζ;n���s�4J�uو2$��7O��)V�5U�nh,�f��(��	��o> ��򫹜�Cؔ-q��ol��rjc�㻍D�P]���t*h*��	Qg�5T���4��}�>q㟃9ɮ ���!c�����M�����Q��D��e���ɽ&�N��/��(wr�K@�`���Ud���%��M��7od�����J�.���妷��E��K4���j���'p::���Zm|��9�-_/v��z@�Q�Z�͡h������{�rqqP��-�
+P���?B�\+��Ӵ5r��Cmnlnӣ�6�c�.����$/�ɋ9o)Բ: �ǵ��9jn��G>�:���ǽ�WR[�D�(��R�[���7a5XZ�e����5>7n�a�/+Է����]�������[�M�����c�o�Tz���*Te�Պ�̵��&�9
[�E�ەs]�����G��;��էBY��lgfk}?I����5�rL�7;R��}��ס�,H̭-����J6m�#�ɂ������Pӣ�-ZGTٓeiVrs�eǀ8�x��+��2pR���Y=	�,�?�w����h��ɍȷ��%�N�Ԯz��u;ڄ{��̠��!���v��8�*�89�ή�M'�t���7M14��:�����q0C�~��r"�-!���7����~�.$�#t���%E�ď}�/��{a�,=P�թ*����d��M���$��0=>��8B����l���+#��#�Umx2�#qO�$�jQ��Y3�G�&-11W�\Ƃ�z�}8c��}��Sw*_���S�ɵ���݁���^�\:(rs�����Hd� �7�с^���������mDa�6ɻRU]wP�0��f��\LT使:S�b[�&މ�f�R�z��5q�d�]A�P?,"z��Y"P?G�J�?1~5��剻�W�❢���I����Q<\�!���';E��~�_c�_�V˝��������M�<�H�NE��N�&���4H��g��PhO�A����"&+V����]	ڧ]֭K��<�f�i*tC�GR�K�=�5%Q����)�\�ӧ@�A�7ۧM�[f�梡[`+lc٢�@M�k��؊� ������=�Μn�(�*��z��q�L��S޶E�̊ѧ��������<(N\3C�wo4C�ʤ�*�' �Czo�h�����l��]�C_���ɷX<��{��a�7gB)�����6�CuQ0:Y�]e�]�~�'8}hM��1S1��a2����j4:��}Bv����~��ڦ�H_"�磯d��/Y�<P�`�����5^�$��=*��[W0�ۅ��H���0�m��1�Vu��9����R(���j�e�0
���a��YzM��~�#
����6�T�^Х�[Rl�~��O�H�R�f�u���ΞZ^s��H�AE@no��2Ť�j�C��׾��9��շ+���4��'M���p�|ܑ��N�i�z�Y����m=kj��E��&�{z���5Nnwѹ��,�c��_�(@�ٷ}������oR`���@�9���մ�����d�l�"w��{~���Cu�a�m�!c�kTqp���9���
����	�Ͻ�m(��:��;}m�H�D��u�����{p�J~G3�Jz㕣Q�o�����02{`�m(R��>�ÚU��Se�7��DU)��S)Ό�-�@�cE��\6i4��z�y�4�7K�sAK�X����nRgY���M��FDa�Y.Z.��.�N�-����҂d-����e�S4m�7�������A��_o��ɗ��݂7'�H�P��4G�CTQAґ0��ޭ�S��P�{N�%�Q�����d�`WY/軠uGN��H�R��RU-5{)���\�×[;�~�"Vi�5�-�����ث�>[�3�s\"}��م���jZ����Z���j\��1�o^��}�a���x��&�杌�;w*r�$��� ����V��\$Dު�zF8O;'���&i����}�,:̧��B/�k}���L{��*m���4�v���R��6:n��� @-�<�.&�!_3�I�Eo����b�x#cES�Ok�s-�ʰ �(�B\1��������I��+⬘�7
S$wqY�Qny�x�?���)�"	���]�N�:&x�uf�:��P��ݥb) ��6~r��C@�mX=�{1�+Ū�[��N�ŭ���_�"3߷����6LaM��e2?m��@�'�l�(m��;Z�d��'$-�<�j��$U�/�/Ɏm�}�����Ez�)[l]�ϑ`���"�f]���l�����i��k��>�b&�w��I����wF�qW�+J
E��
��;3����"v ��:�{�8
A���b_�>���\+/7�*w�iT%�0瘓���~^��M�΂e�2n6��-��NV=ő�I���.">h�5=��Dw2���M�s�J�����/C��[fě��п����C�v���"�\�m�{�i��Q�9
E}jZ��V����ǆ ��wH��̈RA��$;���U�Vi��X
t���}6��U�GaY"ߤ#	�^��d�qߣ ��.)m�P!��~m~ Q�!�2/����!7�hO	�������p"�K�qq�M�M��Q�f���S��{�!cچm0��	qgb��|GQo�:�^�,8�!eg�X�(5с�C/�+��%��?W�	2��n}��'�蒒6P3@v�����Z)�|�qE�M���[�1y�HP��aћc?+]����K�A��w��kJ)�s1���53f�v@�x���^a����Jl�lsS���
�� ��1���nu���iJ��hM麛��E.�f�]EJM����J����tD2OvP4���n�Ճi�:/,3끙E�&������2	��@����8D��{O��z>w�D��Ӊσ���N��c'τ��EL|��%vFSW���`R���c�A+�i0|
�	-n��eDm���;!WȨ}#�r���r~d�q�ԣA��,��Tk8���,�?��旈k�~;�N����={M�f��!�I�I�@1��nεI��۠�H#��5-5,��%Tf��Zq���R��@�f�ߠ��^rnZ7�}ae��-44Q4&�ۤtns��v�q����*�'n�8���5w��xyu'�g�l����8�<��lUa�ț��é�ԇT
�69���m�ܳ���W奭�w���2��iӵ�jR��K����A; ߼��{^~~O�����Htc�id����m�m�m�n`����<�.��@�R��1(
l�'��
���2�tm�6f�͹������9����l����{>䱮o�������H|��}j����A���0dX�.��G�{�S`����`-��!�{����!����c[E~��d����8��.;��t%L'��K�'��a|	f�.N�'%�}���2�Rr�����������E/7�_��4�%���"����RST��g"�Y>:)�o3F�y\*߯�z��Q�{��#�p�O���WKN��?q`b|��x�SC��䖇<��-�l����5������y���Q�o0�a�`�hG�a�,_v	B��e���!3єg]���?%���M�w�>��E����e	=/���5<F-d���=��F4U�|D��EV}�W��[��ź�/fnjV�P��ݝ�h{=	��F#��ԉ�"h��#�y�ֆ�N�[_"���"v4O8^p')I�]�V��k��R��O0�t�6�@��`59�ڬ7�uΊ&�� J�Ҽ��+��[�r��ecP�cjD�Q�_�(1�5u���es���q��*�[�/��Bđ�X����±<�"^�O��K �i(?��/��� [߾�1� box4����'�&�=4\�y�| �����OȻ	L����؉x�0\�� �Aq_���	��l7}���,I�E��^V��Q~3�W�u37���	�t(
�L74ܴ�o�����.$��ԕr��(f
 ��CПp8j}hH�V�n$te�+���i��8SV>�L�w�TI��M�{�w�̔�$
B�U\�1s��K���/F�S��X��S@�����'w@�t�����_�r��
<�e�˷�'�t�iw�}�[�<-9#Ǹ=�3w�輞��͂���Z���$ 2�e�}�j�V�P�w�����	 F���-=C�4��LjDʚep��geTi����a�����r��w� �ܯ�S�Y6Ę�,q�3x^��6G����j�d��z4<i�v�m�x�0�|"\O��v��;�<U]ٔ��d�	�%�&8wt�׼Uj<�ϯ]����c�{0?h��'��I�R%/�Q:�I����� ��jz���t%�erN���q}$�1� ����#֚�O��7��s���>+5+_�/w��1��Q�Nᘌ�0�AU �~�5ld@��c���HV5̲8�:���Y��3-T�~�;��jh�6�:�p���yF�
P�%_N��
"p�<W� ��o-.��.�������D���V�o"����
I�;Պm!�� ��8/�x+-��@���rt)B��p��_���m��/]~�nc0��6����T�IqӁO���bH����A�� �`�.��%�ޝԖ�ĨV��Ōѵ��C�:�<#�;�}i� >#}gA	�f3��.R�ۆ��f�z�	����ճ ��nv��4U?Ē4mV1��	n9�&�	FJ`������id=�@%�����+�S��ҷ1�{���> ��*�\-;s�"��,�ߗ�4(F١s�y	L-R��!�@��j�XY���#Ǫ^?�|�u�`�8A�p�㝩�6`[R�#jdx1h�gQ1\��e�C=��b��W,��h��`�D�N�]f��N����iH��.��	st���X�e���(ZPP��P!&n�T5Tw4}�RP:$�I H=H#�� �UGs��I���֡�`����!�+9����*C�K}��@���w�E��OJ��Pn���~�,��ၱ0݌�
��Ak<�~U=��F1�7���'6�3�g��a�SS�iO>����!�)̼K[!�#����$'tp��K�Z�Ъ3��Py��g �̍��t ʧ��!��:�<���bj�#��m�h�,��ͩ��mvrAk!>𪺉���?��Bw��X6��.IĪ&|��=�`�Ŭ�|��͇{B;���P�7"���E�E�����S:���L��f�p.s��hI�E��_u�ט�MM���A���Ak�>����T��@�(u$u��U�X<"l� ��@�De�.)xJ�& ��<�S�0)�+����N����c`r]�����5��e��^��ϹS�}�R3Q|b�t �
tBtR�wF��.t�\-����iȹ��B�6�� -j�k����tV�}���� MD!MAI��j�;_F���[ɠ�����+oNoR&�jۘ��x�D9�A��E�Ӎ��e�W�~��ΐ���9�I�������}KoE����H�}J�/h �K9?z�Ԋ,W2�{'������r"t�a:o��]qys��T=�]~SY�3��=��4r�O�ʭ`����ҡG��	�$������WA�4��>�������6��q�:�ew�æ�ivN0ݝٔ���=�����%#�`z4++�t;*�Z涻��lg���5wTN�w�Y��>W�$�1?�k�Ẓ�^�W"�}g����i$���5��rB#4e��\�����m~�.q��������S���G߻1�܎�FXv��<1����*ڻ�W�E'����)��$����n�\��}$ߔ�i�>K��Ħ��5�XL��[�C�b��*��Չ�a=b� �_�;� �wXb��>>z�b�W]-i���E�9�B6���e	#)�T��,��1*@Q�.�J��I��mF����������wu�?�[z=#�ω� �7߆�A�`G3���+�O
u�o��*��ʷ�}�QB�#}�
��U��,�z�� ��y���ǽ��<ޥg��/OmS���}�_�9A`4�<5�]Jp!��ʺ�>�,he�.�ĩ ��H"���Zd	��FϺ$�J`3v3���q �=�	Ҁm��d2�|.����}������R�etL%�m�9���1�<aYU��P�䁃0���|��Y!��P�H�69�[�pYˆ�uC)7�`��W9i� �|�ͼ��!�T�]��_�{�5���%c�d��y�"uJꐆ:�v>VB6�2�j����1
�	�p�v��!	��*E(9�Q�;$�[]ǞjAd�8ǀ�:����*�h]�v8I�7�#�b�3�U�̮�+G#�:��!�5��
<��v�,����b�2��u�h�Ji��Zi�<���0N^�K�Ƌ��om��\`xXd��f��IM��@��Ԅ�L����X̄��[)��� �[0�{\�m��~��Oh���V�5�x��l4�8��*����F
A+�*@��R�����`�Mn��<�l�R|�U\�%� ����3;A�	e�ZT'�R�V�7WNْȅ�Fo_:j&`��_��A9�Y����?"���(,�(��If����� yb�C\VF�_<"�WZE�D���v7�	��f���:q�� ա���Ѫ�>K��0��ŬL÷�s���]���#x{8��*�BR�%��ȭ�C�W=*M�W�&���/��̼�!�{�5���Ql|t���ᗱ}�9��wf ,$��y�7�}8�ح~4��fJ�6� 7��s�ɗ��b��t��nA��A��O���6�[�B"Ƀ�)+b&F'P�A�E}'H����1��;���f�:h8�#ƥ�:����S��ii��9L�Q7,ꞌ.d#������\DD���mч�	1�k=]�w]x���D�@�־�������'|Ą���G��|��\a> �y�oS�_U�aG̅���%�@�����`�ĩd�x">\��jn-\�V��@�����ty��&���a���Qq2�Y(z���+�Zb����	&G�IBYh��O���Sv��0�b3Z=��FJ��ᯂ܃L�R1֩<��Ĉ'Ή�avĶ�_"{�AS �7PL����/5w� �C����A]Jo%�=*X	'[�#�L��ϊ�4� �&7��	�m�>��S�S�HZ��v�D�js��pX���,�%��	�yf��ڭ��cݔp�.�B�����n��DrU�%ۻ���7�c��8bK-�{'�Ĭ����C�vN6�<`�D�[
�D`�u{�,ɇ���E�����~V�<�IG��+�@��{"�`��ܜX�K.@u����9�J��eaj?�Č	�,��e<�D���.��C�^rQh��2P��ŖHg�|[j�)�����O�@ƶ5Ox�{i/�5�{B����/�m����by%	��z�786OmӀS����u1* 
"���)8mo�^�"Z���\P�8�*�
�X�ɫ����J�7B�?�z?⣗� �k�i5���?l��UW5v7����U�ҮUϞ
���eL+�ޜ�_F)Ú�vn)�88�m�^�n�`����;�1�8�
��1�=��[�!{��r���c�a�d�%�P?���{�����cϘϢ�^��Fc������3b�:�;�|J8�*�����F��ї7������ؿ���#�lan�ĹlH����~#�i�Mݥ�_s���ԳP�V��[��
Pe��[�Z��׍��wMr�U�،�G�[b�|�n��V��C8e+�^���Ϟ��H!<�\��n+�H�Y��Xv��b���vX�	�����4\���\YHQqߪ��m���c��B��U֊w����~J7|�ئ���j]v������|�	��������r\me�&�2�Ʒ~˴��Z�b�l5�! A���K�ar���ָ���e���/n�k�-�N{6���Ǔ{�{bѮ�[X�@���WE�ٳ������ck��n��,��la��y���r���F oH�$b��Xs��"ET[�������%�M,��xH�h�LyXм������[� (š<5y;����P#��X�Ju05\n���o"�Aop�u��@������>Y[Q����+�K�ؓ��M�����cma��0)S:���dnN���U�ڈ�`>��1+���bJ)s�h�m���"���(�v�T;�O��5�ۿ���L���«f�o�)�f�\W��֗h�p�7�E��T'&�s���-e����W��&z��s%���ӹJb\�<m���z�@�[J����nX�e���}��y�B{HE"��9I%.�3���{&?6��E8�~��w�z��5]E�t#.ѣU��Wd{�Z���3��:re�@+?O O\X~y��K���VUx���֬�� �Ed�s�Ӌ���hw�n���χ���E���A�O�/:��H��8ҽ~M�S���������>�5��.Uϖ٥c��zE��A��O�n��]Z��`��6�xj���3�%?5��(7��7�ӽ9�����f2��K�W�=c��q���>��/�o�$5��׈�g�I��^�Б�0d��k,�i�0�OaZ�S�%����d:R�,ݻu��F�c��L)�^��&/^0'	���L�*���&v��n����!�=C�KH��7�ފ.���!N{�տ��(up��(���p�jw�j�w�H��=��A�ԠK��{�N�!<���[��5O�7�Ԍ�8,�����8��A�]s#P&Z�y�L��,PD��kHޔ+OY���	,/��A��OZŔL:^��:��bE�zP��wZNE	�ͽ��!�u�)�2����>��Q��#pU{�ͯ�G��#�"�/���R VE{�$V�y�ll��`�1"�E�y��������� -�$А(�
����j#�j��.�`4�C0i$(KY���8S�# �@�L�S��P��Y�Lɏ`���Ūw��X��<n����4��l[��,>q�Wmq��4�[�	���4�qભ\�{�nngGZ��H�6�"Yg��fِ����#��e�9́�ֈ	,
�c�i����VI��I�^���$��$shd=�Al�O�pm?�oF9!��C!��8�beP�Hp�����mK
�������Ǽ��7R��)er%�NZP|F�X&ü�<�:�o4�_��χ�9�at�<_�J=:��x>>j�����`P-�p8W�� ��aQ(�z��}I,�@�8X ꒸�t吤�qȘ1��,|��qz$L�N�[�\*F��JSB�ށ�
�&�����Iq�{+�淺d�+�%aJ�p��i�%�U�fp��T���B��ZB�\(I������ZW���B(Ni%
���B���io,��^=4�,O��+���p���bI��+�|����L��Eqa���%V[����4�٬��$�k݀S���4΃؇1���K�}��-@�2��d1R�g @H�����0�^��D~PI>��n�� r�,����i�@�dm�L�$�)3�s�O�Z4�a ­�e��2�Ju��F�Z�@�(��˨�V�I��>�+,}oa��5����ت\��!XR���B�Ey��@L��5���6L��B�2����xK-���K���eV�~!ZU��@��L�z���o�!�*�x^��������,�7���qA����Ň�)K��.�4������@���`ؖK�{fM���R���a;���R���L�1���N
1�7^��?Jı��wsoV]VGvX{}���!�b�W��]<���ţ���w��n��)��i��2��+m��~��sQ��n�C��U��V�0N�<W���D��+����-qQ�Gՙъ�&^�@1���	j��ɓj@sb� |�:hR]�CߡS�t���̻7o
�����
*�FXΝ�s�L�F�1�{�͆;���c�>ٻ����>�b���s�X���l�cu֥RFN�b�?���HO�:Q Z$�AC���/�-"_ת
!�&����ȳ#	�ʠ�8���M.�(�J�iDPUU0�eBT�?]J!'��
�pq)�N� $��)���S+J,[���J
v�����oB�r�J܅S_�����\Լ�8-)΃���чI���6�d�b�7g��P�mX&�0�lg\��Πj�=�/�Ϲs�e!8<r�>?4QD�[n�O*rƛ��a�z|�w��^ւ�[Fc�l`[}������6t��Z3��ݍB��=)��y�Hs�ҵ{ul�y�P�-���օ��w[w�(��d�z�2�ƴ ��UrQ���Ǎ8�N-��n4o�F͚5q�y������^"a����F豕���y�4�H^�a~qXZ$yq��cu���?��a)p��n1�Q]�&P���7���Π�H#k__n˙��T��mv��5�Y�5ߢ���schޅ��r66�m�辄hn�Fw�#p�H��(��Ŭ�BH	��@���-~��(��	Ġ]���Щ��c�j��@|���8U�{���ޓ��3k�X�ǨL�1n��@3W���wg�l�I�c�%̌�#�<�1���.OJ m(�=�eG�4�QD�f�I6�H�ȕn�ձ* ż7�Q.� <I�O�IJ�ɻ8��x�	K}���I��@����-�
��1.*�L��+��/��;��D��9�5l��`/��P����bH�l�sØ'T�!��3"�A*���N/�Sr�2��^�:�B�����!��S^p���	���D��N@#G^7���2%��[A��l�u�XC~%�Og�����Pz~����,Y���х𙠛襕���k��q�^=�Ǩ�.���0{a�d¯��A;܀�us�ك1�k� O�8d����"�t֯Γ��r���%H�,�m;;��z�f���T�\y}R��D��q�����u�����!;ƴo��J9�{���r��-9z�zϥ�����<���g�!K	K%;�%�P�����$p�]�?Iy�2���^�CvՇ�<��d�e�+;��5�K#�h!5���)����W��˾]���X{/b��+��zF�>���;�܊�	\�hF�	g���p��\��A�p���.�(Zo�w��2�I��{%��H����$&���`��w��V�d��yXV�VLurJ
�=N��z��:��,�ǐ`�����&���T�&�K�Sg �@ ! �d%'��Y�r)mA���-$)0D5��z�T8��w��Y���z����O���U c~[�;�Oo��u��ug%�)�+���	8P�7��#A�*+��?��&�]u�v��‣(���6;*E��mǒY��tq��x�Pn܂�@�������ENWA6��:�~���w��GcD�G�[���/�(�r�;h�b���Us@,��['�������āD!��3�����p�hb�9�r�7[vg^�ӛ-�FQ>9>��pY�h5e���=���8��#����ĝ�8�3��D�rA��X�Z歝�	>�G��:��f��Kd�� ��\��f�o����"b�t�5\���>�~[�E�#��>ޜ��p�Oh�����Ÿ�� ��c�l�7���gP��DA�0�%�4x
$���ݍ[j�AT�0���]����s/�>�A�G�p3y�n�å0�&���s���!���M��*�c��@��,Ʃ��V �=�zW�f%�(a����2^�R� nHQ\!����d�Y",e�Qe�9�oZ��������*�K��Ks�r���V��{2=��y >ez�h<��,��i��Y�W���i��駐`�+T���؃��F�$��`�Z����|�����۴�e��l�/G��)7�������`�����c���|`ϙ,~jf���z1_,y���5Lb�CyYnH���RFcq��� 8.Z%�K@v�JD�G�"QtX��5f?|�~p;�J�C�0S?g��A_�w\�I�����Q����3C�e�!ky)N��*�Mۡ�"��Қ��B���lIZy64��k/pT�G��	ZA�L��6
�{������j�b|���i�
���7��,���w9�{�`,��\�tD�� Yoiq��Ѓ�7���~�eUG���>ȰIȼF[��]˽.&,��ק:]fO��Ħ�"�.��r��]����X8�G� ��ϗ�-d�����.�|�Ť�L�����L�.�Z�8]pgؑw(���m�}m؎�Ic,��M?q+((6��
�G�[�o�"(�O������,��񌌛H�P�Z�����y^����-�Cu��$\m���N_M�8#P͢�^���YK���� $G#|�G9 ���Gʃ�ȢJ�k�||��ng:��y�"�T�z��z�6�h���iF;��Tmq!Fxy�U$,�������EG3��f�*9�JL:aF1��az�Sp	Si��	��V=d�D:���2?�,}��%��an���ຄE	$ڙΘy���H�A��^w�>#4a��Mw��f����"vX���D�DN������u���2PpwQ���{�c%��>i�T;%$	� �f�RB��]D�M�"�1H`�g�����2SK��I��&0�")��I7y�{��p��a|�/��A>�'1� �bz?�GT�3h;�3��uTהF6�-Q�)Di<���V(���D"D���G#:7乬��0"N��bv��n��X�H���"�������3��sA9F�XDu��'�թތ.�(�$b`�Ӄ���p�xoEf�!�;W/w�ˈ�G���s�����h�9�����a�{@lQ@�(��-��-aF�H\��Ч2��Oe��7�AHž�S�C2c�5�������_:-)��2F�<j��8;�Ly�B���S�R�3VzS�H��n�e��3����=k'�0��&v� �%<8L�+��0��˻�
@��1�@h�@YZ�_)q��MZ��n>��������(�1nQj�hf��x@��!��F ��	tR@@!j��-E���,�
DD!�!�@����U���U�PkD����M����ZC F�p�&��q���Dg3�5����U�;��|#��_ ���y@N�i�7�k�9��Asޟ$�'���!���CgȋG"&���@�;�ف�f��IhM^* =��X�Zv�m��m�� )�6?����b\�Ğ��}����z����āHtC,��<mOP�|u�l�-�tD�%�`&Tk��D�P�M�#���T5��Q>�q@�֍k��G:]�Q����3�k��򥞣���~���GÀ�&�Qn�������-�]�f�D-�� ��TD�""U��װ��E���V����S��x��2mc�3x��Ss=d�ȃ��4�`D턷�mDW����Oz����Ey���!W��NN%0y��j\�Z(���Oe�b�hiwX+�r�(J�R�i�I�D�~�0ӣ`�f�c����r��1��=I��x��Fz���5�"�[��Ӓ����8�ݐr`��$��e�Z�5�đs��sͯg�&�I IP�q�7���Z�fW?�@獿���#vc0ϋ��gs���HU���$�v�_�����Ǒ��Ϊ�wYJ��=v�f�yk��?uE����:%m�v-�b�N��x����HUj�Oe���%j�8��37���H�vt}�kB��4��A�G]���̉��ٝ:FO69�'`����2��*�fn�|�ԳN�3����2V	�i���P�<���i;����qp�[7������Qe��l(Vx��a/j�]zq�x���j��'y�Un���r�QsTޟ��<�I��΅Wu�%��s�C������G�5��+Y��#n�7�F�Z-�ќq4/B@x�i���W/�m�2�S瀠P�|�v��HM��rZ32���$�N�ݮw��~M(�>�tL�Ü�,�b:;9�q���%�c(ɢ���fEK�Ғ�S�W�eN��kۼ��ft%�w�˲���'��R����h4���u��l���6�@E4�A�L?�҈����[٧�dm�/`�:>�G��6$*.��f�z<o�Yw��F�@�U���͔A3`=0-!�sI�:����Lґ�6Ŵ�ſ]���I{����B����r6�C�lG�D�Z�GO�䝻f���kGڨ��/��S5�}�S^I�^��~�m�o�+���;�з�d5�e1	뫻�g��)a�\�̹����eT�R�9Z�h.���F��X�7�s���i�_U����w�����O#=���	t`� Fp�D�"���X��?�} ��B���Ar�Bg|�1y����(�� 3�VGP��xh�� �z��fC��M�x:}�b��ڞ�&�2jt��ko=��J J��7�K]��Z.�� R�w
$J��\�S�;��q�m�E6o+�+i��
�*2Nr�9;�Z�[k��1k�=8^��EC�nM|�@AEo��^�
� ����w	��_G���bR�;��M7 U������FF�Z&��k�a��v�kE����[�"|��Ka)=s����q��?�����:٧�����y�9 1.����`D�TFY��ş0d�L�GI��(X�!N���}?�(�:��7����}��-V���2y�8��}��39�ݮ�ht����]��\�c���Y^���X7{���Ҵ3�]"��	0�RP[8x7�_Q	c�}�r`q���)�ӞQ������8ڤ��\A	��ğ�)\>����^	�;uYo5��ib$k���� i>���,$
�	�����/�r��ͭ�m������<�^��L4��Hq�< �-�r��R�=<��:T�R��`{�F����┷�aҢ�Ҁ��)���3ҝ6'��P �Ί�,�Z�SZ����-|����	�6س��fdM�%ܴ��n���?�򺱵	�ђ���y���;�;N��$'�u��($l;K?�6�/u\?�iq�zSJ)ȫԸ�ֆ�*5/�{���G�UpR������}��,$ߠ��-魰�]���j%,JH�C4�R?J'�TϺ��o����\��NEL����t+ZqT���!ϊX�r��:_�0<f��OB$u�3���?�va�����01%��=`�3��Gi�-�+�IB�qh�&.�^b��2y��̪2�A��^����2����f��H}�*S�G\3׶�r�Z�*!�Igeȧ3��-�	�g��9N��ӽ��U��Z�O�M�/�-<�@n/����ۥ&]Z�N�*�N5�r��.�=�^IB����(q��u~PO�: ��J*�?[|b;�����ݛ�]f	�7����BT��Z"�ɲ���m��)/϶����'>FпG{�5L����N�Gk3�G�J��m�LA�&J��Z�@Z�18�#:R���z��p���8���X����.��r�K0.i��-%w�O�}�%3���`V�k�e�����ӝ�Q��i&��n�G^�L!SNn�Hm<�&�18�kn7R�r7OK��)`�Ā�N�j�_�3V�"m7��9ϊY�LZ����؈���A=e"���Xٮ �'y���1�.%97��z�4��?߃�e�+'�z;�������pz���~���^���.�����E���ـ��_��0
���4 VvB[1�D�e�+�Df`Q)���J�9����H��6�FsW���З�Η��g|u��HOG(�Ԏ�/�Q"���"�yA*�#�,ϒ,Ϡ�$��I�2)τ�쌽/��x�bT8�Њ\hR�t��c�gqq�R]Ŝ$������q@�b%MQq��ZDfx$����n^x���;H���Ü��L�§`.�j7x�n��K�[�W���7Z/�h�]h+�<��	��KO��d�DΦ2�����i��P"��������w\e���b��?�;ئM�R��Ǿg��E��:r7�A`�����y ���{�ԯ���G5.q���ZS���ꋤ �z�grp�Mi��N	�N���m%w:�����������d��`����n�Z�
L��~��:��c��K��!b� �e�{k߃`�T!]���|[�/�^���WǯtTv�w!��賑˿YҎ���a�3�uNM���K*��Go�2M
��m�a�"|;��7���ũ�ڊ�I�2]7�G�E�Ѩ�S�E�m3���X�X�0����:����bv-�� �J�4�L����;Ȭ�k�"��t��/�����%��<�Z����U6֗0b���}��>bu�[\0O�@�0�D$�)�S�Es�AƐq�jWO!��/?���@fk�s�jB�n$Ã�.�����f먂5 }1�Dc����K��)}O��X�<Sl�"��Z��M���p3��e:a6��z��5�ր
�3Vfs��m*�ü+���ohp��EI:a�Z\�>��k��F��D�St7�Ž�GP�0���gJQ<����;S@�m����v����h�c|O��rO�J����J�Ym�7p=,HE�!�p����U�6�J�~+3h�{�CH�˙�W���Վ����.��0�HV�_'
|qY �ڇ�����A�(*�G1%���EI���<&�l��Cv������0N�?�X6K㹨9��|�Wk����
�+���u���@ɵ@JG��J�2 ���n�cd@[4͙v������g)r��9P������E[P<��y�=�����k{�U���eWT*.�\jQ�+0��+���$��{����N�;�s��Gi�����T�甥P�l1&͂u�)��0���͍�0(K�ƹ�:z3�b$Y0G�I��<�c�3��o���~���Ϙpr��*�j�a3�� 3�9�U,��UBV VY���k̃�������%P���۩��.|G�6j�:9w�SZa���-5����Ӻ�)@�9��nz��HD]��,п��/�<��V�V�ng�������9���t Jx2PJ �k@Z(6<���w��V�R�"��{��J��nٴ |�@6ƣ ���~ۏ�h��E��yo�z�Y{��v��2q����Z慎����+�3���G�+0X�;?�R���`��n���ţ5��*}��..�<��������ZG�\_�:T�S �,�Lp}�Z �{�=��@p��� ^���0hI��Q�s9L�!��5�r�)O����?*����F�U@	X�;��|UD
x'��J ���P6����\K�E�Y���!�pß��,�I�vZՐvL��J������zc���驦�b��e��SA0�j7�l"�[0�J#�Wn�n��
�cƘ7&4ާY'A��CK�B��޶����]}��}JR�:���M�_z\Z�%�D���.��ch�ц1l�]Y�jK����P�h<�ʔ+�-Yݖ$PbvU S��]�cۋ�V�ud�� gnZ���z�&����B8�WA/u��e��hj?49��IuRym0e`[! X<��m���q�0�:1������O�W����-�!��< �*��Y`��Z*�y���B��yU�XLf�G�A��#k�X-+�z�l�C*�\�p�򷗩�]A�@w��;.���w^D��8dj�́�lUX'%o�$�2P h�U`�B����I���p_D�VƐ��!g�`K���B`�8'Ucp���R�}ÆR.�^&�E(�Ȝ�ۗw�Ǚ����沵o�����Z�J$﬿?�$�g>]C��C��C<�s�k�Je��g��gg�+�6��TMζ� ��O�wTo.�G#�3���p1���;���{1�z�̩=&���[��Bw����ؚI,��_��џ"#�w��:7�E�4��&L��OԚJ��{�wTN����}h����(�N�r\�\���֜u�>�p�L�$��^����X�%&�h�k/nm,k�A���)b�&�;,M�o��͞���h$P��!#v�P	�!���>ͳ��;�[��WS�2�-�>�π7����fY����*|�ш�����hv:�V"](/䗯Lْ�����0l�>䀘��;��������'X_-K�x$ѣ�%��o�Ču�gkgNW-��RP>��F���S (Σ�%݅�i@17e�=��ɹ��WW-Q-�U�o~n�����zr��8�����w�����G���c�4�]T�t�t �0���ƒ��NS #e� '��8[!5'^B? �iP��1+$0������qΰO���܄��%M��Y����`F�"4�8�&Rg��p�v>W�@2����'��>��(~h�D�#�
w�6\�sV"l�%��e�pQ�����<�b�$`�z[��݀ï�FvQ�߼k�
����|7
;�v@#t�R(>#D�z�"`�0���F�)�m�Q}��#���A:8`PM�����f�([������CI�KI�:~V�2aF�"�;�8m���ޣ-Նi��{�xXg����ˉD�QA��y� $Pdt H��<bz0�
FܯF=C��`dv�F�6��7�����p��p$�dx���x�8������`��e�����W�07P�]j@o�랩�Γx�@�����LQӢ�w\�&�vep�43����!
U�F=������u�|�U�IF���u��E�0��-4��W�EN�r8��C�BÁoJ��7��X��A�'�A�F����h��[\�K�A�M��J��ûzb�fޜ���z��=8j���� ��[~�����ق�S�4����e�8��	�� ��+�6�C�C��h/��������1J;Y���..��+�P �#��×�N|a�R�AqQ����eM3�
��@�p�m���E?���mH�~p�O����ЫV�S ����y��!��}W��n����/Aj�@aR���|�k���a�b��3>CI�tc�������)Oi("����U�x����L��a]��ȧ=R$S�0�Lz�u����Ono�]=N�a��5��S���}g�e�΢���(,��x�9�Z��Ζ ��Ca�s+5/5q�D�� �`�JCX&��`O���ؙS+oD�;c�����(���9����Se���K��?њ5Μ/��]�N��'�)C˺�qe���L��S!s�A~ѯ
.��b_��[
T�Ί�5�X*��#	��;|/7a��T��rx�:�ȸ�ÿt�>�L��&{ـ��Pj�"��:�X7k��uA��ɥ��_�֐;Fr��ߓ��-;Lo���#^]q�)����k�p";Ν�+n���~�����xF�[���,i�����=Ɩ��6�����=4��M}tf��eIѸX}��}j��j�>�w��Ƴ�:��أ�v=b�cQ7���W�lM�H�K�D1�b�s��,�6O����:6���i4�;���Ӫ+�{��)
K�y�����^�����w(ﺼ���wk�?u��Hʇ����1m+O~	
!�{�7�C�@v��50ͮe�ϧ!���Gd]Nϴ�܏��;�n1
������76���j���BN�o[.""/�{K���*�C��UE҂�ȯ"]�*!Մs]��>K��i`!^gY��ݽxƤ���o���<0,�p0DNu@�sH��$*c\	�T��$-�b��3x�� � �Т@p���M �G��Q�� ���!�s��	�<PB~�\!^�ŐY�k�d�vj�^������u~F�?�AO�E�X��i���!���/��ؓ���Y�Θ��޻�i��ILB�#���}Ӈ� YeƵT-�՝��c��W��\L�O����|�s����)���KY��nvmY�8r�n����;��XLصB�n�� t��:9~z�7���h'�!}��s�E�(��*`��B��g�X
~	���	W.��\S�eU�D���	U	P�^|>~�<Q<
r	���	S/=������Ϊ�SR9�t3�kk�}Z����,삫�"�a��'6�ƾk��t�FFy����$��-������p(�l&�mh��i�/%�.<�QA�����D�Ay�[�8f�.+��-���/�sc50����m�/��"qFS�]L�ٗ��ន �A�+,��kٿ`��B�̌T��FX݉����p�_�q����\��dR����r&3"���}�7�5��Q�� ظ�;jz_aZ��x�1�1��:1�ܴp8������ȹ5M����5�.vg���K���0D�M��bp'�� J�9�X`)�A��Y� ��`<��n_���j��_������?��!_��a̓���8���������D��0{��TD�	��?��L��"z�9m�
p9ā�+ԁ��S�,:PXC���g-�;�3�+ԌqnŁ�/S�����i�Ou0n�50(h4?��50}s-P�ڠ�����Ǫj��Z�^�
(�$ ��Yؠ숲x#L��F�e� p��Z5ے�Ex>b������a�A�B�9Fx��]m
�U���U2�G��u�0r���ː����Ç3����ob���M�p�p��cw���7� &�(8ev�S�Rh*�������,;:q�Z��?z�z�ے�QDM��_��Py0���W8���6��佯��I8�s��H�$/y2߻� �я	���d�m��ub�T��z�`O�z׬�����>���g3R��3�����V� ����S�3�F�+Hc5����������^�܂��1: �������܄�S�)N��ۿ�BV�9��Nf�P���
$����w��f��]�+�GD��2�"��Q�$�bl����-�c��KS��ma+�eh���h�=�:�K��t�G��梻�81v���#�X� gJT��:�f����U�����u��ê��h;k�A���0���n)T48F@���3 O���>#Ŭ�Ÿ<��CJ9�sp�'!O�AOkl�|�{ݪ��ayƴ��|V�  Ӑ��jf�7����1����r�I6z4��_�]�|4�~�X�0>���h���3���{>�4(��b��P�����
���I���̲Q-Aѐ�Fi=�Fg34e��Ƿ��T�+#v1����9c��u=wN]�Wt�ي�]��Z��wӮ�duee9%	!;�y���B�F��%�<�dA"/���Q`���(�Q'
�Rv���>�3/e_T���C,����}EQ��/�2T<�T)�yMpRJ�ʲ��p���:��x���p�%��Q��Oí����kIN��\����!���O��x^+q<b,����W�Y�<6��cΊ���_�]��cv')�dQ��m�7����7}t��$c���H�� �cJݤ^�oе���O�8�H�C.�e��P04-�������sa���j�3'�^t���҇�S��ҽ�[��T��t*�M����4
r���a���6��)� 4�S��fQ��,�~��Gn� ��_����;����j����P�P��Q� Y�"x�"�$�50��T�{�����b��Muv��l�a309o�,�^���t+;��<�x ���n�sV�`��B�����$����~ɾ;\����^��Q��SU�!�� �"��#�����X��z�w�O#�W_�Q�uQ�79k�Y���Y�#dɯ��l���?y ��B��M#k���B�۩�ax�N�.�+K]D�o��}�4'ժ�Q�tj#����<x���{���HR���S3M�{�{Ѻ��qf�G;h"��&Hf��k[�~�}
ˑ�����B�:[;̼<bA�FۭJ?�h����d���ɚR�נ-q�/(�������u�?�f����.�\���g��B|�$����T�g %��
]�ݲ'�,saf��p�T=-��D|��5+^�T��ANI���h(�� �B�dm�R��۩���`�����dא;4���b��?)��l��Z�$��#]�7,�{1!�n���vG@��R1�T�ʞ���UN�n=�r��6؁@I�^���d�͞ꅽ+B>!�u?N����B~>�۝b�ԩ��F�چ�2QN�uV ���dZ	�Փ5��9��uC�Z�����T������5Vr�O�Ջ��&ޚ�Ug�*+��"�}RRq,�#ǎ�19>�(��M����)S�^�\^R���������PoĢ��S,H��>�v0j��Qm��`Y�QY��f�#`��C%ō��ή�G���+�bl%�{�Y��䖪��W�d���(��G:��淋�+�[��K΁�fXlс��B�Lڰ:S��<މ�څ�\w�����YQ�����?�\j��O�z�#�kǋ��-��C��5��T���������v���r���LH�|�_?<b�t�	&IyБ�8��3H���n�Ny��*�&=�;��
D��3�۲�/������g�W<CP��O�=��]-My#]BkibeL�J��L8����::���lEk��f뺟�Y^��^�G'C�yPܳm��''}_�l��;�:T)&%��� �Y��žJ�����������!��ܟ׍k��{C�)��z��J�BI	��.i,,� �Fu�Q%KT��Iiq�LCm$#!WI��qRK��6a�RF!���O>�<E���.��{��
���'��~�,�Ԇ_���2�F`�D�c�V��#*A�=H�>0�ױL��[n{��w�J�rKN8{Dp7�0�vN�$/KH�88�8�����dW6�1��\<���#;�>wĮx�c�t_�&^O�_�9tQ۱�"�L[E�Y�JMD�O���S
wKʟ��� ���L��y:��ւ�bƏ�vq�3ѿ����IԻ����iHf��S@owoI K/�R87�/���	/+�	T|�x�2h9��B(h��;�UJ�;��B��)���]�F�}f���l�1\6�O�3t���نv���9副��+AS�/����Q|2D��yDƧ ��^����6������V��F�|��?���zo���c�6��=�#���f�S��F��Ɨ�\A=��&�w�̈�D��ɛo��@�8��ԙ~���~qm%�W�֕�T�ɔF>�hy��4/&�c���-��
FN'�}��#�c<��aoNwedŶ��yYr&��9z�D�;�X9a!��J�4�>i��ٝ*+�/4����=��dy�ㆼ�r����XRߤ�6Ad�d���V<����}#�.+��F���-���(�
U-1^�Te�	F�y�U�=���؁���t5���� !ДH��p�0��2�"<ۏ_��K�j��
z���^��j��(5j�KEf��� ��FuZ�˾ӿ�]�K��/��`SJ��*s�laaPt�����s��B���rsI<��O�'o�5�igxOK%���󂹨O�l�u�N�?c�F�3s�Ah�{��=��	��J��f���»{Jq����d���-u���q�jNKw��_����-�v.)S!A�!�{�T�����01�%k$��е�$�0���B�r�R������Y��]�3o����iM���M�q�8��n*��&qK�]L�
�#�����A���
�J�-�/$0�,%��f��L�/��W��8�p:'B]9��n솼،��Dӡ�z�����7�/��ɶ6�o�+�R���^���*��g��w?`�#ϱ��n�:��y��ل@|��h�|��E��+��2�u+1'��~u裛,{��x~֒����z���a�%d'�����va����p�j>�W��P����R�*a�0(��E���<�z���N�. �5;#�=��=|e��o G�6�xf�م�{�	�Yl�ᘚ%3��c%���}-�r�.�>��uĸ�-+.�|"�:�C���V���n%NʞY��n{=��4G�k��]������R$k��!v��[EW���Ԇ}};Cנ�o�\�:��K�~��Y��0�gD��HYgT�OA�n�U9���ڧ܊���Q�����8�\(�����9J��l���l���xNh�`Xa-������=i3��A�ɝ1���O �r�h�E�zzR�$6�W�dCiԄ�#�]G4~�߳������U$�`.$GV #�HD�^�o�qgl"k&Cz���]���hʣ؎KjĹL�y"�����TY�f�e��t�g��2�@~$��ojj�2����\ҵ&-����Ag��FA�#V]�Q�Xs-Y2xv��s!fI��{�%���4.!�B��� Q��]
��G=1l���:�㠅��o �pn;8�)L�l�a{SS�{���d�m亞��]I���g�Ω��]Q.	�m7�Gs��'�A��"Gq�k����Lu֔��a4���0h�@%��xS.����Q~�#��]?յ�!�g%���D���Җ�q�ڈ#�Be=_ְ:+a�~�i{�>�Z{�����mfu��Hw#��F��
h]��ҕ�x���.��V4��+�oA~~�.��UJ��:Y�^�0����F]J�C����M�}w)_c-?��>�V�"ƛ��8*�Mqw� ���X�/Ӂ���Ց�����x����d�cb�؉���nj�7,�[aaCͩ��H�?9&2�����aOî�P�!�Z6Ɖ�׽\���3_��%�K�����9'	�C�W�V�	�ߛ����}5�y�Q>m����i�=�5a�|�!`q��p����t���UX%L@�Q��Q�57��Tg.ʸ��?�y�x&���Y�bŝY��G$��w�D�U�>��{U��6w%�w�#���<sG��CVI�_��BD�I��'�S�4��F̗T����A��N~v�$���g�j��E�����Xw�����.B�(W[e��ŕ�|}f=�,���1�1r�m�5���LZc��bd���܏��`%�ҵϏ�貶�ݑ���5�������EO.(*��Xq�}U�:��������� (-���騟�����ci}�g��WF�^���0u;�"�E�[8�tB\�e�;�3��/���Db�v`� T��b-��X.E�[���f�| 㭽/���M��qcW�V*5X0���Q�A���7��3t�ϳYE􎚗�i�p�]11���:d�~( P ���W��[60GBB�����[;��<s͵\x�x�����N.`�g9����kt�!��2��!��Su�Q�l���������Uk0}���]���.���;%��dp`�3x��;�E��fr��}��գ݅/���ڛ�'��0�k�F�(Ny��'����\"�I����d����=��b��E,;�Z�w\�)a�j�0��h���ü;�}\���4��g)�Ic����y�8�����2��gn���-B���j�n����2�	���)"�Sy�ê��	�n&,��6�2�1M��T?����I�]O�b���Q�̰���,y����.��*߭n.�����Y�o��	�k ��1���@�.��ZTC��Kǎ���J���K�'������Q��|�x�/P�Ʀ/�K���\6�ӳ������5��BC[�I�2S������s��Ȁi`d��Q2�!�p ����+
�K]�ɉ�凮A/'I�(�W�cT�����nCm-�9����H�X$a�>h����u�
�#Q���GD�-YUk�Dz���Q����V�T���bx��z�s{�6;�gB����(�.�����|OF���~w�Fb2s�͔#gXYţ�ݕ��k�|�J��t-!�o�Ȑ|%��5���3�9�׊o�QfD�-�:t���br_�;Ι7\��@,z�=�CB�jo��5-�)�t�����ܩ�:
�w��H=���ǋ�iA_���.��Pr�B~vcSI���,wїUrc����/y���A���i�ӆzAX<��e����ܶb����}e�3�%�3�{@������w��C�|�m�	��u�P��T�-ɠ�,�k�D͆�Qm˔�C2;���Y��+��PKD��gt����:l"-�T."`>6���L��st���@"�9��,��f9��}~^W�	�p��n�n�j�~���[������򘱗���J�����9:2+ 4)�������µ�Y/���~�Z[5�)H�]������Bj)�+-�5����k��Z�]5y8�"\��r��u��u��-�JK�(�����P|>�i�d!�8uQQ:��iTǛoy�Z���Pa�����[�G2�<�R���yʹ&ޔ�t6��^�0���¹���=�f���JV(�y�i��{�6ڊ�A%�I���6[�o��z���Z�m�)s�͠IU7�>�"A�n�[����~�@4xw���9�A$�hWoƎ׉�/pJ���k�k��M��Ch� �4p �k��l�g��[fJ����|elj���",FL��EBH���ͤcli�A?��XE��iT��@�J�s#ﶔ��/GT�JU G/��g��[rJC�ꚔI|�4'�@�<>��t3��p3���^Sa��gb.M���)��4Aú�AM �U3���~7C0�_�,y��Hk[�O�P#x}-n�Ě��<�ƞ����>�!�i
7�ӣ�$[X\���[��3X�"��c�Yb-߲�=���КI�����ʮ1r�
������ݎ�����4�a�Hc8�����H���P�%�ۼO�=tE��	����V-�����?�쮌�ַ����2ʭI�0n�m�k��h�F�3�e�7�<�L�/�-�W�!t
�hE��Gۀm%J^��;׾oj��/�Q����������cnS�c}p[l.3����eo�jN�a��p(>ɰ%h�?7��=�^<׳�Ū֓l~���*����ܚ�?)g�CzC�:�2�'���+V�]�L�/��H6Q�n��G��6SL�JX���Mq��&{�'��ocM�%"�i���X0�`��qoB�����6�M8��e�rj��̦8�Zxx9Aś���_�?�wݣ?�_l�!ڥ�~h�\2*��ɑ��.7|���7D.<����l��N'�I?�!9m���B�-�Ψ�b�$l����u�I%��LK"O,8�!lذ���}
���~I�+��/qwj�ߗ�.�������K?���+['BLiS�'���]ׁI�f���C�sAb>!�%9�l�g�I*֨Ye����a_]܉Tq2�s��veTQ�)�z��7��Yr�2�;�����)�f5W�N���P1���[�O,�y���-��8IpMX���k���CG��]l/,�����������P6��jLRe���3� �,V'�K�%l'5�J�*�l��Ռ��:���b�fZT�e1Z���|�	�FmJ���7mS=�	T2��;Zr�#�Q�GW�j�Jr�;�z��Fu]����kam41���C?@](4��yjQ}������t	RUgyk^��,��'#��B̫�D����kE1s��*6z���m�6�P�e�a&ɛ`߾݌(�o�u�Ře���d�~��Q��k~^kb�Fs�57���|]���-�&�]�T+�b����C�"�o)��2��Ѓd8�1(N+�U>�4O��s}c"�TX ���Ĝ��K���֗U���NV����#�d>$5�~�d�O�p�]�� G�%�Joj��{3qL�x��Hg��u�R�,؈��	'�o/#��*�J��<�n~|����J��&?��ڏ�V��彄]���t\�k���U@$��5 �B[G�8TPs�<�Ik����U��]�3�rz���@*�g�Va��D��e�9��j�J�� �r1�\a�<W1��9Ŵ�����L�
=?�ѡ�t�J�k�����{�wP�9(ZxQz��L�#������;\b\U}7zkcQ�>�a;���Ol��s����4y7fp��/��D^���n8�a!�Ɵ:x�W���W-��`p��;c=8*6�)��el�H;�}�hg���2��(u�^3���P7-��@7
�#������gƺ��ƻ�6�l��ٸ�(�fu)�J��k� Q��[�?֓�����e� <��Vg��U�b�aMm�,Th�J�q��Q(,��-�����K'��m�Kۑ�����1��V&�=�k�����ٓ��X< R}0�^�b\�����X$E0��?k�D|U�?[,�ݍܗY�~A�AT�F)�	��@�q�D��o�@�:R�\M�����de�X��ϺE�߂ɘ�����/Mc���A@��W�oX�Y�?�����a��������rw��{	'dgw��jy��HV�*"�O�D�{FQ}؈[��k!-�`��R=�t1�z�@�"��qu��&�t��+a�@�[������gl.������bl���f�L�9E��AL�M�I�qCu0��:����3k�v�X���a�s��k���(�?,�Չ����=�kl����:@��*Æ$�7,"�1�}�o���q)�u�ŗ�d0�h��K�r��ssT��:��BKGe�h	б��]�1�]�AC-R�� �����#n[��]�������b5�_ 0�~��a8��*�@+c�W��=�c����c�I	�7�5���Ŵ��ʆ$�Z O���=o�-�>zkn���+y�M�������g�K��)+a���r��%s1�C�`\j�rp�j��Z�O��p��t*ܓ�@Sﮧ��u��V�Ϻ�r[�M M��:�2V�}1V�W�6����@uO|��?����܄t�a��t��x�߲$�&� y��L�#�Fg�����U�5$��h~T!���ǩ�k�����#(�9�h���8<InZ7"!2�)��Jt褨3j�]���V��� ��Hy��ɫ�<�'���1?�wPr5�Pk�ӊ�i�V@UV� K��6U�:T&��d�l;t��˧��5)�O,�����TCd�TZ��z맚<&����L\�p:$�p&�c��&���������9D�^�%�3���}�Jfv������gJTF��f�;:�i���'/�k�0�c�9r�Db.�/#*�,��s��b�/�0��j'Q�2���۠�슅�0=�5�r��΁M8�D�h}��^���K&�M+c���R�����d���p����:��K�6��a��ȮY�����%H���A�&#�?L)�`j���u�hG��D�B�v��wݒR�!勅A��O���	,��w��9���m�� S�����쮁�D̶diԣ҆���������!确ȯu@[U b��UfܗKB�ܤbuhʣ�7ZS^H`�# I�_IgTvF�)�=�N�P%*���6G}�6)�`q=��i8vv�����	���k���f{�y�d�(����:I�@����c|��*;�/"I�O���ʇ�+B��d\��}4ɸ{���<�5�k�8�NZ��\���۝|��`l�K�K�"Y�-�[Q���|~�ް����R�����F�v�5C$eqMF*�H6�-Cw.���fY44Nw�:[��P�p+:WK��)κ���(MC�0�ᨣ�Y�+�7#*N���t�W�o�"�p"��eN��+����R��]��u	�0ߕ� " `qd��^@}۫�Ղ���F�u�W�\�\�W}��{���5ظ�[�,7��	�s!�\�w�t���H��Qѹ��\S�~,f!¯�BvG��k���p�� �:��;�V[���˷ ��׬�.4^���>oRv<X�a��tNdcQ0��a�E�[۸����*���_�K��S���<��ݜYr���O�V���B-V:���=�Q�]��T�g�7.ڙR'�y\_��h3�:�-�re���y�\S5tGI����bUu�e�nO�y���9;>[�z��"QPn	zXp{��.w���8��0>��6�ч��~�d(��>�b��R�7�b~���O��,*6a�l�O���θ��Ɔ3P,������ql$#�����L]�ip�&�01.��:��聝����7�Uk;X�ù����j�3���me�[d��s�fnf�� �6�9��cצ����Sm�m��7z���s��������=���^��� *	��
�TET*�,*P9���,@��̓�J�xI���ۦ>D� �{�l@>�6$�`}�O�S�_/����������i3[���)k�j��RjF7�L�� 8a/���u!���
w.tlW��ħ����� fV͉�ra���HA�!H!���J@s�яm��':P0+�/c`�9���3�f�yg`����b9���)U�|���� `@ck�eN�J,����0��R���T�VtZ��� F�z�A�éT�d��+q4Q&J��uS����z���_�$�B���\�v���Y�)����7f[�B��h�3zߛ�^�O��_T�i�Da�)�.�`A·츑�ڦ�����ܹX�ē�I��e�j+* ~J��543���z~�
�'�n�î����BYXK2#�Ы�a�1M��%(U�u5P�a\WC'���=�S4R#(3��T�����|����@��"7�������e��P
�5u�ݮnYh��*�F-�ϟDz�Q�-k>(��W����xGuh⭟�>x��:T(��"�d�ڜ*�`� `@Y^�Au�о�Lʺ�X�B�tei'�S�T�p5�,Ӥ�e����A�sq�XY3�Ҏ�'�%�#��x�.V�ʑ�]0vOAq	��ڲ`ץ��V��l�=|z��1S�f�;<-��J?x���2@���C&xM��yu�)怌K���JѨ�8: e�]F�h:�goi%�=>�XT%{���F����8�}78�X8��2 ��`���+}T3|i�E��P�����e,�H�3	�tu��g�w�՞�S����]M�̆?�!� ���Ez���\��4�i�Ng5��)A�VL�ֺ������"	�Fd0+��b�T�-l���JD(k9Y������S��Q�=`+�ooXf0��
6n8q,E2V�z��GV�إO�U��@�N��0&`����1����%�!Z6�(X\�B�߉S搷�`�ތuM!H+ ߌ��"�DE�\T���m���Ug�a���w#��m�b��o�#�d	?��Qi��cX�@���9F�~(iQl-F/[��P�l'/g���}���@�}2>H�E-�������Zh��KU'����\�IH����];��0���^� �ꕕ�x?fL�2��5��<�f�_�3��+��VLo�br���8=
�=�G=fҫ�JV���P�s\#<��u\�8�U�}���txpQ� h"����
���B�O�����%���^*E�����xjf�X��/l&�Տtó�fݮ�:���l{)!�&���c	���ܻ��K�@�gY�n#���ۉw5�H�Zu�[�_��Ȼ%$�>�K���I���~9ϳ��܁�8�6Z�fw�r>�6��F|a��\���I�Wc�̛ĨF�~�Gr8͆������3��S�s8�[Yi܉�d���;�-�o�U5}�s��{�/K��5=Ft<����cr�_^<�Ծ��� 0c9@Fi��L��,-�Z�=F�?����rα���I7-�����?S[�9��-g�7��3�@�2~�Y}N��L������j;�U��E�1~�U�SֶX���bo���%����ȣ9�쩡�Nz�zy�?+�V�/�`Y�b���[7u��T��g~؉����F0�M���D�~�:n���7x���M���f��l��P�DaH�-�/�$	��imע�-�:q�X>W��h��1��[:���	�����jV2e������P����]hj3�ȇ��5)п:�Zs�֫\��} ů?� !�.�<�(��
��&l��#���km>�B(a����\�Q�� 0`�1�ע
�g/|ӛ`դԯ�?����:�Mxs7�(�y��7�=K*o��oх\䙃��mGgL�V�t�-KY���q�h�Y΅�[t�_�&?2	�W,���T{�����󑺂V@�7I5�8L��n�p��q0z\�e
[8�@bQ�5�?���`	�u!%�Ҽ<��v��s����\>�GMg6�����S���1��4�ش!���6�T���-�Оsu3ae�!��%p
$8��#��}���L�f��qh�@���'f�I��;<h[\4)\W(�%�o�U=Y�&<�|[�
]<��.7�Ub�=
b�hq�։��h��Я��;��T���8�Jɔ�g�����4����`0T��h�D����3�$|9�M��zPPH%��F�lbOaZ<bZ)��%:�*fO/FS��o�j'�]�R�bGʔ_9������l�)�On����Ր�J"��>
3<i�K+0��nҽl�����pAYo�4�m1߼�8k��څ@�?���SG�ZcFr��	)ɇ
ŘD0�P� ����v��yַ�u�=2g=�b!���y��=���q�d^!-ضz�*��i=���E�B� ��0!��{����5���@x 3 ����������bZ�TV���*f�@�
��wT�����aAE�<��0F�m���?e�AC
v�Uh+�ʁ2
�>�.Y!6���P�u���o��T�*{�A��ʄvj�	��G�S�9����|nH�y�Q�v�M�:�3@YH��GՈ���c�Vmݛ�� /~)�ļ�gi�!���t-��ޮ�s�����V��O~�?��r��������u`,�/Q�r���[�{�,}^����c}�a��=�3+)9�0�Ȟ"��t~�9ۣ�[sY[��)���M�kMF,�A$�>Ӄ��`�	B�C	Kb��w� ��`_�>0+K�8������M`Y �-lkV��~"��0Ӏ��g�W�,�YWB@�U�%��T�Ñd�G7Eȩ��uf��VN+�Ɔ��Ũ"I.n�-�Ox��ͣТ>#-3f�m���8�0�#���@�i�m�P�,(`���F@D����G	�7�r>p2ȍP��ż[d��)4N�S&
�3VB���5u-��wJ�񄲩H����a,n�n�����/ړ�0���I�ɛ��}��������pRpby�893�p�~���'�~�ɉ�����	���yI<��VO,&jL؞ZO.'&bM�O &�&dL�mp�������&v�u�/K=����vR�FT��ɸ3b.�������]"Cݺs�� �hg���~Ҿ#�%8�W�˔��1,r|Ah�6����TFI��cøP ��z��o}�G7iݗW�v��R�y�X.�'��'O�����L]��N0�����l���Y�~�|���	%�3h]���#�@��_���������7�r�/�"{��B�J~�^����p�*�m��\��ʦ��̰uL��PH �P�}>"M��wr_'��~C��>:�t��ƭ��
ԊYU�ת�K�];�w_c�ACwm�'}m}>ڞ�}?�Ě�ؖ���~���*:X�c�H�rHBf�B��c���(�i"��36����,?�B�8|?Yu����Ť0�TW����դ��a���eα�"]���pJ��5;��"� C/8�L?w���wT]-OU�
�}�GL�Sj��k~˶͐�߉�D:�J������9佌k� DfN���6��r�dH��oE�J�	>iޫ�_o㋣6\����^�\7��ޒ�~�,�:V�Q�rws_{~_���ڻ)/Hߴ΍����b^� T�5H�=E���+\��'"�	�����j���"�N��@_r,<����$��?'�V�6ӗ�Eq�İp�X�:,[�
�t�@��9�f`����+��Hh���r���}v��J���\?�%DI����*V��{������v^\��} ��{��U��99)���l���!f���ipQ�E��PK^�9�P'�KmOӉ� %� ��7���.>Ns�ͳ�A�V�$�e&,p�S�@������\[��>`��-��΁b�X=��<g_�;�8�r�)�	��ȁqe/� �"�4I(򖉧-$�T���洙̄��ϻ������>h�$u���0�y����G������=���rzE���QQ ���B�]��h �`rj�b$��õ�t8����O��t}d�KQ8y��整s�����O
b���9ʁ|(u��$�S0m|C
������A�����֪l��M��B��
��RL�2
�Q�r�G�H��(�wǋ%�(����UX�N$.���G�℁� ��ZΧ7�?�"�`+7�Zе}W��y�ܬ����߀ٖy�1�e��,���L SiB&����;�� �bk��,���K�EX����5�`��sU�ڗn�Nfob��E�A�s:���^~����nm�e�4�o��N�ʡ�����	��i��[������2�^�>ov���Fg�l0�r�~�Q��i7љy�`�A��?��W��~9"x`��&! ���P.2�s&3
���-#�p(V�I"�Ի�H��;YBo�ߡ�Cd���W��k�?#VBr���C��%��k�����V��c�d���a��|f ��L�����\o>Ł蛃w�������Z�̉����J����N��(��zׇ��Fr��s�0��~}R|���z����֏;���Cz"��>I�Qm��8��GӢ!W1��@/��<g��:;�˵"�)���*�4�#p\�PZ��Q�gƜ����='�xc�詿��t �@\9n��ɨ�/m|L�\A�ʇl��\^~��9�Sr#L�:G�p��QY�N[-b�Y�A�y�*M�� ��Q.�,�i���H��:���vME��S�0�?��DpE���V�&��e�����۪Hze�D���,t{�2��-�%d�� �~Pp�hy=[���7ìo����EEٕ�h_/�{�<0��oy:�o�ko�~�\ aV��4"~�<�|��,�KC�t��a��]&�U���!�;ӳ�{����)��;�B{�b^�'"�x�1���s5�k@bS���������89H�ͅ%��>بo�E)�x֓�W����������ď-�}9���/a��Z��
�������K{�}Q�_;��>11'4Z�f9���ӛФ�Z������P&��M�L6�NKh�@B�������wLm,�{�A�cJ?���_�rx�\�hV5����s�8;��d��ٸ�ը�:C�q�E���� �Vj� +�l����|\Q�GA����H�׍���sd� q���(�#Aǹ��^�,���Ҧ+��h4�P�����Z:��ʝ��c�r�����E�Hb��`��-�/qQ�(�tJ#�}O@����Ɏ��`�p��>U��lGbA��R��a��(RzvS�� ��Q�j����E�;E�+п�J�p8@N�Ǡ}�S����~��z�����N-5�ȿ~8���/�2�|\�'�+�Q,������FR�^bu���tOc�E%�Żi�g���b
�������+?Ն��z?݃I�bA��|���{Ӛdxћ?;;_�N�d�D�:5&��nk��!d��v;��B
����ª�2�C�V��>�-}D�R�ꏱ�g���᾿��&^O=^�-���8Rb�cs�xN�%��~t��jS!5�8�,��ԋ``i��d�>�rNm�י-�r��KMu�xj�\A�%[C&�鼱P��"��ݖJ2pߩZ�h�[�# 紒G������o� ��nA������>7\��ܯ:e��ҏ'��n$0�F��d��JG�Pʐ���J�`-J����{���t�к�k7�t�_��^t0���(#����^��aۇ�g�Ȭ��x��}�Y�Zi��/̍w�T
�o�'���e\�t�1�� �^8ޏǮniv�τ�f�4+;i�{��&�唄���q��`F��6����^={�6멋�L�x�x]:Ǆch<oV��: ��t����	 ٻ=��ѳ�(�O���԰!,;V��~�2�EUҼ�EDؐoj��Ļ��>{(i󁘛KJ3�?ۭ�X�}/I }�@��U�s��B&�4��7��E��
}gJ�H(0�K	F|Z�
���Ω�a����
���A�ʴ�jáX)�:a>�d
������'B��Ch���[�#�d�_٪�ӣ,X�=�U�����jKH�c��ȍ.VʒW������m�k�23/�Ѱu�y@k߄{�U�$㋪C7+\[;��7'#(Yƨ�G��+1��A�n�VC�q
�#�现b9��3s�vwf
ILwzB�D�Y�l ��(iv��2qd������\63&���e���҉*�����<%%����E��P�<��rc�x`|ΑV��@l��,�K-�]�L�e�]�j)|�+o�~�+^V���ק��r<�� F`��|�wf�l E2��
 <�S�i�γ>��Hp!Mlϫ������ģ��k{'񑆾���lb���:n^���Y��4���|�rql5h�(wF�D �b?�
l<V�~�}IV���.� �Sn��ޚ�?��lg����fj'�~%��d$[h��Ug�������t[C7��j������� /���~�\6o�0�z�#��Z?��~ F5�.jR���VH;.z�(-i���H�n�yP�:��P�M�:PZ��d��l���O��QR��1�4���!�,��=��͉���="�ZÔ�+Evu�+d�%냍EXc+�o=+�N���U������F�FgO����r��jtqt�R3P�>�y�(E�~uז�\�ʶ '�EM��@p��,�}����3���.>`��,K �r�`��3�(����(nKmn�75iP4�+�akR�#_�[�M����z �Id�
{����͝HV���^�/Տ�.����G�Mzx�����;Y�����xVȣ.f^�����r��~W�{�f�"��+Ly�R��0�gܶ���5��lf�y&VU����/d&�a�ԋ��/7�e1󁴂>K@,ٔ�NIc���2̊��H!�M��d��L٩�eҞ���zו���Lg6�5]��OIynʯ4	�'{Y���+t���nF����6�5R��O�����`hɞ͟�u,GL��X�)o��0�T^j9���!*��۫��Q�Ę'�N`������pn&ESI�
�Y��*��. ����e���6�\~��'
&.8B�'���1��x3�q)�,��k8<��p� @����_�%ӱuI� �^6qz�)p���J.F��~�O�ˢ�l�U��'�.��$���h���Ϩ�S#9a����Z�@�'vW�)�MvN�HMD�K:��S�}���k�O�3�(�k��M�*��A�כHjl+�T ��6T�,��B��#���A�}�!�/�����z�Q��
=8�k4�Q�uf}�;I�6�������/X &$�2C��
k���B����!�.#S�,�>�5����Y��G�6,�6�<�;�<�Fk/o�� 4+}�Mi�ĂN�	6]HCꮹH��_1�S�Ew>�i�}Z�ֽ�`l n_:q�ײ;��Ǌ�����Q[
�ad���RD����Ohl[���@�ཱི}�ID�_XlYN�@�����ub�[&у�]4�)�1�[�2R� �B����"7區�>Y�L�2Lg&�a�$V@}z�V��
�2�d��4]p##
�Qu؀4��c��P��xD	�xX��R��o"�#7p0���/�wi��jG�7v����uޢ8sԡ �'�����j,)�`�M70֬���
4��<����[���&�!����zm�.܃D��W?�B���e�V���y�t�bh�z����<q�]�v�{F���6��X��>T��12+9�op{��y�6װgW)qb&�'��ΞEv4�|�m����s%�(x�"�s��J�4�<"%�p�8Em.;.���K0�����0�7Y!K����FLȬ�(kkgM��5x��X-ƒ��ӭ�"3w��Da��ۘ�$>�'uU����o#m�o��̢%���6HIMȊ&�%�ز���1��5g��%i"��M0�:CV���BO�U�<�@e�5pN�f6w�o��Bi�j�6}��V�L7�	�7$!��yY����`�-��(eТ��u.	�Eh�&�wh��vç���ZL�wY����Y���䨭3R�Eq��7����t��w����W�
�����`�Z}�Ĵx� uG��"���c����#��η�
�y{�^s ]95�,,�	!�/�J^d�j��
y�|�����w�ެa9Vk�Q��	�x��'kEU��\w��.���C�.���	�g1�쒕�c����h���C'Ww�1�(�Z$�\�?��7�؞w��>�_��^�ys4�>�7A!�NE��;���(��U~-�NoRX��dT�t!}��Vz�>���t�%��*Ђ�6��A�`M-��O�ō������t��?��g��*�� �_+SLO?.i�y�Ao�J���v|�X�&-Ђ���m7ڦ�g�F��3[���u5u{�0z
Ӥ�{��yR\}|����ZV�8�!�uF�$�:h3#��9a��*��gU�R�>�̑����@����`��֬��W"s�|h����!ȓ��l��oȖ�d�g�7�@�C��s�w_�'Z�����8޾�C��׬��P��[���P���=A��4`�Yɍ�j,��g�����j��qy�GL����޳3)��>��^ z�7}d[sQ		_6�H¡�V� ����%�K>a��°����@G�����C�h:O߽��0�y��d0O���:[O2
����X�A�,��^H�uۼ�{�`�6L�jN|`B�ѓ��v�X�S=�8�C����ڣW���-�yf9�|�QVX��S�F��ً��}�dX?��Z���K(��	��Zٮ�a��������x��u9kz��M��n��z�*���m^�-X-'���&@�z���J��r��3g��q\[�.�@����؈-%q2�a@�=�F�?�H0�~�;S;��e�f�}6�6�Z�ֳ8��f�Z�ї�(�&}%�3�����5L@G�����(�X�D�>\�l-��r�ų����(,��|����s|����]�<�D [��G�(2S&��3��[��v���E�,]	{�v�z�+m˞�J����G����/��v�N���m�e�4�k--�a�O.�d��d
,�WLޕ����%��e�lAPl��Nu%D�AF�?g��d�*��lA��p׽�J��;W�ݪ�y�ƪ�ʃ�؁��g���b`0]�|�<�=��A�3av}|��xqNk� ��R�쿢4Z:����:�d��z��A:g@!غ0Ҁ�4��E�4&����}Q��b��)���L���,%���h-�~�}X�&�R|�K��x���zX��}HN����)����GjX���h�^�`��(-(�������%@`DvU�Q�k5"'6��i�V�b���R3ux����&��UA�|/�{d�<MOoOX�)T���8�z���>���������Az�جt�6U�}������4>�����YX#e*K�����nk�RU^wq�O	Ɩ �S9Û5�o�vD�(��=ְ/<^�2�^�%O�G����/�t���h(Z�'֓+��&��{[I9��POkbL9�04�	��f�-Bf ��7����h����O��:B�>�n+�P����YM�K�7����=X�G��X:HQ��A��B�oѴk>Mװ���jKȎBK<s���J|�!Zq(���^����߾\cܱJgʕ�\��ި7���j���ئ��|�(���(Ao!��ɗ[��A�N�&����:;>5:}r�'6��.#	�1�=Bl�ϖ�m��]�)�K�&x+�w@�^�8C�<�V��%Rt�P�c�T�� ���������Pz���	eO�.i� R=y�CN�qOx�Ti|�L�=g=aA����Lo[ȫ��M���[���'3��~�r�;a��	0[
-�>�ꄶ%���(�o;�Y6�_Z��r��	��5�+��8؀�W]1�g+������y�S��zKz�B�1�o̵M XK�R�p�2�A�~D� u ��Y=�7�A���k�C�8���Y�
&i[�Ɗ�*�[�p� �冧�|0�)I���"\r��j�(�9u�&Ȕ�p��6O]Zʩ{@N�
|�r3�[s#��p����\�
-@� n�{�}5\�pP91�R���?���;����6���F�a��֞���^d#D2����O��ga�3$a~U�gOZ���h��=���*�#�5��k��;�ec%VW��+���ה�¿dPs+2^��R�ˡ�낇�k�B���'�L`�Cl]���C�d6�b�~M��+-�W�n��g�}7��=D�΋���hh.���Ṹx���ev�*t��e���-L�� �*��R�؍�B"�.=: Ä(-
76k���AWz�!������F���-/n�W� �=��`H`VG�o/[��{�xZ�˂8�����4� !-�lM�Ƨ1���,��;b����� �B�q�a\���T^����!
� F�Ϫ���������}sN?�����^�3�`&��.}\��99��jV�p���٥��.�=1���<�ݚ�Vz�n�'�v�I�	:�D��.#�!v���.Iq���/P�}v�gsP�l|�!F�N]�b�@."��V��|:+�V� kj��b*��CN�r�մ5��o��l�"h���Dd�A��?6@���B6gM�Գ�2�a�%$j(�j�#�����r1���N3eP��o�X��i�YL���m�I��׋mJ��iH��Զ4����?�"�:Zm`�c͛��(����W͎H��/��Nt5')���:���Ǔ��yŨّB���<-���.p-���&����E<���B�&jϩSp�����Ϥ�>�#[mDK�t�Jk�u<���18I`J�J�*�=-�״VI4�MHA���.AiE���>w�P�a��1(�"�g�&��W�ު�Kc|b���|΅r����7}� ����u�T��9�?A�J��{�y+�9�тr��>ِep�2�j6*��Gw �Mv�nw��4�J�+@K��/t^qT�t8yi�ۤ�+�~������S�݂u�+�B��J5�4�녓-�P�E���t&�kZH�Ц���iy�5� �l7¢���]�-y��g�2�ʴ���k��	K���hI^TIcQD�rͺE��C2�G_nֱߝ��<ˠ{j�n�u�.�dX��b�r0������P[�����tV��.��\�*���K���=Vw+����
pX��镸[C�Λf~��w�̾�k$�A��b)�Ӈ�9̓���ع�~�g=_��r�� qT�c����R9*�3�Q���P>���/;`H܆y:�d�\=޸B���u�����4{�el�W�����-	�(�<�e[� l>li��q��q��뾫9��X��<&�pij�%J�4 �+G�v����[�����05�8�-���G�����s��!�+:IXl�Ͻ�z�%��CG*~�0��q�����;W���j�2{s�~�P�'<0~�o�D̖ȷ���9�4%p�LR�B��
�}raX�5��[׋3�\�%�x+O��)ˊ=GR���lQ���Q"� ����q���bC�$�A���U-�wq��آn�2�q���A(�"�M����1��f����.����]��[��a8�����:`���g�زv�%:��O6�B{��d��i�a��K�(������K������h�-�-�^x�r����]�a�K�l�H�Ħ)�������D��%�[���n�m�O �T��<���إ�'hrɥ5�y�ԍ��*e4f����N,Β;�.c8����Ժ�/�#Mz?r���� ��,�Fnaԥ-��.��j9]y���f@5}�]��0�e��W��-+Ӏp�=lإ\	S�+�_1Z�:� ��N�]���c�N�F�}��W
㉇۳�Ij&�[����ʙ���KOH<zTs9�9�DGg�wl�b��Z��WcEx(\�����˕�&� ͢�%c��<�W*dɺ����$�8��6���\�W�'bS�9
Վ�A8��ƏDx�r_nA�;F�mĦ@L�v��|&���8nBW�4RƁ[�C��zIƹ5;�S�)�W��_��h�����P���g�G
�͊m^�����������x�)t�a�b�=S��N���RV�,T��j�tˉ���}�3������Д��4~�ޜ݂zd�o����7�v���L���|��?��4�̬`����<����i��C1|+�v���pf��N����r��S��db^Ԕ��\��;ý��	�F��ڟlO#n���Կ3�ݚ)����Bnn唑qZG�.w�pנ,\\���L]a�m�D�-6�*䇕�k�	JHe��M�����+��e�l�R��pfs�g�'3�D��:V�� ��� ǥ���`V��O2Z"�op&[�NI�R�8!��>��@ؓ�V�����/٘�^$�;��Z���'(��o���u�T8>|m�>�Mp��(�i���qul����lR2a�����I�|{��',w�.�I���'�F3��[���ɪ�Ff�DD�X��qw�Qʜ�k=�)69��Q�^1tՌ��N_�����bK���^���d�U�Z�̘ym�E\Z%Ԟ��}Pn}{FA_�TcjW��P*��$$���<f��9�����)Y����אJ�5�H'��v�Gq���$/�8�}�Ψ�4@-9�oC����:C+��o-��*��5��
��|W�Ŷ@������6s]qwD).c\OV�jȓ�[�Ǹ�R�q�.v�t�T�)e��~�� }\g��A~�]\�¯���?�p��k��?aL+���7o�*�+�5�p~�9�W�:�[�b
�ui����[=e�d�s��z�3��JS=. Itz��%����2��[����2aX�z!�N	�^���p��.�3��$S�Q��=M�?_�)W�z�9�}�o���1���p(H`�NlC�z ��)_/��!�F���JR��H���	������
(���(Mwm� an�`���w�_@)�do�8	���m3≍^�W�I�s�B� q��/�\q�����).mT>gyr���-�va���G��%��[���7,�����4[�ve��]�'7�@.o�̉�E�����3f�R��kr9a����w�J����	�>\�@�p3%������u���[�Z��×�䡇�vH(?�)D�#7�����Ha��s����Xe�R�=�w6�0�=@_����e4����2QV�
V�B,0�]��+�n��.���S
\g�Y����p���L�ƍ�����V#�࿐-ᶵɺ���O{o`UV���+C�~��|$���c�1Z{���SV<5B&hH�h4_���re*w?+BB�)��[G����^x�ٔp+��AY5�Dg��d�O�oRf�C
��-�
�jJ��|a���b���,0���B��2�ɉC��r�\�*�|}s��t�/4��t��� x���i�dҚ��ܞT��*�c��0�銜D��V�0��*� _�h��t��:Yh��O5k�j��oo-������U�չ,��ES�E!d]S�����}Uy����r>sW@�w��'*Y��=Xa6�}nz�/*JW�ԻIF�u���M�V;����Źu����4�a8�f�z�<B�q���b��>����֟��h5u��R�LI�w/��dn�����:E
��r�-k��F������M�mP��S녓��<�E3��[oFS�v�H]UB���A�|ݗ��;=h'�/-x������R��қ�d��H����S����o�ĕ��&a��$Kf�4�3� b�Q�K_h]ɍ�n6�ͬJ�nN19��K��Y�|��I#@r^��xz�~vO��#���d�����-�����������{� 	�N
�F=�J� -yAt*�b�H �rC���EgF�͌͆}���F�������P&6pr�����[�>O�����4�X�&���W�YSB����g�Wt�!���A6}�6mD�x�1��/*k�m������0�8i������tdR}�����U��3��o���?T¿�әdM_Hi��z��&��w��W	`���/�U�//�|=����8N��)P'�+�{d���@�W���� [NfF�y��H��ς�{.�A�!���d�\.��G1��/Ŷ4U�|EV��=iZ3�������v^���[��)B�����v{՛�m�9Fډ%�-����i�1�����1�����hnӲH�y-�= >D��.�ϭ�8�:�9̃3�ҳOM���R,�;!]X綷���ԥ�+�犪l���2�4�(B�s�Hh�����u�B_���{����P���ꔉ����ǚos+�d�cE;��D ����m5�p;�˘.�	�:����������6�l��I�]d�5k�}h�]�&*�څ�ֶs�k�[dRzĴx���#���o�発�T�?妠�Q��O�' z����uN��!��,F�sg�F��wY0�J�	|H앲�VI�}L��i��Q�.d��)����_�i9�Q�^���%�^��R!��]/��m��k���93V�D�ێ-�Ұ����+�>�]�	5{���{t���e�>΃?E�O����n*L����?ܥ�z����g�"24}���ZZJ�@�F�P�]S�"�a�
�{b�� DT��N�w�����i�9����0>MR���B��n�+���zͣ���<���Iᙋ jt@ZS*�OOV���h��g�����Y�WT�_���d�χ��Ơ�����h����1�L�8h�]]4n�j�g.M{u�/�R�U���-�^8%�h��f�Y$$�^�:e�s��`/ۤ�TPQ$QA������ԅn�~ҵ����+D�'��d��$��f^�ǫF�.�P�I�%�=�)I�9A��}��Ն�V����Y`�k����X4�)�^�wG�o�>�Ei4����cw��5���$�=�=3/�uw�¥�xs����آk��H`��Q-d2�h��s6Ƚ�o��oqx{����E/ʸUM��@췥R�J�̟��M`+ie�~�1�h��ۙ�,'|_2'�b;�q�σ��Т�����3���C�A@?y��v�פ���-�Xp�'�m�v�i�&�י��9�0X\хtU�X:EA^�m��r��Yf��I ���V����e]�H�r���\ज़/�i6�a�тI��m5�Ԍ����@�#�0,<�0{�R����P\LY~V0�A��F_���~u׮m�a_�� L�.s6Z\�N1؃qa%�]��^�W\z؂x=��檺d�ooC�,~�V�>���p��T#�Y-3����oE�	��,��U�ݭ�ש!Ţ+����,W_���:W~f�֢t�n�K2��^7�1"�ߞܷ5$�W��V��N3��x8t�$;�\2t}���-HD�����~~vȒu1/��i�_�2)<�y�wf��=�I1���*�A���y��_�u�Q#λ7�s��#�(
A���%�{:�='eDY�K�d�o'V��?�O�Ͳi�I�c[$��6���S]nk�D�}u�"��.>�?\>���u���&�k���م��V�j%Z��i��;��4���ˋ���7�U�1��]�W�l�a�M��G�[�$FU�	�ba��5��<��!v��hiɗ!ۮz2@Ю��bô�\o
9�^mTf<���R-'��[�X�7��qk�Ľ���W�{�Q]w8�6$�=�'�aI����h�l��~`�kf���T�o�p�$��8pHd��>t%!$�JH��H]BV�%���^�ԄBI�n��!|O4:�i��x�WO��}����;�(t�V��(��v�.,�/є�=Mq���D@l�|N"�A/�66HA����z!	�Y��ִ�$����|i���u(�	�W� 
�C�^#@�W��,�,x��`�X
�`��
�`�Xn��F�5�p�M�\\�����Y�B�&����j��TJ{����on$T�@][�9���;	Z$���3��v�I������"�ӊ�o��j���N�4�'s�Ȧ��]�uيt]	�kO7�͗<vQ���T�b��4��`��X�oR��ZSdh%�4�;&��u���6�~"��a5~����� �9�)��4{$Uۀ=i8ϺX`�2lo֪ŏ�X���.�zXO�jI��8D��'띂��C���A�><�d����?N��~Md���=Ip"��$�WK�����v��[��^�t�t����h���!IY���r�{�ԏo�4&�BN*��C1q�a�:6g�^�H2W�ӕ��CT^�é�[Rv� ������"�� ���l.��3��{;y��T��"�_Nq\�<lx=�����^��[��Gx�y3�l�@weԓJt�&�΋T}�Z����T$�'M�X/�sd���������ȣ$����NҪ؞�mH��z�w)O�}��v0ץ_�`�S�پpo��
̬,p�3��r��*��a��a���ݍ�j�Îd~�6m����Z�����8VE��%�؈�o��l�m�@�kX	(��B��5��@�#U�����8�iG�B,��%O���$��x`���l׆�zh�X�\�g�����V�����~,3q�@q@�XN$#���z��FS0-l��,<���*,-�+�Eͯ���o��~.y�j>,��I���l��ٞFW䯧l�ܧVb7�1�aa�z1����O�&�XZ>��aԐӲ*|������4m㑟2�\Ӄ/fo6vg�Vc$�A�n(U��+���L����9!�8����R�6;�L�/��+z�㶹��a���a���	n���Y��G�|=!�)�~r���ĳs�BTc�Jbm����]*k#�?^�1��bB҉�&.U�mD����Z�tp����<f������a��u��K]iح���O���h����;+����q:�U��]H)r 2Ո��l5��cF���]|<	��;�z
>�#@�g��Z1gZ��o�Ǭ�� kD9'��M�V�5����\	@)H3_�!�#����H fN��{k�����ÅP��هi����uA:
��5?L�a���`�J�;�r��eE�Nr�(�J}�%�����!��ּz�a��鳮�[����"�����V�	,��?9nz�|�r��a�ㆃ����э�:���O�	���j�m�j�o�\��6}i��^��8���I�;Ӛ��omP�]�6�yZ�:��CF�4ʂ�g�_���5AӰR#B�<��kww�#y�M�>�`�\�6�V�9��+�:G)����~8�J��+9�oR�)��-���yv<�?�k_Aѯ�e�4�0�i�o���Ny:���+��J{9 u�� ]/{���%�[]�.�R�ޡH�AI-�Ǭ�����P$�q��U���OA�f�k7�5�|�n���E�Qp��;[C����Su$]_w�[�¶V5����Z�����F�J�^��;""���ϝ�o���C���*���}�,���f�9u0~>�X"^��>���s���?�-�`��	�n�5B|B)���)y��:���d'e|��l����.�w�-c��f�y`�K��_91���[��`��ϴo*Z�\�������-F+ێ$btRƫ츖w99��iN��O�
�U���#��3+�=3f"�D�Ӌb� �13x�+�U�]Ʊ(����%K
4-n�	C�
�^�.0X�Ͱ�����E���r��Vl�g�V�������*{o֜����:"nNC,ڭ� �B���������,��9��K����ڿ6\�w!���Q�s@��ի��O�P�,W�����I�0��Z�R�g>#��Z�������IE�vvr@�)`�a������:�zg�)THb�����ܔ�C�ԋ�+5��S�b���XJ��g��g_YF����/ՙ1*�C�P*�=-��=�b?-}{�N�s�fU���#K�Lqo�Vw��z`��,_�Zٛu��M��hm��Vڱf3���z�O:�R�;��S��G;�F���.Mk�l�ƪ��b��
�P�����dKi`>!D݀/�N|�P!�(x[�&��%o2f�cK �X�΀OL"�����lI��,.> �E�g2qFF�ׇs\}�x.��&-d�\9�G3���y�;:��� ��Z��;ݍ�g{e]v#���g��B�B���Ӭ"�I9f�Жq"De��L�������埜��g���F{���+��~�V�O�X1=/�'�F����	%���|(����e��"��>�����C.�����{G�aD��Q��C�}�hZ����u�O<�{�U�I���0lr1��-���aM7�x��*����hLL�� :v�fsˠ����ZH_ɰ�iƚ� ���<Lu���7U�a�9���e�j��"��:��a�R��C%'ᨷ���k�@��V���~�mc�`�>i�o���E�EP�\d
3g�@�>�\��t��z�::�%�@p�_��at�]T\��3�{��-�(��^�T-�8u �0�俧�I��8Y�It�����(_�$���Lp�,ň�e��T�h�<��r�L�� �	�A/D
@�d$
 C� K�0���XPR�*<
`Ձ0�
@� v�Z�A�\8
 ���(�]y9c[@b1$�)�aE�A�D�?.$xWly��\A|�E�?n6)Ҩ��բ]0
t��GYt���-��g[��#��>�+�� ���_��ص����¿����X�ߺ��`�,�m�{�XP��H1�_�[Q �,��E�k��eJ��
=k��!i�n� `c�mI0�� �,�h$����h����N�Dc{��M�G�
��X�p~�]�qC����$���N��v}}�Д�5u|��@�Cࣹ���I!�I�D�Z�#��I�ԗ-��)�Nd!�d��ADd�L�#��+k=٘G:�6Em�[�*+k��;j0�p��U�1Ӆ��QT�u��Q3ji
���$�kGT(T�l�x����J8�iC��
Ӂ�v�=
��S�"�q��-�ŷs�!��N��qf\Z����������٧�n�Z>����,����&�<{B©kUb�6@�$�Q�R����X�"���+c1�i��Yu��;?�#�i��2ӕ���>f���ޫq����D��˨V֨Y���ݹO�:�r�����Gf��}Nc����&[G����ٝ��ٙH�H���NMR!X,E��"�7Z�F�;����b�z5���]��#�Ԡi�3�Y��J�x1C?�kU3�Yl>���q��cSc< �1�=�!!��w!6��<Ha�6�xh}�����zKV=~���">�{\�?_FӐ�Fj�D󸙿"�v�D�#�H��&�����ֈ V�t�+E���<!��L�n�Ƀ��ָ
G!Bt$��>13c�.����#�70�������E��LR"9�
H�ARn��j{�:o���֗G���P��k�W���j��`���ڽ˹�2�����l�0;�U껸af�2���ߛ�.t���	�X[\��~q�N�M�����/�|�-��}y$�{j;P���{u��+�p��^���6��L�]z�!C�3,���������ųD�&�=1� �I�>�iŪ1#g�#��w[O,����e�����^�6�P�
1I���騖�x9�D���5�8e1�̡-Co�阗�6�NH+L`��*=)+�s��0�KDS�(ӒU1���?0(;�]��ƛ�xKf�} ���3(/�b(3�A:�<�ܵ/��3Ԥ0"�6ԨB��mY������ ���uN`S��S�\=W�i�@�3��U"ճv�r)1��V1!�)�{o�{	�V�G��wl���=��sU��MC�����th:}:�ͯQ�]H��JY��x��\�:�c�5-"}�J����JX�q9��,�y��,��}��@��M�X;gun��e�a����j��E���hZb�:��Z�gy�<\�l��1��d-��p�-����͓�5�jE�!ng,F��T�̺�>���mLH5@�;6�}��}�jԀ��v�_?�L=�U��y0~bp���#|�g��ۋ -:�����d`$�ܽ�O�6-We����)?��l6mKJ=���V�sM������ J�p������@`H�N'������#V��J��&��~NR��F/���<q��{N�#~_>J��s�����h@ln�7&����~%�T+5E
T�P>k����N�T�W�gX+�|sr���oX?�|c�\���ݤ?��%�^���e�d��.�D�����;��]+Xb�=9��3V&{A�)⍎[�եC�nv��� ���
b�Jb��A�Pܡ�A%J
(tP������Ae JH����cMWʥ=P�+TRDiՊ��r�A�OB�8�k��� ' �~�����yi�L�;38)E��S�����GVڗI[f��A��f.^�Sv�OOL���]%�_2f:�i���t״���6�\b'������V����VV��}�(R�  ��>켉ظs&`�ʝy|�l��󷡐¾ՠ���_�S	�,���MB{��U��V�C[	W�����AqS�Ze_$��tg�,́4�Y����}�P�0$=�I�]���7�� CeN�!I!��`t����/��E���f?�9�I#6�j�����h��h#����{h6�5We8�qn� ��r���"Q�a?P�5W��U2G�1l�Ƃ��˜|���Us�6#��lF�l�}���MX�>nEn�aA�;���n]��s$g��a`�CgڿU�C�N	��!+Q��sV߫��}�AP]�,�d���T���Φ�����g���e�^%[���z�'���'E$sW�x�<���  tL���z�u2��M�m���_G�J,̡�������`���'#�̶�[��wBî+c��r'(t�`����JR�?���68Ă��5)֝��˂9���A/�k���f�w�*)�@CL�B���͔�����l��>��$w�16�-}��al,���dj|%h���6�o[룯y�A钮��Σ���d��J�b?�B6����� ܃�,�6�U�^�4�SZ=XrVk�s�Q���3 �1��dI�xf��;="V�@�P@T�T!�O� �>u��zc?�ދ�~$#������Vt��z���\�:��̭휊D�����j`����laT�K:���Tî�/g�[~�R�~��v�(�T*L
K��AQ��l���t]��y@w�M��F��X.�*mP(������`�À�Y��`[������
0B[::�|ؔ����Ą� �q��q�(�����P��G��M ��� �p�{`>4'B���R��2'��GC��yq���i�� |�-5��p�]!�z4�$�I��%�OU����QXi�`q�h���בy
c/����/_�(f�ӊ�o|f�H�N'�@��tԸɓ��������RYr�o(7�I1>��.�׈�؂�3�nb�xP��N�g`� �4�%`� ��� 咆���թ`ͬ������D ��!��!�;#dp������O|��a�ؒXa�hc&��8�=G���vsz�w䭧��5��#Ro~p�#���*�>�ub%GG���Q[��,`����	ݜ_ol��S^;A�fF�F|��(�A���Z�-�CIa��(�[�]�`?��g듩�G�)l���K�6��3�4��B}l>�����ZbZ)p<sh��B���93"�ڍ4{��_q
�*��|�~��7L���up����R��h|��dQ�΅d4.�mP���p�f�{X����>�<ђtk��//�wzb��]̇��&�������� މx��|
�����x��T���;�v�X��=�₵�����=&�"S[eR������@?��:k���	M���۠���f�{Ć�����ꏢ/��JfJ�+�0|�5@&-W��(�������M���Uz�gWh�0/��U�ʟ�Nw�v��}�6 �ʠ(�YS�I����T�����r�����b�O	����B�͟*3A�9T%Ʃ4�%ʆ��-��{��`���Rfq�箲_�k��e#��)�x}��K��%�8�lq���v<�q�jh��6���\���s�TM��
T����
�*�߀z�ط�g���4YG8����0���>�R�`��T�0��_A��/��;�,�p	��\�������F��{ށ��T`�9Og��7���=ts0Bȟ3ӓ�e����B��[���gլ�f|�r��n��8} )�`����:@%�S�lS(G<Ф�*[���xjJ���W��ƭ�z�g'���&��Z��t�<g�S�s�+��{��4�m�T�}��
[T�w-ut��qI�_.����[�7�~�\�)�l�q��3���X|����eh�eh���Ǖ��B���J�7�2S�ys�������gp�l��?h�>��L~2���9�̡�6]'{m�{���ޱc���Q�x>2_.���%@��K~ �� .���7�^�� ��pO[�M|��@l�N�I����1 ��fЀg�7��"A��������U�z�'����z��n���A͸r���|�B���!�&���$�EB��I�wo�5̡��������ɝoo��XK5f�*+��!c҆��f�Y��T &��Ro7:%+2�'N��z��&�%1%���Ь�9^�[>�2%� -���t;!�n�h�j��ݟ&]l��]F`]�R�U���ԉ#�X�)vx!ɕ��<��@��C���9"`R`��˃2��`��Ob���<w�����]��+�N�\O �]^�	��tͫ�ϡ$�ڐ<�ݤ�s�����ڧ"�0�Q{Ȁ
I(���_˵�=���˿���7�����M���ߗ��a����tT�D(�
S)�V�S;��D7o]��H^&|����%�D==|Q&^JY6DU>�}�~�-J��8ӄM� n7jg)%?n��y*��&a��_c�}4Ǜ�Q�b��#�!��7�&��^����T��=.R7�s��s�|̐@��>�Hm��O��Di��9R�=��A�9��=�m=M�|'O���2�?	�̩�j@	�J-�P������A;8�?n�y���.R0�ƚD���9g��������T�(y�+�Hy�#	�p�3|7��F�_��A�:V^����M��&�LI����t��Le��S<�a������	6 V�zgZd����^U�:����n��>��Q���Q�t�Q+)�&+b'R	���p�sU�|ڟ�a��!��Y����'�T̟a%�/	�F��I�@|}ct�;H����t�����UNU��`� ;i�4�?��9¥yEf��A`��P��G��t$9�4�t��[�0m��g��<;��j�k��e�;��Yz�b���B��}m4�ڣ�<Efx�HA���� K�����O��'N\�a�]������1w��z�	��n8�M@Lܤ��#�9�ɩ�)��^���FV�(�2�z��+���q#`�·�|���k�K������|K�n&�@�E��M��n�k��z!2W�^!����j�Sd�4ЉX���-l>7G�ZC�%#���M�F���nwA����H���jYS�/��
�\����Ȭ�&���x5m�/
��e���}=OS�o4s<:7�[`�0ub���i1v#���1ϊ��a���霱.Up��$������[�0�"����+��U���g��v�nh0���"|´=W�8��.-M������9(|�&����%�cW��"u ��pb��нP9�5�r�#�(��o
W�����Ú�{��j����sR� �SҬ~B�f��Ӊ���5�����Lc��4��]��J$�҉W��R����݄2W��T�� �tO�S{jS�^)�؅���c=�g�C�+1��?�~9S�f�|
�R��z�K���6-T.A�6_WrE�[�X^m(����3Q�XT�G�%\���Nc�˖#$���
�:jV)@_�3��#���	����*�-�>,}���a���h�ݍ�&���әV�Ÿ�")�	X
�fU��i�������"�6bJ��*)(�Z!͈��3�~�=��Q'1�(} ��\��d*�V��O=!����a��K�`�^��.p\�㈀j�.�"�д}�P�%t���%]���Ss�o��ɢOx�;�5&�+w;�P{���B���
�+���Ɲ��<W@�����⏞+�N�����I�Ts3]�"d�F�ެ�����]A�~f(h��>����Oa|�m�'a�զ��]�&����7c�جf�L�R?9��j�ɡ��N3�S��v�,�qn�X:!r]w����zm�&|�lM���U*�{���L��D��J�J��z�6/?��A^���8;�nގ�g`���y��E�X���V��_�<���Q�yg�&������^:�_67?ⅆ�L�g���G�h��aIo>�0��A���L`i%>�l()���,Q��Ź$���E$d4)���lN��.@=�ag��)Ag�_7/~�/c��F�%G>O"��/Ⱦ<�a'�jn���(M8b����*ǭ��⡦��X����KG��\�7&�T�y#ԁ���ch�������O;SLd�Y̸������w�;���z�� ���̎���gS�������lU�߷��]G?�����b���E��E�	�T3��r�l����[�Qu-E��Ԙ���� ��g*.�5j�E���PP��͊�t��s�Y������N.�{t�����e��z�up:�l��b�}�*�5���nyb�QT�[.x���]�Q�쒹����7=�{�Q�e��T�CY�W 2f�B5dME���8k\�U&)ǣ�g�oڡ5v; W*��>jqE8t]��0�@��s�΀�@+��B�y���s�Zk�E��1nVs���_;�\~b�.Ձ�a�Z%��V~�F�,�֒��5�]{Ǜa�_x�4�|E=Y��r/PT����*E��V�8�}��ͨ��dL�����b�qy�F�fk��}��	qd����EL����m����4���JEI2�R)�oz��Yð��,�3�#N4�S���@p�2�W���0Y��4U���kJ�+�]��X����^V��?Ҩt[�3Cz���PW���!��7b	;��3�2�-�:�x��t�)�W��7U�G޼B=�t���F*L�Y^)���}�X< ��y����3�Ş�^���0y1�XK�FY�,[ gd�����eE!�ww�ru�T��0
�x���Nޅ9T�i��Ґ��ٌQsB���*n�V�t��MS�g�x�'WVs��A�JFzs�<���j��qF/c�yq�'�g�G�fK-���ޟ]�Cx��h@5�ʄ�hsn4�BP���A�`�ߓw�=W�v���r����N�#��)Ԏ��UT�K�3-	�֤o�@��<]�`�$�އ>���fq�����c+�w��z擈xa1D����$-{
���=���a/1���s��I��A��u�#�@��a��(T|���X&�����[��-'����"? pv��~%o�9��<�J$�drbx��B�/�ɣ�x8�?J�%�9�����5"�\�9t	��u"?���k�.�l���5]`V�Ye���""#-��?�&5�f�{j�yU�P�%0�#}����Zv�����[���Z�uA���6~<$:{|f`���q<��c�N���$�{:���J4}�B��`{�y7���<�d:��s
d��!�o=/�t-��;�"?6W�P@���{\>�m����}���
��;+uk�U[����o$A{~P�v���ŷ���NKe���2���������W�VF�X��@�F��3%���q��g	v�]x�U���	_�٭$����x�1��a1�qҭ'��>5������g�o��q�������HH9mP����91����d^���|[�me�V{	��ƪ�w�ə��F$.�K6�-���@�_?u
�p�jVz�cW�H}r�'-=ⲿY�OIc�U���@0[�	�U�XJao��-\�M������ƥM��\q��m�̙'��>�ɜ��NGC4���r9�lZ�F�)'	K ��Q������C3qmoy~("�I�x���:�bT����f��:���b��ϾX��
�=zR�zq1�M;���N��M�B���?al�o��"���������,e���c;���:@Ez>�h�$4�%��AFD��V����b?��/UV������VC�Y7]��B���}Q�Lp?^W�#R��4�����	>�Ӌ�Ԁ^����&�x�8�vG�.��9)>�7.\Ҳ,n%�;��(N���8<��E`,2SK���	�2h,\�HѾ�h!Іe�`�'���k�l��<�C�;B5����͟�
 ��ᓌ=w6$n����8���R��ގRޅ{!9�9xX�<Zv����/�'�7�Գ���=7�$�I.Ľ,�,���̷��Y�XA+�>�p���m�v�u�9e������
���]���v�N���ik��&�2�����)^��o�H��R�:�9�:I,x=D����'�D|���Ƹ}�	<7�@~A�/#�w�V�	6��:�r�ש��'9�Lr��R�����.1d�X�pl%/���5x�o��4m�6����M�@�:����iN����]W;�uo2���Ä	�
/̏�	'ac/��$E��"���&����D9q��m�h��Y �m1��(8>�<��9D�W��Z����@��<��?��H`��g�$���"�����$�=*��|��bȥ�!�Ԗ����CJO\-U�3�e(�����Ȳ=P�'i�;�@�==����_���idPb����`����ݮ}=����^\��"ϥ��|B�\���j�ݳ�2�Q�Λ���}�����hb?����g|n�p��&�����pNg�u�"��Eo�����-X�ΝUP� �
,D�~A����O��k�,mfx]�YҎ���t�H�c�ٗ/<�O��j%AO�s��$�2�@�!G�cT$���|�/��'�c�7N��;v���\��O6`
	�p����~a��9u�^�$�<,D���S��=,�L:%�kf����xα?i给��9ˉ��u�����%M��$�k��!��<H�S��}r�-CMo���)� �"o� �q�^Bj�ϗ�&4Sbh/0��-!���9�!ŕ%��O�"�0�հ�eL�cB�rd`�S��-K�Ͷ�f0V��M4����?�?��Y.&ͽ���D�3���U��E�!$��>��I�^�SzI��d�����1�T����\=c^�S�>sn��]���vA�g4��eP,�-g�%�S�����a��=|O������:�2�V^�h�$��}�݈I]=��{�ܿ��,T���_���TR�T�e�.�{����w�qҔ3{���W�;�h�R��$��B�}�f�SǱ���l��7om�:��0�w@U,�Zw��N�{��WX�C	���rgs����T�Gbf}�������#+��F�,�W�p��kl�0�� xG��r☐DtRpH\���:LQ�>3�a����O[C'�É�c ��!U�(��t�E&C�5~�|&j#�OX�j���<f��-���~g[�]��	�Of���5���r+��~WL����D@L@:�Ľ����M<��ɘ�7�����ov�5�w��޺����z�k�E5��M~�lm�I<�~�Y���0ӻn�w��']ͷ��ey�篏�-���b�|	�����H��4����4��	����r�G�ʹ�W�2�
��K�gLc�7�g���\�5IʔL�E_���c�O���>�=�אݐ��������sr�K�J�w���˱x�#����~��4�3#S����7�JZ��� ��a�k��_��)���Հ�w��Zt�(�5y�������՜k�_�SU�ڎ�s�i����Q�Ý����^�ZE�	4�V��_.UM�dZى4>���q!���)�g���|)��y*b�O���ypzhJ�%�&�X��+���UH��9�� ��Q:�WV<���HP91�p�Y#0m�k�$2�*�juWK.��1a�6wض2��tp,��3%�
jm�*S%1����{	�Aк$��k�s��=�W����Z�W�Q��B�%�ň��ժ��uKC�p(�\��G2�l]�j�䒓�+9;M}��\,Ț �~^��Յ�6�%"��V,|͊U���K-F���T>��5'di��EI!چ0��d� �CA*�2����RwR��5�9qEB�}�P�B�$�Ձž�P������[���R�>'�2���!���<+	�f�;t���'t��N3ac��R
�¯󉣾'�F9��L̄���D&!�Ă�Z�w����:'�dӼ�d! �MWW����.Z�h�A���y��G����^���R�O�Y5+`�f�iE] ��P����HN����R8��w|��w�����k��'�`�Wm������m�Ɩ�����%w�{�(�B�A�e�����*��l
���i��P"���x��E���[�J�ۨ*{�xv��e@�.$𵨉	XSHb\�}�*$���4�9pS&� �?����a�D;K��v��xW(��)�1��11��������t�1�G#y�D?�<'�\��ɭ�֨na̘�VF��CA���N\�f[)*�M�����RJ!r�҈\�/���U��l��@�Mَ���>n�"&�½>��a)�&M����e�B���-�
����k,Д�BӠ����أ��ʗ+p1�u�ˊҺ�BqF˳�
lF�Y�/��0&H�
m(�A>5�-�Y�}��QU�����.-�Y9Wg��ݡ�S���q�V�W��7�H�i�۬�i!�5��El>�HZ���l@��.��/�e5@d����c�.G$i�k~D�/UB(��E�Z�[>���&���t�F�>p	{J��D�����߷?U'	��DJ���s�9��]v�-rŭ�o�$��MS���{#A�a�kqD$�tG4�^v��$Q��`��V��$L�CJ�k;*a�k!�ld�F�1�`͹���Ay����W]��b��K*;�]%�_�֓?PA�NK2H^��9��$�Ok�.�q�i��C.날xK�:?�)���H�.\���rV��;!ٺ��c@^�k0�ka��b���k�J$��Ɨ4=Lb	:�j�ʌ�u���lh��<�7���E_��j
jϽgA��HNN�3�(�)��
fn*Ǒ
k�����D�������
��&v8h�C�UU��n�ȳ�+�����E��|[�v�U+�bhx�)�P�ޏ�W�X��N�#b\�r��ǻ!���7������gj��*��sM�5��}�fg���M'&ɽ�/A:���^J��[�<���a����	O��W��(2�Ĥ�Mxm�9�E<�w�\Q��D]����Op�g��ٝ/bkY�j�%�����y	�^Ey�m� ���6��q$�1�˟�f�ȗ�̢�}^��:�uW��V[��G��5/�ʔ^-7�ϥ�ʨZ�	�o��U`>W¿����q����_��Ie!8�hY\���ξ�|�@?D�4�C�c�|�)�yWKo�i���7��M�jB���H�G�>oe1T�y��F���C�Z�XB5"�BZ�}�D������B�o�>L�����G�����������-̉������l(r6s%x/�qU���$.�ࣥv�����Fr��)+C���O¤��a�h�k���{�Q�\?9B�_�x�Fej�S7Q��������]��P��,%f�\���>�e���p�+�t��S��ʘ�y�ֳ�
�v�@6f���<�W��]������:��?�Yx���,��?�xoQ} �t����;�o�cO�CH�j<���+\<ycW)��f�3�8*Ŝ�}߇��{�Y�HI
���G�mc��dDv��lZ%���m��r���7R$���x�d���m�9/�]Ťc]�������_&�{HZa��Nμ���7����4h_�b�ۂiHJ)Jԗ[���5��ۜN�RHL$?����������<w�P\Њܽ��n�hEЉ�I���Ț�KFrj�����i��P���J6��W��L�+E�gx?+��1��jgԕ�������4s^���ExЀ�dj<럏���]�Բ?Lw���T��R����زS��駶/�l5��As�g��E٬��d'ƥx���fxc�Ջ�),^*�u��A�:U�6�V�g��%� L�3�4&��7o6��KkU�����y���s�ִ�ln��wa��1�Ȃ�����Q2���W�m���a|�;20/�Q�;�h����G��k?3�yQgI��t�/p� 1��'�-q��\�`�bc<6og���<_ܳ QF�����L0�-������@�� ���s��<�E<���g`�ٚ�d"Û%�C�{��BpJ�93u�Ȥ�����4���¦ZѾPv4Ѥ���Y��ޞ�W���ZE�"���hS �挛V��S��a@���u�n���@%� 8��k��k�+L�#&���M�B�e��d � �PR�9c	�
@,}�"2$�p���r��@��b��)4��ti�R�V|�F.��
���l��������K4��$�߶�!���_pqG���+*�pVu^��?�_:�l�
��m�z����7pzs�G����G"�6ͼ^��v� �y�ke��8!�v6�k��>�r�ϐ��L��m�3�� o�����(�������n�xSj�(�w��'4ٺ�^�M,��)�|.�ta�lw�i��tb�0
��Lk8�0��zzp҉?r���!ޞ��4��u��=?:,D֫�ϭA��r��R��Q��+ ��ګ8C�iR�O���G<�8\���&A.�C\k>YA��Bk��?҈s0�E���J44a����pÌ'TH�]� �AϞ��Ȳ/�W���z�ô7Xj���JJ�|�%�w =e*[���V���ƭ߄j�Z�/��Em_�Ϧ��x'E����̫���`5y��K�+�)��\�o/�f��=�9�$s��t�Ū���0^V۩h�H-Qo�8W,)A�i��,�yv	�����)W�oO=DdgY��L�]&�pd������mJ��Ig� �~�Q����?��Z�)Ϛ�v��'o�ws�,�f�Dygs��֟�K���8|9
���y�����>'}(�ؒs�L�v�2t7�ҿ����;,!�5���~�c�Gŕc�6��|���G0��ꡠu)��N��y��-q��3�����-�B#l�����H>V���#g$�o�����ބ��
 ( [^�t�"�����}���Yz�e��v�rq�l׭'��ayJ�9�u�������`D��M���M18lU�D~;�i��&7|�KyK���E񄛉`�����/�|ꨲ�ե����qA^�4�;��l��Ȍ$�&9���բ��	����z�|U4_Z]���x�c���>L�̃��u17}����Ү�~�
i$��C��2��y���ڎ�|�[hqk�ӹ&g���2�o���P��$i �U?�#�3w
+c'[��>](G^B��$�����n5~=�y3K��w��i4�/t��c�S�K`��fH.�*�Fޯ�������|�p��!�����2J��:�́#fu`>�ʡ�	٫v�}='��l?�^���^Ð"c�<��N@��#03��e����Jw�1!ߪH���xW.U�Wr}��w`4��O�z	�``�G�#��ꏟ#=����L���zȨ�@j��Q����2��voᆰ"����s'�o���NUy<��=���3�\�X�wp<KdO76ԋ�m)�k,�?K_�E�N���#m���/>���"ֲ�4�<��ݍr L�����2U���Z^���vc��ԛY���X6��,��È+V�p���U��clJ���2y�>?P
^67˷��a���T�7鋗�������E+̢,t�������F�XRїm�d��⻌�Եß-���Η�57[�P�@z�r/%��\�7n�9�U�E
W�
sGr�V����S����۪Z׸F;3��5�� �o$�����^���e�SU��wH��M7��D��
����o�S����@�+���s�ȿ6���1]wQ�F�/K�Z@�
��ր~Zʪ�#z3s+}$��4��?B]���m%п�@THnV��3��S�V���zwg��t����w�d�3y��I�j[�,l�����踟a$�����ݫ��Şt\�[�s�b�Tu���+1�_�Ѻ!RY��+C��y�W��*-Y�?�hy֣����C�����qw�cA���g�X��#��� �GFt�G?�vz�����Q1�eIß���bu���_�A�6
f��m�"-t�T��!c�Ő1�ɮKb�hg�AS�A��O��_P�M5@��Y�7X���<�_�0_���U���F)!\�}��4�-V�0���/.:/���S����(B�h.e�Q\� �~ЯS_H���Sx���U���_Im ���믊y�J32����}��?�/�H�l���޹�k)���uPw�����v�J7wZ�p�Kh�4����.M�3�6�E>/��aHv��c]�.���}�~$���v_�����]oL�O���l�rP_tx��k��9T�Н���56f�W{�w�D���P�y�G��3��5�����}�Md����3�=)^�j�����*7;��"%t��'��\���P�;�;1��DҴ4����FT#�#�
4��9I��4J_���Kܲ��}�K�U�6K�Y�^����ҍ���]ƙ������?5�����UH�y��)���� �-v`�/z�z�#��u�^��ׄ������`|��	J��r��u�����8���1��!�|ukr?��:�%����0Uռ���gnm_/O��s�糘�������i��W�� ���\�?{1�G?�,��S��Isr��$�e)�^Ч����H����69�6N�'T%I��N�Oy�0�Y�р=ߙ/ˌ�u��E!m�
��sşd�nNv��r�c�|�_
c1d�+&����`Єd��Q����Q<�w����#9f[���uXR��y���F������\��F]/��������o�)�+�*]�}�c*F�4-�F>������e)����K��G�­�F�gj��K�߇5!��єte���p��� O��c�c���`��3�&�
��WWLK���c��WkR����>R��{ӆe2%�c$l�����4U��`cx�5���q�L�"}H�x��Q��l�D0K�	��v3��Z��M�Ε�b+�Z��ŧ�I��nXFr�ud(�U*v���B,ǐٶ�s�TD���T3�S��p�i&���&Z���*O�0�wH\o�a|�k��=�1����)~��|a]8Y��W��tY'O�/`��1�0X��O��>*�����(�6i2����v�,��RP�ɜ��+���ubp��gm��՟c4�=к���<�O.ҩ�%�<���nLZ��t�t2J�x�Be)�,�|�	�B�+.��&%�0�dh���]5���;�Oe�-�伽Qۃ�|�,�2;o哢�E��m&a���	��Wl�����������W�@���~�qAAt��>+�(��6��ڬP�	�p��8�������%��y$�Ӳ�c���������֊qc'h��=)��<�BA�fƚ(�c�f�q�K2��X.E�`��oH��1�E9pf�3�O��qN���V�X"�Qt���u�#:�� �'��ʋ�����>7!v6G�SW�f�yrk��k�|,�l:��(6�JM�1a]����'c�ҵt�F1H�@�M�a(�ߐ�T�s�N*��9Dev�~�դ�B�g��
fN���H1&���/�m�`P���W��a3=�Q��b)لDRa���ʵ�9�l����>^6g�wҒ�e��Fm�]
������]�����z�ڎ�/�L�\�P�}W��P{�-����#��(9"e^
7~.?,���������OP61e��)	������=δ�ݔ����1��,u��]:o�D�H�W)�s���02vۈ�l��_�ʱh���\��}z�۱�ӝ��NS*��i��Ԩ�!Cu5�@k��X_v�3��<ت%UEhIŤ�|`�.�l�m�Nq�i*h�X^9�=�v�5嬷��Q�:�*�U߯�U1*��Dwgs��6�����EAd�t�9�ſ�*S��^X�YK�%�����4L���@r(�YZ��8[fͻ?쎁��V�s�	���I@�x�i'�p�KQ�זMn�TͰ����Y�1W��SF�ۑ��N����g<L�����JkZ�*�{�U	xL�k��f�V���]+mͿ� N\���#�"ܪ�YO&Dl8�L���T��{���+7�d���l�O��4U�#�5m_k*����c��K~ύ�#ivR�T�})O���$�/���b
ʹy^c��t\�q��&7�Ms��j�u�:��h�rG���x�A+�c�^�����ʨ�T�z!e��Z�bQ�39Y����,��g=h��&(���x�<�-_�ս9/���곢��2�
���Q�F
�$��kC�+���g֔��M�Jǔw`������\�0 J�L�:������S��]�Gr;���|��x�^"ZB~ܕt�K�:WG)fy[�n#s��%���� A}ĉ�'bO<�c�X��Ŧ�>�%jƻ�W�T��-��VG��gR���0��RbV?�Hk�a)Z��!IF<�+���&r�5���:�N���Zw���j��
��|���N��R�nFj&��R��D��xx8;/V=Q-�D�770'��m�Z��tI����p�\A�����e��_8�ƪa��⦐�j�-��f�9w�RS*Zk�N��@
��x%i���f�k=�������/�Q�1Ɯl��&�H��dB[��Y'�>�Y&�>[�ȹA�7z�gM��.�����Hi>ys<w'����i��IF<��F�91s��s�hJ�;T���z~%l�vAٻ������n���m�����M�@�0-4�#�~^"e����@JJ�Ut]��q�h����Q��r0Mn��Q�,��cO�5*P�*���U&�[� } >�~���{�Tu�(�����d�����J��I6T>�a3ON�t��Ǒ�L�3��& 0��x��ct�)W:@��p[��N@`�96%S`R��]t��葯b�%�Ґ��b��Z�w�@L��<��ɏ�K�)I���*�x�^`7��:��%GJ)��1N%nQ�T�����=�T�����x�;�T�7t��|	4	��;�vMΌ��@��.�6�?�>���0����?ñ���;�W�+��=��Nd�5x��M�׍��֪?wK.��JhR�u�<8�k�`V��o�d��w�&�R?�R�|���a�[��V���W(��d�FsJ��*�a���O���:�-�Ws��Z\x�8���L(ȃI�R�<�u���G+q�c�s�lF�K$���m��q�Ī+R�i�]�� ���S�ŒX�;'�Va`��̤�{�r7�!5�gE���m7AɄ��V�q���N(7E���b�?;�޶6�ն��<��S2�τ�TV�z}����i}���v2��"�6n�F@Ēi��;����s�>�����O_Ӹȿ�>S�����Pz�9����#�	��	��.4�gX��=-��	���"�K���%s����#�-�	L�~a�ݹ�7s%��dm6�Ux)+H%�W.���Ȟ#Bi�(�r�a�u�=���W��5yo���l��\����j��f�@�Ik,��8���Y�=`Ā�1�#c���040��3u�޷�D5��`�����`�V�d3/W�L�����	��`>��b�E��_��8:87=R��=v�^��%���|H�j��.���Ot���]]b�ˌ��~G4�'�8�DĻ�bڭ!�S���	ց�t�Q)R	bt�z{f�6(��[�����rTG�ąpt=|���G��7���@�B�):xNvߠ�7�Qz�"����� ����a�z����t����sVփX ��߱0n�����+��Zp�lOZ�=�6�L�*ʟE�%C"� $�@/ᐰ����15���Iq�	���� �����P ��B�, %8��<��u��ώ1�ܓ���{�֛���	h P��; �� /	{�)�X�/�Q��P��;������#_��1�Ix�p�i����^�����e���E����iS���}�j���f�SL[���	o�s�}��.�u��l�o�zӴ>�X��I*���-��L���S�Xj�����צ�J��#��q�ޡ��B�	 `@B���l�z�v��a�g�Ȟiw>N`�4l �9����H}��m��ڈ�Y6����6����CM-A={�Q�T-ti#޹m�P?W�T�Q��6��a�'1�ڜ������g�v��<���o"ˑoV�)��?Ʋ���'5�pK�|d@ r��^��ú��3ɺ�w(�T�;�ܔ��"K��.$d����(-z�3;*U�f��1�����dX"K��YqXjh7�����;�=�l�䈊���#ڏ蘿��v����4�#Γӣ�V$2{��^��k�e�\\V�M-�~����T�v�/�!�aI���o���2���;�YU���%�h��U�����UDO6��%�������>������l0��=����Ø�dIm�_�e|��sf@@�%z�D��LB�����S��0�3�ㅇ��nǺ�is�D@�EHg҈%qjS�PE&�G(��˒ے��	x��=��R�^�(}m���Y8؋�Rp}7?ve5�p^ӿ�B7������w��'��&��@�b�:�v
i��]o؋���Y�}*I�d]�[�W��+��>q���1���*�œCş�6͉�1�R�m^��p�x��9Zk�VpMi��K�+�Imk{>:����2IOfˉ�\�R��F���G'%�t�=ý��w�������go��2��	"�U�D�@)��񌻲��w%����dV:(�J��w��k��_O�o&)+J�K����M3Q��r�'��5]{K�-�{h�5�tG��,�y$�ľ*����1��4h���K�}_��e����%MBW[�AZ��^,:3��HP����(<mޏ�B=���`�zf�0rOa�6`k@�� 7n�����:7�'����R�z8��H��w}f=��(� �O0�P5/�DQݣ1��?����r��X���wN1p� �Y��iu���H�����i����Q�74wrD��)�w�æ��yl�T�Q��I�������q9��b�Pu�P�Ӊ9{��!|�����!�Q�Q�RR@/���`o><�]Mh����@�Ԯ������n�Y{��ӕ�q���t�q!���E� ]��!�c�:��I��j�F5K�V��|@�����s��},���9 _�+��JG���.���VP��~�<��k��,{]{���b��{J�J�&;�D�M_)�T�/�x�h>ү��D$t�I�/�j2���Z�.��w�#i�}���߱���0�nd6�L��6��%j���D�ɑ>fC�.5���f�U�.���#`ǿk<	�g���I|`X�ނ᭾N�mv��R	���
EaKYdQ:Q���F�#��7�\{h���3�t:���qμ�����"Z�{�&Fv��L���̗K�����"7�u�a����P��2���}]9�ol�������x@Ծ�,~ ��Fg��nu�׉���I������R$i-�Q
�JI����(䝆fIZ�F�qD��>ݼS`I|?��"�5G1�Y���D�.ڝ����x���mn�C�U�ة���<���I�������@�A]�8x�(5N(���������*���'�pF2��r���z7E��X���gs�[�qa�K�p�����*W��x�74����׃���rįϖ��:������׃ӦL�q�<�{�:{��Q����^�0Չ�`O�ŉ%�Xq���*m'�v�"ݘK�_o��"_/��y� j.CV"S▖��W,��]�a�̈�1NH�����h@z�)	��n�:�0���^�g��E
�eHk�wU�y�
��Y�l� {+~I1������^�`	���&��+���<����Hk`�o�V���J��-�����+��Ӕ�n@���3�G��6hAr�L>iB��i�D(UN�8����A�1z�7,�"o��Akإ�{+�2$���LʘJ�C3DM���c�m[5���4� �~?���ǦMr��G�H9$�iy��t�������)�P�W� ��/���c k�΅�Z��-���.��1
!G./_栴��L�	�s	��ӽ��
_�aSW1��/
U<��]G�/��s��7��aQ@B��]2Z�z$\�f#&�~	��"�4n�8>����\�y�������U�����?z���_��u�����Y��B�Np����r�AG��z9H�mQ��,�c�8�x'J���a!�;��8�V�PG%�h(�ġ#a�(SK��E�_۠�%!6�����!�!��SZ����x��tP�ckI���|�Α����Z!4KK��,�7����=�sòv����_`8��^�H��C}2~�O�h{a��8����Q5��mTr[P��,� ءqv^.0XQ�m3̦\�
^��Z�=�2\ȕ��|Dǅz��<ؙפ��̗�1K�?���%����V;��!��<�!0����LI��C'ia�����K2Q�mSD�wL�}�}ks�M3��u�+d�F�V(o�hj�~0��.�,�#�{���)�CKT�P����vzvdw3.�$:FX͘y{s~�3B)����v0���!BF�<��?���s�u�����RE�42l�jR�saE�����𣏕�j��Y�L����O)>N�C��x����{\�n<����I
�b��I�ݳZ�y��K�Y�ҨW��Џ��XL�`U��7�������"���~�Y������l�
0c�j�6_�M��,��Fdw#/w_4�N��K�[��O��oo�h3M�n���gXĚDCL+Ճ�$�N��o���H�7%�B,1�]����d�Kq�	CA��+�~�g�l��g��^��O��w�qX�5��kW��"����~�і�Ar���Ȩ!p:��C���6'8ϕϪu�|2٧o�~~�P6�zz��ls[�b���I��i��]�|�Y@%�u�}rh�%ϩ���|t?c����Q{��k�Rb��]�
��fBB@Є,�4����!�H"�E �A �t���{z��6,�2��yxغ�{*�K������6B#�a�B�l`N>�u�M7&�^:����Y\`��YQ���q�,�\��0�_8��̫�-ɹX���3:��>�4]��CU!�JA5�K�+r�3o-8�q���&�;�GK�O�1lkiEz�ѳZҙ�,U�����q�}���O��?ê�<����{�{B�ax��e-n�]P��.=:�%�$GR(�I=߫?��2�<E���gF�ȒeYX],�7��/�}�B-��f�3`ώYS#�g�s3*!٪�L}O��ē�n�rxn�zv���pvj��h�t�;DEG����p��G&Y�t���D;�0H@ZP_���;����A֬@���o���w�N�x�9�h9�����V�~���>9T`:����/�9�TR^��g����c��e�!�0<7Y�8�?8���-�p�g1-^99���DT���_��U�;Á���6���K��_�%��cW��Ϙ�w�xՆp`N��(�ĉ8YgFC�9������Ѕ��XG4+
X��&%���s�,�pQ�(�������~��ǉ0\W�
g"Ùѐs<3g���}
g怂�X#�歙�:7VA$�Ό�D�m�ka"H)�_xp~?I;�?�?����G�-�"ȳ��)"�Ȼ�#�+s����FNM�x�X����_B q��\hG2%�.t�_$u����ޭWО%����,��4�:Mg�ڏ�(:Oh`�W̿�?��2tu,���j�KB�u���pY����>k�$Y�ǒ���ɕ|2�`�4�3h��h��#y*�hd�j�I?V
9���'��r�G>`#V����fƇ6�;��Դ��ix�����|��99\h��tp�xJDa�X�����%c��u}Q��,��6w�3RrW*�&�J!By�c>���y&A�֯�:���$��}�xn�nvv$�������{4�ϡ8Dº��gH��;(�Y���vu3oi}�-~h�e�����䆋���S7�4e�� �mT<��q�&�ȫ��?�XiL	���ӊ8M��z�:]��|a�=�y�F<���kH�8r;���ԧN�+�c�;�w�6�39�V�å@; ���T�PH��\K�
(�r8�w)ƿ򌣱`��b듩��Ʌ���C��;8�����*�/mg?V�+K5S��G3�׉�Zd��9]�C�y�bNU�V��œ5�4 g��)�/�y���m�"�-p�ѽSc�B�y�~�,8\b4~}e��f�r�>��Q�ܩJ<(-�l�:^�/��n9�p,(��(��*]��xSC�g?��+ET�T˩�VU�U[Vh�6����گ!k��e�ͣ��<�/9����W���W��Y��q�m���lw�|�u�˛P��u\�)U�E���Ý߳����|�?�����
[F��mz-��K����b,�	����5�e�m�����6�0�V��"o�p����P+ˀ�(����?����'�U�yzY�z?��c�O�w��1��|	�G��Xq$� �2�AG!�����BHa(0��$� J�īL6hAB��HM�DD	�4y�4��$T�ЦĐP��F���l��fTI�$4)��!!N����'[F��}`�Te{�

��Hj^��H�CBq��:E�UPL�Y=pUn���-u��4��p)��l���
��E��&����a���%���jٱ|�(+�@�-8B�c���z�#���C`$���%��V#g�#�ۮwL����%�W��ex�#3~2?qd�9�V�m��]�Ƅ+?vo��-��k�U�u3/��'!-�
���J{u��H�Ó$љ�K�N�7�t���OkI����`p�Ba�|��K`��!�OH]%Q��]X�cϣHo�F*83��Id�;�Αb��b�c{:�sQ Y��S4<�>1I����?�Fsw���ٰE>�I�?����4.x�fꪪ ��Y�)U���T9�|�!4}�cqrA�I��7���c������Ξ�"[1��J��&��e}ؓmG�[[Ռ�	�-�FR>.rL�c�|ko�=J�C��:0�����B1!��(䓚�dA���6m���ɐ����U����\�"إϦ�P$t>^ZVP�)iB\�](�� xہx%2��<�d�pX�[�����Lk�����8ȸ�;�ON 0�z���m9��uw$hG��A��I4TT��J�|\��J7S��@(d^��"
2�>[�!�:���Ë���D�ʀ��.�:~FKT��w�@é�%��J)!ߺ
JJz�Hn�	����������˸�*o�'�Hd�|�J%� v�$N�u14d;3+y� �?��ڡtg(,�ɪG��Z��Hr[!r┌H����I
H%7	D&��	�!�(B^������Xa��{w��/�
'��k����D��A#��}P"!�w���`�?����-'EZw�'�A����k��#����;429�ÍX|~��)�wV!%�Y�L�r<84�`�U�8����nz�J)$?/�+Z��v�'-x������FV� �t15�f�2^�N��,��I��|�}��A1��r%�͆ا|v��fm�u;���Y[���W��'yzTЮ��Qu��SDqr�].�x*j��Cﭺ�fKb8�l\�d��F�4�	Zr���4�7�lx`��������W�fE1��~Ȳ�=?��=����/�>q�%%$
F�F�����F�,�Cm��3Λ�!%�(�û��T=8?�r1TF���|et��׿�	F�!$��O���7�I�
!)� B/\GEi���2��%���\~�&1���v5cJ����17�	-;�n��0��nԘ�:󦡠pq+�_ȁ��m�X�k^�i0D�̺Ma�>����E �`��Iɉ�x8�m-/B���ń����|��IGz9$�(ܞ�Ί$?��iG~������r��I�K���.Y7��`�w���8�L+��l���!UEwB&��C�
%D4��'x#�1@��%�"�?��̧��{��9��-�8��F_���&~�5\�����3�Q�VQ��x��%��=�'��h���@� ��tԧ_�hۄ��&�=���%2�mB?��k5���_��%�����od�E�[�����B�=Tx�2M��!~��i⿙~�S�mq���Зu	<J���P����� х�"��Z�Ʉ�������l��h�K�a��:ҵG�QU�R�J�=�~V��[i���V���i�����w�N���Y'��#mj�eIB�SN��ې�s�_ϼ��.a z/ k��門�YV�)I��f�$���
���z�?�0���	�}���L���
-��p���CC�-���*$���I_'��Y�f��3���3�?�<�P���ԟ��V�2&}�z�l� ��p���tfq�����:~���~�#&�]�����6����&�_��%�[Ϊ� [@�-�|{ ��1"Q��E!�go;ۙw�*�_1kk�H��R��s��%��JI�RT���S[��IP�=ߋdEK)�C�!Uy��0�kUsʴE���Al:Bm�Mir:<��#�����ƚ���;Z5-�CE5$�ʱZ�xԋ��x�`�!�i	�K0l�=D�%�6d�B��n���X�������"��Z��17�� -.��r	@�Jl�>fBr	�����(��Jl���o_�5�ݷ�j������k4H3F��K_�jnǳ޼�c�0�A���=�>��Ӈ��Ĝ&�I`��l�zvR#<<��7֗�+&���4pFBo �N|��<���N�Y��<-�O ���a����b�+Ah�ad{���Z^w�]�� ���
�Z����-73	V$S�|�o��Bѐ¨�B!*�c0 ���*�c@�xݤCͤ����j�c��0��Sz���rA�R�T]؃\�7Q�h7G
 Z���n��"���׶�0��@��G��"�S��
qO$���[�9��+M͂g`���V8��bA�w�n�	�brF�AlIL�	�X1�i)��bnDg������blD���ILƆ���t�ƃA.�� �!�y�bfEH��L�ѱmg������!3 %���t���~ͅ�����#yS��3/z?����Ӵ��]�~�gn��;/�0� 4��:�dR�����;҈́����I#7�G�PE<���/'"�NJ9Ph�x;��D#�ށ��JJ hr�B+�䁤�;�ȱ�?;�w���>�����z��ڒ���ڂnŕ
e�ϯU�F�1��+�=���k��4��9�D>5@�'�J�XF��M��L�6%C
IPa���ռצթ� j��j���5B	V�i�Xj��S4'�d�B�W(U
�\��4��k[Q\�����̍R_��� �0R���6�R�ƢEU.eG_�����.��}Û~/�Ѹ�	�ܽ9t�Ϯ5.�F����+Mߋ��`��e�k~�<t�H-aӐ�6Jg�x�D�HY�]P��ڠ��k�ꕭk��x퐑\F�Z"I^\�P���`�Q��ŝd9!�F���!��#�xϡc���dP��i�vȠ��É:v�f&ʭNU+�>3R0�V�#����
��Y7lmsԿ$k�VA�ٮ8$�{��E9B��O�Ԟ�ېB6&zW��_�NN�^�mzވ��a,T���?�)�#�]B�'5�}u�"JS&ui+A�T���ϵˮ�+Ñ�q�$<C�u}�U&pA���<�f]|�R0NZ�N��]H�B	3~�Y8W�����dN�.2��9Ti�}}��r����
�u�b�UT�d���.٘�V���l/-봥�A�.��z�G��u�
I`|X�R!��ԟ����*Y�l;E�[��u]��KW������Q���ѩ��5}��
J�Ԍ�j�]*�e��{���G���_{�x�n�/�-���I�A���R���vCF�C�la����8B�+k���Ύ��oȏ��|4�����7Hf�j��v�R���8o���I�`�l}Dݖsc�ò~|��)�	���S[eSC��e����_/�v��շ�zæ�W�t]|�X4�!�g�=�A�XM�� V�[r��:)Y|	�M{����Ӕ樊T&��B9EĂ�Q]����������HUc^D�Q�[5#�-�gُZ��V����L�d��OGE��Z%��Khg�*4h��:�I�ds�"�{Z�/�sl�	�W���u�F��˹�#��+��AM\L���:L���� �6
���QV��BY��U=X��Ձ$�K�f�S���K��b���ʫ��s�|9!DvAt�
�#�����̆�Aj��>�\����O�c���7E&�s���8�x��>�&QmEIgN�l2�$��V���������ڡ��f��5:�<�+�8�}~�Z6Ⱦk;���]��"�mАK�ù
h'v96�'az�C��[��#���~�ky�
�I΃?hhg2�`�l�p�u>$�����a7���t]�[=��FV=���&,�L$�0��mLA/�I
_�d�>3�@{{h�򬿂��w�cè/m���_P~!��!�����K��p��뗿�� W�b�!v�j�[g�D641���&w�EI�@�ǘ2rEp�)p�ϐ�E7y4ѿ����Z����)w x��}��E�{��M����Tj��ג���(_����uZ�����2��}��ٸ��!�w���MD�[��'<+��x���	]���i��e6�m�>�^/NF�(�QYM�M�^��-����b�{XRA�	�E�6���%*;��Ao@U�(��y AwaB(�sG"/���U�������d/\<���l�&��IXo��8���[�#:���bi(�����	膤�MHH���s�����T37!i��|���B�bJ���A��^�YR�,�L�m���nܛ6!ᯧ`�d�b�1�H�O\0�!�.يC:�?�gEqI�>Cn��RK�wU��~h���� ���,0:q���`5����r��esp7L7A	�[k��Bk�6�cr�c�)�l,G%tt+d(�x��h,f�]�㝉js�0�������L�B����࿡�fфŨ~��;SU��i;v^�d�s���,bq;�4O�E�OJ����W���*��B�������d�o����2"�:��m�w����{��Q���5Z�u-���.�ڔ�X�og���S�K�dݥX��P8O,���|�G�]�x�"�O<~�3��S�b�*�#m�(B+KA�%�jŴW���K3 ��)
-�(s�k�?���ୠ�t/�߻�G#ȷ�9��Jv{�r;I	������]S%\kf��5[Q�U�D�H���~Է(��~1,�|�|�܇�rN������|�r�4�-符Pl����)��J�����Z�ϗ�8#;'<���{�v�d����~5M�M���+��+�ٵ���)\aIg��\�!#8�U���+��]Ͻ�a����4i}c}V�t�Ջw1�c(�C�I%J}茂_@��y���t�mR�tKҝ���}s؜iV�W�tJ%����Աx�(�M?��;�g�M\`��o���ț�'F.��,���,^��I�БwM�d؈0�Qt��h�S����95Wl�l�*�(mg��,��b8��y��G5�cg�q�����9�	Ѽ��$B���+�H���S��	@赎����,����&T�ZĂ���̃������eU:��&�ux.c��6�j/!n_�1���h��p ;���+�]#���Rka���u�C�y�F�ד̄�'<�N3z��Ȏ�kfi��-Ż�H���T�6���{&֣uz�L�̹����As��S��[���9@)!7X��255����Dq4��ztu�d)O�S�c�"����fQB�ɫo��u͜#G3=���ld�`Dl3R�^��Ņ�??�c�mgJ��y$�(��,U�x�$�|D�}��'C�c$	��w=�w儢�����<���t&\}���0���άm]��͑|D`IV���یd�,0�����ޫAW�#�D��{z��cWǰ�3�asJ�:]&]f��cY-�FY�޲�S]ə���evh:7���� �� ��:5�M���h�
@H��w��K����84�\*�� 65��,.�^������j
�Hw��;���-j��FNz�EZv��?p���"�ì��p�^@��Q�Ϻ�d%A�N�[��J� {�б	V����3������=�C��:�X��������T��Ue7�ȍ����i���<I��z�vLA9K΁��
c����p�^�0�Jyq�2� 0������C��^7��լ�P;/�xSH�Ȇ7�A��1Q�pY�p*]�/�Nt+�xZ�w���}X��m3΄�͋����؝�C�q���֖D̷���[�[�q�����������	��D$|Jc��s��ޯ��m���F��Flj(���4�s�*���|74"�h�aN�(C.��`f����&E�+$kޘ6~g�(f�[��N�o=�53YO�8]��ò#�ԛ���������f�c���d$���D��r�����'�{�ʧ楁��皥�2^�q�4��6X�iWOZ�K L"����\}�� 5�.��=Μ7�����v�;@��ީ���#��[�q`�矪[�<��L43{�+����+��IC�;�9����BA��z�{���&�F�|tdn���`��i�x^�(�����c��m"pX��AzY�u��<-2�*����k+��������#0�z�Kx��Gz�s��u��Iw�:��$8�b��h�u�Dyԗk�zg�T-�����^�4"F�o|���"�c����F>&����Tjv���&�P�}|�nF�i�*.&hUg��L�nG$t&���;�E�1j�%r�/$�Q�y��.`o�LK2,���E��³�WW>����?'�2�3v����պ����7A�!6X���m���#�)��.�C�Y!��mI���_�}��dr#�mNbJ����9��0�G�'���B_r|���p�(�lD2f�o! w!�B'q�)� �r�����elvݥv' �������B�Y�,�>oíV3;�4��1��9*����_e��L�)����m&D>��\�r�r��t�(�����Թy�l���?�*�a�N#k1}�گ�⚑a͝j�%�g{Y���k�ְ�L�3D��+�橤�\��6��k��aK��;����A3(�5� V�+#�轡�?�"�E�h�bw����3p�*�n��g O.@�D�a&��Sdl��*V�G�\��R�K��BD��M'����D=���܄&���R������/�J���T�
ܠ'�d8��7뱖��YB���{��x��s�v*؞F|F�EDN����% ����ь�pd���G��������>��\���!2}7I��u�H��`L�gcX^�A�j7�5��P�wL +ͷ��L����%���ei�b|�\U�3�xV��P��rX���Ƴ��4��D[z�-��V�����l��hb�[h_��;���v!eK�]_�\�/�必MUK穠�Q�'��l��z�0�<ё�T*Q6dH���Er~��Fq:F�ѯ�l�W'��χ2�u��,�`!��i�$��U�\�:L��Y�n^E,:���f=ۺE�U����B��
Z,Ȯ��G�ō͒��O�%e�S����
N���M�C�7�<��ߩ�"�?��)�䒞�1�;�N��9��f6G�.�ݽ���WE�C����OSm�R�A<�v�V�S;�5�'����[P�؟���.�kZ�3E�ۅ^������K$)�66�2����"Rs}�o����aI�4���ȼ�HT��	P�A�iAn
�����_x��][��fbl�jw��]�1��2:��������
d��)u�4��V�	!2*�UHx�h�B,~��w�8�Jr��M�趶\l�É�?{���C�6�dd���GTȂ%ʿ�D/�ˊ���~%H����}�7F|b0��@�^�c���K"���Uɗ/�.[��1C��Lp缅M�ֵb�p޿�n�����s[��~2����2Ĕ��D���L��;Ayީ�^(���Z.+�gG�o�;K�uO:�G���tݘ����p��y�V�̢�0���k��-�c��z�����T��+wfL�.��K�N���$ZS,���㒾�e�"f���t����U�2tc�Vx�?OR�T����tqPKl$4�⤺��Y�NL�K�)��
�F|�������%��]�˷)n�-�1����K�����C��9���{�ר^	�Ѷ�o!p���3�}sIl����u�393I��4FR0�iQ�+C��?�L����gv�߇l{g��|�R.%�7>^����&}Wz���6%Gο��9��������:N59���(Ez�h�=P�* E����,l�|�����^Xӵjw�&c�@���6w������Nۼ�^��r����_����
}����m��(��o�E��p�5�Z|S'����]�N���|~�:�&֝�������|[4*)��������'��nj�+�[+#����������l���I] ��.9����AU~vvFh6��?��G��L�>�::�Q�
Ru2�$๓��H��	q+��s
�1��E�^S2��Vɤjh�Fu���H}�g~ufV}��i�Y�)5�4Y�1�Xm��|�u�P54�x�k�;`��A(���	x�4�+9\��r��<��j��b �й���`�cɠWCH��dp�N]~��m.�E||؄�%|[�*O�}��}YOfA;�����yAP8����0b��X��ݴ����-}��ml��2Ӳ�.>�Z>�f����ͲLŹi��`z5a��8�I��9��+z�J�%_3'~·n=�h�#��=�K�*����;�~��v"V��#3�V�`{{�WQ��"�j�3U�!�,���_�+�%c�I,��#89��7�l�Yd¹Bzi)�C�@(��]6���h��l�Ejd�����|�4��<|��+��@R�qU|�.����'�'ħ��T�/|o�͈�"�+(�n�?���Ο߾��'x��Ȥoh\֗*����5[�^�g#���?t,�ҙhz��{$$�4St$&���`~�9�f�kl��s�H-�w9����0��0j�����_l��OJ�H�oF�)��;i�,L�xg�\����Fh���Yp�������OV���}M������[M3m�T�u�u��^2r@��:XEM%<�/�o�{�/
��E���D�s/�Fhi]�Q��mW� V06?�[Ɗ%.��*��U��r���fP�H0�6�q�vW$���993�� �UE�lI�J	D�f�&��2���^�jj��55JB�ċeG}�m���r.�j�t�dr��t���)8P蘏5!���k̴~1�f�ɴ󱎴�Ӭ8i���eL�D:��`�z����4���yJz�=�d x�,.���Я�MC9�J�1�Z�R��cb-��G�p�n����9��.T8[
��^����з�g���9�_�Dw&i�֢�
�d�1�]Oļ�����\%��+��� ����ƪ
ދ�0V`��5�H�j�-im{i��<e��{��q��쒛S����5z��ֽ���p�p����UO?&Xd��'��l�|��98��p��ƈ$"�X�l��$���N�텸[���Ji�ϫ��÷�@�K� $��"+b������d둇gk��I��20���8��p,A���Ĭr^FWB�>��?^lQ������4tJ�)y�T�氲����^�z�G�����(��}�M��l�cct8�\�af9z��l㊀R���<�B!�[�.x����]�[��[�s�^3s3ȷ�p|�N�����3�M4�v��ߩ1]�9,
�Ɂ�fv�/z��:Iʐ�3�,��LQ{�Z�ҦƽP�l�-j��)��=���{"=���'���� �d{���',۪H�4�]���f������#}C�ωI�T6�ٜ���N�[�ȡ�n�#f��L��������| ����X��3X4�s�z�a��3x�>O�yS���{��L�;-�]�^)��^d�5 '>$��	@Ѓ��^�\��*
Kqa$�$�s�|>ݾ6��E�O���@ ������������9H[b2 �дe ¶�W�z��S⿼1����W�+�Q�T<"��R�%�e���6��V�Gd�2ic5�0u�������nE�\kr�3�0�(��H�i YAڵ늬�V�L���!��S�ɑ���������V�ޏB�ݖ�׀c����s�	ũ�!��$��Ē���;X*�Hx�!؂^�Z�8~��>��P���`�%A��eA؆�I+�+�nVu����%a�G��bs��jz��:s��N���8e�� �l�Jd`��V��`��?���(�V�Y^�-��QK��f(�JmO�֩��Z�����Ԏ��e�I�d�6{�b���h��0���ctH�&�	�h�Jޢ�Zo�	;���]}�%����L*�owo�@��L�c1����L$"o��=�j�Ș��r��{���E��2C>D�5�ܿ��(�xMT?��Yw�t��t@=�ܒDX�h�.�eL�6���a��*�Ʉ��}���M|xB�ϼ�p:q, �I����8Y�9��a� y��o���U�pD3V9_oK�I�x����v�	`�7�ˀ� .�c��<�2~�g���cpџ8����Ƀ�z�G�����Sɢ�ŮP>��$AO�����&HA|z��F�,���9z�ů^�lˣق�����q��:�k/�&��$n-�~�>`�5����^p�V�T�-�:MI~�Ul�>�(Ll��:~y��o�������7���G���[B���3&�u$4
����&�Wo��'C�j�t�a���	)a�d&b�/i�
q���'�f�z �h��h����T1���FB� �S��0�A���ئ(�g���n�
}��"�:xF|T#@&l&-"��e{K���!�{?��ׇ&�@D��f��4�F����Y\��3~���
��۽X�ۼ��]����K�Y�Q@a}�r�e�3sQ�sY�1 wן2N'e�2h�Ld' ����1�a'/
a!>�Nh�AD���0��lޞ�A\��tB
��=���n�N��֤�M��}�Β%�/��1� �6�F�{���40h�>��.�ⱒm;�<�)�f豰���=�zV0qS,py);�2��vDG�_i\�n&�P�7��y:���m�c�1�[?r�u/� 0��+G⯖O��f���V��o�Ŧ�ߟ5U� � C�ק��������&��o�����BLe�u=�xӍ/�{.+����}_HM$�a:����ZQ,^r�K�Nc%3�H��^�c1	RҌ��P��u3+�V{��2��@�4�N�tyowa?��1��{y�
�Y��+�p�h���ѿ��A(�׵�e��t��*��b����3�����3ʤrq��PK�Ӂ3`�虸TxN������
,��}u|�<����_���l	��8لW��p�1~,T��s��C��[m>)�Z\���1���zh$���ӓCʐs D�ř���K���\i���MڊӕH���L�.�ē~Uy1�ԕ��9-�v>��b	��m�Ս'*�p�s
-u�Uڅ�K�5����x��<�Ba�x��\�d�W �^������@wcJc�j�:ֹ�a�"��<�!5G��,�/n�.�����-���5mc�)a��NLn�nݼ/�~ZE�M�V��-T��eX��|�nQz�}��S�\���x�E'ܛV�J��9\�s������/�¤W$�y[�Ì�k��F�ڑ>ߋwq7���7��;ӗm�/ø�}�p�;�J�(A|�qA��ƫ�py�Z,�$������`]�ĐȊ����)���J}��"��q�`��F��|�j���_���hJ�<�PLS�Շ�V$�=I�X#����#���ݡ�v�����;_E���5�S��}�b��d�����jOK��ۀ��itCwj����S�!�U��_�Q��8w�Z��)�$x+n�B��c�e_��ʿ��_�;��g�!�X���XJ���_@��O���J9��O��	��W���4�jph�-�L�i�����Y8Jށki�E@1�Q���31�����7ky̒��謏f��67�|Y�X//��W�GB�I�n�pҰ��y�+z��MJ
�����{���/"3��ޞ����-�M�h���5ꡝL��g)����TW8��Hv�ü��Wo���t���]4��~{���n}bL����q� �!�6�Ů,۽ձU�ͣN5,Zt��?xH���0�)�g��c����<� ���?�`�7K��(���M�����qM����b����Ԩ��ϻ��o�o����9c��0��QK� z�z��^uƲ�O�:��G[�v�m��L)�c�Y�
�)���4��u��K����a�C��t���oȜ�u���#�e�v�'��5�� ��]�0k(�<��v��#��"v�~�1b�#��MpD-���3���p\�U���'��@ܫC�u;:{��7y�a�gAs��0�r%�~Gˋ}�$��0|��&1�A���`�`�TE��Xz�ģ��s��p{ܑ��c�s�
�Yߞ�R,���Y��Jv��7&����o����ҵ�
9K�&�V���;����R�7��B�Mo���P��v���חN�~�'ۻ4����)��=~��HpS4����#��o]���#�x 4i��q��~��`�?��k���n�a|�T'�^66�p��E\�x*�j�0��h���B?<u�/��ג*��m8�d���(����v(Z�gjl���	x�I�a�H�����l�F�Ѡ>�i9��^dZY)i�}�$_Z۩��Xjjj)m�55��5Z����4��|���qȉra�my�'�fE��9~������^�"��C2Y���`���O��q�]�]2�X���>?r��.)�<ҝ���`dH���h~x܇_=��!�]���	��٧7z�	��Nu+���a�I�?Ӊދ�B7�e\�g�\�f!��	N̬��9�s����`�֍i!�}�v%1%��Bu�A����ʢ��f��1�i��#�S���!Ჱ�bZv�5;4�P<���:3L2űw�<����W�1i��~w_�#S8������*rX
s���<���ll1F���`�z'",	&��]H���S��;7�9+�!�B�N��F$ �rO�RؖUfA�]<N��8�U9���g�����v��n�ߛp'��D���}*2����ɇ���3*Y��M;O0���]o���6��u|0�pg�hj�I)�$30C��/�f���c�3L;�kn�i����(X�޺�d+����Θ��T�f6V�Iy���}�]W������_��2��ü1�LS4A�#m�7ig�X-N����Ў��t����|���1��؆�n]���� 0VAcl~�:H�u� 8������|�l��n>-���e4�q�;��`^��k�X�0-` !)��OVk#a�m�f߻-�۳Ś�L���0؝��'�I�\�O�*{���@��^>��}��?Pa�11�aoUx�Y'3����z��c�lYt���n9ɍ)e���g����g5s�1�¶@+l�I$2B��9j�m��*C�Ч�7���0c���m�@���4{�WE;2�:����t�����ž.�yG�0�F��4\K����<~��q}�z"�C7#�XbH>[g����Qmip�*}���H{�o
��ul�wF:n��MPX�\���*�Rk��\O���o���(tۯ�h)��W�Iؕ!x)7�̉������Dx�7/��������p�I��T����O.��אq� bl|AZp�N׾�?IB�Ba���R�@��'�
;�^�b'�����%���yA�SY"���i��s&�����aF��i><e�����Bv*�n���gx���ETr�K�{����o^��&T��Q�����w�;���h�j���W����q܇!��0�N�����s�m�ƽ�*�@}Al�g��Y�d����ń1amZb���Ex�(K p_�Õ%8��+��A�����l�ST������}�E`�e���u�TV�)H�T�[�=8�ί��v�N������x�� ~q�-ed2Y
�cy��!�W�<VXF��CF �	`$�7[�tQ-��5�КӢ�ف���M�%GS%̫�����>sa����!�&^�/��H|GjVo(Y$�#%ٽ��`��w׾��	Kԇ�_|˾k`���.����_��kE�H!$��x���l�L֑VVR�=b��U�T{���ē�����~���Va55G��c4q*GE��'̝�� �LClD��s¦U��2L�Gm���{����;#p,����J
J���w�s���Q��+�OP�$�.�|�>[U�����yΚVb}��2ڕC�C��#��A- <�nunZV|>�H
�EV�t���6�B��+L�c�����'�������<�礫{���)�a�	���O�����;e3��IeR�ص�Lh+��ߴH2|M��<�D��	H�lg���Kۍ�x�Ol]1����O��Ź0Lg¸_#��D�i�W+�������R;�k�U���L7�wI��/z�3���4���ryI��+H�?,���t��o�������m������̰ļ	,/����[�r����O��,k���> D����0�¾���pd�]�d߹��g��d&I�n����M].a�L�D�Hҿ��0��J����[�!��5�Ǽ�P�~1	;�݇��N���~ӳ�3k���Q�H�|tf[
�P�K5�ˁg'o�m�e�$�D��6>��'�7����oV�"�3.5T�V6��e���9�h���7�l�OL�k��HL%�2QҦ�&�&�.��h��S�*��w~�м���Խ���j�����)a�k5�P�Ҁ!
 UU��(~�͔���Y} :6P��P�*kQi11���%-G׶���������K?��GAGJ����Xl�`t{�_��(>ة$~$��
ڮOB�
 n�|��#�ÿ��ڎ[Ba��w\0:�k���]j�]���T����� :�:��pQ�Q��8M�I�$X&�t��bL���3m,XyH������p$<E�����f�{mӄ
M~�v��u\��5k.��_���f�
ПȳMU���ՄSV
�]�!X��갮]��-+4�*�X+���g�~�O҆��yeEG�9N�����[A��[�%ᔳ�;��11��C<o����Wح��? �K|�6r30$ֹ�gu,x�PV7D�����Z��TX�4p�܊	��(0�2lg�ٟ��@��A0n�e���foC�h>+�o����)Ȍ��t��aL�ؽ+?:�޵�Bd�@�۳^?��˄��z�/ \����� �u��$�}�x�nBomj��k#A�������qS�_��c�;͜N�����PC����ji�s�,{;�a>I��2JA�~��x���S4�h�!���%�c+�>�E7���1�~v�|�S�s���^v$��Qa.%6������M׺ր(!d=8",G&��O��J�� �ްe]'N�~M�y	������lp�����8z�v�d�,�+:����$���?� ���ː�X�ә%��y�|3�C��yW
ml�)-��7�)�e��1$�9%A�[�`�:!Nx+���}n��;��վ�����R����>����V�z�������k��G	��b^a���D��}D㏑��e��
3��,q(2I����{��p{���&�}�Fz�J���e֘�T�j(��
%Q��ۚ�w�xD2ъQu�3���)�7Nk~�%��Hs5}yB4Qc�QszI*!���g���PL�BB��+~��<v	�$��e4�_:؆�\*	�xe:��9��|E���7���Bљ�Ϻ��XQ�FG��q貯Z�G��6bmb�����.�I�I{m�N�&��[�Tx�t��|$�q�B��^�V$¢
�#��~�ؗI��*�-{*�=,�N��Z��F�!�wI�������`��� ���N>�������
@I`��"��l�H�85�FӴ�@���j������4����9�Eag��@�[9�8�A����p���nL��m�n��=�34��6{�2�B�%rA��Ljƣ�rK:M��oWi	�4�	vkbi����Y7Ƿ�US��t�'�7n�C�յ��aս)V�G���̎�7��� �PĜ~�kדڢ��½�0m��{���^N�����9�0�
~$�'�'N{���y�^`ĻGQpb���%�?��sQ,�QQ'��>Ȗ������n��
�sٗ��NBM�j"ت)06d�J��!N�h�,gE2!g��!�38�W��["�mɏ��>�YmV��K�Q�ܒv�@n�sdN���bn�T~��e�۟<�<��d�Ax}��tծ|�� 3��W�+�2�4��/+�ծW\� ~�>]�K?+k�͑8���}`�]͞ӌ����||���\�,��55��Uɭ���g�Y׮�T��/��<S[�Cj�k<�6����%u����Mk�z���Fc�f��~�X����u ���5�w7�O�:�Q� ��ы
�bD�b����r��]R-�� 0l`'�Þ+��Pj9�R!�H��ܩ���͸���T�%/����%��/���<=���Y�ƛ�8W��t� jy���N�k-5� �u(]�è�-�*��rԓ�K��k���%3�Ҡ+��v�����\�k,�`F��O����S���W.!�+3����V�5����=_|=�j5܋�|�FE��`�0���!9V�Y@� �G-$����n��VI�_�5^�Q����M��V���λP�b@�ɮA�����D��G.��f8�X�uT��!`��r��|�n
����G<:/p�t�qD�Z���;��|��跪:�>Y�{V�sT��aq��%8V-Zur�Dc	$1u�j�ĭ>q��+�sMc�QK1�)�x�H�*HL\�L�pE��;��z�#J��N��m�@1Xc��8�� �gڠvP��&�kZ�KڠXˈ�T�BZ]E]Z�q+N�%}PE�P>O%�ʘac��D�[�lƔO�JR(��,��6�7�:�O��҂Hm���6;��Vjk�#�,l�c�:Ph����]c��N�� �
���]&���o�(E�P}5P�4��5����o�`���{�k��e��U��Y+)����j%̂����&��ނ�W5Q���ڊ��i�ù��
�K���)�ӽ�9u2���u-G�������o� ���|�	(���a:�M)n��n#����/r�灗6F�E��*;�	wVj��n�cgN�~�i������>ai�nf�M$�euuu��Ļ���~������d���4��Er�#���f@��W���>��4�N��$��c"�e��'Р�&,{�|���G=!��p��Q����RV�Y�����8P�:���U�[ۯ��5c��ErL2�]�l$8{%�Є'~�eU�2�#0�X�0yv���s�-v
qL������BE/#�Xw_V�߻�R�]�����C��d�������a�`3�W�\�ana`#Um#�v팽ߺ��~��t6�*ՊU�o�#~�t��[���4�����Ğ�ܺ1�4B���S,D�=W$�duutZ�Ĭ�b�W1�J��W�R#���s֮"}oj��I��A?s8��,���n`�7V�G�W҈%3�-��=J�����B2BA�2x�-<�I�P.y�5��?E���z��ę�Ԓ��w�i��%b���Wt+���S���i������$Tu�'�&��m["�a]Q'=���1J��h� ��%�㄃��ˬ������q+5د�~��p��gA�,c���A�*x������~�(P\��H��R���7'�XJ�A{��h��9r\�zB�҃D�ݼ���Q��R��ɷQK.m<�*�q�!V�܃Y�v(,~��F��\��U5��>I��,p��	�c|9��@+hJ�R�ϻ@�a��5ⅇ�~�Cm��H�����㬋>�f�rMT�s��;v��i��q|��Ei={g�mÜsu�C�vʶ����fK���|0��I��p�jK*�F`7��߁�U�L~ߴԔJ��}�QaKf��
���ӂ���G!Fi��9���<����]����si>�K�_XT���Cʢ"=D%!N�C��=z�B�E��lxs���!�����֡u�p� ��rת���À.״�b�i��ڤSii�\���$�h�]�Y�_�S�X��ά��M�;y�mE����N���G�1��7�v����mGo�C�{ɸO�W�SS��q�޵[���3��y��N���A�x|N�ycs90�����#�b� hH���U(]g�����>��H�~���[�$�w��oߕ���K��T�!�1��kN�A�GԿ�2��)�b�N��P�-��-��G�[[<���pC�����W�3,=��QI�3��qc7�e����Ǫ�����4y�����!��oђ�AlWAđm�e)sRp���j.Hc��w�>�L�9�z�l������?��$���8����t\�n
\F[0�L��
���;QCV��EG#�	T~^3�$�DP6a�;��i�5廛'��砚9~��Q����lė�b
����Ϋ�x�ܼ��/9����T5���@qJڮ� .�t!)K������ <Ot���5��p��&�k����
�MK9ߩ���3�WyY���E�	e�-,�̖�o�������/Bm�j"<�q�0s3Q�����j�RFO� �m�����)��޸2��
�&;U�������Qo����Y��BS� b&$��E�X��L����w�=5�o$�"^�|b��B��5��VaT�%h�I�s���W�-T�{ �n{��E����4���`��"C[㨄f�A�j$y��u����a��sP��3���w�rz{��+�Y|�X�kQo��h-m��eP4�+�W�@נ��K�p�9����5��@����H�����JV�	�U�!M�s�i�h9��q�w���S)�uc�G9�) U����A�"��%�R�%����Nj��D+=-����$6R����)�(�$�� D)'��T�X�ܵ_���Ǘ.e����9v�YD�b���B
�Ry�pL6y��D���[���Eeŀ��.R�Tφ��D)�H �-��K��ZΟ��b*�h���>4)���� f�W�P� ����]	��.����9�Ua�M��$� �!�g �)8ŉ3�^Ft���M���v=�U߇X�`���x�(?e�:�YV�z �c��u�,��NT.���i� �^UW�r�|�kO*�nYrbd�{����a�]���M����جo���ڷ��}�E@�ēl�gjg���r���i@mVb�z�At�:\0���MBq�jw6[ld��Qe���ZQP�%`j*1�B̅�ŦE},��Y�Gb���b�׃��2��Lcj�8u��v�0�s:4�``��A���0)�M��ͽ6'�IpL��\�[|��:olv���[�����e�
1�#!�q�����W\R&t'�3����Q$��$���	�����M$�S����Gӊ! �'@Hґ��DБ�#!���Q�,7�2Z$mf����`��p���,�c\)8��L�NWҿ� ��9�q����B��g��Q��3�}tG��-��6�a���AZb����0�?3�,\�^���������p�57��ͯuG�N��V�E2�����gI���ϴm6@�:�y��y�"�5����nYZ}���Z4Q�I4(�4Ƭ21gL�FW�A� A�Cߞ��7��Xȸ3�&��a�b��`�m`��a��,�Y���ҽ��JA���-@i�KBi�U�L��`5,�+I!�HY=#����7�	�ݍ����(�g������{��y쐰�,uɭ�=�0�#�_�`D�A�"� W$�Qv���M�d1S���C5�sN�4!gD��Р*�أ�X�0�\H�%HU����@��g_�NqܩFv�_E޵����� ] "W����Q	�NI��i�ť�k�c���5'�7M{^�ޫ�X��X���A����G8�D���mX�+9E$��A�\Bk`� �e���wI�ϲ���C��᧖����\�x�ץB�D����uK���:���7��T%��ң��A�������5�?��$/�$��/�������d&V.\M��P�\8��[�N�d��ԝ:r	�� �����0�t|N�ㅯX��ir\IOѯof���@*�v�������q�v���~�����|B��ۨ)�ߔ����{�<��*M�n��x$s����	&�[���0�l���oؑ�؛=B�_y����l�C4|�C�^�L�e�&%1��E���lO\WzhBG�ˮ�5W���:�M�����cn[x��R����{�c$��d�����m;��=R���=���:O�ؗ)d���j��X1㫵+��_��U���X0WD^6�aYaa�h�*�ڳY{!�V_�N����j^�H3k�m~�c8������,\�O��T�Fex��[T���I����%�b��dBLs�ߦs�F^���	zԮV,�41��+m_J)��[s�N��g�O�NLH_�xJ�@&$J�M톚$	�K��y<8��g�P%�;x�<�6��+T1�+�X
}w)"�ȫ�c�2|��s��t!�tNď�b���C��k}I�Q�r�Ȳ�z���f����z�W�G�8�!+w�����F6Q���lw.mB�.�M:�ѩ����}�vi,`��գfΐ���̖����LZE�!���S�]%K����I�~aOEtw����B7��O�\��Ӂ���qw"��,�Ff�Y���ҫ��T��Ȑ�r(ǂ|t���fY�h\�����6�?����C�;�a4өA�7��D{�w	|��<_�
�I輫ud�&�[���h�n{��J�enml<я�ơ1���B�$��0�A$��0
�Ix%�0_��0J�`�+Q$$PK���Ȣ#���hK��=|�|�V�J\���y	+���F�׋(f�{-�ۗ�I IP�|�=�5�ԍ�E}��X=+����hEƲ���A��服�������E�<�o��T��|��<
�ל�z�a�ȫX^F�e.�b��}5v���q�-g��`"��5�!�!�O�@V�{B�/7���
z���=��j��/��8�p=�R(Y��c��F�����`$�+*F��-y2,�u�3a�Z����xE���%&D��r6�e�RjZ.)߶.?���t�E�wpL=�~�����n3�Đ[�FW�@��G��+������r�1T�Ј����y�����)A�]�\�e/��n�L)�<���*�^ZA�t:�2�a��U)��pK�	���.$<&����Wt����*e�k�b*}�\��@����<Z>����һQ�����D��jԧg>�P\�+R���w���Hd�+`���>^��+g
d��5}�u����Iq-����a`N۪��D~�^��e�ɑ}7�J�3��t�/f��g���I��~|�b�qS�:?��q_G�������sT8��\�ūl����o�~T�vm�^z�g�g�{q\H�7G���Ӳ�g�v�a�{3��K��t2(�{��oE�N�O�ۗzo�y������::(a��A6��s����ǅ����9�c�&���'��I�oH"�l�mnyY��rt�}pP�F�=n�!+�� �q��;�����_�S�a���j���t(�5)��������s��EE�:<	T.�:���H�*�)�J�(�a��\Vz��~�Gt���|��n��bNc�J]��W��Xo�~�7��<��O����O2��"�������g:�s�����D�0d{��KP�,�rwV��^�����*a��%)%�;��w��5س @Y�9�|&��;�<��F�?Q��1�\-*��+�:�FV?���8�Nq�B4ט@~͠��d��bx�Y�P3��g��.�|E�0��>[A�f��ԒD|�+6�Af��;�ߴ2_GA�6BI����j��V<���b�<���	R(Z�A�;�DU8����J&��s��@OC���q�
5U+�Y�Cr���\�)|�"P*p��B��vOXb�t6�������|T��&���Sv��Bj��G]!E�h*��@�AI��
A�a� ���
��#�V�wp&V)d�����݆����u��2Z؉pL���A�����Z�MP��=$�#���	���b�,��
3�
� ���S�̪fS��ofs_��X�	
D\z3S�T�U�����S ��J������I��	<�� LI���4I�j��Q�Nuߋ�7-E�M�5N�{���{UY�s�yw�^uv�Q�l���<�Y~߄>a�.�g5/5��O�̼a~_-B�ܿL�tm��E���!*<��m�BRPqx潾�����9\{�ethpԀ{+5����W'���)c�4�[_#?��JUc����Y�c����n�-^���]���4$ɟZ���vb%����F"1�{�p��/�s�g���6.i����G�Mv�n�@S��'!�4o �V{�&��q����|���\�*��(|T�>֋j�YG
�,�IpJh\�3߇�P��ÅQ%8	1E{�绵�i9cd\N��e�è
����:���#��1�,��>��K�mn��"�ﻧ��?"i������Ne�6�||�I0Z���Xŝ���c�v������T$��7�_�J<Q�����dQb�۠:%���
��%��ي4A�k[���.�3�g1=��$[��=��уદ��QBQC## ��D��'10l�{>Qm�;�� �Κy����b��i�B��R
./:f�Fi�4�e�L�AC@$�@	;����?��@v��ЄihB՛h�p�]}�!~��ýס�8�Y��=c��Yl_�����^_S�����/K���3��V��mB���c�=�2�ڄZYp����f�"/<��U��"k �Sg�Vm�H����"p�i	j�t�3�73��+f�
���2:�k8��}�f���	=p+��I歶u�T�	W+��ew�n�0)0_yH�͛���ů��;&xWsF*���<Sܰ�Ɂ��ff��*���]�xl�yhTd:��pj�[,���	�?΀Rʃ�x"'2��d� k�[Eu������ І�
M-[�K\�ư<����{<X=g�Sp�����,�x���]Rˤh��0�yD��{>�=f-�@[qo�S��m6[�"�p��XV�����a休�l�pNpL@��X���8K 6 �l/��+;z+9Q9�|�rsp���S�N4T҉�	�
8����JJ�%���f��]����޸��D��3�3i����{���/g߭w����>2>O��.�'ӜB!�+�9`Sb���Ҝ�C:oB,��|	n*���%��ς��Df�)���$X��Le�U��,�@&�Z�&�Z=�bY*T< KqW߼Mb!�Fկ��]��^�>��EY:��ˆ`z�ͩ�������L�[�T�)|9&!���ڥ.��:��8<eb�"k��?Mӥ��-��C��6Mm��.k�?M�j8�2{�"uNI�3t�=>�C���<$��)G�N?�)�h��@�IZ��k^1Mɩ���OOPd��uJv����0�}��D$�>5%$D �;����=�7��^��K+��>�����itDQ{)^Ұ2������v7�}QNwT�Q�?;@xrJ�DQ-�D�4O�&���y�_R�r����G����0��GKS�䴂���?ŵ���R�t����gQ���H�A&����}���EG��'X��m�m��@f	-��.g������}x��]�7�V��M��>Tɽ�a�㼶
�U,�N�!���\�o�QFk��>b�����P�d��9���Hɤ��fđ���ǥƤFƐ�2u�(c	�#�&����֛���=*0	��^���suBu�&�G�C��^�r	q�����?:����(U��hl�`D��U!������:8�_��q[Wߐ�6Z)�N�W,�M[�q�����͛F7}�Gm���9u�M��%d�r�#�T�f�)ZI�/J�?�I'�f*چL��;x���E3"�[���}{��yɟ��&�0�s���^�d����R'��g#�\DU�����Z�15�� ���c��Ug�o�8T϶�k9�7�&����%�U@'}�?�F�Y�ʠYLw_��������My�SW��d��X�9Gx)�t.���B�\vE�p������>0������Z�#�����d7�"|g#&"xMuZ�H�����1��N�Y�\�)�%��P���d������5 �UP;�
7kr|��%Wl�`J��C�	xQV&�����͑������|vP|�L�p6ɫm�i���ȑ��a�b���<}�	P�@��bt���^ �x�!�5��EՈ��X�8M�
�
yqJ/2[�hdb@�4,���'PO��\���}�v$��hj�2�r �\=����0)��n��$|��l�=
"C�b�l��K����e�#[���L}���u0�8R�)!Nx6[���h�M����A��/���� ���D!�H�x�b�aP���@�@�u�-�U��4%h��`�=��vl�
��(��+�,� ���Mӭ)�nb��XN�?x�0X��(M�(�>��O{�� ��A����RI�'@]ԥл�ς-���������i�F�*M�8��#�Ἰ!���DW����#S�V<���R�>GDm��)�<i��?h`��� ���d��:���xңʢlN}�I�����>���"�i�Z>�j����3n�og�%b�2�$��r��3�Ek��]a?���_)����7H�,����́��w��<���w��q���/�DG'M�{���'���m�4r@�1���܁~q 
G%�tH��[�+||����]���U�������G��b�7���s#�v��y|;�o����޴Q����&�!HGZsM�H��8M!U�[���
B֛9��k3���vZ���y������ffF�$^LFd'��6�E9sR��6��s_Z��0�a�!�ȵ��V�m��y����e ��2��.r��i��]�����k!��1>;�a���f֭��Ǿ,�5��D��׉���[FUT�"��ظMh.�ڎ[٨��NC�H�q�_�哊1+$۩a�_ft�Q#��{�6�A�Cf�p;XX�2��p'����R���V�G�F5{P͌+ZG�Ց`2��{@%���{���꤮9��a�Ce>$n@�j7��0���paА5��X�J{�i��H�<&	#k��:��ԓ%��J��<;{�-�HR��&Ύ<K���{%Q~:����fO�l��bY�ia�O�>,��J�[c�l�
ăO*%�|�����h�K5�^\���
��jxV ��1b�v�{C�X��L!S�R��)&�A6�n��
R%x���RӈB�}t�����gkp��P�PS���us{r��qߙ���)�E\�JJ�b�K�ˈ�Tۉi�F��:�DZ	���@���Vx���6���l��}Id1������1�i�8�l^oVg���k�y�[T�Rؤ��N���Ήd�h���Yqm�^� ���G�[@�#:Ӧ�@���*f�l�XK��ÅB�d����	|��i~�c"�	�Bo�$��:@}	_��aoPw�
n��+�CSmdG
��u��P���{'��dKS_G|s��y1"2�1���e�tȸhR�Ә��$,K� ��� �ދ�_���vS."�=}$�D5VC���W.!��D��jg�2�p�29���%c}�j0���s�=;�~�1� j�-�·����a��I��^�hmVtg'���.g���a��,n{�³��E��s�͎|aX;�N�)�.^A�K�
8XVvk���~�f��z���0{o���
�c���6�'�В��]�D�f��j%`{��Fw�9G}m^��h��Ĩ�^�(/��٠�'�}��թ����6.�l���P���d��5ϕG�Q�6��sh���9�a��Tɹ64��9�af���/�.2Hn��k�Cl��ݟ�[�3�6�Қ_D��G��c��y}&}���'lZeyb�-��v�$���ZQ��U��M�YZ�w�Q��G�����d�k"+�)c��L��ō�)��2K��~{��k��<z"��I�0�kbd�?%���}p��� KSJuH0��
��ĂA�s�h���r=s_+'�E6l�q���g��q��wE}�F����k;�:���N��ׂ͂��d���,��s��Sy$d��U2C�Ԕx��JPڨ��S�6��f��9֎�u�^Y��.�8np{�3J���I(�i�����O%�5
���
�
ld�J��!�����ԑtK��ٯE��0OG�M�JYO9�����{/	V,*W���H{������#؃����1	���=�~�<0�i��Ɉ�oj=��&�m��Pg}X��� �9���:]sL��wm+��`)�2e&�	�6�d=�ƣ9���k�q�2͇�㶩��8ذ��D�+R^�3A��/RX�{���=�OD�B%~�l&��T��ȍYU����JR�  �M\ATK@�+ۗ������.6�O�nf[q>�>֙V�6UՆ8�D	������R!4�����d�T��v݃�r�Z�ǽ�u���=����]��А���Y��;��$P��m���
%ߺ�.��lu�'9�q�h�Ӥ���-�d��I��8�P���A���ZR�ms��m���+Lv���_�YwB�+����#	{��=+9��2��B�]d;Vy6%Yx�����~QB��!�{�P�q�ì�c�&��>��|=��q	�]�Lhz���`���G���5"�K���e=�lɹ��Z^
e��|���RM�e+��u�&
�P��ߗn�8r�6��3M�Ak�jR��#Vow2GӚ^�ܚA����߱�p��:���5���=��{փ���m.��U�J�{�f�~pp�;;x��F��
?�<l��	1��l0��0lj�E��K�����G ��T���i���8�4������/Ov�}s?����1�t9=8TN�%���\�K���m+܎��ᱴ�����F��!nUn�V�r�W:�!k�u��֋+���v<��]�?QP��D
|�]^E�@��=�y��x6�Փ]�Ȕc���^?�GlC���!�B�P��B����5!�7��'�ӟH��#4���i��;���'�$�ƌ�q�t
K�_S"���4O��p�ln�q�ʆ"��y�$��s�:^D���@@�*=O�f�wW�������g�_�K��D`�����Ӛ�D׼Ȉ�	6'�	�%�-t��|\{�/x߿��yoݯN��K}�;Mt�r:ʊe��*��G���������a?a:��l�ڽ�H��F�a�����Ly�t�N��&ōza"����r7������������:t"�@�d�	�D�3P�����X���!�ޔ��2ο[{��7���5Ax~o����q�K�u]��_��|k�������k�Ʉ��a����w4���ET���r�%�	E��eU���m�&ޡ�3Fd�������O���q�6��'�ig�	��7��C�*�;�o�}�u���O�e2p�빯p
n���Gp�
��v��+���$���r�!*�@`�,�Y�H��ER�S9ӛ���xތ������v�.܆\�B�>4�)%�G�6�YV�=�=��|G���+��;׳~!eTH�Q:��r۫��F6?K�Jz�2�),���f.i��V�Tە$�����
��L�S2��+�G.Pc���sH;�zY���R�9>�oq���Q��̠>gzL��L;2Φ�����)�+�kJW��U��3B���uE�c{HN`8ϴ�~=0L�}z��3��z���U�=Եჼ����&1��{T5�F�n�8/�_WP���R�I�D0	e^��R��и_�m�c�؁ F�uD#�/�zl�Tg����>\|�<Xy釂���[��5����
�~v�l!/$}(��?�G}ԠݣZ
9|ɑ<���0</9��*��pyw*�}�xb�T�dF���5�52�c�d��N+l-|ǛV�~�Jt&���*e�;��*A����婛]V����{m��VR_�Y����~���eaK;�Y�ѿ~��}����^I]<%t�Q�>�f���w�Gڙ�Z�����y"�u!K�a"����=�M���ޏ��yX�7�xo�σGq�_�񞓉5�#��O�m��6���U�Ӥ5��=�maa�j�MJ��x�����s�qM�`�u��ˎ3�����JY�v�|���Y~2�%�~�+O�{L����TD��J��$J�f0��2����(KB�As��ѵ5=u���a2S0��󍸽��蜬����x��W���6ѻ�ٍ��=}�����<�A=*/8U6]������:���S���7��F4y�H�7��7�t�C��dnKre'������uҦ���+B��Y�Q��k-[=>������z��_
x����ģY�@�Ҧ��|J��1q��?9�^�lP����Y�K�x����!�d�fp��3�E̡��Yф����ع�2Sa���<7v~�ٻ%�Ŋ��!TWP�u\l��������$�ؖ3�fJ�k���	��6��,�B�剞���j��8e�xW�N�$�^�s|%��^�K
���E[-��;��F�gSUUJ2"ʼZ�����Ŀ슌L�dB4e/�H�
a�_�W�ҟF9CL�}s��Q��n�x�KKʎ�;S�u*D<�E���س[$13<2�'�QF� �L�H� �M���Ї�Bo $
���a��WP6j�|@��y����&'#�DE֪�pS�"�P5`*_�Om���:
��r%�&�q�Pb��h���~�����n��f�J�J��T�.<��%.La�&�d�[�Yu�ø�nD�����ޗEr;2�TyTrv����$���Tj~# Bw�­C)��DǌP�>|�o]^rM
}�]�m���>|��_=g~2�C𢂃�N��"�k9xPW4��y٠H-��w;z~���v��Ƙ�W�Y�NV]����'�S��A���N����I�북�]nG��qI-���6bY.޷n����[}$M�;ttR>q�I�B8R��n˘���!�ʄ�;��	즦X��MzL�EI]R�HݑD� D���x��M+��V�1~RK�PQ7�O*���(��	����7#��Xp!�~��+��Y{�Re8?P��K~�;E���s4{�BY_�\nn�\��*�8広u��;��Y����#u~~��)6b�Hչr���+�&<�Oz%ʄ�E�l����m�p��r�]W	�>��F�m���aJ�5���zz�`;�V�*�k�#P6��z�2.��[���U���Y>[�����چ���(�*�o� ی�����ϧ��#츎����)VA=9�(��}*D>#��`	~���>�I~,C{�R����rǂ`�6�cTN/n��F*~͒BH�T�� V�@!�d��U\7޶�� 'E5>�'��}��mV%��?2b�����
2�F)�4��7��Gp�I���W� BXxy����|��,���9�ny�R�"���<���jrr�Y����1�}H�fF��U�ۣ�<1	���M���c6_���`���@� �*��"pCG�us�O�z�x#�V��m�
��j	<����tw[a���81ts�9���fG-��7����Џ|���tBpZ��29i��/���']�s�0�:�"I��>�z�À���C,d�6#l|�pg�J^�U��q/�\D�
����XGv���9v�VM	5�D
��Ik�-}
��Ph2��Ͼ:kM(2�?6����+���7��:�_L�>@�����P�)������nBk��xU[j|�\���'5�]ou�3|}���P�Y��z�([�c�!�0���׿�F���%L�~z��3	7k8r:�ǟ�ɕ �}�|����'����(`.3������������d����l�KY�~F���
�o�^���.��u,H������̀0+ߨR�#��<i��43��) ��a}5��ı��T���O���W�9VE9
�1���@���<'k�0p<���֗�=�����ܾB}U�<*�	<�̷a��nk�	�t9����: q!�G��X70%����G��j��CL��D����4ÈI�QtI�Ȍ!�h����荾���|�KN���Ͽ��)����u)�h_��{:軘������EÈ���\�-�جL������*[wU�I��Km,�~��۹��E���E��
}��-~UC`��0���y�)��5� ��!�v�D@�@��*@���A
-��\Q�`%`<Ld]y��	��;�����Y�)��NQ��N�j���QD
�$���N-��TQ�D�#W�v�0@ �y;�u�#T��������"��K�\�t�
��[fE^�
�M<�p���\%G�@��'Wd|�Sz(�$�Qs4PoX�xd_5g]>A=�'xc���햠_��*���S��)����lc�`\�#v��1.�$(�hM�ۻ��ؤ)ՠ�E���xSMC��$(K�ۘ�+2tUC4���y2�2����h���HT5&9�g-&`���"����MI��`%s��P	e[B[�B6b������]s�@��O@��I��E(<
h%W�U�3b`*]~.��89R�R�ڋ�m;Vq��t�.�p� 4�O�i��Y�)���i �@�U�z��(��������uf	jf	mf	q����0H�
���؂��m�#g����������#������� J��]
A����^�T>^��͎_o�B�\�r���ܙ�n	7|�e��G�[��z��C�}�Ze�&ct��7��g�%"��`����.c����7��o�46��G�3~Sv�ߝJ*C~=����Na�[�M�/W�;y3�L]���wl{:'�	L�/�;M�����=��o0S�6XT�@��1��Lqc$˃��A�(¢t+�'EM�Y�$WRQ���2��^]�:��^�<o������*d�[�Pq�p�n�u/2�~-9��^�3��v"���"U�gAj�Uz��N�~�.���ȥ� Z�
�h%<�~�MFDW���*���b5�N�EG�H���m�:}��Y����>�0���7Ǣ�¼�3�@܃njkeV���na�l0�Z ��
t�U�5���A�S�#��I�<]|�R�4��pD��bIW��E;ɢ���%�A�p�ɤ�6kĊ��C��W��$*y�-wSX���O��ŗᕢP�:5�H�_i��I1f�_ Hy��.
���v��@����alq�R ���B��J��p��Jx�UUDQ���/��S8�
�C�����H�R+�aw|F"�cx� �g��!��1��#3�F>�ll
�	_Phn�TDS`H����ܟ���h�A����	�S�H�@͉Z%��}�T�N�eڹ!B\�-aqg"�"Hdߒ��r64�d��,O���x��0.' ��2=h�3ʘ����u8�$�Y���O�A�ݻ겓1��fO��.P�I�7��c��C��4.����'1^�r�|&XlY3$z��Z�9v�yt5������                                                                                                                                                                                                     C;2�  3G��股%i72�b��Q�*&)I=5���I-���*]�t��J8�h�+A��&)G)�&5Mؕ�C�x�����ǝ��9qGTu̯���-�sfnb9�o�`-wAjBo�F�n��XnV�8�����K�be��6�e�fn�������w��~��gn�u��_��aXj�@�$����;�d�d�� �"&<��H����@�	~���! ��@���]v�.?�-sD�v��
|��C@����iŠ��@��%]-�{��_�c���i��G��S ����B�*�ne&��b(1�NJx�82����\y��/�M�i�6�;Cں�:��f�C��
G��i-P���N5BF�vy�N�\�d��c�0�H�H����Q�q�x˄�¼왒Au�o�Ŵ)�TK8i�U���(=�ڍ`����Q4�3F�xP~M�\�.��I�p�N%}�-�rE�.�_����6igI�y�±̓�]��+� ���]���]y21qD_�FV�4���Ѳ/��0�L�R hm{q��;��~[�y���+����1`�G���GAڃ����ڷ4�`�Ҳ�"�J��G��C��~���"��6�m���L�@鉜�L�v����5�+�*zO�/9�!�}9 ���k�K"ZGt�ͥ�O��>�	���鵂�8�ӼI�Nw�;��H)+�J-Q���چ_+�v�+yO$Q-,Ug��rt��z0��t�T-�2�������0�syR�D�x�@�>�a�@�U���V��B�}d?,��Wv ��헧̺<��Bu��\�+���o��ۓW�|#K���iq�8�i.X�;r��Q��H������r�?�����8��æM�w�$_�T����_vCY��^NX�����_hۜl(���]�ķ��a���Z�]�1���#zʒ���O61߭F_;���ꗲZc类���#�@���m����g�T�`��Y��䮇��|�N�y���kc{��j����e�EO��w���y��S��B��A���IM�B`'뇣{RE_�����cn��w�C�1t7֤h���z*o�F���/�7��?�C���v�[���:��<�F�zv�p�����װ�r��5�j�9�V�a��w!�mXv�D��A���-t>�M$ͻ�W�F���%�v��t��.��#Ւ@��4�cj�Ip�e-7wfw���GǞ�&<�E�#f�0F��챰d���J���A���WPT�B��������]��i���嘑���a%z��Kf#���DqC-v���)�k��2�Th�>A���N3	W ��#�Q���G�9w�����H���`�z@uW�$�)̮�_?�_�mj|p%����^V-_��U$e<�؆��ڐ��傩Ojw��D�b���S3!���S$��?�n�i>����o��7cn(m�s4#��|?;���^��t��L�fd]C`����}�$Β�A}���C녌z�#����X�){��.�[Op��G}���ҙv�#�`�D�[5>t���sc��A�	�X�5�c���@��2ՙ�����Nl�`/OD`#��HI��������EW��� O����Y�� ��f�?����Zc��9�$S��>�:V���Kϐ��d�15�V��4�܋8�W8����̲7ۛ���8��������5��}S�[���*5���gX��%sRu���ĨA/�������̣��|��%:_�s2�b��EL3h��G&��������>t��?An |u<�d%1ީ5�L̟w�TO����uFB*��Ty��^NN���8ɵM��u�[1��4d^��Q&�;��o{��l����K�(�,���;�$<n̋�!�z��v��>|��hR/`��j
�j��@��傲�-a`<�\%C�$�=�뼽{Xi���Y�1kb�V����΋�%�D�65
Q�M�(����4��e�;#�k͍Ŭ����c��Ž��p��S�c�2 �%�Z�H�R����u���U07�(D��S[a�	�]wL��S�%���w�/���4�����3�<U���+t��g��3=�Ｃ�?3���,ΐ��eDm�����z�f�}!Uޖ����M6rGbg��mĮ;�켭����s9��iީ�cV�d.V���/���I��צS�I�tJ���*PժٖZj4�O��h�������kXo�Х�F}�)'��GΞR�����NL�� ˲`e���2�����xg_i�����|�#�寥�[����~%�Ͼb���DNWF��_w�`�+���5�W�{�!�juA�*c��wv�>�:>25��6�j����Cɤ�����&Ft�	ȑ=옳�� �n)�d�����"�r&(��{"s�M���p�9����:L�Hz�/�B�ѝ�����1���`�;�"P(�k Ț���xP_��׿KrV�]��7,�d+n����2�!�D��|}�:F�!K�R�Ǚ����q�3�2��X�-�9��՚���X��\L�I2rzAtlS�]H3x�'���D������U3.Q?%�
�	�%��g����y�A���NOI�Zd��y"+�O�2j��IS�j�F����|,RJ¾��N�����O���%\&NOHѣt��w㳽�n�N��Um�W���;	+�`��Y�=i6ğ-{�5a�D͒�����~��@��������D���=���TV I�g��8
��
��L�>֩�����r�6�U�m��J���J[��y%m#���`Q��ھx�������B�=Td3���a�-����O�_���}������������q�(,.LC� ��q?z]c{�#%��D�5��[�\P��r�ŭ�yc�]���^6V�n_�7 �������1xM��M}c����,���/1�v?[���%��vϡ���j7�ݗ^s��D���L0��h7��@                                       $�:��� L�$��vB@ ���"1X�R��b1�5�tY��"��R�Ų���b�YVU���T��b�X���`��Vw���%�K�������%�m���o�Hn%#�+:�T�ڶt�7Η��.�]G!���[��-�;<�U��e�9����L������ng���������Ϝ����s�?;�}����dϿ9���xIK�����5KS�%/�J�n�Up�$f�F�c��Ə�c�,���~[?����#��|�H����(��3�$�83S9�5Sa�7S��9S��;S��?T	�B�TOC��V*g�h��ϩ|������������|E�/�Tt�j>�c�>�I��C��H�F<e# ���fM�+ ���PO��M�O��C�(��1I_#J��M;�[��j:����|k�ǹp�G!���,'#t�n�bC]�gS2�ί����d�X섵?V5�[E��j�k��5�[�y�O?\�4	wC�մ�'J���S��+�����Jgc�El�Z���:������7]�	�&���vOk�%��t��O�"ڧ��gv){��mG=΍�[RF �(6CXm��9�P�C�}� AA"P8[N�P��\��1@�<�������Z�l�|����e��N������d�_��o�Ǎm7�#͇���[�3���>+���J	g���?�1��BK�I��N��(�� ��+xS���T"{w��}���%%�&0�e9}��,�)�0�3O
Q	E
�ѻ�~q.Z�����NO2�,���λ&_L%�<��&0)�i�9��	�~ߑ���O��L�������FE�C���G�#���(��V!t1P�C�u�@A(s{�3��+�6���&dBlH������e��^K��LOC��8�	�H(R%&L��{�r��&��E�e���+\��N���l�>�V���kv+�Ǯ؍W�v�%~�eh��U����c6F��\ih6k]�f�^5���_��{d���f����u�&*g�,U���F'��W,�n��7\k�vo�Ʊ;���_5����,mVk#F��׆hz��ItUyq`5U6ҏ���b}�8'�B��h�������Zp��g�E@ԋ^�YF�6����ܒ�#�����0�0|&�����V2x�~C�9RFl3�;���p�[
VS4�0	��R
aXa|3xR��U�\$�*^*�U�Vu%#��̱��%�[��k�F����b�XZ+ƫ�f�k�-a���i��_���ka��Nv�]�f�S�4Ծ��K��:U?T_7�p���x�����"W�;�O��6:���6��w�+]���|�a��r�f�tԫ���_pݯW�M�Xk�6�.0��i仲�����=ϛ��2����������-7��`O1NAh��q�:¿�Չ	v���*f�Fs���(5}H֥/,�<�h��%����I�����}>C0�sB�J;�i����ґ}�B�<���a��B�:�yÐ���!��p�$���Xvvw!�Y�gUʖ�bu�e��6�T90�(��(��-.Lp+��� _CA���(7
 s(��U V���L@`*�hX��2]�:g��q�3e�e�G�4=��rD(��i������N%��pݒ�v-" l�F)�����C�8�rY���@�t���N��/�J�I��M�ߚ��r��v���\�"����1L�uG��ԙ.�SSV4��h����6���d��F��~�q�����y*�2�^b��^>�E<���K�qtM�����f�8�����~&����6� \�k�����c�s�SeM��b*���{�s{o�/0}e/��Ի[x��X���;C�s��{�g~{���_���{F���s~620�[3�#��&�G�����ãq(��\$�������^�E�:��D�Ɛ؋+h�^%��/w�<�F���񄅾�7Y]�H�j;t|�H�"g:`-�6\Vp��Xț�'�9~�˝|��?�
���"C�)��y���\�c��[Pd;���^�����d#�eZ��sɖ��i}�,"�����t��0�)��;�j�Wmx����fö��-%"�w�}<��դ��;V3�A�c� r�zW����i��s"،���w��5�j�M��cjR�[D��ҹ^\���.{j�=-�~�k��$kÉ�-�0���b�|=L�a��� �|t#���}̏�{z։
6J��X��wS�T�������E��F�7���-�:3k#ȶ��I o2�����C㰳�������6^"0�`�Ø#H$�u��w������/���d�b
�xA�b�.Ed5V�����>)ajM%���wđ�j��؎��U��7�r����!i�XJ/�
v�쨰W2qd]UN �b4�������(�G �o#���L�c}��TH��rRs���,�h�YYz;{��/6��G��ʺ^Eۑ{�;)�����6+��Б�ϊ���T���X[��p%n��C�Ze�yu���Ejnr#ؽ���A�d�+GJH�Z���N�5��/��KP��#1w.����r�J�����^3?^P:��~so��d:��X�}��^n�k�{����~�r�E�"�`;�!j:I"f�UB�\�3��,�
����Ès��*�Ȭ��6����� A:���(j��;� !C����XW���#���i�0X��O��	+�oB�o�h�g�!��_�����?�Cr�W���rd�ߥ�ʿv����y'�湎|�Y�<��Arv.����+��z�d�礖���/����h�X0Ťlcb�}�J	�zR�=c�毥~!��j�P�߫�Nb4y��$���CL��<s�W����� 8!`��':v,*�t,�p/�c@���X��Q�2��A�`C��pr�J,�,\;��Xu#���y۬�O�Y\�����ܢI���LeA2�����w�U��$a�@a �@���f�o	?�b�_�������$�����&��W<F=�+��c-mlf���g=E�x�xV�����>���|�X�Hx2_sk�����/���b�Ow,��Ĩ�8��!���@7�8��$=�3؅�v6R���`�r��gw��ޏ��V�Ê[��F�#xp"G�MO4{�����˟i�/(�*S*=��^ �	R���X���7OB�;p~[�R�^8�������#[�ޚ�X�[v-#z��u��jNj!^�vT��\�;�vfrcyiue۫��Kw��X��v,���U��o��&�θ0�67�=�ڴ��ϲ�{溳�������C8�)7�wJ˹�6M���}��m:�_ũި\F��%p�5A��n~�V�l��?�lWx֭u����:/��i�L��D�s�b���ݢ��X����+��Gu���UG��#�=�P��<��h��M�u�J��͛L�Vm�I�:�u�R����G�s�V��Tn�n3s�v����}��ѵV����S�+��V~�VӰ��S۩�L6f�s�Z�:�I�-�
؛U��WPoUZ�yE�J���ٰVp�m��<
�rF�R��l%i�4*\-K���}�Xl���	We�]�U��69)�9T�k�;�}�U8[^ݻr�UMΈ���`oUN��w����c��oƸK>���j���d�joM�+�<��qJ9z2��Rr��0�R�_ƥe�%�O�g%���
�z[��P�99_/�β�r���O/�,
`��_�M�^Z���'D�3�������hxh�A!���T�]"��E�V�����R�T/բc��u�܍ᅤ͓�(�3�ڠc�
����`�
�qU��Q�W��Y�u�?�j�=\�gj»찺n>��s��R��J}F�u[��V�Ot����K���bjW���j�<�%t}��KJLLK0��1����"�&�sl��������ҭOa�m�jm〣V8�����d��G�+RiU�8Y�s��)�'�J4�3Mԙ5?u�VkU�����3�k6V�o\�[,���߱�+�ͳ��;��itڶ��nw����r�������{����~/��p|%��p�W�q�8>;���whk�㔇�ynj���^��v/����}��'�uN��J!���>N��u�洩O��&Uj��x�*�b&�]�q*4u�˭G������V�3 �oe���0��i�ɕg�����]�'�f��g�gs������}?u����'�,��U|����>�J\���4ѧ!W�*���ǫe2L{��ȭ
ߧ����j�����&p��k i�yb0�>�d�o�c[��Cd��xY�h������w�WZ}\i�lcd/�R�j�gB�a�VC8k��;��� �0���S��^A�4�����}!!D@�94h��d.��+ �j��9�`����E]��`���a��5����~"D݋uT���a���pq��=�rP�,@�.�5wqwqwqwqwpW@�:x{�͵z�Kӥ۫�DP2q&�p+�a0�ȹ0� �a!`VD[�/�C��a�C
�x�P�D�r!�A���!�Xp`�ry���:�``;���C�qT��qT��qUDr
(⫈h�Q�X��%Y
f
U�h�J�����J���ق����B�L!B��!B�!B� L!B�!�!CYƹ6d��t�(Y��W@l1�ύ_LqnA�7�0��8l�!��w�nO_B�oƸ�!�n"�� p0�9�'L�P����rr��i9	^*qJ�ӊW�n����7'��q'!+�tN)_�G'!+�rp$��9W@N����"8���'��!�С��OBXl��b�yK:"z�
�yJp4�����L�b)�C�2�����B�2fd
�)V�钕p1�)WC9��#(J�L��A��J���(KYP)YB��Jo�R�x�!+��"�Jm�$�ͣ����BU?�$%W�>BU�|�E^ǛV�cu�+7�%g�����H��DT���g��$v!�?�!�P&u8�U��[��2a��gy4HbX0�3�W!p/�!Y�Pm�;��i�.��s,˼��$��3	��RQ�Դ��X���Օ��`�j�Mh�[	��{�?ԋ��];��l��K��	����0Q��}��|R��{i����Q��e��yw���5���cƒ�vN���*��NK�h��y뫾��	>�/1{]De�Z��xc���~���f�N!���%S����tm�9�{,���ұO�������{=����FbP%|���K��&�����W�`<\��)g\d���V��i\:�Q��mX������6�]����V*cyAz
#gh�Ft71��XR��+c� �F�#p��81���j��(��=��F�7��pP��i��݅�^E4{���h���t(l"�8��W�Q�j#����9��6a��3���ʊHڅhq�CY�<F�4��
���|]�\�8���5�{kqÌ�n��9�L�j��0�c_�T�TJAo �S�!/B�?!K�������T9���B�N!K����R�)l)yr����/�!K���HR��)l�)o�*	㐗e!K����R�)w��
^P�- �.�B�T!Ks!K���R�)y��2����
_�B��B�w!Kc!K̐����)ub��
Z�
]��-��,i
����M`���jCY�XVB�l X¨d��&#;�H��W���zA���0B�W	b�E('
8�
hJ@�)'֣�)�0*
 ���H;��n�MMN�����O��R�UET#��3������ETTU��5��u
�"�|R�UK�R���a��S[�.�K3�k#r�QD�(��*�c�#O�Ğ<E����W��S�Fo�?���NJ�����k��Yz����󩛽^C�����;�e/֋fl��)��g������T���R;߁���:�=A9E6�aI2��BJ��A�ֈ��V���M2�y�1n�Z��C<��ʝ��?�Q&q�T�>q��x��;�3�.h g�밁�,,q�W(s��$�Nf1Bh-���,b-a�8�@���!
0�s�VXӭ!�9
O��L�L%P�z��h���I�E��{��zʏ�AE���*5+��(J��k:<p�|x$?I?t^hI�m�c�҅����?$�����w2.���gb�/ɥ��p������d��X��>�{^]�yS�T�=V@�������ܝ�f����Y>|=T22�Uh��;��|9����M���mԺF�l�.�݂C����1}�y�=�ƻD���zՈ�rC�J�h����.�K���y��IBCϭ�Y��GpٷZ�}Q�șb=G�Y�} �@��y�	�]���R�\�ּ����T8����~R�G��PO)߻�t�eL��elC��$1�S���K����䜯E<��*l�<��!�'yT��)�Q�Cԓʧ��Ǩ�
}J������CÙZC�N��sQ�2�G��hU�L�T�MȒ=C����L�"�A�i�c�����R�R��q(Q�H�B� � �!���(�␤cjC�����wF��̤1�T��Z�!�5C!e8�r`���ɷX�{�>h��P�ڹP���k��R���>��ߪ�?R�}��#U�iJ�"=[3�y	�rª���_�<2��Y?M���I�_S"���2a�7�0����k��;�H���G����`%����2CIU��a�3���� �xu`/
�j�}����A�P�.Ң�ؔԵze6�k6��?l�3���=�
E^Ѵz��V���{Nb�����X�����u_y�3W+��Ǭ6��Z�fc>��������>7��]ay8k�����q��ฮC��y��g=|8��m�w$����{���|]��7l�7��o�;�����}�|+��]������W�~c��� [���3��w=�*���u�qp�vkV���-v�c��ߴ9�"n.�N��v�7�ξ��s��܃�;�����+�r��E�湻�Q磻��Kvܭ��׃�����v���;A׍�~ؾ#��[��n.w.v�Ⱥm;&�tw�|^��ɧϏ��D�\!� ������L�6��d<�S8����?�ic����.�`fӫ�>�W�^��[����fi���9�o��Zޭa�l9��m�f��Ơv���~E=���l��k�J:.�J�^m~���{���F�nk-�&�<���{M]�����&�P�/3=KXNUY��jF�X��q�����%��&?��eo>3�����Ü�A6uC��^�-�ۋ����`o��n��Ĩ�)p\�/�d�AG��;�9��R�`������V3��E���K���:��T=n�Y�J��q�S۫�ǒ^HlI����|k�Dy �����N���;t�꿛��ԣP�ѵB/!d!�:�Ts���3���عA�V�d��:��r�ʲ(���m��B�^�u�VCXq��A��J:�Chu�C��K�-	Y`r!�C���`�$y�_�s�}�S�/��"U��C�7\]?�n�������j"_�7\a�_��({��OVP���|�n�������c�l��ꭚMx�w��1��įiш�,��\*�����T#đ�@A+��EZ��3��ø{�C��N�-��C(g��:��� �88���"��=��xgڦ4��7 ��x[W��	�
e=��k_��o��﫜\p0,�aBvE�Ig�̓��@]�DWa�MV�Q�O׉�'x�Z���)s�I_���R�PEk�4�2I��W��:��P>������`����<na"	�	�rz�f�c
!�{�#?VI%�ar�1�{iW�F�cW�Y̤�T��֧��s���!�iI��3R��&-_UGf:'2ɕ�#�ң��8���6R$�D2,��{�4��S	�Q6�Q��n�k�$r%�JH�ϔ��$��76��.Y`�۱��_��Ow�|؎�Ѳ��"�������yī�u\Ի.��!`��q����/J�{&w�����y#ۦ"�Z:�nmWE5��#	fd�'=�M%s}� �';��e�"NyD�e���J!9�HH�	9b`2��By�A�Mrف[���1�D�-B{��0!��}�C"�&6_�AJ��t��+�)�7_��	ʕ��I�y9-�F6�,
2y+�Bu�L��m��<���Nh�َR���|�Yo��e[�`�9��G�A�(BD^�*�,�)?"P���SG-L%�t�"�2`B��ZH���I�Xr��Ρ'l�h�&�S�.�����ΌZ˰V��N(�� {��S��a�H��5�)��dI�h쨓~H�6X�1N����4ӎS�F�h���r�F~�$�2�p�96�P���|s�1#�Z��XYNz��^��[$(9INL�0K���RE��T�9NLm�ʄ74t�mF��E�9Za7�K[%���e���Y�[D0��=�!3�H�A�I��Ǵ��)*HՓ��H)�@b�!6I�1�^FO��af^�Gϓ�@$I���S�e�¸N�IL�4;�oSĒI�U`r�uq�ɘD���#��e%��d��-IA���ЎK'T�~���0wl?W6�P�5�X�L�����8��R٦jN�/�]$S�娴�2R�!���D6zGOsz,ڊS�IJe.Y'#h$�u��0�oFOR���K�	c�$C�I�YǉV�	�8�);��ZvD�:��4p-yå�J,�&��Hq$�v	�;R4ו!8��`��b�r4�W:�C{�Y
�����A�M�E_
�����K?�t,2:o�
D:���������q��+Y�<�8qNM�v���E��!'�b�"��:䡟����5)/I�߸LH���4�Ԝ��y���d��{��8�Ns�Wd�R��9��RG�;)*t.���VV0�4�����
���vɮ����eƹ��&"�Kel�JLq
��"YE��(W��Y=����A��[�Y���<:h��V�jg�$��C�2ut�dGˡ�f �c^��)�Ȧ��'ݥ*���sE�M5����U�1(V��y�e5M\jR�󊤏���$da>��"?q-2��'����s�>��4&	�5�)l��ʙ�>I��.R�++rR77vU���QPS��h��S�&L�EQ94�&l2
�M)y�&	rp���bB˒zk�i="@                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                               C3�( 3E���1�f͌��1�g#�1�c����iv��"�.g�o����ny�V�1�1��I��<4�Ê"4�]x'M4�la�Fa960�cM��F0�a�g[��6�<�����>td�*h)���0J".ڬ	DRR�-�eR�R�	OJJz[�2�[�''>���|뮻�����mϟ��������%���*����K���=��qW`�!q���W�b_��[V�%��y��R�w�e���S��`~��^���ޘ%!@����_���{nA��n�F�������T`���`��B�0W{��{�`U{��@�邶Q�������9��q�0Vq�
��>�+�O�7t�m������`��ʧ��V���2�-C�3��A{��ȿ�?���!�h��^��p��'��\&C�!:�s�v��Rio�?�AW�s��,��-��;A��a�j/�q�������|XE�u#�Qy���d��P;�\AAϋ(��]��w��k���Pr���f8��]��w��O��(9a^Bs��-���탗G+���S�{�FF�qm1��3��Gf���h��P<�`,ذ�%���B�?`��I�H��^#��>�."�;1ڋ���x&B`��8��]�^��X��*�0U*t��΋(�zS�P}�_:S��փϪ��w�P9��@���]�f;QR�����J�y����X���C�`�6�,o#�������@Uaر��"�>��C�}��p}�w>Lߜ3��y����(��@����C���f6�@a�1V�	�n�C�������G��SU�EX>
�Rf��y�Qx���'���	C�!͋ ��[��\��qy��~9�O�X>�!Ύ�u"�:�w��+��2{������:sϽ���$���B���}�,tXŜ[��v"�;p��7t��J+bB���f;QR���?	�a��a���O�\;|.��p����"X��[^.ô����$q�G.|ZR.b�.����p�̝?�c����-���6����T��Lu@��J�� ���a��୳&��T=��p��8���v"���*b��0����Щ[�R}T%�H��Z�]�v��8n�*b���u�=`cЋS'�cv�e�qdӜ3�	Ex,�:�p����T���u���w�p�/Zy�N��ׁ|c����b�C��f�rQ��o���V?��f�t���p�A?��]G::!l1���{�c�~yFT������bfm�]����a��WY��Ŋ�qr�.��/�ԿD�g8���0�\)���"-k�}��}����a���{�=���ad������_�~�5�i$���p��Rc���U��q!D!
�)�����ղ�]!R3k+ߴL63Ym�4�.K�U�$�ĝ���Z�44{��)&�)���+�c�r�6$�^���@X3��8��L)�TkՒ\�Ďo��,�V[)iˈ/;�L�nT&)<����K.|��Q
ӓ�{�V��Zٞh��
<��L����))��X���#8A�9���ꉌz\Y�V!����d*R��8ƿ��${<��3#w��֫��������%?�j�l������rr#�ʿD�V<+RbL�֬H�B���q���ù
�w�k�XS�
�	����NtZ���?������Jj���m�D��C�)kf�y�Y�}�*�����B�,vT{)������$�XDW�vh̊�o�V���}P���XqF+�J/��1����k�zVT���qm��/�)8h
4�W- �4�̇ߊ��1	�4���+��*��ej�GfeX��I�g1:�lڷ:�1T�le ���q�M
Q�/�&H��.DcEm��(��]��#k�d6u&�t���C�ˉ��"��b��^[���+ƹ�:rK��o�,\��ծ��-qS�f��~�9�~��_Fq�:�.��Y��iY*=5�s�-�l'���DczDiM>ϣU������|��Ǔ�W��MLT{g$�����	E�� g`=���zR�>P�xn��lAĚ�	��ZTɛ���*3zGD�׾�����z%!��G�/��Ș��XscsH��	̦��bg��W@9�Y�ǽ1��e��Z���;@�����o�IJ��؄e�vz��	g`�.���Tüԝf�Hӫ��<j���1��k�Ew��RI�Ь@�����F
T��/�BU7L�L٬�e4�/VMe���t�(vo�,ֆD����'�����98�y"��GG��+��k�%`��6����,�i}���E2��l�Ɣ�?��g���F����N`��:�a���(�OcjR�,�����������"�1s����k"G�ҧ����̽�l+&��7��7�to�"�(��c�׽]�ݝ{����H�^�E�E��>#�F�i\�M��"q1�efU(>Ǩ��y��U~@s0���6�l����/��B� D_���E���ƶ{���j/�ƴ8����m�k�Tl��`�C��)vN�\�fign��4��-�6.^�$�����ԣ�2mx)v�q2\w����x9y�и��!&��8Q��xu�IJ&���{�u�d��̎���l���:#Fw�|e"/��?����W]���	��iC��B�׊�}��b�Ek�nMk9��#n������G���6����^@�+�rߐ3�\�~2�ZD��\�T���7,�sJ���`�t��8��?�}��,�E�T��������#�D[�6>"q����ˉ�e����;�ƨ�,��{��!q:6�#���g�R���>�7�Lf�<�����Д�zJ����vIv�.y�;�M��cX�@��AQ@�<������T��5Q��fKc(̝�EK�ڥwՍR}����4�PM��HQ.Ԩ̀��o�q��+�dY��㉚.����ύ���e}�����������աo��"J3�&�[(�ia��)Q�F��.��fp�z�=~ me��
�$���.��9͌J����B����jm���6W���d�ػ9PH��?k!�S�~���4;�Z��`�y:�R!6ݻ�_v%:�ؔ�`���C��U��Or�3q�./����1^(h�dCh�de+�%�z��"�A�q�LJ��o�>bW�R��O�0�Î�~��7(�DEҐ���4�}�N�ӣ()��Erf�m8�L˞�VVd�t1����{H6g�m�^��rP;а�����x�ޚ�L�M�7�C����z+O;)�2���{�zoG9��h�z�g3��R�5�V��VW\Eĝ�=���o#U�V�O�:���͞���� 	��r��~�9J$撪�6��z�?�&nwDO�]L�|�%n���i0ڕ�Lw�*N1^KB�C�zW�ɜzc>:L�Lo���O�����.�<&{5i$��������K�r7-G��v]v�$��	�J)n�d$�S��+[���Nq�2����vo$u#N-Fx��>)�,�5��ݕ6{�Ki����=��Kӕ�GA}Q;eF��wM3�O,�Ҷ�����i���0���݇�ˍYL�������S��3��X�*�7�Q~����������ԔUXJ� |�V��Q3���S�lk2C�e��ӫ�R�!|}��rV���Ⱦ��|JM�A Z0��I���ؔ�J(l�e���[���Ӣ(���T��4>����S#�̛:gly�{�f?�M��)���'��3D��S�#�Ye�B�B�.]��y�(�l�c��E��SJ?�Cy\������%�V��:A�9gn��{;��.F\��&�V�/:�C�U'c,����^h�k%C��f��A��
�eZ�+>��8�4�P���Ĭ��l��/���4:s��q�L(z��8�^����]��`���魒���:�a�)�#uG�<�_?f���%�q�2B��|~�]J��+c�HU�O�Ep�-mIpٺ�pᫌ���j[H[9/t��a��K���@hО~}ĕ(1��0[Tq�jϋ�R���T8�+����.~+���I�����+��e�f�1�E-O�� ��Ǎ�uUe[�[���i+Hn9��i�"��*�&E���'з��|h��^%A}��Y��QP?���L��
1f��!�d�\Q�A�ÿͨ[�w��ۨ��*���)B+5��.����_�C~�yr���~��=yݸ��Z�JcJyf5d�*�+�Z2w��ڵ%�*�-8��
IH�iχ-���Ϥ´q�t.}��ӱ8=�J�O�ἴ��$i��۵��&�`�决�?���;~����i�F�*J�[�I.���I��$y��o�������޺��~�9��
ю�:�p��}�"y��c��iw�ϗ�{3bg���9k6�I����x��gӱ�?$��g7濈�?1N�4YkN�4?#�1�]��l����ɦ+�ia������m��F3)k�A�_�FXUӓ����9g��>������I�$��0������o�� �B�?B���+��|�u;1{ǒ7>p~X�
��L-A4������l�k�Ǆ�����7���xe�a�V�8�vB���qR}"�3n
S|^��7�>V�6�3�㖦QApV��D�,��o"X�J���l�4�{��L�톦�Q����qq#U7P�̃�����D��ffC�8)�.s*�3\Ł�U�by�8�:fG�OշZ�%yy��?�j&R.�	Tj����wo�Ɯ,;�3��(����>�                                                                                                                                                                                                                                                                                                  �Z @�Z ��Y �Z                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                     BR6          P  �   �  �   ` �   � �   � �
   � �   � �   ( �    BR6          @ �   X �   p �   � �   � �   � �   � �    BR6    W   p! �� ��! �  ��! � ��! �0 ��! �H ��! �` ��! �x ��! �� ��! �� ��! �� ��! �� �" �� �4" � �P" �  �j" �8 ��" �P ��" �h ��" �� ��" �� ��" �� � # �� �# �� �2# �� �J# �	 �`# �(	 �x# �@	 ��# �X	 ��# �p	 ��# ��	 ��# ��	 ��# ��	 �$ ��	 �"$ ��	 �8$ � 
 �J$ �
 �Z$ �0
 �~$ �H
 ��$ �`
 ��$ �x
 ��$ ��
 ��$ ��
 ��$ ��
 �% ��
 �*% ��
 �L% � �Z% �  �n% �8 ��% �P ��% �h ��% �� ��% �� ��% �� ��% �� ��% �� ��% �� �
& � �$& �( �>& �@ �V& �X �f& �p ��& �� ��& �� ��& �� ��& �� ��& �� ��& �  ��& � �
' �0 �' �H �0' �` �J' �x �d' �� �p' �� �~' �� ��' �� ��' �� ��' � ��' �  ��' �8 ��' �P �( �h �( �� �*( �� �>( �� �V( �� �p( �� ��( �� �    BR6      	     �   ( �   @ �   X �   p �   � �   � �   � �	   � �    BR6       �( �� ��( �  �    BR6      ! �   ��  0 ��  H ��  ` ��  x ��  � ��  � ��  � ��  � ��  � ��   ��    ��  8 ��  P ��  h ��  � ��  � ��  � ��  � ��  � ��  � ��   ��  ( ��  @ ��  X ��  p ��  � ��  � ��  � ��  � ��  � ��    �    �    BR6       �( �0 ��( �H ��( �` ��( �x �) �� �) �� �) �� �,) �� �B) �� �^) � �z) �  ��) �8 ��) �P ��) �h ��) �� ��) �� ��) �� � * �� �* �� �** �� �J* � �Z* �( �l* �@ �|* �X ��* �p ��* �� ��* �� ��* �� �    BR6       �  � ��  � ��    ��   ��  0 ��  H ��  ` �    BR6       �* �x �    BR6       	  �      BR6       	  �      BR6       	  �      BR6       	  �      BR6       	  �      BR6       	  �      BR6       	  �      BR6       	         BR6       	        BR6       	         BR6       	  0      BR6       	  @      BR6       	  P      BR6       	  `      BR6       	  p      BR6       	  �      BR6       	  �      BR6         �      BR6           �      BR6           �      BR6           �      BR6           �      BR6           �      BR6                  BR6                 BR6                  BR6           0      BR6           @      BR6           P      BR6           `      BR6           p      BR6           �      BR6           �      BR6           �      BR6           �      BR6           �      BR6           �      BR6           �      BR6           �      BR6                BR6               BR6                BR6         0      BR6         @      BR6         P      BR6         `      BR6         p      BR6           �      BR6           �      BR6         �      BR6           �      BR6         �      BR6         �      BR6           �      BR6           �      BR6                  BR6                 BR6                BR6         0      BR6           @      BR6           P      BR6         `      BR6           p      BR6         �      BR6         �      BR6         �      BR6           �      BR6         �      BR6           �      BR6           �      BR6         �      BR6                BR6                 BR6                BR6           0      BR6         @      BR6         P      BR6         `      BR6         p      BR6           �      BR6           �      BR6       	  �      BR6       	  �      BR6       	  �      BR6       	  �      BR6       	  �      BR6       	  �      BR6       	         BR6       	        BR6       	         BR6       	  0      BR6       	  @      BR6       	  P      BR6       	  `      BR6         p      BR6         �      BR6         �      BR6         �      BR6         �      BR6         �      BR6         �      BR6         �      BR6         �      BR6                  BR6                 BR6                  BR6           0      BR6           @      BR6           P      BR6           `      BR6           p      BR6           �      BR6           �      BR6           �      BR6           �      BR6           �      BR6           �      BR6           �      BR6           �      BR6                  BR6                 BR6                  BR6           0      BR6           @      BR6           P      BR6           `      BR6           p      BR6           �      BR6           �      BR6           �      BR6           �      BR6           �      BR6           �      BR6           �      BR6           �      BR6                  BR6                 BR6                  BR6           0      BR6           @      BR6           P      BR6           `      BR6           p      BR6           �      BR6           �      BR6           �      BR6           �      BR6           �      BR6           �      BR6           �      BR6           �      BR6                   BR6                  BR6                   BR6           0       BR6           @       BR6           P       BR6           `       BR6           p       BR6           �       BR6           �       BR6           �       BR6           �       BR6           �       BR6           �       BR6           �       BR6       	  �       BR6       	   !      BR6       	  !      BR6       	   !      BR6       	  0!      BR6       	  @!      BR6       	  P!      BR6         `!  � 4           � 4          T� 4          �� 4          �� 4          � 4          $� 4          X� �          (� �          � �          ܨ �          �� �          |� �          L� �          � �          � �          �� �          �� P          ܹ 8          � (          <� 8          t� (          �� 8          �� (          �� 8          4� (          \� 8          �� (          �� 8          �� (          �            � (          H� 8          �� (          ��           �� (          �� 8          � (          4 (          \ �           	 �           �	 (           (          , (          T h          � h          $% �           & (          4+           L0 (          t5           �: (          �? (          �D (          J (          ,O �           �O 4          Q (          0V h          �\ (          �a (          �f (          l (          8q �            r �           s (          0x           H} (          p� �           X� �           @� �           (� �           � �           І (          �� �           �� (          � (          0� (          X� (          �� �           �           ,� 8          d� 8          �� 8          Ԧ 8          � 8          D� 8          |�           �� 8          ��           �� 8          �� �           ܯ �           t� �           l0 h          �0 �          \0 (          ��/ �          �/ �          ��/ h          ��/ �%          T�/ �          �/ h          � R           H R           � �          � d          � \          H            H H          �  �          <" �           �" �           �# �           8$ t          �( �          �, L          �/ �          �3 �          46 d          �9 �          �= �          @A �          8E �           G �           �G �          PI l          �K �          �O x          S �          �V �          \Z           p] �           (^ �           �^ �          pb L          �f           �i �          �l            �l  @          Ь <	          �            �   &          �            (�  G#          p! #          �!           �(! �S          �|! �          �! f$          |�! 3(          ��! A(          �" ��          ��" �          ��" �          ,�" Y          ��" �           T# �          # �          �2#           �N# !'          v# 
7          (�# �R          ��# �k          �k$ I.          0�$ ��
         ��/            �/             �/            4�/            H�/            \�/            p�/            h�/ �            B B A B O R T  B B A L L  B B C A N C E L  B B C L O S E  B B H E L P  B B I G N O R E  B B N O  B B O K  B B R E T R Y  B B Y E S  B O O K M A R K I C O N S  B S D B N _ C A N C E L  B S D B N _ C A N C E L 1  B S D B N _ D E L E T E  B S D B N _ D E L E T E 1 
 B S D B N _ E D I T  B S D B N _ E D I T 1  B S D B N _ F I R S T  B S D B N _ F I R S T 1  B S D B N _ I N S E R T  B S D B N _ I N S E R T 1 
 B S D B N _ L A S T  B S D B N _ L A S T 1 
 B S D B N _ N E X T  B S D B N _ N E X T 1 
 B S D B N _ P O S T  B S D B N _ P O S T 1  B S D B N _ P R I O R  B S D B N _ P R I O R 1  B S D B N _ R E F R E S H  B S D B N _ R E F R E S H 1  B S _ B A C K 
 B S _ B B _ D O W N  B S _ B B _ U P  B S _ B O L D  B S _ C A L C _ B A C K S P A C E  B S _ C A L C _ C A N C E L  B S _ C A L C _ C L E A R 
 B S _ C A L C _ O K  B S _ C A L C _ S Q R T  B S _ C D R O M  B S _ C L O S E D F O L D E R  B S _ C O P Y  B S _ C U R R E N T F O L D E R  B S _ C U T 	 B S _ D E L E T E 	 B S _ F L O P P Y  B S _ H A R D  B S _ H R L  B S _ H T B 	 B S _ I T A L I C  B S _ K E Y 
 B S _ L V S T Y L E 
 B S _ N E T W O R K  B S _ N E W  B S _ N E W F O L D E R  B S _ N E X T M O N T H  B S _ N E X T Y E A R  B S _ O P E N  B S _ O P E N F O L D E R  B S _ P A S T E  B S _ P A U S E  B S _ P L A Y  B S _ P R I O R M O N T H  B S _ P R I O R Y E A R  B S _ R A M  B S _ S A V E  B S _ S T O P 
 B S _ S T R E T C H  B S _ S T R I K E O U T  B S _ U N D E R L I N E  B S _ U P  B S _ V R L  B S _ V T B 
 D B N _ C A N C E L 
 D B N _ D E L E T E  D B N _ E D I T 	 D B N _ F I R S T 
 D B N _ I N S E R T  D B N _ L A S T  D B N _ N E X T  D B N _ P O S T 	 D B N _ P R I O R  D B N _ R E F R E S H  P R E V I E W G L Y P H  S P I N D O W N  S P I N U P  D L G T E M P L A T E  T E X T F I L E D L G  D V C L A L  G E T K E Y  P A C K A G E I N F O  S E R D L L  S E R E X E  S E R F W T  S E R T X T 
 T A B O U T F O R M  T B M P T O A V I F O R M  T C O N F I G S E R V E R  T E X E T O O L F O R M  T F I L E N E T  T F T P D O W N  T F T P U P  T L A N F O R M  T L O G I N D I A L O G  T M S D O S  T M Z F O R M  T N E W X P S E R V E R  T P A S S W O R D D I A L O G  T P L U G I N  T R E G E D I T  T R E G H E X  T S H O W P M 
 T S Y S S H E Z H I 	 T U P I P D A T E  T V I D E O T O  T W J D V I P  M A I N I C O N   D;2�" <G���c�o3����HZܒ��(9]��f�^z��:p�v��޺�v��S_�..�7s���5oE�#��D�Ġ�X�rՈK���w�����q+����7$��3������C��^+sM ��cn�$г1�drZX�,����)����^؍��T�S�mT����ݪYB+Y�hYV�8�U4�%ˎ�������ߟ<�������������ߟ?><��U覑mX�fUN�R����պTi�il�O59�NL�fQ��ß-��˾�-e����+���W���WǇ!��A�5��zӃ��j��ު�vҦzI��φs�j�8:��>�#d߆ַ ��'kq�w���Z��aY��iAH���`�_LO�'�_ 軏4Y�^AO����Vٚ�jXjǔ�s��ȆKA|�V?y�j�Qs�a��d�ʃ�'���a�d>\��a�����m����$]�/$�� 2[!�r����q��t�^B|�A�	���Vk��5�&�V ��Oֹ��D�Kq�0�+hKqo5���z�)�~I��9����EU��J��cBiN�sr��J�@Q�{�A�?���_��������~}ѳ����	n5*9�=��S�;����@����Se�ssBhƦruۉ�M6^}O-C~(�Ѫ��:�6����eq c��F1���d��#ܠ��Q�޵���o7�M�}W�6H��&G���E�4�u�?�;�1Ybi�N�����}�0��{�@������?��$Ol;6#��R�S�n������ͳ�/X��,k=W����{�|���M���e*����Pr:zҜ�-�
���y�aO���޾ڢ�X�s�5˥+����*Փ��\�Օ����˞t~�
m_�|ێfv��εP���;���u��ٴ�=X�ME�a^*�/���ͥT��姕/�`8�qlJ^?'��u]�����~�U.٫�5֋����,;F���y<W#��oc�YO��^j�ws���vl�m��lZF�}m�tR�=�/��̘�τcG�5�q�&�n]�uYѨ��]%�Z��^�}W�c��+*�S�[�r��W��_��zz%(2�zjn&�7�\�Ϙ,��԰l��\W�����f�[už����������yv��ԯ��:�$���&^��Z�]:�>�T�c~P���9���k�h��k���O�����������Z�x?#�{���v�D�.��������EZ�y��/�cVy��3�޵YZ©v�����p�p�ύA��X;5��]�n_��eֻ֏���#�
����*�*����Luݥ���-�d���7���r-r�m�7R,W�-_���2md��Yq����P[��u���;��Xk�U_���}�/T�m�B��Xv��i����%��]=ǵ�丼j�y#��-�:�ִ����wD=!u�����&|��F��gv%�L2�������,�7[�R3|����{�;�|~��^�B>����m2͔}��/�Ë�V���N*�&���Jh�H�%n/��Y�_9�X_Ƞ�1���8�6&И�Z՗����X�k�-���O�,�6��YJ�$�?I�����>S�6�R�R����� |�N��
�8�����o�_F�3��^��Xy��L/��S����J���KWG��j�bF0X�:����Ŀk��� {�E���pI|n�>�vf�lR_Ԇ��|L��5�{�����F���%-}�)e�V,�Z�88 \�ԕ�A�K������������h��v�#��U>�r&6z��,C���\M���z�ە�ܸ���L�?�٢PS�d�}��UE��c���'O���=�M���6��y���-�N�?A>^��3�<�z�|�F������e�`U��\?��å����F���.h�3����z�;Z>j�}��~������o�����������t6ZM���9+���-&����UF�j�V�	�}i]%�]�#�E���Z��������1W��E޻;��oA�j|�P�ѕ�c�m�*�d�����Ufk(��k0��(V��_̋}��2��@��5��`�X1�T&��C����HfW�hB�I�tA��`�ꀩ��E(i�CM�������H	0ʥ�&CsAH���V��#取>_b�\���EB�vh��^4i��)��͜�oF��c7��oo��F�����oOg�,�DQ�f��BTXN8���zv�YV�e�`�[�p�U�n����x�0>����e�V{p^���]Oi�X��	��<g�a�P0����+[	��0�`࠮o���ڒ!��o��v��	u�Un�F��o��g�ѣ�<��;��X6��	94�ICD0�
p�
�� iC��Xĕ�D�%�0��M͂rp3��DT H�	�1,|��>+�5s=�A�Z�f2ӹ��sy8{/�T3�Մ��EϚNq]��c��҇.t��a��l*� بƷ����vP�j�Y���������0��}@�ع��?Y>��6r���m�,6�1$3_7;�UZ4ѭQ�*�-�印��c取>_�%�UĹ���P5�UzU`��r�"U��`A�1���E���{��Ŵ�ȕy���������tA�˄m��Rn7+^��D�'��`3JG2�@J*��Q���p	¢t
j'���D�$�*
r���K6©h�22��%�G; ���,|�<dmsF[A��T�X�2�Äc7��?�Zli�fq1#��P �H��M�,�ȅ�Oƿ,rUD?,1q���KN���XE�ߣH��4Y�S-V��J�\���S���/���,�'��X�Ȫ<��j�,>��6�
����]a�wWN_Pv��
��dZ��eQ�[[�m��J���-��v�

�8���`f>X�c受�a���D�J2�L��UVn��/�r\L^����L\L\L\LE�2�g:��%�=��9�����>X�o\�v�FB�XH�r�]41�����Ȕ|�\$9f��|�f�OFv]%�� }����B[�1�An�g�uЖ��2<�85|Š*��E�ߟk�++�_`���Fg���B�
�>\�xdb�XH"m�K�r�^�4sz��#�i����⌀���v	m#k� 6�X$/�3�m��}[?���]e�KF!��?�k�f�<�S�S��
?|���"
P �@	�
P!�B	�R�2z0!F�J	r H��G&��I*��I.��K0T�Y�Qj�h��)�Q�r�p��ӥOQ�0vU�)�D�	$)*��Q����>X�z�̕so6�IH�{���ӻ����I��?u��_�u��L�~
����Ϋ�E��4KI+u��yw��[$Bx�ބ��p-�HZ�"����Ѭ�@�*�b������/�����������^#c-���m�B:4q�%h�^/���x�W��3+�g!}mdm��2��f�!������9mo��)��+%�j�\�V|�S4h/�h.�M�i7�3X.r���nl����}��jX�c受մ���%[�NX��ѡU�c&�38��d*�$1������{1���
��Y�&>v�Ϣ��ɋ>\���.w���]������d��G���>_�%'\�V�I��+=�I��c1C����$����7�x�9G#o=��)}_=:�V3��.@p�H�%�Ȩm��Ծ��������R���ͭV�[Z���7���:F�p�+Kb�B�#����$"�١��� ��w�P�l��o�͐e�?_�kυE5��ɕ��R�eI.��]I���}�;I�Ό�1����89������h-ϗE��~�X�c�}
��AmBk�Lݜ�2��a����[W
�
�y�7�=�OmH_T��q���e�ڏ�]�^��Bcϼ��gS���O�k}b����A?�YY����?L+���]
�
d˥k\���pݵ7v��Wki��y��co=�������6�(�ӹ�v_&p�d3�4�l��<�
@�Ј.m�A��d�B��QFk%$crƢj���C�mبG웒�I+c5%�$R��4`�L	t��d��`K�a:ɦ�%��M4�`B�T�9�gD�2�x�R	�%NT) 7Q�<�%��)T*��F���@$h�5�!�0B�jURRzeE)��*����U`�W�TSuخ3,|��k,S��N�J�GO�8�n������ݘ���R��'㼣j�܋�~?��|T����A#�<o ~���c�1m�6�/���|g���e[k��I)��l=���/�`��mc]J���|n~�2���j'���/8G�s����c~�,���x+�i�&4���\ǃޤ��;�L.��x_��O	�#:y�7��{�!�Oǔ;���"pe�O��3�$W��B-4��;�4������Q�c�+ztt�gnڵF5�I۾���Z��a��3$�U����&�5GΟ�48��C�@9 ����uL�BbA] � �A�2�0d`�"��D�'����W@ �3Af� �A�2�0d`�"�U&8`�:�`�"��D� �3Af� �A��-���+�]�`�"��D� �3Af� �A�2|3Qa�t� �3Af� �A�2�0d`���Da�V�7A�2�0d`�"��D� �3O�*-��@nW�3Af� �A�2�0d`�"��w$��2�/!�����s�`��Wn�e9ܫ��&���7�KD�A<Aj@�9��#�����iJ蚨)۩ *s�)��l X����aD�
�5Q�S>���nD��D0�
�y��"Ԃ�9�FI��i)����CdR�)�QMPi�L�J�� �R)U�����&YRj��4��?��Q�qT�vƤ('��t�5|�udAG�
�)E*b�=R�����IJ�����EY�P�KM���Ӓ�˫�x�����*�[o^�k���H�pG"���>+ƿ��y�8�����o��<�>3�o�_!=�
�A�0x_�4�E�����W{�y{{@��=���|����E룀p���{��A̖�l����J3��u�>*j�(��b>X����ڹ�+3�X՚��g��Ϋ��ͺ���Ѧ��mu��V���эv�]���C]�����<��4Ҿ��x�{�0!�$I5"U�y4��J�N�I )Y�e#F	�č�eO#NU7�0Q(�N�|�X�1��c�J,�6��^Tfn�Gg�`k��dq�c��r�=�X�[إ|�Ƈ������s��UL�8eZ���h�4b���)��W�0�qp�Q��Ђ]8T5)����R�@�U:
I�,U=c	-	H黸�L��>X�c�2�~PtT�N��4�N����N��X���o.�(���:]4Q��A����5�Y!�hn�~��叢js@6��Tu?���u|t�i�I�M]ڪ�gr�Whi��}u8]����� _��cc}�g�w��8��S?�k@��9Q�U��^�>e��+���abV-��k�k�u��~,|�����x�3�q������F�Y�fM���ӆӦ�ۜ����n�r��U�N3+���߸�i\v,�����qv�l���#�9OQ�4�s����7�W�_�_��s�͸^9��c\&WZ�-qm-��[�_a(|�ȔX�c取#�zF��k�=?'��Ig���\�k�o�ᕦ�u�[���)�V���R���Վ�H�S��Y��+Wi�����O�^�c��g�({�$��j���	,��Th���x�ȑYT4&)JeTʓ�:{�u��T����@�*E ��T�
�����l����/Rj���,}��}LnX�YH�R&k�g���@�%�h��n*�� t\c���@���q�؀v\�� ��AD�#q�>�կg��왲���4���k�vf���]ڏ�,|���������Z��O)����\�l� ��A [6�R��k�鿟�����@�\	怓��,�͗C70d�wE'���DR�	��T��z�>X�?X�]K��:�4뜝]3��A��Ĵenő��B�<:sїy{w��z=�Z����]��ֵ�ޑuo�Ζ;5��Q{s�iޏ�B��,|�������,~��>������g���mcO��������d6�/����xn7��&5?0mL0�6��|�'�׬��0سƫ�8�Eq8�Lp<qes[�f�<��L���r�]8͸����[ݙp�;�B��,�� �v}��س㽽��|zv?������B�6�+*f���/�,����p�v�!F��ٖ��i��9���Yhh7]�gz�U��4�z�_�n���^�8v������œS�����_�|��;]��9S�T�y;��'�z\>T���J`y3��A��s'�]�Ӧ{���+�9R��,|��l���3q���`7���Z�8�*a6Щ�;�秳t�E3:�����,��j#(h@�4(���H: ���3�D�@�"@Q�0R���hR��y�@%hb� (��ɔ�6h��A��*2�q((�\�4�Uy�+�g* %"f� �3��@צ�:��� ą��&L%��1�ԶQץ�(�qR**T��L��:�V��*�:G R�le�@��`O'�#P}~!�4�mzb��TcL	�ͧ�f�x3�@�¥��]"�Z��x�GL1M�t�Q��"H� P��	P>����d�z�/��:Ӫ�4L	���)�j�S�D�F��H�LT��
p��9P@��b�����oW��<�t<o�.��}�S���,�D��.��$t6�	������A �+�^�3[��4�_��o��&R�_�I�g*8?��2ť�"�tz�|�fPo��#�k���?���E/�L$����8�!z�x���`���}�\/��>_��\W����1�$����x��y��o�$"�7�5A��>�<�'�,�X����X�Āz���3��B�#�x��/p�|U�)�p����s���ߝ��O��(���y.�������G�x,O�bO�#o�N��+�HL�w�,��=�X�^��q>;N�Ŏ��^i��d��?js6���_�/��)�a�nVٷ��8��*i�*��M��bjԫUF����0%'zW�Fd����g�<�7{2	\���(=<�;�,�V�{(�Z|/%���&�mc�����𼗳֬+E�랝�!��g7_3�!�5��?3����C����8`χ�\��H��C��q����<L��G��l����C��q���TXp!�a�7a��FbH��C��q�����w$����1�����x������{���o�Ѩ�����݇��ǁ�?��`vû vq����=�@{�|;�@w`����-Qa����BM� �h���s�T|&� ��D�S�Dr.��>��+�ݞ��G�����v~��Q.�Q݉���Qݑ#�GvûCGvH��b�p��4$�բ�`�hƈ^�g�_	��0dg�|�L0gÍ@.E�?d�1��0d`�"��D� �3AfC �>�YX�u��䫰p��fQ.�3S�I�?�FY|&:e�n�,�C�9^���@m�VT�Gt�zm\=��~^��Z�oYW&̰��sFݎ�~�e���tj��v�����'E8RjҔ#�R�Θ��ȧ��1(H
?��Qg+|J��Q^�rH�X�	�� D���Rԝ5pj���K��4�5�'܈UVbl�̉�,���J�A3w�g�w_������>X�r�7Ǫ�� �JFB:�m��K��B4���������G-Y��]+Y!��_�H\��)�`$��vՏ����Q��I���&Qt���dUA��E���[���o��(����k|��*�o'w�B0qV;Şv6�L��L�N*%%FD2tj��L�Nʔ���D/��hA<�	(�D�	�qV�jKK�����$f�7<�B	��!Nc�P	�_�P�gC��J\�D��
p�,}��c���ӳ����7x�ĝ�2�o��z��1���[�����uO6���sKJS(�
��x�<��.۞G�8p��G������Pѿm�������eDƷM�ț�e��@�\���I|��p+�N�2�`�㹣�{���W���K$�/mW	p�{CK=�է���������,u��\�"�'uqm��k��y����զ�;�}�;�ge���R�@֑/�ߺ��~�����
g
�S=ߋe�BSl�eq��>X�>���=l�+��1'�ȸ1���؈a7���G�b~п��T�Ȇ���K�B�*����֒"����H'+����C+����-�t\d||48�^]u@z::��*iۣU���h�2���&1���c取>X�����3�%w8�y2A#ݶQ�H��R���ݳ���1+
��*T�
��=�"��R~�mB��N)��J[ˌЩ(�v�i�
���/�d��f�
_�Z4aM�-Q��Wh���\��EA�þ��r�>��o�!���ZI�������o��q��KS v*�E�����rJ6�nIѴ��%w�c��.�/�do����+䆴��8)s&&$����u8Lr�l�8!����{�>�e���N��]��?����W x�;^7�Y��t0����Λ����
εn�BstE���W$/cù��u/Q��tH�YC�2���b��4�R�u�D7]K?r�G��;s�a�fU����95i�ƈn�g�*V~����[d��,�&�5y�UO�o<��{�H���??���7@�|��8{���̵�P��V��s���פ�ĲVT��I/.	��(ta�����fd�e4�hɩ��)¢�nlP<��$��"���jH�~�p"_��?���i��#�*(�졨M򠃤�N$��Fn���H��R��%.n���-Ϲ�O� )�}ۄ�G��c�� C�:" 4GО�=�{��=� ,!$ 	$H�����ؗ0t�SS��w��R��c�5DJ]\����t^�7W��.������}9�7�;��l��ڑ{k,}+e����n�H��H��g��u��*0�Q�Q%b�C��Q0%�D��q�.�!��m��Vv�*]S�L�YG��ʭʮ��j���������ߟ�y���vXH�?<��矞�§SH�!*�iT�M%Y߉��J��RcbZn��=��� 'T*UE���+�R>>\��) M���3j4J��'��!d��~�Z[�x��9ISW��QU��e
w8�Lbab���dJ->���̵n>���/ci��<k�w���6���Mݾ�6��S3�%o��*����b���b�/��W�_|]��?�wqY�x��!�d��9����}��w�(I�b1�c�E�%��A_|���@��{��򰼃�|_�����o�������w^�=�z�_�|�W���9g��c|M���N_�u���T����I�B�F����B���
w����;8��j8q.��΄�ێ_�?G3-�q�\�ᅍ�s�1���9�Í��$#.���'�wC�<�����|Ê�
�+௃r��R�Ь�e��9�%mqm\4�>������
I8���������i���s���.��6D�+���*
�CMe]MM8�5����!�v�]����	v�2�D�P�@N�@	"�����$9�L��Mߎ[��P��+����q���-��^����3B�2<�?hݿ	�o�>�[�+�r�{�v��O���m���5�9{��A�s���x7����������'2N8�1����Zs4�Oy������"W�+���#��#���J�T��=&H�A�z)S�|�$F�EC��p"(\Yo�;��>�/���4�����_��!z'�)����@�	y��^�r�#\�tk���7q]���1�*��7� ƍǅ���|~$P�P"�̐�F����Wy&�7��ⲿ�(IӪ���C�M�������J�.�)�� ��]��ǻ���!�xE(\,�eeˡ˟������;�3�s�7����UNG-�0e!d\���\�s�w�a]�Q;�%w^�Q��?֚��W�w��}�^^�%��.V}���]��@z �(HA���6�y�Όh���
+����`[夗e������'���2��2��T!�C^PƉ��葔o���PƙuP^-�N@i_�^��P��)�hFk��A��'�mU��9G������3��u�q�N4v��0aa�k������0ѹHe�dK��_��d�r��j���-wto"�.���А��~���t�b�`�ӈ����8#I�eC>�}�w㚿�9Pb޴c�jsc`u�>źq�g��g,G���C�0���|�W�_|�W�_|�W�_|�W�_|�W�_|�W�_|�W�_|�W�_|�W�_|�W�_|�W�_|�W�_|�W�_|�W�_|�W�_|�W�_|�W�_|�W�_|�W�_|�W�_|�W�_|�W�_|�W�_|�TXO�h�ͱt��[�!��`GF��>Qb�������K쯟�W_J���L�
��դ[�
͖� ��@'�Z֧k~t����FA�b�MAw�0�x�}�	
�KγD	Y��A��>:��ϭ�)Tu�b=9����(�)�!���s�>L�v�W�\�`Cn�#g��Әhz��Va�:��;��	�8�[m��MB=(� ϖ�pB��MAo��v�O��է'�G?�i�IH�֌�<d�!�
���� `�u����jP�@��=}DD04>��r"�=ހX����� QB:/�S�<�����fÌp���ٝ/V;��١�zsZÝA�,Q�創���T�J!���#Өv����Ѳ�1����T�ф�\D���5^�T1�	�ߨ�3��l � �_��Zv$.�pLhhtMQn���?��:��6D��ڪD��mk0zBd�&�@.j�ŀc�L�[1��H�0J�~Yv��L6)�-Gz�QHJL��-�iIP6��!�P˾�.�Ǭe^8��&a� (�1�v��m��M��@tP���)�� ���d��0���O�
ya�ﲥ��pp��h|�J�m�;D!�v6:���P�;��zJEP���/,���Xb�c}�e�HJ�����`	�/ G�#�o�2f�p�7���J��Qy�Rμh$��j��s�8*�]�'6�YE�Y�pY�+^��pR�R�]����hvN����6p�J�2�g�4H8��O�
X���"�.�1H�=Q�8�u!/j-��lQgy��|8���1�҇�
����st\�K��&<��0z�l0E ¯+K��r��Qe�d �K���&��	Վ��^?h�?�;	����I�V���٦���~K��@�B8�Ij7q@�8�6.�p(�7H-�ŀ'�<�9D��RRZ�|RVT']��������z��q7ܟ��ݟł�pQ��[�"�8�B��ӠD���<�^��$`@\��ϼ�?�;�U�*$�Ux+4��}$��&�H1�{&��a�k��_��xUGaQ�մ͏�I6�Z"Y]b5�
�K�� L�`/�G�4tJ��
��&0���e�����8���m���x�Ϭ�VxP���B�r��,��Ec r�x��y��<��W~g�i��;6f��!�w��V.�u���=��4wv�R�[G���-�Ei��;e���z8{��b��n�-������l���F X��EkZ��`��O��T�e]�9��eY*�h%4�ǺL������Z:���5�"@��P��n2����S�tD�SU��џ���Ź��l;�?l�[L�uN=yL��]�d� �X���3�nZ�lX��û����8����٭;��r>e
��#�\f�&��.������O��\@��6����'z�~dg���|������,[�=Q����} ���ܡD>=��eW�O� ;�'���,����b��j��&��=�s���&���.X�kyз^��|�OX�_���W����F�\l�4t�F"��Z�� H����6V�\F�\�k�4墛 F �����6����`��t�ƀ4,*�+��j���x��.n ���/(���v��g�{��@�������/�gB��i_�.2��TO�l F�C�:,�'����mK_�r�!�����ذYr��L�%g���x�Z��ZT-R�^�'����%��N���2��X��bkS nv%�/�W������]M�����Gh�T�%��N�G*q\���y�A��\@�r�;�31�K�_�/]��[v�<�-��P��Fty&��M݀�{hY�!~*V~X4ԲA�U��UDb3�Gb�"z���ZU�krrኈr���[���
.�ʑHAj�����D��=l��k��2M����Jlѵ|�����5Y���ř��L:l˒�s)�Om�"�Y��5����	P�
�n�8�ݶ#V�h	s��)�2A�w�1�0���9���d�vp߭�D��C�FHK��`R��[\�xr�+11oNҤ��ٳ��A6}��}����;jF���-`ld��gjk��r���.�?s�9&%e����V���q���6E�gAp�&޿	��m&�dȆh^K�X+ ���C�U�	�ǑK1� �������o?*����8u�P\q�(���/*�6�ZڬK^!� T�[<|�%�d�B�wŁN h��?��m7ᾶ�Aϕf1�nB��l�*��l�?�fuXr�A�����6xɪi�8Q"�ѴpF���m%���͠b��s�D��!��(��5) �7v�k^��=�R����$kY��Ȋm�ܜ�j�Ų��#m�c�c���z2M)aj�� �l�@l���}9xE��X�-;����h��dz�*�Uް1Uڿ�����P:���k�}0M�l䶘�.�,�?�ٖS]���zB�"ÊV��d{^��6���%3���7�U�I@��L:n���B�X�a>*&J�Wh�L��Ku�#��D����)�&挹�6l���q��h<�KJ���/.���x��Ta��� �V��M�./�|���\��瑬ͯmF)�JFK���h����X��"4M4(1\��}*�û-	��s��)P���3�_2c�h��^������L�&���o�풉/��?��s(�	&��o���N\u�e�T�La�$d���� ���d\t����U���8�n�JY��(�͜���ak�6�X%A��v�ʡ
]��m1�&N�t��)0�[����ĜR�{�7R�O��&�P֯�Q�fɒ`�P�rLR���"�MG&��[Fߔ�=e�l�� ���A7k_`k��H���{�n|�r��52dK%O���*�;G ���D��v�����Q���敎��'4�=�ݷ=^��`+�;w�s8:����f��Da�ʵ�څD���UFuG,rb{�.R>�,H
��P.3B��"G3�o��Y�ێ&y�ݚ��e���w$��88��^r��UF4>؟Nc�R�l螓���=�N1��!�����R8�A�/�C\��"ߛKd�3��1;Jb���mT�hGY���|�/K���1�*U�o 4ɸ2e/llP�(�˰5�L�L�wٻa�yԗ�R@�l�A�;J���4��8�����?UٕQ:���EU8d�ɺ3��'d�d�`�Ͷ��o����V�N9}�&�.�^�4��K��(I������O@�������b6+Z�<���0~�m)���/H����ᖀ�Cˠ*��&�8�����Vތ�v�ʥ�V~��b�h�a��Ң�"�b�V��p_jo��3pŠ�Ze�l`��Y>��BP}&��g�r�޼�� �_���`p�h�G_�O��x���mv)J���W�܊����p}���,��w	��y��b�=E�����+jg�ʹ�����`&I;Ft�&r'^`ע%�{1�����2�����d�o-��Y(��H�*���q֔f��XN�(�6:;�:G/&�&_���>'�I�想Z����w+���d���Jd��u�C{R��Zk�m��B�(��4vիAU��f����bF#X�k�f�!�d��$��X;��
�X°Wp�H� 葷X~��3�'�����e5��L�pn�q��?cj��#Gy��m��݀��r
����dU$�ۀ�=4D�+?~Ո@<���,�E�L/[�Zs����57zͰ.�/S���aB:�	�#�����L�/M��h�Y�����"̗1FG�R�]L���Mp�0U8��=[�xñ����!fj��<�������=�ד�i^t���������=iPB�n���)pF��N"
��X���j#xH�V⩐�C�e6HJ&�LF�T ��GM���(��J-��?7���������zt�$��ĕ5�!�D�E
j@�,����O	�����^f��*L�r��(=F:iłx�Rzu�)2���LǮS;��kFf�T}�$��q��3R�g���K�b������dfq�A[=�0d��1���Dr*��Am4ډ��f�0�Ї�I�!�(tq�u4��Թ�+V��r�fMͮ�@�a��q�HOE�$m,l��Ow�p�i�1�R��+S�����K�R� ���pধմ�M|ܕ#�2��Ǐ!,�m�t1��W%�
"JُĐ��?],`�a�Ӱ�F.Q%��0�J�qHb����Ei`u�ck�5�AO����ɮ����OE�5?�-T��35��RY�hR+1闔�i�A�Z����RB�;Yv�h�Jۊ`N�E��7����R�OM�(y(̥�%����M�[X ��jM��-4������ɗ���'��:��0�=�%;�1>9o�`��Q�IUzZD���<-�.n? jAl����� ܞf	"�1�M�4?�3�!|ѓ���&�/�#.ܟ�C�ܕ�j~s��"��� ��c@�L��wQd�E/�&:~S\I��.LwCC�ɤۡ�$�/Z�8��%E���mBY5�v�ǪAKΎ�x�F���ZKI=%�`��V�\�Qc�-�ba�i}��=+�������I�����i�'a?�:���-腩�G������M�&r����s�}�Lo��,�ŭa��t�8��	��On�Y�&F:�ǯu��+�1�$��hs+�������D��B>��o�;>�T|rf!Q��[75�Ѭ	}�����D֡��
+�Z8-��q��XٲkRT�aE���N�����<�%$^��Iy��C��&�)1Qro��91�g�h��4qX�90���wVd�뮿B�A}�3e�!�S`bݎ[��:��lG$zR�ܰ�?��w�����/��4?8w��f��]�
Ӹ��y��I]ft	T�gc��|%�A"v���n{$�=�F*_e�!��V��6V�&G�����!�zb��j����:a�6��G��-u���7�V�k�̰:	��.���Z~,��� IG��ν>|�Ph��v�!�.�/�]$��F���f���G��sv}���Us��af)�|-��{Ȟȭ1f`��nL���	ng~qNrs�и�����O�A>,���q�fH>�,�䪌�=��B���N�y�ZF���P�t�� ��
�r�g BX��Lٰd�g���Y�q53 ��7#��{����D�u+�f2hQ��I�9"hҶ��{e4���E����a���c��2<�#n��X�����G� /�=鬩i�l� ��$��0Bն*�e�#d�O �[��ՓQڕN�ڲّ�����_�|�FξM5Pܭ2d��=��q�\�p�dK6��Jʆ���9Sw�ΣI�@7@a�.#�N����5f�Ü�����Ϋ�����"Ǐ"ߢJ�Z1f� �m7�l��$�U��*��,Y|��9���]�$l�
����Ad���)�	��T���3��U�ph_jŽ�V��w@�b��)V/Q1����_��!₟��P��	n% ��h�^
$�V	��5�-ɤ{��t{	t������z{��l	�D��	�LV�P��l#=�LW3��'�a��T�Z� ������"a�U*�&g���C�Q�|��7��B�4��SI@Q�rrw��i��� �<���)��K,�~��|W3Qv�&+��7�].6�gG�$ĺj��1<�Fq��èU��Oq\�AH�I�A�%����/��B��Ĥ��vg�O>���0�.������x��\"wD�_l�c��B �����Ĺ�LU*�)���l��c�l��O�=�t�~1���*���]A�B�:��L��Wy��Q>M�)�$%��ڂC2zZzEo�[KwVkB]��嚈�F޷6�a8�7p�R��'S����jX������Z���/��m���/�عE�s����T�h�,�I��/�0W��j�ı<��� ��u��ڙ��#8_�h���5Z(�Ajx������?RB�B����d��9�^
�dO�/��];rj�E�>���|���%��U/��;��C-c���-���'�W��ܘ�m`cv2A�`���Ax�0�F�� m���e�k��cn�)X��v;�Yg��E��1�Z&�o�')N¬��p�YI�cS��z�����S��O��;��K@�+]�t?Őfb�S̓��7��OcA�b���/���,
u��H46o���3�k�~w*ք�ze������wXn�q���N!*��QSٯ8D���WG[�v(6���Z�}CM��� ��>���]�?�c:lg��u�/�x�2鋪��dAlG�^^�rH--w�J漉�&נ\y֥�ӤsD��R��{�I^�9�,5[�G���w7{<c���`��>����s��ԈR�o��\��Q>ǻ���C���W0�9���v}�z���ٮl(����̀98�0��93���&�4��a�]��)��G�V���\�F3����.K�6�bu�\�{ڎ�Of�����B��[��s^�o��^oL��=����vS�����nPT��]�S֟x��֙�ݮ�����[Ӈ5�|���u�.hQ;��+r�l�ʱ��
M]�����w���*[�K��n����6%&�w�Η�N�7����Mהּ�����_e�9�t�g�\O!�Tb_l�����;��[���_���\�<wZ��R����}�邺wT�[�K�nӭK@Y�3���\z
�?���>���|�}���\o8NG�W�����|��*�.�	��E��,�J�=_jNJGJOf���Iz����S�Z��j���j���g��%�R=j�	�����W��}#��˅�j��(��,"��D\d�|�%q��R��I�=5���	5nI�����ޏXs�k�nu/����;b�.��Jcd��}7`���s	��t`ꁷEzD� ����k\f���b�I��O�}v�G��́���hM9+u�A/^���N7�
��'W����\��\$��ګүk�7�-�G\�nFo��J�+K?-l��]��˞�Qo7%m����&���l����.\��U�5)
q ��3��bY�)ݔ��׾��b`�J�6���x�^�f����p�������E��BK�:)����h�NXk7(�n�W�������K����{mOw���D[o�b~y�o$7.RQq�����M`���٪qͰ����ʰ��,��T-b�<jX�oruG���i���L��q����
O������ޏ ��O3|�s\�z�/��R����t�'�i�ȁ� �1q܆.̢�یa�tb7�%ݏrG�S��*L���ł�B�#��Vj�I�8pw�����8�{���P��(�n�l]�6m�j�~(X���T
"^ݼ՚�2(�5���ld��0/���+�B��ݪ���g�p�͇��<����5���:'�~%-�u7�\�O�������ꕦݽݭg�O��/X���<j�y���S׻z��4�%�c������k�*���w/EP�Q\����;��(���5{���S+{���Y{U�N'�i�M�|�M�n�vfd\�%�4�/�Ү����-}��r�W N2#t)�5���Tu�Kxkk�o5�q�š��<���6[�X�5э���0\/���p79�3��(���um��\�w���r���^��F�_�Pu��}��ao�f�������Sl���Bj鷾Nv�G�:7
g3���~��8��NiT��>�7�|wF�ք���!���؄X��>��;�Y�b�m��c ���|� R������mu��y� ����{;�z3��|��p²`o۶�$��f���'�\�ڰw5�;�\��Ω���@]Geré�V{[�wY�9�	x}��	;Km�b_��%��&?�T?{�c�B�y헪�;.o�)]��&�r�ow�$��_�`wd7�˔f~�������5&@�6&�=��mby����Ų'M���LK�}(��(<܃�Z� _猄�_�GB�OM_^s�T&��Ř���ӯ_���q��=����H�����,�My��H+\+-�Mνxe��k��Ӹn�|��o�z�v.=e�Xg�|C���y����`����N�y����&v
L¡+�2�`j�m��ms�a���+�)X�����jQ]:����)|�c����޷���C<2�"" +�� A���:�T⊀��NN�8������� Ѝ*�P8p�(+�;R]R�(���]Zj�����[Z��*fm�����w�B�~�od�˽ս˚U^L®��
���Y�e�˻�UM��v���\*�������́W7`�ɱn��*�>���ٹ6^n�;������}��ϟ�=�����'�{��O�|��y��x����xY�n�4A�1ms�(�E�����kn��,a�);GThOo�zx
�_���"U|p�90+�z�n-��g;��&�C߽G�B�?�gqG����Iq�S�x���aJ_x7;��c��&@ӂWJ�+�ʱ�*��>����y��d=,s�^�F�ɜf��x�W�	��]y�}6߂��7X�4�����.>Z[�]�|*���G�����-���t��e�_:Ǟψi�����Ol	H���}ڮ�^��$߁1=�A�u����z��f�R7�Of���y
�*�����o)C��ފ�����υ��{�i9������g(�PU��՝��0!%�hG�z�(����#6u��uZ��N��6�i<��$��~���q]���#�2�p����uFxN��(i��Osr��,P[�߂|�6(����]
����5� ȗ��F�����.@���Z��5�-��S�b��,>E�/�C��v�4\
f�f��OJ��1`f����K��/Juh��=j]�Za�;Ҟ�
e�Z=�(\EV�V�k��$�J��RD����]�N�<Cl���F�ל��9�;Ϙ�0>�!3�*���?T���\�������.�xhr�o�\�w��##yrg��qaM<ԫ6O�ĥ#@���_��:Sfl�F���Ĳ��|�JƂ���V{h��A
�Αح�d}Ke��@jš�}3b4XdK4�d��Rb�Eo,%���hE�c��<�z����Ř� AMQ�g�OUt}�6��}�y5�z���h���g�0'%tO��z0S����lI�Ž��ʼ�9!��vaB_�P��:L�܃	\fZ�K�"���P����\��9e��wxl!�)���|:.%��j�p֝A¼U"I;�pzr����CN'�����tL����/Z����d+��z���y�ʒ	���)=뾠]O�Y\z�Cr6֕NΔ�C�~zk�g̻�;�|FKP|iy3���@~�v��,Sv� ᳩ��{��WD������S?u�탐Tg&�+���K6��Q�W�J���Y��2�kc� ǔ�'��,��b�N���4ԝ*k('��������#XK��F�J `�櫔G�mU�<9�Z�/?�J�7�������\�� ��y��@dP���X�Od�ɽ�*FV��)h?��z�����!]�J�gw����E��i��Л�����ҫ���a��=c�U���i �u��Bƀ�.��4]{��#�ݑ|:�#��X��wȩ�����NZl�o�G�|d̀��Z��=�����D�l7v�PF�S�1��p!�@��R=�}%EW�C ;�А,*����n�ܩq�N7(ֲA��֯��ռ�f�\݋����$�zjɎ�u��� �� �����c�1	 �/�{P=�[���
e�K���Pף潥��A7n���O���!H!^ 7Ä�|�
ի�CsȴB�	����{ݵKa
�������f��-�t(���Pm�pi�3�*9ع
�Aϕ�h�S��t��VAT�NQ��V��I;�0���=�94�G�Þ%�i��t%�D�KY�Y�e��6�R3��[Ґe�����
;s9�>����0)H��.���T��Äbg37�ˣ:�[�]�B�w��4w�^�+Z*1��-��Ji����(���S�'��^�����*�{��cߜ���"�*��iF�C�:D�Xm�4���7:_⥦��P.)Pc^�����΁���$v&:u�	t�������-�?tw�P䘜�4����Ǔ��+��N��$l��4��b}�M�Ɗ@1�,�,�*�$�h��V�xam��V�v�B���V#�G��-�Ho����~�^0�������ڲ�)�J�n|���>�K0G��P͋K@lz���DS���C��.n��������\���@3'���l�hYKw�S��晖z�C�Hz���Q�oE{��L`�B�?c�9�����b},`��� �<���^]��e�,�>��`1UgH�j�����D�?:l�١�)2�" A����2zK����Q	1$6�a[^�8}�6K���LEZqo �F'1�	�yz+�c�w_��������Y�dk������;�{���$9�-	 �.WI�Aْ��Aw�n2��r6� �!D�5�� ��hD��R��$ã������/��X܎9*ݵ[j��&Z����	��ż}N��D]�=�Q�}}(����Z� �UXA���gT`��]x_�%�T�U�	ϖB�I�'Q��^�D��5[gU��ҏ-B��7:��㪶�t. E��VG�dR^[�(м8�c�@9X2s�Ig��H�@k���G�szH�:%Ӌ��F�¸+�e�l�P��Z��O��~^������1�`ڴ�C�+�R�dGeWk���ۈ�x�hq�d	(9ǣ�1 u��&W*�학m�������d]�X��z{Z�|ᒘ\�}���è��Y��=��b��>��O�8OZo��Ty�����~φ���>𵁽է��w��*p�����i( [�0�<#����F{x*�G�IApJa�	CpXU��I�5�R4���Oe%R�o�~D��3ia�C�g,o��3��{��V����/����>�f��G�f�5�r��n\�>Zw-W����.�g�AyQ�ܨ��)�[�j��X/�h����fy}�/[ˡ��)�0����������5�+%��:#Y�(����'�_\��uQ�c)�����M�Hr�=�Zxݽ@VޢcOƀ�\����4����JE�t�p�h�A��6�c����G8	m��iڦ$x�U��[
�������>p*k�^2%��j_e�^��?Q�l�b� l_����o!!!�p�g��n�+��D�]�'�X��E��:*�c{ϗ�?`�w�*[w����ר�e��%9���EU���9�7/���|!��ݰ�x��d�\dzQ@w�j�H���8���m�_�(����OL����p���8�����{������l�ȸk��V�~xE�l�;<��fno1{7��Y�ag�+���IH����c�����cDQ2M�z(��z���@��)��ޓ���Ws�^�����]ʌaM���P�նPN7�w%��?MD�!�L���5�.���Z��]'0�J�
�etiT��H�UkΤ��-��Ve��Q;��˷x��B�>�W�\v��D��$i�˴��B�eUT�;G`!�%�o��(��H�֩�~ˮ�H�ݏJpR�(1^4�-;�n��.�l�ːs	)P�c�;t����eT��6�~?���u��o���M����N�>�[�ב�����&�:3P|�CL�;��2X�m�R���Kh�1��Q�O�����]�üdN�I��.��]��9�u�I��뻯%g<�*�6�\���>�yP��$9_.����-R���Yi�1�*�7I���~������z��bݐ�a�˵�{a�9��s������'.�w��v|-﷍�uzK���O��a�4���������W����+��\�[����tY�޿xN�H�'�� 2��/�;���\f���huy4�8��%4�������Yk2ܐ���/P��s�>�b��2���1�7�_�X�!�ב�E6<%��~���o�}��
�g6�P�b]�\*T��<��n��d�<]E�w����l��<�����o��r'��>?Q����h6�^POԹ����q��|����ϙ俶�M��o�+������D	:�s�.���ۑ�	��(�kߓ��+�#����u�%"����Cߑ�Ze����n`ݟ�6*}���_<�"�igf��K�Y}���薟m��� N�B/Jp�KL��^�U�|1WH��?��6[x߄�{H��8�o�~���Wq�S3����C�B���-bA������V9��V?�<���j:h+��� ��Dt��T/�C�K4(��p�n)���	���N� ~'_����)d���,��Qx��ʂ���u��'}�c����/���o``�˭Xgp�M��둅֭��!:�ٌ�1�-�b:h��T��{��k�y��ې��j���;VԾ�����T��r�ȭ��OA7��CH��f]��/�.:��|n�=�.4�B^�j&	o��T��Y'�x�,{��B�1 m�k9�\�q(�����;��]����&����W��������W962�(9�P��u�G�w����5�;��[7������B�iz)�����ʋ�jE�JW�!Û`�P����|D�V�RP�2�Й!�{��#�G��=��kA��׸�3]B)��a��	o�f���$��!��#��p+��cAH��+CH���>�$��*��W��p�[�qӓz�Q�H�F���N�@LU�b�h@L��?�0����+�v7H�,��f����}"h|&d���ϗ�0 ��ߐ�1���H�O�<�Y��7�M�mA8�*�w��g�;�yv�C�[��[�OM��<�BSָއ��f�?N����;�G�PӐT��Z���<Zw�b�zsƧtw�n<i�)�(֞]��!SBS�?��V)�ħT�Jo��i�a�\|��]^�Ϟ�������s��?8e��,�APX�S3�k�W�t��.`Q�V�;�Ua�K�?�U
�T����F����`��A�ɖ�S��~���
zΧN�B˻����R��^"������c������PE>�t���r�t��}�/
�1D��C[�����3��J�]=�X��ԫ��;�uIJ�_�!�1����&R��^q+��u�4��E>�+�T�v�=�^��£�bc���������h��Es(.Yv��wʟX�����G���'ůW6�l��������$a^DV/�˙ߘ�y'���{��@pm�5��=q�Wۓ�� ����2��(�&
m�.��t�]�d��K"�nj<���6��f����"MB�b�S�4�#>C��	�{Ggt�ω�6}ۧ��9�2R.��nǦ��*�_�&S�]:aD9��+Q������N7/rK�H9�2��2,i�Ly�D���j�~���<$�~�h_&��2r�ra��.���������l2愱 Uy3�ש%I�9r�f�ly���:nS�2��]���_�����5@��S5��Xcgfe�#�[(���p��
�X.v�q}$i�3�c���/��s(�x�������x>�Q3�G��,�������1�k@��������@�z��>t?l��V��z���J�[U�5�$w��/LG"u^א�Gq����>�s�������xf�T[ z��׍�z�H��}�x�=�ۊ$�^ȿ�f4��N�ཽf�7;މ�4U��lߟ��;M�z��;-�9V��P��^D�`���z/�����9��Uˑ��_�M;�W3}�'��#0\}�Ќ_i���j��It���g�v�`�G([���8[�}��ĥERd�۩7F�\���}g �A��)�1n��l��Ƀ�U����T�:�cT5��5�J{�̓��W�K��;���������b����o��p�&j�KkKC�g����� F/>H��j�g�Oڷda���A��_�:љ����<���?;���}�;�m`vň���w�Q���X+f�5G�P�C�!��m��Z�9 0t�h�N�?�W%�W86��d�x���^��a��G�� e8ٯuq<�+��Ӌ��a�A B���������ʁ��h��;ϣa\c?�t�A�ITٚ�/�P�:&����$m9#�.��I����Q�^��{;x�GM�+�b��s�؝Xv�ӥq�v*��$c�.�J�C.��l>�� )m|{Q��W�Wo����{:��3����$��i�$M6ocL�t]�5Z�������:�Ӣa]!�.eʩW_��
�����������^�(�BN�e�\��\�����C�������cW0D��V��`Fh��kq�;jL�V?��J���f��(��3o����W���Zx�(�,'�Le��W��ٿ�.#˸U�Fk�}� ����zO��[���i�����f&Qk��J�_��}�\!}�,��W�T��55��$+F���AqT��Iޅ�ԕ�p>ȯ�eO����2&J�.+��nu="a�Qs�H���2w7wL��_��л꨷s��O\͚*>�Y#������#�o�Z�ј�ڇՄ�2�/� ���/?���.^�W<K𯱥��_�|�>���������ɽ�P5Ԕ�z~�(��qB 	`%�i�D�U���c "��:����|��_�,��0� `�V*M���m�u �\b��*�S�?ҎEO$~?c�\���� '�3��*� u>eN���?ʠ�|��������X��n �ҧ��΁���7�@�Q���G�R�N=�o+]%+�c���P�=K�U9��C��`�:��|%O���S�s��Ȝ�!�|��6 o���N��΍�H�揀.?N=� M�+�=�~|����
��J6�2\�>�s�2�yQ�T�y膖�(���V�y�ƎZ���P`�IQŪC�suz�X�-;$�ht3��%��{��-�fVA4.�Hd��N��^P4O������z:ۖ���H� �k%u�hG��0'�s�`�a~�'�iJ�hl'��a��GÄڜ�D�G ���P�I�Em�>Z%���t��NY��8@9��ET��%�J;�|@�Q�n�u������	�M�H?��(�u�Ee:�h؏�{Y0Fq:�㽶��Z(�&.X_�8dD	�)�o�$ڸ�ZJ����Q��'_ӽ,b��Rs9����h�~�,���]��=<ތP��>8��Ԓ�J��ƣ�P��� Q8T�(��4�o>�+�>@��f�s���<�`���	�jk�P H�r�q��Z�V��	�_,,��w�hk�8���k�'䗢t�]^��ҏ�V�����	�H��j���b�Ga��z-�����$��w%���׷�G���#�%���$:�JKu�Y��GaP��q��_V�GtD���[��Q����L��U���:��!�H�d�Ѡ#э�+��g��{/Y*%����btwд؏���:.�q����֣��ޭDG�H��Q�a��[���^/�rRz����9h����Q��6 ��8�_`���a5 �
"W��Q��I�[�8C�Vy ����	T�Z�gT{6����{����qq�c�ܪ�8���[���JZZ*��z���T�~����c��R��r,��ђ��#����g|��>��|R��RX=ֈ� � Be�dkP2�!�@�_B��ˀȩ�{��2�be����y�ӭd���UV�0dq��#�bF8�FE�~�/;�8�a��&�ӎ�L
�r����������
$DF��iS�_�����;�d�قd��ݝ�4��4�ы�b|h6����	�f��<19�j&��q�يC�kH�ʶ�gM^���ьh�a��I�ɢ�!6��U�|J7��:�za���k	��#���[7��\��Z�%�fx�g�|X��yE�3�2e���������6�V��6�cĶ;�3�]
Ϛ��+f�X���iɻ(c�m[d��Z{��|C�x�~n��F�����R-`5Fc��輯�/�\�[�Y[�e)��h�1Ѻ�7�ĖZiӭa&�����4���3+RF�c����b⦦��W�|j�&�v%�l�����f�%��\e�M��D��]�j�-�c1��E�lōw��b�,��ne�-rk%�l��B�^�7�z c�|%� b0
۪d9-��e�F�A�	XYK6�T�yPx�۫z�HC�}��
�D��7lhs�Z�Q��`o6IlW�� ^b�<Vch��x���8,(.�h[_�&�sW�2�*󱡫Z��c�}*Ϙ��4�k�U{s*+ZmP"3�	z^���2���Ha�L��&ُW$���ͮM�3Wfu��ƼF_N�1��k�g͇�k�˺7l-6�& ��y��P6h��Z6�#D:�����g��f9b�E-m%͍Q+w����+��,���F��{�cNE^\2厍q�r�Vn;����Y�k�,i�1�5"���/�<b�,f�ch+R[��Y\Ɍ��fS��%�����ϓ	�fn\2H��1�pJ��.o���-���Tm5-��m���2�͋�bo.�m���j��%���ύ��� ����m��'��K�s�?�$�*[�b�y���9���(�L�i����_��b������G�_����'���	�˘����P�����T݇����"W].K&$��&��n|ٲ�7�c5��~���\ULC��-��4�w5$�U+��B��'�~pu��G�'`�Cbe���1GG�tʉ�D���8d��b^�8�E(6���6;�g��(�v�[�%�S�Y㦷��pL�	(M_����S�����{=]p���ɸ�9�f�nj_?ӟ(tho�]��p����I��PO�G4�gA9��"�R�t��25���\G6V�U�%
�7�E�@�u���y�V�w@���M�nq秵�trp���U�Ѯ�s���i�C� ��2���f�u����哨9Z��}FCU
�zϱ�ness�՛zM�ÞŲ�	e����~�yV�X�?H�d���xH��̯�l�!}w[��X>��VaN]0�VU��=����{��-�3�k��mmަ�|A���ԫ#�!M�kHt�\�Zc477&,)V��\�����5ɟ�C�	enpj��I9��K3��'Bzt]�E}���M���,9X<��՜�Խm�����o�:����Pnet[M�ֱ6�&���2�������f��X�8v�&�R	:�զ�7{�3E�����Պ-��R'��V&^*���b���W'QY̬��K�s�Sվ��
�����v�c�$���z�E�>1C,z������SZ�����J �U�B��(К��g�����=Ʒ{ }UT��,��˪;�H��6�զ�?k�.U�g)����9��j��:�=�Z]h�K���[�&�+��.��˦��:�V��mS��e�sf���\�=���Z��ޚ�D�R����x?���j�G��{�A���k�K��mi��:_���*���])�W{VuVW6���sl�n=�Ѓ��V�����{E;4�F�KBY��#u{��?�C��Nete��p�k5��V=٤�U�HA���Y�l�����L�5&n� �,���:�'89���I��&�[�fXUY?������KR�C�C���i���T�Teԡe��7�7�⊪������N��VW-��Q�3U}t���W�ϒ��̼:�e���Ak��P*�U�/j+�l��G�R��ei���UIU<_�X'G��yy�\Y\�=�o�y���M� ٕ�Y�ح��m��� ��LvY�z	���H�@�Ȳ-`lE���H�Kp�I*+l�d����E�$P��u�z�2q8�:��$^5����$�')�\D�Y��N�d����'_u�%�0\,=Dfz�Q����&k��xN�����ֵ�zw���]|{��k_���I,��O�㟏���w"������W��b�x��������[�8e�$�O��O��G�_�­ML��u���C�v﷾��s��� V�V2�se�|���8*C}Fev|\u�b�������_�Xϲ;���z�l�z��W6����j���/����,yr��*�{����ǔ�v2؜+����������ܙ�&���`<������b�˒s�o���g$}���ض{O�ᛸT���z���r�z���Z����+��;�䗚1�gw����-�#�մL�B� +wV�6ŻC٦|s��=�����|���Mk�^�B��7y���2��p���V�����������?�i����*�x/�;����̞��L%���h?�KWw��pc˧�-���o�s�7#�G�O,O�n�&��hn�����ڕ��Y>خ�C��<����V��Ŀ�����I��=��]�������}l~^eU���Yp�{i�����~��k������A���A����?������˿3*�Vk�@��YI�-gL ����s9��'�_��� d<�pZ��yZw}�j��
�"D�������oʛ��mW֎试4������Y+�Y@̫�i�
�h��/5x ��y9-��h�ZH7�����	�hn��o�+�����n �f%�tj����]Qo�맽�!���槙��Ƶ^�kP���9�l��|_`+U����R�3���W�6/D^bIb�F�Lz�L�����:���[����9�{�\-]u x�k����@ρ �!��`�5@H"8 / �`#y$���e�ZT�u���f@�w8��*g׼f|�y�X ��7Ə�� �gx���'ⰰ�l;��U�d�N�����it��󿱘���s2��p���
;3�N�f�(�w��]˒?</pfe�f�����.��´�q���卨�[�4�ۅQ����
��yݨC�;*���&fi��	s�����S{n��X���K-䜥q��nq�]y�}�N���b�f��_���������2 *�؟zq�׀��%�ִl�әg�r�?��|�5\2���sP �M������,��^���-Z�*��E�E�k���LV�~��݊��o]s������G�ef0��?-��YT�D��ݢ�ucd��k��zE�,3e �K�֞D��O�� _�+��~R�������d�R&�هR`��OL�G�T�U�bjUN.#i����a�w{4�{~ېǠmH���֋��d��a�]��G�D=y|����r��D�B4�!��Z��Я�L$������v
���k�&�S>�
Va\�����y�/�m�r����hl���D3*��9�
Sp�;�DVv����
�*�I�"��R�i���ß;P��Z�S��*�\ޕ).�d�����G<�_��o�,z!��&NX�;�L�F���(lf�nCQ��'�mB��<�sk�Y��c�@�f.�Y��^�"h�QbrJ�F{�V$�y/�h��5��I���-�7�h�8~����I��X�����R�����s���7'q9	�y�3�T�l������Z��bnJb!��e�����OM�x�%�~�dv�� ��L/@�z}���tx�{��\t�k�S�va�=s��-�[������pA��
�8>y6BG�����鳫��j�PF�}���~	����a��tMw�®���+�:6/{ �K�e�:�Q̀�޼	!n;��N<Ոcy�/u�պ�R���1w�P��6=����`��F'��^�I9�X�c�nr.�,�ľ�����>(cw"���5A��eQ_ދ�B=��Fb�|m��dM6�e���ߕ�����Ӽ�n[\����:В-iq2�X��3�KH�cG� g�r�>s֧Q�-�o�Yʩ��wh΢��������}�3A���`1�
��O9Ph�9�][����HB��cxyy�&���Ikb�A��Ŵ�<�Ea�k�ڊ�p�&QA��b�2��8������3��>1z$�{
Z�&��9��aL��c�U�#@n���YC��7�Y�[E���10�pĐ$NRם���a=�.j��A�B��LY�E�PBדd�8�|����֛	5�2}�gs�]��I����}Q��2�jZ�4����M(�7h�-�ߓ�%�~FG��H�h?ߪ����Y�?W�o���il�S�ǔH]��մ(�bD��O�$���r�S���q�C��c}��J�n>!n�Ը	���J�ao��6�.5����bc�D'0��8��y�?UG�}� �~(�7>/�p��G�h��"���e��P)�y������Y��ș��]�j�uؔ��nAP
S
�]a]��#x	37ؚ;q�Ѭ1��n�$��*ׄ~sg�% �:P������wm�6�^���N-�~��UZ��}���jE���*D����T���o�D]Jx��T�o[��+�G�6��)��"J��s�O�;'͉��B�5Q���h�%�e��oV���]�=.��ڎ1B���!e"珣o�Pd��X�����;jτ�W���LД�-�Td��4�Gp�3"�r سfx��ؒ��PW�؜�j��җ@�U�]��'��6��(�4��{�16�V�m�aP��QR�YL��d�^ ���L����/S9	��F���0����bw��u�����Nɷ�X��6��E�v��)�̊:^�ѿ��r�ul�U�tM�:�<a����iJ�%~G�w�ch��7�,��E��Vvd)0�7����{�{+�ϣ7ѳnl".x�&�ҟ���^�	��w_�`"��'@�o�`G�~�{ �$��bE.b�'�D�lz�]/޸y�fw�p���p�����! ,~�r����FImBTfC�ZOt�e[���"im��e���jsi�l/��F��~h���
�_0��Y�j!�d���5#��4O���-2\����t�7��靤�]�uOŬZ��;�i�)�vY�xٿ>��J۷?�.Է�JN�*uO�u����M�T���M&�7�1�Ȕb��q"�)^�Ї�S��
b��n��v���5k��¬z_�Zқ"(г��2K�
�	#��O���'w9|�A(N��?W�@�8�=|3�Q��d���<�%s�|B�6�'ix?�SS�aL�%,���ilx���=F�:�,/�L�����4i;?1�~]�u4g�P�fT�+�]ndM��L=Oe����o�R�ϐ?]cZ�2��VQ��t��ph"�j���6�r���Ao-�Z<�T������L����l�2�	P��57�?��v-�/?l��Og�&Ԯڤ}��'�L�]=�����Dosd�$���d����w����;�$frQC[�/9��R�zj�'eT�GM�UE��r)��wQ�ۢ�z�I��#v��a،R��ّ1�c.|~X�&��Ԕ$�5�//:� `o�]6��^THw�����J�f��Wi�p�t�I���إ����Z7�j!/S>gށ�fO?��g����9B��ʜ����9�*L�V�°6�~˝^E&#�Vf���<k���b�%��t�(��,l�c�NS"8�^��� ��GH������ �I�`1�n���c��{�F0�D=إ���IB�i�=N�B�gR��K��3�2È�gש�C�d-�����_ݫZ��#��[�DX�Sz�_�r4`z��(P�宅X�5��Ӿ���B���&�˓U�=�VFS�K�.�9Q�[��ĎiDȤ��gPΔ�c�\ۢ.��H|;�������$!+K{�g����S ���;��6��O��M�
{��O�)s�b�F����.~B���K7�0�o�8K���F�������{�lq`魘!���<]��Í�a��P���#�E�,�'COs�Ϫ,��Pl�6D��)����)�ν^����R���lIMm��ah-�m�o��KHy/�4���/0��몾ʶGI��ˉtS篾�4�\�ڤ<.HA�L��$��K�<ͯ�
V7�X�����o,�pr���T��볇wp'�GL]�����!�^�_��B�㘉�-�M��+�߶p�!3AA���XE+��M{�W{�s2
3~�U�{ ��Z�]
�ΔbnN����^��鐲}�e�N��2q�;�<�J:]P��[����`�Z��|k����G�;PtJ�K�
���>" ��ostF������hӟ|WԺ�����;�d�l'�X ��,,�=��!Wr�~�j�%�t׌0u_rVTg�ecQ����OPiR�t�	F��1�7QK}x���A����fA�ۯ��@x�d���gȨ�Z"]	a�:ߥ��v�_���	�⸌km�C"�	0�F�����$��l�q]�@����A���S�w��~'r�uOK%�w	���L$�o:�'���͈ÆR'I�,�4̽��MI6C"g�����#}2%��7�J���;���ö^�S4��v4�v��FP��z��ztr,u8�XP씸��?��Clv�Om�JC�;����2PT+��w/!yD���6����j.��݋h����y��>-ì�Jˋ4�Z���Vw�������qѷ>J��uk���{(��?8e�������%(��_�9}�k<��a�� ��m�}L��da��K� ���(���P���$�7qttm�����s�Vy�%��#;�M�R�~�gZR<��BB<��uk	ߞ3=�.x(X|�K�W�5�!z�_Ds኏�t|�ç?=M�˝��xn}]�+���`',��}UM=��Cj΅�0�^�X�O8�E#(Тͷ_;r	���x.E��!�y?����M������`���
�8����Gؠ�>썪D�$]#����0�m�j���4�S��:�(U
ͤ6M[AŜwy�r��Kv�8.�G�����RƙsZ13�����2j��G�w�N+tiiI����5��V{l���yU�B( �s�Mc��R�EM�.t�%���B��e���S��=\IyU�>5��$��f�"�<p�"X�5%���Lf�7��`6�h�Kދĸ]"�J��3$�y��{�&D܄�.���N��נ�1�,����O(����g�S��I��E�JS���%L���cT��9�2O��r� ��Ұl���1Ṯ�~LQ�B�I1��X͜@��^A4�6<�nPbO;�a`UH��t�ٺk�:y���4��wE2e͔��m��<���ˡnd�pc��	���ۤ�-aưә��/���;T"�Ч���.I�:���'�38*���������v.�G��!տ���6�����~��Aa�t�'���a$J"�5b��������K���Y�� �lI�ax��G��{����
�/���E}qNvfA�����G؋o��ݐ�(���P�䬕~k��ع67��Q���7c�5��v���%�ξkR:��8�lrQS�v�����/��	�Z}�C��.���!	j"f/X�OuD����9H&�4�z�s5�B	#
�u�5g�Y��̮�G��A���Q�Tv���Rfm:M�cy�R2�Nʙ�`�c�ė˲���J~?�WH�e��T�&���k�Z~�m��%��k- ��4���e�k��>9N�ѕ���+74A�F�=n���d%sjU]��-{�ĩzk.��̘Ʊ ��V?ҲN�/ѽ�6�=��c\�g)�?Pd��k��<��_��(9O�a"��?%~#��Q���\J��=���95Naco��X�E��aud1�+A�*��Z<��O���ZD��P~r4*�����f�ľ�԰���{4�o�ʉ5�;R�.B�i�Y�j�pd�6�\ZXPS�����Ǖc�g�h�=S�T���A��2���~�w�y:8�����
�(�HvՇ�ɺm3ӑ����30��j
���JK��CU5,��o�Z#���x�S���`�I���,+��z�P{GWbc�[a:ì���d�:lR3�o��-*c� ��j�p�n�������Vb��Y�q/{y�}ʕdY/U��HVv�+$3��;�g�6Qga�;nF�z3�ɣ��2�)Χ!H���z~�#s�
4�1{�f�ݡW�JH�rE{[���1��5�m����;8=��<Խ��hN��z<�1;.�ņU$��A��x]�`���z�����@=�W}��új��
q��}�����0k��h�k/�5@f�9~p?�l������et���x�@�cq(� �����2�(����d��y�R�{3qG�{�#B샦}j�ؒ�8�*�H�õ1��bO��g�8��Sr3�Ly��	�/��>�7K�Sכ[��}?GXWd��ף�v��'�a�.M�^2��"X�٤�0.�F���KXw %ףW!&h�ӝg�PU��}�t��O�� ����Ln�gC)�(İB���� ��}����� e���4do=�.�q��k��7U�6���Uaꕪ�or�7Ƭ&ʥK�u[V��&׺8�q�O��,��d_X�[�K'����Q0V�x����Qh��A	.B�~|Gr5�Щ�X�m�镱���G-��ДPI9��f	_S �jak$Tѕr7���&�[�0���_�C�S�e:�}︶]�3��ْ���t�U"[�g��+���
5�ׂ�b�u!�ŉ5�r���Ckt����D�ێ�/X���D�!|�4��E�&��r�A�@ADF{@�#�ɼ�*I4R*��
}J���FOي`(��re����#ٝJR��OD�$�\�~���dB���L�=�*��:j�|�M�$����]*��Кn=��!��>�5�]:D_�oI�e{@F�M��5{������'�=3����g�r�lh�q8%��(��y)I����G��S�4������K�����n#m��)�ݔ�<rxժ%�l��Wl��j�)Nh�ol��n���J���w�����TT��d���`����z�s���D(����4��,$B�@�;*��:&)�;մ�s2���6cC-y��$��S'�b�	I�A�ҼU:1Ml,���
��[X���_a�c�e##Sq����m"B�PϴCB?xr��	���@	ӂ�F��$���ժ}��`��4M��� YY�Q��i�`Ji�=~� ������Г[l}S��d����]�-��e�7/-����h1�#��`�\�e#�mZ��]`ԁ���c�jb�T00��'_锞�C�rwk]�d��؝tH�I�wE�-�hTQ�D�t�іRv��<��s�k�.�l+��;]9�{������!mg#�@p���vn�)t��� �]�"r�1B���G�P�I[�vt�����פI	<�i������5d��Q�Ⲍ2�~3%����")W��ADeIy�Hɨ?�ފھ�?!(�����l̄k4J>��S���[�u�v�(�\EN�JXf1�p�.%�BE�[a=��� 7���27�vDh��$L-���O9�q�KcPE��'ĄB���Ս��������#��~9@J n��E14a��Rg����ܗ��������8-¿\�u@�h��I��3������5��Ǆ�b�T�+6/r<.��!��F*��4��"a����0Z�zGo��#�S�\�n�$��[Xȹ��2p6*G�6�fR��<��a��n������_K�%z���m�M�X0%c��"ܶ����Rr��i���,V�):0���h
�Ip�"I72k:mo�"Fd�C5t�����bK_�*�JRQR5�	a�҉���9���G�;f�6 2[��P1���:�wm$6-`v��_6x�5|�}tJr��-�I[�1��[��l�2�)C����JR�'��/��m�H|_e�:�����G�ˁ2q���Qő�U���^Pkz@3uړL�kE�Y'�Lڭ�NM}��/�'q�eN�TWQ%۰(0�%�R2n�?��N���$)�ȕ�nd�\ȟ%��Y�V�@̬�]u�z��dO|��T�&�VbY�,�PK7����B����D"�t�������p�%���0���{c�Y�7�+�/�}/���{d���;�͑!;[�|������g�,��~��+걛�S��w�h��S4����\0���?B,�	y�ޜ�ւ��!S����J׋��b᪭W�6�9����:s5�Re�kzZd���?��x�����m���MM�7kip2���K��r�G�
���X*�f8R:�.�w6[�!X:H�Ea-2�������T�D�l	��d����ŝ���%bz�+���A*�5oZZ�E^I����V�l��@qtp*��jIhRUq�5zʹ4��h�
 �X�F*Z���)�zPK	-�X�
^bb��K�,��I�78w��� p�p7 o ����܁8 �ف< @;	 8�	@& �8�v@�x ���l�h�� 2`e d"� P������Z�}Z��ZY�Za*�`&@�l	�'��<Xp�;�;�7 |�;�7�� `p0'��Hb z(��c�	p 1 ���i�@1�; ���A��@@B �uzQmmni�xT�`�j�}0`% �ځ�o{
����и�Юa���*�
��7�,��+t,.x`�l��"y뀝����e��K{[�.51��B�L8����&f��^�E:D`7�j9��U�'/�tj��?K�[}�S9���vN�R_�l݋���A6�X|�������N__��=u���u/}��)��JH~9ا�~��pBD�ۻ�c:Ƽ��9�F�s]i�#�<k�ꊟ��<+R�VpȨ�r�֢�heQY�S��L�����zý�#�i����eJ�XD�j�Ko��胄��{���^��H��*`��:+�:�v�X�z]�e,D��c�W�F��|��[2Y,��d+8�/e~ajw��dT��]��X}�����ҵ���y�S^�����41?g(]] S��]뛫��+p.���f����5[>|g��\����!]#e�`�r�����9X��H�cՔj|��?ּ̧u����Z�c=�Ώ,�[Cg��|,�ݜ}�����lP"���!cʜ>��%B���Z��T�"���l����"	����M�|�Kٗ��{O�z���DoC�갗ʾhن��9)}!��A���-5D����@V��m+�P71��4�%��7�f����yؘE����S�����H�c�b~ ��3��J��^����P@�.�3��?H�a�j�该R��M��А�\��
[�L3�K�Lӊ�Ш��l�	�,&{GS?��9�m74���G\�����e��-CgU��0G-t�#����z��HE.drEz�G����u��4(�$�=�#B��q���O���l�Z�{դ�ǩ�b�_�e�֮h��q(G��j��q~`����q[T�y������7Ñ}�/J2�_g.��W�ԕ�0P[(���u����!�)��r�R4��
ѭGqE�n��ә�f���@��u^�;���S����N50�Η�/�-Q��47����Ĵ.�v��#`5ͯ�B�<���o�������:���������������.���4���Y����~j4_)ٍ��u��2�V����Wg{A�Aa�*�?���)���E����}U�&� �ꦬ�q��� J��aR��G��#��`�bN��r@K@�Qh� n ($����4Z]�q�˾�-�Lm%ף��OV=��1䙧z��'I�Kq�z���Z�*����y�+>���������Ze���~��{޷�-��%Eݻޟ���|�õ�����9�E��y�A�p����P�cY(;�~��7`�'ܡ,h4�����]���Aw3}Q���j�ѣJ5+T�{g�"FV�MI��#\b�z��u�����e��j���G��OA$T���5�����7���t�R�w�^��u���h�H��f��(�O�L*%LQi�i�cФ���d'?U�3��x�%l�+�M]�����da=\:Jj��Ɏ"}�k�0̋T4A�-SaPX�.A5�Ts����z�A�l{�ޢ��T������s[��Wڧo�������gDLŦx4���î$�2�or�C��)K��l�nB���^vf�~)�ʽ|G�(U�{֑���g�x�U����E������mL~>y�{��R�Y���(Ͽ=����v+S���l?R��\��P�獢@JZ�j�M���o�L+��&���T�����v|��{<�q1e���@�w?#�i"�/�6��1֙����.t��N�sѼZwF���<i���>��.��gZ��&�4ޢ¨�J�H��@�j��Z��:WmHCE�����9'��~`���d�f�f֪�CUbv��ۏ"0�����U,�ے����&c��D�uL��k�0/x�_MN�t�܅�ފ� �K87P%��@
=�\�6S��N��3�?3���g�aϰaݷq�6B����VPiF��&�R,�3���U5�"����ݢ^	v~�6�]>�8kP=p�K�W6��)��ݥ�J�N9��A>���4(Y��U�J�^y3���$M�/����'5�g���M�������g�ʙ��J���N�o?�-q�V"�vi^��8Z�U�J�m��#�QՉ3�����4׉��no��'���b��	��w��.Շ�����m!z�d�]��z���jq�l �:ކ�`ƪ"8�JƕV1ع�F�H�b��:����S�Wm�%N{V0�>0�z[�f�Kw��f��x80��rؐ|K$c�7] 8�Cd�����'*�3Y�L��?[o�kA��>���	�f!O�Ⱦd+����0}�!�-��}+���py1j"�H���-0��PQ^�8�+���Z��-����w(�g�#�Y��Yl���9��4���ܲ���?m쩅��r[�6
�-S���K��f�+9���V��_��B\��Tt�>��<���J�+�[RQ1S�w4܌g0D5��<��uc!h�L*�Gt�1�B��"�ۚտrj��:�nz��iL��  ����c�<t��S�t�������#��6�fak՜���n����bv@�0�9p���Y��l�VfcK%:2S���5e�#GJJ7�q�ĭ;İz"�<134tc��w"B�j�IWc��"���Θ��2�9%���F�[��U��1 ѕ�,�.~�D(��������j6-L5�.��D�g9���b�r�v���&;Ո�
ebd��9 ֳIBa,��t|Rj�O ��[�{ҭ��$ő|~4�����5@���j����T [��}\���1�[QgX�	S���p��, sl�����7��ۮ�2��:����6�=ŗ����Y_���y���fK���dN�9�Ӫ.�ġ�Yv�ƛ#�oE�iVokqO�)�S�>�\�T_��.,D�2�ؑ������m��o\�\�A�y3�b��6$M��E�w��;i�����Yv��'��'�>��(UVGSL�<brb�,�ڌ��/
�,�OF�`zQ61>,˿�Y�EW�wEC����d�
�w��G��C~�n���{7�c��k���+f*��=?�fz��+yk49�n�΂����,�5R{lo)z����^. l�$�ƲS���<B��%\!7����֥�?�Go�)���&��67.I���Y��<�����0.���K�~��&�ҙA����8c��R�+�����C�3�
�ޒ���L+} |��7�5w0����P��'��}_[%+;a�7�@�;�O*��I�&�k����mdM�,���V�?�;'�˥(M��1�x���1�5����aݗ�Y,����H�S�}5����Ǖ���SB�3��|�&�L�R)��ŇQ*w<����QzӾ_�c���Q�)c�7;�
�@|(�28.��DoЂ��E�5a���܈0��r��g�����A��J}c�H	�pJ��N�*�Kk��ر|�֦�Ci��2VPV�6q��Qzm/�AOt6�Cj"��<¹Tnw��_�[}@��L�cT�(���U�L?ߦ�;��Ё&-�lG��;��3x=���Al�==�<���|�!�3������曲a鉓hU��H�5�9�����x[ρ�e�0�̓h��~�V����~��w�C�`���2���U��>eL-��A�S��
|o_��u��/B�� L(3�@�U�h_w�WY4	�<�;1c�i�N�& {<ӿܘd�
�S��@�������h�2��/uR
��}�>a�E�la_|z,W���W@�a�3��â�e���k�[� �1Y��E�>q]���M9>�;�u�)����h����
�AJZ�ruA]�RҰ׌	�Z�c���Y�l�0M��'���H	&ᠢj��oс���_�oE���0i��|%��Zk�ٛ!o;O次�j���Z�^��ޘ\^��ܩj���U1�s�e\�l��[Pߨ�ܞ��\�N@*S��ty�?����E�Z��Yl�u�>���i~��t��{8�z^8H������=�
�r%nS<C��Y�>�n���M���IJjU��M 1�?��#�L}9!ww�w�5y�@M�{�6�]1h�S0N5��wu���@�q�4x�k6œe�~ R�,�����G�l��޻ t�C�Vs���J𮦷�Y��Bf
h!����)S��k����$��&�k����-"�7��:��O�d��WJL�&�'.�A�D�uv�� 7���*
b^��0=���8#��d�ѹ�I�A�i3��Wh<�x�����#�`LW	3��o`�.������s.��*��}��[���i�V���EYm��!F+�$�)|j��W�]�>�XR6Rk�;�dn^�צ:��T�AY!�c�X�z����V2�߇��7\	2��������c��S®�0ޯOu�0K9��a���=9J0�<�����/%	�6����ߋ�#�Q�+n���'��ayҲiH�9�N��q!1��7����P���.�E%��MCrT�Ƹ�<����R7V�#�<,tL���P6��	��!�P�d��nf�!w������"u,��`���D�{�e0�r�A6-���� �p���\�����~b��ՐS����d��aZ)�w���t��6�`bR��P�3�6gd�z�]b���_�*��������&!�mC=�z��&u����M��L���ɚ1T��*�>��L)6��֓���'T+K�q�[�Z�C�>���B��I�^r����{�%�(lJ����4�ڵ~:]G��!Ζr9�՛�yߝ�N�pve�͝BR��5�n6�~�N1#>��בּ�2`]|N.�9�꧍��f׳����!�fRcY��L��*d߇f���C)q��.��Dk�	���#�p�9WF��2�t+ѝ5Xl���X�N��LB��rb$7g��V���7��Fbz�6����ڊ#O�k2�]>q�����G#�5�J�(6S���l�m/���Ҧ�w�3Ư�9���S;y������C�Q.t~���u0H�n9��A��E��$6
 ��:��A���q��;%NX��y(Ź�x�D�ߐ%�)ͧ����m.���w���ٕ��u��A;�l!�
�8)=C>&m��5l��a�VNӶv��s��u�)���xz�8@�WM*���u.����Eq����yz��_3P+y�t�F�W&5���~(�HC#畳���Sӫ�(�����P�]�N���A�E&���.��͘�O�f�0c��v-8>��~&7Ҝ0���u������h�����1�(�o�(�C�����n�Mh��?��a�C�|洩�:�8"�n��c;���e�s�3{%�<�TG�{��Y�7��\���~�{|���JwD+����쒱�._[��e�p�ao��vV����M#��,���d��53�!ܭ��کk�ԛc0KU|�KRMLn�O���TV���#�A�]kJ���0�ٿOp��I����ux�<
#��#�7�K�� �"�����>q��V���޳��2�MQ�����\���gS3*��	����Y�IP�h�uY-#�Ȏ�U�ɿ^{o�]P��j��6�.�����n@��_SQ�<5f�d:X��?6��V������D�m9��-��[TfyK�u���2J�+�9�ާ.��Lux������>������`��p���9qȝt3�;�9��Mk3���ꑫ�����z�R0��HΦ�;�$�<�Y�p��~��� K�����f�W,��uq�]Ȃh�ha����-��f2���NsYi�9�O���(�0ц��(��=rؚ4��(WM���S3�*}ݣ��8�ʣ�G�Y�r��T�k� �-�cU�O.g�Ub�K�ϬW�l�x�Pe���֣��b��05�����z`�Dg^���,Y��5�z0&w�|ʺRS�c�2��y��W�er�����u��l�fJ�Z�6q�c�oM���w�q	���)#/��A&�,?�Ռ��)g�wc��F�P^��q9�]�ALꀊ��Z2��J&vnu��'u	_��eH��ę4f�U�f[K���*z3�<�tׅ��:�puU����>�e'6�F�.��]5]�axa=����?컜IωW�؝x�/VMb�׼��6^�}�Ό���ʆi�����֠	_)�k���͡��/\�UQJ�I��|c��Ç�I�|4��=�\�b�+:	u��î6�q�t�gQeSF�Rq�2:�?��*�������pOޤޜ��z�\�0�
��U��e��1d�6�X�Rf�z�csc�y`��[*�5j�N,��j���d�١���.���V
���^\sk�I߮��U�Wl����y�y�?�ؑ1|���kX��ap'{�?�R�#Ss �\tĂ�s�W�~q;7G����v)���N�[ڇ@x�v�����z��ε|�F���_A�0:��pzڣ[M���)���}R �K��Y�=nO�-��e`,X��<��Y����[�М�1�z��e\���������bt�Lߍψ!�5���/��~�+�3�	L8��Ҹ���P|DQ��j���� �Mq���|�3c6 ��hP[��P*|wX�/+`nP��~�a5Q�"⫥Sy �|��iCv�4k�T�B6�1q�\F8Ҫ���%(�oS�m�12{=���n4���s��>�/Ivٓ���W6�O��s�:��ɫ����M6di�V�p��-��9���u�b��m(h4�&�],|X�f��K�"���ɱ, y8��?ێ��E͓��j�~�it'A����6y�����y�}QbWt�1 ;6P7E0����
�ғ��S�z�ܜ��|z} �<�r`*�� ��b�ioV�ڢl}(���Yq`�����-��{�ڎ#,�a��˫���:I�xeY�X�Ȥ]��O�k��!>�J��/HOqQݑ�Đ*5��ծ��6��P�,�>t�"���>"u� �y��hx�H�!w�M*�q�����r7�Ir�֙D�L�[���ЪM0�Xy�o�L}ga�B�~��t.d�
H��(&~�mp��ٜ�Io���e��w� ,�\���e��my��}�.rx+�z6�!u��
����x���d���ą�[tjK�j�ҝ?4�� z�%����lC�6�d�nKj1� ,��ԡ*l���0�NM!� ���09�{.��9�v�j�m����.������gU;]�V�7�	m˚�]���Y��CN2�Oo�dnO�������tuB]���;k�{w�0�A������~k�H��l��W�+#
ӳFWUd�������x�WMe�$ۑr���Y�k��_^Jpu^��40�����tuH\��ӝ��|��6���Z��y�fb|��	��0�gl�r�K����Y�UNx�04�r�aɼ�C&`���-�{ѻl	��\ɳ�R��:Ɨ�kA�F��<����q��߾����h���Z��//�b����H�ꁨ��/
숳�UUh#
�"Np��	�������όa�ׁzra�/ic�^�߂��*G�T@���_Ѕ��+-w�}���<�@M�>:���Ea��(�7ߑٮ�	4�F���Y7sȽQ����'�;U����}J�vI�u�<�O#�/}�R<X�>F͆�\���D�r��y���[:S��Z�Sc� f�O�Ǘ��l�3�2r߄ڵy��(�io�����lЯa��G����ӂ6��=�н��qw�A�?�tY9J�*Υ�b���49N/W!;�ԣ�5�ǗHI]�ge�Z�-=�����{��"'��п%�A��<Z�9�Q5 `:U|�8 �8S�j�^#�O�l�����$縩��t�]���D� ��ˡZ�u�Z�Fv�u �K����>��+��vځ����D��m��}�Zt��l��(���a���1^��#㉏s�����&G�\�μ���0��;S�������bjx���%>1վj�G�[��N&����	�w��S_��Y�CW1G�e/�S��-�	��'�rc�k�3���gF��ވ�R6V72c1w �|& �|T �6��m���Qu �7ˎ���2G8v@���O0�X��=ߖ�t����ݿ�A�#�@�#�Oi���lw��o��i .�
m�%j�o�W��;����Ou�N�W�63���W���<��M4j�|�Y.�0pw�������b��;�.�Eˣ>�0��}5Oi�M@L�|B*��)��zQ�at�8�B)$�|�K�����G�w��;�b>w�{�R3kO�r��m���u��2��w�6�^�RY�G-���;�
�}�TJ�D��3���v�R��*	J��O�K	��DL�=�|D�c�h�F��*~�d44����~6��!�b�	����^�7��W���B�63{k�7|��ixmi⎴��78��#�~��]4��k�s�����@�@��<тv�M�=;�8�[f���@Jz�����D��}�I
�{~<��N����+�Vo쐚@P<� �DO���~#t�6�Q�ೳ%}�z��ҕ,k���gW6Į�/�����@g��M{d��K ŨpKr/r��&{?MHd��c=KN�V}t�k`�����C�p�N���DUS-�����kcg|>Anvm=]\�n�<��y��Vҩu�s+N��D� ��u��z)Z~kG�Z�����ϱ侔ޓ��LK��%3�AL�>cj0dv�*�� a3C59�Ӽ����-2'Pz���K<��/S��'�3z���jrMll����YHuΖu'�ӳ��6�P�-�Ĳ$�(��XI3�5�㺮=-�[8M�M��t��{���1�v�s&	��/L�"ayqB|#�&f.&�}�G\9�����ٷ��"��p4j{�����Z��
�D+�4WS,J ����7�ܽO;Ȣ`y;�]�=	|#�j}���l�x
mOO��1��#�qዓ�hQ���"�(܌M�N��_Dn8Y��0�e�?���;!��v�/Y�y�ZQ�.�t�;u�Hw��ۏ���8�]k�.�´;3�ɲ�͚�}$	P�o Z�M�9om<�kn<�3T�"��ȵJ���u�����>Ls˿�.����p�tw���cFP��n�JMl^5�?*�����)�[���q�~��e������9��ı+8�>����\)�Y����ˤO�[�}�z/���5A��!����h0�I�����xؒ�9���2Td4�ʌ��$:��և��%�� &P ��PC�u���נ���!�':��[ec���n1-�*yR��"�]ˠ�'%?)C��Q�W��߸�f�L��� �+��C��zy�I}�״g�2��ypξ�*;����(��(�{G]:�c���%�������|�04
̈��}�z�g�cG3m%��/��ٳtd��y'�r	��=�9M�2�2�I/�t�O���5>N�79�a�%L�S� �� M�K<[��8T�С�*a��U��S��S���)��A�Á��	8�'��@�{B�����i��\ �>�*g�@��_�����ʞ��7�!T��D�*�5Uq�X=�mHkq|��2�b�Ã]4Ɍ�WkBЋݿ(��Z�H��^6:P���Qز����ZҸ�MbD���"���|��.~�=���v���oR,��>��	X�ܝԥC�3Ym�	���U�Gip)/�6��E;��f�Q�����Z�S�>O�>O7�iTMq�^m�I�ő6�y^g���x��w���)O5���� ���8�f�"�?nn���
��h�F�z	d�Mrv®�^q�ƒ�X�e�#)ϵ�a�HP�/9�F]���MnE��&+E�����%�NX[B"�*|ہ�����V;��x��	:LB���n�0�`5��`��D���=��-͟�M�9�n�c�h�%6:�����f�׬X��q�� ��3(3z��ўrk���������)�5�-X[~��c��؋���I�c�G�ʋ �~(-2��àSfA�
u�9yuk`O7d�}�ry���卸3.b��m�mM����a[�8��L�S�(ҰwA#S�{j�g��^�[��I��A����!(�e����+�����b�5z��kY2ЁYz�3�,RP���Y���ȣ���y���T��؇�`��?߲�ǎ?�L�(14T.�l��~1n�덯��hE��	�Z��d٧��z�Z����#�-�ՠ�;u��LU>z�����=��3g�"5�P�E��5�";�P�8�l1ʺR�����\nME���9�>00�¬(�j
�5.�����M�>�j�x�`fW��S�� ��A8�_�U���N�����^xC�w��K�	��6�YV�&�74�������&3�U�ٻ���ڋ�mt�C�y1_CwWx+i�~�� 7jM���	>��:�&��p����"���T׳�	Qf����{�V�'
s�dpؙ��a$8��	�\�����@&����e�k(󯗌������@�����쟊e�q���b�$?ֲ�l�����~_��e��_��Į�5��%k�˔g~�eB��'�.Ə�K��'EWֆ��1����:�剄(��oÓh�/g*�µeI6>�C)|"3 Wެy��a��Z��j�t�^��?��\���ѷ����F &oy`U�̵h�W����(��<J{�e6AY��A�}�Q:�v`�1����d�lq�ޅ�����0���݃�?e��R���.������V�����
�a^���Y w�_�R�MZ$�p��<���թ�+����)��P��q�	��g=bؙJbK��y����S��F�u[�B�&��n��{C��0Ray�8��)�r��.��I�����,J��A9x<N�����d��^�1����-�Y-	s�N�t�"�4�������77�2?�R ����<�RH(��2��EKo�e�f߅3�W��ʔ����i;+�;��ݢ.2r[\�g��y��]��9�$�S]F��ݐx� F��]���f�d��!L^�=o[��N���"gďQ!=	R!����8TS7{-���*z���X�)�;� �Ot�ӰP�R�QH>%A��X<2�� �)%�1��9��Zs�rg����j�{<^5�b�}�*9=�S�&� �0�$�Ay#H:�.�Q��D�\���kpgtxDw��5��7"�$B�	�V)n�9��m�g��	�)]��;�;*5	V$�Q��ct(r������Σ�nT?�rFlfEB7M��@�ꧨb���{��Y=]F�gӱ-�׀�X%Eq�3�����N��jB"���$���9#f\�w�z��A��ͅ`S����f��5��h�d2I���u�m���jw��\:8�>r�ؚx(���U���t"������y=�΀Z�(���筁L�ߥ9��hԐ���y���Wmӭ��#*��X(�3z&D����%�JUu�Ο*�)�8�(MPXA��4�2�t�fNG��㆗j����	��oű0��T����O��U�N���l�s��Չ^WO���$�%�Tʼ/ۛ��!�`R�#KH��s��6W�p�eU5g��!��䀂�p��� H���v�ݭ�RKz8,! $T� J�RH"Na`DA�s��vPZB�.�x��L��a�{�3��M�XZ�,��A��'li䗬�#�s�k^!��j�ں���;C�1J]`����lUmJmK.�T�?��:�}����h'ߩ�>� 悠%�"6"�lDF�:��^�]����\�6!5(<���V�c��K�a�10��Z�(r��)���� M��g��c���'  �V���T0�����`�}�
�x^��<�a?��`����t���<��#��:�8�\6sR�[�1[��|�x�x ���t�3���ۤ�:�6*>kvB+n�� �yA�;aT�a���
��ഛآ*!��Rۗ��NЃP�\Q��Oΐ5�Qp�����ϥdF$�-_d=C��9ra������z�&%UV��ȘB�o���Ŀ�$\8�^��9��l����;�]�N_�%�bJi�� v����+$�"�|��!0�;ڳ�I��(��5?,y��0����|��&G[o ��0>\��_����a@e��/���?�$�S�~�߆r�����~�e�a�;�=;���G6q�}2BnyL�Fm	G���g����?rs]]�H����7/_����y4��x�D��H^-�Y3V�G����7ƕ��2��cyH~�
m�ɛ��o!�"~c2�5���<&���=�<#=ͩ��w;������')�0��;6�8��sJ�6{�N�-|(2����^���C�0��j^{�T�,d����"�r�沧��
�OD_�k���V!���8�����?���7S�ҴCV<��B��:�2�{��&�&�"����H���%�N�>��	r�f팀�ݜ�7$�]ɪfg�3:;9��^I������G�I��>������,
�n��<RH���y�]�{1�ML9��E� .&6��U<;b�_��)��ҋ���Lz����B�!V=v?�NO��t�-=�.H#p����uwv�b(�4�G��bo<d ���ѻH��'�7�7�5��ɾ�ۜ��o��űR/�!kip�>1���:�������1bo�Ĝ�@�ަ�6��7��s��^{��=���@��u߸�M�8E�ߐ\��6�NpYC�n<0��"�I�.W� ��fl��U5^$�N���?L�o�f�⯆y|z�B@�`7�?[m�ˇ�fx�$�
4?I�B�h���d��}��s�8[��$ ��[�h�L��'[����n�pIUo����!y๘��59�YC��vXN��qw�ۢF������h��p�{-]��s�޼"sI�7ω���6����<vTī;y�do/�y�K�l��[0� w�:Ϛ�"�f�^DS$�	$刷,��������\��AA~�y�l�ઇ:yxꧾ��N�-J��� �����Ċ?�%�i`<��m?{���Ɲ�>�i�((ד�{�M|�&R�"�GV�W��e�R	���Y2�C؄��SSia�xז���>�mk}.�+[�K� �!�U�2ek�nׂ���R�i3���ޢ��wA'�:�UO��-D�>�-�eem��j]y�9����Gt���� ��B����w�^��EE�����,���~�k��wTQoW���z�ύc>m-�<>sR-ְ����.�;:��z�AtV~��+�݀y"m�����6�홯��O�&�C墪%�m���Ӯ2����QWo6�KS5�Nz�����.��NA��aR��kVz��9"��׼p+�K�?"��s-������'�k���f��)ں�������;����م��9�����#��g�T����}I��8����].�0^K��r�ڬ��4�Q����d�d��D>���ȡ��!G}s7��R��:B���xF)�U۱�A`<����,/F�5�9��鱢od�R$�ڶ�,����M[oR�C�΍Ys���g
�.���R�ɢ���`�H׍s���D]�>W"{�U�����<�%��o�lv�B[�<Z+��X�����[Ӭ���˻)`j����'�B�x9�
]�޹��1�����*M)q4�:ɍ��ϭ8�6�<
M<$�Վ؊x-���nQ�M�fR��=� �Gb�0ٻ����ڨuם�V�� ,8g,�o��F�s�퉨~Oޜ�%�Y�ˊ�U�)&Z��$���Wz�	�{��1��i�	M����*A�$=��['V��$�V��r��^Q�7.����M̛-r�br��ru�\�4}��ޮ�9G�)��Wa)���0巭:��-B; �������p����
×�e���7�7
ϫ��Z��z�35/1��#�ht�SvX6�'�]*�t���^2�.X)�f�=��c�d���d���F\�v�����n�Vo�7��k����������1���ꡫ8�i�����5?V�t�����B��W�xiq"��t�aS�q���M��P�s|S_�$v98������M�"�]���Z�z�U!M�;�9G�� �ocVř�+�܄��SW�dT�a����ܳ���%M�66���W�tt"G����6JV��=��Q�.�ep�i�+F���%���"��Ɵ���mRvz6�o�B�U��D8�y�ku
� \`ՙ�}�EUJ#� �Qޗg_�X�$�����m;/7���T.�$Sa��@�K������$�-��h�vrG_���6��^_S�F��8��bI�؍���o��J�;�g�)��Y�����6��~��i^8��Y��J֋�a���y���h����Jt+9-�枟0e�o�`�O���k{�t���Q9��5#�q�B*a�B8*�V�mr߅�Qҙgb�D�P{��0������9u&�\p�A��l?�S$�l.�Vz'��0��|��SX�@��F(F*��iQzt^��/I���5��dga�q��;H��(�dc�c�g/&1�3�Fg#3�����GPu$ m
��OU�w~Y
�|V�9�sZ�7��Ͼ�;���s�n�)c���,�w�]���؀uk'�q�rH�jxv�p���Z~�96fQ�?�:���8�H��?'8�>�@I��ł��kGuM�Z���d {^��@(W�1�@��v�rF?!o�}�|�`�	�X�C*hl6!�+���B6�S�����^�Z��� W�����j@�ꀿ�����u����Uy[��98��w���I�Bq�rnõ�n�(� ���ͧ �t��۝��V���2~-m����,��Ĭ�R���хV}<^�'y�KD$#�e����'����Mܗ�m��aQ�]����;p��/~b���r��ϭ/�F�p=�D����f�8��P��/_��.�J��<_}�� �ظ���}����u���n���z��|ynB��7�jk�����j��K 5�O���4�ۣ�i��ܑt"?���m��an���=.�#L�(��}�~����l����1���>9��]�Sls���2����]�8A�	
s�v:�����އw�{h�Y�4|3R�*1mit�(��^�aK��� 3�Iy>�r��h�Q{�Y��q�~���}��_.�L��L`f~���"?�&Iv�YYSm�g�Ki:�dT�K/h*�|���������'�����z��J��(}��T��X��d�_%"U���
3
,"�3����(�";��LPlڏǳ6w�Z+�L1f��O,��[{�B%;8�g1��c�h��0'�E�v�ڜ<�'��e�#�[��%���?0���������DSٴ��O`5d7�s���&Za�����b������_[�@e��y����F�-?�9���^�"V���o��ߚ��l¯����� ��ӡUˌd�D�S�\հ#F����!��=�d���LG�K,���σ�A :+��������>T�;��8�˝�vq��O�0����s��M{7�ڕG:Ȯ6������/SX��"�u�v�_s���ud1))�|H!�J��ĆA��C0W$��E�#��h������'#U?4~���ټ��?d6*A#mX�X�R\�ר"����'��f���9�l��Z��fpDb~�`�.���ɂ�˺�s��߰e�&�����(j9�ƫ~b�V�_ŝP�ck�-�$�u`���D`W�3�~c�ź/��^�xI��}8:�K�A�t�}�D�sk�bYJ4ή.	�]4��:�3�����T�t��S+��A���X��QD��H��ɬ���)�f4Sl��q:�E�G['[�i�+;���z]0�a�x���P�rB���}ؕوO��C;ɹJ]�#�KZ�HVS'n$N��������q�\=I�,��]�$�&��^���7�{���\�
���)����fI* u�/��}��� �'$'����"E����@vv��3�d�����#�q����!X`B��Xv��rw$i����fV-�U�H";�2�j=���[�5O����^�$`Q �A[�{y�ĞNP;��Z�{���-�/7��!i��ʈ�cn.\��&������Ͻ
�Z+Y�a43_�n��u����~��u�A�W%�.�,� �:�xc��P�!\�V*g<'��d�+s�9��
O��d;�jv��8�LB���V�	ZX�uv����m���@/ ��-���A?�� � ��%�Ny;�^Yk������Ě-��ٛ�x����$.~� gݿl�����7�#ε���	��j @eq�x���Χ�.G����@��Ob���^��=u��d����MWG�����*~ɛ~*+���Ȍ8�mj�!u�V�G���Z�7�
�H�>X�bN|��x�2 	V�m�$�0��H�	�͜k%����	�/y=e�K���(��s���T��%�l���>o�,���f�����*�ui}'�e��w͖""J���NQ�G��1't�p�G�id�ذ�S,�5տ�5y�<���6f��bڹ�hvr���o^���_��AǛ��)�~�W�`�^�f`�r�:�c���U_a<i�X�x{�+L��#�#�#|�i.+�DC7�<�4j��<�Pd:�]	��q��Z�I�`{_��3}�[�j�؂�D��O�)ovG�AތMOZ�O~-�8�S'�Zp�Xe�i���ڜ��E<�����N��0�o�9�V�]+'6�iƲ~\?�^(�ѕۯ�<k#���	*��,�f�Hl���1Ac��Z���ZY�3+�,W5Ɂ�^��V_Bp����M�0��[���`H�o����g@5�b�O_�7����P�b�Á��l���[=hE��s��:�t::u�I�ր�`Km��P�%������<�`���gQ%a�� �jѸh���m�H|e���Tm?�_�����~����MqM��F�_�2O5^U�ZFM�D��LaUH���4J���&M�D�i����n(X	z�8� ���J�t�~p�`=7��tr��Þ�9�~p�� �Ka!^B�A���\�za:��|���@whD��Nj��n���oЅ�5��sb^~~���v�úQ#ͅ7���b���-�ۭ�}����T��$J��{��;�Wv���ןZ+�_!�j�#CG��&���6^�S�\b�7��Ӣ����0�yT�fl���3jAνنYʛ���f��2��W*�VL��v&��҉d��»z&��)��HZ2����ui%j��[��عIY�=s8�NRњ�j�(Q����h�A�q%	(�f���@t��8��#d�����Y2�C"i!��h����񀕺�\��d�g5����dI����mߔ	#%;V�h��=�m��8��kx̍�P
�����������W�^�m����ӜlUwg�\��.�-�A�N�c���!g��*��	
� ��O)%��G{�P�C�'�'ζZÊm:a�s[(�C��>R�͸�����Qw!0s���� 1N='별�X���J�?�JKdb	�qB'��g~h���CZ�̾�#��Q���[�8���sh���)����Pg�H�8z�8BP�E���}�XC���Gf�����j��˘UA��;ɜH��E�AF����ծ�ѻE�-�!݇Yl���;���=,�=or����P� :�N���[^_K|�"{����ڧ����d�% 	&S;Bs�Ng�����텁᲼	s�p%|��)��d5z��fo[P�}ꅸE[oS�Q(�h>����A`FW4�����ڰ��8�(=@�Ќq��q�<��/�S7�ݏ@�C��y�f&Kl���e5�ɫ�$�3�G䬽��¢�������(��d����E��#u��c]�k�� rs��44wDޱ���>&����O��M̽u�)�*�ʏl&�>�y��{�-�)�.�"�����/�:�#�Fނ��b��ߘ'eJ��bYg��^7^�4|�Xj�[�/��6����-BL����s�>6]`�&tFMZ��� k�Hy(p�􊴔����,�%�T��5� ���RT�tԷD;�d�p����!�~�|dH)oG�f�8�p`�Ho�@��.�y�F����t֬qMb*>��a
�lu�������f{���:�Z�ܮ�z�`�����.9��?<��Q�v��}ӿ~�pv�y_���4�f� ��4���%=�P�6�fE�sa(lp1m&)n�`��wO����ꭑ|Ґujcvk�Ny��b]}��&���B�+@�L�j�۬ްK�pwDC�u�e�z!�y��S`��±���O�I���� �/��M�ʖc����)E4t]��	�^�KS��6�@���)��ԳA������)M��G�����a��~R��	֟x�US�vr�J�h��@�D�r��(�=hA&ݜ�ϑ�z�/lTv�q.-��mn�"��Q�� ZD�n�
fw1�=����R��Y`j���{Z�A|#���_��*BI��/��v�Fc�%U+��K]�=g��|�����TU��QG�׀��kю�(���q�
C劜���ͭ�C��9�M�g]čz<�_���!ͺ	ӡ�`��P��fYb��E�K��w0���%���N2�<�|Z�j��`����[����ʱ��B_�Űn��"�n� �L7����I�%��|+.�Nk�� ����ÿX��}�~������~�ű=�?2�>߂��#�P7-�^{@��вy?e�7N���iJ:��
$}�M~�"�Dc���7$?�=� .kU�r��@��X6���H�gLͼ<�I�q\D����Tj5�t���.��[ՠʢ�L�m�mF�Ɍ�VidB���'�\!���1`��;��r�7�IA���*����A�(�������lP��F�w�}UƝ����E���?.N�{-��ckv�߷����CmJ�LC�A�LͺK��6R�SUhAџL^���Z� �=�s`�Ӯ���	��9�}\���0�V�2*�O��J�c�_;ö���e�_Ql�T~�8�� m���(��"����'��G?�m"2��P�zܞ�6֝T����0*�x�d�"�����	b��r2jh/YЄ�cy�}%l�O!��ߤ=���{�=�^`�%�X:<�pf8a�����F,�cp��� �'t��g@̹� p[>��&�22�o�YA�m,`k�k���Vx#z�"}xa�r}��tΩ�����t.�g��QHyi��7��|�߄��׬��yk�]`靌v]	�7�@�b�w �Mݰ�Q���˻t�,�먳g7gW=�:�������~<��$M���^1��6�T�T�y�bv��w�l�w�BӺo��F�������6��K���o�m2�6#p`���R_4��ߥ��$rv�t���O���G�g ���?�|�g<�Ĩ^%Ϋ��ӄ���2�g;(���++�8Q�������u�/� 
��w�B)�6Rz���A当���?�aUP��>�ق�x�]�Y�_P��`���,�̷\}�)R|G�$3$V>�:���\��,~����գ-�3ZR]
%_(���2���n��i^M;��@�-P�K�`5	w�g����>Ke�P��l�!3l���e�p�����qc��ԙ�U\58�ܔE�@Krt"V��.ލ��S�OFCS��58K�7�D�R��ᵑm�xͣ{s�:��"FR#/�tZ8�i��3C� 򟸈�#&]Tl����D��%xV|��c\�"T�e���,;g��O��k����d�I�������/?ҤWg��7iL�d6e�0�Z�m�J��`��rXIʑ+�`/�Sh��Y%H`�zIH%f;��uR	? �(�G5C,�tRd	� ����x���n⏠�գ����#]�DJȼ�gډe{� 	�����4l���3��d|������kuK#� O������s�<�*����}_y����	�͇�2�����@��������_t쐾*åg��i	�ٕ����*"�v��k�҄���u)��7�hl��׷�ocwr�3lv��da�zT�.��ؙ_�٤��3���c���f1��>*#�:%�<ȗ��*��Fo�mC~|��6�0A��Çx����3�����@)�!�c6�����`�f��/��o���[LªXM~�Ə2�o}7�ǋ��C�u�^�F��\<^"�9u��?�Oa�G�̪0qx���Y�r��ݯc��\��g��@)ʲ��57ޓ�|�Ic�_�2���;�����(�@G�!T��`�Ɓg8W�޴�E��6��W�xOp��԰���~�5Ǫ�Ć���}VϦ̵S7�ٯ��2yʳ=j�8�"�}���X��V
Ɓ�jx`��꣜�T�O��y��g���p��F���:��RS'/V�H2N�Cw�n W�W���h�������b���u��$E>��9��ٷ��.�X��wo~����_�ӝG�'/�y�1F������ k4!RO�"���hq��B��4�� v��Jd�b���s@��s�V-��ɫ�'](�y55�n�@MXн}��ю��ⵣ����T�H,'*lJlF��I?�,�*�.��Pk�kkL�G�653��'�X��m,���	̯���X�����Rlg=�T��fj<Da@�/,���tZ��6էD���3�6�����aY����ֶ�0�׬,��*	��*��30 |ïUfQ����V��+_�A��¤)�zi��S�YN��S��l5����SS��،Z�lX�T?�(�ʎ|mAOaRTd:@��?jC��pP'�1��؎f>�����abnb\�ŹBll�af�Ѣ�f94U�X{`��ZUT�O���%#sV5�%&S���4s/+r�����B����6&E�c��NV@X�l3ne�u<��p��cGeگ^����!���!Uih��Ȧ˯68i�-.�P|c�2�O���*J'��J�2���MiQ�zsi^Z��ڬLJ��ȵl*����b����{��`�����*mV�s�~��T��N�bT>�/k�,�Q`dS=��viiTcI``��*�A��Xvtzk����V��M���(�hlҾƤ�pu_����W�WON��jJ;EfURHb;4fcYI���E#����{}�õ[	޽��lw2KE����bYO(ƥvAL'4R��'��׭,+�:�t�/��yʨw�%����=8ڭit���կd�l���:�_������?I�Ss�-���i��ՙ�A@���`fH`0�ؕ,j�d�lli63�K��	��R�x��`�?bX�P+�2eIc���H�;�.�6\��7�4�1��ܣ%���U�>H� 3Y��c�W ��߈�?A�)�S�.�v�H�?��$U��P�_ܾ��$h��7�����ط`�z`�l�(`��a[�� �h���E����aA��}�Ѝ�ߢ��g��A��l�č��o	)�H]LS���/��*�hT"!�_����[A��p���a=h���C��S��
��T<U�m�/�Mx�	J�	�k���3�@W`s?�:�i������AĪdaiR����>���WϺ���G|�-�id�>s�FM���i�[:��o��2�6�}\4��������
�oC>�j:�_�����h�����8]P>^��
��( �!>ք,.�,�W`�!e¨����u������S=/m��N��q�F�X��]��/����h��8��L�xC��,BW��p(���E���� Q�������D�s�+�� A\HA�h1\�zT�&�\Z�L���y�\��U�T��_2E��T�����F��P(ʊ��vq���|��^4 ��R�P����!����S� ӿ|t@�	�����Z ����B^X:��9�z�.�,��X�}��B��"�go�辺�M�%����xox�7�	E���'j��F܍{(�!.x*�56�U%��3�:q�q����):������:�?82���M�'C�)��^�LP�n{i��zj7�eW�g?���@��a%�`����9��8`�1[�@^�]��`}��!b���u�Dͨb�g�@<�xW��g�с�Z+>���!$�
E�¿
�`���t_0��΍�yF�@apN�0XI(����bj
�t!N���>�oD�y���cHH��"X|S��r�.��k!�<��oH(4j�U:�0�ˮ�I�qW���0��xaw����8P%V]Pl�}�/B~{�'[z;�?��B����36dq)����`�!��7lϭ�t�nn�M�����+�@82���ƭ)��i-ZDʋQQ,�Q�9�"!c$dO�S���U�"� "R�T)Vڶx*�J��J0��	���0��Y�o������;�C��J4�s=m�O��<����7�<�:5�f5�Rw����A�A�^$���I�$j�@�B� ʵl�揟:�}u�w���% G��?sTV1�륚N��U(�4�./󉐵��t�!�)��c˒�}���B
�7�-�K�*��
S�Ծ
JTW:ߔ~�"�u-��,h��B	�x-��'8^��-����y����Z�����6yo�� �j v�Z%7��RWG��}�����
GT.� ώ�!n���Xb�6����q�9!%4"�\�{�w;n'�JT К}L�)c:@���˛�H��,Q���1�]E���q��ۄ���auć�les������	��qt�F_��K���Q
��3e�'i=J|�n�
�0��9�gw�̵���n��-�{	\9V�K��K.l���<K��G��w��Q�7�t����:I��`0 ��[�������קCl/��Sg*<Hp	�����-��>��S�ۤ����-�1�5�P�d�V���,�I��K6qu˿�_��Ǐd������L5{���2�]�s������ГlD�[	���� ���ϔ�7��e)� 6a*NT������כ)�f�L��b>zl zί!��[���+��簰C\��0>��Eg>��n���u(3>š��}r�	���-Q �T���=iJ�dc�T���e;[���2�r�L��b���d2;��^�w��"3|�˭eC�� �k�� �����@�I\�Dm��>o}�Tw��+4�%B"ʓ�ʕ��fUy^U}jV��T�J���7̪�*TU�o�n��Z�!�?��#yfH�VF.�/�l�߯�u�x��l�O2���~q���K^�FSk��)߿�j��kc}O���̄���{Mѯ�/[[�5����X��Xc��\�I�N�h�5;����To
䯎J�ix@~2�_�y�������.>�P�� ��S�v��MP=[1&�~��
F^�no~sǯ V�6���}lÎ��'Mz��u�x���#1kz˂zZ��߃�O�:-!����� ��O�ԩ�7�:��9W	�.�#&7��%�����Ӈ��=��Su��7�{?-�������U�l���睐H/V�~GO���=�h@?�Y�3Ed��ޑ�܁	=�l��r��6SS�QI�}o�_!�j�۲C�Ыr���,�$�y�
�w�#��*�[L��\�0`�a�rue�9RD6�����Ē�@N��a���_\�V���e�-�r_|���ڸ�����=t����������!��w�X�����yb�@��/?�E==	o�|�q� <�uVN�T$OB-{�B,{�1)���b���3����oރ��+��&7��j�+����t�X[xS�qL N���S��5��h��ʄ�#�F��)|�#��IC���G���3ӭP��X��,��߮/{��9W �Y�Ʒ=��;.���/w���qd�\�����Gp*�	I� �}#-W<5w���{����D�Q(�AN���{�[��T�zKδ��8����Ks��ߟ(��4���(���)����]|B��j���M8b0M��"�ƆN������Xn>�!8����EV#д.Pؼ:�e2&a8���+�}NxfW�J_���u�V�E4�F]griσ6J�	��4�}I'�5��O�V���l*`�h	���$�ƆM���7��V�OPG�^e��M�P�$_�r]*�w�Q����Ω�ڀb�	�r�t�a.�t� .�|O���2*7R4�i�l:�Nfo��'��榼��]������$�tʍz�}�[ٿ���%H�?恍J�'�B���R�d�[�j�开�� hqč%u�s[w>�M|�\tD�u��}�p6�*{ۇ_��V ��G��RB̺{WP ��!�sp�xt�$���N�%�/u� ͤ�}�p��� W�+�͋���RX[f�<����h@^������&���G��_޶o_}v`�v7 �D`J@�r_�!>Y:)�n�V1'�C�نo���a��B�]�D���R}��e�����}�#�Q�|�=���-�_��- 
��<���L����p~<��Skxł���D�V_-��@��5�Og@N��UtV6���BAڹ���j�"����1N�����.��/�A�:���.����e��e�1���{Рk���@	w K@����҄���I�����,���B*�l�e4��Cj.�U&$H�ֳ��:"��R��p�Es�Yq#�2¤	�(�IOL�,*�&����5���������k=?7�DOg(�O��P�I���I��4�ah�舱���� +��֢�r��SM5�ћ�C��8ُ���6�׈�'�g��gi<H��J�W���U��G�jp��ip��8�s����W�;�OI����4�*�e'/�bl�!B��b�R��VQr�v���̿}�lȕ��5Ě{�W_;��6�]d?o����3;<�CPX��Òk��;Y�o	�qUZ�ڣp_�9ϦZ#o��[X�~�6�fgܲ����2�/y(�R��9F��?�+"V��<GL��aL�E��$���ȝ�%T+�0�2V���'�ҵ��������j����nN���|2�q�_V��r5A�jo�}����,7qmqˠ�˗�Ne
%�k�k������Фҙ�?N������5s��I�7	ݒ�JF���ai@?��/z��4�X��bA�f�r1���}�3�)�XӶ���D�8D��\"����xF�+W;6��j^�Բ�"l�� .�П#�Ӛ㹳�<���ǘ���S��6��������$M�:���YG��qZ���n�}��=5�3�x=P����`fF�k&����Y��}&U�O��Q��pV	�H�w;� �Э�
HF�3�h��1i�N��#e�s���g��$Ș��8i&:K�{�1)Getj����1GG<�-bz��6ஃ��B�9�֤�(��N'.T>��s���4���n_l{��h���WM^Ʉ�<�˒���#.��9�k�a�
J�.?��t%��(��C=_�`�(fp���,%ݓ0�S�=;3q��ׂi9�a����Pyq�(����11a�I���:���*��R����99	��Ì2v
�ࣻ��Q�^qQ[	Ny_Z����~#0���)4��)=U�T�]!k�Ov6�0�� �;4�fѺ�S���
g�APŁh��X�\pvG��*WX�)��Q��;��F��z$������܃��LOa�X���6y����i���f
�\��2����|Mӽfw$1&���F��TFG+j�}�1���~�9�`�I]`e��Z�4Āp-+k.�p���AMHC?���l�������T���ZT�xw^�mہ�H��5��{os��σ�\����C��79�;���G��0$�)�\�p-��Am���Л^�� �"Ū��Nܗ���Zo�&��\��^לQV�=�_���标m�V!�� iÇ��Xݪ��+��4�#�
����Q�w0�Fi)4��SBm����$��}�����C�`^���o�dz�=��G�u>x:�=��Z���^ n�h��-{�ٳ��:sC��F?-�����г������`�\���Jyv!PϨ�*���̝�*�d<,D���s�ra��B
�@���"F�^x�i�qz�L��+��]��g<'���XgȘkCZ�V6������2u�RC����m���|����a7_�D�J��Z�cLzL]��U�ه��o�cb���T�οH[*�g�#gw�����J���e-��qf(7����O�*� ���&��P;V����V��74��騷�b�1-��N�N�^�zן܎|����ø�9w�7��8���Y׃qp��T9T~��Z�pU!y�}��x��ܨ�կ��dx��y�ǒ�%I�w&=b�<u-�r��_�H�pW,���r����4z�Z��>B&S�C��N�k��-���i�il�e�PV.*������X��gN����`��ZOJE��2>�!���4��*S�imY��8�-d�V�.�j�)a�B�j���޵u��S��_�Xl�4h���z A=9_h����6ش�Ѩ��_����+�+}���.����B�m_,�g>��30x�5��tO/jr�TO�&L�n}���fx�l+q��I���Nx�/�l��҃�HVX;$�l�����e��u�)I�������Aj��zN��)=��GP�~:Ȭ�\���i=���v�m{RF��e�9����Dx�H��<h����P˚ȵ?���xĐ�?�a�-�(\��T�����HZ���Y��Mά0#U཈[s�t�N�z�LS��H�o��K�H�;�y�hA�&p�$qu��G �O{��M���5�0ZI��]���գ<l�)�s6 ��N����� � .o�W��%/�J#:8��f��i�@��ҋlm��!��\��^	�tsį�zQ�.�YI����(]��fj�B ��mTug�����-�/�����a���z)`/���򒬐	`,��$'fOdJ�	ۉ��s�Z	��CϠN]�B
}��kp������9�Mb��.m¢r�G�nM����[Z�b�?�<q�Vyҥ��3��*�����/O����L0�~��-?q�7<�d씔��zT�jp�ի�:�a�hR�z�9	�Z*���:� ���(DץF9(��㺖e��x�t�w�V��Uv=�~��И$O<t%�-�������Te���%�R��]ϗ����A�2Y��Cq�X�@�#x�>`T#��n��~��zN�ui(aD�t��9�9��Jh-ʢX؞����huO;_{,�?����y�sQj��u����g��$��D<�b��[��:&-<ذL�+���7��9��mo��	��Ԝ��c'��~,F��q�p���I#a��EUuUxA՘Q2}N� 
��<��l�!8L�W��s�E^Q_d�{����i#A���\�|�y����K�raڿ�f�g�F�����P���[ֳ�<��Lu�`Ю��y2i9D�Ī�n�N����L�Ȩ�M�'�s�CN#����<D^�R4,��w��[�!��M�o,</�Z-��8V�N@��e�D��q�j@<j��v0r���ƺt��)�|bTޯZ�֙�PO����*�:�c���|���P�_���o9[��ܴP���}.��k�P��S@˧�8Z$t9�ϴ��j鯅~�.9^��#��-=9�ȈM
�P��_�������?<n,B)��㛄��Q���E,����F4ڌN(j^�3��P�N|�z)���H��� �6B�l��2��]�/��}W}�5�$�JMĖ��x
d��=sJK��7�NG[E�ޕC�%"ϻ���bp$���i��a�y:��V�H�]�
g��"��X
�j�D�l�ˇE�NF�No�Y����X���
���ک�2pV�1ɃOB~':{������*[8�t�w���q5 ��t�ʀ��G���M�F����U����&,Z�/���{6}�t�x!�<Sq�ܢ�'�z����GPN,�=<Ҍ�-�*(�~�b��Y�u�|�?ul���	��Z͏� ����m	�4��UWս�!��c��S5�_��e��݅$�]I^�����ߚ�R8���E��Y��,	Ml�jl�a���<t��Fy�q�xF�۲�գ]���ˁ2��ǹ���(��ph>H���BNt�F�%٣���C$NA_���$����Y2��B�a����V���xh�o[�7��/�\�i��!޻��q��l���_��m��h-س�I{g�����D_@��Zb���z����4TN`���m�?'k��Ox�l���G�c5��$m����A�s�������[���|�t*�`���*lA�H���[�qO��l��(�iS�>;�N��R.t�z�k%4���m',�$�;�	C�5'B޴L�jY�"݂�/z��ݫ�#ujt�}������|��P{�ζ�-���C�<-�%��x�w.�و����wV�ls0jno�W���[���z�Dڏ���l!﬈���r��f���ipSHJ��^H���� l
`���"�,�
V�&Xm�ٶ�d����<�b�\���YOw\��$8�V�{�v�4h�i��"C�ĕ�׸X��mֵ'D�)8R;�U��'(ś=y�N�σ��\U-W��
��u��,���3��c�K������Q���xp�&�F�s h�~��K�MI� �S��@��zվ�q�	���s*�W@�\Xf�B_Z,4��F�b<uxA/4r|"��9�m���t���YX�g����ZwI��Ň�sJH�&{���r�<����Ԃ7�w{vȊK	{�,>��21��0�gc����Oc	��j=�38����H���+z���Y�v�D�߇҈�ݐ��_
i$���5�eފ���Ķ4~�%l;�����7���A�	��<�,��{�ޖ9wB;Y��v��a׺�D��y9l�r���iY�?̵ �Z����r(/�Д�]{�0�Q1�Ata߬:S�	�������:3�W[�������?�,��CL�F�t����z_j|;N(�8�HP��q��L�������9$;�4'5F�IM�Ӷ]�J��k�I+����[�<��ar55�,�q{0{GY�����icȞ�n�0�(��d;�����M=lg���w3�%��Gw��~��j��֍C������,;�3_!�a,.5�A���Rpk6O�Jj�g��p����w�d��,�^z���i�EF����}��*A`p���eO�T3���<���Jȅ-U��m��2$�¦�xb�ߚ�5��{��N�9���T��c�"Xo����W! 5�*`s��Z5�t���9���,�����=֒��y ${^e���Y�����e<�|^%�hd�gP�Y~:[��[����m���F� �X4��'��6 �\0J�B��N=^k��OR�U#�9��������VXO��54z�:K�����?�{W	���o�d5����O%Tf���|�|`d	.�*m*ύ�EY�g��<"|�#}vX����I����
v�u�@�Dz�����sGf&�(00��
 �kwN�NJz.��.�څ�,ٔ�=u�z1�Y;D�h��pB�8JwpN���+r+i� q��~��9yda�߳l��z��H��գ��'���49q�$>^~�0���{�#�r��>sL���ҏ�va�>�i��ļ�/�,��!�k�`��6	]I��r,WX�)�t��\�&L��h��5~c��e� F�/^�4��f�����4_�8/��p``
�$܊��41��YDf�Ӗ�]j�Tz빮�1ޜ۩�L��93��yi)�C�@0]#"��*Ō&��xb�cj)�k
��!DPs��澺�D�æ��:�I����z��b^�;�3��ɱz���;?,��0�$�̵��~�_{>�0�/@je��蟱Z����m��6\3߄ )"y���%�V�.ɫ�ƿ2�a\)Dƈ^��{ϛL,�h$+�5���:T�a0��f�#u���t�N�uCY/n(��Ȑ3���Av��^و��O����,Bd����4�_�ڽ��nL>	H��in��[���k�'�xB��_����1��=%o��a�2�.���ŗ�<�v�`���ARv[a_@�WHmx/���Y����V0�INx3ޱI�; �a&����_H#;r���t�������y���v���H�{D�ẕ�!:ށ���XB��6����P�Z�j2���i�5G�W�ê����dRt�k7�Ga����Y�~�̯����m��g�ٴ'���;�!R0KP�fvWoM��h�΀'�oOHt{u�^���������e���D�&�Rgct��_�a+�0�ܮ�P�ۚ5��5�c�c��-/��є���a�Iѹ�e�76��xàb�Fw؎��$v�"wp<29�-�a�n*2�A�Rl�t���'���-8�+���}��pal0-$��4�I��Ϙ�Gy���z�焵]5;�4�yq��)G��<�9���P��{]9���kó`���Z�P0n��7�>���/���Pp��q������NK��'� �U����� Lҁ;��W�vd�&<�#̑}����II���@
� 4�Gv�V6�<u�����jb���{��AnL1mU��L��;J
��Y>a$u��ëJՀ�_�e��s>�^=J��t����U�!Wn3h���n��a�0&$tΥǍ��DN_f픐���yYU�hq�-Rp�ڹ׫�۩SU��Ak�N�بD�\Ou2��'�jd�/��ߦh�S_�d�D��4	;s�c���V̙d�-�t�o�J�-�G7
@��ϕN���z����
��|���3Ea@�n�7�]���˪S�|飄���疇w������9c&�{죧�F�750b@H`�M�� �z�@�B��P�f�|9�ow@M�7y(\�zk�G�B{hEH
	:G��C`\��<��k8[֗Y���/��;���ׅ:[n�	(���[|���g
׏@���R�\i�x&vY���Z^ S�sg>��s�k��Lgv7��	�ܶ�=��ۢ;�Rm�Vv��~���C:���ͪ��y��;�٭����]C}�Oǈ:����(�@�9�Õ���"&��~ɽ	�!�>=6d�{>���HP���$Vʌ��ԑuX��@y(}�d�p�|�5���H����Re����*ЀU���(1TIX��-N�B�P�Y~*Y���Y�vK��K���_��,m%�s�Q�0��~�s������+L�����!�A��,�kn����.���2U%�U�lc��xQ����Z�0a���v��\QQ��=s��,�+�~��1t`�X(N��
_���.���(�b������������Ŵ뒱��ɿY��2�G��qCh,h�a���;����8R6��N����7��9��5_p�܆�X�W���IUO�Es`�G�7b�W����fУ��>��\<@W��P�Z|�]�ր!6��eiQ���F�@,� 0+ �����6.�1MOsQS��o;g�W?�aƏ'Q��g��rs@�8sȇ�3�:�ZKu�{�)ώi���$*�S��"-<�{��`�A�h����d�>��k�s�iТ]��6��w|���)�#]�e'�Q.���.�?' v��/Oˎh��G��@�,�
�{S����L�`p���o����B�����fź>�V������H�ۿ|	��m���be�f-���4�@ƹ	�AL�d=Zx��
ڮ5�[���c�U�d���:I����P�7;D�RkӢ��ܷS� ��|���=�� ��]�A������o���a�Phh;�`UM�=m{+��h&h�<��
��tY�=�����m�ITX�Hs�O^Ϡ��	���z+<yKNAj�F�� ��g�C�J�D�~ؐ{ ,-+B���0ܶ���`�M��k�tRE�0&,F�b�6���֮�6
�o��$T\�i`U� ��fY74,�	���Ҵ$U��ا:�Z=3��cU%���R�d��O&�A���ɕ�.~��'�W��W�(~�YQ@>�.�����f���3/R�"�-gH �E`"���M<1V<�)�&�p[��t��׬E��1�s��s��v<�s%�3a�97e!�}�z#a��q�a��8~�p}K��	?�Hn<��f�����DD�d2/������).@��R=G*���eZ��QF���}�І%Z���}���M�*>����������ߥ�|�)ø�� yx�b�0]�'�{��Жq,a���5�5vk'��GH�S�j�G�rԇ���b0�xR�y��a�ynP�PG��|R'��#+H��ݤ�{�T�?ϕ�#GB�[sLR��m+Uf�����^��h���Ǒ��g�:���㔈�4��b���wK����~�7�v<��B����F��o�zg4�Y9��s|19�2�a4⭘o,�,A���8�@K>%��:����� ���ۙ5�����ѳ�x�k �>$��
�p]�B�`l>�{�i������|Wa��wN�"����1T~��(9ϸ+����8�9�V���U�˲�=Y�
����������	l��l�P������z���A��hi䄋0����z�\�s�
�(�l�E�m�d�g�׽��'���F��9� ������fY��Rr'�D�d��@a֏}��������k(Ss^5d��I���jn��V����'0����@�<+=̢y��M�����-/L1�;[�.Kye�S�~�g������GzF�[F̮bQ'�����Ȟ����hT^�,�۰�^d���S�o.��49pwGf���M�c��.SZ����ۈ�l,�>�_\�9da�8���~����Iu�(�)oEܸ ��;�O Z.`��,hs�y��c��-֫/�U�{�o�ę�:����aP�s��ݸ�`�|�E�5�	S��E�5r"INC)5���o���f2��
��e�|`h�X嵆�ĉ�Anq T���_4�Ӽ-�R��+�=�e9R!]�z�B��L,`���!���|42j�C�%���H܍��tUjwM��(f�C��~GA�X�є��K��>�p����}�+��MY� ��a��$���6� *	����4 F�R��m��l���%�l�EI&�E�,ޑ	�6D�l�CX����j뤷3g�:�u��(��,��'��8���ϐ���4��V^'bk�)m���I�^�%;bW�s�ao��-�L+4�I��D�T�dB�(����3��3!q�?$��޴?��1GP���̱>.o�4�n&�E���g�v�X,�_�լ�Y�(����)Z����]H^j��}f{'ȣ�F���G�8ȩ��#Z��7?�h-��ҝ��3B=C��M)�ð�{��PNT �L!�WȨ�:c�u�&�;��=���E���]��ܪm��t��T�8�;|1?�:����r;�\�o�d���^�D�|��n\���.�l̹����ޓ��7�|P�{��ԋ9S���B.k�wY�!,=£
������w8W��}C7�;���v�Lލ\�-�J�L��et&����UL�lh����H�`T�h�M7��n2�2M�M��0���1!t"�O����h�hu��-!����h4��el�J�Ǻ�`�P�IVwPf�Y-��&y��1���C������%�-����7M�w�B~�e����t��#�{6毽�d�[�T�������̢)�%񯔑���t�)²\�jȇzr����W5�8å�g��y�?8�"�!oWa#��v��T�u��U���)��A�"C�����˭ߗ��a�?����-��ȹ����Ҁ�E1�gj 1���	��R�7�rUB����Tu{T�m�	Q��8����@�#i5I:�1=���ߍ���~�4���@"~���+�	M:r��R��6l��r��֧��@Ԡ{��ۦ^�w+��7��׀�/5ا�J�PE��V~Cd[r+�t1�P҈FO�^=aZv�e�i�53L�5��)�Z|��#8넡�[P~�����N�E�WA&�ր�2!���;c�kEWD�ӡZ ��Ԭ����^���'�;�O��O����\I�N�1~��qMpuC������[	r@Y9_�U�K^;v�Y�]M�@���W�oA��KI��կ���\��*��O��n���_ ;�C6����z�����U�jL��Ǆ~�;��5j,3��{��������]��޾�;��WƋ������%,�T�ۻ�f�_�8Ş$Dv���>
�����E@r^�$ō)
��
�^�׆
p�rf<"�䭴�v��@muᤝ�%��V��5�(�P��|����-��w��{�tRIPnspZ����p��_(+ɱg`����Q�k�[&�+
�a�j8�,�-����E���b���lh�ȧ��,�����Cw����@bsy�?��n{}:��e��^!5�R}���\To �G���Y32����t��"�W��ɶHrI�)�/j�����|V�k�Dr��2����f��u�-I�۪�����|��Ff���v	�$�E}�+$��z�$7{���mٛv�[���{��Q��͉g�ۓk�%�t�E|�Jl%���)��ִ]~	 H%�>&��_���(d��ꞌ�h8��x���F��,!0J��:h�.�[��
�Z�u��6b����nPhG#l�*��xn��`Q}j�������P?V?R��ӟ����4��H����`]���-�Q$r�ή�B�&�����Q��A�J�Z��ÈLm�^�.螒t����N�Q��k�5Ҏ��O<��\���pm����u^�������;1Y�U��+m�ՄpF!H����&�����3�Ңj�g�]��C�s��,p�q�)�2�E�x��ι9�d�n�x)����~h6>?w2�27� �NG+g܉*����H�j�	b|=r$.=���j��z���yRA�+���]�Ke�7;�P�R(X�Iѵ*��c8���Z
|E��n�o��&�o�t�Tw')�2NuV����Z��!s�L�}ϸU[O_�}��E҅X��\
��6�b,h���^�Sr�=&��/4[��w��V�n�=�Hbe<�ݩ�v(m�䨽Ø��qk�h�j��Z�n�_�KD�Ek�)�R*}#���[8Y�2 T�UB�S�|&
G��[�a����fo|qD,2P����1���^�8e&wIl��#����y��ؾ��B��?M���d�.��:�9���v�n�?�d�v���mΎ��1S���nP�9Ųj��SޒK��hQ?�=q�V*�u�W����{Xd�����:g�,�U�\��c���0о�g+�_o^'�"����Ku�v����+�,����<�ٹ���.x�y]�P��]Q�W`��m����)g�I�G��9usԯ�Z\�	P�D+��$�������9]��Rϱ ˾F�$�ۂ��I�r��m���^R������Ԝy��	D���z��u-���ʅ_��Φt�hwWAyc�oe-���ZT��G�q(�T�����+�����)�%��uwia��|�J�|�z��v�(7	�c�[���d��Ʀ���+R���ۯC�?	���#�K�������ÑQ��2�Љůj�;�N`��f,�sx�г�8"q��E��C9>��P�(���(LS�D:;v���F�[d8��'�ݵf��i�Y�<�j��8�GF���:�P����U��Zk�g[�Nњ�J ;��]���#�W��`h�r+|ج-)胳���֣f��(�.eڃ�)9����P�����I�B�_ ���P��,�� j����r_|�Π��zbY��W+o�D4�\}B�x���m�Y�-���F�����y6�:��������}܁�0!��NԳ��F���u:��5>.p��M��{�J �)(�Ǔ��A���ҿێW��*���
�����XJW�+^K���=��)H�p�td�}[�:Z�$�S���K��]	|�l-İ���T���� ��t�d.��K�7��K�K� �ieś�`\����N3O�g��M7R�Y�wL#l�4x���q�$�ɲ��gedlrBq���AN�%�_7)'+��*S�k�2G
�X� w�3U7m�@�4��,�����ɣ_��}椃�g�]+�/�#�&�+�m�
�P�磖B*����j.+��a��"-Q����|��9��[�)'�ʞ>qv�-�/F����nðr��j(���WsV���Tb.�dD�תz,��JG�m̔Q�6O���%�J�o����OH�ey��P�(0"�H���Xu1�W�de�¹�M�]�[���n?O%�JG�E�sJk4���0N��u�^���l�y�Uk}w)ۑ�� ������w+8���~����Qa�P�&J2qA�k�� ��&�堯D�-r���������Q��#p-�˫���ގhe��ݛR��'ߩ�j_�K�M��i����=[��)����Ȃ�C���|d���z&9�{I�ڪ ��z���1��z�T���N�H��o�tx��OK�v߀�ڦr�o�E땂����T����V����Ɗ��k��cD������+�G�>�n�VDR�]��J'�>Ci�x����=.h����[�����,
��{����4�
�B���pK�S�K�g�Z�wR'�yK��gu�3i�w�<��*$�� ჺM
�>�ñA�覉��w{D�!&�J���'v�1Ĳ������7�B��t.�eZ�[�W���\��E{D�4��7`|���i�p�Gb�z�[�S3�/�-j[tM]b�[�z1u����������y��3��u��_�o0��=��S�amc�ӟ�{�����Ϊ`��P�G�����
V�CE���lF2��⌐b��cq�_���%�y��GC��B��}���4�5�M� ��e|tn|L���rx��HB�ΐ+18��[ʑ_���	@�D�E��:�ͩ���{��g�L%��`"[|Eh��NS�nt����67��M\S�T6�n�tk"�8?�K\{��pb��"��R{=�?�  �%U��w3��|U��&X� �	���U!�C@D����
�08Kd	�|w#�S����|��h�h���p,�bq�"��xK3#n���|)�p<�|�p��?�ͼ6\�-0VfX~��9�7-�[,��t��%q���'I�Z�5_{x��lfa"@><���ԝ��Q;�V7,�\�V���68��+6N��!ؕ ��;B���<����<=r`��ӽ����d�
:��p^�ּh����bS���K���0y���|N�It`+�����K���O�R!�qΨ�N.�6�p�3��Y���&���B?�_��_0�$�N"�*�����u��½���꯶4��^�}ع$0�.���l�ki�+�5�x3�ԢUt����6Ҭ9M0pc�D�{7���b�,Z��m�y��D���8��v(��D��@>�7�?��Ջ��tŝF[^�y��μ���N6�E=@y�lr�����?��ڭseI�݅��4����H��M������a�Y+x_%���lkUs��9�\"�oI��k݉�^����/j_��ĺ�d%��m�.-!	�Ė�֌�TG�/���ut'~��	f�?�H�w$�Z����nnm�
Ƞm��J ԟ@Уs���R��D�?��j��4#�0W�Iڈ,|�+��j^T��ߋ���)�M/�:���n�(�"B�~��sQ�Vd_��2���9� �G����f��mm�'�Tdq�-�]�ǻ�p�Sp&�[�i�9J���.6�7�bT	� .�co*@ԟ��t�b8V�n忤l'd��W�F�$�kv?����у����Ջ��b�A�au^��?����S�q̵5��R�ua�^D�\
�[�8�d���p�w%���%�W��8��8��1|���~��`:����"�D�5	��e��X�!�I"1��H
�m"ܷ���u.��í�-J��ͅ�|�9��~�=�A�f6��a��R(�Ns���/�KO#X��:y�Ҡ��1���7f�^�=_��SE���N�����-\��]MHG,�fI���뒶1>^�X]��1$�f�p�۵#��/�P�<���R .�}���S�������G��5�Z�����~R��C���?)Az�i�e5����\�^2^q��d̨!v��'p�.�Z<֑ya�(r�^rM?7Mf�n��]�N��t���Vc��!c)"�m/R3pI�d1�Wu��c���������m��B!�i�[��B:�ዥ�l�To�*��7-
|��Q����
C6n A��H��{'f߰[_M��<A�� yk���0�����GM	��4�FwO%��K��<�>Xq���Z&��H���4�W3vJ\��`��hMh`�3�4��3�>#O	��^�Oþ��r������	���ֱ7p�RF��dBcx��z�}�0�)@'��B��W"���R3
�m��CH���%�ȴ����3��x56���Ϸ��\{w8����"zu����KѾ�O��mp�����V�u��c�jH�wV�T�4�8b�F����z�����C��{�=荪���o�A��2`a�{{�Kt���[��1�y�1���5Ĭ�3����<&��a�L���g�y:��TΥ��E��Tg����7J��P���R+2��4�h�ڃy/r�=�i,��L8��[ݥ�J�dQ�j�%�ד0��蚞����J��tP�$��/fJ�8�O��RjEQ�`,i�_�C��BF^]ܾ�C�����l�C ��Dx�f��^F"+@�z��Ƃ��GU{TE���T�/�}�R�F�h���W�R��Ǒ�|(���(�њW,!������N��2�{|F
�9V'��cbc��q��=��R^l���]_kؑ���J�C��£�GIM��� �s�)�@�խ-��(z�Е��e��Y�fSLO�M~:�\u��Ґ"MY�M���d��p*�*�q�g��H�`��Yj�1{�oh.`�L���2���fi�yy���C����r>';�fȇ}.��i"��Er�����p��#g��J�N|�t���n��q4�M��]�͹�].�P|����ڏ:S�
,�Q^>��H/����k�h�M�!RY˵�ru`Z�W��|���O��Nt4PI�L���4�>ꍔ��Iگ�s,f����|���?0�V�� ����"�"ɱ��ގ9��Je~;����OI�$� ��>WuSti��!@�\q����C�׻Q[pQ�ԣ����gk�.��-�L~Z����\�7K�-�mp��Os��-�������`|�c�NO��D�� �mP.�����G\��wy�����9��{���w��N��ݵ;N���q�ї\�� �fL����̣:٥�J�������I��z\�B�(c�[��׳�<�V�¬e�\2���@��@ܓ��ڤ.P`htɧ�7'����blj����	�|�8�M>7SITc����t�x��%e��A�q݁��%��C�ԕ�,MU�D���K��t�p�4e_I�$ĘP��;L���C�n��ÿI�8 ��a�R0�q�vxϖ���u�#�h�Iн���٦F�4�D��4��r����Tn*�Ad�+���߅��=0�}ޖ��]ɿR-`�>?
X����
�D�N�)� ~@��럄��:Mm�[U��sqC��gHҶ�UJ�r\ѱ��l�BR�P!M>�₺���TO�9*4�a��r�����ɻ�)A种[����Ɔ�1���N���G<�s�H'Yw���j��҉��%�_q�-,E6������P��+���/��*�e�~�Jn�eKҿv!{������X��_N|sT��IÃc�=�I�M�/�!����=9��\Q��I N.��="�h����=��I.[u�et�;L7�9�)
+�GP�Xk��NV�J�ڥ��|I�`�6߀O{���U^�dO�Q��O.B׳<�Ӆ%n�h綋1��ù[Pe7��[���^Q��4
Tq^� ܠO�9�\?k��at(�{���9��w.�a9G�ٽB��7�XmI��4nX[ ; ����N��NYZX�"��ᰇN���T^����>�Z���W�pq�g��	V��!��Q����������x��x$�������@7�3}OGM|�O�Ѽ��[*�"�r����i~5�&�7�ޝ�x�u�����!�ʌC�m~���! �z���c��P�����ba�m/[ܗ#���櫾�����bg���̧7%HD5�נ�<B|�{�:҃�tHa���X��C�e=��S\�mc8�c�`i�N΋�T�G8���TkO�HJ�e��狙y`�����<:M����f���W�0~N�N{S[]�O�Y��o�{s�$v]�"�`�I��O��ZU� ��q*��`��ds-�p��X�%��<��O>�縵�o�zJ�3�X;�����i���>j����R���j���0}��x�1�:v7�M#}�'��b��-���(?1Z���H������%��'�A��}�h�ChbS���l���&�]��1<���n��G�s4��
@��o!qK-V#.#��|�ĵ}�[�D$�O��N��D~��䵿�.3��Z&�m�9=1�$��>���Q\�����g!�o����o�ȥ������z�U�W����]��f�v�㮖�xY�s�u�9�
=�Ob���)��8ܠYC]�oG�z:�龏��M@�e��z�C�{V9!Ơ;9T����N�՜�$���-c���C�������4[7��C)7��n��m�6b��i�	9ʍ6J3���kP�w�٬M� y*5�2ע2��k�N����V�?D��_lM�y�O׵��;<Y��<����\�0 |��U��iL��#u
ūm�J�[D3We�e�,�9-.��9�� �Y������qѫ�h4�K#W|��ӼG�	��7�uK� kϱ�2v(S���㟅���քZ4��$�ּ�˚�.�s�j ,b�cg\��2�>���b'��*��.�����k; ���{;����A��'0�%�	�|8�"v�d���J�D�/3�l��C��BAś)@?s�M�^s�PT��f�+��M��%7n]�\��~e耳H�6��ފ��@��|�C��T���\�WD�8���v�����k���i� m�R=���$�H��O}h=7NrB���I�	Os�x��$GCZm,%#w=L8��H�c���H=\F�ћ�$	��JTBfq����o'�a�>����q��z�!�(�'�.�i��>u��IR��~a��]���B,���$�0�S��έ	}�j�*\���%�?���V��'�1K��pD۩#�j�.�tS!���H�FdkB���*����+�p��rഭ�)�g�)�x�6e]���D�C%LcE�`�D����"*��־%��S ~�,8\C�֚0f��fMZ��<>P|��,Rl���*�2T������sx>�=H�%1-{kOXn� ��GU��5��=W�b����X$�W����)�\�^���o&'�Ƚ�:��i��v���yQ�ʞ]	ɠ:������F%�����|�N
%᷿we4��3@.Vr��y�JU�K�eTUBM��E\����Jy־�J8�&~������I��4-ȝ�^m��ޤ��Gg�\
����(MN����t�H�L0�w}2x2���܄Ol�8V���	�� �|��Dg=��� �!�>����?��9U ��1����*p>�5��Nv�he�$E[�n�w�w{Al+4}����1U��a޸`Ӽ���q�J�ߖ����#� h7Ԫ�Ο{���Ş�@3I������At��hO9n��v��N�},[���)��)&�͞�i/�iu�څ,'������-���Dc�"й�L�8}��W��}C�4�j�s;�mY��'-7	Y蒏���dO�_����+��4$@��e3Q������f;в7�M�SÄ~���)3�<Vkl�z����0�{*�Y,�t��"GsvvJ���tZ:q��)w ���3:��,9�YҤN[����CP���2֊]�0.1t<���8�;r��TE�>��_�Z�]\i�e@��Ϲ��Z�h����`��ĕE[����' |����%J<I����C�I�/|�k��}D#�-!�[p�.:�?�ub�f�P���|/���Ju2��qD����kH���I�śp�Uu}��������!�9y�[� 3v���Nq�(���z�S�2 �£�����D���"��N \�6�O�9��qqMʕOa�f�(@��W����3�Tqm��[����W���hY�c9��C����C�6��d�J]�B|�YH�F������Z�P���X2�a�*������c+-^Tuߴ�|��	���#�|,���!�ZW��:Ȑ�{�e�(k98�F��h��3������M�Ѯxd�� ������u�u��"�ާK�ʉ	��=dXa�8Xa4�~��8x�O'G6�����h�5���f2:R,�ԥlO�>�')X��&�Yk杣�ߝ�}u����=z4I@��( �dH���+yh9g���萓 ��:��.�/�7ix��h�9͘|�4�Z`���P�-�y#��φQ���B䄀,A�N�SV���w[����я�r�ߺY2n�:����^Ǚ� -�����,:p׫�	���!�(����4ۍ�`�0�%��tra�p��d��)[mPW_ ���7��ڲ�2z��PU�m�ݥ	D����{��t������3�H�-<�}���d�������>��p�2�9֠U�����v�#�}����C�_G�8mx[8R�0XS��?�W�� ��łiV,i^R\�	8F~�6x�P|q�[��~�錧�����۲�#>I��X�jS\���!���U�]�MH�CSo.#�Mu�9����bXKjk��9�Z�4b�w仩�a5�)�j�%�P҅�ac��pUs��C˳:v#�sn9a�V)�L;�;��pPr�P�KĴk�P�ϛ��w�縺Y��'_��g�г>��0��޵�1���_x����P��������s��Q�Fڵg�x��`ɂ`�ѱz��T�@̎]�nw'&�<'zW�������̜a��������壪�|X:��0�<�e�Sφj �~ �������p����к��m	%q/|z�ý�^�R�'�U��pČS5�[����sO<�ըbH,�΁rK�-�뤠 ��ŀ��+W�Ł�4�`Rjāp*�BE�6�
Q�@�ȍ�X`m��e��2�44��*7֦� T��i{Z�D��Zl��D����zQ����ޝ��q�q�5���µ��Z��*e�֘|�Tbx��`|jOp�$�������h}Mk?r��6�7\]�o]� A�m�g������bcQ�X��s���?X������ʐ��+d6��p�i����g�m�2���?��ɠ�8Ln�� �Y�mX���&���G������c�	4�����X����1s���9'O��`� 칿�PgI`ۭ�	�V1!�8X^ˋƍ���/h�~���$0�)�΀y�V"'�&�'U�1���#{�FK�>����{x=���'�Z��_`���-8�Rd�KT����6���&8#����c�;'7뵔�@�����re�%h%�D��.���ciG��oI�
�1^{� �,C�Xc������x:̖�����?� f�#����`�ϻO�s��͕h���T�p�{&-vΰ},��.�=ݲuiO�b\�)���}M4ehTתx���i�U��aX�k�u!�5��`��?�r9�Ync'i"��邯4�4�%B��>�uR�#_��T�'\�5��,�?c7T�1��X��	�aɽ��F�a���ꈟ�/w����^ts�ގ4:b�ڠ"^&���ՙ�����X&��bRQ���E�"H ���Dh�	e�p�-��JZ��C*g,F�
0@��ij������Z���yן���@!Z����q]��:��<��*�j84�Ko����vrETF���U�pI?�$Ԫ$"��	i��Ja[$X7k{�t�߿�V�>�?��jh\���
������ix�ϕI`vH}b��&���c���ab3'��V�uvPY�^9�AA�c���0$�vT�ꘂJ�5� �j?h�kt�pz=�ؗĉ�m�Z�x�v�)x�b��f�*�B
�Ϸ,�}�P���1*�lV5l�Aꬨ�h���9д_@�&K��f�B�ט^����ͦ0�HX��BB�*'a�����v��^�v�9�gBr�azh�Y@~l.��I��=���A��D�r^�	b�\�U�x�]��$"�/5���{Id�A���6t'.K4��L�=,q?��4�ʹ!��Һ�^t���=�v'.��hr�?�_�%ޔW��s�P\��}��
B�Բa��%l�5�ϥa��T'.��"�g��̝Ѓ9)F�o:���x������Qѱ��tUTWª,�,!o;�R��Ǖ]5Y[�;M�(�X՟��ysP3B5���]�!�B���*���9vt�{CP�<V&�UiV;өB�|oF���}ƬX���)��TE���
�o)�*��s��+�n��R#�Y�O��A�vE޽r0=�*�MW�A/K��7��YPz�x����e������b?]ӹ�n����@1�����=P�k���[-/C��=8�_@{$�ϋ5���r����J���b�q�҈."�$��a�7r%�W<�z����ٙ����(�ǒ�x;�*Qf���i��	xT�8W?��+ף����`�#�0�k�l"���V�V�8������&*��MpX(�s�10�t�)�X�LG��6IҮ�TQ�VF) �]��1Vs+��ޔ��m�Y��im����A\#���@��7�jI��'��v�	&��"|&��۸�J��o)�5*���l��#��!<ȟ`-��Gy�N�Cw���,`��5�껗P[ͺ=N��T�=�;��%���F��!#}x�[U����	�!Z�-/��`2#��5��5�^+ژ�q]-�XP�i��S��n���Y+�5�k5�E��!,"(DOV���l}��9v*f�OX8��O�D��v߳�[[
M��9��
�i^��y@�"�ur���}7�����41
�DJ��^����Zv���wp��Ci"������s��1a7���뮨�ϕ.�	B�k\��[�:ȁk���&A�߀H��z�����^�v�.�zM�AV�z����W\���kGc��'gl|a���/R�]��u�$��}j^�"�1[��JNfq!�!J=�R��p �}S���m��\1<p����aR��a�X���ޤIb[R���Ӓ��Q�AEiBr��"pT����=��t��d������gk$����js^�OI	N�n��( k��xo�͹���6u���~f�K;�;<�}�NL�V����Mu�]��B�{�=���:�}�f�C?2�n��b,@�W!PF�{pJ�#8�P����&
�&kh��ѵb�)�M�!0�����ۂ���nQіM��8x �Z����>'���L���u�I�8�Eu���6ʰ�V�c6������T���"��̳ut2�=X�:�ô��㣺���e�n�^�)�<x��l4(TQFE=�g� ta�����9q�$7�k�u��+�D����E�4E�V�ة�sS@b������-(#���"t�V}��v߳(�X�svu�#3l���� e�W�T!��c8qb�����F覣�V�Zd�\��C��=dI�؀,U͍�_�j��ۏ��\�-φ�t���l[+{�o��u��3R6��TP
�h{]�i����A����wQ�кN.H�����(��ɮ{&2�R,���`�ǘ�UXO���~��7?�_�����!�_�=4�� {�]�Ns�N�����~T�<?���p�r9�O�5N�b\��<���8I��Xr_�tN��5t`�Ӧ�RK��"Q@Ϧ��h�I�N�(
V4栾��)�1���a����ˑM��<�"��a��i�Ͼ��Aύ&T1���F����NƉ��bh�##OƉ��C�bgBM��LƓ���Ka���4�P�"!��l��g�~��2����3���)��4����pi��~0�"��N��	7�M��TѤ�4���;�AD�� �cx�n����_��m㳲�#8�,�`M��ͬ�-b~3��X\")�k!���>�#�����7��+�4��"ȅ��V�9�U�#�KQ�gN�_0�ە����m�ع\�#q�e�:N�����B�t*K�IIZ��{�TVB����7K�f�[F`�چ�Є�<d{�s��iʹ��4�LL&Gk�G���r{Ix>��]�:��?���(�XZ{�UE��m��<:+��������a�,�X�+�HL�T�`�2o���b�?nKkb5����_�f!t�D��z�i�W�r��D�ӂ�_x� ��b�.\��r1%ҍcu4PK0o����ҍ��o[(�ܬv�V���(b4P&��WVR4 r��7�&u�ޤ�/�����t��@g�������K��>�{��p>峁a�\=���(��j6�u�b!B����Q�?�r�A��\T7�4Ri �k��q&�0q�{�^��T�<N�t,, ό5�?�C� gB����1e���s�)G!q|})����<���W|U��[r�9DP4��\wIh��vB"��>�?<����C A{�B��G�z^����C� z{jT���`��i@|>*�� ��]���kOK�G��f��=��j��}�Y�찺�ԝ�j�8�+���+hHc�L�a��Jg\��ҪX,�8L�e��oǷ;�����yϰd֨�C�Ხ�'d�k4U�;�V�H\��&���G�a}���0��� Q!�:d;��{V��������������-�0�@X*��nx�����.�Q���.)Ue�D��
n,$)����v҄�Jk������dOB�:�'���;��ΐ��5�����	���b>Ԕ.�#��,���remP�K%L_��-HE7����$�2�&��HR*`Y�_T�a_���T7�,Kvc��e�m:�"��E���%m��%��ZY�nI\5	ʉ6@��w�������*<��36�$��b�y|x&��j��JV+C���w��������%�B`�]^X��^g�l�+o��a��ߵ��-5+��~��&e��溲�֔m7s�A�a
�϶'{�ڗ�'��&�K_����_���XER�ӵ���8\8�M %ʺ�XH�!bȶII�d��"�4�e��S^�J�ĸ�Zב~x���Q~�z����MS��:x�Fw.b�L<
R�_jp�ByP1w�W��vΞ`�]lhMd+����w�+:�WCC�j��ex��� ���]���X�P$N>�Lbdv?NL�le�g=M�q���`�C��L\Cn첄odn�طkч��	�ҡ;O�I�Ǩ)����N3陸��u_I��>4���&\ U��I��v�S^i2�A��\�@$�V���uP>��וr��-ٲk����Ӣ/��0����9L�����#7O����?���&P;��:���=����y�t���tlPbl�ѽz�Z\}�؁y;�`�>�L�HT,Q�
C�������-f��K�F��4�0b��I�a�j�T��3���m߶@�W��A(
�b-�G��B��@änr6mE~y��vÚ����%�u�Q���q��e���:pt�DՊ�.:���:h��#��Y�^o�d`�nZ=)閟���,�D���z�sVz0dT�]`S?�z��&J �O���'�K�.>[�VQ��(�
���Ѯ�h�F�@`0N'Kfn;z��i�{$*����o�>�[9�)��g�I�x��z��c�y?^����O� �uN����h_��)�.�Y�>n��wqkG�pJ)����$�<-.���6��'�|'MS�e:5��)r�nx��_��0�42E���"cġ����dL�p�|��_"�ֆ�q�?jÌxE���_	^�TU��~�
���s}�[g��^�L1��"�R���v�yG��o4&��h���v����$�r����Z��xZP��<�輰�p�{{�>h}l��n((L���1#f�n��n�>������M ���N++e��N���R�l��-d�~��8�~����ulm=v�n7��:7t0�µ)wU�<��A��؈}t��HӍ�H�=��
_NC�@_��<�j��e8���8����F�V�\G�Uꘅ�f���N9�h�lZ�x�=���p��G��?��pf}4U�Bʯ�t(�w'�̬Z9l~T�ab$$���)T���c���c�S��ʚ�����3��n�'&�����<qO�/���p^����Ǣ���3,��|$꾩��g��6��ޱZ�m���L�������1PL����v��#+�X��ր>�n��ު7�%�3�tN�}а��T��$\�n0S�F��w��fI�8��'6�?�9��v�5p���pX�ҠO�r,�G��K�}Λ�@Kgz_������9�J�)�CJB|O��`�Ʉtם5y�ϐn�/z�s�'{l�*䵽�{-A�4�~���.,5���ՈVy*j���̾�}`R�~���5D{�6~y��']D]|X���AUEUq)�E�V�8�r1G�3��/���'8��K����>�,3�%��T'��~����ŴIh�WI.|'����2��J��ƞ��R�E͂f�A�E[��9��2��ĜlKԇ�Q�E|BM�s��J��(#_q�ݭP7��p �.�y��B�a{Րa��=]\�~�T���\������@u�蕪��4���Ѭ�O��q����_��7ٻ�ޯ�4�A#?/9�]��@R4�i�=��]��e@ֱ�9ֵ��fK0�v#*��*��$�9���[+����qn`a��α�-ͼ�6�rM5pjz斸JF{q��+R~FMU�Cp��]I`�-��M=jz�ˍ�0�+�\�����h&&=4�α�M�L�(��D=�)T��.���v1ڟW&*Qx��((,{m�1�����B����|�!�IY�YE�sEsS�m�����w[�˭F5�6��8���ƣ��҄���+b*�
���ԁ��;���� �@�c,���j��&�P�ό�N]�\r���`�
0�(�3>0���i'?b2�&�C��dĉ�*�0Uj��:��6؟�ɛ
�Kpx�����΁ך�U�b����1n����=��H��1�k�H�ܭ�)�a�7T��m��BhV(��	���u�0���Ś���΄]��TU<���5k#�C0�=-C�=��;ɣ��|�0���.��*oj��k��ƞʢm6I��3;x/1�����s#
��~���!U��D����U?Rҏ��^JTyggly<�txǪ_p�R���v��ޫʸ�D31w��&�P*�;��cc�9�>p�`��{%���M��Tkц�������	�q'��f��x�=��uw�2�����jl������Պ��`n�m,t����W���YO%���൏4b��+wQ�6�nLivQ�įd��ԕ��#R�.A��h��N�8b
ߞ[�s����e���F��P)����I��
E�$Ɔe�}v>��'�n������Ǽ.�:ٻ�ܥ�L]�/�c���/�'˒2r�S��V#+�b���l�����g���\2�5�Ȫ@��W�f��^��:�������_���n�B��$�>�@eM'Ξ���]����Ka�V�y����4�0��N(����{M�Xe����]�)���ч<j�h������7��R�K�dA����#����o� Ŀo�0L��4hofxme.�L1�Ј����t�[]0-O���"&�Pɍ0�w��E��aɸ�u��n����=���d��3ⷐ!s���\�I<e���|m��N�?.=�˩N%�hϽ+_Ek��+��q��4K��������,B괗�?;~�Ha��qM�T�`&o�^�wq�.��c�w?��E]7�}&�J�f�`�M��鰅�j��aS���z*uo\��=n��^�e
��!�>�������t�����gP���t�7%��۽�8���i�W����W�4�j�ղ �Ĵh�*��<<���$������'���"@j�R�v���d�Bxh /�\"t���_^I0gU��@O���g*2Ԇ^c	r��5_�6>u��VI�)��f���(H��ػ��߶�M�T��T��9�V��ӄIo,&�gŀM+�*yQ��c�՞�ޅJ��-
��6����`%��@4T?�p_7]��۫�p�S�ᮠ���.�|t,�)�IQ�.�qb�jrc��O�B:�߳������8���;�EF?W��JFFg��h�b^r!��d������V�R^����h&���6��LŐ�N���! X6�~�����f��w���n��'k N��w~�@�RsO�n-w��� �b-l��3��65�6n9P'3l�y��L�;>ϛ��B�$��Y�����g��o1�5��сj�|�`�QL�n̐EB�F\'�{B% �DGL7�
ɤ=w��������ڜY8C�%�?C�诜�AK���x����d^T?�����Lw�L���Xʞ(�lTpH�|;�l�K+C,N��D�kKo��-&��ŏ-����Fª���(��\ǆE�O1B�L�]��N�5� ���Q�����>Z�BYfpj���A/�D+�3X$�J��ʖ&��
s�f���/�s��x-��"��Q�VKHcVe� o4tK�
���#�,��)"t����!��hJ�������IG�`&k�ߘ `��V�L�"mXP�����ؐ���8��G��	�;,��[uV
��?B񓳆<�/���YC�l��$��8.z�O�>��)�v�����%ͣj,W��sw����0r��i�P�C�q�E�F��r/9���N�d�ފ���I��?��5��!�z�B���#C`�U�QI�<��Wf�	^�ْ��C�ݍ����R�ϒ�!�\0�?��?A��憊v񮩀�[g�~!�lH��d�dC�R���g51VVR��`첳etM!ա��y��Ҩ��n��)��Kn���;=sjb{ݨݸ����L1�S[3D�K����ć��"�e��=쥤������8,�ͳ��֤�=���,�����h5��pˊ��-.%Ĭ|�����ϳ+_�z*Z+;�r>%���r!n|�^3X�X����B�*Z�쁑���7��?Kno؉�����nl�OOW��j�&��&O������t��߲�˨`��*�8���i*��_���n�{t��}sn���Z����^��^�#ӹb�K���M��Z��.��zJ�=��戚NZ�Y��:�S��L��p���@=/q�╽�o�L��O��@��vE�3z^���߸�a�䧣���/�ħ�qt��W5W��_�jRܚ5�L��BV�Z�zOv
zv�ti��ϱ����� ���b]|��^J�,V�C�4E��L.�Иf�-��3����fZ�>r�@��)�Q}P���k��ߗՀf1۵;)��m��곶q,�O��h�dp�)�Y���+_��z�YR�9��"��-��c��ec��gK%�)�X��o����]��>��'D�.��޶�ӶO���O����:��t8i3�]U�ތ돱��P��#z��M�q<7"KW�q�Bv��W��K̓��f�fv�H�)�ep�k"��u�{rvv"S-�����%�0{�$*(ۣƪ���MA%��jT��R����b��p��$4;S}��򎯸V5l��BX�9�u�eQÃf'���ȡ#�Mj�)�l�L�C#����sF��FmyPu�)�O�}���3��!�i�ә@��i�M�7%<��H��6�~����c������31�:vh
xF�4&b�;�U�]�W�{�U��ǵ�ʽV�P�G�Her����T�e��g�e�O���͡��Rg4��렧��3Y�tq�
�@f��s�oju� �vΠ��!oN��`�rN�\���.aqA����Cy�&	��"����y'J���o-w�
+͜��E�ɧ�s�]�B0H*��Yr��rr����U�oy	�l0��O���lp>��ވ��yȥn�sF���Rq�v,�'s{.s��ﮭ#*ф�~!)xw�<O��`g��D�&����L!:D~/2U�&�{Q�]�Q�`�������g|�D\�%)�L�_ǝ)9c��3��1+;P#Vi^�7?!�gv���r"yϟVN��Le'�e}C���Xo��2io��N��`s�?e�w�(̊�@ ���d�-�B/t�%��P'5�/W��z)(s���Ģ>X7%ϒR2���ˢ�G�RX�Я��oF��ђ�����ܚNh���+ZTP��c��R'�0p�foس��UWI�� J�l�dl$��և�#8�(`�b�3G~�*��?[�$��C��b�|��R�����_��'����`�������\���q�N3}t����"��Nb�|#�k�	hc���n+�pb�|�&�P�A�}����Y��Ȇk�*G=��\|i�=gx̂�.���ۇ�)��L��1I_�mW�`j�W��0pT��r�6���OowF��eJ9
g^Q�.���8��ـP7�����*� �}f�?��$����IvA~/�j��S��\Y�y� xS���0�O-�Ͽ�KU�^\?�`�oX�_�r�)@�����\����
4_�R_�(����A<�.v�*NBg���(	^�	�����[�1�5).ߎfL�cd,d��t�_��P$�x�a�|@�y�*����m}]ڥ;���=��mU����fC&R蔷�x�̍��c\/���K���k��O�h���Bh,��ܯ���W���h#�?�����x*�d�&���b-i�;���'x��!s��L��z�2��LH���B����#��}�dG������y���K���aR���ѿ8��}z�
pldc1V�:� Z8-%���[�p:p����vfb�����[�-	_�)�Í9��.���b���ͳ�@,��/��{X���s�
e�x�Ę}�Sb�q�6�1X�Pk�!� c�A����_��
6��Gem�Q����T1�*��o����� �ćW�E�#�&�7׿a$���uRU�^�]�­k]R{3�
鈽��<1O������\h�����K ��o��so�{�D���@��Y�P�2%��_��=�Ǩ�{ƨ[t���$��գpL6�l;�Q`S�q�~��.Xx��	���b�z1��)���A$,s]�(�ګ�!�'��<��+(h]��>�ܰ4�:ɈN�s������4=�[u��$@�ҫE	Y �'*��Ab)�UE�n�i;�,�5jUl����>B�0>��9�w^�8oE�6/x����$��&�4`��w��9m��ǽ6gϿ*2��/���y��Fl¦�E���/��v�e��cˣ�����u�)�(a[��a���`_�ȁ�F�����i�lT��0d�by$wC��#$�7c?��Z�����C�L��k �@�2��2��"���{�k(ǯX��6����-!m�G�^Qq����ӝ��ܻ�9ߪ5J�S@A�"�:��s0eVQG�c9�8!(����S[�Y�sv ��[��N�M��0F���].�Ҷ�����r���k)8rue�t���ZP�)3^�t4��9������a��ֻPy���n������Ư����l��z�ru������ȸ52ʰ���Őc
��C�܎�D%e�U"<��#,Z/*q�8���P�E�1�&7S��p��h6J�9���ϩd2�e�[�p���3�R��$�t���]�)�{��75��e_&Pø�Z�u�pO5���h�������c���[j2i��?-/�i��[;`jpK��e�J����T�O�	~�`CI�αΒc��wCH��ͣ�w7Z#��;z�G"�'ǰVHI�Gi��j%x�(P�:��Ư��rA��&l�y_A���n���h�����E��~�r�	̅��p�Г��̂߳gE��ԟ�An;�n I*�]��g���s�/x@��l1�<V�'�׏�z7���d���XV�$k᳭B�ǫ0�X(�	���
���X��k�=B�(�u��Q����X�e+ Z�A �k'|@�.(�ZB�]O��fy�O��3����8I�^Q�Tlt;��H����Y!��p|��IRi����22c�#Z����̡�Ҏ�X|~������it\\����K��Q�d�(�'�BmA�H6�#"{�bEf|y�$o%�rL+�Ps.$��� ��9�`-���	GtA�6��z0����e�Ԅ��$�h�N;QĢ�uI�z�Bǲ�
>�Р�[��<W��*�����CG^l��Rf	K�ZK�,^�?��GR0����4�-O\E`*Ukn�P�Wm%�r��/�H�t���#�6@x/؁�b(z��;�r�e�Ub1�4��Yz+9`{�.΀�ӷ<��i��n
3R#�6
���'�2�<��F�up�<��3
an��|�@HS݆�a��!i�w��t�J����g�W9u�
F�/��+�`\�*��zPIMNe�(��5��D�Yq�au˨�@]U(�F�n/?��*3y��J��Z���E�����_i�̨��K�=�:�J���2w����nW�c����P�Z;>�<�Y�	�`֠B�Im������mf�߱z)�J��R"B��~����Ȃf�Bٻ�},w�9�|=�������
4	.����Ѩ��cY�ϱ���G��5Vhw�ff5giBօKi�b��%(��-E��j�P�X��#M�dF�"�[W�E$*-���"&$(�Z�e�d�-�$�����q�������M�2G=gj��uM�\����k�d�0�m �g�Hg+��(c8�h�Y�$��c	1�1,�e�$��&�!K�-�c���?﫯G?��B	������|�|}ݭP't�SϓP���O�t��ծĒ�
��bφR�Ӽ�ʅ+ĵ3AA��y�R?<}��h���yՊq1� =�y)g�i��p;}Öv��[1�lܷ�"��N���$C��łn�y�'	��'đ��{��+�8�d:�������h=e�.���4~;�s�����?�e#e��v���NN�v��7
:���q.��h}��B�Й��)\�|n l�[p�,`z۴p���-n��� ,R��rt$�)$RRRN�Y.� NCV"JI�Hl�^{��,�/���Ke�<��g���3���×_�8�ho����4�t<[��o��ɁܝI����w_��������Ϙ��V��cv=�d�І��|*����&�6o��'��"��ԩ=A�ў`�~ʥ�j�>�����B���y
kitЪ�9X"G(�V$��8�W_:���_[$�ꌅ~��Q�S9քa&�>�}EGBΒG&��<)�&Շ�:��3�o� )}���z.\%�8Ye�̟��4�=aO(��䴄�;��R�b�PS���/�/������Rjǐ�b��:=�mҹ��}%:Dw��,��4.V\����y��EO��\jr�u��׼���¤�݌�o�X���g܈���|��n��"�ġ���ȋ.S��V@��vo�y�^�HN�8���,
ۇh�����	7* �˧:β��F�Ẓ?R��R{�n8���J���ܝ�M`�AJm7���!��7
]O���M�<r�?��|Y�j��u��8j����%#�V�t��tDx1�t~��	o,m�|�g���:Z�g^�(z��3�%k�[�gY�%�s���VwY���-:U4O#��N�l\h�D!]ng-.á�3翩' �]T�Z,��X[ϒ�(�ޠ�o>�D �7M;���[���K�U�p0��AP���˦�5�b#��u�����7��+�%�ݕ��h\XJ��PwGw�1���{qf�` ~|EH� ��g-�����Y��E{��꿺�n��#��a��;�u^��:ޙ��+o�s񕭪��Y���4�����pǰ���@Ң~������n��+�"*��� ��P�eH�]k�?�����-ϲ�A�\���t���e��?k�ޣ�^ԍ�2�Y�PkpZ������߿�IT�_u�Z�a�%n����~-/��)����o�'J�dV�_�fP���s*�٬�5�j36%O��,�鞶 q�?�
j�A�S�H�*�K$F���.[D<v+�H5��}+�fGZm�QQ�8Twӭ�$��q0q��UVaR��<]9�Z��W�w����LUuCz���^���$�fƂ��
�]Z��b���2�k���šl��s�p�+�Q�3��(ƞʖ�|�3�i<|Lt��J���i�Kly���ѹ<dl���4b�(��s�e+���X����<��ֿ��;�i_J�N���c髓��|�/.5�8�Kf�f���Q�<��V�}!�;��cѕGA�_Bg�x��pV����~�=*��!�4)�]�٨Wŭ<R�;�~���b��6�����L|�ؗ��;�=�S�,q��d����1��cKRɅ����B9K���$�ml�6�c�9J9��=�`����e�"[,�*{��☤C�x���l���ܝ+p�]�QЅ��%�ş�×�A2��`ү��$󣓾(`� v
�k 1Wv:������p%��L�f�r�nG>�T�9٧2�T��0�6�|ZJ���Ԭk�hU�A��4Ka�|NY�������!SC�g�Z�g0"�pi���g�?H.�lŜ,�(�{I��kd�gGSL�@��#�����-��+�����EV�s��4�s���2�X�u��c��.j�0a�Z��s��*���Ŵ����s0-��έC��¥*�/�FxF�^�/�^�X]��S�� }A��Y`����06`�p�P(�U�8N�%v�~��uj�g��hJ�vsr.u-�ll�g��__�H��d��Y�Ei�� ,�f7��6�o׏#��4�em�%urN�m|�+����s9΋u$��}Y��˻���:ڣ����=�ўM� �	�}��kب��'������߯.�qnOg�'�^�N8H���نŔ9E�׿�^���&�LC`�v����V����8Zz��uW�$�x����oS[��Σ�\�`V�1�a��'8D�����x.y���Cg�V,�Q�?g����!o��C�MK�o�^�q�6����H��'�ՌFYETR��2W�!9x�<5i\I5i[�_��#���KΒ�ӱ�*8&9�x�� +Ե�6/����MrP8���������@�v[T��$�K��+޼��ͺZY��^��y^6��	��n�Q�*?��6̼�%W(:�8 ;�U�̳�,":x�[���b��/���q]��wJa/�v�ċո���`���L�v��ƅL��yS)���C^�^*u�LsRC��j��җf��ߊ�Z9T�NN3����j'GU�Ɋ_��ֵ�ׁ9l��Π&�p?3��`"Ě̍���Z;�/_*�r_��c!����8{).��1מ�+��w���;���I݁ԗl��P���_Y5������2+��̣��C��(r�M1g	Mv��
�Sn]��z=j�j�UX����8��%�
�C�f�cX����=�ҫ��*sp�
0���,�H6G��\ð�C�O|B�0��{����4jN�.�s��,*XC�4����㱩�y�@�H޼Tׯ� ����9�|	ط�ۥ�t
$����`i���$w<[���]Z�����r���j������D���m��}��кg���t�:�N&?�L����z���<H���@H��_�R�n�'�Fݣ 7s�����s���y�)��P���{7
��a�.��i6�v�NLC�S$�����}��R��3�����D�3q&�0��C4л��n?�+�ʯ4��.C����V=tٳF�g��헫i���F6���t�멵iU���8ګ٦���ܨv���F����3�0�-^r\��0{�95��2�).�����а��)�,�)<le3H=>!��H�T+[ݽ
*,=?�B��~�K��N|�N0�~�Uk��le�g�p@�X�R�{��웺�N�[�b��1J貳[�Wki� �
��^PU����L%�.aw7N�vI�R��p��]
[$G�[����i�+�mP�K����D�O��"F�	ʊY9�31��}��p�n͛ꋤ;@���]�kR���8��qs�s2#j�YM����|��.��t�֡^��R!_7h�qA"�||�K4c K�_��G��P�!#��'8�T5l2��e88��	t 2S+�k-�99r[T��b1:���W�Wf�9��p~'w<��B*]��݄%'`x��(MA��U���2u�������A�o�����	���� X��u�R'	��F��Ly�KO*���.�RM#��Ɍ͉s��i;��
մ��ȍR��a��S���]{���	�e��c*�.���)n��tC���D�[���a�0tP!x��~8�[��G��6k�~�V������8�d�k�}`{vU�� ��y*�����wx�Y�V?�X��}�*�j��Ŗk��ͱ��"����>A�j#`��Z�jn�JF�J��mS[��

�:=uV䂦�u�$���2 ��}�p͡�N��j���Ŕ_����d:��Dp�r�&���j�+g�A��V�ơ�oA,O3^��܎R*��y�����Ck����>־L��-y��9����,�UT�;5NvZ�53�=K���>qE���_HjT:�¤�� ���rR�� ��NK�`�ߺ��)�?�|�&>�տ;�i
��>��!��ek�jA#���Ӧk��(֋.9���c�	/�¤��t_�h�����Op歸C�R�	��r}W���^gnS)9U��"%Ѫ4��ܽC[�jM�sBA�궰����ג�Mi�e4B���)͙�yUAtk�\��X��P���G�|��n�K�hCjS��Jۘ��*ɸ�O��)d}�a����땆��٘�`gtn�tA�Xߛ"ᗵ^dg�֦��Y�f�&�1T���2&w��Zw+��/9�y��#)�l�+V8����Y>ePpϕ|Nf=������:*�[�R���Z1&ƆY~6�ughq�å��g C��YQ!6���X���+f�o����$k����¶m"2r�c��ɕZD
��3a4Zu��;�~����h��[T�r?��d���{$�vvx��l�)+p al����J��Rg�/�\; ��TQ��}�D=v:ʗ��[k��f �[�А+�ݢ�4����v��	ҿ�B.P ��E�q3}���+�K�`�<�5������$��/�؅���5"�B���F�k�)KW�ʶ�-�*L��x|���|�l�7t��-VbE΄
(��h^ �8+A���Ŀy�~�����*~��IVQP��:�֟ڲ��e�x/j�K��K@�w���8E�br� �t���B�2�,ș�������{=��Ѽ�n>p��Y�D(�:-2��LŢ��̒8\%� ���=f�K�=k�[ �2�K��8��_D��:Jʒ�z�h�s�JC�,�袼���"�v�9KQ�'HZE!l��b�0]�	�,��x�(���N*՚��4�<��v�͚Y���Rϒ�za�(�Sвx&��1HS�PI�	_���˘�|�?��q�rL|��}�y<}�V���d����e���#�s�0�"�y�׺�G>qO'r�������?��߮91�~�JtLiH�w���lN[e<��\4�vˬ̽)ҹ4�����^w�Sl)��Op`��rO.&�w�6�v�mx	�n���u���u;IE��7m��>�P��~@��=��.��v�i$�߿8��dH�2S8[�r�.��47��g w�6��R���&���h�X"��H_�_�I�S�0���3�VN� �)j�C�'Sʚ����/����
��e�>nm���bl�)]A9@ٺ��xн�����>�(s�.x��؂yY�R*^�G�]�����zX�����aq�����K,3g�j�7�b_��-<��9�'�8����$��P:��#�s�b�Z�'�����a��~��y�
�j���f��OxG�/j��V��ο�^�����bGz�Fgr6$BN�j���v���A*����^A�^�m��鹛���x� $���ޢ�Ϛ�%����Dz�[������/��R�U���>�8�]ue��{��U�}>��|l{���;�bͲ�97�s���&k�L';f�zG����@���V-4��K��]�6�	>����S}�J6M+�����Y�N����J������*�/�_���Ae�]�^��A�ټ?�HJ�����O*������a�CA��l�kL��[�o�汴Yn�_����>�������9�>�+��n�?q�A|�Ƥ"����y��<���Ӑ]g*�B=�t�,~3��=c�j*s�e\f������HOj�-�W� H+�L׎x������X�_Iw�`������rn�T�����-|���،�l"�g�F�el<&�+�}�g`q��~R��,3�HTKGn$ky'+����B}̶���{1�$�-]��;�zh�Kr�%��K;Q�"� {�~�O�	���!�^C�L�12��r��{G��%~zF��~A�=�Q�І���HuM�����#Y ��8W3 �
��I��ʞ���S+��B�y}�Gx�f�������+
��O	L�b��@'M�D����g�Ub�����`BV��5�!&A;���d+��0o����.���>h��H;۴W[��Z��1�m29�._�����H)�k{�����N���;�>����Ipq�Q��@�z�k���#��S�te�R���������oc/����:J-��+�y"8UM<3���=l�pm��� O�� ����ΟT#��B}�1o����טc��"3����)Q���,�C������2�ȶ����>��6/�������F4�LݣTj;�m:�:r�?�����Y�A��Zp���6r7�fX��"�d��e�^�����	�h���2+��l��fZ���汧��9;����=��z"FpMt���M_��>g����?:�$�%��������P������GoR��%��D�r��'Am�		��n+]C!R���5����t�����y�U�h�ň)���k񪢓�%���_��Z��wu�-�D*���U�����S���_��&$
������d�;A���wb�m
����X$�����k�aԺ���J$�&��=�1e���k��;k ��ԤH- u|Ky�.���E	�:���t��;��6w
.����$�9���Qa��� �<溢�k+��ϔ��ݜ��J2:6 ��O���zGT;Fe�M��	�`�9�&�DI^=�ݜ���gm��s�!����?߂�z��cr�����& �vF���L�J�nm�+3*�]Y�RI�j���3��7s�hq�δYԷe{e�bv>���-�d��M��Bϳ�pG�}iY�w�2���^+��S mȞ��,W��Q���g�1y�E�Js� ң87��C��L��q����J�;Vp�_::���)Gkmi�Je孌��9��&}����o��+%�փ>�Y:8O�E��w9`l��1܍�?O��Nq��Ӌi��$JV�Tt�dJA;��<L�k#O��ܥ��d�r}̭��STE��Of:�Q](Y�yiX^7���)Yy��f׫	���~�Յ��(]�Sc�e�:^����]NA�B�-�T�#���1҇qD�c(;�
�0��@�x��A���_�~q�=�
��p����h�L���na��j�Kp�j�Z�����רX-s�w;���9� |����4+�o��?h��~�A�Zʙ�RO��F��?��;b���w���~}����@@��!x ӪN,pZ\�S�ۭ��2a\���{�nch��[��HH�-wh=#���N<�X&��$]�V�k�x�M����H��(�����.��v'��Gs�yL��2�h�Y���2�j��)b�ɥB"1_J�87+�	��w@a	6�ߙF�a.3�����A�	ڽ�f�u�=���z[j6��>X���)\����7�
�w���`�a��6���{�s�����69�ƌxT��4Q��0rb�7��KǢA�4c�f7���y���e#J|RFR1�Ƌ(���o��<����
@�hz���Xz���bß�č zq��hC��݇�@�E<K�'�4��
�����8kCDH؅$SF�%}ds�,��Z��3�ɋ���p�	@��htb�,�`=P�}8��H8kBDk#�`Y�Xi�]a�|qщ���G	��ȕ�x§\�hd��RNB>o'TJSƙ�(J�@8"�fK�H���-�� 7	��U�A܀(*��9�p�L'�gD��L�B�	�Ң�С�u@���(�S��)����`�d��¬&�Q�h(Ҡ��5\,� T�	e�XD!��8���Q"�? �������V���ED�p2}X(f�Q1hY�P���G ��Ł�D��+�QX/��\Q
hH��g���\�ަ%�FD
��Z�Cp�����H�P(FacW��)���&��"}*j&(�[��2/�Fu�~���ؑ\X�l[ƀ(bh1A��V�0y�f����%C|��;>7a��(��4C_��ڻ���ݵ�KlL��9Hi�f4�6��K�SF0)�`4��S�@5!)h���&G�"�%���cSĹ�x��v��i+�&�'��FS�����쀘��Q7:������N�%qƟdҞjS.���T�����~��R���J9-�-L�t���"�5Z��R*JT�iI}&��I[���U>�ie���|�H&Fi|�pi��}�*R5L�RI��i�������﹨�!l��QYJJhtS��i,���|7~�����m9>� +���?|tY�(-���b��M��c4��b�W������!Oc/��z]��Yӟ��������:}{>��^^��ϖ�E�Q��b��@h#: ��h��q]�5/R7Ri���`�s��p*B^+cA�˳P��+� ��g������wώ�410o��X$������TPd��1��h��(��5�:�4Z����X�4��y{���N���`�j1Q��XN<�C��>puLEnh��7+)LN�G�b�En{��w��>�M����5:	;�kg��
�t�ч�h��!+4�MT��������ha�Y!�C�&���Cp	o��u�`"�h��J��'�R��J� 5��F����a������F����Ǹ1)ԛޣH��*p�@�Yf�K{PB�0h/ARz���w��Lɔ���$��b�fvCN5N��r3�س:�2�"�W"��(�j;(6|t�v���S8��b��4m �~����F�������C��H�H�N	ʺ��N�$�Zs���t��3��
"����Ỷ�d�>Z{ʃ!9�1�����N#L�t�k*X#���p�6-�S/���/��Zu�yq�a�����J��r�`u9��F=��G5qώ`l����H�h�9��r�CD���5"Pz]�xr���&����9ɰSHx��J&��pa��|r#�񑊔��AK��zv
怓3SP�<5Q��.6���|��1jA����~��`���A��ء��docp1��b�>jh���|�Qx�R�9�ȍlQ�L*�Rn�A}N�DB2ݰn�b]6�1_���!^���'IQh��Ј'��X�=xڅ�zAaOR
�P�=`&q�?�ke��Pkb�2a��I�O�P�d�ޮh�8�B�:q�	�Lj@)��V1�_Vs@��tW��7����E���������zf���ud]�
5�I0��(P�a;)��K=��顛��G�v����4�0�B}1
k��Nx
&�1P�Z���¾b�ҽ����3��
ly�;��s	a?*��,�wֻ��(kc�P�jO�^r��IXPS�b0����ж������X��-b�k��'ߓ�����Jv���7��.�D����c�D`����yw��3�Vh�$��L��[lqX�hʆ���C�S79ߝJ'�6�Y�_��:x���;lfYh�1���N�;�4����������>6}݌�ۨ�dV��{i���X��E��޿�ƣ@�G�����\|Bŝ��8��q�I$J�~>1�drY3e��;�0�/�l�i��rN�֘�~}�<�5�IE=el��ʜ�D���-�Ѫjy��Du18rP%n�I��@�9����������&�X�ʥ��|�:i٨w�v��w�s<��i�cf-B�27���@�Z���q�>�P��g��f#r�I\�o[4y�1�@��e݅f��5�g�4�$,J��>FcI���d��J�y����lm� �`�2aAtC��Bw��	�z쇀��WE�_��D�*d�\l�E�����V���5��ƿ��{'g���h�w6��N ��u���Q,�8y[U���/=�Q��)Q�eg�&Ut��c?�u%�|>�y$���n+�c��9��6&���X�l~+�UŦ3+=cW�X�w�t�o�$��n�����'6���^��r�����n��l�d�V�J�o���\u፣V99���r{�̵�O�:
����{_��DMLY��+��+�Hn�Gr�m}���7����\JC;r��8�=�s	ݡd���CS�ځ�Z~�~�{#]��:�|���[��\u�괊�w۞޺s*������%L��5�+�NY;'��De�����FVV9���E��ܜ���0�W�I��}�'�����E�^�S'7��� 5��6z.�ȌHriݚ�l;=��l��։l����Ύ��ؔ��A�t�z|��ǆ�nTV��؝2�Իc"�O���%
�d���9�[j��$��l�,9M�ؤ�~y�j�����E�rd��R�����%�Ae;5���19_�(Hg���}�?n�r]==u�y��w���z;õ1��).��Ke�K�/�Ў��^�'I'���|���Mݹ�i�Z'?�l��n]�t�_s۹�n�ѳx�vg��q\@����Y�:d��)�C벽�c�.dlh���z6�ty!�R��p��ۂ��}�J��Ó���f|�w��<k��������F����ʈΨ������;,���&�D7������=���5��̐L�A@Q0K��� 1�� ȵL�LAV�쥉z��+���v�{
y�uS���Z�E�渹<��]pz&��;� ���yP؁c�t��� QK�AC=uRU@��5#UD�i�g���^��W��bXų��z<쟿�B
�l�o�>_�f�-�v��q_Ci��]�R��^�X�S�~�D��c~�dnӈ��5}��7'��&������q�=x�63��]�s���q���c��_r�XO����:Q�x��7�|��u��o�J��t����D���_�6����3�+��}A#/�3!�/ �o��J*(��_�GNQ�ru^.��1	|��U�L$.���P7��vӤn��o����)O����/����{����BA�<��H�#D���̍o�z5<c��C�bX_:�̚���Ʊ�F?௔=Y�йJ�X�&C�Nn��yU��n:)����������2��DI�t�Ӥ��O|s�q�y���*ȭ�Y��Ix�G�VG0>�jq���#h��)���xs�2u���z+��|�E7�m�?aOy\�0qw~Z^��N��~������<W}]q�Y<����e��*�H�����j�0A$�<�k����z��Y~��/[\��[���Ѵ.a������)�s��"�U��٧I������#��\��:3 ������i�HF�Q�k���򦼈F6�D�y����a�N�C�R��������.B��|L����{�U�K:�h%���ծ��nqfu>�����#�)(�����5���Oߦ$�����C�=����IF��c�����U���o2rِ��Ʒr��X�VϞ���Oθ�{�S�����V�A�3���?��������~�!���i��6��n���q�|<I�迣�{�H�n�'*6:'�����up�ҡ��:ѧ�ڧ9l�HGA�s��H%���(�ln��(��=�3��}�v+�l=��_��]����w��
�i�P��=�wv�'��'~�<�s̜7aπ��O*~ϴb����)c�hy��4�sO?[����v�?�0d�#\%���v�r9'��12'��l���+2�8����O�&�#=����J��Gӟ��������F��/wtw2��zO���ﾴ7+t.@�h�F�(<�bba�xf�|�%*ȷ)�W�
�����ȫy���W��&�<����<���'S�j&�s�����&<ߪ���W�6��[vKqyxHy�s� �T�Wf��4�L_�] �-L/�8�a���U6�LlսJ�~[���fY�LI��Rt\�}�-����������������I�#�7�o�/��~Ҙ�N$xI��kP���O��Q<H�ѱ1��v�y��q�c|�ꭝ?2a���;�χ�g,�y%T�s
�ծ�N'��9�,'+�KHr�^9�z��^�I��ݨ��������qKC�����Ϫ�+)��2�ɗ�pv�����Ϫ�{�59�:����?�i4��7j�N�ʳ67jX}�[�/�3�[������ӛ�&>;������E���۽�6C"��/ R/�������D?��?�COߣ�?��� -�;Qw������]��m��KY�T?V������˱������l�*/�fT���8٣'�>�#7�(������/�	"}z��Ǘ�|�D���A1T���5�B��A<��nJ�E�9��U�5sS�E���8�=��J�(PS�Q��`«�lU��9ل
�S ���{Vb5U�X��<�wC�C�Wf���.�Tf���BP��M���~��ݩ����d%��rO�SV��o�m	��Nɵ�BX�vSZ/zwT�_�"rmjǲ&��ps	��Gc����������S�D���XY�75z�(�����\�C�{@S-�H`CL�6z�R*�%D(�f��I�?�^� �����ʿڗ����-������a�0"9�	�9,��s�#���SkL�B�Ix'�w=p7�-�<7�z��'��)�aհ�����g�CI�B����:�GR�s�_����;j#�}p8i{�>H+�,�����8e@��D�P��"B��ː�?n����U���~q;@ܬ�:�嗉Տǎ�.T�u����VH��](V$;K�\~�f���vȯh��>Egd{�]U�1ϏC�p�6�U��&^8[4'u�.D�+��8�-�����ަ��-��#l%�]JM���><�RC���hV>�� GT�T�X�6n�Rpbu��F��]b膴��L�{�R��
Yy:P�4�ƫJ��{�؆
^����z��j�چ:��{���!�ʌ�����z�z�:�������\R��	�����]��pY��C�
 rp����h���4�8�R��Q�ȣl1�!��Tq�
=A��v�[���W��{� �Ȩ%a�yDGat�S��qeΒU�؀jGh)g�v���^�z<1J8����b��/H�2b��n)3%��i��
c����b�� 莊R([i�	y�I�:p���#|&!��U�NM�)Bs��?0ϑb2�惶!,�(�H-~bu��,	�A"�Nɉ�)F�����wr&��-����`렒%)�6�� ��B:i�;B���*G���*�S��>M��<��.�J���2��+.G�뻢��=��|z����!Zxn�1��QO\��e�ϣ���R4G�;&��-������&�֭ߟ���WhS]�]���Ȓp\a;��S�
�0&�Hd򦷊�N�T��
d�r��Ů�����oF�O74y��Io���b���
�%�#T�i:�U0upWp�ʳ&��vȱ@�X�ò�ͅZ�!)4�_^
zf���Ю���)�����F/���@�"�\s4Kf���؍$�	v�6�����*;P+{fn�Z �[�ʢ����@΅[�I6�������� D�O����
wai� 5e\��v����T��M�PR�U��0�%�3ه>G�)zd���YfQr��TTJ���ć���*"��4�:����gڅ�n/��� ȶ-0q1 �_XJ���9�%�)�0�0����o%YS����}��#J}Ŝ����Aם�ȵ?";}Q�)���~c���))ȕ�v�?�M*���D[0q�T`�,-��A��A����=E �^�q"�N�D��]�(���mN����Qu!��u�C�)�>Vǿ�<�ȭd;~�ҵJ�'!;&�G���TuY��q�[S�f�j�h6�/���j��dg7���I:�
�C����5ϕ�B�>�2}��JטW�C܏݌����Mz�{�;!�����ݮޯV��>Dcj��k&C
���s�WT�$�*����S�iZL��zԵ\Xp�fpk^�^�,4�z�,��=Tc��)�qfa���1+ga8�����֢|*dR��0��,QZX���r<�tdU�awS��ꅞp>dA���"�L�S�(��:�q�97G�#�DĔr	s�p��G�7d��e�܍V�C�b����5�����3��Q]���V�Gu�=�ϱ/���s����1qhM�vj맶���Z�܃�;Z�bN���{|�¬2~T���H��[ZtB�/��Or`���4U��eQ{�:8�x����d�!�w���:)��:��|4a��<*�AI<��>���V�`[�>�x�X�$��F~^hz cζ�>��v������D�h�T E 	�C�����N՟���W�̭l��|>n���AsyY �/�a���a�z�^�e��="��ld��H�H;X��~~F�N�'t�dj��p�>�3(�RZњ`NoS��1@�L�F����ǰ��%��o^����ݠ�aT�j���l# bT¥I�N ��Ƈ����M��9��(g��8V:$�L��ONh	\Թ�\�x?��ȳ֕�Юd7���K}�c	R�O�5�U�A�!�'���jS�
)�m�5��-eթB|x�/�@�;V��uȲ�a_I"Y�U�Y�B��(�G1���ye),��~eñ�Ԗ]N��Ê�:������R}܋�,r�2}I�q�m��#2K�l�x�!z���ڸ5ilf4A�Qeʼ��;�l�݀�#���Τ����ԝ�n��p�Ag��^S�#8T\q�T��V2�����zl$ �;�%Na	 SZ9�^<��*)�Jܱ�cq)
�F|�{�vrR�Q@��|�K�]�+��|؏�,�P� �8M�{���t�,G+jX��,���'Ǩ���l1�i�h!cޯ��Wv�K����"��9s
�Gr��D��Ob6�{�_�Ŀ��4�b�X4�)0�
�f�*x��pZХ^lT�u���aT�D���"<5�8|X�hY�=�)�#PR3�����G.�/����x��� �ؘ)`�;� #�+�E�a��r`&���h�,r���Ryʶ���?o�.V�Tγ"�a��:Q��Lk�+�!u5�I���ſ��L(�Ӆ�/hv��C"םP��w@��R����9��[�=iM`��݊N���<�Kp�ܺI���If'd:=e7c,�B@ɂ5��t�� pI5���t������}(ɦ4t�d�r�eE�W�"у�+(tS
�(��	n��ܓ�N�5��t���1-;�prx%D��!�����.�@]b%g]�&��[@Aa!`&,E��橪�h/2D�w	�Ʊ<�CDX&�.�k�L����\����-p��������h�u j6Tw"�d���}�Mн��r�02�ʔ@,����� p�"��ƞ���KlA�J���r�B,��/��������eB�*�5QRQ� cg0s�
��:�-�s�C �jݐ�+��֮��3�Wc<`�:N�����	��������z�GIN���`�8\��GF��9�_>���G�,�=}#�$\K2r��J�32ۉ;�j�d�H������
%u0�3�Evⓝ�I�/�d�Q`���Cv�%�J#ĸR
۠�Bܪٚ��� pp�@L�8�w�:B�᠗ ���̩M�s��M=j[�?N'��/��#S[:9d$YHl+�*C�<jW�V�.�7k�����đ@�u8�"�v�6�1�����Z�?�[��z����ȓ4�֛?i#�%t]�M8�ޥ��X,�0՝]}
��&`�7�#^E]/����%h3��zю�5J0���=?�X�YfVB��/�e7����RI2�&�]`��M�̓�I��fSPM��<R�ٍ<ryv��c�i�z��H��Uw\�&2	��u_�� 4Jr��ìa�(t�%
A8�D>43�O&���L�JpG_��Vu���B�w]�L�;D��xG|KX�,�9���B{���6��#�O��O�����p�:���s]�!�KG*�8��L�lz��5lJ�`Xoh�%j��5(�:F�Q��󸄕2�p:�{��Y�I#�EF�M�l!���Qm�<�B}h�ꑸ��^>��z�+$����U��:fQ]���IQ�M�E � ����K��� ��]�����4�\���-������w�"���i��r���*�6��zMv���1NGD-���I�D�'�r����&_$��k��j�/�����D�t�Ն1/fghj��ij�]�J�e�o܏�[�����HE7��v��Yw1��%5"��s*,(23Eƚ�X�ЂG����Qp��9��ƽV����B��T�5�m�+���.������!���jk������#
�^&���1���ܯ�Wd	�$��İ�a�t��ԍ��C��?���Y��s�A&�]��xB��K:XKU!��:��Z�؂�牄�)�Dt�Z�d�n�O���˲I�#��h\�c�?�+���U@��YP'�zC]2���C�:�����H�I��jr�^DU��aI�bQ��J�xE�+s�9KG�0�yG��G��\Zna&��m����pZ��#�<x�i�A�E�r<��ϲ1�g���։`F�H�Վ�>qa.ZJ)�6/>�T�Z��2��C��*��\ �c�����ؾ�]\	���	�:b��X�T�$N�W�*�X!�f�*�7ǻr�(g)9A�ac�ɯ�^p	��q'�$�O��@iH��O���/�E�p-Dr�jG�ɜ$�S�� "99$�K��z���P=�H�\��9د�2�����Ά!��6���u��w\%䦀!�'c�����c�e��ۑݪ�8�>$�v�Z%W�ӓ�`���n9 $A����tֽ2�t=���eS�{�5ܕ�y�,��5�R�3���M�=���b��(��Ⱨ!ѷ��cF�3ժ�ޤؗ0	05���m���$Ó��}%Ii|�)�w;��h:��]a���b9\4Au$,)��]d�@��TJx92���$�s������վ��/ԏ�wPG~�l9�_�Ü�)D6��OC.����|��Y�4��gu�Mݎ���������d��m�ke�b��D0�hk���sZ��a�o-���D�е_�o��Lァ=[�Ǌ�sG`X�e�\�% ���Ne��Y(���2�ڍb���r5tʬ�V�6�*���;I��Ր�
��!W\¿�+̡������<�Ey)o�͉Gq�܉�*N���oGw@K��J��q�x���ڎ�Hƾ�,�X��I�D샓� ��M�MxZ�	ߧg�+*�<����Y�	�<@���sW�T��d����\�zW�C�~�N��3O�%*��d�r����Z������Pu� L�߶���0훪���ʢ�t���Y�)�����Y�z�-��$�6Lr�L5�1��`?�����r���)��Qq!�~��Ĉ)J
Q�|:-mY �@ek������!�.���Z��.��"�h8���(9$W�AW�T{��(�%+"�'`@�� ��������5uI���%̈́��v,n!�C�0aY�4ِ�h��Y�~��7�;�	�ۼ��`+'i�r�S��K�t*�t��s��*�P
IGPC �(�Z�nWnl��qY*{�\l�K�����I�U؎�V��M��[�?E#I�q�I����-���x�tk^������b*�5�)�^�M@)N�p� (�Z~[��E���4�k<��`(���=�bn�e�A��r%�o��V8����_\P=`{��c�[4�I��o4��-PJ�Ҵ���?JO"�	U�B�;)��̓}���Un5��F��s���`��p*�s|��r�Z���^�pV��]�
�g�Y�=m)�'5�XO�$� <��(�.��e6���w<�ɴ�;��W %�JZ���i.���#����pI�.��(�iӃn���;HĜѧ���.
��ɏ�s��ð0���c�x�T����3��<���KU\��OCQ/���^���߉�������]��c;݄�������>bwpG�~$�w?�F��q�i�~s詛<��[dt���'OHH[�6�r����� ��,;W�)j���S�*K� Zɉ�QX-��S[�^�����S�g�	�-f�y|�/������5#M�z(De�U>S���3�+t)�o��;�@�K�47O,��
���=dc���Zf���.Q��BM]�2~���rV������3�<=�q7�|��f�ky��L�0���!u���$��k���G������^zۄ狺���Y��c��s����3���33x]t�U	n����/�j��Uhn4�	(�{�=j�͟0
#*z:�_�+M��Ph^_MYi�j�d�>.o���[�ȻV����O1�~8Z�u2��灞�����=Ye����9w��([�?�"]�e!���7�%�!\om��-�ʉ�/^r^]u��z[��+�i����������c��5� Iy���j��y��="ɒ�����LOt�0��rR��P{L��#�x��W�q��#0eھGm~� ƃ��X�Y�+����$⊰��}re���X�/X��.7]�3oß`������r��\;&�EY@�^}�ht}#��{u���/{ɕ���}��a����&Ř2a��'���L�;�N�۾�5R�1�3�B��ɔzVL�Q�d-�*�%�%�2w.ɗ������p�\>���p�\>���p�\>���=���(���J|EW�^�ȼ�,YF��u{��бְ~z�=�[m�y�bWA��z0a��u%}�q�Ϩ?k�����0Y&R��c�3�ɼ<�%�#睪�3O9Im)�]�	�L��~N�����)��\m�|�:�k��;:S��.B�P�tD�&�6�Ue�/m�G��"��Է�АB>J3�{�Yo��y�e���c�i��WY2�O3+;����rf��t�M��2�h���n���Z�v�Q\8h��[m�(D�?�!�NӶ��;�v�W#=�ֶ����9��g����6��^��E��u�AA�!WI�g���.�{]�l��t�G�U�t�G 5���3�r��Y�&�o��(��6�Y׽[l2�� �"�iqy&kk�]�?fg�Q͆�y(o[!炈z�R�O����� �HJ]�@=��{kդ�����:5k;�!J�/B]�Ŭ�tu�m=��Gר�#��u�a=��G%�[C�a��d��������ZeG`�M_�BJ�(5X�s�I�5s�F�H�z.���-�Ej�7�z����zk�{)/߁%śѿ��-����zB2z҃ԙ�M������_��G�����l���\�꯰�+#.��lR�u<������5�잭����7\pw�ђ]R������Y�Ynh�i�Z4�����'@�M��춶������<�Ӝ�����(�uc�ٟQ�v�1@G��Yru�=��57o��;dۭ�g*�\�-ӊO���{,
f��Yߑ�&�]�z�������kwSm��s_=vߞA��Zϗ��q=���;���Iۋ��f��K�;a;{i�"ܰ��X%�<´۠��g��[�I��<Z�ˊ�q��dX�,ӥ+1���\_��n]�R6PR�l�c��9�3�&|�`�K�u(hC5�3� όM��_ޡ,4�=o��W����[�1{tݦ��5r��OQ�q�F%T��}��Ѝz���i���
��>���ؓ_(�z4�yi�/�V�ǎ�F�|�]d�㝗�T{�Ͻ��H����1�)���LixQ���3�ݯ�u�L�y���u�����X���F�<ǧ
��(��d��&��Q�F��M2�1l�r�QzGG>@��k��Y=]ޘm�P�_r�Ed绖��NbCs�"|19,��m���ݰ�E��x}�ܢ'�����\�OQ[`����
�.._��g��qi;=�)@�F�ؚ���y��U�F1�%K�F�����_I���d��,ښ�'Ϯ�eN�����y�с�Y�W֏���YၕYѠ�V(��R�*�����3 ��X�R�K��J�t�@����<\̃I!*T HL3<�p͸�n[q�Jh@DK$� _A��]Z���ߠp���2��se�!=Wz�!���z?�hخ3�6�;&�/N�bhK��\b�Űr%�|�'�I:.�/��?�7��*MA=���8��HM ���\�����2!Z����~$}�W{Fp�x,>�lո-�h��^����7E���EGx�粼�RI�������Y2Ԫm����I�\Pf�χM����C+aփ�A�� ���U2����������=����Z%]��^)�<����m��?�U�w&���6�e���Jq_���R�.(��|\Ŕ�g�G%�_��/Pd�EsN����<V�� �V���=�_���j����Z}���bAk�V��W���d��d�V��-F��ଫ�\-Jn3�?k<�#C�Ǝ��@���ׯ׼	͆���V_{Yg
�Y.�Cx`?���U����tF��8�w`H�U���	��ߐ���F�Ĕ7x�m���-� �p�vNJv�2�w����׻;i�Ӳ��$�@V�_N� �j��,wC#LJ�]�҈+�];���R���DJ/������n�"r@3_;q�Dg��
c�Pef�����qM����_�s>jI4��ˣgn����:�z~B��ݯ-�Ijܾ�P�{���S�*�`���Z�c��T�^�Y�cG�V���9=b�,���:ا-���i6?���O�q̀���H��7rԽm"Ǝ�xQ�u8�`���oB���s����үs��Ժ� ٹ�G�Z��75�{���p��
℟TE�0�.(�R��y�7�<�V߬=!g!i�rh/�]/|�Gv���v�7W)�����&y������}�1��ٳ$|d��v�y�װ8�>j��Mq�� ځb/=RT91?Ka��(�tu'KJ54�Oo�>�\Ѽ�8��e��4���A�x4L��9y1"ÔW�O��vpq�i(�{�rX�wr�q0�qݩSH8-m��@}:�y�]N�h��j�|tT&��<���u���>�SJ����#�%cK��R͗U�v��l%r��q���:�SF��ǫ���cA���.vtb�#OJ�f;�tA��𣩆�b!����T��^3��k��C*�{z�} sZ)������E�"H�t�������4[F���I�[C�!C��~3y{�Z��出�R��`9���ܝ�ϝ�?�D��D�SW�brg��7q>�u�*�cv����5�@�]Ԓ�������t8��p�v�7�)�.^�b�Qh��n,ˆ]:�_���͖e�?&�_^*�퍿�}��=�Y�=&�}��L�z����7�|�5�w�Q��$��ݵsFQ�f��w��*]W=��H9�J�e����O�!���ww
���+-�C�w�u��Ҏ�`WX�~h�(�g������KG}��|��{��Q�k�}������V��s{�:uc�ks��%�7f�{�\$�Ξ�_����;�7NL���SZ����j/[��֌��kz-o�kt�7���R�N�\���i�i�ȣ<�D�߇Flf�~���mA�_0�\���{���Sgz���l��g2,�iq�����sJ]Κ�q�SSp�xHǨċ�5�ʣ�\ARX�|�Z���fcs5e�&��*R��3���V�sm�昮��U�NH��<��\g�;�k�4��Sh��r^��'�|�;a�}f�U��©�	>���}�m�v˕z���<��5-aQ�QR�jt?�O,��8�3��e����u^鸫r��!��~+	����n:�Dִ�N��~1�4_�O)(�W�wE���#�h����ql�Q�n*߻���m��8�n-߂������|��>�y���R{�A_���x�uu�Ո���P��4_�`�T����%Γ}!r��D�q��y�B��׷ �l�N���=��v��y_��qs@Sn�l��F��fk�s�4ou���7����=A�>��J6�Ʋ'��p�p���F���s�b��/�:��O�� (~�);��S
w� �y�~���H�غ��gЯY)���xK�ګ�o|C��b蹒�ڝf�YC=sE?�<��1�-��~=�(k �k�`znbu.t�	��k�k��,��2�[��n�?��~E��ᗛ� ���t����OI���`	G�P�����Ԅ�u�Dp��L�,&wA�.Um�+#m�I�s>{���G�ńk��'<�
Ƙ���"J�ׂer����x�qx�����_�ܮ?����r����qH�����fvQ��co6�6C��u�+���Y�?
�,ٷT��������S�|®d	���Ab5�]��̴�� }E��76��y$h�����$57^���{�tF�	���͞�h�2�����9$���^���K��dr�A��擑6O��1B�H���vF��#���V/��>��8�p�g���n	M?)�P�ϞW�s~$�v0�N}��˿�K�~\�1y�hjt���*;��W�H5�j��4C��ũb=��N{��as�s�F��B���"�y <�v�',B�tC�ϐK��TH\�T	�;^����!��ȴ�"�F�E�R�B�t!��M����=}��/Q�"��r1n����?"az!��(9�_�e)�2�RGW�����ٷ� �7��X<�Ŕ�l_�w��d�{�ǜ���2*�F�fzG~�S3o�c�������y�Q���̰� _�j'��	�HpJ��'�}�O��r�����ty� C.�vN	4����~'�t��
.�X�4[cg��R�h(�39kN�l���d>�v;@�+� |3��|��e�1<�Cp��[����9`���8�|�O���w�B���th_d<���8!R=��9�Ƽ��V|� uI�����_ ��r��w��W�>7�]��9���3��y{�vN	���y�B�lg �~���N�u�(�=c9�>�hЌ����y�8_��2���xk=��{,���^V�!yF�d�����9�w��dU��i<ف6��M��S��5C|&}ޚe�瓛R`L���}h̀�����i9�e^яjQ�MW*z�*�����+�%ᯥ�jV�xL:+�կ�n�#"��WoK��W� ����=_����*氾������3��T�rȦK��
�5Ʒ�N��V�aQ�)9#>��jwB����ȩ�<V�S�ꅵrt��!�j���C [&N�|��Z��CZ�N ��f��O5C���̏�7�T����5՞���]tU��*{_�p�uT�^CJ����b�thI�G�O�Os�UR�Pse�L}QE-5+��
~�W+ǧ��&�
��W��%^'ڣ�&�i��G�A�i���4D�$���jN,Ø�`��)����g��'x{�b�HM��+524�Z�E�l7��*u���S�Ɉ8��ٿL�_�:����^�[�&��3%�z�B>�~��.���
���֝q���n4��5��Y��T:�
%0���N��}�=���*�rZ˙�-�tZ꫾�`�C��K7��J{6���t�W�/(�����>_/���x�!�����G+.�A����n�"�"�+$�՚ +B�֣�șXҽ�U�����å/�������0�%��M���=�դ#��û����1�
Ύ���>H��3�m�
.�b�$J���п��Q�����hKl��q�M��A���E��@p���o�����Qf:�Z��'3n��<}�8�S��[R6ơ�ܘY�Bl��<k�P��[�ʨ�NM��#%��Q]UL[��x,�LV:�	=ɹ"�	�-��q����1a�:UtP/�� 'V�Ȏ�шiƽ5egD���I�SkX���f�es���1a�lV��Dj�<=@ڡ�]UCG�D���$�$�US�"��3�@`l�T±m0'�����.l��E[��j�w*'`|��H���G�l�OC��*�X�VBL��j�E�+�<�>j���7�2Q}�<\�ͼqE�-U�:��\l9���e�Q>��^$�m��xwKؓ��㏞�Ɗm7]>���,����z,ōX�%M����-+Oړi��`m�Eѽ(���T�$A�˰�$ж���՘��m��ˈx+�^���9kb�~�����>V9��{r_��	�'��~������,�g�nY�����z�O[ฎ[K7H�+�}�+
��\��H��<YX�J:���Pw�L��1�(pZ�6lh8w��n�}4��)��Ĺ�w�L���¨�P`{�}�W!#hB|����}g�ۼau�� 5�Z9�����tNx�ֱ4�U�*;�r��T@T��F�N^���t�������W'ӻ�)���h	�������L�}CoDT�|����R�a��\��ϔg�Z�H2�����/�Ԏ���LӇb������Q�4<]��B���͎�V'i;DM��ŎmG+�nU[� �gO��f��m�r��a
Mf���||��ɨi��A7q���.ܺ�C�)W���X �ف�����H�U����걮�E������=t�0k�+!��@M� ���P�Ϣ2�o�juO��s�/�^Ù�vi��C�l��jr-���M�C��Z��L]�ū�rUa[tA,����-��J�����뺆�Qf#�&����Ԁ�(m��W%��X���%e�A��Mȍma��ؑ�$�b��3쫊���A'=�2q���UA$���yt�&)>�_�)0}�Z��[EWJ�+xT�b^�4����~�`�n�C}d�[�a/�I%�̊w3Ծ��'%b��}P}���b�y�ĀP9�w�Uټ����T��� �KJ���P�\�}�f��	1�l0p8��a�:�i�E)@�����@f���h�5�p�>W�
����L���a�em�+��֥�c4��N���ر�d�׋�zb���ئ�~Tt�y�{^�L��x
�n��<(����B��N�Wհc��Z�,ovP*��&Ҷ���C�)4� B�B�+�G���{`�}��B�C���Fv)9F��2���^����.��sWn@@MM���y΅��U��:`�V|�$��ٷ�l�S��͑;[�ɟ1�jngm{0k�/�g�cs`z3[XZx��L�丟��m���U�m:��V�&�w�	']�f�R^���s����>(�'R�Cj8D��-;2�șC6E�J��P�@�ffLm��C��(ehM0(�f���|��&o[p ��:�PÕ��D�6�Ƌ�<ۀ�"
��}cF�j#$�5k�O��� 4�,�l�O�/\^��Ads䐧�u��P�E�A�O^wnq9�-H!�Iu.����0����?�q � m�'R��U��]tf�
Mܕ4p�l�C����	y(��ေ���C����
�|3$W�?3�hB>�bB��lWX1u�Q�T+�a��]�z���hp!�m�.�Τ�+�����y)M�^WKX�;Icm@�#�"���0l��2�S�)����@jHҚ�9�6��{4xbc�0�Z�R2�� ?�U�P����L�����G�A�V
��i𧬣
U�M,�^��̭A/0�7� ���Dt�w=�2]�����ϕ˔�aU5�������!��@��T4|���E��������5�d�ܑ_E���[�yJ.�6��W�����H��+p)"X!��*c����l<z�o�������%�H*�H�������h����jv��>�E��_�G��@ol���CR3�A��>`�h���<u�.�\��HL0Tk�E��\Y
���q�V���Rv)4%�"��|��A�:4�@���M|�3���'�|P�94�~�>hY4z�uP.���^_Dn���[WA�c.T��%�=����<^෎�	I��^;��lO��	�Y;�r,�Zý�vMqg4��0q�1.����g���p��` -0/����!yY�9�zrk,��h-2���
���X5�C=nD1��l���l�5{&sK&��2��:�"��=/h'a&cI��i�U���Е�EM�.�X_cUU[C���ug6?oo
�����~�lr�jcͶ�vUA�,Nm�Պ!�K��!���K�������	\ܲj(���mܥ�u�s��(c����a�ɽt�E��D�Y⚵�e�l�(X�,ȤR&�!hEZi��R�@G2�f@/��{�| ��@��$���ao1�$�X���Dr:�kF�V�?z0pñ����H� ��H남x�h��a�,�͐�mɤ�*��C��ô�:�{��a������]/fB��}l9���\mr|��,?ˇ���܏�cYB^��:�*��,	�^T��%ϲ,��@�L_��Y8����x+�'p��s���܌��Cy�]�X%��@+;9Ƌ�|Xfw4��a�pC�%�,m���3r#�̧Qs�>� j�������U�bm���w�b�D@�G���6B%'�q�O��Sy�)A�����	�<�F�hA�=�rB���U�<п�d@��Zbz:��)��MXڅ܏]�O���c�<:I}qNG�����Z=��4ϑ���݋�b����gdp&�aY�䭡��n/�ڶƱ�T.��ㄠ���{3,-9�L�c���?ۘO��30&$0�ևSp�@�|Wl�< ��o$U$p^����h�ա�������RSJ�*�
�KL� �.F�'5в��9�]�X����w�a-�H�D�QMlK��z�;�]׫�P��,a���.�+�$������S3��1��ͅ��b萌�cx;��'�T�J���H��
˜{�]e�]��fV��A�5���/�^8("�_u�<�TJ�zDD[IT�V�i`,]��رp��_F��.ldh_	����'�'8.A�ebo^(�s]!�qo6� '�����Πc�9C�kVtD 4����6�;:Y��z/�k�:�iણ�Bиy��Q�KzIW�L��	��
^�¯"�nج.�J��)b˦� �,ni\�w�A��,O[�#}�U���5�jS�a�Դ�$`M�~K$C;XcI��Lݺ�=ic��yT"�Ɗõμ���(y�����b���s��06�e����s���o �m�>�xD/�Z�|��~��j��/��ڳH,�
��шP̲w�M.�? Na�.Q�.2�"xƍS�e��%U��xc,�:�'v�EU
�m������ͷٸF4�á��hx⶗V�G��&&�A��DG��<	d���vGx�����*=�z���@�ȥ_9lN.�����E5�30Q���I�N�O#����]�eO�+xq��p&ܥH�(q���:��C�vp�D��j]s��-�O8�,4R�-����9j_s�9�s��xh������K\����һ_8�:�)�/K���蝯vК�=�y�~��2����Ih�\��`�~0�lۊ���u�7�7��7��&�����"��}�f���E�K�lk�n�1X�Юl%�əXQ�/�w���M#� #@�@�%�2]t�s������T����A�9m�C�h� M�`FU�U	��*T�ɱ|����^E(�vC�O���J��-�i����	�x���1k��*���3�\�Q������L��_��_k֭K�>ۇ�������T�
���H�i��6%���S(*�Ί�7�O�\���'��SO ����`(G�o�k� M�s��ށ��0��@���2��~kgN/XH�*�I���;[kq���;&x5�!����^}��r�z0�
u��ɫ�㌚��A��~K��x#����kS@��Nm�n����C��:���բ�g#�X���#4�DȒ��68�rx�b�*g��`����@��~�e����X���~��9���ܚO�`��z���|�������j�oL�nD�#���@�&�h;�K>�U �}]�U`��9j����i*#v:麟&le�ªou`˒'���A<¹ہ��ז$�~h���;����R|��e �Y&�4�k�-#�D�����S����F��y���`͍��7Uɫ?=^I�\���L����i���%�Pؒ�3?��:K��gg�@�4��?��j�쩀�L�f���[���Z�4;�wMۭ�0+p��nӐZ��J �h�" ��@-B���$�����F��4x��7�	�
"�$[�0���	�P� "8Cd��B峩���M9\as�*�$��Tm0u3��=�Y���"fA�uݰ'4B�ʊ �0:��ݷ�!#&��8&�J��O�+X` ޻֝�Ŗ-4��s�����C��](3����hY�v6�r�W��p���ߘ��l	>�,������l���;�hgYb�烃{�������Xf�۾vXSs� f�L��/=�x�h:�x�i��vг	*��_���$S�������5D��/���S���GFP�yC5�>49��|��,1�Ze��A�Q���5_\eȦdb��.0C+&`�<"]�˶DcQ�t��OʐC]��$a�J�F��$�vVp�t/8��a��)����m�-�dԡ�Yx��p��"-&�)u��h�Tʼ\<l ��hH f�T�K.V�\
������AFE4̶0M�� 7��|�B���@��-��KZ��I���^��J;�4��b[�O͈��(�U4���k�^��tq�?O%�O r�~�PYm�<Wt���=�ʀ��(Yռ�b�mknm�p���?�`2n2V�pj���[�M��^o����ÂQ!=���5��+Bovr�	�'a�:�L��[/��]>�I�_3�H��F��B��|�MP�V���D%�x���g���W�̍ܖj�Z�<$��:�Pޚ���Ē�K����Z3b,�����V|Y��v�hw*��oY���S>�9=%'s\�2]}��EE����Yk�&��P���?1����u�֐c`�Go�X���̬&�U��zRI�0�g�hxݙ����ϚIU�����tO'S꫊�VR_��(Da�5�I2]`�5�B��Q���I*��J�3�$@��4;��mџq������'g|
烯�3�ꟍ'r�ɑ�x�6��j%�{�yO�!��@N��s�j��CW�fs89���רXa���z�۝�i]��(���8$��Z�i8ӁSK60QMJ���c��ZO��2�8�u������Na|�|��z�$ؼ� 4��nce��iwf�|��̴kj�G��^���w_~�Wœl (#�����x�cȰf�J!�KM1�G�^3 u���9�&�6�Ed	�:�0L�"��.���O/۱��A���8#��[� H���b�0 ��c�a�+�~Tt >V����2��/�X��h�F<{�j��z�L`��`������@2�ia�1�b[;�=D�q#%�-��I^�:(��i{ѯ�h��}I�����\��9p���ԎƠ�w�E�H�s�E�>MĄ��v8(����8w�6E����k���mTxac���[��
���u�U�z����L�d�w��;`"g��卩��
���A�k�z,��^qne����x�R��d����lr-����nG>��d��C{���c��Gd�~�'�)��Q��*s*�XI����x�M�EP���=�l$́Tےl%��FC
=)V�LB|�R�m�r����ʜ���yn����+~�]��g����ne�6m�-�]x��-6VL��#����9���'n���&�
���x<�s�I�����J�~g�6�7����F�d����<�:�!�/���`'aH�v���>
5��sH$hP����v�DZ�^Mu��U�2�m�ᯮ�������!�FG����������nt�t�멥A��	�}S���k�VKJ��)a�pT���rT�*eul/��Z�U8��M�%�l�`�5GB�w�X��0��i�-����^���*����=�y��T����L��R)���m:��P=�᮸,"QG�P��OA7�%A%F����_���rL�s��M8��zlnjm��r���������R!�*f�%b�5+KO�q{�(�~�Ae�k�/�,�*4���+}�%sI�\�<��PI�j�bR�}���s�,BnΚuS�sJ�'�T��.��ѧ��%(b��p�D�V����V�H���M)B����u��O�`V�S>0��M7ލ2�qP�=�I�J.g�"�2���åS�
}'�X��^Sp܊�Z��Q�Ĥ�pX>�����̨fF` ���-�sun��0b:�2l�!tm �,i�&&�5&���u���$-]d�2"A�!� @��I%�A�2e�_���L��p�e�=I�r��-2�e��-~��!1���HP�q���1�L:1�ƖI��:l�B7�Ō�7���!Bn6I7�77n��یܽ��
K�l�����~��eə~�����y��}��<���w��?w�Iþ��j�ߏ�!:��\|a4	��؎��ibdu�g���P����t�T�"�T�����6a���K�~I �B7��'v�� I���ű����CH�o�� ��J���t����j�%$&4[�CQ�_�t�lf`Arx�D. j0
l,��� ��� _�̡�6Ag�v�ͯn�w.]����@hچ����ߣ|v-{w��G��c?{0���k��P��b�¢��~y7(���1m�V��z�/@�r'�Y��u�1�ko[ð��T�� ��v��Vna=.�3G�Dw�V�������~��"P��~�{���?(�4�BF��W�w���ΈuN�C	���PD��y���P��N��*n�It�J�D�����d�7�taN0���W]���h2LcM�����t�CM(q�T�f�a�-N"T��оB�8�LS�ĲR�|�V�%)��3���Z������H��|�Q|8�Ԙ����,_��u���&��C�}q�d	�;Si�H&��z���������99���svI}P��q͞p*0�9z���ii�O��C`���	R���њ���4���K���ds�0,
a�~v?=�M��T�M�y|�Y�,{L�w)��К8�2���e��{.n�S�+~�|�
��;��[=;�@.#�s���f�ԛ��k�9�0p��R�G���P����I2��)|ga
���6dfy{H���,��R��
�q�Ҧ$�;���̰$V�6#9tvd˟���Nzs�9ai�-f��� �(/Nq`L���d�k`�_��&�3�}�{���^I�����w!2]Lr�s��1���W�Y��ׄ�i��o~>7iz�ޜ6d)D� �%P�i�:��)Gvt(��.��Nh�xOx�F��˻ןu8��ܡ_����'{-c��}?��c������`i��L τ�:k��ē�Dx�/���,��*=az�W���ŋ��$���o�1�$&"O���bE�q�&'|,I I�H\�%+�̲Mz�t�cF�� �0>"o�	��=HS'C�}��h6k�M-�ֈ�W/{4�D� ��hZ��*B�0����ے̲�����kf)�IYSKU����K'#��q-IF,f�y�7���� ���
O2ø�j}� &��&�`���B	1�� e�2Ir���l�w�����B��]������H�*D���r�.�� ~�
�L�G�A�SBcHl����t�	��9���R�1͌N�6K��A���8s��P|�'��x3S��d� ��,H\�X(�X]�8u/	K#>�%���W�*=��I�|���?����yS5��	8e̙�7C>.ֆ��Z (z�0h��=�ȡ���dTe m�I ;�C�Չ��5"�E$�!��
��s]m`l��XH�/k+>����J�w�
.åyr8�u#5�^��L{t"����p����;�^]|�3?B�B�;W���O��O�}��b/�����A�i ��8���
w��:~}��p�k,�{���u���`�4�e�m7�{ǔ�[����>�F:ʣ���Gvݨ6*D���i�h��n
}σ�,���"bpH;+��Eߣ�8L�_$2�$��xu�y#�𩞷{O��&��ax�ᶖ��f��b��K]�v^�c�*��G1`ey/i��p�J7��;66�F�.֏�nO1Fr"�t��-ٰg�HB��
����@U����?Ӱ������_�?X/��3��a�4�=����!��~�KI�c>�H�����v�0���V4T�\�vR��u-r���`�l��g�D�cj�(�#�m�%���2�h�
z� m�P�=���*z��몔�fƦ�9'l-5 ����#0�#ଂ��Y����>�t�]5N"��	M�9O~>���y�T}!	�cA��Ќc�{�rC8��E�1o_M}4c<��ŀRa����u�/�Y|2z`��jZ�Z�+?��+n��]$�ӿsc��S�I_�J�l}�1�+���|}L`�c�m rN��U�
�gF��H�X����еn��Z���?m�K�������.�qgT}�(!/��:��>�S@��h�r��B��$e*�˦�R�����L��ӻ��Sr�!�G_�WWj�c�u��"�JW�d�?/�V+�=T��*����=�G�5i���W��NCB��20�����f�NS�������q��*�[�
��㘀��?ԧ���{��?��X{�D��5zG� We���a�5ֿ��Q�g����&r���0	ʉ�!(�"�j%����6�"�d5
�^��H1=���H��>��L���m ��\���m��=#��I��-C�O`iǫ�2ƿ'��A��D����>|Ƅ~Y�K� ��ٍ���I�>�vH��ƌ���y�����;3窫���HJ>a�s��&��S�>?CS�ƻ��i������"E�#���1b��]]�Ɍ�HS+%�J��GVC�vp>��rևh!���C��S��w9-�λ����톆��e�hh#�����jF٢�R�VX��&���J���Ƃ]�@�B!#',�A�`ʯItt��o�"��	��q`����en�K���8WQP�I`������/��^�bC|1_�Ϝ�0��W�P[5;������U1�t[��l|��U(��.��D��;V4� ��Gс��_��s)�n�$x�-�$|�J���m:�n4����F&@�N�9QA���wp���]��P����ٷ>v+\;a���v=��R�3����:�sF4��LC����;�7*�ݟU��3#�����̶77��"^����\�����G4����؟=f��(ֹIFyz�7Qݗj;��.?%�~Q9R{�/Cm���5��4F�|)|��DF|�(�E�۷��,�=���u�Ϳs�y�������W}t��D}��������c�[T^Ǭ��g��䧡��Q6�0L����NZ��&�
W��FK$
a�!�B������d�l�8
�[ `�47G� ܙN��"� q70�i�	[3ppoo�b��<ǣ��64e�lXЅ���Qq����_T(K�y��v�AKx�D%�p���m[d���<�y���*�,�3|QD��H��������*XBTNNE\]�>�)Vj3�Kկ\,H��
]a0�x�2��՝8���ːX�(y�K3|h����Zn.ev����ƻ�"n�@�b~�?M��\CY6����0=a�X�CID0Ϗ�'!"����̖<��ă�}�8��X�ą�
ʠ��n�����9�|Ҳ�o�-o�>(*lk� �j��o������5Rt�}k��;~��\l�Ѫ�����B��A�c��B8�c��t����X	�ou��^(i�j4'�!"���l��T�����5����D�G8!Y_ڨ5<�%{��M��b�2]�O���fG�b6c�~#J��V��ؼ5lkH������L�h[�[A�f��u��Ae�&�M	cၑM�ߕV8}xb8� dH^��y��@{e]�jHo��8iZ�eͱ�p� ����d�5 �u@��s���E��P�[5���Q�4�߫oZ��J��s�դ�����d:�3��ƾ0�	�FeU-���/n9״��F��m�u��v���b����Fz+e��ުrK�U/���;�G�j2<��d�-E�Z>oǸ-��
w ?v+�!��j�D�eʑ�%�`�\r"��@�Z����י�<_s�a"�&oz��.lZ��j���]�=B��U�r��!�y-R�,i��8��ڊ�� �!��_�^�#O��ۭ�ͫ�kv�	�����t-���$i:qi���]&V�.;�˛��g���<�9�sib(��O.�!.],0���=䷘��̣.s%Ŕ�y�w$c�AxmɃ��?�+�Wkˉ1'v=��;�]{[f�����^�QBRa��gq���3��/5��6}^'�E\���Y�[i���z�^���~P�yWϻ�R���ϴ��L��p�덆M�R�LM�>�*W)�B�֔�P���%52����+f�S9jC:ϡ����L�0X���=�ĖYÜo�n�x��L=�A���� ;	oi�`��?�ɝ��'x97��$��LJUkʋe�bo�}�ګ���_��+��|b@�+����T�d�CY����h�܂���#L�5�3��L��E��ƊwV��[��2"��H�A\|~��EX7MYӴK[�I:���ʻ�<��h_�k�1o�gg˄�tg�j_��x��5L�����}5[�W��yC��X�(�mJ&�,S��l@TRd-�*�<!�&�Z8x�V&�8�Y[�����S�<n�?$����Dr�G�B��E:�P5��hK�J"�t՟`��WW5��lQfK=o/6�f�Sw�l}1�]7E�������э� ��θE���ݔ�֗y	���ۈ�6=��������d�5Gn��#ɑ��g{:͈��2I\���@��W���������ӈ2��!�+���> ��/�E�a��k�}�"C�}g�_}�X�p+dv��ne���|���o@����p��$�M�{�$��p�}��2�v�b-�_�K�������="lya�M��Uk+���
���f ]���_��~��լd	��5Xg_��	�vSa���ʇ�iN��T�%b��B�$2m�b)����1�h�sE�;Q{'B~5�k��.ż2���H/F^o�r[�fK��9'�^�努-��a�*'\J�ǝaM��[����f.KiY�	|v�F�����G��U~V��Gl#����fi>q;���qV�g$3-�����J���N�dNs��S'[,�k00�����bW��6�4\�f���{��y����ZI�¯ۖ�jqu�Z����Ͼon=�1Z���m���l\N�����������m��lOB�j��pO^qŸzq��Xf���p�Y�/-g�����|�����X1��T�F�4����ZYw��u[ ��Xʁ�N���7y��;��({�	;ϔ�����E�@֐�fR�܃�g�̅���<i:R�Pu���2ҵg�F�78���/��$}�'g����XW5ǰe�`#L����Rc�\~�X��<ʥp�
$p�Uo{���6�]�f>��e��bK���[����Q��_�%p-�6�^�m���D�=�������V�78��)9P��K��̧�F�{dD��_�Yx0���W�®���Ie�,8?�/(�N��Z��{V�σw�l��s9%�2�!ƶ��g��n��3<�Nj�x�����MT*��4�e[Ud�TG����<��n���TV3��#ໆ��]��,�le�z7��ϹPtu*=�c�{�S���7���Ц�u���sG�����-�i�����pO>H @�����5���C�	��k1_���w��E��&-�gDֱ4mbh�� �DX�D\x�����]���d58 ��}5"���R2�=Ι-�UŞ��*^��;cXY��X�ig��)�л:���Xۑx6���=�h}L�sl��Sg�7@@&E�`O��i�Ҧ f$�s�����H�V��h�9`�	��w�_���]��v���PE\s�,���0�W}�<�G�(n�Z��r�(���Y/1��Cx
f�p� `����_^#�g�hx3��L»�J_)��� ��ܹp�	{��i���C��n��2��P�/����Gw K�<�.�����ᅤd�W�?ڷT�@{��+��ΆRjW��"�y��UzP��Z&�>Ƿ\r���Wz�h�)<�Y�̃�uʬ`j��ťu�̣"�����(֒�keq\<R_m��dQ,����ȢE=FROr�4�%��.�O�����)��wm��������$�~zPF��ԃڭ���F�q�dѪ���J�Zם��p3��{�Adv��<���J�Q?�)�0`��n��-�9��C�d\t<rh�!���qP̢��x���v�s随/���`�Y�%�*�湼<��Q��!m�� �B�F
=#�Z� ���J;�	u���]���?U�!����!��f�����t�OA1Z�y��!��Hs�U�s�:d(���qV��{7�)����d���x5X��~b��!R]�l�>"�z����9��X��}0V4��'A,~$��N�a[�VI�~]4��q^$<> <G����
#�'��A☧�!�D�>z��.Q�C�	d}���5����C,g\~n���kkX	�8o�%�,Tn�"3s>&
��t�ͪ���w��v(�����ض&8�Mw�ڭR7��$���/���z��H�[d���w�u�G�{�<������ %�*{�ϳ���%�e���4�V�>j
���H��%�p���۠ ������C��>?l�ץ���I�B�"��Tv� �Y��ۯ[�2"�k���_�Ǥm�����,�m�!Y$pA"\	2�qlP"�+H�֋�)6��(&D@$V �B�2J^�<�-��y�Q�d؜������H�����&���t��)�A"h-�l~C8�||�x\-���^�;���QG��S�M7�TC��a�G�8<Q��7�&���6H��'a0U'�yF�~$����� Kj�!�?�Q�|�����U��s>�#�k����b�
��B��%���?�[�T4[K,�� ��) � ��|#��@���# VG�߼|�^S�G�����=s�#��Π���:�>J�g'U��6�Y��c|�#���>��bW�BG���3�)��+�ܔQI��jID�w��%$Q�Q�TIGN�G���V锚%Q�hQGTwGtID��)���$�RE�;��O
q�x���]��'Dy��9t̐Kr��)%�˸5$y�[��2�Svc%�a1%A�. ��1�[`y:�;��є74a�̴9@�72�2���Qe�%̘�Z'b�n��;r������{��}��}� ��7������?~�1�c����ȞL��?� ��H1�c������]q�;�^��=f>Q�S��������L���\�|��������a�j{^%�(e`:p�]6���dO�~v���H��O	��@/��}n�4���w}�ҤF�v�?{�^��5쁅�ې��l,/����\�O�PZ��o��������%���z?�Y���.Č@C��C�+CK�C�?��[��j�q�qtS���߿���B�9�>:=:�=q��9����bWT��Ы"�����z�"����CǺ����C�,�P=�/����>�S�W�~i<~��_̲�k� 19�e�K�{
�$��+T��efF�e�|�Xfh`bhY���S�����@6 A������ �x�O�b��C y f����wC�g_Տ{s��X3�O8�D.�C���)���P�h�W��o�����}O�ޮ��CW��������?W���q}�8����vï��Ä�z��ô^�to̠H?ԇz1���HLPTX\`?��[�l�z��.�������z�(`�y�h�����Cۨ���w��m��nz�&�DI�nES9�;�1��#R�����fA�N�uoHf�����w7ĳGT`Ҹ=DHNSZ�*��^�dgx�����a~�0��`o��3���n����{�1v5G�Զ�"�`��1>�1BC��0w|*��1� ������K� �a��p�4V��2loa>=㡶��MɫA����O���iH�m�u�&/���20v5S6Dʓ�@#�ju���d�DJn��M���b7�	T�f<��:���.���F��Pc�:��%�2��Fe��9��}})1ʛ|�`XAe��u��4NW�"TT��>(ZyӑT��-Z����VR
�t4F�8ʤr^������j��ڣ��e�Rֹ9g���E�N$YU��~�#E:�A1�e`1&�d�b���1R���a�F
`��Vn����-d�K)mx���_DS�����H�F�H2�2+�C�"�o�%HT�X�D���&��N�]�P�)�������T����.c��7�w�,�����B�:��`9����(��3*�+D�S�"�"�ŞA�S�9�5�%Q�O�:�w`����	d��z���̻4���j�t�5k��P+1��Q����=Fuw�I��!m�i�,����uM$r�]k���d��с��5�]c�ٚ��TAw���cf���7S�/���ƱUw���6�A�G/��2�"Jh���f�_x
7.�-��Gu�z���˙��[��Y����R�vt��t�����2�Y���J4W�NE��i&�08~�)l��-6Y��f �p>+&4)J�?�M�s�R�hFd�&�p��k5D5E{���&�&n�վzY2�b\$PS%�L�����bQJ4�6#A�VDD�O5,����&#G3�ʡ%��'3+f�	#��et9u�zm����k����ӝLC�p6�1�������aҽj]gUr�AW���Ы�q���;J��3��Z�p�}Nݙ�njZ
4��2n��J�o�24="���VY��^�'�u�Ko��La�l߄1	�h�7�U6Ƕ���уygk�y��#2_7B���Ad��l�f�#�&F��^�tA������n�u�D�r
����΂Z�КP�%8��d"�߯�Kwn�������T!�S�۪���L��蚢)����l��c�������1�.�д<�H��)6کd�x0UBl�4�"���l���Jթ��f�]�z��]�
X���F�����F����Z��I��1|^�Ge�Q�2S�]6E��V�.Z��'(i����#�?��~�ƾ���Rs�^e��0FBe~m��.g7�ux��$y�C2m�L��T	�w��"�z^�~L{���B���%�1����n�,ћ�Y�@Ʀ�5*d�U�q�/m����&�(zGz8{�@6p�|G�=��'�o��S�0������*@�n��$����T��y���i,�[5i�(|  �˧��c�����+gz�d�*�˥�%����6պx5,�G�m��.�,}�C(��+�R[p�
$Gi���%[�$M�?��(��&f�wK!%��#�rq�i0��-T'X���+����ip�Mή�Ϻ��W)�<)t\�����`�D���ߴhn��l�*HJ���V�P�
<n�@�����D�P\9M/y���m�W_3쓅L��et�ߧ�d#A'�I3%h��x�ז�:�ͺS'�A�,.9f�8)�5�s���'�ilx}�SݴD�Á҈�GI�W�&#�
�՛��f帹��$���`������Rϔ<������|���̭P��)����P�E0�coE]�`hѦo�]&ԑf�;�C]%4=�mt��(�&�Λ����z�����Ѹ*��ţw��V��u�eZ`�aA/:m���R"M�X��+��s;�����q����،��B�V���d�/�e��Q�I�z��X	���ѣ8����� �BB-�'�a��C*�g�SạOr��b���V)�a����:@�p�R���6Z���,����*f��	n1�%�@T��0e��	LeR�HX@N ����Tu;���
*�Ɗj�\]�xH��x S��]7	g�v�l�y�J؋	�
e���~D�͟�ߋ�Kn\fh�nx2UCܫ3��Vt\3H�g9��5��!-,�l�Q��sM������W�z������9x���,��\~ܥ���q����z���(�ȳE�P��Y9j�2�!5���gT1H{
10�Fm�m~�4p"F��><%����nk@��D#�/g���i>�2o���#���j��&$��W��J&��/mD�M4�h��Nh�����q��L;]V9�SkGI��&��?Cpl�O�4C���Y�T�4$����X
PY�G�P���C�P��|�В�밎��5�ӛ��&�������a����e�V�	[���C�/��S�>��]�ҥi��F{��pd�f`6,��sp6��f
V/�eo`!5��'�ib��QG�S�v9,5t��V
KctɚX��t��$\,v�71�Z�S)6��Ub*]bP@�%i.Å�Zwa����b��R�U)0�h�K �3�q�L0���|d�(7���	��l��̐z9���⧠���Z�$�έ�%�"Y0�=�j���D�#�> �tB�0ˈ��m,����W� ��3 �J!�?��7���Q�Mi�d��Łm�j��D���ˌ8A�i�Wy������:��p�}m��P.N�G�6߆��BA� �3��W�o
�������=(,=�p$T�%!��d)��>6�F�c9-)H�N��e���to��еfSA�)��Sgo�f��>h���nd�f�S�],�IN�T[b��;�h�m�2�	Eq貲��a:|�Ĳ��Kq\�j�ݏPG�Ic��q|hUH����۰�M<1���ϵ�F�Űekk'm�mԝ<�>���>�4PB߬f���kŉ����8�٦TѪ!o���xq��3��|"`D�-�,��!�\u(�;HF��4I�=��~`�.�g���%�3KYƙNS��K�ַ�Y�d�h7kV�d��UDi��	��&ƚ�$��ZR���x���Ni�$��G���]������P�Q3�Z<��^���8kM�ȇtOh��x�%'��)[�JG��k��&Hu,ɮz�)4����ۈ��s��2�"�t}�O�6���l8`+���ǼU����"���})��.B�L_�ˎ��L�G(���7�m�U�q)�;s-0:���bū�Zq��L����u�v
1�o��ߡ��]b#h�����Re�:A���^�u�&>: "⒰�X��G�4�=������?�4I�_�!����Q~�ؽ�Æ>�=@��������K����%�D:�?���:��X	�������|~�u��Zۨ^�n�V4���y{�m�O|j�?�{�!^x<��S�_��~5�f��P�r�\���CQP�~NRQ{,�e��Q�ټ��K�LCRY���6Z]\U�G3D��}��z_����V�֨�! �����]B^�~g���r���S����^������x��o���Op�>�uCJ,Y;���i�����Cv�/��)�a�ڮ'��"}k��籞LD *�8���/�/�%��H.�k
z�0�����X�f{w�o[�x�;�k��f{�
�����]�����aEW�knr��yc��7��}�|\���� 9��]k�/��Q���{I!�*�r�� wq?������P��a��g���f[��� �$v�?�����?~�1�c�����?~�7��>����OJ��~��������O���x��!.߉<��tODA����[]^����X����ص�!�?����n��߿���g���?��Rߖ�w�W�_�%�$N����O8Z_E��8�k��:�B�}.i�E���()���w�8�ٕ���@����~Yk�u�¨�}s��O��E��y\b�*h v"�`�x_���`�� ���C����]qÎ���Q�N_�=�T2Y]P�k��;FCjj���/�V�ye녿�������]P쀾�3]J���<f��$yk��s�@���׳�0~vzu��CB-(^�O���@,~;j�����~!?�����k��7�����x��������2Z��üַ��|���h(-t�� �/0�_����yl7up�A�x���>9^sJ�1�Ov�>���Y/ڿ>��w1e%k��*�����F�-�r������Sُ =����ʜ���p}�'��o!U}Am#�������������8�v��ⅿ �xn~�~���@R�7��2w�c�
���x��"���NP�8��s_߱�p	J���v�R�%���왻�
_��O!����FG��U�� � ��es�E����U&E�#52Ssa|����߄a��2��9�^�枺���[k�j	g��P3X�\�K*ྦ�(-��1*�@+��8�_w5�5CD<�������מu�,%�v���m�\TVZTZZQڡ@5��1r�K�����yK�a�V/���ˀ����ț�%�5���0j�f���Tԋ
L
�XX��P�f^�Pf ���EQP�(�ޫ��� �����|�x��4�E��!��巷312�C�Wi��P���$��� ���Y_,;L's
�~��nS�l?��#^S�Q�|�%�~�^_�E��?�<�m�����R��L���}�����K���f�Ț}�p���2e\�n�ZO������J�n��W	A�麹�Sy���ſ�� ��X�9���|���������co,�J8�t_�c��&��Q���u�V��3η��έ����]�ۻ���%�A�6�7P��}����	�?�@��_�����x��V���Wk��W�MEL�~�z��-��/Q��G�]㦊띌���K��B`d\�`�fg�CS&U�ۻ������iU�Q�a�;��h��1����>P�?|��-��ҿI�Ӻ��qe��ƥ�$�>g󑊼MK�$������@�S���[ޕy�;���{L���y��~x2�_�Z��~p����?~�1�c�����?~�70��І�\��:��"�`�D �a۹�I���r!�u�p3��Q	���)�

��_��E�9c����Ǵ�"���Ȇ�Do�����!�#�X<P�*Y�ʖ�E���Eiv;��(��;A�����}��/�C^۱ˢ�9:2;R�##�b!7�
z M�0𻙞6ER�9�����JRZ����&�K��t���'7G�������4<DN�*/u����od���'g��8|Jn-=EM������A��Q�����q11%��s�-1"�?;D*�(Z��Ί��Υ�G\-�����^���-�2�^�cHa�E19S%�n:�� ?��+��ě�x���i��	ov����/y�[��*�]#��i����3=JWcis|����[��%�2i�b�*By�P��*H�T�Z���ۈ u��TL��t������7Θ�C|��Kƿ����nN.
�|��v/��#�گ��zQ�w^ր�6s�dK+g
�~�6�n��6��OD,=��D.٠�a82��0�@JQ��)#��A3�9a�/p���t����y#58p?ef_a��=} Ð#��/�{�fS���ǃ��u� �mS���>{���~�јls�Uu�v�9��v�@�F�s���e)���5D�.d6{�o�xx{{mc��ˀ*B:���Uu)7��Ro�xu�4�'TU��yzE�ƈ��M���n�Bf�PRȲ�RiMʙ�m6$�[�~a'�z��3�U4|A�"DS�-"��8�1f'�eo�������Z~ܸ�¿r~G�k����ln\�P�w#]L��@XQ=���d��M[�[<2I(�=�gj�p[��D�r�Pk��iB�1�٧b����eq<q�W��^�|���Y�8k޵�S��t\u>�~ǓA�Usz��Ր�w�,۝n�n�F�&��ĥ�����ޔ�+�h�r$�R�Y�F������#���&�����U�Xò�,�b\$�T�|�o�T/�kc� E�z�"{�pzt}t=�kŸ-�D	/���	��(~l�Oy���x8�!=?�=�29b��XPBa���1��1�5�ۿ����P������ ���O�܉�3��f�j�t�ݙ���:s@�ƈ��}R6��Ks��c�@`ч���.v�n~S����p�"����x���'���ٙdU-)��g���Q�0{���D�ўOzq�X��o���ҫ��H���BE����/��Y�A��]lH�A��"�'G���d���i"%D3q�G��9�����CPb�0�&�	�h^R�h�����O3���J
)��|f́�w)'6A��L}Uy|E��b�!}K��j�(�1��G}�K�d��ge��w��`�`.kb�m�n�E�b$����	��(1��[],�[��d�eQS-�m���,�!���ٟ�P��լ�IJ�!uR�d�M�qp|v<�O��ܦ�&��L���n�Xf_x�٠GC��;��w XS�IS��	�t�B�֨�΋V�e�����Ď�dd6/�q�����W%�@s�K�2a���[��&�γTN�*����%E=��7�o�u�C�Z�G��Թ#�%M.RJKu�\�$wC���q�s����0��*��	���Lw{0s���p�lI����:0A�nx�>G���w2Po+�9���&t��i�f�H�p�*%�}�\?�����n�{�g	�<~���B�hO��L	���zf{���S9�cМ�1�4sOn�j�%�=mDZ)�1�-���t�j����ch��^fYz���[x8�ƦF�&>��|�;35FW?5D�s�('gu��`쫄�c�
�|l;��
9���C�� {�@@��紅�굊��4�[�a�j�WM����|Ln�A�DU�4�E����CZ`XC��#V�C��e�7:���=L���q��f��k4����vQ�{Y��`�*`�(��(�XK��uR <�Yٶ��驂�Bv^]����RK� ,�χP�{FM?��s(v�U�r~�!h�<��e��$�hQ7�=��p�M��P�8+�/�?/*��rG�����ͨ��QQB���LҪ]�I!)�F�L_t0��[Tdc����4��szFΑ]��n7ͧx5ۨ>���ORFw�9Hj9�S�@((���}e�O`�3�.K�.��ƭ gw2���l����T�������69EZF&L��w�[�|�&�n!: {	��)J�\B�%��f�irN{��#;� �O�=ES`��j�KX��NK 6`8x6�)ކL�(\���YKTF!�i��QM4�����Ǔ���c����czr��(�L ���GUQ'�����k��h�n��K��L�$��7��Z)\��;>��pK4�>�>�&�4�nds�F�X��#w͡�ߌ�,ۿ�9�����.7�.GrF��o^ʼ�`5��I�Tczf�/�pҒ�!��/;�	�Oqmc`J�l�g��֧7ѱ X��^�m��IN��B�^��W�Jب��Ş�i�ho�"�v�o�ѿ������ r��:�~Y�pX"��a����UJ��X�-:�T�QF����=>9Z�rL�v��SS��>�sW�R�&���=$��պ�A�/��ʻuX���B�[aH�����%.��<�M�IH��%j�OH|CP��pq䒢h�]b�B�f�{�g�Ԯ�f��V;�f6j''m�GG	l� � X���a7�!���s�~�S�[ޖ9\Ȱ�B�a
$#tE�k8�aZÓQ�-0�A�}υv�rgH�k��:�K�rҽ?�S�ٓA��mZ瘋eT�1Bg2�ǝ�4���j�)��a��\b�HF�m�e�x��m 9�	
�#�xk^R�ι�(��Q4�������(�����S�O��:��fhȕkZ$��K���>j��恨���j�E�X��m�*<B�\�yNj���n�xB�,xT�~6�?JDcvD�D�<�]�k��$��34P��6GC��\�b��c&'$���1��cp:�~%Gǻ^�%�-���f�#Y����+q�L�CqS�ƭIm�W^!H����jsm��m�,^��2�1)"` e*T���3�5k�8�T����A��Y�]�*[��3ƻ|�W�¬���0�w�t?<=A<�ڡ0�$�
,J�Q��3ǔ���7�t�܅���Å�;�S���8�`ܶ3���j8eH�rX]U)8��T��ö?3�t������C$��ԏo{���N3tk��;?Dޘ�εS=����+V�������H�h���6�.]*��j��t�t_��TU˩��$���?!\���pʴ����Y}�}�q�1��U��r_z�C>��đHxY E�h`��ۿ�����.���I"���N�V�ͬ��xBɺ^��:����;����=�@�T�;�gC��v�%Z/,���o*r���F\DۦZ�q�Rֳ��۷��be*r���k�,/>�l�p!��TƛGEo���U�gj�y��8�4�2�mc�h���}=Vu�^�bKr����'���>�0/�x3+�� _��]�<>��'��u.[�@U(���];`0�5�$�O�+������Ӫ�nsHx�����KR���_[��ZMխ	8���4���U��4	����8�0�mѧ9{q�ӧ|R
��l��:~�_`����7����vxob)X�&���p2|jNi�Յ��?6��y�쮛w�������"!Ռ̈́� B B�! ��E���zB����R��e�z�@�� �RB^��������ŏǛ��z-�E���G���2O61f�=Hs'�u��N�Aǂ���ǀ~��$�� Y!ȕu��h�����L�Rs��|Y� ,~���6��<�e�����+y��>��D���N3����Am8i��	d��5�S���+i���< �$l�s"FK���o!��z��i�1���&�f�h�aao�3���,�_u����_�)�?D�ື�x����w>��#���pŢxM��Jb"s�n��	P^a����)��pW�b�lݯ��L��:�SR%������A��^ӓ��7O���fA��5�ܕ��!���s^q��N��L�ćF<�J�����-�;���b��צ� �M�]�r��,{QI�$�[��������Ǖܩ^q���\ ���i��M1W�rm��<���qʹ.�p~<̬ΰ�ԗdg�FZ���|�!�Z�.�Z�����Z�hZ�P��s����?���秧I��^aL>x�C*6�ؐ�A!u�H�#�:0��ťg�'f�ǲuجf�#'�uI_����I��zϦ�a�;�����%@�U��l(�Qª�<�=1݄%I�K����ʢ��v[ [)������Ṁ�$^��O.��Y2L�@ߎ~[�_n``��d�]/�����وW��R�+�����XO��.�r{��!�e�AH���D���	ϧ0��3o�
d�GR�T$�X��Hy��T�vi��e� ��=2;�M�Z�3>�%��IX�� w?>�\��If��s��|�`�}��`�
f���B_YN��k�j�����O������e4{�Í�msJѡb�[O�/����g1�/|e-�w��X~�j<�(���e]G��N����-W۱k��,QsZ:s�*"'a�e�˔E�a��::��6-Tŗ��{�~r�&諮yDBUe$k���ٛ4�ٍ�wկh.��ld����yv�S�F���.���umTR��GЇ���gJG��]��_֠6�4�qV�S(k��k)�/�`(�)"N(�^��	�Pu*����j���S|inǕ>���=��tӴ�����5�����p���Q���:c��Ҿ�X�����؋�jHʡӞ�O����O]X]z���l�yq@=X�Ц�4��D���9�Y�
�ȘމZ^`}��]iq����|}T?��=��`v��xP�8��W�:���JG�*��k���\��~��
�r��Qbk~!^�s���e�+�߈M����M�@A��ߕQG�J�u5�|Z8�&�Lz�\kE��A����A�A��D��	M�jhT�nK��B�}_�(�T3��&��:���>�N&���^w�b*BV�v{�~�sA��^.���==�_,]�h�5|P���7�,S8��p6A���է��e�Y(Im7ෲ�����O�r
�8��R�%]�ZY-���;[k����MH:�u�7wBɋ��C���S�%
��f�IQT����Z��=P_��p�b�(IrzDiv���'�A�<�	���{Jw&3�}3sB���^�d�[wa�d�o�D/��x�b�>'o�Ww��lgK��`~ᖻV�DUd�E
l}�\e!��K=C�����o#��|ɻ[?�p�ۘ�i M�kr@�u@�k��4xHPPS�עrZfN� �%"S1�-����A��jf	]�(�C���ʛ�KZ�NGH��~^�(�M�Q��&����lk�x�Q�γ�f�{��h*�9�
�ߝW�Y���]< �tӃ��Zy?t(ӊt�
�Z�΀�n#4��R�{�j�pA�)�6��{��{�a���re�����x�'6��v1�:��Pk�&�#��r"V"���c ���N�7��I�YE^�k�SS�Cv<���b��0�y"QA|�4S��q��\�1ԔÊ�ǽ��h��{�D?�r�h�,e|����
U�qCŅU��6C������K>ò�c��*7%֖݄�j:�0x���l��z�kX�����%�#���]o���� {�]�ίL(�ˀ<��:�9��&�{IU����e,�$����V^J��:��Z���1��+�a�D[��牛�����%�鮍�i�|��4}�ʆ%2<
�K�)j��k���[2���n�p���[s�w�U�X�¢N�h#r��5��1�0���<s�K�S�Y�Qg���!,��A�ʿ���}��1xs���+�4]�4�Dj:�J�f�����3hF��t+����VZV;|���-��)�ҏ)�V��~�S��z�q��:oo$A�Z���%~t�߁g��zI;�p�R}�[�/죷����c;uKU�aJ`����2c(������G3>�6�,'�����T���FzN<h}��q��t}��
�hJ���G���=l��'�F�(Jɗ�iK\���o-3�B��L���^�jA�`��>�e<�6��i�`Ëe������bORY	��P�QD�W�m�&�gƾ0,�_ӄ���AbC;����:QU�9�*����V�pMʞܱt1���3����a+Iu��K>�n���[HI��1�����ب���eM&����F�0����HG^θJ�K���#0;^(�U�GL&S�z�[_���J�HeWQ��Nx��F�2����q��G�k�?G�IC�4h_+ι��0*�שZ�\M�۹\�޲�vuZ����2�O�[.1�b\k!Q�?��:X����*.��jv"c�>�����1#7Uh����/#+x�2�Z��������c�lcC�%ٿLx�t�U��דE��]�%�=����+*��:|��X����ǹ����\΁i�1�` #{M�e�2��>�V':��0����]y�җo� ���W�T��?|Q��.q��3�_�!v��#�.�x<xȻP�x�xpȃ��O�ռ��p�N_٥�v�~9�bk�C�%�	8Uޫr�|�����A�b0�ԫ��UH�F�5��E�f8��8�]�>#�ؕ?�D��}ZpK<�D��Ѻ~!�3E��J�w5�hz�D���5�i��[�{��TT�4���Ax,ֶ8���}�.`�V#����W1(��)Y�����P��=���Ѕo�j�d�9_����1��޾�y�_:��;�9�ͣ�3�R�TQ��;f�c���=���+E/?]X?�{^�=��V �wCa���c�aR�ş]��JoIb��=��gX�98���������^aH;�S��8��3M�\�>�Q��.�3g�ae-&�$�œ���z+T��~yHU|4�i.�o��K�����O¹Fo/���L�a
��I�j@%>�Q�J��ꐭ2��	�����Nƀ�Ω���h1z�a�ǁ�Q���5G�����C��ݻ�F�$��W�mO�뫠w/�oP�1��ˬ�U�z�=e�*U�q����I#�/Ͷ< Ծ584��~������B���y~k� ٝaws�Q>���|�W� Ǒ���bN꿬4cI=`����fT��e_ظ�F)�����/KV��=0�&��o�F)���h�gg]^�;�m�G�-RE�z�ũe���:�X-���e�V�2���4���HJ���|`�rպ�:�cO=���W��N�`&u��z.~#��N2׍/�z�}Hڧ�V8|z{�["��`J��n{3�U����[����i�M���&Lx\��:��d���>���,u/����ni��m�
MŒ���Qj�"���0ǃ ]$����ܽ�}lg��p���f\��M��a�����u1�F�(I������5>
 ��ETzw��	EY�G���x��qߑD��0[��?aŗ~3�LX����peb��T�1�<S�����K+4�m�`3��c+��ǅ*�${��{g�E�rL�K��QɎy�=�o�Q�Z ��ٷu�s��zw��L�Iu�;�o�2�z�8��������1+��=Vr�g]��~A�ҶE���f�&�'��r6�����rv G�P*'g�`=s����-^<&��yN�W-�O�=��BU�'&�Ux��(X�Ƚ�1׌�vz6�l䝴���_q���߇�Җ���&�W4��M#:�ǩ��4�ce���Y��]Nv���\�ێ�H\�9��IX2��7�9O�"@`�¶m.��k{�׫����MV~�^�y)��g��O{~S�����=�T��b�9�޻�TW�?�w���~�����x��7�|Kݨ����E �k~���͛iXGtL޵���}հ+@i�a�3f$d������(���O���2rw\�tӼ v�\(>G�k��ӿ������u�'�[�4aG���Pid��8�;L�qg9��D�s_g`5���-!�L���.à��N�q��6墇 )��,�[��{�yWč8�B��ٳNL�J�QA^����J��y�0�N��Qk.��'�Q�p���V�CB�����[{����1����.Zb��{���;�Ln�Isk^��Ӕ}���Da��~� r�Ղ����1+��7]p��r,w���=�e��9 �a|8�1���	O9�V�C� �h]>!W������c�Ur�
3���㗰��@j�䝓���q�h��@�0{1�{"�JJ6����L�t�~���& YJ�}�S\,�?��Y&5���w��R�Mw��@�F˽Z~��%�oV]\}�p0�}�=��N�^�a��؅��;�x�|��.�!�T7c����� ^�{O�9�F���_x9�Jf�d�:�V��o��/���=��ha̿*�e�-r F�nk�e~Q�A$����-?E?\L�˘�fxM�ӣ?@��������&�K9 ⴰ�;�a��%%�d;�&��J9[C&��[���BW�h?�������$�5�L<O���[f�K��.땙� 14j*��W�v{0��G�����ޙ�b�K��p8��ܑ¤�X$U#�ȳ��0�}��B��3il��ߊ	SU}0�阅rl�}q��?�ؖ�B%�KO�H�,y��#�'��6����8�Ӗ��fLfX�x�N���o
�HF_$������7h �d�_�e���|�0��B��Yh��Kρfwl:V�:�'@��[���HKG��E�~���Y��6��-wh��菪���!��)�L��-�;�jP�ɧ��ͷ6W��!�lT�d23��[�CD��ؙ�r�����@�$���[(0�E��|�AW�;���B�C�-o�G/�I ���ZS�R�!�Ie�Ygo��z�\��y���m�ݔ!a��bnb��֚�l1�+�]DB�����
�IL���Y&uɖ�Fw�ߏ�3u�:v\N�}�P�\7&' (�,����('®ݚ�qz�K��HWԳ���#Ә(I��� �6�nw�i�6wV �6@�\=��u��g���˞���̐c�����Έ:fY���1c���ml�̼9�Oڬ+��y������x� �&7�-S�;�|��ME-^�B3k0S��������썍x����w8�̇M��"P�J��e��ewcOxt�A������W�6|�8,h7����Y$ܽf}�F_|ȑ���>,�0�#�l ���,��sv3P{y�̾,:��fKO�eO,������S8���ܬ�:d�����o��}�T���y�X�r-~!��`@���j�*Э��h�'�����JJ��|�2�y�x8F��K�uu��*�|��P��8�b,P8��!3�?FL�g��)�yz/ׄ}2u�>TS���+O}�V/5�� 	���P�����r�̃ײx҄Qu���?��ؑe�h��@u�R�U]���Д��~�]��(�H!	ͪ�R�$��G�`�KG�߸$N�QM�g��W�A�L��$��Ty���tpDn?r���_�w<�N�>�d�j�#�H��ᨈYikk���ӽA�!M@-�{Ǆ�F��
�Brb�[��kFe��f�T$�S�2�%enR�+j�*�>HO`4̩m���q�[���2�w����B����Fj���G;h��|Z���:�D߶c�-�R7^�^�8���h.���0���LQ�%��t��Q6�Q�S���FQ�2�k��cz�!��~v	����6�{!\��W����X�7�P<"��Ȁ܍e�AM��f��~�E�ޘ�.�&�|�����# Gw�+3E�g 9�g���&��2|��`ח���s~?�q5إ*[����e>�����V2���d�J�� �7v��a'w'���p�����{e�U�E+(�#>�'��}��Ծ�[�כUY�o���/�'Z���g)yV�z�K����Ԥ�K�������SNbH�`�hXB<{�RY���a�N��t�ԍ8�)��)~>���F[:��|?E߂��������媛����-'ݑ����`��yy����p�빺פ���� ds�i^��d�����>'�u���{�&�rr	3��EN������K��^���y�J�x�T���01�Zk��W�����1U��;���u��(x�VI{�<*X݃0�w��;�ȡb㛑�͖�M|��]��)�ϻ��2��C�3�x*K��s��]�91;�x�X��2#y�?�=Ag�v��S6���*�>��z�����{T���G����GA�eE���-�{|k8�R����FO`v���I�]an��w���Rw��'�*^kVL�V^YW,�V�7�Ry�w�k''=\��Q��q�%<^v� ��:/a~�휛3���Z�����l=M�^�+Vُ=�-��!��G�e�Y,F���|T�Z���p��+.K�����uG6�%	C&����4l�$����^62�h����~W?��tߤ�χo巸r	�2ߑ�z�B*]MD�,��nׁ��;���L�?��+�E�S��K�ˏ�;>�oN����r>������[����hmq`+`je���"ӭ7˒\�ͰD\�Ւ�B�qun}��?�����qq�Fw���4-��#w�|<��s��,��gp���j|��PH.�||�^@����,�0�KM`�cv���ϧ�g��H!ޡ�򹇍��<.Qsܡ�uGi'6Ѫ�m�d�i�/�R�]���8�͎��χLy� *��п�]4Z1�KHIM#,�8Y��B`*B�Ԫ?쩽�[=!��8��X���Sk��'3檈9<��ބ[�vg��Wba�Bnk�����spM-�4�$^��~TO��4��d���s�;�`)@}<��٫�{�A��u�$�0�W2?�����PΩw�4���􉶼�}���F�8c���݆�oTGoKS24H�ܨ�q�m��c�T��� ;_�ސ��.��˺�u��SQ�T��/�M��"8C�����|Ͱ�mW��IJ��&e�Z�?���m9=S������]I�L���N�Ę]�{ٔ��~�%J�$�I)�C��ł#YVVH��p�g������6���h�L`Z_���	!�vbwsĿ��������)�k�.�yE!�9�Z+���sn�9��1��!V���:-ϱ��5C��+��+�g�A��tg��D6����
�"d��H΄���Hal�e��A]�WLL�8�Ƿ䘻o��'B��_
y��o����J _1����_='����Pj�J�j�"�5�AT�{�K�V���f>���ֆ;5G*Kwcl6��r�(�5���_9�t��x�:�ߤ**@L��wf%��K;�{	�a1�c�$�/�.�T�!��훛~�Ŧ����GU�����J�Dmюv����6�A�Z�)Uj����@�?b��tP�O8�>�FY�]�2Q߀��-Ia�a�@�������t�\=�]hKѨ���> ���5G��'�}������c�D�u�h�r��v�k��Jq+�p�&�N�5e[玬lQ��N����S�%\7
e՜E���Q@�3�.���ݚh���.!_����OH<���-s,���¢�5��;w©[���GC��"�pj��ƤN
p����G�*ϔV ĸ":��PÁ� B�1���y�'bDB���ٔ�7��FNN����t��m(B��9͠9�m�1gz�z3'�K��)G9���(��2 c�ę��ܘ��7���-.������,4��L�^�v�8�Y�^��!�E��.O6t��}��?��Q��^Z��'�=b�b�c�/�K�H����������d��dL-)&�����s-GH	��BС0
zI��Ã������g�,�]���k�����3�
�e��i��Ѕe+���J˕U�cA
�M�dH�d�D���=5YE��=�x��>&YU.��;�9һa߅;�q#�6��n5Q&Px�8��E9׻�0���۶tA&��?Z�;9k&�
�йޮ��.g��0c���|���d���@���J�6�v�D���R�mM�FOv��]�?��}�v�Ԡ�,&�!ly��Ic:Æ鴉�"2���������x�|�g���9J �F.�΀OD����,y�ś͚�eb]�	��O���߹&��^�l��	�=wit��2�4�-��r�@uq=� AA~~�s��'�K&20w��DΓ�p��h_2�qtH�q#��L���O��g�Vj�o�IU�:�2�z_��#�:���|y]��^~����y�?�� ���$���
�K'�;#?�+����)E��a��DmL�"R�!�fvg,�8m�˙3��A%�Q�J$1�*pE�n�P��j. ��DBQ5�+
"�`�8����@B�:"9�%�#(���2��#" ��F1�2�1B��1�e���c<ְ�[<lZ_��w��Ｃ���W�.���U�o�=�+Au��^����)i�)�<���*!�$h�Ġ�4[��Z_����¨�w�4R�Ǻ+�z�����H������?b��43�
����� �R����ū�4�ݹyN�߫�*�$�N��-?&�<���ɨc��[��g�Lٺn��M��T &C¢�f�r��Z�m�R�;/���|�R��a���2���e�>gR]Zt˂���?�3	��˧�-�w�El[����x������ϼo���OZ��F�b�8ƚ���:��HѮ�/<�#d�v#�����L�Y��F����ǵ7�
�`l���}�8@��V������i�I��m�D��
��"�7e�VDL:��^Yg;U�_{H��<z���t|�Aѻ�>,����;��}���\.�`_a8=�F��B��9��t���F�*�@����P�⿰�a�mr��W
�tހ�*��>[���h:Q�4L�M�it�P�t�n$�1J�T=Z��~E+o��nF�!U��MA!t۽
K@ˑM��s5�_̵e��t��٤Ζ�>�y�!�9{�lG�
��(u���otY��J����Wω'��wUW�����oj �_�3h*説���s'nчrJ%�-����>����v�>�ʆ�v�����l#SBM���]� �µS�OE�m�d%�?>�]t��Z�8��n��-֐*��c�C�⼙�T�ߡ-�%��Dw]�k��m�
Q���1Mgn��V�!"�Wocb�c�ݚ��q�ʋ|Y�?A�Eε>o�:�S�X/���t�{l\�3�D�L��6��c7~�
e$~:/����K)����SS��6SW��6_�.L�4}j]s@�5� �]�B"X���f���1@ ���N;C�7�3;m��m,�M�l�B�;�`}�	;�PKt;�PZ42�ܺ�sd�Z[��\Z\"�Fh��E�-���f�IFY���ٿ���1�9�f�3���)l������-���}�������a���s��cF�d���Q���[C�.n*nu���{�W+*��-���c���a�^R}&�\�1#X�o���ȣb5�j���� ��gP�*��g�s �A��nh����Ci��yR�֙w�$0�.���2�D
�U^�.7C�iSD�b��}rv�?ux˵$(�FEuv,���7z�* �y������M�/�{u��I����/��S�� ��T��� 9ʳc�a_ ������|d*�ԳzN��3�x�~,w�#�Hf��8*W���^�#������]w�$	5:nw~X�Fx�Ĕ�`W�����5_Q�ON���h�I5j
2BV�ȓ�\y;�p��e8����4�L�\�d�}Ȧ�\�Z��y�r���d��ă���|Dv�#:9����ۭ�>l]IL�,H�a�'��?"����3P�s;wqeF-�/u"�K��6v)nLdks�|�5�I.Y��ځ B�v�}�nͿ�q�������ٔ���|`����<x$��+d���sd��cU�s#O��d)z sb)��ȃ��S��|g]����+@1@��N�X�Z��ȹ�$���k���.��1��FOg�����0{�����0��wQ���2�]��:�&�k�x�]hi2���C�WG#�
RyM�:�0i����,�)&�G�X�)k�O���x�N���J���&:�q�Q�1Ziƛ�'�>�׽�ߥl�Z�Ǳ�M>��I���ʳ;]7�.�a�BΧ�M5����?a��:�$4��}�j�P�h�i�&-Rh�&UW�#��
V�غ�Z׺<G�aׁɓ-'B���+{�ź5;gajA��c��`�&�&ܘ��'ئ���p����-Ldg��f~�571S�}�6O��fum���i\ٱ��1�(��Š����Z��zn�>�&�[�]�xe���\'sH\ ����e֥�;Z�|�IS�(���sꭢV�M3p�'�2\|�`�t�q�A��.c���bF�//��!!�z��k|�{� ��.d�`�[-SZ�Pp�v6��\���\��� bN|����]*�����U�H����z�pk�jo\:���y xl|��>?(z	�B��?$����5���;�D���V�P锅�˥c�ߏ��R3�I�����;��2���H&��,`�.�#K�i#rwZ����M/�B���/�x��� P��ܴ~o$�<��;b�Q\�Q�D��RKw��}��S�F!T�=�
{�;�A���g*h�En�RR����_b���Ǹ�W�!\O?�l��Ja���Ql(!�zM��6�]���i���>0|E}��O��ЖD��������V-_����z�i��B4B�Fa�I���Z��X�l5��Hp�4�읡i��6�DӘ;]���؎�������G��2G�Xȴ�m)������c���e*�E���.��/��h	���SS*�dH�'��t{r�n�B}���J�}f��$A��.��kar��RHȗ\\�\�ǒӣ�O��
�!�z���1�`�~�ְ:}�>{Ir�=A= F��a��Cn ���g8}b���Ał�	�*^`^΀����ʝŗ�����J,ȞD�2᪯woB�1��H�e4�x���Æ����u�|�4 O*MBK��5Jb],�?3	\0����j��z9��	Y�yӲ��(��!j@�U/�mp.��n��J9(o���+��KL��K�%7�wň����6)�O�𮱄>�����R���CUr��]��"c;M�_	P�tȄ�L���Z�F�ockg�8���=�\�6����\\�j�jtӴL@c�1��44���%*% ��' LO?�y������|U�|*�x:����o��Y��m)�n4�9,}Z5��J[���wo��׋�tV��j�8_��c�n�)á 8-�d���.Q�2VY�¡�߄d�(���s�s}�/��Ҕ6����]rx�gL�]ܳw��,�m0A�U�̍G}��Ӱ�j�G�>*H���,���c��	�x�ݓ��ޠd�5g�k`������j2�_��C����_(��RU�����Ň��qRXSa���h%ܤ�n��ɥ�Aw<:�ɞs�/,����-��b���cO�:\A�C��H�_Y��y�tN��y�q����b�0���m��RDu�8�Q�J-�D��e�^ƣ[�@�x��Yz�\�sG;�1��\FE����]ɑ�b�a�wKF-�t �3r��x�"������#Mf��"''i��r��:���;d�"��w�ʤ�Ny�ђ�5/*�x�o�,���]��0F��YR��m8�`��)%��<��+Aܒ�7jG��Zk�ה�ݓ_��w��m�k��ck�c�_lcB�Y.��:MWT��7�3�ڤ������`R�&��r�p��O���~/�Sğł��&M���"s��V�nl�>�#�e|dr�z|{��N��u�rΨ��h�����lN����A�}�;lg�rW걩�BpIm�ɖw2��t3�$|Ə���x��3�w�Dv����Sr������W�i�����j��:�g������? ��ʞ:~@�7�2�\��V�kπ�!i@x�����>:���i��1,*��E�$&��1'~�ʲ˯��g1H����Y���IW�z����J�ֈ�t��zq;��1�(|�N�w9�3��h���(��z��6�'�r�=��w�*���6ֆF��¥��)�^���-��e�0���ˮ���5GJ�V|0xv�s�f�(wԖɽ�5�2�ϙ�}�|�0�5K�vX�Z��,^�I>&~�pSO	Oˎ�N[��^l�B ���D��vJ��~_������q�*�KZ�-��/K��Ԃ;��7{����s,�L	��"��;����fB��t�~�+��Q��z;co[�i�ݭV��C�[��#s�)�����3�8����(:�.P%�eN�	��������-�e���t�H[}U�P��>�����z�8��Qa(w�86��4�PVʝ���lI���2�)|�bC2G�C�YN�C龏�Qʴ ��zA�@�m݂"ex��'v���g���_6DA�jNeP��q�3����RGW���9�Sw�_[~ы��2�X3���b�	��+��Ƣy�5��PTp���� k,,[��5{�(N|Sa7Y���Y��+EQr����I��E?�"�U�9�����O��"�f-�Y�ٷ\�wR�m@���g�k{�pe��1��Z��h��w�,����� �����Ŕ�I�:���F�Ӯ�1�D�?w�VF�;_�#΃��a��r����2n�ݪ��6���0�R�#�}fk5���wao��n��Z�D�>�p\eZ�ؑ��@����"̉�66t���f��-dN���_z,6��'Q��P�j�+�h�
�����h��(�X�vm^h��+-�\q*�>8'$A�O��	|d��Qy���##Y{�oW�@��;�NS���]�ŝy�G�Q �lϙ��"�ߥ�滣��g¿N�V��-)��2�����K�bD����?}����UÃ�;/GIύ�nr8,��L�*D&� ��ι�>}�k�]7A��T�<�t�<W�AxWR�H���Ee�d��&텄�r���UK�*�I�	�>�t���۔Zg,.8e�ہ�r6�j��#�'i��1<�/;�]Ǚ����X�T��>cdWb �2�El�;�!|��3-���8Eզ�K�FLg_�^����d�vh\=�PF��:t��b��kת�oq�p���~�|n��S^�:�Zv��˸��GHRO4��0���}	�C5�'�	,I�ك9�BW�6����#�`-�S6�����i'f�
O��=�!;úK
c��J� ��(�Ժ�����i�反Y*.A�}R���O���?�k]�ha�/-S5�/D�p���S��X�B�~�f���a�
��8/5g�o^�d��=��WZ\)��ia�9U�nn�<�u�IKA)E�͠T$�������%���@�A�E�Y�6ƐW�6��%d�Ǚ�ry��\�WFY�����<���,��N0�� �25;&?73�R�dPՌB�FqF�ޚ��T�!����2 J�CF�K�:����®�8�^��p�:�7���P�����A�;��ur�,����RT'm3	oԏ%+ҵ��n�ܢ\��%D��F��H�'�}gozt�@	0p�Y�����x�f��)��gf��k^Ra�±��H����/�r��]`���ܖ�~���i�*��i���;��k��2�P��#�d�B+`uKCv�0�-�,9�u�inO��z21uF^n���R�Ra���rFM�"e`�w�]x;	d��HOa�cn�m��ƶ����c�*����q̏�w����-�e}5[��O�:ls�a2�bx �	��g��L�<�<$8�#ƏJ��8hmJ�λׅ���L�f�(A���~��&�I��p*�
R�R�J�\�}c6�.��C�m����7O�'x;̐ӌ��uH��Ze�m�(���_�>��Vz3t5H�:�bŴ��\�}��ۉ:�||�>|����`��!G�!b)���8�E�m��7�Ĩ�F��Nf'��_�9�P�sq���k�:�$t�-ߝ�`��²�@KS):'�I�:�ow�K����p|k@���$��2.�� uJ/m��������2�P�K�&,4��A�v�=?N��*� À�ތ�܃[ߒ�#��}�]�ק�����k�YYi�S�xi�������ys
�:�Կ4�P9�����|���,�x*jl��ح�K�N,ތ'N&!�*�l�}G�X����F�!��Rd��osjs��up-x�7J����In������h,ɷ#6`��{<�"V"#�W���j_��k�q����4��*������g���V�{8�I&I,�+�����6m��3�"򿴛�N�N*�G'ZD �|��d�v���a��dTս��@��z6j{<H.{rcI�3M+�-��ȼހ�XY���u�l̙
��B�c��H#;|���WeYA/�Ô�Ppݚ����S/\�T�#4p�(<�:�����۪�X��6/����	�R ��q,&��>�nEo.@�d|�o `|�p�!�C�L��m�ΊY�LA`;���X��LS�C$�y�Xr�̳y�\\����/�SRm�3�pTz�jߏ��R�7(|�~KPiv�;��Ӏp�:�O�e�Y���{iP~y�p�t���m�	�\k�#��Q��JY���HF��ÒI��]Z�(U�1�Ȃ
�J� &-e~�	o��GT'+e��$�1/���=W�&h��c�.[>n��&9�m���a��'e%W�vʅmn�*���4�`�w��Y�UH�LjJ��^[5�QBz49���%�{86�g��7�����&����7���..�&��a�y�-U�Q�!E��q���$fvG%��{�h�].N�4���i�k���;�o��yrry|Q��y��ۣ�z�H}GX^������� ᎞T�%T���:��bf�z���7����l,�x<�a{�^� �0A�!�\
U�}ijBy{����3��{A��C�jޜM�Ð��5�G1�[�E�/c&F�%�e)1�M{Om�;�7мUM�#Én�:n¬����?�+� �\�PQ��g|�}Pޓ���w�3��h�s��9�6ܻ�.����&;�TF�ki>M�&��=V�2�! �u��j�h2��U#�SN�V��#Ӊ�,���2&�����f�������_3'���� ���B)�{x��k�4����Owܔ^־�F'�z�~FX:L�����\K?ik��d�7C!^��I�s������������E�����} >��G�n!� ���;>���P�>+ݡ|���\��@���DG�"p�R��5ހ�=ꥨ.�$'#!�</��5�k�AP��/=��
r��E��AK��+*��m�mfd��a^,(�H��%�mf4��O���ʵ��B�NbA�t��h��j�6��Q���7G>8�T��X�ƤE	Nၫ+P�;=qLL��6n�~U?}�O��X���~���@<�g�;f�9��Ȋ�DXtN2DPȴ1^5�c�vV6h���7Db��A8��V�:�J�� ��!S{�!���1l��\��i�+����i��O͋S��'�_�*��c�JT����o��z�!�2,,�a��<�}�b��s�����^�>�@1٪o�Y�
����Q�@ō���z]�����Ζ�b[s����&��b8}� s�3�ϋ����T�n��ǖ�i�s�-��Uf&Ke�%.ۃ99���ns��<PK�����������r�
<A��J�2�爊N=�!�t����K1zc�&9nz?V��ѠeP���ɳw�T��`	�%�7f��i:��SWa�('	���Fӗ��W��)�c=��4���B��V�>ީ��Ьg���`��ި�����͒��Fߎtރl��Q}�E�l��E΍�S�$��ˤ��T` !�Xy4��ȏ�{�)�6΄.Vg��˶�D�9�r�v�qr�a��R(��ݔ��̰>8g���2�ﰠ'�>���m���j����"� ��{m��m���0=�&�諧E��t�[$��7C�e�������4�~N�a�B���K�l�������-y)���l׫2��n�����fdJ�޽�����@�+����ЮQ���}X�-��'���h����E�g��4/Ż|��ߤ��F���V��m?�r��RA���� #بY�N�O{ޫ��-�^�?�"�y��-�}x%�j�(��'���y�c?�J2�4�,^�>-Ge�����h�!I�m��`����h3nTR��?ٜ�{H�d��\uLA/3]�v��*����Xb��@Q��'�2\�&h��PaG�����z���a��h���D)��]X�o�����F8�u��I�H=u~�z�81�����Q�P�_A�$l�l��7�����(���wHW�:XɃ�\�W���(���+ۧ�4���ʷS��$�.�}0XI�Qz�֕S=z�Yb��"**Ȋ�:SC�����N�Hd{�(�p�cG���FKd�z\�P<�>��Y���Pt.SV�@���W0M��'`ԡ��&�cb�������h'��Od�373���������5
�ꚪᦨs��D5���4�#�+@��pU����mr�&�8�e{��TYv"�*�m<O��Y9�gHU����l�b}0w�]��_���́��1C�m���f�0j�Ro�n^u�'��I~������+[�J��=�?r7\������'(�QOzm���ى�;�iHh�s^S�+���uI���J[5v̷�7v=4W�O:��RT0�d��V�՜��O�آj�#H!���;*Z��у���B��z?�oh4H���*���z �=z�}0��y������*P�3cy�鮇��E���D-X�҉Ї�*������� �1�C��>b�Kƒ�>v��Oh���I�������M-<���m��d!�P�h����:�~��L�d�> �/�U[iI�1����'ոCz��Z����8��;��Cp�4���{A7��<�"ŁB�`�f�t!�Jʱ�]��p���a��.����Pc'���ڱ�1�򸩟�����P������!»�zΈ��X�������;�*s?A�	�\h ��(w�#�u_3g�ۀjD}敕��F�B=���/����_���������p|���'��=��_�����7F����_�䌜��w�/��'��i&���s:�_�	߷��E.�|�����O������z�쟥=��~W�L�y��q���ݪ���sw�̓�'�����@8��1f�������#����Ȓb���K�����������^�W�����~�����~��~���m|��!����0rC�?�s�W��l)��|�oF��?�0vd3#0 w�y�}������a�k�CH���6I
Nq������d��n1�,rk�����I~�(er����� �~l-jv)i����Q]oᇓZ����=���D��678��@�VD_�)!T� �B�	@�����H�x�ҔzX�F��
Ր��V��[�%ܨ���-THڍl�Z!	ʥUj��2,L�9[�9Gf=C���!=[��)��d���y�������>|��<�������2<�� ��˹�(��h������_�2�ۘ6�����xYB�r����ȷ;�W����(}[�=�[��x���E)GieQ�e����/������A�&�T
A���/�o�GI����HaS�a1C�Y����Ӓ{!1�j"HY�^W��D��+�ܠb�+9#4Ͻ#�Cک��1J`����^+��	[;i�4���Ǩu���?9vDWQ�tD�����.�������t�]5ɶZ�X��.x����}Y��r�D<]<�o\� vx@�_�����}m��{4�Xj�A�,p��>����+!���=���$��^��I��R�!�����-=	�S��2����|�29d�K�qYM�G��,@x��[����\�a��Z���L���h��u��0AR	3	Ҙ���e�(������&���l�%�!C�e�q<Vǎ��w�>�k�Nqa[x�9�Vx���?�k^�b}'$4����� � }%������������9b�k�V�K��(\�t�6��t��b��Z�@=���|wU���W��S��HI�M��}V����|7diY��$!]lY�C	_A.B��j�oW�er;.�U[j��aS�N�6;��ʁ�e]� .6j���f����҂�f�ݿb�a�W�bb�Z���mo\�=��n$DB����#[ٞX.��aOR�[�>t�����Fn����9z����ߢ�����:������4�s�l���&Q����ё�O�w��ւ�uy��{aA����@8�����P	�%R��[��H~�3oo|�lU��hS�`�`ۛhu�:�.UW�1��Z����]$�d����+�n/VUY�Ёlb���J��ǃGՊ~/w����!��&��&�䄸ڭ�)�6�sH�Mޑ����o����fl�X�V�}��0-v\�GZ��]9nj����	���l[���l���%�N�f,�����>/ړ;K>Q�M;�Z�랺7�;�a�T�n~��(=i�Ƕڜ?z��DΓ�3��&��&d�-`�������w7k��p�B&W�I��C�	�֙a@�B.����^��^=��rA�w@%�3�=?�K�[����hnw
��fi��S��ᤎ?�\�뇵c���;
9�7[~��z�+��}A�t/�)�흺��"'f��o�:+��d�w�_�l��2�<7�@t_�Wˊ��Ĵ���f�� ��6�B��x�-�l~���r%2_o�æ�h�m����y578Xl-9�pFk�ڝ�I�r����"��7����?Ѐ�|>�׽U`�{��wͣͬ��<���3<<4n�y�� ����Fj�P[K�z���k>��G`�3dw�a�� GS�1�a��= ����`;޼_oV�[�ڋr�ӹ@���6dX���o
I˪��B��c�x�Q#�	����
�������c��5X��kD]?�䡿��F4ҽ�?�#Aah����l�L4Y!]����:�>�>�>�>��V�n?t������|8��#��>�L��^��y������ژq{g�3B���BK}AZv��*�y�az�r���τ���2	�S�Tc#�p��w�c���C��S2���t����#�yʒ�l� �O:jې�%U2�#���XB4�	��^2��_J���Kχ�.���<��霊ɏOH�A��w��{*�^:�_/L�R�-/ƴ�W7��d��g��m	���2�����6�(V`���.~��P��-~H�zp[�9�~�Ϧ7z�"%z{a~Ɬ$�����xv+q;k{�Q�L�	m< j"���Xpa������)3q� �z
p.I�c"�~P��(�m#P��S���@~sŃ���S8�tv�&,�>�q�������|b |�|�����DA���G��-r���V���D�u��2�Q;����v?4!��'�
"�gu�V3����&���bU�^�ju���`텬6LEH��{<9)��6L)%���Lh�/�N�Y��&�[~�%\��f�@b�ob,��>�������L4Y���G�|�|�|�|�| ���8��|��/=7ٞ/5�Z����9�NW�\![N��I��a#�y2�����/����1�NC�0��c�m<T��SW�q��0Sz���^�ԉ"�
���^����w8�;y/8��j,iU��I+����u�ҳa�&���K��gc�16��W*�{Y�L �r���z��8����|�m1�iu�\�R ~;S��\�jn����@��Ő�>T="���[]JD���A���yY͍�[�22���������19����Rd��de�2v���!���inL�iw��w�9?���s��:�]��B\~`�=UR��ț�T��S�@���(���d1x*Zup��*]K�rޒ^#�ab�*�ؕ��8گ	��R����`\"� lZF�)�'I�e�N�Q:d�ͤ/�1��b:�D�
�ݫ���|�_x���H�-)�rr�7�Q����y�+����Gɬ;�AI��JG�3ԏ�`����������^=����]��N�yk3S�����+-s��k���C��eOP>��g�)��oi��t�"�c�I��'�O�xE��`���N[F�8zwk�JV����Ґgr��Ǣ��zk�N����^�:|�<��	P�nl,ov{;�8�x��D&M�X��<�b�皸�M���VG8:,�½�/`t����;�P>�랫&c��9TA���e+��IbT�[���27vI sDg��,�,��Ԇ���e�Ŏg@�ر��+%U�`��x��>Rt�+��5��JO{]��<"�D��:	�ɧ���a� ��"��^l�0�ڡ�<9�п�ї�s�U�8ٍ_�J8�����2:Dk{���c2��T�S�'��@��K��M�ן�{�������K��ubƁ�U�K�8����}�� 5+ 3|��f�&��.��	j��$��B�MJ�����0���:p����(ǯ���
��o�����8yW��p|��^�}/lS_9���WqC�h�Ǽ��Dй��n|v�b��%���pjC৑��2�>�6�f�6"͹6����Z����qw���ŶX+���g�~ӝ�� eh֫o4`��fZ���ؐ�7�Ω�ѹE�6�3�ǐ�z�F�����;��|6���7���l`]�C#*[8�2M�ɑ�;�[�g{���b�ҋ.V�z��*Q(���7���I�n�U8�6ME��"{�����z��.RC��2�c��%F>�!���\��Ys��£:
\����8Y��'A�RV�-�8�Y�wبuܣq�n6��`����Ժ1��C�-�+�ʁ";���J��9��*\�<&c��|�y�8���ҷ}�x�Q���wl�ҏ�3�m�X}�����i�*�-.
���>띃�Nv������*�os� ��>L*Uz���*b�z�hJ>m���;����{%�8�'����,'�p�����庠�:���um��O���?Ĝť�{|����0�sﱰ�@w0Y����4U6�<K��Mы
�~paT���>�������2/i����Zw�%A�W�x) h��X$�V1�
,H��Q�c�Č}��!I��D�as�s\��ߨ>~As����N�}4_�f�vMe����\�ϰVϺݦ�� �I$M0C2C��f�}����r��ڣy;��Rt��V��0�u���7W�����PV�e:x��
¡��,�<Yhhi��cMJ6O`n�v�}����P�2A�64:�$���\��1�E��r�fF^8��dO���f��ČTTTV����! ��6��&Of�W��D�����>��K�L�vs�7�χ�n/#C>|����G���M�1�|N��FP�&��-��sv.���|�(?�O��k�(�M��"��6a�O��%w��7�j˓�����LxD=C��O�{��� Y��ݼN����W4.���Ϲ���K�7�޶��!�G�j`��'�&��n��ze��'����zWo6�_Ӎ����\�ǬYp����+�����],Sc�Q,x��������s���FK.!OX�$=i#���Q�Aj]kҙ7�'�}/��O�������3�B�,��5+9>� G�ϊ>�eb�����V���s�I�S�A��{�kr.>dA�n�T��r�r��>����ұ�|�IHl�����Ч�O����8�>������R:ΐ t*�\�"F��Ȉ�����#��HL���0i]��$�a����%2j��M��,�y���p͏�e���>���#Fg�T���DT�}�������^MhBJ+��q��$Z&{�
�K�#M/���ʊ�QH���ay���ϰ[��"b�U��4IX��� s����vl,������]��2�=�Pv�F�
L�E����a��,�G3�ε+�sN�1mF�>L�	�0��޲~	�?9�=��I9/�6����}�Qg���՜bm�y����T	�ǒ�Վ�ל�IS��6���[���˽<3�r_�(�Jn9��9w���U�Dك�ъ�R�u����z;����©�"�:�~I|���ҫV��'<���?n��2�d�(��ч�$ݰ��R��
�w�|?q�L4wQ1����u��B5G�W |�|m9v~�W�St��� ���V� ���zΪד�IC^�bS��;��|u$��I��F�	���7gT��^��QT����K܅W�!=��{���M��M�޽sY�ɀsI�>
WI�����}�>0�������d3���v��vN>����w+m|����Ԇ�ڀ|3(�GGÞ>ܘ��)��_����$�[ޒ�Ծ�)��]�6D�nK���π���!ٙL�� ��^S��-=PW*Xl�s���h�Y=T��� ��h��Q��A�
#OLa@��F� �젡Oe��QDX�v}���>�巖�P/�,t����B�ċ�rM�|p���ʗi�G3M�]cp���ܚ,�f �&�2ŌlY�Gi�$�I�ے:)6b�i�Gri���s��9.�y3��]�#�����y�}w��}��]y�~y�����~�|���6������U���`�IWZ�
���j�͞�#����%�����q#��+l��JNVR��T־o~1M�F�D/��)��Pt,Ǳ��O�Z��>! ���p|��dPrpFN-���&��a���	���El�_��|6U�(e\��zY�Y$�N��4����@|T'W⎥�H�E��خ��k1�=d�w��s��J�O���=G�Z��
%�M6�lѭ3����@���JW�9*hB*�nIa�h���Z$N�Q[�$��)+KX�.��n2	 2Q��ۮY|�gm�HZ=�C)�2�f�*�c��D����֍��}J	�r�/P���5
0��xa5VqJ�i7�F��y�ﮛ�-���Y����jy�z��u%����pt���"�Ng"^��J�~E������݇|�|�|�|4�anNPh�����>�>�>���ѥ��RЙ;[����������h-��B�b:!�����KD��l�rp�7��_�x�Hjg�A���b��q�w��V2���0D�8HD�@�����K�`����`m��-�Ӱ�D��������UOߦ6A�+�ӿJ�[/q��4
���1S&D�TA�7?�O��Q�� ���ZQ��\[�q�4�c��A�6
�\�E���#\\�K;.�p`#vqp��W�s۬^��N�1���_�c_i��*͗���8�7�3gF�_�7�Ξ%�����w/���!6�(��]�T���7���1ّi��yM�W=���}6��=��:������ͭ���īk_���<�.���fC�^a���٠>�>
|ybO����q�J�����X�e<7���.)��^��
�A��K�'��R)ц*�E��
�W=&_M#-؅/^�!�2�T=���x�.�q�n�ю)����g{�9�Rm���GC$�.�ztR!�8_B<�b���v�Tȉ"�:=:�
xEZ8�.��96j\I�n��A*+�j�چ,���v���`FsK�����gyI�*��|8��	�	�!�p�b��GQR�qFSǌ��D�p/�
��W={o�>�G^��bTF����8��g9����?���=��7O���<>C�ғ9���&�<3^�	$�>%����؝�W�O����KR�L?z:���:�����M�M�͊�Ή���Ѓk���B7G�JbUX�[093p� ��Fړa~�@������ �k��P$�q �'�#����S}�����3� r(��Dr~j&c��DMY�;��@��l\}Z��g�H���H�N�GbF�ǟ_2x&J�J�,�ۀ|¤jdN!���q����]W8�����fr|��p��o�QsI}���$��T�H��9U_%�x��}Ri�4���>�}y�~P|���	T� �0t����X�	��>?��k��Ɛ��:普1'�Y'�D��^ȗ�򌙭1�<? d+�d�vf�}^mi�H
��}}D�J����<�T�\��b��
!���H�ƅp�Q��pC�'ˢbp�����~l��S����<؋��3�$B��N��p�;皅����U) 
���;�K�Z�i����j�ѕsdcU:<O��eBjS��N*h�PB[0$JJ���_���־Q��U�27\}	<�����������a�%�h\�q���A�R%����<�O�`eus��_�_��'���.]tg>��jfy�����pI��(/j�xQK��8g�mv�@5��tێ������f�\���P kb��~ /dT �9�[��D\�		?$�b��#��.u�>��3 �C�>�>[)l��]{aӝ�~ѩ�|�`\�r9�g�V0&Wg�Xn1
Rm��A����`n�
۟�h&	K{���]�|ali��td�Y��6|,a�C=f���(�.wqX� ���[P�#�Z��Cɹ,csmk��ғ�G��K����Bv����xf�J¼
'�������ACCR �Kv#�/k�T$=AN4���>C��@�|nï8��ʅ���ousuqu�:�y��̘'L���yɉ���a�|��C�0w�K�?K�G:cq:�;��Z�H+���oϗ�4��q��g=��B�c�g���Vi���b�^8�D�ev��\&̈�_G@ ܻ`���$a� 0�:긎\a���@K�NP����8徊��fPy�`/�	�E��9�.f`Y���od9H�YL�_���`�ˍ쀇� W ���aa�R���|����
NI�(���ʹ�����i���cg�-�]$���6���Иj�L��`#04N#�F7�P)f8<���o�nG3��!�(�����;�� �暕$D��&
#�
D� 5|6�14u�K� �7��� &��~���V�M�C�ia�ތ�g"f�ו���k�4��n xH�i/_[Ø,��p�.�sՕY鴛� ,p5w5�+}ӟ����=nW
K��d�D�8�%��)a�%e'�5���Cm�D�3�
��rt���1;ҳlU�Zu�Z��3ዶ"<�Jb��ّ�����B�?���|?��_ٻ����<��Er�.v�uTʆ����`�Q$>�p!�H�/X��~JA���F2��:LM�ȼC��g��f�j�I�F)UE�<��Do�^��֫�[1HΒx}hd�~dD�k(�ݤ*�W����Ԣ�T�ǀ|�6:���R\[Yd[�,����.b��K8>R�趶�'Z�j�>J�%R���s'�Ǹ��;��(G���V^��!�f����ۀ>�;������MG�s�{�����;'s��5ȕ���R��S+�}+i�є�T�̟�CG��6��i���On��5�_����Њ�������JU����gfok��J�f�Q�U)U��I�v����.�mr�훭�ѹm�Zo�,
�s����N�}�#���	���R�&-M��y}z^��.�������Rgھ���W�Y��e8f�l�,��Z���{��z�8Siau�>W)cb�c_�p��7�g��3e�XwE�t���;���$z,��Cq�P�{s��LZ,��KF�ױ4Wk�gα6�Ԋ(�j�M~�.���Vpڜ(��n�ӭ�m6�ٮ�zT�J���
��K%f��7�/�6}���\��	p�V�͎���T�u�{M���ʹ\�[�֝��a٨���M����W�ǿ�Z+�*G�i����o�{:�c.�N��p�����V��v:�9�~R�4
^��Npmh��~�I 6^�G�p�+��]��V�n�o�%�z��ط[Xܫ�:��C���&3?����W��܏#�q�o﮼?t��|�� �W�ӶM^k,=8��ޠ����n���q�ov�6G+U��=�����s�٭V�^�]���}2�R�Q��� F�u:�*���*��5����`:�a�|�dxx=�ߎ����D������~��}���"LHE�3����࢘�Ί{�LG3�N��@���ºl����M���D�h����]3�V;��L�E��L<w�p���f���[>a�G�΅�8��J:��)S�(ۨ=��f��؃��,�M?$lUab?_��K��5�^!���?���e��u��@k�O�E����IE�@l%>J�o�]�>5����r�K�j�=�_pcp��E�a���?��_h��3��>��ij�ڇ�I�� ��zd�C$LEơ4F�q����@�^�C�1g���MG���qI���2���� -<����B�7})\n"�x���`^!� >�>��M4b]ɂg$��)�o���OX�U�rѪqKCY�1Q��<V����x��e�E���T�I`e�s�YqM�&6�vH6J>Et��͝���(�H/_�Z�����6z�"s��EM<��lө`(îr#O=��pć����Tά'�y�<�
<�w�{:��K�C�:�$ǽ�c9�L�κJ����V��dTbC&�3;�$_�5�h�{g[.�ө��c���ŉM��;X��]BD�Rv�r��Z%M�I�NR� ��ۍ���(0a��#����u����(�(��C>7Xi~E�k�岹��y
�;��GLo?�\
n�H��#u0_1���7S�����}�yT��Q�HY��y.�5�f�o�O�$��<�ee���?z��^�E/�WƎ��H����ꇦX:�UD��e���!L?��>��a.��df` �?s�}�Ѱ`0�����A�9���K	��!(@ w�X�H�@�P���	!a�B��XF3�#:3�`�6o�\n?~��y�d��f0����Yf�Y*�kR�)l4ʤC]g3��O���1��%�MV��֚�֚jԄ�[���mx�[QZ�Mm��+�B�D��T�St�-Ů�5�k\�j�Tj�������{�{��{���}��矿�y������_���N�E�Z��[�C��2<�/�ڢ�T���A���{��و�sQ����������q��	u���Ys��"��
%�qda")�kW��':� f�ɉ��
HJ��C1�@h�
�-.I)�M�\0K����?	���4"��)! n�W94:@��`�Yf��NZ,,����%E�W��P�*���(}Zi�m@��"��a\�e�切t�%�@��J��dDc+��@w!Su�����=�6� �C! (�β� �,��a�t9-0EMC'zb��?��}�M!��bpA�w��дc��慮����� ը���\:�H�"���MU��N��Y}	��q-�Zt��j��hZ����e����5�1�o���H2b��!���,`$d�M��A�e�Rz������_�	@����c)���`�B������|�z��8�x�m	1�y�U���HS��	�"�`��c��D�^�ݜ��(�)��vQ�� ������<r�z~��pk�����������ႏ4��q$m	�%��ӊ�C.��g4APd�*~ܟ��CAOf./ m��R0p�]w=�mץ��ތ{ ��5��F��H� Y���v���ӊ�S�۷v��žT'8����И���_��}�yN}�t��� G�SPߴ/��>*����&A��<�_#����|]�fr�L�N�@�pj��L�|�Ŀ��7��y�0���	s�`-��Ն��Xrܯ(�V	�}����-�{���?��^[0�~{��0WeԺP0y����@�](2LX�R��9�_/m�7���:}�nd+ہm^*�R���xb��K��ΥSȮ�y+P�J�2��:��B�(񌘼9�[N���U=ҀSV����S���P
41�5	s�e<��\>����Vw�2���짓�:�8��G�<`��Ai4C\<�X�<�C�b��.�:� ��s�Zd���2�F��)�;āO+�hu.r�`�uA�\7Xp����fד*��ܘ�B���y�S"�=5U���ה���r�Fyp|[���7v�'�gD��Z�X���G4p�8�uH���oJ�l���W�)z~���ˢ��k�I��>�=wdv	�_D��1Y,��
Q �|lc3�E��� _g�5%��[�p��u($п��:-�2�t�W��T�դ�>@e���QN�d����`v�ƽ�v�%����}\)0+`:���bFx��ݰkH����hy�z�h���?^)�®F������H���𾎰h3;/<|U�I�d��PL������3��\7aD�]X�g�m�C��qN[�� v:��%�����i�-������Ƹ4�W�I@M��0jc��,\�O\�X�u��v`�uc�q�ևr8�g��g��e�gZƔ���ݠ5�qV:<�=w�5�gZ<�������i٠5�qN�y9�;V��g�û��\ˏ�:�j­�;��y)�q�\)��:�38�w���-�7`�����Z���J>�o_�����]���"�ɕjk���s@��h-`���(߿T�bA� �i@v���;~�|��0��N�`w�5���b� �8�L�c1�# �&�QP;G��f��M#�45�YZ�X֙�Wԯ���D�璍Z�a�,x�x�l�9�-ൃ��h+ET�K�f`��� 2R�P�p2��w�-^����3Dfɑ�{gx��p_;�UʫU
�1�z��!!��$���7暇��Z�{5��e��Qz�&�aۏ����qZKR�Ha|�r��U�#�5M��$0�w@&B˗���U������w �_�������( $�PK��e�K	��ݺO矿�0a�F�p�w>``+S������V~�XW,+���hJ�! G�
')���eb�,{|$��b� :I�b1F/����� P@!ߊ]��qZ���zT�WXu���P���������/�(����:�󇹠<��bͿ����I�7h�[o|�Sr��i��/�F v���o�O'b�9�����V�����������[��~�0_����N�z2��.@�ih��v\@��0����W��nð]�ۇ_凾�#��B2y��Oh�9<�Hlf�h��\-N0���"a�h7�Fv�^O��Hp당����D�-`erZC8jg�W�aЃH�D��Y�#I��z���Ps��8�1u���h1[������U��E��0˴z�s9p`���'�1�ᣣ�t$�a�WS�0Ʌ�	�V���ɲ���>A�L��M0~��DF��b���j�:'B��I��1z���z3Ry�}=�~H�3�h�S%�{��;�ߏ1&jf�ݵd�d+���'���z��{��������[~���sR��*.A��||M�ntom��G�l�޽h,L�g�5'�����̸����r}�](K${��LX��%����MBh9�\�g��28�rtG�.;�ƾX����DX�9�\�j��Y��r�����~����~��g;��g2y��1�����'zw�x+oJ�i��L�ber����n�q-�xk�f����z��Fj��e�j��M�!�+�wڭ^�F�e��Ƀ�9�d��6��+HEJ����X���no��O�h9�\���T��Ex��wf&w�]�pTa� `��F���3|��[��r�T!a�L6��V]	,�K䒌�Y�+���Ӣ$�.@b�U��9tfl-��6�,�`���&>c��U������dƱb�����'�; �rCΉ!c�����s�J t�e� F��U��@�W��pͻ$T��4`	�p?$�P�zV`�p���F���" ?�Y�c��u����M�`�v�+&`|*�I�j��L�[P�ܾ�L�ҕ���-��W�3
ߠ�u�)@�$mBb���(J�S��r��'������m��
2E}B|�"M�ႌ�E�,C�?e=�㿴D��mS���=�	��WX�"��M�E�U��|CB[�E˼d�=	_k�R;	��	c\���Ϸ�����1�X���Y�@��E��a=\}H;*H��|<����-���GHO�o]���]Ĩ����OA@�Io63{Q��$��7�����eK��1��f�t��0�����<�αfBG�	�tMC�[�I�ν���3��E�K<}N����,�e�=�{����Y{;F&����`������4���{�!�Z�o�����M� ���7��+z��CA����yQ�B��G���á5q'>o_�	�F�e	C�t��W �ND�XO�6P��H,ʑ�ֆް��iŧAQK�35��-OM������ȫ��V����=˅E jV��6#�'�\���W��8�R]hp���k�g�Re}�G����1*��T��[��`|�N�R�/��z^T���_��rS�$�y��wÁ���09S�S���@�ȧ��B-��z�dQ���l��_��'�xA�_�Bc,�m �=�[S�YSz��n݇��L��#����DIQc>�s�#�h��T��"�·~�� E���!z�i��1�1b�_�s2���2�a"DK?M�����Z���d7C�N%��/_�&�����6�I��� ?�Q�#����~�j��y��vV��Y^����u'z�&+|I��/���b�?@��/˒Z�A+�^�u�a4�>?r}���ng�I��S���;���4��C����<Ȥ����L!�z�qB+�>�����=����S��ԫ�T�>
}^���'�	�a9�'e���H�L��F��ŗ��$�Ö��/�I�6�'Ҵ�H��H�AIh_��S~X}�')s�l<�L�6B��D����-B	���'8��s���4��[9Q%@��s�����L�������&�-�职�i��!a��3�PlB������g%���S�tm������%����$�&&��{�i�1򱬅����ğ>��,��_Ȃ��Ll��#�4��t���C����]3�W���FR��{��<�?Z_j�J"���g�zm��cFTx݆��BY8�q��J�΀��߹jҟO�ةA���,�PS���y�K�,4���?��w29!�s�N�C�w�S��R��/��w��������6CtX�@T�d�qGU�F�Z�ˇ޽����|�-�߉c��%��X��c�j���$�������md�r�m�뵔[����z��_"b��{3Ш�~��XX�SFTO��|�_�'���aa��c�+�"g��?�X�t�:D0XgI�M�3�d�CF���pE�l��l�#�S4
M����sG����K���fw3�L�3E���qlOm9�!S�R�D��	�4�ڵ1a�C�K�+۽O��V48�GA���,&`��[Z�Om�����Ǉ�r�<ڬ�A�Pm���I�Vt4b�N+%KA��#��R �l\���m2%�c���-T�d�D���j��ۍ��'[�E���D�Xm��g^#n`Ab�EA���E�0���ǁ�!�����A?xP�X)
2U�����ڍn3�H��','vbk���~�y\X8`m �@�PJ��s��Ŏ�R�X���5/=�Q�wV�9�ERS9���:j�y���I܌�������@�����x0>��:�Gc��ej�gʫu���S�E"H�>x���w��;��k����"i��r��5��Y&�qL�`���2 ���ǽ	Gi�|1��G&�~>F~ᇸ����%�eOU�d�ݕ��yd�B�v�4�ͻ=�P�`Ӳ�ޏJA���"�e�$m�z2�G��H����˹�k�3�Ex��R����b�l������mJ3rw��U-US��oԍ���!M`d��% ����Ԁ��h�$j�*��-��9)"�of�Vv\�[O�(c����Da�u66���.�E|?���%�4����R= ��Zv����g:Z�-������z4�_�Rb՝�)T�"T�hm!N�T{B�o����Ǽg�����0"\����A'�8�����-hihl]��6��%��"U��j��ׯ|g��ea��FKXjiY@��$�4���~��f�bo���--~K���,G0���ߴw�m�7[�cO;e�X�ד�q�t � ���EH�8s��_�8�˔e⯵�j0X�z�0 p�$.6D�5/�&������q���k��wU."$9,�`��f�P���$�&��V��Ė���E�@���?��P<�k�����^��E��Y��>g�'�#��n';6�V��ʦٶSb	��{o:9"݊���I�KA#d���Ιh4�b�w;�����8�r9C�(]�X80.��� �l�+�w4�m��X+������2�Z��_����:(q�����+q�m��}�1k6��RK���5��=I����Ц�uz�Ϭ����a+���;�?zr$ ��F�ax�2~%Kd��2��6{��W�LM��7E4i�V���5�˕��r�n⮆W ��=�n�~ 6�G��K�,[Q��4�\�~mEƌl�P,����f�p�J"}���9��#q��8�
�>@��5RO:��H����^��K�e"���#+3V{�ƴ77F�z>,�]̂L�繀}dϨ$47���I�l���cj�\}���SnjR��u�J4K�Fd�ڜf5��N.@��YW�������>Q�����7F��TVB=�Ֆۤ���Xr(�r!�6�y4�r6�k��~�'�|_6Qo�[��Wl����� ����6���C�Q�a��~Z�ˎ4?7�jԘ��6�����i�k�8��Ib�V�]�p��| �a���5Dr����q�I�#10�KLyDt�f����N��W1>��kL���=ɔ�e=Kg�;�
�{�ЬXnS!�w���|x�tt�Q�bmQ�-~����9E8�����
� p��s��z�q�~���?����=��7ϳ�m�Ƭ�uܑX�9x�IX�9��� p�QG�Xگ�G���V�?dMU�˱X���z�D��BaD����)#ɦ�Q���:,�9-���pXRtR܀9�-�����\��l^���t�9�~�����7�@6Z�g��+�s�?���/����/��ף�.���/��� {�7�U�"�k��x�k�&Y��PD;�[����O�����WH�=�n�l,���6��V��� �/���͟��mF0a�1C�U���� ���M��>VSQ��)�b�!m~ɱ吥y����̠(<|=��j��t�M�5��ɿ�s��ٴ�I��4��<����=��,�Ԭz��d����9K��j���_ƾ����?&�V��8D��n��V7H��/��BآBح��[�#��7��ġ5�V?�a`'J�<^k;���_�������A��;�AP��?��J�3�[���,�]�D�I{<C�y�9v`�2P�&�nN5�E�����NJ� �Z^���U4�O��z�Y�dБ��<�SgOkY����R�u1��Y���a1}�s�~�n�������3�
��DS5ؘFig#�~��eq�dOe�]���q�y)��?i�����9��bZ	����6|�؆<u1' � �~V�N^��3��|F��c��Bߺ��L��[ Ziy���|�kB�\��j!a!�t�Y~����5�u��Ne�8��^���ܢl��QD?
�W����5Ґ-��l_�0wg2CC G>���|���|����`>�0}����>6>F����0m��`1���c�������cC�l|g^c�J�E��UeRm�l��*��T�"�ՒX�,��"ڬ�"�2-ڢ����j�,�ub2�f˸�eSMԱH�B�b�+��n�M��l�QMR�I�h��h��kR�)���q\��,���2��o�/���_8��>{���8��}�߯@�z:���!.�ʪ�µ�k- %>��&V��ak@�߮B� ۭ�<����9�f�1ߡ���\������TƖ�}E�F?o�I:7�tf@��,9褍Ӟ������| �,Fy	^:��Bt�(Np�z���U�δ�}��>��:���?�_��yy�Q�28�b�!�'��ո�6��8�Ap�1�!Q��5��.S{Š�-��*K�j`���	I��Y���K��(^._/������\��]��ӜUAkx[�^���dA�j	t��A�*���2
��̠b'"{�ӄ�@�dn���k�������'�J��ֱh�����Sh>��XR�I<�F/gxk��DGhf���R}O5�%�J_l9we���!���pl9��?�e�/C����4�0g�r�����}7�y��.B�f��7��/KE.@�@Y�>��P$Y��ݞ#pn�:XX}����6���T!���n��nWi�EG4>r�ӯ2w�Q�7AxmߍM��\r���7~��-��+�tl�8NfG���U�t��)�Ù1��c��'��z��#��<(�%u�����|ͨƒmݦx��c�"1�*���Ŏ�u�^!,t}���I�.��_<'�N��O�Y�<Z�?����G����^y��.I�ȯo���~k�%��6���<㛙�yn�����CIh���㇋��mݯX��&����z��K��Q=�j������tB�����[��;�g��@��v�L��,��?��ȸO::��|��+���;����:?�j�50�Y������s�M�5�5~>�U���=A������b�B���C���|׿�9{�7�Y�}��T�������({�x;)}>-�do��'��m�ND��hG�uͭ���Ϣ��>DG��K��|�6��(y����j��˾9rϟ������Û�&����$�ҊM�u"9��K[0Ŷ��=�\O#���xt+�.G:2�fz��}47�GM�j���<ܴ�Tp�34_s�Q�(�e�v�!�%��M����H})'Y�]���v�Ă>�O�Ɣ��FߡҦ�J\g�N|�o�h��Z�.; �G�g3H�y����S���[O��9~H���3�nx ��~�[��R�U5���3���T�%�kY7��6���#�,Yt�[�����<��=���>�"U�U��D|�do)u�g��W�D�kHEba��)~����;���#� TB^/V�w� ������9����+]��uj��|�����Yr�����5�Hr�^q�Tn	�ܷD^4�=���$�4��?�{}[�7W�5��kU��4���U������rW�mk`]�������C�T"�����*]2���ņG6�Lhuk0y�?�.5�h�&��'�t��Fk�+6|�OL�<B�v$e��3����lņ��z�k��#�ݠ/���!��ӯ�O`ɋ`� ����Lۯ����u١�X9�66닂u�����l}�-J��L}G=�g���vxjjJ;Q��-?9���^mzY�+��$?��2��羃T�7C]��榽����(��r&�X��@�-����kҡ�%�/��Mh>��a�?SS����������l�>"��WP��i���WU���W����T_ӹ�v_K�ݮ����/�>�,�	ڗ��~y��<W�\�#fE-�mYI-k-|��L��d{��l��Gk-�z���w��Im�k^�j5�E�/�Z�Ko���G:�R���<���q�8�:W��"�ɲC��#���΂_��K�������c�S�1�O���ʙ���j�3�В�@���rjlnq�2�D���4� ��D�F�]�>p��y�Mp�W;z��"D�B_$}
� ��:Gh>���MU�}l�J�mn{"��y�?�|,ɖ�Ϩ���	���܎�8�	s��'��Er���7ߌ�<��u�`�� �8`~���v����40�s�~�ο/}>�9�Y���0=�u�rh�]�x'���+xA/Y.Y�=|�gu�{�3�ݓ=����;,��^��Xʇ�`,�:s�3����fvjfO�2�����@>||�qW4��#S�ph��E�v�ޝ����}���B�_B�@��҅�i�/���,�Kt�؎�WB����>pW,� �,ݚ���T}X��u���$�n�׌��>h@u���y%BN#D��<xFž�@�pIϢ����9�y���y~����Z�K<7�'�U���o�a]� �
"i�	��-�I�]���@��<:NM�D� 5�>:��y�(�#�l�jl@�(u&���Q�ީ�'�AC&��:�+Xa���E��-;���h���(�V��k]���݈�ns4������b�
�E���+#$>��!]F��QUH�ޣq�;��ؿ�Y��hX�n6�{B8F�@�Q(���۶eW�t�,�fj{8X[�{��x�H�2j��`;���;���6k�h�Iu�0%'�j7T4%�h:VA�S�(��1b����>��h��4A;Bh��0�^��YE��䴲�+^�+9	�өg��q�E�)�l4m���f[�W
A'~E��(�Q��j��Z��kg���QA5��^���A��1c��23�
���F�R�Za��:J��۩�Re�nZ�|��1�p���J{Զ��25|�t9sgo%� ��w:2}��a�wmE�����8q�Q�/yگ���'!F�uB۪W�w���Io��W���>_G�����&�Z�5� �+�-�i�V���
N�����kf�F�q�����.����_xU0�q��[�b6�)�ǖ'��A�C�?Oi/�Z���!�c���Rr��~s���.�!<;)^e�`ʵ�S�@`�e�������crt�]�
�N�����xE���B`�������#j4�,�"|{k�"�o? �z��Ѭ�6���7�Y����)i����m��D����2�3��YP8>����&?��8����}|�mu�x����ae8�9��_ �K�:�B|����1<4O�&�`^�[8$Tk�%�E�R��caH+�g�mQ�ݹ��F��I޷9H��vy������M��b)z.c	���X��\)�� ��:����M|ɞrf�Q~ɎDj�!��X����j,�;!AU!!�2Y�^dI��"� ��.�!.nZ
g�@-�+���ᅘ�eq�*#���Ĥ��n]8uZ����)M\���-W0�� ��v�?6�K�%��1��f eрb�}r䙭n�ť����rʲ�p������3's\}V��g�Ym)�9���6�9����4LO�&!��Wc�I�X)(�:/v2Th�r^r4fiv�-Gx������6��֍SaXL�MD��/nQʯ�H3�T �\q�M��:&�.!B~g5+�~]�f����;C@�b�,�m���k����XK|��V��ǩm�"�Y��U[m;bN�W��NeZX�0_��I�����!�oh^
�|�pm��1���r���&��{��PgMx��WPʍ.o�O*���ɤ�ݞ-'X�b��y��ȇ"��דV��׍h�Q���̙&�;��HʱV^����"V|�⃼a�F�lC����᳒l<�	 ���|���g�[Kꨪ²$j�/�6�>�|��<7�����ƸV���H�鲫�A%N�4T�o�Ȃ,d���r��bfGw},k˵	�<���+}�6�?M���ۏ�=�ķ4�c��"�����bY��G�b�H!K�Y�e������rE�.�uj��|��b�a�%�� ��a���f�5�U"��bQo\S�ŹS}ZN;8�H��&D�u��I%�WS���d`���p�����.;�Ȫk�ۻ����K)��"��m�o�Ic9�����

Q��,bM���"��!D�)���j���7��գ&��I�AI����I�v�C��Ëc�&����=%�8 ni�'=��Z8�|DYZ#(l(ua��(x���^��P�j���m�
U�ū"�`c!T�\�!�Gk���S��e۠��J$�V6&cPUpNT<���@B48����΄�m�s��
�n#6�j��ϭF�$"c���z��1РG�8�A	{=<W ��(h�T��"�Q��V�(Tg^� ⊜�� 4_
��X��DF=�;��n"�>VCx6v�&�
˄��K7pt�n�٢�I��沇Ҵ����d;��-��~�-���j�!U.k��Ԝըп���sS˂Z�Kɠ��<x�����R��S�1�s�1��ɴ�1�穯R�"������C^��F-����:�S�w���Ǽ`���ނ��PK�>+�jDM0���Ԓl~_��QU@Q�`��������R��;�k9���=�tǛ��t1�n��Z�T���C�m	���5$'�b�|�m%r���D�b�
`�/d�ڬN��f��1W���ET�IM�z/^�jʝM���"����Iv�U����S���(�k+FfDH�+<�.��Ggb�ą9L�4}:.Vz �X�#TR�'�}}U���ӫ��?Z(H�/�t�Ҁ�3O�*�L�@g�;@<f��Ը�>�m�H`P�{G���Ǽg���o^�}�q�?Iӳ�/Om����:`�-> �������|g/V�C>�-�4��]YՖ��%~���`��|�G�|�G�|�/���[���&�G��nrlnf�sw��u�GGJ������D��T����T�w����/m3ӳq�Ϧ�qd��������8_qv���������#���!7术�o�~;�O/r0����+�%�h�����q���-i�.�&��S����>L����6��zt	��/ie��#���>�#���>�#���>�#���>'S�Ϗ���t4d���/���XQ�Z-�	H�_I��RqM�K��	�f ���o�()_=������z��J�¤L��K@�m�Mu{ 06f��0n�飫ZbƮ�EKf@����/{����2���5��T[\T��v]���dm�Y��V�25�O�粒�(�^X�,��TW샌�E�USW��c+�I�w�!Q�`^���c��v��[��)=�L����t.�g����.���O��e\d �m�����s��~bS413���?�qxW�녂�1�E��[�eb�}��M�l�.R��Ce,��@��Ed8�e��/H��2潨�*����N63�K�>F=g�HI��td����J��N������,s�ҋ�d�����{���|�;�����?*(��Ds�>�_j�}��9��r Qm >1�I��' �#&�������8��
��SG��|��N�����p�h� @��O�ɀ��y�OI@���800߷˯[x �Ȁ�X�3�g�u�8�A�`�6`n �\	�7�P�JP�;O�4_G�[�)\�!�K�D ��`�b+\��&L#XF�����4� BD�؄܄�oP�	Z0Q��IB�2
t�*PU ��q�q�Z�B��х|
XfL,�Z�!�0�5�1�c�����abC/g��6�3�h���CM����>�9�s��A�é��g���<hy�����������Đē������D�D��P�Q�Rb[�*�>ĈL�L�MO'�e�u���q�{�9�:�N��(\)yGQƊ4�gE5b���J�Q�RaSAT\ ��HU�U�V,V@VxV�XtX�X�YYPY�Y�Y�Z$[n-������E҅�B�w1w�x�y�~ŕ�b�1�X�9�@l7�1��ѓ�������`�T3��*��a��Y��8ָkv5X6>6b6�6�6 m�nn@n�pXp�r�9��8�j6��aҡ����q�A؁�Qڟ�t�3�#�홋cճcl�*@Th�k��G��χ���c������2�2QY�؂��x�؅0���ЇTC6D����h����P���Km�[Um�{k��B�W�*�ײ5R6�7�92:�q=�ܳn�ۡ��6����~
��_�[������pj�A\7D�II	I4��BJ�[�-��t�:K�%��H�7��*��q���}�U�`���VM�'!'����Ɠ�܉.HW&���mr������y+���f�/t:�bn�MmҔ����P�P�Q�)):)W)r)�)�*+*M*ʕCO���������.�WSۮ2룺�	�,�h7�KM�U�]v��K���ے�"��z�~��T�d��`�`�a�1"1F1��љa�fQ�Vc{�����.f<f�g�3�3�4-4S4t4�55A5kkLl\l�m�6�77���M����'��%8���̩���0u���]�q}M߆vpw�;�;�<0<Y<z<���o������yv��މ�X�֊�6{r=Q=ў�^Kޚ�=|,�b����;����}��՟�cϣ�ߏڏ���	h���Y���o~e�F!	!"�fХP�P����t��(��H�Q�T�\�,�1j2�4M�-������0��#������J�8�VO��:`��i�GFzN%�&�*��ڕ.�uK`K֦&'�i�*�O�[�fӌ����?���c��Qa0�l%O��ۜ�����S�
��68k~k�Îa�p��@�!7���(����jT�Գ�T�g�nJt*��GJ[ʫr��&�n�ϫ^U�ը�U�U�+��lR)�V����b�����*��[�\\Y\���qlx���r�J��0���R�"�i��/�/��H?���.�F��ц��1�P�lc\c�2�e�'��8�+(vU6]k5ɛ"ͼ��1���ԙ��.�o���D_"�����&�FM7'�Jѐh��_��m#m+�2�S̫�X>Yc-�˚��{�F��]٭ů��S�l���,s8��ٴ�C��.f�3g����cv9�u���
�N���Q���6.&�.�B�LSnh�p�Ҍ�k;��+��/����L�_?W�T�Hhoz�RWV�Z�ƊY����*Ѹ��:M��c�~��K��[��zj��ǉ�����9ΟN�H������=�p�~��`���D�� )���j��`�����P�!Y!ia����p���H�lI�L$Q�SƦ�t��b���"�ux�]Lb�gX����������t�n
7m��נ������^����N�1#��6��g�7�BmM���c��.��o���"w7��\�솲D�G_$�%���I�e�%�S�f�%������tú���L	L5L�̸��7z9�ɧ����V��y��I���S��ޯ�x������x�{O>i?��A��p0��
�w���E������^�6��Ի�e�k|�
��x�6����jwuKuU�mU��Ǟ�>�6�z���)�s�,���E���[���j�����A�Ą�ń�P������ܛ��z�����=ci� �������?(j�<� ����ts
z/܇O��(^���?�v�7k
��`	}��`���z�L۰�����)B�J����%�G���7?+o�j-�J��t��VO������2E.�o���~p���e?k�˟�l�� Y�;����a!.�8�`�}h~�A,V'��M,�H5�����B���LjPl}�"nI)ѩ�kE���vԦ�^�ң�yZ�5,�I��]K$gxM�����=���#�M�G6���9B<�����-�:{f�&V%�c�Sq��Y�����8�M�m�Il��qL�!�	z�r^Z;���
�0ʭ�%�R�m=&� �,C��7L�t߁��F�Βf�,@ni�	�!�XЮ���������b0�A�s�D�˪�&Zig�V��Lo��`I��Aj`�(��Қ�N��cоً2Y��/�m��$GN;Mb�N����&\3���<����?�\L��&g���g��+ڵ]�c�%����+�9�����F�o���<Hw�&�jb�!��G)�*��ê1ː�.3i̾�m���,�r����8�~�*��d�L�{�~�)�F�hw�5�X���c<�k���&��КmH2Mw2�F�Z��yY8�2�N��r6S�Mn��z��1#W�V��5�3�$�͈"ڵv?��e�D�{�:h�$�12��'&B�?�)��/�)q̨Fh����e{���w�4��W���*�D%�,-�{t�o�BS�����ݠSY��Qu�y�S=~��E^��0���-Stn�՗����N�|H������.t��awcJ��(qn�۞5�-��7���R�n2�RyrX�2���N�3����L˺K|�g���+�*d�(�y��%����#�\t�X�{jD��2%�խ�뎞������!�X.��
OӇ&�͜D)�7�ic�s�ﰮL�P�(hr^Ή2�F����udk	!S�� i	��6���8��^mS|��ϒ��G?�}�ޯ�/�]���6�s?��|?����w����1��$+�op�ӭQ.�!A�F�����rQɫ�O~(�+�]���h��z��TS�uY�k���p�|��H\�_/���%k��c�SD�5���_v�����y�	Q�ks���[�f�� �F����2�c�*=y!��n�ý_ޕ�f�v��wRA�x6�8������%��b�����ev��Kv*�dD5��©�6*�
��������%�h���Z�zְD�ƕ�Mvؐ@��"P�2m�ق1�a�*��n��گ��*һ�V�^���t�:efL�A��#�#qq�؀���GX��Um�`��5n�Z����c!@��E`��g��0�����;��^����X��M�j��㖉:��&1/R����r��n���p=*�/q#r�,R�zY��D��i�6k^��		�V^�ϲ/���Iusy��G�-�%F���Q!�$}�\din���Պע�<ޚ�T��kp$)���,�b��~��1�9�M�(o�����*B��&�9=co	u_W'����-�g�a�K����u�U�G���Rטk|&t�����vE�Δ��{���W�cz8���T���0�Å�g]>��%�(���m��#A1y�M]����Sx$FY��K�#��w��)�e�\��_č�ww�Nc��M��ހj��3�Px�z�{TJR}#��JM�i^/x���c��oT����L%$�S��������7]��������d�RM0�Q+njh/%m�]K�;����z����y=�mpK�sܛ�a�HB�Qr�M'�,��J�+ICͺ������?��Fݙ.�K���&���{c8���~�����r�4�}�"�yR�[*=���M�e=��Tdvoӆi��;���+ű�j����b�}�Q�N�g�,R?�C�R��l�#q��R�7����2��M�]xQ�"�{��8#.��s���!�E{����D�	������N�?���:��Y8�Q_��q�-��)=�#��ܛ/it߀G�<���ܻ��$�_�I�	���4�ʆ�4o�,�~���q��H��T����M��FB�{(�eؤגh{i2w(YA[�m����w�JpI<p��,Z�����]:�����w�����|e�{Z���cR�&Mۗ���{p��||>�G�
��j��mPf�ex:��K�|�Ź�u=��k⼏������|��Lw��)��1��E��a�;�r���/x��s��O�D,%�-D���y~C/�c��J�dY�R�x�v��$?Mw{l]Ӽ��ϊ�������7�^Ƕ���a�2��F%MRE��t\d>j�6��]uYus��_4ίw��f�*ـ�������� �pj�#�X��K�pظWD�%�B6w��-�2݉m�c���d��{�Grћ=�`7I�OK�A-�3L�����p)���}��">�A������S1~����(������U�� M�N�F��H�I#�P��t��%���c.KXY���$�X`�B)�d\���!b�� �����~o�^���`�4n�`8a�귢k�	��u�u
��5�_�y�wXE�����Lp�_N�ku���w���U]���:�G^�ס�D�r�X����u����d�b^�E��N,o���݂P/y�Ùwv��	�"���	�'[g ��F���`�Yx��
�)��G�GgV�o�]�T6~:cOԩl��JY�g��n�A#�4%CC�#!�z,N����ǡ���/�1�����7�93Վ�N%����{_�(��.-Ŕ���F�~��d���6�K"
�d<	��H=�u-q��'�����F69m�t	5(�V�,�[��D�*]������Z[,�R�V����{
��[8�ζ�Y��`��ݳm ��k�r67��%:k�>�*?�(����2� ���F��f��A���T�O�8��<,�Ds��0ח}��/݂^M�Y@���W�M6��X��9��w۔bSy�$K�	0|ј�m�i�Y� �.ϯ	��U��\Ýy�������>��1�PTc�o�3��4D�7W�Q#܌l����խ��K����4#�:cI�4o��U)���W�5�����Q�о7w�~�D���z#�y��Y�\����1��6�����s���aʏ��i ���*�	�iB�[xT���%��F9J���g����>'!rl�}��������>/�^�Ƀ����y��.��[/�*�c>�ܗ��r����z������d��0�:�l��I3� �Xd�$O_��[IM����=Ĳ�
!��\exk]Ϋ��,�e�j�j����ѩ�ɩ����O��#��e��#��Q�R��	T\��좠� ��F���¤0���cyٓ��+A|��g�$S�M5�ڴ]V|���Ik�j���^ш��X�6�>cR��L��5�GH⤋���G�~�K3\�4��PRE�{�v�r�L���N�ι5&�I�vW�Y��R��W�u���x\x���]�6V��1;�����ӵ�|#�e �Y��9�7�5`
����R��I�Vv��66��B��E�GF <�Ջ���'�����F%K�u\wY���镒:���x�ǯ(]H-ﰠ�8|��=	���x�<6:KE���5��P�>3�O�F �ͮfJO��G)���[�(�	�w�#Y0a����9~��w��QĆ���� �-N{F.L|x�Mqb�����ǐ�45�QąG��E�F ��ؐ�/+\�;�y0q7 �#������v<"�ծ$�]���{��>L���N�z�2D�V��75!��{�6y�{�� +�Q�xZ7M��u���K��#/�qy-��/P�5gݣ4b�CZ����8F�Ae1���4�E�ƽ1��j�I��t��	��м��-�|<I�&�c��p#��)I ϸu��N��dO�l���?.9a��8x�u,p�U����a���~� �A�_������^V�6
}��'z|�n��d����]Qn�b⠕�փX�����G�(`t���١Jڎ����39���B4{m!�	���Na��cA�̏p���aI��{+,fB���$�h��H���#��D$�Dܧ%�qv?�|�ޜ����L�z*��|w�]l<�Es��凗Uem&�o�A���*d�]K�;�9�*�N{kU!�8Tfz��	�,jv�|����!��(*v��n.�-�m�O����1A�g�^�$ւ�dp�I�*����3Q�0w�F�\SXY��|<`F�C��
�c����﷧��f<V+�W��Q9s6�����"����#���'�[�%?2���ß���7�r�T���������s��mwO�_8n�I�m+���ԭ�0,�kU��-����,�٥��
���.gn4���?m�����!<��JԶ�_>Xn�s��R�HF췖���h7N���|��]<�D��t橰�iإ:������#���M���NoE�R�=[�#����R��b-�H�z��M5U>A3%�z�ys���ܽXB��
��G�c w&�����0SB�([��)��X��M�=�4p�uvV�ܱJ�:��;���K��ni��΋z�7�+_��!�X!ʛs�tv9JNϬkR��RS^d?�N�u�b��f�[��7�`n���F�^�LHl�'Șb7��2��������A�(1i��/�ǋ��t����d�`��k�
z��yEОۭvn�"�'ۡ(�R�~G9$ ���C>��p{7!���<��Vj�
�xE��E�J�B���x����As���Mb��d(�P"@ܛ�v@YW����q��rCȷ����R�˭��>���g,��D�(x�*�Q�tI1ѽ!�)i�^�A��X���T���Z��	�ڣ@E�	�'�h��l�r�o�� '��-�a�R9�8�+sq�42K����j�!���`�mܣ����$�RV�$Q���ړ�H%6�ۀ��:�e��=ejĭ�5��R82w=q<r&:CǊ�XyN� �o#�#aX}aF�Rɟ�����)u�M�q��&�� ..��]g���w���uf&h�.R�{���I�v�h�w�J��&�ͭ�t��S�^P�4�}"F���=�Յ��\��	��g�Q���*��간}B���=$�>�������)����\���k�rp���k��)-;F�W��WMs��Z/� b�Z�b��K#2
'vcH��9�1�i�j�����,�|�ka���������X-��9�	�uA���>�#)Zk<ʖv*w�g�fҢ�U`�Y��jR,�`:`�[̓����^t.��A�\�A�#ٞ2U&�2��u�rƊ�p��K���C=x�����5��U��X��F�ۊ���Ft\�o��ݬ�(�p	�V �^��z:������>�T��z�~�AT�y�\�=�\�ӓ�|��E��b�hh��"��ݸ�I;�y���b88�����I~rd�� �'�^�%�#�iJ
�aM��^�����op��u|V?a��F��P
.�޳6�[� ��~�'>:%�B:j�i�M�"V�ʩ˔�Mf�ʒLj����`0y�p�zg{��\�q����Sd�pI�x9����H���zq^B_����_�����0� L��j��#�|)M���o��V���T��X$��	+��<�F%�����njG-�x彵Ѽmv��Bw�P;�������PYm�鶎++B�Ҹ �P�,���� �)Z���Mf$M�]����%��=W=�ӊ��Ob��.����%59.N�z�-X�]R���v��<1�o��ģ>�/�mrk}� ����ؗn��$�8�������؀���~�XfM+$s��x|G���28I��=�6m_�I`4�,��+U���� ^�����خ�ё���D�[A&Jxw
�I��;jƗxL��Hh&4W�s[��^-A'�ۊ��<X_���r��4I��=A"�Ĩyĉf�F�ڀ��>ްgPH��u0��Ie������E��΋��OZ�����o�4%7u���k�:��l�փ��x�������w�0��*B�;�m�������J���ߺR��,�|�07�T+���D
��N�����Ġ�ZF�1Irr�]�c��9�m��9u/ t��W9n�¤j�:#Ƀuy��wj��D����h�N/��������ی��?1tx����q�@C-t�D>�P��ځGZ�����n6n�5��t�nV,kH��	*`���J��ۗ��oH�M5�,��y�C�ijt̓eK�-�Hsk�A��gPR�v0��Ba�jV�� sf@��N��;4�:�!a�2FƎD�%��~��y>�4*1�p�T;+�|j���8�ǜ(�w9�Uv%��Nx:�K��N��G��6�,�ܧ�.�L��j��]�ׄ|Э �8|���@OTId���/p	u��m�E��zN��7�QZb�V5:�tU�g�LRY)Ii=W?�	~�������ZP_��L��]�oCH��T�a/[���ظ������3�ľˀ��mŠ����i �/�oސ,����A�s����o���٤�;Nu����`�i�sc�cw"h�A��:�bs�|���?�7
�p�!�qͬԃ��tUľH�"�ne`p�S"����&�flC|g�4#��ˍ#ǱA!����΢�=�V�dI��R�f�GD�c"�L�m	��*Aٟ��*Kڪ��UG����(����?������wp�˧)���c=<,1�0+�S��������v��	D�F��%
v�p����el��� ��Qgg%�DBA_0�.�J�Ñ�5x�u_�}��Y�Ym�p�mQ3���{�t�.A�#�6C�;l�՛���������H���E¢i����Ύ��Dh�V����;�%V��&"��`��hE�}Fpg÷�}�^�x��?��yo�(-_�^�!�ّA���0���X�m�YCN.c�3xI��T\r
��ma-Uj��l�c��B�^=�MP��EWbi*{6��iWf�5,o�D9��*GR��G���_���υ�J��t��^�x4ƲbGL?�c^�ǃ������� 䖊KsB]M�7��"eM�aX;A#�R=� ��,�&�z텢W�36���G��>�Gл���� ��X��_ r�$�
����N��⡡ͶgA��j���^����oΏi��ߡ��R��r���繢���n>���$���lj����\da��������z	LL���p�=�.��3�|�W���x��2Ħ��S�^�����[�8��r4��V0�Uy�Ma�=�غ�1,Դ�\K�R��n�$�ӄ��M7'����u/�wa��H�s�CS��*LnH�(�>�y멙���B�����oiƓ@�틺�ф��1�F8 b� U��6҅���4��@�4��@�����B��Kn���d���jb���׾+U� �pDL]t!�\��`bU4�HS ܓ��;3�ۓ�+��V�p��CQ7�d|\��RS	�XbS�F�N�_�.#&h~u"����x�MFo�~e��d�56�,�EwS�Ԇ�Co؞T�e�Ni�Z���?a�LOkvd"Ȏ�Yb|���A`�,Z�K[n%Io8��H;�"-)P ,P�Y��1�
�d���,�[��.���]9�Bţ����1��2���:��P&;�0�+�w��=]����r�˱7'��v��&��-�x�O��="d��b^u���|$+�1��aTF6���
T��p�*����I��������Ę��޼�{�����.�!(�%�b��_w�>+�0�_�*�w�G߭:��>rw���w� ڡ��e���I���8W�L��m�`������f��P�/n���8b�ƫxA���8x�.|��/Ec{��9����� 1�U귄b�4ze�l�m�k#u���X�jy�`�y�^�ef��7��x$2�����)��N�Z�G׊��t���$b<c,���r�ܠ6l��p���y��	O�*����#mk�äp/}ů��j�VD�慃:�̏ѽ���_�TF�! m����K%W$<�q	�d�������O[q�{�b�=�nr<񜆲z^b�R�������&��R���,	'��\eJ�s]���/�����RP��� r�z��#:�S�7S����R�AZ G�i&jt>�\���oE�Qm�W$�o<��϶4��qt��g�~���2w-�/�=cy `���oI!�$%����hC1��t�Ro�A%l��I�q��^��#�c�-�]>R�	� ���u�_7�K�����
�:���
����SS��m�����/il���u<��J��L��l��K<|����m�� ��{غ��m�����4��4Ί#/���A}���AQM���Hc_�� �R��6�N�i��V,-d��7�uL�N/��k��[\����K��]6��m#b�U���uU���R�I(Y�9�6V�#�K�ٲ�Y�/t�����@Tѻ�IمZBi-�nua1�O˶C�&��[
�!��*c��AS�QOɳVĘgJt���@gÊQ[5圗�p`�oщB� ���8�X�5�ș��⠙���Ԉ��j�s�1ĜX��$;�{���|iA���l]�s�0$�������-�_�"v��1kW�H�q���^G��$�`�By�o�l�.���o��D��OT=%F!��Y��M>���Ǡ��:�����bO(h��~�p^� �96 �KNH��y�9�O�tm�D�cY���� {�P8�j��A���O�܇-!�"eh���a�+m7(�s4gk?h���s�w�K���995q�gҚ�����f	=~;O���_i�kA� 8��`_)� J��bJ 2J�j�#�v�+.8��*�Pfq1\G�y]1��#'��Ily�w^�~:Y�.y3�@V
���D��[����Q`�j�� ؁��H��1h��7��GY���aA��%�� 6y{_&/�mD1�'�'ڥ�U�Վ���ZS~am������mG�iħ̝``�t�����F�G����Ǐ+D{�����^����JF�k��f��U�d���a��~_��ƒ�����|K�����C��Q�>x�l����=����X��O�k<�i�7��2��_�$g�j�x-�r�?��V]����A-9����� � ��|����'�񸟕ě��VaЗ�C{�������ݝ�
���X��7���t+X��J�Y<�'��̀j���m�'�<��X���?k��j�Q^T�Y��;f�f�ee���o��ա�Wm�_���.
�lz�r���m�d�~�mu������&���;��b��c��y���~ǟ�}��g��B���f���ݿ����e~3�q�#Ip@\��S�u05�O��������;�M[��0�ٸ&��'��xt�ڿf��jH�&	YR=�bB���>�O��:M_<0����Z���	�S�f�G�/�`�؋@[���c�xs���PmU�b�"7���0�y���ׯ��xK�E�2�����ж1�g��eу��5�ǻQ��_�p��5*I����ucZӡ���hw7�Э��:K���jp�c�"6��\?�qTဲ�������'�D�L|8��t9EfM��Ϡ	�ł�Q��1)��Te�����=�}�#p�{��j|��4�%pcK@�B�K����B2Sn%�@]>���7��D�h����=k5w��e/`VF�d�������g��)kB��%S-������W1r�}�!$ZNua)xU8��n������p��x������y"N�E��;������U�;Mv�r�/��M3�<�֔R݆���o�q�ϑ��ΰG��a�_��o��o�ƒ��6��b��p�+Ϳ�;u��ے��s�Ŗ��t�4,&
�Gr1���R��(���`CI ��d��n��ĽN�d����A�jᷚN�O��SV�
z��)���$�w�5��@y5���אb"2O�B�(gf���J ��d��1�m��TȆ"�L�F�J��1G���\ˡ��&�h
3����#� D�[��\��O����O��;�e�v��9�w����FW�+<�&�^��4�iE1�\身p
d�&�veI�Arm(��V��+F����T��}���#�N4�V��F�`ڶB +�{�{c�O�kᲧ���]�|�h�M��"�=ՙ"^�mL�;���c�-h4Y�%�2��Ny�a����v�Kw�{�=�����5�r�!:��J�9�;k1 �(fc��}~[�'{��XnSQɖӒ��Gb)β�¯c��%���K��{*��Cn��Z�#*'�e2�A�<	HQrr�#W�n�Fsi��x�!�8<1�ë�N$��ۋ?=~K~�睛�6��,a/*�΂%�$7LK��	��nf��i�Me܀�f��+₇)�w�EGk�xH�j\G��פ�%&{�m�dk[A��YE؎��� �z�֟5�ҥʏ��c!O�A�0��׋l��ع[���L��C��9�����@��m��.٩]��ږ��_�0���%R�m�M�WB;`�u@:�4#G�0>�z�:�yGU��z�[t��Fk4�ŦzK,QOj@�s�l4y�m���B�KF漢L�����XY��i��[�m��G���d�G ��e��SQ��\��jt���J=�� m��ㅭ���sW�����U���P)t0y7L����;B�!Rȹq����r�	��c��L
��U���k��,�����C㛨�apRWzv���_�
s��\���j��̀� i0a��dv����B5{O;�@��^8�V��|{�AGH��%�#���
��(�~M�� ��oE��{����ǃty#%��|�ת���s�l�ݸin��K@1�ax���-����J�w�'�� ��T?�+�ʳ���������R���Jx-s:0=18�K�b�@��b�@��Wk��p�}!�����r���R�fy��	R4�O�2bj�=�A��wz�k 7<�iQ8-���Ë�H+�5WL��9��/�%��a�	귲|q��1��HA��0�fG�2W�+���H1Be T���\2,���.�oT�S��iJ�C�C�8[�q���r�������l��]�g#U�
:"����-����4M�Mk	��6�q �w��ecZ90�`)ib"���u�k�7��	�g��y��>���O��ECðT��.�c�y��l!�6h���vgc$40g�pc8��8�ccl`0l�6�>�>|F��l�����6�6�-���l1�9>c���c��~1���&03U����&�0�5L�-�1�Y	�R�7f"�pܬ7ڌ��!eS�VE.n�F����U5-B7�T���ն�%V�[�}��j�Z�d�`��tR�n)b[�YĥJ�&�S��o���߉�]x��뾻���y�}��Ͻu���[4z��
���-ݱ��	g_^�f�B`�h��l�����z�&{�D�w1IƆ#�KpG��́�.�?UK�H��az��uw�P�)�_���^ϛ����^+6wvl���*�A�SuM�����p;JP�c;�h�'�������83�ˬ�$1M�{�S�r�C���9T���Q���N=�=`�7`F��C&�7-;8�����������v:軰�U�WZc�8�?��r�d���ӖV�w�4�j�����g]r0�k���i�+'���ީ�X��I6�����b�/R���~�w�P�gx�Dws	�{#.�q�c�f�u���Iz֭��5�ϱ=�0����B��A�w��:��VS�����1��M"��
�����A�"��`��m��G:��%��&9�9gT#f�����\�w1gw6�t/���h���U`P0��.pU�KV|��3ҳ��v0��r7�*+#0��6��-�流,��S�-��~�_�'˘	�*�S�9�Q�!"#��fz�,��,1�W/��c�C-��r��LJ�5攒�@�#-Q��pT���@<�-2k����y$�;m��^
5M�(�d�K��vN�=z�~Ǔ������amR����i�4}R/;Pב��c6-+=#Dp�\�Vdɥw���A�ӏg%Ls��k�ξ�2�+r:p��������};'UWhr��@��Q���H�6�쎥��-�����=�uNlp��x�����5�I�d�-�_��Kl�l���iء&<�/RNY�^��dV49~I!	{Q,ڐ�ME�y�d���� ��Հ����<Qlӄ��O�?���ݖ쓇�d�#��N�D�@�����$I��Q3	K^I�a�5�fikBr�a �F��c�T����!���|��N���84i� 5��!sbS�g_�l:�_��1D�Oh����ؠk�:�ʛl�|1	�Z����f"�����#q��`ߴ�}�g�ڝ`�����ф���St��?�0��u�el�y7�$A �b(���T�3�~�9���6���Ur
��S��$���0�%��b)�o0|~O=!^�;B��`ZE��١�����9@��,q�G��0b+q��<	݅���|�01y�$Qu{_��W�M#�X�#	]hE�[F���m������U�lb����7�lYHwJ�>�{��p��pq�Z�Yˍ1�m�J���A�f`br��|"�%����)Q
�Si���^������c��������%�
����Cp��b�^����Y^��ԜOTEǯ_.�6W�t���?�»�A�}M�,�d�9��u�c��6�g�,�c�խF�5Bdʯck�A��؃Z�-�K�o�&���S:�����x"{-
KRXX��b]̈́�:��8c�+�-�ݬ����:�y6�Hn�b�-�è�y
Z��é�������oA։R뎅ݐ�&���9��P"�x�q�`�r%tf;^r���*���,qC2�F_�6�a��  Wcha����]�g�uu�%���� ������툧#� �r�� Ձg8�Ň�ZaCP�=Qr���&f�����6�}�W�?s�E���6�����#��*|�����B��1�ܙ[���VրO3|��u�!V�+�\��b�y�~��h���L b;/$ׁ�I��h�����M�e���p�8R8�+qJ�nŃg ��2,���V��5k�����B)���?�@�:}rw,��M�,,���,�X�	Z`�����ȎҞV��n{!}8�"���PӴ̦I�8֧�Aer+S�w[WB;f�1%�V�2�_�r�д�Q�M:)f��`:(�-�49g��+�2ivk��UtM|�tr.��.%+@��B�A��;ZZ8�"�e ��?s��B�{��zT�sY���7U�w����`$m�oA7?�ʮڀ_�1o�������ӧ��>a�i}�a��z��f��|�T��ޯceRY���p ]�A��>3~�A�ɽ�Q�K��q�?�����}r�g�K���l]�nu����%�үҭ���ݱ}Y����-����'m�!�ѽ�gѯ�{�g��}<O�Hܯ�_�}���lCNv)�(������{0�j�݆lg���ü��-ʶ�HػOMck�Է��5�V��sk��\��/��|����¿79��`��'�����o$������*��Wo���'��D�6�>|jA�)d	�"�;���$~Y����y��q^Y����=sz������ʷ{�E1�S��/5ZOy�m����{� ���Uq ��Ʒl8���hPy�z�|��س�v9�uR�*Ѹ�T�*��d<���#�n{�w�j@���-��i��r�wnxƦ�]�u��M��!�@�os���n����K8)�@ZS���(ｨ�#��Pg���,���`���%�($�"~MN�=���P>��|Q��B�qO��(=˹�|B�}ۜ��`�[�G嗁o�|�5 n��s�a�`��O��I*�Z\Z���~x���owW�\�����ܶ��x�m�
���%7�4��������;w�v�?�8uVD��O%������PSq�}�MG뻒ȑ��(����T�ƭ@o�n�"���R�I%>����u�:�Ew>)R�h��,���k�F�:1A�H�	� S����ED�������P,��$1 �(�>��C<R܅_�q_�wd]h*�s�En�ϲ��3��*	��g&)<IL�bU"e �$��Ӫe9���A/G!ʇ�g�oc�`�0I+���"niϷ��;���i&�A�ޯ�S]�ۥ-rGsN}�q�;�0&��i�|5�8���e,���&�����S�l��R�
c�$i�4ٟ�i,��@wPsp|�x�S��V��d�!!;�I�Jg-)����0��Y�-7�!�6�n�bqU��\��vST�=<��J���?O���/Οu�7��A���_�A�`�@n���No�LmQQ�	�i�.� [���=<g�$tr@������C@L H--��㓀?� 	���&��NC-�=���2��QM��S�8��2�sUPO��`.�O���֣#��?Ӿl)&��=KH~�z��H|�ls�D��@('w�3�Y�9~L��`jF�OJIG'���tpyj��G ۾I�A,�x�V���0R��&T���� gא��1� е'��kS�� #�:�Ly{��Ų�\���d�A�"Iypk�X$9��|����c���[��$B�6$�!E;�����4<�H�NX)9=A{N_�$֖���Eu���3�P&_��xK_@���D�t����2q�����th�C(�\�;�o�4z7d%����^ɸ����I�V��Z��o��z?h�1�.�ò�8%[o�xa����GΗ<�E@o9�o��֑��	I �]-Z�f�A�#Q߃5`i=�{!�#�����ĳZD~��� ���L̀YLL����C��s-��~a<2��##��7�Ky��k6G������{e��dr9%l�Z�mhEX�Q���-(��¿�<9����;�J+KLM�ⓩO�xC�*Z
&��/89:��ܰ8#�E�����j8Vm}(/���|�����u����G�T�����ܻq˝��(;v��^��� �Ŷ�o�ۮ�ZC�-B"Bv�`����$+�0b��,�`��?6=a���)�3��?W=�ض�N��'��ʐk�w����W�������w��Ť�Y�`&�Р&����Ȋ
�Ƈѷ#����nuk�^w/���MG+G�z��e��d����ƴ�N��̐����}=�'�H�A��j:��zJ�9ݍ����˭-��|C�'�W�Kg�a�M3ǲ����|W���x������|zu��n祵S@R٥���-��hݿ��:�~��v��t�M�i�Fb:�O?w�z���F���+�~;m1�Y��#3�ڨX^��'��I�+i�� �������f��8�n��Qx����.�y`�@1MK1���:}�nבu���Lʦ�;�"��H�H��W�#�CGy#��h���E� ��NX��L� �5%@_A
S�����`�,��O*�U� ���&�q��叝�(�p#�_��ymܰ��|�����c����B�������D�g�9����1<����|��w�<�漿�j) `G�>�0�w���&m�xj@��wjj���sx{���:<��l���NN~w??s		;�����!�zV�xqa��ΑMǥ�㝼�Ο)zH*@���S��BV̪7�H����q
�GNya�3С������zbG�{: y`�LK�~~�L��?��`���	��r�|���y�n��������R���1���oP>��]��	�v��e��۾ך��OM���@ۏ ��'��i_�������e��k��k)�CNÁ�ݟQ8��̉�� ����	�O�[�����nxR�&o�����L�J-���1�]�fOf�����T�GD��M
�ŴmZ���2M�f_?��/�{NU<����sg��S2t@�g��e��3�*|���s����g�#zs�w�y3�}�_�ϩr�jI3��9�$֏�{�"t��y����^p>Qٳ�%��3B��N�R���oW(��,�?��֮w��:g(�Q��Z�)ب�dU��Lݍ�8 Pm�5��3g}�{�9b�9�hf�'���+��T0ϫ	�q�u,�/�}|ռ{�ޔ�����C{��9��tыiO���{��1��y߉������s��k���%�vEd��������U�}�N�g�r�,����u��*��$����h|3��J�����<�oz9T{XQ{ZU������އj/�J�����.>~�W|��;D��z�c�;�v�._O>��$t��u��U�qO��?�k/��4e/�uao��/b��4	P��t2>��^+�Hّ%y��˂�^�A[o���{X�f8O�z���;�Q��+AF�C�6��υS�'�x�ȟ'8E����U<
3`zxU;�xg�|�8���]ׂ��P�=�1Z{��_*��^A��:\��k����;��
�g7���O�<*��<3żsȣ�ҾVr�`h�+�S<*��	�燑Bn[ B�T[����ǒ|�{���o���cȡ#�	S�t,ۛ2�@��Rq��QÚ����O��E���`(j@���	�<��Ǒ|��f
��[A�UHjw���1z$�+��t�p��.Py�	E�Ȗ���<�����rÄ�:y����Iľq@��u�?��xȞ�|��<�WL(@^1ߧ���f�n�x�q��kL��;�c��6����	}�,�X������mФ�Q;/g9��}[��_�'?､����{��0�������( >EG��ʖ�{K���p?���c��$���3��i���{��{"�ՠ��k���~�~z\TTO�<�]���WT�¾Oى����tiW�[���*�%����4lm����%�
�⊁<&�ԝ���O�l %{��vh�'�#s9%ſ!PZ�$6�,iǁjq��hL�4XԠ�ys�ۉ:8��߬C�	�%������������Ѩ���"�Px��E�V������x�m�E2��-H`t�ү�wn���H��p�d����ޡK�rP>���	�H�����L�P��S'�x��~��G��x�yy�FhZ9��dȂ�n`ڕ�(f�]�{ȓQPͳ�(&b�}���p��@��سȹ��S(&��H�>����H����ЊV�ީ�8�O������0��	�8۔ࡕ{��yEC�}��D�>IB��N�&UR�;�J&��T��Q߾�[nǍ�{�⃶g�%�98C쨕�Z�p��.�I�K�������$������Q�$Q��U�۳+G>��{K�����/=�ɖն]��T�?=��Σ��hl;M�]�i���A���"�����b�5K�$���C��D@�ϭ��CZ���7��d��py������g�UA˝��
����
���gO�S��Ϗ�˘��l��, >�q�|��O��?_K)�`���o�пZ�V�k����f���%��i�Y������E�7��#C"�B����R��		�q��\H^�K���K����o�/�	�`�ᕚ��k"�>�2����߀`�}@e���[7nJՊ�.�gt5�����$C&Z��N�J�*O=��
o�
��-����rhqa�@*��qˍ��X��c�����m�0��jN��a�4-��h����8��a������0�B�|Y�b,�<֯OU5�YCB��mt�%��*���d���My~`/&N�w����59[,c�:���{ t̾��������`�����'�����LQ�v�l�:�~(O_"�t]��`�T	���0�⭆H�)J:�{y�c3�N%���s�"��3ـ|��~	:�w���C<��e��������P�"��]�Bm���~HL��XKx�,�I���ø�d.Zƹ|�ųC�f�/��Wk����X�Z�R�����_��[��&��QF�.�����{/��խ�'؀� �H7hٖ�݊��5L�ܵW�irf`ғ���sq�b�4��4��P�y���F�<���y�6gPͰ���Aj����6]��M(m�jSn'����yxi�3�����-��,��!���^�� ���dd�z�FF�����;M_�b�U4/5�}�]�㜶��M��b`YB_FU���ɴ��B�}Kl�a��L����I���`z���SҫsdRN��'U�\2����]�
|�&.A$�H�ncgǗ<U��)}&K�	���p+��u���H{�!%e��M�,_�V�S1aj�?��C^UJњKD�����5x�%}&�@yX4�k���׶C=wY:k�0`& E�>b�.��$)Cl,ad�m�b���Ye;Gk�%�W�Ij�fVx��v��n̲�m���0��FE�&6[\ 1��Uy��(1)cg5�!�N��"�փ2����1<`b�(Mx 7�u��78�b[cn6\,)E�t���-OMPV�ݙ*�L[}�e��`�J!�����i���2�8KͶn썘C��|-&��F"bP<��C%�'4%UG=��y35��5D*V�&��������T����,xr���7_~�]L�� ����-�R�+�I���Z�T�2��P��R��y@��YLar�K6j��)o�5 _l�XY�]^��qBw碳�K>�3+��w:l*���FdH6YBQ�=�\_m:�Z��;�PU�Af�(4�w+}�_u�AUa��bȲ���0�0�$�]�n@|�e\I���I�%w�2I����u�ݐf�4�~�kn��:!ި$��3L��.��[m~d.�54�Ԍ�nQd�,�"g^G'Ć�1��&ٹ\�G�ı�e��ѣ����*������6�  x���%�׸��N���V@\H,-�K~3E�pRf>:��6��
�m�"�.�i�kIޡ�M�Ak���9-8�|)�-�u��	��hh�v͂:�����^�WN]���O"� ���\�0�gŧ��������W�3i4Ř���H�ԫy0
&6�)k@�0�u@�`^�:�aΔ[0Y�X3KFH0���aT���A�s�60��
N�{�*�8o�$+������]d���%m5q���"=˹ef+9,�y��%gqugo�q�w�g�U�T���c��d���&r�Su�sVbO��&�^��E92&�ԝL�Rݑ�y��x"���d49��n޹�-|&�
�/��q�Pz���c���ȕ�3���������k��(��x��3)�<
�=����q��!SKp���V߇[!��#�@�5���+��2�w˨�(�Y��/n>s o6YР�ٲ/���|VCV|]D�ě�hp��d�!�
J7�U��DD������FK&&�+��?�bm�M��N�]8��F�p9�{R���;�=�`s���A�=�M2	vlA�)��~���!`N�k�e���뎆�y�#yԪݗ@�D,��w_�X	4t6?G�}�m�em�"��|���L���7"iLk@��z�`8��[�� ��u�j!b<�pLE2��Ibp�io8|��D�Пl�K>^�q�<I�N�J�\BY�ĬE����DW/oG��Y��z��k����G2�s�&���u�~<K4�t�hC� ��
ĚKOcnڈ�Ht1�H٠��Э$���0�\�}gA����β��nC�z��� ��m���G��(@���=)��/VE�	-���"���S4� �Q�3G�*M�a��7ƶ$�C��׸۝a&�޶b/�Py��s�������/�u�@1�N�б��t�9=�r+>��^;�V���D��!�۞�u"X|
���Z�C �z�<��"���(Z��� 2�c��ĭ�IM�~Z�r̠
��'�CS���U[\��+U�x�`�u� gg�[D������WͯYW2LբgT.w��Y�D�@��q��.�5���y9��b��o�F�}H���m�aoU����FF�7��,"ڤ3��e��+���i ;
k��D��<0���v:-3"N�gm�F�4��W����ԏRU���ЉH0��Af��	(�\܁�Cq�5\��%0�O�nq����q3k�h���TL$? �C��V�����--��'4�����<>ZfbD�KQ�6<Y00�i,���dB���md��Cl�v���+}�t�5�mO_r��04!Q�ߔ�-��L�Hyr�$�v|m�k*�W_V��`>@�'��������ݖ<�j.�6.Rێ�"��n��5����$*�>lV]M�Q^�I�b��� ag�$��\���8A�:�@E� iY
n]���9�y��4NV���$r�s�f�"��T��C����z*&��WD�O�P��K��܍ȯ���
�4���u��V�S0�KY��p��_!z���6��"�;`5 �}Te8�d�T�X��6":
�aH��H��2��&��m�T��P����_�ְ���y���%\�:Z���K	F,�ͣ`���ȫJV�՗1o�ɮ�ĎH��;"65YwyR|#\�<�6�p�f/��n�O9khz׫�"����hЍ�U��}T\�٬!\f�H�Q��F��؈�lδ��\���([vX�~ó.�ǒL��hm�<ܘA��*e��}Hzϵ�Yǯ���MQ��v��"�H�ˉ:6�e,�'u��=��M�Zrn���jUq��è������(�FY�828n�i��!"̓~�����RUH]��3�
w�4J�7SW���:Ԯ�n6�	C>t����"��p{P��+3�>�:+:��X��b R�Ighm�ܴK�~��Z��l�7]qy�'!��
�X�Mȟ�:#"�"��.��v����l�Ξ7;h��RN&7u�YY�[\���V�^�cW}Iv��=�=��%����ʂ����IE�Bbs�͝r�]��Y�1Q�m��lc�WB��t�/��eٕȑ@�$A� �5s��S�C�B\�Ȣ� �����hm>͚�K�j6
�X
m��X	��][>�f�H	`DA�"X2��]���L/vr��U��,�yg&AҌ'iе���L��;�(�t��N��*�Y��.���r���Y�p3*fI���ٕfJXJ���ʐ��A��/e�y�2�5NUw{TR��?�*���w�t��V��X��������_���{�=��9�_�s������k���\%[_�^���s=��M�?gj�����������T�G�V<mG�f�ע cx�JH�3W�G�j�kOV����Z?��w�w:�4�3�?�{�y�1��O�:����x�G�R�dt}G��+5�u�<F��h�U>��rv�4E�����M�@�1�Ix�����7�o���:V=�Rj^¡�6�Z�Ur,�3ݼ.U��L�ޝM��)�O�pn��8�+S��>��R���o�cƽn�sm���M~�K׶�K]�#L�:n�뼓�FQ�v#���˦�G�Sv����֥�7�m[��ꞏf{����{�7B�s�ׂε���u�_W�����h3�3��x9�e��m���N�K8׽�/B�;�S%��\oG�:o��{
UCC��3V:����P�j��K��^?�y���ݵ=Z�;ǫ���oV���T�='�x}���R�{����O�9˚��+�nYֱ�z�wf�e���(�(�h���x:�WL����m�.۬w�B�3A����4�?��4�ǹj�^�J=�o�fŬd�_�lz5n�E�x�c㼵D�g���%'s�s��v�2}��e$��yD��&=w��j�]363��VD�
�K/1��nFC�l�/M�y�ߍ����p�V��lÌy������]��g�6���Πb���}������ĕ:n��dz���j$�B=�ЅJ��i�f]�gy<=��yZ�Z���T���d<I�7��^�e��y�K�cC��2؞=W��r�تh����@5I�4/WAN��׀Ӽj���MQ�����:�<�O����|Gv���r�s+�~�cyb��k�ʏ��]؟����!�X�f�P�9,���K���̷9E��*ߐ�u͛���=c9�<엦���=�4k��]�L�7�=�;�p{����V���E@�a3�m^n��~s��;�S�i�<���ts\	��� "t:^g�c��/ːiuMb��S�m34�6Ns�����VÓ���*%�e{v�����(���ul��}D�/;��wG���������WT�������������yT�Qf(]�>�P�r=�O��o�������/�n9N�i��֒�u�(��w���c�i[&C޵���k^����Ɓ���ڳ�����g ��>�F���z^o�c��o�ڷ��s|��k�����:SxȆ��8�ZQm���uӹ�����;_���X�s������^<�����^�z�c/�x*֟���w6��)z�� ���CX���f^C�ٳz�=2����l��&o�m��[��_)��y�3*{��~��}���U���t<'��S}h޿�V��G��u�v������?;�ۿ�����
�{}?���Y��5]�h���Z���?�h�F�Q�3�^O�V�l��_���c�h��v�}�B��mu�n��s�7��v��oײ���8-s�ZU7P�������ULh�Nɽ�����^��p�/�I��f���#������t�^��Ss/_�}�{��w^��*z>I�k[o����Z���3%r�ئa����m:�o��m�gO�ɸ��>=�j�j�������:�W�oT��73��Ӑ&�������9�(���sHO�=����#����=�����?eJgݺqk�JB�����v�;F��G99�<�/=���c��ϓ�VI�ĵ�?t�޲{>t����W(��6|�*��9� �=�;��ı��7�#����cx���+���k<�,9�����?��;�GڟO�(ݘ ��&�ǜ�����ę�נp>}G�j/:�Jf*z��W���|��+q_�RE8��^�=��1������u��7��Q�uOƤx�����
�x"������W��9������<ڢ��;w'�O<��=���[�ג�h/�u��"���p;F�0��RFt��{��#�@���=ƹO�BZq��=��r�r�dJ>����J�T���a�ge��#9�����c��*6�|�/ݽ��f3\��~|5E/�A����:���V=�b�����Cc_������ɻ�-�b���?O�:&s.A���7;�r��b����s�N�־�3��;�7h;�l�Gq9�\�ʎ�Zv��E��6��{�@��NsL��]m�:R��y���ۊ���&
��1���d��j���|���I�k��.����Z�?��bc����_)�w懛
�ϔO8	�c��f3��6���2�k�Y&\d�_@��>](mw�|�)��G��o�?+k����`=�3�ol���$h�h����]�?v�]���o覴X�'���U�uSk��]N�e�|/>�/*k�6w�E�����+���
. ?�E�4���T��v����>���/�QuH=q��Q�M���<��,��y{5��3���]Z7����/���G����~�ߓs[��ϔx��]�z����?�ǛK�G�W�nz|��N>��4L��"�����=(�+{-Ĺu?�sc��<t�v���3(�%��;�u��#GL��.���6�=E�Hc�Y�H-�m��4)�>d��bz)�y]	@�D0�M3�Pbx������B��G�q�Ϟ���kշ+Qe��wqL�G��p�:nN��	�<K��d���A������>f���<�@�����)�Q�����F8ȇi7�m��;p�X��"y�^�^5+ܳ(QO�/�yAn��å|m��ۭ��z�Uf���ͽ�e�{�z ���ʃ��#�/�&�h񕳸���G��>����h֧^��ڑ���R+SA�T�c��ֲ��b<�x���0��s�uC�h��#�����o�v�q�-���x6�R�*@��|�=Z;�q1�L���3��ߢ=��n~+�s`E]� ��P Q|P,�>}G�Q��y�}G�Q��y�}G�Q��y�}G�Q��}�\R��~ʹ�\8.������x�9���s����p��J�HYM+��η� ��VI�}h?������9�'�O���{�' �j���FI��':��$��ڃy>�� 9���?x�"�CWxF�z�d�CV)�0�+B��m�?.{�i(s��u���Ƙ@9Xu��[�@u�H˚.��d��_I��m�w^8|=|׉LwƆ��xh�c��^j�;�&�G��FK1ГdY�$�YraBV��N�+��: ������{@��O ��� ���М�4�Vu�J3X���0����N�+����	�;ϫ���}V�O��9`�!��:~r KVK��XJ?D(��W�s��':�	���@Nu��p�F��CX!��d�⨍'�xPh	�Ny�&}\}8	�0I����i�r5Qr���`?P�Ȝ�#0�+B��
'q��i�4	�k��Q��
�v��¿@�Z`�F���H��z>����3��WgM�
��eyᡱ�}8	��'��@Nu�	=���V�S���![��69[���N�+��<�#ڪc�݊��A��'Z`� �!Z��h�z�:|
ȫ��!_{���ʯ�r�@����<@<��Lݮ�[�錆pNM2}��0'�ƀ���>�˄��jrrҀ�h2l:�N6�	n*`���Td��#�����Ün0�T�����?�
��h���	��%�*�����>)�{Ӵ��L��4' �Y�ƧB8	Ý���8	�Np����MI����o����2v����x����⋝w�{K�%�8$�s�nZŭ�62��8�B�0����;w��p��p��nnMX�i��D$��%K���?'���_sTl�y�N�:���4d O%�5�.D��J@Np��$��-�7�Pf3$���M���N��t���Y�LPM��ťYoZh4@
׺���خj�Ƹ>U*��������P��Cm�C��{�j����Sq<"nkM�^��:��>'Ҩ�YƧo,���s �;f�'7�?�����4�E���i���i��R�P�
e@��O͌��ϳ����� ���?�'n�8N �	�g��:v��8<����p'���q~�mh�I�	���\3Lc$�#4;����l�q]�z�n>�?�b�~ܠ��\s�w��P������6����%��)�)�̸pxV�?X�;�Ұ��Y���s��W��n��q��� n��@VS{Z�՜�^���9e������@�^�5N�
?P~O����[���t�7�\	�KS �T��� U�$�N:��h@N����./�������'v\�~�k^`�����ց-CPU�@w�����͘=��V�n�.+�v	�>������giw�w� �|����}������:}\};
�?���\����~�l�W�z�s�zwH���	6"� ��VL\?���Ujc2^}��zӳ�`�v�U�>��O�Q��w����+��C�Q�	}��o-��B}�O�\�� ���p��W	?-N��PT:3@q�����" ���}�0�Њ��zR>l���5W�?X�RaP��|,�^�++'�Y|e?.",�3
R�A�!D�SA�����1"$ :x� �cF�[��b���|���AE��a�O��ƨ*^�/�x5�I��v{�Vd*<�LEy�Lb�d�\�������0`��g��=ZE������r�-1��4��m2��� �ׇ;�%�H�T�'�T���4�B���i��C�d"��H� A����H�&Rm�����~v_��qM��&bf}��ʝ:����L�G2��zw�B�au��9P�J^�@z �vX�B@.W��t�	#�N�β�|�L�q���CU�CZ�)?#V����#�e�F̘ �D�QTB@�#��|`�kf2^�س1��l(��� �@tt b	���O���Q�A�6)fl���hF������Ё��a�	Y�ҁ������2dy1��ŤF�~0�g������O���%#�^D������"� �"CׇM-1�@g�V��xG<rS��H�E\@��hM�JHSoӫ��p11���x��'�>b�O���Pnk�̎�Q�3(�Ga},A5�w;$H��@
>L�s��,��@~.���i@>��];aW0
\����^������S��ry�b��Q�A<�O�#���t�FS!�BI�}l���F3w����B-D#+�v����J�Έ�C���	���{JJ�0@Ɓ���w�|�OB��pG%�H /b�-���6��e��s��� ���!L��J�S�,��
�n�t���9�L��!�B���z)d���!@gp/L�J~/VЉ��1��ߟK�*0�VqjE��&$}�~}K	�'�:����"Dw,b#�'�y���?��P>#��WN��mGK�8�t�veP�*IgbnH��\��'���S"
V`%b��5tfV.I�'��F��$0}��Z8�	&{@q�,�2:C�L�s�+���a1�k����@.�x?RSdQB�ц�E���W ��Z��d�Z&~Y��zE���@��K���d��U>fw"�%���B���,=&��3���=r*|��K�D���n�qC����\U���H���.��p鵡�#�̂(?�½�C�ŀ�}.U������(��f�m�7m�ew A���O/6�����P~�<qr4G(�/�����"� D����.V�P�!Bd�H�E�%��xD��2������ �� ��a �_^��\��28�GD6�db)|�y8�b�8 ɏ�m6��e�@�����&(r<��'f2�I�>4L���8!<����P!ɞ݁���J�ۄ�@m�T�Ј#7	��&�Ƣ���pn�0{�4q]������v��\ش�C7VƉh��	EJ���.mX�)a;�;hL��R����\�W�VL� xK�3"�]�B<�d=�/�z/HS��\��(��hˠt����a&��X�E���`�?B�]���LǓ�ǽٰ�H0#B#L`x�곟>{H?Z{�𫂌ɼ�,�(J��� �@Y�C����{Ӷ�Y���7�A��u�Q��	���	�Ҹq/D�4�$a�� �������ؼ�%��BL}_:q��BY1�bȔ�:��q��@�C�����`�w
yTQ�m8�@��_�
�����0P����	�!@�]�����G��o!�%`�[�a= �� ����z��pk�G�wvP����t�� s#ܤd�����*<p�
�jM�)<��绰1�xe�����2���B�>Ilu�Q�]��)�k�����RJY���37�3=�p'P�0_��P/ޖ)]	��n�˟�S�+����pG|L��)h$'	]�7k��H�f>~�� U�4�&�$4�t������P'h9��= �]A���#D`E�8q"��J�-�|!����&���fPK��X�Ӣ�Q�n$.�#��R �6�����{��n�خG�G����5HP�����"v4��.�d|�fp� ^ ��"�<{���]0�*���ߙM�ci"���pz_���[����7Մ&W��P�`�tu8�L�:- 99����Jn�
hl��
|QUS��:d�8(Y�%e��	���$���Ɇ��)��&�?��!D���G#B�<˟`F���@`P���}����I,�ױ �~
�2������Ps
�'0Z4�qe	X����;�IW
������ߙ!H]�u���Ƣ�ƽ�&; 8��l"�3�tN<f40�v �[)	��	��D@FrD>� ,��8���-<�
O030t�(,�2&N�5Ǝ;�<c���!�P�9������әNm9�bX9N�� �j�2��a��%\F��F����BN��i �V,�?%�<����;���(s�@i:T�TrA9$�,�%�ć���.��@0H�0�_;<�iq�O���`%�L!t����p(9xh�V�oC�`y���u�)�ܭtN@j��		��m��`)H�(�AM
��v��	� K��%�D��$��	C�.3
�z �|#���;	�L��A���:#`\ �!;��#-t@��M'�(%��_���G yE��`�V�+X��w��?�N�����P8pGΙ�"��$&L(r��!���@p
�K���:l5�0��@'��)H^n�i�~S�A��}E����/(��p�!E�28t�%
��r�Z��k9�а�Q�Z( �P�A2�T(Bj������@
�{[/:�D�[iF�.�
JV ~ '0�*Z��p�ZH�*����Lt̤�@�N�=2B����I�>��A�/�T��y6��D�C�":��	�J�CJ���`��B��-2�fn"|u���E����0nt��t`��n��Yȯ��S��hR7%qC
 ��	�] s�+��T:08�� 	�����[�w�
� q3AOJf�uW��4�ޑ�r�Rr�D�E��m�N�M��V�;�PPհ�\ Bs���.x�R(�/̏*ww%���|楝J`�≠��2���PP[���@7`.�[Pt-u���ƨ��>(u��p&ZAv]��?�dQ�:�����t�g��א�\<��CP	���uZb�π�rc��d�;2��q���
Z�`�������$F� ��
R������b�r%es�U��.
ӂ���K@܎
3����b��?)�#9�u$�~��96VZ>�(�2wÝ���8p9���ojLsx�~��31%"CLZ^��Iܱ�ɤS�ꀰs��r\,\���	"�DiP�l	�I�����2�!����`�$l	�VH>\������P}~�����C(��	�2�H��	��U&CunX0�����2M�yA�_���#��Yp!�8���8k �)>B�A�Ӗ�3�Ot�p��!Eb���$���� �ܐd�!����t�՗��%����Hpďt�"��K�Y�Y��xz�|lA2��`�|�BF���&H����7'��:��{W@�`���}&CJ���CK�C�u�V�$��j��+%2 `p�p'���8�y���A���M���.��nP�`)<�(d��@���y�7\�@��X6 �uŨ�K˨��is�� �e'8��W��EǦh�	�s�81u��������X&L�4�	��"VQ�H�SE9 ܽ�싱�j6d� c �8���^ I�oE>��R1�uḁC0��"S$EIUx� f!�
Z� �G|a4	)RQ�Bc�7Pq"��r��&(@/�`����(Ox��o�7:��4��8�Q+酇�oڸP��9�hQ�%� H�
J��ؚ�:Ӌ�P1��2��t((X�C`؀����$7��OH��ΐt�W�xё�ۦ�Hy���G���q�m���L DP.�� ��I�����9\u���E�$��^C�}!A��2{�Rt���T߉�A�����N�{���p"{��(H���t@��N�h#����h�`znZ#�����S`*���>:D���.�n8V:P ۀ��	�O��Y�!ʖn
G����&���<�����O#0`�t���� k'�x��8�2����%kN���w�WK��06X��~^���>x�i ��q���z ��ɗ�+�:`0&�� �/Xl�X6 ��.T������¿��������!%�TP�d]��߸�4�7����>�e����,0������w_a4?�\9���>��U��u�,B�5�^��g3��B����d� a�����uzh����M'�:<��2n��Da������xʒ例��S���L�_�%Ց��p=RH����i�nD(�('=X�f$��!�
�A�9�,��Q.[c QCc�>P�g�N�!�.�Ŏz���E��!�(��	�� �lC���Mg̓S��P�y�zs���@t ������k�t"����30N�k"��v��,���r��u�r�:�C��F4:Ή��`�9���\3��@
^�hy� (&U
�*,(H.9�1|�1��L�	i0�JE�8���!,��� ���h��D�G.�lSSJ�G �%,���ΨOS��
U �|n	��yB\�{�U�c������+��-�^�0E���=�_:��8�&8(�xLH|�Qr�#<�h��A�Ù׍�8�� ��@��f�ִF�0I��.I )O���AB��.�2q� ��?�jd�䐃��z$�uF�Oǋ�""�R(Ѝsa w�1��A�BBd���
�?����\�&2�&nE2��A�iGP��RR�_.������L¹o�-3��(�qA�jk]'F9��[+�K��X�	J��A�(JX��N��`���q�p� �#��J~�lC7X#)����e��6>w�Cȁ҂u��)�
gz��/t`��� .
��HuY��P�*��R�.��1��]`�@"9u��d��Q��Y]l* ���0�+���t@�&lJT��I.H��}�ILƥ]�z�K�[
8��LB_��Bc@���T��z�H���	�f�ȁ���z{�T%�"�q~�#zTV4���k���`ܐ�#o��
�.KG�R_�J%
�J��2��A��<����z���:o>��>��f�4�*�a�ō�)�m"Y>�1�p_0:���@�b��B�SOiHS ��7��=r�Ԙ� h,��I͡������#���`@eҸx�������!愧�Xk��E~ =�c
(dށD��$�o��f&��iH�RaJ��n�#M�]E���f#�'��#�p��
z�7Ջ�B�Y2G�z@P����	�Z�J~fe�$r�j��E��0��AG��R�,)6+~��P��hH��?� 5��f���y)̙̒���Fw��]3Ta��;�����)9�i���~��n�1H�ʙ`�����`-��b�RWV���}0�'u��[�X���5�k��6`���=���f~��i+%x��A�hp2�8,�"�,��e%��A�fHa������0@���PSBC�H 	�%���ر�TΥM�J&��3_`g/2 ^�M��2r2Ժ4�Ⲗ�q�*l2�rA�&���AM	���u�$Xh	ܱ�l㩼Ѯ��_Z=1��}H�
�/J\�����@ H�	���FMO>��H����a]ˊ6���&�+&�F[�F/�:� �')�y��C�a]���~=^��Ѭ)w6n���d�!E�v����i`�c��D��u�6rO�Ԓqd�#TK��ap�OYa�駔�����tp���f
(�b̔��#�������s�5:y_3��k�;�!�N����G�zX��w:W�.t�/H��h���ԤP�|�&��$
�6sum�	0�sr��3
SQ)f����(��aA#���al�La.U�#�'��;�G?�Zli��R�r�����\�du��P����8L�P�/����=�JH�����G����te��|��%z�Β. n�o��z��&fHT&�CI���9������P��W8p�/����"�	3����3z�C���7a��r���K��%&���c��,�hy���a�\�xk�j��a��xJWp��f�`hZ�t:^r�(3MfI��m45�-J��Ϭ5���@���Q��i��V����7�05�ٲ���E�o4'+�m� �7`v�I�[�t(�i�9\�w��s�&[&����%��	����N �|��0�� ��[��C 8�hNW'3��1:NQ��o�W�N����;���5p@L����z4*[��>��xS��;��5p@N�!��Վ�Dʌ',���cBr�!9_�a1���n��s�Ƅ�p@j��$F���	A�4>q�М�\�_�S|��8�hNW0�0@/~0�����݅��{𫸴�ٹY`L�@����):��X�_1�=K✈ ���ϐ8��h��`l�'z�W��~�*�u9���U§�Wп��|���a����+� 8.H�P_@⾂��S� �1@���V�9��/�fb��f!�'.Q ��=�[u6��^��o�ZAt�W���k�ib���9���jE���l��X�Ӵ�pp� ~{�</�XN; ��4�����]�� %+����ix]�˵q�\� V��L(0\/�8������$�ෆQ��༽�:x,	�&0��מt�R0Θ�f�my�c���'���/�i��BbY�<�n5�fٺ�SV�l�wiwtr�Z��*�&��]�f�0�ɛ�d��U�
��7Y&Wf
�<��l|e �B�%(��q��m���9�'k���^W��xV���/���{��{�~������|~�������#����$	 >[�w )�,p
|�?b��_B��}�Fy���o	a�����8n�7p��G�#���w	a�����xna<+�lz	m&���iC������)��Ku}���a[I�]��7~�宇-�Sjz[ WR��,�ۢ��}����^uv�'S�t�î������՛E#�l���֛�;y�`o����o�����M�^���S`.�������S�o���[h��)]�������W?�w[���ƧO��������t�m��h!�ɯ�+!;�m�u������C*�țe���kt�=_qm~�ڤ�������^�Z���ڞ�������ΣQ��no�/ߨ�|���)u5��wp������� ��{�+���Z�t�S��7��{�]����d�~��'ۯ9���}���={�c_M~��R竹�=����}.��1Κ��1��GO]rV��/Y!�i�Â�������[�w�}]e}'�����a��VV����_�NO���g�����O
��u{���K���n�GV]I��xM������;sd�׆%����/�� m�ޝ7XH��ә��:�6����t���GZ���X����_X��9v�.��=L69'�pu�+�v�$�R�{����GE��t牰�����M��m��\ZI��������螑�����M�>���ًۢ��'���L�.��#-k�ޣ�y���w������v���ԍv?��9�|P��5O^>EQEQ���E�{]��=���=w��\�%��(�,0/'�k�Ċ(��0�:���[�y�sJD/����Q�Ab ��|!����t/�EH��_�S�]C���	��O�w�q��k�o��F�����/thu�/���+x��n��f����������t
���WC{��Ϸ�8��C�K�Q���A�2+ 	(��_B��|Hr�Cm�k��I���E�':�?*�^%�!�owe��F8�����xB���ǣ��� �"<��8^&N
;@Z�����sc��	��O� -<���'���_B�S����,��vI_o�7hL3��7��8�g:悲�p�7�o��;�5�;��a[���xF�3wת ����(���G�8�������{��%�>�� ��%6 ~a#�z�0)��08\�³�`p�jhrJ�  
�`���(;���0��@Ц�tDp�e� j���:2 o, �:����L�p���Na}�@^��1�L,0�Q���þO�þ{�Q6;ߗFk9��l��A�8�#�<Qa������qϧ� ����RK怜�( ~G*�lMi��kmF�p�c��@oS�a�����c�L����R�
N~�EO'(#���<�v�����A��&T��QU�g�J��ł�8��u�wVi}���vp�wB��
��Tn�r���g?`ۉ�!% �ǳ���nMD��o�}t��6��3=kw�tC�A^�p<�`�Y���q�-���=�b�&K�`�j�H����`8���1�@��Z���t��꯼yh�S��z0f
��xA����[
z���$Og�>	p,+��β� Q��&�3r%�`��g���(W������1@F���o@��*v�Yw��I�x�u RA�Hޛ��0 $F�|�K!%3E&�n��b�o��a �B��ox(�Њz Y�2@O�_��A=@�(6�c}�����8�,#-����z��`*������8^�P.8�[����Ԁ엑`��L� ��_̰)���\<>�}��� ������ؑDE�oV[� ���\��,ly�B��\�3\Ksk�|��2��@�Q�-�p_���N\�Q��4�E��Iuu.\S�-��~^[��9[5he�V[*��n���Px��͞��9I;�Cc� ��DNcƺ�n��7Α��̷Ga�&���5u�ٌ]M9-���X���. �{�2�8,� w�C:��z�+�4�1�4��&�lQǍ�U���`ezXj�mȧ�ћ��.�i��,�
�fv�O��0}�����`龬v
/D?�65z���:�!�ߌXy�S����r*O����/��H���b;���[3BvK��JY��3�9��|P�(C��E��Řቔз��=n�Ә7�nz$����I*����ɪ ]�a�Ҋ�(~@<�l��*���"�H�9��YB/��&8�H��,z�ǖm��U$%G�4������������� y�:�!^��_J�v�����mh�����L;���US���"�8o��.�>��H���0�#6����P��>�`sj>��UVݧ��1���&�"/��m�zg�XE:�R���"��r�"�@�`p�������S
r*�T���,fӈJ�Q�L���ٻ����	w$b�x��C&�;5W����k���5��駛�7 �n� �AL�"���4Y�`��)�U��Ƃ�H$����z��
�`c�X�5L��_yf^�����[�1|�q�n�^�0�e{]�<@�nS����z���q��|o|����y �50�S��f�ѫH��Wȼ���<�$��U�{�= ���@��X�ɤp��q9�3��a�@)z�����â�o�����L=�gr�Q�O�و@���IP���f�7&��Xc�w�cC�'����:`��{/��\�"1+*��Ơ�z�ᄱ� J�Bc�U�6-�|>Ž�'���}ݨ��奙����,���p795��17��`�3�9cG��8� e���E��a��d7�70\) i?>��u��2P|�t�C�Q�g�\�����0%{�dČL�>H5��A>���ɲiI4q@�F�^����dɔQ+�mZ�Ed!��2_��M�/N���^�~�^�;dg�5>������Z>k�!�FN�v��^��
P]�?�=O�aUq�RB�t�-�,UQ�.��6O�P��~�h�7���$�Rk6����=��z��[��+�nb�eI���Y,WQ�/@L��j�y�r���-�c�����0���a�vD^��57�������ff�{
�	0�w��@��GvSc��eG��W��U_�+uR�:�����+��@����և�7 �8z/̦����\��h�<e��4_c�ѭ7�<\��`
�����Ћ*��AŨ A�q" #�;�gT��oA��n�e@x�s	!b�5�0$���JA�]B;0��0D�t+��e0 �2-`�'T�зM����k�T�
s�W�&P( 2�H"�$U=�RUlO�@L]�gPI�`(��� $2��1~@��5O5���f�|��e�I��Z�Z?��1i4�"6`& �գ3%㐹� 6��fr���U]�P���w�
k�@æ� �Yg^'d@A��Î(\/d��c�f_>��5إ��ZZ����M=��	7�\{_�R5?=��z��a !o��b���P-͡��دԁ4<������X,�4e�⡛�;��@���&��WSڐ����	�"7���14�짳�A�|#��(e�P��!M>��`ǑՒu������N�Y�k/��q�g��5>` ǡ����,���lU����k�y7�s�s�������~h�d^3r��i�~ƫޔ�m 5�4FtC� p �-����&bq�� g��A�b� ݭ'<���&�����
g���c����3_�s����Ѩ�e�J4���
�i	��[&䵠�q'�`�S�X^�'�@`�����S� ��|J�XE�߁���r�^�o���HwZ���?���x���b���1:t��/�"�k�`!V"��+4����6k��< B��{ހ��J���+5`=Co�
�\�3��dw|�o�?@\�W�!2��~~�	�Q1��7����EO��'�p��r;��즍�%|&�����Q�Gp	�<� M5�<����~�4sFA����"&?0u0uyPv�<����F���0���oV 
2�Ӱ@;�MbC�!�B�y��v�X��f���g2 �0(�#�}AR{�9o�~N� �|��=�J > *�B�b�l�zF��;�?������	vO�@pE,("��;� O�A�� ^z�ݚИ����ޡ �32�1S�� 
(�[��u��@�Ð�@˂��5<�DLQ
.��xH=���r��G�#�:q7|�������{���|9��/�h.�ij)��j Y��,o ��Z���^3��]���A��(���>A|qc�4�ӝ�A��7���P)8\G����������_�WЯ�_B��}
��+�WЯ�_B��}߇���d�����(���Ά9�8 (�,Z��)!�p�-I�ъ8K�$�Hh�%�FE$4b�ţ	"�1Ob҆DO�N-�������nte��na,70��K�%���s	a�����Xna,70��K�%��`�/���s��
��+�WЯ�_B��}
��+�WЯ�_B��}
��+�WЯ�_B��}
��+��8�US33  s*��֏7�C�B� E�����E�`S����&�pB�tB<���h��i�@7!NF�|z�]%�|,E�DiHϡU	p�B�+
m:��A#j:������k	����A����A�GU�W_��C��� �&(Qmμ��QBO����`��E����߯Q�:��s���s��J��s����ľ%�/�|K�_��ľ%�/�|K�_��ľ%�/�|K�_��ľ%�/�|K�_����t�sV/Z�a���ϡ�v=��u��ٯ������D��e�/�l¼Cpgsn,��2j�lζ!�SM��m�����-j��0�j�����a�l�����I������j��wi5O}��=�!G�OH8�~#�ϋ��q)���F�]XU��a���|��e��\��\T�Q�+s y��$�۳�癦��ʛz?�>�˪��R2 9����ħ�3���{��NWWrҏ]E�n�L8���7��v;�&�����{,���Κ�_�w7]�
%+[k~\`�V��|��~ޥ��ʦQ���|�_�i<��Q���ˋ�
>λ��~Z\�eł�c�1�cmD<]h�Em��}hj��%�B{i@~1��Qu����o����u�����S�2����|}gU�(���.%=��%�/�|K�_��ľ%�/�|K�_��ľ%�/�|K�_��ľ%�/�|K�_��ľ%�/�|K�_��ľ%�/�|K�_��ľ%�/�|K�_��ľ%�/�|K�_��Ϋ�l���������^�1�~,8>t���?7b�:2�����T�g���4���T����������-�8 9W�&A��x�������w����)`�� 0� WÂ(O�5]��$D ��'��Z^1��:d�C�� � L�WA`(��D�v&`���L��`���{z�w  A� ���O]��}L� 3���y9΄�4j�ϊ@�Zת;�������a/|���Pf�)�xB���lX
KsdS���<?��[cG���{�, 0��p��l�p9C=�#��b���T
��� v~���ك;A���}����f}:��x�� �A��C�)U��|�Um��|oϙ,	����B��@g~�,����ʑ��.h77� (i�M����jBK���~��F |�O̸O����nN����ߑ��  4@��:J�wu�a`��6m'���~;�[�(�4S23���C��/5�m 0�E4NP	�v��� 1o� `� z��1T�Ax�0��PS[�.���d�8	'���%��H�I���U�� �}b#7����DXr5����JC@��w�h�8��p�Th��b<`?���� �|	���i�%<W	�,���	Z�����G�6^΋��d`@ HUЌ�נ�O�&ˏ� Ms f\��,4O��8�{/��b 6�y�Ģ*���sU9����Cz�W�Ǩ	6i�F�$Q� �|Q;� �\�~S�^@@$Do ���uPwg<D/�)P�	>)�C�$�a+y����3tftM�H@���C �]�^�W����*ı�"��<y�����k�h	4��������@gKE�? �(�lp�}�>��/�0vHm��g��7ץu�`���GP�G♃�P��uh�� ����.���U�K�M����3����$ y��`��+���#�W�Ex! ё���ǿ��{Cb�杠'[�lȂ.����&`A�8�&
O+�'��Ό6x�m�dA�U	��FPv��<p��wi�g� �n8�q��ӵ�{��?��G���/^':�ŗs����gN?��a�,��|�6Gݡ��@��n��R˛{�l�̵��41$Yi�k?7�� i�N���J%Bt��G
���8�3I�>xO��<I�cm�9�l�o���`	?Lce�N�crj�2�� �O�䟖�o6}���/ڤ�r�Vӵ�	�w����'�?�� B^���V,�W����z���@5��T�X	&�l5kP�+V�8�j�K��uT�
�,Αm߯�ra�ƛv���n�a+���ԩ|N�0c^�V�4('<0p�w�:��\;�+5&�{F�O�TJT��L{�+)*��I�F- Ҟ��>��L�g�` �b`V;M�e����H��/p���>NabSF7��,lr�����V��0J�w� ����]_
��{A+	�N.�#�s�>�p8�����
�I���xD{���@k]H�G,�����s�R��F-_;����_�XxX�?�|��1i}`
dRe�#/(�y����g[k�N�s���_K���7%_�*In�|��"�}��{!��LrP�O�4�e~�&4��`�����'�\�΢��0d�DiA�/��| "8�_)tJ3��.��O��c�q�nE�u�x9r*�F����H�b\Va�'��2�u
^?{���:����+6HI2 �:��/�[��lL>�'<��JK�/�(�vJ*��/b�E@� ���G��`9I܁�	jOr�]9[����`S1A.8����#�� >�HT���7J(�{4 ��� ��?�x���n\��� ��D���$�~`)Ն��_������\�C3�z�m)��:�%�yM��F C���2[�����N5�r ��9@�;}3 .��V�z@.*G��f�SKs!6z�=��f�#� O�
΁G��j`l2h`p���+_y���K���b`�A`2S@�I7������?�S�pE�$�Y`��b̀R�Y�h�Ѡ�(E��0�-� /Պ��J1���I�H����8�˰��m8y%��3#���0	�K�P���Jҙh�?�$_D�ſV
�h��1E����,|��K�����<�vf��9 #9�Sp��r>���%IA���TaE���^Ł䢹�BV��r3~	`c�j�2k��4��2�E���%r��'���8�g KZ�A�n��� �}K��J���T��G I"�?'������G"� O���@sN����n��Z�4 �j��m�A�}f  ���|�&�!�,��� $ֹCr@��L9�0?A� ���ê�)Ub�g���vRm t^�&��a�o�`�Y<�����q?�u��,e���?� ۳�&�p��@��͢i��:^ �1�
�p4@�p$ ���T���@9�m[��Y��K:%~���O�e�~��\ y4s;�������h����]�C �H'���~����P֪Z.�?�v��%�"�'M�� -�� ~c���#�vfJ�=��W��`O7�%��������/��l�ѩwd}e��>�����s��`�[�sB��dt�4WO��g��GV�X��sQT�>L�� �G��5|1�DT�E�E�/\_F�|QY�V�:������۸K*�-���`���E�hA�`A��ئ���ҷ��ո�V��9Pӷ��mSV�e����VV6A����54�����bw���ެ[��^U50�v��ꚻ��WU���4o�
IǇ�s��9�_�8x��B�����~&�S�:�Цu_{BS�)����M[\�T�Uܢ�#�ɽ[�ھq%c��{8'y$�M �� ��{� ��V�7)�����]܍u�
�y�o��`����ۀ_��弒k��!�c���/�|_7ԏ��.��;��誷 C�n�D�\��.��6Aw��q̆fh� ���b�ZlV��a��l�2̷,�2̷,�2̷,���fXl%���zץ5��,-/|:7��u��1�F�z�b���۳����!�O�!�G�1ׁ9 A��`hN�52{����BnH�S�Pjh�D��Ӣ�ڀ��6�٠i�����;�����v,�0��?<����1a����2����J��Lb��<�Y@�B�h�!M$����w`��º�Z�ٽ_vPW[w����$y݀��H��JL3������r^g�PD�G4�w �F�+ւ|z�A���1�掜�*$(��?���(&m��w�Ƽ E�o坋�@!:�G<����Gᰳ��s�ؠKDh&F�v��z��A-���?�-��ZuΨ�`r	"��A���$|b�ަ�5ck�L8:�~a����EƋx#@�0nM�;4����b��]q]����&k��<8O"J��&�[�s\���܂�ȧ1��#N*i��Y��ϴh�8N���
�U����Pa�����zA0g	�%���%���u��dl�@�}��yb���,��.��?w��ORNa�0�9=J�R+�!�!yX=`\X!`"�o�[ޘ����zG�3�=���L,�����7��w]d�%�Hwr�F��a�Q�	� *�!��Z��9?KЈ{��i�`��\a�U'T����$�63��`]��|�i�@�Z4g�v�O��(5�����P��$�'���������/}<�R�~�:|��4/�ᶂ�(H�@j��Óh�C��V�'(叴�ġ�@���8�ay&>c�,)�h(�&��2-��#�����Ďo�(]�+�e�`h��e�v�ʌ@�%�V#��8Ɉr^��W�ch��$q @N$bTI�u�/Do~u�@H�-�"%J��	8������	ap�-]�@ Z�b]| ��#⢮ћG�I-+v�Q(Jj���3���s,��|�������-�_�I�M ��c�>���G��]�"� -��Q� �A���~V���8�o���`bUX� �U&0��_E.�Xց|e=h�V`��"�h	�����5,DE��+��te�ҁZ�XN�KF4P LDw��ۯ���Pz`r�W|;x��+����[L�5}���<%V���	�3��\��g;A5*��w�w�ii��E��H: �Ӯ�E{|Z]�������}���a��΋1U���:��ϣ���򷀽��R?��9,n8�Y��\p�/��}�l�:xT��m��!STH ��6@��*�&C�����*���ӭd��C��Z�����ǁ  �N<�$�l:��
��u��ؤN	�;Y{�Q�r<ro�2��vd�Hm�ͱ�J����|m����J�Д��.�����V�r�x�|�B��� �<��ny%�@�'����&2ϗ[��~N; &j�>`�b��4v�� �c�x	�>�E��6 2.�o��[ ���pzX=J����
����	�XъW;���nn,ج*�X|M�y6�+��Ƀ�C��?q�����	�Ɛ�)�����`y� f�a��(��`�Y?�M� ����Խ��$m~�c\ڱ� �G^����wGƟ����
�ڼ�� g�d���d�X�X�@4�{��OE����t N �xd�W���Z� L��۠�\� 9I�N����W�v�a&H#�J�v{�N1��Z��8���8������� GB��	�ڟH�H�i�Ҁ	�1�L�q�9o������!l�	�ӂ��5LzG��|x� �����05nS�' tv���H �����R@��D!��\ ��v�����B',�8������/��2*zL��}g�����̈́�	�QT���H�-_55 �hn����s/��`WS�t�
���:����U�>�˵3��!?���q�q�a������:jU@	�L�?���w�ݖ�`�
�e�o}�O>4߲0�Pg���yL$�}b��$������Ǔ����Pe/��C��UI�*� *Tay\�G����Pc֭��
&[� ���D��џL H��Z3��@�rq��9� ��o��i��/��[�TA �ˠ?��Re�&Y-2��a���$�3���b	o�C�` p����� �[�T��H�c3�w���	�`J&���?i_#����' �>x�6.>X�|�E�&,IJ�B(E޺!�f�1��H�x��L�� ��i䋶Y�x��`� $y"y�x�֙8�z��4�p>Zgv��Ͷ/K�?�j��o#�]e׋N�P(��i����HVy�(�II�vL��M�.r�eJ_H���=�j�`�d�v�y08h�gzZ���}M��>��<�9�X�D'l�0\RR�8c%j
`�>V�[z�@���H�Ofgy��]��hi&��ѝ�.(��n��5�>�������W@@��}?����'� ��W�f���Ww��Q���-�8�<^�N�3���t5Wq����pҾ�qho>��Ks�1j)@w�(���o����xS�b�����9G�W �36�%|����l�jBu�d��WY�_E.*�S�V���Ybi�>s,��F�U:�;�þhp�v.x�2_� E}[#��3/�Y�P�ۊ�����n���1vO��\}��>.6)Mh�(1s��>|���
r·>�?c$j��~�}`� ��~{� �߅�f_L�V�Z��VZ�T�N��6�6�PV.�V?Q>����I���4t��MN�Hya�ص$Ih��RȚ�>�n�1���]{�ب)dK益hj{���%�a�$��w*s��]9������u{(��*ծ��W	��Y���Kc{5o��6�!I�A�dJ�'ؗۑ�׭� (� �J� �ѬŀI�<����{Lz��TdMB�b��{�"�w�:�κT��,�Vҿh����i̽Q�� g�,pޯ�=�+c6O�&4�B0b�$�+�*��E|�!DU���
'U�]Ł"�����
c�����xw��}�1��<�;5�$�T&�np�Uעy �� ,Z����>�i�} J~e�� �����u�L��}�е�@�Z��d�6����o>C���B��ë�@Q��
;�?!�?��W1�ǬG��Տ�p*2�{`=Μ.
"U���I׮�+�_$���@���b%B�ɳ_���KS�f���_`�#g�~�=8/�	� ���'��ބft�qp���n��<	#_FE�Rn���|�:��C#�U	� R3�5X�#�l?:coǕ[���)�'�d�7^��@�@��Dμ	�۩ʓi� �h��@���3� +�E-��H��7[;�Hp�@y��2:��O�8/�r�� ���Y�,mI��
p"��w�C�������|H��F��c�#��z��[��J��P9�т���n )* S��&g�S^bA��	� �S�
B>ۻ�hǾEB�& l����1�I�ف����K�+����	�V�� ����	���x߂�yL<C2��:�D�9T0��D[4�P� ����S=�5�̆�� ǥ�8sVE�?!�� Z�_�`�TD"gV	��/S�% ���A�'ڻOb���Iΰ�fDY�!�&���=��=��3O�	���z���\
:4����EB��/���FpGl�����%Ղ�^!������^cP7����Y;}����Y&f"5��P�����
�l. �y#1Td(�W@3����SV�ri�v�+̉k�bCU{}Ű�g���#{@����ctv��F�8��X������(l%��KG����',ґ����\�$E:?�"4'��]�4�1C��%�]����@��9�������:-%�p1����Z��PN�0 Qb��|���I�����C9��y�
ِ�+�4�*�Q�8�S�>P����^U��� X��������2��-���P����LC�O��!�
x,��,��#}���aߚ � Ul%��@��'$�p����
�}���%��2�as�	�cX5�KA��ۤA^c!C�g�#�{;��xن�DѾ�f��Ng���(�|�d
��4@��?QQ��w�Zؠ��V�hQ�0K�D�o[q��@�r�q�����v���@ � C����P,=��*��4�15��ޠg/�G�A𗥍�$~5����Ma�*<�\ c�ױޠ4��̪
8@������6�
��E�8�?�X�<rt�C�*S=�� f.	T\ [���f T��+I�S��EH<�x� Z��H�)��]����"!C�l���I60�|�8�^fT��.�X0�0���w��@N!/~��b^F2B`s��1���N
+�[G3�
pr�`MSw�p�@G�nIY(��OJ�"��
@����F1�/�vzq'- e	����� �=M��-/:AJ�O��	-�F�N,�D/�g���������NQ�����hQ���Äݷ�����S���O[E�Xğ�~�˾�~/Y�k��錢{���G�{:�@��ۗX��:�;���h�_�À��-�b��l?�3�Ӆ�/�~�`�V`<xI��,دx� � 0.E��oـj�����c��P(l��6�l*�M���k:������������l�A�p�\��Z������~���	}�[
�Q&�������� "���vo`����P@I��([F��E�/��{��]f3�-c�,�6!a�f��]7r��o8��ɒ���w�V#�a&�l�i!+ b�C�	� ��6^-n�q[0X�(�m p� ���d�	z+A�yQe[kq�\ "2{��T��5�Z����^lp�N�R� R�i�f0��c�(6 fXL��Af��O��f��'~N(�}�4����4&6sz��9�2>�a��ǃ` �,?C�(+f�&TR ���5�o��-�D�^vX�� +(�Z�tM#6/[��x���9�a�s�����@�����4��O�X�{j{�%��k�w�A�hy���Pl��6R�嗬�Ym�ֈ4�����~�8��{�F
��6b�埭/��� `���S��(Q���󡺐6X3A��e
7�s{�J�4�;h1;��E�u/j�`���9�W���7teė��Zc�Х ����y���+��u�<'� x+�~�E^�T�wW���hN�_��40�ǲ4d��@x
/څ�Ȧ�l�W&;��7���b��K�~%�w�	�4�Ba�"���ubn�r�.[�r�fJ�������a��W�Z��1�(> ��!�+Wr��ĝ��DHp��y��� Y��_78��S�Z����Y��P?P �i4�����YSS����)�Y���8,��]7�FM6x ԀC<{}�e��'v�i��ܱ��,�G�� T/ к���f �R��/'6P�X! "��̏HYG�B�zU�D+�
n�(��D��8'�׫(r˲6���%�Р@A��Ԋ +� FAK���jq!��-J�=���KPk�C@֯�||xhj=��5f7�T#���[�0P�hT��ڮ� ��'��\ �_%&�N@?� J��ZQj�c� ����h сG��;��@�#���%X���}��G��fА-y��z��i �g�~� ��w���a�Åy�� *k�(L�pE@*��6�-���d�/�
2����
S ���>�(2����{��u�N!a��ar�QsX�AN%��a]J49tIN���t/���G:� *k�>�t�9�lV�K�l��£���h�Z��!����-NRrg��SH{����P�����Y�����A���@�~6�pMA�	��ŃB�%8(+��	%�C�� ���h.���LXb~u/����Q,Ӛ��t�p�;�d �~�av����q���x�7�!�� C��IN�Lr2!j}��&t}xAƁǷ�+X�O�_�RB�A�G��N$�~ȗ��5�����ŉ�<��#�p�����X�	�Tsҗ��p�߰`�9u�}uq�h(A���O���h%�1�\H ��p�K�Mk�������  ��iu�M&�[���5z-�W��h�z=�U�����-�̸��_l��.>ָ��f�)#alXՒұ�Q����A���C�
xW��H��ʐ"�%��,,,P�A��k
R-(Y�pP!jX�;�x�_������}���;�w��R�w����2M�����`Ç
/H�VW�̦U-�2��V��t0�nz���?�,�c�πE�X��� �t��tr]|�QAAz7�_uK�vV�[�Js`B�� ����K���t��=�X�ˀ��9/.��d�5�� �c�a�cU�%��� ˒m9�����#����Q��VR��G�o���=�/ڰ�����jv�:M�y]YY�y����s�6/\�yG!��a<��������^�V�13O�vv����F�R*,-RZ�����Q��`�^�Z��0���i^+��YJv��_�q�`��d��ڣ����yaW�Wo�:EnY�f�A�B�C�����M�J��~��>�c�?�3w}�)P�:�܂�A�g="�la�y��C	ހT��EBܓ��i�����ؚVXc���Ɇ^�ES�^zA^�g��ܖ[op�~)-$,���z8$!�����Uvn������nq�ğ�{�@���4����(���x��?ԯ��^B�����+�`��S[��M�������+���۾Ci�ek؍�W�]c�'	 ����6���i��P�zqUQ#⻯�\Un��1��d��~X*�x{	p�����d�8qt[ �EC�O�V]����v;�@��f�<�En�A,��'Xm��2�2gq�Ş;��IY\b��,*�E��Z���)������p��3UU�s@����[���gz����7�/)FP=�V�P,1ց�
�J�+[p��wm?]�L�=g�[/Zk�57ى�QQ�$ҕ�zȬ��Q�H_\$�e�mZ�}GzZ)w4Q��G��Z$D{�<��2R�X�}sh�i��0�����T�3��Ɉf�����,���v�1
N�_U5�6Ja*N�>軿������Y�	�\Đ�% a��'V�A'���Wi��#��Iw�(iv�li�"��S��H[��,������1&��{�oԿ��s�T���w1Ԭ��fݸ;ǧT%|���(�����#��;�6k��d�����Y\���\��ѽJ9=)�r[��/��z�������L�� ���c��+�mC�đPi`_?֧[/ż&Nl��πǚ Th딴hE�HJ6��-2��&:�>�E�����4�-s�wFL촜d/X�C��qf���"�5^P:yl��	%8j�U�lч���@υ�@wĹk�V[!�"Q��)b/�⏂R�,�|��<��;�8����.J��x�S����t����h����^��X���0���T�%@G(T�1������th��n�8N
/XD�����izS���#�?�>�� ��������T#���V("�312�ǜke�&�(qHK�c�E�����`d�',���oN�_�ί����Т��5:�Uu�) \ ��6���s ˀ��Y�]/a�2�!�=~z��eIN��y𖊾�C�P-/�fIϯ9�g�[�A��@W�}d��\�S�n[���.`,�eU�Ya|�
j1���:%��V�C�o(+�� N�v�c=:�^�DN�3�#S�3�����p"o�2��
�)���7�ۋ�DY���{i� �t?l*�s� sϜ,�_b��,���� f!2��j,��qT���9�+®��xs��iyξwq��ᶴOq���/0�Q�M`:I�V籣�x��������W]GK����f��"r �Z�!@�(ȍ���h��o���[u���̠\��lm��=�8m��jK��\��0%2�=M���r���Z �ɷ�>�E^�v́���	��W����� ��+U����M�} O�ַ�������N�C��)V�&8� �B�a�q>>}r0龭W�.����>�	}\�(�.L}`O��U��Rx��~  |��>���|��>���|��>���|��>���|��>���|��>���|��>���|��>��lS��kW��&��F��� y��&�#�����ƌ��%8���k�i�� ��>���#��0�\>3�� V@���￀��P�@:2��} �pB�������. �;K�}.߈C�T ���|`$����� ϡ&q2>� �� �" >e�
���� �U��� ������� >u���� ��RB�FJ�&J��!1�%X�%(Ԑ�ђ�K��jH\h�V$�R5$&4����U��O�9��)��l��|����>d�!�ا�O��Չ��>c���׎�'�^;8�	1���I��'�DvQ>�	�׎�'�^;8�	�D�k�g����UH   l��f�BMM�K,�����`�jXނ7�4�:a�4BD��sBK%���Y,t[k[��L��m@��d93��s��f}���42�h%�>��x��Y�������he�>��x��Y���g��sWn�>��\|���m��fXe�/��8*�߀��ϟ>|���ϟ>|���ϟ>|���ϟ>|���ϟ>|���ϟ>|���ϟ>|���ϟ>|���ϟ>|���ϟ>|���ϟ>|���ϟ>|���ϟ>|���ϟ>|���ϟ>|��w8�'�ۏ����l�i�a�����wg��8cu�}^���p �]>�־�m�gO�t�_���y��S|1ڦ]�� '�y��yT�� ��1��=�s߀�W�'NR�-� (�.>���=�-� *򵀏��=�{}���^�_=lh��� ����y>�z������o�U=����U��)�� \! �ü�����1O���O��U�1��O�.`��p�����&������I�Ǯ�e�=��?�_���x��ծ��p�LK�@Wd���m���~ G��>�߽.�d}�v���� �^�I�D�]C�6G� �h I?�^�X�}�.��h I}�~��	/����ۼe����O��N�>�ߙa����)��W�]�K��G��ӭ���߀��ϟ>|���ϟ>|��q̦ff` ��5j��@��lږa��tG��h+�
��t��nZl(}3e�pR��k:�t�0�
��(5�	���с��aѨ�P(��흜M���.K&3¥�%:08�)�l�M��D�iH�F�ͫ#f9*I��'#`�� ���%)��$%h�D'L'h&�d.�)m�Z5�_�$�X%l5%�A��E��0�"�dK��mm^��n���<���/9��<��y�9ļ�?�s����/࿂��/࿂��/࿂��/࿂��/࿂��/࿂��/࿂��/࿂��/࿂��/࿂��/࿃W�W!����oܸ�,z�:�#�,{��},�w�n��# z��"����,�G/��q��A����g�p���d�=���n$"��)#�w�>w����{������E�N�����Xw-��pǼ�Ã�Xw/1�?�{�Cﻬ{����u�L�7/c��;�Թ�m��&���`���w#NV�z��N���Mz[����]?s�oSx��%��/�y����sB�����7-�	����`�#F�>�}.G��!8x��o���m��7ϭH7�^�����s7dPo���z����Z����a�!������oDj�/�ˬS��?n���Z!�"��j;�Y����M�BQ� r:61�34������'c�s`��%ٷGG��ý���1tb/)#����ؐa,uD�����ha�K?'΍�lk���zt���zU!��������tӖ��~�#������^�9o ���<\� ��E��v~w��t@������m�3x�ɽ�/��4i�0x]����i]��C]4G7����2�1�������7[g�FML`�X�������z�=���?(�]g���1u.^�U���kA�{c���4�O�c�=b��� ^f*B� ����C���!I3�3����2�gb<G|JN��������*)7��#&X8�����#�jaLf8մj8ń��pG� 緳�W��Q��)�-��Wi�ハ�Y�d�~�¯`En3�fx�<��	�se0;L}E�.
&�a)��9۪���1:0���2=LF]�n�DO�KpZ0s���߀��w a
��{�M���
��x��%n�N�@O�������^��� B�1�L�����GtˣǤc�%�Q�d����{?X��̤f����hdj\����z��n�㘹�����y��B�A�we]�X�{5�?�XyT�\tj�u��5����B#�':�a�F0p=Pw:�Ch�� ��l8O���4��B������I��K�4tƣ�tx����;h��l��:kMt�e���X�0Fq���	��asz��ɳ`�p����p����`4F��l �^w��XMj���St9�kQ�u��Wq�A�:AӤ�A� �$I�� �A��F��;+� /࿂ǫ=;�!�&L�2dϮ���{�qDz�7����T�H�J�@>p��{)ŀ��������	����qS	��u����i��Al����*�1�2�M���3{�˸o�}�
����_p�W��V�/࿂��/࿂��/࿂��/࿃�q�ԙ�w�oǶT8��<�=�ǱW#����v�D��R����2�l��H����I,�q��=�R		� HpO�ˌ�\�e�愭�B�\���hd%�^ɧ��$�r7 R�m��f��<�x`?�(#)��4�q����W��/k k%�D�!s������kM�2ı������r�Ab��Ăc,�lBu����E_�-鋚����پD�x3�������&���1�(�Wr�6d����t�=��|��[��EO�����H��r�RhJd+�q�2�8	����[XbK?(��j͇'�__$f։�OsÎn��?gԀ'
X��A��q]j�y�b��W���W��㓠x�R:_���~x����(���[�Q���֘wt��Z�'@�HJPzu�ٌ�y`% \���%@�!%�_��ޠ��m`a��9:��L�~T��J���c�¶�l����)4}�N<@��I$�~��2T
��%�>B�@C5j !N(�@�(�+��Н�4���4:x� 5��z�#ݸA�C;q��`��� �k��{���H<���U����W>K�� 8��=��Өc��^�%�:|���P"��j�(����ly��7�
��[��d)UToy��J���$����=:�r��_���Kaq��
뺕�k��j��gJ��Du�|���5���+�~�9;�����l�dXw��6�]�9@IcE��p���`�Y�E5;|WLR����h�^M� �叞o	�!���_�M�`lb�rM��@�̣��iP��.������;�o)P+��[�s�y�qb����T��zQ�:P�(�f|�R��t��`�����jj����/�vZ�5����w������T�0Q_	@��6�XyY��8H�$o�ŹYPT������&���]ʌ��r�v6����y� �|Xϲ�L�D�ϊ����O>Z
�i
��k���j��m�6��+�ւ&Iş
BT
��k:gY�H+�=�����'u|��J>�s�!TA4@��=]�ez�rAS>�E�|�Rk�J_l�OG���/�ݴi��od
�8 U�[�[��%  ՌZ�~E6��O��8R��+��Q;���^Ԁ�;q�[�C�i@-a���3��iI'A���'g���,�'RF�E4�@��"7)I5C��+Ӂ��4���n� A0�B3p+@���R}}�m�K�kt����� Ť*��j�Ύ�H�
�	�Ѻw�npl���Rp����#|�����,7PE\��7WbD�E��?b�I�T�+�nO��k����![)�)T��Q�lH���A�f������P�iAD�KP�'�|��-�K2�hۯM񂹄8c� L �����YXB�{�Z9%�9��@Z#�8ygl���Ě^�湲�'D��	x��L#��c˚����h�T/	h�;��oc3?��/���5����-:�[�M@�f�gK�
L%����� ���X⸁�H> OT���?K`sut9��n ڀ����{�a3߶���ż-XkM?��!�ܠ���rp-s�d��|=]`��I��( �3���4Y8�@b�U���m�i�NcRՐ�(9'����h6M�z��`-{�o���3W�$&L0�L�6�Ź���.��*�d�a� ^�Myj�kP�y�Z]�@�Q�SK>Ө��g%-	8��mBmFB�h�J ��I(�]B���e
��7��{�mN*2pI(u%�G�T�:���=�
��@!�m`��Ԡ�n1W�����$�|x�*@ON���@��ԐG�$*���?�,�9���˽ѮW.Mt��:�����%��7[��-��?���}�D@v:� ]�u鼼M���}?�d}��/9�Ok�@|�9�1'&���+˰�_.���@K��)r���Oa�Zc��U |��5]���_�s�i���k�ㅛ�2�,�=F߶��x����R�RCB���1t����e7a��<��a�4�IC��|�B�H�-/�N�nR�Pb�� _Y/�t��q{~k˜��\K�����O;�E��5{x��yT`p雴�[C#2p���;�p����5��i��]�2�c�띾"g�[��Ko�0�ݕ�p*S1z� ��n2Q5ٛ�b�+NM{�w�X{4
�ڕ����lP ;�-���*�<��#��>�Y�W7���?�ZXͭã���K�����:	�vS苌�'�j)'�:�Ǆ ���b���Tv��H$���%V��Ͳ��֦Ak�D3�Q��Vw��Q��k�۸w�����;s4�����B��,a�7y%��������z��0=R�QH��>B���n�џv���T�[�dI9�@�+����mq�xFR}i�z��P=�}���Wf���3�Y��~Ցi �U Gʀ�����O0p}���E��G�̹�*G����Mi�m�j�Ȧ�(�~���N�ԩ�rmu��K�Uo���-��_E�d3�9Flm�=��h	D�:�<WGI#�b�"�<��}��i��9;�0�|� ���ZrF��:��׈sS����~_�k�X���J@c�y�c�I?���/?@�36],o�E�e���%%oط�/�U�Đ�v��_{��(Ĩ�j���O���xێ>�'?��}|NF�W�$L^u����$L(�š�e5�D����+
�{/��[��+7�;v�09�f>y�k���2&/w㱙=�|� ıP}�S}�e�T� z�}��,��e�$��:�8���T�ey^�0���F�t�E���'V�����>b�`8.��}������l��`7�� ��@7���vq#=7�4>��A�dH�>�{��@�����+�S#YS��*�&��Nz��]��d�܄@���}���`�m6�c��E��i���<�H�T'���N ���a(J�7l`��#���H,	���~v&B��+��L�͜H*��_��T�rT�Z�/`j���f �o�P
�d�P�G�]��_2��,,n���/e Xx��ؠu����@.��w��.uS:�Z���uv`�����ueO�m+��
�����I���R�ı���bp�@)���^L) ��s�~5�rݖ3ߓ��uRLi8.zu�#kr[!{h`�� ,P ��}���X�~/}�!	 ��C64N�
&@]�U���;��g]���Ѣ��g����m	j�!�<
ef= ��5yM7���v���>sK�=C�D\" H%�a��� f1Zj��#��Y��1̲k��L9�ԓ��F	�O@�de ؖ#��`�p��4c�R�;�A :�&'�p$b%y��n2���_��d��DI ���b �%�FbƐ%hַ;�-/.��J��Ղ��Wk�\�@n �y�d������\9�cSFvD ��U�݇��ǫ��Y��L0��x�v�X���L�E��MP�a�\�g����h�e��V��Pdq
�023�a���7� R\�Q � 	���2�å�w�ҽ�VY�� Ӽ. D`�@��x`'{�@��(x �"c� ;����d*�u�`�V �� .~i<"E*��	���<�)�Ǚ@�$�U���i��U4�J�����X�^~l��%h�1�*lN\�^#�����&I��BW�	%�.]�ڿ J��!@��sB�(���Z���=B	��<Y@�� =.z \�Yvp��c�:d�@�.@���dv�*����uЀ�p'�8!s�c((�qd=�	D�.4M'%G$J.��l���r{79�� ���e���Dm���e���2��%�t�#�a�J��d��$2�Е���c
���pvY�l4O��2��Lu�a)q�|DC����	&W<�g�;ha\wܜ?iB�ɂ�ArpFȫ��!����cdeu_�����!~x
�dF��B�~X`���
U�`@<(=�'��D������d��5_�	K"[>��ɂTH�� �v�}��` �����{r{}���� ��#~�X�bkChׇ^�m��N�1�7�q�}�m>�!���W�_��}�$(lK{ ֦0��v5$����o��L���2#\�l�a�c�H���n�����G��� �;���bs�lhm�ލ�kp�^3�H��7L�#�xVg�!}{D�c\c�Y�`�]��`K�X[t/�ƺ�������ߍ�ް�W�n�T[�	0��ԇ�;�w���?�6f��r[�����������E�����r����`F�� �+�1��f��I�D꠮�+���~����10`����/�/Ȇ�L@�9��xp~�f�$���S���ܕՐG�P@:)g�(���7�$c�.V���w����9Ǻ�����-w�o�5w����_�A�x��4�GP��1���Ye��xy�VD\�R���v�<*'�h'N��<w|w�O���c�wb�ů"p���v��� �2��w��������տ�<� v�쏭�������|����uQ�Ӂ@�
���z�U}�[s�)X�h�*�/x!u���D��t"���O�����~γ9;q��_�]š	�	ݦ?���puh[Ϲ.If,�?�_HP|�� ƀY��N�1�ΐ�>�5����Ϭ�!h@���w����	�6	_�d\��0��ϯ<�Ig} O����t���	���βꞑm��J�6=�h�����Vb]��`)�s)�/yMz{��]�r$��G�G:�;{���~88�@Ys��zk����5e	���u�U �8@G=�K�1�K�qZ|3��l	�!@��O�f�z�S�MVg!�e�� [�B����w��������M��O%h/�j����.^�oku���A�@��(����);��m��\was������E���zTiY���!I�$*�;Yb�@��i����9��/��D&�[R���"P
�3��fI��?#��N��k��h/�J>�[�������c����;�JB�
�X�N~E]X��X}7eP�8�n���i�4��ic�ۯ3��@��4�OC�����P*�k��o=�A��V��L!0�*P���8�"�	ux�NjΊ~���4%B�J h�e!MAQ�`��������}�w�3�<R�P�v�TП���(�	%��E�+�9�~9F��M7b�R� ˕��(�$��*��:����sJG�h�Y����p�����dĞ�}ޝK�� Z����Rx:6O�g�.���e����Wz����� ]X�w�U��M�{2�v#�/nt���s|7��l���w8��y8WCNwV6���wM���>"�a�[�����4���P?���K�ߣ����\���B�#�}5��?�v��q^���ݢ�l�@�W'F���x+O�ۨ�,U�p�����\NH]��� �Z3`�r �/����,�q��Ŋ�"�� W��}�d\����\8���ݵA׳�PI�<��aT�
�����K��@}�+�(�w#I#�+x+���L3���q�EB�qa���,sa,��E���_"7=W�Y����+�H!��<�8��8*�O&T��T	ys�؄��h��3�<T�H���`* _�^�T78g������@*z�^wb]�]V�]�`��&/���P�G>�>�J�a��e���|`��dHG�PA� ��,�4_��	��j�?&Bt��͖�=YO���&@РRҿ��aVR%�
�J(�s]���Ζ�YB� - "d� �La 36;�
���H#��-��馽�Wu;�NS��nUgx�>�:K_>�J ��{�o����z[|d~���0�R0 �ԙ�b��,�A�4� (�/��2�;����9y�^C+���響�r��F�� �'~�0`01���ѝ[�X1��l����}�����tlgFcgG�`�l� ���0c>�``6��=̒d���`��Vg��S1��gKwl���lȕW�1L�ukz�َ+wbɶ`�$���+�J�,RD�Y�ԛ���LY�\�W���g�U]�H�R�}�_�JԷ���ϽZ�#2�)���]�buj��Y��|����������s��{���������j�A>;������>�#�G�ԩH�;߃���M���' ��������~�/��W;R,	��4ά}�B?@��#��8������O���
Z G��z���9�n�W�%��ެ������Oց��� ��J@��TR Gȫ�i<�È���Oڲ	pD*�����;�( DO�D>��N�*h >0 ���T.�J޵H�����~U�����%@��!��>sЉrW�$*���r��r��V@~��;p��7��R%1!P�	���$ ��( � �sB o9�sFS �T:�#B~[�P|@���?o�ŝr+�
:� ?�E2%C�8��N�L �	G׀#�0�9� �H
t
���::� �ɞBxR�HA�-
����v�JG���ٌ��� q@��!��iS�BS4<)/�:�����_& �x:��<�j!�@�B4�@�����^ �V���� ���	L��	HB�aR�FDR��=��	_��j�T-�3C���`)4���	>H L���iwG����_��j[���D ���*�� ��]D����;)j�� l�9� _" /SD�u� �� eC� P� �g��!K�P������Q�{�������)*j *0��8y\��*�@W^z�����  �qߥ2� ⩄J��RH� \!����@  ,4�iM��*a�|�Je* �*e u^�SD�� ��D�$*P��j�@O��>" I�<�k�bB�
©� 
����@TKaMCɻ �<�� ʂ,)� ��� ?E�~���  �)J��=.��R�o�i
'EuN)���z�,*��;x%{4�^+h( ���`��./3�O���O�T�v\�x���K���� £�iJ9k� v7�� k�'��vi7O��a��.u���	�� �W�랽�.��ˠtW�7��RS� }��1����
��z��$��,*c x �9�9^�o��j:Q§� ��߃e�����/��3ğ7y���uXT� �W+ϓ����=i���Bp��T�@3��y%�����:��tTR�2î�Ӂ���B 84�`?�9��qZ����ω߃�A��0�;<�Wg8�����O[�K�ҁ�߃���i��@%��J}K��'4'<>/��}����`���N����߃��H�P�D�&��
��4���qC����s�}x�*M��'4����N���S�x�4  ����@���s��o2#]�Q�#Bx`��+���^���5 \@��#�̕�k��N��3$�`�N�Q-�L� ���	�9z�<�t�69�v������,*c Rx��@�.~kࠔ����;�z��c�S� �cϮ���ܽ�Rpy��z^�����2YU?f ���#�.,��������Sǿ`�"Q� �nyyq;t�^�%Lk���>n7Kׇ�% ���&��[��@V��ָ^Ƥ����1X�� � >[��R��� vN�p��ԃ"}�)߮Y>p�)�����  	��?.u}����p%��y:o�S���N�p<�_ۡ,���\��w�x��` � �	��@V�n_��)� ;� JW~�g��C�o���&G)��׀ ~���_{�I� �	�	N�x8�"� �����ݤ�(O�����#�׹��W�z�t@|>寁6�8t�uK��6g�i� �7�)��3���Ie�� t�����x��辋�`�i|S�G�K������ŕ9���c{X����	(�d���rX]�v�� oHN`7�TS�F��Ά��` C�p�i D
��wO���E�'��;�)�^����	�ߓS�p"�g��B00]�qQ�4'�*�*��?��1?��	˓έ��|(�@
} �Er�<�N| )��ufnqg��s���T���y�R��P_��U	���c8,�P�t��|��M� +ȕ &�'��� � ������/���� }�B����@��#�Ja�k��m�\��+������� �S�u]=l/�D^��ߴ#F���t�����P�)遆�N_k8Ы��W�)8\.'=���"����GQ���3~�x��Ζ{�o���A��hB�P�'1g&~0�N��zo�-�P���b�6S���_v���/G��}j����~�#���?apY��z���y���6�х�������f�~}P��7�?����h�
�d�"����(��a�rO:��?����_�T�=l�
�K;���;N~2����cӑk���0�$u��U�Y��X�یr�g|� }�@����ҺU�@O�`�T�D��.��k_��XeW�x���A}�_3	���t�^�{��0����*+t�|�,�o�t��n+oݮ��ݧ�V�x���3|3����� �����E��U��������E[��=��))���h��h�'��	���4���[��<��w�K{�o��U���a�S��X�g/�ce;��񓧦�(ʝ�����T�����Z��҂����~����?-\QM�t��;����#�M�v�:"�)�?��=�*+��D�S�D���+������LJ�s���_���p�� ��G֏K�)�Y��$p�h�����UZx{\�%�
$�l�?&�{� �7���=��p�; ��дΉ��.�d	��6eD��/<�>,��W��>���{��
�t�{����!�P�"�-�����&};��I����x�6�0x5}>�f����ګ��ܧv�/�~E$�2Q:+��H?��;�r��3������W��}��U\��
ުUz�<��]�~����$��}����ૃMȫ���<�������Yڦ�+��|M�!`�z�l`������\Ao_�q�<Nwn�S	�����#�����^}����o&%�h��!�p�o��h4��կ���,�;��_��U_�<�S��������]Q9+�u�)EW�a�����������r���;�C�k�
��`�|�42�Y�s;Ŀ7��P��\S�>�)���G���U��6��f�L훵ϻ/\�2M�3絝*��k�{�YWѝ����ڼl����{;�^����;���6���ITK������o��3�y����yY��N�"vé�O��>��o�M�w4?������S���� ��Uxx���gё��鮗����ׁt)ȳt�,���*~�ڿ�p���r�N����Y�D?��%��{�v��rv�_�<Wj���~��'��V?���i�{-�縙�|^���F]��;��ƍ��N��oC����mi�_<���)o��� �i�O����ؗ���џ�o�QhU@�~Coaqe��P�t^�K~3},aR�Kץ��s�q:/��t?�(/�Q�r������"~��d�)V)��c����8�;�=��2��W��o�g�nBw�L'��{�O�6��4R�爳|�\�}����=��H��^����*|7��gf+��~���=o���ʌEE��ڭ��-��c���^�o(Y-W�1��gw������Vi�oW���I���#P����K��q��&
����5j�p�f�*�ry�y�J�M���!��6S��պ=d�\�eG,o3�G�ޛ��m^��ش�%���Δ+�pR[�wx$�C��g��25��y}�4K_�DOM9���*���6f�
<H�H�6	�՛���/*>.�I]��ۋ���E�+q>�\��E��3��ɟ0�_�ί�Й�Q�Y�u�iy�5`�EZc�-^�(25�з}&�j�]�$CQ�	�s7LZ�{栐�}��E"�01`����Ɗ֭������b?L9a�49��L_�$���2�YJ�l�ɳ�ƣVB�w>r⅝m����e
c8;�B3�ē	�A�/\ڗJ��H�=�\2���1��}#�%ڡ�H�3V� �$�������<Ջm*+B!gb\�Z�)�\J�U�v)�*|�.�2$IX���4�_.{D���& n���g<�(i�=Hi"{D��I
��4��WS��n�g㒍���_L�@G��z�����^�.$!��jN
e����𑃶A�/tt�˧2�)
�h[NWDĦ^֘1o0q��im���h�����Ɛ8�*�;Z�Wj����vB��`V�]`�A���"����'�l0y�{�UVEx�nc���Y{&k�X�y��&�p���o@)��xr�gU����9��h�����hD�JzH<�\Mt��vg��,�`�z��˦_n����3_H�f٬5�~Gw���7�Y��B�n��^���|�ȏ�����kd�e0t4�8I���C59I��(<��*F�<#�6��4|0���MVR�I�[U_�1Inn������+w5S7Q�ڐYn5��7�4y�6��=����𵢩�&��NF4���l���ˤ�?�OM:׬���>>����C��bI�[N����I9�Kr�V�=��`y�/D�nIA;���˒N�����Ϋ6���}�3���vQy��VDσ<��Y�����5*�J�'��e�[U7e燊�e:}P8G'Cdh��g5*�ec�&�x���ϥ���i�a��l`��g߯���&jDYY�����k�|�N�9���k��
���Z�1�y���.��B
����֞>�Z[�M��ޞ����M�N�z�m"B�@�-ɹ�BA�vp�^��*Ȍ�����j/S5_���������;P���P�%�î΁�i����c._�S�#7??	o��_@��FG�>N�.n�dojN���'U�f�w���m���A�݂�*���gop�ф�i��itui�������B�������6����"س^�?��tKd��<.w�n.�+���i���<!�r��v��~��#]nB���Sz��q���m�n!#WA��ޞn��9���dr%�S�����-��A�IY�NK�.���M��g
�fE�`�s��Ѕ��_������B'���g�x0�x��Fb���Ώ������	KVy�w�?15U�&���=����{���av��St;a~�|JH���e���j�?�����v�Nna�z`�g7?C�ʎ��ݦ�Ō��Z�#��𲉺K�Q�n�ֳ���e�g����l5���K/�����@�N^u�2p�D�,�2%
0j��,��g���s׌�qܜ��h��㥬&OojS��5�JF�Qp�E(m�`�X�{q�G����'%E,"CL��q��7��}~^�t(R�(E���N�5ϓ$�Yݑ���S
�tƬǅ%P"���b!R�VY{��6b��A�
b�托L��f������`�3�;�Ҫ��nM���in��>g�3$C*	�	�̖�	�F�i
�Px'5%�L[�Yo�m�@��Yf)
�qZ},Y,�*f���|۶��e�d+�A���;rRb�5���$Yh9Qv�!��5'UX'/*�\C9дGF���LB���_��W2Wu���~<��_�k���/��m5݁h"LAE�59�<Gg�<���CZqx��K�D�ĂR�x�e��i-����.�%w8��� �"W��bu�2%yA<�ni�ۄ`Gl��
"����}ΊjhYZ�fu]cQsc�C*��l�ˏ�0(�T�j��̸�T�mB�,Y[OU!��g
X�I�ʦ���V�p�*���%����LwV����pkc��t�$�ڝ�=�������ĭd�������eKF�����}��5&U��uS��s�͞V��հ���A�8�ڦ% �I�>��!s:W�lT�4�$Бę[06d��Z�0h_'1&BB��`m������3;Pvn�[�^�G�O�9MΛ��/��2�,�g���7�Q �Z5�R����@M��$�LZ�d������ы�ga�-��Ɏ?l�% ��}4�C�WsC&79����d�r6��A-ٽaU�$9X���NA��75�о��2f0�����]�Մ9�8@�DA���O�m���Sg�6W�F5;�T��i�z�OoX���P�����l��%y���E_��M¢�.�K�6�"��z���b~����I��ML�nO������� ���?/ Lw}�&\����'�'f��${ݑ~�<qd'��LȬZn�w�9my��2�m����ݍ4�)w4�8���66�6W���G��VW�(�]OD؅%�1��P�'�E�e�R�א���E�W��0&�Ļ����䇻�F��܏T�e�ն�Dc�nu���&�zbʚ#$�J����Bʎz֧s�MF��ac,G�k�1z��`6�n��/�ҫH���@�!B{���1�!��p�V ���l+;'O%!���b%zV��z���3�����Zȭ"JK�f�s���ؔI�XQ�"��e��dxQ5��n�&Ym�䍌�'�z]m�Lt�i�w@���Hp�<2ybq�.T����3���Y��w��	al�l��3Q��GG��V�\���]��sJ]�Y'e�W�1��W<���������y���2Xl��%$6��]˘=g��Ƽ�������mP�FյAwG#/���'��;�9����1�@mof�.�u�}s4�v���)�T�%����=�4�T��c,~�4�7H����`c����d�-D��깷g&W2�ؑt�p���Kj�r#��:-�.�*^��;#��GA��`\̠�$Y�C�[�/�ѲF��*:�!	���Y���t�xj�p}�c_.����Yk�<������+H�B���f2թ�V�7�"xn�+�z	)��o�h�뮉�ӓ�4Z.ҹ�+q[�h�nV�(b��'�iK��ncO���9/�CC����!~�����kĝ���w͒�f��1��Q�DwE�|�ָ� �2l�3u��b�k���������N�)21�!���썵g�ۍx%�w��������e��.��0v�1�bq[�����u�����M羢�{Ŷ�>b\�d���;�:�𧁙�.��AN�9���\�k}Q��@����ȑ��G�^B��8wl�d��WH+��\9y*��t�|���N��Y<��Ѱ���#�+ ��u���_ǯ����uI�Gb?�bb��^�,�]i�@��g���͝!��J�x��9�4CtDFtiԵ�i�X9�Y��`��Yѹ���7I�u;g�8�P^���)�3���\!�����!q�j�6ÎF�V�e�����v����o7q�N�sn�D����Ć/�����H��ۂ�N�����T�6�����F�g4~�Ep�3���ou��AM�����)^&�Ǎ�t��qu���zv��p-�/c�ш?��w����h�`��9���]��땩�Ȭ���].�쭻���АДEj�(��U"��5��f�2�bޔDN�[��!ա�;<H��f%�� m�P���E\�F���\H�s;��}x���ǤL��aq9"�=6S_��#�3���-���q��ťdB(E�K�����skn6&���z����(D,W�+����a��^oGA�M�ZIV�+v�Xz�Cu�����]V�2Zs���x����\�q2�y��������n���'që���Eӊ������t_h���cҖQ0�w+��sI�1��Q�7ʴ��h\V��v����F�ínڎXi'�a�ڐ�31ͮ���Lc:�n�� Ż��;c.G���-$�)eZ�HI{05�1��y�	����!����`��7z��ǻ<.3m�1�}B"�l�T�2|�\���:^�9g�FB�??�$i�4��.;��IU�-9�_}�4]�e�
�2����fY�9i��U�,gC%
���i��hD4�[���@���vU�~�m>����ƩV�rzcrƮCX�F���^��%B�d�f���xe}��+�U�PRv_j�l��Y.B֑�1���pj���� 1�{ny=>c�)�+E��y����с��
�Y�p8Ҳ�E�\�J��%u(�|n.�N���
��	k��y3h=6�b���5t�wh-Ƶ��)Jk�����d��f�A�R�l�[�ӕ�Z�T�J�z����z7Yy�_�m#.����S?.����Y��<���,
6���!O!� ��-��r"Y�����BP�%�1H�k0�T�]YћXV����p��'wul�	�#(������k�5��RA�j
Ǖ�O�4b1�hܛ�+�U�+�*�6�P�b�NdִRL5Z�^�qZ�fF��*QfJ�B��/��/EE%���T\�ݸSJ.t/mC�]�RWa≅|�bA6�.����]����6�9�����U
�y[�d��g��Ì�A�����sgM�"��fw��|��8�gC��H}���_�Q������J�%���+��HJ8y7J�O�:S�xk��`���sqz�3����a@�� ]��>f	K�bP/Y�V@���H_)^N�P���q*��=<�I�:���]��-�'�tތٿ��4��
۽ť�f�4>b�;����|=�1��$��~/f����H(0x��!�F�9���X� �p�h���h��Ѵ�\5ЙU�����~�|'p�Z[H�����K]"dN�W-���PШ4ן���Wv���bf�'4�T)=�z|.�
�+��	*I�0z]Cܕ���,�O-0��Ƕ?*),���W�Rv�+o��C��K��Ƽl0��9 �d%43$Ġ�uŖI���|(XiZ�[0y6�:g
3y���1�k�G*���c�����ذ�A�b�������M��V�o�P���i�fc"dT=�qFL~�2/X!F��b�tg��\'��)���Ȉ�����H���o_�v���ۜ��a�xkqX{�Sv�:�:���=�8�q��^�x[YFv�k.�o"��qY_�W/G�wvFgu�7&�\�-�|iH�*�r8'7�6ޜ�ҳ3�b[��yQ���u-v>r9���dlC]�|�H~z��G�@�f#���$I�|k�e�/�"[N�`�t�H�l��E����P�yY��#��kC+v�V.�cj4����N[��o�����47���غB6�I~)Jé	�HQ���L�g�!�˶�i#+��$Y0
IF�3��굇�eQ#!+'�㖆�A�����7`g�*-�b?A'�r�X9���c��#��O����)1V�
���[*�c�Bd��� X��蘰&'u�&��+��sV2N�Ƃ��j��U#N�+x��ݙ�X,�f���XvoBof���a|5�y�&^2⒤�oyaej�Zn���k!�v�2������W+�=P���qڸα�ZEaM�lq��F�2��UI��'h����s�5#��c�����%a�]�d��뎙#��������K�t__f�z2m|�7�ѵ[��ö�Ǘ�u���#�32��/�α�8�����V�Q��L�L�1�a����õJj�U����7��|S���d����f��oG�Y[&��o��+��Ւ�=�6�i��R�;���T"��3S�᥏{�Oa)䲁T�@�����}N��;?�y�i���sk��1�z�.cJ��î�0ոH_6F�l���5�PPR�Kv�M;�$깞`8Y�����\2�v��mT7<�o��"�oc�d�]���_�	�4�H�[� |�f��}|~��C�;%w:���x#���"E�?��]���\N��X�+���U�P�2i<\f�k�L�f�ϧ-�)�c�����M�9I x���@^�@,��φ��X ��r�0aB���՛6�}��R�\I�_Uǡ��Z��JTL�P����[Lίk�`B��)(�@N���f�UC��pQ$�P��b�e)@�[J�)��RD����e*�X��8n�ٶa�		��/'%[��t6M�Q���6{:����yo�^��AC��D�d�������1��ccX�nC�[×���9��#lN�,H���2np9	{��+��������f��Y�r��d3T�Tm�A��Y�q1'љ�	�N�br��xK��<�l:1�]ן9��L��3� �W!MuH���9��؇g0�1iLT�/�\ǲ4����)�jł��,�n���I��J�+���t��u��AXk��hL.{5�����_��?Rtt٦���ia��/���E�m��ʁ!<��$eZ,���� �Q�z��$��F��21{p���ZhE�1�ئ��X�ny8����5P   gu2D%v��y��IX�W{G 壻ʲ�]�+��wwwzY̝��	4!��2w$�2s$мќМ�>d����hO�2d�NwBL�$�g�y`�l���t�7C�2/i'*��u[���R<<7�t�ZP�vF�ד�^z��X�\Oo������M��#���c����^��Iƹ�	����\X�S�XR����F"�p�6a)��͝SCWw���.��I>�M�c&&�P�>D��ƍ�ρ�TC6���&A�~�Gm���f⢤�OW@8�A����_�-��4��)�jCH�ݱ0���LSQv.Ѹ�SGK��<��d���%�ݥ�e('�{�}ߠ�����5����|������㷅��	�p:Y�rk���8,?�.C^���uE短��>)��GEdc0c�ݢ��M�=|ԣM�Di�:�m�U�O3�¸D������qT��_]w�^-��6 ݒsi8A�/�&'�{��B���٠���v�/B�QS���h����`��G!�_��>v��7J�����������mqIw�=���W,:#��T0�v�T���e�<C�'�C�}�'_��3�˗��'��?Za�]2O�H�$�M����L��o�߂�Ʋ�L운����|������2b6oqD�w~sgv��%��{M�ܢ���	,�٥m�D���/����mUɥ�ed��΂�SQY����(���e0�7d�q+����		�/�kbΓO��K��g+`_qh���;�Y���{"��rл?w�9q���A�P��������y�1����NQ����VI���{�;��6��|C-W�S����ǎ� ��tz���:�#��9��Oq�KIK�����Ǉ�`a���/6���˥���;�֢J^ȼ�
�u�C��ձ�ҽ�e�����՜��ٵt]s]�"��RV������ӯQ��;�gzw��+�.��hm���6�<8<�h>_z2�T�����!m��X�(��Xd ���/@�0��
e��A����9x�V���z�:�ӱ��)*�����V`�K}��Ϝ�4^�6���r��B��8[fDl^d�X����� y��}�F%�Y���ʮ=�x�p��(����	�Mߤ--d푂���a�i�Pp�B�2���˃S��p�E�w�\�G��+��-�-F�J+��ax����%(�ѻ{�7/� ��>�O((�1�XÚ1�������!��f�c3)�:	��Z����YznB���ߍ%@�����`����a_�!�����\���JG}�1j�O���7��x���3�dF��[1Ljb�ʐ�Њ�BD��Ӡ�>��=(wE���#�(�����s39q�E�=�<���p�����ް��*P��&�a�#F�M���*�!��>d��D��TC��5�F�d<�`:�|��?>�F�ң yw������1�X��5��
���>L�~�^�9���f8�x[
�!}f �AK�����ǯ��������w�wOU�|�DB��II�%A�p��I�]\hRT�f�QJWV<`f�bO���k+��y��Y0�3�.���3�C"����i�k)�ts�Y$���rs�o4��\���ZҜdQ'�+TqV�	�d�F�%?eO�i��[5P�я�{C����ոd]�]{Å��!2^g�S��~���t`�{�o$���i��}�6�@��1C7�7�Z�ZT$�RR�����������ȅ6F���얙ަ���nH.�Tc�|
�#XĶ�s"vҒ��w�t%�MP�$bd��c�1zo����Y���k�	&0�͓��>!��*��}� �����l@���nr|�q1��u���;���M����(kZz����BG��K��Or�/y���,���}���8n+��,�b��U!e=�t%��&��k��E"�� 2ޜ�/�Ӟ��m�ݧ�sy��M�z∮�C�aG�b��G�wp/��} ��&�P�Ӈ���j��Æ�z�(a�H[WtD ����zv�#>��C����M�/E�w��� ���X�ڌ�+%7X���|u�Na�r-�8pJ�Ť�_5-%kc�&?��?B�;�6}*�\��|������Y'�E���9ep"��NNUGG�'5F���0Ũ�y�l�on�����%�l�\&�WG{��E��DM��2��)ޤ�|5W�ZCږظʼr?�^����Ha>Pb܈ly��=ID�{�f�1�-3�*R3ay\d8,*Fu!W������{��($_�����0,��7)�U!��vb���.�� !��_�7�9�
޳1�Z��8��"�e�$%[�h筻+�vG�Y>/����M��%!UZ`h-
�І5fu��⨤xq/�4�}K#~\���a�Zii��ڞ����I�Z�9_�dJ���;��xUp�[��eh��%#�
��w8����*p�1b�Z��6��K��e��kłx'#��%]�Q==m�B��'t�����g7M�	�C���齺���X�+�6H	��"�~cTؘ�A��qtN[����ܬ.Md�O����,�Z��I��SK����EM�T����rurj�op�Ɩ�;,��.a���a�x�~�2�q�*rdb�d���h�D�;n���+�WOUc&:�@}ރO� @2��!��qTE�k��k=Q���1�:HKY��>y�b	���e~P��{VR��f�%�^woy��O]t�Y�?�� ���ֹ\LQ}2C����Xz�pQ�iK�����{Z�"ό�|,�8��8�odȔ�]����8N��DǶe�b���I��K�����N�QQ�<KLI+�==0|�7u�+`C�T�R�SH�ິ+
}D$�ƫu�|j�o��}�i~����y��/W aH��`��M��m�"<Y>9%#�	��Qs*���$���6��=�q��X��RȌl��}=U=�Ǖ�?��qF$<�u@N���3C�[?�����g�`�0�[8�����Q�����ayr��Ԗ��ϔc{(��J�k 9����������C�М�v^���.��{�X/5Q���R�tn�gŠ�i�1.D��Ql��T�tW��[Ԥ��U���v�9��^��n���)�/��7n"zᬿF��l���Ll��]�ԥ��
r==!\'�m�Z���9��-���gxL�N��;��Lf�%��A`-�Nz��P�H\T.��Yp໖5Q;���9ۅ�$IkMZ�Kn���
���l��}<����N�Q��x>HA�+).-����{��b�eC�L��U�hĮ�i���f��ʽ���O�9�`�������j��,}�6d�:�QR=���ǰEY���Z��fQ)��&�'��תB�#��;���!��c{��ɍ�����MkÛ�� ��������v΋A�X�6B���|Ք ݃�rT�ܣ�Ai}�Y?����.�ͪ#D��P����kZR_�������H�%VO���#����(1�p��ϋ�k�U�L�D��~npFI��g㫠1�JU�S�7�V/fmp�d#^��=��������琂\���	�U��DZ)��V�a.c�\j�+*�=A�qW�ԫm�����{�8췸�s��~�T4+@\�gg�#?��������l�P�%�dhW(�${/�u��c�KN���/Va<��?	�����Y�6,�r����>!�<��j�����#��$�|5����~��%�Km>jX"Gh�!�����X���FP�dE]�W��ؿ��"\T͔=Ձa�?�Lm5�BG���x��%���rc8X�Q�D�?��>L��m�TT_�h?����G֪(YV7�OX|y���s�a  b"��o|�*�t�D��#%���.ɩ9r�HZi!��;cˊ\.6,�䰲=B
��ͭ�������5ϒ���ّ"��NQ�'}t�Bg9�˕�NJoն���c��Ǿ�u�u5��b��F1�N3��y�Aa���2�v]s�?v��p�)�{�"%B��@��\޴����������[C4��;Z���_2T��x|9����;v&�渓7mfm����|22:)qC�s�a��I����B� ���2���+���
��!�ha`�<���3
����˵�7�c$S/�{|�}�	9�t�@�L!�����}��g�Y-�V<�P�Jp�5O�cC�(�%��\�	"^�S�֝1j	Wf�U�М�G�%�����7K��D�T.�Kt�V��BC�?l�M�F��y�Aװ;Q�Z������Hǹ��aO���E{Y�U']L@{�]{1<��TAM�sY�ZC�m���{zL��"�l!o\Cl� ܺ٩b���Usm��r�����ߵ;󤕂4��Ӻ-�ћ|�w\C�#��������n��th��9 /jxɜ��� �j~}�RZ��r���W�eyk?3x�@��N~ԕ�ۏ�(�U��U��2 ���{�y��^Q@cA��0���� aPI���� �������Ѕ���bt�> ����K�F�$��zk����/*�ɹ���������!�]���C~��w*&��榦�V��wtz5}�
f��:a�._�e�	~��d|Do��
��|���¨�0����pM�&
�j�:����F�&]Z;ŝ)7'�&�&m^o[�-�=�o�>��j21omn�JKc�ϳrSbEq�,X�����0Ս��K��9���s�!���:����Ƒ��sR��$K ``t����ؚ��ը�\��)yCϊB��k}i)U55J��:]��&*�,&�(,H
�x7���[�q\���3>�D��y6����JJ8G�C?h�GT�6�
C8�;�e�������c��(�˯��� ��׻.�\xKX�	T�\��`Un��\������;�@�8*�)7֠,i���,��zAy}���#;��H&�T����8LA,4QW��#�z���g���?$2(k���:���[�J&���b �t�޾6�L��6�/M�Tl��M��Y�������d��(v�Ɖ��/�Mo!�M͹�^t��Ң �
uW��W���܄�ٚ���uT�S`	��Eb.a�Ҭ��@���V��ge�*����G����	S1�_b��~,�щ��y�˹f%�����\j�(�5�%��t��DIxLB��5Q2*
�Q�uJ���f�i+@\�٨-UƦ����+�s��Qt��:���X��a�2�'0�'�k��^[4oA�n�`'��9�[���p����gڧ����1F3��iRw���Vn������2 ��.-Hzb�5s�n�%�r�V�i;��2g��il�ޔ�5���y!���*s!�dKm���r0���.َw��k�ր��������Õ* �ӎ��k�ۑX�:Ҷ"�{5�"��t�9�^�	|�$��ᱹ�����~{�D&>��^�~�ɖ�Vf�n�O,�3�$���M��6y�#�ڇW�F�dݭ�}�Υ�����u����c����26�cUx�<�c���rjm���q��d�\]���9�&��߳���v.�[+S�&�|���,7�-$���c7�A�qV�� �ݷ�$��Ǭ�F��ăhO��������Ȝ%��/���o��n�E�n�0e�&A���2�6&)hRf�(m�k#i,_>����ho�j�:�Q>K�9.9[4��zȚ��7�`)GZr�Cm>��wX�얣��y=�.��m��ު74��x�e,5�b�_�S��K��ưQ����]�X��y�7과*��=P%,}r#�=����G��:��m}��@�=�yvo�]���xOV(|[�3��	1ٚyjYk
Y����ؑdyrr��5�|ݧ�,�<,��;��������Iqڻv�:ޏ�,�	É_����n�d�]�t�C��eΰJ784����o��"��2]�����(��rI��/e^ɮ�����^9[ţ�U;��\���O�}�ޒd�� ���t`9���\)�#���y�ݩӭbu���X���*E�
��|�����tlL�h�q�Ī�+!�F.��ꄻ9+�@�a_�&����y���[	Ig�x��	��I��WO�z���}�-������a��	�J�z�u���	�:�CYh����0�#�f����@�����C �������|�sS)A|�	�v�z�2��Ĳ����N�%��z-��v��zm��֔���Nu����f��#*4�����ΐ��%��0���	IiiO.H�۴v6��"мUG1fqhh�$��i�Ёwx����z϶-�"�c����ߚl��̓ɋRHEd��������{k� Wp�q�tZ�?����I�p�k?�	 1�E{o�`@���v[EfQݞ8M&>^�>�C�ZxQ��/�xL��,��CSj=��c�"WO�;:��'�k�P7��r��X�v�>�*���W&?�m����K����֯�[�uv�uu��Q��9�y��p��.e���]]���$m��`�OD�O��(�5�؛����a�#�g砬���;��f͟L�:���V���{�/���K����#A�#D�m9\P-�'~�;��SD�� WN�Ǹ�u+��/�z��`��]x�"�Ӗv>� q�^�aal�"f��SE�a�t�3�Ќ���.9����j���+�VG�Ֆ�B1'�Y�G��ɀ�3��7m'��,㝄��ܖ��}�Y;a����N����?��.��j�i����mB&_�j�rO=�-�	�2ߣz�������2	V���c�l�"{4����Y{vL��Oμ�ﴪ���v:�	�~��l�Q?�nM�����S����IU��z>�|k��>�)6�[��_���E;��=�
��o<�^݆�Y�i{��Q��N�.�����=P\�P�|��Ml���	9Ki��>�W��_T��;�9�;R����d�>m*�nk��0��v�)7{MR��V2�����[������2��>q6'aݦ^҃��3�"�79C?���Z�y�;_�a '��j%��FV+���ߓ��/l�j�v�s��#~;�ڨzɂ\�ŒB�hi-����Ƽ~Y�EH����z�X�b!��S7h���K��tG�������n?BUT��W��0�5	��i��Q�0ј�R����
���_���Z��.Á^!z�L���k����LE��e��h��s�t��6챩��ِͣzݩ��ΙQb�(۴� ���:z�1%�!�N+��G�i W}��D5/^{�0��e<�p���^�ܽn��Oӹl�����o\�1�/� e����x�F%-n+<(�ǋ�n�6��O����3sJ\H-�73�e��:�R�:�+c�ԟ�	�a:�+�r�K $HF�ZU.�J�fJ�{���N0%�9�8(�4�%S�(��l��l��T����]$_�cٺAد���&P5 ո��M�6�8Y�?U���%d�2�o�(	�& ����#Al�*�\��3�y��=)�mff�D�>��P��;�%#"�.K�B�w�.fWR?> �J�IW4«�2��6>���ǌ�X%�ܲ7:�n�E�%������ g��;!��CI�b�6�d���1#̠�f���ǝ��L��Q��� i��i���[
�m�#����f�s�S��/�(j�w6����G,�G8%�{�3���={�u�j%W��z��{n�t���&��o$�����z��Zs�j����v�HArM	��Dj�)��-'C~�$J���멞QZ�qZ����W�H�/!����!�J�\��8�ʟ�6mw�	%U_�{B����q �h̜i��k���oI�x����	e<ހ����'榍���F|:BՁۨ�ib?�0�$Bf��t[z+��D�sd	&Q��������#��M������������T���2=�H˄������&�u@i�����q��}-'�z��\��#x���z�S@�E&b��1�$�WwSA�0�_��������t�?�g(h�O�Rnj4�6A��y�Ժ�,Nyu�g	���OY��=I&����B���6�&�w�}po&�;σ���dL�%F2���� 1�����������/�7[�ek}�a؜�l6Meو0/���KJ�*�u-��bO��<)fI+�/֎Y�$0�՞"n9�\�W�*��b`�d.��˘� ��CT#9�� ���������$eTu怜���0(Jp�m��v����*M?�z�9GAY�Ǎ4�ZiblN/�Ō\_u��l{W�Dͪ���1�,S�u���۷���-���ߣ$V ��Cǘ��@���ǲ�v�����E5����J��{�=Y[��\��Դ�2t����M��  ���R
H�� �+�\�D���i�f)�qH/Y"/r��٘^��qX��0e^�_�?��ǚ�s���ٛ3��Nlm��B6y�l͟�6{������G�>H����k��'�3�[xV�"�iֲ)��l*&���6��/n7͜7�~�_n����t`�U�"'����ѫ��Q~��v-LGѳl��/?B2�<z.�>��l*�a�.�cD�,�t�w
]�}��K/�ϑ��c~���aƲ#��{���5�Y���H�TF��b滳�λjo���lo�'\[A����v�[�h�7|7�W���M����ch(�ڏ����h|��\H�ϣl�)iK��*q�"M�L���b�3��v�Q<��X B�Ϫ���C�qZF�U��A�G~��&���^'�;�#c�-���2xsu�58'~�/��q�M�Rm����q��ܤ����o��iw��F�Ig����Sl�C��öD�@Hc��h��$�I�Npz�k֧5i��}ysO��Mh��"� 2��=^��+n����?'�|�,�S>J�<p.L�e���eI�hB}�vZ��ojZ������F���Q���tn�Q��%|7u���~��N���?�%~o��E�<( [dA�rsǺ4�&�+�&g�&P�L�;9P��P`��QW�PJ���ù2�%SCN
0ة�ɦ曍�3�~|�;����ao!P0�T7IK`�}i��(�_w7��qRkp�P2Q�HIKm�	��6� 2��ǆ��|h�[�IOoV%�b��+��q���&�o�AE��v]=;��jD�'OK�O�u���r�ɲ�F��;_��n���Y��~��y�O��|���̨�}t��V�̋4�o����%�F�e�c;���
�2'��*�R����������!��'-�s<땣�3\"h�/��H^ݎ�u�3~�E:}�u_�W��p/����2TK����$�#��~c﵏�t�2]�'g^�����ʹ;S��V`��T���/�Vכښ��N�j�+Nt�L8lDe����?������-+*�ӜS����?��� �U�t{Yw�<�ޛ�g'!�-��r�(W=ۿI�Oޡ�d����&=�e�]r.ٞ|�1��,&C@)��������K�	+^OI'mI�4
1ɏPZ���2�˿�`+>����7�5����9G���R���'�g���<"�~JVT�6��ВȿЀ	�s�&"#�D�|�7��^�K;��B�`����K�mlD�^�"��ښ��~�9K��^62>���\d���!X�)山�S��*'�J6�=B�?%�'��۶�ܐTL6����������9f�3W����ZGŸf{'+=a����C$?��A@�����$'7[JpT��Xj���Uzx�������Z��\��x^�ܴDo���>�Yj*�K��4��X=�cZ�)I��#��<)LL,2��2�k�:/f/�}<{C�DD L%����!�M����dy��[t��6g�@ya�}86�m��=ꚟJ��N;��2�䓱Uٶ��sQ�{�N�<���MX�<(���Ƌk�=����H*�����5�=Ԍl���U$˥�oJ���@#��"�Hp�^��B�-�]���4'�J���y������~�
 BlV��Eۨ��}g�4O�79A���wQZ��udi�&��)f�J�Z��	ȣT�7^p=xt����V\d�8n!���Q�e{�d/M���/z#wD�D��� ��k�}h����Tꨢ*�ߋ�嚇Y�u���U�B�"1f��sn��~��^-m{n�e�s%k����lX�`t��W�(_^�_���Euzd}0G6*��8���g��~�[�Ut1�d�G����׫;�J���xID�{po�W���� �Z�.)uZ�����Ӹ��@��L�sU}z�{�IÕ�Ȇɜ�?�e�΍)���(��MBX"^��o��-�L�|�d���� ,¡��9�ȶ�@����a���&Cͦ�*�y�M
>I�v�o���u.�Y�����iK9�;onzӸ���f���aS��/�Dl�t`]Օ��)�~ae"�,c�xp�GO>�7�P��/�ߔ/�H�E(�z�܊�i�^��)�Ѹ��`:Zs�U�̤嚎�QqN�މ�>��Zj�1!��h|�=�#IK�J����Ka����stJ��69(O��
���b��[?��@�<E�YqWl���H��x%�Am��z�j��};Z���#u܉�T}����{5�!��=S�|���*}mw{=�&�����]uI�\1ضu�C2�g��^ ���n��E��.�q#%2�ZeY�9�;�=��_m�����]���ߌB�`jx�m�6���������9�vj��D���{CZkGMd�L��_{��r��j�[���C�Č�Cr9���v�$P��hO(��@w_�"��C��[�cg����3��ZM8���AT��M�c�z\�����B�w�5�.e%}�43f�����^ŝ�C<��5~��ή;$ޅ&�d��oo�|��7bi��R�U����U.�S���i�
6�}ok˙��K��s�컫3ʘ�,�ǖl�6�]���V�۪dd�!��l����_!�NO��xN���,f|]�=*�Q{�h~��.O�`D���A��lqUlUv�I���������v\�&6:��N	�w��P,���
4��e��rWn�sp���z�<7Xw�Mm��~������|���I
0ac�e-z��]PzW��cO*�+*���n4���љyo2Tɛ����#%���SX�cS��[h5���y��3S�l���ؽ4�k��w�ℼn�Yio���=i*�	s���ƲÃ�^����e]_��,���0��̿a��9�q1��9�����mk_�$���h�b��
�E���!�R~�:5�P���QM�s�|��'b�L7�����3h�"a�8���{nLD�Y�q�)~�NOI��y�TS5�{;�8����^�'(M���ҷ�(
d�Z����߳=���h[U)���d��;��5Ѿ$�tEoE�c�8)����
���a0p=\~��}h~	�IUY�2¨�(R�T��;����]�k��;cc��-�wӣR�*jH/딍�h�����~�s\��3D^�eu^-��HjZДX��q鐓�-�J
.L����G�s��;;��3��f�^X������.A9���|��F�]d�-d^p�����β���Xϑ%5��A��1��I�Ax�S-њ��s��=B��e�>._p�{f��I(�	� ��%9ʞ�����b�|�H��v�sM�<��`?�_qS��G�z��}�>��L�a�^�'r2$�i�+�?L�v���f�g��q9�E%d�1�͎�O9�����Nc�G
DC�q !AMY��m�D�����M�W�8_w����L�M������X����������%)M\���xWE}��BԦ�1ni���'���ײ���yu~R����lf��!�K�� {K:���Ӈ��Κh�䅯M<Z�[&�U����ky |����Oݺ*_�n�v�O�M��<`~�3����w�4��.אO��*'�� �Vp?f$?������%� Ԝ�2��+t�|�2-���Z
Ld<���l���L���e��P��eb��Y*_�ӾJ�H}!��K�FKf�/aao[3�5���ݒ�B�|�{
��[<����-g��T��F�j�m������4��,	�3m�ӗ�m0�hr�27�	 +�WPw:9ݫ��KNgk˹j5Κ~���ɡ	��ٱ�#t$qx��E���0�q��Eʤ�����5�J�f����q%���V��g<��:�O����+�Z
������hm�\�.�,:�I�`�<^i�7�f���!gF��8^��N�#R�qj�����1kEf�a��(� ��?�c�~��I�_V[%���w=������Ã6�|�O��㵦�^)�r��x.�W"�랦�i�D"_.���ؓ �,�>y�������F ﻐ����e��Y�F��A��aM���"��Za����1%$f/��� ��#{ӊS��?0���&/`En��½{�C��o��~;8|k�u���7l�(���&B�֒���� �7"��*�r63*�n��M<��S'z���1���`v��-1��b�gq��R_��T�u��}4�&�7h烺���&V�o�۟`~�V�s?�ͪ� g����m��?o�ĵB�� m�T�*T��>�1�[^�T��vH˲�!nr�X���3�f���E���a��K��5ze�������Z_.��Ǚ�8�X���y��$)K0�|�]���m�[܏��]H��ƴ���$������ y����>��?��+ ��'	�������ҷ�ŵ���r�&ś*�T�ψ�t�9i���>\����+�$�����*�E}B\�� ~�@��]EĒ��bg����I�A���p`r��C)	�fnt���@�K�֑{��{�#�L=s&Soo�]�����WYq�\;�cG>�5��뿉W��Zh�M�B�tʎ�F���A�߼��i�B=E�ls��[��tל����t�E{�H	�OZ�}؇6�th�2�E�{�va�<o�)jA������OI��L�,��n+��Lԇ.]\��O�_���:��?J��x�m�-�yê-����{��L�,5L�K��/�1A9���k��+�ط,6�ƛ���4+j\[MF��ʔ3#��onșO�����h��X#��?g���$�ـTq��̯�\Z�~��W����U�,sEbS;�Sܤy�A��ؗ%S�}��Pu� i�)�E';<���T�ӋmœF/3)\V)t��a�F��M��E�I���%����pڂ�5Gl��L���,2Gp����3��M�]�>^1kA�ɫ�*7g��#Ris��qo�*_�� �=�4��p�I�p�_��hL��ń�+��I�o�Է�M}a��Q#�͟|;�jw�B��WwWSٞd@Ö�ǁ��ܢ�����.�[��Ko�$��Ŧ�	�	h����F��t�ms���L/|��C]"Z�0x��$�
�Ϊ$�Ҭ��)v���A�R�0Z�
J����հ&?R���sip>�߿�{r�K�;4 ��,��H�#}�s`��Zd�#������-���$Wo.�Ԟ����~��I�_��c2��3P&���}n�����<0A�%J�{ٷ�,�<݉�q��J>�Y�X����5ec~1�Pg~��C^���A�Ḑ�B���� =Evp/;]���^r�z�ꃡ�H
x҉����M�S�����r���#��}¡��Ks���a�#�3����y4Z�����d ����}-8� ��
�mm���������4r�K��X�+x=�L:��萬ߗ��}����-�L���)�Id�w6E�6�!v�ٜ� ΅�]�{�[�����;�w{kv�/?L� n0��	N9����������B%%��/7��|� ��|�+C �e���{B{��*�M*с
L�4�N����V�w�_�����X&�>x�QP� :]*T�Z�i)�)^]��9��׭�m���]@��ֲ�����2vL�j����B�n7w>y�-v�ڿѫb#�Oo,�ɣ�Թ=X��1K;��=g�GJ"���qBŲ��d礟������������jOk%�}8t!F�Ƣ�&�A�K�6w]oK�[�	k�X�r,&�+7�ԧ43Οb�}ep�����:���l�o�?������9�����e���Id;#){���v�.�3���˨/{��ic����H�T�q�c��$����	�R��溻	��-vM�Z�:_�Gxd�\9l�',��*��:��/E	��k7L����t�����4p1po�o��>[P{a
�3W+[-���%�x��]M_Y���pX��##ڦ��{E~Á�r�u �'��7_���O��n֔���zF,'����X�=\B&N� �4c�΍���A�I{��sS�d9ֲ�-�S��M\Z(�2�Df	��W<������%���76r�8��-�	����G�`�r�
�3�;�N{�hj�=�)\�n]� �pW��<+�
ƍ�5z�V�U��%�,�P���R�����s�7O�X ��b���H��2+ =8o��&@#�X20�������Ǒ1 ��B�S�g��������W�ǻ�	({%�xT��Ls��i�O���� �D�[]	���i���h_e1⌝�_Ў�Ȥ^�s���<�z�+���z�s�3z\Ae��0�����T_(�+�����.3��u����i�����w�L<�J���#l�<�L���)�*'�@&o>#�)w������VI������=�X�#�L�A<��L�n�"�N],�FٲrĤ�u��[u��ٝG�Zׯ])��,����È����5_}	�L�j�Vz���⹢�Cë�K�}�@��&���1,��� �L�.�ڻ�i��1[j�7~��x�4NFv�7^5�]H���7����q���
&n���/�u��  =�7��t?��%�?B@h�l�5�a���/�7�U&�<>É#�c����
�ښ��٩)&�E[�&����)%�c-}��7!#��w����;T�r�aXex�P�q|�ӇT:�iJ�y�K]��:Mژ��+����fm�8ȹ�_,����N�B	|6�dP�d �8��[�����bG}��x��z΄"�{�w�:)���l��/fcMo�Y�Mu�c$���Cecf3�=�iM4�?����������|/�%�4F\Y�:!5
����B�E0�P�^����U���Cv�)�%�|�ת����9]6�DFinP�YV�o}�
7�4F�7lCv��!��|c�E�CVb�#%�-bB��h��|R:�.r��3�׳j��Ջ�����{i\]J�]]�15��3�O�Ϲtp�+*aJ(n�D�v�#r[>�
�vF����	�Ùʑ+ƻ��EW�
B/�����!���9rUB0�ӈ�������p�C�4L#�s��g�>ĳ{�	#xi��g��P��]{J�,Ҟ�&�G#�5�\uh��C� -��V��I�y]���:ݷu}"18u�)���ο�]���١X���m�aKM�څ�p�S�3K!�16+'��"}p}mV1�ł;�����?b
�f����~��c���@��?;�k?x�z\���J��bf���Kyy�,�k@.+���}��l�3�&�r�����D�X�3�z��������b@��e2� �!��w�o�V�}J� 5�����3�\F�he\�a�o%��=�.�w����87���a(���d�db����fޑ���$�4��GC���H����%�:����jLC�K������V0e�us*�5�5st����EX��
�_���� BwP��F]�csZ9�Ra�9�7w����_Y
�Ps��LޱJ�x��3����S��܈�X
��R��9תVבO���;�h��]d�7�����p�}{����g�(�>�T�+f#���,�4�|M�U#���G��u�p�rvg&�2�����r��;Uݚ�S��6��V8���\!\�`�ԶC�V�/=y	Cu�e��a�d�J\��r����i����k�����mRXR`����\�^�q�����k� w�PL��F����M^]Y;Y�Y�����gD09��~ ?�N�g�&*�@p�kb���?�Ƨ�����{˪�-���3�]���^ �'I��Qd�
R��j,���e>M�#1�6/��x����Wy;�&)��0T��ITyV#dX��
!;e�S���ٟ�W�������8|>f\>^���z�m�9z�fOY;	 +S����̵��h�37K������oV��_�wk?��
*&�*��Z!��.��l*Ѽ]��
�_	��f��jD��.��/�rƽp	�"�#k2iQ�[%L��� ��Oa=�I�3��P!M»�]u2�$�|P�6=�I��ɾb(����Rn��q݊��q��!�\!]������z��fh1�[�s��ښ���%��[rQ=S(w���5�!���)+/K������fO�ͽ@�z!��eL���"/�'�	ٜ�*Dp��څ ��w�e��K7o�-֮�*�ci7K?>IG=�7E��S1V�n)���T�'XOwI=��ڇ����'�X�yy�x��ݷK�Dl|��:�	)#ݼ�7�2���i)g�Ip�z~[������ ����) i�D�[��H&�i3��z 9"s<�9�'�DŢ�$�Ns4��B $�"|'���n��?Y�9ag�V���ô�������:``��Ǚ���l=������b��>i���g�������TE4)2� ����6H�z����tE̚������#�y~>�]��vW�0!�K�����\lbO�P�WU02��VY������L����Z�%��$�ȥ��ԙ�a���=.�k.#l�2����P���:~������9`V� ���'ܗ+�ǭ=�[��Z��\��1&��^.�?�l����S94/Y� .���r��W�b��+5S]X訵c*�t��o��ɭJ����W�M�Eި7}�Ɉ���G�aRv��0�o���p3P]��gv��oK����ͼ�d��|����WdI��k	e�����An��c�5�A�V���1�x���䄅�P�Qso�mlp֊|��7��_IW��t��Ƈ��?x-���Ր5�QjUGo
�GLg_��2���ۈP\���k�e�9��m�0�����ɕ%��^@nyDj���j���C5VX�@'�E�Vu#Ḱ-0S����>�P���A��y�P+��.�h��*�����C����x���,��V�_��;Ӓ=�\j�"��#���6��V�����)���5�y���l@�~�BR���?c�:VƂ%*��y�Mw���A��X�`��f9���<a�2����O>! �o:~w�P�)�����s"~�5H�&��/�QaH�8CEOs0J�������1Z����ȇ�Â8�;��:Bm=W����C����V
����T���}˲���]R�`.]�7�¥ϭ﷚U�
�N|u&}S����"ڻ�X���ifY�@�32=_`$آ��Z����5ˈA�8Du5���t�ߟ�~��T��fc�A!�'&?G[�:@��4��a��BE�Xvͻ<��tQ~��(M����|^x{������.�*Y �z�v͢���s��kC�F؁�e0���h0|p�����\Y�w��� �buv�BaE�Z>��O����2���m�-��L���R+dKk��H䁏$�f_�Dy�϶� ��ؑ?2�h"��{wi�[pT<#j�������F{H=�$���w�>�#AQ�F�
��ME­���8 (4Tt1��g�Yߨ����l�A��':�Մ��e��)/U�L�\lʱ�7_�"05y�~m�]έ�t����o��u��&�)�R�����	^���m��p&�������Kٛ�&����wb\���;�f��>�hm_p�M�Y�$���R��ɘ`2$���������?�����cD�<�g1���\Sc?�(:v�k��v�[�k����f�b�!l�� 0�ΧwUEz�Sx1<�%�T�p]�<%���W{I5}N.���@�@|����'h8����Ä&�1�O1�]r�q�o���hl+?�^c拐T���A��A����<�02�Tv�����sn%8U�q�l�k�ll��9��2N��}����O�0�çE*#zM�0Q6��N��/�v����rx�Jr����p8;���pM��̀��@lzs�U��i�����0���:ڋe�p�{�-�������:�ܳ��{�*���^3���F��F�%��F�l��s�<���t��m�g��^۟F��vAi3�R �6���a �}�wf�]�aK�e)�rZ��8�����M���^Yb����+2��✴ ��w�(;˺�z'��Xd$k��#��;��(xߣ�ϟ�ܕ<͝���9,�����4�FUg�T��wxc�"��K"����������h%�����,�E������ë�@����'q��{*�Tv-�ǂ���9����r�24I���N��t��Aov���N�V"�p�j�py���K$�ӃbPE_=����ŉ�e����u���ޖ�[�0����NA�1^Cn(�J��x��ih�ߐ� 8pl���=53�*aM)@O�0�'��q�ɾ�F���`0��dR���K>�k[2&?� �
���1~�\պ�:���; �t����V��W6n*$�})�{��(<�V�y�>�F��w�\lg���r84��X�~C�㚭��+g񕿦HJ��4�B�ڐ��|=E �&�P�<X���uh<�Z2���9aы{dا�:�3dp�f�R���`��H�9��[r��mpH�e������Ԗ���۬|�"�����f2b�D7g	��3&�%��D�Q�V����y����Qe�4���R3�<�jH����"� W���!�s�,��S���F0�}��T����X�>��=��~8��A�yy�cA/���q��2-�����X�H,�}���D�%?��dd����_�P�\�h���.��B-�"�I�	�u�����՟@^��Ҥ�'	>')�҂|���*s�#���3�j�����X��š�X]�����!=�6���W�,|l�D��������^#uS�.������yM�sq�o�Ϲ���X"�1 ب\��vj�ݽQ ���~bC�Ң��0�� p�{�e��tª���ǐe9z�m����(��s�:G>b2j�7U�#��z%՟��8<�I�� ?g�-�p��%�-�a�-dN��Hn�K<�i���?T�����e�����>8tz&�s��̙r~|Q F-}�pu����N
UΈ��,���Ƥ���`��s�(.��-'m�nHl�go�(c
h�/��ŨL�(�i�2��/ر��\18BU�p�dfn(�(B����o���Í�#���,�&җ�%\�Z�."N�[�s�%�ꊼӶ(�&�?V�e�[J���n!j�k��4P�=\k�g��d�
�+��d� ���g�c��� ��T1AI^{1XO�E����3�'�G��g~;	�u��m��y����&���R��� M��P{��]YnOB�:zcsd��V>tգ�?7D�e�vi��	j퀡��'>�0\&C�QQ�Ah��A���Z��#��2��t\��̀ S�t��$�L���0I�1���)�H��|�"AM�z;�	�v���f��g�*��%#�աr��4DX^�J��>�M�����O"��T��5D��w#<��#2F�|v��9nw�g��6g��G�,�0���������:�j��7�����=\p��~��C���+B�l�yP)R�Z�PS�=
�_�{kl��#Ž�s@OξÊ�A�L�|�#%xT%`���n3n!���������n�B̍h���$Y&f�RU�꡶8$0��OEG�Z�
H�+;�����o�Fm�
w��a���-` ��i�"?"�{Z���um�c{�Fu���<���$���`0�zՉ�C��[��E�~��_�Js�V�NC5��Lhã(��\����>��Ny�.�b��i�V�lڃS4I^��<��5�����I8VV�������̸�Gr���3�?�l�@��|%��E`s=�w��1��u[HF*�����^K4�*��H�[-�E�F�;T,/�f���e����i�F��dSޮ�'�&Z;۸0���	�*<qy���_7y}]Lz���I�o������K�:B�����e����x��YI2��jU����-1-�������\�(�"<��Qꬢ/C��&=���upd�Q�G�\'�&96Qw��f�Hm�a?F��0=���e2�y��	�F�|�,p��UD�r��D�ޛ�j�� ��;|U�fJ��)��/Zђ�X����Qu"���]���`ޚr60,N�i1�7��p��<�NQ8�:�����S>.���� t, 66y����P�Ϳ��D�>�'�|�Ҍ�X�A����ķ���AW7SV����]��vv�h�N�� v��/Ś��o$p�~�U����&�PӚh�$�X�W����y���"E3�n�d;rL��
6�v��7��ə�����T��:[sW�	n�ݶ���֠ý�L�-Nڂڝ=��H���)�$
��V��3k���0��gv	g�1�"�m 920��I��2C�DX��j�ɐ�Υ5����7�~�.FkW�r�A)�R'��#�<&y�7-�'��J�y �[� r�#��e+}Js�f�$��GK�x��{h�1Y�y���A�Jmvڧ���l�(�(
�'k`VCjF^�]�}���fceۿ:�S��nq�^�>��HӦ$ߛ11����5�UF�g�3�م\���fo���%V�?��ƬOb���}9P�ǿ�њ�ۚ�N{�)�-��,y#F��=e�����/s:<����س��g�;|rI�Jg�a\�@�݃˅ܶM��P����!�����@P�~�d�VK�ͧ*�y�yg�|���e�ŴG�d�-�v�lJ,.�ri���yEhv	JR3��EnA��:�K@l٣�#R��������+#suo9��Lu�)��"_g���opw�O1�S�ˡ�T��U���!�uZA�d9ٯW��=Dwh�������#O3�]�.щ	�ږ��Je�S*��+kN1|}߂yz�d�~�Ϲ6i�D{Tf�FB�z��m�`*��d}�������9<���W��L�<����h)y���-��9j��r��Ri��=�=��cm��3�xj�䴎�c�Z�76��|rKP��h\:��y�h�V��#�j��=i�1����!��̀��z����R��.����s7qؗ1��n zͱA�1V������/Ljk�#��:v��4� ͆��p� �
�Δs43-l�o���.���N>Xe^��ʂ��"n��az��(�w~���U1���B_��Ó �<ArP�����_�_�s��4X[Sjkes����O���SZ�**�j��<;��2rkP�b�5P��������^�@X�D,��Z���tU�v;��'�1�钶�OV�kF�� �a:"	6qU�ʝn������Q���e;�~��	�����J�2����,'w�@��������캊�/{!v�g�*L0$�fW�Q����У�o/��Xdfn��4�qI;Thօ��*�]L�x�����sM�#�MƘt}�	*��s9�v�-��,�u�,<y���H��*0�Z&�FeL���62��̚Tp2���sW���� ��R)Au��:�4&��g���@V�2�o�=a��k [YjF����2&ad����-w �c �SPҍ�Ǆ��fF�5�/[��*������+G�����L��p���p<��� �#&o��軕>P������Umi�_.c�,H֧w�=���s���d��'�ҭbV� �@����;zI�?�P_ćwD�!ɲ5����_�K�OW���V;YR}Zq��2�	_��,}Pֵ*���n��x��t������\܂�o����^����賠�k��ڄ�"�HN� �I�{X)1�>�|2��C����@�a&S�t�S����Јq/G�nQ
��]`�A�.���9W&����+�]dR�2���[�>�E|�T�i�����7CwVU�n�r� .S+���:����_?�n�g
qG<^?�(Fv�3 �I�˽�»���	Q�
�UH���l.A�њ""Xx����%���
l��}	�d�&��yHED�i�C���d�<-�c�&�#ީ8{��0� i�u�X>��"���վ�+�3��s�yo�~��#�cv�nBW����U�sn�R�_�^��9f�F[2>��������+C1�W��G}9�@:d�'��o�E�A������[���&sbtT
0���Ѷ��9Bw����?����RF �O�S�6j&��RmpG��wtt��4nw����F+r���c��:TN���i���`�PY<��r���T�:���������µx�d8W(��x]�@�������'�����
	ߍ ��ƶ��%u�5~��ŤKP�o)ʄS��dl��#�&T}OE�����u�� 4E�k[f#a����������-T"���L�e�n�ԭ�nK���~���5V���p��[�/H"\n�XJnŰ#���'�W,ȟ�ٱ,�@0���ދ��3ǁ�D�s�-�6�K8ձ��]����c��2�	�1ԦV�ť��*��6)�Qr�w]���o[�d���py\[U��9�ȃR�_����^�u���L���*uR2?F� :[�R<�G�JSD�݀�B⓹M4�TT�gͯQ����t��!��e�G≰;����$��b'��a�1����j���{����}����!S;<�ԧT��AHB����I��S��w��\��z#��wЀ��F�r�
`��Y�+�D��k��J	f�/#�!/�������T&���㸤��@ӿ;wk�h�!����k����?Ҧ@���گ��7^L{Ry4>e��k���꽆�C��E��2L��~�8��������I�M�v�e�xˆ[��W����_�$��$
jV��I��؃e��6���R�Em�u<�)3��v1�^c��Z�W��p?�/��ao-���g���Q�#��E����c��e&0��a�����_���0�x����k�g6�x���N4�Q�D���좚�����6ϑ�!���Z>	�K��T�泜�C���`k���Xx�Y��rS�jy�Y���������l�=��
�?��bZt! 0������z�)}?��!�����#v6�it�PQ��Pm;a�����Ju��ȶ��/�h�t�mM��s�0㐷�s#Zoez�*�A�%�I�	����Q�\|M�ӢE}�K�<XQ��.x�VP��M���w�F�b*H�;���\_AG�-�6��g@)R�3���&�u��u�R��� /]_x�"<w��9�p/�<�%0�9x���u�L���j�����@��a�(|篅rK��.����[//�onP����o��Ce܋W��G�}KV�l��q]n��/V�o���l.�l��D�Π�he�������*K{:���*��$
xwR�2��sw/�&�/�� F��EԾ��|��'�(�I��S^з<tZ��5_N`����%eh�N
��l�>��6v�w� e��� ��U)E��L��)0.n��({�3y��U1����6B�u�˩�<T2�8�����maE.�0Դ�M�	a5��\RAh�
r��PG,9�j3���� �A�S"9�y�T��ZEz�Ś�.�@��.���J-I���w����*��~��d�Ri��Ns:W�������`�/����:��6b��4v`���q��"2��W#�¨B��O�yV�:t#!]��3���7�n�V /���yO���	�i�C�oXD�PB����΢������ͻ��G��U��*��9 ךi�O��?d�P"5�55��ܜ٣6��>�Y��T��s�U�1:�C�UX[l�טO���F�d#�w!��A��q�q����,��cXvI�j)�w�
�ث��I*<�������W�x�i��z�w��R(�:/����$�����k�0Z�L��o�fN�HF�%��H�hB1���6Xj�Q 5����I����x%i٘���L
l�h(e�������-��$6F+��T����9����$:�Ƒ񳯪���Z5��޶M�l0�~U]�Sz�Y�r3�O�Jqo���J�.Ľ�Р@��>(����p�'�Qu�j�����C+�8/�l���*pῳ��Ǒ3,����}���OL]ˊ��c�h-fz����a�qϣ�_�Q�����
,8[�z�?����v]����F�{�\P���p��Ng�h{7_$�r/�Gs=���(�E�:	w޵N��E��x����;=JoY�F�%$ȿc�rI+%#�W�Ɍ��H`�V_� w��qY[)���X@o�����.:��#.��+:XO��z�߅c ̈́*�"��L������d]%.^�>��z'@�̈́�*v�����wa�I��q�TG?z��tr�S�h0`;�[���]�\�+���U�<_���㎕}�.ƣ�~!]��S�%��9��˳C̦:��6߅=.���[Q7��Q۫�g2T��	?!�Kӭ���Y��s]C�q3�}��!��@�i`沵�W�q����8\�e_|���$W9�=�%�ݥ%��m�+�)��8����.����`�7��O��n��Eo�'��P���麱8��c=R^ �1�|��$��]�1� �8/���Ӷ��#Z#*--N&�!x��6����1U;;k���D7")�F\)֐��s������"�ꂴ� �����Z;s�w�bn�9�F'c��zo�YݩuѱN���N9>\#t��Й���S
3����;5�4j�9a~�Cy���P=j��p�<�#r�L���<!�I��D�   �
�f��A�R��Q*�	�E�8�B�ʰ�R�E�I� �`	t��Q.0$���&����G@�G�q9�ù=;����>h�9�O�~�w9�p�������	���}�.zمB:c��@� ����wY(�W�^4c��b�w)�p�5)�&}*�<��X��A:BN)"�8� 
�+���Zh��IH�p���0e]�,z���G���FÖ�<T!�dg�Y�k`��!{�g��8S�#9��SB*��H���v��Π�݌�x�������Ö��w
�����P�h�x �+��*����_��6�|]�j�k�/�}����R������r=l��9]��w�g4��2�b��j��{�_����qyu�ׁb�z�*���������p3�u����m�-�h�0��Eg��`W!g'h�a*���^l,|�\�\�Dp87�Tz)��@���0�&�v��C��"�@�T_��_c�b�,��Τ4)-�S�z~�X����k�r]�
Re��Ku@p�"�<�^�������+u�YT����>?J�'��H*�FS�3�|i���m�`]]����T�g�֭s,��<6�!Y��KBZtm�u��~u�\�i��ƽ��]u���9s�.3ܥFoJT��tu���3�Ϟ+_Jd���/z�*�(@A��(�^0��d��á}��[�z6�f�uYĀ�+�f3o����7������9��L�LIK=p~#���<z��W���dz�	�֩4U�פ�N��s֜�*�$����W�yFk�tb�����>u���|���/d��o�"���$
��7L�	���[붶�$�������#���:�������Vb���`����e%�U���h=;����zX���!����p� ��D�-^;��P�	5uo��q]F����j_�_}�~�O�܈t*0OXn�q�=/f;��B�sr=ny��+������S�~<���P��%�YM5��P,�&ab"��\��-3${c����D�hhw˝`k��ucN9	�ij�Fo޳و�~�����~�hl���$����?��,?���z��@�Ec#���<�i�ٻ��j�F�GO3�$�I�i(R���O�S��.� s8^ZU��i�hN8dI��C�Q�J����G�(Tj�?И|�Lȸ��6nR��\%ɸ!�ҟwS�81*����ȣ?V��.�����yt)�A�Z�2�"{�߇�x�h�/A�o�/���qNA��s�]�JO�=:�uA���w�m
�_��O��wws���'<�YE,��f�X_T	֩���>�ф�@|�[�5��&�ժz���o�y���qJ@� ��kґ-#n���:��(y ���ED���}��&��[���/�.�G(�SW5���,�+U;�rY2�������(�φǅ�C1�3�@#
��O�[:�;<�T"	!�a����^�������p�� b6��rͩ�i���9 �3v���ny��F�򎫼r��o��4�|L�e��Y~�m`{�sz�� ���=�
�8q��Sj��x���p&��\Z�t��/~�O��l�}HL C�Mh�#)�$Ԯ։h7I����{�Ū�M����/ݛR���y��"A�gj�S�E1.����	>�%���y��=�ii��b�����uE��CVU�%�İ�A�G�_E%�*��#h%� �]H�*H<��ϲ�)�3 q���9'��7Ra�ddړK�Hp��~�	0O�A��J�c�&ཛ�������=_���u읂�4`�E;��*�����yٛ��#썔�D�q`�dM�b�4D��h"��f.�S���*?�d
j|Cf��5�FT�6lD����2z����Fj5\r#�mn�e�����77��d�(���	�� ���<�0g1�k��G�X5#y�Ĺt�ω� �;���.D0I��`�����jOn�����-�2�r���)ebw�7ȯ@�d��ׄ� 6$~L��r�t-��U����1�OᰖM9�&?��i��i2f-�"=V����sP����H�;.|�W�a�6�D�gR�JT?_�Lh�資�>8q���E�>|�}�� [�	�����IS�ȓ���T���;"^�&M��]t��f�Ģ��>m`�8t����0ȥ��Ɨ-�T_�M���:�b��=��Gfڿ�"��6a��U�ݮ�]ZQ�1�#�cwx��*�%��}I���ܨz�g�`���\*�F�J�Sr��I귃��R:����ggY|��x����dC��>���\��^�v_�$�I�`���˻�e;�Q�c!Wh�DQ�V���v�Բً�4�N��v:�L<��UU�v�Q�0����f�PM��w&��t*�zU�$��D�>={�i���9�׌6ڱO|��@+G�LԄ>�LB�P��Ϫ^�{�� /a�؛�9��p����|JņFW6�n;&�u����?��w��/��2̖����/N����Ry�k^܄t��Ƿ|�o��%
B3	�EHf�����	�G���+��M�yW5�.�����M)%�Á��C�RȰ�;5����-��n��A��p`��p��ג�_St��`,M�:�
�y.�p?y��0� ּ�U�v'��8\o_[#�͜z{%��:�_�Ձ�T�o����l��,�z�ۂ&�'��D�FB�<g�d�8ͽh�
R�|�L=��1�������/��M���'W�Q��_����#�zK�5�Sx;2��+G�mQ�5�W �'r2>R ��y�Y�V��al�����i�\�HV��EHD�L��Ё-"��D��#xE��p�nrI�k%srG�q��� ǫ�������`��=�S�F���T�:�_�����g�Y����а]�A�;B"�E�SRa���KVUlci�	u�:�^V�Q�I%`A��#�[���0	�ƃ[L�Q���BUǤ��$aļ��錃�ݧ��p�UaZFq��_ݰ���f��ڕ���i+�P�O��]�k�-(�R0�q�K�>K�	�O�	f�����a0��y���m��Ud��k����>�ۥ�4�^̜���\���Vq?Ӎ�� ��gV�]�U��u��e���	���.��]'�GZ4���	�g�1����_��M�2�Ll$��k~ҝB���\Ƣ���MũA�ԇY�8$�t��f��)��4t��O�ؼސRO�9^bnx��5Đ��iR�����.Tv�Ǘp3�AA��Q iۈ�A��Ά�����+Ȧ��� ��6s��G%w�C�rs��՜N$�_��d��c�Hs�+�Z�x�)�����q@�3��� t��`p������H��XII�B$��>Z��f�;$۹�R���-�5�D<�7Ԥ�{&,l�f��Ac�@�+�prVyn�O���pT9� 9��E�?$�PL��"��ݩ�"��,���Փ���mE�+�N+�Z��r���}���ë
�*��3�TQ����'���Dh����'�}��~��呋�՛�����a�]��P���������M��4�����_ �g�3���iV9��cve-���F�=R�/@~�v>�^����1�ugC���j.��8w��}S���&����T֙��-)[=���ʿLg2l�W��P�&0������B#`�Dp�ĩ�޸��E������&��,����oV9�����"��`���j����;*g���KL�luFQai�x���`�mǤL�W�?���p);$�h�m�.]k��,��#D�f����o��~�����W��C�b��b0�W����(�S���8���	��Ct�p6~�����奧������HF��G�>�e�O;7�h��6�>�;�ru�4��}��LQLP\��<_(����{i�p� �'v3f}(`��܅�N$&g��ݚ�[�f�V0%G�wi�2� �B�����Cw�V8�������-u7�߇���[����V9�j��&~x��g����''@���36ӝ����,�(�i�}-�{����'����!��$�����!���x���	���0n���	؝��`�{� $����Hxb����	V���-d�g��woO�Dm&L�C������8�S���%�$q3���*�|s�}<>�'FG���b��6?�'��^.�u��,c��٠��	,8�>�4e�����b'Re�b���[�l�vn�ڲK���K��3� �����Pb��Wkj!w�J �+U�P�aZ�oj��I�Z���۸o�M�$�"q~�U_������GP��B�ιP�Y�z���y8||���{��{ڔ�I���z��#���)�f�����|�I5��m��M-'�h���O}�߫�fA���E|�%�̃/�j�t���g�U�m&�M\s�V2Q�j�EO�nX��ܞ�P9��5J����-B�Ē�,qn<�N�H�@�����&��J�|�.U>�b�n"�"���f5wTG��F�έ��+��Ťcd�JȢ�a1��0��e|���T��,!�_4��MZ`�?b;���7��I��D"�TG1$��=��Ä�X]�Z���+SP��7]���"2��j���̱�s�۔v�m6M���0�������ZZ\���쵅f;��j�3g筝U��>��:�Ծ�'�Zc����gea�&=a��c-W�*x^�T�1m\،�C�`�\ۥ#_zj���l�FX��`�P�P=u9�m���˄��~��wʣ4^�Ƨ��}۲�x�^��.G�����x�2/��)ѓ��9����n�Y�ɶx$=˰��� �̛�qQg`{{��QM�u�DD��e��%�����U��y%?��yz4�U���~��,�W`� ��^��+�����o�W�uk�V����#Բ���i�ߪ���yG�%#����L�_O�q��Y���~��nG���|�q���l�vvw@���y��{����p���6��*M���<���(�6�5�1��NO��jo�+.�����dk��5�<`$�;�xFm�7t,)���	DD�[�A�š���QF�6y��! FFB��&�&���{l�MjCi�^땰���x�Էe��פ�O��HFN�jnҴ�����oq s'j�'Hݱ�Fe��B� -N��f4f�q�EiS3�-q��j�SR���L^�!4~ŕlHD/LM�g���-��������RM}z�
걽3$Fcb��(b���q=G���<��=6��%ڲwe��:��O�����@�ۍ�1�R��|�-�AXq;������4�$�����g�n�OӉ&&�������n�|���BHn^KP���[��CP<h��}6�|3!$+��ɟ�ǮW�:dA3&�vk��!��&ȸ���	�_�]�-o�m�n�i~�"�#l�6=�U��q0"O�݌�\���Qi%&���l�rz]�y�LL0�����a8hhR�+�z|�1z��b?dW6��B��)��Kq��^�|�U��P�׻��v�W��%�iK���E# L��)}-��+ ұȁ9���x���/��|R��s>׻�5�A��zն�o���=����L��a��"[�J�[�J0���)c�fXC�@�Ew�g�K�5��\=���/�Rκ�
��Y��hUO�Cģ����,5�1��P)7~�O�7v��[`.��K�1И���%�T��Jӯ~��l��L��^��Y�\���X��l��x��
6 M��I$-,iXn�Q�W�>DִAi��e�Q�"��j��r�M�I��%,q{��F�|�V{G�IfJC��X�������ň�	�ik�������Yo]��$�TÂ$�:�z;����db=�'��1e� �D3(2l�ߣ�#x�!��}�R	D,b 7�m���	�t�x�+�N!���ix�I�X���Q%��%,�3�\���
®���p�yytd�1�X"3j�� �%�G�Z��d%|�U+1J������"v�e�\C��,to}��%O�w�22��(�����bl8��V���zǰC=[�cS�~^Tn��$��c�*ۻ�z�VQ$�:�����jԻ���f���@(�Z���PL�v��0�O.���.��^�I�p���J�u��v�	��a� ���I�+>f�+����H(b0�z�"��O��:ԁD��ccۙ�WT4�1O���d���GX��zWV��F,*$�UP���9Ȕ�`�h�����\� ]�|�:k�� WT��t��[��`A�ZG�u�ـٽ&`�z�`���V ��_a���<��kVn�����%�<l�K_�H��a����gd�;\�va�ss��l����y�1@������L��ዖċ��c_O����9�!]e�j���N�9�3���"��(�j�?��]�S��9��?0�^�Q�
D�����K�5���in��޽��yL�������5 ���t��,�Cv֤�h
k&��h��ꚠ�v�h�gXG<�Y�f��5���#�j�������XФ���M6�_��_ňS߀�G��������A�G�lCǳ��aH)K��ӂ�iƮ�6#�
W|w��2x�l��B����̪imsi�b��|�bb��x���EeLE�j"�<���t�rז��
Z��,�5��}γ>�8o��Ǐ����X?���V��������D,3�祦F�x|�j5�gm�؆��,T)Q��j]�'kԥ�D$=E.-���TwM}�:�{#.���s�@�_vF� �L/2l����?�g��.�z���9�"��D��D�m�3mr����n�gmb��	�r���*a�;Jg�Ո���7Q
�ݓ�:i�G/FDL0�K�3��`���U�w�GX�j�� ����0:_g������:���C�t��Th)&��ltDE�S�2;)�U$���g�b����� �����%����,x=Ni���B5��N�}s�閩g�g�;��(0�7�>:B�*��X���Y�
1Eo^���a]q�yI�2�	���Q��-Q ��<��x�)y�/FmBq��^�5[�*=u�E�gB�vK0��bS��!h'� ���)�@@�[�҄�ԡ����V:~J֠"�1��t���Q*�hs����;�Fۑ3�9��p�,�b����e�̔YMG�h숳�dBx�l_�"�J��z�Wbޞ��pC��T@�i|Z#yM�a�t�gO1Kޫ�rX���ߵ��X�w���'ݝt=�&:P�=����tpk<�" iP�R������ b1�!����Yrk"����\��]�3I�@yY-�&�d�#�_Q����͐��*]�Ӕ^�BF�^�<ͮ���
��́����X<I�7�D�F�$��F�/'C��������P����1Q�|�+�+�+�6�W��}�m����\��ځ��C��m����@��o �=�T����F�Ds5�����ϯM�iD�r������+o�x���a��1t�*�_r�˴R��(��;%�Oe �s���7�|�Oi�%�s��V�+���ֺ�)/�6�q�`X�]�}�����=� �j(�����Y�o% �U�ˊ\w��57�^�����2�Q7��V,뙴_�s�n�}A�V���/�~-8IKk�O�64�}�^�Uc�����/��(�����	\A�a~쎨6q�^Q�5��7b�r���R��2VK����&�;��xG��-�Ex:)=i��׌?����2��χ���E'P4{ ����eЈ�/�Ȫ���<��s����;X�^���?w3k�E�������?2;
��o$�H��Li���<�=h�[k�2�W.[I-��	+VŌͯ�/���
%�ه��F����-���6�->���ih��0��zf�1�t�P]d�>������zY�-ןծ�2^_ ������6m������i���{�p�������ݸ��Q�?%��.ؖ��κX������js�vaP�Y�W?��ɄoD8��l߸Ǔ9X�RM��ۓ쵮r3�|����ܮU���p�e&�ہƏ�"1�(A�[:�^�_?���Eҟ6D��IU��l;��ïP�BIq�gk�L)��c���ӣ-���E�N=#ؘۉ=;q۲�ۢ�X�$ܻ��ENn��ˮ�P;�ul;\X�R�O��l�{��-��-y�w��.�R��M����'I_�qZ�F���P��ܰZ8S�],��@���x�[�y�x�y@�/jU��a_�|�����y+��� ���~�Ϣ��!����9�v��V��X��ˉ�jٲ������JG_<-��
�r�ak�\r���B��<<+}�5j������j¦���D�[�88E�-������F�(�D�   ���h�HB�=�XQz2��=/D�*��
�_ �Eqd�� ��=-��R�B�J¨��h,���l����_�>l6;J���fl����8!�?qO��Ͻ�H=	3��]�Ē���8wSfj�����]���/$s�<P��-=���K������cf��G�:��7����b�˴�(�x��p����q���v/L�d6e��.ca�4*��U?:45[�`{���7����<�G��o����1\�<�ށn��jg؋>7�޾�Hc����W8F������D����J�Dq��0tz�����mz}[\�\��n�W?=_� ]��������鲖��R>����Ц>Em[z��Aj�	���dٻ
�����\����|���c�����������m��.ytl��ճ��HU<����Gp�%7B���1b�b�5l�\y��������-�;���[�}Ni=��q��Cʗ����Q	hg�����=�������,IXW�pW��]�����ֈh���o�!*����~XLI�c��C�)-��?O{{{/��x7��eQ����cݳ�,M��j��!5�I�gi�s��-�����ѵ輦~�24�)s��l�W��Â`*�Sgc$��1
�\d~���������R�҄ujZ5��_�	��ɣ�%{?��g7,��c�W+Ǖ^-]Wܶ*�=��n��ā��_o��P=�I/�X�����e�8�L�u�ϲ<=�������'�&��,�L���ʇG�ɢ�;v񼩔|��ayԏ�t%>z;ڟ��+Y~0��kst��Wo�����,���[��������s�r���5c����ϝ>�<������dRs���mV67��>/��֡�ʍ�v�Xz��O�>���<x1Ɍ�$P�[��,s�����eS�����P�M�g��Q�bZ�����g�����W���t%I���5Ɏ�C��㨡���yA���~Z��b�f��]�VQX��Ы>B#��+��*-��bU�M�L�Lo��dy���|��"�C>�%��c�����l����AƧ��C��$�J6aE�h��h�1붪2���_�!�C�����g��gVW��Ġ�EU��2|�y ��A��B��,1R��4e��$��L�t��X����Cs/��t �H���R�߇�6Ј��Z�7&�]$ċ�y
�!�Յ��
(�T��(h��25���O��V����i|��"�6TJ���<Ƞ��c�&	��o�D�g	+�Be��t1�^4�еsz;��ǿ�H*���L�H��r��i�q��EIHs���rc���k���_�,;��1�#?Lx�Et;���\�f�qg��� �#��Z*1y�H�)���X�R>b���`$��0�kNHpb;�&A�`!�#�����2��kP��)qu���Â��I����*T[���rZG۬E�
��T7F1؋��R;�*%��'�ތ�4V�׌���0V^����s7$>Hk�Cl�D�_�h�V�4D�0TBs�������Zh��^�g��*zIT?)��|�����V-�f�� ��=c/�π�}_b�O*L} ��
�Bmo�n�3�(,p#j��Z"������ŷ�O�-D��bh#,`���*��<W�DtTk�?���c�A}yPXB�F��%4���]�$��%����
����LfHYSdx��g�^�����8�_?����+��ܩ�f����@�ZK���etW^��z���դ2%���]�Ќ�#��;e���j���<	��L�|��3 y<,���e>8P��!��k���Z�jB�Y�긤����
�c�b4Xi���`B��q?��)�t]�APe�F^���1�N�T
!��-��R�͸�Ex�w���	*�_��;��|Z�4�(�F����{E���A������P	�9����RQO��U��!��(��4A���ZvA=ի�u/J8��{W�yo�,�ã���:p��|��+������
Ś�-i�+����*�i�^��B@��X�<XV�rWL��"� �$�p͔r_��0�Z�S��d��E��/>&�ZCŗc2�j@6`��6��Q��	�/��3�5�ƍ�=e�zds4ٷ���@qHz@��ңhj��^r۶QN"�������O:�W��z-=!��X��D�'�����k�ץ8݇� ��
�`�%I���T,0#�nXf*�|��Q�$ ;��A/2�&�5�Ίр*��_��!��f��T1�(�9p�E�
�G���	�/�^Q��r���!�J~Y��F�Pb����g��A�9*Cm�E���\���� � ����#�_z�/`�����P*`툫�ڜ��lh���<�or���Q2�	E��b놤�賓�,
�u@:��\��.��Z��#P�ɊYZ�ʚŁ�k����_H�O3t�&�M�5-�����!��e7J4��d��QvE�Y���n�,O�*���V^������4�R��PS�Cnx��`_�}�8��p�L�PP��3.�P�Qޭ�XL���2�pÌ��Ec�u��� �;$�<-��FT���_����J�@՗�~,�_�0��"�+�ٍ@%�S6k��+��ޣ�ahAB9A�ؔ�$��2a�E��Td.��U���N�+d�%B��3�c�`��,fݾɿv����]v����%�O �8W#A�s�O���=�r������`gr��^c�,Ww� W\m1]��i��y]/����b�*��ͽY��hT�}�G��b|���a��L���pL�9w�z��[��j�EX~ �-�e��,g@�b.�H���G�0�����Y��B�N=��3��!3P��{�@�*��0��"�"�W���$t���pݳ��&��e܄�H��3?#�E�TN����R��ְ`RY9G,~*<�tE���A�%�Pb�@���z�ʀ��H&�FZ�BL��A��Ju�#���^~U�]S�@I��f1o�w|��4 �Z�M3�l!�=�nt2�f�t߁ �/L%7\<�?i+��r<�G6F�<��9<�ʦ�y+.�-��5�t�\!PB%����)�b�ы֠�-mn��&Y�!�ʳe	N�s{�?3/�S�	<�<P�M�J����F-}�_T-��-��WP�h�tTx����Z���{�N��7}��et^��ӟ�$�b�"��0�h���0:g�N��߁g�Ac]���\$j}ɮ9���m��=3%T�r�����Ӹ~�ϔ����0d�ȷH(��:X�K�|�ې�,D;կ�^_��W�l��KG��.���7p7���c0�ƈ+�':��?�_�
�g��f=4��H*r��0:2v�:�c�S����]zq{a���{P<�,D�����s&�N�3U��<g�h7e��* %F�a�����|V��\�x��E<'��-I��T���[E��x���c���N4\����:P�\���SS=�!���A@e_N��", ���N�f�{_���d�o��A�|�s3�8�8�h<3���iO�
Y��	�i{Fu��뚦���D�.F��(�ľ�\��{��o�`3.������h��ǧ�,���U���{������nd�"Z���6�~�`�r ى�e�#E�J�E<�~���,��>,�����e�g7/T��������h`{R牫*�C�c�=c�d\�����F�����Z��kE����}C+&YP +0�r�����F�J?+����ۿlC���N����2 >��*�0�vC1�����)}�eg^k�T&w����_��239j�E;���aV>�c�4�e5���;���# <�1P����T����r��*?�q�ҎB(�L������F��	�67�h�ѕϨ��E�^�n��y�.;��G�G���6%6�K��ߚӬ��W�F�.�������З̓Q�D�tr���c�=�F�&���.����HP��mE %�U˝%���Oc�ۦ�\�C�4�c}1`{�������O+�&�A�2��� ��*^��ɢ��'$S��/�ћ����I�-�8����I������t����冤����[�yg5N0�i�!�����H�*{�uTҳ�QK\�n}9� h�n(�1�CZ�k��ϔ���cH��(&Y���93#�M�.�-zPIj�XӃ�����2U'�ė���Z�/�&�K,(??�����JZ�T��Y,B���_�j�7��/Y����2�o��/���5��`/.���kǵ�g�~��b���%�S�pL���m��Rw�E��/D��[z��@yE;�THnA�]L��.������Bo:�v^�(�vuSW�!/���ۑ�n�a�:�����Jis��g�}>0���v)sݭU�We3���RGE��;ȄQ�{���2sNx��B��C��6/\��z/��E����^��~�~����o:�ڹdq}c��u��;�ԅ�b���jCY,��1�<�z�I���r1���|�K��9��c�x��~_�-hc~}��a���Jy{#����l7���ms�{0��'�KM���X�)I�X�����(�]-)<�.W̄��=�44$�ud�,Q�$�WUu���ҽg�۝��|H�J�کq�#yN7�;8�>=~d+㻩��+� F֠U�����) ��m'zZ���i�m��3���s�@s�0O��׽�����g���
�Gl����ar�ڰ�D��z6���b���s�6�լ�r����MQ���k�G���W��3���� D�&��.QT��8w#�B�<���Ak�MU�X�>g> ��=Oވx�dz[��7b(��`̮<��M�ѕ�[��(c�+�`7��ܼS\ȕ�I�#��*�bGYX��PYPj���ݿ�ey��-7�<%�G�t`5FK`�*��u�'<Ӽ�䤊s�L�nc�5XJ�B�9��p�刯�Qt�m��[��$�J�P�Ejkl�4�����vE䫖�1�pEgk-�0#ش��]�UԳ�[ ͨv�D�"��Ӱ�0��D��+ݬ'fhC����*�.	bh)]6�D`��2�z�'��
)�|�%�B�c�t����r�V+Β�=wmzps����3E�-�ܿb"���j�;�E�/*��WV��.w����Xp)#2����8�Ւ�'|�.�7V���8��/5��?K�<u��ۊ�ݓ�*QmE�� Q�}�N^�dJ�W�)�.��q���rv��3I�{yv�D�ZjK���O/��T��ٳ��H�����łv�yPQ�� [��B?%6��qV��n�'?���v�� ������F��-���W?A����H����diӜ!�.�������	�땳�'�jG��ði��>k���#V4 c;�&��V���w�2�.���H�����>|4��%u"��3��mk��Qm�bwٲ��ۧ����d>�:d{�R�OϮ΀��Q�9�?�������c�Ae�v����޶}��#�"]sPt�[�g���	
��)*Q ��Ie��A!E�/�\ �'--w���?Y�8̓6t���O�F)B�<��f�c��ڭ<FH�Î�̛��1�&���C�+o�w(·�y�K�T��dY�*b��Y��mpW�<��v�祾�e�r��W����]�IXޭ���c�sg2����R���.d1�S��~R��i��~̷y��	'�E��E0R�P�5@�%�7�u�㜼�Mٗ����R
�n�*=�&eٓ8.`��F(u(��>o��1�����i�S_C8�7�ʈ#M��D�������$'�4��N���o3��Y���P���}��xj�SWݑ�>�/1"Cva`{t=�/HR���5"qn�� ��6g��E�^��\v�t�ME%4�d|�h��8� v$�	=&�	��i��U����obn	{LN~b�!-�\D��ڌ�!yIa�ط)�>f!#C�g�ޭPh��G����\�_sN�'E�ٝ�ꟘW��7Q�ch��]��65�U?�#�應����l��H9�������e	8���vo���n�w�@ov�f�ɤ=�jd��DdWn���;f���og��}sC�.=�c�\�N�6X��j��2�T�u[Ci�k��V� �u(��XV��P%.&��`��첩���i>v�8M�?Y6���G	Gw�MHP��^���+�D��]O��/G��S�,�i-Y%J7�
l�M����詊��cXȰ�޳yRbjo�|-�����gf�<������/�/p��$~���r���Uh�tt�e���F�ֵ�z�މ=��nE��i���E�M
�n���ޥ6����yu͑R��g��hJ���T�>a�h%b?��G>�b��@�I�g`]&'A��_�geT����Xzg��5��̈�v���.
���I�|Ɍ@�W�;�T�޷γZ}��x�y{�5���1^<�����j���EI3���7����&����k�4�U/�	(-F��\�r�'��������@���8�J��֎�]2���$���Pd�	B]��N���\����n ��J�_��/��3������|�j�fX��}R�+���̨Cmg��ʒ��@�Wm�����6�x����t�=jQ����/ķ_y����Ü���D����a]� ��$b�:ʕf3w��4��<�jwL��o��4��Y���4XK�<����õ+ޗ�Lz��S�_���ʟ�o�F�����7^B8��=�z�{ON�7�,���;X_��+�~q��(�δ���t�&k�B%Ж���q�l.i����n�c $��T����|��:Y��V;���{D�k���\x#3�v�ֿ|��I�C՚GCu��U(TNgs���*��#����x��pC��g��0��z'MX�hb�aeF���)��y���O?7�#�e��������V�+�g�{cW5P�r�>�u��vl\�<)��N*���-���r�v~~u_�G�rB����t���MH��-�-�(��4_�>k�b\Lq<��(Q�}���a]~-+M
̯:奪�g��9���t/��wc���w"a��|��/�&��s~�ԇ�c�v���5���?r�i���4�#S�+����z��Ǉ��HO����R��8�+����P�����:W�,��o�Ӵ��?_WJ�������M%�ul�]S����D��p���HT��u=r>���[WG�?c�'�w#��9�$���
��&�cF�	��G/?����3#��W�����=X�R	�i�ΔJ���=����ӊ���_�<~�^[Y�����r��-��o��j���q=�����q�Ĵ��t�j|�ר�ul4�ھݎ%��b�v�[�Ap�5��r�~����eɷ)�ն�������C�S�A>�}-o-�L.�/�"�ռb�E�����ĭ�����MM{�U>�o�7�ZjouOݭ���۫����V-�l%ow�iG2-�[�����������?/5H��oxuN.�0��Y�?���'���! ����������s���|/��=�������5�[/u����~���5v��G.K]�b��+O����Oq�c���T��I��-S���5}z���e݋4������?���͢��!��ϝ���CM������d=.�����g5���h�2��S��}���w��7';��Ǯ#��U�wI&��u���Ƅ��>�a�p�czUlNT���)��2|����������R�w�k"�?H�7OѶirU6���/���5���� D����e9�ț������#�ֻ����7�n��h����t����`���"a?rx]$d���]VQ�}:��z�KŜ��o5�奢����s�Ef��@SBv��Rc���8H�xMw�J�;M�ި����-��5�v���7�ĕ�7��`�d���.9�M��n�#1�ڏ��َ���{�8��?\]q"T|^~��G�I��ߏ���]��zP|m>�q4�'|>(!�iV�2��z6�D2��k*��v<�o��`!�x�$�<�^E:~��zжyc�V2R&"db�B� ��^X�\{�,ï�U�Ѳ�?�|kP+��)�Kk�L��F"
�!֚�}�˔X:�>�.a.]�d�=��w��?�K�C�{�K�{zԽ��nwwX%;}�m�A-����������ApB�vx��*m�����J%Б��
	���S{:������/Za����!٠�U�9�qD�#�9( <T<
'�*���<J��D@T "��PT䈀�"��9�χ��wm-]Z��yu^�����6,�ʺ����oF�U��W�nƯon�L�9{�m\���V\ȵ�W����˼�Uw�/*e䪹�q���r�sdݛ2gf�oЕ�}��Sow%n�M��s�vM�ѿ@l��nE�ޫ蹲gM}��ߝ^�=�ߟ<�����>~|����K���}]��Y|�Ӌ��A=)����e��S��fy�[Z03E8��W�riLAS.��',`W��P��������6"m�r����_�(,�^�ұ
l�t���S|�!���(�Y>�A���6�)�l��Ps}��C�gh�i�Y�z�y�d\�+9G��57�o7,P3r��魙�I�.��v�cy1�MJ�Hz�+���7�����R���3nF����ҔM-}�QS�/�ͣKP�.������w�)�Қ{���1z��3�r�}KjQ�3�9�i��pW�1u�UW�&�Vt�M���$���8\�4��U�S���EkM�c`��#��^�%�^~��G��Q[ڕ2E�tJ�pY���90���5tP0������!�Og�v�Y�]�<\�ՑPn��Ni=��;�DL�E�ò��[ϣ��0#��R>�o�{���Y@���C}��m�e��U�z��5G���i��#u���P��k����Lk���G�����o�jX$v���\y�9aF�[<i>�h�o��]xX�]^�O�x����4�c%S��jO���5PKL�Xϙ����eZD��*��x� ��a��p� mQ�%�j���O�>d.4Ƿ�$��HWL�!q;-��������L�3�1��.W��{�y,N�����$:�2�E�E+,d���lr9k&�v,�P��x��=�<�0he��ښ[5o��S�H�S�D��N�Pҟ~T�m�-h��8k�	�N�[����*� �0�Ea�庰h���K�����3{ޚEo=���p"B�-����I�F���q\�LRn��qt/�.�,*�6$#H;��F/�U�1j�4H/�L��'	;o��4��7��;�LI|��!Wnagj+��p�Ɍ�g0O�Ԭ]�VB_��:	��x���%_I������kM�٬�m���v�_���U v�f�c�}�&��f�����E��4�S������w3p4�%�s��=��g�x'*~~0�J�@FK�g>83�0��4�N���!��,�Cy�4�^��Cp�0.�JpW-c���:�Wi�����$���rdm	��~��[4�^�Ҕ1o�$�����Tؚ.��Ɲ:"f���tE�tʿS��:���]�	��O����c���=�����/1fs�|�{�&���+6���Z�R������Сo8���#:�N�g�SlD����[� -��A��Irm���s�����E��q�k�~4Y:^X�c��fIT&]��[��b�Vq��n�<�B?�A����j�_*l|Lru�E��&Z�񆕗^���51�o�G-13���u�����h�\�R��N
�ė���H�}z,1n8���F���x���]Q��CV(g�W�f�٥AB.��}�֩�����l��	E�������v�~PX�����v�X�z��%a�ý�U�]$1��KA�2�h�|ahэ������:X�s5�H��˲:��&>'��P�*�L���ч�^�fI�[V8-Ab�ճI�� ~�+7����ͬ�Я�;�)�|�.Qn�lt��VX���7U�NO�@�g)jHN�iL�7Ȭ�>�M�� V�����쨐cD:+�Z�Wx5��9X�3y��H�b<Mz׭�\�A�x��L�lU#wk�PZ�V9�m��_UR��Q=z'hx��ZL����ڛ��c�<�;��'a� 懚�&�3�z��M5ܠ�g.�|����
j@�f)N�J�o�^��hD���O��PL��ԟdj��qV����u	x\��t��/�8{���`"�\*ҟ�Z�4���d֙�oڋ�&�UG�"H�S!�6�%a(��ci�;8�6�iԺ��R:�Z2�18��z�Hw�ða��HkwK-�zмUġ��k
P�NjB�RSX��v�v
#e]��Yo�[>?j^q�p�R�oO��y(��
�SZ9��G��&Ŭ�~j�C��c�h�s��SW23˜:{s�A���k14��r���s�[�J��-�V9A�V�L�U!�]Բ���K��k,�Ҥ�"Yz���&l���Jgg�E2�*�w���)��c̕C�݂��g�eq�T�Ԭߖ哑̶{���Ysd�y���Tn�ųdX�۾ܩp��d���;�%�0c���m�Hl^77���G�4"ͦ6� g��y��$��1s���{���̘aq��[̤q��2�n~E]��B2�8äZ�it|��Zq�R\�gܠ[�פ"�ޮo��Q���T�%Ժ=���Y����w�'Tաa��%$l�1��w��IBf��Uz-��V��ܐ�!r�B��Iz�#H��]�����i0OиY�lOk��k&�ҵqI٤dx�$dC<J��kU����Ȑ''�4z�����AgW*T�G��C�?jM����O�9��Pm����ɘ�8r�u�*[�j���!�T�E-cJc������s�����_�Ty,�*�ɌR��[> ���/w�'�C�M�L�f�Ƿt�+م��=Y;"{f�A�C�g�wW�_���F3"���<�C57�/$܌�h����yA�H�垔��p�[9ow��ܶ��0&wG�6ò�_rHtLR,	��c����T���r��e2��}ԫ0郸j�����l\��?��Q곫Xx��+�L}u��#��9��;`Ӆ19%V�k�����n�֧�]��Վ��dNY�'\�i�.+N�G�q�� ��Zf}]���|��k ab ��M4��kqJ��h�|[^%�nF���j1=1��5l��'ԔN�4�0P�
�[��4KmK��i	��j��Phn���+
�b�Pp57Dj�g��U�KA��崏8��5M����-#]��@E���50g�e�i�;�䗳��N�i
�|�P�����O':M9��j�vRnsқ̼�y���쏷��B�H�8��o�#���,+f����(�.�Kd[��eOs�r�z1�+,&_uiP�>�E�S�(�������綾�#/88�_�ZZ��m�;��ο�� 2�,��J]��cl�ت�	k��}�ק�cUP��MO7�K�9�^�`���wI2��׾R�����U�	Aβ=��o��]�,׫n�/�,XԂ�9�p�y`+����j\�������'H�m��Y�*4�ڷrqXU�����`�0{M���s����\d���q׻]�on��֌�(�ei�f�a-����s��"����<�Qd�4q`z
�� �p`?\��`�tW=�i�V#��t���%Q�\�+I�q���Dh,�\&c�K�5��Т\-J27�..d�[#����.�K�Ϥ*���uY=����*��+����1~�_���0�_���;ee�ֽ�+]Ks|;Ѧ�J�8������'k�fI?cdO�(��Z0�L�)�2�A5bm\,N��\�r�NJ]�#���-']Joe���\�-��A!�&�Fh:�C�ggW92ЋZ��8�AP��htp�rb�2�z�RW��2�����}�.�޸�	;<�G|�\|6����C�p�cu8�\�ɾ�c���ϼ��n���s��d٢�pHE������3ۓ���z�ǖ�[���lk��l��2e���hj�y�����R��ɧI��d43�mI���jZ�L�l��|tt�L<yL��g�Q��tK���5V��_;��z�s���m��.����^��S��c�������S�7)B]{��T)5��趗��=5Y�^�{{�¾�vfR����y��[ݠ=�{92O���S\�o������!��j��Gi��Ɋէ֤7�US�ً���p��s�Ţ5F�l���8���(�|$�N�ǁ�Qn�[���G-;�A�	���>�)3��>�OFSd��Z��vNu3Ix:��\p�-�85�x|��<˹�;�M%��y�(��җ�#^j�r�s�f&u7��E[&(�
���[$�Gk*��5�C�cD�麸�Zg��a��y��j��c�&��o:,>�̣�\92�������o����#.kN%�1��x�9,����R��_��=����%Wiǝ��_��]HG�9�N8Ld"����=H|�ȢU�{�r"\��ŧc+Zl��8}ĦQIc����n�	3xMV��%.̫�3�g��}��*���7��Q'K[�K3[�3���(�c��S�mK	MkIn�'�����P���,z��K}�=r�6�K���*SY�c����
����AG����vF���l�����Ͼ"J�h��C���>&�i�>ڰ��My "_�B߯���p;c ���p���~ �XRp�<3�C�~��0����S�6!���{;7�Sm�����.�S�t����E�~/��bN��;;�9KKG�]궴��a��Z�\0��sZ�G��numm��"͝��,�տ���a�c����)�EI���x��#��/g����8~���m���dl�|��
��{o�64-����rK+l��2-��&ƥ��d��$���+>u#�l<j9��Z���Ɔ�u��u-��.��_u��:��q��u���z�¸�ׂW��x���љ�cU�3Ǌ��N�Y�ۗ�=�c�{�����z�<��8���7�|q��O�J����9��#���K���~��q��ڬb���f{�S�6�]��B���wAe��l=���tE���=r�}�P ��ᏻ�O;��y�W�O�0rH!)�y@��}������Ǿ����r���۽g$H����ws�nh���1!T�'���^����?����	�����������e�k����ۑ�7���%��	��2�_�_NX ��@��@X(�������^���[��55� ��q�჏;��'���Sn��j������.G�pZ-	 ==�d�����@{>�e�&��P\nxpZ�����{w�E��&��W4-O]�����`�u���^<���|��K�q�k�� �'��%�0WԮ��~�}10Rx�&��P�k�)o��� � 1t��L@*b��T@+,d��dA����0 `c3�)��3	��� �-���_�22��Z_e�����y�� @:; rg��rĤ���ٟ�l1���y����`�@R���Y j�_DJ�Q刱5�Ë� ���#��eAt�
=ű��_4e�2�u�Y��8ݏ�Խ'>%�@>��Ϭ��r�����@h��u�������y*s�	[�Wlk��=��]����uw�,-��z,e~�N����I��zK���6ǘ����R_����)��Vิ��9k��E[ޏPs��>�T�{����W�œ>j��&�vw9��`1��t��*� c'�y�yceE/p���W_����j���\P���ay�d� 1-`T�h ,��	X� 4�f��?�y�ݵ0v�qZ�+h�w�b�Vj��G���4�����Yʪ�ڮ����w�r���nU�.\��=��m5s���:�N���V�aIm�@-AxVX@11�3�fC>o������}���h= �`w���9�:����S�=�s�����������@��a
�#��ù�[��$�� "��0V�g�� ���~�n��@��	�ނ**\iYZ�yqS�s �
>�'��������%�UUS4��k���8�+����iaabbb����O��� a��O֯��AB�D�p�Z����M�1ϚE��Z����]��-U�҃*)���Gȭf��a�8�I*�߽�'j�i�觤l�8�wH�Z�-]O8���9!�����s�s���z�r��ä5��h��>YWOM]�;5 ���·�J`�03�m?8�	�0��<04:A���o�g[f��M=��_��"���4��rg�à7x/܊=�#���gز��J�-?L*���?HH��ٖ��vM���4̽!1F*�1]�w�^0:��`XZ�}�^s6�'*@00-�0Q	Q���������hc�g� Cl�;:�0�!�Yl�B�+���21����..�IŶc<v��h %(B�����~ Ȓ�-0NT��
��K&� ^�#��k*�Sn��v�~�|hhXr��z�W�`R	���r7i�dN��a4�tphl����5�GV�N/�f^NFC`��q�3��b�<��J�vjFBC^�(����+k7��Nmi�����H��#[*:{��yy����Hm��:��wg���2*�9��m�q�J������ړ��@��耎�J���yy�G�yC��8��k��w2?
7��?�q��u�8@@C�c��_+��8vC��q����c{�.�)�v���o��wp_����G�N�]��c�m���'�mC�������_���3����HR����ps�c\���(�X�XPX��'�XE~C���67_�"V!��X�\Yh�r���� �x����Y�	l%��������־�����z%� ����.{[�Ȅ���F}[�̿�j�7`1P�f���Wd��[^�h^a�7@��t ��V���@N�"������j�������=�1��Y���(��۬N<���k��� ���I��1��%&u�ղm���j�M�H�h���*'�{?Y��Ќ��C
ޱJ�������+�׺:�$ �q�?�`/�[ �I����^�.5G�JO�fyg]=t��_P� ����u���uq���]C��S���	W��D�sZ�v}�Z0.�w[uO�L�ǈc�눊�`u
o�R�
����*?�PJ����� �O-���?�)8J����u\x`����@����/�'&ge�G� ��,�����Nΰ��2/�@��K`@D��)^Wf=��]qڭ�h�uO�kѦ������@�|N��xW��	^�}֚��O�T� 1b��(�@i!@w�^���O��;��S�U}�M���k�b4���o���v��8�>P��9�/�l�X����ZM�P�C8�>�4��C���8�̃?5@׃j�7��C�L9����8 �AІaafd�h��Pn���
�/�g
��I��QGZ��r�30Ù��]���l�^	s&��'�
�yG@ȯd}���J����������i��q����l6�AG�6�qގ��ed�� ��:Lz�6�yV�.�_x*N�|�}�����u�P���7����o~�ڈL�k�ѝ�ȼUe*^�������x�x�k�
����|��d��w��t`�hps��_8Ko�������3������'���_ZC��P�1���2p��-Y�7��pM���F�Y�����j���W���q�C��9���a�v��� 5?�(���ֽ�~r�������:�������f��.�R/������/�w���-��W`W��ϒ�E�Lcń�~�r�!��^����sB���4�/k�`Gf�=F�� `��AT� ���?���N�2O��1 ђ6�]F�~ @g���W0��na���ޯ<��Up���C8��%��tL��2��r@����t�s0m��O�J��i�jd��>�Or�~_�lX<�����Q���̿�������`:��,�F���Dv@�0�`��B�_RBT�b+VD�_���'K�k5���2ö�:���e��,��'>�=7�ꊭ[�㸇y��rn��/��홽�g����\�Y��+���]�-�&�)ٙ����o��@������^�
NC��;����l#T<0DHu���`?]N��9O�zrn����r�+I��C��Hmf"��`V�KpXlR�[�Ȁ���¥�����6��A/�N� ���݊�N�n$$���
Oo]��#�D86:�o�5?/*|�$:�H�)��+�n���r���)�f
/j�\1����X�dW2aQ�̅UMH/��_��T��J(. ��WE(;�w�)�;�I��D[a���sIS�i6�kE~���ݪ���F�7����_��[%G�u5ef�v)��˰UT��T��f����+Ewo���JA��'H^z�F�N����[�]�er��X���Hւ��� ����g��{��Ab�!KQ������y��WqW�j�<¸by�N	��M+��<6�ְ�ɊB���؟�~���~p����ÿ�V!z��T�w]/A*������/�M�	$'���-�1�khhJ�a5ޤQ��a�S*��+��1�3O���A1%bV��7�����#y"��
�5J	��������"��g}N�a�=L���ݟ���@#�Ȍ~�#�qV��7VQA
��\��>��ٹ7s��D���5K
���wh(.�ItW�ĺ�{t7 �]%{�15�z����Sw�V�Tc�P�\_�&��I���&`�B��
�� �����z�����= ��{�|$
��0�<��������:A� ��T>*m�}o�"k�P��o���hf�������DD!c��j�ܰ7�c�
pN���[�^�0
�O9(.c���
��ȭ]�CT���@�b���u&"����6�M�B0.�ꔪ{�������]�u|+�E��e"'�E�į�:B���� ��GH8������gj+`�����!��8"҉Б���#�/���B�$T-ǥ�+�w"���/�E�v)����ߜ���X�7�N�b����������=�v����$��?����#�j`�H"y��X�N�uW���^�)�=0mȁG
���D+��>'�/$C"�Z�ݭi�h1��'���@�����B}a�C~~�b��_�*��!�Qaׇ�XD�����Yݨ���9�I�}_7P͉���Xy�}�z0�rߠ�0�Hv)�頯����]y���+��<"�Ϥx�f|+E�4I;�H��=y�=�ݟ5�**j����`�9e%'p�z������xG������P/I��H��OJ7�蜎C�����`���[�������H+e����(�&"��Ů
�Z��J+�=�:���ݻEHt~1���2��E�zt�7�6��)/F�� D��A�����^X��;���'	� d'c�[�[Vy �'&J���7�Н3m�����䈆fS#4@X�#q�h����=A��A��q��٫5llр؀l�}�3V�Y�٣4f��C��@ Cj�#T-9�=r4���e����k;�`��m���Dc��'Y9m�r�B�>�I��K���p�+���l����mSfF�UGt�AG1�ʧ�+璮T��*���3*���n�gL��ʬ��˥Wі�:n����y�T/���|��<��<��r����߽��[�t2*���4�����E+���X�VZ6�y�b�N�;B�c=H։�P���B��gvi|����Ap�e�X�w�E��]Ea���E����$��ȭS�̅Y���j��#b&`u���u2�E��6F�\) ��5f��HJcM$P��ZQj��z�:�V���:�A'[n�'��x�I=�I�]��~���_��kE�Pڝc���\���҈�s�-����(���ɭ3UW���S�u��Ԋ �擿D�����1%5�N����E�3K����괊��UCED�!�m�K`~q1���$�MpLB�j\�1MJeN�)��X�S�"����O����5�l{� ��TCc7X.�5C	���r�<b�{H�L���ⴱZ��j�$u�_�Pw��'-�ޜ�A?����Nb��_Z���m6Rb���v]�-؎���H�K� �����'��$:�N��5iW�	�K���9��� �����Y���k-�|<%'/�e�l���Z��UV�?5Vď�;h���T�0�ݲ'N(�S(Ԓ��E��f��j��F�I��i�=-�O]Bs�sVP������0Oy=`P�B2($S���q��I���4mY?�����!��x���+�e�����x�O�oj���U��tsS��YO~��'d�'�� O�"X��*�u}�� �dv�0�N�)��8�o��P�gݼ�43cd�s��jH�z�>-�r�����k��6����9��C��x'T�$'�B�#m��H�t�4��8��C��;�	���F��ڢ����L^��
��m���p�w�<��x[ڻC�g+|R
*N����*�
3UŊQh0(}hB|T�l��b�]�;L	�qm�o�f���8F�DN��p-�����`�h{���#08S|r� ��hǃG%��I��<�#����Ӳtղ�B�L-*�]�:�8�!���y�o�H:�p����ACI�N�t0 dX#�����JB'!�����I�A�� �2�(AE��#���NV.(�^8./�����wF���r�q�^Yi�� ��4�е��.��dVRu�� ���w���㨉��ܱ˓6]�T��Yz�R�c��ܑ;z5��\�)/?�3Xf��rfEmp=��Nq�>+��Gs����x�}���.L�DG R'��% ��e���|!̂l�C�G�@�w�\G�t2
Ӥ����75�tA(�ԐJxb� ����3���4�����=Ѭ�?;`�R�!Xխ!��U�N�����mC8o#ęp'�t���q�< ې4t��w��5_�~����D��32AX�i9�v�y��[h9�r�i$ҳ0h�M����&����z����K���)<y#h&'4��E}p̓X���j�MO�o��F�H�0�\26~y����y_I#�r�x��'o:#���B�2��L@��}T�G7�y�O�:�¡
g��?Ii���ࢤV�՘�S�Q�/�!vqUfkҍr��i��F���-�Mͬ��S=���O��ܭ�A|�.T�D��
HMOE�vT�W�.������i[�#b��5�O��8֏j~ Mb�9E���z�s����k9OI�Uǡ;�q�yO�Nu��F�5)ȓ��-�/�Иqj����>=Imu������)���b4���f'6����M_6��{�i��-�b��|��9fB�����/�1�6m'�~_������*I?�#t����k�Ő���[�Q�YT$��B��A��cY�Pb�N�I���
8�����D�U�U<���"j��ct%��JKIw�{������߉�����������P�\f[��|�ex�E@��~�{\�gt�
%j1�A�)�T�3Ӷ�)��.1.�geWJ���YU��X��X���S��Z�l���O������8����m�g�s���o����J������U��:�tD.9aB�K{$(���y����,q�������H��/@ǿ��Bh=!\�t8x՜8�`�(B��������ߟ���DZ�y	�(È�IU�����0E��n	� ����_��a�B���9P0Y:d;�*C��j��#�X���u�o>;	,�'��N�?`��E��-/��U��V�Ř�-1c�Y�S�-,�Z"����a���0I��i�O��	�V��,�j�E��,�c�)��ӑ,��-�&�-�����ЋA�ZH"�
��&̂���
w�. Ys���v��;#�k˾E�)���,Oi�%���;t�{K�5%�R$r8D�-���h�-�Oь%gO�7��o��󫼵"�^d��D�U��=�cw���)RGɩ��5u ��B,�
�o�4&���>x�e7y���BK߄L�P�"�n7��bƓ�o`	�3�-0�&��+��t	�-�gCē�q,(D�d��9/�����M��|hP�7��mVȓڗ���/oo ���V,������ɍ�ɘL�E�K>�J��M(&��Ӱ�o���E�!�}w���M�$v;�C&�уb/��~��ᨬ��T����q:�d��n�O��1���E���9���A�Mrb	���BS�H�a�C�{�`oGa��Aޅ��r��KE�!���"܁;8��k�xBē�k{���+���d2{u���AR}��#���M-[-��[�o�E��Є[��W恳�l����&z��RO���П�{t�n�N���6 �o��+pdp�O����������h���G�s�Ea���54�[�W�/\D\FnhE�zO .~�K�'�|���A~�hN�${�v-p88TF"ہ"��ȹ}�^Ghk#���d��<;WW�iT\�"ް�u:���|&�& Ot���D���'(�&O�J�f�P�������}T ���ѵ�E��W�l�cp/�D�����)l�e�������p\�"��t�Gdu{p�Hu����GI��S��Lw�&����؟e����Ҧ"�& �_ۨ[�r`��'������`��v��\��9��$���w6"�y��E�!9�]x"���xq����{ ��WVUZ�TX�ʹI�zp;���X��W����M[���A��]�"�@�\��Zկ~���"�����r��/3'L������/U�4�2��h�j�/>y(E֡G�]t`�t�1���Q9���'�k@��m¤0��������roj��	�=�ӌ�{6����nU�~�]T"�!!ҵTPbz��u�E�B.��<"�f���� �q<�p�[�{��z�;]�
�߸rz�(�?(�{(E�B/6y��(PyWP"��B/|;��|�'"}'�H���s�v�.ŕ}͛�'�jn~�)��ػ�r@q=R)4���^�XrB�'�{�q,���=C"�� �U�*GjZM��yv\�Ro�����0�F��G��ORq��c�$MHF�jV�Yt���iY ��[Ը�"hi=_h!7(Q$�G��b����&�Z��X��p
�]a&'��tDԇ�� �'�Op�C�x�	��l�>(�+q�v$�w.7�t���jd��#�� ����n�[q� ��[����`N0��5��X)�m&���8�}�)��:�r����$�#8��6���W�R�ȿy^�ʾ����[ߺ�$a�I;�?a�W�9.�>b����_�Ot�D��Jv�J�"�ad0v!��e�88� �0�&|%e��D}l3�{����,_�!�2_6ȿ�پ�[?�˰��Q=y~���C�=��6�	a밆���`��i��R̢l���y�����5�U���!1-�-$}@O�n�1C�1C�1]�|Z0;p�1C�l�QC�< �G�EԬ��1�gp��C�G��t"��Tb!7}��#MNǈ�!�+�����#�M��h]��u�Lv�����v.�b�!�b�!�b�!�~:n�*�b�!�b�!�g"���?�^YAHb�!�y�yhC�1�7`,��I�!�b�!�b������Q/~{ ��ֱ�GS��{(CR�����c�=gߗ"���!�i��(�9j(�Fq!E��˹��_2�ٮ/��~�C�"��������B./��`b�!�b��l��Dh��1p�s�*�����V�"�5���M^�_|�]�����������z�����d�L�d'��F����-=��������؎�~�������>L!
�T�Aw*�^�Sߪ{�O~���=���T���Sߪ{�O~���=���T����.��l��nz}��p�c����Ʃ���NS��;�Ʃ��+��
����F� �j�tUCT��re��j��yb�2�\5L�<�\�b��j�X�L�WS5M�������LճVʦU3V�[*�T�[5l�eS����ƪOo�`��Mg�*r��5�ek)ƶ|r��M\��|�P5����x��A���H��Վ������|��̠P9���*���5ȳح�(5S.U��������+`
�wg�MX���R� �k`u;�ʮpy��]�hΧ�{,V�O̹���~֑��/�Y�?t��)�PS��:��垜��K|��|s���E0

r�S�<���F)Ο�{���Z\�wg�JϷ�Y��S�<H��]ÝN��]m�+��Ot�]��wg��o !]��{����
�Χvx��������R�)����5s��B�kݞY�o !]��=��NR���*xW��� xE��|���-H%�W"����L�WB
��˥�K�W"�ӡ��:��V5�C��(��)��sBTW+�|gz
[p���3P���/%�����P�A��j��z���	j�4jbH=du��A���+�w2�̟��yk�xsp4���42 s*��p�O�`宓���Q��y/؃���o�]���C�c�2���g�m��~�٢9�T�uf�C͢W 䮫*ċ�TlR�f!n2��Z�v�k{-t��2�ߩ�3���BFv�Q���_ي�60�� #�*AIGQ	?�):�m�*��"����\�v�s xT������sB���y
���B����o8щ�L9�R�!�(���Dŕ�����fW}݇�E��OL1��G85�v��d��sB*\!�y�ux�.�37���a
�|W6��7%8���`	_iU^̇=����%H&I~Xd�0)��1�D*����C}��w&�O%So&��;�_}2lp9��Xv���]�@鼽V���������(	�ڜ�9��
"]�15��v�<�V���s8'i�)���o�_��� \�w��k亁��O��p9��gש�̾�oL�u_� ��>��9�Bw��N�2��PLR뭀K1����J!�Q2�ac&�ؚ4d�<- �`�N���q�o��:����4��6�չ�̾H�L��ل-���y�P�4W��S��j�`�[�[�n@n�%�̠�}C���� ::��>�u|�P��[���|k�����ۆ��0����}��D���ê�ۂ{����6·#��sA��� :%j;-'��o�}Zqr^x�D8��]�O=ٷƮ�<e�&x�>v^/�Dܭ6B��(C`|��#���v[c��μ3��s��Rg���JG����ۿT���4�g �C����̾CK�ge���u3����RP��a�⥅
���oB��x\�t�t|C��u٧^;8�c�Go2���b9����!�*p��N�Й<Jl��B�g%BQ��_hFDFNnr�'��@J@�,�ކ �0+�W���d����z�|��fU�����*rD+���Z���'*N��-_OR�ǂ��D��*����>�,!p�i�ퟖg���~5M6]���z�[���R%F�#hF�<����zNL*��mw�( S�r��$[��^��J�GX#����I@/W���i�^����4o�T0vj�b�ݺ����(_�?��TcPL��B�,�wcGA�
��;�
��K2x�0an��V)L�w;\'�]=$�I~5��m���q����C��,�L�t�x�����P�գ���O��)�w�Ӻ�/�)��mS�Ll��j�_�.���^��V`k�F��+ܩ��f��1ǀ�56]�;�3��JV����X]$�`OG���w��򽯩�ic�)����ZB��R{V.�jq[2=h5Z@&hݙ��v�*�[�s��Wz`�ȡ!Sض��&^�"y��3�u���3�{K�]h�l�~�������v��28�(^�հ�)����F���l�l@�h�h:H g���Y��M�N�A�i����L/�N���X��(^h��z��%���>{�,���z,������t=�F�P;����+���q�Lc�i���s$��,rJ�=3ݡXI�3�è�R�`3��fTiQ���@�U�� K��B�!���7��r#��x\����H5�-֗0fm~�|�Į��x\�q�{"��A5�&�^i�0� �
֙<$0�(X"����ɷ��I^�o�<��ͽfcD��˼{]U���5�xD��#fo����W�:�K^��I��]�K	�X %Mߡ�s��U(Xc���x2<�YA�j���������騀�|�ENXl���F:�(���l��A�WY��>�F� �J�0/��ǽ�}Р�Z���дH��U�k�Dz�=l*�W;���Y�Fr�=T��X:1����"ş�����QA2�3p�ez�$�P0���W.�t�)m���8F1~M�G$l�h��N������ó�qz�ȉ5�1n��K��R��[�l0�3)]TGUp0:�co�-��e4ċ�#�)f���9_��,[��R���P�I͆�-hJ9����IJ����������^ #���F���lz��~�r6�RW&o{l���y�a(�z&���3����0��L;�W���#e��]k���d���p�EV�k��������a���1��Ɖn�}2�����WY��I.��
o��b�ar�H�1I ��ݖ���OlͲW�J����4H�Ҍ^aP5*� |���tw�|Q/��|��Gm�8��(.S��j��9��(�y� %��&tH�6@ �)��3ѣeU�y���Ks���x����"Ơ��e�������C�ne�`��=����a4��@����UJ�JL��[D�?e�K��;�\��{.������*�N2qiعhO���!��}ͤ��Cǃ�!Vs0�K�?y;?{Ko��v���k��KL&� �V��2��^Al�f`Zo����6W�t�����|&����rf��`\V� ř�h� f�ޜ�'���V�8{8��\3�	�GN������t�㽢,f�%ج3���;G���s�w�̺��i�������ĴH�6���#փ�J���B��U�K6��5��[���&��mBl�Zف<��Ә��=�!W�\���~D�� ���<&ig5��2�yݲ�V����f�l���ZJ#��L�)~���ꏉ-Ä/�Ne�}�D8۱��9y6g���3��:i� �Q��
�ײ��V��y\�<�6A��>X'U4�9��M�]���eEw�g^�[�1����X��r��ϵ�9��f�'z3�#��%eb��>����6�G����s5��\��okNq ̣a�o5���Ĵzu�� a�)�8>K7�� ����o� ˴���2������LB{x mA6�ց�9C� �}$��vƽ�>I�ʢ�ȦO,S� fw��������L�8Uf�0��^+��ߨ������`�>f�M���������q�O��s���N��0�G�L��@^A1�T��8kA���3� �.S^�Pq��؀�H�M��&�����ͼy_N��5`m��	���0@��l��c������R�/�a�v�3{����w�Q��� ���x�a�Q�R��$uH"�#AO�NI��7 �2�[�(Y#�<XBf>�u錺�%�	�Ȣ큩~0��a�4����+�ױ�p�7Fn��~K1�P�:?�զ�z����C�E����KK.]ٸ}���,��<���nni���%��^�K|�5�Wtj��Q.�O��'����ڧ6\�o����(2��H�������bO��x� �Y�X~��B�u�y5�:vR�.��	���A����=>\	l�/H*Z�:�J��|���@o�q�C��˚{gX��$��@:d� x��3e�EN�x6΅k�{���҃,��L��4���7�dYdHf�g|m�_�/��� ��5+�\�v׿�}��0�����g��+��a澰5y��z���>�k��5��_��X�E"�
W����M�Z]g.�,;:�:�k��!����d3�x�S"�YP�!O�`�~u��^��_�)�7	<5$���Z��yq����Ѿ�+�r�hS@����+��
ڴJ�v6�3�?W*�ji1��3@�t[����am+��x�=��a�+r]���0#7�l�e}��@�5Q8L`�z��$H�_f|��0����_����/�������e-�|�in[BUBLX��`i�/4F�I֩ό�߬�	R�'�R�r[@��`�G��ڱ��6�Q���$3���vuX�A�*:PӋܾ)�y:y
4�JTG���#�B���Q�Ą��)%�3k\���7�`���m��s'1�R��q7](��A?��g�am>`&p��ѣ� hئY����^+ު\�bj�y���e3)F�Ω�|��[Eߞ��kNր٬Ù:��Q�p��##��M6���ހ�m�_�� Y�2�(�O��Ѹ>���/�x�a?I�W� �D���8��&Ͽ+�뉋hP��S	6փ�	��c�Sw�NL�r^l�`zI��&�^pC9��������Z�fo��~�@Tx���Pu6���� � 	�xv���S#�(��у��%l����y�����
=0ƛ,(@�`�N���<���n�6Ц� N���~3��Ƭ^{ٰ}fFsd,s]X�ٛw�p}�- ����~�D�Na -�p�~�b�߬4��6W�������m
�0��r\�~�~-(/�~��$Ox]��0om��/�,0-X~��8��{��4;#��y�]��\���L�[;�~�΅`��0Vδ�k��_���Iў��N�mo��$��<��X;em���+x��Ɇ:�Wo �k�@͛���zf�k��D�.��6�����#���!��m�A��t{5A����G?l��?5���@-����J��f{��0���&��:���E���,��8�sl*5T�nz�����z��|T~�ɬ����̕��Ɓ�A.-P]jFnC�z�Om����x�y+�|6L�%`���nw�{�rFp�p&L�,�kgcd���$"��ƈ��>�6$�z5"��ί���@���k�zG� �/�0����1.�1�܀`*��b�>YX�-��Ǵ{#��+��5Х#V�mXK�Of�Oo��K���M�rs�V+A�d��
�1\��<��l�jȿl,Q��h-��R;Tї���₉���~Ц1_6u)���U��������~�l�V�4��&mh�@���f������QN�;m�K!V9Ec�Xc����0o0#ǘ)U���4|5��k	�(����{I_�AY2�p�"�H .׹|X�0f���w�R�O+̶4��B�K��*�Y�}�
�  ��
/���e�Cg!E!��лyٜ����2��2��e�g�N8�Mx��#@�4y|jSf�2�$����5��Z�
��y�z����4��)j�M5I��
�/ ��%�5l�e|�,�y���۟i�@�qP��i�楣"y�x���� �<h�?b1�K���g����ɠ`�+��oa����T�j��*�5�'��aL�+4���; ����z2��z�+���ݔ��y5{b5���p��v@3��� w�)�]Y|��0��Rç�S�6`��F��)p��8�I�����f��h���8;9�{Xc~��<	e5��7�6z
B�vd���<:�b_�|ʺ�͢��ʻ��lf� 6����n;��|͙�y+��P��0��7�#:������;��Y�QF�+�c�V/\�:���Z<��uR�Kc��E>E�ۊM�� |.�"�Y�>f��~УǖC��V��;��(�#	�u�<yd�W��uK���Hן5��W��~��Q���Ggk�����z�ٖ�F�H�����.�u�M{�O_�X&��Ud���D�hU'���>��~�p����g�LZP8�5"��M���/�xR�������?��:]��'6�j���*2����2̦F@ ����a�1��q�͘ 1�i���dѹ�P��>�����J��0�bc`�`�D�"��7�é����i�J�Z^s������8����t0.aĵr����!4�Ϋu`r� ����$��(�`$����Y��#7E�1H�&����1�����y	��=C��:A�r��������:,fda2��v�����{��=��s�{����y���K���b2��W̚��d0F^������P5mV�ٮX��y�����6	�-x��sJ#� ��i��WG��;[R��%�[(fU���?��!�s�%ʯs�N`��%�rcn�8��q�Kd@݉���Y���EZ��p��J8SX�}��Y��9\�����V���`�w؞�օ�H�)�e�֭�eg��׌aky��+���a��$����iԅ�����4���t�2��3�Σj,��ɋfϱL'ľ%Ќ��lk
�+H2븒�9�h�J�Y�����4cB6�FT���O�TB�9�'�:�{9���Bv����+SP�_�A��!0L��f���I&�꿅j9��� E� �2c�ݔ��\*�@Q�:���4�XE�Vܟ&Í2~�AOA
>�D�zm�\|B���Pv��΂�O����;v6��m�1�!cz�z��&,9�v���Jt�	���ܱ����Y�L�B�6�?A�XM:����Y1q������y���>��r}n9}l%l>�8��ۥ`��&�D ��r�|^�q�A��q��h���|f��B
���1��fXr��f4.�V�u�n�|�� &��ȭ(~bg�֐Ѕ^��!)Xh�:���9��`ǚ@�s��|�t:U^��sRck��cҦ�|�5�
%2���)��ɸ�ڋ�m���ՠf�Ff�n��!���	Z�rQ�� �w�@���)A��hA��:�߇����A8kD?����*)��eřn�����h�jh�S%�z/1�����r��\p�S�����!���?b_������/v@���(@�L���2-�����(P�vAa�SE��^�����I�K���Խ`qM��)�ē���Kd1G+��VCaZ-�*�Qe�x�*e��&z�N��PT�s��Y��!��"`�X��u�0������4��B�փ�>Yf���0�B�Li 
����P�1�6���� B�^ׁws
���*����ok��N.�a��O���8H)�P�OGӾ�+�N���&˩`��)�su�D�)u ��� c�l!|�!B�
�}��z���_��3k7�RFӦ5BAO��O@=�Ѫ �H�� �*Š��$6�$[��"���=�of�3ӧvE��|:m:{��r�Iɤh��G��G��_�H\�xZ�1�0G��V�R�S��jc��N��}$��5CH!r�Zvߋ]�R
:!պ�"s���I��J�ji흣��Zwߋ*���S�� �� 9�aƙ"�v�z��',���zG��_CY�� �(pcǈP"��ŋ��h]�����y0�~��z���?�m�j�q��(� @{<.9���r��������α'�=�B;�Ą�"�$ ��P�sD�	%�eÿ�y�p
ܷ���>C�!X$�P� <�u@r �
�5L�(���z�$6?T�3����Q�o����!@^1HE��`*���qQ P÷ ��7�B%�ϯy�]�	�=�!E���n� xp��
v���@�J�Dq��hc=!��#��u�@"Q��ʲ���M.�G}���D�8DQӧ��^ ����!�%ߥh��� ��B�{��
)�8��c}�>.����U�>C�k�yx���_<aX7�w䑯j�0f1��E7�L���O��}o���냌��e� W�]�1�L�`Nv
4b��ms0� $!;C�8��|����e��9���	�|:;�њ����C�L�P˩NieL��qJ��%�i���fG��"$X���l��	�"��[	&�0�*���ǈ��8�sN�7-�E�YzyO}�G
a�$�"ö���O���d�[G��}�z�������*��εb����7�C�û^��/^�f����x�na�^�ӳe���&�>��6�>�����AA�ߵ@���=�����D�Ø�&�	P��Su�g���8��7�TO�_����V�=��t���v��^O&�z�"p}���4�s�����d�l������I���=�J$�v���3���y�輌k��h_�G�4�&�J�EE����=�p�BV�FT�
�$i�����_l�"ԍM�&<������a���\�Q��Ř�������Q�"����7>��Qъ\T܁ͮ�����xS���>��]��`?Zz���խ��KE���L�y�}��Y7��Ǻdy�#$�]ލc����L~<� }y��6��]�$�P_)����cB��U݉!U���Yn���snLQRN�c	�g�:��L'���G\���F�XĴa,��|�'I���@`[a��>�ǧ�RJ���g����!�ҵ]h�TJ̛�?�C"n�i����t��ꈼ��Ӈ@Qy�C�$��o�c|*���U*�o8*����,�T+M4����l�V��F1�Q�f�/f[�C��(�7��uER�\j �yaw!ؾ���M'js��.a`Pe�ޤY�ڒ�����g�T$b����|/�>�7I0o'֣>���&��������ԫ�%W�������%�$/�a�D�͒@
�8���ݳ����y��Fڎ$�j~�T�e������`K�H�h��΋�(gE�t`gFFg������|�                                         �`a��� ����`�    ������]݁� �/ ��"   ��"  �e  ��.  P��M  ��&  ���]^SP��I  ��M  �]kSW��I  ��Q  �Ew��VirtualAlloc VirtualFree ��1  �t
���5  ���i  �> �!  jh   h   j ��M  ��V  �F  jh   Pj ��M  ��R  V��"  ��V  �vPS�n  � �� u^���   �>�"  �7���׏PQVS�ȃ���R  3��t.x,�<�t
� <�tCI��� �>8u�$ ��+É��������[^YX�        �ȋ>�"  ��R  ���ȃ��^h �  j ��R  ��Q  ���> ����h �  j ��V  ��Q  ��1  �t���5  ��"  ��-  +�ty����3ۋ�9  �"  �> ta�N����>�"  ��f�����t��t��t �,f����  f�f����  f�f����  � f�����뚋�"  ��A  �t��t
�f�f��� � ��"  �F���
  �P��M  ��uS��Q  ��E  ǅI      ��"  ���u�F��I  ��~��I  ����   ��   �u�CCS�����S��E  ��I  ��[uo��   �uW�F�"  PS��u  PW�   �������&  9�E  u$W��J����E  �{<�|;x\;��E  _�W�F�"  PS���  PW�J���I  �2�����F�F����"  ������X� P�"  Yɉ��  ���a���� h    Ë�&  ��;  QP��I  ��U  ��G  P��Q  ��*  ��R  QP��I  ��Y  ��*  ��^  QP��I  �Ѓ�_j0��h  SWj ��Y  j���U              kernel32.dll ExitProcess user32.dll MessageBoxA wsprintfA LOADER ERROR The procedure entry point %s could not be located in the dynamic link library %s The ordinal %u could not be located in the dynamic link library %s R��$;��
�t2а��s������u���ZÇ�  @ ��Y /w�< �                                                 v  �     �  d   �  >  � �                                                                                                                                                                                                         �D$��T  �L$P�  ��$\  ��$X  QR�L$�  ��u
�����T  Ë�$`  �$PQ�L$��  ��u
�����T  Ë$��T  �  
 (08@P`p����            		

Q��V�   W9Jr5S�������@�\$��B�|$�����   ǋz��B�ǉz;�s�[�r�B�|$+���   +�%��� ���_�r^Y� �D$�T$���   ���   �����      � ��   SUV��W�   ���   3��|$,3�󫋼$�   ;�T$ v3Ɋ8�\�(�L�(C@;ŉr�   �t$(�r�rD�t$h3��t$�D$   �L$�j�t$�D4,�����   �|$$��   �D4(�} �]<Ã��E@�D4l|M�u �D$�\$���   ����%�   +���؋ъ��t$�Ët$��f�����ʋT$ ���|$$�L$�D$��@I����	�D$�L$�t$�b�����   t_^]2�[�Ę   � ���   3Ʌ�v;��$�   �1��t"���   %�   �D�h��3��1�|�h�D�hG�8���   A;�r�_^]�[�Ę   � QSV��W��xr0��A�T$��H�T$�����   ʋP����H�ʉP��sЋP�@�   +���N$% �� ;�s���   ����3ۊ���;;F,s
;F(҃�
�,;F0s�   � ;F4s�   �;F8s�   �;F<҃���y��y���   +�+�_��L�D����   ^[��Y�SVW��3�3���h  �V�W  ��0>@D ^�   �����@��:rދD$�OPh�  �H���Pj���   �:���Pj��0  �,���Pj���  ������`  _^�  [� �D$�ыL$W��B��@    �B���   ��0  ���  3���   ��P  ��T  ��X  ��`  ��\  �ʪ�   _� ��  S��UV�kWj���)�����u��`  ��   �3�j�������D4F��r퍻�  �D$P��������u_^][��  �3����������s��`  �1Ѐ��T4$F�`u(j����������~N���  }R�L4#H�L4$F����6��uj���������j���x�������~���  }�D4$ FH�����  �s����T$$�KR�������u_^][��  Í�$�  ���   P������u_^][��  Í�$  Q��0  ������u_^][��  �ƃd   3���  u@��r��ƃd  ��`  �t$$��  �_^]�[��  ��   �^���ED Ã��D$SUV�     �D$$W3�����|$�[  �N����=   s���AG��|$�)  =�  �   ���������P���T$��   ���   �6����N3�V�m�����0"@D ^��r2�N�A�T$�N�N�T$�����   ʋV����N�ʉV��s΋~�V�   +����   �~+ˁ���� ��3�V������0@D ^�D$���D$��d  ���h  3�V�������5>@D ^����tv��rq�F�o���r1�F�V���@�L$�N�F�D$%�   ���Ћ����V�NsϋF�~�   +����   �F+́���� �0  ����Í��[�~r1�F�V���@�L$ �N�F�D$ %�   ���Ћ����V�NsϋV�F�   +����   �V+�%��� ��؃�s���P  ��t0��P  ���P  ���T  ��P  �K���X  ��T  ��P  ��|$A�8;s��+�@��P��;�r��D$ǉD$������������t;|$(������D$,�8_^]�[��� _^]2�[���  �Z @�Z ��Y �Z                y�/ ��/ ��/     kernel32.dll   GetProcAddress   GetModuleHandleA   LoadLibraryA             l�/ \�/             d�/ T�/             q�/ \�/             ~�/ d�/             ��/ l�/             ��/ t�/             ��/ |�/             ��/ ��/             ��/ ��/             ñ/ ��/             б/ ��/             ڱ/ ��/             �/ ��/             ��/ ��/              �/ ��/             �/ Ĳ/             �/ ̲/             %�/ Բ/             2�/ ܲ/             <�/ �/             H�/ �/                     oleaut32.dll advapi32.dll user32.dll user32.dll msimg32.dll gdi32.dll version.dll advapi32.dll oleaut32.dll ole32.dll oleaut32.dll comctl32.dll wininet.dll shell32.dll shell32.dll winspool.drv comdlg32.dll winmm.dll wsock32.dll msvfw32.dll ��/     �/     �/     )�/     ;�/     J�/     \�/     m�/     ��/     ��/     ��/     ��/     г/     �/     ��/     �/     #�/     6�/     J�/     X�/       SysFreeString   RegQueryValueExA   GetKeyboardType   CreateWindowExA   GradientFill   UnrealizeObject   VerQueryValueA   RegQueryValueExA   GetErrorInfo   CreateStreamOnHGlobal   SafeArrayPtrOfIndex   _TrackMouseEvent   InternetReadFile   Shell_NotifyIconA   SHGetSpecialFolderLocation   OpenPrinterA   GetSaveFileNameA   waveOutGetNumDevs   gethostname   DrawDibDraw      	 00   h        �      (   00    �         �       h   00     �%          �        h  	 (                 @                                        
aI�>�  <                                         #		�[$$�g**�y::�W))�Y                               84�b&&�i,,�l..�|==�{<<��aa�                    XD�h..�i,,�p11��PP��PP�}==������XX�6!!�   *         mV""�_$$�n33�r44�����ȟ��ݾ���xx��mm������[[�G  �    V((ɘhh�u<<��SS�ǣ���VS��?4��cS�ퟖ�ơ�������ww�y::�0-        Y!!๎�������RQ������@3���w��wa��~q��jj����pp�l88O    f,,i//�ee�Ƞ��z.,����1 ��E3��T@��QD��!��[Z����������__{    c++i00�����̥��l&%��ZL��ZH��3*��:1������QQ�ȝ����������    i-,4r33�����ȟ��a%$��F:��QA��h��E0���r
��FE�ǝ��������    n11G{<<��ii��yy�{JJ�e!��QD��ƹ��_Q��
�h ��dc������dd��}}��hhx<<e�CC�Ƥ��ϫ��ٻ�������DC��7/��I?��ON�˪����������Է��×���tt)�WW^�������������������������xx�������������������������ֻ�򮈈8    �~~!ֿ��������������Ӷ��ڿ��а��έ����������ּ��к�t���                �����������������������������мӾ�R̺�                                ͳ�
տ�f������ۘ���-                        �  �  �            �                       �  �  �?  (       @          �                                                                  #   E�R�4�   [   -                                                                                             ,  [(�_%%�c''�x99�L""�v   7      
                                                                         
      6u?�d''�e((�f))�x99�x99�a..��   A                                                                          "   C�Q�d''�g**�i,,�h++�z;;�y::�x99�p55�#�   O   '                                                             *   W$�\##�c''�f))�i,,�k--�j,,�|==�{<<�z;;�}??��RR�<�  d   0                                               
      4oQ&&�]##�c&&�f))�i,,�m//�o11�k..�~>>�|==�{<<�x99�Ȟ���ww�X**��   9                                              @�M�l44�a&&�f))�i,,�m//�p22�r33�m//�??�~??�}>>�y::�����ɟ���cc�h22��   F   "                               %   N!�W�]""�l77�e((�i,,�l//�p22�s44�y==���������??�@@�~>>��qq�ȝ�������JJ��ff�*�   Q   %                      "  [6�Z  �]""�^##�o88�i,,�m//�q22�s44��gg�������������Ѷ���OO��@@��[[�Ȟ���}}����ee��LL�E�X   	             RE�k33�\!!�`$$�a%%�s::�n00�q33�y>>���������ʤ���'"��zu����������uu�~??��{{��}}�ˣ���xx��CC�w99�[**�  *            2�uBB��bb�Y  �a%%�f))�w==�q33��dd����������[X����=4��WI��g\�鹶�����ģ���cc�����Ȟ��×��|>>�y::�y::�

E	        )E�m66�ȝ�������jj�q77�zDD���������ď����������u��kV��dP��^K��u�����ڿ������Ě�������tt�y::�z;;�O$$dD                  P�W�����ʡ��ʠ�������ii�����:6��
���������r������bK��wa��oY��~o�͘���rr�����ȝ��ȝ���ww�{<<�b11�                    _$$�`%%��__�̤�����������XX�d	������ �� ����RB����������v_���j������G<�j,-��||�����ɡ��ȝ���qq�m55�                e++d''�e((�HH���������ͦ���UV�t������ ��#��G0��fW���h��z]���o��r��7/���v43�����ę���}}�Û���yy�l77؄TT            g--h,,�u@@�`,-�ś��ʡ��Χ���PP�\	������!��t]��`D��	 ��(��(��)!������.(�|42��}|�ȝ��Ȟ�������{{������cc            g..!i77�e**��VV�ʢ��ʡ��ϩ���FG�Q��
��aK���f��yd��	����"��[Q��%�������1/��vv�ȝ��ȝ��ȝ���vv��~~��llD            ]&'Bi,,�p22��nn�ʡ��ʡ��Ы���AB�]	��=.������ZP��5*��}t��K@�� ������	�o �y/.��oo�ȝ��ȝ��ȝ������ȟ���wwo            g,+_m//�q33�����ʡ��ʡ��ϩ��@@�F	��7-�܆r����$��7#��lS��J9��#�������o�i((��hh�ǜ��ȝ��ȝ��ƛ��ƛ���xx�            n1/tq33�w88��{{�ʡ��ʡ������}=>�A
	�r��;0�އw���l����������rS��3!����	�r �O�e$$��bb�Ȟ��ǜ���nn��ii��ff�����            i--�v77�}>>�}@@�ɟ�����ii�@@�5�P�s!��A4�蕁����������va��3#����
�b�G�q32��[[������UU��bb���������nn        q33�{<<�@@��]]��ff��UU����������MM�p55�a!�o$��K=�㕆����������	�y	�j"!��OO��__�Ģ��ˬ���XX��^^��||������TT�jj        o33��AA�|>>��}}��~}�̦��԰������پ�������GG�v32�f ��.(��r^�Ոs��A5�r��>>��]]�ġ��������������������������ȝ�������gg<        y;;ـ@@��OO�а������ַ��ȟ��ִ��׶������������{>>�^$#�U�p("�w32��JK�������������������������������������ɟ��Ȟ���xxh        �KK���ˣ����������Ѱ����Э��������������Գ��ϯ���qq�Z%$�w>>���������������������������������ٻ��������������ع������        �kk�����Ś��Ŝ��������������������������������������Ȩ����������έ������ٺ��۽��ظ����������۽��������������շ��ʹ�Σ��R            �nn�{{s��������������������������������ί��̪����������Ϊ����Ţ����������������������Ӱ��ͧ��������ű���Då�                        ̰���Ƃ��������������������е��������������Ϭ��ӳ����������ί��ռ������������������ӽ�����&                                            ������_����ֽ����������������������׻������ѱ��ؼ��������������ʮ��ϻ�iı�
                                                            ���ϲ�E̱����������Ȣ��շ������������������������ðǲ�C���                                                                                Ȯ�)ŭ����������������������ο��ͻ�'                                                                                                    з�η�}����ο�h���                                                        ���� ��  ��  ?�  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  � ������?�(   0   `          �%                                                                                            *   @   g"�V�(�  l   @   ,                                                                                                                                                 0   H  �2�a&&�a%%�w99�C�      K   0                                                                                                                                      %   7   Z�N�d((�c''�c''�x99�y::�Z((��   V   8   #      
                                                                                                                    (   ?   e		�Y""�d((�d''�f))�e))�x99�w88�x99�k22�		�   c   <   (                                                                                                                  1   I�2�c''�d''�f))�g**�h++�f**�y::�y::�x99�x99�v88�4�  w   G   -                                                                                                
      "   5   U�H�b&&�d''�f))�h++�i,,�j,,�g**�z;;�z;;�y::�y::�x99�x::�I��   M   2         	                                                                                     (   ?   f�W  �a%%�c''�e((�g**�i,,�k--�l..�h++�|==�{<<�z;;�z;;�x99�{==�z==�_++��   \   9   %                                                                                  .   E},�^##�a%%�c''�e((�g**�i,,�l..�m//�n00�h++�}>>�|==�{<<�{<<�z;;��DD�Ě���ww�k11�

�  f   ?   (                                                                 
      "   5   T
�g77�V##�a%%�c''�e((�g**�i,,�k--�n00�o11�p22�i,,�~??�}>>�}>>�|==�{<<�u66�ƛ��ɟ���||�e,,�S..��   H   /                                                              %   ;   ^�S�y??�W  �b&&�e((�g**�i,,�l..�m//�p22�q33�r44�k--�??�~??�~??�}>>�}>>�u66�����ȝ��ʡ���NN��RR�O##�  �   R   3          	                                             -   D  x.�]""�\""�zBB�X�d((�g**�i,,�k..�n00�p22�r33�s44�r44�zBB��BB�??�??�~??�~>>�{<<��hh�ɟ��Ȟ���jj��nn��II��VV��   ]   :   $     
                                   /   L�B�[!!�\""�^##�{GG�Y!!�f))�i++�k..�n00�p22�r44�s44�r33�������׿���RR�~??��@@�??�~>>��UU�ɠ��ȝ���ss�����v88�����u;;�)�   i   :   %     
                             /   Q�P�Z  �\""�_##�^##�}FF�\##�i,,�k--�n00�q22�s44�s44��NN�Ӻ�������������������}}�AA��@@��@@��JJ�ƛ��ȝ���~~�ě���{{��PP��||�u77�C�t   9                          $  T&�S�Y  �[!!�^##�`$$�^##�~DD�`&&�l..�n00�q33�s44�r44��xx���������������}�������������ж���FF�@@�|==��qq�ɟ����������ɞ���ww��SS��MM�x99�W''�
z   (                    5@�U��NN�X�^##�`$$�c&&�`%%��GG�e**�o11�q33�q33��KK�Ի����������Ϊ��x �j	��4,�צ���������������rr�~??�w99�����Ę������×�����GG�~??�w99�x99�l11�8   	            	   KV�}JJ��rr�X!!�^##�a%%�e((�d((��GG�i--�q33�p11��||��������������a\���� ��@8��cV��RG��}u������������� ��~AA��oo�ɠ���xx�Ś��ɟ���\\�z;;�y::�x99�y::�X               
+^R��ff�Ɲ���KK�f//�d**�`%%�h++�}EE�n00��MM�д����������Ә����|
�����q^��TA��p^��A/��M<�歨��������������||�ʢ���oo�ǝ��Ę������v88�{<<�z;;�z;;�;{&2            *6@pV�n66�ȟ��Ȟ��ȟ�������pp�h..�uBB��tt���������ۻ���JH�|��	������re������fP��nZ��t`��fQ��R>��hZ�ݸ��غ�����������jj�̥��Ö�������uu�w99�{<<�z;;�V%%�X--E                        H�Y�V�Ś��ʡ��ʡ��ʡ��ˣ�������tt�Š��ɠ���on���y �� ����	��	��RF��y`������oY��cL��cN��mY��mX�행�֋��Ǟ��ɢ���yz�Ы��ȝ��ř��ɠ���zz�y;;�{<<�i00�h99                            Y!!�[!!�Y  ��``�ˣ��ʡ��ɟ��ү���{{��SR�V""�|%"����	�� �� ������
 ��'!������vX��cH���o���s���j��R<��nY��wf��WO�W''�q<;��tt�ѭ��ǜ��ȝ��ɟ���~~�y;;�d//�e88                            _$$�`$$�c&&�o77�ʡ��ͧ�������hh�Ɵ���fe�r.-�l ��	 ���� �� �� �� ����(��P>��������������t\���q��������������+&�t11��PP�ȟ���dd�����ˣ��ǜ��ɠ���nn�q55�|HH&                        f++d((�c''�e))�a&&����tt��}}�ˣ��Ψ���^_�p-,�� ��
 ��
��
 �� �� ��%��-��U?�쟍��y\���z��tX��v\���x������F=��E<���t00��JJ�ɟ��Ȟ���zz��yy�ϫ�����ii��GG�[77A                        g--e((�e((�p55�MM�vFF�Ȟ��ʢ��ʡ��Ϫ���[[�q-+�i ��
 ����
 ��
 ��%��3 ���e��(����F0������YC��RB��|�� �� �����r-,��FF�ƛ��ȝ��Ȟ�������gg��������aa�j<<n                        i..b''�II�k==�Y$$��``�ˢ��ʡ��ʡ��Ы���UU�o,*�V ��	 ��������?#�������Z�� �� �� ��+!�� ��*"��
�� ����
��OH�-,��DB���ȝ��ȝ��ȝ��Ȟ���oo��uu�Ү���oo�                        m23,�KK�S%%�i--�o33�����ʠ��ʡ��ʡ��ѭ���JJ�o+*�J �� ����O:��V��yO��jX����	 ����	��1%��+$��& ��(#��"�������w%#��CB�����ȝ��ȝ��ȝ��ȝ��ɟ���YY��oo��{{�                        Y$$KW!"�k--�o11��HH�̤��ʡ��ʡ��ʡ��ү���CC�i**�U ����aP��Ũ��YN��}k�餘��!����A4��YP���_V��+"���� �� �� �n��,)��DC�����ȝ��ȝ��ȝ��ȝ��ɟ���qq�Ǟ���jj��ww	                    Y$$hi,,�n00�q33��UU�̤��ʡ��ʡ��ʡ��Ӱ��@@�q,,�a��8'�ۛ����� �� ��F<��"�얊��~z����+ ������(������ �g �i��HH�����ȝ��ȝ��ȝ��ȝ��Ȟ���xx�ǜ��Ę���mm1                    c((�k..�p22�q33��ll�ˢ��ʡ��ʡ��ɠ��Ӱ��~@@�`))�F��1*��mV�ꢐ��	�� ��.��
��x^��J4��F5��1 ������	�������W �[��MM��yy�ǜ��ȝ��ȝ��ȝ��ȝ��×��ƛ��Ȟ���ffZ                    p2/�n00�s44�r33���ʢ��ʡ��ʡ��ɠ��ˣ��~>?�V$$�Y�z��3)��fQ��`Q��#��B*��B!��Ŭ��^C��qX��?.��'��	����	�� �h�o�W��PP��uu�ȝ��ȝ��ȝ��×��Ȟ��������ʡ���hh�                    l/.�q22�v77�y::��^^�̥��ʡ��ʡ��ʡ���~~�@@�P!!�F	�g��!��;0�މz��r��ì��ҭ�������l���`��T8��)�������u �Z �B �G	��RR��ii�ɟ��ȝ��Ś���TT��mm��FF��GG������ww�                    _&&�t55�y::�}>>�u77�����ʡ��ˢ��ę���gg��BB�Q%&�!�P�i�}&��TG��B,��ï��������������tZ��B,��%������
�o
�Z�G�N��TT��bb�ˢ��Ȟ�������II��HH��ff�����×���Йll                l//�w88�|==��@@�v77��ll�×������|>>��XX�|==��GG�d00�A�U�i# �},&��B3�ދy������������ƿ��:-��#���x	��
�Z�:�f-,��QQ��QQ��UU��jj��vv��uu��bb��^^���������ɟ���{{�ee                q33�{<<��@@�~??��ee��WW��^^��II��tt�����ؾ���ss��FF��LL�n//�^ �f"�t$��E7��~s�����������Q=�������v
�u'&��SS��[[��WW������������������RR��bb��oo��{{�ƛ���TT�w==�bb&            b**y::�~??��CC�|==��ll��XY��[Z�Ş��ٺ��ղ��ٺ������Ҷ���ll��BB��CC�s20�d�l$ ��1+��J?�㠆�矉�ׇo��J?�k	�p��CB��VW��QQ�������������ھ����������Ţ���aa��rr�����ȝ�������mm�|OOL            v::/}>>��AA��BB�s55���������������ȝ��ͦ��׷������ֵ������պ���ii��AA��AA�f%#�K	�k/)��C5��P?��4+�m��76��JJ��MM�����������������������������������������Ӵ��Ę��ǜ��ȝ��ʡ���zz            y??P�AA��AA��BB��ff���������������ϫ��̣��ϩ������Ү��ٹ����������е���]]�x::�u76�P�C�_�t31�~?@�{==���������������������۾����������յ����������������������ˤ��ƛ��ɟ���ff�            �IIe@@��``�ɡ��ʢ��Э����������Ù������Ǟ��Ȟ��ɣ������̧��Ӳ��Ы��Ӱ������ɩ���WW�q33�P�m00�u99�������������������������������������ܿ������Ӱ��ү����������������������Ȟ���ss�            �VVf����Ϩ��Χ��Ś����������������������շ������������������������������ն��Ь����������Q""��``�����������������������������������������������������������������ۿ��������������ɥ�����        �TT�\\x�~~�ɠ������Ϭ����������������������������������������������������������Ȩ���������������zz�ͫ��ڼ��ظ��Ӱ��ֵ��Բ��Ա��۽��׶������ڻ��Χ��������������ҵ��Ӵ���������hh7                    �mm�\\Z�kk�̨������������������������������������������Ӳ������ϲ����������������������ͨ��������������������������������������̥��Ү��Ӱ����ϫ����������||~���&                                        �qqJ����������������������������������������α��ß������̨������Ѱ��������ػ��ͦ��̤������˪��������������������������������������˹�Į��Y˳�                                                    ׿�ֺ�b������������������������ˬ��Ģ����������ӷ���vv�����Գ������������������������������ͯ��Ǧ�����������������������������;���                                                                        ϳ�?ӹ������Ӹ��Ǥ����������������������������������������������������������������������Ƥ��е������ʱ�����                                                                                            ���.ͫ��������������������������ָ��ұ��Я��ά����������������������������������к��Ȩ�sʷ�                                                                                                            ˮ����q��������������������Ӵ����������������������������������į�����;                                                                                                                                Ӽ����P���������������������������������������驖�ű�&                                                                                                                                                    Ǧ�3̰������������������ν�Ʒ��[���                                                                                                                                                                ���è�+����Į��κ�<���                                                                                        ��  �  ��  ?�  ��  �  ��  �  ��  �  �   �  �    �  �      �      �      �      �      �      �      �      �      �      �      �      �      �      �      �      �      �      �      �      �      �      �      �      �      �      �      �      �      �      �      �      �      �    ?  �    �  ��  �  ��  �  ��  ��  �� ��  �����  ���?��  (                                     r
 e! h  _$$ ]++ \55 a%% l&% `** g** h,, l.. z., i00 n33 m;; q22 r44 p88 u<< y:: {<< |== kCC {JJ hQQ nTT rTT yUU |nn vv � � � �
 � � � �! �7/ �3* �?4 �:1 �1  �I? �F: �@3 �E3 �E0 �CC �DC �FE �ON �QQ �PP �RQ �YY �QQ �[[ �[Z �QD �VS �ee �dc �dd �hh �ii �ii �mm �pp �ww �xx �xx �yy �QA �QD �ZL �ZH �T@ �_Q �cS �~q �wa �h ��w ��� ��� ��� ��� ��� ��� ��� ��� ��� � � ǝ� Ȟ� ퟖ Ƣ� Ƥ� Ƞ� ̥� ʩ� ϫ� έ� а� Ӷ� Է� ٻ� پ� ݾ� �ƹ ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ���                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                     ���                    		          B        	77]9     WbpJE[;   C7e>*Qce]J   []7& /USRC`F   ?e$,0OL';^Y   	YeMN)+& :b[h  ]b.LT1"4`Y]  EJ=qP#@[AY  4ein]4(-5hw�m^  ^yw�~tHVwsus~n   y��ymnmh��s       ��~s~�|            ��       �  �?  �  �  �  �  �  �  �  �  �  �  �  �  �  �  (       @                              5 G O C
	 Q \	 P U W b o  d	 o r  t y	 r r c  o$ s! Y!! ]"" ^$# Y&% ]$$ V,, X)) V44 W99 a%% d&& j"! e(( `,- h)) i,, l// p(" y/. 1/ k33 n00 l55 a<< g>> j99 n99 p22 v32 v43 q55 v77 |42 r99 w88 w== x99 z<< }>> _CC [GG ZHH cCC gBB nCC cMM u@@ ~@@ zDD ~KK bQQ eVV pii uoo xqq �  �	 �	 �	 �	 � � � � � � � �	  � � � � � � � � � �" �" �# �( �'" �.( �7- �>> �:6 �.( �)! �7/ �=. �<2 � �$ �" �3! �3# �5* �7# �A5 �A4 �K= �G< �G0 �J9 �BB �JJ �LL �NN �UU �QQ �UV �^^ �YY �UU �[[ �^^ �[X �bb �cc �dd �bb �ff �ff �ii �ii �qq �qq �~~ �mm �qq �uu �tt �vv �{{ �|| �K@ �RB �WI �ZP �[Q �^K �`D �fW �g\ �r^ �aK �bK �lS �dP �kV �oY �t] �rS �v_ �z] �zu �}t �yd �~o �va �wa �� ݆t Ոs ��f ��l ��i ��o �r �u ��r ��u ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ď� ��� ͘� Ě� ȝ� 㕆 蕁 ��� ��� ��� ��� ��� ġ� ʢ� Ʈ� ͫ� Ь� ӳ� Ի� ٻ� � 뻵 ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ���     ���               JC                            >":-                          ""::/J                      J%%%::::I                    ?%%%%::EE�>                  A%%%1%~:::ך/�              L*%%%111~~E:���/J            H1"%%11E��:~:����H          7%+11�����~�ל֏A        *7+1:���g���:����~:B      �D�!:1���Vp���������:::      �*֜�:F���XT`���������Ԛ::      ����Б�kQMOO�ڨ���Ք��ל:�     G���ĆZ^MQa��ۯ��{%���ט�     D"G����[_[s|�����nW1�Ԝ֜�     :D���Zqs��YfffSOl6���Ǜ�     /"����~M���UYd�cd\O6���ט�     %1����~o�P�v��caaM(������     %1����ji�Urw�}eRQW%�������    1:����:p���ܮt]O��ז���   �::~�Ԗjy����ub\
1��ԇ���   �:~����ă1z���bP!���㈉�ǈ   �~E�������~1h��xj����������   �E����������:'1������������   �������������:��������������  �����������������������������      ������������������������         ���������������������              ���������������                   �����������                       �������                            �                �����?�����������  ��  �  ?�  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  ?� �����������(   0   `          	                    ! : G W A U W ] S X d  j  l	 o u  y  v
 }	 x	 h u ^  f" t$ z# T## ["" S** M33 P55 \66 T;; [99 b%% j#  e)) j,, u*( c22 n11 c;; k== r33 u99 z<< ~?@ UEE ZGG ZJJ [RR kLL tDD }BB }JJ d[[ gaa iff okk qoo uss yvv ~}} �  �  � �	 � � �	 � � � � � � � �	  �  � � �	 �
 � � � � �  �  �$ �,) �+& �2* �1+ �4, �76 �(! �*! �5( �;0 � �( �' �+! �6( �3  �?# �C5 �E7 �B3 �F= �@8 �J? �C8 �P? �B, �H= �G3 �P> �U? �A/ �B% �N; �R: �R> �R< �CC �JJ �LL �JH �RR �RR �[[ �\\ �TU �[[ �^^ �OH �TG �RF �WO �YN �a\ �bb �cc �jj �po �ss �uu �xx �gg �ll �on �rr �uu �yy �{{ �~~ �RD �YP �_V �TA �YC �^C �aS �mV �eS �cK �yO �hZ �fP �mY �q^ �p^ �x^ �vY �re �}k �}t �wf �t` �y` �~z ��Z ׇo ��} ފy ��h �| ��r ��y ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ֋� � ě� ȝ� Ә� ۛ� 얉 矉 휌 ��� ��� 㠆 ��� 飔 ��� Ţ� ʢ� ̩� צ� ѭ� ˱� ӳ� ݸ� Ժ� ٻ� 歨 ��� ��� � �ī �ҭ �ƿ ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ���                       /1                                           >"",!                                         8$"$,,'8                                      /$$$$,,,+2                                   >"$$$%$,_,,,                                  8"$$%%%%,_,,,,<                              /"$$$%%%%..,._.,(8                            $$$$%%((%,._.,.ٚ(1                         :4""$$%%((+%...,.,�̝$3>                      1,"$$%%(+++%.,.._,��ق�;                     "."%%%(++++......,��̑���2                 =6
%$%(++++���....��̚�+�-1               8".%%++++�������.~.��̝̝��+!             0	
".$%(+++���������.._����̚��,           �
"""�$(++�����^�����.,����ʂ,,_-          
6�"$$.%+(�����KXo�������.�ٚ�̇,_,,          	��6($%6%�����IH���xz����ؗ���,,.,          	*���Ś$4����FJU�Ӫ���|�������Ś,_.�        �

����؝��ؘP?@@E��㫧������ٛ���̝,.�        �
�������?d@@@EE`կ����}���-����ٝ,6        �""*��̐̐(MdN@@EVYv��ӯ����[+�̐���ٗ4        �"$"̚��ڇ&?MdNNNffw֯Ө���pqF+��؝��ʑ.        .$(64���ڇ&MdNNfi�gMuӢ��I@GG&.���Ǒ˝�        *�*����܃%MdNdj�EMEg@aG@@P�\.����̔���       �	%(����܂&EGz���XEMEh``aYVFF&.�����̇��       %+6�����.%�捱�YEq�Ϡa?@E@Z.�����̑̚       %(+������_&b��@@tY϶VgEPgVF?������̚��      �%+(������.\��EfR�uugVOEFUG����������      �(++������.b��exj棯haQEE?�������ǝ��     �+-,����ٝ.Wb�������{eRE����̃��.��     �+,_-���̖.�s�����sYVSQ����ŀ.����     �,..-�̝,�,�'#m�����hYLE$������������     ,,..�������.�%"l�����UGD&�����������̃6     ,.,����������..+#]v�иl.��������ِ���Ǘ     ..._������������..$%kr\_�����������������     ...���������������_,	+,.������������������    .�����������������ڄ(	%-��������������������    ���̝��������������������������������������     ���������������������˛�������������������        �������������������������������������             ���������������������������������                 �����������������������������                     �������������������������                         ��������������������                               ��������������                                   ����������                                        ������                                            ��                        �����  ���?��  �����  �����  �� ��  ��  ��  ��  �  ��  ?�  ��  �  ��  �  ��  �  �   �  �    �  �      �    ?  �    ?  �    ?  �      �      �      �      �      �      �      �      �      �      �      �      �      �      �      �      �      �      �      �      �      �      �    ?  �    �  ��  �  ��  �  ��  �  �� ��  �����  ���?��  ������  (                �                         �  �   �� �   � � ��  ��� ���   �  �   �� �   � � ��  ���    p     GG     tdp   GGt�p  CGw�wV tw|x�t �|L��� xD��Ǉ xG��F���G��E��w�x�G�p��Dg������x��� ������   ����     �   �  �?  �  �  �  �  �  �  �  �  �  �  �  �  �  �  (       @                                  �  �   �� �   � � ��  ��� ���   �  �   �� �   � � ��  ���        tp             @t             @tGG           ttGGGp         @ttt         DGDtttww       tptpttGxtp     @t@tHwGxtw     @GCGG��twxtp   t4GG�x��x�G   wtDtx�L|��Ȅt   twwG��H�Ȉ�wG   t��w�DH���Ȉt�  tw��DD̎~|wx�p  Dwxt��~ww�H|�p  tH�DLH���GG�w�  CxxdG�lW��w��p  DxxTxG���DGxw�  t��DH�l|DDG���  GxwdFx���De��� DH�pE��D@V�w� w|w�dF��dgx�|� Dw��wDG�Ew��xw G�����dEh����� x�����tw��������������x������   ������x����    �����x����       ��������         ������           ����                     �����?�����������  ��  �  ?�  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  ?� �����������(   0   `         �                        �  �   �� �   � � ��  ��� ���   �  �   �� �   � � ��  ���            tp                     tG                    GG                   Dtttp                 t4GGGDp                G@tttw               tDtttttG@             4tCDttGwt            ptGCDtttt�tw           pDGDtptttx�Gp         Dt4GttGGGGw�tw        CCDG@GCx�GGH|�tp       pDDptttx��ttx��wG      D44tCGG����GG���t@     @tDGGDG��Dȏ�D�x�tt     Gt44ptx�|G|���x�wGG     GwDDtx��DLw̏��x�GG     Gx�wG��DD�Ό���x�ttp   @���x��DDȌ���xȈ�Gp   GHx�tD�DF���tw��tp   Dx�xtD�DLl�����XȌ�@   @Gx�GD����w���Dx�x��   wt��tD�Lh��ǄDGHx|�p   DG��eD�ǌdLlD�tw��w�   HxxVDl��LF\ld�Hxx|w   GH��DDxȌG��DDGH����   tx��GF�Dć���DDwxx|�   w@xxxD�D�||DF�D|�x��   ttxxxtFH����lDD@w���x�  ttx��tF����\DD|��|W�  ttG��GD̈�|llDw�|w��  ttww�G@egx��tE@vV|�W�p  GG||x�udD����DgW�Vx�P  ttwx���GVEȇtGV�����xp  GGx�����G@d�Ge��������  tt�������G@VT���������  G���xx����FT���������  ��x��������x����������  ���������w����������   ����������x�����x�      ����������x�����        �����Ȉx������          �x��������x�            ����������               ��x�����                 �����                    ���                      �            �����  ���?��  �����  �����  �� ��  ��  ��  ��  �  ��  ?�  ��  �  ��  �  ��  �  �   �  �    �  �      �    ?  �    ?  �    ?  �      �      �      �      �      �      �      �      �      �      �      �      �      �      �      �      �      �      �      �      �      �      �    ?  �    �  ��  �  ��  �  ��  �  �� ��  �����  ���?��  ������                                                                                                                                                                                                                                                                                                              