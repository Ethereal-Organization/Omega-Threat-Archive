MZ�       ��  �       @                                   �   � �	�!�L�!This program cannot be run in DOS mode.
$       ���ޥ�����������d�������|���������������Ŷ��������������;���������������&���������ƍ������ύ����Rich����        PE  L �ETG        �  6       �      P   @                     DS                                      Dc x    @ D                                                                           P                           .text   �5     6                   `.rdata  �m   P      :             @  @.data   �r  �  t  Z             @  �.rsrc   D   @     �             @  @                                                                                                                                                                                                                                                                                                                                                                                        ��$|  ��$�  �5��F ��$h  ��$\  ��$x  ��$l  ��$�  �t�F ��$�  ��$t  �=��F �50�F �@�F �-��F ��$p  ��$�  ��$|  ��$h  ��$t  ��$�  �5<�F �T  �=��F ���  �=�F �5��F ��  ���  �u �5��F +=��F �=D�F ��x  �D�F ���  ����  ���F ��$�  �$�  �$�  �P��$l  ��$�  ���F �=(�F ��$p  �-��F ��$d  �`�F ��$�  ���F ��$p  Y��$�  ��$|  ��$p  ��$d  �;���  �U ���F ���  �4�F ���F ���  �5H�F ��  ���9  �5`�F ��$|  ��$d  ���F �����$�  �$x  �$x  ����F �=��F �p�F ��    �=��F ���F ��$`  �8�F ;t�F �z6 ��F ��$�  ��$�  ��$x  ��$p  �=�F �-t�F ��$t  Q�P�F �-@�F �5��F ��$h  �Q  ��$�  ��=��F �=��F ���  ����  ���  +} 9���  �<�    �`�F �8�F ;�$  �n�  �0�F ���  ���  �5��F Z�5(�F ���F �������] ǅl      ��t  ��l  ��  ����  ���F ���F �5H�F �5��F 5h�F 5h�F ��5��F ���  ��t  ��$t  �5��F �(�F ���F ���  �U �4�F ���  ��l  ��t  �8�F ;�$  �U�  ������h  � �F ��t  �D�F ��  ��$H  ���  G���  +t�F @���F �t�F ��p  ��l  �=��F ��H  �5��F ��H  ��P���F ���F �5t�F ���p�F ���F ���QB �5��F ��	  Í��F ���F ��F ���  ����  �d�F +�$�  ;��F �  ��    �8�F 9��4, �=��F ��t  ���  ���F �=<�F ���F ���F 3=��F �=�F ��p  � �F �%��F ����F ���F ���F �<�F ���F ���F �$  ��F �5�F ���l�F ���F ���QB �5��F P��$p  ��QB �L�F ��$�  �x�F ��$d  ��F �-H�F ��$|  ���F �L�F ��$x  �H�F �-4�F �=��F ���F �`�F �x�F �(�F ��������W�=��F �=�F +=��F ǅ      ���  �8�F �J<ыQ|�yx=8�F ����  ���  �5��F �O�w���F �O���  �W 8�F ���  �O$8�F ���F �_8�F ��F    ��� ���  ���������F d�    �d�    �5��F �X�F 3��  ���  %�m=���  ���F ӆ�  ��  +�  ��H  ��@  �$�F ��\  ���F #��F ��8  ӆ  h�  �V!  �8�F �J<ыQ|���F �Ix8�F ����������F ���F �A�t�F �Q�i�=(�F �y =8�F U�i$-8�F ��$  �I8�F ���F    ���  �-L�F �������F ��l  �G����8�F ���  ���F ��  �t�F X���F ���  �5(�F V���  ���F ��������5�F �5�F �D�F ���  ��F @)�F ��F �5�F ����F ��t  �-H�F �H�F �0�F ��$�  ��$l  �`�F ���F �=L�F �5�F ��$�  ��$�  ��$�  ����F R�������  ���F ���  ���  ��  �t�F X���  ���  �(�F S���  ���F ��������p  �p�F �É�h  � �F �5p�F �p�F ���  ��t  ������=��F ��$�  ��$X  ��$�  ��$\  ��$�  ��$l  �����F ���F ���F ������T  ��h  ���  ��t  �z����5��F ��$t  ��$|  ��$�  �0�F R�=X�F ��$l  ��$�  ��$x  �-��F ��$�  �=��F �t�F �<�F �\$�-��F ��$|  �@�F ��$p  Q�5��F ��$�  �   �5��F �5��F 5h�F 5h�F ����  ��l  ��F �5��F ��p  �5H�F �<�F ���  ��p  ��l  ���F ��F ��p  ���F ������5��F P��F ��QB � ���  ��h  �5��F �����������h  ��$�  �@�F ��$`  �X�F �-��F ���F ��$�  ��$�  ��$x  �5��F ��$`  ���F ���F ������  ���  ��t  ���F ��F ���  ����=��F ǅ�      �8�F �J<ыQ|�Yx8�F ����	  �=��F �K�{���  �[���F    ��A�  �-��F ��$p  ����  �-��F )݉�$t  ���F �  ��t  � �F �<�F ���F ���F ���F 3��F ���F ���  � �F �%��F ����F �=��F ���F �<�F �=��F �,�F ���:���F � �F �%��F 35��F ���F     �5<�F ���F ���F �h�F �8�F �J<ыQ|�Yx8�F ��������K�k�{��$�  �K 8�F ��$�  �C$8�F ��F �S8�F ��$�     ���o ��$�  ����F ���F ���  �e  �<�F �5��F �   ��$x  �-��F ���F ��$�  ��$|  ��$�  �=�F ��$t  ��$l  ���F �5��F ���F ��$�  ��$p  ��$�  ��$|  �0�F �=��F �t�F ��$�  �4�������F ���F P�D$�\�F     �=\�F �=��F ������������F �5 �F F� �F +�$�  A����$�  ��d  �����F R��h  �5��F ����`  �����F ���QB h�  j�^���V��d  ���  ����F ��p  ���  ���F ��������$|  P��h  ��QB ��h  �=��F �p�F ��d  ��x  ��l  ���F ���  ���D�F ��F ��F ��=P�F ���  ���F ���F ��l  ��t  �ȉ��F ���  �5d�F ���  ��l  �,�F �T�F ���  �D�F ���i�������F ��F ���������F ��p  ��l  ���  ���  ���F ��������  ���  ����  ��x  )�;�$�  ������d�F ���F ��    ���  ���  �8�F ;��F �{! ���  ��t  ���  ��t  ���  ���{������  ��t  ���F ���  ���F �;������F ���F ��$t  ��$�  ��$x  ��$|  ��$d  ���F P�=0�F ��$p  ��F ��$�  ��F ���F �P�F [����������F �=X�F �=��F G)X�F �X�F �X�F �ы��  ��$t  �=8�F �5��F �(�F �=0�F �5��F ��$l  ��$�  �����F P�X�F ��$|  �3P��t  ���������p  ���F �ߋ��F �D  �@�F �T������5��F �5��F �7��QB �58�F P��$t  ��QB ��$l  �(�F �=0�F �5��F ���F ��$t  ����  �=��F �X�F �=0�F �  ���  ���  �$p  �$p  ���x�F ��$�  ���F �b  �L�E 3҅�u�\aB f�f�� w	f��t'��tf��"u	3Ʌ�����@@��f�� w
@@f�f��u����������������U��WV�u�M�}�����;�v;��|  ��   u������r)��$�,#@ �Ǻ   ��r����$�@"@ �$�<#@ ��$��"@ �P"@ |"@ �"@ #ъ��F�G�F���G������r���$�,#@ �I #ъ��F���G������r���$�,#@ �#ъ���������r���$�,#@ �I ##@ #@ #@  #@ �"@ �"@ �"@ �"@ �D��D��D��D��D��D��D���D���D��D��D���D���D���D����    ���$�,#@ ��<#@ D#@ P#@ d#@ �E^_�Ð���E^_�Ð���F�G�E^_�ÍI ���F�G�F�G�E^_�Ð�t1��|9���   u$������r����$��$@ �����$�x$@ �I �Ǻ   ��r��+��$��#@ �$��$@ ��#@  $@ ($@ �F#шG��������r�����$��$@ �I �F#шG�F���G������r�����$��$@ ��F#шG�F�G�F���G�������V�������$��$@ �I |$@ �$@ �$@ �$@ �$@ �$@ �$@ �$@ �D��D��D��D��D��D��D��D��D��D��D��D��D��D���    ���$��$@ ���$@ �$@ �$@ %@ �E^_�Ð�F�G�E^_�ÍI �F�G�F�G�E^_�Ð�F�G�F�G�F�G�E^_�����F     �8�F �J<ыQ|�Yx8�F ����   �=��F �K�{���  �K���F �C 8�F �=l�F �{$=8�F �T�F �C8�F �$�F    ��  �L�F ���F ��$�  �A$8�F ���F ��$�  ��$�  �I 8�F �߉��F ��$�  �-��F ����.�����p  �   �=��F ���F     �8�F �J<ыQ|�Yx8�F ����  �=��F �K�{�5��F �s���F �K 8�F ���  �C$8�F �k-8�F ��F    ����  ��$�  ���F ��	  �$�F ���F A�=��F �=|�F )�G�ǉ��F �=$�F �=��F ���F ���$�F S��p  �ȉ�l  ��󤉅h  ���F ���   ���F �,�    ��$�  �*8�F 9��� ���F ��$�  ���F ���F ����������� ���  ���F �4�F �$�F ���F ����  ���  +4�F ;�$�  �  ��    ���F ���F ���  �8�F ;��F ��� ��t  ��   ��$�  ��5��F �5��F ���  �5��F ���
  ���F ��$x  P��d  �l�F ��p  ��d  ���F �Љ5��F ���  ��l  ���F ���  ���m�5L�F �������$�  �R8�F ��$�  ��$x  ;�$x  �5�����$�  �A$8�F ���F ��$�  ��$�  �I 8�F �Z����g������F �f����-��F ����(	  U��QQSVWh  �p'G 3�VWf�=x)G ��QB �L�E ;ǉ5�%G tf98��u�ލE�P�E�PWS3��J   �}��E��x��P螤  ������u����&�E�P�E�PV��S�   �E���H��%G �5�%G 3�_^[��U��SVW�}���E3�9U��    �Et	�M�E�1j[f�8"u�}3Ʌ���j"Ë�Y����tf�f��f��f��t;��u�f�� tf��	u���tf�f� �e 3�f9��   f�f�� tf��	u���+���f9��   9Ut	�M�E�1�M�3�G3���Bf�8\t�f�8"u*��u#�} t�Hf�9"u���3�3�9Mj��[�M���t��tf�\ �M�Ju�f�f��t+�} uf�� tf��	t��t��tf��M���v�����tf�& �M��$����E;�_^[t��E� ]��5��F ���F ��$l  �=��F ��$l  �8��QB SP��$l  ��QB ��$d  ��$l  ���F ���F ��$�  ��$|  �\�F ��$t  ���������F �4�F C���F �4�F ��F )�A�ы��F �-�F �@�F ��$h  ���F �=��F �X�F ��$l  ��$p  �����F P��$�  �5��F �@�F �������F �4�F �=��F �d�F ��l  =��F =��F ��ȉ�h  �=��F ���F �������F �E؋t�F ��F ��3E�)D�F ���F ��h  +p�F �E���)��  ���  �]���   ��  3}�)��  �UԉL�F ��3U�)t�F �%��F �-��F ���F ��-��F ���r���F ��  ���F ��|  ���F P���  ��  Y�3��F ��@  ��P  ɉE���@  0�F Ɂ�4  �Sҁu������F ���F 3�F �-t�F �-t�F ��E� �F ��  3��F ���  ���  �F �}��=�F ��  0�F ��  ��HS��  S�Z�  ��Yu�����  �0�B ���B     ���  ����` �@ �@
�0�B ��$���  ;�r�UVW�D$P��QB f�|$F ��   �D$H����   �8�h�/�D$�   ;�|��9=��B }N�4�B S�ğ  ��Yt8���B  ����  ����` �@ �@
���$�;�r��9=��B |���=��B 3ۅ�~j�D$� ���tT�M ��tL��uP��PB ��t<�ˋÃ�������0�B �4��D$� ��E �F�Fh�  P�ke ��YYt.�F�D$CE;�|�3ۋ0�B �ۍ4��>�uo���F�u
j�X�����y��H������P� RB �����t?W��PB ��t4%�   ���>u�N@�	��u�N�Fh�  P��d ��YYt��F�
�N@��N�C���r����5��B ��QB 3�_^][��H�j �E�    �E�    �U�`�F �R� �F ���F �0�F �E    ���F ���F �= �F �M����F �]܋�   �3M�   ���E�   ��h  �ˉu�5��F �m�.���  �UЋt�F +��F �E�+��F �h�F ���F �M�1�1�I�$�F �Eԉ1�1�I��x   �E� ���F �E��M�]��=��F �5��F �$�F �U �M� �F �u��������5��F ��$�  �5�F ��$�  ����  ��$x  +�$�  ;5��F ��  ��$�  ��$�  �5��F ��$�  ��$�  �4/58�F 9���~  ��$t  �5��F �5��F �������l  ���@���3L$ ���M܉t�F ��)D�F ���F 3t�F )D�F �M܅�������E؋t�F ��F ��3E�)D�F ���F �D�F +p�F �8�F ��)t�F �uԉ=�F �h  ����F d�    �3d�5    ���  ���F ��  ���  50�F ��X  ���  ��X  X�F ���  ��  35(�F ���50�F j �?�  �ǅ�      �=8�F �O<��Q|�Yx����  �=��F �K�{���  �S���  �C 8�F �k$-8�F ��$x  �S8�F ���F    ��� ��$t  �
�  �0G ���F ǅX      �5�G ��G ��p  ��X  ;��F ��b  ��$�  �$�  �5�G ��T  ދ�$�  ��P  �(G     ��   �}���   ��  358�F )5t�F �8�F ���F ��3M�)t�F �=t�F +=��F �]�+��F �ÉMЋ8�F �uԋωD�F �]Ћ=�F �����5�F �5��F ��$t  ���������L  �%(G �����p  ��H  �5(G ;5��F �de  ��$�  ��G �0G �5�G �����ǅ�      ǅ�      ���F     � �T�F ��p  ��T  �0G ��P  ����j�����G �(G ��L  ���-(G (G �-�G A�G B��H  ��P  �T�F ��H  �0G ��D  ��T  �5`G �5(G �5�G ��H  ��   ���F ���  X���F ��1�)�$�  ���  ���  +�$|  ��l  ��)��  ��  3�$x  )��  ���F ��l  �l�F ��3�$�  )��F �5��F +�H  ��h  ��$�  ��$�  ��$�  ��F ��F ���$�  ��$l  �-��F ��$�  ���F �-L�F �O����(G �5`G �T�F �o������  +��F ��h  ���  �49�9�I�D�F ��d  ��`  �5l�F �49�9�I;|�F �M\ �5D�F ���  ���  ���F �5��F ���  ��p  �Q�  ���F �=��F �7V���  ��  17���F ���F CT��(  �a����(  ˍ=��F _T���F ���=��F ^�4>�]�������4�[S�]��j ���F     ���F �=��F    |Í5��F �=��F S�������;�������v��F ���F ���F ʍ��F �l�F �x�F +��F HTQ���F Ӡ0  ��0  3=��F ��  �ʁ�H  k�]�%��F j �E�    ��t�����t���   �!  ��x����]���5��F 13�[R���F ��F Ӫ�  ���  $�F ���  ����+L�F 3��F ���  �p�F BT���F �%��F ���  ��C�5��F 5��F P�$�F 4�F ��p  ӂ�  ��  ���  50�F �(�F ������F ���  �F Q�L�F ��F ��t  ��  +��F Z0�F �4�F ���F yT���  ��  ���  �-8�F �E����F �5  ��x����]���5��F 13�[�]��������  ���  ��  ��x  #��F 3��  ��8  ���  FT���  ��F ˉ��  ���  +��  �P�F ���  Ӧ8  +=t�F =0�F ��t  F�^T���  ��t  ȋ5��F +5�F ���F ���  ���Ӌ �F ӊ�  � �=G �=dG =`G 9���4 �=,G �=G ��G �58�F �5xG �0G �]̋]؉]Љu��5�G �;��F ��0 F�M��U��U����1 �0G �M��]̉5�G �M��,G �M��u�뤉�G ���F ��R�@�=��F ��<  ���G �H� ��G ��<  ��G �=�G �6  ��0  �}��HG ��	G ���  ���  ��0  ��G ��$0  ��G ��$�  ��$�  ��$  ��G �HG ��G �-�
G ��$0  �5�G �=�	G �  j �E�    ��h�����h���   ��   ���F �8�F W�}��17��H�F �P�F p�F ���F R�8�F +��  ��X  ���`���|�F �+�@  0�F �5<�F +5X�F �=(�F �e���G ���F ��G ǅ<      �`G ��w�����G ���F ���  �ǋ�G �r����8�F R�U��
12�R�U�Z����F��$�\G �G ��G ���  ��G ��S�5�G �\G ������XG �� ����\$ ����$   ��G �8G �-8G �dG �XG ��  ���   ��G �,G ���  Q��H  ��  ���  ��G ��G ��H  ��
G �5�	G �5`G ��G ��	G �΋,G �5�G ���{  �=��F �d�F �Ƌ �F �%h�F wT��<  ӯ�  ���  {���0�F ���  u�}iS���  ˋ��  3��F OT�t�F D�F GTQ���  �@�F �uS��  ��  �lG �=G ��  �=�G �G ���  Q��G ���  ��G �������  ǅ����|g �58G ��,V�G �	  F�,����,�F     �T�F 	   �T�F �n� ��\������F �,�F �8���F S�,�F 1�[�,�F �$�F ���F [뷉�G ��[�@P��G Y�S��G ��[�A�5lG ��t��(  �����   ��   ������7  �D��������  �f��������   ��  F�   ��G �5�G � G ��G     �DG ��G ��G ��  ��������  ���  ��G ��G �=�G ǅ����|g ��  �=�G �=|G �58G ��4V�  F����=8G W�lG    ������S�΋�G �������$   �-|G �pG ��G �
�R�A��G �pG �D  S�5�G �������Y��G ��G �lG [�[��$   �|G �-�G �M �m�A�-�G �-�G ��$  ��$   �-�G �5�G �\$���$  ɉ=�G ��$   ��<  ��$�  ��=�G ��$�  �  ��$  �-�G �-�G �.  Y�|$��G ��$   ��G ��G �5�G �t$���$   ��G �-�G �-�G �����  UV�5�)G W3�3�;�u����   f== tGV���  Y�tFf�f;�u��   SP�|�  ��;�Y��%G u����\�5�)G �/V��  ��Gf�>=Yt�?P�I�  ;�Y�t9VP���  YY���4~f9.u��5�)G ��  �-�)G �+��B    3�Y[_^]��5�%G ��  �-�%G �����P�-|G �5�G �tG U�l$��Y  ��G R�,G �\$��G �`G �D$��G ��Z��$<  ��G �-`G ��  �	  ��$  �`G �tG X��G �=hG ��=tG �|$���G ��R�@��G �=hG �5�G �`G �@����|$�����   �  �G ��G ��G ���  ��G �Ӌ�G ��   �������  ǅH     ��   ��G �-�G �XG ��$   ��G ��$  �8G ��G �50�F h�  jd�5��F �5��F �p  �S	�PG ��G j��G R��G �T$��G ��G ��$H  ��G Z���l��	��G j��G �5�G W��G �|$��$H  �=�G _���6��  ���   ��  �-|G �{  �<G 	�X��$0  ��G    ��$  S�-�G �5�G ��G ��$  �|G ������TG ��$  �-�G �5�G [�-TG ���������$   �-|G �5�G �H�����$0  ��   ��   ����7  �H������   ��  �%�����   ��  �|G �-|G �   ��$d  �-`G �5�G �=G �|$(��0�S  QǅH      ���  ��G �LG ���  ��G �LG ��G �=�G �5�G ��H  �=�G ��G �=�	G ��G �=�G ���p  �-|G �5�G E�-|G �5�G E��$   �-|G ���*�|G �$G �$G ��G �S  �$G ��� ��   �|G ��  Q��0  �|G ��G �dG ��0  �=�G _�=�G �=�G ��   ��G �|G Q���  ���  ��	G ��G ^������5(G �������	G �5�G �5�	G �5�G ���z  �G �-�G �|$Y��$  ��G �-�G �5�G �@G �t$���$  ��G ��G �G �����,�=�G �5dG �=|G �5�G �I����� �}��|G �=�G W+=�G �=G ����G �=�G ��  ��G �-LG ��G ��$4  �=�G ��$  ��G ��$�  ��$�  ��G ��G V�5G ��G ��G ��G ��G �  ��G �ҋG �������G �=�G ��
G ��G ��  ��G ��G ��  ��G �5�G ��4��	G �lG ��G ��G �G ��	G ����   ��$�  �|G �=�G ��$�  �-|G �5�G ��v�A�5�G �5�G �?�����$������G ��G ���  ��H  �҉�G V�����������G �� ����\$ ����$   ��G �8G �-8G �dG �������   �|G ��  ��G R��H  �-�G �dG ��$  ��������S�5G �=�G ��H  ��	G �5�G ���  ��G ��G ��G ��  ��  ���  ���  ��	G ���  ��G [�=�G ��H  �5G ��G ��G ��G ��  �D$��$  �-G �G ��$@  �`G �G X��$  ��$  X������   �  ��G �`G ��$8  P��G � ��G �@P�-|G �5�G �D$�,G Y��
  �DG ����G �5DG ��$<  �5�G �  �0G ��G     ���  ��G S���  ��G [��G �=G �5�G ��G �=0G �=�	G �=G �b�����$  ��G Y�|G P��$<  ��=�G ��G �=�G �=,G �5�G ��R�@�=�G �5�G �X  �G ��G �ҋ�  �=�G � G ��G �5�G ��	G ��H  �5<G ��4�������G ���hG �5�G Z�D$���$   ���  ��$�  ��G ��G �΋-hG ��$  �-(
G ��$�  �=�G ��$  �|G ��   ��G ��G ��G ����$  V�� ��$�  ��$  �5�G ��$�  ��$�  �=�G �(
G �-|G Z��$�  �=|G �-�G �=|G ���"  ������-�G �5G ��$  �-|G �5�G Q��$  �T$�=�G ��$  �=�G �=�G �=�G �΋-LG Z�5�G ����  ��G �t$��=�G �=�G ��$�  ��G ��$�  �|G �@G S��G ��$  �-�G �� ��$�  �ߋ-�G ��$�  �։�$�  �=�G ]�(
G �5�G �-|G �-@G �e  ��$  ��$   ��|G �(
G �5,G �5�G ��G ��R�@�ȋt$�=�G X�  ����$  �G    R��$  �-G �5�G Q�-|G ��$8  ��$  ��$  ��*���P�G �`G ��$<  �G �1���X�� ����|G �=�G �� ������  �� �����  ��G ��G ���  ��G �������  ��	G ��G �5�G ��G ��	G �������G [�=�G ��G ��H  �5G ��G �5�G �G ��G ��G �8G P��H  ��G �=�G ���@�4G �8G �=�G �  ����H  ��G    ��   ��   ��  P��H  ��G �G ��   ��   V��G �5G ��  ��$  �5|G ��j���P��$<  �`G �$<  �t$�����7  �%G U3�;�V�5tQB u-�օ�t�%G    � ��QB ��xu�%G    �3��\��u���S��u�SW��QB �=`QB UUj���SjU�׋�;�t&�6P�X  ���YtVUj�Sjj �ׅ�uU�   Y3����_[^]�jh0RB ��  �u��tX�=,�E u@j��B Y�e� V规  Y�E��t	VP�Ä  YY�M���   �}� u�u�
j��A Y�Vj �5�E ��QB �\�  Ë�G ��G P��G Q���  �5�G �^�  ��G ��  S�������%  S�=0G ��G �����_��G ��  ��G �=�G �4G 럃�,�G �lG ��  ���  ��H  �֋�   �������  ǅ     ��  ��  �5lG �-lG Q��$   ��$(  �D$(��$  �  ����   j��   ��G �4G P������G X������G S��G ��$�  ��$  �� ��$   ��G ����$�  ��Y�-�G ��$�  �|G �(
G ���  ��G �=�G V�N �=0G �5�G ��  S��G ��   ��G ��P������������G X�-�G �C  ��$  �-|G ��$<  ��G ��R�@P��G �-|G �,G �5�G �#����D$��$  �͉0G ��G S�,G ��G �0G �D$Z��$  �dG �D$��$@  �����I�����G ��G [�=0G ��G �
�R�A��G ����G ������hG ��$  �=�G ��$�  ��$�  �t$��G ��G ��G ��$0  ��$�  ��$   �|G ��G ���  �-�G �E ��G ��$�  ��$�  �(
G h�  ��  �-LG ��G �5�G ��$�  ��G Q��$  ��$�  ��$�  ���  ��$  ��$�  �5�G ��� Y��G �=0G ��$   ��l  W�5�G ���  �=0G _��6  �5�G ��$0  �=0G ��$0  �1  �$G �-�	G �΋5$G ���5  �-�G �PG �8G ��$  ��$  �ы�$  �-G �5`G ���������G �=�G V�H �=0G �5�G ��  �G ��G ���	  �lG ��P�G �������G X�-lG �  �vP��������� ��G ��  Z�5|G �dG ��  [��G ��G ��������G �=G �=�G ��  �dG ��G �=G �|G �w��$0  �=0G ��$0  ��G ��G � ��G �@��$  ��G ��$  �O�����$  ��G ��G �5�G ��v�A�5�G �5�G �������   ����  P�΋D$��$  ��!�����$   ��$  R��(
G �5,G ��G �5�G Y�|G X�t$�=�G ��$�  �4������� ��$�  ���%�G  ���	�G �-�G �/G� ��G �5�G ��$  �� ��$  ��j� G     Z�D$��\G � G �\G �D$�������  ]� ���̋L$W����   VS�ًt$��   �|$u����   �'��������t+��t/��   u����ua��t��������t7��u�D$[^_���   t�������   ��   u����ut�����u�[^�D$_É����t�����~�Ѓ��3��� �t܄�t,��t��  � t��   �uĉ�����  �����   ��3҉��3���t3������u����w����D$[^_ËG ӄ$0  �ՋG �5�G 󤋜$$  �G ��$  ��G ��$(  �=�G �|G �G ��$T  ��$  ��$(  ��G ��$  ��G �=�G �Չ5<G ��$(  ��$�������G ��  ��  I�xG ��H  ��  ��  �|G ��� P��  �|G B��G W�=4G )ω=�G �G �=4G ��G ���  ��  ���  �D$�|g ��G �D$��G �-�G R��$   ��$4  �58G ��(�t$ �G �����=�G �=0G �5�G �.�v�E�5�G ��$   �� ���\G    �\G     �5�G �\G �|G P��   ���  �,G �5�G �|G X��G �\G �I���  � G �G ��G �,G ��   ��0  ��G �=G � G �=\G �\G ��0  ��G �d�����G Q�������������G ��G �BR�������G ]����  �lG Y�5lG ��$  �$  ���   �-�	G ��$  ��� ���	�GW��$<  �@G ��$  �΋�$�  ��$�  ��G �@G _��$8  �5�G ��������$4  ��G �|G ��$  ��$  �$   ���   ��G ���a�����$   ��$�  ��G �΋=hG ��$  �=(
G ��$�  �-�G ��G ��R�@�=�G ��$  �ȋ|G �t$���G �2���������4G �\G �X�v�A���|G ��0  �5�G �|G �E���  �\G �I��  ��0  �\G �\G ��   �5�G ��  ����U��� SV�u�^��ud�   �E�E�H;ىM�r;Xs3���  W�~���u3�@��  3҉U�Ë���t;��E  �x t�EB��;�v��} t�F�;E��"  ;��  ��$G ���� ���3���~9<��$G ��   F;�|�j�E�PS�|QB ���`  �}�   �S  �E��tV�M�f�9MZ�?  �A<��8PE  �.  f�x�"  +�f�x �H�L�  �A;�r�Q�;�s�A'�uwjh %G ��QB ���������$G �ɋ�~���$G 98tJ������u-j[;���3҅�|���$G �0B;Ӊ8��~��}A��$G j h %G ��QB ����3�����������QB jh %G �Ӆ��z���9<��$G t.��$G �p���|9<��$G tNy��}��}@��$G �p��t3Ʌ�|���$G �A;Ή8��~�j h %G ���������_^[�É�G �5�G ��$  �U� ��$  ����G    �TG     �-�G �TG �-\G �\G ��������S�������G �5�G ��G �BR��G ]�|�������G �G �G ����  ��G ���  ���  �����  ���  �tG ��G ���  ���  ���  ���  ���  � G ���  �-�G �E % ���(
G �E E�
�R�A�5�F �b����U��WV�u�M�}�����;�v;��|  ��   u������r)��$�,_@ �Ǻ   ��r����$�@^@ �$�<_@ ��$��^@ �P^@ |^@ �^@ #ъ��F�G�F���G������r���$�,_@ �I #ъ��F���G������r���$�,_@ �#ъ���������r���$�,_@ �I #_@ _@ _@  _@ �^@ �^@ �^@ �^@ �D��D��D��D��D��D��D���D���D��D��D���D���D���D����    ���$�,_@ ��<_@ D_@ P_@ d_@ �E^_�Ð���E^_�Ð���F�G�E^_�ÍI ���F�G�F�G�E^_�Ð�t1��|9���   u$������r����$��`@ �����$�x`@ �I �Ǻ   ��r��+��$��_@ �$��`@ ��_@  `@ (`@ �F#шG��������r�����$��`@ �I �F#шG�F���G������r�����$��`@ ��F#шG�F�G�F���G�������V�������$��`@ �I |`@ �`@ �`@ �`@ �`@ �`@ �`@ �`@ �D��D��D��D��D��D��D��D��D��D��D��D��D��D���    ���$��`@ ���`@ �`@ �`@ a@ �E^_�Ð�F�G�E^_�ÍI �F�G�F�G�E^_�Ð�F�G�F�G�F�G�E^_���PG     ���F �-�G �DG �-XG ��$�  ��G �=�G ��$�  ��$�  �=�G �   ���$�  ��$�  �    ��0� ��$�  � ��$�  +�$�  ;�G ���  ��G ��$�  �-G �5HG �   ��G ���F ��  �5�F �F<��p|��   �Xx�F ���;�  �C�=�G �{�k��$�  �{ =�F ��$�  �S$�F ��G �C�F ��$�  ��$�  �������$�  �Ћ���-G ���G �$�  �$�  ����  ��G �%�G ���  ��G �dG ���  ���  �5�G ��F ;�$�  ��g  �  Q��G �� G �h�F ���F �5��F �| G ���  ���F �5��F ��l  ���  ���F ǁ�      � �5HG �����] �K$�$�  �<G �G �E �@ �$�  ��<  ��G ����  ���  +lG ;U���  �|G ���F �A  ��$  Ǆ$�      ��$�  �-�G ��8���`�Q  � ����U�D$��tJ�T$VW��|$׃�t8�   t�:uX������t��8�uE�N�W8�u;������u�_^Ëȃ���t+�t'�N��W�8�u8�u����8�u8��    �_���^Å�tċ�8�u��t8�uރ�t��  � ��  � ;�uɃ�_^��������̋T$�L$��tO3��D$W����r1�ك�t+ш����u������������ʃ���t��t
�����u��D$_ËD$Á��   �[�PG �=PG    �G�  ���  �=�G �-G ��$�  �G �5�G ��$�  ��$�  �5HG �G �G ��$�  ��4  �m��$�  �=�G ��G ��$�  �5G ��$�  �G �����@G ���  ���   �C�����G ��G �J  ���  �=|G �G �  ���t  �%|G S�|G �3�$�  ;U �x� ��<  ���F �=PG ��G �<G �G �=�G ��G �� G ��<  �h�F ���M���h�F �5��F ���  �h�F �5��F �h�F �h�F ���  �h�F �=PG �| G ���  ����T�}  ��G �5G �  ��h  ��<  ���  �=4G ���=������  �5�G �5��F �7��QB ��$�  P���  ���F ���  �`G ���  ���  �����   ������tG ��,	  ���  %��  �G +�$  ;�$�  ��  ��    ��$�  9��̩ ���  �tG ��G ����d�  ��G ��G ���P  �h�F � G ��$�  �G �=�G ��$�  ��G �=| G �t$<��$�  ��$�  ��$�  ��$�  ��$�  ��$�  �ӋG �  �<�F �5(G F���(G ��G )�C�É��  ���  �54G �<�F ��G �<�F ��R���  �ȋ��  ���  ���@G ���F �  �5��F ��G     ���  �J<ыQ|�Yx�$�  ���e
  �5��F �K�k�sP�C �$�  �=xG �{$�$�  ��G �C�$�  �`�F    ��f�  ��$�  �)  ���F �h�F ���5�F ��������  �J<ыQ|�Yx�$�  ����  �K�s�kR�S �$�  ��$�  �{$�$�  ��$�  �S�$�  ���F    ��0t ��$�  ��$�  �   ���  ���  ��G ���  �-8G ��$�  �,G �=�G �-�G ��$�  �=�G ��$�  ��$�  ���h�F �L$̃�4�h�F �5��F ��G �h�F �5��F ��$�  �}�����G �� G j�k���É�h�F ��$�  P�G ��QB �G �5G ���  ���  �G ���  �G �54G ���  ���  ��������=��F �=xG ����  ��$�  )�9���  ��$�  ��$�  ��$�  ��$�  ��$�  ��$�  9����  ����G ���`��  �5T	G �5��F ��8  �$�  �$�  ����  ���  ��8  ���  ���  ��|  ��G ���  ��G �  ��D  �  ��$�  �5PG F�ȉ��  �=PG ���  )�G�ǋ��  �`G ���  ���  ���  �����  R��G �ȋ5�G ����G ���������G �$�  �$�  ��5hG �G ��$�  �TG ��$�  ��$�  ��G �G ��$�  �=G �TG ���z����5�G ���  ���  ��<G �G ���  ��T������QB ��G �U ���  ��<  �5�G ���  ���  ���  �=8�F �58G �lG ���  �5�G �DG �E ���  ���  �5lG �=�G �<G ��G �u���<  ���  ���  �5G �=�G �PG �-4G ��$�  ������  ��XG �`�F ��G ����  ���  )�;XG ��  ��G ���F ��    ���  ��G ��$�  ;�$�  ��� ���  ���F �E�   ��F ��R����G ���F P�� G ���F �58�F jB��G ���F P�� G ���F h|#  jB���  ��  P��  ���F ��H  C����G ��H  ��D  )�B�-$G ��G ��$�  �=\G ��G �=��F �=�G �5G ���5��F V��$�  �Z  �߉�$�  �T$��$�  ��G U��$�  ��$�  �D$ ��$�  ��$�  �HG ��G �\$�5�G ��G �=�G �D$��G ��$�  �58G �� G �=�G �=�G ��G ��$�  �[X�\$���$�  -0�F �-pG �-	G �Ӌ�$�  ��G �D$��͋pG ��$�  �Ӌ��h�8  ���  Z��d�#�����G �5� G �=| G ��$�  ��G ��$�  ��G ������  ���  �[ �$�  �=TG �=�G ���  ��G �G )�R��G �R���  ��G �I9��%�  �3  �� G �ȍ��F ���  j� 	G ���F P�� G ���F �5�G j���  ���F P�� G ���  ʋ�G �5�G P���  �} �`G �-pG ��G �5�G ��$�  �G �=�G � 	G ��$�  ��$�  ��$�  �=xG �5(G �`G �5�G ��$�  ��0�F �9�����G Z��$�  ���`�  ��P�G ���  ����P������l  Y�I�$�  ���F ��d  �E����F ��`  ����  ��X  +�$�  ;U��y  �5  ��G �<G �5� G �=| G ���  ��G Y���  ��G ��P�����-G ��8�F  G  G �1��G �=�G ��G �G S���  �Ƌ=$G ��G �� G ��$�  ��G �=G �5<G ��  ��G     ���  �K<ًQ|�Yx�$�  ���a����5��F �K�s�kR�S �$�  ��$�  �S$�$�  ��G �S�$�  ��F    ��Р  �- G ��$�  ����F �����5�G �=�G �� G �G �=8G ��$�  ��$�  ��$�  �G �|$��G ��G �5� G ��$�  �D$��$�  ��G �0G �Ë=| G ��$�  ]��$�  ������9����E�   ��F ��Q����G ���F P�� G ���F ��\  jB���  ���F P�� G ���F h|#  jB��d  ��  P�� G j
S�5��F V�  P���  �@<�$�  �X|�px�$�  ���l�  �5�G �5��F �4�F    ����  ��X  ��X  %��  ���  �-�G �E$�$�  �m�$�  ��$�  ������T  ��X  �u��p�F ����  W��G �LG ��    �=TG ��G �T$�(�$   ;�G �n� �0G ��G �#�  ���F �@�F �TG �P	G C)TG �TG �TG �ȉdG ���  ��G �5@�F ���  ���  ���@�F P�TG ���  �=tG ���lG �  �=�G ��$�  =�G =�G �R��$�  �=�G �\$��-�G ��$�  �5,	G ��G ��G �|$���$�  �5�G ��G �5TG ��$�  �������G ���  �TG �#������  �=@G �� G ���  �=G ���  ���  �5G ��G �� G �@G ���  ���  ������    �
�$�  9��E�  �<G +�G ���  50�F ���F @G V�5� G �L G ���  ���  ���  ���  ���  ��G �։=lG ���  �=� G �-pG �=�G ���F ��j �n  Ë��F ����  �h�F �5dG P�XG ��QB �XG ���  �=tG �G ���  ���  ���  �TG ��������ȋ�$�  �5�G ��$�  �=��F �4G ��$�  �9��$�  �h�F ��$�  P��$�  ���F ��$�  �5G ��G �DG �=\G ��$�  ��$�  �DG ���������  ���  Z�tG ��d������D  ��`  ��   ���F �%��F ���F �TG ���F ��$�  ;E��l�  �� G �U���`  �� G ���F �TG �  S�hG ���F �h�F �֋=lG �݋��F �� G ��$�  ���F �G �� G �(G ��$�  ��$�  ��$�  ��G �����L��  �X�F ���F B���F +�$�  A����$�  ��G ��L  �5�G �TG ��T  ��H  �5X�F �5� G ��`  ���=X�F V��G ��P  ��)  �5�G �p�F �tG �u����F ���  ��G �=8�F = G = G ���G P�� G ��$�  �=�G �d$ ��G �|$V��$�  ��G �L$�1�$�  ;�$�  ��z ��$�  ��$�  ��$�  �5�G W��G �\$ �-�G �����5$G S�5x G �( G �5@G ���U���4�    ��l  �� G ��G ��$�  ;x G �i� �� G �� G �� G �M���5@G �5��F j ���  �K<ًY|�qx�$�  ����  P���F �F�NP�F���F �V �$�  V�v$�$�  ���F    ����  �8G ���F �������  =0�F ���  ���F @G �=, G W���  ���  �H�F ���  ���F ���  �L G �5�G �׋, G ��G ���  �H�F ���  �5pG ���F �x  ��D  �=� G ���F ��h�F ��$�  P��@  ��QB ��L  ��@  ��<  ��`  ��T  ��X  �5�G �=G ��`  ��H  �TG ���  ����$  R��$�  ��$�  ��󤉼$�  ���F ��h�F ��$�  P�G ���F �G ��$�  ��$�  ��$�  �=(�F �L$��$�  ��$�  �����P������ ����������̍B�[Í�$    �d$ 3��D$S�����T$��   t�
��8�tτ�tQ��   u��W����V؋
����~����3���������3�3ƃ��� �u% �t�% u��   �u�^_[3�ËB�8�t6��t�8�t'��t���8�t��t�8�t��t��^_�B�[ÍB�^_[ÍB�^_[ÍB�^_[�V�t$��tV��  @P��P  ��YYtVP��  YY^�3�^Ép�F ���F ���F     ���  �K<ًY|�qx�$�  ��������NV�n�v��$<     ��g9 ��$�  �쉽�  �5lG ^�v�$�  �M����  ���������`  ���F 놉�$�  ��$�  Z��$�  ��$�  ���`�N����5@G �( G ���;���Y��G �-�G �0G �-�G ��G �D$�0G ��$�  �������E���d  �t G ��P  ���F ��T  �@ G �8G Ƌ@G Ɖ�d  ��ЋhG ��L  ��X  ��T  �E��.�����`  �H G ��d  �g����5tG ��G ��$�  ��$�  �=�G �L�F ��$x  ��G W��$�  ��$�  ��$�  �=pG �5�G ��$�  �5HG ���F ��4�T$ �hG ���F �h�F �4G ��G ��G �L�F �=L�F �-��F �5��F ��$�  ��$�  ��$�  ��$�  �5��F ��$�  ��G ��$�  �4G �t$4�D$4��$�  ��$�  ��$�  h(#  �5��F h�  h�  �E  ËE���`  ��l  �G �G ����G ��X  ��l  �=\G �pG �U�_��G �=x G ��`  �E��=\G �������  ���  ��H�r  ��G ��$�  ��G ��$�  ��$�  �pG ���F �(G ��$�  �-�G ��$�  �/�$  ;�$�  ���  � ��4R�hG ���F �h�F ��G ���F ��G �5��F ���  �� G ���F ���  ��G ��G �pG �(G ��4��H�E  jh RB �O�  �u�u�u���uF3��}���we�=,�E uG������u�]�;D*G w3j�z Y!}�S�+Z  Y�E�M���J   �}��t�u�j W�Y�������u:Vj�5�E �RB ����u%9=�$G tV��o  Y���v�����uj�] YË����  �;(3E u��    jh�RB ��  �e� j j��  YY�3�@Ëe�M��j�RB ̋F�$�  ���F    ����  ��G �E��5x G �5��F �5� G ����  V+u�;5�G �r�������U����(3E ��t=N�@�uNV�E�P�RB �u�3u���QB 3��<QB 3��(QB 3��E�P�HQB �E�3E�3��5(3E u
�(3E N�@�^�����U��SVWUj j h��@ �u�� ]_^[��]ËL$�A   �   t�D$�T$��   �SVW�D$Pj�h��@ d�5    d�%    �D$ �X�p���t.;t$$t(�4v���L$�H�|� uh  �D��@   �T���d�    ��_^[�3�d�    �y��@ u�Q�R9Qu�   �SQ�3E �
SQ�3E �M�K�C�kY[� �5��F �5<G +5�G ���F ��l  0�F ��G ���F @G �pG ���F �hG ӂ�  ��  ��Q��G ���  ���F ��G �L G     ���  ��\  ��d  j�5��F �5�F hX  �   ���  �N<�Y|�qx�$�  �������P���F �F�N�D G �N�( G �^ �$�  Q�N$�$�  ��G �Y���^��4���L뙉pG �-(G ��$�  ���F     �-��F �-L G ��,���L�c�����`  ���  �5(G ��\  ��X  � ��$�  ��G ���F ��$�  ����  ���F ���  C���  +�G B�ʋ�G �5��F �ʉ��  �5�G �=��F 󤉍�  �=dG ���F ����  �8G �h�F SP� G �������j�58�F h�  �x����Q�T$��$�  ��G ��G �-XG �=| G �L$��$X  �<G �-� G �=�G �-G [�5,G ��G �-XG �-PG ������끋�$�  �-$G ��$�  ��$�  ���F �-�G ����   Y��$H  ��$�  � G ��G �5 G ����'�����$�  ��G �$�  �$�  �Q�-�G ��$�  �G ��G �=0G ��G �5tG �D$��$�  ��$�  �G [�pG ��$�  �HG �  ��$�  ��$�  �=�G ���F �5��F j
j ����V��$�  �=PG �4�F ��$�  �(G �-�G ��$�  ��$�  ��$�  �HG ��$�  ��$�  �5�G �pG ���F �-X G ��$�  ��G �=L G ��$�  �4�F ��$�  ��$�  ��������  ���F ���  ��H������G ��$�  �tG �5��F ��V�hG ���F �h�F ��G ���F ��$�  �5G �tG �$G ���F ��$�  �4G ��$�  �݉(G �����L�������$�  ��G �5��F ��$�  �(G ��$�  ��$�  ��G ��$�  �$�  �$�  �jd�5��F �F���Ã��=�����l  ���F �   �<G +�G ���  50�F ���F @G �50G Vǅ�      �G ���  ���  �G ���  ��G �֋0G ���  �-G ��G �=L G �-pG ��$�  �݋G �w�����$   �5H G ��`  F�H G +�G C��$�  ��G ��L  ��X  ��G ��H  ��l  ��$�  ��G ��$   �-� G �P�F �=(�F ��������F ���QB ��$  P� G ���F ��$  �|$p�dG ��$  �5�G ��$�  ��$�  �5�G ��G ��$   ��$  ��$  ��$�  ���F �-xG ��$  ��$  ���F �=t�F �� G ��$�  ��G �5HG �=�G �|$p��$  ��$�  ��$�  ��$  ��<�h������  �=xG X��d�����ȉ�$L  ��$�  S�=�G �-<G � G �=<G �-| G �-�G �5,G ]��G ��G �<G �-�G �� G �PG �G ��G � G ���W����i����hG ���  X�=xG ��d�����Q��$�  ��$�  ��$�  �5�G �ȉ�$�  �l$��$�  �5�G ��$�  �=�G ��$�  �dG ��$�  _�� G ^�|G �TG �-�G �=@�F ���F �   �8�F  G  G ���    ���  ���h�F P�� G ���  �h�F �5��F �G �h�F �5��F �� G �h�F ���  ���  ���  ��$�  ;�$�  �ca ���  Q�8����5tG ��$�  ��$�  ��$�  �|G ��$�  ��G �5�G �pG �-�G ��$�  �dG ��P��  �5��F j��`  ���F P�� G ���F �5�G j��4  ���F P�� G ���F ��\  ΋�`  ��L  JT��X  �pG JT��G     ��T  ��X  ��P  ��G � �@�F �=��F �tG ��$�  ��$�  Y�=�G �5�G �pG �-�G ��$�  �dG ��L��   �|�F ��$(  G��$(  +@�F B�ʋ@�F �5|�F �ʉ�$   �5@�F ��$  �=|�F �xG ��G �-t�F ��$  ���F ��$�  �����\G S��$�  ��$�  �=�G ��$�  �L$��$�  �D$�-�G �=�G ��$�  ��$�  �5�G ��G ��$�  �dG �\G �=� G Y��$�  ��G �-TG ����j �5t�F �5��F �5�F j ������j@h�TB 菽  �(3E �E�3�3�F9=%G u2V��TB PVPWW�QB ��t�5%G ���QB ��xu
�%G    9}~�u�E�!  Y�E�E;�~P�E�  Y�E�%G j[;��9  ;��1  ;��V  �}ĉ}��}�9} u	��%G �M 9}t;���   9Eu���  ;���  9u~jX�  �E�P�u �DQB ����  9}~+9]�rٍEր}� tЊP��tɋM�	:r:�v�À8 u��9}~>9]��=  �Eր}� �0  �P���%  �M�	:r:��h���À8 u��  WW�u�uj	�u �`QB �؉]�;��i  �}���������W  �e�ĉẼM���3�@Ëe��WU  �e� �M���]�3�F3��E�;�u�P�f=  Y�E�;��  �u�SP�u�uV�u �`QB ����   j j �u�uj	�u �`QB ���u�����   �E�   �6������WW  �e���}��M���3�@Ëe��T  3��M���]��u���u�6P��<  Y����t@�E�   VW�u�uj�u �`QB ��tVWS�u��u�u�QB �E��}� tW�]���Y�}� t	�u��N���Y�E��   �}�9}u�t%G �E�] ;�u��%G �u�'  Y�����u3��};�tIj j �EP�uVS�%  ������t�j j �EP�uVS�%  ���Eȅ�u	W�Ӽ��Y븉}�EȉE�u�u�u�u�u�u� QB ����tW裼���u�蛼��YY�ƍe��M��}����S�  ËL$��tI�8 t@��u�I�D$+�HÍ<�    ��$�  9��$�  �dG �5|G �= G ���  ��H�{  �5  G �=� G ���  ��$  �Ƌ�P  ��H�_  ��$�  �=�G �5�G ��$   ������5|G ���  �$�  �$�  ����  �5G �����  ��G ��$�  ��$�  ��$�  ��G �G �G ��G ��$�  ��$�  �` G ��$$  ��$�  �=G �= G �   �ϋ�$�  ���hG 󤉴$�  �5��F �7��QB ��$�  P�G ���F �G �5  G �=� G ��$�  ��$�  ��G ��$�  � G ��$�  � G ��$�  ��$(  ��$�  �����g�����$�  ���@������F ���  ���  ���  F�=�G ���  +�$�  G�ϋ�$�  ���  ���  �-��F ��$�  �5  G ��$$  �-�G ��$�  �|G ��$�  �����F P�������X  ��p  �  ��G ��G �5�G ���  �ˋ��  �5|G �= G ���  ��H��� G �0 G ��\  ��p  �  �dG     ���  �J<ыQ|���  �Yx�$�  ���w  ��p  �K���F �C��d  �K���F �C �$�  ��`  �K$�$�  ��\  �[�G  ��=��F ��G ���  �� G �S�$�  �=t�F ���  ����  �= G )�;=�G ������G ���F ������\  ��  ��$�  ��$�  Y�LG ��G R�-LG ���H�-  ��$  ��G �5|G �ˋ��  ���  ��H�������$(  ��p  ���F ��G C���F +�$�  A��G ��$�  ��P  ��H  �5HG ��L  ���  ��p  �G ��D  �=��F ��X  ��p  �	  ��G ���F �  �$�  ���F    ��ě����G ���F �5�G �l G ��p  ���F ��X  %��  ��T  +�$�  ;�$�  ������  ��G �$�  �$�  ���G �<G +�G ���  ���  0�F ���  ���F @G P���  ��G ��G ���  ��$�  ��$�  �=dG ��$�  ��$�  ��G ������\�F �����  P��G ��󤉵@  �=G ���F ���QB ��$�  P��<  ���F ��<  � G �5HG �=��F ��T  ��H  ���<  Q���F �� G     ���  �J<ыQ|��G �Qx�$�  ����  �J�j�-PG �j�=`G �z �$�  �8G �Z$�$�  �LG �B�$�  �=  �5�G �5��F ǅp      ���  �J<ыQ|�Yx�$�  ��������5��F �K�k�s��$�  �K �$�  ��$�  �C$�$�  ��$�  �K�$�  ��$P     ��R�$�  �$�  ���D  ���F ��T  �5�G ��G �0G ��G �l G ��D  �0G �   �N  ��$�  ���G ���F ���  ��P  ���  ����  �,G )�;�$�  ������.����tG ��G     ���F �T$��T$��-�G �-�G ;l$��ԛ  �-�G -�G �t$܋t$��t$��ډG �D$�    �
  �5�G �TG �%TG ��p  �TG ��$�  ;�$�  �ӥ �5�G �� G ��p  � G �� G ��p  � G �&������  �-�G �E �$�  �m$�$�  ��$�  ��t  �-�G �E�$�  �5XG �5�G �mW�� G ��G �[��`  ��G �  �(G �e������G �}ԋ}؉\G ��G ;8��Y  �}���G ��t$܉�G �T$��\G �������F �%\G �����$   �\G ;��F �2  ��$   �D$���$�  ��$�  ��$�  ��G ���F �5XG ��$�  ��G ��$�  �-� G ��$�  ����   �=G �  ��F    ��"�  P�=�G ��$$  �LG �=`G �8G ��F ��$�  %��  ��$�  )�9�������V  �-�G ���G �u�5G ���������u؉5�G ���m�u؃�A��G �-�G �5G �\$ԋt$��G �T$ЋG �TG �T$Љ�G �L$���  �Jj �5XG ��G ��$�  ��$$  �� G ��$�  ];�$�  �H  �l$�l$���G ��$�  ��$�  ��$�  �x�F �\G     ��   R���F �� G     ���  �J<ыQ|���  �Ix�$�  ���������p  ���F �Q�i�5|G �q��$�  �i �$�  �� G �I$�$�  �t�F    ��	3 ��$�  �= G �����XG ��$�  �{  [��$�  �|�F R�8G ��$�  ���H�:�����$�  ��$   �-dG ��$�  �x�F ����+����=G �=\G �=\ G ���-\G =\G ��A�A��$�  �4 G �=lG ��$�  ��$�  �\G ��$�  ��$�  ��$�  �=\G �x�F ��$�  ��$�  �,����L$̉�G �G �D$؋�G ��G �j�����$�  ��$�  ��5��F ǅ�      ���  ;�$�  ������ G ���F ��$�  �$�  ���  ���  ���  ���$�  ���  ǅ�      ��   ���F �HG �`G B)HG �HG �HG ���xG ��$�  ���F ��$�  ��$�  ��$�  �����F R�HG �5�G ��$�  ��$�  ���  ���UU��V3�PPPPPPPP�U�I �
�t	���$��u����I ���
�t	���$s���� ^�Ë<�F ���  � G �5�G ���  �6����D �=�G �=��F ���  ���  ����$�  �$�  ��A���$�  �5� G ���  �5�G �=�G ���  ���  �<�F ���  � G �f����-��F �D$�싀�   ��L  #��   ��  +��  ��F ���  �Uȉ��F �U��p  ���   �]��ˉ]ċ��F 3��  �M��:  h�   ��,  ��Y�CF ujXÃ  �CF �0�B 3��jh�ZB ��  ��  �e� �}�-   �E�M���	   �E���  ���  ��t$���������YH�V�5CF �`.  Y�0�B ��CF ��+Ѓ�;�sN�   ;�s���QP��O  ��YYu��V�5CF ��O  ��YYu^Ë0�B +CF �CF �����0�B �9�0�B ��^�3�9D$j ��h   P��QB ����E t*�,   ���,�E uh�  �)<  ��Yu�5�E ��QB 3��3�@Ã=�%G u�=�%G r3�@�jXÃ��HG �� G ���H�������F �%��F �LG �X�F Y�-�G �-��F �)�$�  9���� ��$�  �HG �LG ����F ���QB �5xG P��G ���F �xG ��G ��$�  ��$�  ��$�  ��$�  �5HG ��$�  �HG �L$�5�G ��$�  ���#�����|  Ӏ�  �50�F �u�pT���F �F �M��<�F Ӡ8  ���F �]�XT���  k�>���  �X�F ˁ�H  eJ��-�F }K�؁�8  4o'�$�F ��F ���4�F ��F 0�F XT�  +h�F BT�E䋂�   +(�F +8�F �%X�F BT50�F �-��F �<�F ��|  3��F �-�5�F �5`�F Q�M��1R�U��I�M��5�F ZY�   �d�F     h�   �M��N�  W�=d�F ��E��l�F ��=d�F �E�_�҉�$�  �싍$  �G �G ���G ���  ��$�  ��$�  �,G ��G ��$�  ����j �h�F     �h�F �=h�F    �$������F �5�F �5`�F ��H  _�7��=��F ���F ӯ�   �=4�F =0�F �4�F T�F ���F ���F ���   ,��ۉM����   ����   �É�h  � �F ��l  �p�F ���  ��t  �|��x  �(�F �E ��x  +=��F �=��F ��p  ��t  ���  �;��F ��s�����  ��h  ��$�  ��l  ��x  ��$t  ���  ��t  ����q�����  ��t  �D�F �5(�F ��x  �u � �F ���  �;��F ��m����t  ��p  B��x  �D�F �p�F �D�F ���]r����p  ��l  ��������  ��D  �JT���F �7c�l�F �]�+ �F �-�F h�2��M�  ӂ,  ��,  0�F ���]����F �F ���  �}��=0�F ��P  ���F ZT���  3��F �E���F # �F ���F �M苊   �0�F ���F �P�F ȋ�P  ��   ���  ���  �0�F ���  �=�F Z���F �H�F ��  �5��F =t�F �5(�F 9�V�i���=@�F �5��F �=�F ���  �8�F ���F �����U��QSVW�и  �}���VT��5E ��99t�@����;�r�@��;�s99t3Ʌ��  �Y�ۉ]�  ��u�a 3�@��   ����   �FX�E��E�FX�A����   ��5E ��5E �;�}'�R���~T�d8 �=�5E ��5E B߃�;�|�]�	���  ��~\u	�F\�   �d���  �u	�F\�   �S���  �u	�F\�   �B���  �u	�F\�   �1���  �u	�F\�   � ���  �u	�F\�   ����  �u�F\�   �v\j��Y�~\��a P�ӋE�Y�FX����	�u�,QB _^[�ËT$�L$��   u<�:u.
�t&:au%
�t��:Au
�t:au����
�uҋ�3�Ð��������   t���:u��
�t���   t�f���:u�
�t�:au�
�t���눋�$d  �8�F �58�F ��$x  ��$�  �-L�F ��$�  ���F �5��F ��F �ϋË5H�F �-��F ��$x  �=��F �4�F ��������5H�F �4�F ��h  ���F ��  =t�F 9�$h  �8p������d  ���F ���  ��h  ���  ��$d  �0�F ��$`  �H�F �-`�F ��$h  ��$�  ��$�  ��$t  ���F �-��F ��������F ��$x  �����$�  ��$x  ;�F �)�����$�  ���F ��$�  ���F ��$�  �  � G ��T$ �<G ���D������ �F �G A�,�F �G +�G A����G �5D�F ���  ��$�  �t$�� �F �� G � �F ��R��$�  ����$�  �����F �   �5�F ��$t  �5��F ��$�  �-L�F ��$p  ���F �����������F ��$x  ��$l  ����$x  �$x  ��A�A��$h  �d�F �5�F ��$d  ��$t  ��$p  ��$x  �S  ���l���QB �5,�F P�DG ���F �DG ���F �5hG �T G ��$�  ��$�  �`G �t$�D�F �XG ��$�  �T G ���   �5��F �5��F ���F ���  ���F �;��F �q~����C���F ��l  ���F ��������h  ���ً��F ��h  ��l  �5��F �5��F �����5XG P��$�  �d$ ��$$  �� G ��$�  ��$�  ^�.�$�  9����  �5�G P�5XG ��$$  ^�5� G �5XG ���D������$   ��$�  �P G \$�\$����$�  ��$�  ��$�  �LG ��$�  ��G ��$�  ��$�  ��$�  �5P G ��$�  ��G �5� G �=� G �LG �=�G ��$�  �?  ���F     ��$�  ��$�  9=��F �5��F ��$�  �qz�����F ���F ��F ���F ��158�F �5��F Ǆ$x      �����h�F ��F �d�F ��$x  ���F �h�F ��$t  ���F ������T$ �5XG �LG S��$$  �� G �<G ���-8�F ���D������X  ��  ��H�F ��QB �5��F P��L  ��QB ���F ��L  �؋�X  �5`�F ��h  �54�F �H�F ��`  ����  ��$�  �-XG ��$�  ��$�  �����5��F �5��F ��$t  �9��F �0x���-�F ��\�F �58�F ���F �5��F ��p  �����U��QSV��3�9U�U�t5�9�7vj
�[����0�F�	���~��w��7N���N�@;�r��.;1s(N�V��tj
�[�����0�E��N���u�E�)��^[��U������ZV�uW���   ��  ��Muti��%tV��tBHt0��t!H�#  �F�jY������  QX�~  �u�Fj�g�V�u�T�h��  �V�u�T���  �� %����  �u�Fj�1��S��   HHteHHtPHt+H��  �F�jdY���uj��k�d�Z������Y�  �uSWVj�u�  �����o  3��k  �F��ujY��H���N9N}3��   �Fj�^��;���   �   �u�j둃�m��   ��   ��atxHtfHt'Ht���  �u�F@j�]����u�Fj�P����} �uSWVt,j�u��   �����X����; �O�����  ���&���j �ҋV�u�T�8�   �V�u���   �F@�uj�������pt\��tIHt,HtHun��  3�9V ��9E �O�u�F�jdY�������} �uSWVtj����j �����u�F3�B�����~�U���   ����   �ϋ��  3�@_^]�j8h�bB �x�  �E3�+�tH�Et���   ����   �	�E���   �E��M���   �  �}��QB u�QB �EЋ]f�Sf��lf�U�f�SfBf�U�f�Sf�U�f�Sf�U�f�Sf�U�f�f�U�f�u�VV�u��U�RV���   �ЉE�;���   �ủu�������4  �e���}ȃM���3�@Ëe��2  3��M���]3�;�u�u��-  Y��;�tc�E�   �}��u�W�u��E�PV�E���   �U�H;�~ �u�M�> v��]܊���E��H���}� tW裚��Y3�@�e��c�  Ë]�E����t�}�u��]�? t��E� 3҉U؋E�@B8t��E��Ƀ�d�V  �  ��'��   ��At��Ht[��Mt"��a�W  h�bB �]�S�S  YY��uV���e��ItIt#ItI�,  �E�B�#  �E�b�  �E�   �E�m�
  ��ItIt��  �E�   �E�H��  h�bB S�>S  YY��u���]��E�p��  U����!  �E��M����  <'tJ�Ћ]�[H�DS�t��v�M�A�9 ��  ��������E�����@�E��� ��u���  �E��  ��ItIt#ItI�J  �E�A�A  �E�a�8  �E�   �E�d�(  ��h�
  ����   ����   It)���  ��IItII��   �E�Y��   �E�y��   �E�{���   ����   ��uq�? vl��ы]�[H�DS�t�?v@�8 ��   ��
���� ����=�? v8�ы]�[H�DS�t�?v@�8 ��   ��
������@����uËE܉E��   ��ItIt	�9�E�   �E�S�,��ItIt	�"�E�   �E�M���ItIt	��E�   �E�I�E��t#�u��u�u�u�ߋ��f�������u�3������M���Ћ]�[H�DS�t�?vA�9 tً�������A�M���E���������������8 V��tW���t�9��F��8 u�_^�j8h�\B �Δ  �(3E �E�3��}̉}��E��]��}ċE;E�s  �M�QP�5DQB �օ�t �}�u�E�P�u�օ�t�}�u�E�   9}�t���t����u� T  Y��F�u���u�9}�uWWS�uj�u�`QB ���u�;�tX�}��6������0  �e�܉]��6PWS聬�����M���3�@Ëe��l-  3�3ۃM���u�;�uVj����YY��;�u3��   �E�   VS�u��uj�u�`QB ����   9}t WW�u�uVSW�u�xQB ��tf�E�E��^9}�uWWWWVSW�u�xQB ��;�tCVj����YY�E�;�t2WWVPVSW�u�xQB ;�u�u�趕��Y�}���}��t
�M���]�9}�tS蕕��Y�E̍e��M��w����M�  �U����(3E j�E��E�Ph  �u�E� ��QB ��u����
�E�P�;  Y�M��0������$�  �쉕l  ���F ��p  ����  �,�F +P�F 9���  ��h  ���F �}6  �=�B  V�5�%G u3�^Å�SWu95�%G tQ詏  ��uH�5�%G ��t>�\$��t6S��Q  Y���%P��Q  ;�Yv��<8=uWSP荐  ����t�����u�3�_[^Ë�D8��jh�TB ���  3�95%G u5�E�P3�GWh�TB W��QB ��t�=%G ���QB ��xu
�%G    �%G ����   ;���   ����   �u܉u�9uu��%G �EVV�u�u3�9u ����   P�u�`QB ���}؅���   �e� �?�Ã�����8-  �e��u�Sj V觩�����M���3�@Ëe��*  3��M���}؅�uWj����YY����tg�E�   WV�u�uj�u�`QB ��t�uPV�u��QB �E܃}� tV�9���Y�E��n�];�u�t%G �}��u�=�%G S����Y���u3��D;�tj j �MQ�uPW����������t݉u�u�u�u�uS�RB ����tV�Ȓ��Y�Ǎe�艐  ����F     �O<��Q|�Yx�����  ���  �=��F �K�{���  �k�s �$�  ��F �[$�$�  ���F    ��ed ��$t  ���F ��$x  �-P�F �-�F �E��������F �5��F ���  �5�F ���T�����$�  �5G ��$  �5h G �5�G ���<�  �t$��$ G ��$�  ��$�  �������F ��X  �=��F ��\  G)��F ���F ���F �Ë��F ��P  �=��F ���=��F P��T  ���F �54�F �����F ���F ��������F �����=8�F ��t  �F �F ���p  ���$�F ��`  �-��F �=��F �l�F �P�F �-�F �8�F �0�F ���F ��$p  �ϋ8�F ��$�  �=8�F ����   ��  �@�$�  �5XG �5�G �n��$�  ���  ��$�  )�W�� G ��G �[��`  ��G �J9�����������V� G �=��F ��$|  �-�G �% G �5�G �T�F ��$�  ��$�  ��$�  ��$x  �t�F ��$�  ��$�  �5 G ��$�  ;xG �  P�5�G �   �C  �T�F ��G �G �$�  �$�  ���$�  ��$�  ��$�  ��$�  ��$�  �-G ��$�  �|$��$�  ��$�  �G �xG ��$�  ��$�  ��$�  ��$�  ��$|  �  ��G ��$�  �T�F ]��$�  ��$���<��  ���F �\�F +�$  ��G     �=�G     �x ���F ��\  S�  �5`	G ��d  �3P��G �0@�	G S�5`	G ��H�����\  ��G �	G ��G ��듉��  ���F ��h  ��t  ���  ��x  ��p  �5t�F �5`�F h@  �5��F �5t�F ��   �S��$x  �G ��$t  �xG ��$�  �T�F ��$�  �h G �5d G �G ��$�  ��$�  �5�G ��$�  R�d G ��$�  �� �-$�F ���<�p�������p  �=X�F ���F ���  �=8�F ���  ����������  ��$�  �5�F �X�F ���  ��;X�F �eg  ��h  ������j �50�F j�  ���  �J<ыQ|Q�Ix�$�  ���������G ���F ��     ��������  ���  ����  �-`G ��$  �-�G �E �$�  �m$�$�  ���  ��G ������=�G ��$x  ��$$  ��$�  ��$�  ��$�  �|$��$�  ��$�  ��$�  �-G ��G ��$|  ��$�  ��$$  ��$�  ��$�  ��4��������F �h�F     ��l  ���F ���  ���  ��h  W��   Ë쉽p  �0�F �=8�F ���  �5�F �5��F �5��F ����  ��l  +�$x  9�������1���ǅt      � �Q|�Yx����������  ���F �=T�F ��t  ��p  �xG ���  ���F ���F    ��E�  ���F ��d  %��  ��h  �xG �R�$�  �-xG �m$� ��$�  �\$��  ���  �O<�W�5D�F �50�F j�N����$�  �xG �[ �$�  �5�G �5xG �vP)��=xG ����  �I9�������]�����$�  �-��F �/��QB ��$�  P���F ���F ��$�  ���F ��$�  �-8 G ��$�  ��G �=G ��$�  �L$8�T�F ��$�  ��$�  �\$0��$(  ��0��������F �G ��$�  ��L  �5�G �=��F ���  ���F ���G �p�F ��$\  P��H  ���F �h�F ��p  �5�G ��T  ��P  �-PG ��G ��$�  �=T�F ��$|  ��$x  ��$d  ��$t  ��G ��$�  ������O������F �4G C��$�  R�4G �G +T$ B�ʉ=G Y��$x  ���F ��$�  ��G ��4���F P�ʋt$4���-8 G ��$�  ��G �A���V�5��F �5xG �5G �� �E ��  ���F ǃ�*      ǃT)      ��G ��G C��-   �� ��G ���F ��  �5�F ���*  �.E���   ���   ��  ��$�  ��G �G ��$�  ��$�  �݋ˋ�$�  ��F ���   ��\  �=��F ���F ��T  �-��F �T�F ��$�  ��$|  ���F ���F �-x�F ��F _�ދ�$t  ��$X  �=h�F ��$L  ���F ��$t  ��$�  ���F �Ջ�$L  ��$�  ��$X  ������u�����G ���  �pG ���  ��G �G ���  �=0G =�G �=�G ���  �pG ���  ��G ��F ���  �xG ��G 4���  ��G �5�G �5�G �50G �5�G ���   �6�����  ��F ���F ���  3D�F �\�F ���F ���  �=��F ���F (����E�<5  �E�@   �����  ��  h�,  j@��x  ��  h�  j ��t  ��  h�7  j@��p  �"����=��F ���  ���F ��t  �-��F �h�F �T�F ��$l  ��$h  � �F ��$p  ��$|  �ߋ�$x  � �F �͉��F �5��F ��$x  ��$�  ��$�  �-��F ���F ��$L  ���F ���F �Չ�$H  ��$l  ��$�  ��$H  ������{����쉅�  ���F ���  ���  ��G �tG ��G ��G �HG �XG �G ��F ��I������x  ��F �=h�F �5\�F ��F ��t  ���  ���  ��F ��x  ���������  35D�F ���F (����E�<5  �E�@   ���\�F ���F ���F h�,  j@�|�F ���F h�  j ��\  ���F h�7  j@���F ���F j �5��F ��X  �|�F �<�����h  ��d  �= �F ���  ��F ��l  ���  ��F ��t  ���S����-G ��E��G <����   ��t4  0�F ��G �@G ��x�����(6  ���   ���   ��T  ��T  �� 4  ��4  �����   ZT�(  ���   ���  HG 9��������G ���  ���  �=|G �=8�F ���  ���  �=|G ���  ���  ���  �;��F �A�����G F���  ��$�  �5G ���  ���N����5�G �G �5�G ���  ���  ���  ���  �|�����$x  P��$h  ��$x  X���F ���F � G ��$T  �p G ��$�  ���������V�˔  ���Nd;�3E ��   3�;�t/�A,�	;�t��A4;�t��A0;�t��A@;�t��AL���   ��3E �Fd��3E � ��3E 9P,t
�@,� ��3E 9P4t
�@4� ��3E 9P0t
�@0� ��3E 9P@t
�@@� ��3E �@L���   ;�t9u���3E tQ�A   Y�Fd^�jh`\B �  j���  Y�e� �"����E�M���	   �E��  �j��  Y�V�t$�F<W3�;`%G tc;�t_�F,98uX�F4;�t98u;P�E tP蕁���v<�A�  YY�F0;�t98u;^F tP�r����v<�8�  YY�v,�`����v<�X���YY�F@;��B t;�t98uP�=����FD-�   P�/���YY�FP;d%G t;�t9��   uP�Ny  �vP����YYV� ���Y_^Ã|$�w"�t$�.   ��Yu9D$t�t$�#  ��Yu�3���5�$G �t$�����YY�jh@RB �C~  �u�=,�E u.;5D*G w&j��  Y�e� V�@  Y�E�M���3   �E��u#��uF�=,�E t�����Vj �5�E �RB �~  Ëuj��  YÉ�  �5��F =   �4�  @ǆ�$      ��  �tG��  ��G ���$�  �  ��  ��  ��  �<G ��  ��G �<G 믉�  ���F ��G ��I�@����  땉�t�����t5  ��G ��p�����t���ZT��G 3�G ���>���6  ��6  3��5  5������G �� 4  0�F JT�G �E�u���   ��p����p�G ��6  ��6  �X���4  �x�H�G �P�\G �=@G �G ��x����G ��G �=�G ��G ��G �G �  jhPRB �K|  �=,�E u:j��  Y�e� �uV�q  Y�E���t�v���	�u���u�M���$   �}� u�uj �5�E ��QB �����)|  Ëu�j��  Y�U���S3�9%G VWumh`UB ��QB ��;���   �5�QB hTUB W�օ��%G t|hDUB W��h0UB W� %G �փ=�%G �$%G uhUB W�օ��,%G th�TB W�֣(%G �(%G ��t<�Ѕ�t�M�Qj�M�QjP�,%G ��t�E�u�=�%G r
�M �)3��5�M�� %G ��t�Ћ؅�t�$%G ��tS�Ћ��u�u�uS�%G _^[�Í��F �pG    ǅ       �t��   ��pG �g�  ��   �����F ��@�B���҉XG �5pG �%�G ���ߋ�5�G �=G Ë5�G P�T�F �xG �,G �9D$ �y����$G �T�F ��$x  �=8�F Z�=`�F �T$��;�Uĉ=�G �u��HG �=xG �u�E�=dG �pG �=�G �u����u  �=��F ��$�  ��$�  ��$�  �\$��;��F �������$�  �D$����F ��$�  ���F ��������$G ��$�  �=��F ��$�  됉��  �\�F ���F ���F h�,  j@��G ���F h�  j �,G ���F h�7  j@��\  ���F ���  ��p  ���  ��G �=,G ��\  �h�F �p G �T�F ��$|  �K�����G �Uċ5xG �]��}ȋpG �5dG �]�]܋u����@  ��B ���PCF ����T$+P��   r	��;�r�3��U����M�AV�uW��+y�������i�  ��D  �M��I���M���  S�1��U�V��U��U����]ut��J��?vj?Z�K;KuB�� �   �s����L��!\�D�	u#�M!��J���L��!���   �	u�M!Y�]�S�[�M�M�Z�U�Z�R�S�M�����J��?vj?Z�]����]���   +u��]���j?�uK^;�v��M�����J;։M�v��;�t^�M�q;qu;�� �   �s������!t�D�Lu!�M!1��K�����!���   �Lu�M!q�M�q�I�N�M�q�I�N�u��]�}� u;���   �M��ыY�N�^�q�N�q�N;Nu`�L�M���� �Ls%�} u�ʻ   ���M	�   �����D�D	�)�} u�J�   ���M	Y�J�   ��ꍄ��   	�E���D0��E����   �lBF ����   � �E �58QB h @  ��H� �  SQ�֋ �E �lBF �   ���	P�lBF �@� �E ����    �lBF �@�HC�lBF �H�yC u	�`��lBF �x�uiSj �p�֡lBF �pj �5�E ��QB ��B �PCF �����ȡlBF +ȍL�Q�HQP�~K���E����B ;lBF v�m�PCF ��E �E�lBF �= �E [_^�á�B �\�E W3�;�u4�D�P��P�5PCF W�5�E �hQB ;�u3�_Ã\�E �PCF ��B �PCF Vh�A  j�5�E ���4��RB ;ǉFu3��Cjh    h   W��QB ;ǉFu�vW�5�E ��QB �ЃN��>�~��B �F����^_�U��QQ�M�ASV�qW3����C��}���i�  ��0D  j?�E�Z�@�@��Ju�j��h   ��yh �  W��QB ��u����   �� p  ;��U�wC��+����GA�H�����  ����  ��������@��  �Pǀ�  �     IuˋU��E��  �O�H�A�J�H�A�d�D 3�G����   �FC�������E�NCu	x�   �������!P��_^[��U����M�ASV�uW�}��+Q������i�  ��D  �M�O����I;�|9���M�]��U  ���E  �;��;  �M���I��?�M�vj?Y�M��_;_uC�� �   �s��M��L��!\�D�	u&�M!������M��L��!���   �	u�M!Y�O�_�Y�O��y�M+�M��}� ��   �}��M��O��?�L1�vj?_�]���]�[�Y�]�Y�K�Y�K�Y;YuW�L�M���� �Ls�} u�ϻ   ���M	�D�D��� �} u�O�   ���M	Y����   �O�   ���	�U�M��D2���L���U�F�B��D2��<  3��8  �/  �])u�N�K��\3��u��N��?�]�K�vj?^�E���   �u���N��?vj?^�O;OuB�� �   �s����t��!\�D�u#�M!��N���L��!���   �	u�M!Y�]�O�w�q�w�O�q�uu��u��N��?vj?^�M��y�K�{�Y�K�Y�K;KuW�L�M���� �Ls�} u�ο   ���M	9�D�D��� �} u�N�   ���M	y����   �N�   ���	�E��D�3�@_^[��U����M��B �PCF �����S�M���V��WI�� �<��}�}�����M���������3���E���E �؉u�;���K�;#M�#��u��;]��]r�;]�u$����K�;#M�#��u
��;؉]r�;���   ��E �C�����U�t����   �|�D#M�#��u6���   #U��e� �HD�1#u�֋u�u���   #U��E����9#��t�U���i�  ��D  �M�L�D3�#�um����   #M�j _�^�{ u���];]�r�;]�u&���	�{ u
��;؉]r�;�u�����؅ۉ]tS����Y�K��C�8��$���3��z  ��G��}��M�T��
+M�����N��?�M�~j?^;��  �J;Ju\�� �   �}&����M��|8�Ӊ]�#\�D�\�D�u3�M�]!�,�O���M�����   �|8��!��]�u�]�M�!K��]�}� �J�z�y�J�z�y��   �M��y�J�z�Q�J�Q�J;Ju^�L�M���� �L}#�} u�   �����	;�ο   ���M�	|�D�)�} u�N�   ���	{�M�����   �N�   ���	7�M���t�
�L���M��u�эN�
�L2��u��ɍy�>u;lBF u�M�; �E u�%lBF  �M���B_^[��h@  j �5�E �RB ���PCF uËL$�%lBF  �%�B  ��E 3��D*G �\�E    @ÉM��G �dG     �`�F �U�Qǂx      �}�=PG �� pD ���F � G     ǂ,      � G �XG B���  �0�  ���F �]�(�F �$G ��D.  �B���   ���   ��  �t  ��G �E�}��}ĉ�x  ���G �e���Wj@3�Y�t�B �3����E �4�B �@*G ���E ���_�U���  �(3E �E�V�E�P�5��E �DQB ���   �  3�������@;�r�E��ƅ���� t6S�U�W�
��;�w+�A�����������    �˃��B�B��u�_[j �5@*G �������5��E PV������Pj����j �5��E ������VPV������PV�5@*G �)  j �5��E ������VPV������Ph   �5@*G �  ��\3�f��E������t��u�B ���������F ���t��u�B  ��������ƀ�F  @;�r��D3���Ar��Zw��u�B �Ȁ� ���F ���ar��zw��u�B  �Ȁ� ��ƀ�F  @;�r��M�^脠����jhpRB �k  j�w�  Y�e� �}  ���}��w`�u�;5��E t"��t�uV�Sm��Y���E �G`�5��E �u���M���   ����j  Ëu�j�h�  Y�U����(3E SV�u3�;�E�W�T  3�3�9�(2E te��0B=�   r�E�PV�DQB ���!  j@3��}�Y�t�B 󫪉5��E �@*G ��   �}� ��   �M�����   �A����   j@3�Y�t�B �R���]䪍�82E ����)�V��t&����;�w�U䊒 2E �u�B @;�v�FF���u��E���}�r��E���E �4�B    ��  ��,2E ����E ���@*G ��_��u�B @;�v�AA�y� �I���3�A����u�B @=�   r���  �@*G �4�B ��4�B 3����E ����9�$G t�e�������3������M�_^[腞����jh�RB �i  �M��j�t�  Y3��}��=�$G �E���u��$G    ��QB �+���u��$G    �QB ����u��$G    ��%G �E;��E ��   �5��E �u�;�t9>th   �0���Y���u�;�t�u�����Y�E�;�uo�>���E �F�4�B �F�@*G �F3��E��}f�E��E f�LF@��3��E�=  }��t�B �L0@��3��E�=   }���F ��0  @��5��E �}��u;5��E tV�cj��Y��}��M���	   �E��h  �j般  YÃ=�B  uj�����Y��B    3��-�  t"��t��tHt3�ø  ø  ø  ø  É G �(�F �G �]��G �E��G <��G ����� G �]�(�F �E��(�F ��R�E܋E��M�륉<G ��$�  �����G �=�G ���  ��G ;:�H  ��G ��$�  ���  ��G �,G ���  �=�G �|G ��G ��G �5�G ���  ���  ��  ��  ���  ��G ��   U���LSVWjX�o  ��j�E�PV�|QB ��tw�]܍E�P�QB �M���%G �y���#�+���N����������;��M�r@��t\�]��   j�E�P�u��|QB ��t �E�E��]�t��E��E؉E�t3�@�D;�s3��<;�s�u�jS�u��u���QB ��%G ��}�H���%  �M�Q@P�u��u��PQB �e�_^[�É��  ��G ���  ����e�����G ���  �(G ���-(G (G ��A���$�  ���  ���  ��G ��G ���  �G ��G �G ������`  ��F ��$l  ������  ��h  ;��F �C:�����  ��$p  ���F ���  ���F �  ǅ�      �|G ��G ���  ;�$�  �%�  ��$�  �$�  ��G ���  ��G ˋ| G ���  ǅ�      �������h  �H�F ��h  �`�F ��`  ��  (G �E��=�G ��G �U؋=(G �G �=�G �<  ]� �������=   s��ă�� �� P�Q�L$��   -   �=   s�+ȋą���@PÉ��  ���  ���F ��l  ;�$�  �^8����$p  �$p  ��p  ���F ���F �$t  �8�F ��F ǅh      ��   ��p  ���F ���  �R8�F ���  ��t  ���  �A$8�F ���F ���  ���  �I 8�F ǅl      �5������F �xG �]��� �E ��G     �(G     �G ��G �U�B��)
  �z!  �U����F ���1  ���
  ��3  �}��G%�   =�   t�C�����G �|�F ����G ���$����`�F ���  ��d  ��`  �5�F ����������F ��h  ��\  ����$l  �$l  ��A�F��X  �@�F �5�F ���F �`�F ��X  ��T  �����5$G �\G ���  ���  ���  ��   ��d  �5(�F 5p�F 5p�F ����F ���F �=��F ��`  ��d  �5,�F ��h  �5��F �5��F ��`  �=��F ��d  �5��F ����F �(�F p�F p�F ���    ���  3D�F ���F (����E�<5  �E�@   �����F �`�F ��$�  ;�F ���  ��`  �5��F �5��F �5�G �V����=8	G �=$G �7���v  �lG ���F ���  ���  �hG ���-hG ��  ��A�G���  ���  �=8G ���  �=8	G �\G ���  ���  �58G ���  �\������  3=D�F �\�F ���F ���F (����E�<5  �E�@   ����x  ���F h�,  j@���F ���F h�  j ��p  ���F h�7  j@��h  ���F ��x  W�������$�  �=G ��=��F ǅ�      ���  ;�$�  ������$�  �$�  ���  ��G �@G ��=|G �9�$�  ���  �5��F ��H  ǅ�      �j���QQ��%G SU�-QB VW3�3�3�;�u.�Ջ�;�t��%G    ���QB ��xu
jX��%G ���%G ��uX;�u�Ջ�;�u3���   f9��t@@f9u�@@f9u�+�@@��U�^�����;�Yu3�V� QB ���   UVW�pp�������t;�u���QB ��;�t�8] ��t#SSj�VjS�`QB ;�t�V��  �t8Yu�G�?P�|$�����;�Y�D$tb8] ����t:�L$��+D$��+�QVj�WjS�`QB ��t/W�  V�|��E  8YY�tFu�Uf��QB �D$_^][YY��t$�S`��YU�QB �������$�  �$�F B���F �$�F +��F C�Ë��F �,�F ���  ��d  ���  ��P��x  �ˉ5��F �5��F ��`  �����F ���F ��p�F �5,�F ��   ��h  �s������  ������  ���  ;`�F �|�����F ��$�  ���  ���  ���  ���  ���  �P�������G ����F ��G ��$�  �� G ��\  A��G �� G +�G B��G ��X  �G ���F h�,  j@��T  ���F h�  j ��P  ���F h�7  j@�PG ����P���F ���F �,�F ���F ��`  ���F ��\  � �F �,�F �5��F ��p  � �F ����������� G ���)�����$h  ���F ��h  ��$�  ;�F �� ��x  ���F �(�F ��x  �y���������ډ5��F �1�����   ���  Gǂ       ��@  ��G ��L  �tA��L  �O��E ��G ��@  �͋ ��$�  �@�4
G ��   �54
G �W  ��L  ��I�@�Ћ�G 맋8�F �M�A�M��U��U܉�G +U�B�E��m��G �|$ĉ�G �|$ԋ8�F �=tG �HG �t$ȁ��  �58�F S���V  ��$G ��t�t$�Ѕ�Yt3�@�3��jh`RB �Z  �}3�;�u�u�0���Y�  �u;�uW��\��Y�o  �=,�E �.  �]�����   j���  Y�]�W����Y�E�;���   ;5D*G wLVWP�v�������t�}��8V�C���Y�E�;�t*�G�H�E�;�r��PW�u���k��W�?����E�WP�`�����9]�uK;�u3�F�u������uVS�5�E �RB �E�;�t#�G�H�E�;�r��PW�u��zk��W�u��������M���O   9]�u";�u3�F������uVWS�5�E �hQB �E�E�;�u`9�$G tXV����Y��������E3ۋu�}j��  Y�3����w;�u3�FVWS�5�E �hQB ;�u9�$G tV�E���Y��u�3��=Y  Ë�   �G ��������	G ��j  ǅ(     ��	G     ��	G ��(  ��	G �t��	G �J�P ��(  ��	G �͋�@�A�T
G ��	G �5T
G �ǋ�G �G�����$�  ��󤉔$�  �54G ��$�  �t�F ���QB ��$�  P��G ��QB ��G ��$�  ��$�  ��G ��$�  �$G �G ��$�  �8G ���  �  �t$��-�G �5,G �\$�D$����F �D$��E    ��D$��4����tG �E ���F �T$��$G +tG ;D$��PB  �  �}ԋ}�=�G =�G ��-�G �t$܉L$ЉT$̉=�G �\G �T$��|$ԉL$�L$��D  VW�k  �xd;=�3E t�������t$�(�~jPW���  ���
�OH�A����tF���F��-��t��+u�F3���0|
��9��0�������t���A�F�݃�-_^u���j8h�TB �V  3�9%G u8SS3�FVh�TB h   S��QB ��t�5%G ���QB ��xu
�%G    9]~�M�EI8t@;�u�������+�E�%G ����  ;���  ����  3��}ԉ]ȉ]�9] u��%G �E SS�u�u3�9]$����   P�u �`QB ���u�;���  �E�   �6�����������e�ĉE�M���3�@Ëe��)���3ۉ]�M���}ԋu�9]�u�6P�;���Y�E�;��`  �E�   V�u��u�uj�u �`QB ����   SSV�u��u�u��QB ���}�;���   �Et-9]��   ;}��   �u�uV�u��u�u��QB �   �E�   �?�����������e�ĉE��M���3�@Ëe��[���3ۉ]��M���}ԋu�9]�u�?P�m���Y�E�;�t@�E�   W�u�V�u��u�u��QB ��t!SS9]uSS��u�uW�u�S�u �xQB ��9]�t	�u���V��Y9]�t	�u���V��Y���[  �]�3��]�9]u�t%G �E9] u��%G �E �u�(���Y�E����u3��!  ;E ��   SS�MQ�uP�u �4������E�;�t�SS�uP�u�u��QB ���u�;���   �]������������e���}�VSW�7l�����3�@Ëe��&���3�3��M��;�u#�u��A���Y��;�t1�u�SW�l�����E�   �u�W�u�u��u�u��QB �E�;�u3��&�u�u�E�PW�u �u��v��������������u�9]�t#W�U��Y��u�u�u�u�u�u��QB ��9]�t	�u��zU��Y�ƍe��;S  ÉT$���    �t$܋t$�0�;tG ��$ �-�G ���G �E�}�   �:  �-�G �t$؉�G �D$̋t$܋T$��D$��T$ԉL$ЋL$�L$��\$�\$܋-�G ���  �   �m؉�G �G 뇉�G ���F �XG �u��E�    ���F �u䉚/  �5DG �F     ���F �C<؋H|�Pxڅ��,:  �B�Z�j�r 5��F �D$��B$��F �-tG �j-��F �l$�t$��D$�    �-��F ������[�-�G ��|$ȋtG �L$Ћ|$�=�G �D$؉D$�\$�D$��=��F �L$ԉ��F �L$Ћ|$������ډ5�G ��G �uȋE܉E��}ĉ}܉G �E��M��E�M����   ��G ��x  �U��G ������E܉�G �}��MȋEԋډ=�G �MЉ�G �u��XG �5�G �}܋Mȉ=G �]ĉ]܋ڋu���   ��x  �5�G �M������u��5LG �Eȉp �@�����-dG ��$�  �=�G G��5�G �5G )�F�Ή�$�  ��$�  �=�G ��$�  �xG ��$�  �= G ��$�  ��G �xG ����$�  Q���xG �   �|G     ��G �5|G ���  ���  �|G ;8G ��  �|G |G �=TG ߋ��G � G     �?  �G �G ��4  �R�G �  ��󤉼$�  �=D�F ��$�  �:�h�F �5�G P��$�  ���F �xG ��$�  ��$�  ��G �= G �5�G ��$�  ��$�  ��$�  ��$�  ������   �   ���  ǅ�      ���F ��G ��G ���  ��G ���  ��G ���  ���  ���  �   ��|G ��G ���������  +�G ;�G ���  ��\G ���   �o����|G ��    ���  ��G �| G 9��� ���  ���  ��$�  �   ��$�  R   ���  �hG ���  ���  ���  ��G ���  ���  �=XG ��G �   �=|G ���  ���  ���  ��$�  ���  ���  ���  �  �5\G �<G ��$�  ��$�  �ŋPG ��G ��$�  ��$�  ��$�  �\G ��$�  ��$�  �ŋ���   �   ���   �% G ���� G ���  ���  ;���  ��G �|G �ى5lG ���  �5|G �=TG �G ���  ��G �\G �lG ���  ���  �K�����G ���  ���  �o������  ��G ��G     �5��F ���  �5�G ǀ4      �| G �C<؋X|�px5| G ���c�  ���  ���F �F�N���  �~���  �N | G �=�G �~$=| G ���  �N| G ���  ��������  ���  �=XG ���  ���  ��G ���  ���  ��G �������G ��$�  �-�G ���-PG �-�G ��G �=�G ��$�  ��$�  ��$�  ��$�  ��$�  �=�G ��$�  ����   ��������  ��G �G ���  ��G �����������  � G �<G ���- G  G ��A�C���  �LG ���  ���  ���  ���  �/  ������TG ��=HG ��H  ��5  ��  ���=HG �DG ��  �� ����DG ��  ��G �DG �F  ��G ���  ��G �$�  �$�  ���G ���  ��G �5�G �=�G �|G ��G �5�G ���  ��G �5�G ���  �������u�u�95LG ���  �G �8�F �LG �]��U��}��5�G �]��=8�F �u�]Љ��   �XG �U��G �E�� ;��F �<�  �=G �E��M��]����W�  ����뤉5�G ���=G ��  ��G �	��G �A��=HG ��  ��G �� �����  ��  ��   ��$  �-�G ��$P  ��$  Z�t$�|G �Ջ5�G ����  ��$   ��G �|G �D$���G ��G ��R�@��G ��G �D$���G ��G ��  ��  �|G ǅ����|g S��(�8G ��������G ��G ��I�@��H  �������G ������58G �� ����TG ��H  �=|G ��G �[������  ����=��O��
G ��G ���   �牍H  �G ��  ��G ���  �4G �Ӊ������G W��  ǅ      ��G ��  ��  �|$�8G �y����G ���  �LG ��G ��G ���  ���  � G ���  ���  �=�G �= G ���  �G �������	G ���F ǀ"     ǅ8      ���   ���F ��8  ���
G �%�  ��8  �։�G Y�-|G �5�G X�-�G ��$   ��������$   P�-�G �5�G ��G �L$��|G �H��=��Q�-|G 롍��F �@G ���  ��I�@��<  �Ћ@G ��<  ��G ���J������F ���  ^���F )�vV��  5p�F ��`JC���0  ��@  �	  � �F ��  �L�F     �@�F    �@�F �< �T�F Q�L�F ���D  � �F �L�F 1�@�L�F �T�F Y� �F 뷋5��F �}��=��F �7�d�F �4�F )��=��F 0�F �E̋�`  |�F �F �Eȋ��F ��  �E��E�0�F ���  ��'7�  ��$  �|G �-�G �M �m�A�-�G �  h  hTB �WE  �(3E �E�%G 3�;�t�M��u�u��YY�M���  3�@Ëe���EHt�$TB ǅ����`SB ��   ��@SB ǅ�����RB ��   �M�h  ������PQ�LQB ��uhHTB ������P�"  YY��������P�Z  Y����<v%��P�I  �؍�������1�jh�RB S��M����S�&  Y�D0������f����e��WV�:"  ��TB WV�>"  h�TB V�3"  SV�,"  WV�%"  ������V�"  h  h`TB V�H�����<j�5�  ���������������U��WVS�u�}����
�t2����'��8�t�,A<ɀ� �A��,A<ɀ� �A8�t�����[^_�Ë=0G j�l$W�5�G l$��$  �|$��   �=|G �=DG Q�5�G �|$�L$�`G ��$  �DG ���������$  �|G �5�G �<  Y�`G �-|G �C�����|G P��
G ��G %�   ���%|G j ������=|G R�T$��$  �xG ��G � ��G �@�HG Z�xG �HG �T$�T$��-�����  �-4�F rZ�x�F �4�F j �d�F     �d�F �=d�F    ��������F ���  ^���@  ��F )�v���F �4�F 0�F yT��F ��  ���  S��QB ���F ���F ���	  �- �F �5h�F j����ÉL$�T$Y�`G ���<������F ɉE���  +�l  -ѝ���-L�F �M���  �M���  �-��F ��p  3�@  ��X  =��F ���F ���F �U�0�F ���F ���F P�F AT��$  �}��=��F �|�F �E����F ��$  3��  �n  �5�G �5��F ��G ��G 0�F �}��}�U��U���3  ���   �]���  ���   �L$ĉ��   ��  ��  �-\	G �j���F �  �=��F Y��l  �X�F �
��H  ��l  12�R_T��t
  ������F ��d  _T��t
  =��F ���F ω�D  � �F #��F �����Ճ�����̋L$��   t$�����tN��   u�    ��$    ��$    �����~Ѓ��3�� �t�A���t2��t$�  � t�   �t�͍A��L$+�ÍA��L$+�ÍA��L$+�ÍA��L$+��U��Q3Ʌ���u�Ã? t	��A�8 u�S��   VP�I�������Y�u�uj	�  Y����P�*p��������Y��u�!�E�^[��U����ES3�;�W�]�u����aV�0;�u�tSj=V�  ;�YY�E�tB;�t>3�8X��%G ��;�%G �M�u���H�����%G ;�uU9]t9�%G t�J<  ��t?���^_[��9]�t3���j����;�Y��%G tމ9�%G uj�j���;�Y��%G tÉ�}�+}��u��5�%G �  ��;�Y|F9tB�4��6�A��9]�Yu�E���E��g�F�G��9u����P�5�%G ����;�YYtC�<9]���   ;�}�ߍ�   P�5�%G ����;�YY�4����U�����Y�M���%G 9]tP�u�����@@P觿����;�YYt8�u�V��  ��+E�YE�Y�M��@�����#�QV��QB ��u�M��V�8@��Y9]�t	�u��*@��Y�E������u��@���EY�����V�5�%G �"WP�t$��;  ����u��<=t��t�����u؋�+�%G ^����Ë�+�%G ^��É��1  ���1  �G �ö;ee��@3  T	Q��$0  !!o!0�F �G �0�F ��  50�F �5G �5��F ���1  �p2  �5G d�5    d�%    ��  ��$  ��G ��쉵$  �5��F d�    �d�    ��L3  �-�G �pG Ӧ�3  ��(2  ӎ�3  ��1  �\G ��   ���3  3�G ��  �\G ^T�50�F j j
Q�����ÉB���   �ht�Ht�J�t$̉r���  �j����F ��G     �XG �@G ��G �]��G ��G ��G �@G �]�}�E�uY�m��T$�G �=\G �0G �5�G ��G �-�G ��G �D$��|$�L$�T$�l$��\$܋t$؉�G �=�G ��  ��,�`G �G ��G ��  ���  ��H  �Ӌ�  ��  ������`G �� ����-�G ��$  �|$�8G �-�G ��G �DG ��$  ��$  ���T$�5t�F �~������$�  Q��)ȋt�F 3M�)ȋ��  ���#�����  X���F ��1�)�$�  �=d�F ���  +�$|  ���  ��)=��F ���F 3�$�  )��F ��$�  ���  �$�  9����  �G ���  �58�F ���  �5G ���  �=G �/;-��F �q�  �-@G G��N�����  �@G �=`G ���  ��G �`G �G ��G ���   ��E�    �\�F    �\�F ���  �5L�F �}ȋ71��}��݉0G �,G �-�G ��G �5$G �t$ԋ|$̋l$ȋD$ċT$��5|G �=�G �-G �XG ��G �%4G ��G �XG �-@G �5�G �=@G ��É�G �%�G ������  ��G ;�F �6J������G ��G ���  ��� ��$�  ��$�  ����F ǀ�      ���  95�G ��[�����  ��G ��G �G ��G ���  ���  ы�$�  ���  ��G     �?  ���  ��l  ��3d�F )��F ���F ���F +$�F �\�F �d�F +��F ���ˋ5\�F ���  ���F �-���� �UV�D$�u(�L$�D$3���؋D$������d$�ȋ��d$��G�ȋ\$�T$�D$���������u�����d$�ȋD$���r;T$wr;D$v	N+D$T$3�+D$T$���؃� �ʋӋًȋ�^� �����������U��V3�PPPPPPPP�U�I �
�t	���$��u���
�t���$s�F��� ^�É��  ���  ��G ���  ���  ����������G ��G ��G ���-�G �G �-�G A�G B���  ��G ���  ���  ��G ���  ���  ���  ��G ���  �5�G �5�G �5�G ���  ��G ��G �5�G ���  �6�����G �}̉0G �Uԋ��]Љ�G �XG �pG ��G ���t �E��E�� G ���m�E��m�AE�A�a�G �]́e�����M̉]��G ���   �}��}��]�;;�,j  �}��G �Ӌ}܋EȋM��}̋0G �E���   �}��^  �0G �M��8G ��G �=�G �pG �}̉u��U��u���G �u��E��u���G ��G ������=��F �G     �=G ;}������=G =G �EȋẺE���M���HG �U��}��}���   ��x  ���G �E�    �����5t�F ������  �@W�=��F �=(�F �<}    ���  ���F ���F Z���  ���  �3�$�  �   )�ǅ�     ��p  �΋��  �3��F ��$�  �ˋ5G ���  �G ���  ���   �  ��x  �EȋM������� ��  ���  ��  �=�G �   ���  ��$�  �G �5�G ��  �[�=�G �  ��8G ��G �$�  �$�  ����  ���  ���  �8G ��G ���  ���  ���  ��  ���F ���   35��F ��d  P��@��ǅ|���@   �xG ��<  ��x������  ��t�����h   ����`  V����G �\	G ��  ��$�  �4�I �$<  ���-  �=�G Ǆ$�      ��l
  �= G ��$�  ��G ��$�  ��$�  ��$�  ��G �=�G �=@G ��$�  ��$�  �   ���G ��$�  �1�7�  ����<G )�;TG �t!  ��  ���  ���   ��  ���  �5�G �G     ��  �5�G ���  ���  ǆ      ��P  �C<؋H|�Xx�$<  ����"  �5��F �C�s���  �[�-��F �=@G ��$�  ��$�  �R�$<  ��$�  �TG ��$�  �@$�$<  ��G �(G ��$�  ������G ���  ���   ��   �5�F j@��\  ��l  ��G ���F ��4  ��T  ��B���5��F j@�5��F �5G ��<   ���  ���F ��P  qT�`G V��L  ��X  ��H  ��p   ���  ��`  �	G �D	G ��$�  ���   �dG ��   ��$�  ��$�  Z����Ŕ   �  ���  ��    �=�G �48�$<  ;5�G �p ���   �I��$�  ��$�     ��   ���  ���  �=�G �5�G ���  ���=�G ��$�  �-G �XG ��G ��G ���  ��XG ��G ��G ��$�  �-@G �=�G ��$�  �������G ��@�B��	G ��G ��	G �m  �ˋ5G ���  �G ��G ���  �l������= G ���  ���F ���QB ��$�  P�,G ���F �hG ���  �,G ��G ���  �<G ��G ���  ���  �5�G �����   ������G ��8  j@��\  ��$�  ��G ��4  ��\  ��A���5��F j@�5��F �5G �dG ��G ��P  ST� 	G QVh�  �5�F �5�F �  ËL$�T$f�f�AABBf��u�D$Í5��F ǅ(     ��g  �\G �5��F ��(  ���n�����   ����  �G ���F ��G ��	G ��(  ��$�  �5G �hG ��   ���   ��	G ��G     ��(  ����dG �G ��G ��	G ��  ��   ��G �dG ���   �  �;  ��(  �+����(G     �5�F j �5��F �Y����=(G     ��  ���F ��L  ���F V�5(G �R�U����    ��"  NW�<�<��_����F ���  �=�G �=�G G)5�G ��G ��G �։�G ���  ��G �hG ���  ���F ���  �5��F ��P��G ��G �5�G �&����
G ���F ���!  ��8!  ��I�@���  ���\
G ���  �  ��G �D�����W�=0G �=|G _���l�w  �M��`�F �%@�F � �F ���F ȋt�F Ӄ�  ���F ��t  �  ���  ���  Ӄ�  �=��F �=h�F =0�F ��d  �݃�����u܋5 �F �`  ���  �%`�F ��F ӣ  ���  ��UO�@�F 3��F �5 �F �5��F �`�F 
�-}0�F �4�F ��  ��v�}؋�l  =,�F ��X  w�΋�  ��  �=�)G u聈  �t$豈  h�   �}  YY�j`h`aB �H+  ��   ���,����e��>V�4QB �N��%G �F��%G �V��%G �v���  �5�%G ��t�� �  �5�%G ��£�%G 3�V�=�QB ��f�8MZu�H<ȁ9PE  u�A=  t=  t�u��'���   v�3�9��   ��ytv�3�9��   ���E�j�C���Y��uj����Y�@  ��uj�����Y�*  �u������}j��   Y�,���L�E �������)G ������}j�   Y�����}j	�   Yj��z  Y�E�;�tP�   Y�u��E�P�TQB �m����E��E�t�E��j
XP�u�VV��P�&�  ���}�9u�uW��{  ��{  �+�E��	�M�PQ�E���YYËe�}܃}� uW�{  ��{  �M���Ǎe��)  Ã=�)G u艆  �t$蹆  h�   �\7E YY�����������̋D$�L$ȋL$u	�D$��� S��؋D$�d$؋D$���[� �5��F �(�@�E�-\G �싵�  ��\G ������h������h�  N���  �hG ���  ���   ���	G ���F ǅ�      ��-  ���F ���  ���	G �,~  ���  ��+h�F �Uԋ �F 3��F ���  �-��F +��F ����f�VT���  ���F ��  �X�F �4�F ^T�EЋ��  \�F ���F �ʁ<�F Pg=�VT+��  �  ��$�  �G ���F ���QB ��$�  P�(G ��QB ��$�  �(G ��$�  ��$�  ��$�  ��$�  ��G �dG ��$�  �G �0G �dG ����������F W�=d�F ��u��5l�F 7����F ���F ���F Ӏ�  ��   r����   ɋ��  =0�F �5��F +�T  0�F ��F  �F �����|G     �=��F     �Q������F ��S��\  �L	G ���F ���F ��d  �HG ��B���5<�F j@��<  ���  ���  ��X  ��G ���F �5�F Q�5`�F �����Í��F ��@�A����������F     ��F    ��F �J����5��F �\�F ���F �2�E��4�F )�R���F �E��\�F 뿋0G �   �(�F ��$l  ������F ��$l  ;�F ��������F ��$�  ��$l  ��$h  �-l�F �=�F V�-��F �=(�F ���F ��$d  ���F ��$p  ��$�  ���F ��F �   ��G QA��^��$�  )�F�ƉG ��$�  ��$�  �=�G �=0	G �5�G ��V��$�  �ȋ5G �G ��$�  �������  ��G �=tG Q��$�  ��$�  �=TG ��G �T$����$�  ���l��������F ���F ���F ���   ��$d  �@�F ��$`  ���F ��$X  ��$t  ������<�F ���F ��$\  ���F �|�F ��$t  ;5�F ��������$x  �"�5�G S��$�  ����$�  ���l��������F ���F ���F P��$|  ;�$h  �H�����$|  �$|  �=��F Wǋ8�F �5P�F ��$h  ��$x  ��$t  Q���F     ��$�  �T$��$p  ���F �_  ����d  �X�F �$�  9���������F ��\  �8�F ��`  ��F ��`  ���F � ;��F ������X  ���F ��`  I��������X  ��\  ��F 밋���F d�    �d�    �=��F �G �,t�5G 3� 1  ���3  #`G ��x1  DDgwT+lG ��(3  �TG )��Z�=G 3=�G ��x  ���F ����  j�5�F h�  j<h�  ��  Ë�`  ��G ��P  �l�F �5G �5 G ��X  �G ^���F �  � ����UW�|$�n��$    ���L$W��   t�����t=��   u�������~Ѓ��3�� �t�A���t#��t�  � t�   �t�͍y���y���y���y��L$��   t�����tf�����   u���������~�Ѓ��3��� �t��t4��t'��  � t��   �t�ǉ�D$_�f��D$�G _�f��D$_È�D$_�U���5  �@`;��E t������x u]��P���MSV�/���DtA���t;�������9Uu�A��"��9ut
Af�f��uȋE��+������#�^[]�3���B��$d  �5��F ���F P�����F ���F S����������$l  ���F ���-��F ��F ��A�BQ��$�  �5��F ��$�  ���F ���F ���F ��$�  ��$�  ��$p  ��F ���j������  ���F ǅt      9�$x  �������t  ��$x  �$x  ���F ʋ*-8�F �-��F Ǆ$t      �=t�F ��$p  ��$�  ���F �=<�F ���F 3=��F �=@�F ��$h  � �F �%��F ���F ��$l  ���F ���������-��F ��$t  �-��F ���-��F -��F ��A��x����l�F �E�V���F ��G ����-  ��d  �G ��G ���-G G ��$�  A�$�  A��`  ��X  ���F �l�F ��X  ��P  ��T  �?�����d3  �%�G =0�F �-TG ����G �81  ���2  �ˋTG 0�F ���F YT��2  ��G �XG ���F Sd�5    d�%    �G ��G ����F ���F ��$�  �=P�F ��$p  ��$d  ���V�����F �5$G F�ǋ$G �`G )�A���}Љ]���F �|G ��F ���  P�u���G ���M��G ���F ���QB �5��F �]   ���G     P�E�S��G ;D G ��N����G �G ��l  Y�pG ً�$�  ��G �G     �	����u�P��G ���F �E��M��G �}܋]��5HG �pG �<G �5PG �G �E��E�pG �ĸ  �   ��d  �%G ����E��G ;��F �&P���E���G ��`  �E���l  �pG ���������F W�=,�F �W<��z|Q�Jx,�F ���ܮ��W�=��F �Q�y�4G �QR�Q ,�F V�q$5,�F S�Y�  � G �u��)������DG �xG �=xG    ������G �5G �U܉�G ]�DG �t$؋PG �L$Љl$��G �D$�|$�|$؉�x  �v��G �|$��T$��L$܋\$��T$��[  ���U��U��G �G ��=�G �U��Uȉ�G ��G �]ȋU�]܃��)�;4G �r�����G �U��%�G �pG �DG �M؋�G �
,�F ;E��� �E�pG ������G �%8G ����E��8G ;��F ��L���E���$�  �@G ��G �\G ��X  �t G �hG ��T  �5�G �5��F ��T  ��   ,�F SV�xG     �`�F �5�G �G �u�}̉uĉ]��}�u�]�W�uȉPG �pG �U�`�F �U�E�   ��M��M��   ��  �pG �]܋u���<G �����E܋]؋�U܉=�G �$G �UЋ}܋E܉=tG �Eԍ@�$G �ڋ=�G ���F ��  ��l  Y�I�$�  ǅd      ��`  �@G ���F �E���X  ��d  ;�$�  �wA����$�  �$�  �hG ��`  �t G ً�$�  ��G �8G     �   Q�pG �l$��t$�U�5�G �t$��DG �t$ԋPG �L$؋l$�|$�-�G �=`�F �D$܉D$��G �|$�5G V�t$؃����,�a�����H  �8G ��T  ��P  ��G �=8G ��H  ��L  �=DG ��]�]܉��  �[�]����   ��`  �E��=DG �pG ��G ����R����=8G �=� G ���-8G =8G ��A�C��T  ��G �=TG �pG ��`  ��L  �=����D$f�@@f��u�+D$��HÉE܉��F �]��G �]؉hG �M��G 4
�X�5��F ���	  ���-  �E�    �E��M�G ǁ�      �5xG �5 G �� �E ���F ǂ�.      �E�    �E܉xG @=�   �Y{  ���F �]؋]܋C���   ���   �2����C����m؉d�F �5��F ���F �4�F �=L�F ��F �-��F �\$����F �%��F �H�F ���F �-��F �5,�F �=��F ���U�D$�싀�   �- �F ?����$  HT�X�F ��  ���F ��F Ӏ4  �,�F ��F ��F 0�F V�M���   ��  ���   �%��F �D$��G �l$�tG ��G �Ήl$܉\$؋\$�\$�=G �\$؋=�G �=�G �=G ����n����L  ���  ���Q��F ӆ�  ��  �x�F ���  84&U���F ZVT^T���  �Љ]苞�  +�,  ���  ���  ^T���   
���F ���  h)�]䋞�  3��  ^T���  ]�걉��F ���  VT�5��F e� ,�}���H  +��  �<�F �ϋ��  ���F �`�F ��  #��  �J�D$܉�G �|$ԋtG �ŋ΋|$�|$؋\$�\$��G ���F �|$ԉ�G �ŋ���8������  0�F =0�F ���  ���  ��)@�u���   �}܉��F ���   �M؉�F ���  ���   �Uԉ~���  ���  �=��F �~��F �^��  �~��F �^���   ǀl      ���  �U �}��M����F ��  ��P  ���F �E��u�Z�M�}�]��������(  ��G    ��   ��G ��4  ��	G ��G ��8  ��<  �5�	G ��c  �=�G ���l  0�F ��,  �LNI��F ��F NT� �F ��  @�F �H�F ��l  Q��l  0�F Q���  ɉ<�F ���F ��VT�|�F ��`  VT���  �-��F �%��F P���F +�  �\�F ��x  �F ���F ��%���  Ӯ�  ���F ���F P�F +��F ��  ֨�?���  +��F �e��M�LG �� pD �E�    �E�    �Uȉ�G B��   ������}��=t�F �dG �Mȋ9�Eȁ��   ���   ��   �ߋ}��  �֋�(  �=�G ���@�=�G �Ћ5�G ��<  ��(  �N��  ��	G ��4  �5�G ��G �5�	G ��(  ��8  ������<  ���F ���   ���"  ��<  ��
G �   ��0  �$  �=�G ��<  ��$     ��  �xG ��0  ǅ(      ��0  ��
G �=tG ��$  �g����M��}��dG �t�F ��R�M��E��t�F �dG �Eȉ= G ��G �}ĉU�}��}ċE��E��= G �o����Ű�v�DG �֋DG �u��   ���hG ���  ���  ���  �4G ��G ���  �(G ���  ���  �֋�G ��G ���   �  ���  ��G ���  ���  ���  ��G ���  ���  ��G ���  �5`G ���  �5(G ���  ���   �T  �Ủ5�G �PG �G �E���   ���  �PG �MȋPG �U؋�G �  ���tG ��$�  ��$�  �(G �lG ��$�  ��$�  ��$�  ��G ��$�  ����   �   �XG ��G ���  �[�   ��E���G �=`G �E���G �}؋dG �=�G ��   ��E؋�G �=�G �E���G �dG �U؉�G �5�G �5`G �u؋5�G �   �5��F ���  ���  ǅ�      �=H�F ���  �=�G ���  ǁ�      ��G ��j �5��F �58�F j(�  ÉU؍��F �50G �E�ǂ,      �58�F �E䉲�-  ��G ǀ�       ��G �E�- @ ��G     �E�    �ủ5�G F��B  ������]���   ���  �ŰB���   ���   �����������G ��$0  �5�G ɋ�	G S��$  �-�	G ��I�v����$4  ��Q�=pG ��G ��$  �=�G ��$  �=pG Z�  Qd�5    d�%    �@�F ��G ����F ��G #�G ǅT���@   ��`  ���  ��P�����\  �E���L���R����F ��X��������  �<G �HG �5�F S��   É<G ��G �U����   �R����X�5�G ��  �5�	G �Ћ�=TG ��$0  �=|G �=�	G ��G ��[�@��$  �=TG �5�G ��G ��$  �-�G �-�G ����� �����$  ��	G ��$4  ��$   ��$�  ������   �`h�  S�58�F �5`�F j ��   �=pG     ������\  RpG �G ��G �pG �B�pG ��\  ��빉�G ��  P���  �5�G ��G ��	G ��  �|G ������Z�-�G ���T$���$0  ����W����G �=0G ��G ��G �<G �'������  +G �pG     � ��G ��  ��G �5�	G �hG �=G ǅH      V������=�	G ��  �=�G �hG �=G �ދ5�G �������0�F ���F �=@�F ���  ���F �$�  �<�F ���F 9=��F �������p  ��h  ���F �=8�F ���F ��l  ��t  � �F �   �5(G �U����F �\G ��h�����\  P��G �=0G #�G ��d�����h����\G ^�=0G ��G ��G ǅH���@   ��G ��D�����@����=�F ���h����<�F ���F ���  ��p  3��F �D�F � �F � �F �%��F ��l  �5��F �;��F �t�����<�F ���F ��p  O��������<�F ��l  ���  W���  ���F �  �|G �=�G ��   ��v�@�ȋ|G ��   ���  �|G ��0  ��   ���lG    ��G     ���  ��0  �E���  ��G ���  ��G �=$G �=lG ��  �=$G ��   �2��0  � G ��G �,G ��   ǅ     ��G     �5�G ��   �dG Wɋ�  ��0  �����|G �=�G ��G �5�G �=dG ��   �dG _��G ���G ������0  �@G ��   ��G ��  �@G ��0  ��G �dG �dG ��0  ��   �M�����  ��$l  �=��F ��$t  �5<�F ��$l  �)  ��`  �TG �� G �M��� G �9�$�  �$9������`  ��T  P�8�F �XG �\�5  G �=� G ��$  �5|G �= G ���  ��$  �$�  9���M����G ���  ���  �8�F �XG �  ��P  �TG ��L  ��H  ��`  �;��F �Y3����H  ��D  ��$�  �TG K���^2����D  ��P  룉��F S��$l  �5��F �=@�F �<�F �=t�F ��$�  �0�F �=��F �D$�5D�F ���F ��$�  �=��F ����   �  ����}  �Eȁ�����pG Y;���������G �=�G �u��U�X�5�G �U�E���G �]��]��E��뭉< G ���  � G ���  ���  �	;��F ��M����H��$�  �< G ��P  �< G ���RL����P  ��T  ��G �< G ��H뒉��F �=��F ��$�  ���F ��$�  �<�F �;��F �������$x  C���F ��$�  ���F ��$�  ���A�����$x  ���F ��$t  ��$�  �|$��$�  �'���V�t$����  �v����v����v����v����v����v����6�~���v �v���v$�n���v(�f���v,�^���v0�V���v4�N���v�F���v8�>���v<�6����@�v@�+���vD�#���vH����vL����vP����vT����vX�����v\�����v`�����vd�����vh�����vl�����vp�����vt�����vx����v|�����@���   ������   ������   ������   ������   �y�����   �n�����   �c�����   �X�����   �M�����   �B�����   �7����,^Ë�d�    �d�    ���F ��$  �tG ���1  ��H  ��{  ��G ���5�G ��  �G �щ<�F ���F V�5t�F �$�  95<�F �����V�t$U�8�F �-<�F ��$�  �-�F �I�����G     �HG �U�]܉5�G �pG �u���G ;U��ƈ����G �G �U�PG �4G U�,�F ��G �E�    �   U��QQSV3�W�=�%G �u��;�tb�xQB VVVVj�PVV��;ƉE�tZP� ���;�Y�E�tLVV�u�Pj��7VV�Ӆ�t1�E�VP�������YY}9u�t�u����Y�u����;�u�3�_^[���u����Y������G �U��pG �U��G �=�G �=HG �}�]܉MЋ�G ����Q�������A��G �M���	����G �G �=�G �U���G Y�U���G �]��G �]�]܃��p���U���  �@`;��E t�^����} u3�]��p�u�u�u�uj�p��C������u����]Ã��]Í=��F ǅ<     ��
G     �t#�=��F �=�
G ���$  �ez  �=�
G �ٍ=��F ��8  ���  �	���  �A��0  ��8  ��0  뱋5XG ��$�  ��$   ��$�  <G 9�$�  �2q���싅�  �58�F ���  �5��F ��   jh�\B �~   �E�@cB �}�@cB s"�e� �E� ��t���3�@Ëe�M���E����   �jh�\B �:   �E�8cB �}�8cB s"�e� �E� ��t���3�@Ëe�M���E����>   ���hiA d�    P�D$�l$�l$+�SVW�E��e�P�E��E������E��E�d�    ËM�d�    Y_^[�QÉ��  ��G �5XG ��   ���  ���F ���  �;��F �y^��� G A��   ��$�  ���  ���;^��� G ���  ��G ���  ���F ���  ���  � G �p����XG ���F ���  ��H  �=�G S��G ��  ��G �-8G ��  �=XG ��G ��$�  �-�G �5�G �=�G �|G ��G ��	G �5|G �=�G ��$�  �=G ��$�  �����z��  ���F �,G S���$  ��G ��H  ��  ��  ���$  ���#  ���$  ��P%  ��	G ���$  _�D$����"  �=�G ��$  �ˋ=�G ��  ���   �  �50G �5�G ��v�@�5�G P�|G ^�  P�8G ��G ��	G ��  �5�G ��H  ��G ��  �5�G ��  �5|G [�G �*  ��I�@��G �5XG S��G �tG ��  �?�  ��H  �5�G ��G ��  �=8G �|G �=�G ��  ��	G ��  ��G �5|G �tG ��  ��G �G ��H  ��   V�5�G ��v�@�G �5�G ��(����5G V��H  ���  ��$�����G ��  �|G R�=�G ������TG    �G     ��H  �� �����  �TG �-G Z�DG �l$ ����   �m  ��G ������   ��   �5,G �l$���$�  �5�
G �-G ��$�  �5|G ����   �   ��G ���   =G ���   �G ��G ��H  ��(���Y��  �5(G ������� ����% ��������A�tG ��  �G �5G �xG ��(�����H  �5�G ������G ��  �  �<G ��G ��  ��	G �5G ��G �5�G �=�G ��  ��{  ��G ��  ��	G ��G ��  P���  �<G �G �G ��0������  �|G ������  ��  �|G ��  �� �����	G �G �5|G �`G ��G ��  ��(�����0����`G ��G ��  ��  �����=�G �;��F ��<����$�  ��$�  ��$�  �-��F ��G �5pG �-(G �tG ��$�  �tG ���r@����$�  ��G �=�G �dG ��$�  ��G ��G ��$�  �|$X�5�G ��G ��$�  ��$�  ��$  �@�F �-��F ��G �tG ��G �=�G ��$   �-� G ��$�  �5�G ��$�  ��$�  � ��G ��	G �(G �= G �=G �������G S��  �8�  ��(�����G ��'����=�G ��  P�k�  ��$�����G ��  �|G �DG    j �� ���W��  �DG ��=�G �|G �,  �5@G ������I�zL  �� ����=�G �5 G �DG �5@G _������ G ����������닉�G S��G ��	G ���  ���  �-�G ��$$  ��G �|$�-|G ��$�  ��G Z�=�G ���\$���G ��G �\$���$   ��	G ��G �G ������G �G ��	G ������   �g����xG �5(G ��  ��H  ���G����	��G �AQ��G ^�l���P��G ��G ��	G ��  �5(G ��H  ��G ��  �5�G ��  �5|G Z�(G ��G �(G ��G ��$�����G � G ��H  ����P��G ��G ��$�  �-|G ��G ��$(  ��G �t$�T$�5�	G Y��$�  �֋�G �-�G ��G ��G �\$��-�G ��$�  ��$$  ��G �5|G �����=�G ���@��G �=�G �� ����=�G �5�G �����@�F ���  0�F �tG ���F @G R���  �� G �Ћ��  ���  �5�G ���F ���  ��$�  ��D�5��F ��$�  �hG ���F ��$�  �h�F h�  j h,  Q�d�����@����F ��I�B����   V�=TG �5��F �=�G �5(G ��$�  S��G ��$�  � ;��F �z4��P�=TG ��$�  ��G K���7��]�t$��뜉�<  �8G 0�F ��8  ���F �=PG ��8  �Qd�5    d�%    ��t4  ��D��-�G ��4  ��D  ��7  ����   ���  ǅ     ��G     ��������G ���$�  �j�  ��G �ۋ쉽@  �=��F d�    �d�    �,G � <��lG ���<5  ��G �G 3��4  �8G �LG ӏ\4  �G 3�5  �=,G =�G V�5t�F �5��F �����Ë�I�C���,�����$�  ��$�  �-HG ��$�  ��$�  �-pG �5�G ��G ��$�  ��$�  -� G 9�$�  �~-����D��$�  �8�F Q�lG ���������G \$�9������-$G �쉍�  ��G �8�F ���  ��`��d  ��G ��H  �;��F �)����D  C��d  ��G ��G ���e����@  ��H  ��d  ��D  ��G ��@  ��G ��`댉��  �=��F ���  ��`  +��  ��G ��F 9��!����G ���  �8�F �G �K����E����F �E�0�F ���F ���F ��H  +=��F �}܍=��F ���F �8�F ���  �-,�F �u�wT�U؋�P  +��F �����  #��  ����n���  �]ȋ��F ��  )��F ���F +x�F ���F ���F ���F ���  �=��F �����F �EЋ��F �����X~  ���  �5�F �E�=��F �]ȋUԉu��E��a  ��G ��$�  ����LG ��$�  ;�F ��I����$�  ��G �싍�  ���  �=,G X��$   �5� G �58G ��$�  �
��G     P�=,G ��$$  �LG �=`G �8G ��$�  �5�G ;5PG �B���5�G 5�G �=,G �=�G ���$�  ��G Ǆ$�      ��  �=��F �=��F �=P�F ��3=��F )}�UԋU�+d�F ��F ��)��F ���F ���  3�F )��F ��F �M���3��F )��F �M�������d�    �d�    ��3  Ӯ�2  �DG ˁ%�G ��S灆�2  A&�� G ���2  +��2  � G 3��2  ��<  ��G ����G �02  +�G NT�=�G ��<  +��2  h�  ��  Ë �d
G �@��   ��	G ۋd
G J��  ��   ��  ��(  ��   �K  ���  ��Dj3�F 0�F �E    �E    ���F     ���F �I�5��F �,13l$�5x�F �5��F �4u    �5��F �   )��l$���E�   �΋=��F �E܋��F �3E�5��F �h  �=xG �� G ��$�  ��$�  ��$�  ��$�  ��$�  ��$�  �=�G ��$�  �=xG ��$�  ��$�  ��$�  ��$�  ��$�  ��$�  ��$�  �i��	G �l
G    ��	G �d
G �l
G ��(  ǅ      ǅ      ��(  ��	G ��   ��  ��d
G �K������P�����$�  ��$�  �=xG ��$�  �LG �=`G �� G ��$�  ��G ���������$�  ��$�  ����$�  �$�  ��A�A��$�  ��$�  ���������M����F ��)E�5��F 35��F )u�E���������=��F �=��F �=P�F ��3=��F )}�E�+d�F �E���)��F �UЋ��F ���  ��   ��   �% ���	؉A��$�  ��F  ��  �= G �d
G ��(  �=l
G �= G �l���=0�F �5�G Ή�8  ���F ���1  �5G 35�G AT���1  �΍��F ��4  �dG ȋ�P1  #TG ATqTPd�5    d�%    �8G �pG �3u�)5��F �}ԉ}���3=��F )=��F ���F +�  ���F +x�F ���F ��F �}ȋUЋMԋ=��F �M��F �M��m�����G ��  �PG � G �ʋ�G �=TG �=��F �9�I�=TG �  �X7E ���tP�l'G �X7E ���/  SV��QB �5X7E ���d'G ����uIh�   j� ������YYt-V�5X7E �h'G ��t�FT5E �F   �<QB �N���j����YS��QB ��^[�jhaB �����u3�;��  �F$;�tP�`���Y�F,;�tP�R���Y�F4;�tP�D���Y�F<;�tP�6���Y�FD;�tP�(���Y�FH;�tP����Y�FT=5E tP�	���Yj��/  Y�}��F`�E�;�t�u;��E tP�����Y�M���   j��/  Y�E�   �Fd�E�;�tM�9x,t�H,�	9x4t�H4�	9x0t�H0�	9x@t�H@�	�HL���   ;�3E t=�3E t98uP�j��Y�M���    V�b���Y�(���� 3��uj�.  YËuj�.  Y��d/  ��u����3��VWh aB ��QB ����tk�5�QB h<aB W��h0aB W�`'G ��hHaB W�d'G ��hTaB W�h'G �փ=d'G  �l'G u(�@QB �d'G ��QB �h'G ��QB �`'G /cA �l'G h�`A �`'G ����X7E tA3�h�   GW��������YYt+V�5X7E �h'G ��t�FT5E �~�<QB �N������A���3�_^��RB � W��G ��G �=TG ��G �T$�5�G ;5�G �a����5�G 5�G S��$  �|G Ǆ$�      ��  ����$�  ����=�G ��$�  ;=4�F ����=�G ��G R��G �|$���G �-�G ��G ��$�  ��G �\$���$�  �5�G �5TG �(����$G ��  ������ G ��  ��  ��H  $G ��G ��  �PG �xG ��  ��G 4� G ��  ��G ��H  ���  ��G ��@#  Ӆ0���ǅ$���|g ��  ����\  R�|G ���  ��  �ы�  ��0�����G ��G h�  jd�5t�F �  Ë�$�  ��$  �5�G ��$�  ��$�  ��G �(
G �-�G ��$�  �|G Z���@  �΁��   �   ���F ��@�C����G    ǅ(      �t֍��F ��(  ��G �?  ��(  �ڋ-�G �E$�$�  �m�$�  ��$�  ���  �[ �$�  �=TG �=�G �R��G �R���  ��G �I��G     �;����5�G �5�G �� pD �5��F �  �PG ��G B���   �C_��V� G ���F ��  �PG �A%�   =�   �����������$�  ��G ��$�  �-�G �-|G �E �������@G ��$�  ��$�  ����$�  �$�  �-@G A@G E��$�  ��$�  ��$�  �-�G ��$�  �<G ��   ��  ��G �ˋXG �=�G ǅ����|g �8G ��$P�G ��H  ���  �(G �ҋ�G ��H  ��H  ��G �5HG �5�G ��$������$�  ���%�G  ���	�G �-�G �/G�5t�F Pj
�5��F ��  �ǅH      �PG     � �]��G ��G ��h  �I�}   ��$�  ��$�  ��$�  �4	G �|G ��$�  ��$�  ��G ��$�  ��$�  �<G �D����(G �|G �E�    ��F �]�UԉpG ǃh      �� G �K<ًQ|�Yx� G ��������K�E؋C�EЋC�`G �S � G �5$G �s$5� G �G �K� G ��G �5�G ��G     �  ��$   ��G ����$�  ��X�(
G �-�G ��$�  �|G ��$�  ���u  �VC20XC00U���SVWU��]�E�@   ��   �E��E�E��E��C��s�{S�I������t{���t}�v�D��tYVU�k3�3�3�3�3���]^�]�t?xH�{S�������kVS������vj�D�������C�D�3�3�3�3�3��Ћ{�v�4�댸    �#�E�H�   �U�kj�S������]�   ]_^[��]�U�L$�)�AP�AP�����]� �pG �5�G F�E؉}���G �E����  �E���   ���  P�=�G �MЉ5G +}�G�ǋEЋU���   ���  ��G ���  �U�땉5$G ��$L  j �  �=�G ��G ��$  ��$   ��$L  �-�
G ��$  �ω(
G �=�G ��G ���%  ��d�    �d�    �$�F 3�  ���  �5��F wT���F ��_T���F Hmᶁ5��F �}���  ��F ��<  ��  \DNU��  ���F �� ��$�  �ߋ-�G ��$�  �։�$�  �=�G S�(
G �-@G �5�G �\$�|G [��������Ӊ}���G �}��(G �}Ћ�G �}������-\G ��G ��$  �-pG ��$�  X�54G ��$0  �=�G ��$  �΋�$�  �58G ��  �ϋuЋ��M��5�G �5p�F �7�h�F �5G P�E����F �0G �pG �=G �]��G �58�F �m���$�  ��G ��$�  �-G ��$�  �G ���  ����+  ��$  �-�G ��$$  ��$�  �G ��$(  �=�
G Ǆ$     ��G ��G �=|G �$G �hG �=�G �\G ��$(  ��$T  �58G ��G ��$  � X�=�G ��$�  X��G �5�G �E  �8�F �u�Ẻ5�G �UȉE��u��$G �EЋủ0G �Eĉ58�F �=�G �}؉}Љ�G �   ��dG �]���v!  �=�G ���G +�G ;G ������  �0G ��G �58�F �}̋M؋=G �G �M���G �=�G �   ������u��@G �M̋]ĉM��]Ћ-8�F �l$�<G ��G �T$ԉ��   �R�-0G �G �c  S���  �=G ��  ���  �xG �=�G [�=G �5�G ���\  ��G ��G ���LG �5�G P��G �|G ��$�  ��$  �0G ����  P�=�G ��$  �|G �5�G ��$<  ��G �D$�=�G �-,G ��G �5�G ��$�  �8G �I��  ��G �=�G ��$<  �LG �5�G ������E��Ӌ=�G �EЉ=(G ��G �}��}Ћ=�G ������(
G �   �D$�|g ��$�  ���58G V��$  �G �D$ �D$�=hG ��$�  �=�G �׺   ��$0  ��$0  ������-�G �M �� ���(
G PjP�5t�F ��   P�hG ��G �=,G ��$�  �5�G �G ��G ��$  ����G ��$4  ��G �|G �5�G �LG    ��G     �����G �=�G ��  �-hG ��$  ��G �=G ��$@  ��G ]��G �=,G �58G ���?����M E�G �D$(�\G � ��  �5�G ��R��G �5�G �xG ���  �5�G ��  ��  ���  �G �-�G ��G W�xG    �-hG ��G �=|G ��$(  �=�G ��G ]��G �xG ��   ��G �|G �hG �E ��$�  % ����dG hG ��$4  �E ��$�  EN�!����\$���$  ��G ��$�  �-pG �G ��G �5hG �-�G �hG �5(
G ������=�G �-�G ��G �-\G �D$��-G ��$  �G �5LG ��G ��G �5�G �F�������G �(
G ��$P  �\G �58G X�������0G �M؉58�F ��    �MЉG ��G �� G ;dG �X����=G ������@G �dG �-$G �T$���������=�G �=�G }�}���U���G �]��0G �M؋]ĉxG �]��G �=lG �EЋ=�G �E؉}ċ]��>�����G ��  ��G ��G �9  ��G �=xG �pG ��  ���  ��G ��H  X���  ǅ����|g ��  ��0�8G R�G ӄ$0  ��G �pG ��  ��  ��G ��  ��G h�  � ���Í��F ��   ��  �
�R�A��  ���   ��G ��$<  �|G �T$�-\G ��-�G % ���	��G��G �A���W�-�G ��G ��G �5(
G ��G �|$������  ���F ��   �5xG ǅ     ��L�����  ��t���F ���"  ������F ��G ��  � ��$�  �@�a����=xG    ��   ���F ���$  �7  ��   ���$    ��   ���$     ��  A�k����������U��WVS�M�tM�u�}�A�Z� �I �&
�t'
�t#����8�r8�w�8�r8�w�8�u��u�3�8�t	�����r�ً�[^_��AA��G ��  ��   ��G �xG ��G ��G ��  �5�G ��G �|G ��G �~   밋�G ��  ��   ��   ��  ��G ��G ��%  ��  ��   ��G ��  �|G ��   ��  ��xG ���G ���F J��  ������|G ��G �=0G ��G ��  ��   �|G �=0G ��  �=�G ��G ��G ��   �L���F ���&  ǅ     ��   �=�G ��b  ��  ����   ��G ���F �������G +�G ��   ��G ��$�  �ʋ�G ��  � G ��G ��G �G ��  �5 G ��   � G �=�G �=�G 󤋅  ��  �LG ��  �=�G ��G �5 G ��   ��  �2  ��   �=��F �TG ��I�@��G ��G ��x&  ��   �5�G �����@���dV����  ���F ���%  �(G ��  ��G �=�G ��G ��  ���5G �5(G �5�G �5G ��  ������  ��%  ��  ��	G ��G �LG ��  �|G ��	G �LG �  ��G ��G     ���  ��G ��  �=G �5�G �=�G �5�G ��  �=G �5�	G ��  ��   ���%  ��  ���!  ��   �-xG ���"  ����$�  ���&  ���$  �|
G �5�G ��G ��$�  ����   ��������F ��I�B��������$�  PǄ$�      P��$�  �T�F ��$$  �l$�E ����   ���F ��$�  �  G ���-  G   G �-��F A��F E��$�  �l$X��$�  ��   ���  ��G ���F �Jd  ���  ��b  ���  �Re  �XG    ��G     ��W  ��G ��XG �W�  ��G �܉�$�  ��$�  ����T�F ��$�  ;��F �CD���T�F ��$�  ��$�  ��$�  ��$�  ���F ��$�  �� G ��$�  �t$��$�  �G �=G ��$�  ��$�  �(  ��$   ��$�  �D$��=dG ��$�  ��$�  �=dG �b�����G ���F ���%  ���#  �$�  ���   �% ���	ЉG��G ��  �=$G ��  ��G �=�	G ��  �PG ��G ��	G �PG �=$G �R�����(  �ǅ      ��F �=�
G ��
G    ǅ      ��	G     ��  ��  �=dG �5(�F ��  ��  ��������F ��I�B���������$�  ��$�  ��G � G ��$$  ��$�  ��$�  ��$�  ��$�  ��$�  ��$�  �G �=G ���F ��$�  ��$�  ��$$  �t$��$�  ���Q���F ��I�B���������F ��I�B���]�����  ���F ��I�B��  �5�G ������V��$�  �=G ��$�  ��$�  �5�G �T�F ��$�  ��$�  ��$�  �G ��$�  ��$�  ��$�  ;T$ ��$  �J?����$�  ��$�  �$�  ��$�  ��$�  R�$�  ��������
  E�����
  ���
  `�F ���F �d�F ӎ�
  0�F ���
  ӆ�	  ��0  ���F +�F �<�F Ӯ�	  �5��F 54�F ���F ���F ���F +�	  ���	  35��F �-��F �ߝ�3��  YT�<�F ���F ���F ���F ��`  �������	  HT��,  ���
  �D�F ���
  ���  ���  �=��F � ��h  �xG �B�$�  �-xG �R$�$�  �xG �[ �$�  �5�G �5xG �m�=xG �v���  �IǄ$�      P�5`�F h�  h�  ������5����T  ��D  ��
  ӊ�
  ��F     j ��F �=�F    ��  �5��F ��F W��<������@  �FT��l  ��  R��H  ��QB ��T  0�F ���
  ﾭ����
  h�  jSjP��������   ��,  �A�=d�F �yR���  ���  �Q�=��F �y�=l�F �y�p�F     ���F ���F �0�F �$�F ���F ���F ���F ��F ���  ���  ���  ���  ���  �5��F ���  ���F ���F �=��F �@�F �`�F ��$�  �-�F �5��F ��$|  ��$x  ��$t  �  �}��5HG �5�G 5G 5G ����0G �0G �5tG �M��E܋5HG �E̋U��0G �uȋ]�u܋��   �M���x  �}���  �0�F     j �0�F �=0�F    ��  ���F ��H  ��x	  ^���  1�v���F Ӣ�
  ���F 3��  �-��F w��#��$�  �t�F ���F ˉ(�F ���
  �F ��0  =0�F ��L  0�F �W�����$p  ��$l  ��$h  ��$d  ���F ��F �=��F �-��F �5��F ���F ���F ��$`  ��$\  ��$X  ��$P  ��$L  ��$H  ��$D  � �F ���F �5��F �-��F �`�F �H�F �=|�F ��$@  ��$<  ��$8  ��$4  ��$0  ��$,  ��$$  �5|�F ���F ���F ���F �-��F ���F �=�F ��$   ��$  ��$  ��$  ��   ��F ^���H  ��@  �vV��H  �<�����H  Z�
�=��F 1:�RR� ������F �=��F ��  Z�:��@  ��D  �R�=T�F ω�0  �������F �=G �E�5�G �u���   ��x  �G<��H|�px����ev���=��F �F�~�}��~�u܋v �}؉Uԉ�G �E��  �]��=G �'��$  ��$  ��  �0G �5HG �M��  ��F ��G �M���G A)U��E��E��G �LG ��G �u��]��5�F �8�F �u��}����  �=�F V�M��M�����  �5L�F ��l  ���  ��t  �5��F �  �=lG �z���   �r��G �J�58G �r�dG �B�5�G �=�G �M��m��\$��5�G �=�G �xG �-<G ��G �%8G �Ƌߋ�5<G �=�G É=�G �Mԍ�    �MЉXG �]ȋ]܋�G �LG �]���   ��x  LG 95LG ��|���u��v�l$��T$�싊�   ���1  $�L~��d1  0�F ���1  �xG 3�G YT�u����1  ���   ���2  �}���@  ���   ��@  ���   ��@  �������   ���]��G �UЃ�G �XG �Eā}�   ��u���=�G ��G �]ȋ}ԉ}���G �Mԉu��5LG �Eȉp �@�؋u���  �   �����}ԉE܉=�G �EЉ]ȉXG ��E�+E�;�G ��t�������}��5tG �5��F �7�h�F �u�P�E����F �G �u��M��LG �]��M���G �E����  �������   ��x  ��űu܋F��]Ћ]܋S$��=��F ��G �]��E�    ���	  �]ȉ�80  �$���U��Q�E�H��   �Mw	�IH�A�TV����W�yH���Dw�_^tj�E��U��E� X�
�E�3��E� @j�q�q�MQP�E�Pj��2������u���E#E��V�t$����   �F�h3E ;At;D3E tP�#���Y�F�h3E ;At;H3E tP����Y�F�h3E ;At;L3E tP�����Y�F�h3E ;At;P3E tP�����Y�F�h3E ;At;T3E tP����Y�F �h3E ;A t;X3E tP����Y�v$�h3E ;p$t;5\3E tV�v���Y^Ë�$�  ��$0  ��$(  ��$   _���F �D�F �8�F �-P�F �5��F �(�F �=x�F �%0�F �p�F ���F �-��F �50�F �=$�F �Ę  Ë�$   �-�F ��F �t�F �5 �F ���F �=��F �X�F ��$�  ��$�  �J���jhcB �B���3�95<*G u'j�  Y�u�95<*G u�   �<*G �M���   �G����j�  Y�jhcB �����3��}�j�R  Y�}���%G �]؉=4*G �,9E �� 9E �h�bB �70��Y���u�;���   �> ��   �8*G ;�t!PV���YY����  �8*G ;�tP�����YV����@P�D��YY�8*G ;��d  VP�+���YY�M���i  jV�59E �������9E �@ ���>-u�E�   FV��j��Yi�  ��8E �0�<+t:��&  <9�  F��8*G ;�tP�Y���Y�=8*G h�)G �dQB �����   3�A�4*G ��)G k�<��8E f9=�)G t��)G k�<£�8E f9="*G t�0*G ;�t��8E +�)G k�<��8E ��=�8E �=�8E �E�PWj?�59E j�h�)G WS�5xQB �օ�t9}�u�9E �@? ��9E �  �E�PWj?�59E j�h�)G WS�օ�t9}�u�9E �@? ��9E �  j��E�P����YY�   �u�3�j�  YÀ>:u>FV�i��Yk�<�8E �<9F�:�}��>:uFV�li��Y�8E �<9F�:�}�9}�t��8E ���8E ;�tjV�59E ��������9E �@ ��9E �  ����É��F ���  ���F �L�F ����  �l�F ��t  ��F ���-�F �F ��A�B�<�F ���  ���F ���F �l�F ���F ��l  �5��F ���  �5<�F ��p  �������$�  ��$�  ��5��F ���F     ���  �D�F ���  ��x  �=��F ;�$�  �W����=��F =��F �T�F ��8�F �L�F ǅt      ������ϋm���   ��G ��x  ��G �D$���������`�F ��$t  ������  ���F ��t  ;�$�  �K��������F ���  ���F ���F �D�F ���F ��t  �T�F ���  ��l  ���  ���F ��������58�F �-  �PG ���  ���  �$�  9��t?  ���  �8�F ��G ��  �PG ���  ��G ���  � ;��F ��>  ��G ��$�  ��  �<G ���  ��  ��I���?  ��G �G ���  �G 뉍��F ��I�@���W  ��I�B���&  V�t$��tT��h3E ;t;83E tP����Y�F�h3E ;At;<3E tP����Y�v�h3E ;pt;5@3E tV�ֿ��Y^É}Љ58�F �UċU������  �}̉=HG ���m�}̃�A��E؉}��LG �}ЋUċU��DG �Uĉ�G �M̉M��u��ű�G �[����E�    �0G �}Љ58�F 9E��X����M��M�M���G �Eȉ@G ȋ� G �U��E�    �A�����������  �(	G    ǅL      ��������L  ��(	G ��  ��L  �܉��F ���F 0�F �$�F ���F ���F +��F ��   �u����T  ��QB ���F ���  KP��F �l�F �%��F ���F ��T  0�F �5��F 3�,  ��X  ϋ�l  ӊ�  zT��vQAWd�5    d�%    ���  ��X  �S�0QB V�86E W�>��t�~tW��W�����& Y����X7E |ܾ86E _���t	�~uP�Ӄ���X7E |�^[�U��E�4�86E �XQB ]�jh�`B �,����u�4�86E 3�9urj�<��Y��;�u�b����    �?j
�b   Y�]�9u8h�  W��  YY��u#W�J����/����    j��E�P�_�����3���>�W�#���Y�M���	   3�@�ݺ���j
�M���Y�U��EV�4�86E �> uP�G�����Yuj����Y�6��QB ^]�VW3��&G �<�<6E u��86E �8h�  �0���!  ��YYtF��$|�3�@_^Ã$�86E  3���\  ���F �`�F ���F ��h  �@�F �@�F �%��F �(�F ���F �h  �5@�F ΁��  ��du�5��F p��sT-���ˉ�X  � �F #�T  ���  0�F ��$�  ��<  ��L  ���@  �I�@���HG �  �=�G �e�����}�;;�����=�G �E��U��}Љ�G �0G ��G �>����=�G J���  ��L  ��4  ��G ��G ��<  ��D  � % ����$  � G ��D  �B��4  ��D  ��0  � G �C  ���F ǅL     ��L  �PG ��L  ǅ@     �HG     ��L  �HG ��8  ���@  �������<  ��@  ��L  ��@  ��G ���8  ��G ������G �HG ��G ��@  ��G �jh�ZB �����T%G ��u7�=�%G t$h�ZB ��QB ��th�ZB P��QB �T%G ��u
���A �T%G �e� �u�u�ЉE��$�E� � �E�3�@Ëe�}�  �uj��QB 3��M���̷����t$��QB 3�@� ��<  ��L  ��8  ������<  ����G ��G ��8  ����PT���1  Ue���1  U�d�5�G Y�Ⱥ�XG �`G 3DG ��8  ���F ȉ��1  ���1  +G ��4  ��|3  50�F q�<A0�F ��G JT��0  ��G ӊ�1  ��,  ���1  50�F Vd�5    d�%    ��D  ��G ���<  ���xG ��$   �����G 	�$  ��G ��4  ��D  �9A��0  ���xG �5h	G ��8  ��0  ��D  �5h	G �g�����d�    �d�    ��@  ���F �-�G ���1  6���,G ӈH2  ��X3  �G �XG ��G ӀH2  ��h1  	�DG �ڞ���D2  Ӏh1  ��<  �=DG =0�F ��H2  Qh�  h�  �<���Ë5�G �E��%DG ����EЉ]��DG ��G ;�  �E��E���G ��G ��G ��E�    �EЉMԉ�G �U�;U�������U�U���G �]ȉ]�Ӌ�G �lG �DG     �x�]��lG �]��DG �M��aR�tG W�,G �5�G �=PG ��H  R��  ���������  ��G ��G _�,G �=`G �=PG ��G �.  ��G �MԋEЉ5�G �5lG ���������U��DG �U����m�U���A�F�u���G �G �5�G �U���G ��G �]��M�������$  �-�G �5�G ��$@  ��|G �:����D$��$@  �=dG �=|G �=�G �-|G �=dG ��G �5�G ������   �7  ��$  �PG �-�G �5�G ��G ��$<  �|G �K�����D$S��$@  �-|G �PG X������   ��  P��G �tG ������=PG Y������5�G ��v�@��H  �5�G �=|G ��G X��H  �5�G ������=|G �PG �����W������LG ������|G �G ��G �����Y�-|G �-�G �5�G ��v�@��$  �LG �5�G �-�G �D$��$  �5�G ��$@  �D$�D$�G���������$G ��G �`G ���l  W��G �5�G �=PG �������G ��  Y����  ��H  �G �8G ��G �ы�G S�8G ��H  �G �`G ��G �v��H  �G ��G ���  ��  �щ=$G �������H  ��G ��  ��G ������8G ��G ��G P��G ��  ��G �d  ��  �|G �5�G �������G �`G �-|G �W������|G ��
G ��G ���   �%|G P� G     ���5 G ��H  �5�G ���n�=0G �5�G ��  �5�G ��G    �������G ^�$G ����   ��G �
�R�A��G �G ��  �G �|G �  P��H  �5G ������5|G W�5�G ��  ��c����=�G �������_��G ��G ��$<  �5G �|$�|$��f���������$G ��G �`G ���!�=$G ��G �5�G ������������P��G �5�G ������$G �tG ��  �|G �������M���P�=PG �tG ��������PG Z������������G �tG �"���j����Y�j�����Y�V������t�Ѓ�;t$r�^á�BF ��t�t$��YVW��.G �/G 3�;ϋ�s��u?���t�у�;�r��u,h�KA �����.G �ƿ�.G ;�Ys���t�Ѓ�;�r�3�_^�jh�\B 貮��j����Y3��}�3�F95&G u�u��QB P�pQB �5&G �E� &G 9}u79=CF t�0�B ���0�B ;CF r
� ;�t�����h/G �/G ����Yh/G �/G �����Y�M���   9}u!�5&G �u�Y   3�3�F9}tj����Y��7����j j �t$�0������j j�t$�������jj j �������jjj �������h�\B ��QB ��th�\B P��QB ��t�t$���t$�RB ̋=0G �5�G ��  �=�G �$G    ^������=0G ��H  �$G �$G ��H  �{����5�G ��G �� �����  ��G �|G ��G ��G ��  �|G ��H  ��G ��[�@��  ��G ��  ��G ��H  �`G ��G ��  ��G ��H  �5�G V�5�G �S  �G �|G �,G ��G _�G �=`G �� �����G ��[�@��  �pG �=PG �5�G �,G �� ����5�G �pG ��  �����j�G     �����V��G ��  �5@G �������G ��  �|G �@G ��M����5G �J�B���P�����������5G ��G X^��G �@G ��G 냉��  ��
G ��
G �5`
G ��G �5�	G ���  ��G �-�
G �E �m�@��$�  �ŋ�$�  ���Y  ��  �|G �5�G �5�����G �`G �-|G �������|G ��G ��
G �(G ���   PǅH      ���%|G ��G ���=xG ��H  W�=xG �e������  ���  ���  �
G �TG ��	G ���  ���  ��G ��  ��	G �TG ���  ��
G �5p
G �5�G ���  �F�
G ���F ���"  ���  ���"  ��"  ���  �5
G ��	G ���   ��
G    ��G ��  �`
G ��	G ����  �Q�����G ��  �
G ���  �`
G �=�G ���  ��	G ���  ��
G ��t�^  ���  ��	G �
G ���  ��	G ��	G �=�G ���  ���  ��v�@���  ��
G ��	G �5�
G �  ��G ��  �HG ���  ���  �   �5�G C�5p
G ���  ��  ���  ��B�5�G �t
G ���  ��	G �HG ��G �t
G �G ��G ���   �|  �-@G ���G ��G �� @ j j �E�P@=�  �������F S���
  P�E���E�%�   =�   ��  �   � �d
G �@��	G �d
G �5�	G �j  ��G �=p
G ��  ���  ��	G �c������  ���  �
G ��   ��������  ���7  }e�p
G �=
G   ���  �]  �
G ��   �	  ���   �  E����F ��G �5�G �u��]��5�G ��������5�G �ڋ
G �HG ��  �5p
G �Y�����   ���F K�"  ���"  ���   �QN����G ��   ��	G �G �(G �G ��8  ��(  �=(G �=
G ��(  ��  ��   ��
G ��(  ��G �50G ��   ��  ��0  �0G �58
G �B  ���-  �]�X��G ���
  �=�G ���
  �u�u���v�u��=�G �u����������  ���  ��	G �
G ��G ���  �G �
G ���   ������=��F �(�@�E��$  �식  ��  B��G ��G ��G ��(  ��  ���   �����X
G ��	G ��d
G �s�����	G �a�����   ��
G ��G �ދ58
G �4  �5�
G ��
G �5�	G ���  ��
G ��
G ���  ��
G �6  ��(  ���F ��@�B�,
G �58
G ��(  �,
G ��  �x
G ���F �$  ���   ��� ���	�A��   ��  �5�
G �x
G ��(  �58
G ��  �p	G ��	G ��  �p	G �x
G ��  �U  �=�
G �ǅ8     ���F �
G �hG    ǅ0      �p	G     ��$  �P
G ��G ���F ��G ��(  ��   �=8G �=��F ��
G ǅ�     ��  ��
G ���   �5��F ���  ��������=��F ��G �=8G ��  �5�
G ���  �M����5�
G ��
G ��
G �5�	G �
G ��  ���  ��
G ���   �  ��(  ��	G ǅ       �5�G ��G �58
G �p	G ��   ��0  ��G �58
G �������58
G �5��F ��  ���  ��t�����  ���  �0�@�F����������"  ���   �x
G ��(  ��   �0
G �-p	G �މ-�
G �G �p	G ��	G ���50
G ����   ������)G ��t��u*�=`7E u!h�   �   �&G ��Yt��h�   �   Y�U��$t�����  �(3E ���   SV���   3�W3�;Š5E t@��r����;��5E �  ��)G ����   ;�u�=`7E ��   ���   ��   h  �E�PR���   �LQB ��u�E�h�^B P����YY�}���P�a��@��<Yv"��P�a�����E���;j�h�^B W�4�����W�{a�����5E ���na���DY��Y����=����h�`B S���WS���h�`B S�~�����5E S�r��h  h�`B S�%����,�(R���   P���5E �6�a��YP�6j�� RB P��QB ��t������   ����_^[�Ō   �ÉG ���F ��G ��("  ��	G ��(  ��=8G ��8  ��
G ��	G    ��8  �<G ��   ��G �ȋ�	G �=<G ��(  �=�
G �G �ށ��   �a���������5��F �0�@�F������	G    ǅ(      ��   ��G ���F ��(  ���	G �u%����G ��(  �ʉ�	G ���F �R����?  ��(  �
G ��	G +
G ��8  ��	G ����G ��  �=�	G ��8  �=�	G ��   �=�	G ��8  ��G �ȋ5�G 󤉽  ��   ��  �5�
G �=�	G ��  �58
G �k  ��
G ��G ��	G ��   ��  �58
G �hG ��  ������0�@�F����������F ��@�C��   ���F ���"  ��   �������F �u��u�5��F ��3�l  )�+��F �U���)U�\�F 3E�)E�]��4�F ��3H�F )]�]��]�+��F �=��F ��ً=
G �=
G ���  ���   �����=H�F +}ċ��F �M����I��F �M��5�F ���v���y  �&4  �U؉E �M��5 �F �=0�F �]��=��F �]ĉ�F ���F ��F �u��  ��G ��  �l	G ��   ��  �������  ��$�  ����=LG ���  ���  �(G ;;��  �=LG ��$�  ���  ��G ��G ���  �
ǅ�      ��G ���  ���  ;�$�  �i����$�  �$�  �(G ��G ���  �����  ǅ�      ��G ���  ���  �
���*������  ���  ���  ����$�  �$�  ��A�B�dG ���  ���  ���  ���  ��G ���  �5dG ���  ���  ���  ���  �@G �<���U��WVS�M�'�ً}��3����ˋ��u�F�3�:G�wt���ы�[^_�É��  ���  ��G ������L  �@=   ���  ��G ǅ@      �=(	G �@	G ��<  ǅ8     ��@  �X	G ��  ���F ��G �J<ыQ|�U؋Qx�G �������=�G �=��F �J�z��G �J�UԋR �G �}̉�G �MԋI�G �   �E     � �F     �E�    � �F �]�[��F ��F �MčM    �u��5��F �=��F �U؋��F �3U�   ���E�   ��l  ���e����F ���F �u�3E �%��F �5�G �EЋEԋ@$�G �=�F �E��E�    �=�G �E�Eȉ�G �Uȉ|G �=�G �EЋUԋ=�G ��G �M���F �MԸ   ���G ��r����E����G +�G ;�G �̽����  �M��E���)]���   ���  3]�)ڋE����3����u��u�5��F ��35H�F )�+��F �U����%��F �<	G ��G ��8  ��<  ��L  ��  ��G ��L  �<	G ��G ��P  �X	G �O��  ��@  �5 G ��8  ��G ��L  ��<  �5G ��L  �ˋ�@  �5 G �X	G ��  � G �}ԋ}��  �5��F �7�h�F �u�P��G ���F �5�G ��G �=�G �U��]��,G ��G � G �E��8�F �E��-hG ��$�  ��$|  �,G ��$�  ���  ����c  �]ԉ]��G ��G �EԋG ��F �|G ������=�G �,G �(G �U��  ��F Ӌl  �L�F ��l  0�F =0�F ���  #��  ��p  5j���-��F )Z7��F �KT�����X�F �<G B�<G +E�@�E��E��= G �U��5�G �=�G �U��5X�F �u��X�F ���  P�M��M��u����5�G �M��{����<	G ��L  �	��P  ��$  �A��G ��G ��<  ��G �����E��e��EЉ]��]��}��}ԋ�G 9���+  �G �Mԉ=�G �EЋ}��E��E��}�   �"����}���G ��G �u��Uȋu��5�G �]��G ��G ��h  �@�u��M��3����EЋ]�]�]����G �U���G ��G �F���)U�\�F 3E�)E�U���F ��3H�F )U�U��U�+��F ���F �H�F +UĉH�F ���F �M��u��U��,����G �t����=��F �-��F Pԉ�8  � �F OT�M̋��F �-\�F ��0  0�F ���  ���  3=x�F �H�F ���F 3��  ��P  ӣ  �Eȋ�  3�T  �%`�F �|G �I��   �ō���G �\G     �lG ��  �\G j�\G �G ��H  �G ��G [��  ��G ���  V��H  �5�G ��  ��	G W�=�G ���@P�=�G ��  �����^�;  ��$�  �쉽�  �5lG ^�n�$�  �L$���$�  �\$��K$�$�  �<G �G �D$��@ �$�  ��$�  �8�F ����F � G     �5 G ;�$�  ��������F ��4  5 G P���$�  ���  ���F ��\  ǅ�      ��   ���F �TG B����G �TG ��G )�C�Ë�G ���  �=��F ���  ���  �����F R��G �ȉ5�G �5�G 󤉵�  �lG ��  ��	G P��  �|G ��G �=�G ��  ��H  �J�e���X�� �����  ��  �=�G ��G �� �����H  �=�G ����   ���  ��G ������G �8G �	����  ���  ���  ����$�  �$�  ��A��8G ��G ���  ���  ���  ���  �8G ���  ��G ���  ��  �|G �I��   ����QǅH      �HG ��  ǅ     ��H  P��G ��	G ��  ��  ���  �|G �"�����	G ��G ��  �|G ��G ��H  ��  �J�f�����  ��G Q��  ��	G ��G �=�G _��H  �=�G �j������  � �F ���QB ��$�  P�xG ��QB ���  �xG ���  �G �5�G �4G ���  �G �����   ��  ��G ��G ��G ��$�  ����G h�  �5t�F �58�F h�  h�  �  �� G �5�G ����<  �5<G V���-<G 5<G ��A���G �5(G ��$�  �DG �� G �<G Q�5<G �DG ���V�H�F �,G ��G �h�F �5��F ���  �h�F �5��F �LG �h�F �}��=�G ����  ���  ���  ����$�  �$�  ��A� ���F ��$�  ������  ���  ;�$<  �M�����4  � G ;�$�  � ���� G  G ���  Z���  �$�  ��$�  ��G ǅ�      �  X���  ���  ���  ��G ���  ���  ���  ��G �o  �� G ��$�  ��$�  � G ;�$�  ����� G  G ��$�  ��$�  ͋U �$  ��G �<G     � ����F ���  �58G ǅ�      ���  ���  ���  ���,  �   ��g?����G �54G ����  �4G +|G ;0G ��  �,G �%,G ��G �G �,G ��;�$�  �4  ���   �[��$�  ��$�     ��  ��G ���  ��G �54G �G �dG �4G �5�G ���  �@���dG ���   �)����5h�F ���50�F �O����G���  ��G �-,G R�=�G ��$�  ��$�  ��$�  ��G ��$�  �5�G ��$�  Z��G ��$�  ��$�  �-LG ��G ��$�  �=| G ��$�  �-,G ��G ��G �G �|$�<G ��$�  ���4������  ���  ��G ���  �}���$�  �����G �G ���  ���  �� G �| G �-LG ��$�  ��$�  ;�$P  �W�����G � G jZj
�5��F ����Ã��%<G ����$G �<G ;�$H  ������-�G � G ���G ��G �5�G S���  �$G �,G �� G ��$�  ��$�  �5<G Y��������  �=�G ǅ�      ���  �=�G �Gh    ���  �F<��H|�Xx����  �=��F �C�s�k�{ �$�  ��G �S$�$�  �0G �C�$�  �-|G ��G �������  �5G �Fh�v뇍=��F ��  ��G �	��G �A��D  ��G � G �  ���  ��G ���   ��������  �= G ���  ���  ���  �=8G �`G ���  ��G �$G ���  ���   ���������0  ��8  �5�
G ��(  ��	G �=�G ��G ��(  ��0  �=�G �=G ��(  �+  ��G ��G |G |G ����  ���  �=TG ���  �5|G �G �54G ���  ���   �����G �5�G ���  ���  ����G �=pG �-$G ��$�  ��$�  ��$�  ����$�  ����   �������8  ��G � ��G �@��
G ��8  ��
G �P�=�G �=��F ��G ���G �B��  ������=��F ����ǅ<     � G     �t��= G ���$  ��B���= G �߉�<  ����
G ��	G ��4  ��8  ��G �=�
G ��0  ��4  ��	G ��0  �  ��<  ���F �
�R�A��8  ��<  ��8  �y  �,G ��G �D
G ��8  ��<  ��	G �= 
G �h
G ��G ��R�@�   �)  �,G ��8  �5|	G ��0  �= 
G ��<  ��
G �5�	G ��
G �5D
G �,G ��0  ��(  ��G �5|	G ��<  �=�
G �Q  ��	G ��G ��<  @��(  ��0  �5�	G �5�	G �5�
G �5�	G ��  ��G ��G ��0  ��(  �;����,G ��8  �@
G ��   ��<  ��
G }���(  ��0  ���7  ��  ��  �6  ��   G@��G ��
G �B�����\����$w���������$	G ���F ���  ��H   ��������	G ��8  �}  ��<  �=��F ��<  ��8  ��G ���G �B��	G ��  ���F 	�� 
G ǅ0     �t{��0  ����������F ��$"  ��8  �=H
G ��<  ��G �=D
G �=�	G ��8  � G �= 
G �,G ��G ��(  �H
G ��8  ��(  �l������F ��G ��I�@��G ���d�����0  ���F ��$  ��<  ��y  ��F  �L
G ��0  ��G ������<  @�G ��8  ��	G ��0  �=G ��<  ��0  ���8  ���F O�=  ��w  ��$  �Љ�	G )��Ћ�$  �=�	G ��(  �=�G ��	G �=PG �x	G ��0  �ȉ�$  �����
G ��G �ǉ5�
G ��(  ��0  ��$  ��8  ������@  ���G    ���F �LG ��G    ǅ4      ��G     ��,  ��<  ��G �=��F ��8  ��0  �]����xG ��(  �5$
G ��	G     ��
G ��G ��0  �5�	G �5�G ��	G ��(  ��4  ��G �5$
G � ����5�	G �5��F �=�G ǆ�"     ��<  �tq�5�G ��������	G ���F ��   ��G �|G ��0  ��<  ��	G �5�	G �=�G ��8  �|G ��0  ����<  �5�	G �,����5��F ��@"  ���  �	���  �A��<  �G ��<  �Z�����   ���  ��I�@�G ����   ��  �G ��G ��  �H�����	G �5�G ������	G ��8  ������<  ���F ��$  ����M  �=lG ���"  ��8  ��0  �=t	G ��   ��	G �K����5��F ��(  ǅ       �=p	G ���"  ���  �5��F ��   ��p	G �=�����   �֋���$�  �-dG �5��F �-\G �pG ��$�  ���-  ��8  ��G �5�
G ��0  �5�G ��8  �5�G ��G ��0  ��
G �5�
G ��<  ��G ��
G ���8  ���F �$  ���   ��8  ��0  �<
G ��G ��G ��(  �-�G �-�G ��$  ��G � % ���	��C�<
G ��$�  �=�	G �Ë�$  ��$  ����   �%����_�����`  ��F �$�  9���&���� G ��X  �8�F ��\  ��G �\�F ���F ��\  ���  �� G � ;��F �%���� G J���6&���  �5��F �0�@�F���9�����G �5\G ��    ��  �PG ��G ��;�$�  ������  �PG ��$�  ��G �   ��$�     �=M����G ���  ��G ���  �5dG �-�G �=G ��$�  ��$�  �-�G ��G �   ��$�  ��$�  �G ��G ��  �[��$�  �v����=LG �TG �$�  �$�  ��PG ���  ���  ��G ���  �(G ��G ���  �\G ���  ���   ����󤋔$�  ���QB �5G P��G ���F ��G ��$�  ��$�  �5�G ��G ��$�  �5(G ��G ��$�  ������   ������G ��G �=G ��G ��G �=��F �\G ��G ���  ���  �   ��pG ��G �   ��������   ���G +�G ;pG ��O���������G ���  ��  �   ��$�  �R���-  ��$�  �^�-�G �쉕�  ���F �TG �=�G ǅ�      ���  �=�G ���/  ���  �	�����G �� G �
;��F �%"��B��G ��G ����"������ G ���ĉ�G ��G ���  �<������F ���  ��G C�G ��G +�$�  A����$�  �PG �G �-��F ��G ��$�  ���F ��P�\G �5(G ��$�  ��$�  ��������dG �4G ���  �@�a  ��G ���  ���  ��G ��G �	���!  ���  ���  ���  ����$�  �$�  ��$�  A�$�  ��G �`G ��G ��G ���  �`G ��G ���  �  ���  ���F ǅ�      ���  ��G 9�$�  ���  �g����G ���  �=pG ���  ���  ��$�  �$�  ��G � G ��G �G ��F ��G ǅ�      ������=��F �=x�F ���  ��G     �=�G ��G ���  ǁ�      �=��F �G<��H|�Xx����dJ�����  ���F ���  �E$�	  �m-��F ��$�  ��$�  �I ��F ��$�  ���G ��������  ���  ��G ���  ��G ���4G ���  ��G ���  ��G ���  �4G ���   �6������  ���  �=`G ���  ��G ���  �������   ��$�  ������  ;8�h  ��$�  ���  ���  ���  ���  ��G �G ���  ��G ��G ���  �pG ���   �������$�  ��$�  ����F ��G ���  �� G �K�$�  ǅ�      �5G ���  ;�$�  �������$�  �$�  ��$  ���  ��G ��(�$�  �-��F �쉅�  ���F ���  ��G     ��  ��8  ��   �=hG ���  ���  ���  ���  �|G �5�G ���  ���  ���  ��G ���   �������  �=G �%�G �����$  �5�G ;5t�F ������5|G ��$�  ���F �5G ���  ���  ���  ��G ���  �` G �=G ��������  ��$  �` G �5|G ���  �=G �=��F ����U����=�G �=(G ���-�G =�G ��A����F �` G ���  �=|G ���  ��G �pG �=�G �=G �o����=��F Ǉ      ǅL      �t����=��F �9�I�G��L  ���G ��`  �hG �ǉ�D  �hG ��L  ��D  봍��F ���  ��[�@��G ���   �=��F ��p"  ���  �6���  �F�֋�p"  ��=��F ǅ<     �tč=��F ��<  ���@  ��   ���R���O�@
G ��G � 
G ���   �D
G ���F ��<  ����ǅ8      ��=�����8  �I�}�����8  ��LG ��G �$�  �8G ��G ��   �tG �LG ��G ��G ��F �(G ��G ��  �=xG ��  9�8G �tG ��G �B  ��<  ��������  ���  �=�G ���  �=G ���  � G ���  �   ���  ���  ���  ���  �=G ���  ���  � G ���  �i���  �   ���  �$�  ���  ���  �[���  �D�=�G �=��F ��D*  �|G Ǉ8*      �5��F ��G �50G ���  ǁ�      ��F �C<؋H|�Xx�F ��������5��F �C�s�{�k -�F �- G �k$-�F ��$�  �K�F �-�G �4G ����F ��   �5XG �5��F ��8  ���  �	��G �A��0  �5XG ��8  ��0  �����D$ȋ\$ċL$��T$��l$��=P�F �5��F �<�F ���F ��F ��F �-\�F �L$��D$��T$��l$��|$��\$��t$�� �F ���F ���F �-��F �=��F ��F �5��F �T$��L$��$�F ���F �%��F � �F ���F �-��F �5|�F �=��F Ë��  ���  �$G     �pG ��G ���  �    ��~����8G ���  ���  �pG ���  ���  � ��G )�;4G ��������  �8G ��G ���  �G ���  ���  ���  ���   �_  �����@G ��G ��  - @ ��  �=��F ǇL*      ǅ      �=(G ��  G��$   �*�����G �8G ��F ��G �(G �C%�   =�   t������-@G �  �8G ��G �=(G ��F ��F ���ߋ��=(G ��F ������G �ȋ�$�  ��󤉌$�  ���F ��0G ��QB �5TG P�xG ��QB ��G �5�G ��$�  ��G ��$�  ������   �U��G ���  �G��G �$�  �$�  �:���  �<�    ���  ���  ��G ��F 9���8����$�  �$G �=$G    ��������  ���  ���  �$G �\G ���  ���  ��G ���  �pG ���  �5G ���  �Vh�v�֋\G ���  ���   �d������F �=�G G�؉=TG �=�G ��$�  )�G�ǉ5hG ��$�  ��$�  ��G ��$�  ��$�  ���F �G �-��F ��R�H���5(�F �Mċ��  �M��`  �u���L  �  �u��u�+��  �|�F Ӏx  50�F ��x  ɉ�\  ��p  �%��F �E�+��F �=��F ���  3=H�F ���F ���4�F �%8�F ��F ���F �]���F XT�]���\  ��F �=��F �}�E�U��U��}����   ���F �u����   ���   ���  ���  ���  �H���  �x���F �P�-��F �h��,  �H����F ǀD      ���F �=��F �u�M����F ���  ���  ���F �U��E�M�u�}܋m؋\$ԉd�F ���F ���F �5��F �=l�F �-��F ���F �|$Ћt$��m����5��F �HG ��  �	��$�  �A�ыHG �  ��	G ��  ��   �=�	G �=��F ��  ��I�B�=�	G ��  ��  ��	G ��  ��   �E���F ^��,�F �]�)�v���F ���F 0�F �M���F ���F ���  �%��F ��t  #��F ���F ���F +�  �����ދ��  �d������F ��I�B����  ��  ��I�@����  ���F ǅ     ��m  ��  ���������	G ���F ������-�	G �ř����	G ��
G ��  ���   �5�G �5��F ��  ���%�	G ǅ      ��G ��Q����5��F ��  �I�*�����G ��  �ω�$�  �%G ����G ��$�  �G ;��F �M�������$�  �5hG ��$�  ��$�  �=�G ���Ǆ$�      �=�G 9�$�  ��$�  ������G ��$�  ��$�  �$�  ��$�  ��$�  ��$�  :�$�  ��$�  �G     �w  ��I�B���������F ��	G ��G     ��  ��3�����  ���F ��G ���	G ������|G ��  ��  �|G ��G ��  벋=�G ��$�  ��$�  ��$�  ��$�  ��$�  ��$�  �G ��$�  ��G �G ��$�  �8G �   �Eԉ=hG �EЋ}��=8�F �lG �U��(G �;��F ������ G �}�B�EЉ}�O�Mԅ��8����u���G ���"  ���F �|G    ǅ      ���������F ��  ��|G �������  �։�$�  ��$�  �G ��$�  �8G �5hG ��$�  ���������$�  �G ��$�  ���-G G ��A�F��$�  ��G ��$�  ��$�  �5hG ��$�  ��$�  �k����(G �Mԉ=�G �EЋ}��U�U�9(G �������G �8�F �(G �E��G �����5 G �U��5�G �u���G �=hG �(G �U��S����=��F �9�I�G����  ��G ��  �=�G �5|G �XG ��G ��   _[������  ��G FǅH      �G W��  �5|G �XG �=�G ^���  �lG ��H  ��|G �[��P��  ��H  �lG ��  ǅ����|g �58G ��0V�G ��  ��G ���  � G �Ӌ�G �G ��  �=G �|G ��  ��  �=G �5�F j�g  ÉM����F ��  #��  ��p  0�F �u��5��F ~��T�5��F �}��=��F ���  �   ��`  ��d  ���F �5��F ��X  ��`  �5��F ��T  ���F ���F �P�F �5��F �Z  �=��F ��G ��G     ��G ��G ������=�G ���G �2V  �=�G ���E     ���F    ���F �3����E���F ^��<�F �U�)�v�E�V�<�F �E��ɋ�G ��[�A��  ��  �XG ��  ��  ��  ��G ��  ������5|G �5�G ��@���   �'�}��|G ��   �������|G ǅ0      Q��0  ��   ���  ��   ��G Y�}���G �=�G ��|G �7V����0  �}�붋=��F �`�F �:�=��F ):�R�`�F �0  �5��F �|�F �%��F ������  �=��F ;=��F �*����=8�F ��F �=��F �d�F �l�F ��p  �8  ��$�  ��$�  ��$�  �ދ-��F ��$�  ��$�  ����L$(�-�G ���F ��G ��$�  ��$�  ;�$|  �u�����$�  �-��F ��$�  ��$�  �-(G ��G ���F ��$�  �  ���  ���F ��$�  �����G ���  ;�$P  ������$�  ���  ;�$�  �e�����$�  �$�  �� G ���  �dG Ћ8�$�  �=tG ǅ�      �~  ��$t  ����F     9=�F �A�����p  ��F ��F �F �l�F ȉ�l  � 8�F ��h  ���F     �=��F ��d  �=8�F ���  �P�F �5��F ��h  ����������`  ���F ���F ���-��F ��F ��A�F�=��F ���F ��\  ��h  �������   ��|G ��U����0  ��G ����R�pG �-(G ��$�  ��G ��$�  ;�$�  �������$�  �$�  �-dG �-@G ��M �$  ��$�  �-d�F ��$�  �0�F     ���F ��$�  �;  ��d�    �d�    �=��F ��
  5��F j �`�F     �E��}�R   ��������F �=��F V�5`�F �>�=��F )>�vY��  �4�F ���	  �-$�F �5<�F +5�F ��h
  �-I���H
  2�0���H
  ��$,  ��G ��$�  ��$�  ��$�  �0G �Ӌ�G ��G ��$�  ���  �=tG ����_�����$�  ��$�  ����$�  �$�  ��A�G��G � ��   ��G X��G �5�G ��v�@��  �5�G ��G ��  �����P�%�G ����0G �=�G ;�$x  �ǝ����$�  ��$�  �ы�$�  ��$�  ^��$�  �=(G �tG ��$�  ��G �-�G ��$�  �0G ��$�  �pG �-��F ��$�  �  ���  �<G +�G ���F ���  0�F ���  �5��F 5@G S���  �d�F �5HG ���  �-��F ��$�  ��$�  ��G �5pG ���F ��S��G �hG ���F ��$�  �h�F �=�G j�5�F �B���R��$�  �5pG ���F ��$�  ��$�  ��$�  �(G ��$�  ��G ��$�  �0G ��$�  � ���e�����G ��G ���-�G �G ��A���$�  S��G ��$�  �n�����$�  R�(G ��$�  ���F ��G �0�F �=��F �5�G ���G ��$�  ��$�  ��$�  ����������F ��H
  ZT� �F �΋D�F 0�F ���F ��$  ���F ���F ���F ���	  �����4  �|�F ˋ��F �%�F ���
  ���F 3(�F ���F ��C���  ���F ����
  ���F ��F �\�F ���F ���
  +�F ��  ���F ��F %\������	  ��  ʁ-�F ��#0�F ���F ��F ��  ���F ��$�  ���������   �ݏ�����"  ���!  Bǅ(      ��
G ���(  �X  ���k  ���F �8�F #� 	  0�F +� 	  3�
  j ���F     �E��}�   �z  �=T�F �5��F �5��F �>1�v���F �   R��F 3@�F ��ST0�F ���  35��F �$�F �P  +�8	  ���  Y+�p  �%��F ��  ��$4  �5��F �l  ���F ���  3��	  ��  ���F 0�F ���	  ���	  ӫ�	  �=H�F 3��  ���  ��  ��F 35P�F sT�5��F Xhދ�  ���F �X�F ӣ
  ���[z։��  ��
  3�P	  ���F �-D�F �����  ��p��@  W�\�F ��  ��QB ���F #�4	  ���	  STj �5��F WjP�5H�F ��  �Q���  ���  ��G ���  �5G �=G ���  ��G �5� G �=| G ���  �� G ���  ���  ���  �9]��M�����G ���  Y���  �6  �|G ���  ��G �;��F �4������  ��G �|G ���  �|G ����������  ���  ���  륋�   R���F �:)2�R���F Z��   �=T�F Q���F �9[��  �5��F 1�v�5��F ��F �ˋ�  �:����-8�F �8�F ��G �-G ��$�  ��G �ȋ�$X  �=� G ��$�  �pG �4G �8�F ��G ����   ��
G ��(  ��   ��@�A���
G ۋ�
G ��
G ��(  ������
G ��(  ��
G �A���j ���F     ��l�����l���   �������   P���F �8���F )1�I���F ���  �R���  ��  50�F 0�F ���F ���F ���  �%��F ��$L  ��G �=� G ��$�  �,G � G �;��F �\���P�=4G A��G �,G R�,G ���"����l$Z� G ��G �=� G �l$�,G ��$�  ��  +��  ��  ��h  +��  ���  ���  ӫ�  ���  ���  +5��F 35��F 50�F ��p	  #��F ���F ���  ���+��F +��F ��$�  �~������   ��G ���  G 9�G ��������  ���  ��G �8�F ��G ���  ������}����  �8�F �-8�F �L$��5�G �=DG ��$�  �-G S��$�  ��G ��$�  �T$���$L  ��G �-�G �|$� G �-�G �8�F �8�F �=G �-� G ��$�  �54G ��$�  ������G �<G �=� G ��G ���  � G ��G ��G �| G �5�G ��<  �-PG � G ��$�  ���ʓ�������8�F     j ��X�����X���   ��  ���F ��d���W�=8�F ����F � �F ����F ����3��L�F     h�  ��P����K  ��T����L�F ��=��F :�R�L�F �с��  ��ˁ��F ��>�0�F �-��F l��R��  ʋ��  ��  ���  ���  3��  3=��F �=4�F ���  3�   0�F ���F ��S���F ���  �<  =0�F ������������DG ���F ��X  _�$�  9��s����D  ���  �58�F ��<  �h�F ��P��<  ��G �h�F �5��F ��G �h�F �5��F �PG �h�F ��G � G �;��F �U�����<  ��G �=G Q�5 G � G �����HG ��G ��$�  �$�  9=HG �z���=�G �|$��G ��G ��$�  ��$�  ��$�  �=pG �HG �T$�DG �l$�=HG �G �=DG �8�F ��G ��$�  �= G �������F ��\�����P  �/P���F 1(�m��=��F �5@�F ��F���  ���%4�F �   �TG ���F ���  ���  �9��*������F ��x  �G �8�F ���  �4��d���W�=8�F ��t�F � �F ��=8�F �t�F _��������  �TG �	;��F ��~�����F ��x  J���L������X�F     ���F �  ���F �l��Y�=X�F ��8�F �H�F 1��=X�F �8�F ���ǋ��F ɋ�   3�  OT�E�D�F �F ���  j�2�+��  �����MЋ��  �%D�F ���  3�(  �M����  Ɂ�h  �|@�OT�U����  3�x  ��  ��h  +��F ���M����  �E��l�F �- �F ��$  =)$�0�F ���  �U�0�F ��F ӧ�  ��$  � _�4���F �E�14����F ���F ��<��2��D���XBT�o  �=XG ��G ��$�  �-�G �=�G �|G �=�G ��G ��$�  �|G �-�G �<G    j�G     �=�G ��G ��$�  Z�-<G ��|G �-�G �|  ��G �G ���G ��w���=�G �G �-<G �=�G W�=�G 뗋5`�F _�7�E��F 1�W�E��   ��H  �5�G ��G ��  �=8G �-8G �|G �=�G ����$�  �tG �-�G ��G �5�G �|G �-8G �����GT��8  ���  �0�F ���  %�cb�5��F �,!���  ӯ�  ���  ���F j ���F     ���F �=��F    �����5`�F _�7���F ��F 1��=��F 3��F ���F 0�F �]��   ���  S��\  ��0  ��QB �%D�F 	�%��F �5��F �����+�  _T���  3��F Q���F ӧ�  ���������F XGT���F ���F ��  �l�F �Np��R  j �E�    ��D�����D���   |[�=��F �u�>Q�M��v�`�F X+�F ��F ���F ���  #h�F �=��F ���F �l�F �`�F �b����=��F �u�>S�]��v�u�[�t����	��G �A��$   ��G ��$   �_����}�^�>1�vV�   �0G ��$�  ��G ��$4  ��$  �|G �5�G �D$���G ����G ��G �I��v���G ��$  ��$4  �=8G �-G ��G ��G �,G �,w��j ���F     ���F �=��F   �F������F �}�^�>1�v���F ���F 5�K���F �l�F �5l�F 50�F ���F �%x�F ���F     h'  ��������:���=��F �7���F ��  1��=��F ��X�-�G ��$  ��G �|$��5�G �\G �E �-�G �=,G �58G ��G �m��$�  �@��G �-�G �Ћ|G �5�G �l$��d�����$�  �XG ��$�  � G ��$�  ��$�  ��G ��   ���  ���  ���  ;�$�  �?����$�  �$�  �5�G �5XG ΋.�$<  ��G �5�G ��$�  �XG     ��$�  ��$�  ��$�  ��G ��G ��G �<���Ǆ$�      ��$�  ��$�  ;�$�  �*?����$�  �$�  ��$�  ��G ��$�  �)�$<  ��$�  � G     ��$�  ��$�  ��$�  ����z  ��$�  � G ��$�  ���- G  G ��A���$�  ��$�  �8G ��$�  ��$�  ��$�  �8G ��$�  ��  �-�G ���F ��E���   +��1  `G AT�U�}����3  ���   ��3  ��H  ���   ��D1  ���   ��H  ��H  ��G �B���   �B���   ��   �E��E�XG ���   �x�M��H���   �p���   �H�G �H�5��F ���2  �$G ���2  �U����3  ��G ��G � G ��2  ��G �]����1  �%�G �ǋ�G ��5�G ��É�G �% G �����$�  ��G � G ��$�  ��$�  ;M �=�������  ���  �"����j��D  �J���   �j���G ��G ��G �= G �u��4G �|G �xG �=hG �5HG �%LG �Ë����G �=HG Ë�$�  �-�G �- G �-�G �5\G �58G �5 G �5\G �-�G �t����-$G ���F ����F ��3  ӊ�1  �E���   ���  3��3  BT���2  ��,3  +�h,  ���}����1  =0�F �5G �u�����	��G �A��H  ��G ��H  ��   ���F �5L�F �}ȋ71��]��]�0�F �u�΁%��F �<(���F �q350�F ���F �-��F �5��F �M,ǋ(�F �%��F �  ��H  ��G ��R�@��G ��G �� ����5�G ��H  ��   �<G �G ��  �|G j ��(����G ��G V��G �5�	G X�5�G ���	G �����W��$����N��N����G �=PG V�� ������G ��G ��G Z�PG ��	G ��$�����G ��G ���n�����$�����G ��  �|G � G    j �� ����=xG ��  � G ��=�G �|G �������H  Y���$(  �@U���� ����=�G �5G Q��H  �5 G �=xG �5G 둋��F _����F 1���  �5��F �|�F Ӯ�  ��X  VT���F ���F +��F �z  0�F ���F �]�_Tȉ]����F #P�F �(�F �0�F 3��  �M��X�F ���F ��4  Ӈ�  -r��3X�F ����t0�F ���F 0�F ���F ���  #�p  0�F ��8  #=p�F �}��=��F ��B�>�=��F =�F �E����F �T�F ���  �+=H�F ��x  ȉ��F ���F ���  �  �E�    ���F     ���F �=��F    �O  �=��F �Uȋ2�]��d�F )�R��  ˉ�T  ���F 3��F _T���  +��  d�F �M����  ӏ�  ���F �%d�F ���F     �h�F     �h�F �=h�F /   �z  �5��F ���F ���  �S��8  1����F ��  Q��   ��QB ��x  ӅL������  ӌ$�  �T�F ���F ��F ��F �   �5`�F �f  ÍI��   ��9����H  R��G �|G     ǅ      �������G    ��G     ǅ      ��  �Ή�G ��G ��G ��G �5�G [��G �   ��$�����G ��  �|G W�����ǅ     ��G     ��H  �� ���X��  �TG ��G ��G ��  ������ G �TG �%������F �=��F ��5�F 17��=��F �J����5|G ��0�����G ��������V  �Uȋ2�=d�F ):�R�U�����0�F �u����#�D�F ���F +��  ��h  =0�F ��d  �E����  ӣ�  ���F �%��F �E����F ��  �=��F �}�=0�F �E��D�F CT��x  #�  ���E'U��  ���F �- �F �}��=��F 3=P�F ��  �U��U�ʉ��  ��D  +�  �  R�hG �M�GN���hG ��$�  �-�G Z�5hG ������   �2  ��   ~T��0  �-$�F ��H  1�$s��  �F 3��F 3��F ���F �T�F ���F VT��H  bJ�F���  ���  #��  ��  ��H  ~T3��F � �F 
���  ���F ȋ�D  �FTPd�5    d�%    �5��F �5��F ���I�@P��	G �=G �D$�=hG ��$�  �=G [�����S�hG ���G ��K�����  S�]�^�����   ���I�C��  ���G �rL��P��G ��G ��	G �5hG �-�G ��$   ��G ��$�  �-|G ��G ��$�  ��9���X�T$��hG ��	G ��$�  �\$����H�����G ���F �G    ǅ      ���  ���F ��  ��G �o����  �֍��F �R��   ��o��ǅ      ǅ      ǃ�$     �������8G ���F ��  ���G �E��� G �ދ8G �5 G ������E�    �E�    �E��}�   �  ���F �uȋ�]�)�v�D�F ��F ,�F �5��F ��h  �����  NT0�F ~T�]��d�F ˁ��  {�∉��F ���F 3��F �O  �(�F ���F ��F �$l  9��������x  ���F �8�F ���F ��p  ���F ��x  �;��F �������h  ���F BI����������F ��p  ��h  ���F ���F ��F ���F ��x  ��F 둍��F ��I�@���������  ���  �$�  9��y�����G ���  �8�F ��G �= G �=�G �/;-��F ������-dG G��H���u����5dG �=DG �= G ���  �DG ��G ���  ���   ��E�    �E�   �M���%  �uȋ�=��F �]����F ���F ���   ���  )>�v�uȋ��F �]��=��F 붋uȋ�]�)�v�u�������<  ���F ��� ���	��@�
G �@�����$  ��<  ��0  ��$  ��   ��8  ��<  ��   �F��0  ��	G ��(  ��8  ��$  ��<  ��	G ��   ��(  ��0  �
G    ǅ8     ǅ(      ��0  �t)�=��F ��(  ���$  �*�����0  ��(  �͍=��F ���"  ��G ���G �B뽉��  ���F �5L�F ���F �t�F � �F ��t  �����  ���F � �F ��p  ���- �F  �F ��A�B��l  ���  ��F ��h  ���F � �F �m���F     ���  ���F �5L�F �5��F ;5l�F �����5��F 5��F �d�F �T�F ���  �8�F ��t  � �F     �������F ��l  ��F � �F ��t  �t�F ���F �5 �F �5�F � �F � �F ���F ���  �����|�F Ӄ(  ���F ha.�E���\  3�  �}����  +��  ωE���F 3��F ���F ��F �u��5��F � �F ���F +��F ���u�+5��F �}��=��F GT3��F ���F [�6?���  ����U����  0�F 3�F ��p  ��$  GT�-d�F 37�C���������  d�5    d�%    �5�F �)  0�F ���  ���F WT���  ���F +t�F ���  ���  ӯ�  ��  ӏ  �t�F �X�F ���F #�,  38�F ���  � 󤉝�  ���  +D�F �8�F ���F 3p�F ��+��  _T0�F �]���d�5    d�%    ���  ��  �5��F ���p  �% �F ������F � �F ;$�F �������F ���F ���  �d�F �I���0�F ���   �%0�F �5�F ��T  +��   ω}ċ=��F ω}��}�{T�]�ˉ��F ���F �0�F  �F �u��5(�F 5D�F ��@  #�F ���F ���F ��F �]�XT�pT�-��F ���V�}���   �=0�F ɋ��  3��F �=��F �  ��$�  ��G ��$�  ��G ��G ��$�  �=lG �����  �4G ��$�  ���-4G 4G ��A�G�=G �LG �,G ��$�  ��$�  ��G ��G ��   �=|G �=��F ��8  ] 9��kT�����  ���  ���  ��\  ���  ��G �=|G �tG �54G ���  �;��F �jV����G F�tG ��G ��G ��G ����S����G �5�G ��G ��G �54G �G ��G ���  �G �q����5 �F �L̋LG �-`G ��$�  �-G �-lG �-`G ��G �4G ��G ��$�  �LG �4G ��$�  ��G �C�����$�  �%4G ����5HG �54G ��$�  ��G ;3��O���-�G ��$�  �쉅�  �-�G �5HG �Ë�$�  �Ǆ$�      ��$�  ��G ��$�  ;�$�  �:�����$�  �$�  ��G ��G �8G Ћ�F �lG �4G     �x����=��F ���F ���F #�x  �]����   _Tȉ��  ��  ӯ�  ���F �F ���   �_ЉM����F �-0�F �-��F ��qm�5��F �u�3��  �]���d  #4�F 50�F ���  ���F 0�F +��  �5��F ;�ǉ��F ��  �0�F ���F ��T  +@�F ���  ӏ<  �l�F ��F �5�F �5�F 50�F ��  =<�F ���F ���F ���F ���  �-@�F {T�@�F 3�F ���F -!�+�E����  ��  �M�0�F �p�F ���F �H�F ��F �\�F �H�F ��F �p�F 0�F �}����  ω��  �|�F ���CT��J�΋{T�M���0  ӫ\  �%��F +��   0�F ���  _{T�}ԋ=��F +=P�F �MЋ��F Ɂ��t46���  ��F #\�F 0�F ���  ˉD�F ���F ��F �5��F �5D�F 35��F ��  ��5�
�sT��T  ��T  C�{T�E̋,�F 8�F �l�F ���F ӣ�  +�F 0�F �}ȋ=t�F +��  �	�����8  �=�
G ��8  ��0  ��G ��[�@��G �Ћ�0  �+��<     ������$  ��
G     �t����F ��8  �=�
G ��
G ���$  �������
G ��8  ��B�<�F ���F ��t  ���F �(�F �5��F ���  �] �����  �<�F �T�F ���-<�F <�F ��A�B��F �=<�F �x�F ���  �5�F �5<�F ��  ���F ��F ��ZTP�E�BT�J|�Bd� �F ���F 3��F ���F ���F �@�F �5��F �5 �F 5h�F �Kd0�F sT���   �;�#���   ���P�x�F �P�`�F 0�F ��y�EeP���   +��   �u�?��0�F ���   ��7q��   �-t�F ��mP�\�F +l�F �4������F �5��F ��d  ��x  �=��F �T�F ��p  �5��F �=<�F �n����-��F ��$�  ��5��F �h�F     9h�F �G ���5��F ���  �h�F ���  ��  ��  ǋ/-8�F ��$  �쉖�  ǅ�      ��$  ���  ���  ���  ���  �|�F �=�F Y���F �$�F ���F +=��F �(�F S�=��F ��t  ���F ��x  � �F ���t(���  ��p  ����$�  �$�  ��A��]�����p  ��$�  ������F ���  ���  ;��F ��������F ���F �h�F ���  ��t  �(�F �=h�F �] ;=��F ������=h�F =h�F ���F ���F ��l  ��8�F �=|�F ���  �T�F ���F     ��h  ���  ��d  �5��F ���F ��t  �5��F ��������F �8G    ǅ     ��G     ���   ���F ��G ���$�  ��  ��G ��W�=D�F =0�F ��F �B0�F S��F ����Jp�ƋJt�-<�F �5<�F /�y0�,�F �j(�Z�Z`3�z�z(=$�F ��F ���F ���F �R���F ���F ���F 0�F 0�F ϋJx�H�F V�rl+rD=0�F 50�F �e��5��F �|������F ��I�B������Y��G ��G Ǆ$0      ��	G �pG �tG ��	G �5�G ��G �|G R��$  ���   P�-tG ��$8  ����   ���(�F �-��F 'I�����F �5(�F �v^�qLqT�A�y<ρ�3r�Y�yT�ú���AATYT���F �IX�J�J\�J�jh�'9>�jh�TNV�r4������F ��� ���	ӉG�8G ��0����  ��  �|G ������-tG ��$  ��$4  �-�	G P��G � ��G �@P�-�	G �T$�5�G ɋD$�|G ��<����G ^�|G ��$8  ��$  ��	G X�݋5�G ���������F ��F �%<�F ������F �5<�F ;5��F �����5��F �h�F ���  ��l  �=��F �5��F ��F �<�F ��p  ���  ��l  �5��F ���F �-����|G ��v�A������  ��t  �=��F =��F 9��Q���|�F �5\�F �58�F ��p  �5$�F �5\�F ���  ���F �|�F �;��F ������p  A���  �$�F �$�F ���A����p  ��l  �����F ��l  ���  �5|�F �5$�F 넉l$؋�G �tG �E��9���������XG �E��8�F �G �	  ��G ��  �t�5\G �5�G �\G ���  �5�G ��v�@P�5�G ��H  ��T����G �=xG ��  �dG    j �5�G W�������  ������H  ��  �dG �c����|G ������K������@G ��H  �������  _�@G �dG 듋��  ��  ��FՁ��F ���2��   +��F ��   +5��F �]ċ��  0�F ���  �=��F ω]��]�ZT��d  �]��U��=X�F �}��V  �%,�F ������F �,�F ;��F ������p�F ��d  ��`  ��h  �5��F ��  ��$�  ��$�  ��$�  ��$�  �HG � ;��F �7���XG �HG ��$�  ��$�  ��$�  ��$�  ���z}���XG ��$�  ��$�  뉉0G �8G �XG �;��F �����A�0G ��G �0G ���5�����G ��G �M��8G ��G ��G �XG ��G 땉�$t  ���F ��$x  �-P�F �-�F �U�$�  ���p�F     9=p�F �\�����x  �5��F ��p  �p�F �p�F p�F �(�F ��x  ��l  Ë3�$�  �`�F ���F ��h  �,�F     �  �5��F ��\  ���F �=��F ��P  ��  U��U���   ���   HT���  �=��F ���@  ω��F �\�F 0�F ��`  ���  Ӡ�  S�h�F +��F �K  �E����   �E܋MԉJ�5��F �u��}��r�<�F �B�5@�F �r���F �B���F ǃ,      �M�E�}���  �@�F ���F ���  ���  Z�M��u��E�}�m䉓�  ��,  ���  ��X  �=P�F ��   �L$܋T$؋D$��  �%��F �����d  ���F ;��F �����p�F �p�F ;�$l  �¦���p�F p�F ��\  ��x  ���F Ӌ�$�  ��X  ���F ǅT      ��\  ���F ��P  ��T  ���F ��X  �5��F ���F ���F ��`  �����HG �LG ��$�  �G 9HG ��~�����HG ��$�  �HG �58�F ��$�  �-����=��F �5��F �=��F �u���3u�)5x�F �U��x�F +U��F ��)U����  3=�F )}���F �E���3E�)E��X�F �  ��l  ��h  ����j�����`  �,�F ��d  ���-,�F ,�F ��A�G���F ��h  �7���9����5��F �5��F ��d  ���-��F 5��F �-��F A5��F G��\  ��X  ��T  ���F ���F �,�F �ދ�X  ��P  ��\  �=��F ��h  ��P  �p������F ��3]�)]��E�+��F �E��E�+EȉE����F �]����F � �F �x�F �E����F �  +h�F ���F �8�F ��@  +��F ��F ӈH  ���  #�F ��F V�u���   ��(  +��  ���F ���  �����F S���F 0�F �^  �E�+��F �U�+UȉU���F �U��
�
�E��]�E�E����E��}�Z ��3���U�|�F �]��=��F ���F �u����F �m����F ���   [���F ���   ���F �L$ĉ��  �T$������  �|$Ћl$ȋt$ĉ��  ��  ��  ��0  �-��F �5��F �D$��|$��l$���`  �=��F ��   �%x�F ��F ��d  �-��F �5��F �=p�F ��Ë��   �5�G �P��D  ���   ��D  ��G �H��G ��G ��G �=�G �E��(G �PG ��G �=�G �$G ��|����G �%XG �ً-�G ���=$G ��M����F ��)x�F ���  3��F )x�F �E����3����5��F �u���3u�)5x�F �x�F +E� �F ��)E����F �t�F 3 �F )M�� �F ���  ��L  ��<  �PG ��G ��@  X�PG ��R�@��G �ʋ�,�����G ��  �|�F     j ���F     ���F ���F �@���F �=��F �U����F �Uԉ=��F SVX�m苸�   ���   ���  ���  �T$ȉ\$čU    �5��F �-��F �.���  3|�F �x�F �   ���D$�   �D$�   ���F �T$����F �
3D$����F �E�    �l����-�G ���F ��E���   ��P  �}����   ���   ��P  ��G ��H  ��H  �P���   �x���   �P��|������   �\G ��D  �n����H G �� G ��d  �5x G 5( G 95H G ��T���=�G ��X  �=H G �8�F �= G ��`  ��   �=�G ��8  ��@  �,  ��  �|G �J�>����8G ��G ����  P��L  ��8  ���G ҉�@  ��  ��8  ��4  ��G ��G ��4  ��8  ��G ��  ��  S��G ��[�AS�����Y��G ��G �U�����$  ��j�\G     S�5\G �\$�5�G �\$[�������   �=�G �=�G ���F �H G �;��F ��]���H G ���F ��l  ���F ���P^����=�G ��l  ���F 룉�   ��G �|G �=tG �=�G ���A�=�G ��=tG �|G �%��j��G     �5�G Y�|G ��   �t���   �|G ��G ��G �I����5�G Q��G ��G 볁��   ���   ��  ��B���8G    ��G     ��  �8G ��G ��|G �T�����  �|G �J������8G ��G 뽋�8  ��L  ��<  ��I�@��G �	G X��G ��G �lG �	G ��8  �lG �m  ��$  ���hG    j �hG �=�G �T$_�=�G �=�G �����������  W�=�G ���A�=�G ��_�$G ������=G �G �=�G ��@  ��<  ��G    ��,����=�G �=�G ��L  ��������,�����L  ��8  ���G ҉�@  �f  ��,�����L  ��@  r>��<  ��8  =   ��  =�7  ��  =  ��  =   ��  G�   �=�G ��8  ��@  �O����-hG ��U���   ��G ����   ���   0�F �}��=�G =G ����U/��0�F ���1  �M�u��u��2  ��G �5�G ���   �]����1  ��G �Q�}����   ���   �q��2  �y���   �q�u��q���3  �U��=hG �u��]���x2  ��@1  �=PG ���3  ��G �E��G �%�G ���ڋ�=�G É�L  ��<  ��8  ��I�@��4  ��G X��4  P��L  ��@  �������<  ��8  =   ��   =�7  ��  =  �m  =   �=  G�   ���   ���  ��G (G 9��_����5�G ���  �8�F ��G ���  �hG ��G �;��F �������G ��G �hG I���������  ��G ���  ���  몉�L  G��  S��   ���  ��QB �E���l  ���F �H�F ��F ���F �E���(  �U��E���QB �M�OT�U�0�F ��,  ��F +@�F ��  �$�F ��0�F ���  +��F +��F ���F 0�F 0�F �E��E�+��  GT�]���  3�F ��x  � �=��F ��G    Ǉ8      �=�G ���   ��L  �=��F �=G ���G �f  ��G �=G ��L  ��G ��G ������]��uЋ�M��0�F �v�uЋM���   �=�G ����4  �5�G �5�G ��4  �  ���F �uȋ�]����F �-��F ���   ���  )�v����F �i��L  �5��F �1�I�F�d	G ��L  ��G ��L  �d	G �5�G ������L  G��<  ����8  ��<  �5�G ��8  ��  �E�    �E�    �E��}�   ������]��uЋ���F �0�F �v�U����F ���F +,�F ���  �U�0�F �=��F �=��F �|�F 3 �F �]���  ���F j
�S����\�F 8�F Q���F �l�F �t�F �(  �<  _Tj �E�   �M��h���_�4�E��E�14�W�E��ቕ@  ��L  ��  ��<  ��D  � ��L  ��4  ��b����<  ��D  ��8  ��$   ���	�$  �,G ��4  �
B�,G ��L  ��  �u���S��D  ��@  ���<  �I��G ۋ�L  C��D  ��8  ��D  [��8  �O  ��8  ��L  �4G ��8  �=4G ���@�=4G �؋�D  ��G ��   ��D  ���F H�f  ��[����G ��@  ��$  ��D  ��L  )ڋ�G �=�G ��8  �pG ��@  �ǉ�4  ��<  �ʋ�8  ��L  �5DG �׋�<  ��0  ��G ���;  ��4  ���DG ��4  ��G �DG �a����=�G ����4  ��G ��G ��4  �6����	G ��D  ��L  ��  �4G ����@  �ڋ	G ��G ��@  �������<  ��D  � % ����$  ��D  �G��I�B�  �=�G ����G ��G ��8  �����  ��D  ���F ����L�����G ��@  �=�G �,G ��G ��L  ��,�����<  ���  ��   ��<  �K�����4  �  ��L  ���F ��D  ǅ@     [��G ��r������F S��D  ��<  �	G ��G �4G ��L  ��@  ��D  ɋ�<  ��p���������D  ��L  ��4  ��8  ��^����<  �׋�L  �x�4G [��<  ��D  ��L  ��@  ��L  �	G ��<  ��@  ��G ��,����4G �0����=��F �9�I�G���`��D  ��<  ��T  ��L  ��   �˫�����  �  ���  �ܛ��ǅL     ��G     �t��=��F ��G ��G ���$   �i�����D  ��G ��D  �=�G ���=$G ��   ��D  �=�G ��@  �=�G �$G �=�G ��L  ����@  �  �tG ��L  ��G ��@  ��L  �tG ��<  ��G ��D  �tG ��P  ��@  ��������F ǅ4���    R���  ��,�����   ���L�F ��0������� G ���F ���  ��\  ��A����G �M��G ���5t�F h@  j �   �D	G ;��F �*  ��G ���F ��\  �=xG W�� 
 ��\  �=<G �  W�j���F ��X  ǅT     ǅP      ��G     ��H  ��G �xG �(�F �G ��L  �����A��� ��G ���F ��I�C�Ë�G ������L  �$$  ���F ���   �XG ��L  ��G ��D  �=�G �% ����$  �B��<  ��G ��@  �	G �XG ��G ��L  ��<  �:�����D  ��@  ǅ<      ��G ��<  ��P  ��L  �����=��F �9�I�G�������=��F �9�I�G��������=��F ��G    ��h  �=�G ���  �g  �������O��D  ��T  ��L  ���   ��5�G �5��F ǅ@      ��G ��L  ��@  ���D  ��<  ��   ��@  ��D  ��L  �=�G ��@  �=�G �5�G ��@  �O�&�����D  ��@  ��<  �5\G �=�G ��D  �֋�<  �p�����P  �=PG �H	G �LG �PG �8G ��0����D	G ���x�����L  �=��F ��G ��I�@��L  �������@  ��D  ��L  �5�G ��I�@��<  �����=��F �9�I�G�������=�G �p�����G ���F ǅ$���    ����t  ��\  �Ѝ��F ��G ��h   ��\  ��G ��T  �=<G �H	G �5xG �xG ��X  ��G �� 
 =�G �LG ��T  �5��F �����ÉX�F ��$�  �=0�F =��F 9=X�F �B�����$�  �쉍p  �(�F �X�F �8�F ��t  �0�F �   ��0  �=��F �$G ��0  ��!  ��0  ��(  ��G ��I�@��$  ��	G ��!  ��(  �$G ��$  ��	G ��G ��0  �$G �5�=��F ��<  ��G �	��G �A��(  ��<  ��(  �   �c����F �X�F �;��F �?����X�F ��F �@�F ��F ��������=@�F ��뷋�8  ��������0  ���F �������G    ǅ8      ��0  ��>����=��F ��8  ���G ������0  ��8  �ʉE�pG �M�M�9M��6������}܋8�F �}��G �}���  ��T����=L�F ����F �0�F ���F ��F � �F ӠP  �d�F ӈ(  ��P  �F �^  ��(�����G ��G    R��  �TG ���$�����G �������  �|G �����������TG �=|G Zǅ����|g �58G �������}   �=�G �?��G �G���   �5�G ��p  ��H  � G ���F �	;��F ��U�����F ��$�  ��X  ��p  ����V����P  ��� G ��X  ��V�������3  �r������7��O�=8G �=�
G �=�G ���   ���%8G ��
G     ��0����=�
G �I�"����=�
G ��j ���F    ���F �w������F _����F 1�W�ۉE��pG ��G �5PG �u��;��F �6���� G �5PG �E�pG �M��E��������� G 뮉��F ��p  ��\  ��X  �9��F �NV����P  ��p  ��L  ��H  ���F �=8�F ��G �=�G �T������  ��t  �t�F ��h  ���  �=��F �=��F �;��F �A������F G���  ��$t  ��l  ��t  ����������F �=��F ��l  �t�F ��t  ��p  �=��F ���F ���  ���F ���F ��   ��t  ���  ���F �F 9�$t  �������p  ���  ��t  ��h  ���F �58�F ��l  �����=`G ��G ��G ���G �CS��G ^�����4G �T$��dG ��$�  �0G �;��F �������$�  �0G �4G �54G ���6������4G �dG 룋��F �q���Q���F �T�F ��p
  �W��D  1:�R�,�F ���F ���F ���F ��F ��0  3��
  �$�F ��F ��  ��F Z�
�=l�F 1:�RR��  ��
G �4G ��@�A��(  �p	G ��0  ��	G ��(  �?  -���<0�F ��82  �H̉�0  ��82  FT�8G ��\2  �-<G ��`2  �L����43  +0G �HG �LG ӆ`2  ���2  ��l1  3G ��d1  �<G ^T��$3  Ӧ�1  Sd�5    d�%    ��G ���2  �LG �j �x�F �   �x�F �z?���=��F ��  Z�:��D  :�RR�Ս[��   ��d����
G �4G     ��(  �4G ��
G    �DG ��	G ��
G ��0  ��p	G �������	G �p	G ��0  ��(  �4G ���
G �a���
G ��
G ��(  ��   �=
G �=4G ��   ��d�F     j �d�F �=d�F @   ��������F ��F _����  1����
  3��
  ���F ��F BT��D  ��D���3��
  0�F ���
  ��0
  �5��F rT�����0G ��G �5�G �$�  950G ���������$�  �8�F �0G ��$�  ��$�  �u�����d�    �d�    ��G ���2  �-�G ��G +��2  ���2  �t2  �G �HG Ӧ�2  �-dG W���2  fq|����3  ���2  2�y����2  0�F jd�	����                                                                                                                  �e �e f f (f Df Xf hf xf �f �f �f     �f �f �f g g +g 7g Ig Wg mg {g �g �g     �g �g �g �g �g h +h 9h Kh ch qh h �h �h �h �h �h �h �h i i !i     @i Pi fi ~i �i �i �i �i     �i j  j 6j Dj Tj nj �j �j �j �j �j �j �j �j k  k <k Tk dk rk �k �k �k �k �k �k �k l  l 6l Pl ^l nl �l �l �l �l �l �l �l �l m $m >m Jm \m rm ~m �m �m �m �m �m �m �m n n (n <n Ln Xn fn zn �n �n �n �n �n �n �n o o 6o Bo     ��������    \�@     ����    �N@     ����    0�@     ����    #�@     ����    ��@     ����    Q�@     ����    4�@     ������@ ��@ ... A buffer overrun has been detected which has corrupted the program's
internal state.  The program cannot safely continue execution and must
now be terminated.
 Buffer overrun detected!        A security error of unknown cause has been detected which has
corrupted the program's internal state.  The program cannot safely
continue execution and must now be terminated.
        �����A �A Unknown security failure detected!  <program name unknown>  Microsoft Visual C++ Runtime Library    Program:    

          �����@ !�@ ������@ ��@ �����TB �TB     ����N�@ R�@ ����K�@ O�@ �����@ �@     �����@ �@ GetProcessWindowStation GetUserObjectInformationA   GetLastActivePopup  GetActiveWindow MessageBoxA user32.dll                                                                                                                                                                                                                                                                                        ( ( ( ( (                                     H                � � � � � � � � � �        � � � � � �                           � � � � � �                                                                                                                                                                                                                                                                                                               h ( ( ( (                                     H                � � � � � � � � � �        ������      ������                                                                      H                                      ����    �ZB InitializeCriticalSectionAndSpinCount   kernel32.dll        ����R�A `�A     ����    5�@                     h ( ( ( (                                     H                � � � � � � � � � �        ������      ������        	
 !"#$%&'()*+,-./0123456789:;<=>?@ABCDEFGHIJKLMNOPQRSTUVWXYZ[\]^_`abcdefghijklmnopqrstuvwxyz{|}~ ����    ��@     ����    �\B     �����@ �@     �����\B �\B     �����KA �KA     �����KA �KA     ����    ��A mscoree.dll CorExitProcess  runtime error   
  TLOSS error
   SING error
    DOMAIN error
      R6029
- This application cannot run using the active version of the Microsoft .NET Runtime
Please contact the application's support team for more information.
   R6028
- unable to initialize heap
    R6027
- not enough space for lowio initialization
    R6026
- not enough space for stdio initialization
    R6024
- not enough space for _onexit/atexit table
    ... <program name unknown>  R6025
- pure virtual function call
   R6019
- unable to open console device
    R6018
- unexpected heap error
    R6017
- unexpected multithread lock error
    R6016
- not enough space for thread data
     
This application has requested the Runtime to terminate it in an unusual way.
Please contact the application's support team for more information.
   R6009
- not enough space for environment
 R6008
- not enough space for arguments
   R6002
- floating point not loaded
    Microsoft Visual C++ Runtime Library    

  Runtime Error!

Program:    ����    o�A     ����    &bA ����    4bA kernel32.dll    FlsGetValue FlsAlloc    FlsSetValue FlsFree     ����V"A j"A Sunday  Sat Monday  Tuesday Wednesday   Thursday    Saturday    Jan Feb Mar Apr May Jun Jul Aug Sep Oct Nov Dec January February    March   April   June    July    August  September   October November    December    AM  PM  MM/dd/yy    dddd, MMMM dd, yyyy Friday  HH:mm:ss    Mon     ����_�@ c�@ am/pm   a/p Sun Tue Wed Thu Fri SunMonTueWedThuFriSat   JanFebMarAprMayJunJulAugSepOctNovDec    TZ  ����      @     ����    �A     ����    $�A     ����      @                 �c         �f  P �c         �g 4P (d         5i lP �d         �i �P �d         Po �P                     �e �e f f (f Df Xf hf xf �f �f �f     �f �f �f g g +g 7g Ig Wg mg {g �g �g     �g �g �g �g �g h +h 9h Kh ch qh h �h �h �h �h �h �h �h i i !i     @i Pi fi ~i �i �i �i �i     �i j  j 6j Dj Tj nj �j �j �j �j �j �j �j �j k  k <k Tk dk rk �k �k �k �k �k �k �k l  l 6l Pl ^l nl �l �l �l �l �l �l �l �l m $m >m Jm \m rm ~m �m �m �m �m �m �m �m n n (n <n Ln Xn fn zn �n �n �n �n �n �n �n o o 6o Bo     � CryptEnumProvidersW �RegConnectRegistryA � CryptReleaseContext � CryptGenKey � CryptGetDefaultProviderW  � CryptSetHashParam RevertToSelf  �RegEnumValueA �RegEnumKeyExA � DuplicateToken  �RegRestoreKeyA   AbortSystemShutdownA  ADVAPI32.dll  AddFontResourceW  �PolyBezier  BSetWindowExtEx  �GetTextExtentPointA �GetTextFaceA  �PolyDraw  SetArcDirection .SetMetaRgn  zGetFontLanguageInfo LGetBkColor  /SetMiterLimit �GetViewportExtEx  " CombineTransform  GDI32.dll TGetScrollBarInfo  KGetPropW  �SetWindowWord y DdeInitializeA  � DefFrameProcA RegisterClipboardFormatW  � EnumPropsA  �ShowWindowAsync /GetMenuContextHelpId  � DrawCaption � DestroyIcon FSetCaretPos � GetClientRect �MonitorFromWindow � EnumDesktopsW PtInRect  U CreateDialogParamA  � EditWndProc �ShowOwnedPopups uGetWindowRgn  �ModifyMenuW  AdjustWindowRect  USER32.dll � InternetOpenW i InternetCloseHandle � SetUrlCacheEntryInfoA � SetUrlCacheConfigInfoA  ` InternetAttemptConnect  4 FtpPutFileA d InternetCanonicalizeUrlA  a InternetAutodial  WININET.dll =GetCurrentThread  �GetVersionExW � EnumSystemLocalesA  ^GetFileType 7IsValidLocale � FreeEnvironmentStringsW OGetEnvironmentStringsW  �RtlUnwind � GetACP  �GetSystemInfo � FreeEnvironmentStringsA �GetTimeFormatA  7 CompareStringW  4 CompareStringA  5IsValidCodePage �GetTickCount  `UnhandledExceptionFilter  z DeleteCriticalSection �GetVersionExA vVirtualFree >GetCurrentThreadId  VTlsGetValue [GetCPInfo �QueryPerformanceCounter uGetModuleFileNameA  yVirtualProtect  �GetStartupInfoW GLeaveCriticalSection  mGetLocaleInfoW  kMultiByteToWideChar �GetTimeZoneInformation  HeapReAlloc D IsBadWritePtr OTerminateProcess  	GetCommandLineW �WideCharToMultiByte {VirtualQuery  GetOEMCP  �GetUserDefaultLCID  GetCommandLineA iGetLastError  HLoadLibraryA  ;GetCurrentProcessId SetEnvironmentVariableA �WriteFile SetHandleCount  InterlockedExchange �lstrcmpiA SetLastError  
HeapDestroy InitializeCriticalSection sVirtualAlloc  UTlsFree �GetStringTypeW  vGetModuleFileNameW  HeapFree  �LCMapStringW  �GetProcAddress  wGetModuleHandleA  �LCMapStringA  HeapSize  WTlsSetValue :GetCurrentProcess HeapCreate  � EnterCriticalSection  �GetStartupInfoA ?GetDateFormatA  lGetLocaleInfoA  MGetEnvironmentStrings �GetStdHandle  �GetStringTypeA  HeapAlloc �GetSystemTimeAsFileTime TTlsAlloc  � ExitProcess KERNEL32.dll                                                                                                                                                                    �H�ʭC������z����        c=�	�pn6�7u-3�c�EԢ                                                                                                                                                                                                                                                                        
+�y	$e4��6k���	�#7�]>�s�.%�o��C뮕Q|6���ԛ��x�_���;��IU��aM�\��,!ȴ�&7���;����^��C��Sv����u���1]C%�s��)�|�j�^ǵd�%�]j�Xz�]3��D�����H��{�qH5�~���@o�OG4�^    s���D`�S���cw)h�1��dM�Q�^��XԔy_k^	*h�'��z� �sNF�>�@ݜ�G��8^ы�H��6N�"�P�9���G�g�1Ԏ��2�sc�h����'dܕ�-�v��wP                                                                                                                                                                                                                                                                 ��(���	u@��޳b�4�pΌjT��]�Z6髥�mHwQ�����(�8��ax�Q�}as������4�+ì��TD���$���G����Y�=���]��'�N�WW��H�d���.�ӂǜk�^P)�[
�eV�g8=�f��R��!�H�I��r��b��QWZk�B�!>��հ��1(�eo���B˫�$p�X7g!�p�zMA��dn����t	�{��|?�UK6	���G��vt>IsoN)R\E�[Tw@,�����\9M}XE���׸}���{�?�!}�c�Mi$�ԝ�����E4�u�y� �]��5�Z��ԇ7��P�Q߼2U�[v3&<:@�T$�8p��߶g��_0���y2)��=������nw{g���
����j�<����r�������ך���%�)v��J��}+���坴͖�)c��:����^�����R�O�	��&��Y�k�(u6X���a��~��+��4�Rڴ�>,��|�GC%؍�$�Jf��e�Q��uw�`�E �ǡ���^���(�0�݂��p��Rf�O�C!rŅe�0aST9��f���7�N ��H�[��������G�-�����su�&��,��>�w��h�MB�)la~Y���N����d�ٸ�/j��YW\c-lǻ��Z�r�GQ��Ad?A_��6�}��SA����@}����̻&U��׶`����$�_rE�K�������$��&�[��L�_;)�Nm���:i��ä[���ΐF�9������ :d��C�[|��>�E�E�`�>k�-��M����S�f|�CiU!�ϝ}
쁿�V}������+�X���6w�_sP�a�%�橢Ǖ*lի��j/҉�OI9�����;%�kXZ�e^Q#:�FC8����>0�jCG�!:�fO�҉	�Xa~��E	}�Rl���듵ƄC�A�p�+wڮ�� Q�0��J���wr����t�"@ �|k<E`�,z�T��;�d���n�ޔ�`'(ސ��W��H�4C��p��)�&(�f#�L:u��"��**?W
��@����R����0�ܔ�)�lm�{F"���3/V5�}E��N�$��B���e�6,47o���2�Neg"��$a��vW�$��i��v�f&s�@�FK43 ���<���գ����\��gY�Y����,�v���1u�^�?�~�3���<� �Xx��⫭�T�/r �]�9�0G,�7�bk�qOʿ�5p�3�(�Ih��,���<�����ĳ��.6��r���:�M�^�$�	��sZ��� ���)J&��yiH��f�MLu�A^k*�*�U�p6F������� ˛aW0zt�X�ɸ���	�ӊ_�׺R�7Ȫo�v~����1�U�n�-9�iT�u��`[�aOhP��gP����'��Uw��=3.�xx�g��!���w>q�BT�#fY��U���(z�k:S~�ɲ���F�{�@�.f@�3�Ƈ);�>d�H��`99V�|�11��M��X�;�Δ��qO&�9�D���u�v��d�:m��{��8L���i��(?��FA���#�&��/ ��#�c-�d���l!���:���)��#J�m9��2#o�W�4a�}Wʖ�K����.z��M�F@Px��ď���	п�4�b�C�w��W�&��5��j�Yؙ�=0�U���q�,�u-�1�<&Q��	r���i1ysV��fw�Фz�c[*���3p�W� �_��.����k�n�$��=v9�*��F�hc�)p��OC���iV��m�}� F�8_.a,�="�J�,b�bS�\�,AYQz}�ێ��=��;Ʉ����R���ҭ��P����ս�U�����\p�4uk_Z�6AJ���;��.yޔ���ex �b�Vi��s�j�mQ�����iʷ�X�2�R�J7��KY��Q�I��&�LG���e��2�.H��Z���:�%�D��^���5MP�/a�}�=�/���o���H��w�+.�P���c����z{y̟���E�-�#��[�I 2�o��S�u� 8�9�(ؑ���Ռ������ރ/�P��I�4�����2T�y�iٔ
e�I2<�����P�;��٢��L�2$�� �V[icGL��b����2��z����M�,�kF�~��v���xZ��@FʎWk��!Z��#��o�PU�7��S�x�(L�T��T���N��{4����d��vR%3���&�$����:�D2C�=$���s�6qy�WQ|��`L�@'�y�cb�u|���dz�o�J�|�浊�- �@�Gڸ�}��>l4'}Ū���1?�,������'�֜Ȣ��ڨ6�8��ם��2P�Y(_`:�äe��.�z��	���V�	6bAY,MG� �[Ф{�E�xY���	�����zNFL8�L�ؤ݆�����;�a�:���5_?B}�� ���!ǌ�5�pg)�3͹A����[2F����������/�ǪKP9�;0�.l��x�Mo��='�m���u�����	Dd>T�<����+�m_��!;o{�!�a���8���U�e�D�I�)P`m"�5����0����<b�SRBv�8�[՛F[l!�bI)�����S2�e�ϗ�0H��&ؾ��v�Vx��)�V���Z9��K�Թ�l���7�ⅰ��*ai,�:�1��m����AW��`%���iQŹv�O����5:�ݒ�H��`�v�v	Χ1R-�F�]��b��*DN�����v��x"�Dے��}㔳�J�G�gz��. m��m,���]W����{���ZH�q�L*��Q	l�f����5���m�t�YE��᳓AJ�0��|og��7�l%������x輓�&+�Kib�l�i��6k�.v��APhh9�P������p%}x�Ӯ�"���k���9�Xk#��ڰT�S��Hk� �ǌ�6r��/�e^��}K&(T��l����M�������ե���m��H:!�0�\�oq{x���z1O�kz�9���V���9Io��w��\��;a�Uʁ?�Ը�#1��7/O�!2o��)�ym>옇uF(	��i�e��l�4���2ę��=�,�?=d!�	�@�T�Ux��7� ��I�^����r�(�����)���?��ukY��]W=0�V��
x��X�d��u�N�y��Y�I�'#KO,��a����bBQ�7w�`.p��Q��=$�J��c�H�6�C�ZL�'*Վ��\e)�z��I��Tc��W�L:i�LK��|ȱj��:e��'R(��0fGp?B-�s_B�s}.�od�
IG�P)V����8j&�n��=�����NbҲ��n5�ᢕϙ�Ȉ+C���:M� �;�G ��6*{/��I;��05؎�]�l���ze
5��6b�����HԚ[j����m���X�U�ό�������ٿ�,��ܬ}
շ�_J �W%3�cA!P ��!	�s��-�o.{-����~.i +�dq���Cș&R�d�g�e�Ǻ��@�X�Y�9�Pxp��_ݟ
+w�V`������{����\l����'�]����E�l_�Ӫ{���H}�j7���a���yQ$B���$��d� Ws���C��V�2���2�$������Nu���Z����1��'=_��v�/�_�u9�u��x�h�`�^U1d�]����f�X��L&Mt'�L�6���D���[)��R܈"m)ѫ�O6_�!�HT�  '��y�v�nΚH�!r�9�ǹ�b��c    `��^t�mؿ��9R�˃� AG3�-O��f����%M��p$n�u�M�G�I[�����V��Su�w#�饥ֺ���0���2N��Q��u!\QJ���`	x}e�J;J���j�0V����4`:ק����5    '�	uK�k󳤿�8��D������/���VQ����d����ʺ��&����WsxO�g�~07�s�2ԚZ���ܓgt��˔�Z�+o�	* ���R.�߸[F�0��K�;�Q\$����r	��P�o�����
������$7��KKhlM�xI��=���Q�#�����wYl���l�J
 �������7ӻ��#-�
JI���7�K!-���U�;��t���q*w�/j���3�;bP[�� ��"�@e�!�nM�
E�|_sܧa���%����M#�Y#ڎ72edS^F7A]���9	�B�,.5_�U/�3 ����^Ԏ�lsJ�>�h�'r+�RA�� ������v��l��"�%��.�-1����LР&XC�B������Q
?�Q,#~�B�����"������k�w��-!�2��w�{�;*�Dyē���՝�ݐba&�2�b@�/�zI����j�_��`9�����%��|�y�9�4�Tp�+☁(3&��C�7�20)��gЕAgL�#��� ߾4CՏ�Ŭ�0��,C��h��!Z5���Hk\ʎ�	2e��7��Fv�Np,Ef���@�F�M[3�9�W�M^pO�a�]p��
>��f�*��I��
g@p�XN�K+,�1:�z�C�^�r�����.�>1��^m�W�v�M���$�AMA�*T��Ep�����&�@����ӇA���ڍ�t�i �������W���>���C<���G��Ӈ�?7����ߥ�#�V�V��g?�e�:�OI���) �lsjO)�q��g'0�������?�~|�����MRps������,zƥj�֭��|��#t��%OY�V�(.��T>A 1��ׁ�^� mS�o�&�Iix�E(�E+5���U��b�r��2$��opj�R����)-���V��G��xlFOX3I����?�w~T�7�c���aJJ��Y	?2�I��s�@��ف�]�{aL���=�߁�S]\D�'�vOK&��Ԗ]�� +2�.?�LmL�� ���薫�P��7�	߉�V_����w������wD�����CS����a����a�<�����Զ��|��u�/c~y]$��?�)�#sDy�G� 5�CAr'����)!�����>��SM�.�� �W���v ������H�r�}�6�؏.V����վw`�4:�[�E�����ʍ/�i�_��vsµ���
����wɟ���]�CTY�H��p.RjXH�'�9��y'L;q���ִ"�&�#Ώ�3pzN�q+%SТ��҆.#I�-����i�o����<	�F�~�!ͤ���~�=��c�^�6ˆ�5�@e�q2*�� �\�~bm�?F/3�G		ld�4�����)�<����K�4Y�s�&�1�n�Ae����n�;���z:�'��Ӟ���$h?�4 W�Ac���0��Tm^G ����0u�)˔~5m��٪�@0���'�?���(f�D���v��~jN^�ժ��ұI�_��\3��jJ�7p��G�p/���ѴG�iqb#+�
aT�P� 9	������d�"4G��q���vgP-&!��Q�/�׏MLy�W����Gu�HN�V{��@~B1���FbU]Lfg�lu-7��6Fv.��O��dĽ/x�E��.L8�r�F%�.��͊��3���X��D�2[.�-��a&ѲXJ�^��_��]ѭ��]��L�$�O��~��	so�^R��͓3RDѧ@&Ҕf��t�4�4�DÕ��^��!�
��r5�i��<��f�TCa��QKH,|/��%�Z|�X��ٯn��E�d�#�O��E�L+�����}=����>��qÎ�h��&^���,�MO�8[�~%���'ڊc_��`�:�����\1ӊ��!Ė��0Tf�)
���ꈣ�k��R4ak5��#�˘6�j�,)V�+>��K�-���[�H.,���3� #�$�A����A��)W>�a�U��L��n��H��<���D��f�q��6��t�{��Пc��4�8�|~A�+�ێ2�bit�*�6š�>.����P��I��d��h��2�9g�H��<�?�Y��P�^_w������3�MS����A5�2���4�y��)`iYO��僡`u�$�?-�gY�R1�n�֍�R�!����tEfٗ;E�)�(KO!�\�=��� 8�/=�ɿPG����]����v����-�u��1�:Q��	���9���G���
�����H#6�?��h<�Q�2ѕP�,۷P>�����OT�w�惺j�Y�>,�<�����#�{H�����-�����sBϪ�qzn�L�l*A�~��,���HiS�;�x��)�>�66��"�~`0����./�{+)/�%�����N��0��mF}A����\���!!5"΋&3/C�~�ʶ�i����F�}ӨY3��c7�5b��R:!x��tˁt��*EsH�T�l%Iߴ�Qf.�R'5�_=��P&!!�Sg.q#Yr���fDgE�#뀶��^�i]u����g8� 9Ԯ�I4B��D4��~B- q�~�,������x;2V���\��Q89��Z��ޟ��(�#���Ǿ]�ڞ�b�w>�C�D�;E	�Ab`�bu<��)�.��ݏ0ۺ�d�@��}X���FqA�J@"���]`7+ݐ��ol�2�USY��k��=��頇�_�<z�`�՛�P�;	N���En�c��+��-�eś��M�]�0��_�6�Z�t�J��Ef�نvyN�9:}`0@��+]��Ï=�@8���I�$�����A�����?O��,�ƕ�Kw�eE�7�������#�j�qkp�����ȧw��}(��\|S�A)��|˽�m���$�03Ɨ�j����E����H��L�k�v��:��94�6c������nէ���
S�;G$Jt��,���,A�W�(�-�4�!%�R��q	��SS��w�:��`~�Pf(4�(e�E���o�,�6�M�Q�<�ܿ@k�OAb�~���sW]hg��$+�0��0��z������^�c�:[�}�FѶ��J���	�Yh��X[=��+���j	�YF�6 �ƛޞ�0�:�Ն�j�U�"IT<¯�R��Q&^7:'���R�`U�F̵����|=�6+���  �S��	dF�z��r�O!6j�!�T�^L���ni���B`����+��U����QxV�{@em��+���>�HN������^6R������%�*3̛ۭ�XG�?�����"=��04�R���g�1���a�.�8O����W����\⛺S��J��n��������عOouÉw*u��i�?h�����M&=h%�X�SaVے�
��&	;��7^�EX:������J�X��\MfZ��@���'���~d'�1�ăh��_)y<�`\�{����д�܇���SRU�"޹�� �j�	K��cvY#�@$�C`>�@�{dH��Ν�d�-�Rj5��=+g�u!̉�μ�u@p���S��@
��#I@�����:�<]�hWۜ�}Yg7rUfvhS)G<�t�N�2�w�)�� u+/�҄���Dfg�
l�����%��^['˙�C�Y�Wq!U�1h%�}�����]��������뗩*�z�Wa���W�5��U������ه�+�ݪ����ِ���}~rr�]tt�ZY���,�BU��Vn�C�_����u@0Mʙ
����3C=@g�g����b�L��f���!� �}�QT�ߏ��'��x���v�y���
y)���7��|�J�KE��g�ݨH2��Z���-�ԩ�m@;����X'c
��P�}�Hg_� D�F�����@�иd�����j�#m윍��&;Ť�8����W)�攭8d���� #T4�fA��ă����_Ύ	�4��HX^4��#艻�
o1ӕ�7ǩ����ߠV�{���`Ǳ9m��(W��t�"dn�b��~xQ�rJ�ש��h��ı7K>��X���7��\��G�(?M�D��}�����*����8��oa��8���T���}�x<Qy� 4��5���*K�^0H�x�I8T�V==o�Ĝ3��>=����/��^��8��s}�Lac�@�����9��=��QPޜ9+���W�|���_�3J��ₕ��q�5&̢G��ժ�dL!s.���h���bS�,H:���`4�s�����6��L&�T릍�$�D�S�*�ͣZzXI�y��FYkO��{iU��v�
���ԌW�eu��U{��n��î��!J������^%�&��t�Oi5�pE<��k�?Xu����"��5���'�\,�Q�f"�0��Шd����ƙ�	�@�4��8��ݗ��߃�V���2	7T�S��:h��əή^Jy�Kw��|���[�0��f�B�u!Xe`4y��b�	f�Vq��?�A7�L�F;�ܛ�#����#�t�Cn��#J���W&5�*����ЄpOLmu��PR�_��(X�&��-����F~Iy�z�V�DG�T�87l��T�H|�]����&�8�s�9�6ԧ$ֺ*�hd�I� �C��g `2��88�(�P�	��G��׎'���?�T=����Ji�FR��so�~cO�.0F��ƪB�1"�����B����>��A�^�w>���^��&�\`X�8�K�`iz5ۘz���p��*a(��FmYOk�-��;O�����&��Aw�ZA��>�D1�P�W]=�b��Z�'��F��H�ۜ���.o������9��,���o_V�&"{�	SmC�n�?���Mk��ЯB�S�����{�2�NU���,x���W^|���?�Z4Ͱ�{�G����ĚTvu������C�����e�Fӂ1�SVi2'�B����''���`S�N�Rl�f�N��됏�/� ��f%�sU��ʶ��e'�����ޑW�(�+�U��N~Eᵣ���D�-�kw��cU��vq���OX�8O��a.Xu6�P�d*�TZ�������k�i����q/(�4z�J�����C˽G3`��1S<��9txR\_m� {1�X1F�=���izQ��"*�"�"�������[�
�ҘJ�#$I0~�&Q���,
�V��p�s��=�Ɲ,}�
�МC�nk3]��W*�G�����o�_4#��ߧ�H��f.t����>;�Z'�V^킨�(8�����X�UMt�͏��N,G�y�1��.w��4c�ľWS�?^���������j�������rӿLe��m{3�H�x���l%�r���p��Y�s��\1r�ba��R��i��y�����c��w�Q2�j��:4rP�M�����ȈUBX$�&��%���)��~��1���_/_}͏���9�%�i��Fݫ"_�:�G���WtG��^5���[���*f�W?�/��`&���B��gUJ9���R@����c��(W��k_$d�q��9$(���ENL~�N<�3A�w�l�˒�E��o�������^�>��W����IzFO�����]ٚ�����	�7��P/���.H^[-�)N�U$�w�����ʷp�r�x/.^qH�C�Hw���f��]�|�76E��S�(��d�>��b����oCf��g����_ٗ�]q{����`D4�g�w��������v������k<������7�ȼ���Xk�8~�2���!.�Nls�M�M=0����z�m��zb#͔���/�J��"R�5������%ˌ�5�V<S�Hz�J�\�G"l&��]�󰏟s��ƔV��ZF�{����J�3���<�F�|�{�ǉ�ɩ⾒<����nn�ukIͭ����k߅ S#�XM�AH �ZKc�rej��kڤ�lU_�j�'�5�W���9p�ps��A��s���ٚ��۴�y��!uZ�%>|�����r�J�[Y(Pb�}'dX젼�=�qwD{>����}*T�+k@`�ǰET���_,ݔ̲ع�9���K�l� �ń�Oy�H��ΐ��DAZ��pD<~x����$�Zw��fC�;�H�����݉'ڣ���?|S#��L�o��u���P�q\}&�`i��<��m:Б�ǫo�c��2m����A��B��r��Yn�8C��kw=P˃.� a�U�4��4G����CMH7�|ZU�0�x�ö��8�dwU��0U�~uu������K�&�Xk������-���Qk�����w�ʼ�Kے��I��\�29�z�F*��Yxw0��WcZ���
0R����:���Gt��=�;�`'��T �A�}�H�v�0 �CN��P"���~<�'�8�YO��%\�
j�vy�>L��C��U��
�Jr�������vBp@@@)�Q�V���N]��
�&���X0A����4NHO��i'椰DQm���M9���`Cs+"Z&��u	MJ�y�='��BZ��&M{�d&.�Vl9�z1�eL���T��8�W���Ճt��6�Z�U�����/�Vv���]P�la�T&��g��v�w�}�t�X�
����k�h=��"��>iW�	�y�G��p�Q�w�~��nӅ�xp�C�C�>�5�`I��n��*~偽1\펠J)�N�9e� �~+[)6����<�cM���`ؙgPj��_��s��u�~��y�y�U�D��`[v�]ʞ����i��j�pRZPdH�~�C��8g��T�o}g��9��̆�+e�f�\�)���x�� �?�5���V>jA?�r:����8A�D���䳈�M�蜊����er���9�����WX���~�l�QnԔ�x��A �Q���y���ἆ����2�U02���4��u{o����ӱ�_��Ԯ?Mo����(_����Y�.(+�|����T��#� [F��L*�5.�Rm/��.��,�Fm��X�T����u��n��ӈ��)s�~{��G�,�>.�fɾ�1M�\�`�����w��9t>�"��Ĵ_�2�a���2E`��)�uX?E����d^A'���Mq���%rMe�f���F���XG5����0����c �I!�>�Ɲ�X��]�Ǜ�~�`1�V���K�E�i����jbn�4��v�lg����
N4�>��n�6�N��4Z2�d6m��zu�y/�݃�AI��1�E9���{���r�y!B���=��l�b'�Gů�8����v�+��*c54�U�c˕dnh]��U)��/vO�m�j1?�]4Hl�D��c����J�]D���������0��B/Rݼ/��r�Q�)���4�g(RzM/x���53�ȋj��_n^ZNυ䨁�st���.c�OLk���A�&��x�X�B��r�=>N����Ǝ�{9*�7	�zږ���-�}ݡrtY� bR��=�v6;�Jw�-��!9�_��I(�i���8�o�
h�D̂4�m�'�o	��]��Xf�mTT��$�|7#NIڦq�����
�i�Pz�y�0�t��/��e&{�	�ޓT��!˵���`��j�e�FO!Y� ��:YJ!�L�54��4e�'V��'7jH��n�,sVP=�����}��5��2�܅x~��,�#�:�Y��Q&{�����8��1��nׅ��*پI����&ǮC�S�D@����W�zC{�+��V�0=�)�L.�#��6ߏ�w��߲�2����X�>D#=����P��\G*D	��y�� p E����ݡC�Gor-f�@QRshn�x���G��6�<��B'�S���>(M�Ha�rs	�9�4�,W���ф�c��N ��]�R��/��c ���gF?Hj�9�w��6g�(G�ڴ��~,w����������O�z]�|^��a��͆P��a�w�|U��y��&�mx�m儇,��5e3�C��ܖ�O^7Ǡ5jm�S�o��V�4sZ[ζtFV������x��8a1�i唅Xv2�o�dn���S�����]-�[�*F?�����_ܡ-ߠEP�GH~�?@�����-�9��|¢�B/^��t�&fr#ס�p5��s`UNz��m�>Ő��ۊEd�e�x�Ec��5�������ܜ�ܚ�iY�ﰟ�m@��Q=t�y�0�[,���,8�s
򪺡�Ȣ�mvi�C���X�{��c؍!�%����>�|#��çE'�����)�ԯ��q���8	0]�z\��/ES�Z.�dBbp+L��i���2����%c0�}�����6��
w��U��������>Jq�<h$�-Q�� ��z��a�}scG��Fbz�dM����l�ZQeel۔�ih�炘Jktm$%������CP�I�z�,��×��oc��,��W�r�Z���H_>O��d�aF�o�I���;�N��,�.慼�e!�wT���ܼ��Z{��l�g�E�z��mrw_�
��ޕ%���R��Y��q�qr_�~X��[�`~�~�x�pũ|r��9���w\ՙ"D�(��g�(
��
h�D@4���U���H�7�?D��"�+\�9�f���Ѯ&�&^z���"N��D#����`�S:,�~����,�Y�GU�芡��|����*Y�f$*����G�BKTAͭnl�H�@��&lbJ�
���	��c|��KZ�����֌���NQ�@�U�p�e :ɒm�]��X� �`�x\s�D�hFN׀`p�#��VdT�H����<��&�Kf��c3rp�#��R���D�t�W�m��Mۄ�Y�"��9`8��G�%��=ʮ��u�0\�f�u:!�����۲�c���P5&�'>Y0�~:{��'L %B���Y�yӿW�	��9k[�ve+����a!�:�+%��C�v�Bm(ؖ��٘;�"���ڙI�q�.�(��Q�C�u��*���(�J�qt	��f�= ���(�s�*rj�oq�j'�G�He�����Ӕ�]������7ă��I8�W� ʴ�(Z��UR���v! 
���[t�@ߒ�ئLA��C;Jh��H�Lp<�Q<���*�����.+�L>��t;w�3=/Y�!����LQֆC�COɻ��(o��)����AN���c��N��Ae�_�ω�e��2��^U��-?"Ůp�������p�˨���+��X�U3Ҳ��Ơuy�~Ŵ����EXeuB�L>����^�Z4���fǷ ��~I�R�ˊQ�n.���Ht��ś��$z#��|�y��/�8��̆�f�k��c�`���s�߿׭�.���-@
w[J�^W�f��VH���bz�0��w���yz�°�7@�,����q �!ͬG�f�!��]*��Uj�N�j+�09�+[�\����`]��W況���;0��0��G:�Y���NF����1�8�N@ 3�rc�,���z.�l�M� b���2�?4:�!����C�
��D!��C�cWԳ1V�����l:6�:��Wݭ�)��#�A�.����
��Y#C"�F/���z7��HN6���]YZ;R���y�O�������ѯ���y�������07�jD�t,����[�u��zԴ�&,FdZ���u+��R�[�Q��uB+@6�HΎ�Ed<�yu��I&�cf�̰����a;�2O�\����ͭ>�4��v �H�Bxw��N�;|�e���ij
�J=�EcR�-~�ZGwcU��a�� Ez�	�b(z��*�\m�)
K��Јw�F�>��6�(�;�Bx_%���,��eΔ�>M(2�n��?�ڝ�+Y��֞ץ{ Ʀ}�[��_ʤ9$w�!s��h�vT{��f��5�-�Q�P���5"|�w'{�酛�>/ED��sA��_ec�cJʶ԰(�$)#��G�������ĵBھ]
��\D۝E���x{�J3���?�y��C]��B���R��c�*�V�E��p���'ty�v��ˠ���˚
�ɳ�Rn���.:�}�9g��G0Zu_1Ng�A��Z�s@[z�����(��ʧ�H����B�ۮ�g�n�	t;w�msߠh=�+��.f��e��M`j<�^��#�ߔx�i�	*њݹ3��E�Gs��[�?"΢�EX,�*���FrU|}���8�5�<��Ǫ�Cf�瞴�Ī7gt1Q���/��%���fG��R�#���@$^�x�>�\�(��١����<[v�`��&�zǌ�E�,���PzB����6�
X0))�O����X�k:Ƣ?��t�`�?<�-�:;���]s�c��.�#I�[(��4��q�Bq��c���� �$���E����J�VlWE>9j $<��f<c�K}�}�V�T
��#��A�J#���H��&�M�웼�?'�4����Hm���d�h�?�J�J3�@{	H)�'&qp�v�@N�����^n+/���<,����h���&�E}��0����G���iʮ�O�����=v�[$�J�͂n���F��N��h�e�Ϲ4R{��M���Z���i�yj1�I\�}j��I�&-� �Ч��n���9ld|�n����b̐q=_"I�� �����PUd��o�@�:R����WY�yb�.��vGw�/�Q���^��P?���^����b6A������m�{n�w�B.	���@��X�͎��ꮂ˯'!��R�r�D�;S���ԝ�b]쫸k
���ޢ�)ʲ~C�Fv9�g�@d����t�q��K���Ѿ_�;�4na�i]-E�?��˓B�0j:��mN�iTqe¤�m�Y+Yp�jF��6��={ں�ҩ�,m����� ��b�z4+r���;0ھӳcQ�	��ǴJ�y��3��e�'��s�҃���(�����?�I�\[�_s-�܂[�[z˗���� k0�\�+dU��NI���K��G�gS9b]����r�$���J���?]�qB{;�M��YH�`���77����$��  ;N�wGn-���x��(�|ŕ*�Pcl�!�陱�|,Ν߹J,�3��
OK#ckeх�І�G;yr�_�������i���G+b(��C������Ā]�=�m������}MK�njT��Kh_	���F���Ȣ呆96W�����lf$([݂L�'}�;��F��x_�'�Sb��̈́�=WNuF�âJ��4��$5->o>3g���zK��P�j%��*MV�</o�K+lIB��&>��~�Fttdis������a�[bx`��u}��Ū���C�f�ߌpP���Ё{��wZ�9�Ө��uԢn�f�y������Ȗ}}�<	�?��茂t�y&���Y���8�jF����K����I��ac"__��O|d�q�Z�mY�ܢ�����a�]���.}B�t/��Ƥ��7�_I��O;D��j���ݫ2VW��5���H?ꢺ��-�`�|@��{��m%�Y�(��|++d�3��'wf)���E�%bh�Ir�8�Z�,/ާ��鲮����,I��@��ߊ��_��K+�uh�|`��[iݝX��%����1����
��Eg���vE�k ����i#&O�1XG�ű=�m�)�mSQ5�y��\��҇����%��d�mߛ��fҘZ%���wf�G7��Jzd�<*H��܉���A���}�Mr��?)�m���Y\z���Ӎ�qfͬqAcu�7)E���������J�9\dY��H^����`��Z3ɋp�^�K�B�p�,�z�7݅MJ�N�D[lQ����_�L:k{����,/�;$K��U�� ٻS3pW�����Jk��o�� ��I��<��#�ҳ�U���%��Ҵ[3�5̹l{yuܾy]w8�7�-X_O���R�����ơ���В\�7��k�2,�-�+:e��z+0�木��<�1��ݾ�I{���7#�$����4����~�}v>:JX�Ut�ɷ�,F�ug�['�ֲ#�;@
ۀ�L!MX��f�s�zP[��2�~��tk>���tC����\�@��Ad{�
2�a:�U�]���6�o.w 8�+!c���à�)�EH[�_��r�ǟ\0�F��.T�И�6�����NU����Is�XeFT��k:��R(���&0��C�Ur�+{R����R�4(x���쥳�ծ��4P��w�O��ѢI+���QR�l��VY��
�ă����Hj��f�\n�)�0��j�ƃ�<���:�Nj-��;w�d��t-���%Xhb�Q�D֓R��ˆ3����z,�1���}�\l�,ܴ F|�˔X�]�� �r�X����K����%l1j��-�p̦�)����i��A�#	[�*�����儸��$%�?K[$�_g�>e�_�v-�1mT1?@��j�ZA�avyH�,B��^�U&H".���k�MzC<>��0�/3~�7"��n��Z�q0�g˄�{3��ʎ�*9�	)k+He��Y��� ���Y5�`|l��'Ń�޸kS��:��o}��,��lI&���Ss#%�(�����_	��d9��sV���Q��so:�YН�f�%�7x)�&-!�^��$|ж��䄹�Y��]=W���Ei/զ��4��M5٠k�����m�|��4����C\TG⠱͑ί�oY���jf=����6��B�q���f7��`�(���AM.�F)�&���2vea3��#~��u�;���3�O{�@)VS���۴ޞB��7�{������Ɂ��ax�Q�zF�zw|sl���
���^��^S�,|=D��Y�ȼ�C�?�0�N۫�AT����	�����L�a 
-�w�-1�yW,�:�$9�E���F�A��b��;/޷�"��[(D��w�E�`�̶�]��n�<y�ұ�Ҝ)u�k�XLJy�<������R�O�ro�����U�ѓ��,�Z��[Vg�E��8�dɱ��Oꈉ^� Ub�C���>���Gʅ�̺�<�ylmr%G�X�bܣ�-�����l3-9��~u0�M��[F��u�I����W����Q@;�]�8TD�Ǉ���B;��ʤ���M�+�!C��7�����JR��#�[����4K<����I���n�RL���}8���N������j��PK�}p�B)S�mk։E����Ϟ�ؐ|�mW�d�ۋ���Y;�;�F�?��!V�H�o���Z��6��l�S	Q!�ϑ�%�1\U�W��8'�[>j�W���W78E����g��:�|eĵ�tBT�wE�*��7�߂�D"�����F.���a+�)d�7�p�����j�vYi�47㼳R9ڡ��>Ʋ��o�(�vgd�i���/��BQ�w����1��k��r�$�v�ۖ��i�d�v�~���FY�P�>�E���@��@��/����Imi���܉��S��_�I����.�D)�������9��>�[��@���r{J�_�s �t":4q���+o������c����ҫ��[@kջ���������Y�y>���\�:!�튙'��K�O�Yt07��xG�4w�k�ނM���ұ�;3���t��WP�2�dZ�u�-��v7�$xk���\B������/�s7:��=�'�o��8��� ����-AB+KF�!�v������٤z�[{mb �Q\ʟO��׽�o2�X��ަ�@fX�h@�Q���(�uU ���W����0�����w�L5����4R��sZ �l���ꋽ�{ )�_j2��eՌ���36�$WG��.����qZ���!m�g{݌�Bu�K�-vH��c��5���$�em��Nݍ��ͮ�QE�n�G-�%���Dp����v��F�=������&�� 9�i�l�}ڨ�d�� ����v����!�dU۝�v	[�a��S�of�j�5�?���5���H|���f��ŵ`�oCX�v���0��2#�W��tʳ����BW�%5i�Y$�'�a1,X���k�^1�)��'�.�&\�:�3�A�[(��C��)��S�����j����w=�Vl�Ϗڕ�����9�EuH��$3�Eo�uP�5'gܝ��!�n���/'6 |(��>w��p��n-�b�6�9�����νc3a��K��Wg������aWq����f
;��H�Q�g��f�-c��F\{�-h��"	����d�3ō|�0��|��E�����J#(�V���U�p�"�a���p�)���ǲ��E,]t_��&1�B��w�#5��$!�b��4mJI���Lc9쐯c&�h��n���Db܏�g�<J�j�-�����9<����
{r*
�)�;u��ǋ��d�چ�8+~۬��AQ٣��@���y���~���$ɫ�mw�� 0����N b��:B��o��l�I�c�oBZ-�����3mò�u���Z6?���b3;�ͺC2g���%����bt����K�����\6p>Y�`��T Oc�M=�C������0����̵4�
]A�4!�w"
XТ4���Q�X�)Zh��<L�G��}m�`���L$]���F�ὔ�_?B�����R̚V���*�_"f"��w�J^AQ٨w#��[ל7a[�J� 6
1��{������M��B��l�@g�3K���֙j��9�$�4&���u�U"�n����ٵ{�*���cQ�!�]6�V�Ù�f�hw�G��;�w6�9+����a\9�	Q����,��\����J��_q{j`C�Qy�dC��X���(춥i�j���_����5M_v����/�)�:�gK�Y���æF܏�'�
�)X�OQ*A@]B�g���1bkC�Z�R��ŵ]��pW���Վ�ĉ���#_�B��� (M���5=�iUU]��U����&S�t !*�	�	K�7N�L�	i����]�c|yA7:{]�P�ǣ��L��B�WҤN�}�^�RT�[�x!�m�� b�Ԗz����ʩB+�5��(ӷ�S�y k���O�{-!j56����D�M&zV˟,7�<��$'�Ȕ�f�䇮��a��R����f�d_���5|�E�`�D!~Wh}��:x�8��������2�:�M��~��M�#�Zt�l�\|6��O���?��~[G�k���Isjj{�X'�.B���d1�Vo���B�;�ϗ��"��mz����]L8�+v�}�3�}������fZ!��T.}���& 8�z	"4��ܦ};��%(��'�}�B7��.�ѻ^�״��������N?���?��y��(T�x�\�Ҟ�V� ]\*�y
��N�jD8^��PG;��P�E�3�m���Tk����=�/Bt���� ��Q�0 �	x�ɟ�|Zk�!Z��Sz��t�,����xz�l��r>�mr�>by�н\������9��
Dt?e��Y)���%���q�Zܸ=���)�Ϋ�L����K��&�R���f�<�d��)�w��΍��%�)����~�@���x�n
O{l��e��
Лah��k��j�|:F�kݳhk�N������k�����ר�e/vb�i0G8H捞�0���{��3�T:�=�����K9{�V�_���^;�Dn∙x�K�ل�e�;���SZӚ���6ЮDM�5C��
�~�b�4��Sg>�\ �j�e�yvS��Z2��D(�!(��Ҷ��"���'�l��T=}̞jMɥ���`�]Ar)O6��`��#4$�d1s��;x{k�+�;�������	�v�;n=�˸l�	���҅;q���@�*�Ǳ�a��"��tߤ6�ET�I�>��A��~��!���W������b��ϱ��U6�f�◕�P�Db����,M4 ;�=��Ie���
��h��R֦��Qe����`4An�yd�Rͥ>wd �=:\�W��A^�m��(��M/+���TL(,y鋮3�f���CO�'��]=bp:�_�jý$�8��]}�Gϗt�%��R�uq��NG���Ԋ:�VX'=�|�ӟ�� �������7�����+��)$$��_N�2hBǋ���&�fY�������M��������M	��8��R����&9�Ce1�9��i��+K��݆�o���i�������ł��(<WܒJ֕/U�`&�����N�J���@��Q*��
�|�a#��f>,�q^��*�?H�O�4��g`?�Ȼ2�b�1��������$brY�Lz���8��:w�Ò�x�q�s	�~�z:ΟP@�v�uy[r�޹Q���6�nJ\%�l�q����`��R���)I�"�G�]��l �̐��c�����N�u]e�]>�Hhs�
!�j�af�$�������MM��^ܧ�E�R��Ǽ�_���BVg�QS���j�vT6�~%������y����ʼh�e�Y�E��݂�%~ c�Q�m�� �^pM�$WL� ���ߚ=S%�>*�{dпe@T�aTs�@	l��9��a�=���l��;�f'��a���.�L3ЖR�n�?���K
�;�������L��?�ƚG�_6��AƁ&��R ��N��P	SӬ�2�"�����#�������� �[�*%��p(|C�D�k�4驙>�#���e�ui�Q�2�����}w �e��)��5`�L_��vv���pv%v�����U���腂�Zsh��'�7{�a]⮂��ĞQ��d��3��l���Ǎ�]xo�<Y6���x���բ&��4�D�,�x�c�?�����J(/:����p��׮��pC���w��E������J���{�^��g�-�	����Y��W3��4[���P���C�����k�T�ӶṄ���ݲ`&��8i9���A�ۇ��F�qT����O����H8/��=R���	�Ih1g�[D���+r���7��&�����R�
�G�%B�\�k�x���RAٜT<���wDO��O����֟#�b.��0bݴr�mh��ݐw✰�y��Px��\�֊_U��V���?xI�g�S�=�E�N���U�x[��m�ͱ���8$�IU$��N�H�Sf2K�vF�3�Ȉ���ʿ�H eu�=W��0c!f; ��Hy� ���M�`�Tf\�
2j��+�Yچ�ܸZNYEV��4��d��6����;���c�ϻV˅v��&C�X����m��ꐨ��&����B�X��2�i�j�KE$P@�6,��+K�i�d��;�,:�|pM�G��ڼ�g���!0i����Q����r2�`
�/��A+��;��-o�x�Z�l+�d�kqz�Q��$%Nؐ-�����^�9^kvJ��5k�m�V�.��ȏl]S!I���Y��n��k��� ���b�K�p,��:��J��z��7��UN}'�z���Ue-֚�5�50�7@GI(�9mA��(|F�]?�6�[$��M�S����{��\cw�υ�7�Mi�ނxA~X����NH���:˩0�u�Qv��W
��{b�L��-�ah&cCKb��[ݷ��IS�04����{;]���7���gϼ*��H�L-I��FA�Y���؄��,$����=;�6b�P�x��C@�?L���(f]������3��tScW���_D)����)�\���ѳ���x�N�wOx��@qc���k,��M��*�UV� ���l�Sf&�9	�=;c0�>��H�>�H��u$!���(.8p�:�&��9�e0xm@��E��#��B�>�tؗ+�-�q,�_�)U3�@dr�����g��cSG�w`�@~�@�->�j�"��W�w��<�ϐ���7C���o*��#.	V#��]������FN�\��I���Z���E�X��WY�DՍ�K�>@%[��N'Tut)`@I�з"�j)�Z ����O)��ۣCI:��y%�V�)^!<�h)I^�f���Ri���BUc�M ϊI;�#GjU��v�lT�Ŭ3~-b2���R��j�9������9��i��%��E*$h?��s>;��"/���s��;\� ~��ȃ��+�1�J�L�E:�L��$�MY� �݇Y?]^�����R�>&0O���VNK�e���Wi�Ha� �UI,�(��i�)p)���~RƮ���#�����޴z����Q��6P=�}����p}�|j���@*P����<ɢ:���Xy�\�TۨT���ޞjE�Q/#�_UC����e;<���$�&"�86L�o7�z�d��È�Ӝ]�����ݔ�a�FA uw�Mw��c��wB�:{[��Gt��,+�		J���o�rs����d����E�d0�p�\	LZ�u����]I)	�����/l1<ܝ�d��{�C/��F�@�?����Hi^%��2aB�������?Ţ��7%\�D�|j�X6觅ʣ�{L��`����woL�~���I�j�J`��w�P0�ә�m���g�:n�z���O��Ū���7���zz�KͿ
�y�t]?g���öе[7)<nMg�;�Q!?�L\��<Z�ݲ�i�2Q�^O[D�Y�^n�c�q��:X�t۰r�X��y��Ů��$w!�Z"Đ�<���AZY�o.%�u@�����j���u�}�L�r��\��j;�r4��[��z�z�x-W#[� �8:��(k�y��Ð��OX_}lfY)�.��y�ρ#/�Ϝ��t?a*K�Ja��5���h�%�Nr��|���M �r�������$���r*ț}>G�m�->��]:����J���*[��\��81o{�C�'����\m��ٯu���C�:h�� $��1U��~b2����y/��;���K�4r(4�����=fcyK��ױ]A^�� ̏���X3.��?ô�'6�`���s����?1t���,�e9�!��
1��0�x�hB�U�����!U2x~��Z-����)�k�k�����Z�#d�y�x�w�>cܝ�*;�#�x.'�獳.�Zlg@�{��y�g�עףx��}�i?��y�$�I��#�����h��#�kH��܆i&}(O|kGV1�'\	a��/�,L���bB���ׂ���pAq�o�نR�f�"�PM1ޒ�w.r.�(�B�d�ɭ�U B �(���r�\ڎ�,�.[�K3o����`J�P_=BfG��m!�L�FA&�AWm\��t)�]R*�t{������g1�ӟ��	��Ci�+���>�6��Cro�c�?��Z�`S�3�*Gy�u��eG�~[���-%H�JFGw�S� ^G��;k)7$ ~`.�������:�����q됂�]m07x�d#�	9����M���Dj��S���7�[��j��������W��""w<O��<K��n���+�+��~I�%���F������m�΋[�*�,_�B\���<����}�٧�I�w4���dX�IX<=�oX����ڎ'�J���\�<21�����a՞w���?��"n#3���k7���6�R���E����[��D#��(׻a�ޠb�q���e,B��xIG��M����9�O���������.��cۃo�"�DG� ���e(g���U���ʣW�%�\
�l�����26�"1���S���������f����:QZ�Q�i�򭁳n(?υб�3�mf�A�;)
��,p#�U<h����lpʊ�^�'a����}sP�3���(�=8��`+�{���6|��@k|�����o�E⢴�#!}���ի�{�`B�eL�K�v�?��|�J�'��4z}#�3��h�+�$�!��xa��6 IW5N?.E�{DT������d?T䉆�	�0�>N!h! 0�.���\q�8��{@�oyi�Hۺ��w�h��{�NZ?�N`�%\<�cR8>�u�YxS�w�k1���{j)�r�W,l�e;˪�Q��s'����>�>V2n6f�#��@�1��x�_}�2]��FC����L��?<�}��\�ڂEM�-we���QPӝu��[�{6x)�+�pqC���pR�P賄�S�σ�I�Î�~c�B��zt:ܔ�y?I內4��{!�JMVjꋐz�@F��V��`�&?�K��X8�_h�,��k�C��̌&9��Dm�C���
~�LE�A��ܼ���-�Pa�5�p�.��$bo�0o(�:J��%>Ո>��P�̨m��K��%/Uϵ�3LK��`&�%&���wr��*Tx�
A�x������2X�N����s�9���ȯf�Ȉ��n���Ʈ�yk��(�n=�r�YC�?���n�*-GE��*AP?���Я�L�[ZxP�k|�;�*�#�
s��������(w#WiTY2�z��Й��siLdp)� ���Ѻjx`<4���KA�2VúnC�(Q���6�u?�?	��ˌ��+Dҕ����G�;/���_�K�Gb=]�����g�/��e���2�����gN��&ޱZ[�2&�ǀۛߐo�Xed��.�7��1M���n��wCv��/�m�ȏe���iٶ�u�}꽕��kM�O@Nfy� �9����ഔG B'Yy�vv~������]`�G����,��a�*����E㗈�8h��7N8�S
{f�C�N�C���=�lT?�ՠ_�ԛ�R��m$�
4p_.��ge}wP*�w?AJyH�+�C�½��JC�4oy����RW��D_bD�@�.s����q;Q}�>��3����������_���qk�\W�b1ja��i@�E�!%tL�͟���;\s@K�Z��1�cQ���{z��脔8�j�k�����_�.��8iE���,�b}�aH�o�l�ܑkXf �p�IV�����2���be�={2TL�T�����W�|�p~'�G���E��s#�����4d,�[��d����z�sKg��ݒv-���u�����4���}vQ�5�5����IU/#e�/NK�dl���.�	.h:d,N�>E
vs�͛f��l�+��Lr��ku���x]a鉧eN���qG�)��� uѽ�J��b�2�����ً�m�䊭���V�~��!��<+
�*l>
���^��"X�d�H//���M�{�pC��O�N����e���!�ʘ�'Z|-���1&�y �0D�q�{� %J����Ooe����M�(iA�f�X҉�
�뛏�0^���.��/�yȇ��i����M��y�0{s��8��3n�{����ҹ�6�af��[Q��?2����:U3x��_����#6��b����m����D�R3�\MvJ�c��
�Z���m��,b{YI| ��)y��'?$_=����Cy�=!��5�Z�r��~_P�B}c���&=�-��<�}�}]�ǮOU힢P@O�\ANa82��9���M)o���'B>$�S���<$���\�`=ts�S��M����{�%!�("U�)*ӅIR�6�O���0�?g��v�_���=(���O����d�IMIK��MP ��3?e��DI�K���`����b%eX9`��T��3���ߎ�ro�~������[��ߢ曃�2��$G2@(U��f2J�iP	:1�f��u b�Z�nY{Q�j�g0^�V�h"�oUy��6�pv��É6��(�C�����j�yjc��Q�$����"��S�������Y�["�*� X��ލ������@�������ONƸ�f{`��(O\\ˑ0|���k�~/��H�/?R�] ���9;Gҙ����Y�Df�ʈ��<-�6�r.���e�Mt��i����)���먝�|�1�z+�aΠ�����:����+3�j�r3��H�8L�v;l;t�޻x�� ��W��¬"�h̀/��)�iT�w#VQ2/�.Y,ٕ"�i�l�($�|��/�(� 4���	,���G�i�)*5�y�ө��,�:xy%� ����8 �G�eʫ~��f&q	_�G�7��eÂ�P��8����%��u�P-�o6��o5�}��z�DfP_$z �������	��u�3�̚¾�l}O�S<8��߅5��f�#;��/��(k�����?�q���EA�MGi#��_ ��&.�`�L0w��)�`�	��,l[i�1o�`\�߫����x� ��!U>W���F�=ػӒP8;�}��TD'՛���K�x�d���I]R�]�En�e.�8��[m\)������18��؁���`�T�E^'�2 ���>�p>��Ђ�ک	 >#[����͜�Ϡ��!����T��if���px�e� wMcH,*|�����ݮ& ��;�������Y����@V���P\W6_gA �|``��%��QOk#>�觥�����q����X�[��>�ڊa�>i��G��^��hg[����>�655ɻ���92���YÌ�e����f��_;����v�M��oE�O�䔺�HJ��E��mD��I�>�d$[Q�XȚ��5�������ٴ�����jw �K�c��= �6��	��(;.��/@D)u��}�f$+SNe)����u�}��=�к�G�۰�qzrM%�9���� �� ����b)�4D���P���9u�f�Z����~�$Ќ����f�+��T��i�7_q�-��"q=��/�����8��wø
�O�����$G[+S�@�(%d�x�G>���>�X����Ư�cHo�d����j˵�����AW�5��jpL)f�4���5�<�)/�)Y��ru���Hf�}� ���-k�}�*�e������O\�	rw��OG�)cM^�ե��H6�B��`��.��ߦ�������K����+��wyQR���5'��2UPe����:�~�IpM���5�nu]<J]X���O6�@7��`uy:҆�'2�c���e,�a�Z�d[�[�"��i3bH�5<����9�2�����=������k���]������}�y��(!���3�Z:��X?���&3�<�d��\��"���T>R�hK��9-�K�?/!a
g�K/�����q�2�ޓ�Zq�@{�}1�p��䊂�1!�~2���gѸ	��V��:��x�Lu���q��	�>~HU���m�w�<��4}*�)�݆��;���eá�m��o�B���(2Wa�;])J�)�Y�Z<Ψ+�G]�n��ȪBd�2�72ڄ�g�f����GL1�wZܝ�$H��D���3P���86��63�D��0`��ȗ`Z�o���Z��e_�h����j�ʷʙ|��~c��(�r�%�[��T;�6�1���]���A�)��Nv����ɵ?���R���I3Z��[��k�Wb�}Ɖ��M���36��y������뗍71Η�B����_y���X�40����ϰ��h����ar"�O���U�<2����f���[�(��:��v
���r��%��[H�D���(�-fF�_��`��)/���V8���Rܓ�/�֢�^��))�78��xR\k�ZD�L�Ǹ�h�27�5�>6�/�C��H�W���+D׶���Ȁ�ܫ��2�i!X�`��p)Xx1n�&Q���6�ʗ�:M��R�	Ξ{���%e�����X��\)c���u]�	~�L��S"���m#�a�[�H	f�*���0l��n��lg�̔�#�lu��-�	���v�������3���º&��lA���2J*���sg�شq�n�$�y[;Zs���if�6=��l˭��D����*�O�}떚m�n�F�O��M��������ٳ�fd�!�� ������v�����ض��˞+= [��X_�mxk Q��QS�n����ZC�hNA�и�}=>��H�����G���󒷍%
��ס (��@��oTQ@�V����=P�ۨ�1y�~����B����p�b���y���h^jp~�3��5�N�+�³���s�4�n�4�iH���	���a���Z�{����wSy�,O#)��4jLw��%�o+�O jh�{�!/�ޢX~�o�߆{�#��1�����t�v�ѷE���&]��)��]�������EDhd5�q��%Ș*&�Q��'�
0�	�9W������}�3�!c�j���*bpq\�6�d�i�����{%�J`�n���9{��8��}���2?x]cM��x�����O	�!*��GkL��Eh�y�yOݰ��G�0)�Z��p�v:�L�VT)W:(�?�z��~.�P����j�_���X��]�H����������d�#x�ZY#{���=�+�!��*y���f���&�N���7):T�)�����j,ٹ��^�Z�0��,hkb�����8K33)A\"��'�M�zpt�-�'c�3r�'$w��kh��C_	�����H�[�S�ec�c�S$�p�L�Y��2*vꎊ��18�t}�_��U;���r��'�]�y�>��cdib�!����Mb���ܽd��4qo�lN�:�����Y�M���;�pi�!�{�(�f�C��-n����~��q����
�C�y�Je�mO��M�������B$��^����l,�B%��m�x��i�1X��#k�f,D:ҝWR1ٰ�V�@��џ�ċ�4W��a� ��!��~�wMD�6�K}_!>%
V��*T�(�)|��9O��[Z��.�ΫQ$ʙ�no��7ʁ�?���a�?�>h��ۈQ�CPzCb4'sƨx��WA���$��(���k�i�{��n�Y��_��������+��>W�}�m�bD?l_f=��e�1���[Nz�ߧp�}�\_����"4�tWP��~�N&
��8(��F�g�+M=�b/���o���!����sc��X1<���������;Y����f�m~G��Z&Zw|�D�3��S��8�eV��a�0���� k��8:�Q!�~����3xjAp�>O�^dL�ph0�$w���xا����>�Q�g�h_�/
ߢiJ�9�����$1Bֵ5"��y�g��6�;������S��Tv���,��0T��%C��s�Y���mI�e�)8�n��8h�dC�1�[k��ಸ��U�lڦ�|F{�|/���IU��^s)���胋H>�&%�j�K�t�����8�S� ��U����-��i��!K&�gdM_��-�c�nUYa^W�b�T#�y'�5�.���Z�M����?�/v12�5�}g�G�f��gD����x��K�B�).�8[~����Q�%?IjA�UC��+V�V�u�8B	���{�[��8���� {�<}6K����a�� y$"s���m�_ ;f�@��by��)�����Ռ�c�;�s�r"��L�������*�/�tU��K�ú}���`��@��We��������eC��#�&	���#���{R|�p5e_u��i��de�y�D{H���O8k؀� ��R1�ْ��[�X:�	�-��������'oS�{�U�J�ߐZ�PԻ���A��z�s�pa����/*^T�vB�{��fj��\GH�s��2)7��L�b��W��[�j���c�+�2����>�p7���I�+���]����+vtz��t�I�"�rH�dcF��9����ҩ�����$!y7e?|��F��.I �K�n�^����bZ������;��<O�m���=�D@�#<�,ڱ�o�L6�<��HS)3"Q��cE5>3�J00w`#�1�awm^�Sa�]ՠ��*�	�N��@�r����RE>knXZ�Q']qW�<�C`8Mz���w2�wa�['��P����9�`Dݏ��P�������J�׭4+aɐM�G��:�f�������Fe �
���?ܧ>T�;rh�P��]�Ya�[�
$�-�$�u�R���Z���"�23sh
��&)�]+������~G�|]���zH���Ƽ迎>��
�����{V����Y�����xQ�k���i�7��K��7��.D��W���:G�wp���LN|#��`�vEF^�eqp��)%c����1���f`��%��$SHp�K���^q T��׽N��Q��G�O�@�z����KM^e��9��ϒ�S�*�*7�­r2��L!���Y�	�o��*$��o�`bJ�N�ʀ�%�fT��ޫ|xp�	Gqd��&�z��!�^�]��(K�J�ZX���b�d�),CH��>��Qdx����u�~wѝu��z��(Z��Z�$��*�w�cn�&���şg$T���	dh�'�� .`�9'�؁r����q�b�ꭐq�w�������y<��T��"З��f9��B9Pr9W��I8<�Z�*B�a�>��*�I�I6�u��
5���D�"��5�jX�F`��E`�����q�h.s/�ެ�<d5g���3�J!�z��߈�&=`W�l�lV�|�$iL�N?'�[�T�C5����c�CR����0�
^F�T�c�p����d��Uf�PeF�Jbz,���9g�E�ස�S����F?&e�z�����8�}`�ب+�;j��x�iݽ�%ħ�g9h�����t�e4I��>a��g�z�\ �g�J5�؅Ɯk�?)�+A[��u�� ȥy�G'Q�3؀[�55X
MQQ	�)�\�CLKB��G���2�}Ҧ��ƅd���^��ԁ�g0�vւ�;�~�5�[�r���Co�;��U�gG�zkw@��������'R+�	h���yw��X(8�鷴�G�Wo3TP5����0=�����8V��К�Q]oܯ�zP�O�km�D�K�	DЏ���}?�Å���}g��2��N~��tī��T��5�=ѹ���\�ݒ��n�QR^�{��ś-�u�7L#(q�-GS�A&�e���#g\���Rf�XY���Y���|����ּe,Xs�vG xw�f�\�rN:�]��E"�8/���T#](i���3�8d:�A[�����y}Pw�+��*���N��N?����L�T'ͳV�6�I��;�î�l�#�.d�`CG0�������4ے��K��>�Ґs�;�iV}:G���`���#�LQ���ǿImD�\8�v����wF\N8�៘AZ����v���s3p#�(��],�u�~����aG���˶�Z *���yE���-�6��,ٮ���-s��Q�7����ȅL��z��>��U�TDi�5��-���]�0$Z�E���㧴�Q�(ĉ��x��f�ʁ��u���4XVE�_��1k�p�(�w?./�����u��`9�.�AԜI��3W�]��v�)�v�����o�S��X[�/4V |�.�Oڳ�g; �C렘��)w�v]������s�QL�PPF�Z0iC���d�U�xst�h�sa�`�B����~e�^�v��H�mU�1d�ں����'�����iU�b�WB`��x+5����B�z1_�$�I�|�t_2JӸ�:K�&9���G�8ٽ�ܿ�K�ma��{�M�$"ɜ�M�z�:*�
��+a�c�녹�ت�0�R֛�>�{AtcM8F�{|�D�}�v˓�D��i�I��i���S�2��
��I�� �`�
�d�V�ː�ތ��=��{l/�ѐ"y��Y���Ff��@�����@'�k:�ɡ���8����� O*���Zzo%�يQF�_\���*jF���JI_N|�XW��V���^���ލU�c3��4ܮС=��m�R~EMd����HXCE��v��g1���<n�V�W��X.J�P�MXp2 ��b�-�W�c�|t7N(re��z��*�aM�;i(u���� �7P�}�6sw�Kb�}�ʠ+���5g1F����J%�7\��Oh�a�9������| ��oZ�U��k����w?��'Q3o+t�����9յSH�1���|Ѐ��C����7U��C�ec)2y������N�Kh���`>�B`0���Eh�EOD��}����c�\A=���0�����(�P���7�!�x�~/��{�M�m�2!��s�6�� ��T��qU �׏�#gf�����2��>�[V�jj�L����LN�?#�1*N{��[h��;x���4E�t�y쀨�A�C��f��N�Q�pej�B6���Br_;m��\���.郔�L�����_
��~�=�p����*R9KVG��Q,�vD4��j�Bxv<�=��	�B��D�Ӧ���q7
��/��F�'�'Xʴ#l������u���u���"QF;�E� `N|�%���%�x�Z0�?(tKeE����jl�y38�HlΨ��g\�c��d��� Y������:5�8\q�� �~���	�F"�,���)ٝ u�}�+�X�DC�R�5�&y�hc^٢(���Á ]�lxY<�ht���o��W,��r6�V��3P;��3e��weL�6	A�t8[p}7�TхiDJ��R����0ػ�7��F�z�?΍e��pV�m�Ҭ�$� %4���>
��%#��Л)"�e�D��p�G����,0(���hnӭyw��(�+8�7����]��B��*T�t���_���A��Q�A�r�]p/h}M�|���s�8�ǳGf��T	no}� \�g�x����EX�Oa7�H��&��E��xNf��^@�G���dؕ���q�g���<�ʮ���H2 A�F��Um"ߠ	2��R����Q8�~F ��v�-_E�������#m��k3T�7BZC�����	�r�U����>��mW�Mh�ݡ*#+�xeǓV���� �}cs)�,hz�`�������R)���=}VS@zaoF!�h��A�]��E��D�f�n�xn6�W��;�6�[y�*� 9	�na�zɌ;L�̫y����@��ތBk3Y��%�9��x�? 7"�﫦_O*r=�
b�D**�o�^�`ȭ�%��6'�[��Ӗ�
���U~U5쀄$C�ɖ��,�����^�gm�3�����%gC�p+��%���]� �3d᫏T���Vc��Ϗ�Cl
.��?��WI:kb�C�`~�Ç$'sY�Q�{���ơ�U&�tlX�-ӱ�)I�P���z��5�l`�3�Z{w3��&��qw�H��NfS��A�8b����2� �RL�b�l������e�����n�5s�'� ��-�- ��F�p�]�sR��"��DF��^��%�9'ۖyNha
����+��h�NM���2!ֱ���&q����Џ�w:DCyKnb��lN�����w�M�G3��#{3����p�K�X�_̡(�ۡ8�S����!F ���u���?q�2'�'�KE2[��Ji鹌��gJ(u4��-�ȣ�/<k���O^D9i�y7t��e�k����A(s	}��+c�H��䙯�?n��#�5�!�ELucoP �V`��y�i.�����H5(�i��Y�=���D	؄V��P޾��	(�a��8f6;d*�E?�Xb����6�d덦�^��(UȘ�:���l%xc�� !��7ፃ���jm������#�ZY.:��B���U�Tp�f��G�o��ߕ�HGD�㠯�|
Y?ۄ4�[�em����K���z�����F��NӬ���~}������g���2���	�IP��iy ���[��rK{���iZ�	�Kg�}�LEP��9OAs�F:l��:�Ӊb|���<��a�M(<�ԐpȵC֨�K3��u��<�g��M��2U��?��Z\��b��s�Pd��Ә��U�(��PxoM�,[��N�1��3��O5u'^�[�M=-��M��WAвb F�D���!g��f+�b����ǝ槲v�|7�9_�WL�̈́8��}w�~9����ZP�Y���+
&�;=Z�c�z�V��1h�l'�缾R�{.�M�2Q2�OqP)6�d��L?( ���#�*X�2��oO��D�u�q�ZKR���g\n���	�C]��l��d��ri�R��R;�ü4�7�E_��D[C��H%M�<�ʐ�=��N��f)���s"�<���\?�jp&�`'�ߑ�L����!XKN`=O��2���s�݆��<�_d�:кW-9��pS�3�A����	�g�/6����)�T�4��dp��.�����p�Ӯ+�:.0c��\x֩��s�����.�;�_��W#��H0db5zj�&�Zpz5�� ���ˈ@�5]V�=x�9���W�<��bܪ1�8h�����t�t�6�C����U��6���Eu�ŝGT�\����9ſ�c���00d��c��UY���&V�k��z�1r���ґI�.�LOM��>��3:Vp�L��2M���@�a~ncg�s#�q��mYe S�Ԍך�s衵mO$iU�D������T����<�	uf��D��j� );��r�.bFs�(����������b��ȕ|�?�_4��Io0�22AC5���
�����1|�|ݾʤ*��M6B]m���<�F��#X!�p�v�j2�xj	��A���+��h�'����\��qg6�
fH��qe�1_0�5Z��M�/I�U��`��ir��qE���@O��<�t�tr_ԯ]��o+Tۑ��e�4����ܶh �4�?'�l&w8�9�7��H�m�9D��h�ޡ
V{�p0(c:�
�ʺ*�Y��ǵ��Y�����Z���=:y��U�����!U��5r�p�2B2 �gt�58�ʠ&/N֒э�'I{�@�C���9��_��¡�H���.-�ݵ '�)R�X�+��97�k��0ι�4�΁lZ�r�!!���V�d
�fu�/��O*�"5�X:��)ᤩ��"
�>�af3��b�׻�#-����BT��U�	Z���%?����l0������U ��7x�Fs���.*��_R�KK��b t��}�6ysD�E��i����0X/�;UM=1�'�-A�s �����rc��-բ�ŽI��ՠ�L�	���s���MX�r(�%�+�E���dEg�v�<C�_��&�z톰?Qܐ�} �~3��C�w���1Y��9B�]���vƘw�N�	GK��猁��z�`|�6��L�?���X��豋J.���[0x-9���i' ezI�-p�����Q�k�C���������i��rk�����6j��d�\U�LP�e���c�6��t����ZH�eJW���a���O<wӷ�Z��ƞ�@`�^�T�sѵ=Z�����_đ�eJQ�R��!�t����񋃎����6��J�c��\�쉧��	�5[�k"��`eƊv�i# ��QG�X?�+7Qa2���3��w�o�<�R��R5��z`�p
}tu����r�"4��� �9��E���5��|J��_��zɽ=t�=4�}PKI��ٰ�9��	_�rJ�N�P٘#&=�V�cW����m��HOK��c��j�k4Cy.<�Rx���S�D~ۇ�G���ɨ�&f%ʫz�X�<E��<�td�t6�`%
F��b�
3��"m;a|�<Ut��_��9�乞v}���lꊋ	G9�䘻� �Tg�<�����pn�AH
uKa�E�wk`-�C�W�v�+�]r�1.�}���e�ްW��� ~��C˶`���RR9���jc��W3G���m
x����T�D�7A�˺o�j���G,�G���4iz��i�Ù���l�������R���ඐ�<�t�P���5[p��O�=���
���f�,%'����5r)G���ӧ���sIǑ�Z�����|���M�_�
���rw:�UvB�^	oQ���`@�Q�@������\5�oЈ�g��=��4�j�:�7.����H���K�]8����
����T�u��0uQ����/aJ���KѸ�$������%�i~2��i�~��:@w3�)��;?^�)���m����Jb��pq�b�|NѸ�I��gg)eq��5���3�ӻb�K�`n��6)jy[�j�e��Nq��%���{��h�T�cUu�u2Z��+I�4YԖ?b���y�"a�DM�Z�E5���\�Y1b��"<�O|J�����/W��:�����u����T�о�@ԝ��T�D}��?��(���
�{S�h[S���i��:l!CRdkF\�+A���p�1����ƞ�f�&�6!
hK�"�E��;oOu�	��wb5f{fj��T�
��i�-pε�L�J�"-P|Q$7����|���'+`" ��p��;��y�x�o$G���1K���Nw/;v�5���d���3� 8��V��J�����qK4�D��ש��i�ȴZ������G%��8�\`����i>\�Y��r�r^���c�x�[d��3c� �ad/�@V���b�6���&1"'�)���"d� ,/�7a�{'� `E�/�Βb,!q�t�ȸ�{���~�}�R��#�&�Eb�?*T9N*���=+6hA�2��H10X#�%�R	�(4�%c��8?��x�)BʹȆ�o��rk,�{�lۉ�a������kd.��)+���}�P���r�F$��M��)���vL�m���$��*s'��^sl���i�Br<L��i�D���pQH�3+����h|��(��ڒ�׈��O�	ڧ��2�6�s`Զ}�!@�C����ə�L%�h&�ʣ�>�{��M�p�%[�N�
~U#�5$X����5���٘@Un���t�Z)���/7�D�Ur��U������PP�,�_�/^���U��v�N�=�t
�g�������-tY��	��)�H�.Fr���lk�3P��
S7[�]�;�m� ��_�+A�K�D+���F���/ܔ�j��ҙ�_��.!b� KM�#T�
<N>%���rr0�M�Nu��Mx��FQ���cڇ��C!&Ւ�8�����bp�O}\3ˈFu�B휊	�ƿR�ܫ����1f'>#���3N�O���"'|�f#�U��Sɰ>��O���R�D�6�����u����3Y#�x�l���xLhh&�wz��ڄM�wF6.�)�ơh�HeA(�����A����h�5�Z�ZVų� ������vD�����K^	��WP~�qI��۹�g�2��b.Z���<�Q%�rq�.x'}n֦�e�#����М����r���+�1�q�0���i��x0�cL<��ωf��1r�����3������]�f�۵�4vt��hruu�+��4h�l����"b��]�M�^��K-��+н��{�~ �"�LQ�W��y��6w�wC��V�VVn5��/g\����-���~�ҡs�2�� v�7^�x�s�r>������W��_��r�>Jh
�w����x'J����5��V.�e�H�QK��UG���l���"U7i)��~~���ݡ��� �u�D�V���s��}x�� y�����ք�)�{�Nr���	F+�ԗ�^�Y4�82���yW{	�F?%��� ��D��u�U|D)�G�\}��8�^Q��0���Yq��{�����&��h ��͂�.�������!nܫ��'߱yN��ԓbȚ��5eե.iicbk��*(`���&�g\��+�u�j)�v
��S4H��3mT"���4�Ւ)n�1ܦ�7�p�wL��J�.��Ѐ{��=�-���S5ԾW�-F|S�]�!�z�d�� �a�;7�}�y���d�xN��)҂>I�hp�eiah��9b�jB�iW!h/@�!,�R��ȢO��ݳ��PQ�!*�I/�
�z·M&X[��:�}Q�kן��?�'���9�ʍ�sH!�$Qي]���-������T�o��c1�5c0�X�.��Q{ZH7�1ʕf2ʓo@����L�#躻��*7VCh����4�fʍ1��Ķ�?�'��\�_^ܡ��B�P}�u'e�s�� ��40'���Œ����ɏ����4Dz�Ke��c�A��%�P�����'n%xG5��h�z�{��W�G��Ŕ+�6�J� �ۼ�-���u.L�Z�<-�𦡆3TVj�|BM{Pc~_BZ�)S�5�ш�T���(V'�4���,��/e/
!�:��W��w,[�]8vV�̭�j#8�5=Mt!��n++��-���gzr|�hq���p��S|5Ò�hIǺ��{�/P��X�R�a$�n_�	MU3�� $�$٥mZ�/�4��z���&��1�� ��h�7��̽M����bi�:"�2��r~.u{��������j뗊K������̭�д�S��n
2A�D9(�j�ٷ�w��c�xR����ǭ��p�0��=Z�Q���L�]+�u,ևi��t6��es��L���Si�Z�gv����Qh�b�������	�Qד�(כVY���0�J �=	t�dus"XJN��}	F�1���q�W�;&C�G#(K�+�p�^�St���oE&��Bb�\Q���5�9���8{�� X%�{�T��c�DǑ�����zSH�_�^�Kݗu�B*�P�Ԍ��i����.b��g�n�kk��U��-�㜴�b+����祉i�?��s5�)Ҧ��D�ρG�n�t`��A��2ؼ�)����0|[���Ԫ,q�Q�*��F�C��rQ�9���N�؞:��P'I�gvڷT��Ιygт@�hcPW:T�����GL����nN�,�Ȥ��7� `�C��V�KP⾶i����GV�tt����3G�<8ޛ���[Tjb�;R�����(e�9�V2tɇb��#景+J%?�(����:Exo9Au��
G��+�v{ paY�q`g�7d��T�
��g�Q6a/�{�������:��ϑP��w��,~������T:���p�e����}�VQ�
��J*������<���'�=Z+}��wތ(���s�'؊ �h�C��\�c����
���
MOc�QXM�Y*Eڔ6�LZsI)ڰ�һ,k�N��B���ύ�~��nT>�t�0+4������Y\a���A�&Q߻���x=��;N�M0����=`'���>���	J׮	�Uu���X��"�4D��mh:2�r�v�TM��T����Ɖ��5����9بt���垲��v��V��0>���`�K�雂|Ry��؎r]��BD�K4�-)LD��W>�,c��
�Z�T;,%h�7��r@Nl�ڣ�pV2��{�h�-p�M�	�F��Vτ��b#ݘ�|�GO���8P4��"�)<=���3�&������x����EN:�r�MT�C�P2����w0Rg>=Ae�d������֐�t(G�/$I������#�?�v��i�[/��.d�Ԝy��!$��Ʋ�B#��Z�7�&�2�Tj���n�ѫW�K��K=�#� �K!�K��1�x��J��UCԒװ~�}���1���j��� _�/b��2�P`�!��(P�(����?�j��<648=es��+5/*�w6w���i:�j�eÈv�@�qi;|)Ơ��t8�����4�:�¿5���|j����l�aX;��2;5Yu3� ��$�����Ok�pK|_��)V�q�/p�gf���1�
k�0`��I��PAxm�w'ـ�g?=�8� ���R���.�S_�s龽&��2	��� �
Y7j�����jb	����;Q*W|�ğ_���j�����5��ސ��R��(�`��B	bM��hfq���=`J��SН��y��R4KNʜ��ǈH��K���Z���6ݰh�ۻ�hh�9q�"�1FqgB�
l��~�cdm9j�[���"��, ����&��$����{�N��Uu\�k� ���]�%�4����~�Q�����O���?|~�cƵ��Dx��, ��	�
B姉��_s�a�`��<�cv6�{J��p�S�8��+��I��g�qfua��-��D�l@c���}����t����F�o������ˆj\�a;mb��I`0�S���q^ϑ��;gn��"�Wj�YQQ�9������~�q2��jUu���R��'w�Ҕ�&��ϕ!��T<�F�!9F�	�{�䎽�%!��Y.8(3;Q:�%�X$��ET{@p;�5@�'L�{n�N�X߲���̭M����}��X��������$����� �o�[�>[	�F{$�s��z�G��sVq%��D^���7ȖE[yCBâ��t奔�%	��Wb��>B)�sv��cd��L����t��`��������w��'��۰Z����~ߑk�ϫ�WrX�V,��5�e��[��!I�YM�0<r��<yQB�6��,��� {X_��������6,�@��	�r=�]�g�����z�����*���Ql�t�oN����.8��f9����a����!�K�����HW�Ź��L����q��x��l�y�3�o�2+K��P>[�H�'gFn�z�z)(=��<R��L��#����Yj���e/�0��jL#�ݏ�$�]�2����L��O&��\���*˽J��S���9h↍�I�By_w��ɸ>z�5:��F���������9Ɔ�D8�������<�I�_z�q�c���X	�w���V"�q߱�dM�д,�DP����C���|R^����\�&&��Hrq����
��i��s@�\�zc��Y/9�oImXY_?o��E-׼�n��v���P�H�T��(no�S�%:y�c�#mFtL�����f�X¸$"�Y$R�Y�e��q�'=��L��\f�V��y����>��f'\�b��'�#�I���Z�)E{d_��i�@�g܈g�����I��A	/�?9JNUZ[{rE,�59��U�V���D�b>S�t�:�>�����-J��5��^4z�I���-�`�z�.�J[T|y���Y�[�q�60�n�&�#����,�4ᩌ������|���h[M��:�/J�	?F��cř�E`�K�x��cx޼��q}�</rp��
_�~SD�P9�3@����Q�s��}o*4����G���54:.T
��D�"PT��:����5�O*�����t�PT5�s
���y%���4nj~�-aG�1l^��1-��1f�A\��.F���!6�ݏ|O��b�X�-�R� �_d�����6�S �T�%����$��PC���f��݋H���%h�� N�-��8�X�~K2H~�k8y4/�|_G�w��$�pH�����>�䛩$�bo�m��&k%����x��U�݁o�,lJ� ׮ܺ��u��j7��hPg̀����&OM4[�U^��'�����ڢ1���<�������I�?."1:��a�	�tM0<wY���Y�2Fj��: �@giA	J�;�r~�n���!���aFA����IKReq�6�h�˦���씎t�����M.gr��&��߱��9-
	��������N�M�e'�\8ulXMi��lrv���V� ���P��Qn��|�q^-�őNf򀺥|�/	}g1�bS#9���vA1]�"�%ަ	���g�¶,�ԀێZ��N�
�N��z�߭������ӏP���˒,��|�4/����O�� vߏj��w8�U��H>�νb����VO��85naY����|����VJD��p�B]@.S0pN�N*���5�v�f[��gU����_�/���?ud�?�����sPTH�)G�2�@T!��P����C�|����z���F��Ag��zXH;�c-0Av&�8�sW��S����:s2��q8��/��#��D�I����p��~�㖙$V�7�����T�8�V��6z�;��)Rd�����IҎ����Y�X�����	n�� K��j�_�Ҳ�����,ԴH;�I,(V��h�L�}&���/�U��^`�B����!���q>�m��F��Ʋ��C@�'���BǶ0,�����q���|��>zFr�������L0��B9A&�&>�	��>2e��oԥP��\�+K8��Lc^6�c�%0���Y\t|G��W��+Sy�~��b�KUC�u�LoX��� N+<#i�}���@M�^U����ڣ(;�}�s$ n?�"���G!�H��K�e��U�Σ��lb.�]~I]�����Ŏ���\��q�q��S
S�J��3�|�C�W�����7�!�w�G��@t;oj��-Q�	��V/��i�4 _��%�Kq����@n��y��źXv|��.}G���b������	T���<#�~��m8�.�2�uO�,�j�����wꒈ7>�J� W�}o5FIomӂ���Bօ�خ�60\<��&P^lֽOR!�%������Hm �퓈s�j�D)�X
D��?;�ע: *���L-�36hR�a�K	9���=�6*2E�̕RH��a,�i�r޺���Z�E��һ�M���S[���ˡ?zaa�I+E�W�	H�Cpr>�s�:�U��V\��iϯ���h�`n�,Չ��0Tr��7B��o^C:�=����&�ۧ����n8:F6[M�Q�|흛���C�=y0؉G�=%����{\�No�0;K-.&��@Eͩ��j �\AM�In��o��o�:.����&h�^�I�u��0�/�?��l-���T������t����,���#��`W��� ���m�2����cN]�=�|�5���?1��hSm��������n=�ma���8�&t��A�+#C����������ij����U���p�$��J4��jKjxVT�X��C����͋~����b0��sLz��I��o����CQ�`�՜9��
���C�ۙ��Kb��u�o��,�լ?]@�h�"!4}U��Oc	K��b͏���Zk�d�r���R?L���]46@v�y��ɹn[�������5є�;���|)�AO4Y��Mgz�#�W4T�'��mR`�7��4���L�v�G0s<���3L�n���0���u�;x�I-�"M=���:��j��"F��#��x����=:g����w��-m�	��T�aa��������q�y�h=�D��v�0�_��P��������g���d�u��5��Ha�O!oV %��"�&-��j&�n�s�; Z����'�bI<"0UL�!C�W@}`)z;�x/�-�@��~W[O��`�qJq~4�}���I�TY�+��HmP�KZt&�~rW_KL���V=u�++�A����Z�����b��"�-[-�I%�t�z�$^BQ�����:t�׆�k��DPBk�T&Z2�3���{�F0)L`"VQ@�g��J?��؞7,��R|f_�s-I( L,�A���"g��C�r��,�Enh&���o�䜳!ݵ��=�N)�#�	ęwͲ�34 ?|τ�6k�[����k�&�Zy�w�M����wr�\� N>��N��$��ǚ�g�p�/9�/�ky=m��z)�r�"���M/g��:�jz�7������O�Q������i����Q��ϛ����g�d�v�ݳ:o0�D:I���T��A��u�J������G�������D��6�
ܗr���
g���+�&���I�ěq����6���0鍹�`
���B@#�V��\�W��%l����svl�D�%�,���4Ey��8�T�m�%(�˩��q2J[4>�;�h	^�>��Խ�����Mߖ�b��Ly�ϳg�yl$��C~y�|-��՞�}��hK��!�)�Q¶����֭�,1w�[Dֳ��s4��X���Ï�b�|zKdXnƔ�)n���:��F.�)-.{+x���R���j�֫��Ymhc����
Z�K��2@'I�c+^�A��Bȼ�?�dox��ӃZ��F�dI��
Y5/�	X���f��*�ZaU�s��/
���k��_vl�MWڼ�<�ϳ�u"�˦��"�� -�8��:LЮ?9?H��;�����ptٿR��R��|�۵4Em{�*S�7x���H\�W@S��6� ��"��J���2~WE}�^y������q���%m��9�h�D���f�]�s&�����:�x���QJ��3YsP��\�Gf�J��[�)ףA���RO��_��;>��bT�L���oʩ!��Q�,��ɚ���߀1O�Y��6N8���"�@��:5
�)n��%�����k'�)�����LhzuH9�^��Q2��a����EU���ܮZ�Q��S���z*D'^����( � �߮
�Y��
n;Afdd��bz�ీ-U�S+�XQn��}�]<B/2�
(��#�� �
��:�-�o�������G�k����*��a#������Z�%W�9����h%�_)4�X5���f^��5�b����]�+�gG��_NLe�DIׅ�˝��\la��j�:%yI0#�Z�ڀ	�@A���,�m+
�*��R�ˊ��k���,CDޛD����Y$���e<:�����FYoLoo�O!|ʪ/�v��:�g7�� �r,�]�T�A����3����dq���Zi���<��C5c�I��Ze5�|������JQ�Q\�n��*�ҫ�$I�Æ���G �*�H���_��f��2D`��ǣ�Og����ۄ��ٛ.��1��q�J�����vYh;7�l{"v�:���"-y�v^q�̨�S�RrU%���X�Q|��)8,�|�X7�"��,�����l�6�{��9�`��m"��Q~@�V��ʇ\zH�wK���\�,�=��Xy�V�x{�t��_f�G��\�ҿ���V�®���Ƈ�	�5yN%-�?��G	H^:W���#o��3����r��a�[�83�QiB��-�_��џ����K��-��0�}C �>&l\��"ڌ��v�#�YR١���O�Fm���
�xw���!7&F�8��:.W��L/YL������ԭAq>7�O�A<����|�Z7����ڽh��L���gT��_���T�ߨ�:��e3����`����+r�%I*�eTb�7͛� �!��YZ
��v��(��@I�2]�$�\f=o��9%���S����z؝���qR&5|�c�?�bߓ2�d_����c	���?�q�yh/?�N�/�c�3��(�E��H��S%\B�L��. D7ac����)#?,U�%ԫ7���5�;=�_P%pam�m��_�;�_�E.�mZs��Bֶ�*��ad��L���ȦP�}%[钠��Ȓ�7�ú��a�EX����5�e�zeQ�z̷%D�&�����P��OR�]{eJ덃�{�!_܏�J���S������k_�A��k��(�ͬ�X���
\;�� �ǴR�KD�D����`ouUFgD�J����W�2:}9P{6���v3&��u�E��`�G�����LZ����c]�'�`��A,S2cf�&�8��\k[�;�7wDa�L�QҪ�qtFL�K�������dM��F��=?��AM��9<7W鋚5�Ǡ��Ꝼ#��f}<��}qz~����� ��9��_Ü(_��
��fWU�+���G��n��.����)���y�����lBی�y���}7\iKCF��1rx,j���/>nVS�O�+#߸�R�@sm�-�]�+p�o6���u��f���O] /�Ɠ|v��<@	
�e\8�elEc��w�Yf��䀢̊�(S*��h�|�u��=oa&�S�-1��p���3�s���l�`��m�z�Q4�+S?W���r�y�*Y����`��p�E��i�*�� {�h<�N6!�A"��é��z��CT�י2h���0>�c��f�����B�|��Ts��g��֢��E��v�?kEZ͌���޲���A�t�XxB��h�)���Ԣ��J��G�;�yy��cq�(�x�<��0�@�*؋��*vp�G#�{�û�o���M#*N���u2���a9�.��ϚT��&),�#�.4�r���-�*&q�FQ6d��(�d7?CG�}zN7��= �N�t&=�M����@�YU$��>�żd��ک$ΘL�mI˥q��;�Cqzv�Q��m��6@�%�"��4nD��~�cǲ�,�T#?��5�(�엘���cQw��%������7���v/��`�Z������*N�4!�^$�M��r���S��s1a���Џ��`u�/���C!ls8(݃�.�9��f1���d��iRI�zR!��g��f�jcl���r<�C���ˠ=� E�
��bO�ϔb�w���g�*ol�2���&����HC6LL�=.e��Jz���Y���xִE��oX���j]ܑ��El�?4t,���;o� ��߭��4͠ٴ�g��iE���Ǭ	���C�L;���;mt�'��l�#۟�m����X.!��䫽�nȏx
9D˴�%�$s�F�D���-1Ń��;�TE{�@2�?��i7�#���a�_�E��G��b�bґ�iJA�8y:�Ixu���6VM;�4����7����jP��{J՗jy�W{@���4�qf"ߜDO~�r| ﯽ�_�e;��%�)$��~C�2��@���A�b�b�c�79}� (Bk� �Pܺ´A�`��y߆}s4��-}�y|s�
e�Z�V�|�v�r���DejX�=��7��nC�R�slb	�gF�s~=D��(T�Ҫ�U��_��AO���di�2�`�ƥY	��;�D�8�7����Ɵ���)>��)�óvro�Q��t[��ȁ���aVȬz����q�'(���O�m�s����^�
��_�#\�E�%��G�[Ց;��c�;j��1W�/.�w��/(������Z�&��.kK�ׯE�Y����YW�-ҫ8Ɽ�<�v�M�wU�ќد�P�q�[�����H�k) �v���U*+���3��^ef��>�o˘�d��pfV�*���h��q��\C��,�H_z�_�N�����=���,so�^,,9���W�o���2�������w���x�f�C�M���B-�^f�PR��>�b��= I4;hy��U� ��w&�~`�����rQ���4xk�4��*t�3��9�f��ĵ�ڛ������{�+&��e��F8�%R/�c�S.���7}'������}Ѓ��H���c��+�ݴe�Q����ionmm�8��d����]*�ֵ�sO�pb㡩V�P��TRK�\$T	*��ҝ�~�E^�MB�	zEg�,���l����X��[��vk�[]��+f���e�d�E��ʟ"-i�*a��	�ʈ���wd����"�\�=5�Դ����ui,�)y,�祡���L���4�ͭ)/޵���9����F�M���"��Y�ђ�&��Q�3l��tI�~7U���H|����m�A駬JBZ��l[!�t軂/�:��
�AWYt�4�.�3�ZH;�	���kt���<*yO,Q-Wt�ly%<��=��2���䎎	�g�+K�ٕ�/܁��k�=]ќlS2#���-�#�0�hM��a:8ޙ*��M����n7>hO��!�����>w�S,V�6�����Qj��<S[��˭5�Q4�U`�K�䓐��w�g��1*�,����a3�M��G����tj����kR�}ʍ��~�t2|5" D@�\�<���Dh��P�!8�Zv��᥉�G��o����i���r�Ü�f�A�5Љj-�a�x �Ucޏ���l7b���-��?��0.<����u��
p������vJQc�Pǔ�D�?>�6�|�?2�t�Vh]�������O����q�S(����v0���!���,S����m�:T�3������?��P�����%�D�ú%����r%�Qso�2�r�ͣuaL��`��<�ͦ[K��4�nr�@�dg����L�`�\�齃z�S�ێ�����܏�'S(<[�,`�P��j�es"�'*��0�N���8@�u'2�k�G �:��BM� jY����Tf�4(�%a%*��̣C�x��NS�
����dl�ɣ�p9�NP�_��l���xؕ���r��qR�?I��A������ftP��=t�d\S=^7w���_�����2�mj�G��8j՞�D��}�YG�P������P���H)_̼�U�No��lb��U�@ʋ�g �ts��5��s��ŶQJ^� �:�x��{����eEwf���)��=5�+ﰎ8�=�bqh�˻ ���7+�����Kd�SA��d@��t��s�-K���Z��5�]$��<�Ў�r�u��r�_,�`<,��O�(�=�~��Ь7�M�'*���PN�+{Z�3����p$ ��N��I�@ԩ��\����������bj {�BB&�Sf�*4'�vԐ��l���QW�&���{f�@�VG�SY$߸̓�DÝ�%��)\%��C���j���!X�b�ۧ;�?�]�η�y���jK�I>�\���c�v�Un���vj7&�H<m�S�I��s�<C��`��Qh&	�G��A�"�V�4�Ē�q�(�2�U��3�##�',�8�
����>w��9sf�G�hAL,�^Zt�������{J�Pdܰ�v����V6V��#SsTX���&^rA�M�>V+�ا	����fJ��"�^)br�-ρaԩԑV�U��% �H9���*�ư�}8��.��ڷ:�YZ ox����ӝ��k-��Y��2Rf5�.l�ծ�x:���٪d��VQ�B{���bb��t��(c%=��o}D$Ae�6��p���s׍�&������C	~����Y{l2��c�
�h��?���A+�'�`R��/��'���Z2�=&P엉4���-9��w��pT���yz�L�����Uf�.�GΣ�q`�m�̠�����^�Krל���n�	��լ�����~T,��lái=:��tvzn>�u��dD���g�j���a��*��r.������J �A��(a-~3r{�U~֜��>�T[���=9�b3��8�0�T�w�)��o9hhE��P��#ٕdcw~S�v>��l����(NHzFᧁYR�<�x\\ձ� �p���O櫶�#���a�	�$����4��Y��=�Q�@$��&;���#Ě��b<�Fhd���|����KQ�o�Z��c/"��?���Yr�;S��
� D+�#-�J �\���ě�[|�+�/����#�nki�}��;�W�t�&�%S�0%��d����Ib>��AL�E�o��oS2�럎����Dľ.71ԫ�h�:~��5^�i����	^��n2�|�!$�h!8X��u+dW�o�?�Pa!�>ꡗo�jN��5f�P*�YeY�i��Wh�_�	/���ͬ$�1���G���	��H��h!x)T.Z��ם��1f��xs���&����[م���xo� ׅ��}�?qܒg���п�w�+�9�0�M��0�V���tW�2��:�X��%��B��q�N��;U\o��%B�cv,,N#Ɓ
ɕʒEY*X_����*�'"6!�VG~�$�1��Q C|�uo4�(Z�H7k��@i�4��Yܸ��5�/>�f��'����P �-�I2%��e�(a���˦��S�Hq�Tp&C��㦫��S&����̫:q�[����L"��W�&OI��HEhNq�Ub��8����^߽��Hq)+J�*��H�oKl�>�(�lP&5Tnh��f4P�Uls��zȖ���1���A�>��u�]- �)d)Q&���4ɡ��1���l�O�Do���� H��_N��I���-��u������7�]�cO!"pA�i]z)?*�!��9�d=T	��0��_��GǓ���W3&B.c� �)�Q�,h���K�k�({ӳ/�f�x�!T"N<���;�I�����ݺ�g��tU�x,���}�[
�p��j���@�ɹ(��ᅦD����*�Zi�?�PM]|���|E"1;Q��e���} ����K{u�.��"\��,R��C���� �cVd�Ԉ\���"V���V�{�0���۶]/��ti�'����Tm5�Pd</�A�)�����DM����i,D����g�/�x���G�)�>��Kgn��H�GgW�*�����#�F�V�+Aڇ1��x��L�$
{]`�.,
��^�����!���?Ҷ������<��c"]��)�{�� ��HXU��gV��usES�z��V��=(�,yo���8'$ZW�e�Fӗ/W�H���6���S��,�1��迉��eg�~�9�A���{��#�VP1����X}d�m}x*B쾃GF������),�^�/��7j�\��!�YB�r�|�z�f�L�#���ǂ��*Lf���V"T��0�HB�ck������M\np�\=�_��AӾ��U���*wS�H�X�����-4�Qa�%=!a�o�V�8�u�/�w5��V'd*1z�ܿG'CL��"���y��D^I�h24 S�Zs�A�=HP�K� ��q�v�d��6�F�	~=)@�|5�c�:����*;�D���W@`u�ҏA,̼&ž9��C`����e���ݺ�PR�Z�תbW�Z\ӂϕid,=2�/��z��Ti�I�i�mU�G �b0$A,g��)�^�[v��O�j�=nR��j����q����p0!� ��h>�bZ�8	�T���ہQ�f��=���6�28������6��ܛ����M8�80l˝��Q�cb!0}��f���d1��yv�Z��7Ib����n|t�JaY�С ^�;���g��� ?w�h�K� �m��Q	���W�Ky������_�TGC���V��F�ma�Ԍ����2�h#�ʛ�K�$��/~7�I�'S|�=`�Y�B�w�	�־��Q���٢qe�X�Q�G��ݟI�]%lD��o5�����S'b�U�6�龩N<U؀12Cc(�_h��8���Z�u��}��Ӷ��2PwH���FJg�n���{b��#��F!����̔KX�
�v�2��4ٽ��Θ�-�v5��>͂����ã5ߡ#4�CvG?�D���68p �F)�o�e�a�?������Ɏ?p9i�Cn	�R��)��/���EV�2����C�������m	����3n�6発2��{ܠ�h�^��*���%?Hk���%���(�P������wm�-�_(��K��-/I�gȺρ����\���I AB&���� ��D+b�q}�����
)��K舜S�@Op�5�?�hÛh-�|��Z����k���y����=�E%��Y�q�j����O�K2��r����w����Uq�c!r�j��k�k���Y%pX����(��,�@��-ϖ�&qM4�s¹ܮ�R*1-��{gf>3�ys(w���z�_ʯ��	�y�qf=��\��?�ߖ|E�Q��OZs�����6���{3�4��z	�S9��B?F0s�X\aߘ����rv�JԈK?�o��x�g���;"�,"�~n��.���q�*��"MAQ�R���a[WNj���{L~r/�5w��G��fNU� ����H=$�>�HQ�3��-r�w�F�J��!Z�?��T�y,�5D�XB��B��-���0Df͊-����Fd�e��_��Moi��h1O����N��G?o�{���F�A�i,͔��`ą1��G��U��j�'��6i�MQ]�����{'�JƱ̲��\���@�03 ����,���T�[�["$�ޫ
���F�8��70��e��`;eg����6�}��4]d9i�p���Z�y׋^O�!֧e�]T��������$J�������Ul8�	�ˤ`c7NP�QF�2���w��E�}���q����>�.Q1�1�ƻ��);#���UtD�!�>њ�&�I�4�g�x�
��fe��GC&�ȍnb*
u�T�\�fXw�섘^CI���E'�,:�~�7Dkõ�;��u�|&�Fw�2!���d{A� ��z���Xg?�;Z�@�R��
L��P?�A�/g�-��A�nleW�c:w�l K��߃i��}�@+�Mp�������t�CӯG^߃oѥ��*z)����{;
�C��ل�97%��P��h��4�]��C��b�^{t.��!u�y�J͛� �<�ePEN.�I�,����Mh�	�ۚ4�FR� �֫���.�����3B�� �A�����_$� Z[��,F�G�z{b�!g" ���2�-pƼ�2}��;OC���u�J0�%?��+�U<-���Փ1�������h@]4*�D��F�74Ι�4� �Aq�6蠪mt��ڪ�:�`�-ͣ���L�l�2��-��G*�u�U�E��p�h78��	m�;� �-x���w}�	��w�g�D]uwݢ6;(z]/:sl�B(��4�X�N	�Ds?�\�@���\���<�Y"�����;�bXvΰ����ٶ�s�RO��|v���{��-�Տ�fN�\fr>��X��">�b�<�)�� ���{ɨ�����V�ŜN�0��0�\d�	��^#5� �XYa���,qr}��9��_)zB(L�ȗ|V�J�ί�� ��~x��+�h�۸8|���0 ��F�7G����ل����>_����lij��MZ$��ڲ�qgOS@ͱا�L��2N�c��΋jVCF��__/	��`i��A~c
�O� �$��.���˹�?[���᡻&�7Y��x���9岶��O���c(^U��3W�C��[H��(�����K�y���s�aK*r���NC����k@i{��Q4�K�h����d*P^8��K*z����/aX��{j,���^%��9�j3��O��2�
�T��k�E�E�V�#Img� n�40+����%ت�^Gr��ĵ���C9S�g|9�T��^�r1�6ܲ\?�iq�������؜>�0am���is/���}���p�Ҳ;޻�ʜg(��K�Z���m��lcM�%�Xq@��n�읿�(7QV�sfT�+Q�
K���G9���T�h��%�ri�^�����c�����l��� e�K,����J� +K��>�\�]���oh�w5�ɰ)�EY�#���a�\J+ cp�oN��N����21�rdZ���ۯ~|���u��oI���b�7<���e����xɾ��.��@�+,�g"JG.<T�m�2�i��o?�<�����G1Κ��c9����g�VL��^i"ʉ>�i� �ϱ��T�!$�3�6_ t�f���A�^����V��T�����'�68�`�逊+�� ×'��m�5\�h���+��^g���G��{,B�R�gi�>�t���@�2ֆd��Y"-���1"6Nfi��N�}b�0���1m=Hc�	P?�^D��[FPؕ��/��4\��a���uķ,�Md7G�7s�@�X�n3L�d<�c2z8��䟳~�~��[�P��\�7����1m�;dFtYGA�ϴ�]��R��������t��!3w.�Kl�&
�˼P%E|bZ|ts00ђ�V
�l���J�Z�oum��a⿺��m���M'ʪ��A~W_s�m����0���G�c��l�˄�P��Ď�ܿ�z��9Iw�VW���H��˴��~F��Y���7	�#T�逦�_�\ɑ;��W������~"Od��a�"Wx��l��f4`�g�q�ԴU��j_��_A��Wy�3����2(ߨC"t�h��N�������4���TЗ���J������{g�G�h\�	b�梢�
9�7��t[���מ���b���xx�(�[5�z
����^�����)TB�7Tɀ&;S��
B�
����UJ���`?b����`�����F @k��7�X��t�V��5�9-ҪwZB�<*Z�澾����޷�&h(8�6󳭬�{p�D�&���)��{�S�|��Ԃ�B�+����a���1�ʮ�z�	�e�r'Mh���^����*+o{�ѳ����: �a����:�I1x���_���<_D�r%����Ν�,xPRi-g��DЯ{�~�ڨ�f��9L��T���s1J��ThޑO�)��ٓA�\�	�c�֔�����S�ʕ�L��K�RtD����)���/��yl��B�O:{�	�(/�%w'��O}K�kD,������F��FK��P*z�����̃�z��="��a�"o`�AkNL	yt�d^R�$�[�bo�)}A2�c$,����]�I��jA8]� p�hnꜲ�8����5p�;ޝ$���-O83\Gh�T)���(:�ȗ�������PBoT����E�d����_m��:��K3�̬�V�LyK�x3�	[K��~����i���F�^Nn�5==+9
�}�08�B���p_��0�!���E*��W\��8�E�Bہ|�0u�3�n��_��f�W�޴����N~M?�W�>�>���RL�B���Ld��n�2�T?���!W�x����_F�����h'�F�xƱ�XwI>�Ӓ��F� e�(��U:�_|�(�)V�����F�?��'b�\f�^���ز���OT�bV.���U�������Q��o/��D���ح�,b[�����4G���g���bd��Q幀EaK��������@M��	��u�x+gՄ��W�@�s8�Vފ�c��;2?�s�<X=�Va�KQ5Nm��`�ܑ�	�?=I�&ʋ�k�d����&�s[�8P}O]� �݀�V��
�ݑ�w;�:dMSMiR��A6�|�ia ���#����4Dc�#�m�O�g����'Q?�����%��R��J^(�)�fm,e���;Y�@�-�	_�Ӄ?�4�,�/�ۿg�����7T	^�+YF��#�#݂ӯ�p0�����ߊ�3]h�(�_B�BXS�F���TOz>�L�>����!D��u�<�:	�yI����y 3�ܟ��@P�s�S���1�D�p�K��?���,@��zv�{��rc����1x?�M��Eױ$�Ǹ.أ�/+�Ț4�hG�W��νlz�R3vT�ݑ���j������ �Z��-�7�Q,��X���P6�8����G�� o/
�=�F�Ds�^X�U���S_�l9V�Q��+�,6@�1!�o^��6��L��7x_��]����v�g��0��7��|�9�YrO|�3�:+0j~0�ǜ�9�okbu�2\$���n�yD ��<l(����qX
���	tʰ��?��=K�㭑��&��Y�Iā9����i�25�ʆ�<��,��Ki����<gR�_%���2�I6C��N�����iz���N�G��EM���ogx�Ҽ�6/��<"z���L�(ܗ
3^-�,#�B����	�@1��F1��Xb�Z�ty!OȽW�"^�1����]a�9�c�n)8�꩚����9��5Ut�זS��6Ӭ,�M��U�3���}w>��wgqV� �lΆ���L�q-	��%��� �T�ƾ������a�M�H��_9���6yk��. ���q����yDE_kD(
���,����=�|F���S������Iɒϰz�SXoa����D�l)����y�,%[A��$���Uj�RGX���1�P�Osg����Ds,�	��4�,1d�=��ӵL�V��UUv8���s��Z"����?3	�n⯪��&
pf�)�X���6xVDR��J	QɎ�oI��X''zb��JUn�NY^t�7$2��܋4Z��9��~�-o ˭�'c���!�ULq[�4�	[�n[q�Y���]߱&d��d���1�o·;�[i���j'�k��J %Ť�����L;F����*��MY�^Ȗ��3وö(�F�T�d�U�J�i�+�q�c��µI��y�0��[�m�!�P����F6��m���'�uB�֟���ְ��CaG��§_�Ⱦ�ޛg��ϕ�|D;�/�x46��T�����*�Rw�
UL���]>�[�U��l�E���If߻�j\��4{[�!g�{���!��R�v�26M!�e�@�;��k�Nqhՠ�7�2��;u�6S��[1�ׇ��m	7A�; ��:���p@VH��n��#_v�8{����� ���F�%�r��5;F�t���f�Cmu����0�я����g�O4Ҥ�_mV�0��O�*��L{��j�H��H��al�4�\v,$w*�>�ݵ\O�O�����]�7|�1��9��7��a �������c�0������Q8,t�2��?��1��Z��f���/,�<�J��`L�
�E��(��$�C��0�9�MQ�(�P��}���u�Kh�	v��uE�]3v1P�jI�"稟]F�HUҠ�D�=-�4ϧè~qjz�����9�� ���
d$ʗ5������a�lzK~Vd��u���DEoɽ48�f�w�J��
> �B������w���l�]�"�E��<��3~!�M�<�fU(Y�↽��-���+!d��y�Sͩ~��q��`���#Q��o��%)�����C�k�^ѡM$�hG�!N=H���OZ�KÝhk=��$�pu�������>0Q�FO��e?y󘿑�����(Rv狨����XTV���"�ny�I ]ƚ��Z���m�7(�h�w'ޕӪ���V]�����>��]�>�l�2y�X����+쩬��>vc��H
m��ٖ�`���KWsy��&��}��2я��:SYX�ahJ��@�S��NHS��2E.;��\V4�df�D��
ƕ%{

���� $:}f�3����O&�s�����~�=c5���� �2��;������<��F�k�@
B�y�;=v^r�;����JeP�ݹGz�y�'\��S7�T���w^Rs�5^ç�		c��fx*i������,�䈰y4]����w��\�'<������� ��7��W�_����V�M�#տwj[z��)��a|��<�j���W�7k�G��ho�u�4�<��8?�$�`����ȱ�.�Κ4#6������R��dQ/>U�����T�.���_>SՌB2[�_?��+� �2�����~L��w� ^A�*K������w��@��)a���Sa����{Ւ�2VhZ���&<))<��@� ���r���h�A2\���@��Z%�i����@1��KAt?M_�׉� ��%��O�Hz�ّ@��OR{�K��jU,\+� �ڏfz���@XOo�C�귍
N�����~�m�f�q��?l��C1�Y�uX�����=g:��@a���0�Η�;��^U�ɹMC�7C�?,��2h,3H� ��C�>/�|p؜�'"��J���"���'�|h�|�%F}�uK��tcbl�����$I3:Ds/MpX�"<}��	MKĒJ��|��{�i�l(Փ6)�ZIv�qB6ai�;�j�%%_}�����t����5�����a�%�H-�t6[o�1��?�K[0�.��)��rX�b�?�Bf�9�3� ��"#Q�Qv�l���?��1^@�pq�g����i����&ʎ���a� w�m4�:���`�zo�.�yO�"�$뾧����:i�Qhj��Eg�v?��
��f�C�JV�V
��r���N��V O�`��+l�4	�#����DX�f�h�1�XQu��]"�s9�L����!٘U��H��=��{�}���2�¶BI�,���ٻ�%�ul]���'�kY���� �6�E��:��o(C�7O}�vW:#넖��"�IP�_��h�9S$�D��Qm��?Ɗ��;V{�󔝢+��|Qo��%Q ��8K�����\�	&vQ@��g�������m[�967ʁȐ�HzמɻJL��?as197�6�U���E�]��l1S��٢��:��>��(f�����+�̈�mZ�m��%�amnU6Z�Z���y��H�7F���������/�d�t!��i�U�q&E6��A���VevT�b�?d.��2�F:��_:2��TL�7��]�I�lh �#֮���_`  5ާ �~jۙ�@�(C�R�+$��x\Ig��Ra�php����Md�(:��T��RX�j�����Π�~�Ր���e�v� g{� +�gK���r��6���t�a2�N&$"���>�����+��{ޭ�7��̀u��+���[n�B%rD�ԫ��B�/@{���*-q�?����1�ȭ_LK5�%8}��	I`2�2(��;�)�=�΢kc��yׁ0vb��vW��p>�.>L�s������+�Y�rw��A����1!K\��-�G� %J[8Zۆ�,#uG�c�\m���WwNm��b��\�f:l�)��Sf��{�ك��P�p�1�1�]K�kMw���䱍("zJ��z5>�*��K_pސJ��W���ʻ��إ�+��3�;UД91��9m�%K�*��ѩZ+�����Yu�@�,`�b����9c�s:M�l �����m�9e �<�=��^y��KU�3?φ#��:fd�)�͗����澜����J�AP�FC��q�N����qǢr��U�mS�M�]L��q/�3b��S�6�s����� �����8,�1m:Qf�.�O����[�BDv�j����<e���a;���ކ�d�EɎ~�=���E�(�ĭGDG���� Y53ŧ���e i�����궒"�i��I�T���Xnh+!jch��s�G:[��b��³�H�PhpW�Fs\σ|4�(&�|@Nw���/�J�>�`T4Yߛ+�%���T�50��C����Ϫ5�3�Ey ���[�
���N��	�W=hBM�y�S�F ��p����u�%8����k�^"�7~������1�@�\?�G1�w�,b�]��%?V�v}�#�Y/ŉwgE�'+�q��%貲V�]�q��K;�s�G _����o50�z��\e.pg�G�e#Ț�P�d��Տ�}n]᲍+&�O9#�~��0(�>�ڨ��x�v���I]��.};�r���GT	D�hR�I�`Э�h�E3�w_�|���i/xg�,'�_е��8[��(yr�z�J��q�+^wU<C�UB�?7�B}��"��إ��TE?b�0���qc���u���t�𫾋TS�;��;3[�y�T�(ˢ����3���4Q�����M�Ҹ��C�T5�gܜ��9�8�7x�ak�3�2��t,r�|_�4ʄi�H���+�A���gc캌��U�r��*��S���'a�R��C�P�@��	�D���H�Įx�z��5�k���yhKM��z���H/L��-s�{�UL�	���[v|2�:k�m`���q�!ƅTdssPũX��i��d�绗�z�8O���Y��y�9��&�>O_w�*������dV�����9��h����@�(��q��YB�M2!�^������F"�K|��;�m_��Lb`���l�abIHSN}�(�rw��BZ������Q����Y��9w�jսrݻ�@�[@?�.�^J�P��@/$���UE�Gx�eo�.jR���z��:�4�@1:q�,�}}Mf J_�u�*M�ȵ�`i��hU�?�j-�f9i`˦$�_>]X'�� zs�O���G��~�7�Q���`��{C�N ᪍.��X˸��E�9��P���w_w�V���L�w�]���"�B��mŀU��J���a5"�a�6�����v��	a'��%��S���Sg�� �X�W�DM4�$�oh#�����i̥�Fbo�Z�.�E�<���T	 j�e8/�D_�f��sr�lR_`.��_��oc>�����nֿ��-��,������z�LT�ӧ��r�i/2�N��{���O5%Մ{HL�O��xΞ;_L��(DB��h���&�-N4�=�6�2Y��s�e˪��I��/��()9�m�L��{��ݘ1~Á@��$���j��w��8�r��-�$����@^�W��܂��$���L5]X��Y6�(ҙ�CL�$_�˰�ځלˋf~k)�q0E$�e�a��#-`��z8�L������C���$߂�ʩG�/��B`:��d:�}~��hKp���V[�n���f8wE*��m���k����
����"�%�'���3�:NW����n"�MP���[yU������N�=�y��z��3�V��f��H�ܔ�&�W�;�
8��y��x��<p��n��M1�f�R;(�4GV���v�R'"�Nty2�JC}�0�Ε��*��FD\�Kc�e �����y���vu=/���n( �Z�ߞ�1)�p�dr��GD�x�C��&��*,�����Y���Ky��SgT�I�_^���nd��/�S���e�D��{��G�����$aD	�bE��P/,F::��8D�g��\����	N�c��_��\R����&�+c-��ڕ�+[ \X�T�{�0S$�6�)��ݓe�+]e�g8'��fP�Kt��5z�k
q�%Ҁ�PK�=�'np�O1u�r��I�e�n傷���{���{qsȦ�?H�^�#�xR��b��#b�cm���09	m~��A`��Â�6������h���D�n&؆��woWWVP5� Xm�؍���hE�9�.��<&����2�${3d
�?G+��	m�� ���X~r�f6����@�"ۢ��ᐹ�ۡ��!��,��Q*Z�kβL%���8�´o^խb��>}�����7�1�"����#_����u+�=�Bb���C
c�?<���~-���D��P�26��?x�)�"���R���n��"�3`�)�������ƺ��W��<�~MFHY�GZI��{��D�r���Y�K��g���m�I�9mY��}R��8��#��E�8	O�-�xRcU9
1�"�^�Ӓ5�n$N>ŷ�4�^v����e�u���Y�<NW�	)A%�B��%
��p*��u��N�G:��d3tг�Fk^'*�7��G*��Ѩ�6��h��vJ�w�\�������� �C��T�ɩ��;��1Q�;��g?�z�5�}�Zڕ��y"�x�o���}��i%�2�$VgxY�V��	U
�UW�Pi��?��+U��=�.�4��Ap���4��p���,Pٹ/"��\��{Ʉz���aN�ӂ&���5u�#�Q�WEc��ʿ\3�m(���b�2�EoR��Rg�7,���y}b�fdろW��$&��^��fG���'���B���1���4ϭ�wk�wϽd�K�k�0�`|B�p���^���4�:���r�t����y(L-X��l��>W7U���;�oP�f��6A�1��YjLs@>��T�O��#��§C�d
�,c@�
) # �?#�{�A�\�b\\̭��G<׫ǁ��M����}ș�� �w��r� ����'k4��:$���/���ޜ�c�B�w�M(��:X	HX�=�p4C���)v����G�1KA��|�� %�Y�g�}kqu�Q��׆���};��*�ag��8Z:�^�`��<����La�'Tx__R��qQ���#qC,� �'0���g�����R�׹��^5bx�>�h����L��[��c�;R���E۔9سv	`T�=��iK�Ϛߊ��� -�1{����I�}I���OޜOR����3 �{R�#i �E+�q���v�St�:p<
+M,�x�o�����U��sj��9��H�Y����\O{#���38[<�y���:#���X �S<��;᭜�e�:��Vd�g	�<���3
�]d1�cr��HaRg�0ݫ�)����ٗ_f�|�T����bG���d�ˁ��{�j+��n��+��@<y��X%�&½����t�f֥�"+���7i3�s�`���
*�^�1~���^a�_AǺ
J>N ����q��t�̾�$Sv(�݅�J�XJl�|�EA��µ�Mim�L��	&���k��n�Y�y���æC-���h���-e��[j)g��̛�������]_��,����ف�ί9��
���O	���W'U|���P���ODP`��d��8���P�
%����n��`�[����J�t��>���Ηi��kc��?dƚF����ЮLZ"������Ŷ ���A��r��V)Y��Y;F��G�1��1����hC���'4�!A F1
�m���0�Ρ/��g��0!��[�����}
+#�83̥L����f��D��N�k��T�Y�Eɳ�Z�{̎+j����do��l�Gգ�,��=< D*ҵY�ِ�X��K�5�J�͝�����4�N���C�[�Ű7�UQ�*0���H�kX���A}|��T���v���פ�w2_�Aݙ��V�z�<I�b�<A��n��v���Y-+��E8$�ރ�������S�v�A/�C9E�a�I���Á�2��lR����iQM���PK��(��.�*a��ʾH���~^�'0�X�<G=�$>� MaSL|;ժ�g���?(t�@/����Y�6V��t�לTRY����ћ�慬9��"���cQ�����tA�#e'��]�Ιlݠ����5���F�����4��|�#��}$�׃6��������_��ڳO�T�������G%/� h!�Ƈv�,?��mFs:�Xm�-&X��F>u,	\+v#?<��o��Q�h��ފ��6����Ík�4 G
i�3���8��'E��w."w��zz�SZ�ѿ?n�I��X��1v��:	M��P�� H��*�5�֝��>k3�u�nb�M��y���`Ba{��a�ϳg���f�@:�3�_O�'��%�@)4H�[�(�?O(4�o�S:���5<kK��HKyPF�WH¼��e %���j>)"X�v�����m]كu��3��"k�5k��v��̄+Z��5�.n�]ɛwsjQ��h��=P��}~�i%��Cԛ�夈a��k�~'�!v��O�Ua5d���,�^��l�\{�2���V�����0s7i/ ����ft)�� ~Rv�����Z?�ݗ�n�W� �H;3R"�ue����ᆙ��+fc:����#��O'��/o����X`U}�9���`^�؅]��\i�
�{46G��-�}~��˞���)-����->5����(�ф7H���C�#��n���NT:z��N�F?,)�P&�/dSI�~aYc��ն�~ˍƷ�Cω���u�V����ZS�l�J���NM&���wU��>���+mXq�
'���h4_����S�{_9�(^�2G���nɱ�T�^i��+���R�Лˀ�[��'U=���CG$`[kV���o��v����m��ZQ�q!-�I+�REU0��*��ʃ�U6K�����I����#�b��tM�[9Z}x�#`D�Q�=1�GK���	�9ʸ����gz���Xm��g�z����)LM����/�M"��`av\>����W��}v5=�=K��V��5��b5�T�},k�x'��f�AȏA�F�2�I�Wm�������ֶp}᭪΃엝O q������Ӟ���N���g�^�V�l�qx�f��5��~�]�3!q�mO!��!5�E1�܆.:��鯺<��8��d`_S�e� ��|�콜o�M6Y��=��g�ܗ"��/E��lJyo�C ��N���n^OΦhط-��]wLx v���&�1P_��rK�r�uxE&<�YP�������F���	��z4��6M�M��g���) �م�n�����2�0ӫ�k�*sa�!lR��e�p����c�{,�!?���j��������r<���u�����E���G8]/�&���+�lP�7/��ԑP���k,�v�0f�рҟ��������ϡEh-�Ռ#Ϻ�٧���p�F��n3D�t���ٺ+�c�:4~{o�
��@���H��u���6i!WJ� �T�K���¿�OR�%��������� !�Rf?ja+Apn�Ѻ�eԃ���M�M�F=�k�՚�B[(���6#��SO�=�}.ð�DVHTׇf�K*�F����$-���[�we�����D�NH^s�7A��9��q~2n�u�\B��#bO��ke'�Z�o��t������2�!,j����t���<��B�٭�׻us�V�.�������g������������t;�O������s	|��MV5ئ	9g�ˠƎ'�&�D芞tC�f'����+��PQ<�{ɛ�V��O��!kH���b���̓>so��uȒa��C���ze��>Mxb��!�v8���d�g�g/�5�V�kC�h��� ����nS���W��O�\����_��́���G{/��^vL����=�ǃ���f�uR�#-e����qfw��5`aB����1C�i�� ��MZ���_zt�DObۍ��9^\0��$�4>�&�E�c��Z�V�D��IJ��3+��_w$+�J�M���� ��n�c|s\Z�fP:6��3�����R�bIjT��R�����6e�&�P_����\��yY �t���qC��,+1��Ok�������K�'��h�x`e0U!Stך�5�Jz�� ��� �VҠ\��Mz��VÌZ���
�!b��\����ڠ�:	I��U��C_��V}Q�5x���+���ǤX�]��B��F��!�a�!����!�f���(M@�\���ѩ�Y�'�L�IĔ�,U�<��Ri�۪4do�y��8G_uPg; ��� )8�PC'^n���d
�|x�Z��2!8�q۠��۪t$Ћ��AKy�d��+�}m_K���%����� z��.��Jߥ�X�K�Ĩ`d�}D)\�힚b�\�Ұ�.����bg�v\�E�1C�c�4U��`��9��7*�9r���O؟�a���)N7���y�x�Ȣ�����6X�*�4��f�X�F�EOp�7���yY	����yɒ��_�Mz�ej\��ݧ:p�qb}bu��~yTS�	��n�kZ���ك,��mx�Wbu��� �S�5����*@�p��������?Ѓ��
�R�"��E�a�������H.��l�43ƙ%�(A	:Y6_�1#� 9�� M*����f���w���?���ژҢx�)}�����K,T
�d<֍��@\�P���mmP��vI��_���T���B���1$Ȅ��d��QU��?u���� �JC�^�/��dc����ŏ�-{qi�K2b~e�h�@9jr���Բ��"��������k��5�h�����RX=Åu:��gB�6"2��ȨI ���@�t��C{�!�%��{'���.��3���AtX���m"���LтAۢ7J�i�9�����ʻ������p]*:H�\,��Y���Aۨ�DώT�V�Q�J��<�K��>���J��sQگ�T��&������CKVp�⃻����TE�E�݊�Q%?��)��b����9�1�*�M!�e0��� �Mr���
�sD^�tȗ����4;N����J�N��n6/������/�L��;�{��1�E���Q;�y I���>��hNo-1�����oG�"�_U�}͒c�u�@<&�i�eZ��*D��u��c�.��b\��rgx�!,���>��C�A���o�cY��<l�����ǲ�{ġD�����O�gءc�&`Ƥ�>N�ۗ}ۋ�?8�D`��ǕO�K�'f��|�&�Su$�e q)�W2�cQ��p��M�w��U\p�����8\zԛu<�~���ĲK;6�0;\�����F��G�j'd�i�||v ��Z;6mt���Β��QLo�h��R��|qf�fl��1sH$V��(>�C;��5� "P -HFa�#X�9?��[I�$�.E�6�Eu��"&s��B�0��5���i��Â����m��ae���psoP�.�����(1E� s�v�[�}��Պ��t�Aȑ�+S���a�����;��=���j�F�GA������d�F�r�����?�U���҃<� H3_x�e�r�s�^I�P�}66��t�i����L(���$�L�4������X��kYtK��(ʌ�)i.���m���M2�'OԄVRP���
�Hy`ꕖ<������R�7���#<�<�|�hq�$�I�Ș�oH�`��n�Z�'�h�f�T<�tj'���Zs�BΞE��^�����G�֐(d�� vC�u��l\BB��d���� ��{��V�6�;帶V��=p49[���T��X��>��embNG���r��t�B'f�^�,MhH��ر��)�Q��Hّ�7̸�U��V̠�������X�u�|6��X��=&���*��Y��`��\q�g�8���2��k�p�m��;�]J��4ѮKP�N9k�ͱ��	:���u�S��b��0��R!�Y�������l
MEw�:���G>�+vuVO�T�U�'���H��(��S�Zpm�g�
���%�ɮK$��F ��3H{��R���~�R*�;�"�<j��*q����||O�S�����'W��ysh���I�.i�@(\��3��ge b��fJ�и-�!�5���D��0��2�@w��t���O�`��ﱘ�$G�o'�T 	��?�%pz_�מZ�2���ua�}�(��������"����<g��f���P^��,ç�,�q��Zgy��U��Ǔ �sk��ɉt΂7�����i���3^a$WF_/���Ω�����ǢyRb(&�@�:	<[yQ� L�$wB��n���dcd���p_�����픋��=9p+�U�БR��u�俁�G�`ݠ���9�V�n5
R*��˓�����{c,+�N��b�8N�Ȥ� xI��٨����?�$:ߨ'�A�Ij �U��F�}�汝�H���b��dq����� ����|[�h�=���k�o����b,4�rLU��gPq�#�i�u�Ͳ��ڕ_P��=_��嶷�H�Z������k1���P��`�!�l�{����kh�i',5�W<P'L�g����������N��k{��9�(�9Э����\ݺ���![9���<T�4�����;���BS����?v.����d)�X""�~��M�XI_���)���[q��E�fDs�5����l.�_�9 �BA�Tiu�Ϣl!���9��ƣ�6��
����yZR�o߰��o=j}W�N�^��J��i�6l)e��%tV���͝,��N@���ӆ���7	�U��ј.E�����2cF��ҧ��[+푣?�"*m��jS�숹om3��8yY��%O���=�S��(Eiha4w|�_�6��,�ӯ�5��1>�g�/E�q,I!j������Nd�C�բ�@�������Y\�1^���	�C��՚��gf���/s5�������<�7ӣE壩�^_8l�����m�X1���,�	��tJ�?��0��a���+����Jb������ �C�(-�"��p�<J���S�dog	�N5�Nn�NZ��2��I��oZ���!hOY��ֵ@��GIA6�i�-�=���]�1���g씘-���<2@�tB��H���oP���O�Y�,����\\-�
��
G뮠���(.#u.��[m❋�,�К����3��al���­?�FEYKOdL=�w��USh���̣a\��P�1�����t��f8"�ˡ�[b�l�oL6u��Q�U"��4��yrc�u���*�;f!*���s�h�1��gH|T��@
2B��7=q���12E�Q�sk���������r���u	�_vep��O�	��^���?=\�Y']��{i��#�b����{�o{��
W` �I���ޠn����&(���.�X[��Y��T���u�UI�lW���˻d��I��1!�A	93p~J��b[���F�A����b����W��V����Ow� R?zZ����ߺ]
�$�R�s.�&c�}@M^4�?������<Mb�@�߉�b�|���]�x����a����@��OC����Q�.�0��u�e�:Fy�Zs����X�Cy�o�G��.�7������.�՜�%��:�˷p��O��Z^r���u��"/�[���-�6�s��SY����j��~����)�Fby�/O���7l����4����A�����ݸ�<S_I�9K�
�x� ��ܠ&H��8]L k��խa��}���8�W%����7*Qy�Rd��Gc{�4e�&��+�\�h$�A	z�����.,�%p����{0VwTbbY���1j
�+�n��/�(�P2�9zaL[J7�/K0嵧��$���ˁ�������o���l�	u˓#�5�j��S�����ZW@���y�X4�hSi�˥�c��g+A1C�Y��H�p��T*��� �=u#��\��,R����([_q�M�RMz�4WCἄ�b�����lH$��hc�t?���bdF3t��fdT�.H���8����b�w�<_�� �B�v��C?���M�bq	��ۄ�DT�@?'��C�	ML��pJ�9�p���M9��BzȼXw��ݶ���zVn.*���W��P �W������F>Z~���΄k�c�݅���i�qW�|�������n/�nֳf*(2Qt�+z��^����n �f�+n��pg"���=�
���aKF�R�h�H<N�����z2w�| 3���_<�`1K�FOlw��]�uŷs<^nKo@ȋr��cR���ǢZWLR8fUMi~�XġI���^�%���^�r^�����k�p��J��B\p��mHkgE/��'p�T-�_�����~�.�'�R�$�L3�f��y�*�"������ŭ���|3����7s.*�u��*> ��/­�v��Ϣ�|۶i���s~H���j�|,��䓃���=��^��p[w�|el��{��'��WZ
;�Ϡ;�5�o��Ǽ�!��5�.V�\�5�&�^K?lm4����,I�\�N}�I���Rl�:�
�v���y�ݧ-� ��<�>���w}�H���k�q��� �Y�Q����_.n_��$��#߻z�5��86�.�?���3b�[eNB=2�h�+D[�=+*r�g&j6�<��m��D�� ���������|�l(;ZG�x ��&�� U�z�ו��6Hk�O��M�RE[��X�L�q���-M�,��~�b�+�P�aE���;�0����w�����ҭI|!-÷�� D7Aފ��ի�2��B�a+�U����2�eJ�9i�o |��Վ�A�g�TP���S҄p�Ʉ�M���r9^�1i��%F�p5'�R����C)�y�;�|�B[���PwU.De�q�������d��%UE��V�H&chb��o%63��J��:9����r��t�FS�N�-Y�"F�_K��	�e{0�c򇞺ղ~)��>���Ԃ�(Zy�p�c|����I�kk��h�c�O�{�Q�>ߵG���棈/�C�} ��o�O�h���s�D���SO�u����Xt�ཥ�7h?q�1�wF�D��X} �Z̿���Ȋ�F%~��y*���&��~Xн_3�e�fM����Vg��/�ѩ���
�*���|*k�;H�`����5�8'mܸ �w���U����7)7O��c�0��a�p�|R�#E-�S���עR3+4��]��^�M�Y�n`������Qx�M��f�.rh�E�^��ykF�I��e��::
LW:�cUj���U-�#2��H� Tܘ4�_�8"WM>�����U�`.�Z��5�&\r�[�
ׁ�3����`o�P����Xǌċ���$I���g~��O	`;��u!�����dR�e�I�*ZM}nD?N��ɢ�t���ب>(*��%Q��)>��AE�3��/��]�T���Q�6މz7$dZt�{|�Uy��i�C���}}#�i��ɓ+�Z�@F�Ò�vE��Qά�Z�8����n$yZO:�<&��E3t��	rm�l��Ԍ	�(MN�p��ʨ��лA�8�}�u�5ok��i!+Ɔ�J~7�5��x֬�ƒ���Ö)}�1ńc�k��2�1*zU+�$��� �H�Z<Щ��?�E�����
��D=������ҙ�����ǜ8�==v|��þ�ӣ����"8��-���U���(��Eh���KF��-��ߑgީd��s��L�{J%�y�
dⵅ?.Qe�ݙ�|�M;�ʲ�@,H�>�ػ_�ht���#u��;ɍ��v0̑-dÜ�j�N6f�dUh7y:v֙t�1�B!U ����[��gNzC��b�}b�'H
n��� ��*	�є1��C�}a�oz	��Y��$L�4F* #V_Gҥq�)��s�"�$�3#��ƣږ���{2u��G^�6Jy�Q��xFES}�����K�s��LBZ���D���4~���{ﰧ��
UMErt�J 4c6Y`�!S���5�!�瀿r�"8�����&�m�%'�-���v��� (��� �&�`Q��������3|y����k�8�����	�
.���)@���:0���U��=�]���7�G#�jc��$հ}��Mon+��`m��'�E�kK��I��H�$��7ݲ�)�~�֥;��|��)t�]0
�]��u3��7����$�hI��.y��m��	[�����L�a B�4}�I�겞P_�aQ�K����`=i�����O��)���nk�g#I��IWCe����Ơ�Av�y¼>�O��*�ŧ�>�L~���l$���FY�G?��e�Nk"��vE��=P�I��V��1�X��y۴T�"P
�D�Y��e����Ѭ.'�)]��/ɒP4� [0M�R��}��)돋��[*�C1�A�����m�4^�Ū�����	;�ɮ4����v �v��,n��@"/��(@t ����hH�yH�Z����T��t�J=�����,Y��qq�
�Y7��3Ǌa�@�-C�H�L�~w���Pň<{W��@���Ɔ��A��>!\HƏj�瓦P�uM��3���qrLMь��s��VwX�T��Y�[��T	.��E���TA��+���>T0>)�\	�.)/9a�&5��#:`N0�6�*~��ʰ��:Z[r��E{���7Q0e*���v�ɐ^����1�8�)�Ą:�/5�
ź��:CWJw��p[��#�C$�N�y\���9B�2�\n��� �n��|��Z�_ljz,J�3zO�{ �_�V��q\���}lC��M�zx�#�ʵ�=�'�M�Óm�����b|���p-������e���p�]��Y)�"�~�_�Eq�D����U��G|�g������aYh�W����oyr��/�e[��覻^ھC���w�i�bky,�^��0��e��Ց�H�a
'���҆�@����R������-�:WF�q���+A��ʮ4Z�ty=^'<s4!-�� �0ڇ�K-M0��D�A�S�L���3$!ֱ�Ү�J=fj:�AM��kZ.\I��=Hv
S=�p��f�^톰e�gI�E���?,���V �v�֒{;6��s-�J(�����q��2Im1���J�,�l)��f����~C�N.����'�\Ĭ�>*A����j{wl��'���t�mָb�&��5�;Q��ݯP3H��T0ݨ��+»���Z�]�Pof%�Ad�b�ʸ]fh
���������y��S�v=�;��@T)'�M|:����ـj�wLuZܾ⩖%~5HC}!),E 1�&����,�(J�HI|Y������"�5��� �A6�8�',U�����o)�{�q!����r=�����y�!%I�=� M���]���O&/�	͔ W{p]�w`�>��uxe&�=�wA�r��w�8�0}B�jRHD���<M�I0s����$& }6���`*G�����@���o�X
���c����o�u�\-un0�a�B�&)�jd"E?�k:�i�Nx�O����`�D�k,��U\�	��)ֽ�P!W&/���b����㔸�s4�>90fE�0 �nƢ���
E���
���y���ZY�W(�)�����{����wZ�F[��1z7��s+9�\���->xj@x���c���*��l�qs�1�Na��̐ET!���L�-/�(z����w7�'x��_����v0����]S���h&�}�A_"E/�o��b)���"���T�(wf�4X_j�|��d�j�	Bn+���Z�%��)//�q�G�#saBL�lɖ�jH8"���g�=w{U�����"��L��(0ԹH�q�^A
u�!�~yJ���]2J\�#�!�}���X��$88dS�:IJPL����al�����B��l[{�˰NNZQ),ʯ1�#�Ls-({x����E��s�@YU�>6�q=%����`�;�^����vW20�H�'�ԈO���!NJV��e�5	�;�}i���[�|h�ǕZ����>��y%O=۔`��S��s.����]c�9zff���])��? �V�?!$�(׉�%GT�4�  f�`R��͒Ju
7ʮ;��sK3WU/�1r�l��*bn���4��`�d��؉x�"��Mź+ߌ�-��h���sS穿P�}uD�168*� Y���3���貖kI�p�����h���ՖW{�]4���I��:�
b�����3甲��F��Ȣ=����j8R��SH�(�ƻ��i�?�Q���f)��;�:/��ł=�埅 t�kp�&�]�-�uKg#�;�LϺ�]��hߣ4��So�
�҂���l%1._��V���[�'8Eq���.���=�u�8�Y�ŻB����2�rw�p������M`��*���qhLX��*q��$�cYي�N;�ʈ�0´ R��i��F�.�Ya!�r��_�h����|c��pߔ2���w�9R�$����E8Z��O�-Wd=�m;��%��
%��`�k��A�o8<��C2�G~��2ͺ�[��uX�����������`$}�������h�X�N^{�7ׯ���$(�6Gɻ
�o*�	�BU�U�X0�u�7�/g��UW��2�0�b��ؗ�awb�*Q��s�����&d��f�M`^���z+�+mu������3�픀h����>�x`1:~��}b��[��6��W��x|e̩%�y`�m����αƷ��&��E���5�t3�ے���m�?�5ʪ8��;����D�i����ln�S�sG~*E�CݨӢ�Ƞ�~���F���/ג肕'f_�w���� ��P�������OT�-B���� ��R��g�@dX*Y6F\2X}���b�z�1�����x��Ы���gSs���W=6%���ݿr�B�(�w'�wI��+�.���Wx-t��I����V�{a|�$ק��ޜr�b
0~|(�,�-�Q���J���_&�I�S��0OLY5����"Fǜn �.#�/y,g��.���&pR����A�Bṛ���+�6:{c��p�W���Eֳp�[���K�o��i6/W��3��ĳ��s�&�8��Z&�h!�Hz���Weq�x�s��?�d��L0pS���"���,ʈSG�㑒 ixU���4� 1f˱_�Z�,�X��G��죱�IQ�O��ɍ��i�ͫ7��a��	A��l3@I��~�	�y�
��Dڈ���4��Q!�`n���p#��*80 h��v�]@/������9���q�:C`���H1���0������K�/\9�
��C�?�
�#���^�b!j��KG����1�H�%S�������ݞ�|������"��U!�no�ji/H$ѐ	�=���%��1�sQ�@��z-�7eQvÈ3����)�NH:ɣ�  �n��R��l�x�q�ڡQ�8�`!vEy�r�j��<�V��6�������Q}G��K���V��2������S�1���3#u3`Px	�Oc	��TOQ,H�C���n�1ߘ�q�ģ���Z�҄>G� �sR�Cq���KۗT˃�Y�i�Us�3X<?�x��#j^+�M�j�:/��/ye{���,ehtW���|��'-v��*oG�M�|KQ2�7G^���`K��!P�2�@E���V\��_�r�xY��� �?�<&�?�T@��v�[gU���PG�9�M��V�rܠ��Me�6RZ����k*CX/(����������6M��#��F�]�t��@W��)�gqz�-m�1���B܂�	)��c|e񭠦�dYտ���v8��5���~����,��x�9!i��؀$ ��A��!1�o����&�\�M�3�*7����-;��!�В�W��*�˦ ��̔Os��mfO��;�M��)\�Eŏ�dTț�A��t@k���΅�a�<+j�����:��/0e�˔��ۅ�>G��I�jȪy��}]J�� �8�y��͂��k��G��Z).�\M]y�U<�nVI,��<m�ǵ��fk
/-�6���`��|G�Ax-���?#�	u�3�S���"4�\Ձq��ն<�T�r�LG~!)6w�8?0e츪p�p�)^$ԗ�9�(RM-���~����'��<��3'�jr���_�㹛vF������=�ou���*������`Y���iN�"ʁ粼� �9��D�O��0���)�"|�w�V�U]������!m6N�h�	�L��H�.��n�7a��]1��s�N��[,8ͼW��;��N?�l@R�v$�+4�_�*2�#B��7il�9��eɲ�M^���鼇���>}�h�\.�x�2H(���N�*x��U�ثE�ZG�� j@f�ל��Ӈ=�==];�r8�#��ϰ�'�GL?���(��0M�c7'�&_9\3� �}fD3����R�W6������o�/�H�E\ ��i��A���n�-���Q��0_���	'�c�(���4AI,1��?J��6c�b5�.ǲ�%�㝰��3[�t�ּ���}������T[CY��s����1q�'62X�����e	c~Ʈ}��w�|�e�&9���Á�栙ݫ��A-��I���D��Ԏ�i���W��c=�~�x~��u�4֘Ӥ��9�p�dyN�=�N��Lne!���������TO�d�X��pt�7��Հ��f?bO�;T49�\ԧ���!duX�H3�) �n�]�ʵq$`b���ЈNi>/z����b2�,��V�b���n��PhtѪ*04�#,����%5�;t).�z|T�K˵ެ=�	S�-.?��+3t�W��_l����=Cig�~�>d�|�F⋝�hCOܜ�����&�8��s�Fj� R�`~z���ն	T-Ҝ
�zػBv��'�������,匍n'�y�ܲm45��I�5��))�r9�UxuCͳ�p[?��=J�<꜂��c�e��>I�� ��poT��yC��Y5S��dQ2\q�����oCK�72�1#�����N�m���R����e�;Qr;��� W�0�O�QY���X<hr0�Yݚ�X��쀤���.c��{��}`/��h�2gH�3�lHPr����c�l3?�|q�u+�u)��xOm��*%0�[uO74�&������>Q�k�  ߣ�#�4 ��N�6��_�׌��:���ʅn�jZ�C�k.�SE�~�t�z3�	=lQ�60C|�C���5"���=K3
 1躿�1�bq�vS���Y�9�p^��[@�G�;eU ��B�!�~�J7p_
#)����`�՘@$�]���S���:��E��E��ӆ����a�?�?� V��l��t�������v�,	T���k��_ދ�xV� ~T
}� )����!O	$����R�,K�P��潜qy�G.#?[�*=FФgiQݛ^4���=ퟔL�KC>�����V�U��){E:��_����� ��}���h:uä?�'�]ɥ��[��8hR�Yw���â��k����
���V���l18���H�_2�@�*{P�p�ȌfK��2Ŭ��G���S�W/��a�%�9a�/����a:�q!sp��+�6{�]�j`�����>����fu[c�i�H�T&��E{���:��{s
�a�(���FA�C�z�Ok׼����C���~����\)�����1�Ҹv��t㨇��>��c�S����)TW"EOҤ���2�[�\n#h��k�26��OȷX�]o=��γ���g~���������k�S}q-p��D�++�?~5#�A4`l�nu߾~NW��rE��/�Z�,=��힯`v�TN�I-�>�J����+��j�y�%���kB��"Y\�K&��v毭6@���0m������b����\�'�(���H���2N&�V����-�9�a���^� �z���.����������Ԙ���y�݋U��6w�d���{'�)�y�e���*�;�����XIP$�H��ŭ�'.R/(--�Sǔ��:�Ze%��6����숞8���VLzZÖ��bkM�����yPq�!�bN���\+H���N��Y`J��gC��{��٫+(%v��9']:YiO(�bS{���kTڴ.�D/�8����������U�#��*�6�&�+�@}Ňb���O.��~�
;A��NB�NON��#���66>b/�E
����@��i�k��&������cX����~s�Ԃ��18��l޴�6A���y�4�\�˷/�u�@y��!t��:��X������o���ni��l�)$����69�@�*��+�~�{�������l���w_�`��#�0�yxl�k����!��Z�O�5GdF�P��0ܛ��
�./���j��+FU��������P�,��i���Z@9���<�EV�b1��R�ﳠ��(uD�YX7	R�D�Z%��~F�﯂ 5����a
Ҷ�/���L͇�萊��������{�@��6���R���ȎOe�E#�R�D/��(�Q|~����� ��9�Z�04�rs�W.�3��#3����01޿�La�>�Y�I�b�b`W]�m'qfo���~�wSa�����Q/�Drd��H1��EJ��V�	�$���ڜ1�w�Q䂲�>�_����Xs]�b�k����b(~�XK�` a��� ��S۠>�jz�n�v�yH��ε���Ŕ�����Uh`�zs%؞KVV�;��e�P=F@�M�b_���&9�׺<�?�����qU���a��kB���^�{����sZ�(���?"o�R�|:$���>s'斚��&Ɣ�&Ɵ�C#?�D��P�������f�5V�,���ߓ��/2���-l��`M|��c�����E؅1m��@*��
�TR��c�{�xE�(���χ�4z��^jګ&,�eĭ$oom���X�Lߧ�� 7'�qf��Z��d��W$������J���1$8��/4"��_\D@vaD��`� �z��������L��c�*���q�0J5�ˊ��"!�!蔶��X06-Y�ҧCX} �Ob�����\f��g��Y�v[	)��3)�[2hg5�[mi'4�hq�w�|h �S-C@�"�PЙ��!7E�H��[�hn�U`M��/THV�m���2'���fKI~J���%��~����K:��q+#�f�@LR`&���=�KJ��-�6Z]1�8:�v�ܛ�<��MS��y��!h&��U�U�+cVl��r�$?dZ�i��8��#����-k-�yWhN��|	��#���h�t|���^ܬAay�jJ=�_�ٍ⇂~�Í��c[�y����9Ts��:�����y��.�\���a�gҮ頴r�O!���(�ͻJ�����
ֿp�ꟲ�����S����6�!���W���Q3���QM4B�D7��l�qXAW��@[|2�8���kDv~���T�M@"kn��E�a��ڇҞ=X0u��"�׹���/q�V]�~F����]��7j�+�К��ޯ���@qQ�KԯG�6�7��[^,��e
���R��2?u'KWX��*�zKC�oE�����Q.l��]�d�=0��	�߇̻"/z �C�uy�W�~C�h�Z_M�T�}��4�9��Yi�ƲS0=K�S ��(��&��Zʀ~y�f�ទ�툘�,�V��Z�����Irjۓ�[(��>�5>�\���p�@��׿��SlR�NA%O��p�^��t���)Ӂ��"_�[���|e�xׁ�)7M﯑���"{eC`�o�`����˗I�`wr0�̚M��bա&��Avw��;���Y~��f��SJ{>[jc�Y}��V���>��An�D�4m�&�f;�q�f�h������V��� Υ��,x�sc��s��(���Sg�(XP�a}�^^�mr�v��<�f��Fbh�Ǟ���z�͢��pD�����Sݜo��Vh��}�yfitSsa�dL�༎MR�a�p��ŇM��u`�C!���kI���9���q�vb ��\�괙S
���y=��]�F����e�]Ȑcy
���5>"��d��2��wuo�*�|��8q���n�Z~?���բ$�12��n4��u{U���5[��B���&�$�WA.��,��-�����!��?�{�t0_Pc�|�+nr�D�!��;��C�����3e����0�
�	�I����`z�I���U��s��ׇ�لU�|/���{�`�>RIX8�	����2�hΣT�Mk�u�,0��9����Z�b�6}����IA�8$��Q�L�S�N���+#�6�9����e���F���瑱��{4�(��
W]�Kt�2�|24��1�:��܋�󟑉�m���{�[�>�������e#P _�%EHX�_U~,��ʝ1{YO=|Vy�v���&��N�����һ�~���c�3�b�nT`�H+���ԺӷD�o�L�o��ْy��E�wb|�4��&lk�`(��-����i1�Nl$�]�������H�Βgmv	r|��>	�	8�2�"An��$�ߟ�[������e>��L� �;�gAM��w���1�����p��J��=*MG�����tH���t��"}�I�:������^���{zΌ�]A(�U�C�AJ�6����o1�J�[�{�A���	�I�?�@$����Cʝ�\�6�����[,4/��� v"���J����z�⿨��g�[��ٿyݥ�gWWS:3����Z�6�e�4]h����[���l�P��V�I� ����h���:�������N������n���W�}��q����?��M��"MW�(��rF�g����-�y[pY�=�EC�F���boD5���/J~<��%d5�v��]_D4[�h��o�-�i�(䵓="O�T���.J��ٛ#�tL�:<��b���	3�q5䌸�0k�m7{#t�0���.�=�׵�=�<ùW��'���Ř��b8�X���<=�a4�b�I��J"7zp�������A%@���5pH�Ɣ���h�T��I@�h��A��}:Rٔ)����R��oZ�  �;��\�g�?�y���d���'��=�!�y ��0k$}t�k�E�Uiݯ�)����w��^V��!�mY'b�t��mW٪�����f���i8���bONK�X�����-�]���Klj�`ana ~��t��J�	�����9R�3�ĉ<;��k�>���,��ӣ������[�0���y�KZ���H��OYp�8�򧻗A�3��aTSJL���|�[]����	=�-�����`��-��8��ľ�LE �?�^g��dx5��F��|`�N��7���eBg�AA�B�2��3��c�h|I⶘h}�b��M}c�L���g�n*p��9�P^Fn��zg�k`��f����WRi;�4���b@lh�R��G?�;l�zHf� bhm<��F=�:��rG�V��JV�D���m����]�*�K
��S)�Û�{#+�jS�ˇھx�XΐnDa�ti�D&���-�B�t�����o`����/S1���Ò�u��$����N�BNo+O���-�����wj<����� Y�B��W��+8���Gh�iN֬��|��g��������c����@9�C���mŋ��TJ(GH�pɩǜqۂ��\����u��'8(�kow��bn��.}l���M�ug�`UHv�y�ۛ�r]���+�B�I|Կ����F��	Sg4���L��s<2����A:iq�Ģ�6�ab͜����8�z�e�x���������!�\�<X�.�jk%�}��f�_W�F19��.>��W	��4��-=��V���p�J}FKu�e�M�T�u�g=�լ�����,Ǉ���b�(�s7�z�>?�H��&��3�Uc��m7G|PS��P��j�S�� �n��pQ4�=@l_2G�&�;(v'C&@�����|ǩ�����h�mk��t9 ��	ߕ��������R��P��=���0�n�f�98��Ϩ^��O�!ޭ�N��`�8�m
)���F�����c¯v�7���i���ٔ,	=�k������Y�n^虡���ʬ-�O�d���d�n���z#0�Q�����3��]���Jn���3�� ���q��B:����t;�#�/��ov �;&�7�ܝx?�)�g_���s����'��L���pAB����I�G�R�;#uﲟZٌ�/�bL:�NY��Q��)S(�D�F3��y
�@.��T&�>$��J�Ɯ<T�wXf���Ksʅ�C+�&dg���C�ԣ�է/})=׼HY��������EK��P[��~9tßQ�)�B��3-�c1��b?L#)m���dP�*z��[q[�IJx.Z+aw�V��]��>����	W��W�Z�%���X�h�����{z��,�?�$%_����.������}���Q���O,ΕF�]d��jU�F����4`N2W#e}>[5٥���w���|���3��]��hbm�Xu���![�h���㨯g�tl�󹬦��9�%�:J�p�j�����G��[�>�Y������X�O��p��'0�Z������V�&�G���������{�6��v8���s�!6��h#x؇���\(J�����Q]Z�OQ��{������2�,��M��M�V�c+���&=�f����]��M����פ�<@�6�se���h 	'`�]�����-��BN宱u���?\���r1����1������"~]b��Z᳌��ԡJ>!��+}	��j�D""��|ġ|r��Ef���.JԚY&x;�[,���sw6����_�� !�و[�������l�;�W�pϩ��lĉ4$�NZ�/����9���黷'R²�n�մ=ą*�%8��Z� O9Fjpx�KtX�Z�\����d���RU��	��\�P>���Lj�8K�-�x3���ˌ��3"]޷!��gv U�J��J7��
X+�"��ɾQ�:]�j6��������w�ky{�E��9j����A|��+�G�BAx͂����s�P��U��� �Fx����)Zi@��/��l۵iC�@S�J9�9�NK�BB�����K��H���܉�U2�,T��&ܼ��b<d_��I})�߸ Ji{��=�O���]�:)v_I��;H�G���ޜ�|��L�"���e񣻝ϝ�GN�"�&�չ8�y_,`kg�yQ�β������@N�҆�[1|U�ٓ_�39�֯T\�{F�xE(�X�x$~�b�����=�aEU�QW�/O��D���ʣ֭A7���~
���xu��&~����7�h�%�Q�>�����(�LS�|{��m�Z��B�����Be��g�z2��4�UQ�$cc���aFC�'��W�5g�%��_���0���؀�V����h���7�;?6IV�����x�����e�O�փYZ׽}��ڜ�+��'W�� K`��/2V�03z�l�:\��W�BO�-�hl�m����NI�â��GO3� f�SNp�'�-��|s1=�G5�%Y3p?�R#���B4p�$��^�,Z�.2����ӆ�ҪB  �H��|�����E�ct�@QEmtq���(�>�D�Q�7�Nt�dI5�M���a@Md�Z�X��R~�χs:g��v��B�.�	���8�	��X����ع�)a[��̛����Pn��Y�!i�iE?M��ek�9zq����*}4�lP%�Ng5H�#��������ye%x鶘O�|'<=�Qr�wJZo1�|���M�3)/T_��+�V��#R�r������]��^�mh�C�D�e$�x�K9l��o�Mc�)�g�9#���U�/��I4�k]L��X�t/oV�DNt��M�c.l�|q�p)Z�vѦB�34Z����������t2:徤�OƊVq��Ln+	zZ���QZ;�O�N�m���O���P)&.�2�L�NI��JY7����YO{V��?���U?��.ćRVS%>4�0������{M�c��\N1Lr�X�}��޺�VLIQ_���I��뗤
lu{U���9�f�O��\/��̟�j����{n~�dӭW�б�V�ich)#�y��p��2�|����J��j���c���Wg���
�t���/�a_ة7Kl�g5����L�`-y�?)>�G$7�v�S�P�m�Ɏ
�{�?�/��zI��Ǒ�T�FU��9�(�����S�R6�F�@�jþS.�hX;�8�
)½�I������?SH$�$�Z��!4�/5�'B�T��,r����|޺��i%wv0-��*	���1�áx|������/�aF��Sd�q�K��f���L&��\��;��*Nm�2B8	��D����!2HKa3ڶOjMM�ILW��l����|��㚄�����a��)�$�qQ��71����q���s
+G7QH>@����D��L�w��X9���s�(�z07���
���K����*��07ec�a�e�b���~���z��9�[�P���5%ꄮȩ����ԢQ�lrX�D��kX���o�� Β�ٱ�s�O1߬�R�ѹ��(.٦Q��ס�2:��t|� �E�8d�Mxq��������\Yə�*�%&Q���}�+���NT*�KI	7�=�ADD�1,��rD��h8x$�����Nc��]]�{E������t�]��b&�����$	���_�;�hnp�ˇ��P�˚48ߧ�?cP��nc|`�*�8��#;7�`q�ir���?@�qYr{W `{��1��l��ٶ���--�c������vP�wr!���S�G�knL��eNt񕍔��F�֊�x�XAOC��s�&u-���&�]�{ĻF	 <�N}׫���`�Zv��.ڡT�R����+)�=�BvVO��kxL[�:�,c��&�bG>!B�T�N�fbMf�&�]0�м `#�u��Avk��͠y�*Ŏ���=O�j��ϫ����Y~h<����G���v0�NG��A�����DxpJ�.�݂�RM� �1�T���7[P�|Y��QepE����Ul0�§A���/׃q�6Y��x�t"<�"��D��
���AS]�%�S[�p���Yt�fT;��Nc��|�h�[5T�xsz�<{���\�>����Ҁ,����v�u���\�ét��6�	[r���K�4�)���>hGĖ�'�:o'J�\6�J~�L|I3���
��ǈ.O��?�c�{Nw�?�{�'uU-��]#"�ut��_t?��^eV^����8j-�Fi�	cc��n�Y��3�@����Ff�$��͙7��y:����vr�� �}�ER�������� �ɠ�}�v7!0�~Zk�d�6��
�x柆ه���% ���r�P�|j�Ö��[�I
^���)�;��f���-]&�C� ����t�?X~����38.�xj��^�?>��1���2�^�,w'AADxT6�j#�Y��°����
��y��g�[�� �a���u¾*�To���-;*,t!\�}�6��dhQ�sU:d�4���)�Z򳜰����p��m�C������aSG2C�X>0�7wM���t��t����0Ѷ�X�	*�,��q��oo�u� loH�=y0a�p��(<������N���L��g�����`t�P%WzU��7j���P,�O��}��9�fA��_~���z����K��V"¶��[\�2�����&)}�T�OG�C���Me��O��p�R`Y@u����e�M�K�N�
p���W�y��'H�&�9�sl�γ��׌f�|k!�Z�u��pƹ��H|Y���2�f)�!��i�)�
�Юj$w���u!��_�t"��NnN��v���{MV��k�[�񥑡�'��mFP���eS���B\�rBn������������wg���qP�J��(i!�<��p��p^d8�V��{���.*��v�G�N��~H��C��D�D����=���G��Ds�!K�������2��2L~b��#k�Nz�"�)i�NJ����(�N���͕i���K$q����e�3�<Ǖ2#`lB�i��"b����D%�x�Z���͞��V���i�[����"�a`X#y����h�s3��/���2�A%h��+���i+ynZ~_��kf�9�w`r�4�-I5V��ѳ@.M�i���|MN�8�"���?/��i��Ln��4��a/Y�{���"�PoO�y��mX�t�z�#,��WD�>C|v-�%��,:<&� ���74�"P��k�}1���!���&��Jȋc8��g力ΌcC��B���t��K{@w�6
�B�bd#�V��3�Z\��V�G��e@zp�<��}��j�?<��^��,@k�v�6��P�Vj�>�,�����f���=�������Ocma�M|(P&.M��xF3MG���'mN2e?�"�"�Ue9��9E���nu�d�)�Z@�F^ш\#ġiYz�h�����Z�:f,u�� ��0l��(z���5�7˪���2��gE�?�V9|��GFޛ��4ک�VQ�>��JY��Ѡ���{�]��,z�K ����~p|�]�/�*L���0H�2wq��MfǼ/Z�;{�ߎX���Kl2k����5	�#ҕ��h����%��$7*�������N�iC(��YDEA�������A�<_s	��-����E�T5U���%q�i��)�:����M��;9�}�y�}]�pVF^��_nq�٠�+�3�l�<�i��D���7���{ёo�U����M^:`i �s���L�>ڍ�X�Y2l���^i��b����-"�(�kx�g��OأV�x%D�4��WĦ�L�?���1��C���Yt�f���JǨ��0����"W#锇Б�<T�G���Ӵ�2�;�Ij��ػ�Q��-1v����>�o�E4`��&�)���HW�J6u�&����gJy喷�Dq����5h����t�f5���o胙3�����j�S
��dN�m�N�࣏�Tч���X3Q�
��IX�@+����o�VPD\����E�hg5�@<�R�sPx��h>���^��8�@�+1�����[v�>��c`�QBQl������e�nv�~�x,����w��U��ߴ͝<�͈Z1Y�>�.�VT[�$���U�A3����t�0B�2�d��ݑ:Ţ����#�u~,�~��{1�o�Ȅ�Ed6��#t�:�D��/���RpÎ�F�'�N�p�T���D�ԧ8���|����T	is���4��|���/N���a��Z����TMj-@ߋ�蜿5#�C�[$i���� �~o�F�;D����(.�b�6�J9�e�6f5�����I�o���!��p���M�2������;�TH�n#�݂�������*�b�HR�F����\ÙjGDׇ7�����9{ß�vdU��)tMb�t��z���wq�y�W%+Fh�����{hAy�xM�ue�l;���N4���gL�"��ap��Z�D��J�����=������nVV߸��iZ��U�J�v�}i�hP�ԑ�#քY��1�ݞ�^�!a1U��kB�'w �*o]e�,���u[�'U}�a��ABzPccz֡�Z�	s�ŢO�[��K)�d~b��&���.��T���8k2�:Eę.P!��0��oz�i���;�}�";�E�6c2ޞZ�n'E Aү�{>h�m���0�_d�s�}f���S�́<��2�����jLo��[`]_���b*����l��`�\�Ý�qOAͰ�\dz"�{9b&�+IY�&dzn�|tO�W~�m�#HA��d�[� ��7��+�����X������ߥEf[��u���Yp�� T!3	��۠d.��9���4i�]�WK����m��ٰ�.ޥC�S�ܙz�����ZXH�n<p]���>����a��[5���p+���M1AN��V�UL�K��ӣF�j�ӛl j�!^'x�>��rv�Ye$�S���"HI�F5@�5g)o
v�lf7��	�d����xs���c���dL��a7�,;M�k^-���=sU-
��w��$,W�+@\Y�豑+L.�	�3�����w���=I ��s#��f1�:�;�*�=?K}9�$�����z _��Ay���A�O��Q�B�ۮ�}�ں`	i���Z���s߶��Q8*���Io~L�0�ܵky���ƂVCR���~��\�]>�u򂌮���D*�ַI�N}���|��?��/�$�`��܃�KF0�[�����!��ziM����uC�ݴ��<1a���3��=����Rp���H;�0XX���)Lh%�2]y�K�z�Y}���4�����O��1��u:N}�q��I��WD�P��O��O�Z�)�r����&��ް?�x�ي�F���V\C��j�<�5�)����P���H����u1r���IA��ٺ6��*C�(��D� ����*T�Cud���x�S��� ��F�v�t��_��e��iK���V'}js�R�Uw����đ=�	�L�&��#�-Jv@�� ���/��>'٩��5tcñ��o#	E@�?�f<דk��jG�^Q�=ys^����m���F�G;=�!��%]�dX%'�n�tMa�X�Uj
�X)��8[v��s����;�bA39���eG`��I|�X�*�]�)�`�范�u����M,#L��A���$
�Q�K�܆}���$�im�E�	/_Q�o0��C�bo�󖥨dhT�6��S�y�)C�#8��Lf�9&���ЯMϋsa��/���y�S����}������� �}7yLa�a{ 9o	��E��l}7��636�ʢ��T�,�k4d�þ)'���Ѩ�.HR�6[���y���>`1��o�A� �q�YŸåbS��(��e��MU вj�9��e�wnp,]B9��rnJ�ʞ:#و/&�',3]9�	֯�:�o�t`}ԛ�7�H !u|X�7HS�<rS䃑n��_.�͖Sϗ�l�d�clS�H�6�QNR�:����	��Xw��>��#�gN��J��,�20ݿ���1Z��_{?/���8�[l>�C���(�՚Z�3�-���u�"�[�*r�.�O�y��ȕz�u��Q��/���.#� ��B�L�������>�gX��(� ?3
P�Q�d�q��~r�eF��9�� a�Ȍ�O۔�9n'��z��:\f���{�o�\���@��2�C�΢8������
䊭�`_�[�9�8+T;Zu8���`�1��u ����#��6�g�% XtR��T����0p�}>ha��Yo��0�\��4�{�'��\S���b��y�\�/DLI�ߊ�u}d�o0�r�������5��E:�?V�iM>(;r�ȟ�z�(��3ߺ�ߢh���z2�ڬ�WG�LN�2S�N^4h4���S{��K��S��v��)£�K$�K��rA/?��3���#KV	�p�1��\�o�좋��lt��_e�� �ݻ���Q
�+M��Z�ѓƠ��R%��ؿ^v��,�8�ӑ�@k��gx��(nӧ�#Y#	����N�ދ�E[�����uB�>���\g6��!��L���YK��y�:j����wA��T
�qi��^ow,�q��P�?����ܢ��?3��UN֦	Q�7�/;| !�Զ�P��O�I]..Α9�_�{����>_:i��`{k�4n�jM�NW�Ӽ[�qy+$�0|��?#�N�4���`���4�j"�~��$d�H�������3��GaCw�"ώ�hR�����W;�~uMwi�o����{�+�T���qG�=���bB+��k6��w`�7����%W�!�g(�%�ɌB��5��uE���˯*؄�ؚ?@>�?6��NF��˅��`ܰa��#���`43E7�P�P�qý	�q���'���ܟ2����ٚ���XUkh���4�22��� �S~�#ˋ����3�<���N6BQ=��dc�`).�vr�z:�������Z{<Gd��mT��|��d]Y��}��dn��/�(f\�eqpa�����X���b\�M+"������h�n'�ۮR3���Z��(`Ϩa������"@��L����q�w�m�9�y����B�]�+^�<�@c�O-Ĳ(~vk��8)���)�/vkuE�˵OAu���p�uM���"��Ne�L�4���ܵ�H�9	�q,8s}�K,��ڜ9ٮ��[��,�V0������c�y�+S ����S!cHw����0��%�
l/?����)v����ELV~ђ������Q�V�'��f2������	��w�,71����z����Z�!eN@���qy7���ɔ����_w����9�������=�D�>�P`
��[���)[%���i��^D�c����q�7|Ъ��}o:%�u�/�IԒH���g�.���ϑR�?ޗ���g�[�����'��(��2�݌�6�e�%��Z�R�P��6�äS�L��� ��/���b�wi�i� �6�VK`cݗS�G�.�ܳ�H�(9��8V$��u ��F^~�	�uM�;���.w�O�l�QP���K�D��[�z�G��m?���9���1d��9;N
i�D��;�S��w�U遘k�u�w�Sܯ���'����)Z6$��uu�!􉲰m8|���4�(}�l���ɱN��&sH�Z����xs��S�qO�Z�\w�����,I��S��Ȩ��z�]�ō65�v�T�*(d�*�Cz*��V�,�řIn�o��UE��0*���x�6@�����&�ϥ��"^�~�����#�',�Eӫ��v�B�5t��n��w�\)LN���/\T�X�E䮢��cU��"9�"��lT&��^`�,&h+r��dbc�mD훫Q`�CP��1])Z9oxw�H�*z�O�� �Z����VI��fD����0¯پ�P�n��2������� �V�䃀W��ײn�.=�Eb0.�����8ja�E������N~oM�L���gc=�B��!�\07�7�<�ùxɄ7Ż��:�v�n�9\���h|���#�htV�M�A����$"��4�!_���=wv����38�U� �V"\B̿� \�}Z�n���(f�%�޵��"w��+��.f�#���5)<epDkA�x��<v7,`�oCܾ�(�
8��3���!�m���w��}�@����S�9�����K����_#}�Z�S���������~�|X��k#�:�dZ��΃%��~��M��"\��$mR�Z5�85b�>^C�g���\�q'��Yhg]�*9��8��0#����j�ƚܺl���]�Qq�3N*O�r��x�7>e�A^sj�����(�6��H
��I���
8.��UȓQ-�&;�A�=pb������oHr�\�W�'6_���H�������r�z	[s�%
[Ԙ��I?�������ljsȓ\�C�ф܏�D�>���|�IkR�co��LF1 ꜧ-��{�����*��Ye{�'�2�5�z���\O����￉CO	�!�,��H7�6�'��"�@�}��� �O�f�:�F��鶲�@�[�Ζz-S����Q-Hʌ��'F��w��T���|^9Az����5�֐8�"9�3n���d�����MC�=Mn����<0���r�OC& �<5�S(�}	�)��k+��\<��
�0f��<��q9ɛt6N�/�g���{4�a�slī��a�5�c�����j~�T�f��;{o9���aY��60&�� ����é��,��YE�i{?9s�;n�.F�AV(o. ��#oK�j�;GT�or�r�cQ���-!KS��5C!�����eT�+���5����م
�CM�'@_lm��@V�v��C�=����h�Ƞ�i"���Q��%��ĕ���l�h�m�5�+�~lf�M���vǲ�}�#Y^0,�.��������XD��l����Y%&u�ׯv�[���M1�+�y�Yhٝ�x,Q�o&!�y��*5*89�8���7����;� ��Q���a��Q��p�qi�cD�3�"�븩�-���U� y�óí��^*.��@�<`���E����8�|]�G`�Q��6�_2�!�A6��"]�z=�9l=U 0���E�&�P�,��?�G�Y�B���RKf)��x�.�4�~�E�6�-nVT��s[�Q��[� 4|Mw%�&T�G��;��w�
I�3Kr��	<l�����,�BY��>�l��"v�h 9)}3�D�9��10@k8��4�
��]�d�eA��,)e�?g���y��i,u�zL�Ύ�����*�J�F��HRv9+��es~����ub�^b~[�U\+�+�#������3���B����Q�z���_0����yH��#�KP�:��ֿ�}
�b�Ul�#=�T���)őй�V��3�r.��5��L���k�,����EG���\�Y��w�*=I�3ub��\e��n�S������g��X��Vvy���rz���tŔ����8�#%1��Y˺ai�� $��Nv���c��T�y��-�d+�P��@�C��pT�n]���u'.QA^Y;�	�!5]�w9T�1��5'"�C��hxv��Wm�������V���ы�O����f3<g'�%���dy������X�\��Q�����m���N$��Ek�t6�0�|���ƝA/{U�~~Rt����v9h{�"����k�$/mtX{�VE3O��U�އ���J�JN0U;z�Q2�	��0AG��J,�����ԩ���w�$�'�ME��_����%AL�eHKјB�^��q�nH���]?�Eb�UX��P�K\��"�����SA"���W�U��t��) tZ�Y���)w�Bn" V�����~�֬gR������\I�2�� ����}UX�0A����ǫ��H�<t�.�,4��W��R��R
�|�H�Vy�*N�'�w�������#�p���1=QAV��QSb�bW(o��(A������\x������ا�<�Rŵ�s�o�#��~~"ݾ*�BP�W���ߑ��_���y�nڏa���	G
$�DZ�ک�ݦ��;��E�����U�Xo�ϠQ�ʮ�gTMM��qp(N�q�"oA�|��N�>�g�c�+�E�Ys�i�K̂s��&s��F��G�*j��J:�����:�5��U=Y<����R�Y��Ǝ�?��;�"ɸ�3$�ظ��Bp�E��+�<g�kWZG<�/'� ����g�ʳ�r��x~� Ж��#�~P�fe�GP%��D�ͦ��ʓ(�_(Q�����(?0m��aЀ��%�ǦuԆ�8���+�u��1!"av�@GH%U��叕��XIƜ�Ue?�θ��N_{m�^d8����E�$�_�2��}�ך��x�a}��S��&����X��bx6W�uw�YA0��(G�v��G'���cF>��B/�ĖwMQ�z�����}|������g�i�b1G\1�A3L�<9e`K�t�����C?�)UC	7��&��j�c��*jD{�.����O[�>"���=���$�㬺�$���
� ~��֫�1VeW�dF)6��0������+16��y��"u�*�Y���h"
�'�PRG�r,gU�����Fi�(g|c�-�5y�:��3-�!�?m1�>�|rA}�J>��)C'��d��%����� �m���xoS��,ڤ��0���Ѳ�ZlÏs|iK�׫��g�`bۮ����9Y�,e�6�ֈ� �c�r@�E�bd`�kɫ�+��s��tn��cq(��)p"����G��J\��*'���A���S��!z@��:��❫�����3��G"��a�/)�%Fsꌦ�}��"y �
%�`�gtxMb�Ҡ)�[����tﭱ�D��<�&�o)}��!4�C�^�zSɌˣ��?�鱮Qb�ci�ỻ GX�)Sr5��G"�.�H�D�}0�1�pu�-���;>���爯�#3�������c�9��*G�1"���.U:GZ_�����#T�Y)�����A�l�;3�խ@������7���<ߡT��E������鷹���X�M���Wջ]F�����F-pB�+����e�ug�}J'uϔI�rf��TKh[(͘v�f;�`��V�+��K�`�F*�a�����yV����u�"�6���2.�2��_тmU��sU��i����+d\�� m��,J��#�7��oh`���t,n��M�3v^vd�+�$z,��}>�M��j>.ھ�eR���&e����Q�vg5D�����G�ӎ�4^a���ӥӵ4"�*:I�t�g�9�ˠV��)�O)s�J �?�&�����b�����]=_��Z���~��pBn�ϲ=�J4��@eX2����j��3��~�X��m�l��"�>�L��v��iAw7�Z�!��L��(C�>'Ps�ƣ�6�8�f,�'ֶ������!���Q�|_]�V؞�M2o�+�2�^���nc��у��W�1Tk~������/݊�O�.��M�A�9$p�-ևgb[i������<j�:^Sl3���<���[M��iA���n��0t�,Q�8��s�S��(ߩ!m����2@�DzڼF!��L$ً-NIw�k�d:�]`pe���x$},�ܚB��>��(��a�;݁���Fd�R�;uZ�bOf�Zz�N��ȧ�n'F�����7��>7��D-����AJ9ц;<DH-X���ۿ+���3����5w�̓�����h������U�D=w����O�Nv��N�>�E���I����Q��V)g�	�1��Y����#k�x�+�4$72�g�dA�N��7@�W}J2�m����vT�Q\�z˪�� �da59���l�H$W!��cK�z��`8���#�(�_]X��m����V	�b�#��V�4����"�"M{;U� O��8�x37��aFZ�m���p���N�w���ь2��B�~�[s����U�Lމͨ�=��
,t�q��6�i�v��7�uc��it(���.��F\���+`ݑ�]ÜT�+��M��s�27����w^��p�,|s�q!X�Yi(4K��^A?����Y;�^�����.ё��ʚ�.qY���Z��"T��!����(���z�'�����k���9ujRw�9��3i趻U��9��7b��V�V5��W�֪�o���q�na}.X}�QZ��SPp�;���4�0�#
��,NM����U#��|ͪqT(�vd�/`R�佭W�ā��k�|1��OU���yL�W�
~��X�1�!I��Gڏ��^��]Ԋt"�h�Y"���x���W�sX���{#b���z�^Twg�r:?�0)��i���ҷG`�f�HȄk��f%iM�9?��F�)��gV�J>v4��H��c���~�S_��ȝ5���}�x�g�m��Y��t��44@\\kր�`��� E�]�֟��JN��W�h��ɜV;��Lқf=�|qZ��P��t���X{���,\���O0O�CR��=�ؙ� ��ɪ������	�&����z�3o�� FE���$�G�f���oE��n�����**J������.�1��֧Q<��$�z� ό�Q�Y�W�U)��fʘE��.�j���2��6��˻ǌ���N��xpsY�*��ϰ�Z]��)¡=ە�[�iӧ�=C�,��k�bo^F��쏧^�i���xz������=il��|����D��(� �yYbZS���OE�1R
�g��T�[���@�ȕ�N)��3Dә3P"� bA_�u������k�q����n�eD�����s�m���;n.b�g�N� �����#��
��P�:<W�onX0	TR��Ѧ��`�7d�nG��@�'��PAk��y��^pc��ٵ|�0g�ˊ��H*O�O!{�))���	�1jw9Ps�1������!j�I��@��
�^�6Z2)�����yJ�j@1�%�A�q�C}1�yO"/�����M��,:��$v����Є�^,��E47K����7���Q)���l���l�[3� 0�
�\")U�m���̛:)b�_Y3c���Fmd_֖��:#���R�ƏރT%�?7���PG�y|a��.��^��3�˨ܨt��-Zr��)�n�\7���P�NTu:cdS�������]�9�BЕ��6yO�}4%��H}}bܛϔG�4!$�vB��O�|�V�ҭ�`���(mi!���|�C��VSgW�#��j���7U�z��Mwc>��N�۶�D!S�V�����1�7�`L9�}(s��ts��'�]��u�js����"T���~B Ѹe�m�]
���qݮxr�Ҵ9��Ÿ�7Y(z�6��P�/A�i�)���u&L����zf�B!U"�xw@`�ެ�˧`���^���A  (��B=jTK�~t�5��ɿs����77B��:�����9��2N�Sj$ޤ��
�f�QVR
n�Ɔx�J��{g_��/�¶�x����p�<aӝ�g����P�XQ�����yr���-��ݗ^a����|b��+c�֏�ċ�4��T�ǺxF(���&�7�qL왟�2�'hӹ~��(��ya���)*B�������]wud��}��N�4����\�g�^��+���[Qj.<�[�*�IR�p�h�S����`�vs����m�yd�LI�ԛ�㥙|@B�;K	b`�.��^s|�}v��O��*��]G"a�j�HS�u�����tY7�MX$����"�`ʨ��$ls�V����r)1� ��L�ڮy���hL�M�*���zJٷCօW���d)�vx����V)A���TzfK���s����<����8��%t�(��*�y�Fd�c�����&$s�0W�z����cC��5dL����F�,^���}0߭d��U�٩���ZN�HYI1��:���0U���`p���
H�����g(������TIHӠ*�?d4C���������f�' �ә�c��_�s�=�2[�(M��҆��;��7�
|��f��⻞�?�^�H"�t)���x�=I�L5�r�Qn���Y&f�2�w�-G��K\�n��mH��'�3�j7e_��K孢vj�nՃ`@�Γ�{�c��JI(�ø�Y)y�黚n��%�&�F ����$gɮ��Q��2!55yU_�R�����CnP�F6!l�]���N���ho㺱ߙ鉢��1�~�޻��7��=���CF���ť� E�4^n�&��C�-�jy�2�~	I��)&����bSpy�H��ǆ\V��U$��4��U�~�O����Ka�}�4�,ֿ:˨JB��+n_�uv�&�Jm<��`8��wi @�
̢͈$.h��~2�}O�R=���S��6A@E{��_��!2G�����V�1D��ЄP���3�5��l/+���SP����l.��N����^x�d��w�_�LOԊ����Z�R�nzU>��hXYr��-���C�V�������1��{ݓ�O5ۻ��κ!B W7�����V�'��G=�H˽Fy�x�cn�N�sz7L]�\�(�L*�}�򄶾�� �����i��^sG8��\ql׼}��C�y�)�5���w�+�اpX�s��l�������ҡ6�BS�-_�_���Ɇy�W^w懰��l�^c-�D%��ř܄$u�kɼ��,g�Vgc5��&�I�ƽƯYAJ�X��=E�V�e�T�ж�S�`ܢ�;�\Һ���f/�B��� vh	��"T���D���S=�#�$)�۔��̫�]K���+V(��^;Wqc�yRL.6��a�}���9 �,��K�
N5~�z��Xj
4�p��e�>���$ $T�sVHy�&�2^#���~_ٜj�����!K�׺�W�=��םi�(������v�Ԯ چm"?�؆�\�p�/���3b�t��R�U�Ȥ߮[h���^{�KM\'�]yw�S�+��r���mJ�ߣ�]��bm��1w� 8b��h�k��}��#fY�Dnur!	�ψ�����K!��Bmtg�N� ��0(�z����8T��/��'P������щ��"��b.rm�.Ί��:t�͗Ù Uܚ�2	c�����B@����=Z��$<���֛h>ޥV� �f}5�v�=j��CP�����¿��O٭"��s#P�������׮�U^�}{	<쭜/�p������)S����Ki����]�6#G8��t:��y��Z�_ߔ�s�O��W�j���5|p;j�|\yb��$�V�(\���������b���uϔa�Z�u�^��PG՗WV��&9*�pO@��m,�JM��+�F���N�8��#����h���52b$]!{u�®�U�����k�S��i
��&�%���P�9���0�`H���!k��w'���*Ul҂�iQRh��xG�.T��j��jJ$% �cL�ʻ��m�����&R�G��ץi���%}d�������[���p]�N7�|��
?l�W�'��C݀?60��<���*:\|@����?��xSR�VvG�U���84�OKǫh��T�m7zN����$�u��g[����8��#Z�LN���zXi�g�OR��U��<����>Z��A���EL| ��nzHa��٤g�~���] ��cz����Odj�/:b*�^��]6{ʷ�F����"V�!G�WW�m�7[8��/4��]��'�Oy�)�=>���wM_gxo[F�C�d�A��ϼ�����+ɫb�xX9V���%5����z
�P���+[%6 I�D�.��4#~fɣ�h���/�O��P��s�-�h��z��_oX��0�Ť�z��9���8_���& 7Էc�����=�{,V��,�T���l��f�o�n627��+�>����Y��J���<�=؉�{r�����^rO�B�%ζ[DUkt�t n�p.�h��t�߀���U?e%9>c��3����0@�����9�gN���Z�qw��B�6�8+�>�i4u��*[*f^�B"��+����!U��`Е"�o��2��m�r�J�#�FU ��^������(����Yl'�Yń�F�<@ϡ/O	�%��rqJ�v"i�̊�6L�)���g�p���9���v����6��K��4׊�<,�򫳘~��tD���VS ���	NF����� 7��]p��7˓����Q]#�Wb�bq֘�h)Mk
;���䘞S$�c=�������2����L�c�1f���'��+\�+��k�2��/���Q���X��|�
��7��X��W�.�N�@�Բɫ�.y}cٜ�4`�Wݝ�PB�d*3��3H���g*�D1�d���;qX�]�m�a�o�g�޹�s���ۊ�8�ܥ���J��㠢n]uϪ�{ů�@�~{���/=ʹ��%�5���n#��LX����k��#!%�af�)��ӶB�Oq�M�<rA���Y��� 4����j#��f��@�Qh�$yH���O~�{2��M�=8%�?d��ٮ�,"K�*�1��)H�S��՚�јaBO��l�7M�c*X��g�����g[�%��B�>��uB�B�{o�B�w'��X�b�9Ҷ�c�����8�r�o�Ƽ�z�v���Ej���<Z�Eѐ:���\�T?@&�TU\쵄	]�V��ſ!���FR>�ࠤ��_���ZAA��Ɵɚ�����"$�[�{}�M�IaƗ܎VQ�	x9�8��Vf�#cѝ�B\+�������觽o �@|g4L��6�R�]oO�J
��zO��P��ڒ��]f}��5�n^��4@�՗�����_>v���lD�뮐�[S���co�a�h&p n�a;�����Ed>d��� ����������*/��>e��}��C�VJL�� �3c�-@�tc��c´������������e*\��V�����H8��a�W�����H2&$Wǁr�#�Jq��/��'�j�0�2���ĶI��Jk��I�8��7������,&���X��!)K|y	`�M��wW�J�(��\���@�2��d�
I�|[�^9%�� ���1��i�P)�F7�P9	������O� ��VfS]R+��ZhϜ�§�b�T:���.�z ��e)hi�X0f�;�R�"|?����c�l�\߈�yTѩ���-��q��e�Ɩ�x��(A��-D�I�G�b��=������K���:�)_�Ԟdg_�A5@Di�������I�@������1�%��������k�l�A��d���}�o�l��6�j��ן��O�|�f4"�ʬ��Oȟ�9q�_]6���Z���N�Z����M�����M�O��d��'��j��T��Ҫ}�.�w���f���۾(�{w��}��kR�|��j�}����'(�5b C=�ф���S�iɦ��ꦅX�:�5~��B��4��Kl�x� ��m/�pK����p��s[b��k����uF&��`�R��K�y�.�y>5%�td���;�3���L�L/���(?q+���&�'�5�=l���oF�nx̲}�ܜ6���JCl�R(�����m���8P�P��L���[��Psn�E�H$�H��:�20��w��[E�D�mk�g���T2��Z�O����\���g��{�)0a��/���坔��5���i��Ȑ��.��v�-'�]N/r��Ό���ӛ�h��-�# 6�J��Q�Y�;~Q]׆_xI�����;�s�pXkm����D���-�e��%�b���w��z�1ΉK$�.�5���c��C�,<H���cg�]�h;�j]�p�?]A�:���J���[���[�q,/a���5�cnN�7���c�!��7���UO�?�-�z5�M�Y�$�.G��7][���̏�@�V[�҉Hvgx������#K�����3^��u��F0Y�ۣ��}$���S�@�=�쳝�3Е��T1�L�R�����Z�-@�|�h_D����;羜~u�[�Y�d8���~y��kFۭ�D����|��$޼��]G:
���;�0�{��7�O�� J.<�HQo�aa">z4���7����t^���h�Vjz5�_	�BA���]��vT�<�qR�:!�G�G�=�p��̟�U�Acb�8Uy�5һoG"�J"�(�g��It2ޗ��LM�Y��ҙ�Y�G��������,PI��轶["��R�q,����vgoN�s��I�,K�!gt
(D'�a��BO��~`���=�.�2��d�]��&�4,2D�"�,��WԖ6�2�5��a�3�+��`�A���Ns!�@��F�����<g���m����*����7)�<���vت\�5y�Ϲ%��,=����ǳ���{<I����] ��Q�2W��蹢l�1�"N�c��s<?�d�B�<�rK����9-���v��ʶ"�é���+��˓ɏ:��lE�E��g1P���������^�����W/�gT̘����-w�6�f�<������'���%S7�����`O�E>��t������HE��q��!�p�q7���0� �q�&����vW3o���|�nV|b�����'P�'�b�2ᢨh��J�A��M��oH5}~ٚ)�0gt�>����������~���|&E�X��SF����핵���]ɴFj:\=,�M�G�V?G=.�D�[�@���KQ|y7��٪#EȷRֻ�I=�-L�W��W� �[YwБ+t?D?l6F�o�P����p<C8Z�a�,'N��Ezk:NC�Z�X�N7��<QBp_^G�ŀ6d�|�R��L����\K"�-�	��S�7���w�썐1����"k��>nA��I��"����l�p������ߛ}��e�9�J	6�uM���������z�z�R���ݿ!NI�aM�M�H�Zn��q^o���=x�!��$�����xbn�:�튑De�_iE�bY��F/�	�ȩ#�b���u��r�\���U�;h�e��굾�0�f��w�����"]G�h �`� ����n2�}����ǲ�|K/��:�o�b85	�E.-�|��sa�J��'�]��9�iJf�p{`�E��T"W�Pq(��b[�9�)�U(U�I\H�=���>�F����<�hS;����������Q�q�ï��V�o]�V�k�vk��'�tOO��-�@��?���]�#�ֻ�D��;ׁX+Q>\����E]3N�n�g��Z�x���b�|^>�� 0R���z�/vT��F��+�?:��'Q�[���I:n��$����Up�c��U�Q�%��B�V���ڨYt��*���ѥ8�5�Gh-P��[FY����Yb'㹜HNX1���Qi=�^6� s!a�/!�Fu�����2�U�Ľ��T�9�f2����TG�x�z `� #�X�/MQo�w+��p�`hF�e���0�~΢4ʆ�d��B�bU��	5�@��;���l�����sҼ�$�wDf���r&���`���V����ʺM��d�� �®�w�Yi�mLs�MR����hA�^�q���_5�^W_c�oF7�Bu'v��|B׾0$�gL�E�(Z���4Hɋ'Pl��7l�b�:1h��t�U<�1��f��{��$(x.;�fk���uT��G��}��~��5V�Y�11�z����i@"��rtl�d� ��k(<Ң}4cN^kS��F,�G����-j�=����g��,e�(!j'"�:<_Y��|h8�������ug���(���P�nһ�� f�SAJ'$D�����)K[�(o�[16��t��c���`���eD+C�Sa�,��Hq۫�/�k��irǙl/���g��I�?$�~^�S�a�:I�����[�J��ƭy��ҁ���-WS�0�$)*�����ϩ�8}ie;���5���/�.��E}E*�����}�=G��N��;��RP�9���]p��jY7s�-�T�Đ�/����b�0� lzC1y$����4$^��������MP��t��t�� x��+(H�����A����j�-��ٮ�	��'�Dբ��\��r������a��p
T!v]}�\m�!jm�K��u�s�.�[-��?f��ō��/Vd|+��j��V���U�S�6��<<��pz��B���ެ���!�}<}e�S�`���+i�&=�*fV������R���g��k �����C����F�t.�rB��*E^j5%�;#�_]�������a��D�;���nM���:�GR���Bc�#'����Z+�=q�8���4�溓Jm�:��VA�����*�y�X!�����|�������6�Ǫ��Wa� j\&,��ө\�9�O=:���\5�.X�'�;ʔNQc%9���j�aǞ�N��k��ORI�o��G�b��*���Meu���It��-��q1���Uj'Jx�!�fo.+l'�@�S�Z�J������'����cs�YX�3_�+���|��n�LYx\�wՃ	�*aTxyk��'�Jm��u�*�]�`?� i4k���}WS�G���sf[j����a��їI�� ����Y�.d5�;���۰�~��0v<�k����� ?��� ��z)A�R\�;�2��hrU�6�����M#G��<��_�&'� �8�d,a�nm� ̱f���2w{�*!s ��7��NT���
tش�� ��X?4쥋�[��nk��}F������Β�8 u �x4�D��c�p�ݞ�&'��	L#�YV�o�j����s�Oes<.�ѥ ~���fR�3�it�������I�k8(n��ض���w.t�t���i|ٝ���/5����6~'�R)Bʂ�S���~����氚e�?��f�:��q*1�k�C4�R�-���jƠl�p�|YT�!9q&G�l]�����ekM�j/�Rw���˾}�p��̒lJI͆��B��pr�/�{���(��U��� ��a.�'�G3�b��A7��1�@X��7O�w���M�K{�b$H�������|��G7��9"Ҫ�Z7_�L�)V��&���%%�A��h�li�}}�����. �����v�x���s��7q6:�E�z3리�J/���|�-��Vc�ڟIUV�����ݎ��ࣰ@\i焁E`/6ē�~��u��o�f\�
	b��3NK��������k�c��y��7�$��]�.]NG� ���Z=ܾ��R-C��Z~ý$�E���vE�`�D���(�;LJ�Mې�O�V��$�~G�6"6���cWw�x�3�|B:)��/�ƀ�2^`�=�<�Y��V�������8�7�q�砘CWT��V���ݞ>�Tq<`7����i����dC�t}n(�~�6بM	����1�2�b�Z�(���x`,�@/��n �31�������T�����z��k".��k��
qč����q;�N�j����ꑝ�k's+�0��/�JX^YUcF5��ƾ^�I���;ـD5E,9?)�r׍�1��͕h�i�F�"&�kX��wm0�	Лg+r[:�q-����_u�YL�YfO����)6@�b����N���7ob��I�kz�,�9g�^��_�.<ch��	ick��Z�2r��U�)zw�!a��,/c�f�Z�E�IB�y����ŝߒJ[G㞆����K���4���3�y^\�A�5&��!�b�f�a �S�^&�&��£��0��Vʲ�~l�ڿ><n�n���jB�
�\�:��Q<m��@�Ys�oт\�WՁ�#b#�|�'~b���%B�ߛ���-x���	K�{H��u2ږ��n�-Ŗ�%4�9��խCqnG༎�[����`�x(Ǆ�"PN�L���̶��L��{�h�7̇��_����$@Q�&ꂜ���!���zO9��:� ����A�* ��@<�	��-��j��{B�+��ƛ��-�/����ܿx�=��[}�!58���ʼEZ���QB��D��޵ʟeCI�Ƚ�[m���(X.m�E���NLA�I��`�\�hhXh��N�E&��ά\��4��۳87�W�UN|c��&u�!ȁ�*$qPr���"�������VA�o[��LP4��KA	7jd�o���h���{��8����ݷ�D�fT��i�rʮo�@j
�<M��V�&D�]�~���=�|�ͼ�p�9ƨ!P|�����GCp�������ɴ�&�� ��<q�C�t-�%�+�K`�h־�bq��M508WF^o���MQw.	W��8��=�/Aj���'��[!�
q#�H�GÖ)^N����9F?�{��,�a�����r����TP)r8`n,��F�4Z�]!�6�:S��5�T��-J������$�QE��lc>*�Q
7�%�_�	��&2�G+f20���9���q��B�b�U�{훝΄�h��½�HD�
�ȌLFz�݌I��6`�ͩ+���eu3����ۉ�ck_�Oڭy�APLr�&��f�ڲ:G�0���,5|�B�<,y��;�Z,��N ���G��ЍT�?#�f����k��FQ�J���gtbjӯ�'OWC����g���< =�_�R�;.d�΅u������I9�h6�ai��%������#��j��4p���q�w?�@�<���!�K�9����yàɕ�f��:�g�W��ǧi�	�?��Y��V�V�%�¡n���*]P�bz�0��S̱��\�5R�~������x����!����_�����"l]/+�9svfmHE�}�7h9=e�{|�/R���x>-��eI!����������G}9E��[����]������se_�>%#������lo�Iy����{;r��R�^��CL�A6�ǙV�A�{���|�:-ۓ�&����㢊b/����i�p��<��ç:��}�)�*��xP���'��2\=�u��9�P��w�a�?���n}
6�!3O����K�Q�cN��4�`N��h�0;iC.��AC.�v�<�t��=��n
M�a�Y��~<nPFli=�/�PA��'�Z�w��8�~h�dc�v]�̺Df�$b�� �r@
�ˏ>�py�"���N�ޅ�.���=c�f�Q�tє� s#�Ӊ+񄗅���U��9H�2���"�.�.O�`�� n�ݹ��f_�:w�[˚#���"��N��aM��Ig���}�Wb���_JMYN����q���	��EA\�r$���6�(�뽬q6��?���K�F�fE3tڐ����ݘ��p�a�8�{G�Љ6�����Z	�� :z9=��@GQwG����U���lb��J��ǈ�8�z�z�圅���.�pZ�8�ٛ�˽14��0)ZH���"�E���"p�9�\�-�qd�mY� �u��fר"4t�$w��o�֓�≶V|&`4�����;��ǚ���l��*	w^���y��5&��S<{�8�p+P��]ҿcݠ���i�<�؆�-ʫ����D����fs@N
�������}5�m�E�=YGO�.c%Ū��N���@ev�0�4����Pw;�D�˖����ǂ��#S��Oz~�& /����C*��h�}����]&�5=7!o��XY�)3 [psؓ��f�El�n�"�q��S9�����ҔʖZ�Aoױ �A���l�Tk�]ŷ�x�(��)mZK��uG�8�6?�� N��N���|#F.���P�a��;@���4�������4@@xm����H�H������Ϥ �'�z�k�A��ρ�h��&�{��V��Y{%��t C��B�݀�#I=�~4����)gܯ�9��כj \�s�s����_%6.�0mn��AJ����9EǼ�>�b�;���^������#�����o�Qq��\�H�&a*��3'�LPU5MM���nEoN m�_Y�g�`���&n�3�|!�_({7�P@}XBn���$7�a	p=�Q��f����ѣ���t��>&���&�3�au;�x�pGbȦ��2ik|�%=��v֮�y)cאk���d%�E;�R#K�>�0Sڕ���0�g]
��M�6��
,�u2�憽����2h���8��<�?���!7��93���|ExTOL���Mj)��ↆ�LA�u�r��z\���MG���'t�79H���X�KP���VB���y$y��x�#��v��l2p��G6P���Tm	���u�ā�S��A=4�����Ex����3D�Ҏ7z���g,3�K�\�&S�M}?�Z�tv�0�w>�;6+I�]=�_�Z�"��!�܅��~��� �[c!��+�Z�6˿�@:_
�P>H���O�>����k�������#�r|L2I�˕ZK
�{�K�N���A���0��d����ڏ�,�-iZDrO�Ҹ�U'�n�ф��\�z{h�p[������ |�`����������ZF�7���兠#H��иR$	"����=�7ĳ+��d��a�+-�v>��vw��xi���65
ii[ZYMI��?�v�"�=���g��)��Gؔ��<6�YW�|��o#���O�l�lJ�X�pQ�o��5;�J�{�<�-1A�]0#3� ����C��M݇GS�Tz��JmN
��ٜe�Q��@r�3�c���v{�S�]�n�+�I7-r晐�kt�u27���Z���2��}�ȫd��]#7�wm���5����D6���l�t�Ƨ�����G�j�P�k��о�r���!�s�&L���t�'����RT�˯=��T��/�U�����9f��O��P�jl}M��PN�[�&hR
W� b�k9�y]T�M������]�X���U�ҭ&�&��.��D�̿�{�㒭���g��"���7�47�"-����}Tg֤�w���X恧�y.	
T������.�[wV������7|���{�k�������GH��G�O	���E+Q�v��A�[��c�P���co��[�T�q�h>�b1W��: �-��H^��!���37hr���΁9�!�J&v�J�ae�����=͗���k��mhx�ti�ׇ���W�p+D���P��H��7	��0���%@�kr)�g���R���~���@��T�.��~ܱ*��;��d�A�*����.���s`��R���x�	׾�:[�ZS#����1��Y����sҌ�z��F�a�ױ譂ĥ]@�����,�i�5s��T�yU�+�
��|��?	���K�&�
����y��Իڧ'H\���U���U�0^���z���O���Ӭ����o���*�+$�'?�D�'Ӱ/���<�"L#���(�?ɞ�sR��I��K(ʓ���a��Ng���6 ㄢ��B����X�M��"��?��)�,8��f�O�_,�K��]-[^�h�h>%������¿����~��a�vѮ5S�����U�}��w�)!*MUE��+����]��&
��]�ԡ�z�_�̍�G��-�7��������[�#m�ۓ�̟�[�]q�N~ا^jw������}��vP��$�}��_���1xM:e�Xc��2b3)GО�Q$2�A�ƓU���9F8�5�\2r^.��[W��O�����?�y�%Q�v<��N�R{��v�m;����)�<y"�L���bm�cY�:�hd�D��"�/e>�kI�T��:� ���S2���*��j?�o_.yQ�>	w,O���I�G��f��~�c�n�T��p�m�NQ��-VRv9?�P*��VY$�}�y�����ڱ{w����S�$\�U��b�*]cX0'J����R�����9Dѽ��v��쥛qe�FZ����Ѕ���oɀ���0l�D{U�]�i�g��1����F�^b��e4s⒬�u��,�Nͷ��j�"�*p�	ʽt���Ž������ψ�w6�1� �����BxC�QC�WUE�d1C1�`)��z��Ѐ�ƌ���P����Lé{r@��&g�0˔�J�[�mf�qXhT=�����g�u���Ϗ/���R`�����A���J��b�_t�HD�3�����b�G��#��P��
�*�";; A��5Ϸw�>��c������;�����)-���-;�u��Rw�Z~��%�8�#��R&ťH����Q���G� +��n��S\�!�Ҫ�сc�x��HǞVT��sY+N����*��Y]�
G�C{p�Z�@'���c
t��d�z�N� ��k�r4���S��ߖ�ʪ)�={��8�HD\x�n:p�%\ϊq��H���*F;֤7�@�T�(��W�29��OW�G��8����1��R��爠��-X��ٲ���}/
e
���!�wU��A�d-��k�!��"蟘	�m����&F#8N�
-���`Û���	���O���Ι�� ��^ގ��j�KG@Ay}g8@4�����_�^+���|�O��T���j�q��A�R��o6��/|h�	�R�{��ٲe����hD�u=�)�Qޅ1x�qC��������j�m_0���J1�����,%�쯥� gv����]�o'{��ҟl(Q�(��y&3a���]���=%ںZ{�Ѽ)45��C��LwDVN��ݑ8F���S����(�q�ψ��q$x:�pvWY�ڿ�w��H�"�{�HRS�ޕOG�)�.��"8��sn_Ӓ!9��q����z��Ete'�),�T�PbɊ�Fc+�f��{r��x���C��U���̖u�B�W�i�<�3���1������e�c�H���ˣj��<��6��)�*�^��K�Kr �nƁVzƑگ���w���!=���H���3҉zN����B�v��ġn��q�a���>F�5���:��R�Vj_���wZ����g8Y�N�pġ9�a��@�D}�=ZH��a���9��E��\4�&߻HI=2uBS}5)�g��]?�}��Ӊ�!���,�b.�\�>�)�ߒê6@̦�L�z4w�a�̩}L�heҊ�˻:�aR��7��hL����Pz���A���2��i�<��h�Ѻs4}�A�*���8m~�KM�]Q�4Xd�K@7�u��؆@��:g������R;j0�0���D�Hs̑����4���D}l[^���F�?�iz VU�:�0v��w:���,��2���� ѧ��ш�"�}�2�(^q�p���ܽ+x'Z���lF�����}�Q�&+4Q���q�[�C���^��>dͬ�/V��ъVN���Z���|��$͊U�ԲB�CNܧ�g�$l��i׶���� ��G5?�V�M���}����0�*Sb^@^��3���&]4LO�wK�p����D�T�k�.�� v3bө�хG�+�M��P�J���t�i>w껓Z��ѽ��2�MO�Ӵ?�n��k�E�A��h��-���߁�'u�#��;5_`��-��	�jk(@��cr��"k���IR*�����d)���3(��;��j]b�!���/C��OsWjS���d�Թv��<�Q_$�� ��E��QΥ�h���2�=͙��v�I��`qP�*����RB�-f֑qgy�Y� �.d� h)O�,�"���Y.o�k_"��=n@Oa!k/�{���ƃX�w�D�?�Aykh��r�1G�[k�T���f��/�����s�)L�?�8GT���:�D�-���X�w����;��r����(Pf
�m�Q�k9��0DQJ��8��WV5¤ ��H��`�G�9b7s�2Z���ܬ�PZ���	9�~�v��k������g��f�%��~��cN�r��;p's�kQ'7�R�ڳ$݇_p��3�6Y~�~v�D*@�d����[ �~J=B�̕�e!��rZ�9t�,DE�f��n���Qu�l��U�-#ȇ	�
�3�݁���?T�$`Q�K��7�8����o��!��hVNA_�[g����N 1S2���KN@��9��;��u���D��K#Z-�qݘ�.�(��^F�.e�\'B�4�'�y�^+�y�~�&��C<�l����u[oRcV�b�΁��J;���P\}�H�Ї}��Vi��N�M(qF~��l
�L�h}�G�����E�/����f��R&�w�����Q��1e���/بS�oq׎�x���i� 6(���y�F���7��)��!�S �zF�_E�g���f����t!�eȡ|G_|�Q����f�BY2?�4^�6�_H�e
���.��N��Z�fêѱLל	�z�=�p:X[��MQŉ�g;�m��{�"z�T�
�?_�@��g��F#���T?~`��4�I�;���uA���8l`,��*q��_؋r-|��\�+��%�j)|
�B�`���96&=?�ġ�?�k�%���Yo�B��6S|�*.��%|�a��@n�"�~V����Fk�WE�'�b!nb�����_�C�rL�(l�<�0�0�v�C�;r��'�X�B!Y54BpO��<��י�5X�ͩ:3[r�R�58��.�J�����@a�TM�+����
*)�|AI�&��ޠDp�l��n�?w����<���%���B�Y�a"p�n0���,ݻ^�qJ\�Ʒ�&��'�vtk�����EX7ԡ4@��״0B9�����(�UI R	�:��`�z�P�S�Y��V���Ϻ\�h�0���|KF��=->����+I�TuV��i�1���#��ģ��ldk>h��iC)>e~�C�8H�U�^��������$��1�
P�w)ْ�.�r����ә�@�]xSf�A/lAF@�<d��9�~E�4 e��Eɬ�{�-w�q�� �R��H��y�����Q�����DM����T�Ƈm\w��q����0\��H��Ow~3� ��[�8�M�?bk�/�E=���<��?����)�mſ�ߐ��b�J[��3?��M��x�"�K �A�<M~'<7,�q�n�?�=��K�����
�"������_�nl��޺;.G�1`�k�WP����K�J�7�*����ǱQ���l/�0�?Pz�e�|Y���}�#L��3riZ�Z?�xCdԑ>齽>M�pX5�v'�T(N�P�x��Y���3��J5��]�<�wb�Ĕye	�P�HN�����S��(�&�$f<�I�©#���J:p|j��BY�m���-qq�l��V޼1���?d��ZL�<��>�~�Sc�M��`�cK0.����i!0��1&¶(7�`	6v�����'�q|�%H]fE�4�OM�k���ذ��E�_��M����+9�%̪%�#4������j��b��Aw����.�Ϩ���$�b�Zє����.Z�i�z���%���,�o6̋�0���C�1�ӂ!����l�U�E��/�*e�������~{+�C�Z�<w7��t~wH���A5��x���`1�U�#�������x�P���vR�Js��M�,&��?�5��q�R�ր ]psv�Mö׵�"�{�1�D�W�6[w����"���.��{�` ̨q�%������l�yB?�>;�~^ӂt*!QM�=���^v#�]Gr/�Ń�:9.?�J���M/�$��4��
��u�D�Ƚsu�P�C��eY�`�\:���e�K}��������<a�f������\�0x�G{��K��/J�mŋ���S�k�;��$S��"�\�ʿ�h��&����xfG���8����R21��S	U��
vFW��[�ֵCr?��uwi���5P��űx;���G{TB�U��C��^�O
Ti۟��qC������T����G��b�k��5�<��t�����p��7���ba��х|�|��0�P����7�e܍b6D'��]�*�i���k[A���~MnVc����DiV*R%�-���l��66��V��,����f��+;[(%[�n����K��AC�;2�v����s�K�h4r.*��g�P�I]��!9�y;���0t
%f�؆3�+T-��h�z�`�3ό�Z`qhcG�q���J�ɲ4��B�^�p቉@N7fZP
��m�K�%!|�3�+6��M!\�#�
3��"e 91�>w���C_�=�7E��C?�hğf ����-��Z�juӳ0M��rD�4���%�u�niR�1��+ Z��4oG���w�m����;�q�s[�jH�t2J���N���Ǜ�_���ܮ��"���Z���N:��2~�[��Tm�dt�[�D�3&u_t�>c���2�?�*���$30�7�i�v����!�R~����+�!Ŋj)����(� W�,�]&r6}��EU��z���޴�|��' H��!����h�[+Jvx����],^U��p�΋L}���}��m�����aT҄V�pk�G�V��n��%���I���$�ټժ.:���I���*њۯ�ċ��,�:���(Q�U�N�ҭ�M��J�"};1J��m/#v�Ј*xƖʓ��;�C�&#J'�\�%��5w��U���H����pH�����
�z%�W������9��<��Y��֖$�V �o��M߲@�∺��>_��<�kB���� �8sU�P`�&[Uu�3�{<�����T�!J񞆆:���W	��&b�8��-��l� �)*����&1�JY]�ϑoF۹+���"5;�r�1��P�9wcl5�rkF��E����*{�$�ݒ�a���Z���qQ��{bg$*��J;:��)	�,�wɈ?_-��
���u���tN�X�s4�� �4h��l��G׷�Ip�u�Zs8��QJ�r�	���� �b U�%�i������E��`!MqL�o�9(%�=�J��+J���1Ħ�kp1�d�\y�<�羶D:6��w��b�W�Ku!�G��_�l_��F�v��ܔ�BI?zu��4�V�;��.�����{�6ғ��s-��o����Q���r�6���l���.z8��`�F�eЃ�J�-N]e�<���+��6��07���_~>qֻ�{�2ĵ�srv���岇��qeU��iwE�nx���,A5J�ϵ�G}J��,���>�3�I��-�N�L��ݡzy�H�^Y�AF���OH�m���k�>y��޴5WT ��/���cR��&�YT�vA�M�8W8J13��p���a��1�U���3�[��j��NTDD��T�2�)�{Nt^?����N!�wn��g��eGA�@��'GDe�RKQk�,\�X�ٻ+��x���_��nQN�(��4�ѐ1�F�0�����`���Ap�2�76�cH�z���-M�~2^����6�!�=-�N1z��z!h���gg[J�O3�V�O��پ��Y��F� ����Ƌ�֙0�dA���9p�~��LN��g��d����K��4��w���vHZX��tNO�1�Ц�J��t��,�T�g��У�vPl�^���|��o��H�b����!X�>�l2���=��.���Jz��'M�������s�<�M��~�.I����G4t*��@M�����A��5�?�ZȫXp�Dծ�����J�Ʒ�5,�NS���w�J���os{%�?�8��Z� ._#L�����nޝ�E��Z8ʲtĆ�,�@�0/Pb��l�y������6���+n>���
x�b}7g,X
冚���7DvX�o��߆�_q+`�BR�y��@��$������P��VQ�
9�mR���"���{��mO*dq�����"0�ؙ=�uOB,�I\~  �x��kJ� �?+�(��=i��CA���`���t�7�j�����D�&�+W/rT�v$Aĳ=#��0�?��~�Y'���+c�)���v���Y��qj��7-P�G����?�uP���=d��Ws~�q#�z�z�[U܄u����� w���4��hj����Pk�뚌*H%���-��M��U0k��l�5%OXC��K�]9�S��;�Xg��ڼ���åU��#�z���g�UQE"�ҵRai�w~}�:ߔdq>�F�4�V/5`�8[��3Փ��GDu��*Jc��w����rE�/E�qY�����|�*!���=�^�c��mF�*�hz���+����m�~����b��L���˷�LO�����
����J�6 �����<�Q�$u�iT�\���m��ǎ=�l\�1$lZ�G5w���T��O�X�$��
�=��Q��EF�GkW��t��r�
��U��F=�]�h�ܡ�S�|�%���^5�و[Ϯx���|J~�%9��M�n�Ǌ�olB���g�s��<h:Q�4��;�}Al'Yu;�?rsJ/����:/������Q�zo�/4�8��-�3~#��4s����)��ٳ�
깍'�ͯ.�xg/�� ���|�.�v���0�A�o�}��K��A��&�Ŝ��`7�36o�=�.{��^C*�0p
F~TB�Y�m�Yᨀ�5�m+�#��«���K�e�(@��jv:�)O<����m�؍���:���{�9����~�$>r�$Xu ���M	~�иJY���'F(pz��A��k��uVPL�O
(a���=����+G=���OkX�gr�<��N~�lR��q���ɶ��1U� �=Ĕ�Kи����qxV~��@����N�H��RYO- �X���-�D2��펚�Ğ�N��q�?�� -�����ǒ ƃA����a�i�Y�$�t��m���zp>�ɪ*�V��]M�z�M��|���9�T_��N~o�z��q�U9�])��%Fpm�,��/���������X���D���:�X��M,i���U�B�>�-!����sf��,���h���4��=��Dٙ�&�!q֐ W���Q
e.��3¯Y��JB��%��z��V���� ͔�P����Q.`�CFFZ\M�9���Pt�ܙ�ʄ3e(�ɝA�.4��q�EI�@`�D�	����@�uK_Ӵr�f��/+���)�͊>JH�0D��@�@3D'���Qk��������!Ps-�F����-�>	s�&�/S�L�Ӣw�mt��vW)�9�	JjC��d�%� M�,�8��Sa���,�y�)�eU�����Η����Y�I���N��^�� �r��\�t�q�;
�[�b�KO��l@q�}1��ؾQ���U�Ͽ$�<z{��k�ez��V��mfjx���kO��g�hmpT�[-��_~;)�+�6� �;zp_>��HC����
� �PI���!�=�o(�6� �(;^��� a'#�>�ឩY�%�H����Ư�t�#�3�2��[mQ�Ĥ�U��&$-O�E��ҿAi�M���SVjn�A��J�����\�|8�a��%��z�e�qq���A<X�ԭH�rT��=�1�O���� ~z�z
^'�u����"���N�೘x���� m�ZH�>a��L&C�(���z�n���V�r�c~D��-�5'&J����ãK� �u�%ѡ7h,�j�iU*�[��Z[��4�5��Y	k�*��'Ǖ�c���
��&�$9�_�N$��Hg��T�����f�ZK�.`�{Z[>V�B��Ϫ�J+Gjs>��PdH��Aw����}����x�7'�,E?�Q���M�G���]� �����<l����'6� g��Ћ�Կ��"�!1�T���/�TJBd��J���V��|��K.�$'����*��J��l�8K��d��_r9�nָI=�bT�~�r���m}��,�/i}��i�����M��`�v�B��Y��俢�]r
�L�g\킷��s�brS�vhgz�Ω���� .�ˈL�v���������x�]>�3
.�y����(��b�%#�氩�g�W�+�悎1�	�O���6�ɳ8( �R��.�oi��S�.Y�@r��@����PW��%
�f�)�W���lz�-�F׳�O5g&�4End�Y,F�2lh�%T�����F'�֫HF�I
�H`�ZI��cI�GOŁ�f���lN_O8�J�t��n�D|
uĈ����_��Dgjrh���l�BF(�@g[Tw{k�7���j�5d?��P�B�Yd8��66+���Sb�緆���Xݶ~>��V��� J�I��uL� 0��������O�}hb��=���B�<�O��ѽ1��{eo�����灱��4��E�y?d�$��0݅�:�S�;|ht͚辛����d�˛]��(-�QDJ�k��8��(�','�*�X=l�<�'W����'�t�э�Stac��r��!!
+M�FA�VHt�5ȳ��RX����oE��˽����y|16�K����>�]c�!�K�$�h���PT����`��~���$Һ��i�i�$$w�/-�t�'�C�[��?�LV�5�`�]�pZG�Ǫ*�^�|��۞�I�"�
��9�u�M�ƊC��'[���1y!3�dcb>p�"�C�A�UEX#�yI��x[ �I7�� Bc��-ڌ��,Śa�u�wV�:����H?�&̂a@G�w̒�;�b15%1j�������#DcW�̞=o��`�z����j.d/���cl��i��)����k	]�'Ѓ�篟�I|�t����+���؛~+�X	��L�c�d�g���g��L,��:蹔J�;şT8�I���)z���W�Z�=�{���l�\�`��?o��T�،��O��;��o�'�һi�z��m���#�~6ii���bZ�Ե/e̕�ݥ �2 M�b{t[����S��zr�W�<W��a?c����!�ڪ2iѥ]
�Yv��UT���Y�cO�*q�h4ESRċu��'��pC��q�aT�ɦ��C7�#\��Ȉ;�-}�$x*I�.�Dߍ�ry� TȾ�9O�w�3�h~`��'ן�d�d��U���c{��~�!M,=����u��������i=��@��jK��Z.G��7��V��\j�8�Q���4�@�U�MB��Y\�˿��K�J���6�D�����P=�rna��q��ȴ�;�Ο�z�r$��pPԓm/.�	ke,��X�ޖ���� 8���j|Ī��}�g�Awݨ����PNh,6��uEL��[���W{nyx��,�����ozR�sL:�3�����W�4�0B<@Ӱ?�sv}��;w.9i�� �<?q�|�(L�Cp�y�d�W�ջy�������Ϟ޼���v`p ���K�������Z�zK'��
�Bq��hK��(�2�
m�����Ѿ{��}L1+��a�1���iw�G;��qT�P�oq_��S(t�f����|���^�<�;I�Fk5�1��\��A�On�� o9���@B�_A��';f����4Ђ�.�94ڰ[��3r����2Z�:,�3C�?�-�9V�g�e4Z�zp�ZQ��Bp�z����Zj�}jR(���J�� z�H����#��l<=�н=�G�A�����j�=�&����^f(q6��85m/@��U�[R�qV�w��/���ĵ4�U���v�4�<ʈ@�n�����+q#]���[��d�,�8�v!��q:~���y7�I&�heo���S@�yƏ|M�+�����>�W��Թ�Y������;�S������S���H�2d��_��dE, �!�^�)�j����ˉQ�M����<1�_б�
��U��4L�&�v�^����/��{W[Hcܮ��u���d<�����P5�C�5�E����:���Y;2���a�W�'��W�b�y������Q���e*萍��ϥ����Uf�.��`!���!�����2{1�^�I�mހ�'AWs@}��=��0��+VL�5��l�O��I.&��:f�hY)%�s!eH�G�g�G����W!�_*Jٺ�u�;��>�v2���(�ڪ��P�֋�{�~�������!$P�Np��~]�FK�������"4�
Jw	}����&�/O*����.S�ᯂDl;)���+��ڢ4��GK��I��F�1�6�#�#I��%
G9+Q����_�xNS
�z�x%"��=�:�k�S$�I���$���-��+ۼ�������O��]�
?��ksO2��ɲT^�.��� M-��Z##�I��d�^�v	�+qR(�Y*u��B����o�c���	�t�`&Xy�dLk¡V*%3��މ�/�*��1yed;�ȅ�b��V�c��w���Z�iq�U�(�Sŀ���֒�2���-�6zb��k�F�+�gG -��|Ƕy�d;4t�l� �t!���LO���+�"���X�}LL����j�H��R����������ҝ�S�x��`��ǚ����\�����Ӽ�+w�\[���Y0�ߟ����HV?��B��E؁�'�B��yB�/A��M�Si��NWxL/�°`h}(]�i37�z tY��� �8����%�I��BX��U�����Խ(�gLzT����fp���AAQq
��MY�T"w!��h��<"��s!��%����\�ଝ��-l�ɼ��,�'v!�����AL����,���h@��2�$�0��XiY�q�[}�6h�f2�����U?���Y�!��H�a��;���> �ncP�(Y�_Av7�Kd���C���n7|�Ȫ�IPo��G��fh�"`����rkX틜t��N1&�>�XJW�[|�Lk.	/yL�H�u�6lqԥW�����/�:@����R�B́�^��l<�YѪD�Ps���[?u���)@u;#m/�5*�3!��w)%�n�@9L��BL(�U�Ǿ�x:i�qo��0٘�"�d#�S��ѭJ����]�uk|v>s���%wU���f�L��"{wv��-�(�L�c 
,�����&�ՉPM��H-)�y��d�/{5Fr�.���,<M�̗2�H�I������&�ق�՚�U��S�#���]���r�e)��P�#�� +G �_�K����Ϸ7�W���	����G[.��5�_��sh�L�>HK3��tZ|�`���A�$��)J���#~��cF<���t���7�F��qv��:�N``�
#en�[�q����='�.�Ʊ�����#��@�]�K���ʴ��纶_{8�/��z���?<Ry�<*I����v@�\{��4����~�ƅI��U }^�"��ey5��O^>���&i��(J�l�����Y'�ڻ�9��m뾩��\�=�����+h椒/�����P�R�As�Xώ�x��UJg��<�$�/�@f�oRR_nM �,����˯C4�I��֣�����-Q��Y;��e�� �����`U{��+�o�zH�_��<#���7M��Q�2\�g-����ܦ�4��B@���m嚚��*����Zc-�]�%g�=5?�s���w�tAPޱ��|\F6�bC8���
��Yt�����]\z�S�	D'i}v�����g���`�׸�.�U��#I!�@-���� �$��3�p��df��=_�	�չöV:���TԶ?cd��'x���r�|��6!��	�I�v6��A|���^��|��@'�� ���5{̰�"iH���*��򶥾�+\�A���ד1�v���Y�Ma��;3rNp%���?��q�nțy':��mw��h1������w,'0Uʍ�15����|l&-��{w-���,f+���X ���yI��W�OG�5�D�$����E�����&�AG'�I��&���f�K�7fO��M�%�ѐ�J��]�d0���J���RM
1�M�Y�#E�Q�~si&[3���r�ּR�E��]��q�K\z�0Ƌ��H)�u٤5?;�bϘ��
���W9@����P´��\����P�[�u�֊�a�\l2�Ǖ�Q2VB$��X�p��$�`Ru��K�4�~~��'���p�V��S�O!�XL����vZx���{.�+E��;���E^$;�|%!6:LЧ��]9����@m�+�0ALG�kC8n�;H����*���e�c���n���kW���w�a��g���DgM|C���c�,E^߾)-U�>��L��}:O���&��ԃT@�2�Bᱽ��АM��5���Ya�?+�;%�G��.Nܽ�dd$��b�1���3[���@������Mܢ%���2:<FÔ�+�(x8(K�ϥ����y�P��&�n�+�,/�f�p5��qZ��U��,�'�}R�TV�᦬���'�^q ������z�dE�V2��}�6��b���8M\�fg�)�_�p
�Qy�(̕���I]qa�e�~E�"fBڲ�Fe�_�1za~-d�M��W��%Z|��K^��ѹ���0K���J��JB2�����,Y�AWMY?��!�u�&g�FvC)4�Py���p���*�6]�(��RږA���uAcc�\�#�!'l?�;ެ���g����������^-"s�\H�m5䀲�R��0*k����/��D��6�H��.��ʴY�,$v{*Z�����i��W����<t�(�����l4��]�����!Oف�'?��s)��`�[El��E��x��;�}�U��4����Q�8�b(.��H��oJo���l?騢��	��l��sg�x�{v{!��z9|+�1Y*��=�s1'�a��� |_�zDɥ��癥�|%;m���d3VoD�[��s�m�6G��v�љy����s�А���4�t�$�_-�H���r'i_������[s�m}�p/��g�'H���ij�G�7����DK�Ck�%�����L�xytm�Z�Y_B��]�#t���n���W�����)c�Gg\�U=�j�ۘ�]&*�?i9P�"����\��8�\�!KyA�O��u0dn��<.L5��/�V�-^˕�M�ã��oъ�k����Ա���d�8EƢ�{�?��3�,5j�yHt���9b)��`�R�~�-}�X@��Z���6����JQwb�jȲ�k�	��g݅O�&N�ݰlbb$t�4ܤX�~"Kyj�d��F��4�$U�O�W���̯y��y�.(2�@<��Q����fM4�Ui���	�������es�*T��\ǉ)�#�	_���_��ȻA*�������XDs\�ڕ$��,����}�Ou$���P�+%��:Sr���u��ԟ����j��~���몐��J��@�_}_���y� V���Nlb_d�����1K���=��Mw�0�xB�/N5��m3m) ��1Pf���L�������,����� H����ծ�Ĩ*YQ�d��k������8,��<���lG�);��Z������z��)��!�x��T���΀ס��~�� 	��\�)�du�Kķ�φ=�"SG�8f����њu�3�u%yjM0N^��J���+�@�oQ�0����XQ���D*5hȪThRl��%y;�
u��^�� ��
n������q]���mlO���3�o������aҵ�(�ĥq�D2����p���h-���:�J��8�J��{Ǉ�.>[]d"��`=P�d"s#׻������K"�Wy>����ڠ��TO��n-�1��Fu~���,��,����g�l�ɮ�I2�����`Zŵ\���c���.Λ��.�JR���P�n�`]�p��+V�(=�Ӓ�xR6{��N��y3��0��ݚ6\�?y��C�a�ȋ��CU۰�1�FTu�}?<���5��9�3�ح��`e	�1&/wh�q��H��J�+K�!���#b�.��Q椬�C{kD"����ޮ
��u��Hd)u#Iz�=
Z:�[%�c��l��5�Q]�Q7�>)"	nVy���1�9��Vl��D�z[���� ����ݝ���ݪ��#G��iO��xNm'	#O<���T?Wi$�B�i��k�6�� _.�^��Y]V�٥����T}��g�1�D۸Ek�ӌm�_1�ζ~�5nl?����h3\��(�N�;lI�����&���,+�Gh�&��	gtrk�2��]�Nu$`�昏�/;>�qjסU@J�ՀPd��I��>no�Q'����!�|]�i �b,�%�3]��ޱ�>&�;���ɟdJB�lY����٤^<Ps�:�b�!��V�}���g�g�.�G� 5`k)	��ֆ$��it)?Bd�L ��匕z��4�;T����pF=�Bw0 �K�0F����Y�����jS�n�4��}�y=&������kj��פ^a�4�nm���D;��5͝��&`I������+|��Cv��r���FV��gFg�Y��-G�t1�`V�����4�VWo��􆵆T#���d-�_��xQ\T�d�;�т��E���r�c�=�>��zR^��;�F��(�!d�=��2$����w)1ũ�jy/w�ckͬU��^�rs?y3���&Mu�����L%t��)�CO-v"��3x*6����ci��g�ݼ{�hx!��L-	.}N����U5�c��+Q�R���~����s��ȵ�h��Md^������+�sn�rq�sX���K�1��K5�������Dʰ���$\3�����nM��l���܂D�zhh��_��ˢ�W��TD�&\r]��Rr{��G��̴�/�W,�g/�}��Lι�*ŒKK;�冦.��9B�sL�����X��f��v�h9��͛�Oo�����{y޲������Xh: P�,�J�<�K^Nw��UJ�z����H)��Q�e׺lϋ�).�<���"��?�cUY�&�7���J�������7d/S�j
����)%rs���o](�6f�{�乪�g��2�S����P��U�X�?:F�p�<mg_��v��Ѱ��#�Cq�"�Y��#prH��o���U���6z���G���\�����SK�2}(�+��Q�Ċ���l���Z�|�k-�������O�� 82�u����P��_r]T
m-tؓ�U��&�Y����F�S��
G�M�3쨏DX�.�>�]��U]y�ڷ����I?�����D� ���=R��)���ר��00�N�CMn�bj]=�p�r����q�s�p�$�r�c$���J1��P`9��LdGD4M5�4����kn�E�k��f��W��U�O��<LX�y�)ۋ��s��z�/����ś�3�@~"� �����.Yu,ߗݑ-�L��?{#�ƒt������ږ��=�R��G�Y/S�(� �w�2����z"ӆ|B��������zP��(��Xjb��Hq��ˤ}1��E ע��~v����KK0���<sP���s�헪���PE�H`h3Q�[|o��h� .�D�tuq6��dԁ��������Tf�^�����Q�������f
�h���:Ϸ�Lg?�G81�f���GJ���
X���QSw��%eaʼ��!%�T�@\��J\�M��w��u-G���u%��D�g#A��m��X�{��#�@�3P����l����'s�����^ /I��]�hF_ n��dVC��A�$τ��i��� ��R�ӝ)@3����s3G��&�	�Y�6�>j�)/��C�(�D�5�G����|���c&4�W�����Q����~���Ҍ��G2�K�4���@���",����ř��S]Ré�+�`�����!�&91����h��b+��|�
3�4H�Z�f���휉L*�p+�C�%;]�z{���F���?ۺ���+����N�|G��vng���1nW��Ķ���q7� 2��&���3-�;U=���Q��ȹ����XP���/�8 U��0�rFJ���B=�\<{�m���I�d��8�uS�/�]z�U�q�<3Y��N��)h�B����[��k�.��D;-��p�5�Ʃ�n��:�(���M�'�`�U�� ����t��Uj~�$^2.E�FåX,��j���������b�R�� ]=��?�AB�StPCD��ᢚ����x�)�p�c0�����p��3k������X�4Wy�}��u��A7E�&�r�k��+v�c�{�B���^�ӟ��n�#�sH�����\��z4feK�%�����b��%A���t`�FT�.w��k_b|�'�>~g7��qu(���>�/l���εB�|��4�8:�!� 	���i�u5����
��81���!q���t"S��S�ަ�=;��$�"�ۍ�"�d�Sjd���$k^�c"�:������Ž:R��b?xO���i����q�O5� @8}Y�yQl���\ ����m�~�
G�@�K�j����m*;,~�c�6�zX������*��-
�Z~�� tȬEt�䥈����IP���6���%4K�:<2-��z��>e���;�roA�$��q��:�������̾��F���Cj�t{N�E_��^�#L�Jv�F1N^`.�;A���\)ʝ+�<����"��[�CX��L8-�Cb��D��[�W��(�_��t��A�h��3q���b�����HWq:B򆨀*� ���e0�:��Vɽ���v�uv�ރFSc}�:I �����I��$��|��dw��ԡH�N�Th�/NQ�<����:�:��S�Kd�W�"�E-{I�BXۼ��[j���������k��=���u�6���]=�Fm?������ۗ��h�����I��1�nw�=�]�*ޫ���@��2S�e��b�SYN�}��y��\jd��1�CZ�����T,����DneJ|Z� ��u�����oUƽn��v �����Qǵ����`+?3c����'�ʇ���W��F�e{G��H��9Vܱ�ݗ�������$���x��5�41TL�`g�W�f(1[42�h�N�zw�QRq0���KV�G�Eӛ�P��zgc������k�)6����	�K8D�x��(�-Fz����hb9`��<b��G�SƑ+M��׋ӳ��׍5{�&b���F��\��/��E����q�Lz7Q�Vi�t�

dSXaC%����G(���m���R�c����
��#tmG���[�����{2�P�ˁN1c���F��H~��v��k��{+�B$q�W�����⁂�Ei����N7��8�<�V�`2��w�u�\H%f-r�X[Kg��}1�VLe���ڪ�jC���F[��b�ըñ��s����	v�#�H�sy��`�V�9�R,{K�
QĮ�WJ�ז��V
_sX���q$J������V٭NØ���3R���D-�6�_ϋ�� @}N6{8�|`���4�6!�η���)�P��_����ӈ�+s�rj��0�����k�d?LݬLXS�>���� ����Y�_�,�&���=����]����u�{�/��e�V�Y6⢦+8(5���Mq��pH���@.�P�\X��(ga ��6	x2�S9��QC|o[= ��B��K�q�?���ZƢ�S�(�K��J���������xs5g�_�-Ц�� ��Od0_-ʎ�Z2�u1q ����a,���$�J�R��*s�� �$*j��opeKWHX�w��ck˪�M���.�wGc\������������;d>�z�r���ݤ/��C��X��Op3�t,�"�,:>�SW�1[��hN\v���4�5x����s�5xg9���W�۴Av�@��=mC�%͕$nn�n*�- ��pT�HMb�*�Y�O���W7�1gL�|����	��fT}pȧ;w��Xe��^)����Upwç��p���i���i��:���.��%�q�ݼ��x9Gʐ���!�m�[��t%P!uF7��?`��ך".�Ń��3���qql�O�Y�dd8n�0�{O���p��>Q�`ʽ<�WVU��~ �}D�	���jP_�6����0*#���xp�HV_�(%���Sa��jP�Z����O��m�mb���Ĩ�&�]��� ��j��u1��o?3�����r����s�G
 ����bP�߉����P�XZT�1jqxQ��A��R�
u�d�<7x��q�x�Ә�Ss{��$��Dp����~��š��(��iH{��%cuL����p�#4O�e�l�	,�[�}I^tʯ��bw3�>9ۿ��G����)���[�;B��q}�/�5��4��)�v#�C^��?��Z��ǵ>�GYcM��J��c�u��߻^>6��n�[=8?w�RʮB���(�Z�k/��)�%jt�RQ*�W��;��KL�G3�B;Aex[�c%r	b���>`��#�אqy�sk����'�wH�S$����?���v#��b�������n~��m�<�y�@Kk��5�h����Yl��A�M��*˸z���~�,����J�el�m����/j�5�J�2IⓈ�z� X��஗�Hg暏$�\���VڠkxDw����4JVY��ɏ-�'��BP�d�h�"R�~k�����We~0�a�����'��ۘ����5+ �ZW�»��j(�����q�/���X�����A_P]�r4�l�A�}���b����y�-j!�g9�&�%Ra�BL|N�R�3�q6��:w����fA���_0C�^p%�
0�s��ȁn���S��� _�H��1���,&Ql������7�����'����}�+��&V������W��:Sp�X#�b��ì���`��Q��}5�/T���m�� ���N��B7dL4�&6�i��	���oI����Њ����B��݅�"�M�Q���/E>4L�j%H��쏧L�FV��p�M�Too��B,�2�싳�y1�>����ޮ� :� 5���g-�()65fMM��<��Ξ�����,���d�s��g~�N6BWA��~GϹ���B ��k��6�Z$���]�vI��p�E��X�%�D���Q��no8cq�c�x�4|�f�t�C��z\���b���%�
z��h}P�P�/Xt�LF�f����������������LWס�>�'N�-��U3���H��w �G���>B�!�X"�<Թ�-�|R�Fw`|���f���(�������bIK�Uk�U�@�IN�J����`���.��lFɱW	��cEV@CL����m���ڱ&���dP��/��-=6:>�#y3u���X���Mί����6��W�g��h����=So��hJ�̏�+-^w��[�����RxL�ЬO��5�2�\�x�R�N_�#}��0!�ҟ�$��5����ޢ�ә+�7m#&5l��dE�o����Uk"�O/V^f9�A��<��v6�tˤ��o�^��rs�BI2��~�[��0�A����8v�����3��J������`L�s��+������� 7�2v64�*A�o��*�=6R�n'�!!��9��p�=�O�F�Ciх��ixY�Mt�.k�xAjU!d��c�0�h��s1��)3{� ��#��Q*_�/V0Ж���n��X"X1j��F�!h����/�N�0�un�3�=^�<�)U�pz��H�h���,�D9���_1<�\V�a�sݚK�ڥ�:��h��n���h� �S�-� qj�+/�)�{֫� ��KZ�;a?΃��f��Se��9JQuآ(���N�݋�����#���q�~°}�k�,���΃�H�\n�6�q#�gۧ���9�촄?&C"��U��z�$�WAt.c=�}l�������Vǘ��ݫ���ݐ:Gb��i�LۖԼc���ϫ/�����cE.���^)r�������W��X
�ހ�m�l �ƛ#Nt��}ܮPxt�,��I��}���vV�]΂w����}l�a^�GtgR0�S˃x&\�i2�ݪ��^NTf�Sl�[�x����z���A��.�׌����E�e��.���j(6�N|�-~�E��ڡ��
����@�#��ƙR�j7H� ���8�e��3iB��
K�B`�Y�/'Y&\6�ۜ[N�M
����q�I0Lմ�v4o̫�7y�Ut��/�����;����$�7�>IK�2���M�8�B[%��P�d1�Î���P��WRW���}&�����g�fcoF�M�M�9Q��yKe�JQh����.?U%��J*��7�#�������#Y|���%|�w�xu�(c��U�O��i�r���z�Ŗ�1�QRؔI�< �P� c��$�>�Z$UG��U�@ 9T�jPi��.��Ϫ���cE4mHH4�8
8�"�����J���ݍ�����\O��>��?��$�S;S�5�c
wV�[-�_
4�>�LiZv���
8�GE_d���N`�w����0'����(n�V"�f��~r3��u'��	O�D#q����P)�$b��A��FVn���g㌤=����\��}H��AS��iEZ��V���p��(=���1T��-|~��EL�U T&4r��bm��y��H�G����|�dr�}#�Z���c�M~�8���1��S2�(�.�p��� �;u}��86�<���@(��r���+#CN�ץ@"�Za��y��7���J;U�:�Ⴃd�	<�*��K�Z吺��oḞn�9�'4,!�����c�9gNU����x���2�5/c��<:H0:��n���;���� ����1�E����D�a�m�F�!m_䜣;�Tu\	�M�~�W�c�{� U�!�KAG�D1oc	@�Z�7����^�] ��\�as>�j�3���v@4���K��Ȕ�zm;L碕�A�*�%H�����������o�.�]3�Q�b�Q#��o$@�~���H��,@�&3/i%B��� ���L�9�.���2y:�cm�$!�HD��}.��K%���ä��bޫ�1�!�O5K��o�F��ۚC�{J�lO�=y~z3Վ종�xc�*��hM��M��N�Cv��x��?(K l��.� �����"s�'�'�E��aH�A�����狖e�S���+��P��K��6]�{Ⲝ����w5-5DX����E۶�V�bg̏Z��$���V��}�&>h����!ߘ�kZdʕ[�3�ܒ�	@�\�?�q?����t���Z�M����~Sn����ga�b��'��V���׎6g��	e�wu9����`��(��=�k"8��f�)[��( ��Ah77Y1�U�Z@S-d��@�(��,*�K�JO�eA���u�K�r�a�.��J��bd����J��i^�4�&h�`B�����WZ<l~�����	F-��p�lUK�^�_f�6>* c�;f�o�e�Dl@̀�B_�bj�_�/�ӷ$:x �iKz�%c�}�Cn���1�ػ~��d��������-i��95`���1^��y�pT�E(���2Q�d���dq;3 �����۹��E%��`���]"�_��:Q���g+���?���s��r��U��0ʢ=�~!��U���Nk����X�3�F�ei��>�>$�G���|��P1!������}2K8��(]ձ��.�n+lR�F.N�r�������$èZ�����	6�۴���Ȱ�}+}���2b�-u
�zgJ�5�R���Pg����j�A.�U�NmF5�]�S�V�5L���Zi�^]�v��4o֧�?�Z��RG�c���~�yU������>�tTO�ҟL��ȑnQ��*��/4x̳��u�)����X̆�q_�H�>�ً�g�G�j��t������ו��#�(1�����6Y��'<pn����3�"�A��*r�JP�W��v(���ĺ?M�!�Z�hܝ1��tb��I��]��Ns��#6�+A��Tsw:��|F�$��Z�p�D��]�0���P�f�n�HC���.�w��B)��#`-�$A�E�r� G׏s����z���
d��+ǵ��
���sPkxD���U�_��ǁV���biȈfՠ�5�[{�;��ܧ���A�� [�;.L�ݿjfV�&���ܧ�zV(�|pʃZ�����5������Dѻ�l�ǳ��&]M��1��Ą�pP!
˸�{�����]a;\ .�)� ]�t�ea{�$.�#MM�.� ����܍�x&��<*n��cr��CJ���+ܴ%ne��Q�*�6�O�Fُ)���ϴ�T=��"&��! �	Fʣ-�hV�ܮS��5�اyH��xm�h��{�y�0��}�ôD��ߛu����  �J�(~�8ڠ&���9�Na�q*O.�h�O��v"t��t;��[�$DQ)��߭���
y�l�H�)�
U��E K��H�������ۏ����v�D�n��	ܾúf2<�z?��e��UT��晉��$��l�κ�vd?�' �0��>MbG����v|�Ԇ�u4P�������]X�ِ��,Ƌ����K:@k��v���b�Z�9L�Mum\#�2�{f��p�Dm�?Iώۧ<�r}�.A��87��fVZ���I6��F$��lؕ�#JIn��n#�O��D8zn��x4%�TȪ�\�QN�l^<¤[���k)i�1���b'H�&�������Q��ԣ �5tp	e�#�z"�T��]�?[����R����m�=C*��M`�	1��ƙ"_�������B��]'4��Gf	t'�B��s�n�֡0I_�?a|�%�v£�j�ͺ�B��P(�>ld�8i�J'�lz�5x\�pQKS� �4�������~�p��G�&}��I������y٩;�ֹ�DjRX!���E��0�&�Y�~��7�sz7l��z,E-Ȫ0Q�-�eK�Ͽ�:�~��M��4T|�VC����-l�7Pvsa�B�Nw:^&�@��/���u�0/e�h[��.�A�e�y�C��~\z/����	�	ᓯ#\�?'uЃ"~��植�`�kD!���pP�Ņ���F�����U��S��$��F�·��z�f��A������r.:�s?���!t-�翩�G��[r�K��"�Z^_���+ޕy�J��H��_;C� ո��JYKc���؟��β����)r�u��t���YQ�A��½���$Eɹ��9=��{\6:������"����|1�m5��x��z�/,~��������u��e�L�GaJ�zH=N4C�*Gf�4Xۙ��lD0����ن���xЁ�;�8J��HϣX��ES�� ���h�Nw1-w�0ޭ��L���h�7+�އU�l��/.�?O���"������!_�n�57G"k#Q�Y��}Z�Nq_'�`���9�aϽ����d��o�u�W,a��F�[�
̏
�!'1;~��XCc1~���{��vv�� DA'j�|T<�nַv�:AU�n�-0o=�d�Fa9x+4C����D)D��2�!��,���}��}��bKC[���� W�$ʑ�F
W�� @Z�ݰwHf�o�
���X?�s A}��&�l�z1�u�Qd�h���G��'�8�=�c�5�1_;Qy�������gav�=t��qL��N��^x�~D�x����{���*ȱ㖒�OSe�-zaf��h�Vm���)������C�
��H�]�wXx/��8!##9��ȊBC�dGo��ױ{�|�8Z��x��5�A�tD��m65.�{=HdYi
�����Y�!� �P$]��>��	'4��+d̪*�X���;h�޳���@�Ӻ��wt��`+����-{{4��j��r.�6 �}M���� T��盈
?	�J4}�_�8�SM8��VN��t>�c|ޙ/_׷�7�{Q@߃&s���4^Ѕt�0�$m�P�U�=�S����M���a��^}�g$��s�wx*CK��]�{'�غu�\u�/hd�f���g�PK�d$�IY��$�����IWwLnǣ�����V���[%o3>!c&(\�[!p����'�C'D�9�q3����
��!��<t��z|m��7��[��a��0���hu�*��~+{��ZN߉lJm�W�؟��N��z8�5�K��il��b^*^�V������!��A��C/�5m��6r���{����N����`�d�e�'�5~�������ٴU��gdiK��޹�c��nLr"(ˣ�!5s����*O�_{>I���0R�Sy9
n��@G�FʰP�_�-x��=��vc��3���+�g�\t�ӟ/;�c<���,a�
�,-P�r�A�J����ڦ�hp1my�I���)}v4�T�05��:�D�#��I�䈦|I.H�)3O�g�7�����]�)S�ǉ���r#�X~���5T{�[�)*C� �(��xE/򀓈.W�2+�;<d����^�G������i�^5t��iF��)M;3u���;f{���W��Tm,n�O�O˿/�6�F�'��#�[�<�o��K�+�R׵I�����4���Q1W�
H�c�Yv�O�h6}������XKTC����fk�L1�5�*2W�d��Θ* [���|���~cH�Y�[ou���=aj�\�P��V7p�-LpQE09��2ʸ$���W��X���M2�&��W�޼CC�����v�a��Eރxj�7�gG0J�]B�0H���@��m��i���Iдkt���	V��[RJz-`�?�_If������թ��ɓ�נ����������G�~�C�W�������YO���P��*p���5���BY\u�I�K�m����Qt�|:9�i{�㉯�z2�#�)���9�e"�>���A�Ы���ȩO����5��4�����j3�� ���,�WQ$N���u
H��� _����������c9���g�����.'gW!Z%#B��a��4�X�&]�c� 6��j�d����.-����&c\��<���n4$�(s����YͽĂ��ju
b���}!�cL1�ս��G�Dl\8%t���25�;mn���H'ŌA/({�h����%Y�I�ÿ́�ޱ�p� �q��T�kߠ|�s\�*���Ï�K+�]X~+Πh�"wK��4z'U�P�i���cHc�N]y�
��C$�;��s9����� j�UP��cn�ӝ��q�*��%�Ш��֧v�f੦e�o(�E�ދ�Y�j��e"tJ�[ي| HL��g�Tg�'0��=2ѓ�w��x�����&������;#�t��C~��8u� ��5+^b���9�0R,u釜#��ϧ��6Z�t^c�3	N��m�g��?�ٱ`ɉ4��jc�%Ҹ�q�(F���s�d��f�;��v�Z�Q�4�[�����d�r܀H�h��XN��&{�|��i���5�V�Eiқ�6�N䄩�ʀ������Za1/ֆm9!en���{8�(xU�;A3]�(�r��A~^V�󉚾��#����IA�}X�����+�gA�AX[��g��B�.����g|ߖƑe!��`�>���#�V�t�uZ���V��=%��Oo<r5zi�q�'�C��	�z���璜�����p2�к*_��'?w��7���,���!�/cO���E�5�]�Y�J����j|������跗/a�v���tl3G�&�����^(�솊Oc,곜�/dM��	���S�:D�;���5�{�"�	�
-/�������LNi�r�e�?��#�Z�]f��z��s���@AF��g�p�Ug��~�]]��sX��u�Z�Qf�E�3�����&�ȏu��w`���|P��r�n�ac�q�������zBە�;ᗻSIWcO)�̈9��1�P�xL�)@Kk֤���j#�˘�Y���a��Z[��Xe5���͝"�%J�.A�����K�лq��r8����N��6;Jxh1����W=*e�?��BE̿ ��>���@1X�̪�"gi����]|��~)������SN�%JMs��W	8�us죐1I�;;F`�P}�E�)ғ�gT� ��'���&�ʣB�2DF3�w�};�.^u�>����%9������&�kQ�"ⴎ9����:�^�.=���$�=e���5�K6��4�!���\|�[�~d��9��5�D��X�����V���d�-�`�cc�8S��9�kG��A�c�;C����8tp�N�{��r�$�c����:|v�w��̿� ��G$}�|-ك�%��^5Rۼ���  @�l�-��k��3����F1Е$��_�"X�&彉������	�/�/W9�t^9�
%�I�#��R#���e=��#�q�!]w�gc�2^�w_��s]��� ���aT܄��s)��|�]��SJ�D���JF�(���ê>�U�W�ă&��42���
i�ۏb��~OO�@F��y=U����[o�5~T�~,
�/�0�t��C0D����O<���sE��3n�t�y,.�w" ���'��0��E�aV�5s�O�%��ΐ޷(�p,�)��ո�
��� '����-/ڧ�g�r�?RP���@��5�����^���i� H� $�f������%8s��l��C`���#�V��U){�ݦ�sw_�d����ε8�����S[Y�DNB[�G�W�xȿ&~i��C��L�!}@T(?at]�Yُ�5	#`_M/]��1���#?�KT�����B����__�_Y�*J�y� "�����ҫ�j�-�@���X9���Q i)-3����Z�X���%X*/�ֿ�T- ��'�D.K�W��߳K�����SVE��i�
{������TcL�(k��V�0Y���l��P��lĔ���w�w؜�oz��B��*�d������g�l�Fh�������U��9����� �wP��kR°ƈ�����|T��n���E�fy��1�,YV�p��Ҋ��!|2]��m�,?�i!bZkA�#B� x�E�����g��lՃ�ȳxm���Ip7�[�z�91w�S�����y��oa��)>Rܒg�x�L	��Y2���X~5�M��)�H>� ��}�p�am�a��`d��������u��1�6�Yt �g�H�j4�н�$�*o7�"uV��� ����H=Zǋ�g�v�;S�u���A�jVp����&�+l��NR�6���~�̼KzNK%�`���/�~�ifo^��*	��:�t@��rq��ƒ�6���<+������wЮ�=���{�̪<�.���-�
��������a)u�i?��ǖ ��1�ق�Cpиԟ�F�������}������^8X����@�Nҥ�.Hk��"1R�&��{�}��ަ�Q�L�2�#�,0��j);/�]�͞<��YlmuK����X�xTG@�]��s!>��:���VwH�q@U ��*��x�ZB	s,�7�X��m��<�Wpm,i�����EE������cm�͕����	][F0�F \.�=[��k����R&��~ V�%����j�	(�U�'�Sѷfӛ_���ËȾe���n����l��e|�J��BZ�l!|%���W�}��i���^
�Ȇy��5цEZ��M������?x �e�c�ͶP�*Y�)M|'��LQf�V�\ڶ�Q�����L{�I��]r�DpA'TL��'��N���ɫ�V����i�e��X�|鞕��DG>y��f���.{���RWg>��.'��?�la��8'��B��F�u�T�ծ�q�bS����u�7}0G�M-��5�A!h�x�<�ܸ��\h��]�7�@�#���)�!��t���=cp���	�t�4�#	��(-Xܰ��r����#OfТx]��-Ƅ�� "��9dc��!�X�Y��R�1��m/��?��>z��v��H�A�\���B�6�t���ՃB̐X��]�G"�^��G��ݍ�1��o�V�˟���W�3(A��b)J���s�h.ʢ�-��iM��+b�W��m�^R�ɥ��^��Q�JE����O_<t�/��ׄ���b�Y���ɯ�Ew*2Q��{r��b��#��4�ȟ�FQ��j�@�EZW?L��@.z�J((����Z�ƞN�8����a�d��k�����ҏvZ�A�\�����߮ �I�vj	��O��&�����ˇ؇p �М&E�Ԕ�j�[�@��uv�G�_��v4�\Eb�m�����Y<�
ŀ]�!��6����xm�%�Y[��nw:<�	��Q��|D�g�I����kx�5r;j����6cW-3�â�a ������;ک����+<�n&��G�
�V���7h79)EL�j(�o7��S�i �=��^�5t�Z��Kb�{1\L�i9��|�~/r)��]e����m��� �M��<�|9A0�]�Kp��u~��k-�ʨ�ݨ�n}k�5og�6��q7ۆ�\�9�9��(s�Jy� �mr�ԽsCB�����'Ԇ@y��`��l�s,��G,"gĠ�V��ĉ��)�8�ʆF�x��6�B�!�1��&�׻"�y5��m������d{��V7�X�h0�M��@k�E1b�k�p�w.��FdQ��j�8�+�����c?��
B�(^�W,h��
yXT�4?\�`H4"�AN�{�&�ȍ2j�O�6Z�N�룜�SH&��%?��[��ͷ�N��W4�S�ʆ�O��!U��# �`R���P�Џ�kC0PT�9��Y���Ϛ���r�Ǌס�$t	�"�r?�O�x��¡�^c�g�0̚��b$`�ŞM���!�cA�1�"�UI�p�ov�e+�Է۪�tj�!��Y+�������u2c�����r7m�M��!�"3��v۠ƴ���6C���ba��3}y$��
C����]���]�� �1�y�jE�(�D�y��w�8dP����ݔ���܊�ӌ� RՍ
�+�nm�H2f2lu���]���f��W���TC�r��=A�x��'�4��|d��bY�ǧfC���05s�sI��r�{�wC�讟`QkSW������XQ5�Z;@��+'�u���cLlyʅ�n��.;}=E�Q)�T��b}�}FW���+���3.�@�i&�Û�*F�uv��UAF��'�d���$�S�k$�*5u�b`#q����Na0��2|�?��v,����5Q����`{�)R�!��*�`�-9�4Dp��w$��jևpq�@W�
wx�B�%?Z'F� 6{D��FUo+Fԝ�0��.��y���_�?�R��S�a��k�=�ߧ�;A?�%�J��1\;Q<T�8�*M6�'��M��ۮ����w7TR�\��^�Fw.��c�i�+k�I�)�x��\����$y1�hd��Z����/o�aZ(v�uO;s�)Z$E�o�������mDȍv�CI��-���76��j�3�[�7�os���9`��3N�ۑ)!�D�2̊1x��Mº��L8R�n���uN�$5�[0��ǒ`�b_?a�\��*�|�A��2&OO�������svт}*�W ���)����n����D�kBt�G�a+4���(� ��b���O9&��VA��UY?���Wٛ�tM���@źq����!������楔�}K��.��v�ڍ���/��ߖƮ�nG�B�Ct��)ky&����z�Q�^LХ�����"L���C��Կ�BNy���e�r�xa $���p.{�dDj?Z�:p��4�it�a��nP���A��1QMh4���_µ&�뗐��]Z���i�����#F#��F�rհN�#Cttwzm�ZYrK*��O�[�訧﹧�6��+=o`�q����}�
vx�r��eR��
�Y�ڈ�:���=q�<�<���:�/�2ѿ�^ �~D5h���<b��x,k�T�?�vQ=���~��ڄʢI7����˧ī ���PE��Y�����?��e�k����	[�^�{��Je�I�|� ��i\�W�2�~�/i�_��.I�h �G������	�d#�5S,a`�LWkK�����Z��S�ik���o�ӑ�А?C�Y��Wg1�O��),��Ξ�������]���3��<�z`��f� ��l$\�5Sϴ{�\WɅ��Qv���Ij��4�d����KL�3���30.�aa�"F��Ϋ�᛾pH�+PD�'��t��k�����NGŚK�v Z"S�g��X��^�ð��3Oo2b*)���^�n�Ok�P���98�~��h�y��S(7����v�S~�7����Y�y���u�_Ą��ުu1���oO_�Z�>!�E�F��Q3z���h�^g!��B'c)UJ��:A�U���G$�I�xRo��r� �̵"	��Z���2d�Ȑ���˥}���m�D.Dگ����uQ!ZF��:�cf�Zi"���ct�X��������kNq,����@�<At.�0���1`\d�^Q��[��`2��>�C'�{�w�.Gҡ8%y[�{y8�kd}	��,�Z��<ˀRT�����J��XP�(�(דF��4�ơ��������d�(@ܣ	�W$q���?qF�	�K9��;����l����Y����t�� �LY�]W+�E�Vm��6�x�V�.3�A��Eb�}����c}>!>D�M�{;%P��W��]�`�Pc�+�)z]�� #GR�%\l�1����.����A׹6�� �q	�@�U"D�h1�>q��E�$.��.*�Z��$=����V�sw9m&LL��1���;�>���Û�d�#����oX��+?�@J[=:u�Aui/m��+v���7�𸅍���.
��ދ}����X���U�PM�9Ov��:f����/s��������q��iq��gV�g1�^��r�&��Y��r�a� ��#�c�4����$����p�[� �M�(-���"�WZ�Ԝ�y�����tֆ��!���V�~.��p���4��̫����j��M�G3.9N��;��c�$Yx/!�?����O�(�R��|����yy[&����c�BN�"#X�L��j�y�
��fp��3���)�1�W�Ek�O�캴�E
�&,��N�,H���oD��.���vR~��`�]m�C��wI-!2N:��:5/@�rW�uH�8I@13���*�0�ă/��B�{��e� <��l���\�����4�q�)������}����-w�q�s��H�C�vSt|���7���̷Z��M9������z3>�ս:�\<�)39�s���7;F��F��ɻN�\��~W����:jH",��v_�z�\v~ _ig�^��>@�U�j&���4$��ϧ9�V:�@(�*�$�3&�˕�~	|�m�l�c����![y���M5,�a���J_�%�L1u<��d"����
^$1����xS�8� �n��u����Ю�F�����<�X� Lo ���!t��y	JOsj�����f��3H|�Ƃ���=�8�=��n��p�1�^}�b�>�o��X�r�H�w�q���]%�8Z�.[�07H���Q�mcf`���';\�te0����[�:�éf�yuhQ�iK�`~|U^�=-N@��j�wP���0�PFt6��s�������I�=��F�áw� �6�t$��&������ə�Ud�X�69Ke4��۰��,l�<~�V=���.��mߣ3��;q�$IdUYJ�,�;�#���"X��_>%q<������H]<�����&�� I����N%d�Hh�}L�*����fF<�ᦵ��l��̀����G<ǷCm�Wr�A��4w�\�<o��l�)&��m�������?�����ۨ �^��K�8ȳI'���l�c��}���X��.�0�=?l�=�"m;�����Cz�	L�sc֑!"��8�
�8?����MM���a֡V�osw��fΣI�\�5mV(El�G�y�养"ӄ��i��~[3��倊<U�⃎\�2��}Qh�r�!\�n��T&�EU8����J.��/_�[:��I�&�]� ��nf<>mT���Jk1W����v\gX�B��eT;�,-�kk(�c�L�ԟ���?�2�
V ��DO΃��,��*��
�=���5�?ߟ�G�r�LKZ���H\�&�~�y��r/)�s�����P���z�?!�T�EyI`2M��������Z��(�B�CŅ �+��t<�q�)��e��Л)�>�9��ZQ~Jk�D�`��3��5Yf�e��+�O��$�^&�(eU�������4�A#gM,�EG��_z^���ԷL�Oi��R ʇ�o�$����>5!�m�fz�y#�FXFt��Ub�K@�0�7�G��eW\�j��4�uW��@ha�O)es�b�Ǫ�o�'�W;�m6�?���Q��YB��4#�K���'���]�R�)���ǢK��U���9!s�Acs�G�+��>�/=+)]�/�V�\Y!i�/�B�d�Ԡ���!�=[�F��U�o����)	��yn�]���2��?�1�Д�(�T��f�D6Xƨ&�E��p̃A�
�g�Ix
��~��_��V�ܰz&r��G8�C�>�7=�?�y�o�C���̫�`�9����]�+�5���%�7��Π,�7�������:r^��
R}����Lĺ�Bro� c��qT#ŅU�l ?����G�]��?N�mw��!�>`O��}&^L�D�̸��
t�'����'Xv�o~y7Q�oHE`��=~��n���D�b�C�-\̀��<2c$����!q�+��:�����X��u�3ⷝ���ۋ�2����ު+
lI�mLB@`]��v���B��M
�lu�bN'�cC�O��i�|�3o	w|,��h���ϳ-%��?��'d됡9Q�����PQ�Ź�>�G�.B��0����e�$�
 �%�S�|8;�;b^-����Y3����{���({x��mP Vj�09j�ݶ^ A���;��e!9\e���ˋ�Z��@��vm��̐�.��������� e�3����E�^���ڈ�y���*��ݳM�y ��qVs������"]3��6.�w���S?}[��l�����ù�@u�W����U��۔7��u��5 ���W��9ܷ��}�mI��e��r��W��*Z�����I	�bt�E ��C2���/�P�|��t��)�O�F��P�kх������	{�����)z3���&M���ġ����/<�)�ݠ���/��%].�LD��?���j��Q���	��M�cM�d��s�n�ܕZ����:�'{N�����Jy�u�@���3��"�|�k��]�d�<��Aa�K<�¦5r�xz�ae���;�Pl��%�?"�Fl�i�G}�@� !�	��&`��s���e�����̋7�|N�\��E[I���X9�h˘��[hڗ��M�9,��}��Ur�ȀJ!�:{&ء!�M���M� �/�3w�������:f ����1ŗu{إl�mz|ߎ����0��.���w	����0w��9���PF*|s� �<�j1�5���1��Bz[��7t�d�����/Q��+���|��	ʷ=��0�,V�?xdu�HPoG��QG=�N��v����ГCjNy�� I�v�.���{�(	~a�ǁ���j�̘�f��*��Po��A�\���	�T*s�hxY�B>�qۓ��h���o����d��U��N�ʠ�-�>ZM�U��`*����^qS��9���Y�:؏�������ӣ���I�؏���:A<�g	��o&u��0�ӕ��/)�Dʤ�5��$�ƽ�Nf�א��g�#��k�˪
+þ[qG�t�t���٪7�vq�(�az�?>�v��9�����!筿����D�9���z�x�ͼ��X��
�'������bNqfBj��)Y��5���U�Jj(%�P�{���tdr*��ق�f�5?$� 㗼z�Y�����>�C�4��g��"q��}:�p&�*t�5�RH��$Y^{��'��l5�m�Gt�_��-=J�%G�ɧ��}��ŰA.4Lh7|��%�\V����O� ����s�'Ǩ�PO�3�6���kuGtX�"��	�z����B�x�K@x��2 -DNo�����DR$����ɎL����~_%w�e,�/
 ?]B�{��k�\��SǶ�0���0%������lR�&mE|�%���/l��|M��o>��%A�HAR����l�ACɍ��7xa����	�t����D��>/����:X�q��棛l�!u��}
Q�D0���0�W�saG����ѕms�@�h���HcB�����g�⸞>I(�Y�X՛��l��F+�԰��c���.:?�v�G��ټ`N�Ӄ3�ԉ���gi����	3۠I�<��]C=�7��F+E^�
�ȝ �����Asc,һqcY/���u|�[M粥��=%1m�<��A��)��
��_:��;F�$�ו�=�5�.�}�1E�t�PB��T)c������ҽΟ�W���L�a�V��4V
����l�+��F嫾��M%@�U��R6��eWj^�eV(J�f��@�����xhB�dp"�Sr_���:�F�:H�v�x0#���U�"]p�>��2|
��LKC�]j۪dgf��ȋ`N;M����:+C�!-���Q�����a�������ͧ�/�O�X\d��gT��4~!��ñ��6�Kՙx��U&�'@#��=B�?Z���麏b����6�`�X[JX�5'��Յ2���A���˩�P�/@�S"�W^p_h{
 6n�]�w��*" �"�����}���HGt�h��Xl�d��ۘ�}EDF�)�B�o�e�˦p>I��[�ν5ZZ8lW;��i�Hgt�&��H�'�fϢ�9�d��I��bbQ�	�N�Ŭ\B�����L��GY�#b��+�)�љP�����I\�x'�h����݀_E����uq 	���<p��#H>X�ş��:p朱�O�2�e�	TYs����p�AF��>��
CB5����G�Q'��!ʰ�~��۔Vְ��ʨ�u��� ˅*��CN�Yf�"�luX����LIU�f��<d�%�����:��d6���(�}�<|-���<6=��������@�`Cd<1�O\֡����<фLZ-i΃�A}D�}H�3ڮj���l&��(���o;6n��5��%͊��w��r�$V1�]LF��.c��dO���"v�
{]�R8���Xn�����&��$2:hs���o��7��YEf.�O����&Na���:��@���\�ҝ�<��k�)�ȀT�6ZjQ��ZXn�C�2��#�i�k&*��ӭ�b7s��w�8Z���U(�i[�o�m�e|��%�����?����G��ί�9��#�Nv)Lo$��㦩�߾�~߷�t=?�e2}��������Ml5�R��^%���� /Ɩ�M3��o��#��5z�'2��	k��w�Gs�\"ߩT=���������I����~~�o���Ԏ�Km��MU����w��Tp='�
&�HL#�&{�H�%�LC���V7-~5r�|�K�QL��FQ���S�`U	/����>fI���_�SP�MT�c����*��/G_G�4Oc���Ԝ�/6/�y�ݺ��H|L��vy��u���4U&��>9��v�m��8S��'�}�H�O�E�2���'M��K#"�\�@G��϶�(�;�g��5�{���� f}-p�F�,.bx�ǰ�{|����Ŝ�ٵq���ޖ�~=i�:�Y[M�ˌ�?�3,�bJD����?14����+=`���Q�����2$�3~�]�l�������: ���Ҏm��t7�G$�����.S�j�r�f���h-g�p{�u�Ӊ�& X�U+ͼ�|F�3��A���o�3@{c�,�߬�Qz���$��|^%�߽J��nZ�^-����v���*b��\�����j;�%���u�,��;!�yУd�6��Y$no#����+!��	��Z���ʣQ����������Q���"��^C�V��;Ϻ��*H0үu�Q����z�Q�J����0/�	7��f��a�w�]�����OŽ����Y����m�QZ��_!Ȇ�hOpo��L�ڝ�K�Ԉ���W�\���o4���O���*��'�AL�[G��&�L([��C�m���EjU�_3<���([��ė��u!���V�&�h3q	^��R�K�bj֠Td;����ƪ�Q�.���1�I��T:#%�8r#�ݪ��� v��+$�&9���BP�X������:P}��2�7��L>��-�"�S���k����[VƗ#���m���$�K��#��� �@��q�	�#�I�	g ;�U[�;i��?Z+��V0u����5k��2\ Ѕ�	+���&�i��j���D���-�F���53�����%���*H=��O~�V����P'-�%;)�D۴{�a.��Q9u?DƁ�"k�i��fas�s�G�O��[W����L~?�q]� ��xPm)^�v$��q�70{���x͒O׹��R�*�e��(!���!3#��
Ҭ%�K>.���� 0ڪ�
�-���Wv
�2�|Juj�p�P���,��hS� ^x�w�To%1���HMcå֨j!�Z�;���o�T�Ńƽ�_zj�>�k0�jz�5����%>[J|M,&M�� 3Ճb��V�#6JI��T��`���y��QrEȥ<��2S�B����&����_�����P�ؗ�A�*��`΀+ˌ�B�Д����%�j�Ȗ\�;�����D�������s�$����O�=���6x���T�(%�zEB�X&��{��G�� |�7��&$�C%��9N6V��q0�s >��j�p�~���i;��!)�c�a��p_���Xw��,��,�����`5�ΤB�AR'��;��n"4�aN7��.Zҏt61,���x��&��6�����Ϩ�"�s[�N�7q�LD)��t��G�Ջ\AOH|��r�]�on@��6yHz��d�_j��ޅ�M����ݩF1�*i?��d���ac�Ha�j�0,F�	|��Q4Q�tI�t�HTS��	3ǔ�Z�����{��B��f��e�/��¡�F#���ۭ�:�u	�uBq��%磌HVڕ�hLy�A��1ΌA|����d4�H)�f��m�$OCe߄��.P:����@��"[[�4;�,BA��N��zarEӏ����; �w��������uœ��΀`Ǵ��_pmgY�����.�q�N��w-�H�R�$�E���q2Hy^/��?�_�s�.��x����V�5���at��e�͇Y�>QӾ(%�O��|�R]Qv�����f�ڜT"4>tg�a`VJ4�Q������ϖ&��V%�K�z܎EX%���-�(���F���.^_O��!n���OUD��3s���DۉPd��Q�:�c��5t:>!G�$�_kd&����r����m��[3#���k)�J'��./ɱ��n�Ip�2�Pp�;T�IX*7�
|+���
��.}k?�
+_}�����0��NF��?�m�)�In���UX��C�l��ɴ�mM~޾Iv��j���.�R�4��e��&H0�T�]����,��%h	l�m��m�=}�U.����Q�*�$"��/6�+���� �
Uͩ�31�a���B��|*�Mll��GS��&��X�n�ԇ��Oa��#���'Yk&�O��+��@ʮ���8�����>yn��N��r�!��<I��3����Ce2�Z��07v��.�O6@��;�ɢ��/�@�1�{I%����a�s?��:�s�k�C���k\ ��Yr��	��H��RM���.v�6���E+�L��N�����l=�bP��mV$�j���ڐ3B��=[��e��/����kO�������P��sp�Y�(��K��Jk�;�PK����ylֿ�Dp�X��ǯ�G�ײC��vG}�վ�Ϣ�j��� -Α�_�c ,v�.��-��L�~f��M�dZ�d�M����_?�c��/��c�dEN��SGzY-��T�A�$�94*��Y���B�.���Q��~�*���]��*���JY]�
 ;N����^q"��}18���Za�̼��Ff�Z���x��F8�_�;1�A��.�;���rA%?�f`B��;��}�C�ɍ&���2U� ӗ���A�Ջ�-��qU���䲫���� �#<��>y��t�m� ��zH��������Dݟ�ޫ��|"�m�eC�Rz��pP&��P���s�Lkґ-���>%�!����-j'����::���ͨ��u��0w����Ls�r?W��#�wA�k���K�[�-y��lZַ*�	y%��y�f�d�0�_�$���� ��S͑<���s�J�o��|�~� �Ďb�L�C���p4��&o`�7]�[c	=���3�]����/?qbKe?��;r���$��{����M-瘉���UmA���lNB?�꿒:L���9_�4�=��=����?r�ě٪,wV��O����nb�"�ֺ�B�ҳ&i��;�f��B;��/n"�ON_�f�]c^-�x|R7��c�
��Y�!�#���	�T�ג�/�J�[%F�c�Fmπ��+Z�H�&��%zBf��t~�}���c�õ=�.څȷ^[�?���Z�!�Ƚ�E�'o���SK���3�8޵�����4`Ȣ�$�G��/M��3N�F�����T���X<;�b����z}�bP�6g-w�+΅�z8�wå�N����4ԞgjQ�a�����$�����kǅ{n�.O[NZ'}+�R�(1��q#�ė��'�f����MO�+A��k�Nf���WT���[�Y�ӊ�T�
\�{ʻ[�k�[Յ�-MGt���2Đ1��bG�S��:B�i�09an֝F� ��Y��QN�a�,��\��ׯ���R=��iS+�*r(�L4�l��@R@�!�}%�z��V�ɓ�TJ�{A�K��3�RTN5�$}�U{�۾�9r��oN���@�mf�ϋo�����\)1� Jv�������仉|��B:�i���@�qU��r��4ܖ7ݪK0�*��LG�� ��dC��^yý$�������C��Q�Z��"��#��^? ��N.�X����Z��8������+B�ju�\Ɨ�2����of;�}��R�p����o���")�Z.���v� �j���]�e-0 �8�;zu=V�V�c�׎z����ԁ�~�S~z�	�L�9�V��?cg���`��tWV�Ӭ�U#�+��i9!����xJu�G��	`��$�*��
5��7?����vT�wR0=��i]4?�vW�qB�ۄ��
�%5��5�."5���C��S'���.�,���^�u#2����,�����<-Bu����3\����\�R[iυ�(ס\����W�V@amHIB��g<�Ѡ�Y�������1З����̀xw5ɂ	op��'����-����-��3�����}�m�� ��AK�&%�2j��%�s���7�-b�bH�f�>%���w�׀El�����CzÇ��+��=�O�j��'��)�/���1���k��"�iG+�����z�ƀhaE�X�������K������|�~��ɧ@!��~鸂Rt%w�y���|8��t<�|�7��2/���kI$�=D�Ž��I���O2��{����>B�.��Ki��91�_G���؍���us=��MU��I\�4��P��jh�@����c�^%o�/��M�	5K6��̴{�49q��k�^Be��#�Y�E<XV�MK�b9���5����]�ڄ �&�R=���%��ʆ�e4\Ѝ�����o����~t�]����;I{ƾ^ݎ%�Y�o4pQ���\s�Gݨ�̐����F��U�j���A�)Ѹ��탦�5�v��V�U�t���6]^?���i��'���t��ԣr��G�,���Ϟ�F	m�c�%2K醠l�a^�M�U�լŃ�����%���M�.�eI���ɡ�t�a}=!cs�B��v�B)���`{DT�Y1��V�jFl�l�3����RE'��	/��E;����2g�E�4}=�)�4p��p�`�Tifv�5�<̻S a7���`$��Fu�1�y@nP�q�K�{��e��K���H�S�
����o�瘮�}f�l���k��W��}��l
��a��AU���*`��+Mk�"�UH��bF�F���+�ѷ�b��+��Yl�p{m�'�8$x�2j;e��;sf��῀����M��wՋ6Y�0��&�!���-��ػfG��Vt��fl����,4�������i�-�T_!W���	M�Z�����I�K��B������PV	�̪g�C��2���r����@~�����t`�)%"����3m��ۓ���P*\�8m��(3��@�B��*zbY6����F(�Xa���֋����z���&�#͝�w� GIe�v/)k�APA�r�!3~���?�� ٔ�`&�#[2�b�zMG�c�
y�Q_��'Ȝ,���T4܀�`���G�E
���R��ْ�L[�R޳P|q��ڠ�*�p���*�&�0���ا ����Љb.�k�l�w���X��V,�bX�z���Ⱦ+��0-���b�8sj#�)/J���|ZH���z5�#��V�]�ݫ���d��Z� ������Ky��
=x����i�%��)�-�,��T���+f�l�V�Y�@	�f��,��g0wf�+W7݌;�Q�q��6z����"$3^T�.�v�j��:�KW��6�-yV�ُ��%7��?�},B��s��}Xz�B>E��4gS|d��˯�g]{3.�L��Tv���1O�|�ۓ<�.��J����لB*������ ӱ���i?����%�g�Z T�Cۣc�u��r�T�GY|�j���HQ#?(^�(�dG5�Sj��jr�r��tw^%��k��2)f�A��O?��(��Q���*#IWq�L`�
z�HK��bܖ�jY��C%"wީ\��6����Pr���&"�3�_v�XI�����ȍ�O$�i�����ԩN���1%"kQ��>��J�v��kꅥ1����@�7�@k��e�$O�o7�g5��o�Dŷ;��x�$s?�=}���¼8��	4��W�>[�Ⱙy�wV5�b=��b��o��^�QEu4+%�׺�ɷ����F��]zC[���l�X�|E]W~� N�׆�m��vʊ�/�[����5H��QK���6m�O�\��<u��>�,��z��� a�z��=��V�Y2El�w�(��~0�E��c�`�1��y���ul�d��f�@��c��M}*W��w����)^6B��,�,�N|y̢�os��5;K��7�D�*C[���3�K�'

q)��5#��q`��5��UtI�u����d����
!��x�;gn��n-|�����T�#�>�V�3?�C!16d#�	6E�!/�Md`���H&��Ē�5��`Y�ĸr\M钱������nm<�X����WbE��Ow��ʥ��Fe]��l-�� 76G���B5�:�?���F��ǥg�hƤ��o�]��,�^�de`X(sa�t(J��!�$Ǉ����E*�v2��s�����q�x���T���+�6AE�QǨg�{j��R��]Q8NeN����gUE�6���K����9^B�;�-Y�a��y�5�KQg/N��.���
�q�����d//��w���u�p��n1T�3����lO��W|���׳K��l�1?��i�G�~�jɠ?�J�A �9c��M�E��ۡ��p|���3�6��ʀL��8[�^�X���|�k�Qt�8*Ut����۝��0yL��ͭ,�g�e-��l}�m�|xb䍑����P}�Z e7�QB_
ց��QО���N����Jy3��]� j�=�9�Dߍ���&p?�t�Ҍ6殹�y��%��d��n�)�X������lx(+�`�L�&�7ϋ(�e��w�"Wg-��5y
�vV,�f��jԡAw]O��g�lF�G�YmZ���%��0�3~˲Ra��a0���)�˪���L���n�m��Xyξ���]�������xw�kBhM����g��v�
��� �2�����ʣ���"��y�����ɚ��GJ6���ZU�T
1�wC��3�d��'!9c�p�0�B��GpP\/�-�?��Σ�����t�������y�]O,��H�����u ak�͉.Ȅ+?��/-L�R\f;>�y����,G������:R�͛}o�sf;���2,����
������{>(�5�����:ޗ~(
M؊-^��s���0wDΖ�bQ$(��ǏZ��G�1�J���U֭K|�{�I"b$�t+�v��6��P�j�jߣ���+��v^R���z@- D�B}�&���3�[Ġ��T�t�����9�+/?���i؁�r�ߢi�ß����kZ����a(�j��<�y��#�X&.����"��,p8�A��-� J��;nQ��׃9�4�nzB����	�}r)v=ԕ�T�X�"�.�<B��e'�WlًT��k����{�{<��m&q �@D�	r;�s*Hh94�տ�t���2�(MlܔPA�-3�}���']֗u0H*�Ouwi@QR�����}w�(�:�Դ���y��H(�#Ǣ["��Y�����0V����4Y��F�1�Z�Z!�ڎ��-N��h-5�w6K��f��7P>��Wr�)j1����k���O(Ї%�u���_�X�	$-�Wn��G�ɬx� ��0QFĦ>OTC��#���t+�A]A��Q=L�@"o�b�!ؚ�&�˞ B��[t�q��) 1�|������$�cF&_��������A"Ug#�t���8M5~H�������t�o	���|�-�#�m����z ��(�_O�M��&�C��E9�?gu�F+��C
���1�l�����ѤME�q_(�Q3G�X��#��%0Yh?j����<�y���>����S��åO]Nh����z��^��8 ������	QN��w!Fk `�M�j[��d����+Ȗ�t;�^��2�m�����^1���q[W:@�*�^M6j[j`�A���
T�r��Z�n�w�U8Ev�������pԷ*�$��|Mf��d�w�Y�Uqit��#��2�{��ً۴G��sP� z�����fj"�f=i�SOZtN�_���Ë/��d�B�i��JN�Fd3�Z3��B��4°��Ρ�E`�s������+�T2�~��:L] �"��`��?�x��">��G�7�B�*2V�Ñ�L%�,<�=ڥ;�^�
��k)�Q԰��y�Eo��i߂c�jC]���ޅ�6<B��j[��Zh��@�����2Ż '����P���ɒ�st%�X]i��N��]���׹F%��7"��.{P� &�2��O�C�M���BQ�5ihv(<��TRY�4�9����R4u"�O.�Rf'�d��q������2���H��P���h)��g��S]������6B���GA��ƃ����Bf�F�����{��h����CtH,�sj�O�X:��%x��ŉق!�����_����3�$�Qv���{�۬�9x0]�ӽ��`��=�MP�Z���M���r��\�����#�9%}�R}�m%{ze��*}u���}T���J���1)����	���/P�l�;tYUp����Ѐ/Ě�[^^��N_7�a�Q�?A8��t'��I�4�JpQ<`S��_@���L`1��� ���LU� ׅ��ײw(6r\��ʼ�>H�C�)�u�wё����� ��V..�Jy)���?aǈuE<�kb5��S\�7�
J��a7`R��s6�sW��I`cQ��������l��l~!�����ݟ�;.�5�y��lM��<�p�	lUPT�,C�.��:K�]�}k����O":ʷ�z3�#fQ�扲��Z����*�d��,��6�����T�4{Hz�L��Vb�,��&\����iP��%PcM�:�,��:�H?���Z��V����>|H�\k�(��Pfi	���P�^_24 a���,R�����zQ��5��2@��/���ee��D���hL�E�E�~N�\ �VOG�b�Z�Y��z��6�8�؃L����X�r�M���?,㼉ۅL?^�����Z�7_.�/��8�z�بg_	|KA
P|���g�ӌ�r�t�����!L]:�{�~R��-�f< ��%��=��L1��Tt�א[2E�������܁i�����~/��k����.deq���I��R-Ƭ �6�{\"	�Y�ח�:�F��K�ZD1 >����w���@j�����71%��X�w�&uXX?WL�������(�h�,#ӧԸ?�Eksn|�Aí}�h��`�D�rR,����������l�Gym�{8j���1"����i��|7C`8X�"+]ӶR �V���*�O�(�B�1 t���I뎜�#⋏��͐3cEN�����WR�û���}��6�y�� $
`�&F�Z3�Nn�>C���@c�y9��5�i���ɿiE��L�Olz�9��)�	-�?k'��0⬎��8ݠD6��[�N�eӲ���%�j!f��v�@�ؔH�)�8���Uo�/�(
�@Qی�5m{'=�b[х��G�o~��o�=�oq�!�r(�1U���X�9�m�i�~"�*���P��Iv�l�l�m04����Y�g�ϊ8+Ս}h_͏�2F��Z�\�+�/�ot-�b�P�1z�&ּ�����>��:E��]/�w)����}��UFBHg�Oy�4�?[Ŕ�XG��o��yeE��N]��B����j�����	S��:�y���$���ꪧtE�Ŭ>��y�{}�F�L�������U��� )����hs�p����b9��:&K�_�ްK��T�x���oti��CQZ0J�(%'vͫcD�U0��Ӭ����J�t��.�&.#�e��Q��]�EE�4[���_�Vu0o���\	73����+H���B��ܮ�]�uW���5���˘� ���U���e���UFL=h��X���_��H
o��9恓�k��ZOfF�`�'G3vx�ѬX��[�c���Z�C��_D(���ܧ��g�	]xP�|���{���A#g�mj��X�wS����a���E����Cc�)^^�+�����n耟���ߌS��5(� Pi0G?/.R���r3O�����I ��b��-�&i��55�إd���f
���H��㖱vd���f)����n�۰����/Ш{t�Fw|~��_;�4(�����s�H �o��SN>|5�צ �o����g@�C\͒��#��|�,%b��JR��F�6�hU;�R�fK!�KS��u��vJ�&[����|͆����r���׆u�R�Z�'zI0 F�B��fH�
��!j\r�q3���� ���M�$6�~��iN3�P��G�}؛;�R�>Q4,}�U�YDA{�*,���� dqUݚ��{�^\�����U�h)Qg�6��&jM�I@�T8BkpY�v��,-WB�6LS*�E����e��ϥ�a�y��b_c&tM'b�����E�纂.Z6���ݵ5�Y�ܺYB�2%�?3q�`�'��k���tB%_��?)���b�Cp"�<B����6��`��}%�v1�dd����<���Kİ���|�uԚrɅ#%�]�czD��ބb�u���y��U��TT���g8�-�f��6茏F�]I��wf^t��9Dp�ڭ���#���H���T�g�/z�e�SGaڬ�|�W �^��m�EG��͹)�Q�toL��ɠ�w�Ӗi�J�y<��b�H'�Mh�F
5�'��c:A��F~Ҏ�$q�5JwO����;q��aϧ�'�!W<�&.S��
d���ڇhϗbm!�.4�D�iqW��4�tDn����5q!�s�ֲ��+�OwiM!K� ����!��c�\zK�z��u�?�����5F�x;�=����=�.̃j�u_~������?�5@
=_T�F��]�=��� k�po@�)W�q ��|�>����v,2�^��Şp�jNaOak��t[�Bڤ�wzP���L����ּO[�"P,˃8�.�ɗ䬥U�S�
Te3VNW
��fk.�5ǚ/�T�������%L�K<j������*�pA��H9���Z������(�����#B�P�qeu�B��9~a�����[#$V�8{v��us7��E���iv�I�l� r���1֜A�s
#D��_��.*�P^ǣif�-A9<XՇ7@1f�I��àHr�㡈��C���P�霂lab�{ � {��!~9br(T�t�u2��]�<;�N�fI�}<����h%FQ��2�Ż� �aT�Er�/^H��̡'i������U��΃�ћ�7�<:gxס�Ŏ����x��aa7��H�� :���j,j����sY	X�U���2D�[�4��s�%qk��gWS�qv�M��+�/�q��1�#��6�L��d,=��%�Dd��x���4���L�քq[�ML��jj���{_-�>y3q�[���WA�,o1����Ő���S}2
����
�`{�ڔ����V&�yȳ��ob�)�הT�h�q�5���-l$�i��z0ĸx7��#R��� ծ4%n����4R�w<
�拨n��WO���F��b����c`��Xa=�^h�	Q�bM|XO�0vt�H�Z�����ǰ�e���3��P�i,���"#*G���y�煍D^{�T��`\��z�ʇM��H�˓��dձ}��G���Ȋ&R�<_�~�)ٛ	=�ʽېo��4Lz�1/�|G&�W{�<�y����L���ΰȊ9��'5�-I�)8(���N�������z%��q
["�p�s]}���B��e�6�,�%^!���3��/��:�>����<�Q>�l�<�eH�f,�^��[�.���j ���!�0��?�� Z�9[��`{ �A]���4�1#�~�����Ӝ����F��rh���X{ޖ߇���ߙJ#B�0���a����.!��%ZzMco����Wtk5�r���YV㹌aK��#��T�'磔k+�����on���F��M�����0�M����zl]:E� ��U��ݔ�t0��h�?� �C�Kv�(d������4�jqh�ݬ��s��	�+d$���yS��bo��L7+| �*譁�v�x��Q��+�ɡ�\�^mtdGgޟI#��"��U�V� �9���sm���Ҵ&�檤JQޑv���؜��̱c������Í��xO��/\�	Ni�;�� �]W�`�z.���B�Ԝ&���.�	f"��`�Nlj���Q���k�A��CGf�����fD�嶳�K
�z�QE�}�LP��sǓh�8�g����[�ۉ���D��J�;��VA@4u�,���P� �k�����
t�B�Ku����������P�    �k�!����@��&?Cs �FH�|3������Ȝgv�/�W�Xc�]�|"LV�PЏ"N����"֣����qS�����Bbmf�(�z=6y�&u�
�PD9�W��#ږAbM8d��^��iɱ��H�*�4<[a����Q�����3�*|</9�#(��B����������n�_�E/�)�x�?iҘ��!0<
�Cѕ�c���z�J�T�q�j��h��Xa^��aߒ8�ۼrz��tD��v�KI��¨��iC�i�#�Ŷ�>��?�b08$����R�e���6�)C,#K�v{���Y�����Q6��Ԙ�ɂ� J�4�G�nl��V�F✽�[j��R�g��XU�qg�����-��K�j���Ӹ�+zV�q�m��o7B������sA+�$���-�Aa��$�\4[��J@���	�I��j���F0@[u��*R�=DN��-�L~z(D��wB�U�(� �,T��?s.fLE5�a�ɓKz��E!�RV3���t���-0g�m�į3=�"��}n���Lr(-�_ԋ��:LNQ�] ���f����s�K�~&��§���a��,+yT�vBV�'��!����Jꊾ)�B��Q��5�*�X#(�W�+��UbQ�L^��5�6i��	i�E��6�������                                 	               	      
                                                !      5      A      C      P      R      S      W      Y      l      m       p      r   	         �   
   �   
   �   	   �      �      �   )   �      �      �      �      �      �      �              �����
                                  �  `�y�!       ��      ��      ����    @~��    �  ��ڣ                        ��      @�      �  ��ڣ                        ��      A�      �  Ϣ� ��[                 ��      @~��    Q  Q�^�  _�j�2                 ������  1~��     �            N�@�pVB rXB .   43E h%G h%G h%G h%G h%G h%G h%G h%G h%G 83E    .             C                                                            83E             pVB �7E     �3E                                        C                                                                                                                                       C                                                                                                                                         �         �       �  �       �  �       �  �       �  �       �  �       �  �       �  �       �  �             x   
      �`B    \`B 	   0`B 
   �_B    h_B    8_B    _B    �^B    l^B    �^B    4^B    �]B    �]B    0]B x   ]B y   ]B z   �\B �   �\B �   �\B                                                                                                                                                                                                                                                                                   ����&�A    ����   ;   Z   x   �   �   �   �     0  N  m  ����   :   Y   w   �   �   �   �     /  M  l  �7E �bB �bB �bB �bB �bB �bB taB laB xaB �aB �aB �aB lbB �aB �aB �aB �aB �aB �aB �aB �aB �aB �aB �aB �aB �aB �aB �aB �aB �aB �aB  bB bB bB bB $bB ,bB 8bB DbB HbB LbB XbB tbB 	         �p     ����    PST                                                             PDT                                                             �8E �8E ����        ����        E��0�pCd�l�)0d��f!���2πK���3PI�ap����U��~��r��"J�Q��g�x���~&O1�vAn�.��բ�����`������jm��(�1E�ّ���^~��AWή7[�`��{�x:<�ќ</1�q��Ss�?d��V���N���ܧ�1��艬Q���t{5c�K�"��(H��R�S�獁�D�{L!�y>��$�F{E/��2HU��f�P0���`K�Sg�c 7-�O���(]`�0?�x���ߜ����kq�8�h�p��������G-�P2Ў4���ْ�[�o�e���D+.u��ʈ���{�Θ�2)n��j��C��fGf��<b�{�";�Nh�9���3�꾺�����|�rA ��\�p�.��'0�ڹ_��-�  �sYt�l<�	��A���91�D�mqS�<h�8�i��@�R�����u���N��UV�x�pw�9����zǸ�%�OG,�5Q����z핅&?����E}��l	S͗L�v�j����+[�V�̨���kx�Xhz��zTu�FS�c�
g���]x[���a5Q�♶$�۟�ps�?I��-�W���|�#���������g�y�W�u�߿����� &5�y$��ې�wƙ�0c>3�����o��M�E���k_�!~�]S;�l���&R�����󕏰�hӪ�7�Cs� %!Ä2�c�e�8��.5���8��N2}�"L�!\ �N�׷���(W���)+t4fV운�d��r��P����b�E����\#���kj7�vX|�w�v˟O3�ވXM���޹������Yj��BT��kݍ��\�U����݂=���zLI+&�x�ɚ0�1�0аP;>6f��o<��5%cr�l6��*��'�"o6:v��ʟ�x��Ż�w�i�� �-�&��)3
��덵�!��qډ~K�����+t�v��xZ��h��^B"�,�?~�'���dt��٭|~��������h��r��ܻ<�e�=�,!g>������51p�
��+�q��p$h��|h�:{3� ��י|��Ś��<����L�
ʹ��
�%��f�� �;2Es�f�����3�T�Ӹ�/�t�% �),Q��L��e�|L��u9QrS$Mpi����� �%�)��t�Д�oO�A��YF�fj��E.����{��?����V.P҃&�G|��!�o-��=W�g�9Kt�m��� ��o���S��l��Ub�%cn%Yt�XW� ��J����+p��B���&�[�VD�nYO�{�M�PJ�w<�z�$�}�J��ߎ쀃"��R8xJ5�!EO=?�1q���g^�zip`Z�8���C�}V�W��-��Y>@�;�Sp��#�0����6O�R~�mL�8���y2��~:�����)Ņ�'� F]d'ہ�k;�#��a>�k�Rk*r��0H��KJT��O���	�\� aOy�J���������}�~�hT�	�x��w1:F���?��fzn[;2���{�f��Pr�?r��Ke| 3����̃�k���ٞ�R&�T��\R�Ɨ�e.+H�6E�eHh�(�M��h�;���pr�M��t/I�[8�Ui�Ñ����|i��3�j�ӿx�|�)���C�_^�gt��zر)O�/�
�n%�}��.���Cۅ�8���Fv��k��,>�n��7���|=����̓����F�e�g�=�8؟�iX�[c��pԎ�����r'���/ω�����K�(M��a"xL��v�S3f3.i��}���M��2sO�Z6DZ� 3�XӅ�K��;�?IL5c�I&�&�eNT��O%��L�ƏWID�)%#f�(��[�	8!$s����A���[���k��B�$�S��|�@zt\����_�Ee�쓍S=�a�H��;G�_-\����dϊS�(��f�)��_Fm��h���|H/z$5K��2�7�沥:�b.J�'(|lY �0��^/�(%T�+���R���)x-"ɡொa�l|���B�r�^)�,�i�g�w�>���3�&�  ֞˶��:W��R�n����ӊ �p�s�Q�q�����>�� *1�␇�8�rBV|A�ڍq�/�Bۦ���6�\^�a�t��(O�,�$�Q��WAr�Hi�4k�ncq��UE�RʔPǊ��*]�L+�oTP!z��j>��t�3NCc�I^'c�����.l�B��E�$,m����;e{�.U�X}�s����c�vS�n�U��d��5A��Pq�?Ƞw�U�gc��*� �N�mo��Oh���������:w`[A��"�o&�(�U�E�A�r^l��apg�	�,An`�I�E,�7���ٛ(���;�����FK�l��yo�B��vR> �`����������)o�k��&�����d�"'��L�K9�4\�����LEn��99��������k�l���B@�	��nea�8��4zYR¾�7��w��l��)��oŅ^C�4��'2���R�1��c��H��Dkf���:/��V�����XW��&�3��>�=XV�jV#�����2��.Ѧ�k��8�鰰�P���&����53T��0��="a����n���>�)�A�������T�����:��y��}�<�Τ�ܹj�<�fF�)W��&�
Sػ�M� k�7�ǭ#�,I�H���j�Ul��)Jl��w�|��G��[*K��? C]HƉ��1�V(�w4������Dz+�@�\R�X��X@ ����q��腊�b�˫г@�%Q���O.U�b�����ief離"%]z�	�̨E�aHX���[k⥆�ʍ�e�M�<�ib���&H2MrO�����&v�~�#k �-$�#��n�E:p�nMͧ|V,����c�sn(^4y�T�5`E���[S�9"Y�/��cJ �(z�r�����G=��0��C)gCy��K����qZH���#�ĕ�U�����Z�u~�@�����2N��a<���]�����\j{���ʹ�����,�s$�o-�K,���v*w���{?�i;���ZP-l9�Ũ9F^{�˟p �sdS�/˫E�W���p-=����!��`��!�s�)��L�3~x����r�В�s+�@'{��ϯ7$^=�,,?S���^k�B�x��G�O�k�`.C�?����j�ܠR[�T/x,��nɢ��#.�`#�Y{P����9�?�����G|��!�x`�Xp����r�Q�+�2a�j�� �����wJ�rJ0�ʽ�d�����|;n����g�U�8�G8�d��ž���a/w�qD�.ߑ��,nҦK|?���e�u6s 8a�i[]��"áhH�i�M0�s�:�%a)������B ɋ���tP5���{�e{�@��5~/i]+��Z�L����A377aW�E;��!m��I^���-h��>؀��]�N+�/�Z�T��K&�{��IH1l����TMm`�m��h�����%��S%j�\�=
�*�F[�?��	lו��ķ�N8:��
�Ww��L���yT���b��pS�v���m�0�gr2�_�~�h�Xe�W|@����tD��S����&~>W0�F�E���𥑥`+
���AP'���7��7����eD����m�Qs"������ס5��a~BI�������z|ν,��Z<Q��Cİ�Y)Mzao�ѝ[��x��H�"��n�$bۤ���≫w ��x���+����\�J���u�Y��r`�
��N;�v���%F��y����D�Rt�n�Y���힆�xW/���k�?���48��op�	��Mx��3^�)Q��*Y"c�`���(_\�))B��H���ӭA>�n�|��Z���Gb�>�! ���������&~�*���bm�~i�W	zZ�I�2�k5O����ř<<'yj6�O�����=�����kA�?��m<�C5I{i�d�ӣ��@�C5���.���I"ݦV����*��R6��z��v��Z���b8�xL���[T��eM����a��=��y|˺�4a43j����~��-�ݧ�'7]97p��X�J������'䶍���)  ���U�P�V�n��q�d�uq�V�Ia��l��] �(MՌ�k���2�����I�?0���T�S5��\$�ki�!����q��Yd�x�\R��%b�(}�q��1���苝�Zr�KKD��T�{��N��f��~�Χ{_
G-O�U�X�[:�>܉�%I���?Ҿ@������?���W����� �$��G���/=֖1��N𳦘��rB��D�!�}%2��T�}t�F�.+�+I�X���$E������J[HlK�Me� T���.�fwk��^�F\�3���s�[!�M�5��5��m ��Q��h�P��-�$�,8����\��!�v��ra{"��%d�z�~����8Q�P5
@��C�r�#�U�i�e��
tq_�>�<��p\�k����Q���6|�bŘ@�8}ԳIV�Jؼ��#B���>[�*�Qjf
}�b��J碌.q=�6�(>"��(s<�0M��;h���.k�[1�]a��{/�x�m�?�+��ȍ-�eߘ�v)��Ccۮ+�qwI�-�p�7�%�@�@}\����zd�U��v�(�����!���v�Eڈ�[�(�����fA_�P�Nx�7�V#_�Jo�*�/3��lW�����t�-c�w� 7����1ל�Sb
�;B��)��a^��2D���ި�l�0_��ѫ����gn������� �Iޥ%OЇ�l����;3p���٭�UZ�<,� #��r ͎���_~X�M@���_ޘ&�.cw��2-f/L���*���_硐'����rI��/�k�;;��|�t0x<����d�	b쉌���tH���lG(��an�z���3��a"K!z�� �ת��DK.]�S��m�d�C>�m��	oKGe}E��\,X=В�EՖfvQcE1ܿgF����l�UH
��dҾyp*�Z�qQ�_��XkN�����ԏ���Ԫ��[>wS�
gcdeCK�ߦ��V�*����?��"I|�T����?�
������h�7�+�,�n�\{i�\��(N��2�n����c��k"�i˄w�1�YS��=*h�^2��gu@C�U41s��� ��0C鉌�6�"���L�W\Fw�Q/� q��},�02���tX�ψY��=�bu� ��v4��D7f���n��%Qvn�G܏5��j��鉙�����]�!=M(a�~���N41�)��7�� �8�t��fXaM�w�7lb1�8�Ě��!ҝGb�;j���40G�Ӛr)��?���I&�OVm�]�yEI�ޏg^�fC��ѣ�{�1��&�`@ �7Ej�^��V�rBf
�B��͠x��9� h|�ʙ~H�}O��,��ܲ�U4򨣊�!�k��Y�i���v���)��x�,ު��/|���4a�o�(��Ƨ*Zo�è�@���z")?��$�DYR ��1��ԪGmﴻ���Ɛ:� �����?nd�m�-�_���Z;���~?4=kb�������^_ �ӿVI���V��*2�`Kt�� ���&�}T�������q�!�	O��+�8���uL*t!�Ң����y�t]��Sc�?
w�wU>a��\��V^y
ί��drÔ,^KӪ��k��D~��@�F(w�(��{p��.�.l+�D�F��T��v�CPɸ;���Y��𵈅1 �ZhP�v�%C#0�Z(Y���?��D���k~x!��#�仮L6���q��N�VC3�w��X�$���L�&w
(|�;e��-�z�8��=���|�z:.*�Հ� n��
C��Y#q0h;D�|J�d���b�@~���P���w�d�A-�OG|V=l��w�FVdly��X۵yR;�@����������`�NE���?��;զ��x��Pn�ow��1�+_ԑJ@qN&�^S���%2��%�H�eľ.^k�iB</>�[� �� ����7�Ն>�Ί3F��q�H̲��%�+�W��y
)��,4��X��t�B
�j��#V���.؟v�ź�55r���{'����_L�q�uÖ�јkU�5��ۄ!����yD��.�!���>��묐�h|c&�ܑ�Ivy ?l�u���K�����hA� E)u�(�r$�ۉ�֨���9���{��|�����E	��ߓ	S4K��C�F�6�I��c�4�C�jj9G������Ç1W}B��ok�����4�FM�y�O�s4�j<�U�����|/�<�{���J�a�9���K�����r�
�[Tug�����,��I��W��٤�*N6o��ƃ<|��bԨ�]�@��߂V�^���;f��aM&2��:��x"�-b8?Q����r/	��nt�.Q�3�G�.�P$�.��Cn��}��=e�p����e2�����Z�!܊^mi�����@K?�c���f�MSq�<�MΩ ��`�I�=Օl� Ʋ"�jY�{0�%4�����T�V�J�bƔ�`��]	��������U �
�P��A�_;��c���,�3��D�+�[�zh0��l��h�|t����[=�q�D@�Q���i,e�ካQ�6�tnh�B_�qAsO�$/�q���k~8���K�ab�hP�4��	v��c�������겲���gTj}Ty)Q1QGu�XռMx���Fj�"Uʱ*����خ+�<k�g�&Ӧ3���/�-3�ƔI�pn!�f�p+�cC���ݙ�zL�g���������NI��i`i������=%��be�Q3�f@�IH�6/�`����p�ϛ;��C�Úi3�05nm2��k��W��,b_���Dt�p����L�W/v瞯�I�?Į�:y��NTh��
�p���G���?)��8 �Y�s��:~�/��/��:�|1د|�}V�Yeh�ו���)����>���?�����zTε��8��^�Y�]Zoƞ� D�(�B�KC�TBE��I�L;�t��\{ʼ��n�`�d�~�/˱��v.��:�p��?�	*is��;ߩq��P��L��ut+%3����-٠k��M�:���\��x�>M��.�&Q��T?�I0��"��,�@i�_�n"�}�!gsw�r�IK��}��mT�9�Z�]`{X`]r�b�N��>s�N���9(�c^���2�j06��l'm�J�f�&u��_��,����s��F<����R�0���sY9�KiHzu!C�i�E�M7��W�f�W�)is �ϡD������.���9����6�*�:������tA[ya.���:m[a������%��w��ĺ����i�8��C�e!zaŧ��k��\gg���_��u��3��e�"ْ�n�^��g>����&��1�M�-�o����Xץv݌Ӄ�*U	�#Ķ�~�4�n�5�ȉ�0҂�823��G�>���O¥v�F#�_JdY7��+=����|�X����QV,V���z��z�r �\D���g�T,���㣗3��&�ѷ�ƾ��A�K�AN�\a�2���)f�.�l��3�$���@V�ͧ8j/�)φ6�?B�>`���5x|��,������;�,�&�D�;�Ifl~%rͪ�hm��b=������:@tϹ-�=ڈ�>cv*�V��F�݃����&3;�c�&*#�ݮ����D�񼿺���a��U�,�J�ѣ�9�!�����r9�0�ܖ��R ���.^����$]p�Po��C�������Y�KP�M3Ё�=rO��3��۬/�T�2��Y	6�߬���b~�|���tu�%G6�Kލ��b����rr�~��T���]�e�����+1��`�zVG�)���Q��mO͞5�QG��f�=��rIBƐ(h����-0*UK(Uh^���D�ֻ�Jn������%���l��y�a ��r� �]S�z\+��|����;A5���x�g�!5��������D���4q���u	���r/`u�����<�W�ND�$j(���R;��tOk���!��_o� 3Fr�r��a��^:Jd��"F��@�@��Sc�Y�������s��6��0x�I�^����3�h����ݱ+*�<���m̶37�@I�b�Z�v�����ĊX3ev�3�Cw����`������iĮ1>�ag�t"=��}�ѵ�J/�t���1�nY�b���9R��������N����]$1��y+�/�����&�S���W���m*���"8����Q���<�z��R ���t>��.���7���v8�g˱��_P7�B〥��ʶo]e�&细W��S��.־]Ԑ0iR���WD���/��h/��E�һ&ueS�U92'Dy�7p��
���f���9�&ezQ/>��� !�N���Pg�1�����h��W?�9�͒���־�-G
r�Q]����G����Χ��
V�L����Y�qo�+���@�M }�rG��3�1����M4㘼�'���ˉ����� ��kE����F�$��BJ��YSWeI�"�`�g/�Ǆv@�
�Nh��vh�L6P�+��ӊc4�o%r�����|��)��m/��;y�����/�����Or�����-�����M���dc��p6Z�����&�$�ib�M"�y�2���������!L�cct��y
ozėa�?�I���BV_�}̿9	��'i�.����d�I��A�{xYv��mP�_ݝ<��+���s�n̯Β�Rr[!q����ɡ[#�!d����EZ����P�ۨyDd�X$��V�<�H�س �|��o}�L���Z^� �,����f��b�r�g���0gP:�����	!���žu]�wk8���՞����=HU��O�S:P�"�͔EgLc��f��s	�%�LL5��*	�Y��B8;���|�VeA�24.O��y�y�f.6r��Ubv��"Nu���˫̾j@��x���0� H�לR�vm�2a�=����gw@ͳe�gA�E:&U~��6"�dp�כ��z����m=�#N�[v;�ۛM� $�.��P磁�*���QL�&��$oӮM�hvC�`j��,3/�$c��3TT�%��L4O�c�,n-֡ r �l27��S�:k������Vc�ż��}F�8<M۠�vST���]%.�cPz2����F9/q~��������K�f�P�fu�"�1����J�S���E�=��_M������°"����Z�;q���8��`���']ͫN����OgY�9k��7F�Ɖ��@.ʴ+kﳕT"�N���cP�(Vy�V��A�f-�s�:�=��������^�c���v�"L���!n�F]Q<��7Q���ųb}CSk�&iMN���>r�m�鳓Ejd����	)H�^ F�MQ�N�\h�+�V���=G�I
���R�!/����W�n(�q���P�ߥ��U{s���,{t�}�-/�r���5�r\(�N��|�j�'OZ� �ݵ��� @�D���@!.3�#eN��9dj1�1 ���\*S�bn�Xb��^�p�b�d?��2b��3cz|�y�)�p�M�
�8�?my��B`�� �ɫm:U�U�3���0g iIE��B�'�2n9�zC�.H�`���>�rg���{�]
�^V�`V5��0ǭI1��H:�8������b�p�K���*}�
�k0ˎ���/���W�
��L�a̴hn�Ӧ�U����X�jV�M�����iZ
�>_9�ؓ�/�����/�ZG�f�� �J%<��^Tg=�����ă_�˂�-�Yk�t^�u��k�;#��$���5jw_����ůmC������׃�]�/�[�\�Qm8Ȏ�5z�q�����qٔ�}��.�7҉�Y��O��0隉�����ڄ�iU36�r+À�����ͫ��>*o��xN	6���Q��P���r�o&�!��J�����ig�F�� ���^�7�z�d�&�u#8��Y砼�"�>�+b��������З�����Z�]Ì������+A��z�`4�(..�w��/��\k���Q�:(�H��@+����2�?d\#�[�}>$A]�pI�e�u��'�\���ȡ�|?V&�f���gƺԸy�l��UC�#�a������)VO�q�����*�L
J��
��i� ��L+h����|�u{�r��`�׼�Ac�h\r�J��b������$L<�f�C���zf|\�"Ų�m��F�<BJ�,��Z�2J��e�����I]{�1�R��� �4��m��)�k��~ ��{\ ��>�{�jE�� 36.qܛ޾=��:�:��-mɋ)����|��Y^
tD>���^�ߤY��}�=�X
��c��%�B��c�D[�D�N��d�������%�*ޱ.aq��}�@z"9�G����1x*A�V��2"u�\AĠ|w�!�)��"�T�eIw��s��`��Q�"�J~�R	FH	k��C��f���A#�%L]�������4�>E���]����yl�����5��J�kP�l�j��3�o�4�{#�v�3)Cz�1�,+�dLb�X�R���qM6nb��Ѯ�������3W�:f�I��*�Q���!�
�_<S�l}K=���Z��-	�y�(�l�#���+���%�koL����-�R�5A��l�Mʌ���ٷ���-�t��Q5H潓�A�A��O�gǪ<��]�pT���F���ؽ���o�3�>�Xr�-ہ�u�E��5���T�@Mcga6��%���p��lM��]��#F�_cq��`<.Z�Lf	O@��hv�-t�rP�k	B�h�OJ]���qd �gOOQ���[)>L>w�
.�ո�#�\���;�C�5kC���Q�jh�t�39��|�8��!%�]3�r�M8�<>����]�{>�ϛ.ݓqH�KV�P�n�J�?Y?�T�~�?��*R��TSP�r��0X�h�}�&��3	r6����Ga���V){�����E4@�w���c��3���F��/��hz�{�Ւ�"�+	jjR
����"Z�d;ќ��:I�*���5_��`�)�~yc��B�P����-Z�N�V��U�;��&Q�����>h���u+{����B�j�'W���Ņ�}�_+�*�Ĩ�s1��i�È�S���q��7�����&�Ηx8�go�ʂ�N^J���u���ĵ��P������l�*v�n�`�I̳�ϵ5<1v�waʊ	~^̟P=S7l���W���FxR�˖�'(I.57M�#�B�$oX��=�Kz �L㉯$$ՠW�k��R��f4��R��,$RFR-���3 �)f'[h! $���!��j7p�2 ��<*�3�L�?mԕ��U?���<n~��n��󧼼��Kٝ_
ʲ��j¸'�"��u@����7���4s�����yL�i �o;c��o۠ x�BlB��_���<�*��S���򳡤�'00x��~�Upۘ�|��X7��j��"���*	�x�Vݚ�������cyX.. ސS��j p�$&��7��$ ���9M�}Ϟ�W�!Ц� �OL�2Am1&�%�v� ��:�����߶s��R�2xD��Sc��8�
)3�\�m̻�����t���q�F��d����˺�Ƈݶ����"��
Ѥ��
W�6��N�MV9����q��Pu;^�uMW}���]?RPS6jw��Զ*�O�^ 8qӉ���:���T�4B�Y,[1 1�סJq90���`ب��C�(j��H��о,�&�����2���`���k�"  �-�_^M�D��g���ȅ� UN��;�΍]�o�Z�T��=B6�+�"1�q��v86�\ªR=C�Á@"dn�N ت�k5�{�R�e�&��'�	�T:1w�Fh.��.�0�C��q٬�˓N��0�&�}se��,��?�a�k"A#�%��k�5�Ks�w��/���UYoʴv�1�U5x���/I9v���� J��B���΢Z�CO%h�(F��"�+Su�<����ǡg�_��ꖫ��Ӂ`�K��H��+��fg�6�gRU�ڐ���M��^X���3�>��/�z0,ɬn�x��׭ɸ��C8M����#�\�^L�2�ܱ��^[
����l�0{0~r���ȁ�}�V�.��]Ԝ$v���a�A�I��g�a��uȫ(�5m��Z�v����|y?�+EOuk@�){e��a(E  ���<x�Xg�eq:�e�����
��٧If�,0*2;�*w�i
��D�z���	tRƲ�ɗ�u����޿g���@*5l˻����y��c�/�YS̟�o���Y��8�lΤ�59f�,_��=����"j�o1
�݅��<)_#�3Cz�]�w��P��)�~FH&}w^���E��<&���+ˉ�n�܃�.d��j�阙<N��.7���k��6��+�(�Rg~���rjݤI��D�	1��	m_��F_�\B�����(�o{7�7Y�ג#[0��!/.�Es���$�t6l��{�o#�����x��������b�}�ǧ�vûZ������Lvt!q�;C�O���V#|X�ٹ��p�T�&�Sj�� {��ʒL�8Ip!V'�N#��&Vts����pT��̽[��4�^خ�6~2لU��������s��$�~�QN�j�'0+F_.7������yt]GY�1ij��P�x릷l����e���P� ��Y�>5����~D��N��*J���ZAR�'C�Tս�)��]�𘚎�Ĭ�$����o���LHG��C�r@�RߤV�6=�����zA��M����J�C�-��)���o7�v�e��l5��T@`&��%�zE����EfL�'+�q�]�?$�C� �}��x���lm�Y�^�/���<�?N�=7��1>ZcYjEb&���<nE@pf�V������*4�B,�"�Z�����Y|�]+(S��?�t���s�|E�bT8����J`M���p~�F�z��mӇ��@�j��%����	�ց�W#�E�M,^�H�}�
~a�Nv�N�,��54�x-��w�Z��;���uq�^�糴����oEԆl�y(��B+ׁ�^���J��{�1\����B�,Q�(�O�"�l��)E�߳��%/�F�.2�Cß�!Ԉ|M���YD��8�q[<�F�f����Y�$w�V� `�G�,N1��;��Ns~�i_D��OU�P��c�&fY����
F2��)V�xk�(�D��'�^�}uzJ��hU�����#bɋ�žE�ڡd�p ��q����L���]�"wt%��Zy�n��;\7����+����ո���~�zᳲ��~!"�C�(%Pյ�[�J��Gv�0񜣳}!�6�\���ko�N&ˏ#�&jṘ�Ae��7{.��u�?�U̹SN��M�Qˎ���M�z��ʙ����5r�)f,�;s����W�� e&��PBMM���f��V�TLۥ8{��퓧n�c�� ���70��rq��Ce���p&���J�>r{h���,"#��D��	e�t訵�%��Ui��$���s��lN�AƑ(a��帇�bN�0W��Em�"��%�^/s9s3��!�[�}Y=�_�rz���f�WH��h|�n��;��W�{7���:~��%W�-�X���͝f��|-Iz7�|̽L>���	��;;1]��(��MU�e�B��Օ�Eó%v���?^��$� i����O��5n�6=�E���O�xן`�A8�2"Akt-�b�EO�B��
��[l8,լ�5�͟������d�A8��EA�$L9�*�r!�%1;I:���1�i�Xr�<f_uTl���v���W��ѯ�ex%��z�.�1�.ޓ��NBE�/�������J&T����o�����>�V�L�8uH�R����g�C���Ѩ���9K��W���Z�C��m�|&I�I:��Xl׽���Θ1��X}�bwg͍�z��Ҿh�Bݣa\Z�˅ �{������������꜉�#�<�8}K��7+��z�9��D��|?��/�x�?���[UV/h��Vկ�#M�x��Ю�(�X�PQ�Ԋ��"�<8�v�)���g��tr��!m첒oR��J'��WA��FD�8�Bb?���U�  �^2jrW�ϳ�P��|���|"s��Bw�89�p���>Z�����)��8yNc`��8�'S�|od��"�%I�%�����Q�B|߆/dc���c�=�J��1�Y/�����j�g��xK��DZx**.�G���S��!�բ]�Y6�#�A0M�H*aCHJ�P�٨���UAO�QY�X�˯�r��xƾ?�ܢQ�lI*F�����ꤢ�ҪAҾh
X\�N��ߚwFL� FAmNx᫔��՝�9Ì�7(��lYgA_�!^�a� c�\�,�B�ۥ?1�=��)sX�딞��Sm���+�4Ğ�}�K� ��>��̢w<Q?��ez�~ZC�1+m�7�:�}�D��A+	�ue�8�����E&�F|��Đ"C7]V�,�!�Y�Ǫ�:�4Z�-���q2� ��[�)��R����c�[�
(io�^����]-�k5=��rTk"���\��46�&bv�ܸwj�v���
��1��[���x,a&(-�6��(T���$3E�����uٿ�+��U_W��
��<��S6�<u�p�IP4�֥L���-�^��ś���:B���;�m�P#����s���p�SՂ�A���z���WQ�`���D���EZt�=�@�OX7�CҬ� \��9L����b'S4[�2>�r��(q^)[��H�5�(�o�OיT�`V����緤�)��r��EG��E�՞��C9Wgq�K��H�~�W�!�t,���,U��=1�r�򔈓���]1b��'V^k�W���~6��0a��;� �0���j:�P�tc��fX�Me�,ݎN�0�ف\,.}�?�r; �"��[�9N��� �ii�vx����K�%\�6s�x��P�@+��p�O3�;7�'0�L4�̀Eg��2� ��.��R��<Erc-��I�p��Φ�Oj��RbйϜ$���cAR�����@�Pw$E�ؘ��z�Kg�ȴ�������Q.K�b�ݯ�h=������]�b΀ɍ�{uX�%�s�m�.]�v�"��<����RR�?��î�n�h�J^�@x<�N�����Z ���0y�\N �V2;�{L�'�{�$�^�S1�����U`b�����'~L�#!{�����Q� aK���g2a1uyu�ܓd�ZB8>U�?�$;�g���U\�����5=�Qႀ��s���΋4�! L������Ӧ��P�E[)���҃�ɘ�j��v�<hY�A;�_G3�&�7�aò�v:f�폸����o`Z��r��ql�,!Wm����$�V���s���
����!�s�R���xѱ֊vuk�"#8Q��6�]ղOz��o,���H-�Y�G��%eK��$�́�}�"��{�l[�l^,$C��}}̬�Ϡ���ߖ:��KV�d,�5�F�w�'��0휴��"A5t+�V.�~�K&�'<3�CYWE?���?�l��qԔ������-���&���:�O/��P-���Eu�|~C��}.s�5V:X+�7q
�ݳ�	}�0�|�杇��;=�b�j Wr]WWӅv#�)��I���<�Ӷ9�AJTÒ�ZMn�Xq|��W��ζ")���X��p��7?�uP} �@��E7$x���K��v�V�#�LJ�=�A��J�����˶�T�^r������<X=z(k��Nѓ@�'�Q8����)���8eȈ�"�@��$��O����s�_��&v��F���2˒	����/�+�3g3�O��|%e��'_@������Ma�/1����f8rזQ�	��܆�WpE��y�J�F��"k_8ʺ�����\�^�8�q�nd]��n�M�-ҙaθ��3� z|]����.��#	GvP���1��5��߫S߹�?pn�N�$iЍ�AT��M-�O�� ݊�T����d�ޱ"���<p�*�d�2�S�{"��8BS���&ٛ�g��ƚh���>�R�U�Ɏ�z��3�5���{�.���\C^%�&�W�z5`/yt�g�ae#/�a!�1,�N�I����@�flV=�>��Xx�@J܂E��ɐ遲��4���!��p�C<��%���E���G�Ӡ_���n�zڮ(���;�WM�1���J���H}�J��gȿ��6�J�����96,h;�8�)H��p���4ڱ��I«�My����l]�uE����j��S���Ah>�]�t�"����6W���9�U'c���/p�;"X��m�[�s�Sᙊ�R���v#y���!��2%�[���P^�ٔ��oܐ��T�lh�a����&!�g���侀��L0���qR�h�t�G�D.���,�4D�>���� 2.#^�/G+s �W^���Q��Xfl�Z���u_B�jz���Λ��:{� ;����4���Ҋd�x)t��e��\�쭿�db�� ;Y�}���/ZF%�L�+1ڥw��*+:������ĥ�D&��3���n��I�58�e�(�Iv��҉AfH���Zl����c}�.A���u�B�{��*I�r�&�uX��fٓ�;CK��sd�j�v�g�හm����C@��D�/��)ZE�4���)	�o���w��V�<���p�K
f�S�]����Kl)�ɕ���o��f�
!���x˷�p0�&�KrC*�~O0��v2R`����I�5��P&M���DP?֯�N�팧��
?������?���)��"�R��bm�#�c�*[��{�{�X�8�gA�J/�Ie�-��)�d�Kn��5�^�g֊h�]����[�J��y��窾AP���x��N!�r�ڎ���Xk��?�[�,��h��l��T||�+@�0ξT�ɺI<��Z5Q���-����/�9� �x����n���DE)a�gȲ�HX��!|������\$:�݌��H��1w^`z�a��v�n�
�>�uL�����Ǫ�����xo�.2c�B�)�g�=�O������t=�h����.�ة���p�t2���n��bE�ד�E���&k�)<�l?]�q_B�gs5�%�CG����{��������g�vM�><U�n@r�ʻ��ov��+�(?-��ΐ���T�3WU<�nx����@�[m��*���C�#�,pP�v�D��0�i�HE8�@R�&T�����ȱ�8�ΓV|�1lwś��������F}��uwC㍆��ί���U�}��vDԏЩ�{��<�Q�);L��1�坺��fy1���%��|Ia���fH�2�z.0�����D�[���@݋�=���Q�
���MY�_:5;>S� �.������	�(�⧴���Ƅ�
?E�Õ���(��������*
�Y0�R�h�-0�����8Aߢk��϶-�_(��zdF�*V~�i۩��%c;94h`3��qum=U���U%ڧ;��c����0������봨2&�y
9��o��{{�����:����4������EIv�������)�De��Op�_Pn��K�r^6U�T�󷱰��
H�L���zO��pA�s�̻�K�1�s����b����.h&�jGќ�1M\Tm[n�~X�����b���|�(N�8ϐ>��E6���^�xO��4�f�.��7���ڪ�~�ʄlc����..����sM�z��Y�Q�E��c��P�aͦ�BN�kݿ��8O�z�/q�Ш�
MuUC�ĵ�4�/��� �D'��#LE�������А�̋���Vw�}	����=��� �nR�-j� �!R�3�}� �5�P/�i���He�֜�ϑz(��2RB���*�d�j���[����J�Y(��X�Z�u���^���ZvR(�JtG(�#�#E�n�0W�|93���+�U�mn.F�96�l�������1o�)�đ�/U�����O���\n��ٙ	��$�-�Zk!���N�F��:�����O|��}�5��&$���x�i^�d�A)7N�b�U�`�&��K�����։�9���������ۉ�� �����Wu^T*�z��b�����뎎sW��@���	���u��̝�C���'���v޻?3�O��Ys���>�Ρ�?n�<暫%�򂭃"�Rb5kL3�%
k|
��B��'_�Rn��G�=�4�6G�1��N7-Y�wLr��n��5�=���W��q�Kr�C#�|O�OGZS�}�����l�6�	����^R���}��O�}���0�d��iZ�I��''-LNqWݶ[�j�r$V��b�b��$���jo�o����S�{O����^fl~��A�7�	��`��\�4Ao*���t��E�\��w�����E�<f����{����3���&�B+��$���ՕT~G�~S�H�MWEla=�Ӯ���6X)2���`��
�b���=a�W5!@���?ڪB�0}AZ����n�
�Cv2���5/.��m���xG��P!���,�EQ����0���J��:}8�.�ٲ��{�ٶ��\"�B�����5��&��=����#(N���cᗨ��[	z���W�ZM�}�铌+�U�Ka�]�$i!Tׇ6��Z���/�{N�_��t)���aS M"&F8�<>嬘���W!e�g)i�T�t]��_U�*��@;�y,�6t� �^�3��J���	����K��8癸={���P�SUo�ֺ���%�X���
:i`)��``�I��}�'�־(`�L\�^`�U�|5	_y� @ /0>�]���y�s���o~��h�1��:.�g|xsE�b)�\�tN'��O�n�o�����!��e mj`�T���w���i �IS�G��g������>w��s�*؍���KL�)2u>jw�>cXX�JJ�OH$���c�WA ����t�?�V�C�+p_s�z0����ہ�T��;��
G��;g�:r��I���E�1���"��W�ns]XH�&G��$P��yp��ٿq���2	pQ���X�����bهS��[l�>:���-���rA��'�.�B� 2�A�l���. �Jt>����+a�б����Տ9Q���h��q�!��v64#��`��ڼ���U�!Q���ձ{J#�
��D�vZ$�:���6�����o/����4E��Tۋo���^+Y�x�t����R��;�o�еM�w_,)�X'6ӭ��W��g�uƯ�/{��0JHT��X"��!�یc�է���)�ZIW�3Ph/�I4���[�cG������;/�o�iH54�}��O{ɩ�r���_�yu^�si]��u�e#H��O	�M�
ul��<�I_	P��_��������C}4�s��(~���H�8R]�ys�w��k���c碭�%|߯�K��׼�$S��q���>A���lSK�Gh�����u�+���z6��j���!����i���2��:�؋=�AG[�Y��������f���̂���<|l�/�p=���V֫u��
s������+9��t�[en��ku-��;��_u=�|�$¦�a��H�=Hʢ���������L�r�ǅ���(�s�//�����_�o�<�/�����Ic[���vZ7�	V��z7&o��1�9n^���z����NN��3�����dq��^�ݮ+�r���vs���)Z�}���'�F.5M $��qD�����N�a�L�e����,NGs�Ao��xۥ�%��K[�ؚN���k5p�qZc�[�9#=�j��ӊً1Lu��}�Ŝ����{ڋ�[��v%�ѯ�_���4sp{�(n*4���w[S��Z��a�_@��{ѵ�ee���^=� �S��A��8�J���C�ؼC���zĭaD�7�C�aP��f@��>ɜ{�h�����Tfa8^I����-k��$~m1���x��Ư��> H�<��-t��xdحtu�8�����AjC�F����ꞹz�<8̆�&�bN<M��v:V�o��T�
_.WJU�ª
L壟[D�S:�,A��4v�8yK��aYN� ���q�:�:�=���׌ y�O$S�^G�l-}�UN��z�[��-):��sSJ���)ͨ^ͩz p�?#>OG3ǁ�o�rD1��ķ ���د$�[o�����-~14�ZWVC0�v[)�����BDz�)�rY#��)�:�	<_Qv��p���A�B8��=�)^'��5�����a6Lʭe��i]��a���סQ��};L"����`GW����˧���8(��L�e��\���
��t��/���Q�3�f���2ծ怨_h���1���F�.���l�����j�
�cu�:��إ����X��)6��H��jw�A��4��q ��Z��a*�� 
w�Q�ǁ��}/�d���s���)��"ю�'2�(�J˭D�/ hk�s�fڏ,Z���hG�B�>.�����xsǡ'Ľ������_,�B��3�R��W�Z�w�r��O:�㫦2�|�-��7�n�xV
9?:�S������P3*l���ɐJfo���Y�$Vk��8kO]9d|�=7�KD�c�Nn�O�MFh���Go3���𝿬
8��)S��f��h�P����b��y����/��?�Ŷ�w߀e��Hfk2n��f�]���fn�����(���"�P�u&�k h�ЄǴ�{J��^������6���w��M�>�4�>��;��P+h��ޕ7���Ц�� �?��7�I�_�Ru��4�9�������^G�<)�P���$�� �p_�����8���T@��7��yN�̴��?p���/I,�z/2"�@[�ǘ�;̨���5�\��)OdGO�p`y�w23
�$��C�&�&7�����_oL\uP@�����Y�@�@�B�����B� �(o6����P7�~�3���������
�y31��T� 7����H�-���^U���W��ŖՐ���d��D+LD���~���[JH��ka���*[�d�PYy,���G���\n �]��0�V�*|dr�lN���F�<��l���3�ԥ��Y��8����td�՜�X>E��1��B*`�&���.w�l9�L4����驂�6˚�a�a#3ix_Z1��5���1��F_`x���cA���������ҀLT�~�1��E��JJy��4-�Մ�:�;3��?&�p���_]D���3�B�Z�#z�U�{Xk�C�S����{j���{�1x!`m�a��K�.��"  x�0hh�9�pf81z��L�f�U=�w�$
S�Y�B;���f�Yߒ�<�H�Y,v�N��8�"YM���T1�\�I����:^�DŇ�pN]2�[�Y��i��������1i��~{`m�Z+z|��� ̚�F����s�K��=��[4����G�\�%��c�Y��Ϩ��>*���T���8&�e�j�0|%
�U�@����|���L�{ K�՜�v��U�'dNBV�6��ˈ�Þ�WNW3���k��
$�Jc=�E�	 ��}qȱ�P��z��2�#�	��w`��/������hê���%��%�pʉ֦ʌ_4�\ى�0�̲�F�o�AH���Jmp?��O�j}F����}���<�"gw��aJzh���c]�D�C��}��E�;da��� ��h��>�f/.Bn�	���s~t th�]p��--��y/���Ϊ�U�U��׏���C��״�?!����7V�R3 ��~U	�2�l)��=�fh�W}�SG�-���T*l��Û,_J�m��\m�~���*�(=m�l�9ݤ���%�7�������������HQ�"&���	K2��F�Ó�Q�t�綘B�<�i�"���e�g��{݊���>~���� �}I�2�a���+�pY��H����������&"M����u��N����Rᇿ��
L/-2��w������7`^b��`u��v-a���tȮ&]^.s�*)~ˍ�<�{�I�ĺ}����J-��x�ӳ*�W5l;gs��]u&,�vR���w
�OPR�:����+�=r�INCd}�1��*��3i�۬���y� CT���`U�=ax�2A�G������,xt�WR�JK�]�WgO���Q�|-�
�F@�I^��t�7�6�G�:��P����娟�WG̊ʉq-�#:��x�"#��e�-#���a���Qn���0��� !�vo�~������q��: uL��dB��K��e/�����J$C��*:�1��מ۱}͞,� ?�hD��J�c��v���*���`J?��U��N�NJ�mŽ���a���,�с��1�ꏷ<�`hG Vs#`��q�ݕ�����C��T�C0%����E�FrL0����k�);i��T��yV�|fm�~���]��c��̼���&�$a��~�6i��8)|�o�Xd�R����]��CfZ�V'��į�e��u�,�v�?/���U��1�6��k�x#���I�"�h�f����KK-U)��Rs�`���ģ~�X�w�]�X��ԍ�����Uv�+�*8;�50����d�˦�/u!Ѱ9����c��IY�#�Z��!&Z�㼇��Ҹ���\��m5b�XQ9��}�Ͷ�u���hb�zڞ ��w�	�g�[��B�8Q �o�j0~Xe;���;$%H��y�7�|7��vI:-!x���#s����h
���}�9�Th%3�A���!���� �K�ި!�y�x���H��o��4
��_�,�R�k��q�֮ 6|Sx+������No1�کôI�);-� �M�ں�4�X�*�h�ko�@HX��N8���.@�0��A��VY�`��s�C�e�p��qa�
JG��w<��_ʽ���k�t��R�B�yj"�u�ߟr�����"�\��#&r�q� ����m5�3���e���ioU%���Ic[GN��`�OT�}��+�(�Uĝ��I2���|�!�e�g)"�R(��Ɠ\¬U҉�'�2�x@�!M�(���[H���"�"WV)n����O3�CMa�^6�n�*VoSsę���i�(]냇J`��5}�$�IUL��'�8|�����0Շ4'*й�w^�F��T�9f�H9��)x	\�Ұ������rO�V�irR0�<p��t��W�����.0$�*5���7li��/c5a�0=��NAr�B�]�))Tz
�U�q��-w��I&���C>�0��zUA+�:��w���u�{�Z��Fg8�,7�s�E+��q�����:z<$Y��VUW��E�Y_U��aD�/>���i��`DvЖ�|QN��ϕ��:�7�`ȶ^ �H�G�wTz��v�8{��r�t�mQ2-I�pb9������Y
4�=�GK�K#9D��n,��:��Q��ͬ9_��V�.�%ߍI�O���^�U$20s��������i�ɵ�l�b�l:�����֥gW������NNOQi���J����"~�v�����B����(xW�5��uU�l�'O��T�$�D%�NV���1|�^H/z	?es{�*"p-�!t�#PP�/\CU:`�$(�#n��̔��=9�7h�	t��
�S0텾ד�e�q�}*�1xC��y)�gو�8� N(n2�n�Y]�j�@߈~�����'��0as7ǘ�aV���1+�:f��	�-�}�BI>��֘O�b��wHQf�
س"���@[(�ߣQB���tPڐfάR���A,2���_�}��+q�^�o�	9��Rʪ�q�N��LJ��v�M�4�o���1�4�d]S�6��gdPtE��G*�W�_|�Ò�d�S�J��lo* �z��8�j�j#�9�<ȿw�>ć���&�:��;$w��p�J��cP]�K:�QΉlq�����A=j[Z"�h}���s�#�e�ؼ��� ���������.�f;"?��&/�:����Ӳ��E���F,X�+K8��S"#i���������<�2��-i�����ג(���ɑ� ��ß^&���&AUY5�ET��t��5-�<�0`<ݽ�>���WS�T̸�Bh���݁-4LS4�Zr�CzX,=�
b�$4���{�}V��O�3}��b�T��)d�b�A�dD���O*����e$�'XK�ۘ�P�OPcچY���i�rG��[4�U>(f��b,s��k��G�1s���<�N��P�w��Z\5E����l��S?��^�e��.f�M4g�<��P7NA�K�H����&n������c[�����ri�;�%`[�5r��}��p����⽞U�x7���kwI>����up��g���U[k�N�o,ߵ�?��|�W�j�z=���!w�������1n�$�&`��M�v���M��$�0�ln4a����x+Ӭa��2� �1*�}rGW��c
�:�_��O�d��(C?<.���ȗ9�K� ��g�6x��e����X�:���E��U�g{�<5#�e�`�q��n����}�w�Sߣj�l����n}�䣖~� ��ثӿ�Iݤ��1���(�VA�՜K�y�N���_ZnS�:Or���<��Eї� �%�}��4��U�7h�g�T��Ǿ�դJx��R�i<�
���%�0�(�%(�H�g�m9�6���a�3u�(��Ef��n��LE�G�Մ��G�}iU{"n�G����q$�.3=�*uD�H��~d��3�)��t���,�o��ǗZ���.yKݯ� �}1>�'�gR��N77����[;��?��m�/HJu��>�Zw�M�ݟ��n���K�Ҥ!;�l�H�"o[��_�66#b��-\`ߡ�I%7��29��n��bC�a����y�N�JI��D�ig̀��|K�e]����䭩쪩f���X���r!F���ڨ�'�TV��{W���X�{��^�)�?�;�e�����&C��}���f�8�+���VИ��}$� �ٔ)-4��M{�wf�f��$�9!g�"�*M7Dwx���_k�����u/��<��{ F�;/�VT}��,�~5'��`�ʈ�D�4�6�+-=_��6PA�TSF �r9T�U))���U�R�n.!ث������`X�H�*��}d�2��x2�)~��7T�Gt|4[�v��5�)�¹M�St������b�D�����Ԣ���g�ᙵ�L�GAo���2*�^M:"��hY!F�(��T��!�	�9��WH�ٟ[#\Ӂ��I�0�	���wX��{���"���P:��-���ܵN)Kk}Z6�����N�v�7�k��;�S�传�,a.�r�h�bL,h˗g� (M��O�3���*���cP��N`����g2����k�Ϡ]�R���C�!�D']�϶����9�=~=�i'L�����E[�e���n=�hs$���zbS�3t=�&��f�"�:���I�X���"Tv��ޢ���sK z� K�*�C�Jd,B���vlX�~RLL�l~�۽$xХ�0�!�tR�rs�ۮ���_�[ܭ����u�/?ʿ&�"�t�h�ߡ�e����-a�ă��:�2�%�b��]��$C���\r��"�9��_`�Mw{���$�1 7s���<ڀ�#�����c�t�Y��aN�Rp5��!�P�tŜ��	�6G)�pr9�co��r0`i!L��������ժ�����Uf�8�����A��`�l�|r�It�/�Q~��h��':z��9� ����<�Gp����;���]�+�B��sUt(ܚ���v�����S�SD��ۿёk���(���g�����d�ۖ9��Yg�&On�s�H��T8d�Fo!2��H�)�?�!��Lcr��^e�c��=� Ͻp7p���y�@0����<=;��P��r&I�mQ�/b֗�0O��i��Mꌫ��J��	3Յ���d)h%>f7()j���� c'��.��Wy��ߺA�3�K�pK%PHo��d�2�ؕ
 �;��3������H|�h�̀P��M��Ja��u�ֵ��aU�D�W�������艰���%).�Z��?�ƢCI!������(`WD���'�|]�@OpA�gǵMx�]�h֗�l���Q@~$-|s�r���٭ �*�Tw6n��n�`���]*�o(��7�g�l;z�g�s��Y�>S'��l�W��-��B�s(����yU�nm����`Wѣ諣�����/�t{g|L�oː���7�t��/�4H�5��|l�h
�TBKN�i�t0X�mr)�M
�>͹P�[��&�ԮQI�c��Ioj��8K��N�r']ړ���D�,}����i$W!x�7]��iA�?��2�lg��)�j��&�}���6�v�(�'���@�b��<�R�w���������2s	����%�	��������Xq(E���B�Gl>WW��4?a�I�ڬ�A͂o,�1�ک�PkZť��`���/�ǼBdg-�"[p:�8}�5��f�|{�â��}��}S���=��DS4<-�j2����͛��}��rR�`��H���d�[:�${Տ"�"�g|B�m}B����YY� t�~?\V�X�$k���ϥ!�$��}���iK|T�j̑�,1	�h���~zo��i����#i�]>1�7��U���"��fWŽZ0��>�Ѥ�N���9E��&��X�8���{R<#�����׍�_��9��t�R�2�A}����lK�1�����*\�
��<4.��8���T .�������ya3/O�[�eY�ve����l���M��E�뱮���k�͓��ӯ%��1��yԵ�Thc��QIʍ���S�^���8�e�J�c�L��K,i�[m��Php��@�2!�9�P��S�PC�q$����n��-HO'*W[�lY�~"�`"�*l���<�@AغN��BIⵂ�x�Q���unu}�I��R����ߊ����hw�F�4�^�p{w����N��y������VS���B���+�E���V����{����n4|i]�v�����qJ*���
W�E�t�f������b?L"��f���W�ɘ��k�+�#�|:U3�Ҥ���g���z(��� {:ƔʗK���>�^\�&X#��o8����O��n��^�&�uk������;��C���]����L<�O�2f��" �6}�R�b�'��}���M���ה��ɣ���2��4�#Jz�l8�C���N�o���oa�jO��[LW��'O9n§�fjeބp��vJ�t5�3���mrQ"}�>iw���/��\x~���@��[�1�m]j3Vw�59#ف~U����h���o2�C�|S����f����'[R�d�����I��-?��������[P�T=��i���rK��f�'��l|-lNwl=��bE�8
"_��Ł}������0,�p�$��ͤ�;w�x[B��6�*��/s��{%�����Y�-��;��2���;'�qF7��w2�^z�
fP3�3�{Az�����:|S�l�ũ���1.��ِ�ͬf��wZr0�M��Lk0[���<�(�6�������-ڏ(z�t����l����"��]�y����	�E>��\�"���Z��	���6Wb -����
檈L��Ӗ#����O%#��X��m��4T�W�y�k�%�?~>Zd��1a�:��wY�g�\�I��ӾF:�� �!�)�{}��+�a�[-�|�v.m���NB��D���7��M|5J�D5�|��Ϭ�R�I�����Rn�^&{�\����941�@~�<�LO(K%��,	;���q#��U�	�ڼ{&���o`����z9���2��'���'��?�:�R!�8�?��fkw�S���|��+宽��D��0d���IP����v�=)��!�`�J�O�p{��.n]�>#��7M��Z��"��T<�I����8�u(b�f�)�g�W������43uyjN��:��!,�?p��_���AN��(�%Nhk���䌿�şS�x:�"64lvg�I�����P��-��<��9�<
����o�v�~���.K�����:���5jaYC�m�E7i�0C�a���X������s��F�=F�/�0b2�qd^ ~r�\�/ֻԬ1)*��J���c��T��"0��Q6��om��V�\K�<o?�
yp�Fc��(�ON](;_�M��G�����\sd���}a���ör�7`����3�E2W�������;�(����I�?ak�YL��t����E���8L�5K�Yq�g�,n{Y���9��3��
dP���z���;i5&�?�R�|j4�e��9�U�67�½�vL���b��#ܓ���k x���U�/�3�v�=u�Tu?ǖ�!J��D��Ԅ�� �z�������lx|����
NI�b�L������hBc�W*���g�����r��h_R�mL����{  ~�ع�e���� `��Ym����5`��J��v0s�1�E�ZQ����w
��p+$R�g�2�v˟��I~�;��ѹ�����jWm����j@De%b���у^�Z:�s�R"�3���*q�e���T!CQ���c����{�+D�8b�������~@�;��8�]�ۀT�.j�;o��1���ɂyVi�a��DC�B�r&fO���4"����eOa͆���ɮ�bi۠f,*�9f�dV��ˍn���p+����s&�ǵD|��`�.��v|�+���)0����̢teL������e��S��<�S�Y�o�XsF٢mǡ��%C�=�а5\�f��#xD?����8ɍ��J�",
/hǦ������>λ��E�Lƞ�jA`LĴ��r��>BLj�:-�)���2ZO���WO0���D��t���&��E�\��Z���]��wB���p�(�JH��smNހ��z�=��
�lQ���`�Fy�x;Q5�z���J9Q��J.1��仓��]�;�B�:�t���.bY�/�S�wr�k��-BE�f̢>�t����%QB�L��;@	 ��nqi(g����$%چ8#Ǎ$U�lcx�pשh|��x��#�uN�2�!�)m�M�3��PHD੣��ř�W��W?�&vǏ��A�Q���`w����IK���C��L�MR�{��&Ŭ���7 "�FSK�#�h����1�����<>��N�}��4{F�B��s�y��lR~��gF�ٖ�3�ܞ�W�Blv읓6�b���I5I�A�<�ϟ��!>���3�X��=	�y0M	��pM!LAf^����������sB�(A���/0��<❰69V�}ĸ
M��[��ŷ^ʒ���IDRmV4���=��`��:� �l� 	y���RPA�#��U����~c�r�ٺR�c<�ſ��96hW���T��l����U�H=�ݘ�'٢��%�(^K�V+�KOC�t7`'�@�-=�����3��;����,c5 ��䝗q!t�)wԌ�����kV���zU������L�͈�	�KN�Q��f�5tl4�����A�-�����j-��R9�t�е�*�j�`2E��������������nI�h���3悈 Ӻ�2��u�兡��W��	�$X1UA(����P� �ps3�`�61��-�Y���aͲ���Nۇ��DH�wF�)��l����J��QG����M��H$�"��eɸ�羏��|�U>&|g�:KP���Vj�ޞu�z96��$��fB,�Q.4=����`C:9�x�P# ������Mi�V��Gp"�v{"$@~����
ң�Ej�f6�����jC0����3-�QXdꤒ��o�J�tbǆ�G��#,��T�F��g*�@A����?L�s�z��Ǆ���P֢���x\�unǝ�'��W�v�o/U�	��{�*f�����`�^a�#,l�lOh
4�a��̒ː���V�5�t�JǕ��N�2����q�O�&7JEf��N�d�d2�YC��?)q��˔7	��������I7�Ia�>���0��Nuo���a'Zz���i��*bq=X���0�	E��t`ҲK��`I��(��;+�*LR�Zv9�	�<���'�Fce�J�����/�	W6DH�밐�ف+�e�P�]�K`�C��\V���smi]+��0t	+*q�R6�Fi2���L��k�֠~>a�1x�|���ϹX���Ȍ��셁0)j`&�� Lt��a��_ d��Y�G�,?0������t��e�PY����ݬ	-ͤ�o�c���*����l�YN�<���;�CAVxk��$U#rZw�ߛE>����w]@b~Ġ��CO�*��\���Bwq>x>=����V��l�s���E�������ݒ�L�;(���P�c��,]�K��>l",�t�!�� Ω������:=�Y��Z>[W��dt�����'B�1��!��~���`�E�ShT�A�u��>�&3H��&c�K���P�7��ҀS���Ź%%�
@2`<�د���ʀ	��:�A�j�e��C�R�)1���t֝A�x�>�kC�[���o[��9k�`V�F�-"Y�肷�6���)�Y��i�[��ӓQ��G�6�l$ ���	����.�oe����+�ѧ����1��ʽ@uMI�_¨RB3�� 8�(rv9�8� n�s���TK�_`AƮEvWM�Ӻ���~	&�g�C��P׉�-���Zb)��5�.�u88w���?&���~��)θ'9CD��w�-�ɶ��t�Mc�s� �-�j4����":�,���c��F�g;��!�[{f[�b'}�*Ur$�-;�1����ྚ/;Fl[�z�1���q����X�K(�-i4Ϧ��X�x��uU���X��>�ϛ�]������ū͵�'L��)17_�."L�8�0��˖��&�*s��x����Wۍ<���8Ȉ���������Zq���a�ţ���cLr۴������W���HCJ��z�d���ȼ�a(ʰ��,��������[F`�I�f��U� ���t=H�{���5��\K+��~Μt5ɛ���"�hī�iM�
=����p^h,��F�V�m���N2J&䧶��tb��"�C�r>搄p�g��65��ˋ%��ZD&$ROe�y�Q��r"�� �S�'���>�;E��_O�@��{=ŀ}�A6r_���>�M��Bx쇋0*���j������]/H��<BƓ�<��{�=�kk�e��c�s�x	l�$����oۿ&o.L������?����;Aj����vB"��z!1�ӂ�
.��~�{��l���a0|ő"HĠ���ro�lWKWHF�j��"��{l����|�k^��J����Ad����ڇ�j��B�+�;p0c�xnnyϓXx���ҋJ�E}<k>d)���;T`��)/:�Kr�j��O�6��[�$�4���~��_�����.a��|��,5"r&��l	qi�S��Ͻ7����Ō���/��_u⬼�o��]���}�5�'�VtسJ_��E�N����lK�7���V��]:�>m:Ms]ut�>��Lo�~YhZ0�4m�حD�(�+�F�!��4��~�1��-�!���������|�;��Z�j���Wޢ兡�H�әk��"��ղv��������  � ����1�#�iþ=��IMKSx�n'�Q�L��[��1�>���p�����zϭ�}Q$aI̽�F����1�˃�ȧ��X��lѺ��
��E~���8]��Uf<2C/�}��$6��Q�Ӛ��UA��:��������:0勳��r1D�pD���s_�It��yg�s+�T�|�-�3��Ӗ�[�1f_ǀ�� C��6�;���lwJ�\U����������8S�M����u
������'/�D7j��"��;��ic����aK�a��|U����v���iIx��;C`�Rޙ7��~��C�1��N8T��I/��O��nUSp�٥1B�ی�6��uq�)8�w�Q����*ʟ'��(Q�j���<;ǭ�m6��`@LO��NW'��~�)J~�6|y9��=O�����JСF�;{J�n�Jf���PB6�	�t���=P��Sb��}���I�a/�L�6�崈KUǦ)�7�����Ზ�L�9ܾ�QrY��Ѕr�`�i�?�	K~/�5M3���5�����H=���L��E:�8ƅ~PҢ��I���SF�}��Fym�7�P^���!���ڍ��]�D�����5C�tE/����`%�\��
��N�a>��c��Y���j�V��L����~��X���7Lr1C��Y�M�l�f�O]H�ڂ���;�
I7Fr��(�W��W?������̮�f�c|�J�}k�λQ�
9P{�ʪ�V������ߘjho��%����lBs��D}?p�M6���%`~f[�_t-��K���(�H��|gۣx,w�q�CÖ����V� 'n�\xx�{�� ����Y�Y[W������'��'dO�Dcj,J%m!;��K���'=ǡg�Y��`���#��c~N�76CEN_!�e���nʥS��~�a%�)K�
J�&�^�����F����1���$�w���(ǜr�$�r	����sJzp�cJ�(B沭|��!��Y�<�z��=KU�A����Uβ3�Z7�n��H4�3��v����7l�q�>�	T1ة�^8[�V90�HM����v���`Q����8��	�/���^MԢϲV!kMA��C(�Q�����?��6�.焭K[e�+��n�WHJaMSP��R�|�D����p$E�u0@/6��z��|�n9,s�Uf/Υ���_Kz��Kvʅ�O8m��v
�8���'k��y�)D1�ryW:�=�j���{+7Pa���(�i�$�M��V\��� /�Պq�A�)08�(TtBqY��'��376���?�SU��:�^��==Me�z���~��l��'���'�������ap �rU��ú+�^~���^-��E�%ų�� +zR0�n�dE*���52���)�!m>n��!��7X���ҡ��n���Ra�����T���;�2�p�	����-/4=����0BL� �FEO�N�q������e���kl�.~�(�`)8/} $����F�ɤw��Q���w ^��|�{7��{�.~�$��P-52(_Z�6�&�L\Ce㐺7�E����H�=~:�(Q����,�]:� ����`2����Dc��`��O�*?H����"Z��zˁw`��_��� ^�>�    ��������y�    L�5(�ת_V�3�+8���-���ߘ���<�3�ˡ����>�I���/��Ei�Z�x$��W4;X;/�;*�3�hm3a�^DB�R*@K o.��w��؄��Z���y�	eI�鮺 Yn�D�Z8�c�a���^Pu^�U��    �W��3� �Q+_�|D�0���/�����M���鈮�l��8��w~�<s���\��%a������VJ�����:�F8`�[k�����X^�U��[��7��(�<�^	e�;���񁔝\����k���V��G�{�9�h�y��,I�o�J㏿����|{���[L��z���P�L�"�q�"��Ga�"���ԝZ��NY=�l�:$��	 �j?9h���[E���b+#&;f�[��C�]"ȯ�����_�    �̭��2����^EnY �I���\ �$<a��j0�jU��F����c[@            W�ᯂ���`I�k�*g��6    ƫ���Q�C�����S��;R���BP`�e���t�-�
���l�Y,kL�.Y����~�i�        �#Ԇ�NCJ)1�p�%!n:Y    JBV��&��i���l �D�WE	�h*dD�^���e(S�lߜ�:,p�9�<�����sb��I܏�Ύ� l�F��E�����m$u��d(6�ƛ����}��Ul�Ƅ�V\4�%{�0w����VCH�S�����\k��pa�+�-!���)���`�SԤa��ia�z��MJ*���>��<;6���p���fe���c�p�^�D�ߠ5^y�	�d�*q���.?���������Va���c�\�g��XLw�nD���i(n_��@Zؼ�B�w�7R��c�m>���Ѧ����Y�!���}|��K�Wl\��zE̬y�%�w"�f͚#�>�U�<a�b>h��j��{�#3~��dm�˥����D���s�gyG���T��9�N��7�� �̜�mR���2x�J�����(q��Ӥi��v�2��5&��w�0u�X��*:����T�����:#|�tV9�=$3�Ј]��W?���J-WE4��7�ܣ��K�#��B�A8�S�֩{`�76����8۟Ƴ�F�Y>=�8�U5���<��n�)m��g뜸�T�
�4g�]X'f.{#��(�N����҆��6d~�	p�o��u�f��X����\[�,���7�-�p+���T�)i>�����NEs�ڣ�߇�K��_�m�b�I<K�|h���-$��_����\�_��G�G��.�M)��k�ޝ��H���n5���X�4�
��ю�6��Bp�����l�gyr`��8.��5�S���0P:��.?�t�S*�{Bbˤ�~�坭s���ڃ���V�N� �Y�6.�<��Y��I�v�n�� ��sR!��!��X�2��0-��1ʖL�q"���s�}��o�Ԑw\e���Y�*^h)e��b�<��.E���5�4�̏y~F�Z�^�5S�����񱌓������[Ѯ'��٧�� �o)�����v�Lb��֦�̃[l�&���"��g%=�?�u!F s��Sf�	h�?s5f\���s�n�pD���>��#����*}����ڀ���ˮ�ք^>ŌLwJ���������[1�Y>U$3��@�y����5����*d�B����FO8m��3��A
~��Mr����.!-fȧ]n�|ؼO��u��x��FeE���-ꕆX����m�Hl��>o���	���� ֆ+��
���n:d-�b$�'�s�T�����}(S:����}�%9A��p؆ �GX�C��J*���M�`DTA�.S3�8��3`ͥJ���N>Im�F����:
?Ǖ֪����Mh�e���r3 �~EzY��~'�XCQ0��QE�8|�w�1��#=�Vwy�Z�U?�w���n�a���o� 10��	�0����{/����EĊ�P~W�	�SknpV�&.@ƙ�� �!��7YV�X�;��oL?����2?    +���D�r��g���֫���9�@�36�� ���m�+
�ͳ�Jjޜ��^t�5�i����2͙yD�R��w�p0u��)+:��XpT�O?Ol�:#��rV9��B-3�Q/�[�:�>��6�VE4&5g1��g���>��B�M�9�SqD�{` 5��P,ӟ�L�G�Y���8HE5a�<�L���)m�a�G��� 6g��U/f.m)3�(������=-^��6�k�	pE	����e�ƇK*�����,��Ѭ7���.�p�➩Tb�m>����NGs�`[ۣ� ��K67�m�%� �I���|h���) ��[Q����mև�G<���.�״�k9��̷9��n�����Y}i�4���
���w�{Jq��H@�l��� r`K&9.�1����0[�xR��O��u�{B�jͤ��Z�k�Lgr8�ڃ�����!%�Y_��<�s�I����w�n�aX$� ��P!��m ����7����w�	1�i`�q"��}�␛Րw����,^h�e�^ �<��x�+�ʇ6�3}~F��^��`���+𱌧���E�Qb������o�An��v��NbЀ)ۄ̃���&M&�"��l%=5�iՁ��Qw��&�	he>>s5��^��"��n�rDAI��>mP��~��4m�����ڀu��ˮ�҄^�?�Lw�����"����0�Y�I&3��������o1�,���<�`�B�����y�i��>�Y�������l�.!�^٧]j�xܸK��q��|��BaA���)\���z��Hl��>oS�	�\�� )�#�����a0n��b� �s�S����/§z,W>��Ƴy�!_J��u܂!�u	\�G��N`�����gLPh�0T7�<��7d��N���E%Nh�B����>;ÑҮR�������e�C)a3 ���`X�T�$�X�(=��׺�<|��s6��'9�R�R�Z����wS5�n۞��I.� 1�E�	�4��������gDĊeW��FSkjtR�"*D9����U�!�#�QV��:��H
p)����3�u#�.���<)vazuu���e&��VR�J�DESX�k��uj��A�yd	=�%�y�R�Z$~)	>�٦���$Z�m����N�	' fnhr"��Mɯ�T|���1�V�sX���3*��0H����c    �ٽ������c���y����5�=J�cn'��n[e�+oCg-JA���+�����2�d	�X�{q�}Ró푥��@     fQLA��!�KS    �e@A�l1�+�Q���g��d	�\�u�yV<�	�ގ����K˚�3"����[�:�(�B��r�d�m�1��Ʌ滜.��%�[5؈pC �nW}O%T:�3�pd@��BV�1��h"���jzx�ɟ����b�MD�~1?��T�6O�)�=����%G�H�!�!�Ə�L#{0Si�.xLm�aIMY:�L�,���Y��j�э*	W%`ؤ)�3H�3PFf��(L��V���#�ǳ �(�}�\xfu��G��¬�B�J@\�;�^���p�G��	���9D��Ez���&p��c��u1���;�Rh���<G��5�������P� ���q�{<p`a����Sm��I�&f^(�V���!�~p�A4�d��ֶ/ �[�'5�N�m<�1:*΂w~��]5��㸥�)a���4�����ݎPO�W�:��H!F\7��+�Q�m�S���P (��>�R.-�f4մ�Ђm��C�>F�4�]|��s��I�x�5�2��t��}�u� %\�S�k��rTl~�Td%:�%�yOqS`6��n��`��[��4n��R���%L�5�$y�$�ts�ʇΘnQ\:s+�\狙]I�iMʫLz�i�|��?���3kUc��d\$�9wA�ьg��A�ơV���@��Q���@�p>��>q\���[tκ2D���HVڊ3}�\��?_SN	j��~>[�Jr�%�xպy(�]�����`�p۶��g�NG<�{�+]r�E�^�*����5��hB��u�N9�_�O2e*(��R3.��L��0TE��������'��2���8:#0.��u��b����)Lr%�W���q�a��/�o�x��1��{y��Z�2B�dZ����O�ERbs|o�!��/k���@��Z����I,<X6�̯]�i1�K_�8���j�bm���.sŎ�(��_��wF���(��m��g�EXQml#�p�yʁ�6cC!�)����~q~sW��6z�m u�+��yQ��=�ɆL���G����Θ>A�]/*9��L�-�Dt'L���658
n*s]�= �L��ޙ>Y�;��zϝ^w�Q��v����(O*[o�ſ)�Ck�R�nƟ�&�1��T/f�z�Fބ��"P(,6I($	&*�I��a�ʩ�엸����Đ�ۏ�o���Y�.���ʎ@��S�����cn�$N�C=(~G%ax2��
}��[����Ĩ�	�q�9ƈok
ц{���CŖ��R� )�c�
�~����u7d>,�.�.^|�5�j�e9QH���M��=r6U�" �������S���|���d� @��2#K	!j�u��̃�f�	�H%�?�X�$�	���H��#M�NП�M���-�H�'N��o�+�3W��t��)i��b�Er���mz|��!�mn=A/1ݮ�.�R
Q6TN�2:�4�h%N�F�SQ~ig��C�P�Qd�k8�Y��b�L���Ԣ��l�U�^�?�d��*��]].ᰈM6a�(�/�?��@�- eѠ_�ކ��#����ә��H�趚R[)�]��~~��SQ�8��v�m�u\�ش��ۇW���<K\�zJxkb�������h�I�����a�Pܾ!����:���`�w�;���B�KM ҵ-p��ۼ}¬ܞ�MJڐ�=��u�s�q�5�B�|F�``�bdܣ�s�����c�ݡ���K�w���'��&]��x�E(�{"6C�C��zH�ay\ �*ЦA,'�yB}��
�H+ #��7 K�'���-��/�u���7�W!����@��j�1'��:�&柦�x/���P���&n�{1��GE�dx7Oq����%�@K���T_ˢ5W��1�D�"P��cp.�N�mW�eP��q�o|�&0=��Q	�h������}5�G��$�W23��L�	u���Q�ז���>�(�I'��l�v?eز]E�l4��>=Q��S�ƣB���lx�ﮮ����.Z���Y�h��Q{>�x^v�5v[I�ѓ����J�����ލ�x⏨o=>�z�����~��8r:(��^��lG�:���x��Ξ;�'���@[FLf�6���Z���rQAY����\៫<�\D3`�g���uA��#!��ݢ��R�� s/0�4�"���Fc���-��+5\���PV`'+c���U�i�ӵ�e̕BWY�N�7�|��p���{RֲQn)��h4a�������+�R▭b��0����ӏ�@�3�=��!��2�
t3‘�gڧtx�]ά�r���ia!�O�ZdZ�G^*ӎ@�Ua�Y����0��Ƹ�� �K��%���2Dp���%7��#�"pӢ֝,a��2Tt�➧��^�M�Tw�D+����xb��,{�K�k�]�Jvl�X��ݛ�ƴ��m��N~���\v���d���[t�5|�����Rh[��dk)>ߐ� V��랅����F�n�H$���	���y#D&?��pm}���e��B-A���n~�vK��3��#�*Vi�[��7�#g��zX�����ug-����'l�wq�3�:���d~o�	��Y����IE��
uI��gYj���˻D���UM���5������+Z��Ì#m��L��$�H���4h����z���+�ޫ������'Vi�DW�ֲS�2L�Vyv 9Ȓ���[��ʅ���g�hoGjH�Q�#iH�}�����3��El~��"1��Fn�)_� e�K�XAר/#Т�=����)���gM�,���Ì�H�_�8�Q�sݛiC�������)#��މ+}���A��\N�SlCm�(���+_��q|7����q���}��e�76V��YLc&A���M�g3);��Y�>O��}���S����F:�.�s�%U��	�Ĵ��k�h$=&�'9:�f
5�y�J;PmD����1�<ͭ�1f���h�I� �0��uY>�xQ�Ω���� ���B��GX�9e����iZp�>G��q8�R�3ݧ��c�V��eo��P�T�c9�K�SnƜ�sRv�?�+�8/p���M'BE�C��u�&we��=��4�� B�d��K�Q��9t=� H�!>2�6		W�EY4������!N� ��m(�Tދ����w��E�2�Q
�赒���@��@Q�Y���浀������Ek����ؾ�U`��E[�����}aW�:
�Xº��i�۟�>��c���E�VG�6���;�o�9ɩ��;�W��ڽ?K=��)�<T�)�y����ѭ���'\r0ބ����`t"dԈR8�)�FJC��C?ǖ�?i�c���j{�p�^�(O��U.f����9~��[��D�l��&%Y���d�RQ �/��g))Ŏ��Ā)�V�<�wa/�	��}�r��Y0�ԌYL}�JP�+��~�j����V׵��Ư����@���0��R�{ML��}S뮷L�щGw�>So+�.|}�[��
R���bU�mp�e>	�` �ǜ�)a��|��G�8ɓ�w&G�����4�ހY��$�ڝ��ȷ��d�k�0oA���~
+#�K�\)�F�'�"�:��\)�m�f���&�ý��n~��QT�u>�e���݅I������k����H�rM6�i��ƃ��hr��z_�@N�~�@��BA��\�'��裑��G��lX|.~�A^�i�a��7�2)�|�	l����	b�?0·񕛆��0|h�WU���S�:�J��8{�˯���B�j�ܒ,`��0M�����Nî':MX���렀��`#ye����I��ڤ8��/+����M&�j��q�R/Í����<�+2<�t����E�\}�]�"ν(�V5��5ʢ*�do�����R�PZ\h�{�9�{�Y�V���hWbZ�}	w�y����|�S�Dܔ�(S��>&ߟU��l��A"�dź>`:��i��.��'�aRm��O#�m�8��alO�8�&�L�PJƤ�Q���۱=8u2{� ��ǁU��A���m,��i�c�#=~hj
3p'%����z��T��������	l�/%X(�qg(au/
�VW��q����ȵ�g�Ro�ڴ����-��)c�A�B�;Z�Q���G֤��gK0n$����ݚ;��We�5��n�y���ӧQ[̏-���Ƒ�����^V�Hϑ�v��q�h-A����z�Qq�����#&�<aq9��:x��͑�e��E�Rs��B��=�˲�C�`�jg�	�*���/�'E�����$ 95}�3��eC"��A
���fYeD�D��m��3�1l��������MM�����*|��M
�h�־�.V� ]��:j������h�a����׈a�D�:дh�����(�4ea��܍9�Gu�$�Ѫ���4h�a42��>ޏ麻�b�� ���I&A��s
�Z�;b����̌��W�'}&��/TU,u�'�4~t:�p(OLf��fAny>����	�UMI����[�����2�S�ip�?ܓ2��U7ߕ0�MO�a�����R�f��|Nt]�7A�8^�Y`x6���ˮHo0���j=��
�]\����]��@m{���l�w�nZd?�6�z�/�%I?[��ⶼ"W��6�Q=��~����@�؜ޗh"�@�;X���Eedcl���'������n�돻�긹1�>��X�4�E�_�%ya��FA`��&��R˭n!�|���x/7Ѭ���\����M���ω�}��mf������ׁ|������'z����&���M�q����]Ķ>�ay���f%�Hߖ�G,>��ڼ�B�N^�F!f��sg������-���M�~�."Zp�b�ǥ�������0Zy�=i=�Th�'^������C�������ō����ε=m�dap�'��n����Mʮm����$�l�=3d����_ �Y%A������m(��[����!u���(,-1EM)p�#���8�a]��6/D*«�q��r�.n���w�e&Eb��$AHaV߾��ϼ�g�'6��O�_O.�1v�Q7��ꦠΊ��ဟ��&H�`����V����?�b��iRO����ٴ�?9��£�0ďU��c�D��zp9�6�j��z���Сd>'�߅�M�%�}�f�ƞ0T-���>��d�?V�f��$icTɩ<3����$�bz
�h��Sh�j�*2�| -�E���^�
�)�@�D}�u��.�j�?��9W��V�^_�O!AR4�:R� ͂x�z�������S,;���x�
S���@fQV�.��:~���2�ޕ��f����cR��~,��L��NnΟF�5���ς��]�8��2�����D��--F��֫s{�o|��^�	����o[��`�9A8�
��5^��^��G���p\�=�P���3�?C��T7ځ3�;���},>q���(���TyÖ{�v��[6v��1�U���0���Q��֎�b+�6�ѽcx?P���.?b�w�_ A�@��^$���v��a�����7H.zb���h4�/>���CK �W�`��!	�#M�-o�g��K�����߲q��X�}���-�� ��h�>�b���`�]n���͹S�ϫ�3�H��p�Nkf+5�D�g-�J^f�,�8��9�qڹ8~�	���x����*\B�<�X�Z���q�y߈�����*�6�e��<�W��!�2f�=�����c`vPs�iF���%�t�7��"�cv�Xd��l�R2>�
O;��z��y�*��� ���5�M5�v�]7̦�|��H@�6�S?@��`L�ː���5�U5�֜�g��n�S�i*�Ǿ�^�coG��\9���0�,;����:	-sKa��d�����y�}�zc��p%�	���P�����Q���D(���:v �T;T��ߞ�I��%Xj:�^�=�6����/��d�/3���#���3�Jz7��5*�.��l�_S.��z�ޜi}�x8:0����$�Sk/���VX;\+#�����a�{� :yF~�M��փ�n�͝���p��F�0!Fל��HD������A����s8���a;򀅑ZQz�Rb~���Me����ߖ5�J'$�#�/!�݆22��x���+D�v
6Q�|!.�T�����e�Į��#�����BjL���0�̰{ fD̯����M\��k�%V�]~�꩘��V�?��R���LC6)��x�$�Yd|�,sЉc2m��2��AX��\�	�	/p��`�:�Y���} �C��@mSs/RpCh|Z�G� ��� ��i�_�X��X��S�ql�h!uC5�kk.��	���5��� ��ۉE�,)����,���
��^;�JI �T���[K{��vMu��5&5"�y�h�4����Rg��Hh ب,��Og���g���=��[[�h�war+�!���bPcv?�f��ŗ��)��L���8�TR�,���^0�d��S*�mZFw�䫶�J��%�s4��;���A��w��)*uѐ�Ε��:ݍoA����C����O�V(Y����}�����×��%LhK����jT������+;�G��C�L5W&l�+��h^D����>���Dp�@J0��ǆ���ۡ�܆3(�) ������>���G�&�&}#�v;5�|E�f�#���Re�:���Z�bd\��E� T�%�s{o�_�̚�ѹ���uT+��aJ2�(���_��ex�nM$�O�É��\t^/�?�wі긟��+��Piø �=�^".`��] �f#�Ԇ�1��JN��"]^x{�~
��ms�����N1q�y�������+�k��L�'�"����R9$���Sc=���1����V,�����6�a����<A���֌��#�d�a����>94�/�=+�4ZU�?����0!d�Ŀ��Hi���n�G29Ͽ�+���jd���z��:v�Q>��$�6|�ƾ�^��f����ǋj��ȟ��%�� �E�+?�.ym@����0:!��҉�-����L���w����o�4dח"��:����)�>_a��Ƈ�k�ɲ�p��̙�xǟ!JW��1��۹[I*k,�1&�e9RE/��ou�5լ��5bzv��Ҹ���Z�O��OL��ڣ����3���&�Z�����y� 찬~��w#*����H0��:ށ�~��߮RP�=���h��ّ+>T���Ș��=H�B?DSs��~����o�2��'�}Qu�$�@N�N��)�e�W,B?���s�9GG5g>
u�q�f��S~Ψ)�m�,��� x~�&��p ^�B�Ee�u<��6=�H��5O��9�G���"�ާ���"��J�N��|�a��ʫl��b[���15��`��*�3MK9S)ۊ��W����Y�qlF�L�鷹4ǿ�N�qu?(�����<ۢ�zS޹�κ��*���a��\Qv��j���� ��%�|�ۆ6�
!�k�1Z5;a�p�D�o�֮$p�ߋ�Lf��!��0ǂ�|f8A�N�Z�&�*���"o"@��
�g+�>�]��Pǵ�J���r��EL.^la»����	��^�����7Ћ�)dM��ڿ#;�XؔB�g�&��$�j�9o��do��ˤ�qA|{W��r���z��� �B�r�����Y�G��(-�p=�W2lv�,�D��h�d�y�w�䦼[Y��ޠR��q���@�7�z��.�!�n9n�T"�#L2�H_�i<A��>O"Ǔ���H"R��>��c��P�1
��2�z����M�CRےD��;��IE"��nJ�"�?�r*İ��H����� 0�+J{����ߎ쳎 �M��V��ϗNz�8�(jM	/C$3Lr����[T&:B�-=�.2*Kn�������H'�}a�p!�'�[g���{�,�N��2*^��<c�9{�2r�����g�lr���ڶ-������}�(�
��c�sCÏ��fNS�����iq�Nu��Z�d�&�ӋC���"�z�I�qa�o�?I2����,a��/Fd-x5ϒHļvb(44$1����#6 �y�~�<��<+N��{-<+3�1��Kt�qZ�{ؖh]Q�x�-r8бT��
�s���[�E�iT��+|8�p-0kN}R�fKj<{'��g�4� \RT���jE�����+4b�����m�R���/Z4��=Ef�x9vs.�入�0�d����h7�Q�'<���5�]��冥��\�,g@���(<�B�wgoO�J�'���^��-K!��2�Ƌ@h�W�d͛Z��q�XM����B��+��C�IN���-{w��9�a�:�Dk�������=�JK\�Z�g��4��	�,�6ek_a�O�k�6&8�GB�:^�l�f�g�~x>����["M^��I&j�&�%�WŉId��K���A���9���������9�rdI^V
��<���������,c$_Tf�-%��n�]T�^�RN�������X�{�z��
U��D�Gc��#q��V�v�W6�5pT۶:`8���T�,V�)o<�Ϧ.�6�~0��8�G��pdx�~8�ߡwr��\��1����H�l��n˦�h���1�%���P_�-�:�Gh�R���Qqf(
�J����C��Wb)A��"v>�D�|&��^O���=�A:��~���.�����h�)��7��o:QX��!��ǭj��-[ ��9u��;`5a?ڙ4�L;�=��{o��}LL�T�K�xX1��?�4�,6t�>��Q��!��!� 	�Ny:�2?�iA�_���эqi+�����5��1C�,�q׶]]�p������f�=�&߃പc l� �9?�ޛ����r0�Ik!08�o��r�͆3��A���k�c~r0��=�]y��b�3#�E<�����������J�NnK����)�`�;�Oȉ���xs_g�t�[��N]��DU�V�������&F�:��w�]˼�0]"���$���zw,(�x��$ڽ~q�<���M˪81!�u�>D,�d�$y{o
�87������β	�����l7.Uub���L�}�\L��>6�����F�Pߴz�@�]d֣$?���@Fm��|�о?{�acow7e���=�)����*�����mF��y�4k;A.��!��4*k�;� kZ�߫sq�+�X`ԥ6_c�W~��,\R����sп�gd�b�/&�Bl����8NXp��.���ތ����Y��7��E͋���O!?�|���1s2<^S��ͻ���v��ZN n�޲C����k@�$���>9����8�{i1{0q���[)b0.�At� h���N�Kmz��`Lvz`^h�
��+�˜��U�B��N]���eJ��F�����!�A{�&�5}�>�~ٶ3[���$�ɽq*К	����Y���$oo�/Ȱ9��Eݲ��Y�O�`�Y�����837�[�[�>�W&���ޫ�k��͛�(ms�O�ف���"�Ȭ�8���C�P�VX���d� �Əqv(��"����.5���0��~jX]��,��ETM���@���<O�
]����"MM�{�Y�G�� �!�;�?D�t�,Ӂ�ϏUK��ڟߥ.,���h��n�-��y��H��e���;x��J.M��bb�Z\-nQlo5��k�>C�<?<g��w��J���Ԇ�`:�!]�����M�!�7/�
-z25P2�jaF��^��
_�!1�#!��?Et�,�
H���w�m�F������%_#Ǧ1V�h��Cy�]�5�dڮ`�w�i��t��o�ˑ��JG���`?,B�eTv8N�4o;ާ��C�rk�Ǧ91-6��Q�·Z�)ӷ�W�ή?/�ƺ�����=y�/=Ǜ�祄{%Z
f�[�����շ�3�/���4s��u��Y���R�4��ʸ��v9���?!��a�3C�Z������TV|8�r�s���/B6�V�����#�uClUF��%�ɿ�ڀ#�����	�d�4��F���߫OQp�u�k�
�H<:sMwg�4�G��Jء����D9(^���ϼe���"@��VXFZ�6��c�W��H*�"��x�0�'���ϥ n=�T��!��:�A��������4�:?�=�@��6���ϲi�lI��{�TG�a\�ۺ��+D+��*������
�6�W\"��p&`�rB���¾�I�qs�>�(rON� �����LʓM={��Ӹ2�P��ey�Z�Da$<f�N{�c}���f��,��6�,�x��؁b9o�/
1�]o6΀�,�8������W��5��l,9H-���@|B����x��  Jݦ�`D삛�ȁ�7\̯"hY�����m��,���� �G�����hL��r#ﻚ����c+�&���0/c_�}�~)��R����p�y%Կ�謪�!�APzr�Xj$Y�����	�'rb�@ᠩB��]*�LG�B�Ҙ�l�c�����5��e�~u�V���._4g6D��!�j�?T��*p܆Qh�3#�����A6i>� 8���+����.A�
 vG{����[���@ꭞ�x���jj��f\�S���#Ǚ�M�ޞ^8��ED���W�]M{�W����n�X��X,o���?P�P��ƾ�Ϗ5�z�+T@7W�y��c����=����ۍ%Y�Ջ�}���5|����!�Ћ�W���v:�X�
���?X>_�N�܍#�*�P�:( ��i [�U
6M�������u�>D����S���.�����K��J�}R6.�n�3z���W俺i�!�|����ԤvP�-����(x}��)Y��Ҧ�_Q`��aWQ�[� XsF��L�LX�,�-4����v��KrOL��-8Dz���@��}��f���o��)r��⏤Dg�:ӄ�v��	����Iѻ���W�\S�GO�{����S��{�~�pO"�T.備����i��(����5����rM!C�����Se�Ա8��0 ��Ge�7���3q�*Z��̢����1l>��nj�pԆ�K�@�h���h�^Ԛ%#.y�8t�!�:C�g><0}AN��������?E���b���T����ɞ���|�3*�Y�ꬺY_�B�B�6��V��@C^r��tC�	��#�0ax>2w
\H��ج	�Qy��_�q��I��\Ћ��[�;���N��l���cF��։���(R���^Z��;����c�ȿ,)�t��B��1hM�Ⱦ҆�Љ-�<�>�Mh��fg�y��CK���I-� Ii� `�JQN�khh/�ߛ�Ӌ?9 ���VH%/�4 ��1,��S�
L�%6:Ǣ�H�CX=q�Biw >*���tC�M��U�|�ȗ'�%�3��7���S���j�eŚ��RB[i���D5تe��q�f�@j��z ��A� �z�ԓE�{GkAv?���n�C�Hlѫ�"�?9	��k~)��<�j�^뎌y��������y��=G0�ҝءR�d8�}�7�'�&1�"��N�B%*�9���D�ޢ���D����ܝ���i�W�@%15�r�f�v4���U��X�0�ӖZ�aϹ C��U�ˀ�{x޿����_��E����.���?��:��{�^��&[�W5�q�_R���^�u�����>����М�Ĳ�tO���^%
���fY�<e��D���!��.4
� �d�4�m�^B�0Ml*�2%��y�?$k��q��Y����� �P��14�i(�����ҚW�>.F��4s�;ﴴ�K�}lg
k1p�lɖ�iZ��H�E��|L���#C�:ݑ���+��b�D$��,4�ݒ��%�[&��(Z�in�'� (7���Z�M��(Z6��@'�ѭ�Nd�mգቕ	�&a��P@��ⴭ$~��>��ZX�Y�ěnXt7R4�������b�x�HE�-~���d�k*���������*�����X��<=�%y}��pg���pb�>w���?p���9�l�\��qu�n�ub�n�R�/ں	�'�wz*N�jDoV���
��������R\�W�����I�O��au���E�9oEۙg�����q��GK�(Z�q��=�`����3�9��]��$��pLC���ZL���o�o���y�f����Z�m��������9������.n~QZ�Sp3�	����s��IӉ����K%CT�y�ɬ��j"��)?t�s�+��;����|�����m�!�.׺�jAm4e�����D���Éڡ��o���V�)��ES7�X:�-��}��ı���0�.��g���5�p�:�eB������狺La�)Ȉ]^��ހS�.������-�~Xo�5q�uN�Ю�K�	=K�������U𐥋����Ť`:�����ϙC�S�p�9/�V�ycmU�6�<]!Zɢ�g�:ɩ�]���<�)�nTf��	��.�њ���*�C		q}��(ly����wp�<L�D���e�QD'���/��#@C���^g4��tqؤ\���$�5�t����O��tP �JV�F���M�^�Nv����� ����-E0e��k��]�x��\6��G7!�F���w'pl��Gvo]?�<�\�Mz�ys��7���^.w����&�= G ���S&aLg��E�3y?�(��d���/���C��um��0��Q����)oU����W��m�g2-������oN�6�V���l������MX���������/�
8��q�p�PC@�7�ՆX��i�5�NǸG����}���; x�d��n����8���S<'�������=ZW<@��g{��~��h�PJ�=>���J�+�#���Z��[��RP�� e�>�a�':�z��$�Ē�i?��*2Pf���-{�R �,�^Jv�������j^w+�9���K�j�B���L�G�`5��ţ1b]�Tq�>�a�`}j5�|���} ��
�]���"����<`$�� ���9(~��/���ξ �}˛ƔMi�h�0	�:Q3@�>��P��9�b��`�@�'6�1�ؼ>b��ؕ��c�<|��6��M>�+��̼PĠ�$m䣚����Iɷ56>S4N�Vmm�[�rp�6��C�_R��@��V�?69GR�u�-�\՘���,-�_�S%*`�9�ô���
W����lD;D 
o<Y�'Xr��"���L�UF�ɔ�}0I3+�݊&�֙E��N���w�IEQ���WBh��M��X���0!�&6�%�=	,c{�4u7����cu���x3��j��d:�D;�����Y�Od� ,Y�6�Q��a�R�ś���jxE���v����>A�����zv̑o˓	!�Y�2���eڦ�L~T�D��aΛz��.)Lyȝ�5~$	�S��O�RèG��i��P�2I���Ui��ǭZ�Z�G�T*�To��7&����2	G�O��m�93��8\�3WNw\w0W�I�~ET��;5,�S �}���Ks���4Q)�����;pȻ�B޶%��}�7Fhd$�r��@��dJ����%}�Sp���:�63ۼ���':��vRQ��l�,�?�����d��56� h�������B+� ��ڿ;�K��\�q�~����`�.�9y�>`��C�$������_ᐛT�yqlDC]�S��-���2H0�ROR	�����޷/��Y�I�W�t���RDph�?�o�@�f���;�\���{*d����!���VXb�d �c#��s�v=)���R0׮f�xf�ڠ��6�e}��KO����57QR��r�vk�o��1O�5�}��<(+ϐ���o��ww�������R���I�:Xw�o�ݪ2?((O
��[�C��1�W���ȣֻ�S��28ۆ$���m�斂��o��*�>����A��8��*t�^ǻtR�D�	�,\��-ZRq0��L3i�?�����ejsq@��/eoR����q��͑��?(G�5ݒ�e����H�Cs2�`��7@��Q�ȍ�)�P��a�W�g���jl�����*�=(`cF���+`�/�̴e�a�OO�������2ȉ��?>N�L���)��'יN� m�&������>z�r�a`<E�2?;�J����jG��<�r.�JNٵa�E�O 8�o����D2}-����y�"E�Ak�=��ӝ��#��ϭ���l�|�p�s��U_#8���z�Ӷ��@�I)O���4�K���Q�
�
�����o�U"t�tb�+���g�����ul���R���`�azV���R.�H<�Bw����~.ĤEN9|��r��䮬�de�e<�� ��2�:=���HH���t�V�WɋQ�[M�E6�x�=W
�r�	X4o��LEBvH��[��~q��:����iƑ �	u3L��p���c�9�x�i�̛z�����f�Y��/��n�7�`�:K��[.�T0��<�U�4�eI�����°��R�Kp��|��St٣��Pl��)��_.�(����c�|���0�i� �H]��� �2�:�֯�%�6��xA#aC��3�zuﲡ�pw�Ȃ��V9P�.�O�vE�kHf����s���X6"g����LPwBKEb룯v:�S/F�Ie����#��=?`m�y�Ta��ɽ��t�b#9whR0e���9����!q�2�Q�{ײ'�<yT�l�w���'����1�T��ڌ�.�P(4]�cKl����5��'�9�-m�:����Jʎ���o�(��0:�{���oα٠���
��2U����rڴȿb����L�X��شz'餖�O
��KS�e{cr�f��f94%?B����t�6� ��z�1��z�J�%��^�����B�;[D�[SzMcq�5����a8KJ�C�G���K�uY=��3���:����vauR����Ac�v����/�;��Q������U;����ƭm��-���(���".*�<�������=uy�j���Q�Ⲁ�i �B��ӈZ8J]IC�V�\cC��M΍Q�-I��ڧ�ʪ�K�bhG�F�1"5��J��i�C��\�S�236�{L�s�qRN�ԁU7�b?��t
�A?I:��r�-�$
� H<�P5�i3t#��K�c�jY�s�)��.T90�\���FgĄ��]��~�����]|�̎jR�6W������P�됎q?��Q��\ 6a��dH�́h��\.��Q�H{l`�Wr��$ح��� !��o���Nn�i��G�f��T�.�Ûn�rB��-B�31-; T�����mK����+�M����k��.RX ��ڽ���NAR!alsG@H4�} ��SƴV�H4���ځ�u�W���r2ݡ���v���s\F�T�_����j���4�\�1�_�߻!�4��V��n1��1qN3��?��x}x��
���q7�Y�����a���t�KFR��jݵIؖ�0	P!��ͳG���%�n���QL�Ф���*����9>r�՛�l�����բ$�jp�N��e�L��y���F.�Q�����]I!<����_Bhpl���4�Pru]n5V��S7O��
�t��{.^�C��e�)��Q���ݓv��`b#83q�0�,q�39*��0�5��Τ� �[�������C��p��a��ң�m�=Q2��8 J�qX2�\���7��).o�����c���"��Uh���AT#O��i��R�̑���,���l(@l��P��1M�`�-k�vO4f
�J�� \�^���k;���I�C<�7�����;�]�
p�\	P^fʆ]+^�������,��%Ώ�` � �<|��;���9�@|�֕����f٨�)���r{^�����,R�Rp8\��С�i��4�j4y�ɱ��C�	MX%M�gsj�m�C�-g��%��_�d��6��x=g��-�@_�/��I\$�i\zF�nn4
(=�f���"�̅T���,����*ӕ�M�D� ��?��"�`���^^aEzc˳0�a��z��3�^k�L��r��e��Z(bE-$1r>�V�ki��fa�΃*�}#?���y�fE�	6�"[H��,��$��a`�Y=4��ZXa����=��54��+i�.���M�Uv�~%��ȅ����.[�{Zq8!1z�m�'E��e��p�Y�]�{�dR5�Ȣ�ǵ��A����"@���cp�yr��\;�����.�K/)P����Y�G1֬�;Y��.U�_N���"��&s+�>^��I���?1�ճ|k'Wݿ��7Y1����Ա���a��g�8��ٱ�A>ݔ#V������G#�J��:"�/_N�<�d��� #ҵ�7�i�(�t��.��P�u�m�.�	#զ���7H����FۇHW��tNj1�.�7�qe*�FT�=�
�R���.��|�R������i��ìZ����h�d���ƭ��0aI�0���4���d��Rcr����&������U��1��@.Oh������ޯa��w\�M�!���;��=ǝ<Z��xlIa6��<LL�{X	Z��L���=D�ﻴ�]\$6>�]t�(�gDdD���`���w�5��`��֑����euԍ�������.���_��Zw�' ?��|�� ���e�'�g|s&wn$���z$���)R	.G�j5��a��`,�Y HƦSQs�o�[���S��9K�>�\$�è�~N G_���C(E�gZ�־��C�6Gz��0�g�&�ak�Q�֍quYfd-�aǱ�O(��y$8�O�wwL��r�,��`4��rg6�����-о(�	[�q��~B��Su�Sy)_�E5:�0#���.�ƿ�He�:E�g2���S	tH�k�N��u�έNR�z���*6��MV��pʨ3�{H|?��Uc�{{ۑ�;uոa&���̎Ғ���d���&�?��'�g��h���
e�b�l�r)� ��x�� {uJ��I���L���&{�Q��x�=�BP�
[�r"/���t��B�@iY�����G�����0�u�V-ک�Fh$�^�����=�m��q�d�)Ů	���g�W��ͬO�!�VS:1�GBݔ'�qۉ�����Xq��)�Ҝ;�"��qyR����G}��pR <���yF,*��������O�O��>�H��$x0���5�l�Xk�\�vn���f(���P�B~|0e�O�DpW5Ax$ �*�s��|i�Tr)���^��˼j]�To$c�ئ��&𔽨�9ghv ����o��Z�~��B�ܔ;�}���ȁ���$!УE@�[��@x�����N���w�Y$�=�	N��N���#�����odHH��ګ���|�w:+I��A�}Nx�*�}u�����F!���F�IN�;���*�R��Ӡ�e�iJs��*h����zrV,E&�FF%)A�,������D�@�t��}Co%�֕L�U���ғ����?T���aۙh�ۉ4_79n��-޴��bФ���7����PC��U`7���� ,����$����JQ?���C�F�P���o%���ۼԼ`��p�t�c�q�0d-x����0Nqx�F�˽��s��CuG�3C�j�p��f�r�O&d���Ӈ4�C ��s�_���:9xy��~�},C�=K������E��}Â��L�8��lD��D�ϝ�ą�(�Dt]�u�C��ͤ�]�+�<Pziǖ�Z惲�ݡ�[�EԌ$X�;�s�����]�^ �Jwt�{ ��zjo�
�sKKB[ �8Նk����A�M�폗4N�L�6�(]1��N+P�[���kv
x��\.����UÌ��C��%!ֶ�1���{���jX!cb~ �Ϡ琢^70���9r������M"���S�����<�N�7�h�]Ds<��|� ��������	�&��ךi��-M��M) �l�q� x�q�6�����R����H��biü�#�'�*�P׾_��ߕ����ǏJg8Q/�0��)2XP-�{��mxb?˒�As6=��7�I��H�r�����y#XET��'%�lU9]{��U˨�є��W	�F����Ò&g��T.{mƩ�0��ǂ�1	���,���N�h�Hy�G�I|et���Kg��wu�s�m�O9��l�`С��$b����s	�m�l�]���Y���BƨcQ�A��<����(ەiAӳ��NkWf�a���&�>p�q���z��G�˧�����ֹ�"B��-��.��!`yfؘO�J���w��Z8�'^VB�j��Ҡw���ӡ�qq)��������W>�v�?�D����҅���%	4����7��Eea�'Ȳ��@t���c���U�I��!z�Z�F���K���₅e�:lcYf��e�D�;/�O�դN�����Cv���f$tn�L�A��HH�4/�{X!�u�=D�I��:ݍ,O�pG\�'b/���2� =[Y�H� ]�z�=,`����W�޵$�/��(w, ��Ƙ^�Kw�Z
�,[������O��.�\�,�P7��_ԭ����Y�Z�g9��>
�5�t�(s�C�D���\E�+h	J:w'Or��PB�~���d�i����gzm${�Wo�+��j�d4f�R���ƧV2�`C��Qz_D0�h�� �dlk]�FI�����<Ƌ3�(��?٨sΖx:���z�3M0��PUK�˱��;:Y���[�n������K�ǣG>�l��<e��1Е�uNUM�'�
����o��?� ��O�X m��������5�e���C]��`����jy&z>�ǘ��xcE�&��AL� X�[����K?�,�1Ѝ�.%����C��hTF|on��<���݉L2S�{A�?g�����;�fz��,Ǽ�Dά����B�i�D��x�=��ʢZ�H;p�>Y�'gST��)��xH:�wڭ�,L���+#�'����C��jҤOb(yAh�Q�,2fY���E9�G���SL{Q�����n)�t��̡���O��FV�5i�&�ԘG�q׺���7���.z%���	8y�N�k����C2��E'�%
rA�(OO=��
'*OU1J����S�ٷ���G .��%��w`�0��	���(	/��7�%ƹO���̯8Vp���3&��i2��PG���C��a�zI���
G!�`�%ږ��E���ߺLs������/�'�J��z� ��(����;LTN��W&$x�V3�%��1@�[�R�I��.���+��%R��A��n�ϒ�f�qud�6KY�|+����m0Ѕ�l����t̆���d���v1�i+��L��T�����O%ƻEw;�U*��ci����B�f�9&�Ö��g! ��ΏHhN����+���RB5K���,�
qV�3��&��4�df�����d����蚓D	awY�R`L��E��Ҕ~�m,�������A o��PTg���i�<��q�����f��.#3�(�3c��+MI+L�}����r �RL�Qf	<���'V�Ne��<z��1E�a�_ĐrCsH��-�lz�|�������L�X���� ��� �01�˫I��Iݏ|�ZR��]����$8���jG��Źy[���-1�۝��� b��Gǝ&�I�jH�~���>@4�&��&=&���"ڇg�K|,�V����=�Fa��qo=��y�0k�5K[���UмL�,��ͽz^�n��=xi�◭<;����F���Y�{�҄C�顟�4Y�ht�!F��n��_6?4D���Uwb���g8���]$�݊�_�TQ�i��v�<��;���(�1����'���%i�OU���Q��4����S�<���F�TXQ�W���3[#�pK�lP�!Q��uЪ6�'���������^�x.N���挱<c��ؘ=ۄ�O��{U"�#�\s�2��(�.$�,��F=�݅G%�Au���6��[F�אuKř:�B��q��#��4U�,>��m���7���@O�����K����W��@"���ԙ!t�0tqI8<,)�O��#Q��z�S_��!N��̦��0���f��+c������+�n�}=���$�y3�-���2�z"MdՐt"��.(`b���>�2�kW�f5�z��8�q�.�ow0��D�Vx@���.ܝ����vZ(�4�w������2�V�*I�]=1�+,E�9&[q��-����F弰���	p/���7��ui��D�EhW�)�Kfƻ�?n ��R�W�C�n��aA��`8:�e�U��w6w�	��4f����b��Pbj*P��� Tp� �����.���:�������7>S�^�tq6%��m4�}����P��:`�Lf�����s��{���0S�
��P?6��~�x�|S�����H
X�&{z�\(���Q��|��h����+o��v幥��^���td8.?_	G^Q���N�d,�9	��Q�/`.Ԡ���u��N~�{l�������+T���o��

|G�_��I�g�|E[F����, ֩6�W����c�_����n�?��O�jm�2�����'[XKaqV(�Irh�i���O���1N�ǣ�&��rP:8���)�WE
�C7Bt���Eg�i��X]��6��4��i��t.��G?�^��e�!���v
EHb�9��=v>x׻="6e�K�۸,�:^�B��v�9)�5����������u�-=[�@l���B=�V����\���h�/HZ�o���l���P��\{kJ�H�����E���6_�gf��Ĝ�"W>k르�I@I7���Ǿ-f����8T��׸�� Gz��@$��f2{D*����������4Ά�_�q&���^7E&��(���(P��� 6ͻ&�4���R�l���q=�d���PrO�ڐ;�!�h�kS	SR箑ᬡ�&~�|��\�=7��
��c�C�v󛗌KNS��I3G��B�w��N0;��R���k'�ά���� �Nq*���������Z	5T$׾F���R�Y'�;���Hr����� '"U�����&=Ñq�b̚�*#�B�;~Xw{|���6�e���W�n|���"�D*�a�Ry����*X�0�E����Q��R�/`�$���1��@�/Yz�m�(Y�ꙷ��Y��Hcm���H���c�����>$��MX(�jy�Y1ב㣞f�t��=rc�W�K<}�_0����G��2z��H"6��F���n]xF�� ���Fx}���82P� u���pt�Vx��	3�$qK�B����̡�Ÿ�����ȭ�N�6���Λ���Hru
�z}������0�)^6��Y��#����5�"W{���e��m�T��Ѱ�,�H����'E5C��'���d��r������P��}���[���"!|�̢`��0������h��#���^�dB�e`ܐ��lr_�\C��8�P!����a�w�\���J2��;^)���8}NHm�|��ཝ���Y�t7��,ds��� ���0Z:����=!�_��͋�{���ff�t����/�������d�ý�^J.j3�ivu	��ìDg�_�CY(U���k+U�Ѕ14�f���������l�/isr�	f�;u��&��$�w��M���e�8��L�s����4�iK���DO�?4�,2�h�i�[�<����� ��V�!� �QJX�fԿ���oĕ�7]�(Exb��	��M8_�����+"7�c/�}���ʥ$��"S���go�|dԡ��r�7"@(��J��Հ�>kj7=f� F��&2B���>�l����G�l���w��v�.�����#uZ��#l�\a�ս?�k�b1 7�ꈒ�ϝ��	�_���9�3�萪ӕT[�1�P�[�\홰W|���F���4y(o��ܕ������#ҝ�R܃�y�'m_C�H?_;���|e��Q@��8UqW:��[x���#|�c����$��70q_�߀��󜱔
�˰��b�څI����'�vҜgI�����4�}��ߩ�������|�p4t2��$p)
de<��;��́�mtS���%�"����Ӽ�/�l�uN;7���Q0��kz24��tZ�ܧ�)OY6A���!�\��镧@߀WJ�u3SFw�RR��ɂ��u.� .$�M��o�V�`� �cKu�>j��7�3d�δ�&JL��_I��ZS�6����Le*��|���Q�(�d���pM��!�Q�0����D%��1�S�B���F�ė�1��B���n��t��� �n��Th�U͘�ޓ�P�h��Q�;op��Ep�x?�LbV�^�=Ps�%) ���1Y�����Ґ�����U�洞M8��]���2�n{�+�Ez+AK}K|�버'�vP�ɽ�z?F���T��҅b���g�oOvD-�),7��Z��?�)롟�dw7t-ɱ��@u����-6�*H&���.��y)��̶�A�l��,�;|��w�s&+.��l`ys�\���Hw�Ё�h)̋�D�����w�<�h����ƾa2fr�����"�$��A���
Z�.Ĵ���z��,$֕�K���'
��G*��aC�)�����oj���|�V�Χ>�<�n��N���-&�l �������%�qe$���W����|1ـΩ|���g�!�{縉�\�"��]�w���z�
-��/�|�"�	���u~rv�G���IhX���wIE('Fu����L��T���a�~��7�y�ko�xu�|q�{�A�ł�������q�k����K(�2�Rw9����x��u�L���T\��{���x ����Uy�X6L&��w�%j(o��B�焔��[a�HA��L�E�R��Gt�"�i|	���f^�i�L!�p�|?5�s��S��1�e4���/�#���)
l�h)y�/c�M�˲z������J~�)4@װ��bh�'�m��fL���>S.ZI�0������U�C�̸9l��{}�!���iH���^����TV_�Z�M�騳��q.@�j%8���#�Μ��G���(�օ �tTY����2��Q� ��曆�g7׷��1>J1�5<'f44�ȅE8���w}�J�����>�w�����rS/M'�/�sHw9��&�.W.M����[��_-����n���2$P�=�a��eT
B��|ag#D�����Z�Oy��3.R�����>�b��jNg�Y���s�����F�@k�a�
ȰDFg���ny�
)%�H�_e�6�mգ���@���b#��H�/��Ɉe!t�=O9�4��v�i�<W�gweQq�r�G�4AU��d]���$'%l�YN��u�Ȝ��rl�[�l�����7��������߰kv7��Z<Q�R�v0�t�&�M�;�xz��#� y+t��N�p'z��/��f�h$�ƽ����C�5�D��Ƭ"� zG��)v�3g��\��&� �:��D��8 ;/�h�^W�{}�anͶ��C���Ӆ�"�G)I���<1����9T�O�"2��,9k�!H��L�B���T+�ba�%�ڇA-&�$�v���
���@@����j�[�s�+d���>-J3&���@���൹*�)8~�U��0�67/2�X�H	?��V����)9�1m
�?#@29�qCm����3a�� �0i)Z[~���;жN���ye�K����k�SZ������p2�L������UȜF�x�0��ו5�[$8/QzQ>�50D4�)���ӂf��=�"tQ��|�I	���fhC@s��>�
u�ݖ�;����HD�#���)h�	��U�|6����9��!N'e曷EO3hf��hl�ta��W�#Oz+���[8�Pf��DA+C��q��͸޾�/��˙������My���UN�Ұ8�{�����7ϔ��`.=��31M�Kv�&��9�r� u��mDqC]��.&��9A�7X���W*ӧ ���b��ܣ�J��R~w�o�XZvS�C�p�l�CZ����`��*8�ø�I���4B'��N�>37�=��j+�7���[ɱ�P�ѬJ,Ɋ	6�88;T�Ӟ��ӊ���j}N��l�w�?�B ��G=f�kn!KS��?����z�ձ���ڂ-GL��WKvŲ� ns�6Y-�^n5�ȡp�d��d���g�ӹ���پ�͆���a��>�v!�^؏_-�&K�*|����O�����@�5~`8�R��rd�&u���o�2�N)��d��W��\�Z�D�����r�X��^��SX�vj7(-������-Eb�垰���5�_��m��O��/!���M��l���dЁ�C˙�NƝᅅ��l+z)I��!0�K�_�rU��IA,��U���>7�����n�=�_�� ��0֔��5��F{��7k)'���X�z�#��؍�D��u������ȣ��k�#A��.-�/���G�G.�W�Ewa��ݘ0d!����:��HL+�ơ\uw��h�DD�g�
��j�6�W��$����V�tv ��b|�@��k���(l��l���j:��3�G:}v�$j���ќ3�n�,\�Ig?1�X]o�?YyFw�(i:Cq��p�>o�&7�ʡ��T�^%�7}�T`��{C������1T~�dj��Ȓ�Ul+�ǚ`�2�M��'ɽ� (��q�3�Tllg%�x�������"��3|�[	��?�L���WR��;N �E5��8,)��;|�9x>
B����X2�MG�sH�\*dVqUO���9iEJ�􈢿Hl!MHe�n��,G��# ��M���f�^j-O&�u#���L�<�HY@?���C�W�����F�=�+)�u�U�F�r�n���������m�5�����p���Pq�u!�;�F���Ҝ5��i��i7zR�H'ǘ�,���V�{���V!���BN$���J�Ja�;=l�����'P��Kq��bo��Tb�𨶴�8za�"�p��C�^I�O82���ɶ�V�.�1'�EjB�v��R"o�xL�_Ԟʠ�UjBb�~6��7-R��&��� TFɈb�$&Ъe���q�~�v����Wii��A�隋��U�OjV�G9!��@;�y)��	�gSs\V��x)3=�{���j��fg���TB��.�u�;;��F�u(�5�JZ����PÞ7`%n���}��U^�V�"�������l��� 9���0�����|��l���E��Y�L�e�>�˱J�4oW2/W�(?��A��F�,:􏮛aPt i9�A5]�>`����U-@�H���6�D���Z�_�:^f	��+�s��<��l�[Is��׽�*i��-fG,@�,`t50q��7^B.>X���tؗ�l	L��/�_�#|����}�Ii$Ջs������3\-�vt���= g&}�M��G���V��1:�0_a�yX������H>�2�����@l��0[V~���9V���v�#T"���y���i)������N��x9QԖpyPuV�#j۰>����t9�(&�V+�n+{�W����ƘL��r�.3j�
�@��z��jcgia$�o$��U�y{������X�M����x�!A� �ޫ9l��˟�}.#��0���X�1�n$."�f5�v���:�d���������1'qͪ�	f	���wТ�5T���3I"�'/�Yid���Ƃ۽�����A%Wś��9A���m>�lV� �6`k�*4|���Hl	�?uR�e��T-v��zNW>L7)4V�V[}Pص����]�?�'�x��'��~�ܰ���d 8��n,�ݳT�V~����� X!��g5�*��e�"#���k
O�+����5��u++�3x~6M%,|<A����*��+��L:4s�a�0��AS�Xѻj���]Ψ��+��-������(���W��J�h�D��!R� ��O�6hl��,`�A�x�f��S�nD���\�#N�4��\|����0C۸��w��W�7R�9$QȪH�h�5�bs\��D$cy�Q둞ō������v�So��,���v����d%�օ�KG���l��ޚ/�z�9V�W`�(���p�ǜ�Y8W�����I.��c\7!����a��1EQt��Lj@W��i�`J���ռ��뢽��O�g2GZ�$�1*�-tꦲ
NO4�t )��a�y5�`�8���c�=y�K0`�ʛ���A��j�2���<iyL��'�	�0��R�ώ`���{%_���7��X��:�$���A�j{56���.�@�"`�tK���+y�?U�e���P6���I�I�Op]&R�wC|�X��7Kq{'��2�h���W����S��Z�K���3d�e�7�L��a�r�}d��[��U���C�����-�Kj���W3���|�̳T(�Uv6����Lr>��'9����������,�P�L ѯ��#�k�:d V��OL��A�5����]��ĪO��KUv���2��<�Z�1+Eg�<�!��dT ��aZ(���_�YNYO�����F��� �ɪ����Cδ�9�S�+
b{Q��*K(c�2c>�[P6F�'��/T"s���_�!�J���&f2�b�/�"��[Ƿ��.�֍v:���;�x"0U<s!~,f��[WS˞�Mv:,��$��$ʟ̧��"�P��m��M$���h�b�_���vQ9B���V�Ff���ý�У�r�����<�h����h� �<���Q��y(���k�.�Y~9?'��U9\{N����L~�~�X7:K���{u"h�x�p3V��x ��˟B��@C�*
��u�z���~��i9n�ڊ��m[ō���O��&Ǥ��Ak�ߞ&r��dv���B�YJ �������\�R������ �չ�+n�m�f���Q����ň�.�}�1��Q���R���Z�	���y�<9�EL�/	A�e�d?���Z^�o�
�nM�J.|k�����|2�b�4��&e�P���W	� B�Q~~���C��u����,6yR)�Ġ�WKı�����<Ѱ��_=Ʉ\���t�\���1�'�^+gM�nHc ��H�zg�����wM���I*>��[�ڃz�Z���<�&�m	�3��s�[�*	�@}�
G�s�t>�zf�f���_��@�&;������x�KU��n��t�x���>�i`�s ੌ}�h��rl���*Y"�aY�=`�����]݇��G��WA�F����;آ��I�l�d��.�6�9�J�;?�OC$�]�.��l},���6�~��_��U�g���v��v� �Y�NbSfҸ�vۇ ��P�c��b�H��$�]�Ncp�D�$QC���
6��A!��G�!CS(�H���Q<�b$����Dia�:�����g��.�O���Sa+�G�u��;)��1�r�u<27>��4p��B`w
��5(��ؖ=7�WD<�a��p�=1����V ��(֜RP�7>����')j��x����u�`b�p���|�L����hL��9b�=������Z�v ����ɛy�%<L�|�d���l��z	aR���� �x䳌��=�nד�5X1�*V�B�09R��zN|��E�y���/1J�a��qG�C-X:�^b�S8y�Ac�,~ɜ��l�����S�j����W��s�d������C|,?�0�o�#�����O�u��o�}}��o/�r���Fn��2��&�֌KQ�������)AB���_���gN�|O�Y�V���?Z�^<DsգGJ;~�:����xe���>���F{m���6�NP�N�o��}5���u�4���a�?9�'�m�S�t��C���0\�2��z|z�j��2����񑞚CR#�P�������MH'ϙ���!��B�^��q���r�t�����Z�v�Zb������FA�d��r҅|:�g�����"R;y�K�G"*���uQ��E� �Oi���㾹媤�9�"K3A%g��-�����H4eq�C4Q�5���w8\��I�XA�FTh� �~�ɸ�ۄG�L����q��P�Gk�����烰`��h��ο��C�O�(l����c(�4i��n|CɎ}�h�l6����R���b{���}��WE�6��x�2Oc	���4��R�)�k0�䛙����̃*7�fE�x\�ء���:�}�aJ����2�K�9�O�*o�x�/����}l��`#g�2h�Yr�p�-�n4L��9P,<0�	���!d"��q�EtKTZ	��-��bA��r��ɟ,�$r�j�x�{�u V� �����;�k�^�PƧ�(���|a�[��%X���GL�2��I�������a���i:����F��>AǂdF
�Z� +h��8O��ۦ�"��A��,���`g�T����1��ͤP����P�8�W�v�"&+���8���VJy����?���m���.�B	��o3N85��"�xE�k���1N��/5����4?m��]���nO\j��.�lUB`��V"�Ǹ���Iv,���F�8#�Š�Al0�^�hJkA|ݔ;���ؘzUOJ��?QJ��@���n�(��]��ˎ�VH�u׾U�>Y?�7S��}\|�ִe�]�g9��%Y�&�\d��������TH{��#�w��!KɬP��@ܮ�^l���H>D�l���3����_�TØL\�{�*��i�g&��T�Ԋ>��|�(��"�S ||Ũ�(z���JN�,.���ŀ�0	>zH��=iG=vNm�0m�Ȧ�z%1��s�/YK<8� ���F��~���M��D��c ʲ�6�;�B�^h=���r1/G8�)p1�s�9=����pQH4g/r�l/æ7�PȠ��sj�
��[��_�
�]֗~#P���U��a���[Z�
0�#>F���-�y�-����I�*�z@�v=2��iK�ǫ���/ڒZ�M�����z<W�t;���F��'�{)�A���t�7iA���o���%1䑴�E��<���+!�!��d��V��,%B䭴�#$Jv�+I�2���WD��o�u;�nn�#����,���Y�~��Sä<�βd�z�.��5�R���7�6Sl3��Z�Jvq�����g�Վ8<�{�Tj�%M�:'��uߜ�8u�F��՜��?C�yYE	�ym�E�M$>�43���i�+q�|b���x����2^c������o܆�\E�[�ݵ�|�6`bGqX��B-�	4܈^�Ƕ)T>��F��WedJ�^��-'@���k�kXZ���GN;�󔓼�K�|qy���,��N�Em�=@$N���/�A�5c�yAt������P}���J�����L�,��}���͋6
�g-�*�/��    ���3D`�Z|��V�����m���r�A��O�v9�J`V8��(E���R�ѿ�$
�^>/�M�!0L�p�    ����M���Y~�Bd}����*JL���������s�,8���2���=����1�J�ί��(��c�D���ɓP���8�4�*�S�U�6�ܑ�    � WÏ��x��k�M{*���"y���}Z�i�<�q��zU��B����    
�!�OЏ?OI<��Kõ�1B�}�>p���َ�/�����΍�����}&����XT[�ԙݔ�xtKL�'?��'$ט����� ����F�R�+��^(����*>c\%�gUp�ɘ�>p�v��7Z��ċdgr5/\Z����^����.O�%��'_z��^�L�`�9L�rc*�.�Ĝ��^ǤI/O:�Yo��4+�uŊ���
�2G�Ⱦk�C��m;fb�~�2�d�����2dx�9�L���T�8��2WK���F�~
C�h�?
/|\�M����$V�.�ʷ�,�JƲ��h0{<�"҂�ԾH3�S�0:?D�Ë������̢���E��dJ1,���5y�L�q2�rj��u
�f_�ÇMU�te׍4��J�RCU:\);�`o3��Rb1�U>V�����:���z�G���ȭ��E,'Rm�Ͱ�]!�
���`Us����͗�P-�bc�+P+�s��J��8݈����d՛.wbag��K���"��v��%��^���d�܌�Z.#���l��F�m_�� ��o���Z<v-�̩���(�{�)����ΡuNw�K��0�yoʩ�sy��C T7W�n�ŚHe��gn�|ݳ����yNf&��5����0܊��>4۬�s!����S�	ޚb�z�O����]${.S�v~U����w6~28]ue*x'M����]�O6���2�#�#?O�҈3Y+F�sn�8��$@�l�����2���.����&����yp�4N*��[;To��b�[��^r3�ۑI8}���`��v��k�=	_�>]�=T2q�^�D�g>�)�����$��I)֛����1�le��И�[��9/Tyw��f��8dz���5u�֋g�"x���Wf��&IM�L[��t�q=���IK��^k��8^Ļ�B�	� ߲�>�9V��E�@z5�ʆ��)����,�x��L��D�ԡ\�'^���L�-N�ϲg�bG����:;���.�vSy�Lb�1�9��vJ�P��i�
O�����`�Θy{Q�&~Y/�t�L�/�`p��I\M*oЂZX�;�P�+����on���3�<�:��.s�C#�Y�r�u{��&1�ۻU�^�(�&��7lz����k,� C�k9<Mv9����!pˎ�z��Y��O]��]���4=����ӂ4tń_��]�n(ej�,��+�*C%U-N�a�b�,1�l�����vG��/4��:��vbÊ��G�
vpqI�>�h!�m�zQ�:f.�����^�U%�}�AH�$�Ȱ|�V�-
�cc2�d}�`��@7�y������إD����*c.�Wj'=9g��u�"�j�`W�0��l��='����a��oK���$�Z���rhc�<�'��3��H�p?j��os���;=���3Rt�S�7�`@�H�x@�����������-i4?O^_���§r@)��d<-߬��bZ3�6[cv����o�?>���L_6����ҟ=��Jβ�Lg�ςZ_�Z��"��(��ܟ�-�S��z�.�t|�e���:k/8�b�fxT�`����4;�ճ����Z��j�������C�CPY��)�y��A��C��`��D��[�K:�!5�hC��`�;��"���QP��i���!�n�S������JJ�����1$Cg)������V��ь߮��[ �"1A6����7�<����^ٸ@:yX/�l�����q�P��F>�����;�>�x'��B-/m�J��*�xݱt�����܍ |2�O�K^���IŠ��|6�=��U����[M�n���g������~�Oϳ�ܐ\�ҁ@m�A����wj~]��+\����	�H��Y�E7L5�k|��ԋC���"���[Q��Q�x����^�a�Rn�-��9�'���G�}�#����=J^cB �/��+||b%/�rm��˿�~�C�E�q�-�D�K��(�'�Y�Z-i����DP� ~�몺�mw|�Y��$�T�{o�:��irl1�ٔb�,�7��t���@ތD�iBV)�<!~{��jON�h/�zm'Oԧ�z�x�ߵ���$��m$����
lT��@�֦j���^8LgF�e��'3��ʷ,Hn�1D��c �iC8>Q���Bw�&���8�A0"�I�z?0�!�޿/��ܘ!Ά# VE�x��Ψ��Yh)�Ά��;AU�4��� �����NBo�Q�5�o-�^9a�V�,9�����Y�@�u�E�</H+�q�8�	��=U ~��I�1��kz�kG���r��?\�S�rl$>4����ܛW����SC�������l��ʂ�UFb�"cq���;��cwH1�I��e4O����R �;���D"z��U�D��O
̬}�t-����|@�[u,�)]M_Ш\p{�5\4���[W���2��D
�ƸDkn�Ҏ�wc�o�?>�Z�'�#�m6Nz[�
	|W�d�#m���������{Tj(ٞ������WҼ��+҂8m7���rzu� ��s#O�R'��E��2u=���]��Nא���9��V�,l뺳��t;���wd��w=Y�����vY[���%q�'�gP�$��
���%����Ja�)xV�h���?.�a�V�"�����[�`��kfk���o<`"�۲K
�:2��B�v�:��*Pԙh���:���3�\�(�:���!��"��qTu��Y<����gF�i�,B17�+Z�0fTţy��n*\�N.q�Vی;�;uV<$n�[[޿�~=I� C
7�y���ˁNڼ?��B����X)ck�)�����A0�� Z��k��[=�x�:�O�	�_�EW{
$�y��m�-�����1����,�-S�d"�RKt ��y�]맋rm���i�n��,�a�2#�/�̗m4����c����9�'��L�@��GB)WP�b]/W�oW|&3��[NC��z�G���=z?���Pt�AuQ��ʢ�q}�8�q��p�V/���Csڦ��k�&b�0�|E�oK��G۵�Ҹ_Mi� � Z��	r��0N�u Bc'�e�G6 �еd�m�"�(����ݺ-* ,���h\]~-�U`y��҃ڢ�;<���}�������)�`k�t�����L�$��]FJ>E����Ui�^G$�#���]ܚ��0�k�H���ҁ�^�Ψ��i㗐&t�����Ee3T�p[Vep*'`���V4GT��#��ެ/�Q���d����n��A;Yn��v���)�.y���5}��0��W�M�������1v�'��Lk<n�f�?ӑ�[O�� -)��!�v���.Z��9[��o[��F$��;�܊�os4�r˅8��.M�T+ǹ��(c�:�[Nl]\��� (̎ȼ-���_'�%E��������t�� �yf�4B�auP��.�VQY(�`�)��-�P.��=⪌���r���b-��A��!B@�I�ݥ�&��k
��<�Y��Ԩr3g���m� [톶�ظf<�[d�UҍMˬ���~i�z)ȋF�-�`����
�����'MBq1ȦX)^��ԛg{��)�+.�/��P�o�� �!ց^Di�l=s��Ô���鋀�o����QT���<�M�[L!Fg�7�Il�'��i�oJ7��}Qw!~[:�g�Ki*�`Q�n=�Nv��[�4�l�d!A?�ϙ��'�&Ct���SG|��T�g+�ݡ�Lt
Q�2?x6��o{�t77Gu��ގ����=96��-�l/��3���IO�j�^�H�u�=8#�m�ΫbM�#ഴn�]s-���K[�e���J�cV1���lξ�L2�)tΣ�#����bMb��Q�^�]Pr)�5Q:���u`_�} �x,�	��	d�^} ,�´%w���᫶���s���]5-�^h�	����t�j5 XN��E�'S���GQI)������)��mr�o��q�8��o�Pyأ2�ظw�A�+t?pX�$@���@#�lB���l>ˠD����"h&�[J�z89gC�v�"(��`W\��lV=4'�)���<=o��gM������Z�ExvhN� K ��3��H[Wr?�ʳ�o����;����$���S�Lϑ���H�$��������-t ,i49��\_��ç�Ͽ���a�i߬	̲hS�j5[�����]�?>���|#�����1H�l���Ib�ź_d�_�j��.��"��ɕ�%�T��h��(�	|f�k��z
�|!�
�q4�-X˳��(��ֳ��[��[�j��Ӎ�®K�J���)�T������`���Si7K:��)5�v��m�6��$���_W��n���/�h,]�����HJ��z����Ag)Zz��nV���s���ؤ��"1r�����;�&r�^�_ًI��Y/� 1���ΎT��������H�>�"^��fr�2�mEؽtu�9��j+����ߍ�*6�O|�J^Ѩ���"������=�j����"��n���R����_c��~`��L�ݐ\�J�K{�J��|�lx_P��b�������F����T1D3�Z\��NρO����<��j쵶����Q�p�ߧ��s�@;�"���-��ɝ�5�&mݠ�/��`bB ���"iw{ �`��ά�D�E�C�z�'�`�A��"�-�T�R%oW����IO�gt����rd���Y��0�R�ke�<��uzF=��j+*�2��q�2۰b��6�IN *+.�B)pZo��1ax�Өh/�v|4Iҡ�|�~�ӳ���9��c/��l���@�)]k�����OgF6�e���'3Q����l�1J��m	�n[?!V���Le�4���*�S>0�[�v*?�3�̱=��ۓ/܈-QM�u��ɯ ��l~!���ro�;Q�H4��)B�����B�ʧQܰG�,�^��W�+h�C��=P�x�V�v� a9�v�>���Y0f��A�%��H}�gN���.�~?P�_�fe!K(�ֺ�Y��h�BF�������j��̄�YuK�z�~9��	��k{M����s,H�������6L��}G��X�H���2�/�z
�����5P���Yu'�%`E��vv|�3P?��o�Z���͵�D
�9�Akn�Η�P�s���Z23�8.4l6���
yk�C�u������>���\zTj:&@�����Ȳ^�|
�*҂Ǒ5���ghN��,��sܠ�R(�U�!p3��[������,����/l�E-��t[���~���w==T����ĉWt4v1��W:U�8(�F}�۟�
��M.? ��Jm�!���h��Y2�'@k���!�"G%���J����kfz=>�o<f)�5ڲK�}?2�m�N]e�.��" ˋK5���Ź��뿁�#�(�uä�$/��"��Tu�X<����aD��m�9#���|p�"����yaV�n��N.J��.�;��9}#62K�U4l��'.Lg��7�t����C��M�#����N/ia� �������1��M�c�E�}�<�x������EW�c%�y�����d���1Ϥ���'�1�vg"wFMt ��\��&A,֜�z7|��<��3f� ļ���j2��<�a��$��4�4��Iv�K��ME	.RY�SJЬ�oWp��l�OC��[�d��J�lM����[̋��|P��i��i�.�v��w�&�o���cʎ��f�
� {���3> �gYo}F۵�ڳaLnq��8�&qT��3�r�_�/N95�j�I02���Q�k�^����̱'/ ���cYV{9�HfE���|ӣ�<�V�e����~.�Ftf򪢥����T3>oB��~�FJ�漡�� l\�YB#�L�L�W��ȶ�]�s���-�^�����V봍C
��4�^m;C�lRY`q����P/{+0��˯/��u��d���L�nw�C=�(��vrS�)�����5�:�2���7�񈦚ܟ�7 g�)��Cg)r�h�5^��ذ�� h"���f�w�z�.Z��/t���o���F$��!e���1�](zN��I��)ǹ����'��8�[a�sZ��5/3lɼ-���Y �"B��������}���/lk�"G�oN��� (�;�b�'�LĘ�-�B<��/𸗌4�F���d���\��9eQ�^�Э�!��*����<����݌t
?a���`�劻�аl5
�Vc�]؄Cœ�֒ez�eq+ȋA�v~����
��Tj���|uc���fLv����d�z�vh���.��r�OJ!�!~�Gi�s|�H�Ô�4苀�g�5Ԏ������<��_֕�)����Y�{P��?�
�i� �p Rw!i�v����Kig�iQ��[�Nv8�]����l�r)�B�ϙ����pu���W�Go��6cc+��]{<[�8_DN�n{���"Gu��؞�3���;/ ��+�i5ȉ?���CE�c�n��p6��G��y�b�6_b��]�y��R��?�P�Nj��,z��g�@H����y_��N4������
/�8�*���|J9Smΐ���+��2Պǒ�-����ڡ솲�i��2���t��֮XD�`��h�A���    f�!�9v
�� ^wR�AZ~Y��n�.j��J��&��=�j��<����yz>K��$�$2F�&���chO�oA��iv茴AO�jrU��x�����+���cل���A� R��x��B ��b±S�W���f׬�0ky��ss<ߎx���`��ر{�y���!�l��aĎ��d����s�'�j���-�*��d�^�H�%12�݀�g�_��bY܃'Q�o����LX�Y�J�~���q����e��-��걥�{�=��4��丿@vÃ���ؓ#T�xǤ?����"j4{峓�U�8`G*,��$���k�y���T*���zȇZ^k�����f+
���Y@`��{�v���D�!�0MWY�QyE���=���EtI��g �D0u��c�u��}�/|g��mcE�PR�	Ik��O�۳"}�����JW ���b�&V���+$��U�!�~�>2�2Nx<�jdawxM��<�yu���&X�4�n�����Cm<��g��n>��{��k���=Q��D�����,�f	��W�V��o5?�J|2�~�F�Z�����
Y$i`�r�S!�����7���	S�!X��rf�]$[�R�]x�Jt���PQ�Ż�vv��A-<,6�V滌�<�����)�K�s,<�' ��rW��X�W�I�
�*ƑHh8��oOq����pW^<³����p�[�CV(F /�̾��ث<��n��~��R[h�ɼ5�W?"�H*It��v��x9W���kBT�>(6���a0PihϚo� \7'���$��t�e���YW�cΈO����E��F�s7���+DA���?c����}�ݱO9��U�R�n?�#�/�-u��R�3�Xҥ���Ix�Oj J���~�@L�.U���VS�@��r�<B������ڡj�'f��%f���ӑQ�oW>6�2F=�3(�V��^��P/o~�[
�ғ1�f�F������(�Q�?q#j�L���/�)�z``�7ujz���"��Bi����~:����L����Q8=o���N�pL<���܏��7ü����P�Jc2���@O�%)�������t�#AU7SL���{��}GZ=��q��PHaOY�ɔ�� TQ�IS��*z�D�`0���"�i �y�/#<�ޟ��i�cY�1-� '��������h�Ϥ��F�Yh���Z�
=r�M;�sX�u�!�^�y�j��Ɉ���P��2v�E��񯎜�D�!�2a�03���������F0�n '��M��\�Ӌx�
}�?�'���$��b����Tg�x���:�p��(zܬ���s�h�;,��D}z���h�%I�q�}$��y���Ѐ삋���b��[ʝ�Rz�;$/�mu2ǣ�m\|+�����K|�� �r6���4�aB�{�31�.!�yp̗��/�X˅	u���d.�_6��,ޯ�w��k�����n:��W�i2�p�	}$�Y y�#����"�2x���6\
��<�d����6t5SMi���c��%-A��sJ:^�,D��58�g��;%%�T�G���^0,��M�ͣ���
s�e<t���8���+�0e�C��p`?�稼�JS�A��jk�)���ۜ]���t H;l��1�GĂ�W�j�sXSw(U9�y�W�Z��@��ĝ[,�c>�E��}iؒ⣎G1�����?Qؖ��*��:�����#�K��~3�ׯ��W޸o�-��[���L�4٦�Vw�?
+B��V4D��(�~@xtq^�� ���"�}H���I�ʢh����Qc�G��[Y!����}3V�o�lV[p,]F����
4@�]�V�)	>u6�dL��[ �&�J�\"ri]�vCL>:7챸<~�O�-�=���Ѯ��&��Q���ƥ��]_�C�!�uXjĢ&�
!d�����N���c�����,�hd'�0��3�;x^O�L4�-���Ê����N�Ѱم���)��;'QM.:P��j#f5��D��!�J��.E#�n	#��FV���A5G .�|�9��Ch��������$sȫR��
<{�4��6_�������i�~C�G�!��;qH%z���n����������ɳ����é���U�R4t�I}ԡd)���~.���ktBp��n?TTkW������]��F%�~�����%�7�o�9��p�_��F�]]����V�\�����<�T�\�rd"��%�+�-���)��
��D�V���ݞ# ����X�������s00�(V<�\�)5��9�X����0�BMy��`h�s�;>�[.�iǢ��<�{;K�ě�[�Q��u��0ע�ꖴi	O����P_��zT�۪�v�2�3��v�����N�[H@�G��"�p����|��m-<{Hq�SZ��˽�y��er�6��
�:1�Y0��EH�����a���,U������D�f�X߼���ق�`�C>�����vVk���ɾR|����dqh-�az$����-�_��8a���^g���!��6���"6���2K;xG��t��#�������MQ��X�¹�h�.1��2s�0�Q�5Y��/��Y	�������t��}�`�bF;���4���
,�v>C;6�?�%�5����gb�p�]�)g�5g?�8�%�Y�St.=5��ӗT�9E���sy)�Y@ӨKjk�����I�����\�:,�RIy`yt`:�@���P��!W����o3�\U�
�1%F�0�,C݅��Ŧ���~�s��c�����4�UL�[��0������7�X=#,��@uHEr�aޱ�^��L=Mm��5Ofd�@�7��;�ʅ�zOS3+���2ҏO�//M��P�6A�����pԮ� =����Q����2���2"wF����q�Xj�V�L$3N����2��*�w,vdr9�^�ϯ)q�ޠ���hpխ^�joF�u�c��e/�e\���!��ʟ--��1T�kpI�.�j�[tT�^O�Y��?��L'<����zg1D�k>u&g���h�vG�c�f���*�cycl� ��p�ӝ�ըt����;g�2,qf%����^l�(���F���ѭTJky]$��Q+���q�UD�W�Loфc�3�ڹ I�@y*�J���ժ�.�<c!.�6�����m�f�n3E�)��t� �����#�p����/e�pW]���;O�1�\�H�!���ö���P�>78Ny��)}��S��"�m�ڑ}�Rԙ�����$�N���~�/�}�� �(����3�M�Y�L������p�I��"5��V`�������Xȕa0�[���(���~qr���p	�J#}�W�VT=Tm_4��L��_�)����~� $0K�+��j3d�Z܊���4)�
R0�"�	� m�T�ƞ0��>'�]Pկl����f��ށ�/m�� ��͓43U���eY�I=���k�����E�_7��-�d�3Ψ��N�Xͫ�d���0ǜ�(�ޚr:�	-n+�^�Rԏ�O��$s�+��������,��W(�BG���$�I�9D9���M[����!�]��N�GQ��C1�3�,��Y�	?��Ðf��H��*`�#�����Ɖ����eD?��,�t:�9�Y�s�P�����G�E�/X�O���okTn�9C�U1��kl��NB�z�4�Tb� =Qߖ�_��rsj����I�֎odG�AS�2|1R��v����%�5Ʊ�-B�oq��Msg��(�h��=���*�"u!���4����B��l�j�ɌY"���(a�]���9�!���ZC�4Y����W�H����M�;	��=ѫ^=�q��?6���A�,D���_�����X~��/cy�@@)���	+5S��D�E��QH|�j����	|#�����R�)<�b�{���H��u�q������ ��x���J�Й�U&u��%��
�A��}�Ib&ݘ�O���_:��)������'�ھ��rj^�^Sz8����F*oZ��Q{Q���@��?z~w+���^�M�?)gd�^4h��"qx�*��O���t{�)� 0"���ll���u"C
Bct���!�B���>Bt�tk��q��gl+#A�S+a̍���^��}p/���,�N�CU��&N���̢�K(Ù���k[�3ӵ���d� ��)D�"	�4�%SwJ���{�=L��Z&,4�lm�=/�<o詿�E�c:
���l�&ڿl�_�	%�����s)���Β�bT��!�y�oaҾ��W��Wa�Cnׂ��x��a�i�z�~�0C���&uۜQ6_�m���R�TW��mٗ�IA^����9������Iz��8L�v�fŭ�ߖ;J#~¡�xvH0�^���篆��ʌ*;�i���H���|�!|$�x��>'?R̼b���Q��;� �'��s�m�S �B��3�3�����NBY9��Xd��u�5� `�>�)RNsb\s
�A� ;�E1OR=���;�V+���`��Fh���Q��b�bXo�,&DC�%�F�P��[\��,G���˰����<�J(��6�)rM�����)z{�ڰ�7�{ho�V�b��8_zfN�0�Z	��u����^YA���.���9�wr��#cq�4Ab�^�n@T�G{Ɯ�K�V�^�v?X���_��hj����fq�m`�$����^;H�<��G�Mň�9G��Z��X���O;�#I!M9��Mb���h��Zk���nA�!�DDK��<ɑ��X���*�Yȗ�Q�����q����e��X�3����a3�w�]"?B�T�!�bJ(z��~�� ��[>g���~��@9�`�	CZk�3C����Td���ܥ^]Q��W��V�{[�;��0)6Ԧ�r��f+p�-Q�p�p�[��6�1
��Q�PS����r�͋�efO����!Y�k�wQW768��J��z��SeN��oڪZh�&c��|N(�0��	�Rw<�N��{��O���)���s�ȫ�FC�(s���G��q���F�UR8�W)����7��{���cDi�������Ң�¿��RX^�-����}�i	O
��Sy<��|#�`���eٛy�S|�v��S$:�/���wh�D�9�L���k| })�Z�)�a<i#��˾��En��69GB(���Y����_��l�=�߃�_*l��;�Of�pT�A�Jԭ���d$�5���\���?���Y0�R��x/�1��$�1�N��ߚ�eyzj�L���m0��U�����0(9�A�k��!ή\p��ց����V�#���?b�,�n>?2��d����a*�����T��U�@O.�����v	��"��{����`�aTɇc۹�T5	����r,�8�����]#Rq������n>���)���Z��&W�� �\E���<_zҮg�
f(!�CG�Mx��
�U�}H�(��rG�9�đ��a&�g)ENv�1w9�spD�����Hq�� &���P0	���F�݊�l|F�	��涷2��h�e5���ଚ12)��Y9N9ʿ��[Z5)�D�2��ce����8��p�譩x��t'�~4���|X�f�8�p'�����JaJa)'D"�:��VvrH��z�y�x	+��Y'�'�$���{�����7L�Ql�,#�/>n�,k׹-�G�u�-Y-_{^ ���{�����b�k�i�\�b��ޅ'Ѱ݇�A��;�92FRO�ͥ���aUS���oZ���e��E�^�nho��4�.�C�v��lf���=���@}�,`v�G��E�4t�{�t]2x�Uzs�I�pn��0�ANv6�7Bӵi�N&��>V�a��:r`�#z����'���s:��\�Ap����q`�tNU�ɈDA�9&1��1���C4�Z�8�Az�(H�;����oM�;�Y���{�Ű4hVL��z~���w�$S�~9�T��n`ԭ��dO(�1gޢ����K`�K�B.^W�9eb���`^�ú�r�?����-����
��V�թ,Ֆ�7-� �Ak7$ �`��!T�� �y��TS�&����J#�T�������t��ĺ��<�Rr��E������[g���i0����k�fAx��x�)Z޲�kO�g��ic�:���(&����S|��d�o����}�X

va�ue!%4��:,�9��D|:���_���z�.�7Qz��D������Փm�@$쓚#5�r_HH�?�i�E|�k�<�{i7�8̯C�L�oNWM��?��-q+>R��"e���FK:ɔ|d�.�_'s&�f N4%����q����oU4�h��)Y�^��j��O	8Z�aH��hy�?׉��#����ߵ=���X��"�?��ŝLP���0�3kCP�T���pދ�J�&hԇ�w'd�u�ƁΎ�N�I�?�!�d��b�H�']\"`�f�I?���+��:��p��d$��Z����˼��ͩ�6�����~&��ʶ� qv�2<���CB1���L�d�,��2�qZ�4�j`G�qp��?v�W<.H0��R���no���z��Bf�ֺQZ �פ��<��dm�\��C���/�x��{�L(��CP%��ei&Q��Ӻ��c�L��t��I'�vb)�X��V��b*s�������E�F{�m�����$��}CX���j�E���E�"�����k,��/KWJ�Bo����'�:�)�:��ҕI����[b�"���@ܕL�L�4a8�C�<��"�?ˑ�a"�ϬM�v���l5�%�h����K��>�g���}�uz�)�%Of�"}|��ʫ&��;7��Ij�y��ڬ�I�~O(��Y �ؑE�Zխ���$�*�"~�$�M76��>	E�2�R2��:1�}Y��%#�u�H�ʐ�^7�Э����2ON?�;Z{��=b@.�Ʋ���("�}���5-�?�RG�G!'���6�.�̼�%�}���	Y�ϙ���6����.�VOka=*�<&���/Ó���9�v�j}�;�F5��EMŦ��F�\�Ǘ�C28E�����c]�UN��.;9YG݊�P�n��~0�p�#�j���������BLȀ4���z��}��IoC�l-��m�C�D�Z:U����Y�n#��o����6M�ju��"\���k�ˉuj	�_�E��p���eԧ]���A/���p����})07��J%�-�s�}eu��)*`?�f��\���`�ߞ�;�ys)�6��(I`Bͦd(h�T��/�=����-�\�_�`�Jo� �n�j9z-�G�	�Q"���K�W�!�J8J��Vxc��9��F�*R%��@��7$p��)�����,�`+�Cl�q�
��H	9`RU�xs>v��!�2y�dk�ś�'�>�{!��W�k�A��\�:i|��׮�ةV��2>����K�
�y�+y{�揪^�uN$���X"������qe ��F�Μ�p����|ͭ��+?�y�D(k��9�90�^�s���Lv�Y*�ꓦ.��C>�\�����4uW��P��	��B��4�CV�����K�NYH*���[�(څ��HmϹ�,r�-�/y�F�T���������#�*
޻8�ga+�Yk�|8"0�+����K���N� ���ǔcv�ڪZk)7?}�6��c�j�L?i�1�����D�0HL�H�M��9�"z��_2 ���k��tj6e�e=��<����7&��G��P0�$��_2��N�ܒ�>���ݴZ�ĸC���QŶ�4*�[p/�T�	�h�s�����y����a˴���N�R�Ȇ���~X����A�q���Ep��ֶ�G~H��i����>�i�n< ������<)�����a�8�E��5�bb[˔��vJ��׀�43�%�1pX��%�>����{T 0*�y����jb�h�ǐ6X�X\O
P�$�J s���~=�ىC����E�����A|��E��]�#����Iޖ���d�b���mU뵶8̂����^��j���1R���QǄ>�x>\�G�J���d/��A\�g��b�d�6��
���I��|ز�<Ƥ�_`Ӯ3:D��Ok�D5㵗���-ȃ�����[�lx_�����"5
y̿o�=Ҹ��C�d�?p�gpT���0��x�� 榶^D�V7���	W�d�C��2e����;�[�B
��w0"�=Hz��@9Y�y
�;�dP�ʊ����RJ@1�Fҁ�m�~2GP�u����Ӆ���1�%��I�T[ХF��z}n��47���L�]y@V�@����&g9��\_3�f��4t���?T�$���!ͩ��lT��aWn fM�����3�[K���$�R�m��wPU<���"7ʺ���#�m���ǂ�i; ��'�`��=Nj�+˻�����I/�Ϋ�Am���	*����6,�Ɗ�À�(�K��v��ׅ��#;�����b�Ca=�:�?����6|�i��ȏZ�i;0��O�B�!�u(ᷪZ,�sI��@�KT��MOn�@��i�Y���𐱚�y�,	�B H[x�3Lܸ�t\Q'�:�5�v�c���o��v�����&[ԣ"Dݏ�yZ#�R�=�!�6�l0�KjeH�>>,�!#���B���M�>K*�;�Cݻ8��fG$]��z���W�uG�S�=h�\\Ķ�6��Z.i��y5i���(+��,��v: �S��4|��p�C�����+�FJ�|�*"2�p���+6]|H?u��(w��x�^O���I���I0O�wB����}��+���z�B��\���������@f)2<P=�A��� }`��L��Dxa�o�4��̫����ڵ��z}�?�r���P��7/�X(@N��2��tA�x3���VJ6#�j�:�F��d�4>x1���.�������iv
��#x��)]�.#F��i�n?$�#e�k]u���&���ż�����tN\g)���S�� ;"�Cϡ�}�o��;L���|M9X"e��[��~"���p�^���v����Na��|Y��G��Iq}�53P�D���S��#��&����	8���dK�l����T�P��¥��bӊ�G�{�):u�)b6��Q�Q���ݸ�U̯TN��%�#�2٨)��V#��!-�� ���n�ҧ�X �0��}�ƈ�nϯf��4^���bG�����R>��"�{AN�7�OU�e��Gy2ٻ|��p	���N��Z&%5���Hw+��O�ak�j�|/!������ui�$�\�=d&�l?}��%����� G�-�G;��GI�Q�����`PQ��=� >���e�m�c�W�c��d�p��C�\Ěƨ�Ŏ] i�8�1��zZ3�A�[�8��WY�lqF���藰U:x�~`����4���!�Ū~�zp�"e���D�?_	)G��}�a�t��Ë٨Ha�#W2V�w�f��)Z�7�Fu"���!Σw�:'x��W;V���c%�cvs�	���B��ͿZ��`棱h��;�2�#UƑ�u�B�r=���)�@���lg��駊i(�3�	�a����N�$�
m�A���"�0��"��2��Ti�F���H��s<3�����(k�!�]��w5L��.r��[0H	te��"KRi�o�τZ�w�G�F�3׀D�Ֆ�[s(*�|�;˗9�1}2��3k��-$L�`���::)ғ�������
!��OY�c�ͺ�:���$ݳu��	�S�Mܙ7���!��UƢk
&� �\~��g�/pj��H��n�+��L�{��������	)>lw>/��W�\_p��'�w��?��)(�bmV.&�A�fu�xY���x�C�e��̲�־�$����y������e�en�w"��և�Wp)�˴�}H�?��" o>o�E :e��hm��/�lJ<�R�2�}6��<�H'��x�p���00@����c����s��+�df�R��(n�����ve�QNؚ����3��7�S�!DkX����S*��:��#�%׺�iQ1ض��R�iU�����������ɉ�9i�m8���$=N4T 1���d�ASǴ�b(#�� �/���e��z�8�ח\�����%�f��~��ףR���T�yY���΂��h��>�g�eD�R�[&)�d���F�.w�m�|hō�ejT8�l��U!_���3��Ko)&�c�F��[�υ���o?{~���(�y��q��b�=�a���j��!��cC�ՏVE����ۓ��?$�J�4 *�.6��YD֛��{�DX^��7#��%�� �R㵵f��¢M��jc�zQ�#�Z9��.7�`��zY&|��-�sFQR��l�0�������d�U?�c������ S;���*ޝ7�HU��|C ��X�S�a�.�SS��\/�~�Z/D>���.�s���w-u��s�sӦ S ���ץ�/�*@��1L���I���j0Tf=��Sc<� W��7q�m�00}����?Px�Xε��_�t�>>�%0���,J(n�ݴ��MG0!D�< ��y���nL{�Mu]��6�~�\`�@E�1g��.m����G#��#
�F>|���G�j�-�	��Ղ��*uc�uq�$u�����M����������7���F���g�u>j�Hxs��ܻ�/`\C����Q@ϻk��
r�LDN*��O8���ٺ�;�Q��V�/}���p�����ޗcb��Y��J���~�?0��On��7���<iY��b�L%�Su�9l��tL�$����tor��+ѫ���t�Xmo���z�q�邥��|]����F�G"����{�:�F����:
�+�gX#���V��Fm�.�Y���{L!氶&�i��hbuA\�汾vh�C;E *B0����N�ាYP��`Y�^�(0��\�o���Y�䗉�N.���������������E{���h+M��Z����qGMί�y�b�?��?���2/[@�G�|��t>�M �uAJ'`�B�ǹ�)�2eSʰ�-n,7_9f2�6��7��L������JdM�tc��6'>�����4���~����6�{a����S�7@f
	H$�;򅸐����tVu��e��sURd=��<"l���]�5?rR�Q|v��0z�,Z���qC��0�l����䶃���v���"�6@X�q��sO$G�������4����S���pf��l
�<W�N�T�FW��p��Џ���H%G����HQJxWuv�E���8ѩJ
��Ā`˫�'h<<��Jנ.m���� '�����sH ��eqY��ꛤǿ�L�f� ��(��ׅ#y��dY�ƨg��l?�o;X��xL��NdG���4H�m�8�	�M�n��ؽ��|vs���o\��gy��gI-8�;a�����;��S=!�0�^��ϧ��t㪤��ȨǊ���d|��V��~��^2����ފO�zRD���	����R$:tܩ�W0�����{T���M�O���.ڰp��� �G��`Z�W�Q�Ey�S����<��3�v;�K
�T���"˚�ܑ�W	�^:�����^-��[�����4�Q(}�����Q*� Fo��~4���˷�O�/t�ޙ�C��˫��M�����c�( �9XR�� �Bw�(�BI����<+6�9�d6a���^na2>����0KS�'�(L� �$S �q�d�Cx���ƍ��a��6[h+G��u��qZ����S�L�j���� NH�.�p��i�D��˴���@,&o�fe�~�C�VS��|P���-���ᑗ�!�w��^��	x!����������2�F���ϸ��T2��<JM�;񐜒G������K#�sM-��	�[K#��3�����Y.ic��O��8�5E��H@+o�P
���R�Q"P҇:�8#��sb�ˮV�$��
"��5�7�s����*�Ƽ2�ߩ7��n�e�~�(�m���)o4Vq۬k1��PD3�aZ.��B�/��՗JVs�+�8��p	��{�@���*�`�� /*:k�+�d��ט?�d�Vɸ~:��(y�5'M���*L��z[s��>{��`�^�T\��W��A�p6�h��0pz3OvO�.�A�y��?Q�q��!n:�#�r�!\pDe/�+�f���"�L~
~ k�6g�+���h��d��?�ɤ�9�t{V=��,�[�E@_%
�~Q򳣨]r����&����I=�7Z52�c�[<JŜ'Y�w��B ƃ\۰p 5Rt|�-�st�$8��?��=�Q��<Jc;[��3=MV�(bQ�C1�V� �Yt.r�������g�Ñl�rH�<�҉�.�o��m����*����΀UauZ0��h��B�c!)��V>.K-Ԭ�C*�|Ng8-@پ�!������3��ﻊ�v��s��1�Kx�<�g��Ie#�s�\�����]@��^Z+()�W���$O�~���O�  �f.�?z�2�U�!��_�W(������f'���q�RO4"̸0R�\�4N-�����R���nn�Y�%`�d�;���BOi�+Af�{}n��f|B��va�,+]��X�J�V��7JUZP����'у i'&�_j�d�����PIכ0��d�n3��猻"����{�4YS����F�B��� ��i�YGAT����*`���T���}\�ۅ�&~W���d�A�d��<�������fŅs��5V���,��������;U��?G|q��b�_J�|��4���F��b��Dc�j���?��S�ћ��{�%;�x2�s�t:��Y��v�c�
6� "F����Jۏ��=�Q=SK��~	hS{�����r��k�R�=#Ԃ����X\�*2�=���4�K`��w��e�>�o�g7et�'��R��Lv�F��)�.S��8B�瘔��lXݹ����S�ůՅ���������଄�պKv^TxR{����K� �e_�[2Ht+�U��w}2���i�snj�s����I��\=��@�m}��2�Ԡy����*K�
c�j�����ۉ����\�P�K�t�$�+�Wy��.om2k�]wJ�6��2�%
��7���ޞ8��h���:bx�����\zp5s>��b�W�&� C-� ��J2 %x���lw�v�b�}��.����'�JѵہD��>z�LB��t 9^��;A�	��?�ǳӲ���F�M.zCo�sЪ�A�����L�������*��Q\�;>t1b���M�h�2RB8EOw�0�������V�b���h�$�-�τ5��Q�L2S�V"�b" +���{��"0���N:�������A���ǠjR��k�dg�I!�r|6���!R0#M���3�]=-��AT�,ܢ&�[q��Tp�L�-. j����o�C<՚Z�:��[>�H1J�5���(i����Å�o��g^���ǿ�ی����
��Y#�HU����I�)ςf�e��� 嘀�g )�b6s4%�GK8�����߰�ᜰ)��	���ڄ�2��=��m:����j�������|t?��4塩��M� C�O�$&�G~��bp �mbe�"��w��Y�c��-&e�؆���Y�<���R��}��F��;jd�mꀾ���t��v1:�v$�{P�'�y�b�������x4�C����j�LZa�?�Q��cw1�ր�=
+��')F􀹝VL��6�ОT�.�ui���OҼ�:�X�=�4˱"k���*ikȻ[U���M�����=l��/lQ�'K\K�B��!��l*��ov��;��)ss����=0��:�D�W�szNJ����l'���tP�U=�h:�C�>iЕ���I�(��q�)m���s�u��s�2T�t�W����q.`*.��r���Hsg9�Q�	�e�
������!SYi}v��reO"Y�������)��菶�W�Ù0�ǝ��#}o9�Q���t9�����O�=2�q"��k���{�weE9�Z2�)1�1]8P��a�/NԎ�������	��'"�����B��ћ!P�����t�v�[f)�"��|6��+Si���tN�A�-z3����`uP��;���	=~Vo瞢+�_�u�s(&C�^y�Nd�*��n���J��L�P��(gV��9�׫����S�
�|t	��"̇:xN���@,��{G��8�)���@x����8c�-�q�*�#c5:I���ܣ+CwwlaZ�]�/Gu�	�'�U�=/"BMK��iOb�����*��p�lr\���q�����yZZʣ�J�R�NoSe.}]��֪�N���DV��5~�qvj�딅Нv=�
��)2�aփ*W�uQ3��l�/�C�i�3���3
Gx9ˡW	e�jdR�a���st1�+Þ�DRt����k�(��\�4����Md�O	G����U�ލ��G���_��u(F;3+���Z2YA�;���qK{��Y:`�
���1�J�����]�4PÍ�`�j8,��}����g��v�_ꦔֈ��C���/M��}^�Lp��A�]�9�@�)(���s~K�kI���Wn�&"��II�V��c���N�٧c��Ɍ1��,~1&g������ؚ1���O�<��߅��b�o[Zާ�\���@�9[b���Q(k�r�5���R���`j4�e�ϒ�G�O�|�}A������^�B8�~2&tˆ�A��w�?,C�1P�p[��PɨF�ƙ�_������wy.+TQk�OÆB����6 ;���(�wƬ�.#M���X$|&�*��v $�}���s����ad�ޥ�g�}�[<�_�=�g�f�?'�P2�N-�X���e�[�5��'81 ��e�[y,s��"�Z=���s>�7��%2���Y4.���ټ��;�5S6�Z���	������3������N<��g��e9�/�l��ZLk��A�!����N�ɀf����]C��"�1�C�2ґ��\'�i
WY{�!��WZ��nťs�K��t����ՅV3��������ƿ*e��{����Wk��
n��tw��cZ�#TV�b��.��p���
q*<!������ux2
�j�yC@)�g��d�E���	�K9�O�2��b��>)���H��EDW��5�>hl�o�Qd��P@C ��M������4���"qq �y&	�
�5)�ݪ���S�k,yI*g����ކh;�lh̊ͣ��n\��ȳ��,���+��L����ZUA����!`��'���B�s8��t��Εº�I�2���)&W#��z��i;��`(�|�Mf,�`L��ϢIF)�}������aˁR �oeu�	b��A �a7�rʁ��Q�i�<z�޷��qUG��O���wn�#��4��>�ߴ�x��)q��K�aߺܾ/�f)�1��B�*u���ń��J�5Ⱥe�fEE�lOR�3AJ�F0��MX�;��e>�l�/Y*8���Mݯk���t[���{��kᵧ���'�M^�щ����kPJ^�%�L�2��x\eu���d�,�
�W�3�V�J�#�l[z�\�����᫂��oʞ�ʞ�2��u�^3���j��T��/�?���RY���� ���]���:~��y*���a�"��j�]U!�i�p��n`��q;�	IQM/yF�_�O4��⃷�� �"��c�5�Y�v�������if3��4���:���Q<e������9Y��(@o�l��y�3�D�>�p\{����7�j`8~����jN��$Q��}C`J��\M͞�\<�ʰ_6	��B��%�� M�&�d�2��N�D�{��#�
q]An�
��#!:)�@g�H"���ĂGz���o��p)�0�p���M@GfS�%:S��HؕUsBDI1� ��&,H�W'S猶��;I�0U�t���U���5'ϭ`��J��Aչ��G�=������S�
J��6MT���(�כ�x!;"۶��Iz��.S(��(�}��F���6�'l=����K�G}�i
�Y>�O��M��sb�1����d��^U���֢i�\@��S��K$ʍBma:A[����e/%��ᓥ��!���K��'�8G'���
j��㧍vu����,N4?��{;֝9T�.nd7ë�ƪ7gխ�vlb����ug����c�$r�'gY2�!=RQ������]�
+��^fLh�u-���1�B_S��ɫ�R!��~���0��M�:��@:g\�Id��-^L/WGF��7Kӟ�	�.�����/�B�Ԁ�mܫ��])dӗa˻J� t�0�@�wȹpc�iQ5�5j(�Ob��T��3��̨Zd�I΁W�d�X����lP��M��^
�����s���Z��*�EѼ�*]���� �am5{6�ʧ���Jϼ����&�B�ۤ��CeHT�=eɐͮ���^�7QZ�#5��XO�h �_���Ӆ��=ʓH�]�*��t��v��g������͠o~��Ʋn�Oll���ǌ%z�4��;�r�Մ�$���g,D�N}1K�������F����:��rq�(=�BE�2z1+��@R.Qژ]7�¤��XW��bS�lv���|+��y�ӂl������U�S|�_X��*��{�aX�2a0b��?x�qG���N��>�����4@���7�e�222��	���4+���`�h5|�	�����\�
F�)/[a?.�P͵q���(�V�7�|������i~��8�s�}^���nG�\���M�)Q�hZ9�[��
}l����c+WnJc��cDH��E`}������-B#<���Wp@������F��7� p,���x�QB[��!S���D9E�2A�&��Y�!X^��%�%�o�& ��Xcu����L���c��d�Nhi����Flyw���'j���+��H�(^ʷ�F0Ӂ��cU�t�5dy�wI��� ]~}%c���d��Z�u�Ț��uځ�4�h��phV^݁�����L.�K�V �|�@':�'2jK����3��ܞ섺�y���e=U�zf����4�P���f4���qq�ԭ���!�(��,�`���4�Q�yv��NS�5����L�ye4V�D�eEfN1�pnt�2��d���e����B4Q�0�7B��_E�
��Q�Ҵ�ڢ���W2Ȱ<*�E|�8�;�G%>�R'0���t�yrx�+�����.�/�J\A�����zv%�mJn��\� (�D�5O3ʸ��</Z�1�Z�.�-���F�9��wA�R��l��t;4�z/;����^���x��;+O%����K�Ϗd�x3�X��TH�u�������G&�eo�TI�e�*�"K�X�"��.h蹌i��r�5]�U74a��8o0BǱ��ɿ�[a��ƅ���'sFd�Y���+9(���wNMe3�u�՚��dQ�fc{��,���Cx�p�x@q<m�ډ��KJ��7��x��~�|�X%���4�i$����&���tUw��|'�\t���}"v�F]�0͌�gr�� �Ɨ�5�d�J"ɲpx֯D8[�8Q��>��cLw<�_��&�����x�Ǖm�A��)Bf��ٸ_�P!.	������ż��e���������QS,��E�#�+j��&�w��i<O�{��H���5[���QF,%qm� �r�8Q�*��2��k�#fZdp��2Pn��z�&7�Ɂ��%�}*�Mݛ6��z��MJL�qN�������i��Q����`���'fd�*$B�o�ԍQ���e���7G�7� ��T �.���-������h�d,g
E� ����7�Y�� ,�_�ҊU~l�v��^�h:ϰQ�Z��e�������-U�+BV��Xi��Y! Dҙ[���5� .\��;F�v�O��oV�i(��$��:c�x�?T̫j��G� /��dD"q�H4K�w,7+�Z�{,E���Ic��`��y���Y%�GN�����:��n���G3�)��#�m�� �e�[���UN��͊'C��Q�zug�D�O8����+������n�;��ٕѺ��pލ�B��6�@T[��h��6:xS>D�c��x��z�3D��+�j"�b)�Qj����ƪ ���(OpMp�q"���8�a��������s�@�e�fvy�;�U�� ϙ�	)���ѾK��P�ml^�3��s˴Z���#W�ܙ�b��G�p�%i�|	6�)��:��+�g	gp���ϔ�MW⥜��{�����䇢QS$�0��i�}�L>��g��]m1/��X���lps�u���n#���Y_��%�ߛJ� ��a���K��vU4̜ƅ�T�-S���G	7i�M�ZX}�hʨ�BU=ܣ�ͼ��~<Vu�Ԡ.-�e�`Wת��^U�Q�>�r����iH���U�h�
�=V���,�_h���-b�"z���)&��w�����`$��:����B���ͪ�0���<{��5�~gq2�8�2LA���y}�!c�o5z�c���*H1.uҸ���j���:�W�[�Lj_���)������l')�9���~�mp�rp>�.i�۽�k�S���/'��5�:���N�^��u|��V������[z�}4a��w�{��y��L�o�v�U�N����꼺����n�t'�\�����~����3RB�i��I.Z��������3��A��y)~i����b*1 k��W�4�*�jW��yf�*�X4����ܱ����K��,,���L���W�Z��c���FF��������ö|�$6hFJh	�ۮ�m9>�q����^v��~�K�D�s�e� |����+Ϳg����=/,A:ruǼiA�#�jRm�9���j_��GW� �?��-Adq@`#�M�;󻫓0���cY�*��mb(�d^h���c\y� ��e%а��yRur���J�������I�պ)���T@�'rx�����V&�'B�b9�7�l&��'�΁�*��,�i�ϴ&�%U�C�ծ�VR�[4��n�.mL��KYAE��A|��}��OO))����a�x�[z�=p��<�jtw���UVDS���y!\�*n�ӓD$b6Q=�X^� �	���9fD��5X�<:��R�Pn�������)d��G/1�ip��
��T�ܓ�C�7��Y��؊����W������@����)G6R�>��AՑ�<���M�ϞݼE����i����q%���.������.:��_֡�V��s�>ʚ�["�ĺ"��%�pɺ�~�@-�Ur	[�<_���,m�#�4,�:Q���]S��n�T=�t=C��*��6p�|˭��Dp�;.令j��,`5�l0t��G��G$�i�L��N7L����.n�,���Z16��;J��!f
���ܟ��J���er�^�7��d@�J{X,�����ź���<O-���%M����C��09
�W�0�~n�2��{\y�B�2.z�t��I/3��(Bȹ�����7��`{��Ů�m�I���l�8=����V��!�QE/�L@�Ū�`�Բ(�p�{iG`̇����+q:Ս�XA�fơWВ��6l�гxF"K��2&W��f�йܯ9$�7f[_CEҔa��?�<]Ͻ�� �y�G���Y].P��8V�^h��]�<��5���D��ySֵ9B��>'�Q$�Я@T���zv�8s.�V�̃���t�B��!S��iv�`�M�q+�¾8��޲�!hl�r�=��-o���G��z3�ml�,4Gkm�|�D-o/��$9Ob�[����	��b����*	��Qў��T���C4�@������"o�6Y��}��}O�6�~xШ7Ky��sv19��@�v���,_Ԗg���.���'E8ko�gB�`G̹9O�>�q��n�5S�u�h���7.X��j�QR.癅4l�R�!���y���v���ح0�$��"����WH�5��1I��7�/Z��C@%ٕ	a�Y��#��.}'u�bC�HF�H�ћ:��{�D���ѽ2������)�&[|Q$p4�,���v������n���a�Sz�U/�+���8/h[
��_Pڄ�f�e`޲"/����)��N2O���'6��3�1d��R|.3��f  ���U�1��R<s�s?�s-�4�R�vN#���+���[8{�l��c�!L���(-�F��4�l�0�H�ql{`�o��4�댟F�!s,�"�'��T���0V�=���h����Ƒ�H���vZ��([���#�^��7�[�P/BL6�4�'_t�৮0��ˠ�j�}��v_Q���谭�/{���q�HCƻz2���u��#oV�����Q�[�e<�3U14��t&�'�@�V�z�`X���y+�q�b��j"uP9q�{r�@S7}�U|=�Y��L_�b/�ݼy�J,#�����\�A�VI���o�Az�U;?ؕD��a˒��
ikփ�G��
�G�z��p0��uz��,���e ����9�ᘱ��n݁�_���%�:�6�'�G��v�tc;����о�3W�'k��S�f��M��.�	E���XS�� Llf��kZ�`��u?�HtcF>��sP���
2�in͍u'|T�U�mk�R~~(��rR�N[����g���<���cɚ�N2�n%�*�O?5��A�����{�Ò��dx,l!'�.b�8�ib���)��7�G}���C�aR�G6�8B\_���i��ѓ�;ގ�C\�Ó�⅋�Yo�6�z�!���w��5�
��N՗�c������Q�������闵NѶx-/z)\h^|�V}�cw,+Y�Vw���
>9b�\G�>�Jߢp�Wd_v[G(���/���J�S�O+ԝ*"��x�Ih	nyt��?P	�P~���hx�ε�]���d��|ɯ���?a2f�-����h�6��#���A}5Yk�q��{�ЈH/�^q�?C{�8�L�=�w�5ž���p�d��2޺�YF@+u��V��?@~"�S��%A��
y��|��w{�m-�c����Hks�o~�|
�:�ߥ�-���vp�2V��a������o�x(�{8jD]��"h䴁�XH����ڹc��-��U �<q�%��ҫOI5�1�~�� :�fl'��a.�R`A�k�!Ї���=�u
$�����;r~�������_}�� SH�[��
��K埼RQ�8Co �HO(g<	
�㷎��AN4޲J�����*��X�k&{)k�"HojY8?sr*�D�NEs� h.��
��.�a1O�2������wo��T|���ULg�bd�	{ЪI��넝���gr?�/L�����[@�nCmw���!�v�^��F�` ֈ�Y���ʡ���F�]9g}�
J��M�q�~�|������[�_F+�gV�@A**l��/U���fCͥ�ɯ蘴��Y�4�N��ř�7�'���[����P"$���O���8z.<R2h1�۪���:��L����=��Ym�CY�u#�s+���Xg^�	pY��)7����w�ۊc����Obd� ���u��nȚ5����d!��)�,��*���e��ɐ@h�!K�~E��q��7ׄ����tldʿ���Y,%��\YvG�� �2�!�
$�d��o�o��I�������f3���a�}Ep�s7	"7I"d�3��0Ck��0Tɞ'6�&BE/u�`��|�6�!W��B{7C}+g�����k��k�q�Ǐe�o�k-��(�	��0|߼�h@3�l5��{ŗ��W�kOIv�v՜�$��.����|�ʉ�� �eJ��i��]�O2۱�o��[��]�q7EV�EZ�O��%E6�yw���5=�2û��!�l�z��rc��9o��"�#Y	E"��|� ����;�Q��>B�쫓|G/�.
O�' ��Th����C��;%��/�<<�#����ؐ	�J�2d�8J���UD��۽�.����l�����_KU��2d%׵��w���Q�Ng7�H| 0���.�eי�E�� у,�����s,2�!���)���xbm������1�1BJ�.����P����1w�`OD
a�*�UI�j%���}��/n 3GI)n�L��.(�|�!o!#�^a�4@�c�K�'v}MHE�7|b�4^�okӧIC&K>t"�ۢM`&�f�Hq�BSFE����"�yۏ�����uv��IHG �]*N�z�S���`WKq��KB1�"�g�+��*8�	�0�w�7X�]lgmO���0 ��H�������=s����2�bK��}B��E��缣���,	��D���I]<�X��;�w�%�����D9�DW����Od�рU#����fJ���^�����r���9�������w9݊����ޫ� :=s���f�{hܺ:(e�;�Ȱ�x���%�t���z�A�3�O���AP��[+/�1��������V�F��MA ��;����X���"?��D׀3Տ��{z�o��RUkP�����NZ���A�'��}��W,��A<^��jT�5b'���5
��e0rh�o��C
�N��eN�T��3��{U���q�޹��e.���(mi����w6�^�8r���N`����na���59o#ې.��ܦJ)��
�����NB�f��P�3'$�m���n��n�2��YQ��/*����Hl��F��=�ێ�$+ �;��JBx"�F�bR��� #}
��7�j�Q��+/��"�!�%l�P��|o1P�]��ޅ��W�VM�*���r+N��]�M�8���4�+�.$���ޞ3.��|���ݎ���l)�D����Z��TX��� 7z71�S�I�Nr,
oU#=#t�S�~o��՚����N�ϏFZ��t�\�Ǘ���$��%uYaU�K��t�d+�]ơ�q�63����}$��v��c�x��GLR����]��@^�"N<�ۛ�Sh���Xͥ�W���y��`���=��z*i~�z^Ƀ�`�`��*�H(c���K�2ń[vᅧn��ƙ�F���-�̉��@��c����Ja�y��P�J�;�Ǫ�43�>�v�A���2�%!¢�.������S�
d�<��ў���0w̍�|m7P��냁,�}rF��u��0\K�.��WI�X�O�֪��a�,ͼ	�nVO�#�A1?�TπX3���=�r��U���h�7�=J��ؐIݪS	o��R_e_6�ćܓ�?�D��LaF�/�nZj'�4�Q,��_�8_B��aQ���X�ːB_�8w���)���;���~����R�J�apny��{���&���R_r_��o�T�t��;�eF�(M-�����):������$JЇy�z[�8���X����QH�:�S;A{s��aRKR����B�0�����
~�.k�@���!m����-�!8��������P�]�e�fSz#\>AH<���;[�|�G��kibՒ+�`@��W������̧q����2�W�x�c�Q�;?��:u��Ll���x�O�U�KzF�*#� ʃ�X��@Q�IjA����/��gI9����cD�ģq�</Q���x#�h潤>7h�~ڢ�Rղ��Ц��i!��2Lˉ_Ju���n��V��pM�A$F��!�#�-/ꑊ!�Y|�sy���[�I���)�1)��-#}3�u���(8!R��V]�����l���纋����*��'�|����R-G)@ؗ�������h�[����[w<f��ts�H�#
��\q�gN��E�x�e��&txa�c���M椭���i���� Մ��� ���sq*�@+z#�>Z0 ��G7��,�S�x��w�̚ݺ���l�Gt;W!���Д����w�OIČ͡��kW��ݺ�zL2/�A��沜�(w�.���h�ӫ�e�R�c\�V��c�O��AWa���}f��[I��𤿐/,z�1r�� |ij�8�m/��`?�77�8F�N�8$k!�&a),���0Ƃ���@���ʜU��� R�vP��S&l7�~�.�5�!h��͖�C(z�O@H�ǵ�2��jG9�-��lzź{^��ߚe�[���Xս��Y�,���K������&���sO���s�ˣ� q�\�،R���}����2�����{�V��� /��~tg��iyf��ޤ٥���@�:O脑�x�+�)x�((o��+y�,cvm+��V�ǡX�c��H���t��7_�.��20�0ZO�d E)}�U&J��-/��A�.��@a�H�#��eW�x�zLw7���Oʷ�<��+�	�X��5��t���ve%ch|[5v�^N�WN�����\'<���g��MuI?H!� #��>�1B�7J�(�<�^_%vЇb5�� 0V���[�G��f��2�Sq��������`��8��
�E�����]��$�1tw�7���8�|�f�]�F :>�(��/s����WZ��L=������p�!Y�t���#>�@��� �j� �\=[ߤ{	/D=ѱ�Z6�K�6�oזL�7�i%$��_�%1�:��V3/T�Sl�K�(��W���tG�K����Bt�w�b��~rK�[��~�b7M��xg4����q�9.�O��$��F��A������1iR�R^.��"�ж�����{?-����t<s�OuI�kN��7FQ���4M��Kfal�v�rPAct#��t��H�"x�񕭶F���ܰ}?o4 �E�3qd\*�櫽䟂yqТ9I9��'`��C����,g>A�J6#ogs��"]_A �^�M�v�Pfx���D�Q�Za�f݊�&��KO�\[�H%BS�GhnAV1��|�@�oR?*��B�h��PI��u�r{a;�?��SWy�<�P���\"ȗ�r-Qi�k����ܡ5-���2S�T��	�G�	�]�Q���$�� ڻ��r�іo0�Xa�G��:,��s�
������p�)���<���[_��7���:� �
��+}�B*)�1������ɐA�%��x�^���8������*�bJn�G����4侙���1_�PD�u��~
q*ay2���Ԫ��IfZ�䃹�ÄI�j�Eh�FЭ}[F2��h�beP��cr��S���5^��@����٥��_��� 7�X�����[��i����D!�#� �z��i �Rc�  �H�04T�^����峋�Q6��Rz��k�v��T�V��e�f"�o��Ḧ#���iWi'��)"	Ӂҵ��
T�'	E
����7�,hQ����J�$��l-��O��Tp���1���}�����q�?��r�G��Gl��gI��ݑzJ��=�jZ�,�-~~���Ch��Q���to���s�f'ۯ�'� ='b*��1���9�4���t�w^_g���d����������!:���^�N9���u&�==��$Ԇc䞮 ����oJ�J2��c,�?��ަ���vR�̚�3��tΩFZdQϋz�<Rj�X*�ܘ�!b��@M�!����� '�y�4��(�5pF�-b�6X�0s�@\��L;���˃Q>e(��3�맃̚t9�p#,b�,9�:�?a���T�|����0�{��q�����=ƍ�E+FS�gk�lvR���� EJ�b|�Y���
�����b5�%z�o�����`7��b(�N�7�4�@8��j�~��8C0�ԧ�v+B���z������{R/���M*=� �R�w�xP�ʼ@\=�<-��Ѻ�c{���?~�l!����&�ڇr���K���}�����O���7��������[Q�l����u?�$�L
xb�M�����O�k��t��f ���W���G_F@�5���x��=e.���Vp���c���2j��A�w���[��ی,���Z�����$is��<�A\܈��9<���)�w{ E ��1f�W��C�~yf�77���Z�k4��Y}(z�#O��A�ɘ�9&�����&E��$q1�1D��5 ���:1Q�T�b�u�c�G2L�ww�a8W Ȱp,D�)��P ?u�"��ZuÈ$�p,z@y>�R��_W� )�*@G#KL�@^�QI[�L��['�������]F[���薹��-�oZ/�(��}?^�Ș�JAm��b�̳#͍���f x����%�/���������n�9�R$��G�W�7���A��o���a��(b���v�|Db���[���B�˛P}���n���>2��m
R�&���$��D����aF�6�o�,��4��뺅���d
�y��q����z`B�N�o[.Y��j�%l�$Cv��A\��kV����U�����n�x���yb0z��`�'���,�]���p��mo��S����D7�\,��=�m�H�,�v���Go�CݹUV��n���F�p@W.�u�I���cR�QR*yhq�y��V��dg�<��ݍE�I���i�	'��vnYӲ��\� ��˥g��v86u���? p]�.r��	�D����2)"e�p���߇Ǵ�j�MJ����ꐞ�QG��Z�x���=�k�>|�m��E�J����(�굁G�]�U���:1�cW�Ksε�۔T�Tx�;���"��+�I5.2�,��	����p/�%Wߌ���s;��
�㋮W<_UW���'{;�i�}���NdY��
P�jL�KG����+k���w���Ȭ7�l��� T�Y��AsU�j�c��l��?����OԊw����w�����Î�qX���׮�9*O�n����Ԛ��#&�Ov�
e"d%\�<�C3�����W:p]�Kg?�C�������
$�i�ð���.����֮x���%כ1��yQ$�[xtג�a`)�d�w�� ƽ�`wv,���*�~��K��y�w`�X�s��ej�m��D�7�-��~kQeQ8t�>�<b~%R�;F=�<_%�T�عI��������eh��^�4���_&EʲS���Y�R9}j�o�H�킐�� �D{����;"�Esd'�I�����P��Z���ݢ���E�-o�m� "��>��������D?�W��K�i�c|<_N/��5����'��hm�����(R���Eى��˻��k�G��6�\���X�|��Q�fճHn>�6��T��ė��O��n�2S�{e!�,���$�ZHגS��������ޓ^����ʤ	$��d.��}+���#>�ssD�� =��ꔺ��9�N.�:�/�p��/�kW����]Z����Kxx,P&��E�gtYT �?s�;>�YW����]�� ^�ҥ[�F̓	 ����V��>6�a����;x��������N��sT�ˤK�^�qem2�3�Q]@m.���j��܉&M�
�_��̺!((M>�i6m�G�����n;�S�d�#[q��՟�/_�w��J�}��uh��2b��jѡkLڻt���u}���p�;ݰ�x���M��G����E<97���m���,�� !r�J6ƺu���+��>Xt� ��S���9}��h�Ʒ��$%B=�xgnmZD��Dχâ�g�Z8��Q+���Lں�T���f��4�n1�$_���>��45����Z������7̜h�,.�{n�<M��y9��\Z*����8�)Ev������0)�Ө#�`��s���Td�ދ�5ƹ�J��ߏN@��������`c"�O��X�Ȩ
¨S��B�-�\�)uݨZ�{s~0���<Z�d��&��~�%�h2&�@(qOn�(]\ �Ă��MA܅�����r��T��γ�R�7��-�[z�,Wr]���+SnV`nG��1$"{�H8���ɀ��-�n�r�uS=d�u9�l�gO�ep��w�|T�.IBT*��1� �jP���� ҿf20!�f���ܔE����y1�r���m5��Vbji�A�4�\t�1G*3��� 77<,��������j�ܭ�J������/�Ck�oZGWVlO�%}C�d��=�==�K�g��F}Ł����!��:qC����J�Ya��s�9��a���ރ���D��eQIu>�!��A��7F�	Ft������{�`rU,Ñ���������T���L�Eԟ��<�r��/ߕ�ڑT
��X ��2��y=�rSM{�~�j��6����b?}���֊��	�/J	�]Z Î���)B�J�k�n�r���o�N�$v9��#4�~H��5�������[0�C�sh@���q��gG��.�%՝���K .2|V��V�_�u@�D���\��Y��ϜV3*=H0�����7/�es&f`)��EZ�9T;�p��q��-�g�� ��gf��w8T��H�/�o�92�	LV7��W����dcZよN.уg\;5��9V���)$�R�a�>�"��/�KQ�(���WY׺�4
D�|������{��(@{�!�ͣ��wq�����Et�~�˦kъ���UHì��+��TM���o�q./�-3>�$�">|���0�+����d�`S �0�M�⽨���'-�q�2t>i����wW᚞c�Ql��
�c�C�:�����ve�����-������ �Qja߈*��y�#%>1a�J��L�=�H���\�BM��o8�۟Q��4���D������Qt�2g/2��Śq�H�Ķc�4<�F�X���ڒ�jW��e1���h�YȬ�����\!.���Q��!�K�we�	���Ol���^nO��e/Hb�3�K���g��%Z�߁J�e��ʤJ�Rw�K�r�P	�,A�ʱf��/m~f� Iɭ�>��e �l�*E�3�t4�~�Qϧѳ�ib�K������Yy�6�^@͙k�I�7DBAoS��f�r��*ꡑ���?��6�ʁ����K���&ϸL�K��i@���#�gT�ݕ1����aX�_��k*s���Jtm��q	}U�,-PT���-T�J.���������MLJ�-w������t�������ÆZmv������>a�xt",�BYQ�;�ջ*�Ů�7�(�$�e}ϴ��4Y��(Ω�mv�C��ƙ��q'�P4q�\��W,�4�f��Z�C��	�:�������b!���Dal刔sa���$�sN.P���z���,~��'���[fm���'�R�*Ŷ�t�kb����+�<ve���n�"g�{e�o�q��乯8@l��p� �,:ϳqǑ�*����6Q6�A*��ZC��&�u�z�m�z>�=�=f��]����8�]���~��20�#\�h������ПDRH��)(���<z�D�Fި��*�-z��Ҙ!����$E}�ݕ,;�W�vp$-������{�|[U�Qy)gډ�	#h;�sm��X�&�]�Yǣ��wD]�_^ݜ����`|p��2�X"O��eAٽ�҅�P���qq� ՠ���u4Pɽ�f�c�5�������Ip�|��d+��y%������C+U֯sA�z:ae³�w����y�jA�ȟYq�f[z�x�k�W�oN>aud</��7�Zt�鼊զz��I�A�-}��[����Y܁��\�`� �Zk��eW��YZԑ� ���MO�!�����ءx/T��������~Ed�t�zK��AN�Z*�dG��Rz���]&d��D�.��|8B�������UEP�_�	^�`s��j5��+�vU��קsV�5f���^$
�_�H��<�,��r��&:_A��9 b�V�6�V�����4� ~�T�mb�#cS}��S0��L6*�u����j��/��׌�ٰI?��-� (�gJ&,����؍?f�ޅ^������_ �c/]/gL�ˤ%埛�i�h�G�
��%��|��|�wb�*�i���ڣ��	N8̑��q�~+V�����|�U��DJ��B�
4������uSM��kq�r��
�gѱ�Jl�&*�-�E�����!*�du	rN%|�3E�`�7R�d:B�������V�Ĺ��wߗJ�r��������8^�G	h�T����&a[$��d.MV�&ЁIV-s_�o'���2���$��y�����1γ����P�� XpV7��q���lb��L��*�<��[��Rxҋ��Y��8�0�|�w�IߓW#�Ǯc�/--�]$��s�d:eE��N����Z�5�NJ|���s��V�Ц���u�䋫k��(��V�_��ϣ��?_H��(��姦�OH����]�����X16�;L0���|(H�Б��H�2�\='��؛-�^��l�XT]W�7� !��i(�N�j��;3�.d�����RE�b	1�NFky��M����\�Hҧ�R�N"���}Z��G��ӣ1��"�^V\�����S�d	���G'�/��B�BV4B�E�x�W5l�M�#L�v�sag��͋L�{��[e,����x@�V��F�j3��;ϓ�������Pb/�4��1zgf�e���!�[�n�T����a� ���0B�#B�Q4=�e'أj�9���?"@���Ұ��ƌ��W�� 2���"�#6���%*��D����lE�̺��G�0l'{=�� ��eS1�;]]�����;����o~�k�IpT��i�U5B��[�J��i�.����P���ɕļ�+��Q��>�S���Ȳ�L�S�d�FfQD�Cβ���_�2�{5uh]l���w�7�`]!SG�k�n1�_S�'�e�̷l��/�0ǿg���P,i*SJ�yv��jp���փ,�6+�:Z������ya8XOP�T�o�o+J#y�0uh"�G�(P�����Ul$~W`z� ��`��L2j�m�fWxv�d\��1D2��!=���L��� ��a�a��
65�e{(�u!qbم+Tp��FP��}��.w�:��tP묻Tl
�;��m��Qv3�y��`$+%�7�>6�X:�hP�Ħ@�7��K��������FE�L]&�'��e��y�F>#=)$�ebZ�g|�`RA�
#l\L�E�jȩp�~�������ᦆ[�W�9��JJE2�Dk��k��A����9D� ��)���nA����í�����QD��5>|̐pfqa@Q߶6N�3w	�b���-�]:K�\EI���P�w�s���ۍ���e=+ʣm�Ih�
c�
+1ox���H-:�+TϢ�cΏ�-Z�\؍�9�8詎$�B	�$���ʄ�������ySv��Y1� �Ttg���m�B�!jg�/�����M�E�09�n�7p֔*��$�C9�m���W>RmF�&[��l��=���OS5�e[-^�λ��n���>�
��^n'�0���ˊm:L�ah��w����cލ���>�.��jN�S���ɬ������.���ֲ������nh�eN���XN����(S�x`�N>`�C�˕D��GR[-3c|�M��D	��l?i�(�������"�WJ<`>������K��˱���9�w׽"���r[�$�XW�Y~��2��И!�_ds4�ѧ
�PE]��f����Wl�i�j���*�N�����5"�J.1?xaRJ9��ဘ��d�wG"��p�(n��e?ՙ�s�l4M!�;����[�`����H��[���`�,�\��U��;_���V��tD����2�)O;ק�n&F��3mRZ�y��x���"�8�f�X7�5 �R��ǯc2W(��]7@��ׅ��0hK�FԳ�o��f�z�ǐɹw�%����>-���5c��Ѕ���1KSF�E��-u�QZW��Q	zf�|� [_�4Ǒ�j�졸ͭ���ïԺ��4�eփUk�������O����Ѝ���m�k�=� �)��E�|+�u��ծ�l�kR1��(�;a����ƃ9U��@�ԧm��!��@��t�"R�T@���;1j�E�!89��U��P4>��{�RR��-㞶?�Jn���11g����8���  ?6�E�`,��{�%����7��^3!�6�Ze吀�Ĉ���>�ܨ!�8�D�9�%F�&ˁ�+L�jgI\���3�D���NWG�2�V�1�_�I����4����.n.�֝���0��S��_(�U� ��/���;���un��(>Z�����͏���g/���z"&���q��Z��v�	S`�o��M�^���%kGPƾv�j������o����볾�߳-���}�u�ۻ͐�h?�;�MB�J�A!l%�\÷�H`�����A+h:TM�Er�f��񱖦��U����W� �xإt��c�8����qÀ���wr��Z�k��or�	2�6I�u�p̭�"��:����a�����~+Q�it��E�ҷ�EWW9�h�'�3�Z����r��ִKѦ��%�E�e�Q�Q��3��[p��`,�9�;6@�5/�&醃Z�4`t��q�H�hr�z��+�h���t��(<"ь�9��]�Q�^��~�tJ��p�d2��E��w#
�B�V���(l��:�
�Ou�Ì&�}:���i��8���7��'��A��?@E��g�%���I�w��4�8��]q���] �6q�]�ݯ�x�5Q%m��0�'fh+���=��h�Rt�`=��oE��x`y��'��"�F %'H1�b�mׅ�U��8K��W����ݮ�F���,<���Dʙû�]��<9)����)h���sKu������5W�~�ң��Je� V,���7�g\7P�@�9sGn)!2e��P�+b<3��0����*Gq�a���c2=ޟ)���	��3`
�a���籤�t)M,��� i)n�
����d�	2vt��rg��b$�8��5�Aٷ�ȢX6ye�C���_�(M�@��_	Ds�W g�
���̊c;\!x�)��PC�����O��Zѓ��X�W+��Ev6��(�"];�!���)x��|8�Ԓ��z��ˏ��~�+_�0�廆�#~��������G�Vf��]ee�w2�;������L�x�+d֯�1���P��r]�R���͛H0�7��<��? ���lǆqR�/�_�����/�D;[��+}ذ$�i6߷���ώG�s	�zT����Do��HECS�x@��z~lJ��8Y����4X�� Nu�o�sX���i	�4�1��Y_Mg�6t�b��}UZ��3�^��K�� ��]����#�N1�`(�B2�{�Il�r�]^/�P�r�E� �ʸ�z��5"/���1�$e�:����f
���yL�^����\c��6 �t��3��os��c��4s�0&q�p��P�]c]T�ǎ����Ð$xB�n���|8U%)Z���S�L%.�h�!�|�� �?��ΘL��9��~���P��V�N]}�SkOY]�0[BT�]
�0��y�!�t ����ΰTއ]�r&;�m(4���vO�q���XQ�Ǟ�1l�ר��MF+�!�+r��I����)�|���g��S��"�ΘU�x��G�e[�l}�E�hӡ���q�d�?�h���MU����f|eC�݀<(�t�Xx.}�D��D	�����U��\A��`�b�S^�B��g�S���ܴ�PN�f�ul���O�� �Ѣ\F��0`��{�X�A����$k��� ��>q�m��K��?�<�%�
�(�ΗV����7���~�I77�%�К���������S8���w�S�Ƹ���H�L+���!HlA�1v73�)�累Lw���**zp V�����~�
Ų_�d�@��t�0���2%�����'k'�B�T�x_cL����g�>��Tw�71�2���Dy8I���{p�V�wS0sW�HI�vfQ*@Cr��"}��*�^���Cnլo{J��A#j,��tq�}'6�,��ѻGDb�ؖ�B���9s��Wn����z���07vx�$V��7���Y��"`��J���r^o_���M��� Q��v��>�	M�1�
��]��ZSɔ�����n�H��17�����t"��x�S��\nR�o_��\m�&�t9Q9[<�ў�!&Bn11$Zj'��g2�Բdd�L�g�#��^�$7�R������]�� n.����R�����Q��_Ql�4
LU��D@�C����Nm���ёv��N�YV�?� B�m�	�l�E�Q#�x�N�չ9g�����w�����SfǲA�^Nx8>V�{�$��                                                                                                                                                                                                                                                                �.e�K�ze��ӥ!��Qe#������f������#�k����⌴�e0�|ۑ�;�1/1/�<i<P�w1�yY�&I*C�]emr4E�J��S%c��O'�|���	bq�,-p�-{ �ݗI{�?a���t�4�c3:^bF`�1���鼱���� ٩j��Vϣy��v�d0��7.w�S�D���Wl�	u�O����H����z        ��    �g�    7(U��������Պc���   �u�46�m,�S    �A�U�V���	   3��      ��N�1���B*��a�Q            wh� �0�q#:^��Dx�$�J�*6Nm: ��,    ������	n���v��쫨���    �A�    K�\                _���    	           g��   �@<p���g   zI��w6\���]           &j��f�B�   �$�    ���    �D2   �U4�J�:B0��   �1�bxe��        SZW�39J'   @(� �L�               Iڴ   �b�    )�~�       �N���t�          �/e�           �o��    �Y��(��&       x6��Y����L�    ΀����    �i)�z�ӷH�k#�N$��:�UZi     �{��$��*    ���f��f��        ���c}�I    ����    u�0�    �|��h=����m}K��q��`    �YOƦP�Z���:    ԍH8_���wy��    �eh�,LΝ9�7rIt/%O    	   h�j�            6�9��`4          w��G5ۙ�=�~    �n~E�ï�Pǋk�J                  �gΟ����i@    U      �d��R��Ox�v 7�!Kx=c�7w����d0�bs��    "A�s�!�0=�����y���	   ���Zjt�        )F���(    爓��'�?                h�[      0�e9s��        �=�I    �>��)M�;"b�    �҂�KU            F���m
+�WĞ�R    Ɨ�@�냔ci�D    �q�u     a�    0p/�    E�    �H�����   �%��    m,$.Ԗw�Ց�<IH1A;K            ;�|�   ��|�    _,mz�@��                   ���h:�Rյ�B�7*޳��=0    {=             ���      �"&B#���   PGU�-yح$�м��Qe�U   h�^    F�bv�A�        �X5�;����   q`T�                  ��   F��HNg�    �}i   ��:�⹒t   m��    �)        �R�    ���t$j	��{������H��o��,-    z5O        w���xoH���g6�W�a��[�/�[�   �tˠ   i�,㿿C               ����    �A��L��            L��B+�        �--��
        
   ��DQ�B    �|>���l�G�          ,$�X    �w�
       S���� v��=;�C	Bat�ֿ   ɣ8N1�GP���DT�PY���WV�4f��K��~r��,���z]�5�f�~gs�Q���
          �`��       �,��}�{�w���n��      u�H��\���K;�lw�T���L�B�FS�          	���   �{����    +����           6�v$    �q4<        �CH�    孨�>�Re#����   ������J�w��8g>�Gá4u    7w\�   Kʞ�               i��       
      )w*m���yRb�N����x�U    �뱵    4�%��NK ���-            ��"Z~c    o��	   ;�.�   &�G���'l    C� b       ��u|_�m             �[M�P?�[Y7kr����!4eq   ��|p                       �0~ժ劯�'W���    J��        ~�Q�          ^	?��icb��%~Z��   �&t����    Ў:��ɛ� 3rZ��ـ�g(                       
EO                   !"    ���*��6]��f+        �P��            ���k,�&O�A            �("G+_ �2>��Y��    �Y     ,�Y��0}�       �    �Q �|Pt	                ��-           �N�       	��   /��u㸠                �t�z���            _�Ҋ�6�        ��ڔ    u@�4�Z��       ;.�o       �.	�$��	        d�v�y�                  ���b'��rE��K6    ��P�/��        0-�$*_��       ����        �B�(                    Xka���6
               ^�X�����,$n       �jR    �.:	                �n=jb6	����bJ    ؐ®    ��R��    _f5[��                              �)sy                [��                   7��фo|A        ^@    
��T�륞o�ch)i��	c	   �w�S       ������                 ��:ت��u����7n�ƕ�`�+g^��O�c����V�*�0�$#�i        �6pM       ͸o,Ի)t    U�
0�             :L����լ}�k����    ��    �O�F    ��-Mf�g            4�H�5V�o]�F���<_� ���            �a��                         	       :��M�m       ���           C��M    �0�EFÖ        ���M&;�`J    ���    i2�E�f                n�    c��M�2�%���n        }83            �U�T    >`H��@�               �MX�                ���f    ��Q���/        ��e    ��MS��G�               �Ŀ�                                     �p            ��	��J�       H̡        ��p            ����    uÄev�<*        uts0                       �	�m       -��            ����&��5Gpf	       ���                                 ��b               o�^���(Q,�[        k���`4�        sǫ�       ��7�>&Fm    �k��i��iD        T��j            b1��            ��Y            ��B��%    'k�'    ��`�                    %�`        �����y7�                   �_�                   �cç]8�r�̥                    	   ����UbMQ           	��c        쬰�    �=�        ��       �
�w6H)                                      �Y2;R            �[�W    ����+���    ,�A�              *��#y{�z     �                                                                                    ��+�e�?n                                                                            �%R            �K�                           � �                                                                                           �*p�        b�"0                                                                                                                                              ��?N                                                            �"Fh                                �pi�                                                                                                                                                                                                                                -�F                                        �i�#                                                                                                        �oO`                                                                            �+r�                                       �6                    !���                                                            �?�{        ���                                ���                                                                                                        na�                            gci�                                                                                                                �~��                        
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                      �q�                                                                                                       ��                                                                                                                                                                                                                                                                                                                                                                                                                    �(�                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                7��k                    EA$d                                                                                                                                                                                                                        ��)                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                   ����                                                                                                                                                                                                                                                                                                N�	&                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                   ��
�                8\j�Q�7�t                �էK            (���    ޿�\            ���        W��        .9��   0��/��:    '"c�                   ��}   }�&    ���)��                    ��o��X�    �Iz                                                  �Gtz)�(            ����   4Pn,        �VY6       �5    Ά�6    j]�(�ēe            �?{�    ��>�    �
�            �ݮ
tc���V����       �H���l,	   �L�        1g�n               w�2:    �e�                ^�n,               +)(   �$�   �7��N]4&�&��%�    ��M�tE`                  ����           {�B�          A�~+    ��B݂'�W�H�    ���x    5i�            �Dx            Vx��    @               ᅆ�                    I�A�    �j+�    ��            o>��0b�S���ڽ    ^�* �	���Dh�@���9��vV��    �):h�1�^    'sD��'����j     M�c���)��^�<��       �/j    =�鏐��G��]7���n!c�X�q    79P�ۑ�l�e������\�    �u�G���7�Rz5J�� lЂ�2:���yu9��
:�1�LP$�;E�̬ZKg�!�(Y�|���t	�����X����    cUZ��X�[鏍����h�64z"!"�"i��R    �Jj%�(��    �_�2S#v����oKlP��:�J �u�^�h��������>���k�n�5�`�I8   ��L�    �	�?'U�ֹǵ�R ���U2��]��<2�G�2SaGA�7���2@	�@��
�0c�    ���}v9X��Y�z\4Ĭ�D�]���zSf�
�I�ǿ���#7q@��ӗĳ�*%�$�YC#
���I,>5    ���<N���    �
�T�&��K5    ^�^    .%�H1NL�        �ڱ�]IS��`��=���	v�)����    9��j9�Xz��<]����/|    &_������\+WfeE    �<�e��� [Ӳ�-�?�nqQZ&nq5^�>��nt!�hW���]�3k˖�(k�$�    -��@�V߷��,�D�����c��`��+[�C�S�e�w�@��3Zvͤ뒇��� KJ�fq a�#q    �g��&1[!���	a^>u&p_��n'�Kԋ;KM8��OǱ�5F�yPx���ц�'���	�V�/���ƀU��|�ؕ���,lG@�+3��+(۔�
����		����B�V�/�Z,����.��`\%�cQt�͜��/p���7Z����`�b-/X^��ZAՙ�.K�!��#[~��Z�H��e�9@�g.�*�����ZàM+K�<Xo��0/�q��"��
饳6C3�̺o�G��i?bf�f�6�`�����6`|�=��H���P�<��6SO ���B�fG�l�;�q\�I����ۦ�.˖H��,Zֲ��l48�&ֆ�кL7�W�4>;@�Ǐ������Ȧ���A��`N5(���1}�H�u6�vn��q�b[�ǃIQ�paӉ0���N�VGQ>��1�`7	��Bf5�u.R�����.���Z�W���ة��A(#Vi�ɴ�Y%����dQw����ɓ�  T)�fg�@/�w��N��<ٌ����`џ*sfec��O���2��j����Z����`�؈�J*'���|��B�}����k���J8V1�ܭ���8��-����ʥU^s�O��4�esֹ�w(e��GPK�j��Tu��cN�lٷ����}JF:��1����4�����:0$Ǽ
�w#%�Ҡ��s�v�n�[����Y *W�jnQ����W2z6MqE:|#m����Y�K2���6�'�?/K�֌7]/B�wj�$��{ D�h����60���*����2����}t�0J.��G+Pk��f�_��ZR#�ߕM i���d��j��o�![�:Y�9Pm�Z�
@�G.�-���� ��Y-ҟ����5�Lu�Ԝ�G��=+Lis� �b޷,t~���%q%���K*�	l���sr�:�eE� S��X�=1��Y�eg"'�V/��V���n�%�,���6�^���l^i�⎤�Ѧ��p�P��D��� ���p�r���X���o�vSڻ��>w���2:�rWA�\&�)�	��Zf0�|3��Eٞ~cҪ�%���\��E_��:e�@�D��L2<��PE)!C��~P��t��C"�	2��;�&4*�~��_�o9�u�>�}O�?�.�ӏi�V������'@�Ń��c����h9<E�I                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                ZF0v��..�I���T�d̡>e)�H
$6d�zD��yӦ�s�p紭�D��8���vrb��a���1�� l�jȌA�����i q��D$:�����Eu�YQpn��VX0�!�4s���RoXԬ~����Tc��xi�#�%)
��6-��`�긧W+hb��mi�~��IN.���:��8?2���t���ba���g�t�Z�@��_�_y��l�"y���&7�w��������^i����
�\́�7ڬڮ&�tj��`v
�.&�LbL��(N ��T������3
�qi+��ׅUZ���߈N�HQp0\s=V3os�C��2�Z唠�\	β�4��R�{jP���I���h�g#�s���N��E|���o��|s�=Kb:���,Y,8�JV�95� WC��qx�mr�{*>��"���+�~ZB�<R������©��$    Yo�?�1ө��!��y>�'�8\�G�������8g@	9׫c���JP��#��~�'�%�E�����iK'�)|�b�Hw.��2s�EجM�)��@x8B���	#x�2��{�,Q�E����f�X"�%"�qլ|VA\�o6�����x��
fT �H�{�=��X"~:.�)`�ww��Ś��`I2�c�.�s����B1y�'���R͹��@����S��#�n���g�%�P�e��l"q�s�=^�������hCլ�c=P�C �f��l�P�6�m�r��[}�'>�����rɉ�fu!�L���)Ls
49h�eZE�l^#a+#ٳg�[����8ȯW����躶Tt���wJ�t;8���6BG��W��86��͉ ���ʙ��^,b��(�����t��%��&;����l ^�B�c�E%�������{|�s�~!SqP_�B�ۤ�U�
Z[��P0qNu�`v�6Z������p>��X�$&���#ˀ6��&�Bk�1��j�ڦ�"E�;�SIV��D�
�L�K .�b誜F]���p�?Q/SV�>�!b�&B9�pt>���+�Z���'&����[!G�is��/�����6a�����U��f�'�ֶ�/:x##�,s&�sgM�8q��Ea��K(� ���a��$d 'a��i��Ƨ�ҵp��U3Gø[���mO�$�0φ�V�m߬�׳��|ܴy�(�            =�@ ۠@                     �2�xі�"����P�_{r��F�@b�����@8X޳�(1��(�3f����{;h��k`p�Sb���Yn���������C��1	������@i#�<� 6���U���wc���u�(:@̶q�b��!c�F|L���\�9N�� ^�{B$���E^`0���YG��x;��b<qR�#�K ��r���,���ցȹA/��NX�����	���/�x*N����^�O�Jݳ��JA
�*�bT9��|��rm�ľ{=U���C���}����jx��X����0�'�0�CSxYa�v�_ ���#,�1IX���+Ы�t���֌*�2�j�J�Ө�p��f){W)�D����/�{H�]�]� ��*�.v��LGz��g�����X���ya��*x��ՠ)<!�0��� N	P�͝C��N��`�����"���+"����Z�ӆa����x㥜�����C��#��� {�@��x�$���-����͡1r;j���������6���e�Õ�eX�����J+�Дa���=j��� ^DqS:� �YZ'3��|���}E8L��.ߥ4��~�3��g��Ehn|�����e	��PU���:]�M����9�C�_GHٴ`+^�mSܕX�r~���'�@XJ�z(�V���)�j��?�p�L��?j����P�0<��Ù�<V4��$�����0,��-Ѝ���Ѓ�٣u�96�n�6�G��+����ci�w��h��.�m��I�EEjWL�I;����y%8��J�P��ʊ�ꐚ@t%���܉t�Bþ�B|F���,63o�I�5�H���\~�ݖ�"��lu�u                                                                                                                                                                                                                                                                                                                                                                                                              (  �    �   T �               p  @  �               	  X   h@ �               & A h i e n d i e   h s m y   � �& E d n e l   r t h s h h r    & E r t   e d b     �& H r o y m t   h p p     �& E a i b s r     �& N l r u   s e t k w e n o   v n t e o a e i   � �& I v r e h   w l h s h b w a   n i g i r u e    & H i o s i f     �& M h h   f d e h   a t n d h e i           �& H r u t   w v a t p h i   e l l d u p g     �& N r d i i   h k t   e w h     �& E o i c i o b i   d s t b n t e   w e i     �& G e e o   e e o     �E & o r n d n n     �& C s f w e   i l h t i e g s     �& W h n s p   e d i t p t   r t f   � �N & i a d   n d e p    & M b t a e a     �& O e e v p   o g a n p m k s     �& S p n   t i i t d g n   r i l n c           �& H c q m o t t a     �& A t z a p e w i   d i u s f e     �& D h l i t t i d     �O & e s   i o u s s r i i     �O i & l e r r   t a c u e h   v e w n o t d   � �& N e e d   e t r   e t m t h    & R d n a u l w     �& D c e o e i e     �& T l e   n o r e c s a h   r n r a h w     �& F e i e t t   t w n l   t i m n g w           �E & n s i   g w t f h e h m   � �& R u m t p g h s   s s n   a n h   � & S n a e     �& V a o s r   v d e d d h a   � �& T h w s o   r e w e e                  �  D ��  � ��  < ��  �
 ��  � ��  � �               	  \  lE            � Ȁ         ��    E t y d    M S   S a n s   S e r i f      �P    I� >  ����         @    mZ*  ���� L i u h e   e a a l e e a      �@    � \ � #����         �@      $ ���� L n l      �P    hG  7 ����         P    > K Q ����� E h e e n t e l   t d n u r .                    	  �  �F �          � Ȁ         ��    N d h y   d r h s i v b o   h n e i   r o l    M S   S a n s   S e r i f       P    W � }  ,��� S k s a l h   v c i g o r t e       P    � � R  ����� U e r v   s s a o r   e r t u b w o h   s a i n f .         P    ��   .��� T e n o         P       /��� O h a e         P    j 6 7  0��� U l h o l t n   a s r e n r i      �P    � � � � 1���                      	  T  dH @          � Ȁ    	     �8    E i g   a u s i g e s   w g w h e i i   i c r w    M S   S a n s   S e r i f       �P    � k $  ���� T o e o r i         P    � %  ���� E d s w   e h r i h         @    D L  ����� G e h   a i s e h s r   w s s y   l e n i o b n h .         P    B #  ����� E e o a u   r c i a o e   o i w e n d s .       P    n	  ���� T w t e e   t p r c         @    g+  ���� A t a t g f i       P    _    ����� I l d   r w u t d   n n y s t r   g e y r .        �P    ?E / � ����         @    h� G  ����� M r t i h r   a n t ;                    	  �
  �J           � Ȁ         r�     P n s d n s    M S   S a n s   S e r i f       �P    	 8 >   ��� D a t t k a   h c d e       @    q � !  ����� H f d   y a s n e   i t r   t w r u o a o .         P    � L   ��� I h o h s e t n         �P    s � P   ��� H h c o   n t e o h                      	  �  L �          � Ȁ         J�    E l t e g a w   h a e c i a e   d t n c o    M S   S a n s   S e r i f     P    } � I  ����� H d i i ;       P      ����� R d i   w o s t c   h n r h a e s   a u l n .       �P    � 7  ���� G w e   t b d i e p         P     J�  ���� V d t   l i e n s t e o         �@    � .  ���� S a l       �P    } � -  ���� P l m v d        @    � E�  ����� R p a .                      	  �  �M �          � Ȁ         b�    I l h   n l h o u h n   l g n    M S   S a n s   S e r i f     �P     � �  ���� I s r o e       �P    
� T  ���� U w t e p d   m r g a i a d        �@    � Y  ( ����          P    � � ^  ����� E h s   h s i f m i m   m s r n   r w n i n t t .      �@      � 2 ����          P    � 6�  ����� L l o a a a   t r t .       �P    Q �  ���� E g e o u                       | �   " �   � �               	  �  �O ~          / H h g k d i f h   a o m e s g t o   l o l n e l   h e s h c d   h t i u h a   i n d n e f o . 	 A n f h r i h s . 8 E w w w   n q e o o a a t   t t h l c e e   c r e t p i d   n n b s s t   s u e t i   v c o w c d r t   s p e ; 4 C w g a t h l r   d l e h i e   e i h r s t   l h n n n   l c f h r   h e r c i s m   e h e d e o e n ; 9 O r o i g   i m n i e a u   o u n   i h s r r   c r e o u a   d s e h s e t h   o o t t   s d n l d   o r n d f . S L d a i   a e e l t   a h i o   p n u e s n l n   p a a n n r c   x t m   o t p   o i c m e i h a   o a e   u r e i l h e p   y c e e g n i   o a o o n b s   o i a !                                  	  :  JR l            U c t t   s e o r   n c r t i o n a   m a e u .  S v o   d o h .  L i l i o i .                                        	  �  �R f            T e a e .  B t s e   u t c   s e s g h .  O o s n a r   e t o i t r p m .                                                                                                                                                                                                                     