MZ�       ��  �       @                                      � �	�!�L�!This program cannot be run in DOS mode.
$                                                                                                                                       PE  L             � !
 L   >   >  �     `                                                                 � <                           ` �                                                   ` $                           .text    P      ,                    @.bss     @   `       0              �  �.rdata   0   �      0              @  @.data       �      B              @  �.rsrc       �      D              @  @.reloc      �      F              @  B.pcle              R              @  �                                                                                                                                                                                                                                                RP����;��ϴx]XKC�ԁ
��Xc�ԓ��/�s�o�{���]�.޶(ő�;HAv�!XՂ�ySj��d�I�7|	Њ��;����I�h9�x��RY��Uk[e�b����S�����cL�[c[�$\�>��[��%�f+�?x�{0ƃ�c\+�@V +h��@�o3��r��K�z�UJ�J�ާ���H�1��%�&�ڐg]y��n�bM7h�/*�QR*T�*B�C�@Jɥϵ���
�J��$u�������vdey/��!S�Jc�\�����ub�X���m�r_ U�*=��,���3� }�!r��aƸ������H�C�S�1R;'�1K�:W��ͫ��W�:e}�Q�ON�����aŗ�%L58פ]$@��ĵQx����)9�Nf`�D/N~(QױczO�/�.I���P�����Z7��7A88��B�%&�;<��?梎Eh3����x�{���A&L	�ձaU0N ���f6�|c?�\�:9(/Ԩ̬��_�� ���{�Z�݂�W�3&����W��q�潸�9���X�!2��ªUx�>�N^�'�T���AgE&,�hn�]�r�.�Ƥ��.ߧdN$�|Eƕi��qIV�y����{���E��� ��;���)�����&܂�H.�I(m\�:A�ma����/h{L��#�
�C�⍬������*���
Iޡ� ���1yo<���Bk�
Z) ����-�=dL��&?�[�����]�1�ђ],�zdm����i���88*���o1]*�h�%.P������|��a%����*��AxXڠ�(�)��.U,>ǲ��p�]�3�D���Y�k��\WW�w�/;�[�_8-0a���0��_�BS4�B�-�;�ҭ��*�l�:k��~o�ZIlm&�Z*h��6�yUe����C�g1��NHOl�0c�M��>s��|�%�!6?�U����R�{j�<����}Z��ic��Dfo����zw�C�U����_^�gT��^&��ɺxQ�6�u���b����KXU����!̪��k���[X�53��;R�%ˌ�_����Wΰ4Z��R����*���5�3�޸�]����W-�T�������^i��ʎ�܁k�}�ɡ~y�0+Ӟu��FI��ۻ���-�چ��+����6�?f�AH�jOu0����F?ͱ�F���æ�,V� �B��������h`�u�-��&�Z�k�-����Q�L`��|BAO��D�x�|m����O4�Q����<�E�F��}w�g/��U8�9�&g���o`��X~�eOe��xEcN"`�oFY�@ТцO�O*Aq�\��3��>޷z* =����k���J~£-�;�?�6�#�����8]�<a ����o�tn|��^To������ɟ'�)RIh�L\��ߋ���mi.�o�RG Hq
;��{g[�._6�e,��!���7�S����^h?��m�v��®	�jGQ8���CR;MpN%��,�u��|o�,�gQ[�9m�}����(V4�E�u����~Fm�W����1�wuo�F�E��V�{��������"nQ��`
Ҫ�L�q�Gӗ � �
������
�nM�1Y�$�}3'�N�?�h��v�T�����%�������3���ߍ���c)d�iS+���41��dM8�u�f�"*��7�}�i�#�SX%��T��������=cg�&�������27Fh��o)�8ݙې9�؎7]Yef �Rf��[i74��d�js#rv�s����V����V����]���j%3h����W���/��ӎ�'�_v���j	W =��6�5�U�*XJP"$i�ɽ�x7�.�7�{r�eU��>��cq�l�l 91�����Ԓ' L�N���=�[��қ�voF�F�<>�n�Dv08ؤߜd4�nG5c_C	Z�/�\���[�� !^�	�$88;���?�����sP?����㫭���gp+��{[��`B�L]�%���{0�Һt��șO.{'D�3�4�^E �΅�Oʅv'�D#�o>�x�бɐ��٘t^0��W[9��a]����-Yxp�h�Ã�� Q$:L�_} ���K�ϧ����)���(�E�#؞�Z��b�����
�}cC'{�U�L�>�?��L��$��U�̨y�����#�E>B�����v�6o���h���y���f�v�l��u�A��uٸ�~��(���2h���O��m�wO���*�(�EdK����)��2�~5���q.���^`��~�9Z�	`�3�+��-���4w����=$���ވ�!��zQzv���2�Mua����� 8�?,�c�K�bɌ%&�����F����ʝ�~�����xOm*�ȸ��2Qp�g�W$��xEG��Da��蛀z\��I�C�{樸��,?��먁�~���>�ͯє�����i���p���J#7X�����pUD�)��=����Ssl�$H-��G��󍂹d��Q�/W�����..�����zk`�8�@�7��aւeq�b��љ�I��!����q.��[ĵ���yd�:����ڲ��VKM_f+�����ˮ�(=O'ї>u�a�ml�~B���H1�|�ϑ�MU'TH�a��y�gZ���"5��C}�Xk�DFC��a}/ȱA�>���_����֪9uG��v)�#�A�Ҽ�P"֤�w����hb$p�(���ʺ]`��$�3�@ kL��-ݱ��~��<�����8�?|�oVʖ��B Ѭw��~�Ѭ���m���f֛Y�gt1�)�6�k����%�;j�k��.(�����
3�-KIH4A.���K��٨���H,�C���_߿&zYZ{bz�_�z�I�/ű����~}�
~�%��Q�������a�D�������gk]Y�/���7��%I���2�I+����QI(�?�v�@�b�~<&��1 ���B�Ԫ�&�ǵ�<�h��sf�b,Nx�-�Eeꚾ\z�6���Ʒ���&
K#�3�����䣱�&)���7�h�&h��|-
��6�DSoE�*ޯ*�
���O�ǵ��t�������Sn�������JPmR��:��XP+�Җ���	x妣����۸�I8�N�k�4nc�K��-�V{��m�{����!+7�Q�F��\&�jktz�؊���@�Q�ʬ��fU���=�ɭєbs�ێxT&����f.����-�����&�]|{���6u�^8�X��F�vJ&h��,���������h ��K�2=�_е���e�n�!���%Iz��p+SY�K��ˉ�EM+'A���P߫��ݾ��Z�HoZVQr��:�Ѳ�홯V�Q�l���Ƅ�Fj�(w��<��rv�f�Ot+�CX��xפ���o�x�,Ҙ�p�M���-Oc�W�@[/n��*"�Nv�}��"ᤡ�������6= 6�!�`���lȘ�h*e�Fs�3�>[)�Qq7���ے��h"������$��*L�����"o����t�T�p�aE-x훠�Ε0r�ӟv}h69��';�f�˳h �.���9vd��O;�=m�7:�lW�mr|)��X� 8/���������ۮ�-;+�`Ӿ=���4S'�@�G�8�}�����x ��c��hKqMd2;�;F��;V��b\�|��S���"�EO�9V�0t͆`ؕE'�����=�w>�t�ǆ6"F1@�+� !�h/�ߺ�.�q�E���c��uʩ^��k���Rd�"+s;Pz7wr�8��#l�!��~��%�)nA�`�^7t����!mq��"j���Wh{�/
���x���#<�;�oh�N�B���>g*�lMaad�C��I�f��Ha|K#�RHi���{���0�o�@���o���B�U8LY>�@��� ��l=��UWX5�����L~[�4����3a��K{sf�j��ߝKZ��&�۷����0YK�EQn�u��,k(Ҳ@IT�j6����u�ڡfr)ƎV���2���&�����ˈ��q�T. �q��(��:U�FZU���D9*�
[�"
����� i����[p�ՙ�L�S��b �A�����Z��
G�5I�>���B-j�t����+a���^�����U�E��7,�A7[81E b�ֶs���]P *�b�7I�`5�lӯ�Jf�q|[�Q��\�eA�m˅�Ws�/ `���+X�tu��Dhx�'ڇs6�ν���g9[���
ve�6N_�S3 {���	ȐD�?|�t����eQE�Vt�Ě�+�O�'ީC�ؖ����A���S�2$�:��tq9�#����q�-T�GS���P�0�Pr,�cxO�i[��7Nƥҭ�����܃�x�Uxr�����OP��a�f�Co�m��N�!��߆��\H���fH��DT���q_i��݋��x<��|�X�K�׉�|��P��>H���`�i���bu�͜@�2��ө����-�}Ge�Z��E�zOv�EFQ�h�����l����q����U�@����)T
r�NN�]G�
X.3��7*$喅	�<aw�]��f�ZU%X���|κ����W���m%�(ġ��\���I��$� �;�ѥ�N�D3K��R])�.�o�g/�r(����0���<�i)Z�G��5Uռ�[,�~/2��D���GGU��|��?�	�B��
*�����d��ݔ�!6b�{n������=|F��
�d�����#��s�럀P�0#7�����T���O��f��"*��m]D��K ���<Tq����Z���O�#�M�cYZL�+�5��wv��-�X-��R,ut$�^hm���s���:�w��Z�
�z��-����d�$�B�E*��V0�P���r��kf��
��c�ʑr)+^Ft[�#�Q������:����^�iz�r��?��v:�ωD���@��m��?�c�<ðg
�A�%V�V;��k��0E� ��Ju��zfҀ�J�B��p����/_��Ɇg��S�w2}2=Y]�C��u¶s�.�/��P��M`QWϔ8|x�X4����Mbs�g� m��V�G#��2�0b+l�/��{��L�d��elw�v�?[bP2�����I�N�G�Z�Dڵ}�f���Gf�>,i]o(�e��E��D`��^��u��+br�
��#�AL��Τ����n)kw��Q��1z݈$5-�fAƖ�F���e�����rЛz�&���D�y�P5���4���2�A�>���N��'��`��6odG� ��y�Y*Q/��K��$�M�!v����z�=A}�d�������` �
�ۄ��Z:֯��K�Q�Rj�w/�#x����W���ɸĖ�k5	�pfj�Son�6f�z��Z9�%�t��V�#�z
��&;��p��S�P	O`>R��x!U��)�Qo ��E4%�"��V�}�ܫ*��23��V)r2�!-���t��V�6����aG�J�;\�k�*:�-������{p��a>�`��zP4�d�p�7��m���$]���}&"��&�V��=��<�So��(% ��@���˧��f��Wy��  eLD���پ_h��!�
m����{�K.�e�[����6�bJ���.��+^ʩ�K C�=.}I�[��0CB'EM\��'u�&�p�})d�ll���M�~���y��=��֋��}�h��AߤC�@�����l�k�Uʆ���BQ�k��������!�����e����>�'�� 2���n"{�8R�^��$�<tgY��$v�ZW�w�٩�g@�T۬O��S(R���C�J��|]�z����ҵ1�?Փ&��h%�֚�����H��γ}�D�7����b0��)
?Z8���0��F���"�j����K���/�א��;���]�&D����S����ȡ�5��n en�{�f$��g�!�4%��˕������)�7�д��$T+��̎9;��#�0��Nײ���G�[Hο�6��A0�Q{�-����A�U����i��f���cf��^}�޺X���$Gs}/�q4�h���oE}���N��{��VO�<j�;��<����e	,��M�fo�^�Z��&f�9��&�/b�X�	'��셇�e���!�'�	�i�DO��|�3���td��C���ܓTDj�oKm� Jy��_�ČO�m�_X��8�����pq���>�|�cFcg)� �� *��\��$b/��n���𜂠pv&6���Y@�F�TU1+4�,>�rua�r�*��qVY֘Q���--�c�'�;?�qA��	/�P@J�.Y+�6ia�Qc��+���vV��T�k	|���$��X��&:ȞO}�¾I�,���W�P��Y����p`ȃ�7P\<����L|�G<�"ST�C��eV��5xg��=�N�*�d�_Iu�*��^rIP��_�}�:ʁM�_��{�`�=	v���$�(������ ���d��A�2d?��m��f�Xa'�Ԡ�X�������cM�z�W�0î���XCʀ������=�0�xnXwb��<&U�Lk��wAKr�-n�Q���ʳ�8�[v7B��۱�+U���^��.������G���3KR�/�F���T��KF�̔�oQ�D6�2mji�1���J���Y֋��ޢ�.,b�+����X��> �R-�_b�m.�ٻ��Ժ�1F����x|M�dV����xytHmy����{�.Ԁ�1�9X~��O�z�G	fߌ�~n��SCǢ�("\��Y����c�n�ZI����27���yvxS�{��]6���x�U�ʼ���Q������)�����@�xr�'K�ȫ23��d3�?<!�";��f�5�����pi�m�fV����F�Qt"_d��u�?�n���oC�ag�FEbř�("��R��m�_�&�,��{��ǽ4�MMGk����-7n�6�VI�6RE����,z�Ͽ��jˣ��.�F���w��䈭����_��q�>���_G��7&zKlՄ5K^l��J�� �d�� k����+m�&��[�Hz���$�,84򾟗����g�O!�e�:��uЛC��qi�wP��3N޷�zz��� D�l���u�̞�gǽ�Q�<���"�V���/���J���.��QPܑ��](p��2�9�jٓ�kVc����º4+o姽s��x�c-�+<�(܍\Q�dό��g�0�P���$Ro�.m�Gw�#�Y�
B�H���It�1\�Ut�{�tꧼ�k�L�(��Н[ʮ��i{*?I|���jw��C�hܬ�&�y��K���:�͂�������N�����jE.J[�mjI~5|��G�S�@���Am`���ťà#�@�;�$�g�U�d|�<���a�z�+�>��H�5-ŎV0;�����T?�ߎ  ֮8V�j̢��<n��E��h��tX���-��7�8�;���#b<E���֫6�ddc�ʀ���Q��T�6�O���l�rk��}%C!����ՠ塚7¤�-횃�{��,�P�����;�DsR�����{�{.V�;�B쨀���c��B"����*���o�A�34:��r���\� +I�>|`�R
e'�.䛳7���«�a�TAq��~�;�L[�)+����tB١���tJ�w�����đ :B�H�����]#� O0�GB�rFl�}zQ/2W�sN��ʀ[	:����,�)��|�afH`�p����G.����y&��7h�n�m?M���[׃K�!��[ˢU�~��;�F���V_���9G!'�g�B�$��3ȯv뤃-n�$@�e��>�m�9�ړQw�|���k�Z~!�*1�[d��^[��n����9?����T�c��^y��?K�2Z�����^ֶ��d`jk�E-̷c���Si�a�6�cՆ�-�������qY~�M�.H&�H;s���+v�� ׼X���h�����g���Ƿx�+�?��O1#�3�E�{�P�sŠ��L�yGÓ}��A+��6�e'S��g/>��|�4"�@l1�6��u�]���횱C�|��`�������ԩ�X�F6�U��J�'�B�}�Ǽ�0�5I}[�#&����̗���{� 畫��=E��?�eV[�#2�1������r���^��w2=�(#��Ah�5������sJVI,�f�t\���qw&��s��y��8\�ɑ�-p�>��~5hs�!���2�����s�*]��7��R���o~����ZA�F���PjILe���eE�ʆ�nv�ۮ �7����PG���*�Fu��%���m������O�X*z	�bp7�ѝ^���%�9E����ڣ,�v<����Z�Y�n��ɼ�rU�:��K�}���B��3O��3��x�~4� �8��*K���!g6Wi3��R�}��8�yR�e+��$��)��_�'jt�H�6�c>G��3�����6��ɚ�T<ڭ٢ēD��2֓�L�5�WS �dRR+�~���o���o�:�O?J�3)����.q��#����m�z�Siƺ�3�	�ktyj)9���Z��9*���{�*"�Ś`3>u��!m��pQ���/S���A��+Cv�h�<��e;gh�SՓGh4�6�D|�*$�w�֋o��6E�a$�l��oo�6�uh9�@W+L���#�[��5���c�	�R��FU�(�A@w����1�;-ܽxu�V>{�`�o����+n-����2A^���׷���	<_d�ڨ;�K3��EwLR]�{n���nW�Xy�X+�d�^/=n�=A�7�Z�6h)��#�_�s$��ǩ�"�:��Ǥ��n�����:
���T�W�A�T'�T����&k��}Q<Q�F9#gu��1fq\�e�ti*�|��AQ%��A��/�m�i��tᝠ������=l������?�w�ۡ��щ&����A��b�o��s*l��a��s%����π%^�V�����2��U��ѩS��ٰ4 �U�'~�P�ʠ��ڎ;1�_�5	 2��6A�tj���G	wH���y&=�=�+���dƕ�d[��/��JP�rA@��k� ł�
�w���{\���^����3���S�Y�l���x�+�c`��T��l%���C�$���<���;��g�ᗝ�^
�.�*��1.)�/�C��a��"�M���v*)�{,��i��BlX�ԩvl���F,�a�b�!������k���%��ҴUXF)������{�Yý�}l|�v����8T�<���m��~�,p���1��{g?�kðw�g���7،�y��i���mY��+D�h!MK`z�2)6����-���X=�]�{�����BE�d"��$F2'6�H��]�KtǫAlm��׏N��#�Zޢ�6�U�u�4��p���z���k_�c�_gf������@�@��c�[s�w�~��ņ�-�k1��Y�I�G���(yޠ�h�`���I�ϊ�G�Õ��Nr�R��(�iٳk�q3^:���pPT�oToy/�6*O��K����t.�k^�N��MT@��	Y�~�5�&�+����A��"�T�V�jg �7��L��h��% ��
�U>��`�%��a���7`ת�V
�=��s���G��}�լVp�L�L?�n;��,�)Qid&q����&7�e�����
�w�U�`��9�N� ��q�_���0��?��p���}s.kPB�(=Y��a���c��{:�NPFe3�g��:�P��uS����F����<���g�WR���O��t�A��N�V�c�Ap�`�gnO!�(jW��|�1��j�ݨy����.���p|��e5.#V<���2���M�p���F�zC];R�p��y�P
˻]���YӊEV���΂+!~��#�.&ܻ�sS���X6��eI�t`��w��Śm�+ȷ#�1���۾����_Cҽ-��Z�"u�dd(:���9��:�� D��,�����v����[$ۤp!r� ���!F=��������'Ąs�Ѿ.+?����Wh�(�ᙐg�n�ԫ<S��:,��r��Zߺ\M�.o�j�!�`� cQ�d4p����j�l�)��b(�EmU����;��Ҕ�d�0��齖��&�@�W��	<WH��("�)&�ו��P@A��b�6T��#E�ݐ���6��/߳9Y��@�X)���ִ�3/�8��� 첂�?0�CΎ���r��l��ٲU
 ���B�б'ķ�},�B�ִW������j3�_(�Ca������r�3=QXȞY ���[���Kю�+ߤa�^2b-��Z@:��v�r�<�tXĂyG�
��S���A7���в�2�5�6Q/B�{�0�i'�|�0�Pܩ�|'Q}�K�L��L;��^V8�B��'U�-y�&{���M�{��ھ�~�"���@,ݱ��®�6[��sh+�P�ֻY����/�Z+���!�HPrGτ�.��u-�~}��%;c ���E��yE�S#"  ��C
���wSV{r[��Ԙܡ�t�Q����Ȉ�fy�ō�^����>��]OHz�˓p�i���x���7�x�PÔX�!��I��f����t��:���Y�t����C$L��M��Z���l�ؖ���l��}�-��V�z-+�q�U� .���u��������B�>p�-+O����H�i���xb�����x?Ô/�!��B��=����t��	:�J�������c
C$�������/�V�l�/Ҷ��M����-���V��~+�H�U�w�����u�M�������F>G���O���AѳiZE�x�H����xs�Ô�!�C�����cmtײ�:��s��s�"��:�C$���̒���-�l���������+�-��	V�(�+�hU�Ζ�Ә�u���Ľy���h>���O���˘	�i1��x��r�x�+Ô�2!��E��������8lk���͝W�;ցx��f��lO�O`Z���Kς����0��l��%�8�.&۠D�K|lsj�d�e��l>@̱��`���`d�k��؈
#$���>�4˓�}�p�ڟ��Ő֭�[֒r>P1(����}:����S)�����N��UiC]�8�Y���,��*�讃��/�6��ro�XR��Ɲ��Vac�|u	����P�sq��F��t�.9�#��}�|�"�e��ΒÒ�94<���㊶�����b����6	t��iɲA�}�������8-������nҗ@�ԮQ�߶���G��Rc���Y��wX5��
���P0��7��,�ω�G��W䔟.S�&�bq;��x���N^ѽ*V7`���$��A��iSC �$]�Z�9�.�8�#Zh��ܴ��<�wl���Ct����[�he�섂K�������K����9���2+�>;��V
�H$�>b� !�����D�3�./4�BPe1�����d�n�D���.�z���|����AW�A�9;�3�պ�����#��A�7(�T��k�� �R=j�5�4;��d�L�1��d]A}�L�V�Y; ד�w(��|,i���������s@���-�l���~F��|^���re筆�k��fz�z�撴�5�x[��p�MhL{����P���G�WFm�:����9�ũd��&�p0�/6���H�[@�׷�r��ѳ�jW(�D�6pQ$L�lې�:����"��+����Ш�e�YD����;���c1�#Yb�������"XOy��9�,��ާp�	T�uzo��1^sR�f걕@t��)�H�
�l�E�o�(!�.��9'�zyb<�'�i�Vgd��o��p�ٿm�UR����n�_��c��O~u���]r�vu��s�.���x@��o�iN,�$��S�m�e�5sn_���8 �y�1�����E����w.�BFiFz
|�E|�>�brF�C�!z���0@�n�WZD�?��Yߺ�f��i�h{�~.�A�[��r>u7��T��V���3����j�1�l�&��)����ę���� ����J���ć���Yvw�]�	������p+���9;&嚑�^D� �j9zY��j&����l���F�^��5>Njv(��[�fl7���;4�'Ph`���,W��S(��jx�*,�F,@�j�ax��i��[]o�N��\�ӹ>�$m�d����i��5���STD�],�����jv?G��;׬q��T�NgAo���߭IO��Y���%>�ߋ�C���Rl
oXq��Yͥ� �_����a1�E���+�9��UicA�xi.75�V?��7$�"�fs�M:���\0�>x�(���:@�^����+Y���g��E$�*�u'�`/��8~d��^�-�~db����$q|V���d�%q���pRb����l˶8Q��!l�x/��b�%{}���I]�9V����2�r��g���^D��
�܈���k�4Gi���Q!���0��+��s���O'�v�SV�x���y�R'���&L����bB��|�O�� E�嶺��<n�{[��H�=�>�3�MO��;��m�a���b�g>9���?đ�'v�ze�GHJG��4�ĥ���/X�֖�Z��)����s/���<a��{bM�	�1*�[�wE� _ߜl��YNI�o�0yG���:��MS����s�o]eBV]f�[l����������^Q�w��?�A��e>���A`7G��-UG��M\D�$4�-��P�7�n���X�p��z����A�1��\��5�o4i���565��O�Z�t@��@]@��OTG����.V͌q �8�9�}7�#�����ҳ�dǾ��R��؋8��|"'LgyYWr+��L�׬L��L��fò� ��#cY��]���U�7�}-��d�����&>]&�y��9�*H|�Vܰ��' u_���|�a�Z+h�G]���vd;z���M����^������RK
�Z��n��m����Zh
`�O�X�x B��܁�"T���y�;x��%�Y�M���|pd���=��`*%�򚻙��|�F��1T�I��6�� ��~�;x�t��w&	5�v���7�*������R:�v���ͦ���ZZZ�stk�6��QA�*#P.�-	� �Ʈ6�M-L;�@�ܤ<���/��:��0��$����e���+a��Tt�g;�^�o��^\�Ez b�9��)^�P�WjK1,	K,��q�����jvՂ�郪C��M����?�,� ��HT&�n�����Fp:���|M0�5�����e�W$�"7	��a1�O�G�w )1�5����,��0S�y��^��V��a�9�.z9��"�qޤx�Ry�i���q�M�[p��MY�,��jc��hE�i��#�L�,��8�p?KZ��=QՑ2 ��}�Z�z�d������Ʉ
کK����Ȯ~�h#$�Y��s)jEvok%�B���:�L�Vfef���p������:Oq���>��e�;l�~l��U���=��aт'�oO'{�X�d���n؊�T~ *�&^��_}������ڃא�Id����qc�!�p)�R(��}��
f��=���{㗁���@NU�T�<�k��}�,��[���ha�z�0)�	���ݒ��L�G#�i~�V�,eƎ��H�VO��0�c����Zw��F��i΃��Hk����������'���̭胪Xw,�������9�YM޲���i�re*��OE����"�,����_�{��A1����r��T��ѱ^�;%L�	"�'��BX��뿧���O{��ay���w���W�F�:`�:��� � S&����׶����6�SC���L�Rͮ.��5!:r�	kzAN$ݏ�?x���7BRSA�Y����F��������a��6]�����n��[g����zɅ������W�;�	��5�/	��x 7nh�n�?.��M%	%�g�/�uM�6X�/�K��z���z��݋�y��-�T��۲Fw���f��y�����#�"]X�T<W`@t��I��s-���$�~�u���-��i��	�de��N@��a����,��GW<��w+v���v��u�D�[��,螽��� bDB榎�.��{g̠��d����X�2(Z�۶�t(��FѠ��D'�6EW`�4F�7y5X��Rw�O����ߛo���C�c)̃���<�k�_��)�Zp*�!���5hN��T��_���3�Ǎ2�l�Ι��I��f��bIV��tx�R���ۑF��5��ڂ�T�#,��s�_�U�P	�Cy�כRqvn'�RU������U#���g�ZƧ����`�yր.Xby=��8���W	��M�+����2�5�g@��ko��B��h�AlX����1�SV�����U,�.�vo��%`^���zt/�Kz��3]�����{���5�7�8_8�'+	dk���cW�i.I�/����4}7�D��f�DCJY05`f��D5�
��F�9�H�����tp0���O�+<C������J��0�ͩ�il��o�����5���\%�	�� �[M���@Fe�t2��� ��q�t�����S�����o�K��!V�c,:�!^��ڭ�F��(��Ǟ~�e��V��uN6��Y{4���&��r|�0��������fR�7(�*j���$�g?�Q�����B+���:#������?�J��Y�Ξ�AƷ�e�����d/��g�����o������Y���L|����Wy� �k�t8ղ|�ӻͨV��O�8�A*���M��z�&Ķ��g���Z5��u5s�t���We��l�t�{�ʍ��m�ڹЀߋ(�p�����ķ���V�����엽L>;��Ĉ�����Y;�����in4+��8h��w����_��jv���{w��M�O^֑�8�`��<��4�u�ĳZ����!�/#��ʐ����ǽW~fK�eŒ�y��'. �þʞ���3S�s�a��P�@��T[,a�@��Us,_Jx��%o��2ֽ�~�I�=��M�;�ӕ��JꜤ=u�Z�:3�brL��
�J!K��I�@�W��K(��<�(��� RT����o���{p�3a9��P{�����Tۼ̪���U���J�
�%�Ι2Vne�2[��
X֑������<�j�u���Z�Q�����/��ʱ�W��h�W_[K�'�Œ���7$'� ���+�@��3���Da�i�P��p���T[M��@�Us��Jx{B%o��2��~��=�t�4��;򧕼~�꜅`u�8Z���b����JB
�Fخ@9�W�σK(8A���(����V Ru�[��Ą�\��a9P{2ͨ�ӄT�����L�U�CJ��$%��i2V�D��٬���+@;�M����Tk��V����NzEb0/��aza�Y�z�	[��^*L��H��fU��¶��HR��nZ�j��Rlo ���T5����`�[_�P��mcP���tU"��i0st�.�D���߇S �w��/S8 �K3 *���}���^����s�0��u����Se�ˠ1���T�l]�J�wB�ymz��dQ�{�\rr�k�&nv~��V����Ɗ��΍x�v��z��[���_栝�Y�ЍW2P�}I/<F7���H�544���wE����%@=���x|���^�V%��=;��x��X�C�Ӭ<�6�ȫO�/���b�+�����(�)s҃����+܌�O�'#��o�� �{�ok�Ui�Ej�@����{��Tj
�n�B�UW�"g�҇���q�
b��y����a��}����rZ#��ѱ9=�����H��v�#�vdU�5�^V5�=��y�N<���]��0-Xn�����X(���2�XW�)�j�Y�#��S��]+1����v��J��\'���= ,�o?�$�R#*϶	��>��"�%�B!�u�싨jB|~��j�d�.k8����վ�͔eС�AsLMΡ����m���s���)+��y[ۄ;� i|����?ur6��Fţ\���䅣�%��R��� ����fw ��8�2�Ac7ؤ/J�A!����-O;l�Қ<��),M��;���_]����Aq޾,��YP�� նG�q����?>+X�5T��bJk��P���B�D�zIN�QYK\�O��,�;j���t.~8*{%1fs�໇MWe����'��I�(KY��?��?+���3��}nY
�Z�d����v��։n#@1�,�U��ۆL�ދ�m(U�a���mm��(="+h}i���8��TM�P�x��L������>ˈx/T,�c˩����-�� (U�:�xj�T}V�����j�&���	%����J�-��j��:��1~Ab�aѰ�T��d��ECS	"R �9L���>���v�ƞւ�[2�9���S0�����A�d��ö��VF%�S'�9D��4MSh
֛���+�-�B�k��xs<����f��>��"�2��,լ��k�@Q�ϰ�!9�a�&���|�?�(eut����.��v
k�,N�u/�Q/��0��|�����Ŵ}��`(����Ʈn�:]��*�4�ӟ�"F���] n���R��s(�
\���$h�b�)���v�������}�;�D���!�ezc�a�D��y�۔�n4% �$��Hh6M�L]�6�����Ⰿ���ѧ�*�w(z�_?�,?s�8��䉃E�8$�Y?�y��{�̮I6j6�ƃsqS0xC��n�ُ��zH�v�kG���!���B�7EY�k�5�d�1�v��� �dQ�Qʿ��#$�7s�?��<��H�2nT�h��ď�\�ξ�J�nl�)�(o��Mn8�+q��	:n��'˜T��Hk(�|	��,pX��IPw�Q5�X�Q����X������y� ���nA�D��n��/�<��NrMnQ������:�ځu��2,5C#�h9Ψ���mlB!�5�\4�(a�E ��;
%�٦�����!U��F��;��1
��{��I�>��\�}��n�Q5k͈��/D�n�a�T��]��N������%��cz���ֱxU�u�C�i�������(�f���Aə��O�$�!�YЧB�K��r�/�=@�Z�ބ,��'�-�kV�Qh�	�",���_�#��XYD�UKf�C<@��ɘ
Mꃈ/�!nJ���|E��y*�q^�ɇ�K��7�"���I��ۨ0�ޡ֛,�"��ٝ�)�N|)�,╺��"�����"I	����K�+>�����˞��c��U��`��� ��	W����F�?������W=ȓ�Aet�p�)T������:�?	8�]aB�ѽT�����Z�vz#��A���~��8��a%����ŧB;0mx�R'Uº� T���@����7eq�:=�d����l�t� +aI�$A�ł�W_��y=o��tZ����RԈRІ#{�X#5T=K ��7,��̹L�w	�(�f'���층��V�v�����S(����g�Co�~bĸ�Ow�u�$��$J�a�
�^�O�YtH���r�	�f������F����!|A?�s�XNA�*��3�?���eS����ho(]Z�V����i�&V���^�"kNQ��U�N�0��V�����i;�����#��9��0��	'����nW{���O�� �3���.ޱ��J�Or��lLxzH
ۃQ�z9}}�|�ݘS��`	�BJ�2t0>��}�)�<D�K��@������i�b�	E=�����&l+���ߵfQ�����.]\�ZASn����~J�}�ʜ|�Q֫!����P�M�HA�V_���_�V�X=�v�+U��Ci�R�D�*��g��.�N��-�.��o����8qV�SzP􏴊�Y�E��i�E��H/E�b��欯���E�I�H����@�}�x�OG�du�������+4�!�����Us+�u[�m�Y\]A��{� ��T�[�T��k�y�c���;��*�C��5g��ck�������Df��<���h���B?�%�fZ��E�A�=�l��Ҋ3P�F�\1��%��*khOt�
��F���!�+LꜞG�ݎd�����!��@g֊�.���s	q�L'�`l�Dտ�d���o�Na�#���rBG4�G��=�l�r�!�C��_�\�$��'�N#��U�5�C���Ǧ�쑬�W��Ui<�=�,�^D��?�ڙ�l_p���ȾjG���>��;�"��zX� ��)�hI%g�ZQ~�f�i�3���#��M���b���/�ې%3�ն%�>E"LSۼڵR�%�R���nk��}�_`�L���
�_﹓�g��6]�'9�E�eAR|��8ҁqWJ��۩Rs5y��"�UE�n��ͮ6��þ��,��l
�W$���]���c)I>T��WJ�"�ג��2�Mޭ��Ŏ�=�����X>�f��,ڗ��SH(�QyD��;_�r�,��R ͅ���v,I��%�RBOt:V}.⛿Q�T�zp ͪeI�1��~/����c��e����`��k>��UX�Ƚ�Ap�{�L�;aʙ�9�uwnT=���b$�n���P�G��EBCt��v�CX�A�{�����9V���Hwy�ܱ���w�*[�%�"v�����e�[u��ybWo�c��21^N�����`��-��Z���%�r^1��M5��Q$&����4"�2E[�ˡ�b�[�4�|��0g�k*�R^l0�	s�<j�vok=�c�������@�TG��3�oN>7%Z�&����Br����Tފ�S�nV����\o��/�P�_y�Gp@hd�S�G��:������#�i�l�=H(�WY�O)�X�@ě8�B�?I��"�\��G�h\?�J�"k���]��N�/�S����|����Ws5�JCl]g7���7��j�2��L԰e6�Mhw׬���������T,BH�:J�׸�r�(�Nc��";��u�DϨ���S PE��AH���xU��ԏ?Ǩ����s@��
0;�m�� ���c���i:ҍv�@�k��}�ן����G�`y� ��!w���Us/��c��=�n;��P��ǊV*z>Ql��-�Yjr�`���Vf�M���b�&�O �띋�s�x�"؊�'R�x���(���9�4�H(pQ�]��)��V@�7��0����c���7�拳�5:M� �q�ќ,R}OP���ʜ�5�)���HQ�:gM^ˎ5V������1z��r�4��
���3ZPoj���9K&B�v"�������y����A+�`�t���445�s*%��9[����:!z��93�pPzl0�5�?ABs�wZ;H�雰�w1�V[��/Gϊ����&8p�P�o]$�7�.��x��F;,2_U����:  �@�  XX�	   V�E��'  X�=D��  Y��  ����0  !u�E��E��   �M�����  W�E��5  j@�5L�4   �<3T�Hx�'  =���   �d   ���  ��M   S���S   �  �_   �+��h   �   ��Y�e   �3��Ð����σ~ �_   ���_   �F�W   1��G�H  h��P�V�=��  �A  �@3P���9  +�J��D  ��  �E�P�L  �M���  ���~���  jh   �6��  @�  ��L$�A���  ��QS�O  �5\35��K  W�}�S  ���Vj^�t$�/   �F��}  9��  ��hP�a  ���   V����������  ��������E��   V�   �f  P�u�l3���  ������U���@�} �  �  V�����   S�l  �E�[  ����������  QQSV�6��������D$����Y�f  ��T$3��
���������!   ���p  ���U�1����A  �L$�  3@V��+5��   �@� �@Ð����+���   8 �~  ��  �4p�{����u����A��  �������SU������P��Q�G   �  ��  �|$�  �t$�  ����   ��T�  �Y�]���%  �A   �Q����   2���d��5��0�   ���E�P������V�t$��������E��p  �Ð�������U��Q�}����5|�5x�5t�:���VW�����P�   W5��~ �~  �����h�����hF/�����������J3Ɛ����B�������   �����QÐ���������C  ^Ð����9��l  ��   ���������������1�P3���   3����G  ��   ������  �a����U��Q�P����������E��E�}   ��  ���  �t$����W�]��hP��   V�E��]��l  �e �G<�/   �}�}��#�����   ������U�b���Pjh   �5��  �t8x�D> �T���P���I�����9^�)  ���   �\3H�H|�����E�U�g   Y�'������}  ����X�U   P�!�����E��S���i���V3��"����a�����Y�  ����SW�H�x�������#��"   ����  �������Í���Ð�����������^$�N������f�� ��� 0  �j����U��Q�e� �p�������������D$�����4�W�Aj�����@�Q������� 3��������]���������   �~��Z  �����`����V�  �U��Q�M������e� S�]�6���P�u�p�)����������A<�a���������N�����^Ð�����   �5������q���^Ð������               �@  �E��E�� �   �����[   S���_   G�M����������h����1����   �6��������C   �;������M������F   ������N   ��  �   ��d   �؅��G  �E��]   �83X�8�8�f   �M����l  ���������Y�   �P�����   �E��   ;EY�   ��   �:   P�A   �8 ������:   ���h����4   ��8a�%8�-   ����   �j   j@�n   _[j�s   h���V���l   j �`��������   P�>  �   ��   �   J�I   �������H   �E�E��L   ���R   �6W���O   X^�Ð��������h��b��B   ������G   Y��  j3��A   �E;F�����?   ���P�F   �v�F�O   V���W����K   �M����U   _�E�P�����X   3��j   �E�M��V   U������   �Q   ���vP�O   �� ����_�G   ��   �������>   OY�4p������:   �C���_�5   ����4   W����S�=   ^[�Ð�����19���G   �E���C   ^[�Ð������������������   W�����P�   3��L   �-   SW�-   H�   �Y   �   �L���_^[�/   ���/   j�   ������$h �  �   X_�*   j S�+   �Ð����+Ί	�������   �  �E��   ^][Ð������3��
   �W  �   �   =��E�P�����j@�6W�   �E�j�����Z��E����   ���F�	   #�@@�   ;Ð�����j   �v�   ���e   ��������[   �   ����v�����PW�   �u�֐����+ъ��   �������   �E�H������   �   ��9^��   �U�Mj^�   �����������^���jX_�   �^  ������������Y�{   �   ^[ɐ�����3��������������P   ������E�P����������������Y������~����u�ΐ����+M�	�������E�H�����������T������   H�����H������M𐐐����������	��E𐐐�����E�P����������� }  �����Y�   �����@��   ������   @���   �   �����@@��������   �}�ϐ����+Ί	��E������H������u����������E��M������� ��E�������E�3�������} ����������E������_+�^�����[�Ð�����          . B V     �         � ` �         h h                     �          . B V     } ExitProcess KERNEL32.dll  � GetDesktopWindow  � EndPaint   BeginPaint  � DispatchMessageA  �TranslateMessage  � DialogBoxParamA USER32.dll                                                      <�� �ev05       P   ,  U���      `   @                   �   0     ��H��!      �        �B���3     �        ��@�3     �        F~C	�2                                                                                                                                                                                                                                                     �J^wÃef�05   �.�    f05�De�R^w4.� ��  �   ,4�2�5�5�5�6�6�7�7S8Z89n4�3�3I64�7�3,;�;A7�6�7�2�9:;*=F=w=
7�455Y3�2k3�:�:�;�;<$6*606�2Z9z3�3:#:(:-:�:�:�:�:�7&9,929�5�6�6�7�7�2�2                                                                                                                                                                                                                                                                                                                                                                                                                                                                  =l7e0_*Y$SL~zGNOK{Fu@o:i3b-\'V!P~LH%?$zIxCr=l7e0_*Y$SL42�1\ϝ����K���