MZ�       ��  �       @                                   �   � �	�!�L�!This program cannot be run in DOS mode.
$       O��].��].��].���!��Z.��].��H.��z�ȸ\.��z�޸\.��Rich].��                        PE  L 2�yF        �      p     �           @                      p    V�                              P   P                                                                                       L                           .text   �                          �.rdata  ^                         @  @.data   PY  0   `  0              @  �.data0  ��   �  �   �             `  �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                        h����ˎ  �8��$׊�4$�D$?��� ���ЊRhg1��Ff��(��f���s� T������ז �����E �E覃 �E W�U��� f���� �I� f��f�U ����4$��$
f�l$f�D$�d$P�6� ��
��蟃 ������Y���Y�f��^���� �  ���c� B��  hc���趀 ��f�E ������M�����f���ƛ h<����=� `��\$D�$$�t$�d$H�� �ւ �BhH���蘖 ��m �$$`�d$,��  f6��$�W�`�d$0�~� P`�E �4$��D$:�d$@�  �D$��t$,�E �$�D$�$i�d$0�x   Ȁ�@f�E f���� �訕 f�D$\��D$f�E �D$��d$X�B  �`�t$�d$,�� `�E h�aX�d$(�� f�$��E `�D$�hoVэd$,�ӊ ��t$�h*�P��$.�d$麊 �� �� 龆 ���Q� h
����̌ ���f��$���<�ç��f���U ����Q�f�$9h�(ćhN���d$�[� �Q�L$H�$�$��t$H�L �t$8�E f�$�^�d$<�1� hp��W�D$���D$��t$�t$�E `��d$@�<   f-���D$�X�sf��f)��6� �ES�T��d$@�   h7�d
�d$L��� �������f����壍GP�V� f�E �t$�d$0������L$f�`���t$�d$8鑉 ���u f�<$�������4$�d$�S� �����O� Uf��f��
R��f������V��f��f�Q��h    �͋t$,��f��f����f������f��f����������f����Ĉ 4�藋 ����ќ���    f��`鲋 �\$,��d$0�� �t$(�E �T$��4$�d$4����������ъE ��鷊 U`�����f�f�� ���f��f����f������`F��O�~f���f��4��o��� ��� �$xf�$�t$<�E �t$�d$D�|���f�4$��U�D$��E鵋 f��f�U �f�7f�E�p����t$R�M 藋 Ɉ$�A�������������+�5zz@z�Ë�$�H����%D @                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                             �!  �!  �!  "  ("  6"  "      !  <!  
!  �   �   Z!      �!  �!  |!      @   �           n!      �           �!  <   �           T"                          �!  �!  �!  "  ("  6"  "      !  <!  
!  �   �   Z!      �!  �!  |!      �QueryDosDeviceW �lstrcpyA  �GlobalFindAtomA � FindFirstChangeNotificationA  �WritePrivateProfileStringA  xGetLogicalDrives  KERNEL32.dll  o DdeCreateStringHandleW  �InvalidateRgn �TranslateAcceleratorA USER32.dll  2SetPixelFormat  � DescribePixelFormat : CreateFontIndirectA �GetObjectType /SetMiterLimit  CloseFigure O CreateScalableFontResourceW GDI32.dll                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                   �c���r�
��Ȅޙ�������ܨ:�& 3�)D/2�9;>E�GlMP�WY:gbex�oq< z���&��o�>�͞����Y�\�ڼ�N�����������������:�6�F%(+~247`=@ChJ�OjUX`adg�npszy|ʆ1����u����6�������
�m�������߂�������P��>
d�n�)��33xB��OB��SMf0�[mKie~X�s��;�O�x�����a���6�D���ۉ��b�.���I��c�i|/�<��'&\셽&�AǇHАUٙv�{�x��}s��΁�ϰVة��/mp>�
J7�S�(_P�jg����?�����J�M}�/"%+�~0j6O��DV��V�F��\fߜ��~�	�~�𒞑��������s������������ZY��������N	�\�3B�"����43��Cu3_���{b���-Z��{~J�L��ڽ�(�g��<�:��C��W�W�M��Br�J���a�QY\���"(�&)�sVI��)#TJMۗzaܗb�x��}Þ�hN̉�X�[띶����;���/�V��-k���!�Ec�����L���I�r��e�.1�}B�͎N1}�RU��v��}�w.�g<����_ʜ����*�.�I��4�)W )P��'4�qS(��?L�H1r�TG
7(*�/�ZE�0*� KN|�{j�.�eݐZ��{~ȫ��R��$�ê�3��z4�H��T�Z�b�\�X�*p��1�x��i�l�	�z}��&�1��Pz
�"���A�$qh�3�u���O���wtO��+�Ȼ�8~�oż�M	��N	�L�hU�qf�|> �F�ӛ�֩kF-��14�*�:.(��;�AX_^a�0�u�4�!}�Vp��L���q���86B����H�����U�b_��v3D��w)_�Ce'��	)-03i�'Jx��NMSV���of�K�iEA>�pv���������;6(����;���N%��i�i�i�"���t}d)�j0y�!+D��9Kq�Z\���%"���a�p��Q� ������ٴ�+ɯ��A����Mz���b"�T
^,xk�C�t+�^(N�l;�+�|F�vWō`~ҝo�g�~���r���d�̡s��ز&��1��:��2��A�B�^'���i����-q��	�c1S�*]�N<��69<ʓ]�"�T��~�{�ڐ�䑳r�����*��7#�+6H1��DA^.��RXb0|o�G�x/�b0R�p;�/��N�z[ɑd�!֡s�k篂����v���h�Хw��!ܺ*��5��>���6�E�FIb+��Z�%ija�o%�וM0���{D0�G��YɔfԔkݥ|䯅�ߎ����H����֭��w,�� �=�D �O��\'�P�m5&0	i��G��V+��&�b<�-03��Tz�M��uɞ�|�=�o��̚
����΍"��3�:�E.���R>�F�cL�2�_�yI��X!��$�a2�qC�qD��Y��bʼkՖh�%�_�ۉ��œ�T	Ӟ���!ݾ,���9�-�J��F�`$���o3��~�?�O*�#N���I���#�!8�2�����`��/L��mp�v}|Sp����$���󥾌���E���1� �&>�=��M���q�M�����^Lw+=�wZI�̆id����[�^pbڍ��Ι�B¥������m&�ò���u��Ϻ���4�/���R��x�+n�N)\^dg&!3%�PW1��byE�vL�W㝀a�gߒ�܏�~��n�ɏ�\��,r�K��C�۪z	��
0��Q�Z|6ccZ��P��.u��x�7:ʌgb1ԐRUWςuc|��q�5�ހ�p�����������6���C���t��[���z��r4
�D8��j]�����������!���J�uh�S謇z��W�(x{�׃���b~|���m��	B�N;�W�,cS�l$�T�GC�/�VW	�	�I�e+v�q+��?K>A�FIMPR� �gfehkm���{��C�¹���2a���t%�A/�)�P�����]C���w=��A�)�[
�]a+�m 2�v3��@�"�fCF�M��_^��S���dƄJ��ђ���.#�1�'��M1��R�R�G�d�c#�c��?��̃3��L�w)�82�=;T��I[�IS�c^�kiA�N�F�v}��Xu�x��'bp��E�C��6�]���t��r/����������Y�Y�e��225ŀ.�ьE��xqZl�ed�o��h_�}��q������쟱/�����缿G�<�X�5����i&Do��R�>tX��w�&8�$�9�<�E wT��Yk�3Ommpjg��Qj������`f�4��'�C��6�j����N�j'��`���}����f�#=�o"4|��z�ozb��Oac��]`c���r�w �#�����嗩'�%���D��-�"��������?�y��sH\;˛� ���ˍV�q녅��-FG�@TVY�G-sik�5��
�o�����T����;���6���S�g���3-��(5��J��=�Y��\��adl�'�j {��7:<pB[9�Pb�S�QL�mp�<�EA���z��"�+��܇�u�<�����N��d6���y9�K;����l:\��@f�W�JřfΠo��x�iI~gil��Q����ȃ��-�4��?'���L8�@�]E�$�Y�sC� �R�
���*�\5�sF���wA��JʜkՎh��}�~�;����}͜Щ��k$���5��� �1�K��Z���k8�r�x:��B݁L�=+�|$'*��Lr�θe�B��p�d�փ��晷r��������2ǝ�Aڬ�R?�Y�_�h2s�y6 �O	�[*�M+��<�n9_��~L�<ČWˏh֟q�*㭀�x��������
Ɵu�ղ��*��1�7��@��K8�T���`����Ix5���Z�Z)ch�g��c(NjM4�4h��&�fGJؖW�d%fmh��y�9~}�)ݼ�� ܿ���R��r��G��=۶+^���U�q��d�K�sf�!5�%(��V7:ȅK�l��d[]Ոki�o���}��NK�-U"[_��+r �<�ܿF���]��,�V	��b�n!��ko�T�(��ޠI�'!�HK���c�(K�lo]w�;琇��\�_�����<�B��N���}��(1�U�u��P3��^`�Z�k%�gJ-g�G��O�X�տT�ߋ��j�X�0ut��qҭ����������A5����E�Y���e)���Z���N���Vf�@3![=�14�@�OMSO����#lg�n���}	�
G�������+�0�3�@�5�1ʵ�e��F��Z��c��m��SX
���( �#��*�9<�	���\W����W�8n晈c�1��[x�.���d���?�G��Q��ʁ��i������B��?l�o��
!�z6H�*U��\�VY\G��hkdIÞ��C	i�R�;�梴�2������R�ڹ4���H�����f�QTu�u)�kF9��14�~aP�ӕp[:��[^zU�vy{�p%���"��.�/��:�9�B�Ơ��H�dN�c�Z��k��2�KNX���['*�e~:L�@M�T�Y���I�dv���z]��~�M�u�Y]������t�+����>�ߓ��D��P(1�h�b:{���\�!3�^���9���0�@R,�Wi]ԅ�uG�r�x��Xˇ������Ϥf0�;��\��ճ�o���b�X����^�hL�E�=��d 2��3S0�7:�7�^ԍ_�Y�$!��X�s����}p?ݑ��%k�۩�w��L�J��Q�����8<R�X���.� ����G�\�hK2}��z]LgCEH~M9MXZ]Kz���������Ѵ������0n&���$��Q��j�:<l�D�B{�y�RX\��`$n�,��(A��6H���RҗU�^�D(ehV��s�*ρ�֘w����'��2�����:�M�UϦ!a$��~����d�E��p�
�М[�c�r�i47}x�K��:�Y[^�L��mp����
N�p;����+����Eʩ$���[�8::����y��R�� Y�'*n�2�q/��36Ɖ3*z�KN<��I�G^��'7�y����{\�~�I����9�฼�N������c �?o�G�����!�S�R}�ݕ&Y��k<G���Ir�Y���j�v\��}��IMQ���­/�ι;�D���?��P�����?D}aTXY������"%�p6���B%���ILORU��n��w����šЮ�ں�+fk��@��<�Z�>�;��5s��}'����V���	��n�tj69��
ON:MY\,b�5�p���{���������/]̯��?��P�"��p,��n+s�|��Q�]�*)���&k:w�L�Z�V�bQD�eh���|�j�F��ߑ� 쟱�*Э3��?%��'V�/�����8q�=@�j �C�T�K���D%(�{)�p=@΋QVU��O찋rU#�vy�~���\yV����e���&��F�����V��Q��Y��0I���z+�O���&�C��K;�fU�M�xg�ELfiWq�5�=���v����"�+�ހ<)���@�=�ZO�b�%e�[�w�}�?6�v�J��D��e)닍����Ew5\ۗz]��z�[����{�?��o�����#�)�(�9���>|9�K�HD�mpZ���CE�zQ���	�/�x$=�~2D��5?XʙM_�C^�)c��63����~p����u�c��5�;�D�O�����Ā���v�)k:�NAU0#�L�oB1'�b=�W�9<�I�K�Y� �s�-�p��z�A�s�����{�Y��-��+�ɴ,zK�$$���`��d��:�t����	�Z5�� #&�C���D��S���\UVY��i�-Yt�?y?���x~�#�,�5~>+�E��l��(]ʞ����� ����#
�e���J��76�V·I2I��MY�j`���`�^�s��Q���� ��'��r���<�O�K����YU�+h��/~I%΋ˇ��� g��k�B5�F,oVu���]�%��)&��X�Vm�g���޽���"����6��/�I@���
�J�C����$D�	S�.�]8?qtwP�,/krtk?Q�32�}SV�\cce񯒍��h�����������6�=��E�Mה��@�&�"�3����.!��� (-.1�J9�L�A1ޣRU�䢅x�iX�݆a� ���R����.n�����A��կ�SI��a �m=�v.�KJJ�E�g���g8��9��{+?BЖO۔l�����l�<�k�$u�������]�����/�M	��]=��^���u�yq�z���;2�dGV9,/2��buFGIb��Wi�覉���u�����I��CF����8���B&���[��+E^I�i<x6��k�N1Dc��FU~*�U`6OђDV֐sr����e�fޑ�:��������eWػ��Ӣ3���B��.�2����/�S� zC�}��J-0�'J3Uu(:��e�8l�BE�9�<H]`�}�/�{�1̍�ӠV�"b�����&$ͨE��T�.L��W�t8A~��tG�O2-���D?&�2��9��:S�D^�T���ꦉ�j�y5f�|��n�H��\�d�Ⱥ��$�θ���KJ���O�c"���]�M���R ��OU$��1477<?�.�cOR��v�Z��rX��y|
Ʃ����|�_���4�Ӿ�/��O;��#,��C��m�j���*���db�j���Q���A���0T�QT䦁xKf�lo��E�D��ܷ��p���ۡ3�2)E�M��V�R��[�?l+�g#26p+>%}�`R�A"�M<�~Y\#�DGבts�樃~M��nqÞ�k��?L�ټ��������⹼B��X��J?��s5ڦ(��G?����_:1��%(��@��:=@��]�ܞypC�dg�e�wpg�Ѭ�v6��(�&��(�=���>=��B�!$YX�"]�<G�;)P�R-,�~cn��*�03Å`g*�xKN��~��𲍌W�x{}�Ӯ�x�˙�,��ȓ�ᴷG	�ۮ�n��Z�On)�:z4
a4XX�(V��,s����58;�ADԖq`;@�\_ﱌ�V_wz@�ˋ��"俶�t֪�= Ρ����')Y�/b�:�8q�B�g	�p y�i�i'��4�0�;"��CF1�|RU�f��*��\�b��㆘ۉ|2>��0��<��HѬn2���C��W�� C��J��`8�bpP$'�z8�h<?ϒX3��TW# ��R������z�l����b����8����9��T�\�(�S�*=A�;����L
m`&~q�%(��"O>A�����XЃf�)oV�wz
̧�qd���Z���/�-��k鼿�G���$*.e���V:���k�B%$�N1Tc��@wB%({��X�J=@��4h�UX�i�ˎ�p�?a�ԯ����-����<>�۾�TV�$���-2��7@�|�|5����Bi4'*}/�N!�bBE�]��WZ]뀾�m]��������`��Ҧ��������:� ��U*��K�p.۩t��[�Аך`;2�0"�ML�OK;>̈kb8R�䨃~�{��������ZwZ����a1#��[^adI��X�'�S��*�����ь��	��[�oRq�6�U(hIL��}袅|������჏���������g��հ����������	1�b8��v���� �<�����(��9��469�7AT��OQT䦁���/���v`㠁�J��V����k�����=���Q�VL�(*_������Q�S�]�[Z�lGfrg�#7�b�-JKMP��}�obe�j�Y��z}C��֖ ��,r�����:yD��<�Y��c$�n-�w/� ��D!7�C�4[&�[�7d���G:=�^���s�eX[�NO����Æy|	ԛ���"&�賦���s'��J����PO���S_rl>��J�7�*�Ռ��h,��5��!p*AD�֕xj�m맊���� ���ٌ���S���¥�!�<��FA���@�\�.��\�����W"���h7`��M|O25�v��)F�q�sVY�v�(�~�����ϓ�Q�Xټ��! ˽�;��1�M���f��.e���r��:50V�](�Y4�v);�)�}^��+IIL�K��vӢ�b���1a�[�p�]���������;��FỪ��!*()ĵ���nT�z` �L�S6-�aB�%������@?�D�oZ�EV΁lK�ylo�;�=���v|� ��e礨6��7��GI%���B��f-��_�{@��@�U�*��_%��mP3��k:w�h[�h��zi�O�m�t�>�M��������do���y���H�ʹ ���0���`��;PW� r�t���W14�7@C�)�Pb�m?�bt��5{=�Ћ����֌�'"�y���v�� ������շ��r��8�3�t���	B�ؐ}��w ,/f,r��CEHɗ�4�[m�J�m�E�'V�Ei���T�����x1�����C����ۅVl���}���8�
�JQI¤��Y(�8m���v$�K]SVY\nfnl�u,xz}��(����P�����L����$����XS����-��:9��|���� ��9q�/S�:���Ta�9�Ζ<�W�Q��e*�Z����z��ip*,��$߁�0���'�E�����[��z>��r5��R���M��b5lo�ctw�r$���;�.D]��Rd�Q�,u-�3U���ä��sޚ�����<���P������f�l�FHH��L��HHK^�u��i.�:��Y@�P�X�ՓX��Z�j�*on�E��@n�	����� �j��q�IʕR�R�I��2k�q6�p����T�dcC	m���&igS��GI�CFINښ8��t�jl�����_�F��q�����������@~5�Q
��� ���o{���6PtWB|�_��Q�iz��18;�AZD�Oa�f��CahkW��x{�����!ި�hk,������JE����]���7��6=����N���k%�2��M�),�*�<ry�P�O��_�W�j�k1��\��}��S�����.���2�D	ǈ���Y���e*�k��2z?x4�uB��r0�2?4�@C���eX��M�z�\�u�	�zm('��!ܒ��6����仾L���&��a&�/�<���~A��Z'�Y�j?�i/�����*ǋfQ�i��/�c��gu��oru�����QӔ����Y������4�H��I�Օ�g'�c�&>�s�Ƀ�
�e�0{_o0�5�~?��/E�PSU�`�ZM��nq��~�O���V���e���-q�8�-��@�E�%$��?��<�{���~�cee�k��9~��*��=@�6�B�\�cF��gjX��}�:ò��ۉ|ѝ��3���M��I������i/�h�HeL�f�pT�M�ԨH�y��8B�gG�KKN���T^�(�􀳄6|A�Mژ ۉ쇺=��;�������Q�.0����6o�m��FLPf ���m$m�j(�{,/���c�@�H�a�Tf��Z���vY�z}�֔w����+xҰ��.�L9�S�������n�g��}��N����;~�����<7��,�*A�;^�W�rvl�u�~���s_ޔ�b򤶨 Ӿ论�9��R�G��P��&��M��L'�d4��|�	��=02[�@R��7�=`�Y�lKǽlo� Ń	ql�䍐��" ��ϰ*�G
���c��]"�+ƛe��z=��!��-�\"{��|�5�8;i�hS��R�}hGb�hk����?���}��霮̪m;�A�A6���Y%��6c	�lR��x^�_�\�����+�j0fsA��F���7���vi�d��xv��psv��]ȻTUո�����e�+���(�H�` ��d����9��GIJ�f�	uc�\����]03���Jh���[�2ciA9q����<	PѴ����-�!���=����T���f3��<�p��y��QRV[��b(6{5����� QD��ڜwfAQ�be�j╈vk:g��Y�(�Ŵ1��|ֶ�F�����)b�h%�q>�*�|���O��n$Z�*��\y?��sq�`�'ũ$��)��psS�Q��N�S'ǚ�)�4n�"��T�` �֚���g��҂�f�pT�M��;���,J <�E��	�xKNڍ)e�a�@�����}u[̖ؔ![5��0j��y½0�W���H���"�Fd�1�w���Gׄ)�)˜/2p���K���T��aGa�%�r��=�@Ǫ��՜�"e�*n�6OT���-�!%�����>w�CFKQU�����B���-0��I�G�>O՜Nd�^adv�psv�d�	j�������&� 0�LJ����]�]�S�K���t��JT��Z�ՌCQჅ���76��oFEH�N��E�o!&�3r��w�b҅�Mk�̣���O���D@����T�O�L�j��y���,�C� ��M$#&d�c658��,�ǃS��]\_q��knq�>}�q����'����*���@=���E��?H�"Ȩnl���x���>�f��
�|+.��5>�\�HVUX�]v�k}�7��<������2Ǟ��.#�1��:���������`�,j�͏���y�	��	�ޛ�H!,/�.�{E�18LPSדe�k�o���cDƏ�+�����_"䲺Cq=��JƮ���`�"�n4�q��:4���5�O"�."�%��m6:=������N�3H�cgj�i��~�����[$���4&����}Pf����(e�c������}��^	���%"�`+�3�Om��,�GKNa����hgj��A�h�gK���Q���3�j���I��=ҵ���g;�kQ��y�Sr������%$���C:9<��T��Pi3�^p�&�H�0�|{~��(������0Ы�6t+H��J��%��K��r�F{�w�-��L��C�),�4�C=V��K]�b�J��&wrqtw��kƱ��U��b-�����	�ש��\�\�R�f���9r0�o�DW�5�ِ���14w�%��FI�G����iL�mp9z�|
Hm14�����������Q	��L�J�����;==���y2��F!�
��j�o�q/�r<�x�?BD�WMf��[m�e�h�v�w΀��܎�V�*�*h�1�.�K�����h+���	��~;��W��\_g|�l0tw���*�9Kq7,V�MP���(�n�i{Vrwz
�{���P��*n�����Rö,��a�W�/y<�ݰ���h��h���W$6��;MA����p�b��_qeꏵ�t�y�㦕����V ���.�ͼ��V ��-�7��l��诎6<�����5ۂ<�z ��8���=O��O��Xj椇~Q�ru�ߢ��
���$����F����w'�ɐo�蜦��T I���K&?�i�*<�&)��VE8��̈kb�_V����fxj�U�x�@��*�ړ�[�j�tS��̀���8�m0��c��^z6
�T�V14�q��iLK~����@Cӕpo:�u[^���>^���&�֏��W�f�pO����|�������VR�'e��+�%y+|��R-8����eHOz��:�<?ϑls6�qWZ�o�������¥��K������������<z1d��;�E)�"箍5;���%�rg��iDS%]���6H#P�DGבt���'G�hk����b^���س�}p�����ν;������Te���WW��W�`�D2�Ԙ
�W:Il���y.1��^m(�bIL�����F�*���w�y{��v�j�� d�i�7�5���6�Tɸ2��jW�k��f��o	�P�2an�-�t&�+58�/-o�Ÿ��VE�[eh���i`_8��ו؊鄀泌8����ֽ�K�K�]�9��9r�p��w� �O2d #%>x�3E �/@CJ�Y��b栃j�i�V�svye�t���˓��������@���*9)���I������l���R��v�G�x,>��#�)L����W�-�Vk��`�t�>��xj����	��r���7�5yľ3�M�X�X�OU
���&c�}t�r������%5z�)6�>D�@0��Gc�]��fQ���`;~{9������Vޔʪ�����E���Q�&<�.�����m����"Y�Qz�[�\�&i�n �B�N�~��>Ւ\\j�%he�1tq������O�^[��/��'��>|6�2�Y���������Y~>��_l
��l�$����J14"<p ƬYLؘ]㟂i�m�������D����]�����`)���8p�����>�S�M� e��&�mނ�����^��cfkq�v �w%�P��=Ou��FۙS1�(�l@�/���?�xЌ{��Y��kht��5��NB��&]��\���ph�OQ����8��Kh;�!cg�=��*�BA��;���j�[�p�7SQ�tw�e5����ࡀr���7����տ�S�Q�*04J�?��G��x����=z#��u�(+��<�x��_�:�[^d$��8X�y|Ǎs����� ���7��@ ����;�7-� ��mx�8�A�}L���o�"4']c�nX��͚DZe��T�Ե�ckoru���;�Ћ��˨Z1�嗢�s�:��5�Q����]�i����u4$��P0�L<��P�V/�;7�:̙Cʉ�S���^夥n�M���������i)qe��n���A�GƎ����த��t�6��D�Q`���d*������&�$;�5ORU�#�ew�����a$���'���$���������>��Q�� �� {�����D�
��x�Yh���!G+-0��]lAQ�KNQ�~`cfj�����A�3����ʦ�0I��� �D�~�����e'�X�R}Q��dg�f	�r��>� #&,����\_C��=�qSVY��i��o�_�p�;������Ũ4�Ѹ(�!h �ճ�6�5����Ig������vo�n#��&8�zU@��@CӍpW��rI��jm����d
���ҵ��ķ3��ϱ)��5���A�>�=��5Ѕ��z�����H�jE8�I03Å`G*�_KNޠ{rE�zfi��z����l��� ⽬�̼��9��E��0��C�������r.����{&%��;�3}��S:�|_J̐kZ@��e\^�ig�2�u�=��zt������	;���/��H��C�_#��6˖q���8K�u(�����fI0��54��)�/R���B�s�t�9��n��u�ۤv�ڳ%�%l/�$�:�F�O�A�\�a�V�![f��J�	�b1�!$��5�I�<?BЉc9V��x�&�c�Ñ�M	�˭��(��-k"����2�L��[%���lY�s)ln��Ò�#����«�"��O�+�Jw�\�O֞kAc�~Pm��y���	Ѧ����-��2p'�D�J�M�C�_$�b�X�tI�������Iikk�ك,u�(+���[>�HΒmTؚY㧂m�r����ċ�N����A�������� ��{OC��[��'����*P{�L\��� 	 �kNA�G9�6��J�E��f�T��h�c��z�:�����������"��6�&�}��������b����#��v���	ɖD�+��J8rk<P�:�QO�e]��fs���͘����L���\���d�2�0��7�����"8�>��U���t�t�j�-��K�N1cl�`C2M)+.d3�?B1iK�Z���c|V�q��9�����ҵ����q���1o'���%��R��k�;=m�E�C|�z�V�K\w�u+�n��03�$�/DG�N������e~��s��vto����#指̹��9w�}K���R��%�O�o��a��F��L/o�r�wz���1��6tҿE_	�U�e�%�u��5�o
Ƃq��O�^[� ���!Ի���P�ғ��/h�47?�d��=�N�6
�C�f�8(+��� �A@Bk�Pb��G�E\�V����ȣ�m���П�l2���3��;�8�U��,�Q�����ڀ����`����[�mHG�qTKP�?Bp�o^�KՋ�'�]吇�����7���umD��)�Ƶ�8��؟���S�ߺ����(�f�{7�/�Q,'�2��dG>y�{VY �ADԖqh;Dk\_�p�����bP��س�}p���/�A����i���=]>�iJ �{F<�R%�[U�g:�pN��R9�xb�ɔv���UX[�x �/Ak���B�tz����S�1p����D�ON�������j�_Bt�snH��/}R�W��E�'*��{5��͊@��5Xck�>�w�x�U|�?
�r�ݏ!l'f�l��<;Ӿ��҄�Q�]2�P�f�\��~��zQ�Pl��M�|���s�:�O�2� SV�DYdg��t��@�����#�'�1��=��1-��U�!a%��IQ��w6~>]��e�h�mpx�m#~�%�_@C�4��UX�]�l�8Utvy	�zm���ܢ�ie��7��)ܿa��ڵ����5���s�y1��PT�w*��a</�R��-0��8�cZ�3p�TW��"of��[�a��>LK��䝯,m(l4��BE���I�\�X�il#5� 3y�{֐Uagk�۶�&� *��:~�?QoO��Tf��W�&)Kp��s�w|���Z��)b=��0��*�&� �Μ\1�gQ!�q��t8��Q���j�����!�q��%*��J=�v�\�G�T�R��ģ���sj��SU��"`!�2���L!�ك�ީ�!���4c�^�U����#�۟�#i"4�8s�<��(A�@�Zd�#fm�h����$�h�ل��}*���}�z��C�W$�����,����6|�~��*����@8�Ｕ@�?Q�M�1Y��E�fēf�p����n[k��\���/�v����Ԇ�Q��K&T/]r��l�1�ǑZ��FU�-nrlH�7�L�N�\[^`y?�n�6�9ρ;�������i4:߶���c��X�V��]�v���D~8��i�/�`k�#�m2./H��=O�I0;�QT���l�1T��uxf��D������"�-k6�wE�#�����4ɡC��{�O���[!~pt�#*),�
��;�ATGJLeK�Zl��`���u��e������
���Ĥ�-q�@������V�355��n2�W�G��҇
�T7ܧ !�L3хd8JȄgN1z�RU�fa龜qo�u�{��։��i�W�_���4�2��;�*4ݸ�2��� �Db�G���j	�S6%�}H7)�8��]p'��HK�R�^p�󵐧ZD�{~��HR┦��'���8��*�1\#��eQ4t6L��_��[����wM�oJ]WE58Ȋe�/<ZPS㥀�JNukn�ަɤ�nɯ�� ���1��ݿ7����U�$�����-@y31H�J%<�l�hCN�.1m�N� �GY[��UX[]�x����[1�|ɬ���ƅ�����?��c���Z�&�H���R�{5KJ�L'6�'��Ow"4&Z,E��:L�2<&fDޠ{�T>K�vlo�h��Ы�u���)����8��������S������l)�%�e�ޜ��@˔R5,&�!#&�pSA�91��J��k{�]_b�(��p��|������䖨�a*��ʼ4h���I����$����c����yHNQT{.Yx�v,�Id*CA�8J�0~9��snd��_ad�ǅ���ɋ����y4��o��<���PB��W�#&f >5�`~@v�|�	\�V9�k�eHz�tW��ɋf�0ʓQT�"Eبfi�7Z�{~鄇�-����򞷱���> ������Y�5�����t6X����Q,{� �lGn]�.�9K&R�GJڔw��飆ٸ����_���2�����������C�/�����^ �*Š���w<���9�Tcfl1't&8�zUD�:M@C�Ҩsj�WC^dg������
s���֣ʽ7���EB��������/��9��|8
�@	Й[6)iqn �KR,EK�:L��	��ud�^��4Q�`qt���U��{������ǭ��	�Ϳ7�����'��>�\��d�#T�Z5<�( #�uPg.B;>ΐk�5@]VY髆�PRxqt������t�X�[�������`)�������A&��3kW
�q�p�G"	�K.;Ԡ-$�3fv�%��C:��/�����T�c�Z�bU�vy�
~�Ċ"i�-��7��4�A��TŸB���>m�FF�����<�
@vb�eG('*��w2�-3�Q\v�asgh�'�v�G�p
n�:�����3�> �ʥ���W�`��\��{�����Zb�U8Kjb&)�}F��b��/��PS��h_q�lnq�ơ�k�������.�����1��$ ��X�0��[��9v8^��y��K.m`�Z=�o�iLs~��[�=@C�֐s���߂dgj�������L����$���3-�S���KE�W���#c] ����;�f ��!�	�k��H�*-0��=O�-�iNQ�f�(Kܫlo�=`����Ru�Ֆ�'g�ꫮ<|����Q��"��+k-�Ҵ*���H#r���>� #&(725��b�DGJ5@[VY��hknYXz}�	���}p���13�M��������UW�a���Š���y;m��V1x��!�qL��<7:ʌg�1�WRU姂�M�jmp���}�Ѭ�v2������9��ѠN;��T��#c +2r,6A�;AP�J-4_�Y<Wn�pKr�t69�*ƉKN�?Ԟ`c�����]f�~�Ӯ�x��,����Թ��G	������b$�������}?�

�Z5T�% #�uP_.?;>̒[�N���ak�Abgj��w�����Sꖨ(�����)��u��R��S��m'
<�g��G"Q|�܏l�fI\{�uXg�ʄg��ٛv}@*�ad�2U8�vyGjFȋ�� ���9���2���T��D���o1�V����L'�h)�"#�2�|WN!�!AD՗ra<�a]`�q��� ]�@���yw�������)���y������ҙ�³����T�Z�`�}�,�/�r$6���|_ZCDF_��Tf�]_b������v��҄���䖨$�����--��-'������(��J�s-BH�с�{�-[F,! '*1�+�ʄgZ�԰Se�C'cdg�1|rꝌ��i䘪*�Ƕ�(����{R�*�&��$1������I��N�h	@ס`�i#�M~36�<CBE՘JڙSB�Bbe2/�;�������=�V�Y_"ɰ�9�
,��v������h���m��v��C&�݂H#�ڝd�F�)��P�^�/\��t[�b��c�(�a\�'{h��|�Ja�k�k��1�1�(��|���N��%b&�˖`��}9��]���Y�ܓ.u'@��5G��DC�̲[Rؾc^�'��Y�_
y|
􊍐�^	���=����͗��J�=����Q e�\����lede�T�e0
r%7��8i�|xPy�^p�g�lƥy�fd����S�!������A<����1�������1���#�{��D��Ob��Iz%>3E�3A�fԏ9���M��b�g�^�u��tˁMo�V���l1ë8���O9��	F�S�<>n�D���i��2�^#I��1����87��,�*A�;^����RLĤmp ԁJj�����Z(l��5��>��GܯXF��cU ��β��JMG���g	���p!ux��/�B!��BE��ri<$]`����:ZW�{~So����!ެ(��q�ѴB�N�&���+�O�o�T��)��P�˃��"N,��72��,�GC�R���ze�kZMPnnq_���~͗�}�����(�,�~��S�$(a�-�X���J�����
�Y&i�_!:�{/A�/ǃB��I�7�(X[�%p��}�r����mOe����>����0��O�,.0�.g�3p� ���P7lzos}B���q��(~�=�)n�r�*7�KN�S�!��m��4W�zx{	y�����$k(硐<J��D��N��F�X��k,��L��OR�t����������삙2�)#tUDGI�TRk��`r�+��]�������k�&�l�����0���;��E��eZ�p� '�p���)���
I�#�of&�w�>t�;GŇܟM@��ad��n� �qd�]����^����毲@�A��T� �6M��o2��T����
�Pq�a% ��!$��r8���KB�T%�XjE�_eh�W�]wz�JJ����'�-�1�;��Gī�=��U��2k/���a��U��]�	ax~�G(+�����ɵhS�8O�Y\�a�gߒ�\j|ʭ�V��^�,�*��
A�G&PY($b9=i(����3ÇN��_�p(��"%(f�@��:=@~X��RUX��]t�jmy|�܏���a��������A���1�V�լe%�p-�Y�8z�	�Äe�\�mI�|��#a
?˚8��ڡS��2�]Z�g� �w�Aݎ� ��'��2�9�?��K �S��]+�c��$(+p�t�R�W�P
Ucp���*�i��6H:@�OI$O�bX3�&q��74s랁�������d#a�Fk8qu��J�F�_���d_I���9�t^����	"�c)Oߥ�*-09�CvŷEHK�S�!��P�i�r�{�����v�`��(�n���@��P6��O�D��O�j/���������Nmo�,�uH+��!�|Ag��L~M<V�R�)�e�}���|~?����_����0v�����E�Nђ���c!�@B���s�J�K&��^A$�*)��#�>���R�25RU܂_��lk��7{ӳyݼ^z��Ӿ�1�-��+����K��I�][�,����t�A����p4���-6�<�&w.N��Na�e"Fkm>[F��r���eSW"��.�!���
���;� ��W�j)�u�*k��0ٔS�A�aY�8��wCq��B�DԽaߎ�d�+�o�qH���I����o*��p7�+���Q�
�^F�R�4�x61��my[�]:X嬔=�2�4�ǯdF�O&���"��T���= �y	�~��Z�a^#s��|yJ7�SH��a #j�-�d�y�p���ik���@#!V'@��5G1[�PO��D�BY�Sv�o�����������������z
���8�� ���Q-��j�_��h�	e��d?&	x%),����!�UH�N9�Y\#�m�o����	�L�@�ߺ��yA��9�ػ|��Q� �J�h#��\��e�F��0����E�m&).1�}CLG�L�w^�M�",n?�r� ��	ɎғzI{��,jl��A�MK������07nc�o�5{�,��#�v�f��>�'U�q�6h�Z�Ex�\���Z��Р0��B>��̓���"h��@��1o;��/�L	�M����������׺���g^����O$=�i#"136�%~���4j`�Z[]`�u�oru�č���|�6�
} ��==�����ޤ ��c�c�Xhm��~| ���PA�%\N�-hn�6�ƋI�PK�OT�Z�d�-j�o$|@e�����ڔ�,*î��=��EE����Y���A��2[�o-�i
��%
��r)+.0�c>=@,�JLOV�!Fh�gj��o_�}��������S�1o��D�OM����`�hh���|�ߊd �G�$��?"!$�2�1359%+BEHJ�}XWZFAcfi�� >��4�o.ɐ��������a��L���L�WU������j�Jd�y�)tz���Bx�<'&)��/���]HGJ���P��h�+P��qtbʌ>�	���aȰb���n���N���ʹ�^�e���L��2-�v��� 
��6�`%�:��X;:=�KJyNR@^Z�hgj���zy|�@������o')�#�B>����Rғ�������k���w�W���!�`
�$),/�Z=;pAZ؛Oa[Z\�b{Y�p�8�o�
��� �{���.���"������'��^]��b�]��2��ZJ/er$6�:.��<;��5ҐU���A��be�v��Ρ��
՚"��'�l��	A�G�Ͱ����'e��R����f �4 SZ ��w�#"�i?�("�pCF֚W:��[^�$�}���ˤԱ]�`��ʹ:�8޻A'�ǲ̒��d�=���Aye�Q��mb��wy�%$�3`�J:�9b�M�HZ�Z�HP�j��s��������������'��q�z�}�Q�O��(.f�f�>^�pq�p�Rs�c':�#&!025ň6)vJMӐR�]ob���vY�z}C���Z}Pq��/o���|q"��-|1��]��%���.?���Fo�s#~{ 2X~.1�D6�AS��Pb� �_qL��mp��uĀ��d��O�����������	��W�#'C�I��Q�G�r[]�Q�b���$'����i<?ϒ03�JSV�a�dv��WZ��{~�o��s�&��2�e�������R��c��.��=}@��)�X���p�('14ň&)8?ILۙn�Ԥ�ij�m�x�
�[��������+��7���, ��P�����*j-��\��E���	�]���!^^-���j<�Oӎ$���&C#cf�5X�tx{�Ҁsʻ����0�*����?�C�5�2��i,��lX��<�M�H�Y�Te�`��$�+=��F<?�	T�9ЈZ]��aT`�ux�Yl���� �y�ʚ��8���ڲ��N�Y�%��H��t7������O���_%����72��'������Tf�����d��x �u��Έ�┚t������`��U�!�L���6���g��bR�Rrt�߇B�);-�X?"�jCFԐsV\[饈k������������(g.qc,���;۾D��M��V��&d�d��	��������Ռ.�eH3�4��f=<?�H{�<V���%ji��^�\s�m@�����혱����H��PJ����(C�����\E�	/�U�����s,��-),[�8;�S�TPS>�_b�jj���x��̂�����晫�����õ����)��3�yT���c����Z%l�f1|�r=��~I���U���a���m�ORU����dgj���y|!���� 6�0���5K�I���J`�b���_u {���t�������*�H�jՌb��4�78L��CX�<ޠ{�#��ujTt�uxdl���r���\�'�����~��أY�̷����=[ @X�H�g�\	���t�.b(m�_M�Z��=�Tf�P�cu�9V��wzܧ�܋�ř�)o�������-���<.��n��
_������ʁf��'z&8��:�:=��j�LOR�@J:`c��l��D�׃�pcڑ�$&�H����*��������N�D�)C�G=��y�ܼi� V�t�e�Cv"4���69��fMIKN�<�o]`��h��@ݰ��l֍� "������ң��
%��W��PG��45Ϗ��OIdKZ���z��C��PK358����GRMPRk��`r��uwz���ފ�`}�瞡���ݱ�*�)�-,#��_�� O��v8�z%�7C*�C)+��%(+i,�\���DV֘s�=�^a��� �g«��ݸ����J<߳�C�v�t����`b�����q/�����S}0+��<�!$w�936� K�Ҕor9N|Z]��!lor]�o}�������ȓ�����I���L8��ˎ�'��5�X�kG���y4��5�p�rMP�i8;�@t���WiD��eh���<wz}hby���	�ם����5s*��6�V�9H/����1��|v���T� olO��c�2D-�@C��pGRUXC�Tcf��Kvy|�jy8�����(n"�����NP���ӾF���r,BA�;QP�.knk�Ex�����7I$�EH�M�x��+��j|W�x{fذ���� "������{ϱ�
��K�.e$��A%��qs������@(-A'�,s�'�Ї3E�	&��GJ�ݗz���0M-cmp�j�Qn����Gv�� 7����� ��R��!a�)0M�:?xN(�4�cf�����!Xf�x[RƜgV�c��Y�N�q䥦�{�^����ϲ�۾�#���0&����E%���S���`_����*�*��b-�L��K1�+�h�UļKCEH��iV΁pbڍ�n晜zNH��Ѵ����7Ҧ�'z���2���T�:�O��X�x��j�v),
^[>+f�$9�j�\IM�gIJMٯzmEydeh�����bz惆�۶ɀ������'$M�0{&�俸C��q5y��W��L�nIT'36��d+FIL7�FWZ����6�,�w�d&腈ڵ�$�\�����+m����Q��o���ln	�����Z���Z}0C*�l1��}�?�5�`w*}cKN�cEt���ي��c4����[~`{��0���8����DDѴ����i����T�Z�^�N m�c!�[>mp��M /25�#��DG��;�\_��+nqt_\m���������TU��6zŤ=���5�$�K�%Ȁ���r�`kV�V1t��~��L�.14��ʄgv���vAX[^���� �������ڵ�TƠ�1q�b۵�I�������f(�}������ �h���B$'*�#58��f5HKN9�GY\��T�btw㎨�����䗩)���Ҟ��D�����_!�������2�l����I,PX@gY-?�`�GF�wK]Q;�\_�(��{��b]}�Nq�⒕ ���������D0�� �?ӹK���k/
�'�f��~1 ���{�"+.1m�^Q�Z�)�SR��r�j𮑄^������ʙս�֪�$�@���ZO���Y��[�e�D�	+K�J>&(?%��mHo~25ƈcb-�:MP�tv�asu�rhqt>������u+ߖ����z�t
�7���C���A���r.����Q��M�ѝ�,Ah.8]2��}CɆL�K��]\���a�6p�g����Xt͖�������'��G������\��<>���Az�FN�3ITdz��f&�(�s-��ǂ<�E�N�YW1�`y�n�r�{�~��+ޒ�����
����}��R�X���w ��8�b ���H�	j�mqu�a�z.@�Z�|��D�>�Jf�`cf�'ssux��
��aPܝ�����3q=��1�ȣT�^�R7<��u�?s#X]
�Ԡ`1�9��D/�59;>�͵fL'��׮�r�4��Є���ߑl#�&d����A��D�9�ͨ_�b�W�9��};��uW	�Y6�ܓ%u'�0j�(]ΔQ�V�b�e��tǌ�֗�]��� i�7�@��� =�'�Z����[��u����h/	�PY�}�a�03��<@BE��RRTW�hdfi�~vx{1����C����+U����=g���Q����.�Q�md��c��y����3�]!�+��8���`�7��j�5)�VY�Oa�lS��tw��	
����m�%���ڠ������QR����e��[�Cׁ���W4�fhhm֡�4 "%�g�2D�"��CF��fTs_adO�ps�a�Q���v]�g#<����5Nζ��I R� \]����p+'y5+S��#	�WӫN"4w��t�8;��MIKN���z\p�&ކ�����	Ll�0���\.�-p��^���BH��-���'`�^��eӒ���LP�C&%Xs2�u'9�/e+~��CC\��QcU�d�Z�/���vwy��Շ�󶩘 ^�-%��4�G��P�V�Z���U���0A�^�B%q�T7*is7�z,>���?�B1��NQTײ]v��k}�3�d	æ������&Ǿ����%�N��:�>����<q_�.O��km��u�&!y�~����5�LDJc5�Xj�P�\�w��}�c�ބ�u�ٕԬ�3�;�������� Y�b�.ɨ���F�-�y�Y�.�d"��/�n$�9o;&(�GJڝK>FF^a�s��=9~}�rџ����.񛒚��F��=�[���<��q��`���K	T�i�f�'*�~(�'?BюT�g��h��^��||���Շ�r╧]�)q�������UA��-d��������T����lQ�#4'*�0769;T��I[�����O�Md���|c]���}�����0t�#�����N��Y���c����u$s����
�
e�����>*��PK�B��M8LX[�0M��nq�_1L����[�&��g�ϭ��D�D�9�NF��Kݍ���E}���xZ���u�H%��21����,��֑G�T�c]vظk}��n�d*H���WT���.��lv����J
�S�\��%����b �n!|��3��-���83��(�&=�7r����U�j�_��������:���,���&Z]�����Q���fR c�bG.myQ-I,#�h8B���-t��rwG;ɐlz
8U��w�.�b�1衣ո����� ���(p��¶B�K5V������e�[�wc�?"7�Cd�]9��F��!s96��ȇk��T��e�6��-�j�T�Ѭ�y�!���xN��2��,�I���Q� n,|73%A$'�M0+�8gB9)gl<0�z]X*VȬojQ׻~u`Nn�����̟����C���*ɼ8��̟�J��I���Vt���nX�V����F*8����Z5�� �%�uÁv|�kṙ�_䢛������Eb{����Uj�#a)x��_��>|������\��>~��k�w�g�+�7x{�S�U�*�<!s95">3�KH�T�yh\^ad�ޑ����z~��H���|�`)����r���A�ò�X��/g�+�i0[�P5��Q
��xQa"��p1��t�B�D]۟Rd�Y��iځ��z6Y~���o?���혱'�.r�|��~�����z\��������W�W���	�Vpvzʙ/2�E/�BT���SV��p�o��oy�)���w��)��﫽1t�Ǽ����K��_��[���u����!�� �h��p,>��[JLqFҐsb��nt�k}����Cæ���[۾��	��s���!�ы�<9��e+!�/1x]��G*M�u%�_B1\'*-��f9<�A�HK9Uߛ~q�#ӷ2�u<C?J��Xq�����+t��w'�ɐU�陣��r�n����|xO��SO�/�w�Q�I���c�B�`�O�.U��o�	�+�͘����14��ŋ������$g�F ���ׄ��Z��H�8���f�yU�Ї7jm�fID���Б=@+�LO��L����o��/��	˦�ps�����K,��S]:��3���V��Ym9t/,���r*��0��� !_��7��6�9>}�N�<8�^o1K	�p��;�D���r�V!���-��6��,��Ƌ��'`�^�A7=AW4QL,׌G�[[��Pణ�ڵ�D��Ή3�ڕ�����behs���v�	�*܋��晫#a��
�'ٸ1��:���%���U�qP@����v��@�rtt��j$���^E(؜ILږy\ba��V�Tk�eȁ������蛭�0�ͼ�m����ÝU
,$��DkC��x2G�ԍ�*!e�_B5t&?��4F�4>ˉlW�~m��e?��y{~�ˮ���m&�ò�����GA������I����88��u�k��s& ^b'y{{��!�:�M�82T�SV�T^�t�v�9�{�h�މ�z� �)�1�k8���~��S�/1���5n�?C�g	��N�;��hlu!�4��0�?"H#BEԑW���naq��ꌸ���Ĕ�Ф�$c��oue�~L�X-�	�2jW�q8�|A}��Z�����%�i7��i9��L�QҞO�[�_��"g�o�c���=������	�%�(����q�0�M��C�[���Y�x.�n
��(��f�$"-(A��6Hƃ=ǬRM��^Yk�-ehk�y�̂�[�>���)�'���4T�����?�W�
��Y�vJ�+ l>��E��v(�0`�>�-7Z=@�N�V؞�\Zd�o�-��~������ٕ�Ӷ+ ���5v���3�R��H�Z����^�|��F�	<�H�,�8�s+cF�;v��C}L�?ٮ`�i�!�v�eo�ux������$ᛡ�6������L����Z�799����B{�L�qz 
�%�*�/��.1��C�X�:L�W>f�_bMJmp�����F�������­�����>������"YM��e�k�o�y6�E�I�Z
�Z"i�m.�~.1�~NƆW���YX梅h��^��z�����Lߘ�n���+�@��L��� ��i-��p6���Hd�P��a���.�#�C�v;�?��D~3jTW�\u�j|�6���@��I���������6���
��M�RǺ����da��a`�k�L������b�k�t&�4Ƌ9ϼ:��aU��S�^���bz|���#	��l�u�zB�H!�Q"�ZC�]��f��o�x�{Շ���db���m�~,�>E@ΓQٔ:�@�ad��UXVx{
Ǎ���ZV��(�1�7�ֹC�����X�V��_���AEnG�v~�E	�Y�ə' !$�h-�qÆ0'Z[HKه��T�NZ$nq�w�	�x�rA���$�%i�8�}�������_"��������{@�a�Q�2c�_%���0/��$�"9�3bNPS��髆q.���t_*���D�����%������E��>|�GP���	���di���EA�j�	��76�f��LK�O��^Q?�j]4A�UX���l�h��x�ԯ�y���-����<��ȣ����W��J���+h)�f�_�O�M0+b�d?2	9*-/cÅ`O*�,JMޠ{rE�BehWt8���~�Iً���������3q)�"]"��V��!����\�z<�U��W2���k1�������0���`;�\_�[�1��~�Ehpf���"ڞ����8~<����:��V՛ל_�q7�z�*0�4B�H�]�^o�k,��9��%;EHהN���i��8U�7uxE�NK�}{�������:�@�z���!�`&��-0o*�v�A�PJ� ����ۧ'�-��H3�|;�J-NQ��і��G� Cc����u�W�����0t����N��A�"�����=@u�إ����U��|�鄄���@;��0�6]����W�VP�qt�u{n�����$�1�.�A���H-��\!Ϡ"��q.�(7�u��)��iv 2_�{�2D�>�BFH�C���Z^�9��lp�����H�Q���fc.l��:�ټ������E!��д�������I���3]����8a$6��236��Bȭ'N���щ�1�<W߅x{	�؋��������~� ��.����^��� 8���8�I��V	�� J�mp�)y�0�58;��C\Z�Qc�Q[�Mw�stwĠ�ֈ_�m�+���$�<��7����"��_��g����}<c�g����1%(�ri\�9R��GY��hW�j��7�0X,Px{�k0���Ċ��)��:L���;���OP���^�j�c1nS��zw�@�z�Q�Y��J�)��~;��T�Pi�^p�&����w����������9�9z��Q�Y��b�^�g�Kx8�p"��X
#�e*��|�;��1c�G��Ct�S��U��d��F�5�:�= x��z��� ����!�-*A��N���_�`�#cNw4��+:/�L	��["%��T�3���U�Qj�_q�'��|��x�����ݙ���(e��C �K��W�S��\�@\����D��Q��h�fV����3���m�@�FVЬ�[�^�m�q����~�^��%�v�S���?��胉���\�(�3�o$�>�y�i0oH
���j���4�w�:�M���U��N��W��\��� �u�釋�唭# �"������=���\(��9AAH��C�	�� ]ʏ����`B�}�����.�YIՔN��g�d�d~��~������D���؛0���1X���H�L�
H��8�)n�z�� ���%���!$'k�i3�-K�SҼa]��h�mc&i4�㜰k������Y�gڕ�0�'�A�E�Aƽ�b�f�$(8b��*=� {a�%���Q#�4`6�-BLGJ�g��i���|�{��u����<ڊt�#��%	���:�>�� E��A�[�_�!f��b�|�>B�;N�V�M���-�;�2h:R�Z1U�R�Oi��������	�����������J5��-�D��?��W�����)k'�h�	��z+P!�)�#�U'tw$|�@U�C���-�?h$Ht�i�[�l�P�����آ��d�A+���}ڍ�� ��[Gn��6��� ���K�a�;��47:�X�WMSN���v�u�^q4wr�p�u�����(�,����(������ׁߒ��ס���>3���� /L�e���Mj$f{-�R�!?�
HF*p��"�0-����m�]p����e�Z��������/���J��M!a��Z�4�D����9ҏb$��g��+-0���ōJT��V�b���`c�h��v�cD"��M���ß���������j(��܈r��g� ���3����df�lm���uP3�5�?QϘN֠W�d�m�z���<���س�"�c)�ȫ��v���G�Ɋ���H��h$�t<�}5�MN x+�"��+"z��0�O9�TB�YK�^=И^a�r�5�w�oj.1������"���"�=��i��Ʋ����d!�@B���F�}����-_ei���ED�v03�E�/*?lKN�/���q���v�ЃŨ�u�ﺭ'��s�2l���G�G�Q���\����pF�;��-�N��X;6��GJ8��258�Eːk]ڄk�g�����ju����[5���/��0��*�A�8�S��$�S2q5}�#��VW�Y4C���!vy�rUd��(܎ILڞytC.�dg����^R~�̯���#�Ļ3�������P?���^�� �5���(�C)�Q	`c�\?N��wxx36Ĉc^-�~NQ�~�H�<hk�������l�O�� ���z��n<��/�K��<��E��S��\��n����D
b�f���U��h7�N��kr5�vVY�&��v��9\lQ|ʭ�z���,��t%��$}�� �T���^����"i�fb�Y�H+]�&�hCZ�u.1��"�jCF4]�V�� �bt����[(�|�ԯ�yޚ��f��<���>���B���ə�P�o1�q���d������d?N�%�25ƈcj-��NQ�Ά�d󭐣�ğ�O�r��������ۭ�,��E�����Jݡ"����g�H#2������G5)�T���<Nΐkj5d�VY飆������_���հ�zvl��.��ҕ����A6�U����1j,l���2����4^r���hCR�q.1��9�HB�m�Ngq�\nW'w󱔏�	˦�pb�����%4��s�˾�R�VL����L��s.�zg��U�;��</�Z*�QD��]L��EXKN�<}\_�fh���v�¥�ʑ�Z#�������"�ܶ�B�8�T@��,c��ٝ��x6��m �	&8i-S"_�8�<4�_b@Yk�N`�}�GT8gj�������k�Oӱ[�/��2p'���6��Y�_�b�Xݬ'7j�ƌE'�ͅ�Z<�u��O:���+ȾK�Mk�:�Z]�f�6����C������ʽ�%���ƾ�O�X�Y��>����y7�UU�}0|�B-7�,/f���N��YT��I�O~��r�l��Ԓ�x�ۙ���������H���_�+ƽp��=}8�I�t�M�^���>"��j>58ȋ1,BLO�ADR4dg��y�r�h\ʉ�ߍ�zp��2�|xżM�K��T9��06:��{:��C�m�w[�TԬL"(���9Y6�=@����FQ��c��3�,���j�:Yj̋�����-���9�5��>�!>�6�@$���p�������ÓM�r��%�u;��4�e�_OP�_�l�n�pp�5�6}�x�}xw��,��6}�����M�����c�=??����H���8�b����ȆΌ�q?��}1�̉S�֕E��g��[������{�ѧ�ݕ,��6��C������*3��2k�i��BHL�P������f�/.1�6Â4к�K̈́�.��]��bm��r)}
�y���!��ڼ��o����B�9�N�E�$#+d�d��PRR����� ?�beh�E4N�/2�=<��1�/F��V�i�Te�t�u�ႁl@�\�'��g��<�:��Q�Yֽ����q5������f�&��p�&���.1 :n���Аaݘ^�(�JH�kn�B_J���֔wte��)g2�
r��G�E��L�]���06:P��[����Zxt�����!�0d*6�E(�HK�J�WZ�ՙ�j�����{􊄝ޒ��%k+{�	b��:�9�L
�!#��a,��j�j�D�~Me��mm��x�v��t����c˒<3EnTW�S�)���q�F���r [��"ᗍ�1 ��G
ȫO���]���m����{P�@�@��$PU�5p�+.����K��K}��?B�`be觡���|y�����#a�h��7�Cħ����Y�WmA��p1���c`�Z���]�j�{�v�ǂ$�ӎ�R�Yk�IKil�7�DgL����X$l��3���4���(��?�] ��f��R�AY�V��P���)��#�5h�B�<?BҸM�Gc�]`c��m�e���M�וx�b��,��8�}�+R��P�����,/n)�u�@��:��SV�P���g`#&�y#�6:=��FJ�@ǵ�]ɟ�WV/<vy@�����"准Ol��1p'�#�L�����'g"�3s6�������1�T�����l���-0��ǂ,��4�UX�U�O��ps�t�j���Ⴢ&n��6���6���N��F���0Fo2�ӿ�������T�h&	��),��F!�ADӐF���#pc����oSo�͐�!g'w��諮��
E���l���	���=5��L{�TT�X]�z5 mqr���V/2�}C�ΏO2�zSV��o��x����	Ƣѯ�ۻ�,gl��A�?�"-�-��<<��+�,����fQZ%7g,��j�{х6
� �~ԑW��v���4ux�W��:b�X��#��2�:��={2OzX%�六���� ~9�J��V
�W�ے5�t��25�< +Y�,F`TW�e�r�,�z �g?j��VS�!r'��������NA�WC���������~9[�Jf�Yo�u�z}�1�D�/Α?2b�SV�\�]��<YJ�z}Ђ��]z�훞.񟒆|��D� ����V�K�]�Z�=��H��7��c���Xh)�i��[J=�Gy	7��|g]Ո{0tp[�{~E��_|��&n�����/���@���&+��AC���F�}�Y~��e�e'*�u+��
'��HK�P�_�+H�hk��m`�J��ϕ�\X���Z�����V8���CƊ��]�3�3l�j��AD��OTX\;
AF�M�[S�1bx��MT�K�ǖ�E�*�Q��j}>C��w�.��,n�3���?�㪠c��\ ���n* �:��F�ʘ	�؝��)�1+�������:���P�Ne�_��ࣆ�����\잰0����P���K?�R��U��a�V<P�F��F!�I�Y<3n�hKN}��z]p�.�I[�9�7Y\�'r�4W�yx{�Ы�u~���)��Ő�y��D�����_!��������e����?��Z5$�1Z #��5�y\K)T�Gיt��ocehkVz�wz|������
���<��-q������6�U�������p2�״����N����^$~����=4���1v!��WЍ��d�h��p���m�Z���%�8(��:������}��/d�b}�.)O�s�\�I��:����(:��369�>AEH�Mf��[m_�~h���v��̙�X��|�>���0�.Ա7��(��ܷ!���i�B�mi��n��G��!�&�xS:�<ɍhK�5:�VY磆i*sn��c�i��������#������3��B�7���� +bW�7I�.����?Pq
s�X1�t&8�s%�Gǂ0�E�PNg��\n�\f�~o�x򃁚�ݏ�����f��;�h�����%^�*-59�]�y�D��A	����S�u�E�rE�@v�F�؛I<s\_�&�o��_�vi�P���\�ea���6�<�����>��G�����r/�M�����|���vz�U�o�.7P��EW׽p���]oJ��jmȧ{��UѤ�!�'��0�5��ƀ�K��S��`��L���w�F%���}g�jI/�,���j����E�p_:X"Z]#hg��\�Zq�k�����ែڣ�4!�=�C���L�K
^$�g�m�s�y����j~`�b k�eHGz0j69ǌJ�0CrQT䦁pK�1kn��s�Dɏ���{�^����6�<��E�H�>���,2i]�%�n���S�r	2)�� ��5g*�GñB�D�5��VY��jeS���x���b����嗰6�5��6z��or��Y�355���<@wk����Tc�g }I(+��@�ǋL+�mLO��� ed�q�sŠ��Pڵ��٣�4�Ӷw�����G��(a�-0eJ��AGK�7qPs(yR��$�o%���s?B�@��ņ[m�o�h?n�m�}Xw� �)����;贷?}5�Q���W�N�k'� �c�~F�T����)]�s�5�q.�D�<�S��J�b�X�ʽ�l~p�b�C��їY����mj�� ��&�*����;�'��y��Az�x�O�Q��H�a+!U�x&�r:=͈>�ٜB=�S]`�r�X��y|�}pT��$獈*l��:���}��R>��*a�gׇ���MO���R���e�bF#&�-136�Ɍ:-H�MP�V�U�h�iport��΂�������ꝯ/�6���}��K�$��Z��d�j,�s5��K������BdjnMvy����6HȋI,��LO�N�Zn��hkn���
͋n�g���_��.����= ������Y�<k8����#��CF�?"9��Z��J�cFmx����:=�БU4�tUX誅�O2or��K�Q���y<њ���3���=��.���W�&d��G��>~?��"�X3J�x� �sNU��8;��.�KNQ��ěH@hk�9��¥��ژ{�[����3w}�ʥ��� _�i�4��$��= 'R����rkn��͊0BTu>A��בt��%�GF�hk�����Kk1ꌏ��%���/s��z鶹O	��Y�$����q�Ԙ����M�V10����qLC��69ʌgn1�QT�����hz��{^��~��ƌ៩*ܢ���^a������';�7���d���GQ�D'.Y�\��� ux�����:L'�~HK���~��/�Q��ru����Uu�����	�2��֙K���C��="b��1q3����PS�L/.��g V#&z}�vYp�
�,<MP�!A>�be����\j=|ҭ�w|X��+��ǒ�s��L�0w,��aX��q�'�H�E�C	f��!iL;�0�[N��GY4��TW���t��u�rꝐƩ��v;T����.rx�Š^���Z�d�/�P��~8BM���;l$-2$'e�>�lȲIѻV��@?]`c�Ӫ����¥�o/e��!�����	��A�騧@��
�^��V
=AU�Q�	�K&1�׈R�dG:�:�~YX#QvDG�֔wj���.��o�\��}���P�	��+�����\���I��V��m6��m/
��&����v0�N1$>�is�fI`{�}Xc"�BEH�s���I5.il����dD����ػ�(l�(௲	H�R��D
��j��F8��C%�r�ei}�y1�sNYG�8;zT�PMPS䦁�K�+kn����f�F�����)�l	����3����R��b%��nJ�������^``��k���oJ1��f=G�D�wF5R�b]�ꮉt�o�\;5|F�wY��]���2�0��F�R��Eۡ"������MJ����	�I�9�5�=14����L�4�TWF`�$��q�<9�ki�z)�����0�������|����#]���
|��A�e�PSvk�a<'3�'*�tW>�ɋf]0XAPS䦁hK�*kn�Q�|�Ы�u�ɖ�)�ƭ�8���G	�߮.���`�h*D8:�SG��N)$���(��oJ1:�47n=�BF��tw�Հ��጗���	����۶���ԡ���:���D������^ �����y;��¾ �N1pcl1ss&8���9R��GY��v]g�a#�u�3�z�Ω�s@Ɣ����6���\��O��9�C'� �x�����6A�_BE�sN]�7�$�tEHؒup�Y�h𪍼�܁��iG*��W��)����8���G�'V�%eU4t6$�L������Z��h%(��v1:=ΐk�5PUX髆�Pb-psơ�ktH���ˆ�c��:�����~��U�	�����p2׼����M(+�ژ�hC6��-0�|B���+��Q�|g�RcێyX�Ix{�K��׬�/^*dk�����3�GG�����d\�����������)�,�;,0�6��<��7��S�n�Y�y��Z˩{~�چ��b���+���9�����WC��/,i�����~��2��ޑ�X�9�+-L�6n�I��H���:��"�$ih���e�y������ �S#|�5x�����sl��*_�]��-$j�n�SZ\�Y������"%��RA4��adC���؞y��m�'ߊ����{�ԯ��!�A������-��F�W��r���,
�h}a$��3���&)(�58;�f}{&וx㹄{e~��s��s}�����Ȓ��*h�<��E�K�O��]�c��������ć�%�+�� ,���dG9*;�)�=�9@�L�tfV�%ӎ�a���p:}�����:����%�V���+�?��A�N��R�]��X�0�3�s?�K��cF8(�'s�N�;��p�F��z�Z�adgߊ6���|{������ ����'�~����GF����]X����_�;5	r֖9�!&')Bt�7I���i�KNQ��~�`cf�,�.�{~�/2r#"��̒	�.��:�F4�.��>֞N�M�1a2���F�j�-p��u'9�Ӎ6H�)��IL�KA[�^�d��r�I�|ڇ�t˦���_�����>��|��0�&����ΏB��K�?"IT�����W�3��:�7:�(��HK�ߡ|�F�gj�H��x���y���)��%/s�B���I?��]�)i+5�l���v!Pmb��6q��eHw},�W~��W�-?MPߛ~�믊��3~�$C�����ݏ�'����7w���ִ$Y��^��̧a��~+]N �l/.�c>=qޤ�0����buC�]��z�\_b��km��y����ˑ�,ퟱ1��� �-��KA��ͧW;���*��sqJ���2%(�zU���?Bѽp�ߙ|����mps��|~6������ܢ�5���8��0��B��ST��Tp,J|@Z�>����rͽ���T�Z�h(�;r�C��ӏr�ߣ~�W3]:�1�@�s�Վ��Ș���8��(~��4��ܷE���a%��B����s&=��V$�Y�"�w<���|_R�wK]�zl]n�ikn�z��S��;������2.�8���B�����כ����.��}y����%`������J�3F��ACF��Se��-I�qjm�3��؀���]y����%c�-����;3���S���@�D�=��v��Rj����\���� P(!$��tWZ�B`�i\6Uܔo㡄w�D{�ux{	������$���(�Ʊ��I��W��c����l�k\|:<�	��/���q�j��b58>�����$g d�kn�:q����XP�'���hr��yA�U�>���E�b&n'�y#��6�����W)�[$$tOn��j9��gYI���K�ςu��"2�t����Q�s@���%���3-�?����XJ��[��U\��p4[���!�	v���䴶Q�369�M*�JM���~q�Qs2���yc�:�����$Zs���8��(@.�4�=|�νږ�6���^�AN �T/Z��;fy�%(�{Vy B�@C��qcS��[�����zq�񤯅Ϙ����(檭۸z���
�J'�H���1��/�����p�tX��p,>�yG���I�pρ�t]v��k}����d:��ty���M�-���:j��K�"U�-������s�q��O��TW_vk|U�6�w+=��i�w�����]U�m鴺�������t��Տޔ,������E�F��C�%�P�=���F�����^����?yV�5.G��<N�F���J���g�|�C_x���qM,���&�)��;���<���wk��09;�8q�o��v��q[&ouy�L�;�8J>�h��M_Rؼras�m/����æ�+�ْ�����l��²p@ξ�����Б.���o1����e�	�B�d?> �/�25��̎i`Z�GWWZ����oru�cJ��
I�3����/��ý6����-�12���}T��:Azt����R�T/2�����J�,/2gG��DDG��TfX�az�o��7�Q����T䖨�ɣ�"���;y�C}���$;�?.@��s5�9n��T[��1�l�nILj�36��d�FIL�aں^^a񳎕X�bx{ϥp/�����0������]��D��2�(��f(.�|��;EP��-�h��%��1C���@R��o�QTW�꬇�Q`�ruCf�s���� �ȇ	`��;=�O�������_a�k�������E G��
g~�DS�uPS��:=����q�SVY�쮉�S��sv�9�#���¡t���1�ҕ�ڶ��7�U�$�k���i��W�M��M(K��:�`Cbu�oR���9�A��M_��\n���mps�ȣ�mȯ��_�f�����<���q{��W�#�V���r4V�h����O*I�z�q�!#�N]�Z]$�DG����{]`c�����]F�}�C�-����)��ݷ0쳴���u��V�� ���q3����ioH�[!�����[.�Eſb�DGJ���Wi�G�gj�5���}�հ�z���.0�2����]��4�>"��s��O=���	)�c�%�cF��0~g�9<?�V�L���|�^ad���q��aK/��O������-��͔�&��H
�<�L���c% 7�^���DK�~!�	\�^9<
�#&��T�69<qQ�=KNQ�Xĝ�~Q�qt�;���Է�,����a��=��0���_!��ƁW��z<V�d�bP	wсe�^%�V),Ғ�9K�	LlI�PS��h���knq�|�e����� ��+%�/���V����{��W��3J��y;�=q �V1������L�.14��?B����v�X[^�񳎑X��x{�>�(����$������i�Ω�9��#*c] ����;{=����3�Q0��*-0��]T'ymHKM�xk�لwhx�<mtwd(���ٴ�~�ğ�2����g��JӮ���b%�����z=����U3�&�O�������Ňbq,J�LO�}�G\gjY#\j,|ҭ�w|G��+��ϒ�b��F�ڭ}����g*�˴���B�ĳ�Z(����rH��36Ǌh+��KN�C�뭈0���wa����粤W��
�1��㲵�@~8��A��a��d���v���*��t'�Rb��O#&z��o�;>���UTV�dv��[��ϮY�����
����#�6��)�G������G#��`�U�.%k�o��+�O�"��M\�1�M�;7�F�H?I}Oh�]o�%�s����ck�9�ܚ}�L��.j	xżM������'��W
��?����B%��n�q��#�����l�GY�ܞytC �dgԽ�����~�ڌ����-�������
��F�;�X�Y�S�p���	/L�S�U0+����hKB}�ZM$�eEHؚul?�_b�h���t��ς�J��)�Ƶ���Դ��b���Y�����Q�W�]��gT��DԤ�A@���יB�|_b����tXY#�������s��ρ�I	�蔭�𢴒��p@2��jmpsX��'g!6?�3���_#�u��'@v�5G9�dgE^��Se�誅�O9"orƄƩ��v���*�Ǿ�8_��E�ѬJz��^�;=m�E�C|� �3��Y�nx]���*(;>����F@SV����a��n<�om����������q0n�SxD~�� W���Rek~<	��8
�5$/�p$6��?|s�V�(z
��ZY�r�l#Yd��qk敌���� 2x����?��:�V��- ����/B_��r%������cF-��21��&�$;�5p����\륈����^��~�D@ݏ��ʜ����:���ִN��Į�T���g�\E~@&�'	�S6=h�k-@,/��]d'��GJ��\�)EzHeh�Ӗ�x���Fα�
����q�2zJ��N������W��1N�w1`�L盗
��l*J4�+.�+�����}PS�'j�g�nq��
ħ���z�*��$h��:��ʡ����U��$d3s-B�<2Q�T����
*-��"�KCF֘sr= 	]`񳎕X$x{Ω�s$?���Ԉ`���3rE���L9��ҾV���r5��f�����bdd��o�kq���.�s;�������o^�L�^�X�^�{�r Cc.Ȅ�𘓁�'w-�6�ߖJ����j&��i/�j��C������gii�p�!��14�AȍhO�U�Y�]_�+�-rq�Þ���¿j�U����5���0��D�!H�\S���^qht�jۆJ%�p)�|1����K�wX8:=@�X��[��sIl�.U��d~���s� �����co=�	F����H���)���ww�����.e�$��H+*-�x2l����ׯX�����jil�0�|{~G
�����\ţ��������?}4 �������p����������:��8'&)�3�;>��_NMP�m�&֌�v���~}�˅� �����/u3�9Qֽ���s��V�L��̀���{�������4#"%����@;:=@	�VPORU@�`c�m���@	��� �ۚ"#�������x-�F_�������P'eJ��qV��z<x"�k�� �� #bo5�@�Ŝ>-�*MPݜb�/K��kn�m�z�S̆����*�11µ��E�"����'`�^��g��p�LRV5O�SG�]
)),�@�E=�hS��t_[�@�q�=eh�ԂKv�t�C���!�5��e��-������b�b�W(Q�A��G"��*�Z=,o���03ĆaP+��KN��rI�il�����
Mm�h��!㾭�2Q��:���>��8�A�J�$S�-]*V5S�
�kFh�(�W}"46�h�7I'D�u�L^ޠ{nẼfi�����Ii~c��ߺ���M��
<wE��T� %+/d+����~k�͍�;
����m�3+�47ȂYd��8�X[��m�F���~
�s��
�������/u�>3��D�M�S�[���T�"�a�}��K��"]a'[�0��:�>D@����\[��P�V�����
s��]yD���-��7}��L��Y���&f!�2p��fv��J����b��#&�z��;>�FՐ:��&Bm�be��s�w�}��؋���w��/���^��B�7�3�\�(f��
l��@~����X��(��ꅇ��65��*�ϼR�;8[^�f�kn�B>��� ��t*��(������+Ż����[࿬�������}�VX��^:@�	���[k@�>��Wsv����S��p�QW&i���ե�Kp���Z�ݜ�ܳ&�C�+�R���K��a�;av4/=r#ƒR+|�� q#�J,ES�:L�Ύk�Y�Y�#�&,��� ƛ��Х�S�\�*�/�6�B�C��=��Y��r�q,�=Xq\�|P�Z
#uf*z�'&�xS6D��j��`�k�9<�"��3�Z�<�A�F�LRV�d'�-�6��yG��V�\"�1hY�s�?ڝ����J�Mf�@3%�xg36�L����]X���]�i�t�6d��ḿ��W�����:z�,���8�޵�v��g����D|��2^���km�!p�#�>�uC5�D>�IG�ZP�_B0be��w�7�{}���N�{F��/�̯��\����T� #+/f[�o��#{��6����5+b�T�4�h7a�?�MHOJ��b֕d�ւ����l_À�΄�d�<w��4����]��J�$&���Կ�����)����
���b���<#"%{��=��źHƫQL�Q�b����Ӡf��Y�	���n��U�Ҁ�����Ⱥӥ��R�G�c �!�2&��n5<Vz.H��6��" W�o���7>A�G`J�Ug�!l��Ignq`}�A��rj���᧍���1�/EK�(**�����M���B{�y�RX\�"��5��(�;��:=��%�[ޣa�GR}hkY��Će�]��ܢݧ��~��8~>������X�]�Ŧ���wd m�N��K`����j �.4yCe0�F	���B��_�d'�R�Oru�{���{�v�s��(�)m�<���:���W��X��m*�JLL���U��Z]ei�#��d-0�.8��A�P؛I<�u]`���mG�i����b~���2����Z���5�Sķ���iW�8;z5��L����` �s!>�47&N̒K�VO�b�h J�jm��@<��ʭ�Z��5��l���9��,��?����r-��s0�!(�;�!���k��A[�v0�5Ɉ:���Se��E��n����oI�p7���^߉����:���+/�����L,I��=�w6��o�x���]i�-�o-��(369ǯVH�C��`Z�Y��y_��8�`i䆐��!L���� �42ú1N���%�0�f��n�����A�X����P ��g,�4�/���i��PSVY\_��pn�m�7|h�����������,j!^��B�ٳpY�t����X�ti�p,~<x5�[��!��;+�*@�{�C��,L?RU�6�j�fympv8z�af���y^ܖ���1�Բ��"�(��<�̠��7D�b��U��i��R�6ƒQs�]��-�-}��kǄ>������S�bhknqh��D�v|��&��5=��7�H�3�\��m���j��e�1�q	�R���*fy%�4�) �jADԗA8Z�X[�m�40ut�i�녌���#����G�,�U�!*����i�fzmH�v]	���\��^-��|6��+[]LO��u�o�9�6���������]�����@��0܎��2j�5R��'��N�Ɂ�� L*��10�z]@ʒMӋR��?��`c(ml���|z�i�/��R����������w'�N���v��cR�f�[��˓���v
������~��0���C�K��Wić�fxj�y�������J������Bǹ�M��R���d�Ⱥ���z7���[�`��\!\vbuK�03E�QE�p[�aC9cf��x �z	˦�іy09��+jn��C�V��׵�qc����л��PHv�a�^���d!w�Gu�4F��>�M�FUTWZ\3�&x�grux��Ո���������0n&�~������YT����.I�N���VJ����S��l02��,/2��?Q��.KOR�X3�"t��nqt�d���܎iX$a����)²Dz����E4�_�����yt����r|�#�(o
m'*-��G%z�q�I�Ng)�\n�$ۘ��r�{�n։�Q���0+a���C �����),>������?����Y�-oo"4��<��58;>�AG`��Ug�\3���52� d������{����Հ�n%�@�F�O!�X���g>�� x=��$���>I,�[�m�r4jA�qȖLJ�`�{�t�h�k2�y�BM�����c�ټ�8����d��S�	�O�k(�HJJ�� ��u(�zrO�':������/��դNޥS�\�i�e�9��	Z���j�*ᢑ�ur@��������V��i-�C�j���>!Y������,q�u.�E69��LKщT��Nԇ�3Ws�ECf�솉P�֦�3m�w���K�,R�0�-f�d��m�I�E ���
�v�rM8��7:=�hO�Le��ZlG��gj��|�zpk�\��������0t��;���!݈�'g!�NMM�E��� ��`�b=(��'*�}XG"��BE��[RʂZ҅lOBkor�9�����yWe���.�6�Ӻ�HZ��O�(X�0�C�I��]��]������L���ؙ�q#�.,�WF!z�AD�Z<��I�G^�X�sux����u�,��'w'���q�G����� ������W���2�w�O2Ad/	q$6��K�8:�eX�J�QRkŭ`r�g���u��mǪ���z���&dp ��
��G��`�//b�:�n.�q�f�{
�̈́A��R��{���4�~aT��B4�TW�҅t�j�>�Na�"����e�������6��L��^/��577���=v�t��{�	_ei�\?Fq�))B��7I�\��I[�Xj�_��mqH�;���㎠Lɝ��K���E*��K���< ��ۢ.��{;� &�292d�k/�p$6�D_3E�GnBTЇY�TfXq˲fx�m�@�{�������8�˟�"�5�h=�첪�M����d��g�^�6-2+�����b&L�nIDC47�<�gbH�d��^ad�����u�Ω�sH���%e����<��أL^��U��`�V�$cA^��A$'V�X3*�c� #WW�2�]P>���ޠ{jE�rfi���u����ֱ�{�3�����;��ˢ#b��V��x���[��H�����^|��]8'6�"%(�SJv7=@���lZZ\_�򴏊Y �y|ւ����������l.�Ϫ�j��^ ��Ÿ��KMM��X�R{.�W:)�(
l�*-�x[B�KF���v]���n��ec��>���w��"���1���'�C�d��ݸ�_��b��E��J��T���3*�l1{�*,�WN�B>�i`�N�TVo��dv���vt��ς��S�U��'���̯p��E�C��L�]"�^B��=CG[�K��Bbe�_)��v2=25 �oAD�
؅˧Zl��t�oqt�
͏no������d�3=���C���R׶v���G�K�;��A;�]�	���xC6��3a�Ćat�.�YOR��_qcێ�oI�9�����T��*��ґ2��� {!���>��Ҭ^�S)p�U�Lw�M�O*-�t��%7)�TW5���k�R�`��e�𲍈W��x{�I爚����r$bk����)����ǿ��F�e'�g��������y�Z54��:�(+%�7�Gˍho�0M;\�[^X(i�w����ex������h�˾��������I"V�K�E�5��y;)���W�W:Il��'*�}Xg"��BE�S�V-�誅�OypsƄƩ��v�`��*��Α@I������CvX�c 2�0���DM�#��^9H��#&����8;�*{�JM��~�H� hk��}�@Ђ����fV���3z�S��JϮ�f��b%��~��x�RTT��_�]�����	|v|\"h�A��ʠkn�U��i�e��t�はU�蓭�����霮��H9��<*��H6��B��Uh$�S�K���v-o�_#Ϲd 2�-03zF����Մ��Yk�Ո���x[TS{~Pp47���Ɲ�����:�������;�PI��M�5�_���u�k����Ռ"���V-0��;>��X�Lژ{��kｐ�����DŨ̊�W׺�ؠ�)����5�����B��D޽���=�W �����=�ah�&����+.�%ÁFʈk��PR�a[�fM߾mp����G�г�}�/���;����k��2��H�����]3�k �t� m��1�7�iLg~�B?BƆ��SeX�|��o�����͆��s�ޔ���+���B��@�F�O�5 H��,0m���E��2@tn�-Oo"4Z �158$Y�DG�NYTW穄�N�nq ���k����Ǖ�ӊ-s��<�<��OO���7������8��������F)@��5\��AlA},/�r��?QD���[�΋즉�Ն�\��}���|؝#�	��� AĤ!��Vƹgl�����w�Z%m��k�N1Pc�]s!� f,@��9<?�.LLOQj��_qM3glo�Š�j������(���qi���qB�;�0���Y��H���z7S6A�gBI��.}D�8;ʶit�T���~�S�ݐ�ZP�{~ɛ���Y
��U��4�<��
����Q����f"8".,{ ��>|/n �* �6�14s��QF�q��An�ad�[�혧���	Pt�U����|��A�?��/ȳl�����P4��'kU�?"��.�q�e@MqL;�w8:~aPv�LO���f�IW0il�3���� ����╧#�Ŀ1��ϳ��˩�.���$����R6��55���	�Y<+YeH��ϻ>�:$b/DG֒u�⦁�r1}�s�w��Ep��������6Ѵ�=��FB�0�F.B��W��`�ؑF����AO2u�Z�iDK�mPW�9K&��FI6�PUX�z�C�r�<\s�}�ҭ�Vֹ�o�����=���y��][��\�\�ȷn,�m'�w�/s}���o�{� ��36řdg�@�j�0�b�,L�mp �FƩ�_撤�,��1o@�����>�����W3���v������d�il�f0z�u1�E�lN F�3�ڙc�fZ�uâq�fܿ
ҌW��]�����}�`���b'��X��]�N�B�^�Dt�]�V _gl�(3���}3�	0b��Bl�Cdhkn-FΏ9F����������;��>��?��$&&��*bN�:q�w痚�Z\��E�"@#"%�3�B37�<�oJIL��D�BY�S���{���g�O�������0����?ģ����U�����l.	 v��t����g*��*��&'*�3��]L�F�ؚux?�c`c󵐇Z�Bz}Ы�u陖�_��5��͜�&��N:���U��e����z�4��+"Af�Z5(�\�`�f���,�OɆX�
K�#�e�X��o��uw����۶��;С�4���C�۪`���^ ���<|6<c*ZZ����.u�wRM��<?Вm�7�WZ�ᠥj|��ux{h����ݸ��G���4�=���M����[O��iQ�h��!�y�x�?)���XV��#,��Å`W*�MKN�D�e꬇~Q�truk��ʔ����('��,�P
�_!���,���x=�F����W2Y�6�y�mP��_^)/�ILO�㥀{J� jm����h������"ܿ��1��ј�F��J�U�$�n���s5�ʊ��W�K.i`�b=<ã'*-a��^Y(+�HKܞy�C�cf����^/��
H��ٯ�*��
����lh��U�V��,����{=W�z��X3*��!��9��158'�͒Pؒul�Bp$be�����w�o��ֱ�����5��A��)(����&��l1�m��C�ؿ��T/v�4��f.qesVE�GɎLԏe�;[^ﱌ�Vrvy
̧�q� ����±/�ν����H5���V���1��3˕`��K�E�ҕ	�]+��!�m3�������!���}�Q�f�/iX�����������]�,̯�~�?	8�U�[���:��O�Dr<Dk�Î��m�w�ow�?���$ӠEH�9�bZ]Ke�)���8�jp�����"�Հ�����B�I�Rú9���l1�s2��O���z��d�&�e�t.1�0�=@��ՒHޣE}�B�c��l �U	�bg����9���p	'�B�H�Q#�\�d�0n�ri�ڏ����I�	�$[cv!�4���9<�;�HK��3�m`��uX:{y|hL����|c��1��B��-�� ���k*�t3r`�B�KGT*�v�Q$��3[xB���Z�Ӑ>�TZ�i��Qo6�]KC}�K���ۥ����6�,��������`����e�p5��q��
S%�\&�e7al4���}i�P��SS�b��Jh/�V�<vy D�Tt�����g��; �F������a$�żr��w4�TVV���Q4�Z0�&%{���-'�?B�9��Qj�_q��B��[�A{~I���W�]��C���=�;��.��B�`�,�0���y��`����S����������43��(�.Q����L⹅�f�_��z��w��z�ڎ��b�*i0{���$�G@��$�R�J ad��@0:�yq�A�ޥ�k�),��) ��@CҏU�[Y�P豝�r��o}>��Ș�������(��pp���P�V��\3���*�`�<Hsn	c����{"%��*'9<+Ey	����^I	ijm3�����������#ۦ���B?ӿ��J�D��	����DD[�>!��9b��si#&��;��
'��GJ�9��Y\���,�p�5��D����Zd�Ǥ'��t
B�B�Q�@�W�L��A���x��Ą���-���M���m7�4�_B@Y7�N`ᝀc��Y�q��~}�n��� ^�`��2k8�8-�B:��?Ӻ�����t0�z�p:	: �D)R&8�;�8J�8D�R�\ƠYkӠ��jmpr�	̀�
H�1ߘ���f�2ҵY;	��/M��>�\��d6��-H��	<"nq[��cΰ~7I���u�XʜUg���_�Yށ���D�X+۔��������9��@�C���+3B�6���?x�v���X^b�
�C��9g��y\G�T��^M�`�X�g�4P�psb�ݏTt�R��(�ż0��ěj{���9���Y�Xk��h�D
�$]��A�fI4{�}XS"��BE֘s^=�]`��h�?�Á	æ��s"���'�Ļ�B8��@��R�*���.g�38>Bw>�߅���~��N�	^�),�zV��*Z�JM��Y�w�e�o�yy����������n�3�t���H�!!����X�R�d �b��G��K&	�����J-+`1J��?Q;eG+]\��Q�W~��wnh:h��ם1T������;���N�7�����m(�9y4�E`4q��nzq'*9�89Rt�GYם^�[C��cf�-�] �w�KG���������/��8��E���UB�^S��l�.�x�~�A�*�{χ'� �����"��@ϊG��GSl�as�h���v��<ƃPM䷚����6�1�E1P�K�@�U�h�����^�{���/�-Fi�m�;V),��A�1�O�2�RU�D;�dg�m~��{��ʹ�������,���s8.��S�*�N�n�l�u[�����	��q�Q��}��/�)t����N�Vg�bt�%9�t��	æ��۝|ޓ����6���wG��N��\]��F�L�>S�T��A$;V�Y�2 T�w9��8;̎ip3��SV�\�d%.�p���S႔r������)����8���������Vۺ7g��n0�}��f j1j�a#��"%��1�9���Ԏq���hG]gjm�Će���۶���'�������*�+��^�-m0��l����+�N���e@G
�*-�3�;�t�GY�;�Vh袅����|[�q{~��ؚya%��-��єF;��H
��"���@�F�J�K����Z��~��o"k�gB5�(,/�z]L�ωl�ޘ{������Z�z}H�UxX��*���D���Sط߷���q4��I����K&-�.��fAP@�+.��\s&R�FIڜwfAd�ad�l�q������ٛz������4��ԛ�G������I%��h����|>���ԏ	�	%�f!$�x:19<͏ja�G:�Z]�񳎉X��x{�]
�	�	��'���6�:���3�D��A�S��P��;��H���_}� HW\�(YX��`>�iXؚu�?e�`c󭐗�ğ�i�A��ߺ���*����&Vv�!�ӄ�0���18q3ش�����z^d�`;:��%(���:��x�K]��㥀����j�������հ�z2����/o�B�����L���^��g)��s��D.�Ԏ	���!� 2O�-��C�>P�Ӎp��=�Q]`c�����^O~�ԯ�y4����3��Ϛ�l��E�T��H��Q�ʳ8��~@�|��[65 �� #�w9��8;ʇM����9�� ���k㖉wl<��ڽ�a���6�4��=�� 6�<�B�i���R?��W�^)
�5$��f'�	.14�G��kfOPRk��`r�񯒋���ħ��L��(��RU�4c���B?��?C\;,��fJ �9Ni�m���`C>&(+.0�Jʄgb�K�VTm߰btf�}�A^v~�	H �������6����+���	��P��a:���HqU��D'Yt�x��%#�B�C�}`[�D�OMfة[m�[e�"��yw��񉌥#蚬������ǥpH!δ�9�b��1�]��wH��dff��q�&S�vy|.�YH#��CFQP���L�a�����������O������/�-�9�������E�A��Sq���F��TW�G7�}�K���14��<�[яd�J�a�ԁ�k��t1�9��EL�_撤�����4�2��; ��U�U�K���3R��������b�5�$�k�l".036! �ADG�^�T�Y�h�4Q�qtki��}�҈�
�)쒍�0��
B��� ��W�13�����[��6K�4��`���j�]�n*</���S&�OGJz|TVY�d"�i{�w$x��IFE��� g�����/m= �.çr�ʹ�+�����s6��������y<�`��!$���3�"�+-�KN:_�Z]�W��@���Հ��cvN���(h����?��PE�Ƒ�����l'�8x3�D���p������q���25Ɓ;�D��STW�\u��j|��U`�8����#�|f癧�������P��G�B�H��\��e��$O���Yׂ�y$6yy�47�MCwI�LRky�`r�+Vr�vy�[�tw��������	�1�������L���6��|7�Hc~Z�Z�����@�03�Ǌ+��KNߢC�cf�� [ �{~�hs0��'�x�@,�����C����Z��b_���Ԡ���P��Z�G��1�6%$'o�258�G*�JM�<��\_�*u��v Gc��S�d�%8��3y��7��H�"$�R��c�:r�(6�tMf[@ɔ\��$\l-�'�{<��'N�Oh�]o�l,Ou��z�	�nwޏ�\�#��5�t�����-���.��h4��o�TV�Y������!"%{���I��}�DV�s�VX[Q�׉�4���D�~����BD�j���Hz�<����x<~�I>�S���!X	��н}.��K�.03������I[�x�[]`��èSJ�Iً�ﺵ%���1��X~>�p��Ɍ4��_����U���#��v'�D�&),�6H�eGJM0�Wi#�)hknU�x�D�N���z���e%�s�����̆F�����<��g
�����]�Ȉ+�/
*-��[�=@C.r_OR޴�p�k}�3<������<?B HJ.���:N9\���,���`"���͈���t2��c		�n9<�bEH�B<���!�Ǟi�Z�VWZ�Hou�qru�c��7���~��#Φ��1���>`���C��L�"n0N�����C&eX�Z50���"�uP�&8;>�ѓn�8zLX[즉������{}��������+-����������RL����0-��{��r����
�	]�_:5��$'��U<8:=(��HK��y�\^aL�lo �Ā��p.��$���
���B��p���]�1,lf	D���D�~!�	\��9!�,/�ý`KCEH��9��Y\�'r�4W .wz�Ы�u�E��)+�������7��MO����ҽ[��qs�����$�W2i�6�*,/�_�)p<ILݗzѬ��<knq��� ��������������C=����!��k��c��t�� ���N�P+&�����F�(+.��9<��j9LOR=�]`��qsva$���ײ	} ����3���f���N�2]W����5uo����M��*%�� t��Ql469��*��JM�c�%H�hk�����f�5���������'��>@���îK��bd������o���H#j��j�fA�\+.�y\����k�NPS�����fhk�� ��~��n�����%�ͥ�� ��M��E��V�����0p2�~�����(W�����LK/14��?B��p�SUXC�cf����a��Ω�sL���'����60Ӯ���NH�*���&fh����֎���M��*�kh��#&��<��!��AD�ؚup?n_b���gruxc�����k�����#��;=؟���� G��_!�+�b��uL/*@�C&)�O25�O,��"(+���|_^�����VAVNad���	twzegڅ���ڠ&j񌈙��@B�T��Ű����\��d����"�-<2�H+*�T7*�`C24��.14jʼgz��}-姂�����svy	��m�(������� ��,��.8�FE�M ���<�};�8}0;*l1L)�T_5N,�CUяrq?p�����;�]�j}�l�͍���"�ö2��ڙ�4��C�AQ��bmiZv�F)�P^A0�2bpSF�>t�ed�dڜwnAd�adg����󞥋�҇����(�ż��)��A-��G�<)Y%��_�T9q5w�lI1���.���ʈе�R�47:����m�ORU����gjm��*� ��p� ���')�3���:��ʴ��Qҵ\O��g���uw��������\��� W牋������1������Y�^����v��P��і�*�2���8w.�J�P���L� �����~;���acc��f���I���&� �BTԖq\;|J[^��l�=Y�ey|C���Oꖨ(�Ÿ�����C���R��!+dK�G��B��� ������r�tO:��9<͏ja4�TW誅�O�orŠ�j*���	�%l�k&���'ͷ/�����B��K��T��S���w��L'��h*	��),�x>���'�
_Nܘ{^�($/t�03>{�?BM��NS�!���(��D��P
��7�4��.��4}��y��2�U�_��lG>D�14øJ,E�YTr�A��ad�+��d�����
�����+�=��;y�K(�����$*g!�6v9���o���P+����8�oRAC�>m�+d�KN���c��QU�������ԯ�y�����3��Úw7��N��\M���&�;�֊����\��k�[�q3��25�,�Q�L��9�Y\�#��\�v���	_������������8��!�JϮe[��`��1�z���w�Rq!�	?�R5 ��A,a�=o>�9W�ƅhW2��RU���J�.�7������ٛz������c���U��L�'E�A�Gp2יh����yBtzO�e@7
��*-���d�d+�KN���q�dfޑ��>x�m������]+���䴷H
�ܯXF��c% ��ja���b����P�wyy�	��90�w=?�fI
ON:jY\�N�mr���҅����i9�䠲�~ֳ�����|������6�^��B{�GLRV�ݓ�Vg�k�(+�"�.JEGJ��oZY\�b��߂��늹���ы�#a�१�����.���M����春c�]8f�{�v�-�!�!"%1�487:=|m��B�NW�"�e�qU��y^�~�8�Uy�P���.t4s����L�R��#���ڪm�������M?1~tW��0�5kt58%�BEH�T9&Y\�+�?�6��tcnX���PZ~TT��0x6|<{�����y�W��|���l9�u�{�����������������:=,����\���)M;�mp�>b�8��Th _�.x��]�;z�t��P�V�\�b��Z���?z�����	�,��>)(+�8pa�I|n�Q��a�Y]`�'���<9�ۦ��s_��]��)��2��1��"� �1�2j��y���;	��V�3�KL �kN5��>9��.�,C�=�XZ]���h���v��mՈ��X��y؃0n%��-���AU�H&���t.[2���R�J@�sv�oJA��z6H#P�CFR�Wi�vcu�>�u��Tˇ��Wږ�������2p�:ƽ���nM�ӕ����<v0.EK�qTu�p)�cFax*��F�@CF֘sb=�]`�����[��{~؄������Ʞf���?�צn���Z��)i#	8x2,GKN�G*-��b�~ �kNi���;>�	T�9
"Y\�+N�nqt�ʥ�o��#�������> ���9��Y���T��t6� o��y,�U8Sj5�v*<��H�=�h[בt��Xq�fx�m�s랕h\��V� �š�������\-�ǳq��-�����KMM��X��H+�� �I4��36ŁdS�X��D�Jq�~���J�
��؂�8X��)�j���y��̔��MM��b1�kb�_tqy"�����߆�%l6,�K�~,�*&�KN��b���R��{r�>�ɓ�[z���%!��4}��J��W�S����a]�3p��7�V�;"ATR_)�����$���5ԗU8k=X[�"�vj��Ŏ|��n
Z��"壆���:�Þ�0��#!(���-1�T�t�z>�/���	`i�@7��L}03���LCяT����_ܣ�oè1��}��S��ԕ�%��1�m����N��O�)\�M�j0���BKG���`$�f+��4��s8�DĐcF�\�M�\^]��R�Pg��ī��
v��X蚬XZ��-��J��.%��6��@Cz4�IM�v)�R50g�n"%��;�� ��@CFz �WiD��dg���|_x��հ�z���	����_Ź����(2��w���f#5��Qok�FHo�(C
�*-d���GF�M���f�c��;X:^x{
����|�!j�&��&���C��O�W�Z�Q�Ap�I���L����Z]�W-��n	�),/�JƁK����9�<Y\_�nQ
Mqt�?�ѓr���&鷊���<��E��T�R��),k&r�=�����w!�"�'�(�j+.��PȋM�V!�TfA��ad���Yt�y|Ȏq�U��&Ű2���>������S������%X�q��|�x�Zu	�<���鄆�213�^IˇjUןZ��_��cێ}X��x{A���v"��`X������ټ9�Ą��OΛ��7p�n��w�PVZ���t�B-$��E0��ĈcNЏ[��Xj�����;q�c�h���׺���ާ��&����S��Z�̳��n0��� k����}#U8#�aD/apD��h�����,�XS�lꮉt�r�_b�l�݈�������Oٲ�D�B��=�Y�?�/��������!�K���1x$�;� �c<?�>H�#��W�f�3O�or�����J�������1�	@��h��2����d��/���f �=R�I�c(�Q�i/)ɝP�38˚DJ%�q�TY�ep��{�B�y�����^ *��ޭ<���*���\��� �j9ۃ��~;'D�����u�0P�o+|*�}C��PM���%"���v�s��������-Ȝ���H:ݱ�C�l����^!��_�U�y��,��#�	f^��w{�x��|5��<?+��KN�[�!�$cێu���x�m)��!㾥�>��:�ټ}��O��&^�d�b��q�>~B��#���m�p��"�C��-��MH��[ߤbE�	ehW�q�Ǣ�l�l��ƕ���#�6�>��
�5�S��"�(`��g��=}?�ܣ�Z5$�8�"md�7�ÈFΈkR�8P7X[쮉pSp�sv��q�T���)���Ѽ@4�G���=���b��D2��w��?M���P+� �������94��)�'>�8{����WzU�ux�ZHɬ��Wػ��f�ʷ�u�����w��+Z��)����x2G�I$�8��d?6	��),���c�̎ih�6_bWZ꤇������`���ֱ�{���%��(��jz��M�������k%:z<
�ڟ�W29�6��!-�UA�|WJ�ѓn�8cY\즉������b0 ��س�}�	���*�ǿ?
���M"�"Y������n��o*�l-�7t`�b=4K�'*��L��aܰ��FK�n�g�vw�|�����_!㾭�>��@{I�!���!)a�3l0��8���H	�H�BҠ���Ϗb103�!M�AD{��ˁ�g���sruˆ����R���+6����=�=~�;����),g�q+{�F�����\�lG6D�14����	RMӐ֤]oa�tj�xv�5ф��O����!墨�$�¡U��K�ڔ_�e)�q�u�}>��F�
b�����5{��^|�;M�v!��7]�WZ�3�납qsv2fW��|�����!e�Ь��l���)��#[�<� ����5F�
e�r�V9.3�v(:�tWJ�L̆i\��Pi��^p�^h��tM�|� �P����*�k��a���K�I�� #?�E�IF��X�S��w�O2%e��!�N�-?��<N�,�%LO��!D=dg�z�\v�|ˑt�W���,�2�2y'������2�Y��n��A�>w�CFKQ�V �W�0fs/�� �s-�p�L���_/��X��l[b;��KH�z���*��ů����9��B����,��j�_�i�J���b(��#&�zH��;>-��փy�Xj�_����f��z������x2����V���5�S�����k&�7�b܀;�LVz 
�	��";Y|0B��Cˆ0�2L-RU�KJj�jm���bz낅٧z����/�yvG�M���A�U�h����c��Q�̈́#� bZ�-���3���DC�7FQ���_qc|��q���į���NR㾡+��2��=�D�O�Vߘ��4m�k��BJ�o������t�Iux���+�:L'�%GJ���Y�h�Ny�nq��Lis!���F��*�j��?������P�L�a���Xx61�Os$� �.�ץ:�s'9�=�{H:r�C���g�K[�rd;����x����Pң�����tצ�+�<��:�,�2ͤ_%�f�q/�z��{��J��Z�Y Z�9�a񏖘 �B�mTNg��\n�\f�|�NŠ�j*�W�]P���� Ӿ@���L�U�%&�P��H����0�C?M0�*�_B%�?Z.@4+;>�E0d�PSf]��R�Pg�a����\x�6��,�ۡ�����B��T����`�h�#+u4u ;\�Go�S��*��_�.A�]@�kVڜwjAgbe�����Ie2��۶������)��F�ޭȪ��a��0n��z���G"�E��c�]@K���,>�)�<?�
U�ܖy|��ew�U8�ux�C��Zv�/��*��ƑD��E��V3��`#�"�u���)��?���V��~�胅���B9�������ul�C�/�ҍ|W�wz	Ƅ�e��ˮ�p���5�?�����T�՘b�^�\�x����諮�E2��,/2��<�:t�O�I��m�X��m�g���v��	��"۠��#���1���;�I�5S=FbEi�Pn�x�x�	q*g�I�+��P�)r�<�D�.H|'���a���iъ�[u�K�=j�r��������~:���L ��������s�v�==@�	��#[�`d�c--��ZQK�dDGJ������%ji���f�����J_Z�m���.�7��@ �����Z�(c���2��@�*�o 竮���,���98��-�ҧU���e���u�a�z��z����t����!���N(���A6�!!Ф\�Q�:<<�������v:��^jllm$'�,2�|F�L������@97`c�`�u�t|����s[j��]���2/��/�b<��U�J�355�t3�<\^^c�g���6����W�0*b�JMܙc�h�A�k�5����Gȫ�����j����t��C�׌���4��]eW�N������>�d~!�D?w��_�I?�&�|GJ�#�Ⰳv�>�r�?�J�ܧ����[����ߢ�;�鸂��S�V��d�3q�Ԗw��K�����b=,��'*������%�QL��F�i�*؅�U!~vy����`|u�������8޻ G-��.�a �8p�&4�rV�W��\$e�a* 9�{.@�.ĂG���~ܢ[�&Ԍ���WOwz	ǌؙ�[�c	����䱴�0���N��U�����Z�T�G�/������su�! x��*�$G�~��K]P���k�#ehk�՘�zC�'���MA���`����0�����Mi���A��m���q�Ki���f]	�O��/+.�M6m�+�'KN�̮뭈wR�ru�	˦�p�̐��"����� ��@������4�8�8��l.	 ����~�tM0��<'!�+�/x4F:ɋfU0��PS�P�n�4Q�Iqt�c�̃��S�Ԝ�'����Q����!!T�,�`�`�Ul�aF���X��<�8c�?X��(�>;��z
�޲}h���Y��y{��haЈ�ؙ�Ÿ�q��%S��J�S�T��9����t2�PP��V����1�cF-x��5Gǉd[.&%NQ� Cj�cf�y��u�䁂����䘪*�Ǯ�L��E�Ѭ^.��`��/JK��~@
�D'���� ���m25�@̎iP��U�WY�_׊}k���y�ͨ�r����&�ê������޼����Z�2�0i�58=CG���X8b�&�!3��.1��K=VX�K]�+D^U%fܪ�����|����┭�*n�5�F�7�0�5���O�0�O���u��k`�o���8�)x�6X������Y埂i�O;'or8}|
Ʃ�ޙמ���cc��t��F��U��W0I�>#�w?�u�f?O�
�^u�b�
/�2Kɍ@RЖO2V��]��lQ��ru�?����֛Wy����ޓwL����K��R��79���<u�s��I��^dh|�l0d+.�m�<N�ѓna8�.X[즉x������
͗n�(�� ����7���]ӻ�M�M�[���z���K��A��f	��"�"��7=�xj9�(j�HK��ͭ�~U@Jux	æ��ҵ��'괋�D��=�"�Tٸ���j�j�x:�A$�n�d?.	��),��ZH<��.�KNQ����oN-�nq h��7���uH�� _��5����E�5�6��S�*t0�@]�I�
�Gm��(+��]�Ewώq`��}l��y�z$u�����n�
��X��ϥ=���LѰ�-���N�n3���Y���J%��n�f(��'*�~H �?BюT����@�#xg�n�sŠ��PM�����(��� ��?3�F���>��]1�d��u���y�ܭ6�����pw����/2��-�A�PJc�Xj\�k�ak�v�`U��
N�Z��_��̳9�7ݺ@&�Ʊ����c�<����a������&�j�b�d*쁺�3�-h������d�.�Ph@ps����n~B��\����@��?N��Y��[��ty������T�V14����'�c�2DĆah+��KN�-W�뭈{RBru����ײ�|�Ü�0�ͼ�P��Q��[�&�^���9<{6���M�x���E��4���\58�'��GJ�ޠ{rE��eh����`�ހ�����"	���0v�ڳ���	��%\� �A��w:��(Y��acc��n�l�	qt��4/���G��=MNPSV͋��lkn�|�s������R~w���/��6�<�<��P��*q��e:�l+�B|g�HK ������-(�I�y3%_?�bMLO��dC��cf�-�y|ڄV[�\��1�:z��>�»���S���ji���q,s�t��N0��#0��(�S� $ �DG��M�/�(�9�0Tl0tw t���[Z~�o��0v�س�E�E�;�OL��cb����^�z�6���:��U �*\�5�}7���UP��E�K�����q�Ăeh��Ԋ ݓ!٤8��A�E���B��������z7�{��I�Z���[j�V�y?ֱv�ґ3ݢ`C�^cfm�P��A�J���u�b&��h4�5ո�~5��?ո���82MtD�ܷ4��\_��_ y� #�w%[t:�$S��aٞ\?�-_b�d��y�c�
�Ku�����o��3�����=�Ժ�R�SR�����eW �Ѥ��[�M瑎��,�#�vZ�7:ǆ2NеV�Kjkkn��o�4��I����?I�� 3�63��3�P��A�b'�Ȟ���r�	H�K��V~�[�#���+�v� �?@C��PbTm��bt�Y��by��p�9���#�t&#}�#��F��h)��\���eJ��y6��x� n�e"�6Hx+=�x2���CUG�:Pi{�^p�Y�7�v�z�m���ޑ�ސ"�� �ğ�g��R�UR��R�N�u:��2X���J���y��e�B./2h��R̉?I�T�&�]oJ��jm��bb�@��ч��������鲵��H������{�����@��D��V�>I/!ZP[/A�w9R��GY�s�VhŤ�df���t�a!���O����X����4���Ȯcee����^#�g(�n0�$�
�M��R�Z=�?N"4�w%�|F�͊@J�U�k�hKYKkn����G��xe*��"f��(.-ػ�2�N
����V���� &��,/`���t�7IP$6��SZ�m_nBTJ}؜w��`eXV�������Ͱ��ټǟ���X��F�����VB��b���'z>$������Z=8�岬O.�36��@��EL_�qT[nɹcj}ؒry�瞁���+���-�����"�(�,����=�-0/�:��C�w�>g�1��w�i��3�R;truI[M���[m�2QH�qt�.l�
�=��I%䊤��޲ğS���������Y4��p'&���*,;!�?MP$6)�_b6H�jqEW�y�Tf���cug�Zp��~��q���^[�)�%�����D�B@��?!$+A�ń���w,BG��
���2�%{��1069�?�JH#��@�b�@�k}��vy|灄�������򤶨"��� ��#"M�҆�:���\�٭V���O*��l�&!�_Z.@���X�R-a�MP���i�.Q��qtc}�A'����V!���
E𬾙򃹼K�͏�b���M��B{�G�JU���Tk��F #�o0��I �gADҐUۡfA��be�~����`�lm�/�Fi������P�4������3�� @���Z	�$cgk4nw);��my�^ǽژu����cjc��x�~����yu噜%c��%ƴ/禓��R�Gݠ!������8$�n�y�;��f��.�}/:��;B�_A��d�a�'K0kn��tUi~�������.�ewt	B�@��G�����e�1L�����EM VY�R5��mf�(+.�= ���DGJLOޛa�#n�M�1�5ơ���Q���������|A�?��F�?���*04H&����!I��	#: �8	!�'�.0i�j>P+�KN�d�"adg�����y�g-���/�Ę�(��1�8���F����	���d�h.	v6�w��L'&�L|%q�bEH��036Ƹcj���OaG�Yr��gy�e�;��8����	䔦雴����9���Ad���4o���hb����FC� ��59�`$���,/2��G��hJMP�Y���Ehkn�;z}������!'¥���80g���HF����]c������?BEH�q��.�i4�u);~0I�>P���MORT/���&�`svy|��f���#�T�,��.pC�V�����U�TS}o��v"yy�n��"
KY<?�/��N.0391u�fi�R���/H����rux�}��׋�����+)�s���B@����RP����ig���yw�����#�`Y�gV]W�5y\_ǅh_�	t�VY\_}�l~�����и���ћc)�2�؀�
����7�V?!�H�V�r@
(�4Z%|?�H`�=��#�I�yp٨FԽ�}%[1�7�q���v筷U����h��)���ߥ|���Q�� =D/�����Dy��P��m_D�E+��&)��?�!j�AD��=�C�^`c���J�� ���R�{~g����������T�����k.�r��,I��7��?�]�'��}-?�4M�BT�
�q��]���Mk�mp�;��C�
������%����;�y��R��ޟ��j%�6v1�B�=�N�I�Z�U�f�!$���u9<�.h�NQ� CX�cf��H[0�{~�Xs@擖'ꀋP���?��`��2����fa����;�DG��H�Y�T�e��p"4�w� 8;���IMP��-�K��kn�9�Fi����#戇%���;�����S��*��k.��(B��>�O�R��2��("�-+�&6J=@�V�O�U�PGV�gj�a�;��s��كz�횝.񓒪����-(�����.��<�n
��|�Wv'�O�`�c�d
&(+.t9<?s.:�NQ��$�ch�p��uo�g����q|F��!L���������&�(&��=v�t�;}
P�bhlK�� H/2�]ߏ�FX3i�SV�$��}��4�v��Յ�UxH嘛(睓�7.���U���RI��c����w� ~C�3�o,��U�y�=���6H�ޕEW�8ȥX[�USn��d�e5$���V�	���	p���;{�������\!�*Ŏ���Vڃ�����B�f�7� "%�x*2��%��EH�O����bt�5U��uxg��E�~�|����륭#�8��N��j#���Q�m2��B����B�K�G�E+-�`&),�W[�>A���g���as�	�p� @c:σ�e{��tÊ�H���{.�+N��:�0��l�ς;����/�R����A��(+�"p/��dǔFO��WY\�IP��psz���.ݍ�c��젣���pA��x������K�j-���>��E�Q�	�`p�d�uۆ03�Ǌ�+�3KN��HC�Ycf��x��}�����Y|�.~6�k;��}��ݸ�"��l/��~@��0w�t�V���}e/2�tȿ1W��RTW�L����:��|~��o����!��R���9��ż���R��Y���q,�=A[�K�SV��v�l*h�%(�t��	&a]FI��>A�^a�?V��vy��+ڊ�`}����/����+���:��S��[����=@T�F�����	��^rr�`-0o���yE�@7FWZ�!�ۓl�g^Y�~��{�
����õ��5y���5˯��	��W<?�c�D��Z\yfo #&����L|>Aҕ�A<ƫ\_�Eݒ�i�̉�V��ٚ���(#�(��8������[���[&n�j�t��2�mmɃ"%�	�47ȋ5,f�LO�=Dv�dg��ms�ff���t���(녌�����¡�������3<>>��Az�v��Z`d�~"��,03�9R��GY*���V����i���s����.����������=2�F���T��@�5��p�x/�}<��ǎ�?�	���(��3v�Tt7������F�L�hil�Z
�z}D�)�������50f���
����Z1)��I�;��}x����RޘS��Z�k�|���6:=�C��Tf��`dg�mG�:�6����i윮񣼦���9}Ȫ�/,��%��je����?�
PL����
f�"�'@N�5G���AEH�7FWZ�!��2�96u��Ň�ᕧ] Ǫ� ��)ܿ��<�ݓ)aT0��?vj _ZX]�҉=��|%7�,���U��I[�Pi3�^p�&�u�q����o�+������a���6�4�ð�����"(,M�	5��p��?� �QqG�b(���|k1�H�͆@Ҟ]�V&�Sc�d��t�Ǹʛ�ܒԵ#�&�������m�ŵ����_c:�<'li��j.����࿚ّ]z4��`·M�{M����QI~�~����Ð���ʧ�� ����m���I��F�R(f�������ߎ{���QF� ����$f���\�JN�T��]�b{i�p���;�l����ۑc����9������W��]�V�!����e�c�O���a~��J9�047�FA��6�<�L^��cui�������·����㜮�'����{E�P�q)��h-��@�H��� �bX#ىm�f�^14:���GYZW�^a�-�p	�mrQ ����!䆅he��9��E �.�4�:Տ1'��͸��D�?�P��7��$��	ܭ),��>�$l�DG؛5<Ƨ\_�ETֿtw�ml�׌���D
U���>��&���j$��A�K/�(�KA���+�xm��p�(`��9K&~FI�ݘ2��N���R��w��?�א�}�ĝ��4� ��绾E��V���]��k��
r��EN隅	�`��k!$�x�9<͐:1�QT�2I$�il��ba4ˁ�Ж���c`�.�,�Ǩ����!B�V�-'���k><���e�=Ԟ]�f �zx1C���@R�3�SV���dv�,��;�:����T3�ᚬ`j�f�-��ڀ'$\��R�4V�F�9����v�zj]���un"��~0B3&~FIڕK��O��h�r�v0�ȁ�nδ���%����׬�6z�G���M��!_�]��v9���C���Q���[�i
�s*-҄�;M����U���bt(2u�9���y~�����򡳑�/��3�#��׵�8�+��l/�К���?�P���J��h	�r),������4�:UUWZ��[f��gr��ҍ��I҈ 3����L���A<��������1h#�4����OI��f
^��g�b싶}-?�x�=@�V�;��[^�4S��sv�<k�ԋ�ڐ^�m�kC㶹��M���֐�V���g����uq G��K��"�^��v�o4��� ���R�(�0β-�.9{�H=G��^�U��(z� {���J!����������qH�|Q�c�mQ�J�r��)'�M��ę/� ���VY]`�.���ZxB�F҇eXQ\���ni꠬������V�:�-��1�Y0���ob�lP�I�i��(F��7U��̙7����_5�X,8y�N�h�y�a��^ܡb�}3�LoYB�¼�V�ךe��(�����G����I���6�at�$�v ����DV�4I�TW�Q�+~���Ra&:��~І����3�x�X������>�] ��t(��hh��gO�x��d%h�k���,/��8<���I[�VӰ^p��(W�3wz�\��PΓq!\]g��o�
M��%p��Y�^5�i��B�������څ	�^��d�"v���147�ˆ(�ג��Y�c�g��^Y��y|��-�w志�!e�2r��5��G���J��^!s��(��v9���@���Q���X�i
�p*-0��>PГ�42TWf�ew���G^N9~��|Ꮱ!�F�h`�����H������;�/��o2�Ӝ����B�S�N�_�Z�k�f�w�r܃�~ȏ�ʜJMP����]������~��݃~.����5�b�S㼿F��\WQ���1q,�=}xb���R�U��z�����+.�� ��@C�5��UX�'J��jm�<_���Qt���(�e���@E��	��Xe��!��p3m��9����}	��Z���$'*{69ʍ�.�NQ�?F"�fi��g^2�~��7vBۖ�*�w�RU������)���] ������u0�A�<�M�H�Y�T�}�s1tȉ/2��H�
-��MP�EЪeh��F]��}��r�%���!_�5�R?�����T�����S�o��b�����z̖���ow�s�v�47��EWך�;�[^�	�l~��cb�<����擥%蒉�c�����L��ފ��?4��s6������f[�]���!�n3�~ȈǊ̔���KPTWC��cf���'��������'�|�3.(���H�TO���)idF���>~y����S�N _��d t�o����M;>A�Ր2���~\_b���+���}����<�#؞���83%���MH����"b�.ni���C�~X�X���0z'9|x�7:�P�5��UX�'J��jm�<_���Qt���&f��&��;{��;��P���P��e��
e��z��z� ���&���4�'*��B�<?�1P�QT�I(�il� �x{~j>͊�!����T?B캽��j��`c����̀0����F���Q��/ #�r/2��`>AD0PS��_beQشqt����r�Ւ�&)ˡ������GJ���ȴ��hk�����08�����
�FY�m�Vq.1�&f�FIڝ7>v�^a�_V��vy
�on�ю�"���馩:�G�� ��/سmc��3b�W�v9{C������I�*��*�5�<?+ǋKNߢ�C$�cf��4[4�{~�,sDՓ�'�<�T�?B����j��`#��z&��x;�܊>���S���V���#&)�w58�̞DGJ6ƘVY���ehkWܹwz	H���VS�!��������!���+��Z�b�.IbM�mC�;��� rc'�RTu'9�3�z4��CTGJORVY��)�dkn�tvP�˅���������}	;v�M�N3��*04k���{:�~a	Ɲ=��"�m'�� ~C
�����a(�/�-��<�=I��^LW��i�ࠣ�w�v~پ��MƎ����ߡ�m�w<�k�gT|E��'�-w�;/2��T����ܚ_��y�j�n�y������x8c��"f�+��zH�F��%]J��8q4�ve�� u��m Eܦe/	.1����wD�bM�Z���`�}hSr�sv�=?���M�����N�h�r<��ſ�8�-f%�q.����{�~#��f�g!��A����I(Zx6��Q�B׻6�yXBU�K��Z؝d+ki�x�y��䚈���刦�p�������j	�b����a�)����E$�\z �z��`e��]�=��l�k�� ہ�,�"��D������M�F�6��z=��R���Mxm��p(`ĺ�9K&��FI�O�^�G��c���gb����Tw���+�ﯲC�����[�����s6���6���Ffhh��k���(+.���"cWBEL�[ߢd�F�fi+�w�	�z*�02�o!]�0��>7�C~W+�%��S��c ��m�h�{��*�AI�)��[�fܑ*}�G9<�Q�[�Y�fE�eh�_�>�q��̖�P �_ݤ5ը�7��x����E��9n7��f�q~h����S�}��D�&��gd�����Cˆ��2�RU�g���41��~r�����U��Ȝ���g��+{̿P�N��'-1j%�N%���E� � �
fiF�l�Q9&8{-Fh�;M͐:ґK:�Z]왟�n� �Q�~�����X�o����m���D;�M$�V-�_6�h?���X��3���>�b�&e}#|1��.�25$D��D]�Rd�w��dv�\��M�z�}J������`�w����7.�@�I �R)�[2�d;��=��(���T���Zmsw�(\��4Mw�BT�֕C�`����41��k��w���ߓ�蚳m���8����KB�I�\؎d����t�45��AՂYQ���,,.1���:?B��Kd¥Yk���k}�r���s ��?뒤$U������=����yQL����&زG�B��{v����P�PG����~%7���058�>�GQTW\arfh�k��`c`Ń���s���������B�@���D����.��t7�{��6;��U��FSX�p�q'758;ˆ��Lek�Zl�"ى��9x�
�G�񁏒����������������L�4���9��I�NO	��U"4��-03�9CFIK�N�C�IFcil�s���ρ�x���䘪*�1��Z���5������i$�5?�	D�
��w'����(�c�t�-03�8QS�FX�6TTWYr��gyk�j�C�}��׋�璫�젲��/.���?GV�:���1�H���~�RUUR}�&0g-�p�$\s7:y<���USV��_dg���v����ٍ�ڐ(�e����������T+�>;��4��y4�EO�T�Ї%���&�1*s-��6����Kd��Yk��\v��psv�{��Չ�吩�Ʞ����;���ĆPŸ����H�R6�/��'����.��1�z �r�r:<?�Є��UgB�[be���r�~�B����������)��� ��Y�`��#��%�e�n��X�� -"}(A7�6H�?,)Ҏq\��g���sp�8�Cʭ�R	�!ȯ��Dt>�M�K��\)�e�k5�?Czj��x�<����"�\'U�p*347:ƽ/ώ<R�aW�Z�&(Jqs�nv@q����[$ֳ�j�q7ps����O�����S��o!����zw� zȔQq� �n%��킻�%PʏM�\ٚX���l���x��i�
��`ᛤ�����=4�F���Z�����&�r����v�2ɒD!A�?ߥ��*,q�.�*CD�3}ݏd��k�,�;��pw�?Ȏ��ݜ�gd�2�0���/̳z��e�c��^�"�TV���I�Zd�X�5"<<-0���H�B[��Pb�F:�W��x��kҔ�B�$߁���~���:x/�B�����O�ħ`�����DIMQ0���- CڤbE8��QD�78Q��FX�MfX�[m�_mil������Gȫ����%�ɐ����Bn�����O��>�H,�%�}���և���0����|"g�6D��x�hYґtfe�_beg���tyz}��ڍ����%MP�������5����"��1��G7��"�.tu p�z^�W�����3S0�7:�rܟ@E�$�j袅|�i�X.tx{��̯�����&"���0�/z�.�4����*���[�v�F��N��0"j�#6�w+=95Nx�CU�Jc��Xj��ߊ}�1�����ˮ����ꝯդ����������"+-/�6_�������N���LaxGp�ev�y7vo:=Ή7�ڝK>H�^ad���y\��|�yt�̔�(뙌�䬯z�y�#�Տ��8��%��M���:�b�O�0w)�d�I�,>�yb�AS�({�Vh"�A��k}7�Z����L�s����a��
���&jx�3���B��[�P�(h��jځD�<?�Rs�ޫn,�f/2�=*2��7�=`��^ʉ�tW��wzA��Ҙ�!h��M���h���=�����DQ?���g��o�Ig���
���M�׌*<��9K�N<�K]8��X[�o]�l~�x�{��C슜w''��)��﫽n{��*�.�޹Si��k��1��H]�a��u��#d 2���/A��>P+��KN�T�\���hz�T�w��郄��֒�$ߕ�0󱔿"��F��n��] ��{��u8�ً/����d��d��>tWb�8���I��xL^jc�0]`cЍT��tw�A�BL܎�������9y�g�N����(��)��u�X�]�琔
a�Y�j��4g+.m0�I�,� LO�>Ny^a����U��
�o��to���)i�����@������X�<-,(3����NQ�C�T��U#�"�!vy�s%��%��ILOQTW�JI<zil�7��57ʆ���Ę���ߥ�9���g��Q��w
��i,�͇"��SUU��X����
fiq��,~�-/�:��CU�6c�VY� r�)lork}�ɂ�����䝯�����W�������X�k%�_�i�r{
Cy_*�!��-?��n=@�f8iR�][�ʰi{�q�{�~��nп��\��Z\﫽�o��L�г����S�p2�������E(Z������qL3j69�JВmX7�*WZ륈o��?[��{~Ѭ�vMʖ���ɧ��F��U�S��,26mb��t1G*��N��"};!Z�,/�ىl@RнW��H�!a�h��r��\~�:GKm��Lb�`c��8��m����|؍���f�1��X���$D���3X}+�~>��:;>�r֥K��V]!eh��Y��f�����������5�=���J�?\�'
������'�����&Kp(�)$%(��\�Ċ<�=DLOۚP�Ms�[nps�y����Ӑ�ڝ�%����=����I����]�"��m����3(}�zq���s�,2�.��6Q�K�zT?��N)li%nrux��B�r�������w��9��$�����U����bQ�����En�G�`�]�b�&�2u1z,��3��.�W���_n�?hkn�{�����W������䩶/o���C����S����g�*,��w�����NBP"��"��49�:tD�J����B�K�=��["m�sv��w����ك#��)��2��Cܪ����S������
0�|9��'��#� +�3:�6�9<?�0QW^�Z��X_cfi�2�G1z~�����������7������I���G�Y������:�h��N��3P��% #�E�|3 �D��/W]<a�k�,Wt��e�9�Ɖ������/��6���٥5�����_$Ҟ��f����u���L��Y���0k�4�:}ú4.K҅��5�N�$Z�e��v{~���ӡ�%���~{F��R��^&2jS#�jiQ�x?A�Hn�2S�5�/�}ln�u�I}�ViK/� �#��/�:t�>�p���Y�q��+�<���A"T�]�c�a�\�.s��4�{�e�T�3�^�.���� �>ADV��ܛU�^Y�s�v�Ȃ����ͭX����&ߵ B��.NK��L�hh�^�MM��Q�u(	�h�=,�I8*����F�?X��M_���T�Z��}�w�og��ό���n�����&�;��6L�A�� �g'�j�_�|D�N��^�]X�*��w6��7��HʂM�L��_�&�k�p��yc�	Ɉԩۚ$���(j� �hҹ�!�#Z�`.+�+l�a��qn��D`'/w|x����{�-M���R�\[�j���|��}��Jn�ѯ&�-%�8(�A��J�Q�Y'b�k�vr4��{!��L#�[�^5�P��D8��_�%�EH����溅l�����w���%�������}.l8��-�A�ò7�&�O�޹j�t4�h�d�S|�աa*��*�/�J8�Ύ_��W�\�se@�/����=ȫ���V��b��۪�-��E�4�Qк�`&�i��`�}4�2s"L��L��&^��Q2� �=@C�
��\�![J��(V���}�אz� �)�-+�;�C	�H�$&��+��T�q)����8�	?�`d�7�� �``�O:�>y�D~�<:a��%�i�o���w����H�Q����.�2�:�v��A��M��*_.�h'�q8�|q�r��S��qs����uJ-@��9<?B�ӏra��~m�ϊy�O����y�r�ؒ`ᛡ���7��D��$f���ϕ`%�Bj�����LUWW�S�YH!�iD+�=�2E8;kATGJ�Q�Vi\_�Q�,�Q�xI�ɐ�U�� t�jp>2��J��V� `V�֐J�z6 �J%˘\7"�%�fI,"�D7�4!�	ԐsZL�rb'�xjWzV�D���ո��]�1�п=����U����e���>w�S�W*�S6�����9��-32�?�re�N��pd0�z�ƙ����α�	���ò�������������ƪV�����B���FM*��F)Ύ*^�qD/#	O58;>ʈkZ֤wb䠃zn(��ț�tXz`�����!�¹-����s+�G��S�����k'
���{�)�MzR�`�Ӟb=0�vI8�rU@%0$X-�LRO�%^Α�mݠ��O���帧����л(������������3�7d�����~�	nm�(uwwX)�tWJB��X�ӟraK/Q7}cfil����ҥ�α��V��-��å���׽���R��^,���\x<�@#6���ע^A0�s��Ɗe\Ҟqdޚ}l0M6A<XBL�U�tzwR����$_,��¤���+����B�C��Y�7�{�Gp�����z���;.���^Ei�*[ORUY#w*m/�V�pux%K�����ػ��`�4���@�������X�^����p��/|��V!�Z-�V9$�����>��065�8B�ul�"複z`RrC熶ҥ������ڽ����}9w|��|��ߺ�;��I�������Xžh;!�|�NU-?$:=� �}Qc>@�^a͆�o�\PE|�IB�����l ���ٱÞ|�����F��B��Q(��� `�ƐC)Ą$'�t]5G"�BE�څYkF��fi���w�d M���Q��Û��q��uo����|{����a$�j-�s�z<�}�M��Ȳ]+p�&)��_7I$�DG�
��[mH��hk��y�f�O���SLFᝯ��
��,�ͨؑ��(���#����L��[x%���
j�ЊM!3VX.1�k?Q-jvLO��]oK~�jm*̧{�i����H
ř���Ц�f0�ɥ���ǄV������|�� ��U#��G!��s/A
e<?���M_;�Z]�k}Y2�x{(����v��X��N���'��V2��P>��FJ��BV��a���m�y�*�%'D�13p�=?��IK$�U Za`cX�mox�y{�������������4*��R6��rB�ېN��Z���f���r	�~�!#*�-/@�9;Z�EGr�QS��]_��ik��uw�끃�����4��L��h'���1�˦?���K���X��d��.pJ|d���)+��57��ACڸMO �Y[�eg>�qsZ�}x􉋔���������%��
1��$=��DI��\U��a���i�u����%'��13��=?��IK��UW��ac��mo��y{�텇����������~��|(��t4��r@��nL��[��zd��	���!#�-/"�9;>�EGT�QSh�]_~�ik��uw�������������� ��&,��<8��TD�מO�����g����|�h�)+~�57��AC��MO��Y[��eg��qv}|2��4�����������)���4�Ǯ@�ӦL�ߞX��d���pV}�%!$�?-0�B9<�vEH�YQT�c]`�iil�ux�������������+���7Ľ�C���OE��[u��g��s���� ��),�C58�TAD�^MPӏY\�behk��uw��,���������Ϥ����++(��*@0����;MPOOLMc[df*xjt�v�w����T�X���7���C��LO����������ޢ���􅈋���/'02�B�CGK?BHV���aVU�jp gy|{{xy����V��]����������QTW���c����פ���������		 "�*!&�6-2�?E?�TJHLY]c[`��oumr���#�����d����DG����VY\_�����������������ת���*4�#587745KCLN^ScSg��euey
�}��T���147���C���O�¹�Ðܔ������|����� �!, 2�7;<21@����DNV�dZX\i,x0s|�xvz���'�����������z����������lo��x{����  �� ���$$�-%402���67?CCMTNY\�Im]bm\iwy}���&),/����xpsG����¾�_������tw����������
����+�):4D6FJ6���\eb����Qzw{ozlV������k�������������Ⱦ��ѽ��jmps�y|��������Ѧ���!'�,&8�-<=����
F$+R"07^	�<,@NV�LZb�Xfn��BIHK��������̕����������� �	ȿ	�'$��/6-67HENFK
N`cbb_`vnwy=�A���������_�����pg����������֚������ﲩ�������%�,/..+,B:CE	UMOJ\_^^[\rjsu9�x���G���T����f�������������ؖ��������������������)�����<J<BE=Tcdj^tlhuqJ2bkdcAZUZhP�������h��q���������o������嶿�������	��)1*8CB�#,�"
R^ KL7t{B<<IBHHNSL&),/<x������w����������٨���������ʲ��Ƨ���%!-#2-�������&UW`T`i%OwqiA*##))"%(+~���Z=@Cf��������nn���䭖y|��������ɬ����!&4;�����BEJX_=UearajkC,t�Bmn++e�����c~��������t���Џ������݈��������
���##3%��157G=M����3bdmamv2\�~vN7���������d����q�����v��������tw���������� �Ͱ�'".��������@FRVZ���gh]mbbxh
����TZ(+��������������X[���לmps����������  �# % ����?=CC;>@�ET]YbcmZiaerjzv�v�!$'���������EHK�QTW�������o���{�����������
$#,(����GELDKF��]b`XhgkcgwuH���&),/_b8;KKDGwz]]VY\_����nqtw%b��䭺꺾��� P�������#'+/37;?CGKOSW[eimquy}������������������ɂ�����������vy|����摔�����㩬�!1#/8@����+5VD0 %,Kvy;`SuY�7<�z�UbJ�|T�}dj�l����ʆ��`c����rux{�������ϙ���#-'."$�	�3����MNR\d^p-fqtTU]Z�����),/xy�������PS�������k������������������"#).$58-/!:N<D�����?H;A�
9�"#&(,�1:7:{�C\IL�RUX��ձ�����vy|����4������������������������������#'+/37;?CGKOSW[_cgkosw{������������������������#'+/37;?CGKOSW[_cgkosw{��������������������������������
#'+/37;>���KOSWZ_cgkosw{��������������������������������#'+/37;?CGKOSW[_cgkosw{���������+��������6EKAFQT����Z(alo	ru����U���369<������ǂ���`�ϗ���ux��������������$�)+$����&)(
����8b^_sttvtq1U���@o��������>AD���������Ņ����������������
����(0-=D:7<���&XNMc[k]Jbfz*Yyv{�����(m�Q�����c����RUX���ɺ���������� �������4&2;+6<�,)*�%QQP\e�8nf Ku}Wt�\�����M�����_�����q�������il����������
��#* "�)=5E7(%05:O_f\Y^�Bqrxl1Xdc=w��Im����;>AD����������eh���������������������"!+&��78=NOL����3WadNsmu~r�3i�}���H�������@���������~������������������	����䯲��'3)3/@C�==OVJZ1`b]cduug}{�gvdgj��������������T����ǽ��������������������&/8?����������`Uelb_d:�v�����#&),������ADHJMP����׺��ϓqtڽ�����緕�� %)$9:4<8�/$:';1K6:K>PJT[S\^oi������n��������������ʷ�ad��pxvy~��������")!*,��-9?= ::P@VL[V1��">!O'*-U`hgn�BEmKNQ�����cfi������~������� ����+54$8.-���
RF\[K_UT��8rgqmn�PF������,/25t������M��������hknq�������ì���

�����ⶹ�����	������<V��G��X�)k
0##"%��.1�Y:=`�����RUx��a���m���y��ą��������������������5<��=���J���J���j���c	��!�'*-�369�?BE�KNQ�WZ]�cfi�oru�{~���������� ��)���9���5���=���S���Q���qkgs|���� #&)����8;>A���Mļ��\_be����twz}�����������),����50<E����L\��XXei���pl}����%���1���=���I�ºU���a����psvy���鈋������.����)5-2����AM��LZ[�Uk_�aqiny�!����0369����ǜ��ű}���؍�������������������,1-� )@&8�@ORQW!����LNUYW������V����r[��������ʈ���ҕ���ղ�������Ҙ����!!*�82*�/ADCC@AWOXZj"oru.jv|z=����������>>7:=`�f�l������Ԅ����آ�����������ʽ����������������8@)L%njp	1�7�=KVyR���0369v�BEm�NQҁZ]����loru��������������029��=F(JQ��;LL@bi��Oqx-o<6xE?�@H�)t������������ſ�����ľ��������������

㶹:
?����;?KTLLRQa��_y$,}0;;}<lj�Q+.1TW:=�����������ڷ������|���� ������������(��1��:�ODT[QNSdX]h 5	44j}A!����0369������NQ���������������������������� �i��%G�;��,���8�K=5��IA⼰�$r�8,/25jmnAnu�ŵSVY�_be�˗��ث��鮯�����������*���%�--�J1X\A'C;B76ems
a5RHa\Nv��Y1dejkpqvILYR_h}'-���Ȝ������ ���������������) +11@@A19%vDe\gmDm||}mVua��j��[[TWZ]������������������������$��-�����&����SJ��Wee�ine|p|:�|��^&)5/25E;>AN����SVY����hknq��̻������ЕԼ�Τ���н��������������JDT�RTT�e\pew|}t����%���1���=���I���U���a���m�������� ����
"17)99=11LRNHFFagARhllaa|�\�}vv��k���~����������ǔýӭ��߹�ژru�������������'��0��9��B�KT]f"o(,x16�:@�CJ�LT�U^�^h�hh�qr�x�̆ҍؔޛ�����������	��ध�������;��D� MSY_e!k(q/w6}=0
8]w������q�������������љ�����������������"�&%#3@-A?5;KX-Q[MXPVfs>bchskq��_y��g���z���z������ʛ��֧���������������	�˥�����������0>��gZFU�7r^��O�vX�25�g��p�JM���Y���e�Ϛ�twz}�������������	���)�&�A���0J�HWZY&!lor,oi~};s��H"%����nfi���t������ȍa���ݪ�����������
� թ#&%���8;>�02FD>SRHWX�\knm:25���@�y�����X���e9�����z}��Έ���������譁�������� �"%� /0������GR����Zj4��/::MV[#&)RRbhqv>Aj���ĎVY���գknqМ�}���댏�����
!*,��������76!OF[VQ]fh\le$Zo��|���"%M�h�47:=h������������ڊ��ז������������% '&1/ j����3O7LI[EUXgW_Wshcoowr~�}����������������ĳ������������������ ���
�$���0*0<39E;CFQJOD]WKai`[fu`ne�xot�|�������������������PSVY�������q�����������������&���#��,��D���� L������k�LW�}�'"%�/10�;=�G�LWRUn�_ad�km�w"|�������`蛝L�R����d-������>ׂ����]��$I��Xm�n�!�x+-�7�<GBE��OQX�[]��glwru��$ً6�������f��\(���5��d@��^L��TX��Pd���o�{���')8�35R�?A~�KM��WY2�chonqf�{}�������������� ��$,��B8��`D�݀P��\���h��t��#%"�/18�;=N�GIh�SU��_a��km��wy�탅������*��B��Z)��v5�ͮ?�ٴM���Y���f��r	<~X�!r�+-��79��CEƺOQ��[]�gi*�suL��h�������������'���3��?��2K��RW��jc���o�wЃ��')��35��?A��KM��WY��ce��oq��{}���������������*�Ŋ6�тB�݀N��|Z���i��r���#% �/1�;=0�GIL�SUb�_av�km��wy�򃅸����
������"��.��4:��JF��bR��]�����$u���!��+-v�79��CE��OQ��[]��gi��su�*����@�B��������+���7���B�ռN��Z��f���r�~d�� '&)3/2�M;>�PGJ̈́SV�g_b�qkn�wwz����	������!���-���9���E���Q���]S��i���u+���
��$"�,+.��7:�QCF�bOR�l[^�gj�psvy ����:����`� !"(�����2D'?<G"QZV_��z�ImeqV{{rw��|$x���������������TW�]����ѷ�����V��������w�,6:;/0F��a�(LVRdX<bhdC�Tz�{h���l���s5;�������ƻY1`��ܿ�������Ć������!�(317A��:�OEDZN<aaX]nqB�gt�b��x�����������IQ�����Ƹ�����vy�����������! .�~�E9G*ANDCI��8�G\nRnkgwp{wy]��������y�����E�M�����������ru|��������������. 558.:C&=J@?E��,�7Xj<qqtjv^��z��#�,��������DGN��ʬ����կ��������ǉ����! �(317A�ѿ�!BT9UUa\W>famsqh~v�W1"u��p��������FI\P��̞�����Ѽ��޽�������	��7�&891E?;!=MFQM,���AbtFuvyp�yd���{'�.w���������������Ťfidp����������󓕚�	�#��?�91=>D@���IYge_ma��gwq}���&������8;6A�������˽��e+n��������ǉ���
���?�.:?C2@LBE�A�3Tf:pdrDskoax�{z��(|��������������U�[�����������������������*.:
062Ӣ�HRVWTP\2����Ghz\�sZv���$'�-u����������Q�Z����������������������f��
�'$(')0+
?;A=/GNI�B�ChiiamfYp}srx�c�������������}��������hks�������������<��,/��-CB�7�!BT)OUQB[o]�^Gyon�xc����f(+2{����������͙[#b�����������������	��$./59:��F�>P+QLQNO]8icseVz{u}y�Yq"k��q���������K�R��Ρ��ѯ����������ˍ����� ##)����8><3I%@QTENO.��W�PgtjioACZ����#�,������qs����PS�\��ֹ�������������Ø� �'/�( 58��X�#G?K4KXNMS��K�Asih~rV|�~]�&o��}���������ŷ�X[c���Ѷ���|���		�)'-7����?E;=K4J)WZ`W�EBRQKU?A@y��!�)���������E����������fi@p��߿�������י���
�"6ý�49&M@PZ:HVbU8n:��Zpudy�p~���n�p25<������ø���_og����������������
�%�1���0B$9IPFCH9]Mcgh���Swo{cVcz�����l.1�8�������Ż���^a'h������������������ )***)9@638�ً�&JTPbVG\lsifk	JU����t������~�����HK�Q�����ȹ�����ݾ�����ΐ����&-# %���%I9MR4IY`VSX9mnkFn{{o�w�a#*~����������őS������������z}���������	��",��>IL���?cdHlm?�]��V��j`"%+���z���CI��Ę��̢dgwn������Å�����䦩ð)*-
2;���)MN15YZ4/���MqrUIq~Pkcjxews[���9��t�{}|���Z]*c��������������Ɩ��������� ��*�8G=@����),"3O:L@ZNHe��~����,/�7�����G�O�������e)m��������F����� "0�h�:,<5��K�IVGU\WS�h�gtesx�}clrbtyV���47�=�����������a�h���������������C�-.2 *+3C��?�%MVJZYSe7cipeKgwp{w�g������������E�K��ȼ���׵������~������
	� ��/�7@4DC=O!PRUOPd4��Q�Jy|{]�y�l������p25�;�������������ٰ�������߉�� �"&*���F�9B6FE?Q'HZ,[^]^]<��S{�x����u��n�����~@C�����������g�m�����������	�ϣ� �"�0%)62��?IDKRFXTU`c���snyr���u"$T.@Aa:LcmFX�yRd��^pɑj|�v����%���O���qͦ��ٲĵ��l���������������������b	�n'rz!3V�-?F�9KF�EWF�Qc>�]o>�i{2�u�*ف�卟
�
���	������!���-���9���E���P��\�R�y);��5G��AS��M_��Yk��ew��q���}��ى��啧�񡳪����	�ˮ�׶ ��-���8���D��P�\�h+�t%71C=OʘI[ڤUgڰasڼm��y��ԅ������읯�������������(��5��@�L�
X	d'p!3{-?�9KB�EW2�Qc2�]o:�i{6�u�؁�䍟����B��F��: ���&��N8���>��nU�vazm#�y/��);��5G��AS��M_��Yk��ew��q���}��剛�������	������!���-���9���E���Q�]it+�%7�1C�=O"�I[*�Ug.�as2�m6�y�>���F쑣N���V��^��f��n(��v4������L��X��d	�l'�|!3��-?��9KƠEWάQcָ]o��i{��u��܁��荟���� ������$�����������C��sf�F
�"Q*�.647b�A�FQLO�X[�dg�ps�(|�4���@���Ҡ�{񬯳⸻��ǵ���Y��7?��_��9� Arw3�#!$�:-05R9<|EHCDQT�]`�3il�ux���{���E��j]���@��20���M�̛���\���c�����"�a�w �Y),�e58�qAD�}MP͉Y\�eh�;qt�/}�%X����>����@4��8��������,��3!�顦��AA���
w���"%��.1��:=�FI�RU�E^a/�jmP�vy!k�����ʖ��æ��[����?���_��֤m��c�����2��,�u�'*��36��?B�hKN��WZGcf�kor�{~gb��@ٓ�2���m"��܀�����ƒ��Ҟ����>��r4�����i�4@#&�/2�;>�tGJ��SV��_b*�kn)6wz�׃�ߏ��"�������ͳ���¡���V�ڀ��擂��X���>3
J?)�"�q+.eQ7:R�CFV]OR�[^6gjiLsv����勎I������'꯲��7������?��}��x(�����G�*E'*in36
�?B��KN�r Zb`ci:loI�x{0 -�����虜�&���S�������������	������!���-��TL� ��),�58�AD-&MP6Y\[�eh��qt�}�SH��
���Tơ�Ρ��O��j�����E���+����O��.�$�i��%(�?14r=@�yIL�tUX��ad��mp��y|%h���y:��������𲵳n��\��,<��U���b��"	��.	i�a!Ҕ*-��69�BE�NQ<Z]�sfilru��~�w�疙����t�����N��ɂ������?	��	���UG����&)�b25��>A̐JM>�VY��be8�nq�+z}(���*쒕�䞡/MS����)F��S���b��]2��_�������
�D�P"�\+.�h7:N�CFUORmx[^Ogj8msvjy(���������D������C��sv���e��n��r%��g� ����h@$'�?03kJ<?�HK�TWn�`c��lo��x{�����吓s����è��v�����ϳ��������v����c�� #:z,/��8;ϾDG�:PS�w\_�hk�[twnڀ��;���M��>v��j�����˺���?S��>��� ���X������(+�w47��@C�lLO��Y[:�eg��qs��|�R1����t���'ک�]���ԉ�ıQ���D�ܴ����H���C� )�	A�+�!$7�-0>_9<��EH0lQT38]`+Jil|Wuxq���M��]љ�2J���_���J��xk��Z���Me�����%����(`����&)��25�W>A�cJM�oVY��be.�nq�0z}!0��Ò�Ϟ������d��iN�Ż����������f�����
A�H0"%��147:=ZFI��RUH^aI�jm�1vy��������� ���;���^��R;������SG���a��B���}���#	&-?!O�*-��69�"BE��NQT�Z]��fi�Tru��~�1���cD��BZ���Z��i�����������6�����5��Z(����&)�#25K>A�JMv�VY.�emkn�<wz�샆�o���G��n���z���<����Ɗ��`���0�����	
iQ��"�K+.dp7:8>CFԵOR��[^LBgj��sv���!��"x��1�������C���O��i0��I �����!���}"�V���'*��36�e?Br�KN0BWZ�cf9�or`e{~�����\������=���c����������-��j�������+�k7��n#&�/2�e;>ǑGJ�kSV��_b�kn��wz����V���ܛ��᧪
	��^���ϻ��T���Wk��w���c����
Z�8>"+.Od8:�$CFa|PR��\^��hjI�tv鬀�]Ќ��Ę�Ф��ܰ�=輾}D��� �������lK��u0����6z'*�36?B��KN1WZ0�cf�_or��{~�l��K��㿟��t��q�4�����Ҹ)��y��c������A�P0#&b�/2�m;>�GJ>�SV��`bȖ���w�~��������˽���#�j���I�=�,
;���$�+1>7]=�C�I�O�U�[yb�h�nKu�{Ɂ�����M�n�������˾�!�/�;�^�$�y���B�ju
���#-)G/_5n;{A�G�M�SSZr`�f�l0S69�?BEi{��:�p����L�a��*�9�������	�&�Z����B�U�a�lL��w&�,3$94?�E�M@T�Z�`�f�lrxEQ�o�{���������*�x����¨ȴ�\�hڞ��ת�,��������(�	��Xr"�*1�7?aE�K�QX6^ld{j�p�v�|���!�9�W�f�������ع����S�fׄ���������
�H	n��m#�)�/�5�;B#H�N�T[!�'*-fcsi�o�u�{���4���)�7�'�J�k�����:��nջ�������������# B&Q,�2�8�>E$K?Q�W]c�j�p�v|b���ŏ�:�Z��������������� �ٗ�]�q���P���4�H0FRo �&�,�2�8�?�E�KQ&X5^_dj�p�v�}�!���ҖO�l�/�°��R�X�5�h�z�����������
p##A)h/s5;�A�G�M�S�Y�_�e�k�qw}'�N�p���1�S�fil�ru0{~�ڷ��'�9Ͼ������!�-�;�G 
4?Wd%z+�1�7�=�C#JAP\V�\�b�h�n�t�z�r�������۟��C�w��������Ђ֓���0�m����^�#3J!b'�-�3�9	@F�L�R�X�^d�k�r*x�����ݑ���0�O�r�7�y���;�\ϔ��$���������3�K�`p
����"�(�.�4�;�A�GN�T�Z�`�f	lr4xe}�������<�p����_����Ʋ�c�2�>�z��������I
_{�"#�)�/6-<nB~H�N�V �&)�/25@kZqhws}����
�{����� �_�������P�p؁�3�U����9�DWd�f�$�+�1�7�>�DK0Q�W�]�c�i�o}v�|������ʔݚ�d�jm�svy�N�f�����	Ψշ���.�n����p ��Ly��&,I2�8?�E�KQFX�^�d�j�p7xL/���������֤��ѱ2����ĺ���1�h�H������#�9To��{��`���#4)�/�5�;�A/H`NoT�Z�`�f�l#r.x��􋣒Θ��������JÈʴ���;�X�n�����.Yk{�!"'�-�30:!A�I�O�U�[	ag)n7u�{$�t�L�RU�[^a�(�]���"�4�A����m׭�������}������	!'+-�3�9�?�E�K�R^Y�_Xfrlr�x!~-�8�E�V�a�y����������������������,���{���
��U#�)�/�5�;qB HdO�U�[�a�h n258�>A�GJMg�����%�5�ߨ�;�G�����<�^���R�%�e���U�t�
R`l#})�/�5�;�A�G�M�S�Y_"e4l@rmy�х�;�H���������A�p�|ȉζ����1�<�t����*�У��`�����!+'x-�3:J@zF�L�R�X^,d;kXq�we~z�������R��������������&�@�X�r��������*;#L)]/n5;�A�G�Q�W�]d`k�q�wO~1�?�N�\�\?be�knqd�p�{��������������� ��2�=�p�{ 	:��"�(�.�5?;aAsG�MVTZ4a�g�m
s�z����������������,�B�X�pť̰�����#�j����3�Wc	o��".(�.�4T;�A�GN!�'*-qc�i�ovM}}��������>�q����>�s��ǫͽ���������������(Z� p'|-�3�9�?�E�KQOXm^�d�j�p�v�|ǂ҈�����&�:�_������Ÿ����� �)�4�?�J�U�`k~����&�,28>(D3J>PIVX\�b�h�n�tz,�<�Q���͙p���ƬҲ޸���[�i�~֋ܠ�������)�6�i�z��
��#B)�/�5_<�B�H�N�TZ`*f>m\sgy�҅�3�>�c�n����o������������#�K������.AY%�+�1�7�=�C�I�OU[,b8hDntm{�������řݟ�`�s�������/�@�M�g�r�������EXs��%	,�3r9�?�E�K�QW-^�d�j�p�v�|@SGI$ORU�����������Ѱ䶟��ĥ˱Ѣ���3���$�1�H���
��##0)q/}5�;�A�G�MTFZf`wf�l�r�x�~�%�7�D�s�����ʯ۵����b͎ӫڿ�#�{���� r����$�*81E7R=_ClIyO�U�[�a�g�m�s�y2Y�d�p�������������м��������"�1�u�����������P����Hq}%�+�1�7�=C!J.PHVU\jb�h�n;t�{��ҋ�W�g�y�����������������#�3�E�\�{������� �'-3#93?CESKcQsW�]�c�i�o69<�CETKNQ(�Z]`�gi�pru|��������îɸ�������������&�0�:DNXbl#v)�/�5�;�A�G�M�S�Y�_�e�k�q�w
}��(�2�<�F�P�Z�d�n�x��Ō˖Ѡת޴����������� "&,,62@8J>TD^JhPrV|\�b�h�n�t�z��̌֒����������&�0�:�D�N�X�b�l�v������
����"�(�.�4�:�@FLR X*_4e>kHqRw\}f�p�z���������������ʿ�������� �
���(�2�<FPZdnx%�+�1�7�=�C�I�A'&                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                          �������<$f��f��,���   ��D$`�t$<�E ���d$H�؂����$��4$f���f���1  �T  �D$��  h#n}����d  �EP�d$0��  �h�URs�t$�E �4$��d$�}����d$P�x  `f�L$f�E �D$X`��d$D�Y���f�$����D$$`�t$D�E ��d$L�<�����f��(ƋU �؈�������`6�`�  ���4��)  f��@O��`�E T�d$(������/   �$�t$0�E �f�D$���$�d$8�  ��  �4$�E�g  �l$�\$��D$�4$�$�`�\$(f�D$���d$(�  ��D$�K  f����f����0؜���4$��h'���������`�l$ �  �����`�D$Q�E �`���d$L�F���`�E �`�$�6� V�E �$�$$�d$H��
  �ꜜ�U��D$�E���D$4�  h���E heQr�D$� �`��E �D$��d$4�
  �\$ �Q�$�D$�d$(��  f�ϝ��|$(f�ދt$,��4$�t$4���d$<�w
  f���ĉ�f������f��f�Ԋ��  ����f��(� ����f����f���f��f�F��f�Q������������f���Q����f��f���(Ü��f�U f��	���˃��  `���f����М�8�hT9�20�f������f�f9����7���f=z��*h���d����4$��  �C  U�l$�Y   h���f-����<nf���f)����  ������f��f����U ����������f��_�|������<$��f����  ���������  �f������=  ��  f���E ������U�  ��D$0�$���   T�\$(�4$�$���d$,�  �U W�1  �����$$��D$�  P`�����`��D$ �l  �И�E `f�$qk`d� h;� ЉE �|$Q�$�d$H�  `�D$���ЉL$��E�4$�j����	  f�E �D$��$�O�W�d$�R  �4$����  `�4$�U�  ���  ��f��`fE�������ԍ��0ȡ�  f�W�4$Vf�T$�d$D��  �  ��   1f�҈E f�0��U��~��`��4$��D$@�8Ü�\$@���f��f���W��P����C~���  ��  ���E  ��� V�U��  ��  ��z��f����f�E f�����Mf���!  �  �;  �E ����̓�� E�  �t$<�E �hT0��d$H�c}���!{���:���W�`�����8��$k�t$4�W�oh �(Z8�8���М�����(z���ʋE f��f�ыU�����  �  ������}  ��D$�$�`�=	  f���E ��f���f�Uf��f9䜃��*������}  �6�`���D$z�d$8�~  �E f�������`�d$$��  ��f6� �  �t$0�E f�$��D$���d$8�=  �f���    �E ��U�  �  f��f��/��f��k  `f)؀����f��f���4$`f���<$f��f����{��f�E�D$ǜ����f�d$`�\$4�f�<$�t$�d$<������d$P��  h�|���$ǜ�$`��t$$�E W�d$,�  �b  f��E������E  ���݊Mf�����`�����4$f�E��������D$,�)�������d$0���������$���������  ��D$$`�\$@�D$��7
�$.f�<$�d$@�B���8�`f�|$-&��[������$��������f����`1�f���{  �$��4$f�����f���   UT�d$��  �Յf��1���  ��C�E[1�U ��`�E�
  �f��f���U ��f�E S��̃�`�t$��f!E�l  �  �f�E h�!FRT�d$8�F  ���D$$6�f�$�t`�D$%��d$D�%  @�E ��f)�f�f�U��
  �f-�Ĝ�f)����$�  ��-�����P�{��h*cY����x����,$f�$U�D$�f�E���D$h�T��t$�E �f�$S�4$�d$��y���h  ���d$�R   �����q	  ��f���O@��f��)�f��f��0�f�����E����֐Yf��)���v��f����f�E �  f�E h(8o�d$P�ey�����P&��4$`��t$�d$0�  �Q`�f�Ʊ�f���m����E �D$�U�d$<�&y��f�ËE f�ԊM���������`���4$�E�4$f�$�D$���D$$��y���'w����E �f�׋U`�a���������4$h���	  ��R��x�����F��h����t$��dz��f������1��@���-&��[hV�5f��
`�  �����f��
�f��f���f����f������f��fʍ��N&��<f�֋��`���,$�|$U�U `�d$D�%x���� ���<Z�U 0��؊E�<��Ƴ������������f�E h�bo�d$4��w��f�D$f�E �$$R���d$�  ����  �  ��  ������_  f��Q�U f���7�ЋE�4$��  �t$<�E V�f�D$v��t$�d$L�~w����#O �m�.�f�����������f������v����D$<�����t$�E �t$�d$�  `�l$�����Ę������f�E ��d$�w���������t$8�E ��t$�L$�d$D��   ������<$�,$hVG	�V��D$�$`�\$ �h�|I��D$���d$,�����f������M����  �4$f�D$~y�f����������2  ��f���  �x����~  N������f���l$�����f���   �̉�of��f��f����f������f��u ��f�ي � �������f����f�����u�
f������f��������������f��f�� ��ʍ�(��f���������  �����Z���h�q��`�l$ P�<$�
  f��L���`�u��U�,$VP`��D$$�������{  ����`�������� �����f�E��������؃�h�z����4$�4$P�4���h�SE[�F�����`��D$ ��t$$�E �d$��d$�d$,������f�m Q�d$�u����D$0��'  ����,�f��h'���4���9  f��f	�f��j  ���  �$f�Ef�$h!ղ��D$�\
��D$�$  8Ĉ$��`1������f�1����T$(�d$,`�hD��B�t$S�M R�d$4�  �2  :�q���b���f��������$���D$f�$C��t$�E ��d$�5t���  �M�������7f�U f��h����8�f��f�E��Xf�M8�������"����4$f�$u��q���d$,����������`f��h�@��d$(��  0��f��f�������;����t����Ѓ��t$�  h�gHQF�  ��`��������1���1�f�ЋT$0�z���������!�������`��4$�����f6� �  �����T ���������hF��&�f�$F�t$Th���f�E ���d$L�s��`����(��t$�  �D����f�E �,$��$$�t$�d$P�����4$����f���f�����T���f� �4$f�E �D$tV�$�8g,�d$8�����Kr���r����E ���4$��`���������է�E  �f��8��U���Mh6���4$�������������  ��D$0�`���`�������s���$�D$3�\$��d$ �<����`�$�l$ ����f�E�  `U�l$ `���D$@�,  �E ��d$��q�������f��f�E f9������ъM��!U�4$�����8����4$�$�  f)��$�`��P����t$�f�D$��f�������h���fʀ���f��f������ ��f����n��R���$�o���$G�$���d$�E �D$K�l$�$f�$�d$P�Cq���t$��t$W`�d$<��������f��(��f���f��f��f������f��
��f�Ff����f����f��f��	�������(�f��f���   0��D$@f9��������   ����`�E�4$�$�q�������D$$�n����d$�`����������f�E �$�d$D�vp���$F���f��'���\$��f���1É$�$����`o��������4�`f�Ü��o��f�D$�����D$������f�U hJ��E���N����Om��f�$��,$�u`�U��7���� n������������t$,�E V��d$8��o����4$�t$@�E h쩄�hO�˙��t$�d$P�o���������Z�������]?f���f��Xf!�_��[f�ݝf��]h��-��t$� �t$ �E P�d$(�jo��������`f���D$��$�d$,����8�` ������f�E �4$�$�$��mQ�d$�%o���\$��D$,�m��'���g���8̄��<�����������;���������������9��������D$8�h����n�� �f���蜍d$�������hz�K�4$�4$�t$�E f�L$�d$�n�������5m��`��k���n��`������ɜ0ڋU �Ń�f����f��)��d$��8�f��f���
V`���$������f��ŉ�h�Cg�����   ��d$,��  h���?�d$������Uhd����T$f����*�ʄ��M��������f�f�����I  �����\$@��d$D������|$�4$�E f�<$�d$T�m���t$4�E �f�L$�d$<�m���hd�w�����V��������D$$��$�Z������ĉ�Ј��T��0�����<ٜf)؜`�o  ������/����$���  �/���`����������#�A �`WA����  8���E ��+���Ğ�Uh=�&���l���������0�h	��f�f9���t������4$�  f��f���f�U���Hh� 2���h��L ����P���`�����f�D$��4�f�D$��� ���`�l$�-���h���"�D$e�t$8�E ���4$�$Ǎd$H�vl�����h;�Af��h���xf�4$`f�E�H  �������h��"��_k��f�$Z[���y����k��1(蟋E ����f����U��2�M��i���������T�t$�\$h����&�T�t$`��d$<���������T$�E �D$�f�D$�f�D$���d$P��k������|  f��f�U�    �4$f�E�`��D$4�$�����������h��(�������������`�`�d$@�$���h�\`���f��1�f�$�ߋ|$��t$f�D$������������i��`�l$�\$��D$�%�����d$������W�T$f���|����V��D$0�j����E�t$R��D$4�����f�����k���^�aI�fԍ�C�h��Zߍi�h��WO�aI�fԍh�f��W�ZߍW%�jb�aI�fԍ����&�貍h�cR�WO�aI�fԍWO�h�e��h�d!�l�aI�fԍ�2�����C�i�_�d��aI�fԍk`�e��Z��Z��鍍l�aI�fԍe��_�X��aލi9�bs�aI�fԍk`�cR�P'�辍d��X��aI�fԍjb�d��P��a��W�W%�aI�fԍaލ�C�h��b��it�XO�aI�fԍd��k�V��g��a��g��aI�fԍbs�_�Y�X���C��C�aI�fԍbs�\\�Y�g��辍X��aI�fԍb��d��P��Z��cR�g��aI�fԍ[čk��&�P��V��d!�aI�fԍP'�b��XO�_�aލP'�W%�k�it�h�ZߍX��ZߍcR�f9�i9�jb�WO�k`�^5�貍bs�XO�^�h��it�^5�g��貍h�^5����aލWO�X��a��i9�d!�g��i9�b��PY�k`�辍XO�Y�b��d��f��P'�WO�^5�b��^�P��XO�X��V��l�[č�&�k`�h��d!�f9�辍it�WO�h��f��b��ZߍP��h�X��bs�cR�e��jb�l�h�V��^5�鍍h��WO�b��g���2�cR�it����k`�cR�cR�b��[čaލaލd��d��X��k`�i�h��鍍W�XO�f�d��a��鍍jb�d!�cR�\\�g��f9�d��^5�X��aލaލk`�k`�a��辍bs�a��it�g��b�������f����������z����f��`hkb�f�U�������\$(f�t$�$eh��A-�d$,������������D$�����+����c��f�<$��D$(��t$,�E h:wߜ�d$8�if���E�y����>   f���\�f�1T��S`�l$�-����k����$R��������UP�$$`��D$ �K�����҄��!�`�E�O�����w���#��w`JB����w���*��wJ k���w���ee�wZ����Y�wb\���Y�w^�b��Y�w`����X�w]�,)��X�wc��6�&X�w`�(��[�w[�0'�][�wb�T��;[�w\�����Z�wa��!�|Z�w^�w��]�w]$����]�w`��"�]�w\ /��\�wale�T\�wc�<�3\�w^��{��_�w`�[>�u_�w]<����^�w_~8��^�wd  ��^�w_gpa��Q�wb���RQ�wd����>Q�wd�h�P�wdT���P�w`����S�w]�^��S�wb�xP�S�w]�3��R�w]RPy�_R�w^g_�1R�w`��-��U�wa<a��~U�w\>z<��T�w\+��T�w\���
T�wc)���W�w^���KW�w^ b��-W�w`t���V�w]R�d�nV�wd�k��i�w\��0��i�wa�� �i�w]f����h�w[����Gh�wc8o6�"h�w]��Z��k�w_)^=�fk�w^<Z{�8k�w]!���j�w]��m�~j�w\�D��m�w^��O��m�wb�р�m�w[ ����l�w_�h��Hl�w[����/l�w`�E���o�w]����`o�w\Q�1��n�w`��y�n�wdBvK� n�wbCВ��a�w[U�Ea�wa㩼�"a�wa�M��`�wd�ߏ�o`�w[q~��c�w[[�+�c�w^�&��{c�wb1����b�w_�X���b�waT2�b�w`�v���e�wdK�����w[�-��]��wacL�:��w[$.����w_J׾�p��w\��5����w\(�?����wc������w[����W��w[��\����w^������w_�f ���?�ED���_I�C8~�b/�n"r���A�O&��L28HpH�~]N�6^�(��4�).�6ѭ����e��f�����\��#���>Ӽ���H�NN�?|O�[s�A/��c������}NE�Ov�S������>�b����3zh��ZX�}LUr{~V�̨Ch��:�H��5�t2e��r��K�Xb�V@+nԂ���#d�n����F��U�M���{� b9�5��f���6Z3��a��S�\��.0��o�Y�Z�Zᆐ/'Tϙ������Y|,*s2��`��W������rs������*�o~���2�t��o�`�wZ�r{ۉ���"�f��Ӝs$'.�t�v�0V*Xn��t$(�P�t$0�4 ���Vf�����NZf���t$�f�$<�t$�  ���6�&\��9��[�$�Y��Ut�j��7M�rdE��*犇Z�|�?�
��[0� �B��U!]����D&��Ֆ�-OU����<���c쟦I����R��=�P�2��h��!+��9xI��'&�Ǌ+�=����9j��8��L"���JPd������M�1=��x_~q g&%-����_��A�|^dcY�Wk����#�����H�e�h�ǱV-PoRj��E�rC�ydO��F��φ�D9��>� P�����=���S���9����T��4������*�UP]���A5�L�3{��u�>W�Vg'E��ϙ����S�_��-yT���+��뜆q\���n+�D'k_7�+�,���`{��o�q:�@��?�.�y�S��,��o��x�Ouz��]�)�짛G��8Y�l�0dR�xR׵�Ea"���'?�OI{�l��jg�{�qM9���kQ[��[�4�6�C���P�L�(|�%Fl�|��v ���vm�?�u4˄X�!�����`�ЎbsB1�k��tw�tHY�9}>�L5���8�]G�SsQƕ�����W̮��;1�I{BmY��/z!��a ���F�+z���h���o�l]ຉ͍�N%ۮ]�����Oܲ�� ��N�D� ^)�n3bNǱ���5�ɔ2o�2�)~������'����Sx|؊�rN I�/�j��3�cO�]�zQ�$����1c�^y��x"A)^����KH�WeğV=�K�C�K�<�������\��Մ�;O���^Q��]D5���Y��*�� ��J�d��k�����X��O�x�OzDxȝ��r�о:�c�&���� ����, ?>5�<���^�VA�˝��lx�ֶ!�OM�5�e՞4�� �^�p6[���U|M��k��ٷ
�ک�2�gv�4��Qi�A��s5�6��Vq�+L��D��әI�e��d����cq!�]�Y���)��䙼��+	T���.�꓇e@� Tv���Y\��N|��!I�9᨟���^����YV��
v�u�뿀���j�.|Q�_�W�u+Ưn"F��C�������
�� ��9��Ց2�Y�Q��TÂ������b��h��7��{=��v��tz��:R�\A�����(^W#��<%0<Y���`�/")����
\�u��wP���bD����,�D)�:�cj��mT2��`V̒϶\P�	�51E8�2�/la`�4���1�28k(����vu��A�,��=BI�G���d�UT�C�J�c���d�K���L��S�'��$唯T���L�clSL��,_t2YX7��ԊO
�617����s�.��$좋y��@�0%���x٠[
� -�����%{)u��D�>6����-Y���x^��?�0�A�/>�R���B�~\j������O�����WO"�+��}={`�bL�E��V41�Vl$�s�p5��f�D3Bq�]��㊋o&L�����A��m������������%~�\��M(Oݢ`�Z3ſ`j��F!گK�*cT���.�:��$�t���+u-8�.9�L{�L��L�&�vj
����|�r_��Rf�<Wd�!+jZ�N�u��e��N���A���D��p�^\�NRf~(KI��~a�Yty�i?~�bsB�
E+�o�:R��B�����S☽Q���<� ��죂*���x~)�S-W"��w܇>a�ͬ+u<S��2[,��W��;O��90��'\S��KVa9���x���2Ms&a�U���f�y�p�ky��<sI����B?Oj�e�ݸG���t{��ؘa�)T�繻�S��G͖���h�t���z��T�`�ap�e����G��{�?wPh@6��r%:���2��	Zxw�h0/h3�ȹQ�A��9�s���N�/��y����KD���sK���%|�}��
�h'p#����'�g��dG⫚������E�1���v�Ez�D�U<�ZH��"�Vt���l���Jy�?>���$:�3�KZ);"����r!�_n="��I.��2��<*>QЧ �Ah����z�($m�T[R<'
�<�c��ZDU\�?nv�Nߘ �G���D~A,bp܂C��g�,Sw� ow]�bi˲dQ$�7�Q�Ja/j��/�|�P������\l�4�}h<�(�+���v:Y�G�3�6�/V�4����8pʔ�dS�]4TN�
�V@ ?@��$-�g�M�\��p��e/E[���4���>�)	�{7T�u���ǐ'�:nH��}��P��p�I�;�<h��:R��XW
l���S1:J$�C\O��B����4,ђdGn����m#L3�n�WV�q�8�2T�p��q�s:Ӝ׮�E�U�@h=J7�z�6Qz���B�? k$�΋Xѭ\P�� 5������״}b�,�..��� LC��/"�ܤ�Tgp���\+���
�ޭ�S"2�.<�h^�@Nd"�?�=��`�"m�o�o�<�j�b��S��`��4ʌ�cZe���0t��� *	H!�����!�Ц�B���BH�l����ˊ��_�L
8���(�{���WE�Nv��i]X'���u}�Jp#�S
�9�7O��gQ��U л���7L"w:�l)���6Ⱟ�iO���F�f�z����r4�y�I�m�q�ߔ�_�S���b�H�>�l*/>��P��������v7�/9*�� �s���i��j��n	@)�_�.=�_Z�f[��.����z���{���+#\��zD.�FBbV$���ﮍ=���Uӹ��;i�]{�a�Q?��-����R��-���e��b�0���^�(�ʱ������������vWB���Dٹh��-!b�Dg�y�82��(7�K���-~�2�^i;H��:�U�����D$E�8��T��k<X�9��XN�fy�C-�Y8�X�Yr���耍���j��21��Y��6'갱D����4�gG1�TG�WE]:��D�{�����bE�xz�}6�L���@*��Ze���r� �����l6�2��L�2Hw����+�pp��2�Z�0��m$�
oJ�q&3/�V��]�j/I,��?�+r-�,U�d��8���/�"Ma|X��uI�
C�@�v싉�fk��_4I�w��,c�}��	��L��=�P31�Ƅ��;?�C�h,+38�-!���P���0����m��0ӌT $O�������С���G��moSp�y9�_�$���5�"Y��*>��Ȁ����ə/�_'�6��W�5{j�w�[�1a0�{g����!eW���Q��L��w�4+�q~�]e�|�0�0 ��#�(���h�`;�q�'%���{q�{)�l[��x�6}�,xl�X�b�,{��b�i�/��.-'�M5S�q�)����V<���DkR�$��^\�m=)(W���Ki�~�u]n��>����+�����A�	�o��F��1(XV��n.�-����Ugc	���-����Na��Clü��MI^-Lk��9�V����V�J�bϼ�Uq�Ⱦ��1��|�~�p�*���Y,�m�x�3`qa^�����Or�Je��m�]1 �!uD���ϼ���En(B]��T�c�y�H�Ȍ��G�tWn��Zg.=	VI���}J5���B�Ȱ��f���I��܇M,�Ek,� '�1�6��(F�r(��2(�����u�L��;��-,�j�`x��U~���i�z����S�I���~V�ց|�&./q��.ꅜ`d�ۧ�N��6���HgM@6ma�Z��y�aD[��9S4���_��c1`@m�9�+�_^��B&�0�ލ��S������^���QT��ٽ�7y �~uLZqHQ��?*0ޜФ��0T���Ѭ�]�3�#�z�<�M�R-�3ǅ��T���*f�{�ј�I{�/�\�SPǪk�+���A�h�8�P֛jC�v�8(m~�ڴ5�y|+�g�$�s��BT��xk���PC�<V�j�D�T_�gH?�8�Jl H�Y���8ب��i���J7r�램������!2]g���(�A%��o6YgO�6Nݛn���K��dA_����?X�q^m'*VJ�po�:� ���vVE�8��E2��FY�=��8y�n��D�����7}�H�ޕ^���.���|��C���[�S>!��V��ɒ>���Kp%�k�)��9�N�9<�'w�^w
U�hS6�M ���4�X(Vd������?��2��[�w�ed����h'�:Й�m�0���aO�o�����H<�f7�����|�N$�g�,��^l	��q��4l�:�C��e.��t�.�Z�(��5D4K��R��Q��(sfmV5:ڛ�iO��9B��P�7x��'O�s��۩P,~�K7�!����@����r�۽ �}�dS9���C; ���)�|ߪ��FZ�tA�]>�yt�{�k�B��*VY;5ҿ٭����PkF7�B�|_v��J�h6���������=��y�!BQ��7j�6�[r<g*rI�n[�Ș�'t������P�8q�<��¥��K��I��	e��[}kf�N��ot��c�]�	���C[�T�Q�A[H�z��EI:ɤ/�P���砠�|߂��G�� ��޲��p��׎9���#"� N"�{������ID݂8�7��4ֳc�@�|�7Tg�E�[�i�Z���d1dн���&[CD\�\�H��[��Z=��JhXn<� �|*h����D$����W�������t$�  ��򩘮�����/�N��� oLG�h��-���T'&e�5C�H`������R�pǀ���t$��|$`�t$0�4 p�Bu�c�F�������I�@ϵye���/���ă����F��j?�4F�@L���(# -��k�)�OJ���M��@V��
��y�J%���>�V��]�c��1*�D�zS}Q9Z&��i���λؾa�D���KAˮז�Ż�n\}UF�B���(�{�6�'�d��H��Vm��?��/�����݉��ddE�*�߉Ը��Z;�F��=�'�LȚ�Ѓ�g������Q�7�8���R�#�����ɓH��MZҠ(������A߻`��j��}�7ІC;�ks�O����ܭ ��s�0D*�i�:d�%*���(!8{���_�8��	��d�����L}>��R�!i�mWػŖ����2���V�l�!��ν#QG�#�'%�ǅo�ۀ�(��UT��<��E���!",��bCj�R�	H䙠��Kڑ8`��E	��6u8���O��+��٫��|s��3���њ��n�4�e�mڝ�"� m��eĐ8�y���fx���T�>E=�(O��ʹ��s��\��}�_�K9'Mnx鑖�K�:����!��
��P`eܔ5�;�=��O��Q�n��gv����Q���1�	Q�0�A���Z���7 �!��UF���P�8s�2S�h����p^s���ƁKD&���"��!�R��gV>���3��}��A�, �@��(8�o"V�H��<}��V�o�՚7� Q"g%�7�Eh�p�{s\=X�ܫ%�m0	���)�]�����f��3��"��_��8ᨗ*�
�X7��,?QϊQ��2 �P�YY9R�1�nu�v������|��^��r>�,�WĭD�Ex�c�M��WoJa��36o�k~�R��~�5�����[�����Qe�~�c ��?����E����:�ũ��!�_u�Rlu�&���>�&�[P�t�S`��MQ��]~ '�����YfE�&
�������(vt)�-���q�����KH+h���a����.���f0��=��c��LM�a��&罴��aM�Š_�q�j������G�pa������M������.����B�|� v�1p�n�yM8Ihd�k*�_�6uװb�ȏ��[�����Ћ6,���\{F��ns�(�q�H��8��8�_���@�i�L��D��L�χH�;l���<��K)�^}��y~4�.��(5��OZ�jjm�Ph��(�lK	�ʻ6 �v�_B�����z���LN��ܳ/9M�d.�������\�1����F����ɱb�{+u��v[<��T���k�������/4�^2Y�$��u�����g3 F����o���7ZCl�ጞ��&ֵ��,#�Z�K����gf�������-ĽCe���P#��fA-A4{7��j�9ϴC�p5�bJ���A	�]�YH��-��o���
�*�ʸ;,W:�0?��c�^��$T�����'(���n{Ɗ�(�D:d�e��XYc�q�Z�<���Z�6�!h�ƾ�ŀ+���5� �}�>߰�͉��������%��R�����q��ِ&���϶��I��գ�wś���y������Q�t$Q�ù�g�����lG`9�����!�H  �u�+�9����2s�-�,roL��Pal{���g'��"g�5by��:��H��s�˚~�8��2
��$��֌F�RۊU�W�Qt�a"���T�E���Wz�2o�����{�<)�N�'�pq��m(�Qo����qȘ��$�V�?���QҳMM�7���m��,D��t(��ƅhOE!�>կJ_T'"9�kw�L��[���VZ7�b0���R2>no}/{D��Ѳ�.�rL �$�������6̽��=X{�~�;7��g�<�(��*��+����J�W���~�xw�>����-�la���?g�})���4?�Q4-DB�oxW�#5�M88��t�����f���IŻq��i�-8���w�V�$��t$A`P���Z!f����U�1�P���D�_�f���5s������ș"��v�t$,�h����$��t$4�8 ~�t���hw6E���c�?5��ޭ5+dޥ��Qg`i�/7�Z���=С�o��/���-�+@(<R�t���}>L��fM���C�Ɉi�<�`��z���j��g__e1TZ��/4���$��P�Ƶ˫ RO�Q
�����p���Z-r�'�OI��9�<���Z@H�q�X��2����Y���s� ��S�0��Bo��!��#�&�V�� ����|k[����`��&�gʁ�X�n`/T��ʍ���P�Zo�&/z��h����K��#7�c\!�f�\�{��Ú_���9We�k�-����s�;4{���鷫��j?g8+b��Wni@>��-bN��WZ\�n���]
����[S���n�����d�&�<�H�+ݒq�{��m\��ZBa(�B��5c!'U	e�)4gN���r�8��%$��&���1'�ʁ@��Z�于�~��)�s�g���y�{I�ˢ}Y��j�ʛ��^C���b����;�=�qu��nN)�������������X�����B�@����m���u���<�V�fEd}¯ ���1c����|�V	kIm�vLjy	l�uN��ٗ��������V�5����j��g��}���LX�uH���8N��[bLԾ�@b�Qr�]����!5,��/Jj�`�T��"��e���߭��z�-~H��"���V/by�Ӣ�?'35�yҖ�)�������%p��d��ndJ���Ndf�v{]gzqn 7�D�R���>����YÀO����Qp,��X��m�]����4Ҷ o �UG��̄�7�#�p��B�:��eô�v�;�;k���
,hφ�i��+`x��5:��F]5\�$��yܟ�{���gÉa��Gc#���א`�">��X�1�:t��`�������� �[R��J���e!���_gj�'^ڠ���KU��  q#c��N�^6��l^v�R©���Ļ������X�Kz�jO����k6]w���?�d���p�ƱPȠ�.��.�C'Nrkr�o0�}hSio�4��D�8�x�xc�������"Ȯ<�6$��m��Ϲ^%��[2Z�s��[C�ǽ��zQ�w�ռ�YRB��?�b,��Y��q��P%���#b���bS����-&+rVa��>�mz����)��P%RqM�~�5�9��l.7ƝGj �:�4���qt��ħ�,q�� ��F�=�\bJwaP�1�ۊV�ށ�+4������>�s>A䓳"m��ɗ� �s��$�M��^�������l�7���]�z��YX��d�0�	j�X������l�G���q9hJ)��3�	��E�i�œGe�o���D["!8W��&�̆@a�:��������#���T�e�e�&W�<� Y|��+G��Ȍ!��ǃ���X$� �z��9~uB<�˜����1��ὸWkd��^@5O:o�V� �ak<�[�=+�d���3e�&�v?~9��V�~$���ĳB�9�H���B	4Uh���B�Q�*�4��Xa�A���J-_r^����/��^��5)D����BZ�:R]����3%2�x��z�Ӳp���f�k���d���y�(��!ȟE������.�rp���x�d^��R ԍ a@���jc�Cs�{���`��t�¡؟�����\u��m��i,����!�. M��;%�?X��7�_�1`�_ch�C�dr��>m�����Q+-j炻RePG1>�f��|��hr~�CI2/����v�3�;����h�iôLkb��7r���]��頺@�xG�(?@J�:
�/P��)����uo<��W���÷�:J;%6Ž�F�����H�Ӳ��Rp�7\��0��$ ��=�ПU�����F��G�O*#Z�($A ��W�����$��،[W<���H'Ō�BA������9���զ��lE�B�*s�z?B*5-&?�cO2~��m4�ӯ��a�����-wO�|]�ٱw}V�z�*p�e3�=*�����@pG�xbM�r�H��}�3�0%$�V��>y��w�}4׿�����$h��^���G$"�
�8����1N0�h�8B�[4����E�
�P���o���yo5Sy���w����',LmI�x�i�Dc
��<�Z�]o�s*|j~E9R����c�5>��#�݉�"Q[����t�};1�A>M|6A���M�/�:��4�o&
Z
+*����g:9Kr|��B�-��(�S'�h6R���7�k�8/��]��s����bzIē3�7$�rѡ}43����S�?>#��F!П�T�J���>m|Ռ��)�A|�&/���@�%�t�w�l�>=ν�gN�E�l����+f�I�Wyϼ�8D���%s��P�]|���������lH^k�������&�w45�N&�X�3��>=��%,�R7ݐ��Tl��ר&�e���)Z����
�0�%LZ�����Qk�lj�����0Q��e���/zEO�2^��K��)����`D��a�G�5:�"��h׳s;2�2�w b�)g�����;�4Vt�5߉&�Q�+FUC^��#t��p�Ԓ"�;fC�n����oQ�%�f��:�M\��3Գ��'���L;�`���;�K�B��&�M���;,��Y-hZ.%��hXU�����Ɠ+�:y�E��L�J�D��~B��Y$�7S�P��􇄏bq������#��Pڑ��V�4s����mp�+��A��`��C�G�%c�&&$���ʳ�I��z��ˈ�������/�����K������b�^�$=X�%����h�r��α��?�,��Ydq��0�����kS�=�D,Oi�n}���(�C�]�DQ�F����W�Cqg5�/�]s���͝�}�����"�����|�Vdk�!x'�]�m���u$c<�ӏ��*�;��7��Uެ'��h�s'�v��?f.̶��r0��
�刭.*q��ޒd�$h_N�J�Y�X�e׳d�}�~����y�dc����z�nt��6L�y���<e|�e'�Dh97>?J
�Կ*,u�
Q�� T�����W�ts������jsPH�c�'!�~Y���ܥܵ	8�T�A/"h6��T��Dg�_̬�.�����g�Q�-�u��Ȅ�����Y�)�����􂨔��M�մ�� L��meU�Q{�ę�(�~Cӽj=�}auNUT�MW�Vpc��|�"�h��I|(qx�,i�K��K�Zo~=��������M�ìk#��ڢ�'���s����[񇅃�W�3.�����Ц��FS�KΩ�RB����]4�QP���x��%kd�;/a�el�q����
s��w���d�y���yp�_�D{S���c!�Ib�L�a�~+������F�&a�ǝ�Ѯm�êA�����Y�N���F4G�-�ӂA��K��������7Q� �rC���(ߖ�2���t�MlDL�IƽaU����O��ake?��SY�:E!�P�}�J�F��2l��T�BAU"=���(�8�C��"��yK��_<�x�`,��P�� �Sms�[���I���Q�#z��+d�d�X�o^dY�7?�t��֒hړ4�/x�s>��� �3�Tn�����V�����{~o�[����Z���7�i>KKo���ߨs;Ȝ|ՔI��%�Jr�`�vY���4�a����u��.5ʑ�#ӣxp�<pv4+���/j)@&���/�lO:4в˱�^�Z�!�ej�N�i^#V|/r�]N@�� 0H�f��<Ո~��k	��`X�;7����ȋ��x�~ӹ�G}��A�?/���Ӹl���ؔ���ҋH�̀�Ajƈ��H�D)�%��ȱƖzŲ��?bQ�^�� ��)*�v{�(�jmf���q�u��u%�&;+(���G��ڡ倿+�M��Z�G5�'��y����N���SMI�i��$��Dp�vʿ�O����
��r�;�ci��vv�N�@;����g�P�r����l�P蝥IJ���񘌚l7ӏ�NK�1�?nǗ�Z�gq�fs�ޚ��8*S]�v�`��o�����:O��ڴ��X�S���H��W�/�J�tD������
{��M#f�65���l6/i�tw�u��	��� �X���L��W��v��So�;wXo��Tk�P�j��Ne(G'��_�����U�DÊB����%"�~xuUTp[���V�|Kz�$>2@Ȏ�J��-�=*5�Ѓ1�l��u�NyM�t �o1�>�B�HU�CB���5���ۮ1(�����B�et������TǱ��3�|�$���M��������v�/�ܳ~�)
"kJ�X�W}��t���]0��H�~���R�蠁(��.�5�����ꉖ�FѺ���K���V��*5�7 1����:�Ah��u��A��nU�F��S������v��=�Pn���}ZU�XY�5�EV�b�0W�`�1��S!��2�$C,EO�sf
w�F�^��
�%(i�?|���R3��N�50G�J��f-�Fz_*���V#O��B����W�
��Nn��t�7f���M󜦉� -�~�]�����S���x��oSE�ua�=ZYU��������EH��i�@��Yh�͜o|n��%�Ԩ�?3|�δ�7��tY��>\�ScjXL'FEx��*F�j�[c�H��mp���2)�v��;�y��2Y�@� ^0�iu_$�Hɴ��GĤ�i��/���Ҽ�X[3N��� ��� 7�SI}���&�B1pWf<K!XL���ꆉ�%�7����)�<�iY�^m�@fm:���g��`�W�y}����f;�C.UѶ���pSh}\1E��df�M�r�d�$%:KE�t��*�*����w��5��o�'� 
��7B����1����MW%ҹ,��M�/�3<�L�C��c�̜#��iw�-r���{�B��)IZ������a_���FA����-5Tأ��T���⍻)��2�i�G�k�r��W'6b-hPaX�;� ��ΰ���M����wqA.a��F�e���@h/q(��҈��٦�N=�!n���"�0��Y��VQ �?s�%��z�5�t��z"��� 9]{��ŰId���% W�[~��&��v�����Q\��=N����L񈁦���VT#��x0�/�oFM�3���N����@s����^���<��d��>C.�%�c�>76���b�D��5C�
U��Gs<CY��nS��PY��6��͆��= _8�y�_���?����W@��d�0��-��,�1c��(�6v��oĢ&�W�p�g]�SMm���	g�i�s}BWf�xY���'^=���SѥJ�U���g#Vp�웜�$�x�Rx~DZ�)���(�n���;�vX�Ο辰	��M��as�&�1A:Ko�M���O��`Y��Ry?�-3�X�Ήv�0S��2��W���v�9](>8i
i��������c���������.ž�j�C^e��N���׿0?k��٘a���? �K���,�S��y���ns��%k|�BIL�0l�y�$'6b+:@��3u��ýP΄����7g�[��f�}z;����_wUf���KR�q��?���QNz;/�� �N6��;(�V�0�~�8P0�Q�%�<)|������|����)���E���d�BAҜ�C&э*2T~bm
��.ۃ���{�@?Gn���,�qFe�/&I@C�]����{̢�y�,��pPl����~��x�Yo�>�^fjw��h�ڌ�����]� ��y1=�/�zd��c�2%��! �a
Gι�x��a]H����{��_�u���,]n�Ѐ*�K2�6SȿGr7��LՖ6q{��3�L�t�$GF�["yL{V���4�T�)�n;��Tw,��F��
3=����0�?ܷ�
��<�^�����y�_������5�	o��ҕ�����|�b��޹8��%�?=�v��{r �&o��|�of�9^&�8�	��},��A��ω��������1��8@���4K��f��fu�\����$�Q1Yxsd�gFU�C��U �VY3��t��K�\�/�dRe��{��R������r�{�(!d@5x��r����W��3�	�)��9�p�g����̿����]�*#z�C��
�%�J�@��7�iQ[����������]�=D�]"a�l�|^����E�H�c���T �7�<�aK���ޓ���<��ZS�x���X�\�,,�Dtq���A��G�9�o�=��C�(����|�#�s~�6��S�8�u�t9P�TA/	/����\�E?�=*��ơ@8�F$�]�@V��[:;İW��#�����a ?f�q����f�.��D��&���a����(���9L�{ުU�c?�	̓6
�+����1GL����4*��y65蒦��?g(��9$� ��c�pn��� �9tb��%��)ɧ<��}�[�^�٢��2#Lǭ�9t3�U�ŪKy��TN{g���NJ��wH���ٱ �H��A��~���mif��աF(&�����*o$� �������YԼsb�Z�j�3@��4�϶M:xC2�陼m�)I@���>�)ms�P����*���󦡟����k�]C�6Y�;rr�3�JA�<��)����x����7�^w� �U_����9�Huu�&���#����7.\����~�E�iF�ӵ������[}�&�/�;��W�L��6�$��hW�<C&}��()Oۑ����ȆR�j�_n��L���i�0>V�S��ُnYc���F�fĭ�hw�����i�@ɳĳLU�p��M�O0��~�CVa��f��� ���Ｉ���f��<54o��/�h0�t����j��Z��|C�Wh��n07��T�A��* AR]|�]�`	H<�8$�X�9e�����N]uB�u*J��rCB���iܤ�@�^������߆��N�B���$}�2>�@�s�B_W*z�F�w����T ��)��?����uF�	�V�M��v�ş�{��9��Xs���{���J+뾛Rz��e�4���K�`(G��!��Hڱ2$ǒ�o�}$���F�����	���f�$a ��>��$�������f��f���(�����V����kf���wE  ��ے�x_f���:j��� 6o�]ma����ܙwU��vUL��H�Z��ql�x�[i�O��z�?Nz�g[�ΡL��M�JI������fR}�-���k_��14�Zm�%8�����I[hvU��֪;�M:���?Kؔ���u#d;����.�����'B�-�`ꑀp�0n��f6E�>L���\d�n���!��n����m�! ����Mv2i�BB7� ���u􇂑mR�Q�xVo��	c��F���b��b3b¹:��(s9`5��*��.�H<��E�If_���Cq�ҩM�Kz�[0ۆ&a�T�O��7�,HWWN2�l�4�t�w����`_Ʃ$3�}Ec��j���͘�V�tK��J}g���P�E���.c��)Ha �BqY����?�+a_�)��j(�<{��(�:s΍��91R\�P6�NQ�oG����(�Q��d�R
{��A�_w��X�LUl	��
���<O;�5���u���?��u
W��HuS��YJ/V}y������9�y�~����|�B��86�`���-�["Q���т�::�o5����_4+�uܓ��0�F�O�s�M������%n�=�%׊#Y�ͺ�/�)4�Ӎb�j4�\�b�����$�f']w�m@Sscu`"��_/&��nڿ@p}�h�w	خ�}]�����Lp1 ���|h�wfGU��ng�V�o��^ /!�9��k7^t`�V��?���?�*�!D��6��io�of��8ҍ�9-ļE}�ӔfϘM�h�p��-�)��[���*�^Ĵ8~ũ�����H���tv�Ԟ�7Bh���\O�F�- �����q�����Ĩ6I�>��F��9�P !����#Kt��_X���5��'mc�{}�h�3�sW�C�{��G=���[9�e����0�}�ӧ+I��>����=/��]�߆C�a�Q|ypGo5;z�[���0��;�{��0O�-�&C#���7�gi���. o&d���Ah˚#���@����ax���Pq�
�����R���p���>(��D�U֍C�k.P)���B�Ŭ�3ez���o�u�c�n�ƒ���Z�U�JﮧZ�(��F4=I��Y|7��]s)�!�=��GE��g��I�g�휜�$���Y��,�������3��@K�A�hi@�����
��W����L9�Qxc1	�C����9
,�l��,�뙎4�\qm�%kN�>�ϭ"��kҜL���5\L�jP��lox�VDÖM�V0���Wvܪ(lrȎ� .B���~Ϲ^=�h�#�?�"�k�CkP���Gƅ@�����#�ߜQ��=��opI�5��-A4�;o��/����t�=qsx˦������ǐ�� �9�:�815��>6�/
�� �#��F0��M���j��tz`ͭ8�X���Et__SSS����*!���/�퐚+nXCN|��#�|T��Ck��ڋ�eTK
AH����ű�8�������sX���f�3��s������κ]J����^}��CFIU��}O��ru�����~K������YLPtFI5�1_�L/\��Q�l�d?AK���<��q��W��l�g ��&UN���|y&�Œ���I����;����t[�V,����d�����O:n�/�z��T��O`0>�2�*�
].R9Q�K<$o�������~tE��Alo�fr
j���I�?�7�L����v�\�`u��X�aV� �t�ǰ>�w#	�(��^�l�D\�F�|M+�)Uxe`?�4��5�N� fu�GD;��=ISN��~���9ä����Ch]����.�%�����&�<j��zӵCꏞnG�=\]v�jå�G�O�n��ڀ	�2�T��-Œđ�OV�Z�&;y��P����pS�L�Ww'\_�rk�EtS�� �E�����������6�wZG��d�Fh���}�F�=�F^��0�t���Ӎ����x^
퐺��"��N]l�sd�2[��05�C�D���� �w������t�M"�+j(K��'���Ue���u	 okV0uI�<c7��#o�D1�N�����^�r��������%����a��u\TJ�B�>2sN�WL��'��2�`�N�;�p���9@����qS�t�_�O /c��B�'eի{���%�x�J3�m6��a|s�HK����"�d�ú�(�V� �b#4�<ͣ�ލR�5t5Z�����tL�z�8t��h�uk!�dp�؈�ł�%bm¯.�^� n��/r��ǵ ;�� ���BA��O��i��M������&�H�bn���2PTu}'�
���߾�Xq�r��i�:Ѯ#�i~��Z���Ia���I�9����Hb���M�Njqb�ߕ��V�
l���C�E�_9��P��թ��E�'��?Ak襥t27*���%�׮����]�i�e;i�U� �Fsx0�I�j�i�t|x0�*Y �J9���=�:��E��Ao��;ę���w��٪���j���e(�v�l�p�t[���A$�����hvD2(&�(N���s  #���q~���_)ڢS	�~�5#�>��7.�,+R���v5k!]j�'�v�#����b����Ib�O�^�k���8{Q��g8�Y"�k��-r�348�3��Aj+�]��m�����B.���dq�R�q�F� e�p�k��ۅ�d���l��9��(�fv��mRQ]�G�3�d],�Ţ����&0[9�1|5F%�3f�agUPX��G͠���LFc�4S:ɍuϳ�|0�1���Nת�VP�Qh��$Ul�ҚW��fq8�d�t?��1�A��l��0�[�*��I�0'��l�Cf����!�����f��/�������|�n=F�t����6��9�J��O�ſo6�mTDq>�NIX覼2Xn�"�ޔ�p��B~vE��rL�On�l�*I��E�X�� �����̓�K`����?����&��
����!�V���-�9�0o�`)������\6L?�P�
�i3c�9�+}�Z8x�h#�*��x��G��A�R�Jyp�>=X����I�b���ζw�-j4L�����Bůh�i;�U�Ǔf�#���4��5�Y{��0�,;��q��]��&��u:�Ǎ���A]�2��%gI�46����/��m~�O˂1����jyp��R�@�(�x	��k�	V���yf̍���h��M��>�-Q���@g^�db"�,�Ug�x�.�jwz[t������� )�����ăp�s�W��5,&�v5�|��KF U�t��x�.�suH�	�-XMņ�o�m�w���c�7s�|�#�ٮ&�ΤV�=���'���GJ�j�Ͳ��}\6��s�i2�_�|�#r+e�`I��x���rMw���/�2UB/�M���W&c�U�t��	���?��ᗴ�(��<����Ŋ▙|����^�Z�v��p��2�hZ�]�e���ޔd�B�Rѳ��q��_;�����!,����m| ���uĻ�E��R-ܾ���sL�S���ɒE~�h����;W��F�E��lG�J��I����Du���r��%~�!�Hb��e睝��>l�t��9Nc[:����ϊXC��c�g}='��p��1���X������+iL��LBl�+A�q�~FX0���rUA�x� ������uV���ݖ՘������f�j�CH@儽K�s���� ���5t/�V� ���Ɇ�)QܓW��溷"�!Xa&�i��:� p�J5q���c��F�jvR�kP�7
�n�	����C�_�
b��Q~W����Gұf���;��]�5�Ƭ�j6{�����ȿ���2&qG�gD9ֈ�b���
��X��'��q�d�����+J+�,���W�Y�/6����el;^��Q�G�(�y���j��������}�N��,cc�[��L�K@�{0!V���32m�
ۂ�B��a\�����gP���Kv� �B�E�A�~«�>,�=�7p{��ul� M/���sL�E�+n�+�~C(��?�Rd�;�	[4Ñ�I{-�5X+d_���.��sʔ�F���쇃�_�7<��h���2��/��=r���:'�������(gh��2�!��ס��epA�J�m#?�F��q�0�jH�5�Tӧ��3�(5�k��6}
3�Y|.�1���tɄ���7�$c/��	x�%�F�L5�	^�e��>/_L���󳨆�7���BCam�`�Q"�(u��ya6q���/�*[E�}��f���s���i#f�[ɺ�g�^��P���M>-�/�a����oS��!�.	Y�^����0�egD;2�T�4	5�сjvn���ё̽A�Ƅ���"䏙<�4n���"t������^������(A%>�-�Ͱ� N����'A���.퀌G�}�6'-�N�K;LV�����-p�]�	Y�G��1���$�M�U:=�Xs4�<V��t "��j��;SB�Ya��Ӥ���j����i�n �6q	���u$�׷x�����5y��u� N����M.F�C�3tlfF��7��0�G)P7������f�4��!�%�
�ωV���[`�ԚQ�GnM$�k2Ώ�2�O%�HK�3�g�����i\|�����N�u=x�a�w��U���� ���ek@����mmk�S�\����-*�D1a�.���e�$�F��,%�Ϡ�\�N��/�\��x�eՠ�,�a��h�rݺT�WG�
����yB�>�\�'�t5g�|_&y�:�(��g�qЈ���#cy�C!6-l{z��.�ȟ>}{�s3��/w���G^��s���O��"��{��p9�J��Y����zFę��]k8@+-�n����H���^K�T� 璤y�rr_T�n=dO��冥�6�;�`W{���\݀���/���v�V����8����R��^VU��Y�~L��S���gl� Z_>I�VcS��� -���71)����Z)��-�l�*����a~d��TJ&Ʉc	E��7�#b.w��_m+�/�c�>�7OY�AQ,��Y�(����X/w]Z�WY�V���������R�♰��<{BѠ��!�T�q}�Sep�6��~�)p [���g)R�5.U+a�.Y�>�P;K��#�笌�@����{�B��#mq� �f��]�L5���|@_�/
7�+�/���\�U|�?F�GN5
K�W��r7�@e�-G�p()$'�����
O��'�����S���4�3V��R��%IBYd��j�@NC�� ����O���s��8왏1��9���ׅQ���)�[���0�m~3����)d��R�~a�d{:�(g-�{�j�dd�W�]�l�(�"�g��95�N�����6����z2���,�#T�[fm]��ZQ��e��-�Tr7���6�!�Ł��Ļ!�Wh_�.���}X��`�-g�ѻ�C?��d[��'�]Z�Ӆ/���5E�8��pg����M\�=�m��v�H�+�$�)4�Y�_�B���.RA�P���[Գ�/jU�	՞͵E�i�c�@̼!$���G����8ˆ�y0�A�B�A�G��G��{���?�L�l����-.}З��Jj�э	t�)����觮ut�z�>\�����̶�M,�I���":�b �R��R���Q�������U������=Q�[;�.'R����Bqy��Px�.gxm�9�;X%{`@�Qp�$6��`GNϼ�tT�y�d+��kuF� �M&���"\r`H�R4J�8��B��_��3J��������	�:�h�����ځ�&Y���\bW����`���K�\��Q�x}S=��`�x�L��Fa���=�E�b��L�^�>|��� z��^��Ļ�Q"7f�<������l�\nOp������������;�}�N�p}[��b'Ժ�O d;*����$Y�5ov���J)�ii��%֫^��
1�����
��K�H[r�'F%�Ҫ�j{* ۅr��S�u
/�9���|z@.���t�N�whd�(w��$P��˩�̜���/�p�5/��F9�������ʾ���I��vic��7���`�:�h��{�iпřw��E�P
��އ���+��2�B���d\g��y\�\�`C����Ϋ�5)J1yB<o��SF1�k�)x���s��p�2��pf -w[��c%f�D�o;�{w]��}�����d{:b�f���/茁�m�a8�BmN�Ζ��i�Т���SRb��cm���l���y�`)���R(�\Z��}�U�q�����	4�^��bF�!h^S���8�����wic6I)�Q
��1����?V�{YgN.<���wd)F�
�_D �sX�`���AV�C������ֽ����\�\0�_��j�YLw?�6�_h��u�z���f��<>�ä��ZT�c|��3]�lYq����Ɋ�1���s�[���I��[��/
S��5���9�Nz�	�_��:I(��;��p�� o�j��(���@GOl-����Pl��鰟���⠶L���t�6 :)�H�n�.D�picy�)� �л��h����r��fR�\%� �m���m��6�c�N�]�rh��Mh��}N~�o��(�h��D�2�D�s��fF9��OŞA#��U�~vr�v�a��� �������6��ಹ��WJ�/R�	��o���,1��^��!�	�SU�'l����y����t�K�Qf���hH"�I4�ryl�����D��U�����?n��s�md���Ɔ>!��ӽ�G�XO-%�H�:�Cc��>�Y�No�-�j�Q������zΙ:���t�5W��<��=v��x��c���f���.��:�x����qǌC�t�{S�rU�m��榙���;:gj)���(�����t-��������o���Xf�>�(��(V���6��h~�}�s����������@W���z��L����q�<N��)�I ��MD�"١��-��]��w�}2���dG�h����������n�gE��6@�U�d�������e��*a=�2��o�B��!���:����"�1��D�=ۂy�r�6q�{�k�פ�W'�H{+V �{rm�>^���iJ��I�7�xǚld5��$��<�z�*�J�}��D�A~)�h�g�r0��G�4Hv�+���*KaL�b*���8}�T��8�/����48x�L�N	�K����^@+	v�Kj��i��:i��k�[�%�\�kt�oo����d	f.`�-O&�%oF������ V�]�R��5��-�i�jђ�߷it�����*�������1Z��� q�,�E)-&E��k�+��n:*��f�r�J|p\M�@�E>W��_���'�8�k
u��5%���{��ǼZ�>�8*ƿ��a�t�_�ߕ{�GqΧ����5��v�8��?�i	���4�NC�Ծc���M�K���Ű�e�jO�/C�I�ﾼ�(���� -��%��E�-eŐ����TU$��������Iu�iP�@淚���A��iC��ņr`A��qć�	D��'n��S��X�я���N$��o0g�p�O�5'�u��Y�>N����*m��(���<$
#�x�]�ٜ;37:]ٻ�9v�Ҹ�\
�^��@�a�ӻ���1h_�u$�c?�G-��'*
	c���1<��a�'���xw�:�~ XK'Н*6�>���V�k�7��.�bdY���5��ڡ�k�&��Xv�TRj��U�!+�0���-�s��XF�F������TS�sv/�����捋-3+)�%�!7=�q-��!�v�4+�����$���q�������T�������ޢ���5�]�X����e)+0���E@N�T����Q[�\��2y>�V�8�5���7L^l� _|�����LG���:��Ot�j��vUL��i�b�V��5n���> ��0<P��-v�Yf���+��4z����:��>q�cst6�0zir��P�6U�dq~Lo���C� ��e��̡��ws�ԑ#ԦD4����w@�{<�md���SQ��}�@����ڶ2[l2��ϋ�)���r�d|JIt����a�k���Z]���-H�Z=Tp�������k�3�+a��..^��v֧�y�śُ�s���)�g��kK)2�q["�"��?	Z9 �N-����8�_<@!�)� �o�6Ɩ��fbX��wF�dkJ��Ne�|M<�rP���a�d@L�Ǟ[o!���(�_����ՃP��}��os��KDQ�a0N��݉rH�Օ��.�Jg���&@yd���߀�\�ohf"���6/�9�:�k`�Z��̫�K0�	�_�4���ۨ��N� �WbS�ɢ��y��4����E���Q�B�+�,��Y�:R�sj�ku�q\�:�ğ��vG�(��|h}��Q�co�Fwa�@�j�	�_w��z�PЀ�#;��pDM����F7���#�/��kBA���a8�kr6r��g����T���C�1[����&��&�O�����ǲAM���rEl3�?��?P?����FZ��^3��s��Z}�y~���O�NL��k<F��p9�xkqw�S��&n�N:���B��`�5�&��H�Q�'�q�pC�D}�3��P��sb�1��7na��	���6��0�����L� >�������'�q0����@*h-ĩ@{1�����y��4�k���&V�x��+ўP����Vhm��49z�V�u�3+ʳ�?���0�/]�k>�k��r���6
�7�����9�\��]�^FAI��!7�tWi�<�;�@WG�?)JI@�WE�Hok�˓�ˇaN\���bh��=���^�e�j{z�F����v˒t[j�~�r�/���"%)u����A��K�}�W�v��(م��<���do�C;�~�%�QX���([�:^�^�a��
g%�:����q�L �;���7��M���jӈ�gha=f@��I6��`��6��1?z��]T����!}��ZY�-�\ɰ���a��� Â۞n�z���"򤉰�&��I�ö��-�q�9���������M���C��%޾�̈D�zaH*��|'�����9�C��Y�cZ�/6h���[�b�~��I��n[ď�b����P=�WR�A��^	�����}G���W�و,iP��~�vD��s<��=�3�,�|��G��0�hxݥI�/PT��Dg�_ɝN�G���o���E@6ӱI�
S~��|��a�/��ݞ�?�����ް��O��뱉�n�t�dih�.b��d�����]��W(8pQ+�?��aM�R��y੦1z}�8���͐I�/3��3vQ2���8�W����s�|W�n`����:�@T���S�fM�� �[H�4q\��3����rC��[t�h�}i����.N;y�l��8����x�:��;�&c��I4��i�0��{���|�W�C^�r�f��:��.}9��l�
�5�/�d<�6w3�C�z*�-���%H�oS��qv�ݑ�ܐMz\��l�_��6#�ϊaM �7�[��*�q(�-���*��x7�Ih�ٱ� r��V���7�]��N�)�2��{;xLED�N����@��I0ۨx��§�ɗ pj�%Z4D�f5�`b�B��KŲ�bv�[e���c5�_�M�ð�������;��7}�lK���ⴂ�Vyq�$���ҫ]}pk�EO���+��4��>(���yW�t���rg*�9(Y�1����"<�s:=���1@�ߴXX�=��
���&2��Z	=�3��<��� _�+�7�P�r��@�� E�9�F��\S�N	3���)��~�
�}O���@���tԎC���P5�#2�EwH�1 ��hcx�K�rQ@�����c4��#w�d�9|Q��S�sb������a<��;�.��3� $����?�i,3a��D6�8��(�hb~"Dt�iݻO|ߪxW�@�2�?�ahKbyπ�� �q�#���tw�$���3[��D�n��A�4���O�N4_ z��ν}��el�ږ��1���z�Է+����ʆ0܎�� �� �_��1<lP�Z�s�=8�u���{K�*"�E�F�n`DQ�P�����~�E�P,�
9k�<�.�7j't�e*�<;�����`z��H?�8�d+�`�Xu~5L+�(\���X7��;��/�p��C23�S �u*�1)v24A1Z)��UC8����c,��;²�m����ԙm~�o&���hPE6a�c��v	��\%��g6����^�0��˟>��@�3��ƍ��AЁ��[�`j�aU&��8�W���1�2���ҁ�����DTn��t$,�Q�t$4�8 5-2f!�����A���� '�8��t$�   ��u�����d��}����\�"�xW�hR=ylG���@��D���lG&~��^�N-��*S��g��)@I�^�����Q�H�qb+��P�ܬ��O 8�`���\�6U��]�3;��'^�Ұ�ˢ�dT�Q�l�Ի�*1���&���	Ϛ�?@�MS��Z�O��S,J��]S�#BwV��]�e�Gz���Q�9��0w���� ����363ˠy������}��� y5��V�f^�oU��ܥ,+�i�i2IfI�oņ�=<�.qdN�ݫ~�ߦB���c��h���_�rX�����>ZJ�\��F��3��.��4��qv��������m񣷆�6����J�t������`��Tz�bK�AFy1�!{+�\,ŃT���%P=���=�Y����.lI����E���p�L��ٔ �`k����U�Q'�CY�]��g��nf!jA��/��Cv�Q�R��N��;�ِ��܃AO����h���)��ɢw��k��}g�h9��>b-F�/�Q�f���K�ɞq1[�4�-��:A�KF�%�)�yr�a����Ɨ�iuR����.6����KXfE�E
��.#'6�>�  ��� 6<
 u��Y�z��D}��C�{�����U
�'�)���9�h�Bؿ7>�!�H�Lw�"��Ж�q$K��P�����;�n��a�:៉��{}z��"�#C��]�e$³M�w$�g�@��;.o	�E�6H��u�����&�3x��G¹POsl�V@��V�T(� j���̚Kl�e�O�6-�O�F��j���������oEA���������(d�wn5s�����`
�'����o��^8�5��f.U�QDQv��c�n������+p 8w�A�8x7�ckj��H�u�/&1r�w
ǽ�1&��}�����J��ԇ���!��o0�y�c��[aT�	k28j�*)�r�d74���%��Kpj��J����'��"�|����=���7e۹'%[����������3Ӣ�ά}MQ퓴-�(��_�]��!Я�Ǜ�n�ߘ��n���w�te��v�|ż���˶	O���"�2�Lq����K��!���_�<��͟4O�_(Mk����#0}�{���Hi������G��i�o�Hd[��7���fl�����ބ��5a��ѨU��t$(�  ����&��鴘�����Ձw������3���4��d|� ���M�7�&��rS6����S䬅D�n����^/�� {�)�7eK�Us�MkA[�4�
Qp�>�ch�%Q/���nIĘi�\�6���b�M>�'*c�k�Os�b��{/SE�]���[�q���ʙ��:���ůT�I�RI�;�%���xN� �<������������]�{��SI�w.v�\׻������K�4�,.e�d��]X���O�Ky�eo�|�b�8��tC��̅U2鐔i�lI;��{O�&t[�35�-�{g�P�U^��VCA-�P�lX=�V���LNǰu��+0���f�
�8ͥ�p[�'�O��F�9��+b����H�,:xtJw��RIP?�~7Q��Ű�Q0 w���>��+�`�G��2���
t�������R�����^!�6���(�j��l�������5=��*W������Et����h�Nܓ���*�~3�*q-v�]�5�y���9#�hI%�ց-i�ޯ?L�2����
�0m�X.��,��6��6�,�W��6�7�&߉>@��챈��(7��X;���c$��2�r���h���WϞ����E<����Q�};9O�s�o���<�����&���|�!��t:���i��q0GG�I޳�wP(Y�X����x>�H��F Z?�0�/L��9 ���6M��t=|i_Y�i�TVf�C%�3�I�Bae��0~d�����Y�e5�~�L`Y��Ⱦp��5]�|��C�2gٞ�	����	��H�e>��P7b�@���5���y�T�����8�_Jn��VW��S݂��(y7���?��A���	\g��f�Y;o]�b���WY��}�F�JE��)%��8s�`3�ʰ�����l����NÃ5n��O�5�c�m�[�5[Z!:=��I�!C�����2}�A�$����^Ml��
<�܋ð��`| �y�|:u��ʊ@��V�$D����J��ܲ�f[�*��B%n��FݳN����`�Pk�Q�'^�R�]oخD�a�B!�# T�k�T�~Q��ؽ�b������,��
$�,K�kv5�*A9��>$��0w�6:!���ԅ�/p��|�ef�	��s�g*~���z���H��8���f�ּ2C?r��;�� 51z�Y������Q����w�T����fu)L��LtY�[�;�G4�� ��<Q��Ym�C�J|n)VF1���Ƣ8D,�!S�G��F�8y��y�\��q����r�&���3�Z��2���g�xiD�䙉2d8�2G����L��C�Z���4�6�[z�zُp3�&,	yM��vV&!s��N�@ba�����
��t����W����������*�S��������Φ��?���Ͽ������GF�N��H��9�N����0�6.����u΅�.;�$���*V�
�� {~=H�Q~i/�M,Psy����v��0������8{r>]A�f�1��ܭc}Td9�{X��`���jU(����,LI�p��r��2h�c���$!m�v��
���u�`t��@�M�:3jQ����J��]D��S�"�	>��Lc���	
4�VL���PJ�۬�`5
�^��f$��h��JQn XJ�@�����Ϊ��n7���#�j;-)�W�"�nF� ���s�������.J�}�`��B�r�ZL���	e���$Y�r����d�Uxw�����n5�lA	'�ί[gbk�҇�pb�ONi8��
���n$G�Yah��(9��~�x[ ���A6�9�q?�fkKKz�D8{�(E4{�"'�,#Ӕ	��]�pޓ�Rj2�_��}�A����^d�4�x�~�9N(�qi��O�<���/{����C�*��"wG����ZHd��v��w��@0X�=T_���?�n�/3�.���dͷG�p�
�: ��s�8CJ�h��ƍ5�-<l���}�|3���*u_���s�t�Q�L����ܧ0�~���ֻ���[�{�G{"(v���vzQ�>��>�ͮ��z�z�ع�;����t�䷡H�tĹ��f�Q�j�֮�^��o�ޜ(09cr57�x�*yC�F�X�H�|�z#�h�Ӕ{���)�:���{SZ��.�|��^��E�w�JE���Qa���t�����۔��(�Li�W��h�x]�}�v�H~؉�r̷A�k[�̚uհ����}���jaeDes�}�=�̊��]a�:2K��'o6�ʹ8��߁�L��B|;I���)�BB]/��jW�=������p����w`����a.��y5*�Y	4�Ͱ�f%�IGݦ�\�lE#YL��s��V2#5�[*G��|H,�
D�\D�dv�_y�mNY�e�EZO���}b�ENSY�H������@}�hJpA�iG�� �j�s�v}���@�o��	�G-�j�r]3nXR^�œ7#�2F	��e�=xw�tː��Tn�?3޹X;�~��(���ڃ�Vn����譑&ED�)�	��cz91���]�K����-���	�ƦQ��AH�d^˩�3/x�Ƶ@���G�Wv� ���KX)@�5R��U8���3���I�ʢ_/߄K�?DsH�$�>�|gP���(�"��_�<��a�������C�{�x��u��oc��}H�aJ	k���7��?�2����UA�n]8n�<���O6.Y��	��t�Sm&����?��c\7�.L���f%�'g�>(N�~�N0(�äc��-���N��䛟)h���e,��8x�)��-l�J�i��G��b�������K���(���@'n����w��ME��h�	��Nx�L?k��
+:|��0�����^�H����]�]�=���3&<6� *��&�tk���k<����H��ݒ �Y"M6��qT�!�8�j�I��r����u��<���K��o�}��`�
'�ٸ� ���q�EnpFU&e]lh�U�QC�p��NFɲ[���]<s0�^�:�JH��˚NG���9`@uF2������a�P��σn��)O�Y��#�#����s�v0��]-|��bq�ߘ�%P�o@�,��;/(g��Y����:�N,
ׇ�f����͍!\���臨�CS	~���A����V\:0%�Z!�2O�w�qx��MD�6X��ғ�O �p
)�"�n
�-�d�{��ǂ����Y�4���k�Sz����#���(�l����>r*8sYH�y�����+�g`x�*�jQ���]״1��9�	[`_6���r@Sg`�w���6-�ndvn@�a%Lo��5�R��E�2Cf,��z����cS*�4��w��G����C���弓K�M��NS���mNAi���,���pN�3)��k�ı��l'�$��H�-��V���r���r18���]d��Y��3�#M�CW6nv+3��Yv{��zqj�-����3Z�-0#-��3���0��b@��r�Ynj��0��Z���r�o5����L΍e)�k̻���U�i�ض�VWn���X�((��X��uL�2��n��k��Q��r���e�4����F߮�Ì1R$�A3ED_,j�l��|�� n�w����"���@ݔ�/�Ά�f�
5�3��S��:�����5��R��Rέ$_�2�Z��� 7�Q�k���~ [%\m_�Fah�n/I��[��wt_� �� �Jm�D�J`W3H-�(���r�l�94���-���/M�Y��<��+^��݄7f,m�]�|^t�}�,q��H�s�ɿgr���2i��U�N��^`Uh�9X���⎡�<�#F�����,�I�הs�1_]�LQeӁ�m��J9��Vz?q8��������!��08=ˤ9�`P�a��pJ3�+���)��'�W�Uv�c7����X����+R*�R����^��*�@��ݴ��MLjH�����vMu���>�zgfh�_!�~��A0d�������h��&�<��>��4r�֖w�e�ydx]��0w)|��n���	���m4���L�X@���$5NŨ3Uj�p��f���V]���BDQP ��jp����-�`�/Qf^a h�4�(�|��48�<��!`W^��b�G?�ٲ<BK1.� ���)��zI �E��iy�"�e���1�I����7�c�o*�ȇ���+j@g��os�ƹ�a���j�U��~�4�j=�^���W�H_=�����ԃ�$�xIFE�L���\c����w1O�W/6x������lvG�?r�߱6G�"2v�O҅3�lh�Ux����K��;Zs����H1��1�yU��ߺ}�\u��򳁢�n������ �5xzG�	��z�&�Y�YoVd��o���r�������Y�������/H�Ĳ)]6~ՠn
aT��;�	�s���ܽ8H|���dT�	�DԌi��[��`�_��Y�|�~�b�P���0�/z�Ӥ��ׁ��޽)r��P��Iv���5�VP���Ar�(�����G��#�M���=P/��2�P����Zr�n��l�Ez���d]�Pɳ��VG��A�kx]�ې9��!�1��ݬ7ɒ��N���[�9��tr���J��Y27�$�x�](G`�����D�d�H�2��&J�R�
����=�-�~�����mL��F��Χ�iƢ;����K?��u�7��BI��pi:���w��H1��P+8ԥ	�v�3%�(����?K�u����d�XCLW#]XI,8��e���7KXfE�E��T#�8/$n�g~�@�LdV�)V��@�;�3P�3�;��RS&D�K�j,�'��q��ňzֹk|�0s>�+U5g����9���Oَ執p�3��O��o9��'���-J�͎�)n��7'8��^ʷkۓ=$5t���5%2H���^�a�
qJ��l��*_���� SG�-��Z�l���'��^�y@��3�bm1 9�P�wD5p46�4V����/�6α�b?����W�k��c�Y	kh��t�\� [�$t	�<�`bl�ܟCSi}�ZÂ|9'"�Va�ΐB���nF[C �4���+���~ �K��vU��[�;p�Af���=��9��*�"u\J�.� �*�W�L'�@���m�S��$��_-��Qb�G���&����w��E�Ӝ�E���9&�#,���7��C�W��_+v�9�;�q"�K� �����/&�Ckdw�2٥*�c����3Ȕ"��.��+�n�:j����MT�Q��S?:�@��Y���8�o�R�����c,pp��|�8�b�m�;��	���r�P�	;5�C[OX�,�b��a$�����2��o"�9R��Lfl��xMD��(Z�I�@���p�V�`�| ��	M]#��$�r�L�:�V1����~�.i:ѝ��9�n��x�[��j`����u�P��E�L���宿Xd-�1LX������M;�Q��
�<[j�pR'
�T������t���7�i4}�"�/��YN��J����G�ة�ԑ1��&n���Q��4+�}�D�s��7d�"�u�0��O4;�u�[7+�"��*3�7Kbƕ�W@�M�e`7���d;��d���G�3-ۿ��q���m�f-����ow>ו$����d������w=�)�h��菇#��]:(ih+t��t$H   9ށ�,N�v��t$H���$��t$P�T ��V:[I�`���&3:������I`/�D�J1�@���켃
.>
y.�O�rk�r�nj>��Пq��=�X��g����!�֜��6�z�F��q�G a�)$/�M����iJC�U$�"��U(|4⨜q��t�"g�?1Z�y�+�	C�MR���5�U	�+q����L�RM��l.�@�.vޑ����K�Nv~�ls �&1B��9;�q�h�H���i�H��!ddM�ZjA���K�v���S�(V���흙䩇n~o#���[�>7U���9��!��?���^�[IY�#�Qh�����o��?â�������@k�l@T������Q��z�L�����^�q]݀V�:�:YwN�]�^_��M��]�ݞm��M�s�fc��ꉈ�V�i�@��	����N��h�T)��֐����ykc;V���Yf�Q��Im8u_�;�|����
_�s�����>=���zӾ�F�8�9�<���gQ�r;�"���ݜ���*1��̝�߄���j[1����P�lx�{��,!�AQPV�������n�6��#B�����b%�j-i�%�Am�d����B%
���_:�Y��g|e<(A����:0��\�,~�i^B�@�F��Y����s�c���ab������%��4S>SGs��n���ZH���[�}�e��~n�l�.A�E��]�G��r�P"��� m@�<�r��J	φm�<H��Sf���|�� )�}�T�=VY��j�P��W�Nz�x�6�i�
�g�SbZ��*�*Ѷ���vP�S�ݠ �uS� v�3�F�*'�\�P��N��y�w=�reu�R�p�l�l��Ǿ�yf�\��s�<�}�Tw���j���l�H�7ArZs�u�����C����8H�;]ԲpA��� i�ɬ��;���&�ݙ��6�ѯ�2�D��b��(���-Z3�3��W�T��x���,��� o�'Z�c	!U�s��FOn���r=���@޲���+����2��T�$�/��}��hT9�k� `/O�3�	t	5SX-T��X��S,�Ly7�@cJ��!rԻ֫�]8�[ e�`��<�����h�J1av�5݁��R%3@�{V �`|�O�e&�_�o�Y��H��2m���bY����]u>�ӕB�͹�_r��4{�}VS�Ѓ�ĺD^��}��Dud�5_<Qe^�jda�7]���S���߮p�C��U�_�ǇG"����	uB���۴3�F��۰㝛���)ah�Q����~�p{,E����!@A��"���J�=����D����1 ��m�O#�h���7�O8H���I�r�2��������ߨ���1�Bf�P��,��O|Ը�!#��+�����M�Ͷ���g��4��F�4.�Q��
i��&�k	R�
��DU�>Q�iI��R�f�l%N'������u�"V�d�n�w�Gi�<�t���.9��Y�6�fCP�+V��w����h k�Ö�y�)L���?n�!�+� ���y2Iox/�I9ui�XL�8��ml�.��g�A�>�\�4ZYs�[���`�^�w����b�J'߆�E�ѻ�t�u$�J+�nC:�R.�1D7w�
��QHÒ�Q[�t���y�5٨1ȋ-�$V*�whR�v|'�"%�H����9/.�R&���)�T<J��0�"���rA���^����	  w ��zQ��FR��s9�^������l����^r�6ʑ�����E<ųB�B��p�uJǻ��\�2y��]~or�H
�d�j��t�J��Ut��w�h�p�������P�.�>&��{=��"�y=r��.V�S#����!�^�9�W�E{+�Đ;ƌ�4�x�,�b��X�5d��cxӄ��9,!�(�y��/����[P������,��_�l�t���8�SO�<�0�u��Wjl*+[��,�W��<)�ʧ?NX�F.�4���r~�~R�����E�$+���6cW���J㐷��{�}Y��.���)쇎�Z�7S�K�>��զ�L��c�镩�@�If�Y��h쑷���*�-���ӽ�ܟ>RK��+�B��N˕�wz��U-��K��I�r���8��,�l!n����b+Ŷt��03��[�v]��٧C�}�i]�~r�hw��eZ���Q��/D����ɈWF�|Cj!8�WZ��p����1v�-��+&W1�����s����)��sV��R����T�x�D�T�
���tyQeȍ��(H�8�m��7� =pY�,k��ɷ��šj���r��j���*�
LmM?��{R��&��wi	\	���u&ɯ)�_�g���_���:�'���3jѢ�1e�nyj�-�^��!r|2���"�u8�u�@�^u$�8���m!;�B� SѼ���E�Yp$ �&���v�$ڵ#��p׷�`\q�"�W~�T��mK���ܤ�_��l\`3|v�v�f|��/��1KTA:��On�+�:��x����4�5X�m��j"�S�ɉ?�냡���On�^:Y����k��ֱ5W�`�ǫ5���eL��[�v\��'9߀S�~�af����&h��Ӯ�7�f�O�d^v���ˠ�o����q�ʉ[��"�����W�V1� W[T�>�D2�;��)-p_6��Lou@�,� �Rq�q�yZu�p�E�9��de�t̏-�y�B�)1!`|��.��eKp ����I���gԢ�n	tk�Ln�%���\���,���@G���r�?%�:�N��I��W��u!>�4�����?�Q�ǧT��s�]������sH�H������P�6�m~	�c}<�B�j��%�^9�ɋ�yHk������	�,���ӌ�����0@��i��р&�/�B[��H��Q>����J+���i=�������a�6-X��b�-J�_���x㢵0R�=_�r;�4�^~�d�y��(429�;����z�q���W�V h�E����/�7�~���m�]�k5��va�k㏺�����a�5&����aB}����/&���X�fI�)j+�+���>P�uq�Q��7O۠/;���E	��u�Px��zL�N�5������:��,�HB� k~y�c{�f���,�fG�+�B��)|�J���g�Dg�����A�z�5 �U0����SV#�7d��L�nX�%�g��ґ�����$�R��-��!�[���g.��Zepۺ���R��#��u��(�
�5P���w����?<���Ȋ�e`p��E�����\��A���(al�4��m�v�K�n�,�	��c�4WeHhվ�`C�}یQ����CY,͐
m\gb��5 !Uꡇ?��#��� O����v�0�I��Y��+�u��71|.І��d�D�>i"T���BW��,�(�?Ȳ���3jP�X�y�dGn
X��e�U�9����jҴ+*2�Z���p^to;
���y�A�!���؛���I���]�[��8������L�EM//���a9a�sV��F���H߿����p?"��_,��p"�*�������I�� K/�2���d��~��t0�y��.� ��3?)�{i�qe��M��ص�(�t�܊#u�n�4� Ҷ#�H��Ay��}c�#flX�*��ߞ�S��GF�0�sJ�a��jH�"�{D۱?⪕ �U�u�E���G6�cSA��33
#�8���g�'�AD�b�r(��[D��6���b��9D�}�0�Y ���Ԓi���|���f��Z��Np��&	���^~]g�'4�"!�٘F�Ӧ���m�� f5h]T;��O�e$�2��7�|��~?AX�BB}zU�6;}0M3��	�����qP� ��V���n������'��Q�aUo�h<Ti�f��O��7}�>N9�ul�-?y��_��:Ù�5��@��q���?�$p����%��x��L#�=���n/����w=��Z�*�N�3����i"�����=���1K['WM u��<mk���#�7�ʏ���|���*&ofI�?�f�j1�ƎT-Z�:[Z�c9�j�#�]��n��r�.�BXnB@.y�2(������ D��$������XT`��%���f��	��R���D$��a���8����t$(�   �Ɓ����!�f�,$5-a��t$0���t$8�< \��ʣ���'�,���k"�ԾP��C)S�Dl�p)Ai$O��h���3�Slaeޔs�}��R�� |'E�B�'�Z�	<Gi�<g��P�0���k\��+���4}&4mUW���J�� %��l��N`՝�7�I���k	�����'��=�6՛h��ie�2��*�/Ry@�}�� ��ß9����)�NxJk�d鉊0a�2��x���Z����ǋP?ao�� V�N�<A�=�\��,?�t#=(j�Nڔs� ��ᡎ3�J	3^�]0i�<����(����O��4�ڃ�1��	�]��)�bo@�-�)-�q��/�J��6#?�m���;ZU䴥�����O��I���!��{������Axr�G �T�ZC
�W3|����t�/o�ρ���:f��ù*�A�D����:�tWԿG�zs��
�dI����k��9_z�
�\b����}�t�\v����Ӧ� ��k��WfǺ��e\�6���IL6�rH��P�B��ɞ���%fqP(~�Z�l8Ԛ蓚�=xI��CeZz)��X�����juKD��cSR��RĢ����d�B���}9�8q�:�d���:wpgy[��OJ��韢���o��7n@����B�6�����}!���6~�,r��ǀ��6��Fu�'�(��"�Ն���lVl6�_ �O�=��nn�ҏx�#Kޖ�P��R�57|�|_��e\�\��쐉�H�/�pⴂo��Bֶ�+Ș����vN������]�#M�<��`_�-:*��*�6��G�e�}#plܴ���e�l�G�o�IQ/��R
�y�E�#KR	�K�f�buP��}�#B�@V���퍫FE)��L}3+�?n{A��X���k<!Tt�O8��^�v��炉�"�X��v#�L���8G?l\�R瓟��	�aD�]Lw[��u92YI�	�v��ov��i�HYC�x�j䐠Q�F���@�!����A���S�h9\���+z[�>��.�s�����y���qP���2jG>�(�݉�����*;t1W�8h˵�o�X�\�:9=����NߓR����QZ�K$��$K�@x%SLI
��x�����7Ш�/������׆t/	Ȟɤ$���
s���I�{��EZl�l3�9FYCT+ѠD�g&���Ws:1��ge�!�[��9W�D�������tTE/@����ȆM�9�6�qz1ܛ:�_ }��3�'\*�ab�9����+�~����d�>��{S	Mk�|-!�JcB�@bR�UNme	��ƚ���[_�<�	���3��/��cm�W��$���Q���|�����ωL���<�j���ű[���!�=3�C�����=��t3�kP�`7o�PmugNt��W�l���!�~L5��
�d�y ���	�N5<�9�c��t#�i��Μp1�B��I�j�]���R��j��BIX�\g݂&�����V���b9��?�O ^Z[���4?���͐v�[���rK.�x�P�
7��q��	i�.�"�ʭZ�S�Ң<��D#?l'��@�>��d\����~nZa7=��]�ùJ0�\{���C4`U@|����6Ҧ�F|�D���9<ծ1�;�ةd��S72Q�LR����I�cX�^٩���rx-�	����1R	���MDߌ���q��C���e|�О[��5�C���H�*����<�g�4�V`�<R��(� Q��M�=��΍��ӸYV:�;���n�;���ӽIa�?f=~o�¨��k�I���%[iW��!oݣ�?�з�ԣ⡡Ҽ͜�n������ǭ��ń��$#2ך���if|r	� ��v���j�(%^���rIT�!���� S&�ⶸ���%�V݉��J�E��] s�m� w� �g��ttJ��}xi<�!�k� ��㑗U�r|�jQ��'��W�;�F[<�֥M�Q>����)�y�����_�2�l��뜧^�D�J��}�b��n22��q0�f;�H�݋N��ˬ�h����(&���y���k�%� �p#C�U�#L�B�ϲ���ݫki$(';�<�c� b!�m�'����U��������G�f�I�2�7j ���	�?w	(�;��6@�i���X<�y�>e1�E��VV�e����~W���F� ��s�/��w���D� ��3X�z|�;TԎMg"�R~˛�L'�Ay��Ph�_]ֿ���۝̩A��Zh �`hJ2�785�ea��1�-�{Xk�V��aƪ��Q_�h��&!1H����^�{�T?Y��눦�hT������3��3@���QPRs#$]��M�Ro���������ғ�z����Cu:?ϦuT9�O�S9��i/���M�x���bocڲ��1Z����ۻ����=�{��/~Sڵ/U�)���8�'gȑ��ܧ�,���5�1�o&���X�lGFf$���܊��t��.Y�5��:��x��1��@ۚ�&�t�\�|�x�.��Bᰐ���T�r���b]�5����j� [�f71%Ԥ	<k��N|
@�������]3�Y+�C:r�c�+���C�b�n��XGV����Z���@�P�u�\�צ!��.�,����9@��>u�=��
<���`�9�y0|@�0�d9:"A��h�2����Q��&.�ͩNg�?#v0�J�]Y�a��#�'�_�@|# )�6580ѻ��.լUgh�-{��yNfp�+�(X\��C�)e�Ļ`�JV�����u�+�էԇ]�j��]=}�<����j�"kbe�4��3<^�N��X9����x�q��#Lj�3*�����' ݇�N��x���=�V�+e��/���y9<EV��|�5�?E���m��Wn�G�1�W4-9���Z#v���6�{+����]����x�c�	<p����������}���~ʹ�٘��[d�H������'�y@9������&�a�LZYh,qKџu���L��nĐ|�N�8���x�5T~���n���S��1��Ϊ�9����r��~�PJ�Ѵ�w�Hkj�xqp��Y��%-$ ���r|��Q����<�s������S��(���
��MJu]�ba�� [���шI�3!���x�u9�nd�rP�1�Տ��������b1B�+"��m6����u'\���@���p�63l!p'e���{.=���/�KMb��p�&"��)}�T�$ϗ,�+���[���J)��z%��)P#�ă�Nd�
a^W�%�e:	�
�����s�W��!ղ��g��y�k"�yh����+SA(5�{���I�SZ^�6�g���kNM�J��@����w>>Ϲ^�ݮ����G����UT5)�l�^BI�-+K/ixq�$���\�n-{�����
+�>H���]Q�j9m1̔�N+�X�x���um+y�u��]�!W}xdZ����M|'�$�$�^L�������7�U��r[�� �_G�����3�0�JP��bNk�m#&kl{�HoG��{��{��~%���)8���	��,�Q�]��:ܓ����R5��*���5N�qx`��?B4�੠�	
��d%Ty�w�	��|�z�A���j�]�{�������(�"�V1���3)�]N�J+�uR�1�-Kn ���=��Xt�9oE�q
��GLےIQ��6�k���T\���ڦ$)[G�O�="��l" �J�19Υ�^1!D8�o��4B�I���D$}�<���1Z�U�޻ǭ"	��m��2��fM᧌+�8�au�O�"qѲ�4�"s���.d��Q7�wP�\����1�8B��)�_�g�R�e�CBj�JZ�����v�K:=uJ�hY��J�ʫT)��{�1���OM��9�=*֗aD�L�L�4)���5�{�����~�I���ĸ���4�#N��R�;�%����H*�G�z��9`!Eb: � �-W4`T��v%)<H��R��wl�+�m�
�,�
����f�в��h2�.J���P�Krj�[�$�������pE� ͞����e�UϚ�z]+yffG>�/�M���~��!�v�E�_vS�뻤ۜc�Ho Iqi�q$Y��:����<8���uX0����-�L-cg/;��cDk]��n��i��18�&�F�-����9�t&e���Ƣ��k�M���\�b-z�i+WB�f�T�)>Tdʎ�_zy
��k��"��ځ8���vPV�w�b����S`l���)��	�,��<a��pH������y
���1(�"���+L��׬�K_����a�M*�'4����E9��0�0A�����OGF����'JMtf�u=J*%��[MW�9������#��B}$��)�%��_�YO�3��?����[�s�Y|�Sy � ���K���"���b��<�L�����#_��������p�4�6A�]��`�,C˄����弮d*#�aޠ��d������}i�SP�T����%�ӌt�����t8f����i�1� ��I�Y�`�M����'h���I����!����[��1���� j)�'��>g}P1K�裂��܌���(�!�4�޸�U��M�浑Z���>|��ntj�KC|K�o�v��.�R;��
�f��6N�Vj�_��X� ����])0�N5,�JQ W-�6	��+�,�^S�+ֵmޟii� ��D���(#D�p�Jt+\��h�,� �e/%%v�(q�\cΣ��y��[̹|(WLQԕgF����-��-/�	�?f�<�Y�թ�^���\x�Z�1Y=Xd-���ŭ���7�C�P<��-7|~�W��I&�Ļ�I����|g�$����ʫG�^6���,o�p�"��<:ݥs�n�w D��G�+����j"јu"Ŋ�S�����K��q���~�����y��8�"��o7�H~���yG���(�!_66�\�b����A��ݿ{Ė~7�:Q�WZQ�k���kNU}�M�#��?c��D0)_�G��l9�c�7WVip���V�����5��@�������~��L�F}� �bL:@P��JQd��#�`��:BG�Ց��'br��D���c��7�AU`x>�l�/�e�q�1N"rjs
�ϕ`�:i�,����i.*i+�+27'��Jy��_o�(j|�@憎��b8�܊���2(T��@�`�'eg����9�������ɨoΥ<{({A�'w�K�&�U���7��5ǖ�81��֥N���)@0���^2��9�'�'?sz�N1�t�w4����X܆@k[
�������uOEpP{���������a*q	��˜���=�^�9e�\��(���%�4�/�{l%R5n�a�[�Mr�"��<�h"倆���{���a*D��QW�����E�H����RbJ�� ^�hY�ъ��L���%�A�2!��E���-~C>Z#N8��/��,6֯x�}�l�ӲL�b�VQI����_��
q�jTխ�ϝ�t�#���,M�5��VM��xw�}T����0#=j#��ok1�T�l#�~=�'����>#�2�{6���`����	����d3`�1'�XU���_��f%���m��L5�C�~;�v}wE�f];eo�$�N'"T��d��p���0�2
����� e�qbz	D��9C�n&gQ��;�X�l�I�륊�r��1kB��xU6��K�E��E����D�&�%V@�M��]Wp���v��K��[�JmX�9��UZ(�ѝbQ7����R��h�>~%���VbPb^©g�� �ʸ�7�Ȍ���� X��H�����QQ���ϓzP�ᲁ���:�41l�.��y�bz�wl#,Nm��	�*��X�^=��p��j0�\Z FDz��\[�`?*kL�ө8nLqQv�QWvmDúj�T��0r�۶�/B�;5��%���X�C妗�}0��N�[���_y�e���Y���s~�P�01u�����Z �@L'g�vܥRSR�7���E�vg��#�p[�Ԩ8$y��_z�bwO�j��w����) �& n�n�q��ZmKr�k�n8,�� Ϯ�fs��x��#!oěj�"Ѩ8���{J�I��-�,W��DF���NM{UL3R��f�r��|z�&\Z`V���v���|��_bb�2V��i�B9XW�����(�.�8W�7�u���Z])��_�E�n��Kƀ�3|�q�6ݦY�o�`s�G�Ų�WBr��y�&DUO����y�[讀�Z/l�Bx
�c�U�z�7����N*�3��th��ט�f��j(s
W�.�� 8i���s�"?j�g�۴#I ��	k��26���n� �� �+Y�Hc҃�bdXE��O�1��G�1�`q[ �H�n�m	+��,F��=�ܪ���=�#�%�G��e�޻���{ʷ	���U쳩�3���S���X���3d��*%���r����� b�9�r\ݵ!)��A�>���}ܤ�J1�0�$bx���f$R�K����|I[�0�"�H��tY8~'��6~295uz϶�d;��ȗVd�l6�iT���m��D{R��9��0��)\��1�5��ꑹ�/f�k���P��~S��|�"�u��gꁷZ�\?=���.�؝�<�[P��lIT�>�4!Dɰ��C�-	KL�����2 �MQ�!XR��ٷt�d���:&���P�\�6��0V1nlr��i��8����6e�S���^=4z� ��Z�B8{JY�.~N��<�\<�d	���;ry�˄Y�V�T�c@�C����^}č[��ʚxGZQ;"���M�~^�YFk�пZ��e"���"{!���պ����vZ��zY��U�	?�8���`�gF�@F�����]����{v5�\r �
�����̇`��D$����j.�S���Ҍ�5;y�`�$Ł��jzf�����x�6shR~l����L�� o¬=r�~{!��!�t��eÊ�@7u\˻T�9W^�n�et�4���$�2�V���?B}nL҉�05h�U�tll�l+rM�+��ø'��#�\[���;�{kR���ay=`��x���+��� yX�|���ޜr�?�fE�ov+�j�Y��%]D�R	y�=3���K����������c^�2�ڢ��Fј'�E4����>����C�P�|(�~�I���!uJ�y��;�����˨�b;،X/mx��k�{���6��VsA�k�,�� �x8�1�xxB�Ƌ�e��n�jF�p��A��!�4e��H�"[��↙��J����f�62��OaDK�&a��Ab3�/O���Ag��޶��נ��gQ��Ӣ+���X��U���羵$��xV2�N��h��\~�s:�iO�c�6��c�d��٢�o��za`=�sXYPڻ r�D�9}{�:����h���g���5X��"g�!Ú�G_#
2A����5�� e��K��6A�ѕ��ܟ�
�oFQ��Y��S��� ��K����0O)1����3�*t^}�i�Zp_��60�Ei�	at�%�5�v����Kp#!~C$ r�Zj��Ә`U�=6�����;M�(��V���.YR����3�$^�����z}���6�V/�̠ af�@,}��/
J�(��s�z���m�ÒX�@�o����a�XG�Vwj/�pڛj�����A�39��sq?�;��:bN/v�:���Kʁ/%d[��p6�&�'&@�̏��;���}M�:Ye.����j�����]�e"���	�}����%�V!qN�Y$g#�^���|�8�T�aV� I�yI��޲p���X=((����,z���:Y��(���`�[s�횹�ĭ:
��6= ��i��KS4��'��}�� �eq:Yy͍f��S>[��O>�cM����VF��,0�����^�AUwha��t�����-[��#z�����-X�,!i��T����M!����B�A�Cc��շ����F��F�υ�����
���O��S�叿D��@@W? �9��q��N}�ֳ�VT1��y�6�_����[�Tp��\���k��7���t$N�p����k����Zqi�t����|��[~$�=��N�>�/���ٯ}�G�+iϪt+���i�)�!Q%�{u K���Cb�H��$�.�]��D�:Zf�}}�	���_�<��.
$�`L����	��tΔ	Q�0I�(�����6_��*�z>#��3[�9NWn}�5��8g�"��Q6�d�O��
����$^�촪�Vtj�NqYZd�`Y�h��9n�h[?X�ڙ�������u,5�R� ��:�a�������Q�����%_+��^���t����A�.���u`~�������������~�)~u�N�И�?w���-�E갠6�K:����E���O�v���p'X���ٔJF�ۀ��C��m��`kƍ��
��H�	�!��d�Vխ�܃\��0_�H7!�r�ڔZ��z���0:���2�m
<�1���c�Y_UZ��>o+�����̈�o#��.T��/K4���<�*1��zmPoq�h��&o���LE��I2Y�xG.��6�h��rvpAxW.�T�j��_.g�/��T��F�j��|Pb5� ���@T�N��1*1G=>��\�0-��d�v��n����|di�S#�����5���1g	7}u�\#�hu5(��m��d��/	6V"+tܞ^�Zq�r<��N�YT�)~D��H�B��)�=);���o6f�J�Y��'��4)�}p�E��h��\�%v��l�����{�Tf�>���ۤ��}#���4��׋�{eP{4j����9�nu�`�v]��B^\HD�x�Dn=���JB��t�71�N]�p���]���Q ��u���:r7�B<��BD3x�1>�y>P�Lp�]��hվ �*%DT%$�{azY�Mu[��b1�x��~�o�@�� �+�b�r������eg�E���t���ޭUv�𹾲"��/L!��M�X��P��p<x?=$�\vqO�5:^!��T��W��G7�l2� �����3�T�!X�<����#�0�?�;�ֽm�x&����&/�}���0����y���̥�#�ʖ��&m6e�D�����A��:�\�}���6E�<�-�.�����,&2{��
;
�ec����4�b�N�){����:��Kol0��"�q9��݋E�)�0�� �vp�d�X�u���0��E��I�����Q0�' #$'>�뢆4�{�u\�E�h/IU�(���,���,��`�5��3�s��3��s[�A������6Q|�.Y ���{+@�����9�g�h'���9�u�I�;I��+1Ld�y8�N崴���h�R:�gA����h�l���FD��S8Ǹ�����g?������'���E�9%w||��������	��૵�y�g�;���lc4%A<�y����W��O��lX�Ő&K /��UcI�e;��̓�9��6���At��R:�O�����ڙ4Ӣq�G�lG+p�T�Ƽ�� v�l@G��V~�u�$M���v���q*�2����6���e�Z���- ��nOv��"� �]�6e�� z�)�А�['������p�ҕ�ߟ�u�fi�̔,G�ra��O�LP$Ax� �羊�Ef�7�s|3�8����1��>9�w��r�Wr�`Nt�8Nlh�Trx��#jqp������waz���0&��u�ϣx$m�Z��=�շg~�|����ѻ����y�˲Q ���(���^ ��&cz�&G���-�^��~|���ȱ�ᮔu/�{�s��ۂ��I��Q�$���!8Cʗ�שR��j�^�
'�{���I,�v������*�n�
��6�I+#%V��d��$f�����:P5h&���S���                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                  