MZ�       ��  �       @                                   �   � �	�!�L�!This program cannot be run in DOS mode.
$       ���si��si��si�ld��si�Rich�si�                        PE  L �G        �   p  @     �     �   @                     `    �D                               � <    � @                                                                                                                  �     �                @  �.rsrc   @  �     �             @  �.idata      �     �             @  �vv2      �  �  �  � .DLL        @  �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                ��rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rß��3��s��2ß��3��s��2ß�3��sf�2ß�3��s��2ß�63��s��2ßʚ3��s�2ß�F2��sB�2ß�
3��s��2ßʲ3��sZ�2ß�b3��s~�2ß�3��s��2ß��3��sV�2ß�f2��s�2ßʪ3��s��2ß�3��sR�2ß�f3��s:�2ß�R2��s��2ß��3��sn�2ß�"3��s��2ßʂ3��s��2ß�z2��sr�2ßʖ3��s��2ß��3��s�2ß�3��sJ�2ß�&3��s��2ß�r2��s��2ß�~2��s��2ß�j2��s��2ß�*3��s�2ß�:3��sb�2ß��3��s>�2ß��3��s��2ßʊ3��s��2ß�.3��s��2���}ß�mÞ�r���r���rÞ�r��Q	@�}|"�.m\��rÞ�mÞ�rÞ�r��^�M��rÞ�rÞ�r���l�� -Þ�rß�rß�rÞ�r�V#-æi/���r�>�2���Þ�r�t���2���2ò�2��2�d�2ø�2�
�2þ�2��2�~�-���-Ê,�XOr�W�-��s�X�T�W�-��s�X���W�-��s�4)8"���}�(("#!Þ�r���rÞ�rÞ�rÞ�d���r���rò�2�
�2���=Þ�r���r���r���mÉ�r���2Ú�2â�2��r��r��r��rÞ�rÞ�rÞ�rÞ�r��]�m��^�M��r�.�r�6���ư�~L��6?���rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�r���rÞ�rÊW-�*�r�.�r�f�SRC�axCa�oV>J��rÞ�rÞ�rÞ�r���rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�r�5�rÞ�r�rT-�z�r���j�� -Þ�rß�rß�rÞ�rö"-�nn/���r���2���Þ�r���<��2��2��2�>k-��2�:�2���2��4-��X-��2�7-��7-��2ò7-�~�2�r�2�f�2��2��:-Þ�-��,���-æ�-��-þ�-�~�-�X�[�W�-��s�X���W�-��s�X��W�-��s�X���W�-��s�XZ�W�-��s�X���W�-��s�XO��W�-��s���i�� -Þ�rò�-ß�rÞ�r�&"-�*m.���r���2���Þ�r�\���2���rÎ-Þ�r�*�2���r�2�2Þ�r�.�2���r�2�2���r���b��2�V{.Þ�r�^0�<��2�6v-��-��:-Þ�rÞ�r�V�-�~�-�ڥ-Þ�-��-��-���l�"�r�Z3-ß�rÞ�rÞ�r�j�2�Z?�<�3-ß�r�S�2ç�2Ï�2û�2Þ�r�2�2�J�2�f�2�l�2�r�2Þ�rÞ�r�V�rÞ
0^Q����ʥ�,m�V�rÞ
0^Q�#!�ʥ�,m�V�rÞ
0^Q1���ʥ�,m�V�rÞ
0^Qm���ʥ�,m��r���rÞ�rÞ�rî�rö�rÞ�rÖ�r�&�rÞ�r���r�-�r� �rÞ�r�t��%P�2xSmC����s��%P�2xSmC����p��%P�2xSmC����G)a��
F�Ȗ��vo�
Pucb�w��L��rÖ�mÞ*�ʯ�r�AIIF�{o�Z�T�%�T� �$SqDr�BV�����r�>��#��rÞ�kÞ�rÞ�rÞ�mÞ�m���rÞ�r���r���r���r���r���rÒ�r�������5��:����������������=������5��������������;��;� �;�����-8�z,8.t�=.k�#�h	�P !Z ��Z�\��Z�\�����r�� -Þ�r�n/�~/ú�mÞl/�`�2Þ�r�����!�������������+������3���������:���?���������� �����rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�r�
�2á�r���h�� -Þ�rß�rß�rÞ�r�"-��l/�c�rþ�2Þ�rÞ�rÞ�rþ�2�V�rÞ
0^QmÞ���߬b�V�rÞ
0^QmÞ���߬b�V�rÞ
0^QmÞ���߬b�VmÞ
0^QmÞ���߬b���rß�r��rß�rß�r��r���r���rß�r���rý�l¾�r��'�<��<��rß�rß�rß�rß�rß�rß�rß�r�V�rß�rß�rß�rß�r��r�&�r��r�>�3��r��r���s���rÞ�r�n�r��rÞ�rÞ�rî�rß�rÞ�rÞ�rê�l�n���'�<��<d�D<��r���pþ�r��r���s�=��Þ�r�>��>����rÞ�r���p��r� �r#��s���rÞ�rÖ�rþ�r���rÞ�r���pæ�r�:�r���s���rÞ�r���pþ�r�6�r���s���rÞ�r���p�.�r�&�r���s���rÞ�r���p��r���r���s���rÞ�r���p��r���r���s���rÞ�r�������rÞ�rÞ�rÞ�rÞ�rÞ�pß�r���r�>�r���r���d�� -Þ�rß�rß�rÞ�r��"-Êi/���r���2���2Þ�r�B���2�[-�Z�2��3-�Z2-�.�2��b-�b[-ò�2þ�2�}-�~[-î[-���2Þ}-Ú[-��[-��a-�&Z-���2�^`-�Z-�zZ-Ö�2�"|-òZ-�>c-ÎZ-���2��Z-��`-�"U-�U-���2�`-�VU-�f|-úU-�V}-ÖU-��U-��|-�:T-���2ê|-Îc-�T-��2-�2-æy-ên/��'-��2Ê�2�rb-���2�&b-�:�2�6&-Þ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�r�V-,���-ö�-�R�-��,�f�-Ö�-ê�-�z�-�6�-Ö�-Ö�-�XW3�W�-��s�XϦ�W�-��s�X���W�-��s�X[��W�-��s�X��W�-��s�Xg��W�-��s�X���W�-��s�X�F�W�-��s�Xs��W�-��s�X7��W�-��s�X�I�W�-��s�X��W�-��s���m�� -Þ�rß�rß�rÞ�r�f#-�^n/���r�Z�2�l�r�r�
I�<b�2�`.��g-��g-�~x-��2��2�Rx-���2�
g-��'-��2�d�2Þj-�Zx-� -�j -�N-Ö-�6&-�j�2��{-�6z-�v -�z-�Bz-âz-þz-Úz-�� -Ö -��z-�p�2�:�2�(�2��z-�v�2�*u-�2u-�u-�bu-�|�2�Bu-Úg-�B�2�Ju-��2��$-�Ru-�H�2Â$-þu-Òu-�.�2��u-Ê'-�&t-� �2�t-Ê -�nt-�Bj-���2�&-�vt-���2�"�2�^t-ît-���2öt-þt-Êt-Òt-Út-��t-��t-�N�2�T�2�Z�2��t-�&w-��t-�w-�>w-�fw-�4�2ö$-�Fw-�r-à�2æ�2æ -��{-�>-��~-��h-�&-�:-�b-���2�g-þ�2Ö�2�v-�J�2��o/�rv-�d-�b-�&n/�~d-�jd-�Nv-�Zv-òv-þv-�
f-�b�2�
�2��l/��2Þg-��'-�f-Òi/�v'-��<-�-ò -Îd-��v-�g-ì�2Ö'-��2��v-��o/�x-�^j-���2���2��v-��,�^�-�.�-î�-�ʴ-ö�-�X�y}�W�-��s�X�a�W�-��s�X?�W�-��s�X�U�W�-��s�X�Z�W�-��s�X��W�-��s���k�� -Þ�r�2�-ß�rÞ�r�F"-�>m.���rÊ�2���Þ�r���<r�2���r��@-Þ�r��2���r��2Þ�r��2���r��2���r���b�B�2Î{.Þ�r�^0�<2-�~C-�
C-��@-��]-�B-�\-�2_-��\-�^\-ÒB-ÊC-�NB-��C-��X-�j]-���2��:-���2���2�"�2���2Þ�rß�rß�rÞ�rÀo�3��r���s���sÞ�m���r��rß�rß�rÞ�r�@o�3��r���s��r�V�-�"�-Ö�-�Ҥ-�ª-�«-�z�-���-�B�-Â�-�B�-�j!,ö�-�f�-�&[,�
�-��-��@-���l��r�Z3-ß�rÞ�rÞ�rÂ�2�Z?�<�3-ß�r���2���2���2�'�2�;�2��2�c�2�w�2�K�2�_�2ó�2Ç�2Û�2���2���2���2Þ�r��2���2�f�2�l�2�r�2Þ�r���2�V�rÞ
0^Q�(!�ʥ�,m�V�rÞ
0^Q)���ʥ�,m�V�rÞ
0^Qu���ʥ�,m�V�rÞ
0^Q9���ʥ�,m�V�rÞ
0^Q	���ʥ�,m�V�rÞ
0^Q	���ʥ�,m�V�rÞ
0^Q����ʥ�,m�V�rÞ
0^Q���ʥ�,m�V�rÞ
0^Q����ʥ�,m�V�rÞ
0^QI���ʥ�,m�V�rÞ
0^Q����ʥ�,m�V�rÞ
0^Q�u!�ʥ�,m�V�rÞ
0^QU���ʥ�,m�V�rÞ
0^Q����ʥ�,m�V�rÞ
0^Q%�!�ʥ�,m�VmÞ
0^Q����ʥ�,m���e�� -Þ�r��-ß�rÞ�r��"-öi/���r���2���Þ�r�j��<Z�2���r�Ff-Þ�r���2���r���2Þ�r���2���r���2������Æ�2�Fb.Þ�r�"��~M-�
g-��o/Ê�2�6M-���2�RM-��o/�^M-�vM-�6[-�vf-�nj-�g-�`.��g-��g-Þ1-þi/�"�2ê�-�z�-��-�Vf-æf-������r��>-ß�rÞ�rÞ�rÒ�2�F<�<�>-ß�r������röf-���oÞ�rÞ�r�f�2�z?�<�f-���o���m���r��?-���oÞ�rÞ�rÞ�2�<�<�f-���o������röf-���oÞ�rÞ�r���2�z?�<�f-���o����"�rÞf-���oÞ�rÞ�r�r�2�J?�<�f-���o×�2���2���2Þ�r���2�"�2�f�2�l�2�r�2Þ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�r���2Þ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�r�&�2�"�2�f�2�l�2�r�2Þ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�r��2�"�2�f�2�l�2�r�2���2Þ�r�v�2�"�2�f�2�l�2�r�2Þ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�r�^�2�"�2�f�2�l�2�r�2Î�2Þ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�r�V+mÞ
0^Q�!!�ʥ�,m�V�rÞ
0^Q�%!�ʥ�,m�V�rÞ
0^Q����ʥ�,m���o�� -Þ�rß�rß�rÞ�rÆ#-�Jn/���r�*�2���r=��r�bD�<�2ên/�b�2���2��2ò�2�i/���2�.�2��l/��2Þg-��'-Ê�2��'-Òo/Ê:-�Ji/��o/Òj-þt-Ö�2�"f-öt-�`.��g-��g-�
�2��'-�*&-��'-�i/��'-�v}-�Bj-�B�2�2!-�^j-�Jj-���2Þv-�Bi/�Fi/�
g-��v-�&-�Bq-�*u-��q-�Zi/�6g-�:�2�2p-�p-�np-â&-�f-��8-�F-�;-â-�Rp-ú&-�6&-�~&-Î-�j -�bi/� �2�>�2ît-���2Êt-�Zp-��-ò-âp-þ'-êp-��
-Òg-�F-Ê-òp-ò
-úp-�x-Âp-Êp-Òp-�-��a-�6i-�J-��-��-Þ1-��<-Ö-��&-Ä�2��-ò'-�-Ê�2�^-Æ&-��-�f5-��o/��o/Úp-�v�2�&!-�>!-��-�j-þ -��i-��2��z-��p-�g-Æ-�>6-�4�2�v-�B'-�v'-æn/Æo/���2��p-��-�s-�&s-�6�2�ns-�r-�d�2ø�2Òu-�'-ì�2Ð�2ò-Ö�2þ�2�~s-�-��-�:'-�N-�Js-�p�2Âs-Ü�2Òs-�
!-�z!-��s-��s-�"r-�R!-�^!-�2u-ê!-ö!-�!-�b!-�n!-�F!-�
r-Ò-Â!-�&n/�B -�b-�B6-�~i/�vr-��-���2��-Ö'-��o/�ni/��2�ji/�*-�^r-òr-Ær-�T�2Ör-�H�2��r-��o/��r-Ú!-��&-��!-��!-�. -�" -�o/��!-��!-Þ&-Î$-�.'-��$-��$-�"'-�R$-��&-��r-��o/��o/þi/�"�2�vf-�nj-�6M-���2�>M-�vM-�~M-�RM-�^M-��'-æM-öM-ÊM-��~-ÒM-ú -Úg-�"n/��M-��o/��M-�-Ò&-�^i/Òt-Út-���2Òi/æ�2��i/Öi/Üi/Ê�2�r&-�&-�f&-�N -ò-�j-�^-�2L-��-�L-�bL-�~L-�^L-þ-���2�Rx-�"�2þL-ÒL-��L-�|�2Ê -�Bu-�vt-�Z -�bu-��L-�
O-�&t-�jd-�O-�rv-�
?-�nO-�~O-�JO-Â5-æO-ÊO-��O-��O-�x-��t-�"N-�.N-��t-Îd-��v-�g-�u-��{-�>-��h-�&-�:-�
N-��O-�b-�N�2�nN-þu-�
/�t,�X�}�W�-��s�Xo��W�-��s���r��\-���rÒ\-���r�F\-���r�.\-���r��]-���r�V]-���r�]-���r��B-���rúB-���r�vB-���r�.B-���r��C-���ròC-���r�fC-���r�2C-���r��w-���r�Ny-���r�y-���r��~-���rþ~-���r�v~-���r�.~-���r��-���r�V-���r�-���rÖ|-���r�R|-���r�|-���r��}-���rÆ}-���r�~}-���r�>}-���r��b-���rîb-���r�b-���r��c-���röc-���r�nc-���r�&c-���rÚ`-���r�F`-���r�6`-���r��a-���r�ff-���r�h-���r��i-���rÖi-���r�Ni-���r�>i-���r��n-���r�Fn-���r�:n-���r��o-���rúo-���r�ro-���r�*o-���rÚl-���r�Nl-���r�l-���r��m-���rîm-���r�jm-���r�"m-���rÖ-���r�v-���r�*-���r��-���r�-���r��-���rö-���r�n-���r�"-���rÚ-���r�F-���r�-���rÆ-���r�-���r��-���rþ-���r�v-���r�*-���rÚ-���r�N-���r�-���r��-���rî-���r�-���r��-���rÆ-���r�v-���r�*-���rÞ-���r�Z-���r�
-���r��-���rî-���r�-���r��-���rî-���r�n-���r�&-���rÞ-���r�Z-���r�-���r��-���ræ-���r�-���r��-���rÊ-���r�F-���r�-���r��-���rî-���r�j-���r��-���rú-���r�F-���r�:-���r�� -���râ -���r�: -���r��-���r�Z-���r�-���r��-���rö-���r�n-���r�&-���rÒ-���r�J-���r�-���r��-���rê-���r�-���r��-���rþ-���r�r-���r�*-���r��
-���r�Z
-���r�

-���r��-���rò-���r�-���r��-���rÎ-���r�J-���r�*-���r��	-���r�R	-���r�	-���r��-���r�Z-���r�-���r��-���rÎ-���r�F-���r�>-���rÞ-���r�Z-���r�-���r��-���rÆ-���r�~-���r��2-���rÊ2-���r�B2-���r�>2-���r��3-���rö3-���r�3-���r��0-���rþ0-���r�~0-���r�>0-���r��1-���rê1-���r�b1-���r��6-���rÊ6-���r�j6-���r�&6-���rÞ7-���r�Z7-���r�7-���r��4-���rö4-���r�4-���r��5-���rê5-���r�5-���r��:-���rò:-���r�� -Þ�rò�-ß�rÞ�r�6#-Þl/���r��2���Þ�r���<��2���r�*?-Þ�rþ�2���rÆ�2Þ�rÂ�2���rÆ�2�������~�2�6z.Þ�r�� �<�<-�j -Æo/��h-Ò-�6�2�>�2ên/�v'-Ò-�nj-�Bj-�Ji/�
�2�^j-�Jj-���2Êo/���2���2Îd-�Fi/�Zi/�6g-�
g-���2���2�"�2�g-�g-�Bi/���2þ�2�(�2�vi/�^i/Òg-�Vi/Úg-Ú$-��$-��$-Þg-�.�2��l/��2�`.��g-��g-�"f-�4�2�
?-�*f-�v -�: -��-ò-þ'-�6f-�
f-�Ri/�f-�i/Ê�2�:�2�rf-�b�2��'-��o/��o/æn/�B'-��o/þi/�"�2�"n/��o/�F-Òi/Öi/�~i/�x-�bi/� �2��2�x-�i/�2�2�&n/�*-�bx-��2ò-��|-�rx-�Z -êd-�j�-�B�-�ҧ-���-�B�-�6a,�2�,�ґ-�^�-���-�ޜ-Ö�-�
�-�r�-�-�~�-�R�-��-�ޔ-��-��j,�.�-��-�F�-Ê),��-�R,Þ�-�:?-�
?-���b���r�?-���oÞ�rÞ�r���2�&<�<j?-���o���b���r�?-���oÞ�rÞ�r��2�&<�<�?-���o���m�"�r��?-���oÞ�rÞ�rî�2�6<�<�?-���o���m�&�r��?-���oÞ�rÞ�rÊ�2�<�<�?-���o����*�r�J>-���oÞ�rÞ�r���2�<�<Z>-���o���a�.�râ>-���oÞ�rÞ�r��2�f<�<�>-���o���b�2�r�?-���oÞ�rÞ�r�R�2�&<�<�>-���o���b�6�r�?-���oÞ�rÞ�r���2�&<�<�>-���o����:�rÎ>-���oÞ�rÞ�r��2�v<�<�>-���o���m�>�r��?-���oÞ�rÞ�rÂ�2�<�<�>-���o�����r��>-ß�rÞ�rÞ�rÞ�2�F<�<�>-ß�r�r�2�C�2�P�2á�2���2��2��2��2ç�2û�2Ï�2���2���2���2���2�3--�--�o--ë--÷�2Ë�2ß�2���2���2�/�2�k�2�S�2�--�C--�W--ÿ--Ó--Þ�rÆ�2��2�f�2�l�2�r�2Þ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�r�z--Þ�r�f--Þ�r�--Þ�rÞ�rÞ�r���2��2�f�2�l�2�r�2Þ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�r�*--�>--Æ�2Þ�r�^�2Þ�rÞ�rÞ�r���2��2�f�2�l�2�r�2��2Þ�r�>�2��2�f�2�l�2�r�2�&�2Þ�r�f�2��2�f�2�l�2�r�2Þ�r���2Þ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�r�N�2��2�f�2�l�2�r�2Þ�rÞ�rî�2Â�2Þ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rö�2��2�f�2�l�2�r�2Þ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÊ--ö--â--Þ�r�N--Þ�rÞ�rÞ�rÞ�2��2�f�2�l�2�r�2Þ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�r�J�2Þ�r�v�2Þ�r�b�2Þ�rÞ�rÞ�r���2��2�f�2�l�2�r�2Þ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�r�.�2��2�f�2�l�2�r�2���2Þ�r��2��2�f�2�l�2�r�2Þ�rÞ�rÞ�rÞ�rÞ�rÞ�rÖ�2Þ�rÞ�r���2Þ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�r�a+	?��r�YE��L�"�n��r�J�2ß����:Þ쵙�,m��n)��rÞW�-��s�V?mÞ
0^Q����ʥ�,m�V?mÞ
0^Q����ʥ�,m�VmÞ
0^Q9���ʥ�,m�VmÞ
0^Q���ʥ�,m�V#mÞ
0^Q����ʥ�,m�VmÞ
0^Qյ!�ʥ�,m�V'mÞ
0^Q��!�ʥ�,m�V�rÞ
0^Q9���ʥ�,m�V+mÞ
0^Q�!�ʥ�,m�V7mÞ
0^Qa5!�ʥ�,m�V7mÞ
0^Q-���ʥ�,m�V7mÞ
0^Qu1!�ʥ�,m�V/mÞ
0^Q����ʥ�,m�V�rÞ
0^Q�!�ʥ�,m�V/mÞ
0^Q	���ʥ�,m�V�rÞ
0^Q����ʥ�,m�V�rÞ
0^Q����ʥ�,m�V�rÞ
0^Q����ʥ�,m�V�rÞ
0^Q-���ʥ�,m�V/mÞ
0^Q����ʥ�,m�V/mÞ
0^Q�!�ʥ�,m�V�rÞ
0^Q�4!�ʥ�,m�V�rÞ
0^Q����ʥ�,m�V�rÞ
0^Q�3!�ʥ�,m�V;mÞ
0^QA|!�ʥ�,m�V;mÞ
0^Q����ʥ�,m�V;mÞ
0^Q�Q!�ʥ�,m�V;mÞ
0^Qm-!�ʥ�,m���n�� -Þ�rß�rß�rÞ�r��#-úo/��rö*-�F�r=��r� �<�--âN-�BN-ê$-öN-���2��N-ÂN-��N-�^$-�>-��-��-��-�v-�v4-�N-�*-ø�2Ü�2��2��2��N-�"I-�Bm-�:m-��$-��$-�:�2�l-Ê�2�j�2�vh-���2���2��:-��2�6&-�*u-�Ju-�B�2��2���2���2���2��<-Æm-æl-���2�*I-�.�2�Jo-��m-�H�2�nt-�>I-�N-�"f-�g-æ-�z1-��6-Â1-�.1-ê;-�'-��1-��-�>-�i/���2�'-�j'-ên/�(�2�vi/�N'-�`.��g-��g-�~x-�I-Ò-�6�2æn/��h-æ'-�Z'-�BI-�-Ê�2�^-�Bj-�vM-�6M-æI-òI-úI-���2�4�2��I-��I-�
g-��I-��I-�2H-�H-�rH-�RH-âH-òH-ÆH-ÖH-��H-��H-��H-�.K-�
K-�fK-�BK-�^K-òK-ÊK-ÚK-��K-��K-�2J-�
J-�J-�JJ-öJ-îJ-�Bu-�Rp-þJ-�rf-ÆJ-��<-ÎJ-ÞJ-ÖJ-��J-��J-��J-��J-��J-��v-��J-��J-��J-�&E-Òg-�Rx-òp-�.E-úp-�6E-�x-��r-Âp-�>E-Êp-Òp-�E-��a-�
f-�E-�bE-�vE-�JE-êE-ÆE-��E-��E-�:D-�bD-�BD-�VD-��-�b
-þ�2�v-Ê-��-â-�f-��-ê	-��-�f	-�-��	-��z-�p�2�Zv-�v�2þv-îD-�6g-Ê:-æ�2��-��<-��l/��2Þg-òG-�n;-� -�F-�bF-�vF-�BF-�RF-�^F-ÂF-ÎF-��F-��F-���2�2A-�>G-�G-Úg-�jG-�FG-��E-�~A-�nj-�� -�-�;-â-Þ-��r-ÂA-�rx-�^-ú -�:@-�^-�*-�*@-�Zi/��v-��v-�.-�-�J&-�vo/�V&-��-�Fo/�Vo/æo/�@-�@-�f@-�v@-�B@-�R@-�^@-ê@-ö@-Â@-Î@-Ú@-��@-âG-�rA-�nJ-�~J-�
I-�bN-�v}-�R
-��8-�>9-� �2Òu-Ö'-�T�2Â-Þ1-��<-�v-Æ-�*-���2��@-Æ-���2�"�2��&-î&-�B6-��-��_-�F-�b\-�d�2��_-�&^-��'-�6^-�
^-��&-�^-�ji/�F^-���2�b-�0-��0-�V0-�&-�V-��5-�N^-��^-��^-���2ò-�Js-�
Y-�jY-�Z�2ì�2�ns-�r-�N�2�2-Þ-Î4-�-�$�2�*�2�0�2�6�2�<�2��2Æ-��-�v-�j:-�zY-�&-��2Î!-�n-ò-��!-Âs-Òs-��-��l/Þ-�o/��l/��l/�n-��l/�*o/�.o/�2o/�>o/�o/�o/�o/�: -�:-�F-�" -��8-�F-Î-ò-��-�-�2L-�L-�B-�~L-�bL-��2�^L-�FY-Îd-�Fi/�g-�Bi/�
�2�^j-�Jj-���2�>-��~-��h-�bi/�&-�:-âY-öY-��Y-��Y-�b-�j -��z-�|�2�
O-�~i/�jd-�O-�rv-�
?-�^n-��n-��Y-�i-�.X-æi-�
X-�VX-êX-ÆX-Þ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�r�"�-��-�b�-�&�-��-��,��+,��-���-�>�-�*�-�"�-�&�-�.�-�6�-�Rb,���-Ò�-�j�-â�-�ޙ-�R�-�9,�6�,�>�-�:�-ò�-�r�-�^,���-Ú�-î�-�/,���-�"�-ò�-�-Ö�-Â�-���-�f�-�.�-�b�-��n,�V�-��-�v�-��B,�Bs,�Zy,�,��,��1,�"�-ò�-î,���-���-��-Â�-�֢-Ê�-���-�ք-þ�-�ڦ-�~�-�z,�6<,�F#,�RN,�D,�V�-�Γ-�J�-�f�-��-�R$,���-�~�-���-�f�-�:,���-ö�-ÎV,��4,ò2,�&�-�N�-��-��-�X+|�W�-��s�XN�W�-��s�XkC�W�-��s�X'y�W�-��s�XB�W�-��s�X���W�-��s�X�)�W�-��s�XM�W�-��s�X��W�-��s�X7�W�-��s�X#t�W�-��s�X+{�W�-��s�X'x�W�-��s�X?w�W�-��s�X7?�W�-��s�X[��W�-��s�X�n�W�-��s�X���W�-��s�Xc��W�-��s�X�e�W�-��s�X/~�W�-��s�X[m�W�-��s�Xo��W�-��s�X7X}�W�-��s�X1�W�-��s�X3�W�-��s�X�l�W�-��s�X{j�W�-��s�X���W�-��s�X�8�W�-��s�X�D�W�-��s�X�G�W�-��s�X-�W�-��s�X��W�-��s�X+k�W�-��s�X�X�W�-��s�X�{�W�-��s�X��W�-��s�X���W�-��s�Xϣ�W�-��s�Xg�W�-��s�X?X�W�-��s�Xk��W�-��s�X���W�-��s�XW��W�-��s�Xb�W�-��s�Xw]�W�-��s�X���W�-��s�XK��W�-��s�XS��W�-��s�X��W�-��s�X���W�-��s�X���W�-��s�X+S�W�-��s�X��W�-��s�X���W�-��s�X/=�W�-��s�X�i�W�-��s�X�\�W�-��s�X�S�W�-��s�Xנ�W�-��s�X�o�W�-��s�X�_�W�-��s�X�J�W�-��s�X���W�-��s�XӤ�W�-��s�XOK�W�-��s�Xs��W�-��s�X7"�W�-��s�XG!�W�-��s�X[��W�-��s�X��W�-��s�XWO�W�-��s�X�q�W�-��s�XC��W�-��s�Xg�W�-��s�X��W�-��s�X[*�W�-��s�X��W�-��s�XOH�W�-��s�X��W�-��s�XgT�W�-��s�X��W�-��s�X�	�W�-��s�X�Q�W�-��s�X���W�-��s�X���W�-��s�X���W�-��s�X'5�W�-��s�X_A�W�-��s�XJ�W�-��s�X�E�W�-��sݞ�r�bm.�z�-ß�rÞ�r�m.�{�Z/0OQ[Qn�����g���g�6#-Þ�rÞ�rÞ�rÒ<-���r���rÞ�r���r��2ß�r��9-Þ�rÞ�rÞ�r�b<-���r�=-ß�m�colÞ�r�*�2ß�râk-Þ�ræn/Þ�r�f<-���rÞ�rß�m��llÞ�r���2ß�rêj-Þ�rîi/Þ�r�n<-���rÞ�rß�m��llÞ�r���2ß�r�vk-Þ�r�Rn/Þ�r�z<-���rÞ�rß�m��llÞ�rÞ--ß�r�Rh-Þ�rÂo/Þ�r�F<-��rÞ�rß�m��llÞ�r�J�2ß�r��f-Þ�rÞ�rÞ�r�V<-���rö=-ß�m��lÞ�r�F�2ß�r�J-Þ�r��l/Þ�r�^<-�c�rÞ�rß�m��llÞ�r���2ß�r��_-Þ�rÞ�rÞ�rê<-���rÎ=-ß�m��lÞ�r�Z�2ß�r�k-Þ�r�vn/Þ�rö<-���rÞ�rß�m��llÞ�r�"�2ß�r��f-Þ�rÞ�rÞ�rþ<-���r�<-ß�m�colÞ�rÊ�2ß�rÂy-Þ�rÒi/Þ�rÆ<-���rÞ�rß�m��llÞ�rÞ�rÞ�rÞ�rÞ�rÞ�r��>-Þ�r��>-�&9-Þ�r�9-Þ�r�9-�b9-�r9-�B9-�R9-�^9-î9-þ9-Ê9-Þ�rÞ9-Þ�rÞ�r��9-Þ�rÞ�rÞ�rÞ�r�v-�v-Þ�r�fv-Þ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�r�_-�_-�j_-�r_-�F_-�N_-�V_-æ_-�I-ö_-þ_-Ò_-��_-��_-Þ�rÞ�rÞ�rÞ�rÞ�r�$�r��v���|�O��r��|�bm��y�O	�L��r��|.:m���b
m�+$}3
�O	���|!)#��|����P��r��^�M��r���r��� ��� ���r���r�3������	������!��������Þ�r���r���r�������3A��4�[���s���wL���J��6���ư�~L��6?��H|.���xb�D���+T� �$SqDr�BV���8�M
��`82R_y>wU�(U�~�>#��h)=)p78�L�^�<g-8�z,8.t��b��r�4)m�-8�Z�\#�]��r�r?-Þ�r���rÞ�r�B?-ê?-�k.Þ�rÞ�r��C�"�Z�r��=�y�2W�r��^��|�^m��=�y�2W�r��^��}*�r���wƘO�3G�j�����#��s�M�^:"�\�Pi	�b
��O�P:5/
�0�}��#w �r��?-Þ�r���r���r�.>-æ?-�k.Þ�rÞ�r��Cø=�y�2W�r��^�*�^
�rÈ=�y�2W�r��^�$�V�r�;�b�^�r�(�V��rð=�y�2W�r��^����r�����=�y�2W�r��^�$�V��r���`2�^�r� �\�L"�W
���|�^�o	�M��r���r���Þ�r�(�V?(�Q
�O��r�"�Z�W��"
�O�l�^�r�"�Z.P�\�r�.�X	�^)bm�'
�|
�Q&��0
�P
�^�M��r�0
�O�l�^�r�"�Z(M���Z)b,M�b
�r�8�M
�`#�Q��;�b�^.P�\�r����Þ�rÞ�r���bÞ�l���m��d#��r���j����S��n���Þ�n���n��m���m���m���m�*�Þ�o���n��d#��j���b�e��S��g#��rÚ�m�t�mÞ�rÞ�rÞ�nÞ�rÞ�Þ����r���n�"�b4��mÆ�n���#��n�)�b�
8-���g#��rÚ�m�t�m������rÞ�rÞ�r��rÞ�r���Þ�l���n��m���m���r���Þ�r���=��m���n��d#�����r���bÞ�r���n?��Þ�r���n?��.Þ�r�"�n?��jÞ�r���n?���Þ�r�h�l?��
?��l���n��d#��ß�=���S��n����m�r�n��d#����r���Þ�r���n?��
Þ�r���n?��fÞ�r���n?<�Þ�d���n��d#��r���b���n������n������n������n������n������n���
���l������l������n���r���2Þ�r���n?��Þ�r���n?��R�rþ�n?��z�rÖ�n?��bÞ�r���l?���q��r�=i?���Þ�r��n?��Þ�rê�n?��"=��l���n��d#�����>=��n���`���r�+
�Q>��r���r�'�] ^�J3�Om�N:-�^:-Þ�n�k.Þ�rÞ�r�Ao�|��O��MZ�:-�V���]þ�r���r�0�v�v�M�r�N:-��:-Þ�n�bk.Þ�rÞ�r�Ac�|��O��MZ�:-�V���]þ�r���r��M�� _
m���r��L�I��25-�5-Þ�n�nk.Þ�rÞ�r�Aw�|��O��MZ5-�V���]þ�r���r����r���r�#+M
�Q�_*�M�^�r�F5-�R5-Þ�n�zk.Þ�rÞ�r�AK�|��O��MZ�5-�V���]þ�r���r�3�^�r�N:-��5-Þ�n�Fk.Þ�rÞ�r�A_�|��O��MZ�5-�V���]þ�r���r�#�b
�M�L.m���r�4�O�s�^(K��r��&��ͤ\-C�m���D���r�N:-�"4-Þ�n�Rk.Þ�rÞ�r�AS�|��O��MZ4-�V���]þ�r���r�
�Q>��W��r���r�/�Q$�^��r�V4-ê4-Þ�n�^k.Þ�rÞ�r�A��|��O��MZ�4-�V���]þ�r���r�*�_*�M���r�N:-��4-Þ�nêk.Þ�rÞ�r�A��|��O��MZ�4-�V���]þ�r���r�'
�s��^m�N:-�67-Þ�nök.Þ�rÞ�r�A��|��O��MZ7-�V���]þ�r���r��M��r���r�#�W7�_�M,�~7-�J7-Þ�nÂk.Þ�rÞ�r�A��|��O��MZZ7-�V���]þ�r���r�$�^*�M��N:-Ò7-Þ�nÎk.Þ�rÞ�r�A��|��O��MZ�7-�V���]þ�r���r�*�T7�T3�O	��~7-��7-Þ�nÚk.Þ�rÞ�r�A��|��O��MZ&6-�V���]þ�r���r�#�b
+Z

,�N:-�6-Þ�n��k.Þ�rÞ�r�A��|��O��MZj6-�V���]þ�r���r��W
��W
�r���r�8�Q�i	
�p8�\�Q��râ6-ò6-Þ�n��k.Þ�rÞ�r�A��|��O��MZ�6-�V���]þ�r���r�7�O?�P
�L-
�Pm�N:-��6-Þ�n��k.Þ�rÞ�r�A��|��O��MZ�6-�V���]þ�r���r�0
�_.�\�v�M�r�N:-�1-Þ�n��k.Þ�rÞ�r�A��|��O��MZb1-�V���]þ�r���r�4�O�
�\%m�N:-�Z1-Þ�n��k.Þ�rÞ�r�A/�|��O��MZ�1-�V���]þ�r�!<�y�2W�r��^���r�N:-�64-Þ�n�"j.Þ�rÞ�r�A#�|��O��MZ�1-�V���]þ�r���r������r�	�z��*0-�60-Þ�n�.j.Þ�rÞ�r�A7�|��O��MZ>0-�V���]þ�r���r�	�y
��*0-�v0-Þ�n�:j.Þ�rÞ�r�A�|��O��MZ~0-�V���]þ�r���r�	�m��*0-ö0-Þ�n�j.Þ�rÞ�r�A�|��O��MZ�0-�V���]þ�r���r�	�h�^��r�*0-��0-Þ�n�j.Þ�rÞ�r�A�|��O��MZ�0-�V���]þ�r���r�	�x!Z 5�M�Q��r�*0-�:3-Þ�n�j.Þ�rÞ�r�Ag�|��O��MZ3-�V���]þ�r���r�	�x(M�l�Q�r���wƘO�3G�j�����#�L�rÞ�r�*0-�F3-Þ�n�jj.Þ�rÞ�r�A{�|��O��MZ�3-�V���]þ�r���r�'�],W
��N:-��3-Þ�n�vj.Þ�rÞ�r�AO�|��O��MZ�3-�V���]þ�r���r�'�]+M
m�N:-�22-Þ�n�Bj.Þ�rÞ�r�AC�|��O��MZ>2-�V���]þ�r���r�'�]!P m�N:-�v2-Þ�n�Nj.Þ�rÞ�r�AW�|��O��MZB2-�V���]þ�r���r�'�]�Q
�T��r�N:-ú2-Þ�n�Zj.Þ�rÞ�r�A��|��O��MZ�2-�V���]þ�r���r�#�b
�Z
m�N:-��2-Þ�næj.Þ�rÞ�r�A��|��O��MZ�2-�V���]þ�r���r�3
�q�_.�^&�_

�O����r����
����Þ�r���r��rÞ�r�N:-�-Þ�nòj.Þ�rÞ�r�A��|��O��MZ~-�V���]þ�r���r�-�N

>,
�O��r�V4-ö-Þ�nþj.Þ�rÞ�r�A��|��O��MZ�-�V���]þ�r���r�$�_$�L%�W.m�V4-��-Þ�nÊj.Þ�rÞ�r�A��|��O��MZ�-�V���]þ�r���r�$�_,
�O$�^!�r�V4-�-Þ�nÖj.Þ�rÞ�r�A��|��O��MZ-�V���]þ�r���r�$�_#�L�r�V4-�N-Þ�n��j.Þ�rÞ�r�A��|��O��MZZ-�V���]þ�r���r�0
�_$�^��r�N:-Ò-Þ�n��j.Þ�rÞ�r�A��|��O��MZ�-�V���]þ�r���r�'
�y�X�Q4�Q����r�0
�p
�t(K!�r�~7-��-Þ�n��j.Þ�rÞ�r�A��|��O��MZ>-�V���]þ�r���r�'
�h	�P;�K.m�~7-�v-Þ�n��j.Þ�rÞ�r�A��|��O��MZF-�V���]þ�r���r�3
�y	�s�Om�N:-þ-Þ�n��j.Þ�rÞ�r�A��|��O��MZ�-�V���]þ�r���r�#�L'�Q��N:-��-Þ�n��j.Þ�rÞ�r�A'�|��O��MZ�-�V���]þ�r���r�'
�y	�l	��N:-�
-Þ�n�*e.Þ�rÞ�r�A;�|��O��MZ-�V���]þ�r���r�7�O%�W�r�N:-�N-Þ�n�6e.Þ�rÞ�r�A�|��O��MZZ-�V���]þ�r���r�2�^>$�L�r���r�'
�|�P?�L��r���wƘO�3G�j�����N:-Ò-Þ�n�e.Þ�rÞ�r�A�|��O��MZ�-�V���]þ�r���r�2�^>,
�O��r�N:-�>	-Þ�n�e.Þ�rÞ�r�A�|��O��MZ	-�V���]þ�r���r�/�Q2�^m�N:-�F	-Þ�n�e.Þ�rÞ�r�Ak�|��O��MZR	-�V���]þ�r���r��]��W��r���r��S
�L��rÊ	-Ú	-Þ�n�fe.Þ�rÞ�r�A�|��O��MZ�	-�V���]þ�r���r��P�^mÊ	-��	-Þ�n�re.Þ�rÞ�r�As�|��O��MZ*-�V���]þ�r���r�.8,s)�.w*�r���r�'
�v�W%�W=�V*���r�b-�r-Þ�n�~e.Þ�rÞ�r�AG�|��O��MZJ-�V���]þ�r���r�'
�h	�P�r�~7-Â-Þ�n�Je.Þ�rÞ�r�A[�|��O��MZ�-�V���]þ�r���r�'
��O�Z�H��r�~7-��-Þ�n�Ve.Þ�rÞ�r�A��|��O��MZ�-�V���]þ�r���r�'
�s�Q�r�~7-�-Þ�nâe.Þ�rÞ�r�A��|��O��MZ-�V���]þ�r���r�'
�h	�P;�M�s�^$_��r�~7-�V-Þ�nîe.Þ�rÞ�r�A��|��O��MZ�-�V���]þ�r���r�'
�h	�P#�Q.m�~7-��-Þ�núe.Þ�rÞ�r�A��|��O��MZ�-�V���]þ�r���r�'
�h	�P;�K#�Q���r�~7-�2
-Þ�nÆe.Þ�rÞ�r�A��|��O��MZ

-�V���]þ�r���r�3�H7�_m���r���<���r�25-�B
-Þ�nÒe.Þ�rÞ�r�A��|��O��MZZ
-�V���]þ�r���r�3
�h	�P;�K.m�25-Ò
-Þ�nÞe.Þ�rÞ�r�A��|��O��MZ�
-�V���]þ�r���r�3
�h	�P?�L��r�~7-��
-Þ�n��e.Þ�rÞ�r�A��|��O��MZ*-�V���]þ�r���r�%�]

�Z�H��r�25-�b-Þ�n��e.Þ�rÞ�r�A��|��O��MZr-�V���]þ�r���r�3�O�P2�L7�_m�~7-ê-Þ�n��e.Þ�rÞ�r�A��|��O��MZ�-�V���]þ�r���r� "�o!�x��r�*0-��-Þ�n��e.Þ�rÞ�r�A��|��O��MZ�-�V���]þ�r���r��W
�<����r�3�W
*�^�^!�r�:-�
-Þ�n��e.Þ�rÞ�r�A+�|��O��MZ-�V���]þ�r���r�'
�s�^ ^�J)�P��r�b-�R-Þ�n�&d.Þ�rÞ�r�A?�|��O��MZ�-�V���]þ�r���r�$�^2�^2�J�V2�^��r�N:-��-Þ�n�2d.Þ�rÞ�r�A3�|��O��MZ�-�V���]þ�r���r�'
�s�^�Z
��N:-�2-Þ�n�>d.Þ�rÞ�r�A�|��O��MZ-�V���]þ�r���r�-�N

>$�L�r�N:-�z-Þ�n�
d.Þ�rÞ�r�A�|��O��MZJ-�V���]þ�r���r�3�S�o�b�r�N:-Â-Þ�n�d.Þ�rÞ�r�Ao�|��O��MZ�-�V���]þ�r���r�0
�N
�[
�_��r���r���?Þ�r�N:-��-Þ�n�bd.Þ�rÞ�r�Ac�|��O��MZ&-�V���]þ�r���r�.�\��*�Mm�N:-�-Þ�n�nd.Þ�rÞ�r�Aw�|��O��MZn-�V���]þ�r���r�.�\��"�K�r�N:-æ-Þ�n�zd.Þ�rÞ�r�AK�|��O��MZ�-�V���]þ�r���r�/�Q.�\��V4-��-Þ�n�Fd.Þ�rÞ�r�A_�|��O��MZ�-�V���]þ�r���r�#�b
�P�^
>3�S�O��r�N:-�2-Þ�n�Rd.Þ�rÞ�r�AS�|��O��MZ-�V���]þ�r���r�2
�V	�O?�P
�L��r�N:-�F-Þ�n�^d.Þ�rÞ�r�A��|��O��MZZ-�V���]þ�r���r�'
�w�W&�Y.må@ao���uJ̉]��$N:-Ò-Þ�nêd.Þ�rÞ�r�A��|��O��MZ�-�V���]þ�r���r�'
�i�Z(K!�r�N:-�* -Þ�nöd.Þ�rÞ�r�A��|��O��MZ: -�V���]þ�r���r��\>��W��r���r��x)M	�M"
�\�O	���r�r -�F -Þ�nÂd.Þ�rÞ�r�A��|��O��MZ� -�V���]þ�r���r�'
�v�W'�Q���r�V4-Ú -Þ�nÎd.Þ�rÞ�r�A��|��O��MZ� -�V���]þ�r���r�'
�v�W%�W=�V.m�V4-�&-Þ�nÚd.Þ�rÞ�r�A��|��O��MZ:-�V���]þ�r���r�'
�w�s�q���r�V4-�r-Þ�n��d.Þ�rÞ�r�A��|��O��MZF-�V���]þ�r�~7-��-Þ�n��d.Þ�rÞ�r�A��|��O��MZ�-�V���]þ�r���r��b>��W��r���r�0
�~�i�^!�r��-��-Þ�n��d.Þ�rÞ�r�A��|��O��MZ�-�V���]þ�r���r�%�b(Q�P�Q8�M	�L!�r�N:-�-Þ�n��d.Þ�rÞ�r�A��|��O��MZj-�V���]þ�r���r� �\&�Sm�25-â-Þ�n��d.Þ�rÞ�r�A/�|��O��MZ�-�V���]þ�r���r��W
�r���r�0��L?�Z�^
m��-��-Þ�n�"g.Þ�rÞ�r�A#�|��O��MZ�-�V���]þ�r���r�,�[�P�J�V��r��-�>-Þ�n�.g.Þ�rÞ�r�A7�|��O��MZ-�V���]þ�r��-�.-Þ�n�:g.Þ�rÞ�r�A�|��O��MZF-�V���]þ�r���r�0
�|
�^+
���-þ-Þ�n�g.Þ�rÞ�r�A�|��O��MZ�-�V���]þ�r���r�0
�~�t(K!�r��-��-Þ�n�g.Þ�rÞ�r�A�|��O��MZ�-�V���]þ�r���r�0
�r
�J4�N*���r��-�
-Þ�n�g.Þ�rÞ�r�Ag�|��O��MZ-�V���]þ�r���r�0
��O5�W
,��-�V-Þ�n�jg.Þ�rÞ�r�A{�|��O��MZ�-�V���]þ�r���r�0
�l�b
�~.m��-Þ-Þ�n�vg.Þ�rÞ�r�AO�|��O��MZ�-�V���]þ�r���r�0
��O �J!�r���r������������?Þ�rÞ�r��-�&-Þ�n�Bg.Þ�rÞ�r�AC�|��O��MZ-�V���]þ�r���r�0
�|
�O �J%,��-�J-Þ�n�Ng.Þ�rÞ�r�AW�|��O��MZZ-�V���]þ�r���r�0
�p
�t,��-Ò-Þ�n�Zg.Þ�rÞ�r�A��|��O��MZ�-�V���]þ�r���r�0
�|
�O �J!�r��-��-Þ�næg.Þ�rÞ�r�A��|��O��MZ&-�V���]þ�r���r�3
�_-
�L���r�~7-�-Þ�nòg.Þ�rÞ�r�A��|��O��MZn-�V���]þ�r���r�'
�#�r�25-æ-Þ�nþg.Þ�rÞ�r�A��|��O��MZ�-�V���]þ�r���r����r���r�3�^�}
m���r�'
��^2�^!�r��-��-Þ�nÊg.Þ�rÞ�r�A��|��O��MZ�-�V���]þ�r���r�3
�l�O/W"�_�r��-�
-Þ�nÖg.Þ�rÞ�r�A��|��O��MZ-�V���]þ�r���r�'+$��.w*�r���r� �}
m�V-æ-Þ�n��g.Þ�rÞ�r�A��|��O��MZ�-�V���]þ�r���r�3
�|�P?�L��r�25-��-Þ�n��g.Þ�rÞ�r�A��|��O��MZ�-�V���]þ�r���r�-�h�y N
�S

"]
�O�r�~7-�.-Þ�n��g.Þ�rÞ�r�A��|��O��MZ
-�V���]þ�r���r�'
�w�\)M	�l�Q,�N:-�B-Þ�n��g.Þ�rÞ�r�A��|��O��MZZ-�V���]þ�r�>��N>ͻ~x���8P<.N:-��-Þ�n��g.Þ�rÞ�r�A��|��O��MZ�-�V���]þ�r���r�'
�	�y
�l�^!�r�N:-��-Þ�n��g.Þ�rÞ�r�A'�|��O��MZ*-�V���]þ�r���r�'
�y	��Z �^.m�V4-�b-Þ�n�*f.Þ�rÞ�r�A;�|��O��MZv-�V���]þ�r���r�3'*^?�O%�P&)w	���r�:-î-Þ�n�6f.Þ�rÞ�r�A�|��O��MZ�-�V���]þ�r���r�3'*^8�^�W$�_!P�Zm�:-��-Þ�n�f.Þ�rÞ�r�A�|��O��MZ�-�V���]þ�r���r�3
�y	�o	��V4-�-Þ�n�f.Þ�rÞ�r�A�|��O��MZ-�V���]þ�r���r�3�O�Z
�P$�^2�^��r�N:-�V-Þ�n�f.Þ�rÞ�r�Ak�|��O��MZ�-�V���]þ�r���r�$�^2�^2!P�y	�o	��N:-��-Þ�n�ff.Þ�rÞ�r�A�|��O��MZ�-�V���]þ�r���r�'
�y	�o	��V4-�6-Þ�n�rf.Þ�rÞ�r�As�|��O��MZ-�V���]þ�r���r�'
�o�b(�Q
�O��r�N:-�z-Þ�n�~f.Þ�rÞ�r�AG�|��O��MZN-�V���]þ�r���r�3
�o�b(�Q
�O��r�N:-Æ-Þ�n�Jf.Þ�rÞ�r�A[�|��O��MZ�-�V���]þ�r���r��|
�O(�S�^7�_,�r -��-Þ�n�Vf.Þ�rÞ�r�A��|��O��MZ*-�V���]þ�r���r�))^ �X�M�Q�r�V4-�b-Þ�nâf.Þ�rÞ�r�A��|��O��MZv-�V���]þ�r���r�'
�n
�q���r��-î-Þ�nîf.Þ�rÞ�r�A��|��O��MZ�-�V���]þ�r���r�'
�s�^%^m�N:-��-Þ�núf.Þ�rÞ�r�A��|��O��MZ�-�V���]þ�r���r�?`�� _
m���r��Q�r�>-�-Þ�nÆf.Þ�rÞ�r�A��|��O��MZ-�V���]þ�r���r�	�W�Z��W��r���r�!�P�^!�x�\*�o	�^$�V3�\�r�N-â-Þ�nÒf.Þ�rÞ�r�A��|��O��MZ�-�V���]þ�r���r�!�P�^!�x�_*�o	�^$�V3�\�r���r�	������������������rÞ�r�N-��-Þ�nÞf.Þ�rÞ�r�A��|��O��MZ-�V���]þ�r���r�3
�o(Q��N-�z-Þ�n��f.Þ�rÞ�r�A��|��O��MZF-�V���]þ�r���r�)?�W.�z��r���r�'
�o�b �þ-Î-Þ�n��f.Þ�rÞ�r�A��|��O��MZ�-�V���]þ�r���r�%�V.�\�^�r�b-��-Þ�n��f.Þ�rÞ�r�A��|��O��MZ"-�V���]þ�r���r�%�V.�\�v�Wm�b-�-Þ�n��f.Þ�rÞ�r�A��|��O��MZn-�V���]þ�r���r�'
�w�~�M��r�N:-æ-Þ�n��f.Þ�rÞ�r�A+�|��O��MZ�-�V���]þ�r���r�$�V ^�X.m���r���<Þ�r�N:-��-Þ�n�&a.Þ�rÞ�r�A?�|��O��MZ�-�V���]þ�r���r�'
�|�^�M�L&��N:-�-Þ�n�2a.Þ�rÞ�r�A3�|��O��MZ-�V���]þ�rö����kÞ�r3��%#��s�
8-ß�rß�rÞ�r��m�.�m#��s�:�i#��s�	�rÚ8-Þ�rÞ�rÞ�r�6�r������rÞ�rÞ�rñ�rÞ�r��e#��sÞ�rÞ�rÞ�rÞ�rÞ�r�j�e#��sÞ�rÞ�rÞ�r�N?���<z�e#��sÞ�rÞ�rÞ�rÞ�rÞ�r�J�e#��sÞ�rÞ�rÞ�rÞ�rþ=���:Þ�n���n��m���m���m���m���Þ�r���n?��Þ�l���n��m���i���mÞ�r���r�#�b
 N
���r���r�/�Q3
�I	���r���r���������<Þ�r�N:-ê-Þ�n�>a.Þ�rÞ�r�A�|��O��MZ�-�V���]þ�r���r�0
�^�v�K��r�N:-��-Þ�n�
a.Þ�rÞ�r�A�|��O��MZ*-�V���]þ�r���r�7�O$�l	�W<�U��N:-�b-Þ�n�a.Þ�rÞ�r�Ao�|��O��MZv-�V���]þ�r���r�7�Z
�����r�"
�^
�M
(�\
(Q���rî-þ-Þ�n�ba.Þ�rÞ�r�Ac�|��O��MZ�-�V���]þ�r���r�%�V3
�I	�L3�O,��-��-Þ�n�na.Þ�rÞ�r�Aw�|��O��MZ"m-�V���]þ�r���r�/�Q3( b�^.m��-�m-Þ�n�za.Þ�rÞ�r�AK�|��O��MZjm-�V���]þ�r���wƘO�3G�j������-þ-Þ�n�Fa.Þ�rÞ�r�A_�|��O��MZ�m-�V���]þ�r���r�3�M8�M�^!�r��-��m-Þ�n�Ra.Þ�rÞ�r�AS�|��O��MZ�m-�V���]þ�r���r�#�L8�M�^&�_

m��-�.l-Þ�n�^a.Þ�rÞ�r�A��|��O��MZl-�V���]þ�r���r�1�M8�M�^#�Y	,��-�zl-Þ�nêa.Þ�rÞ�r�A��|��O��MZNl-�V���]þ�r���r�1�M8�M�^3�Om��-Æl-Þ�nöa.Þ�rÞ�r�A��|��O��MZ�l-�V���]þ�r���r�%�V"
�^�Q8�M�^.m��-��l-Þ�nÂa.Þ�rÞ�r�A��|��O��MZ*o-�V���]þ�r���r�#�O�l�Z
m��-�bo-Þ�nÎa.Þ�rÞ�r�A��|��O��MZro-�V���]þ�r���r�3
�h	�P#�Q.m�25-êo-Þ�nÚa.Þ�rÞ�r�A��|��O��MZ�o-�V���]þ�r�25-�J7-Þ�n��a.Þ�rÞ�r�A��|��O��MZ�o-�V���]þ�r���r�3
�l�^?�H�O��V4-�&n-Þ�n��a.Þ�rÞ�r�A��|��O��MZ:n-�V���]þ�r���r�'
�|�^�M�L�r�N:-�rn-Þ�n��a.Þ�rÞ�r�A��|��O��MZFn-�V���]þ�r���r��b>��r���r�/�Q.�\�o �Q��rþn-În-Þ�n��a.Þ�rÞ�r�A��|��O��MZ�n-�V���]þ�r���r�*�T�M	�W�i�^!�r���r���=Þ�rþn-��n-Þ�n��a.Þ�rÞ�r�A/�|��O��MZ>i-�V���]þ�r���r�!�N�P
�s�Z

�^�rþn-�vi-Þ�n�"`.Þ�rÞ�r�A#�|��O��MZNi-�V���]þ�r���r�%�O7�_�~�r�~7-Æi-Þ�n�.`.Þ�rÞ�r�A7�|��O��MZ�i-�V���]þ�r���r�
�M���r�N:-��i-Þ�n�:`.Þ�rÞ�r�A�|��O��MZ�i-�V���]þ�r���r�
�M

�h��r�N:-�h-Þ�n�`.Þ�rÞ�r�A�|��O��MZh-�V���]þ�r�����dÞ�r3��m���m���o�"�m�&�m�6�m�:�m��nó'�X������+%���#G+�G��pW΂m��(Þ�r�5����rß�þqÞ�þLÎ��n>m���r����
����r���r�5���������7����������*�����)��r���nÞ�m���n7��i���Þ�r���Þ�lÞ�rÞ�i���Þ�j���n���r���fÞ�rÞ�r���bÞ�o���n��i���rÞ�n���f���rê�r�cÞ�r3��i"��s�	�r�d-�p�H8ua���1aX݄����#��sÞj-�X݄���Ɯ
Ք�g!N�m#�Dr�R�m#,�s�V�i"�qr��̶���ß����ß����ß����ß�U���ß��#�������&�î��&k���V����<��M����<��}����<��y����<��u���=ß�l#�=�y�2W�r��^���rÞ�r���r�7����������r���r�3�������r���jÞ�rÞ�r���r��^)�Q�S�{�^�r�1�������r��Þ��J�n��m���m���m���m���m���m���m���m���m���i"�V�	�� Bk-�5zsW΂m�<�rÎ����g#�����m#����g#��>���g#��:���g#��6���g#��0���g#��2�"�g#��.�&�g#��*�*�g#��&�2�g#����6�g#����:�g#����>�g#�����m#����m# ���
�m#����g#�����g#�����g#�����g#�����g#�����g#�����g#�����m#����b�g#����f�m#7���j�m#/���n�g#����p�g#���r�m#���v�g#���x�g#���z�g#���~�g#���B�g#���F�g#�����fÞ�l���n��m���m���fÞ�l���n��o���m���nÞ�m���n��i"��r�	�r�jd-�p�H8ua���1aX݄�0������	������?�(�	����rÞ�r��r�&�'�*�!�:���������������-���������������7������������#���������������������:������:�r�����������rÞ�rÞ�r���r���r��r�&�'�#���:���������������-���������������7������������#���������������������:������:�r�4),	�(!w��r���r���r���r���rÞ�rÞ�rÞ�rÞ�r���wƘO�3G�j�������wƘO�3G�j�������r��g-��g-Þ�r���r���r���r���Þ�r���r���
�.�%�"�4���r���r���r���r���<��� ��� ��� ���r��g-�`.���r���r����Jvtp�}@�Yw)�|))~\v�
���3f�SRC�axCa�oV>J�^;��x|z��~�I=�=�y�2W�r��^�2
�O��r��v���l�Ð=�y�2W�r��^��l����"Þ�rÞ�r���Þ�r���n?���Þ�r�2�n?��Þ�r���n?��nÞ�m���n7��i�&�rÞ�r�"�^;��mò�n7������n���b�&a-���g#��rÚ�m�t�m������rÞ�rÞ�rÕ�rÞ�r�"�nĞ�m��i7������n���b�>a-���g#��rÚ�m�t�m���ò�rÞ�rÞ�r���r���r���r�-8,|-�<���r��l�b<�^�r���r���rÊa-Öa-Þ�n�`.Þ�rÞ�r�Ao�|��O��MZ�a-�V���]þ�r���r��l�b(�P
mÊa-�&`-Þ�n�b`.Þ�rÞ�r�Ac�|��O��MZ6`-�V���]þ�r���r��l�b?�^�^&
�_mÊa-�n`-Þ�n�n`.Þ�rÞ�r�Aw�|��O��MZF`-�V���]þ�r���r��l�b:�S
�b
%^�M��rÊa-þ`-Þ�n�z`.Þ�rÞ�r�AK�|��O��MZ�`-�V���]þ�r���r��l�b(�Q
�O��rÊa-��`-Þ�n�F`.Þ�rÞ�r�A_�|��O��MZ&c-�V���]þ�r���r��l�b9�LmÊa-�c-Þ�n�R`.Þ�rÞ�r�AS�|��O��MZnc-�V���]þ�r���r��l�b8�E�rÊa-æc-Þ�n�^`.Þ�rÞ�r�A��|��O��MZ�c-�V���]þ�r���r��V�r���r��^)*^+�I#�L!�r��c-��c-Þ�nê`.Þ�rÞ�r�A��|��O��MZ�c-�V���]þ�r���r��^)*^=�V"
�L��r��c-�b-Þ�nö`.Þ�rÞ�r�A��|��O��MZb-�V���]þ�r���r��V��W
�r���r��^'
�o	��Rb-âb-Þ�nÂ`.Þ�rÞ�r�A��|��O��MZ�b-�V���]þ�r���r��^)"Sm�Rb-��b-Þ�nÎ`.Þ�rÞ�r�A��|��O��MZ�b-�V���]þ�r���r��^)�M�M'�b
��Rb-�*}-Þ�nÚ`.Þ�rÞ�r�A��|��O��MZ>}-�V���]þ�r���r���Þ�r�Rb-új-Þ�n��`.Þ�rÞ�r�A��|��O��MZ~}-�V���]þ�r���r��^),_)�Y
��Rb-ö}-Þ�n��`.Þ�rÞ�r�A��|��O��MZ�}-�V���]þ�r���r��^)�O��Rb-��}-Þ�n��`.Þ�rÞ�r�A��|��O��MZ�}-�V���]þ�r���r��^)�Om�Rb-�|-Þ�n��`.Þ�rÞ�r�A��|��O��MZ|-�V���]þ�r���r��^)�^
��Rb-�F|-Þ�n��`.Þ�rÞ�r�A/�|��O��MZR|-�V���]þ�r���r��^).W��Rb-Ê|-Þ�n�"c.Þ�rÞ�r�A#�|��O��MZ�|-�V���]þ�r���r��^/�p
����r������������ ��������r���r���?Þ�r�Rb-��|-Þ�n�.c.Þ�rÞ�r�A7�|��O��MZ-�V���]þ�r���r��^/�s
�b
%^�M��r�Rb-�~-Þ�n�:c.Þ�rÞ�r�A�|��O��MZV-�V���]þ�r���r��^/�n�^�^&
�_m�Rb-Î-Þ�n�c.Þ�rÞ�r�A�|��O��MZ�-�V���]þ�r���r��^/�h�^��r�Rb-��-Þ�n�c.Þ�rÞ�r�A�|��O��MZ.~-�V���]þ�r���r��^/�|
�^��r�Rb-�f~-Þ�n�c.Þ�rÞ�r�Ag�|��O��MZv~-�V���]þ�r���r��^/�m�O��r�Rb-î~-Þ�n�jc.Þ�rÞ�r�A{�|��O��MZ�~-�V���]þ�r���r��^/�s�^��r���r����Þ�r�Rb-��~-Þ�n�vc.Þ�rÞ�r�AO�|��O��MZ�~-�V���]þ�r���r��^/�m�bm�Rb-�
y-Þ�n�Bc.Þ�rÞ�r�AC�|��O��MZy-�V���]þ�r�V4-��:-Þ�n�Nc.Þ�rÞ�r�AW�|��O��MZNy-�V���]þ�r�b�����nÞ�rÞ�m���iß�rÞ�s���r������rÞ�rÞ�r���r���r���p���iß1Þ�s���jN�����rÞ�rÞ�r���r���r���c#.���s1Ba-��s۟�r���rß�r�#��������Þ�r���r���r���r�,���*�&Þ�r���r�������Þ�r�<�y�2W�r��^���r���r��r�J�r���rÞ�rÞ�r���rÞ�rÞ�r���rÞ�rÞ�r���rÞ�rÞ�r���rÞ�rÞ�r���rÞ�lÞ�i=��rÞ�rÞ�r���rÞ�rÞ�r���rÞ�rÞ�r���rÞ�rÞ�r���rÞ�rÞ�<ß�m�F�lÞ�i=��rÞ�rÞ�r���rÞ�lÞ�i=��rÞ�Þ�i=��rÞ�fÞ�r���rÞ�rÞ�r���rÞ�rÞ�r���rÞ�`Þ�i=��rÞ�rÞ�r���rÞ�lÞ�i=��rÞ�rÞ�r���rÞ�rÞ�r���rÞ�nÞ�r���rÞ�bÞ�nÞ�rÞ�r���sß�lÞ�rÞ�mÞ�r���r���mÞ�r���rÞ�mÞ�r���r�����������������r���r�:�=�������Þ�rÞ�r���r�4�!�7������3������	���� �����r���r�4�!�7������5������������Þ�r���r�3���3�-����	���������Þ�r���r����������������Þ�r���r����������������Þ�r���r�3�,�	���"���
� �"�&�*�r���r�������	���� �������
�r���r�������	��Þ�r���r�:�r���r�:����������?����Þ�r���r�����������r���r�.����������(�	�����Þ�r���r���r���r���r���r�:����������?��������	�������
��Þ�r���r�#���3���/�!Þ�r���r���r���rÞ�rÞ���r���rÞ�r���r�:����������?�����������������������Þ�r���r������������<��������r���r�:����������?��������� ����
�r���r���r���r��������������������������Þ�r���r�������+�r���r�	�r���r��r���r�� ��r���r��r���r� �r���r� � ��r���r��r���r��r���r�����	�������	Þ�r���r������������	Þ�r���r�:����������?���r���r�����������	�����r���r������Þ�r���r�����������������	�����r���r�/�����Þ�r�#��h)=)p78�L�^�<g�];��W:�r�4)�n,�r�
4-Þ�r���r���r�Rw-öw-�Zc.Þ�rÞ�r��C���Þ�r���n?��:�r���n?��r�,�N�l�^&�Y�b�Q��r��-��w-Þ�n�^c.Þ�rÞ�r�A��|��O��MZ�w-�V���]þ�r�)�O	�Z
m�1�M�r�2
�V	�O�r�)���	���	���
�����Þ�r���r���
Þ�r���r������������Þ�r���r���2���r���r������������������Þ�r���r��r������������Þ�r���r���r��������������r��r�3�#�$���7�-�0�)�:�!�	������������:���	���������:�/����������4������	������5���	���������
�r�l�r�&�'�%���?�&�/�/�!�&�?�!�!�/�&�%�,�)�:���/�(�2���!���%���-���������������7������������#���������������������:������������
���:�r���r�"������
���� �����r���r�"������
��������������Þ�r���r�.��� ���	�������r���r�5���	���������
������	����r���r���r���r�2�r���r�3�r���r�0�r���r���r���r���r���r���r���r���r���r���r���r�#�#�-���.�)�#�r���r�:����������?��������������� �����r���r�"�r���r����
����������
��Þ�r���r�5���*�.��������������(�	����-Þ�r���r������Þ�r���r�!�4�:�r���r�3���������	���� �$���
���3���������/��������Þ�r�'����(�	����r�"������*������-�����������Þ�r�'����(��������r�"������#����������r�"������*������!�����������Þ�r���r�3���������.���������������)������!�r�������������������
�����Þ�r���r��� ������Þ�r���r��� ������Þ�r���r��� ������Þ�r�������?���	����r����������������
�����Þ�r���r���r���r�7������	���� �3������
�r���r�;�r���r�=�����#����������������������
�����������r���r���dÞ�rÁ=�y�2W�r��^���r�=��;�r���r�=�Þ�r��=�y�2W�r��^��{�G3kQm���f���r�������r�:����������?��������	����������������������r���r�	�������r���r�7��� �/���Þ�r���r�0�)�'���"���/���"�rÞ�r���r�0�)�'���3��Þ�r���r�0�)�'��� �%�,�-�0��Þ�r���r�0�)�'���%���.�-�,�.�?���8�r���r�0�)�'���-���*���)���3��Þ�r���r���������Þ�r���r����������� ��������)���r���r���Þ�r� �r�:�%������������%������������:������������� ��������r���r��� �����r���r������������r���r�������Þ�r���r����������r�	��������������Þ�r���r������������<������������Þ�r�������������	����r�3����������r���r��� �����Þ�r�0������	������?�.�����r�#�������r�"���������,�����Þ�r���r����	�������
�����r���r�"����r���r�����������r���r�3���3���%�!�:����������r���r�"����������r���r������r���r�3���3���%�!�:�/����������3����r���r�:��������������Þ�r���r�3�������r���r�-��Þ�r���r�.�)Þ�r�V��&3[m���6���r��� Þ�r���r�,����r�����r�3������	���������&������%���!�r���r�#���
���,������&������%��Þ�r���r������r���r�=�r���r�'����-�������+�����������Þ�r���r��(Þ�r���r��r���r����&�%�$�������)�+�&����r���r��-�0���/�������.��Þ�r���r��-�0���/�����.�/���,��Þ�r���r��-�0���/�����&�%�(�2��Þ�r���r��-�0���/�������)�+�&����r���r��)�3�/��r���r��.�%�&��r���r��*�/�!�%��Þ�r���r��)�,�.��r���r��"�!�+�%��5�"��r���r��"�!�+�%��"�#�7� ��r���r��"�!���2�)��r���r�� �5�!��r���r�� �5�!�.�-�"������r���r�� �5�!�.�-�"������r���r�� �5�!�.�-�"������r���r�� �5�!�.�-�"������r���r��,�!�/�+��Þ�r���r��-�#�/�%� �2����r���r����!�,��r���r��/�!�"�3��*�#�#�'��r���r����2���'��*�)�$����r���r����2���'��0�%�'�*�2��Þ�r���r����)� �"�#�7����r���r��-�*����r���r��-�*���'����r���r�3�����Þ�r���r�/����r���r��/�/� �2�)�6�����!�%� �5��Þ�r���r���r���r���r���r�?�r���r���r���r���r���rú�r���rÚ�r���rô�r���rÔ�r���râ�r���rÂ�r���rÿ�r���r�N�r���r�<�r���r���r���r���r���r�G�r���r���r���r���r���r���r���r����/�&�*��Þ�r���r��"�0�%�,����r���r��"�!���3�)��r���r��/�!�&�#���*�-�2�#�0��Þ�r���r����/�&�5�!�%��5�"��r���r����/�&�5�!�%��"�#�7� ��r���r��!�5���%��Þ�r�������	��������� ����r���r��"�*�-�9�����.�-�5���%��Þ�r���r��"�0�)�4�%�/���3��2�%�2�&�%��Þ�r���r�� �%���2��2�%�2�&�%��Þ�r���r��)�-�-�)�&��r���r��,�0�#�7���%����r�j�r�&�'�%���?�&�/�/�!�&�?�!�!�/�&�%�,�)�:�*�!���"���!���%���"�)�3�/�0�%�.���)�#�,���3���������:�/����������.��������������������!�&��Þ�r�%������1�������r�#���������� �����r�"������
���� �����r���r���
�4������	����4���r���r�(���
�rÞ�r�|�r�&�'�%���?�&�/�/�!�&�?�!�!�/�&�%�,�)�:���/�(�2���!���%���-���������������7�����������,���:�/����������4������	������0���������������/�������r���r��� ���r���r�7����<������r���r��� ���r���r�7������.�r���r��� ���r���r�7�������������������?Þ�r���r��� ���r���r�7������	�����Þ�r���r�����������������:�r���r�:���������3������������#��������Þ�r���r�3���
������������������$���������
���.����������r���r�!����r���r�3���
������������������!������4�������"���������Þ�r�2�r�&�'�%���?�/�*�-�3���%���?���/�#�2���&���2�"�:������
���:��������������������Þ�r����&3[m���6���&3[m���6���r��A-�*@-Þ�r���r�3����r���r�-����r���r�2�����Þ�r���r�7����r���r�2�����Þ�r���r�$���	�r���r�3����r���r�(����r���r�$��� �r���r�-����r���r�!����r���r�-����r���r�(����r�@�֏ӽ�vD��}���@�O���{n���8P]#��nÞ�r���m?��r�#�b
.P�O		�^"(m��-��@-Þ�nêc.Þ�rÞ�r�A��|��O��MZ2C-�V���]þ�r�~7-æ-Þ�nöc.Þ�rÞ�r�A��|��O��MZfC-�V���]þ�r���r�#�b
)z 8�\�Q��r��-�^C-Þ�nÂc.Þ�rÞ�r�A��|��O��MZ�C-�V���]þ�r��-æ-Þ�nÎc.Þ�rÞ�r�A��|��O��MZ�C-�V���]þ�r���r�3
�^"]
�O��r��-��C-Þ�nÚc.Þ�rÞ�r�A��|��O��MZ.B-�V���]þ�r���r�"
�^
"]
�O��r��-�fB-Þ�n��c.Þ�rÞ�r�A��|��O��MZvB-�V���]þ�r���r�"
�^
)|��r��-îB-Þ�n��c.Þ�rÞ�r�A��|��O��MZ�B-�V���]þ�r���r�*�_)�X.m�~7-��B-Þ�n��c.Þ�rÞ�r�A��|��O��MZ�B-�V���]þ�r���r��]8��W��r���r�4�sm�6]-�
]-Þ�n��c.Þ�rÞ�r�A��|��O��MZ]-�V���]þ�r���r�'
�p �\.m��-�J]-Þ�n��c.Þ�rÞ�r�A/�|��O��MZV]-�V���]þ�r���r�#�b
.P�O		�^ �Vm��-Î]-Þ�n�"b.Þ�rÞ�r�A#�|��O��MZ�]-�V���]þ�r���r�/�Q#�S �M�r�~7-��]-Þ�n�.b.Þ�rÞ�r�A7�|��O��MZ.\-�V���]þ�rñ=�y�2W�r��^���r�#�L(�Z	�bm�~7-�v\-Þ�n�:b.Þ�rÞ�r�A�|��O��MZF\-�V���]þ�r���r�3
�|
�]�_"�b��r�~7-þ\-Þ�n�b.Þ�rÞ�r�A�|��O��MZ�\-�V���]þ�r���r�%�O(�Z	�bm�~7-��\-Þ�n�b.Þ�rÞ�r�A�|��O��MZ�\-�V���]þ�r�#�J2.W	�P��#�b
)z �r�#�b
m� �^?�M3�Q*�^��r�7�O�r�&
�Xm�*�_.�O�}
m�.�Q?�\�^��r�+�]��r�"&/l�Z/Z�O�r�0�_�L)�O�r�#�b:��0
�b�^��r����Þ�rÞ�r�)<�y�2W�r��^���r���������r���r���������r���r������� ��Þ�r���r�������Þ�r���r���	��������1����/����������N�Þ�r���r���*�6�r�3�#�$���7�-�0�)�:�!�)�/�0�#�3�#�$���:���	����������� �2���#��������������������Þ�r���r�"���������
�"����������)��Þ�r���r� �/�"�(�'�*�(�'�-�"�1���2���7���9�<���>���;���5Þ�r�"���
������$���
�����Þ�r���r�?�������r���r��� ���r���r����������������Þ�r���r��������Þ�r���r���������������
������
�������r���r���>Þ�r���r������������>Þ�r���r�3���3������������.���	���	�������r������rÞ�rÞ�r���rÞ�r�$�r�3�)�*�)�#��������(�0�#�-��7����?�����4�������/����������
����r���r���������������r�"������������	����r���r�4���������
�,������+�������	�����!����������r������rÞ�rÞ�r���rÞ�r���r�"�&�*��������������rÑ=�y�2W�r��^������rÞ�rÞ�r���rÞ�r���r�7������)���/�����Þ�r���r�������)���.����������*�����������r���r�������)���.����������*��������r���r�������)���!����,�����������r���r�������)���!����,��������r���r��������������#�����r���r��������������"����������&��������Þ�r���r��������������"����������&���������?��Þ�r���r�������)���3�������r���r��������������/����������?��Þ�r���r��������������/���������Þ�r���r����������������������������&���������?��Þ�r���r����������������������������&��������Þ�r���r��������������/�
�����Þ�r���r�������)���3�����Þ�r���r�������)���5���.����������*��������r���r�������)���5���.����������*�����������r���r�������)���#�������r���r����������������	����rß�<��dN�H=6'H��}���uo��(y5�s����#��w���Ua�H���s�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�mÞ&mÞ�k��|����i�$�V��.m��sß�	>�*�M�r��r��Þ�������%��.�$�s=��r���rO�^m=��r��&��m���rÞ|l �r92�Pr?��r���rO P
m4�mÞ�r0��j���r���rÞ�n�2
�O��nÞ�r�-��������rÞ|l �r92�Pr?��r���r\�^m?��rL�����5n���r���r<��rß�<��4I|�V�"O�`���W�eII��!N'V5�q�#��w���Ua�H���s�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�oÞ�rÞ�l�$�r6��r]��r��(P<�����YÞWgÞ�kÞ�nÞ(m���rÞ�h�$�V�r<��rÞ�rÞ��8'��r��?mÞ�h�*�^
�r���rm�I��^�M��sß�iӞl�m-��=�����r��Po �r6-8l�#3
�Z�o<��r���rO/w��o���r8�r��|kÞ�n"��r?���Z�r��d��l���r���r\��s��m��r����o�L
�ß�rv34�Q�T*�7�L����r*)d���r��)9-��rÅ�rÅ�r�p����hÞ�rÞ�rÞ�rÞ�r��$nÞ�j8��s?�rC��r?�.b�s.�#�h	�P !Z ��Z�\�mÞ�&}��
Þ�|��jÞ�I<��I<���m�r���rÞ�rÞ�rÞ�rÞ�5{��rN�rß��ÞldÞ�rH3�^m���!l7�L�w		h	�P m�w �r��r"#�;��r���r���r��b	Þ�rÞ�rÞ�rÞ�rÞ�r
��r���kÞ�nY���5��i�"�Z�s.�#�h	�P !Z ��Z�\�mÞ�&}��
Þ�|��jÞ�I<��I<���m�r���rÞ�rÞ�rÞ�rÞ�5Ӟ�rN�rß�Þ�i8��M!�J��o���r8>�r���nÞ�n���9��d��|�^m4��r=���,��kC��r;��rß�n�"�-Þ�rÞ�r�"�-Þ�rÞ�rÞ�rÞ�rÞ�rÞ�r�
�-�"�-Þ�r�"�-�"�-�"�-�"�-�"�-�J�-�R-�R-�"�-Þ�rú�-Þ�r��-��-Þ�r���r�zS-���r�"�-�*�-�6�-���r�RS-���sÞ�rÞ�rÞ�rÊ�-Ò�-Þ�r�6;-��w-��w-�F;-���-���-���-���-Â�-Ê�-Ò�-Ú�-Þ�rÞ�rÞ�rúR-�n�-Þ�r�"�-�6;-�F;-��f-��@-�R;-��w-Þ�rÞ�rÞ�rÞ�rÞ�rÞ�rÂ�-���-���-���-���-���-���-Þ�rÞ�rÞ�o��z8��r���r���-Þ�rÞ�r���o��r8��r���r�"�-�>�-��-��-��-�b�-�n�-�z�-Â�-���-�&�-�2�-�>�-���-���-���-Þ�ß�mÞ�rÞ�oc�P-Þ�rÞ�rÞ�r���r���8��mÞ�r���ocS-Þ�rÞ�rÞ�r���r���8��mÞ�r���oc6S-Þ�rÞ�rÞ�r���r���8��mÞ�r���oc>S-Þ�rÞ�rÞ�r���r���-ß�mÞ�r���o[2S-Þ�rÞ�rÞ�r���r���ß�mÞ�r���oc�P-Þ�rÞ�rÞ�r���r���	8��mÞ�r���oc~S-Þ�rÞ�rÞ�r���b3��!ß�mÞ�r���oc�P-Þ�rÞ�rÞ�r���r���8��mÞ�r���oc�P-Þ�rÞ�rÞ�r���r���=8��mÞ�r���oc�P-Þ�rÞ�rÞ�r���rÞ�	ß�mÞ�r���oc�P-Þ�rÞ�rÞ�r���r���8��mÞ�r���oc�P-Þ�rÞ�rÞ�r���r���58��mÞ�r���ocS-Þ�rÞ�rÞ�r���j���ß�m�JS-���ocS-Þ�rÞ�rÞ�r��iÞ�e8��mÞ�r���oc�P-Þ�rÞ�rÞ�r���r���)ß�mÞ�rÞ�o["S-Þ�rÞ�rÞ�r���r���18��mÞ�r���oc�P-Þ�rÞ�rÞ�r���r���	ß�mÞ�r���oc�S-Þ�rÞ�rÞ�r���j��-8��mÞ�r���oc.S-Þ�rÞ�rÞ�r���r���ß�mÞ�r���o[�P-Þ�rÞ�rÞ�r���r���ß�mÞ�r���o[�P-Þ�rÞ�rÞ�r���r���8��mÞ�r���oc:S-Þ�rÞ�rÞ�r���r���=ß�mÞ�r���o[&S-Þ�rÞ�rÞ�r���r���%ß�m�rS-���oc*S-Þ�rÞ�rÞ�r��im���1ß�mÞ�r���o[�P-Þ�rÞ�rÞ�r���r���8��mÞ�r���ocS-Þ�rÞ�rÞ�r������9ß�mÚ�-���oc*R-Þ�rÞ�rÞ�r����fg����a8��mÞ�r���oc�S-Þ�rÞ�rÞ�r���b;��r���ß�mÞ�r���oc�S-Þ�rÞ�rÞ�r���j;��r���r��-���rÞ�oÞ�r���sß�nß�r���ê�r����ß�mÞ�r���ocfS-Þ�rÞ�rÞ�r���j��2���5ß�m�Ω-���ocZR-Þ�rÞ�rÞ�r����fg�f�rò�-ß�rß�rß�rß�rò�-ß�r�2�-ß�r��-Ê����98��mÞ�r���oczR-Þ�rÞ�rÞ�r���h��b;��rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�r���r�J�2���r���Þ�rÞ�Þ�r���rÞ�rÞ�r���rÞ�rÞ�r���r�֩-���rÞ�oÞ�r���sß�nß�r���rÞ�oÞ�r���ê�r�� m<��r���2���r���Þ�rÞ�Þ�r���rÞ�rÞ�r���rÞ�rÞ�r���rÞ�r��2���r���Þ�rÞ�Þ�r���rÞ�rÞ�r���rÞ�rÞ�rÞ�r��2ß�rÞ�r���rÞ�r���-Þ�r�S-��P-��P-Þ�rÞ�rÞ�r��r���rÞ�r�"�2ß�rÞ�rÞ�rÞ�r�VS-Þ�r��P-��P-��P-Þ�rÞ�rÞ�r�.�r���r�
l���r�L����rÞ--���n���Þ�rÞ�Þ�r���rÞ�rÞ�r���rÞ�rÞ�r���r����K��7��r���2���n���Þ�rÞ�Þ�r���rÞ�rÞ�r���rÞ�rÞ�rÞ�r�J�2ß�rÞ�r���r���r��S-Þ�r��S-��P-îS-Þ�rÞ�rÞ�r�.�r���r���r�*��K��7��r���2���n���Þ�rÞ�Þ�r���rÞ�rÞ�r���rÞ�rÞ�rÞ�r���2ß�rÞ�r���r���rÂ�-Þ�rî�-��P-��S-Þ�rÞ�rÞ�r��r���r���r����K��7��r���2���n���Þ�rÞ�Þ�r���rÞ�rÞ�r���rÞ�rÞ�r���r����K��7��r���2���n���Þ�rÞ�Þ�r���rÞ�rÞ�r���rÞ�rÞ�r���r�&��K��7��r���2���n���Þ�rÞ�Þ�r���rÞ�rÞ�r���rÞ�rÞ�rß�d9��r���r3��r��2���b���
Þ�rÞ�Þ�r���rÞ�mÞ�r�
�o���rÞ�rÞ�r�
�ra�n�r
rM�Þ--���j���Þ�rÞ�Þ�r���rÞ�rÞ�r���rÞ�rÞ�r�
�r5'�nÒ�GV��FǯUEM�W�--���n���Þ�rÞ�Þ�r���rÞ�rÞ�r���rÞ�rÞ�rÕ�rÞ a��r4��f���3��r�J�2���j���Þ�rÞ�Þ�r���rÞ�rÞ�r���rÞ�rÞ�r��r��&�nÆ�j�o�r���J:�����m��2���r���Þ�rÞ�Þ�r���rÞ�rÞ�r���rÞ�rÞ�rÝ�f�r�r7�xe���v�r�r7��lÞ섪��f�����Z�2���r���Þ�rÞ�Þ�r���rÞ�rÞ�r���rÞ�rÞ�r���r�&�y?��r���rÞFxƟ�r�r���r?��r���2���n���Þ�rÞ�Þ�r���rÞ�rÞ�r���rÞ�rÞ�r��rC��C��C��y�r���"��nÞ�Þ�rÊ�2���r���Þ�rÞ�Þ�r���rÞ�rÞ�r���rÞ�rÞ�rÒ��E�oa�rV�x�r���rϟ����rÊ�2���f���
Þ�rÞ�Þ�r���rÞ�mÞ�r��l���rÞ�rÞ�rÞ�r>+�r���&�����������	Ϟ�:;��a���rÞ�r��2������Þ�rÞ�Þ�r���rÞ�rÞ�r���rÞ�rÞ�r�
�rΞ�rñ��
�rט�rÞ�r�!@�O���
�r�r+�--���j���Þ�rÞ�Þ�r���rÞ�rÞ�r���rÞ�rÞ�r�
�r|�&%� ����r?��lÞ��K��y�rR�Þ--���j���
Þ�rÞ�Þ�r���rÞ�mÞ�r��l���rÞ�rÞ�r�
�r|�&!�Ç���'l;��lÞ��K��y�rR�Þ--���j���
Þ�rÞ�Þ�r���rÞ�mÞ�r��l���rÞ�rÞ�r�r�r'�2����O���O���r�r�2����O���O�����rÊ�2���j���Þ�rÞ�Þ�r���rÞ�rÞ�r���rÞ�rÞ�r��rC��C��C��y<��r��oaÕ�rÞ�����r5��r���r/��2���r���Þ�rÞ�Þ�r���rÞ�rÞ�r���rÞ�rÞ�r�r�rÞ2����S���S���r�r#�2����S���S������E��rÊ�2���f���Þ�rÞ�Þ�r���rÞ�rÞ�r���rÞ�rÞ�r�
�r|�&��lÞ�nO�"���,g.��rO:�x=��rR�Ξ�r�r.�--������
Þ�rÞ�Þ�r���rÞ�mÞ�r��l���rÞ�rÞ�r�
�r���b��r������r/��j���n_��m����W���;��r��ve���Ê�2������Þ�rÞ�Þ�r���rÞ�rÞ�r���rÞ�rÞ�r��mW��dŞ�r�mW��dŞ�r�mW��dŞ�r�mW��dŞ�r��rÞ--���r���Þ�rÞ�Þ�r���rÞ�rÞ�r���rÞ�rÞ�r�
�r|�&�����xe��mk��p���mÕ�rÞ���mÞ��K��rÞ--������
Þ�rÞ�Þ�r���rÞ�mÞ�r��l���rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rò�-Þ�r�J�-��-Þ�rî�-Þ�r�&�-ÞR-��R-�R�-�>�-Ú�-���-�B�-�j�-Þ�r���-Þ�rÞ�r��-Þ�rÞ�rÓ�m�퓯E��`����7�xe���;��r�-a��n�r��S�]x>��r�9r4��n���r�Z�2���b���Þ�rÞ�Þ�r���rÞ�rÞ�r���rÞ�mÞ�r��k�
�r|��3�)��+�rW��O��)���nO�"���,g+��r���r�r.��rÞ���|�<�--������Þ�rÞ�Þ�r���rÞ�lÞ�r��l��l���rÞ�rÞ�r��r� �r�<�r;���� ��y�r#�xa����<��rR�1W�7��rC��7��rΞ�r�y�r3��rÊ�2���j�"�Þ�rÞ�Þ�r���rÞ�rÞ�r���rÞ�rÞ�r�
�r|��3�)��+�r?�p��,iS���;��|�6�r�v�m=��lÞ��K��y�rR�Þ--������Þ�rÞ�Þ�r���rÞ�lÞ�r��l��l���rÞ�rÞ�r��r���r��r���r�L�Þ쬑H����rÞlaÕ�rÞBx2��r�L�mÞ�'$��K��Þ�R��Z�2���n�&�Þ�rÞ�Þ�r���rÞ�rÞ�r���rÞ�rÞ�r��rΟ�rÕ�rÞ2�����W���W�����rÞ ��<l;���� ��rV�x�r��+mϞ����rR�Þ--���b�*�Þ�rÞ�Þ�r���rÞ�rÞ�r���rÞ�rÞ�r��rϞ�x���raT�f��s
�sM��x��rR������
�s4��f�� ���r?��n������r�|;r����--�����*�Þ�rÞ�Þ�r���rÞ�rÞ�r���rÞ�rÞ�r�
�rΞ�rñ����r�&��+� Õ�rÞ���j�h#mR���� 	�
�r;���� �
�rW���3� a���r�����2���r�.�Þ�rÞ�rÞ�r���rÞ�rÞ�r���rÞ�rÞ�r�
�rΞ�rñ����r�&��+� Õ�rÞ���j�h#mR���#� �
�rW���'� Õ�rÞ�mÞ�j;�f1���r�����2���r�2�Þ�rÞ�rÞ�r���rÞ�rÞ�r���rÞ�rÞ�r�
�r|�&��mÞ�}�����m7������v��8c�����xe�r�v(l�lÞ��K��y�rR�Þ--����&�Þ�rÞ�Þ�r���rÞ�lÞ�r��l��n���rÞ�mÞ�r�>�o��r��l������r6�r��r:��aK��r"�2�Q�e;�f5Êi�O\pW�Q�e;�f9Êi�O\:;��a���r,�2���:�2�Þ�rÞ�Þ�r���rÞ�rÞ�r���rÞ�rÞ�r�
�r|��3�)��
�r|
�&� ��
r�rV��W��[��v�����x=��rR�Ξ�r�r.�--����"�Þ�rÞ�Þ�r���rÞ�oÞ�r�
�l��l��l���rÞ�lÞ�r��l��lÞ��7�)��
�r|��/�)����'���W����W��������.mÞ ���-m7��n�
�������2����"�Þ�rÞ�Þ�r���rÞ�oÞ�r��l��l��l���rÞ�lÞ�r�
�l��lÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�r�N�-ò�-�ެ-�f�-�J�-Ò�-�b�-�*�-�گ-�
�-Ö�-���-ö�-�®-Þ�rÞ�rÞ��7�)����r>+�r�����
r���c#�����r1���� r]:�iÞ���?�rV������s��n��2����&�Þ�rÞ�Þ�r���rÞ�lÞ�r��l��l���rÞ�oÞ�r��n�
�n�:�o��rϞ�x���raT�f�#r
#rM.�ik�����r>��s��x���6?6�ic�����r4��b�
?r4��n���z��m?������rÞ--����6�
Þ�rÞ�Þ�r���rÞ�mÞ�r��l���rÞ�rÞ�r�
�r|�x=��rW�d��mÞ�p����rΞ�z�������rq>�e�<r4��f��<rb�r	.�p� ��#r.�--����.�Þ�rÞ�Þ�r���rÞ�lÞ�r��l��l���rÞ�mÞ�r�.�oÞ�r>+�r���k�hmΆ�r�PlaÛ�K��/���K��d@��b'��r������r"��o*�eO��2���jS��y��rÞ�n������<�2���f�:�Þ�rÞ�Þ�r���rÞ�rÞ�r���rÞ�oÞ�r��l��n��n��rƚr���j>�iO��o�iO��
�ra��f�rB��~=*����r�ᐦ�;ri� ��
r�t���r�T���;r��r�Z�2���
�6�Þ�rÞ�Þ�r���rÞ�mÞ�r��h�r���r���rÞ�mÞ�r��oÕ�rÞ aÕ�rÞ��������6Ϟ�����p_6�4�r��r��r?����7r��s�Z�2������"Þ�rÞ�Þ�r���r���mÞ�r�>�h���rÞ�rÞ�r������rÞ�rÞ�r���rÞ�r���s���rÞ�rÞ�rÞ��3�)��
�r|�m>+�r���j��gI��r6�;� mW�fN��r:��[�-���r'h�d���r����:�����q���r�*�2����2�Þ�rÞ�Þ�r���rÞ�oÞ�r�
�o��l��l���rÞ�oÞ�r�>�l�:�l�6�lÞ��7�)����'���$8�����m?������rÞ*��� ���4r��������=o�{e�
�0o�����m;������rS�3rj�;r�r�*�2���
�:�Þ�rÞ�Þ�r���rÞ�lÞ�r��l��l���rÞ�nÞ�r��l�:�l�6�l�2�l��$m���nO���O��mÞ�y�ra�f�r
r&�h���W�;��r�x�r���r�<�r;���� ����rÞ�f��mS�V�xeÞ�d3��r���E��r--���f��Þ�rÞ�Þ�r���rÞ�rÞ�r���rÞ�mÞ�r��l�
�r|�
w��l���KM�8w���
rޒ�sa���S���<��r?*�g?��r?*��
�8w�����lÞ�nW��mÞ�vH
rޝ�nW��i���=K���<��2�����Þ�rÞ�Þ�r���rÞ�oÞ�r��l��l�
�l���rÞ�mÞ�r�*�o���r���y�r��$m;�����mÞ�'��j;�f5���r���d>��r��r���d7��r��r���d7��r��rÞ�j�o�rΞ�r���r���y�r;�����mÞ�j;�}-���r���2���r��Þ�rÞ�Þ�r���rÞ�rÞ�r���rÞ�rÞ�rÞ��'�)��
�r|�m>+�r���k�hmΆ�r�PlaÛ�S��/���S��?��7��c#����� r1����r�~%mÞ�r�����m5�r3��?Þ���2�����Þ�rÞ�Þ�r���rÞ�lÞ�r��l��l���rÞ�oÞ�r��l�
�n��nÞ�r>+�r�������r?����� x�rΞ�r��r�l�rÞ�rC��l�-?r?ސ�c��r?>�<�)���r'��/[������r7����8�n��������2�����Þ�rÞ�Þ�r���rÞ�rÞ�r���rÞ�nÞ�r��l��l�
�o�>�h�r���rÞ�r>+�r���mÞ�nK�{e��~=��s^��Þ��K�{e��-���y�r��m�� ��r�r_�/�+��b���6�� ��r�r_����!��-r?�����g��l�����r"��r/�--�����Þ�rÞ�Þ�r���rÞ�rÞ�r���rÞ�mÞ�r�:�kß�q���O����
�rW��jO������M����
�r;���{���7��j�h#m���(��r>�o��r!�y"��mΟ�rÕ�rß�mÞ�y�r;���������r<� �����������r���2���f��Þ�rÞ�Þ�r���rÞ�lÞ�r��n��n���rÞ�rÞ�r��r�r4��r�rɟ�r�
rΞ�x�rj�x�ra���r
rM��[��mÞ�'�d��r5��r�rP���S���O\~�ま�rV�x�r��mΞ�r�r ����r!��Þ--����b�Þ�rÞ�Þ�r���rÞ�rÞ�r���rÞ�rÞ�r�
�r|��3�)��+
mW�.W����-3r:��&���r;��&�� rq��e��s4��j���s���n�*���?mW
���=W���
r4%�jÕ�rÞ���mÞ��K��rÞ--������Þ�rÞ�Þ�r���rÞ�oÞ�r��l�
�l��l���rÞ�oÞ�r�*�o���o���o��0r`��n��pɞ�rÕ�rÞ ���rÞ2l����'���'��
�pɞ�rê�5����<�r?����rÞ�5��+��oÞ���rR��1W���#����rÞ�M��n��j���r��n_��j���r���J�2�����j�Þ�rÞ�Þ�r���rÞ�rÞ�r���rÞ�rÞ�r�
�ra��n�r
r���r�P���<r ���,r4��f��,rb�r��"����K�����S���
�rW�g��r��rÞ�-Þ�nK�"���,is�����ns��s�����=K��6��<r.�--���2��
Þ�rÞ�Þ�r���rÞ�mÞ�r��l���rÞ�oÞ�r���l�.�o���oÞ�r>+�r���k�h3mΆ�r�PlaÛ�K��/���K������r��r4��j��/m?�p��f}��ry.�?>��7��c#�����r1����r�~(mÞ�r�?�rb��n��������2���6��Þ�rÞ�Þ�r���rÞ�rÞ�r���rÞ�iÞ�r��l��n�>�n��o�.�o�� m<��mÞ��=��rR�1W�e;�}1���r���y�r��dm?�e;��>�
�rW��j;�f1���r<����m;�����j�h�ra��j�r
r:�����rR����j�h�r5��n�ڛmÞ�j;�}1ß����r���2���f�n�Þ�rÞ�Þ�r���rÞ�rÞ�r���rÞ�rÞ�r�<lÞ��ڛoÞ�y�rW�x�r> ��\��rR�1W��_���rÞ�v��iÞ��]������r7��l��mS�I�y�r�	lΞ�rç�P��mS�I��^�B��rR����mS��^�����rÞ--���f�n�Þ�rÞ�Þ�r���rÞ�rÞ�r���rÞ�rÞ�rÞ��3�)��
�r|�m>+�r�����
r>�9W��7��e���6W�iO����m��rÞ�Õ�rÞ�mÞ��S����� ��
r`���r
r>�qj
rM
�_��gW�g4��r���W�����Þ--����f�Þ�rÞ�Þ�r���rÞ�lÞ�r��l��l���rÞ�mÞ�r��l���r9"��O��Þ�O��rW��O��rW��O��r��t����~*vr0��mÞ�O��r?���rW�O��r�yr.��mÞ��O��mÞ�y�r;��h��mÞ�j;��.�
�ra���r
r����+��mÞ�S�r��l���2���f�v�Þ�rÞ�Þ�r���rÞ�rÞ�r���rÞ�rÞ�rÕ�rÞxa���y=��r��r�l�r2��rC�xa���7��rΞ�r�
r�-5��f�������r�:�;��r5��jÕ�rÞ�-Þ�nO�"���iw��?���nw�<W��&�
r���r�r�rÞ�>���Ê�2����b�>Þ�rÞ�Þ�r���rÞ�lÞ�r��h�rÞ�����r���rÞ�lÞ�r��k�*�o��sM:�x���r�:�mÕomÞ�����k������+C������rÞ���s>�����<�m?�������s"��ƃ���]��������rÞ--����>��Þ�rÞ�Þ�r�"�rÞ�lÞ�r3��$��s�n;-Þ�rÞ�rÞ�rÞ�r��$#��s�n;-Þ�rÞ�rÞ�r�"�l���rÞ�mÞ�r�6�l��r9���������n[�oa�
r`(�f�r
rM��O��mÞ�'q�y���r49�n��rV�ig���g���< l;���� ���r�6��r:��O���'q�y=��rW�d��mÞ�p���rÞB�S�����=K��rÞ--����r�Þ�rÞ�Þ�r���rÞ�lÞ�r��l��l���rÞ�mÞ�r�:�lÞ��7�)����'����Ξ�rÕ�rß�lÞ����
r7�����sɞ�rÕ�rß�"��� ��2���s>�i�����n��{^��n�>���,r�������%�ᐦ�	?r�r�L/r=�<K��2���Þ--�����f�Þ�rÞ�Þ�r���rÞ�oÞ�r��l��l��o���rÞ�nÞ�r�>�l���l���o���o�
�r|��3�)��
�r|
�&A�����m��ak��mW�q'�����4r
7rV
�ig���g����r
r''�n_���_����$l+���c�����7�g�����7?;�rb�3rj��lÞ��K��y�rR�Þ--����f�Þ�rÞ�Þ�r���rÞ�oÞ�r��l�
�l��l���rÞ�nÞ�r��l�>�l�:�l�6�lÞ�r>+�r����#r������xe��s:��,#r>*�i'��T���n'��/ǜ�m�9ǖr��&������m1
r>�sN���Þ�jS�4!�D�4g�Dlf��9w���Þ�~�r������u�6�r���rÞ--�����f�>Þ�rÞ�rÞ�r���rÞ�nÞ�rÖ�n�
�l��n��n���rÞ�nÞ�r�*�o���o���oÚ�oÞ��7�)����'���Ϟ���
r����¡m0��O�����,m������0mܞ�n�������3����
r����¡m0��O�����,m������mܞ�n������~��rV�q'�m��c3�����r1����r1:�O���rO�r�rÞ--���f�~�
Þ�rÞ�Þ�r���rÞ�mÞ�r��l���rÞ�lÞ�r��n��nÕ�nÞ�����r;����>����rΞ�p>�ig���g�I����k���O�!�O����� ��
7r4��f�� ���r�6�h�>���2�x=��rW�d��mÞ�p���rÞBpU�x=��r?� ��2?��g��r?����;?�r��rÞ--�����v�Þ�rÞ�Þ�r���rÞ�lÞ�r��l��l���rÞ�iÞ�r�>�l�:�l�2�l��o���oÕ;mÞwÞ�y�r���nÕ�rÞw���y�r���Õ�rÞw���/��r���f�r�r?�w���y�r8���r�r3�la�<�r3���� ��r'��/W�����r4��j�� r���Õ)Þ2o����S���S�v���3��ra��n�r
r������rÊ�2���b�N�Þ�rÞ�Þ�r���rÞ�rÞ�r���rÞ�mÞ�r�
�l�<MlÞ=�� =�r>�x��rW�g���r� r'~�n���������s
�s4A�f���n������rÞ����rÞ�mÞ�no��k���r���nW��mÞ�no��k���r9��:;��iÞ�y6��rW��9�s>��x>��r���r�
?r�H�"���KV�g���r��rÞ--�����N�Þ�rÞ�Þ�r���rÞ�rÞ�r���rÞ�lÞ�r���l���lÞ�r>+�r�i�nÞ�nW��2���n_�la���<�r:�`��r;��o��r���$!�nW����>%)���9���=��.m;�*���
��r"��o*��e��2���j��|��r����r[�r��s����
�)��������2�����r�Þ�rÞ�Þ�r���rÞ�rÞ�r���rÞ�dÞ�r���l��n��n���n���n�
�o�2�o�"�o���o���oÞ��3�)��
�r|�m>+�r�����
r>6�9W6��7��f���6W6�iO���6�m5��rÞ����nc�����rɞ�r�
r>6�9W6��g�`����o���k�����7�o����4r�� ����rÞ����`W�x>��r��qm�� ��r���l�� ����r?��r���rÞ--���
�N�Þ�rÞ�Þ�r���rÞ�lÞ�r��l��l���rÞ�mÞ�r�6�lÒ��E��m?��nc�����nc�<S�����rΞ�rêoa�<�r?�lê�	��c�����KM�8c�oa�
rޒ�sa���O��iS��mÞ�vI
rޝ�y<��r?� s��2?>�g/��r?>�7��rf�/8c������lÞ��S��Õ�rÞ�pɞ�rç����rR�Þ--���&�N�
Þ�rÞ�rÞ�r���rÞ�mÞ�r��l���rÞ�lÞ�r�>�o���oÞ�r>+�r�i�iÞ�nW��2���n_�la���<�r:�`��r;��o��r���$!�nW����>%)���9���=��.m;�*���
��r"��o*��e��2���j��|��r����r[�r��s����
�)��������2�����r�Þ�rÞ�Þ�r���rÞ�rÞ�r���rÞ�dÞ�r���l��n��n���n���n�
�o�2�o�"�o���o���oÞ��7�)��
�r|�m>+�r���r���r���rC<�r7���_��fP�y���i!|�r��rÞ�lÞ�4��rq��i����-;r9��n���=W��>����S�?>��h�
r��s'�����O����oÞl�;��rR�?9��s��s���r5��rß�����--�����J�Þ�rÞ�Þ�r���rÞ�oÞ�r��l��l�
�l���rÞ�nÞ�r���l���l���l���oÒ�KM�x�r���r�<Wm;�!�� !�r���r�?r>.��O������u���u���r&���g�aç��
7rɞ�rÕ�n �2�����w���w���
rɞ�rê���r'o��S������w���w����OmW��|��rR*�1W*��K�����r?��ns����Pm;�'��'�r ���O��b���6/�--���>ê�Þ�rÞ�Þ�r���rÞ�rÞ�r���rÞ�rÞ�rÞ�r>+�r���mÞ�n[��Ò�v������r0
rH3�-�����h�u�r�����r ��&��{��lÞ�'2�r9�zÞ"x�rΞ�r��8r�l�rÞ�rC��j���!��2�o;r����8m|6�ik����#3r>:�gm��r?2������6�m7��rÞwe���rÝzÞ--���:�R�
Þ�rÞ�Þ�r���rÞ�mÞ�r�
�o���rÞ�oÞ�r�:�l�6�l�2�h�'��rÕ+mÞ	��r�;r���r�?r>�i��mÞ�y�r���rÕ�rÞ�mÞ�y�rC��n/���/��mÞ�w���s>��9W���1��rR��1W���7���W���#��h������xß�rV��0��rR��1W���#���<�r?��� ��sV
��3��rR��1W���#����rÞ��E��rÞ--�����^���E]��x;E���4mÞ�rÞ�r���rÞ�oÞ�r���l���l���lÕ,m0����$r
'rB��nw���w��������w�aÚ7������rw�'rV6�x�r��QmΟ�c��r?*�9W*��k� �������w�Ú7����� rV2�x�r��Em?:�x?��rW2����rR"�1W"��s���rV2�g'��r�]mΞ�r�rV6�g'��r��mΞ�r�r.�--���:â�Þ�rÞ�Þ�r���rÞ�rÞ�r���rÞ�lÞ�r�*�l�&�lÕ,m0����$r
'rB��nw���w��������w�aÚ7������rw�'rV6�x�r��QmΟ�c��r?*�9W*��k� �������w�Ú7����� rV2�x�r��Em?:�x<��rW2����rR"�1W"��s���rV2�g'��r�]mΞ�r�rV6�g'��r��mΞ�r�r.�--���:â�Þ�rÞ�Þ�r���rÞ�rÞ�r���rÞ�lÞ�r�*�l�&�l�
�r|�x�rΟ�rÕ�rÞ�	���rW�f��r��x�rΟ�r��8r�")��(r ��_��>���r/��>���j#9�s>
�r<��r_��s��.���x�r?��W��lǫ�lÞ���s�� ��
rV
��r'���_�����s�� ��#r.�--�����F�6Þ�rÞ�Þ�r���rÞ�nÞ�r��l��l�
�h�r�������r���rÞ�nÞ�r��l���l�"�o���oÞ�s��'���a?6�g�r6�m8��rÞ����r��>mv&�e�9m;�-���y�r?�i�����r0����6��$m�7���6��=�{�r��sV�I9����<��s:��`��r;��s�$�rÞ�?��s��d?���	m����4�r�z�s9����b�����nǦ�r���r3��r��2���"â�
Þ�rÞ�Þ�r���rÞ�mÞ�r�
�o���rÞ�oÞ�r���n���n�6�o���rÞ�2�����*�� %��r?*�9W*��(��rR"�1W*��7���W"��k��n�*�%�
7rɞ�rê�Õ�l0�l�� r
#rV6����rR"�1W*��3���W"��o��&�
;rɞ�rê���0r���r�
;r`��f�+r
+rM.��s���
;r4��n���Õ�rÞ��
7r4��n���Õ�rÞ���mÞ--���:ê�Þ�rÞ�Þ�r���rÞ�rÞ�r���rÞ�lÞ�r�*�l�&�l���rÞ�2�����*�� %��r?*�9W*��(��rR"�1W*��7���W"��k��n�*�%�
7rɞ�rê�Õ�l0�l�� r
#rV6����rR"�1W*��3���W"��o��&�
;rɞ�rê�Õ�rÞ�mÞ��o�>����������
?rM��o�����6!T�y�rR��k�����6!��y�rR���--���:ê�Þ�rÞ�Þ�r���rÞ�rÞ�r���rÞ�lÞ�r�*�l�&�lÞ��7�)��
�r|�m>+�r�ɛmÞ�nS������<� r:
�`{��rT�J$
�s^>�Þ�K�3�����
r�4rH��2��/��s.�*����{�Û�����=Þ��S��s��g ��r����6���.�!�&�)���1���nS�����r���y��2���2�J�Þ�rÞ�Þ�r���rÞ�lÞ�r��l��l���rÞ�dÞ�r�:�l�6�l�2�l�.�l�*�l�&�l�"�l���l���l�
�nÞ�r>+�r�������r<�r:�`S��rW�6��=�K��ÞbiS������r��a+��r;�`���r?
�h-����lm4�����r9��0�����j[��"���nc�����r6f�g���s�,rr����Q>�y<�U��?rr����Q
�y<�U���r��a���r�����m/��v<�r:�`?��r%�m���r�"�2���&ò�Þ�rÞ�Þ�r���rÞ�rÞ�r���rÞ�oÞ�r��l��n��nÕ�rÞ aÕ�rÞ��������6Ξ�r��r�n�q6���o��lÞ�nc���Ě�"���&���r�$r���r��r�n�q"�������nÞ�nc���Ě�:�������rk�;rr�#rz�+r��s
��rÞ--���.�j��Þ�rÞ�Þ�r���r���lÞ�r��l�>�hÞ�rÞ�rÞ�r������rÞ�rÞ�r���rÞ�r���r���rÞ�eÞ�r�6�l�2�l�.�l�*�l�&�l�"�l���l���l���lÞ�r>+�r������r"��o*�eO��2���jS�����mC>�����rO�r	>�m�<rd��nS�la���<�r:�`��r;�4��������m`��rÞ����,m;��-��rV�+s��B��s��,���('��nS�la���<�r:�`��r;�s�#�r�����n������rc��s&��r,�2����â�
Þ�rÞ�Þ�r���rÞ�mÞ�r��l���rÞ�hÞ�r���l��n��n�>�o���o���oÒ�G>��7�&A�?r_������S���7�#-��,i3��r���n3��s6��m����5����sג�Gǯ��S@�S�@�[��f���r#��s>��s��rC��$��r��yË��˜�m��l�r�
�rv��e��s4��b���s���s7��n��sS>��5��y<���P쾔r�r��;?��s2����	�sK���r���G���=K��r���2����ú�
Þ�rÞ�Þ�r���rÞ�mÞ�r��l���rÞ�oÞ�r���l���o���o�
�rΞ�rç��Õ�rÞ ��r4��f�� ����rÞ��W��lÞ���<m?�io������no��sr������s������mΞ�rÕ�rÞ�*��}lÞ�b��k;��rv��n�|%���n7�#��,q�&�l���rv��n�|%����/�#e��,q�&�n��$r'7�/w��&��?m|.�is������?��*�8i�r��"�*���--����ò�Þ�rÞ�Þ�r���rÞ�rÞ�r���rÞ�nÞ�r�.�l�*�l�2�o�&�h���r���r��r���>��r�ᐦ���r�Hve����3���
r�
r֘�'����Y��ꁆ�rɞ�r�
r>
�s���������r�ᐦ���r�H�mÞ��7����������rÞ ���r<Rm3��������rV>��O��mÞ��S��lÞ�W��p��������
rɞ�r�
r�-Ξ�r��r�-5��f������rV��K��rÞ--���ö�Þ�rÞ�Þ�r���rÞ�mÞ�r�
�h�rÞ�r���rÞ�lÞ�r��k��k�
�r|��3�)��
�r|
�&�� ����~¤���rq6�e��m?��Õ�rÞ���
r���s^.����s7��nÇ!���sV��w��yÜ2=
#r�<�m?�e���s4��nÓ�m�S�K��*l?�*�
�s>��g#��rW*�I>��xß�r��h�������w��p�rX.�)��rq6�e��m?��lÞ��K��y�rR�Þ--����ò�Þ�rÞ�Þ�r���rÞ�oÞ�r�
�l��l��l���rÞ�oÞ�r���o���o���oÕ�rÞ�jÞ�n_����r3�le��;r=��rΞ�r�
rl��)���rÕ�rÞ ��0���rÞ�oÞ��_�9s���Þ�y?��rW�����s>��r���r�
rl��i���rÕ�rÞ ��0�Ϝ�rÞ�kÞ��_�9s���-Þ�y;��rW��?�i��)���n_�1i{Z��Þ��7�2+���qU2�?�s���lÚ��K��^���rΞ--���ú�
Þ�rÞ�Þ�r���rÞ�mÞ�r��o���rÞ�lÞ�rò�o��h�l���r�
�r|�x�r?:�g$��rΞ�rÕomÞ ���0m$#r>:�v���i�����n�����
�� r���j�*��������rÞ���
r�ᐦΞ�r�
r��-�����<.l/�����
�s�����
r���r�L��w������;�mΞ�rç�u2��6��m3��6����K��j�����*�1���rÞ--����â�>Þ�rÞ�Þ�r���rÞ�lÞ�r��l�
�h�rÞ�r���rÞ�hÞ�r���k�:�o�*�o���o���o���h�rÞ�r�+�m��r�
r>>�9W>�x^��rW�i[���[��m4���1r
r>�qj
rV�*Þ ���0r�6��
r{���e���O��j����>���
r�0��
r��[�����=_���
r{���_��P�����
r>��c�����=g���
r{���g��=K��d����>���:����5�#r.��r|�3�--���
ê�6Þ�rÞ�Þ�r���r���oÞ�r��l��i���rB������r��s���rÞ�iÞ�r��l��l�>�l�:�l�2�l��r�ᐦ���r�Hve����7��lǫ�lÞ�R��S���S��wG�B*�k2�K�a�K��S��mÞ��S�����}l���m���3���7��lǫ�lÞ�Ξ�r��r�-?�x�rW
�[�/Ӂ��rR>�1� _���rɞ�r�
r���r�LaÜ|l���m���S��mÞ��W����ޛmÞ��7���������6� _����8oaÒ�v���rÞF�;��rW��K��rÞ--���Ò�Þ�rÞ�Þ�r���rÞ�mÞ�r�
�h�rÞ�r���rÞ�lÞ�r��k��k��$m�x�q���ig��%���ng�'Ý�!�=����
'��	���������3�xe���y�r��%m�u�rΞ�rÕ�rÞ�j��}lÞ�b��
w��rΞ�r�
�sl�!m�	�s���r�
�sl��s>��hw��!���rq�����mp� ��u���rÞ e�0�J���y?��rW���?��s�)a���s'1�/3��b�<9m7�I���sd
�s���n���r3��s$��p���v>�--���Ê�
Þ�rÞ�Þ�r���rÞ�mÞ�r�
�o���rÞ�kÞ�r���l���l���n�:�o���o���o���h��%���rÞ�r>+�r������r"��o*�eK��2���jO��y��rÞ�n������������r"��o*�eK��2���jO�����r�5�j���n�����r&	�r<���?��7��c#�����r1����r]�iÞ��y��?:��7��c#�����r1����0r]*�lÞ�v����.��r"��o*&�e{��2���j����r=��f����>���&�)���r_�#r��r,�2����Î�Þ�rÞ�Þ�r���rÞ�rÞ�r���rÞ�eÞ�r��n��n�>�n�:�n�&�n�"�n��o�*�o���oÞ�r>+�r������r"��o*�eK��2���jO��y��rÞ�n������������r"��o*�eK��2���jO�����r�5�j���n�����r&	�r<���?��7��c#�����r1����r]�iÞ��y��?:��7��c#�����r1����0r]*�lÞ�v����.��r"��o*&�e{��2���j����r=��f����>���&�)���r_�#r��r,�2����Î�Þ�rÞ�Þ�r���rÞ�rÞ�r���rÞ�eÞ�r��n��n�>�n�:�n�&�n�"�n��o�*�o���oÞ�r>+�r��ye�^�'G�r0r�r3���Û�j��:$a�;��m$r��r����������r$'r?�rϞ�����r�;?�rz��l��xe���_��0'@�r�im���V��*����h�r�r���K��h��*%��eÒ�p�`�l��r����&�m=��m���c���b��m���P�B�xeþ�y�8��Ýxe?�rϞ�����r�m=���;��r$�w��m�����r�r��([��k;��m�s�2`��~w����9[��l���r/*�2���.���Þ�rÞ�Þ�r���rÞ�rÞ�r���rÞ�oÞ�r��l��o�&�oÞ��'�)��
�r|�m>+�r������r"��o*�eS��2���jW��y��rÞ�n������������r"��o*�eS��2���jW�����r�5�j���n�����0r&�r<���?
��7��c#�����r1���� r]:�iÞ��y��?2��7��c#�����4r1����8r]"�lÞ�v�a���6��r"��o*��e��2���j����r=��f����6�����1���rg�+r��r,�2����Ú�Þ�rÞ�Þ�r���rÞ�lÞ�r��l��l���rÞ�eÞ�r��n�
�n�6�n�2�n���n���n�:�o�"�o���oÞ��7�)����'���"�f,��r�r	"�m6
r`��n�r���mÞ��[��lÞ�?�s�������Þ��O�����r�=�m�� ����������_��p��~5�.r>��(��rR
�m0�rq2�e��m?��"�f,��r�r	"�m0
rV�IΟ��#��bW�I>�x>��r��aW�I>�r*��r;
rޝ�r9�rd��y�r?� o��24��j���s'�w��s&��r5��rß�����W�������--���2���>Þ�rÞ�Þ�r���rÞ�lÞ�r��h�rÞ���������rÞ�lÞ�r���l�"�oÞ��'�)��
�r|�m>+�r������r"��o*�eS��2���jW��y��rÞ�n������������r"��o*�eS��2���jW�����r�5�j���n�����0r&�r<���?
��7��c#�����r1���� r]:�iÞ��y��?2��7��c#�����4r1����8r]"�lÞ�v�a���6��r"��o*��e��2���j����r=��f����6�����1���rg�+r��r,�2����Ú�Þ�rÞ�Þ�r���rÞ�lÞ�r��l��l���rÞ�eÞ�r��n�
�n�6�n�2�n���n���n�:�o�"�o���oÞ��'�)��
�r|�m>+�r������r"��o*�eS��2���jW��y��rÞ�n������������r"��o*�eS��2���jW�����r�5�j���n�����0r&�r<���?
��7��c#�����r1���� r]:�iÞ��y��?2��7��c#�����4r1����8r]"�lÞ�v�a���6��r"��o*��e��2���j����r=��f����6�����1���rg�+r��r,�2����Ú�Þ�rÞ�Þ�r���rÞ�lÞ�r��l��l���rÞ�eÞ�r��n�
�n�6�n�2�n���n���n�:�o�"�o���oÕ�rÞ�bÞ�Ћ��rRړ1Wړ�����{��*���v#�n/�)�<l;�1�����$p"���-ƕ�rÞ��
/pɞ�rê���rW.��'h�nW��n���v7��n���vV�iW�$i���v�3���O��lÞ�R�i{��N��l?�����������nߘ�*��lWړ���"�
+p4��n���rÞ--���?���Þ�rÞ�Þ�r��rÞ�nÞ�r2�l��$��s��8-Þ�rÞ�rÞ�rÞ�rÂ�$��s��8-Þ�rÞ�rÞ�rÞ�r�&�$#��s��8-Þ�rÞ�rÞ�rÞ�r���rÞ�lÞ�r��l��lÞ�r>+�r��xe���_��0'n�r��rÞ�rß�7[��rq6�ik�{e���n{��1���n{��;;�7)��r���n�6�%���y�r?���K��lǫ���m�����
/rV�$7r?�rϞ�����r6�m5�,rX���Þ�r0r�r/���Û�$��4Ξ�rÕ�rß����� k����r�r/��*���r/��*���j#9+r>�r<��rk�'r���mÞ�n�����v��=���r �imW���K�My6�`��~w����9k��d?�����m���r/*�2���&���Þ�rÞ�Þ�r���rÞ�mÞ�r��h�r���r���rÞ�lÞ�r�6�o�&�oÕ�rÞ�.�<�rÞ1�� 1���rÞBs^��Y��$r`��n��s���r�
�sV"�g��r
r�0��
/rV"�v���s$�s���r���s4��j���sǏ�sɞ�rÕ/mÞ�"�Ąse�� ���?��g��r?��p�^�f
��ryN�v�~�x9��r?n�g��r?n�v�����??��s���b������m�N��n����(rX���
/r�Ê�2���vº��Þ�rÞ�Þ�r���r���oÞ�r�읳n��n���`q���r������rÞ�rÞ�r���r���r���r���l���rÞ�dÞ�r���l�^�l���o���oÞ�oâ�o�N�o�~�o�n�o��o�<�rÞ�� �<�r?�	�� 	�rV�x�r���mW��=��rR��1W���S�����rÞ��a��"m!��n�����n��������
r`��f��s
�sM��[��mÞ�'���[���<�r;��� �r���Õ�rÞ�mÞ�yß�rɟ�rÕ�rÞ�mÞ��S��:����W�����r;��y<��rR�x�ra��n��s
�sɞ�rê����rÞ��[���<�r;��� ���rÞ�)�rR�g:��r
r4��n�� ����r?��s��l���2�������Þ�rÞ�rÞ�r���rÞ�mÞ�r�>�h�rÞ�r���rÞ�rÞ�rÞ��7�)����'���Ξ�rÕ�rß�lÞ����
r7����r�ƛlÞ�nK�"���,io��
���no��.����������fm�� ��(�lÞ��	;r���r��rq�e��s4��b���sb�r������m��rÞ�rß�7_��rq2�io�����s4�����s���j��iO��o	������m$��s��
r�ᐦ�	+r��s0��W��i'��W�Äs'����ۜ�dW��g��r�����mA���r���s��--������.Þ�rÞ�Þ�r���rÞ�hÞ�rÚ�oÊ�o��l���o��h���#�����v���rÞ�oÞ�rÆ�l�2�o���oÞ�r>+�r�������j<�r:�`K��r?�6��g�rP���j<� r:
�`W��r����
�m#�r��m4� ����v<�r:�`G��r%�m#�r��m4� ����n<�r:�`G��r%�m�r��o*�eO������nK��a;��rQ��S�\:"��o*
�eW������?�rV��7?�0��O�����lmÞ�����j����K���O�0��W�����mÞ�n������nS��c������r1�r��r��m4���r���c?����� r1b�r���rO�r�s�"�2���b���Þ�rÞ�Þ�r���rÞ�rÞ�r���rÞ�lÞ�r��n�
�n�
�r|�pΌ�K���(��'3�nS�����y�rW�ik���k�a�<�m/���� ���r�6���9k��!�� ���r���r�rV
�fj��r�ig��lÞ��o�����<r
?rɞ�r�� rV�ik���k���
�ra���#r
7r>�qj
#r���rç�n�6����Vm!��y=��rW�d��mÞ�p���rÞB�_�����=_��F���s>� ��2?� ��2;�`#��m	��f����[��lÞ�R�l� ���9� ����r?��Þ--�������Þ�rÞ�Þ�r���rÞ�oÞ�r��n��l��l���rÞ�nÞ�r�6�l�.�l���oÊ�oÕ�rÞ��rÞ���
l�r�iÞ��]���rÞF�>	�d��r��rÞ��l���r�HAhU�����6���r�	lI�y6��r�H�����r7��y>��rI ��[�Þ섕� l5��f�ڛiÞ��]���rÞF�>�d��r��rÞ��l���r�HAhQ�����65��r�lW�hP�/�'���
r9�-����T� ���lo�rI
��K����!|�lW�hP�/�3���
r9�-���iQ������W����l�~e�� rH�y*��r�l5��r��rX����rÞ--���b�"�Þ�rÞ�Þ�r���rÞ�rÞ�r���rÞ�mÞ�r�
�l��r�o*�eK��Þ��O��mÛ�O������r,�r�o*�eK��Þ��S��
Þ��=��s�g<��r�����K������n<�r:�`���rW�?��(s������r?������-���s8��B"�j�$�sǏ�s��eÛ�M��r�o*��e��Þ�0S�%�������@s5��B���s���c?�����xs1B�r���rO�ws���������rs�r��s�s��Ss���m���v<�r:�`���r%��"�2���J���Þ�rÞ�Þ�r���rÞ�rÞ�r�&�rÞ�cÞ�r��l��l�v�l��nú�n�r�n�>�o�.�o���o���oÞ�oþ�oê�o�Z�o�z�oÕ�rß��� r`��n��pɞ�rÕ�rÞ U���rÞ2l��������M�
�pɞ�rê�(ß�f���nϝm����띚mÞ�y"��rW��x?��ra��b��p
�pM���㝚mÞ�'b�s��n���p`��n��pɞ�rÕ�mÞ U���rÞ2l��������M�
�pɞ�rê�ß�f���n�����r=�]��p:��h��
������_�ם���p2��l��p>��e;��6���r=���NI��pΞ��'���ם��ߝ����p���ם�Ɏ��MN������rÞ�r��A|L���ם�E�r>�e;��>���r?��e;��6���r���r?��r�J�2�����Þ�rÞ�Þ�r���rÞ�rÞ�r���rÞ�rÞ�rÕ�rÞ�?Þ�y8��r���rÒ�v�PAj;��r�l�r2��rC��mÞ�;��r
�-a��n�r
��[�6��<�r?���
rɞ�r�r�r;�����2h����[����
r�y�r7��mÞ�nO�{e���y=��r����E����`W�;��r�~���3r�����퓯e��`���~e��q�8�g1��r�9�`Ơ1r4��nÒ6q1������r?����퓯e��`���~r��q�8�g1��r���rÒ�v��r���rÕ�rß��s��m��`Ơ1r4��n�
r���r�� r��r?�����r[.�b���r?��b������`Ơ1r4��nÓ�m�퓯e��`����S�����r�Z�2�����Þ�rÞ�Þ�r���rÞ�rÞ�r���rÞ�mÞ�r�
�kÞ�r>+�r������r"��o*�eK��2���jO�����r�5�j���rK�r	���o,��nO�la���<�r:�`��r;�s�$�rÞ�?�rN��jN��S��o,�8�g���rC��0��K�����,m����r>��rc�r'��w�����r"��o*:�eg��2���jk�%���r�>�.���r�Ψ??�r~��j����:�����r_�'r&��r<��?��奞�u������r?�����rƛ�sa�%������8?�r������Þ�r�rC��0��K�����,m�����O-Þ�r���rK�r�oc�2�����2�Þ�rÞ�Þ�r���rÞ�rÞ�r���rÞ�eÞ�r�>�l�"�l��n��n�:�n�6�n��o�&�o���oÞ��7�)����'���Ξ�rÕ�rÞ2���������-ƞ�y��rR"�m#�(p>�O��b�
/p4�j���b��(p"�r=�;i[��n���v7��n���vV�i[�$i���vx��iۛ����nۛ���-�v:�����r;��ě�ğ�7��hÖ�EǦ����jW*��K��o/��r�(p>n�O����
/p`�j��q�|w>"�O� 5Ƃ3ƞ����m��8m�� -���r?��r5��rÞ����S�--���F>���Þ�rÞ�Þ�r��rÞ�nÞ�r3�$��s��8-Þ�r�	h�9��rß�r�n�$��s��8-�b�rÞ�r�	h�9��r��l#��s�"�$#��r��8-Þ�r����<��r��rS��rÞ�hÞ�r��l��lÖ�oÆ�oæ�o�V�oÞ�r>+�r���mÞ�ڞ����m7������v��8o��"�G������q����m�>����8r�ٛÞ�no�����y�rΟ�rÕ�rÞ����8r���sV�f��r������4x=��r?� ��2?2�g!��r?2�7��mΞ�rÜ����s?���ß�lÞ�n_�"}��,i�����n�<_��j�2����M����_���Û�۞�j$b�/_��*�r*��mÞ�����r;����>�V��8r�֛h����Z�� U�
r>��9W��gמ�r
�s>�qj
�s>��qj��r��s�� Q���r?������r7
rx"�p�
�mÝzÞ--����:�>Þ�rÞ�Þ�r���rÞ�nÞ�r�
�oú�l��l��n���rÞ�hÞ�r���lö�l�2�o���oÞ�oþ�o�
�r|�i�Q:�����N���Ny�
��Ξ�rç���✽{��a��mW�_�;Q�B�&�r6���
����?�_%7��.�����Ni�✽{��a��mW�_i�N'a���r#� A���rÞ^�R�_x�r��r��rq�_e⠽5��b�⠽�>��?�_i�N�l�_x�rW�_y=��x=��r�␽�o�r2��rC��m�� q���v�
���~�mÞ���Nݮ��2�����N®�
��R�_x>��r?�_i#Q����6?�_%7�������N�✽{��a��mW�_�Q�?����r���a��j���
��R�_��N�mÞ�'7�~�r>�_g
��r��rÞ--���q�>Þ�rÞ�Þ�r���rÞ�lÞ�rÚ_h�rÞ�����r���rÞ�oÞ�râ_kê_oæ_h�rÞ�r�
�r|�pΌ�K���(��'3�nS�����y�rW�i����a�<�m/�=�� 9��r�6=��9��!�� ���r���r�rV
�fj��r�x���rR��i��mÞ�n�/ic��mÞ�nW�����s
�sV��7�2x������������7���n������&�rÞ ���1mΞ�rÜ�x=��r�
r7S�j��rɞ�rÕ/mÞ�2�9�sq��c��s4��b���s���s7��n���s��87�Ķ�ǰs���_������>�
�s$�s:�`#��m��;;��sƜ�s������rÞF�[����
r�0���
r4��n���rÞ--����>��Þ�rÞ�Þ�r�&�r���iÞ�r��n���l��l���hÞ�rÞ�rÞ�r������rÞ�rÞ�r�A�rÞ�r���r��l���rÞ�iÞ�r���l���oÚ�oú�o�Z�oÞ��7�)��
�r|�m>+�r�� ��hm?����
r�r�?r>�iS��l�����m,r�r��]�����km;��zɞ�rÕ/mÞ���-?r->�2��jm3�xe������Û�W��[����*=��,rǏ�s���s7�j�$�s���r���s4��j���sǏ�sɞ�r��s4��j��sǏ�s���r��Ps4��j��PsǏCs���r��ps4��j��psǏcs��Û�������
r������m0��[�����,mJ�����O.Þ�m���rW�r&��n������r�/r"��s6��s朣s��Cs��csV��r/*�2���
�&�:Þ�rÞ�Þ�r���rÞ�oÞ�r��l��l��h������ o<�rÞ�Þ�r�
�l��l���l��n��n���o���o���o���oÚ�oÊ�oú�oê�o�Z�o�J�o�z�o�j�o�
�o��h����rÞ�r>+�r��)��rا� Þ��~��mÞ�y���ra��f�r��rÞ ����r;��r5��rÞ(Þ�y�rD"�r=��~��r�%ml�r��mÞ��7���y�/p���r,��rÞaÇ+�!��?��a?�gx��r�m6'mT��K���m���%�4!m�zr9����b���_��dΞ�r�'m���aI+��7���'��r5��rÞ&Þ��w��mÞ�w��m���m �x�r���r�#ms�#m3��r4��rÞ��w��l��#Ú��7���'��r:��rơ=m��mE/�r=��y�r?:��7���s�/�Þ�lǫ��o�El�� ���r�?mh�ri�r'x�r%
3rW��KH.�-���-k��p�1�rÞ�~�
3rW��KH.�-���-���r=��ng���3�r���r��2���
�J�Þ�rÞ�Þ�r���rÞ�rÞ�r���rÞ�lÞ�r��n��o��r���cÕ�rÞ�1��r
r���rC<�m/���� ����rÞ�S���KmÞ!���rÞ����2������&�
+rɞ�r�9rɞ�r���m?�9W��O�`����{���{��mÞ��[��3�#�s��7���rÞ9�����9���mÞ^��9�����FJ>2�q��A��9��-w�rÞ�2���Eɟ�râ�c��?�I�io���W��x*��r��sW��y=M?��sΞ���7���S��3��rW��x=��r�
�s7��f��rV����S��b���~!�s����������'9����l��s'b����=� 7���S!n���(��
r4��n���rÞ--�������Þ�rÞ�Þ�r�"�r���nÞ�r��l�2�hÞ�rÞ�rÞ�r������rÞ�rÞ�r�B�rÞ�r���r���l���l���rÞ�lÞ�r��l���oÞ��7�)����'������r��rq:�e��r;�������S��mÞ�w�Nl�� ����r�Ω�S��8Û߯��jl�� ��
r�8r>.�9W.����rR*�1W*�IR8�??�8rr��T8�J���râ��'n�r8���u�͛Þ�~�!r������'I�r8���u��jT(�$��cW��F'��v����/�lÒ�v���K�y�rW���3����r?�ll�� ��
r�8rV���3��o��gT�y=I�����/��lÞ�R��r=�hl���cW��F'��v�����/�lÒ�v�����y�rW���3����r?�ll�� ��
r�8rV���3��o��gT�y=I�����/��lÞ�R��r=��r=��y�r��f��r�8��i!��r��M�--���.�F�Þ�rÞ�Þ�r���rÞ�lÞ�r��l��l���rÞ�oÞ�r�2�l�.�l���oÞ�r�� -ß�rÞ�r��-Þ�rÞ�rÞ�rß�rÞ�rú?-�?-�b.Þ�r��?-�bb.�b>-��?-�fb.�b>-�J>-�jb.�b>-â>-�nb.�b>-Î>-�rb.�b>-��>-�vb.�7m�6m�5�\��;�S��r�8�\
�L��r�"�_�r�)�^�r�?�N�Q��+�O�r�,�]m�"
�\�O	��3�_�r�3�M
m�&
�S$�^��r�&
�S#�O��#�\)Z�b�r� �^;�Om�b>-öf-�zb.�b>-Þf-�~b.þw-�Z3-�Bb.� .�))m�
)|��r�
4�_m�
'�Z��+�]��r�
8�\*
�O��rÞ�r�
8�\2��
8�\7�O�r�
8�\&
�Xm�9�S��r�
+�L#�Y�r�
+�L;�S��r�
+�L4�_m�
+�L'�Z�� $�b�r�
=�H&
�Xm�
=�H7�O�rÞ�r>+�r���:���m$�����(k��
��m7��
���v�
�[��h�6�5���m�$r��;��
ۜ�r� r�x7r��r�ҐuN������
�)Y����O���������ro�rk6�P��$r���B
����7�s㞑B������w�J�eS�4����w�j�7;�KmďsbѸs�������Z��z����m4�r��sH��fW�����=��j$��/��&�O���j���J���	;
�s�6�Q���v�����4r�� ���r�sF���;��k��m&�S�5��rk��R�����s➑B�����7ssݞ�B���j�B�w�����;3�4r
��s��Cs��csF��g?�sI����Y�������<�--���n�j�.Þ�rÞ�rÞ�r���rÞ�jÞ�r��lê�n��n��n��nò�lî�l�
�n���rÞ�eÞ�r��l�6�o���o���o�Z�o�J�o�z�o�j�o��oÞ�r>+�r���:Þ�{���-;r:��>���=[��cW�x�r�����[��m������r��rHy�~=��s^*���_���!amÒ�v���rÞF�{��Ξ�r�
'rV����/kÞ��vl7��r���(�iÞ��	�s���r��rq2�e��s4��bÕ�rÞ����s��Bʜ�sΜ�N��m7��N����{���vlh�r�gm�Ϙs��
���u���m{
rt��rÞBpU��x=��r?� o��2?��g��r?������{���vlh�r�~i�Ϙs��
���m �mi��vʾ�i㜒�:� ���+5�� %�
rHy�-���-k��p�z�l�
�s}�q�����ϟ%�
rHy�-���-���r5�rX*��Þ�r.��rÞ�
���r;������s���Þ�q���rÞ--����Z�Þ�rÞ�Þ�r���rÞ�lÞ�r�
�o��l���rÞ�hÞ�rÒ�lþ�n���o���oÖ�oÂ�oÕ,m0�����s
�sB��n'���'�����/���'�Ú7�/����r'��sV��x�r���l���r��r?��9W���� ����/���'�Ú7�/�	���sV��x�r��ZlΞ�rÕ�rÞ����}l���m��n��mÞ�y�rW2�3�/������/��3���sV��x�r�
�sɞ�rç�מ 	���r?��������6�|7r�����s7��r���s:��`w��rW��xD��r���f���mW��g'��r
�s4��n�ڒ�k��rΞ�r�
�s>2�s����������sV��x�rW2�3�/������/��3���sV��x�r��elW��g'��r
�s4��n�ڒ�k��r���rÕ�rÞ ����s��s4��f���b���s>6�5� 	���r?��������6�|7r��r�--����æ�Þ�rÞ�Þ�r���rÞ�mÞ�r�2�h�rÞ�r���rÞ�nÞ�r���k���l���l���nÕ�rßa�<^m;���� ��rV�x���rV��Ѝ��rR:�1W:�x=��r�rV
�fj��r>��W����4r
7rV���e��rR:�1W6�ic���W:��W����
rt��rÞB�c�����=c����m�� ����r�n��_��mÞ������
�rR��O������g���g���
rɞ�rê���rV��Ў��rR:�1W:��W��i�n�����n�<o��:�
r���rÕ�b �2�����g��y���rW2�ik���k�!�
3r4W�b�� ���8r�6���
rx��x9��r?��g$��r?��v����7���;��Bʜ�hÞ�nۜ����nۜ�B������������rÞ����r;�������
;r7��n�$gsǏsb�r��:���u���U�V��v����Þ--���n�R�Þ�rÞ�Þ�r���rÞ�oÞ�r��l�2�l�>�l���rÞ�gÞ�r�6�l���o���oÖ�oÆ�oö�o�V�o�F�o�v�o�f�o��o��rR��O��Þ�'�~-v�rÞ�l���lÒ�7��r���r�y�r?��Z3��7��r̞�7��r��ta���Ş�`Ξ�r���r-��kÞ�r��r��`���r���r-��kÞ�r��r!���O��?Þ�'��~v�rÞ�l���lÒ�7��r��ta���~��y�r8��ß�r���qB��~=��y=��r8��ß�r���qB��y��r���nÕ�nÞwa���~v�r7��e��oÞ�k7��r���r��Þ���nÞ�k7��r���r��Þ�F=
r���rç�ޚ7��r��ta���y��r���nÕ6kÞwa���~}v�r7��m���`Ò�7��r�ސ`Ξ�r���r-��kÞ�r��r��`���r���r-��kÞ�r��r!���O��lÞ�'��~=v�rÞ�l���lÕ/Þwa���7��r���jÒ�7��r���l�s�r1�_F�恻�v�r7��m���b���rÊ�2���jÎ�Þ�rÞ�Þ�r���rÞ�rÞ�r���rÞ�rÞ�rÕ�rÞ�mÞ��7����r��rW��y:��raV�j�+v
+vM*�x��rR.�^����'�m?.�i#��H���uV*��؞�rR"�1?��is��H�
+vΞ��'�yß�rM��w��b���6/�_mΞ�r�
'vV��p���s���r��mW&��7�/k!�%i��<vV&��7�,5�����p{��ns��v���m?���w��J����Ŕ�nǔ�"���mT��y¤�D��il!��{��lÞ�R&�x�rW&��7����r��r$��{�oa�!�='�m?.��{�oa���
?Ǩ{���r�
'vB��-9��??ᓪϔ"I��,i�������ϔ%��r��lx��n����%��r��lx��<?��{���nâ����_mW*�g3��r
'vM�Þ--���;r��Þ�rÞ�Þ�r�>�rÞ�oÞ�r3��$��s�;-Þ�r�"@���gÞ�rÚ�$'�s�;-Þ�rÞ�rÞ�rÞ�r�.�$#��s�;-���gÞ�r�6dÞ�m���rÞ�nÞ�rÒ�l�N�lâ�o�R�oÞ�r>+�r�������r6^�r�
rr7mh�rΞ�rê���� m�������r6^�r�
rr7mh�r59�n�������y�r?�e;����K�?�k�/�+������nS�la���<�r:�`��r;�s�$�rÞ�?�rR��?��7��c/�����r1���1rg
�h�����r��n������nS�la���<�r:�`��rr��W�� ���r6�����rO�r������r"��o*�eO��2���jS��y��rÞ�n������������r"��o*�eO��2���jS�����r�5�j���n�����0r&5�r<���?��7��c#�����r1����r]:�iÞ��y��?6��7��c#����� r1����4r]&�lÞ�v����2��r"��o*"�e��2���j����r=��f����
���"�-���rg�'r��r,�2����ú�Þ�rÞ�Þ�r���rÞ�rÞ�r���rÞ�dÞ�r��l��n��n�
�n�6�n�"�n���n�:�o�&�o���oÞ��3�)����'���d���r��s��=Þ��3��gΞ�rÝ�fÞ�y>��rΞ�r��r?��9W���(��rR��1W���7���W���W��j���y�rR6�m�4r>>�i_��mÞ�~�
�sV���W�����?���?�����_��y�Uy=�@EM2�m&��rÞ ����rÞBi[����r��r�� ����rÞ^�g��dΞ�r�7r������r>��g��mÞ��[��r�� a�
�sV
��+��rR��1���?���������KM�8��dΞ�r�#�s���mÞ�nǜ����rÞBs^��J=���ǜ��!am���r?���;�a��@s4��f��@s>��5��j��,�ǜ��!am���r?�*Q��ps4��j��ps>� ל�2?j�g!��r?j�v��r�ss���W=���ǜ��!aaÕ�rÞ����kϟ����l���kϞ����r>��l���d?����/l�� ����r?��r���R��--���r��Þ�rÞ�Þ�r� �rÞ�iÞ�r3�lö�l����#��r�J-��m��rÞ�rß�7c��l#��r��h"��s���n��rÞ�hÞ�rÞ�k���lú�o�z�o�j�o��oÕ�rÞ���mÞ��
rV�[&��K��oÞ�R�x�rW�A�⁻�� r�l�r<��rC����
r���r�
r��-a�f��s��sV�����=Þ�3� ����i�T��S��lÞ�n����m�������|�mÞ�y2��raT�f��s
�sM�����mÞ�'��n[���Þ�y=��r?*�-W���M��rR��1W����)���rÞ���i�nӜ����nӜ<��B���lÞ1�
�sV��iל��ל�lÞ�nw�M�������;���ל�2��7�;�)�πs���r�
+r>�� ��2?��g/��r?��7��
m���rÜ���";9��s��Ss&��y�r?���L��r�[s�� =��lh�r���rê�^=
�s9�-�������|��� )��,rq��e�s4��f��sbÀsV��hP�/p���ל�B���sXR���
�s`��n��s
�sM"�i�m�h�Þ--���Ö��Þ�rÞ�Þ�r�(�r���nÞ�r���o���l�*�hÞ�rÞ�rÞ�r������rÞ�rÞ�ræ�r���r���r�
�h�rÞ�r���rÞ�nÞ�r���kÊ�lÎ�o�Z�o�� rM"�x=��r�"�iÒ���rΞ�rÕ�rÞ�.���s8��m�o�r;���w��mÞ�k��r���r}mÕ�rÞ�lÞ�k��r���r}i��,r2��o�
/r���r��(r2��k1��r���j;�f-�y+r6��mÞ������<�r?�-���&�<�r?�5���rÞ 5�9�sV��g2��r��rÞ��+�����9+��2���r<� -���rÞBx?��r�'rW����mÞ�nS��j�h#m���r�L��3�clΞ�r��rV&�x?��r�
�s������r?��rXEM
�8+������O���
r���qB���W��cW�x=��r�
rV�=���Þ �����O��oÞ�W��K�DoÝom��r[����rX��j���lΞ�r��rV&�x?��r�
�s��mÞ�nS��j�h#m���r�L��˜�lϞ�`W��S���G�r��r��g/��r̟�G����O��lÞ�W��K�DoÝom���s��g/��r̟�G����O��oÞ�W��K�DoÝom���s>��˜�l?��ßJl?��0��rR��1���rÕ�rÞ71�
/r4��f���r���2�����6�Þ�rÞ�rÞ�r���rÞ�mÞ�r��h�rÞ�r���rÞ�mÞ�r���o�
�r|��3�)����rÞ�,���q4^�f���q�Ґu&��f���q>��h���
r'6��i?���?���������n�����5lW^��#��n��i�
�qɟ�rê�]=
�q���râ��'��ns��n���q78�n��vV�is�$i��v�̡;��L��<p��;�����=?�e��<p{���O���
�q�Tv'��R�gd��r��j�⓵�R���Þ�n7�����n7�)�$KvǏ{vV�+���BN�)�$vǏ;v>.�>?��j���r?��n�
�q>.�*?��n�$+vǏ�wH"�(��B.����<p��������=�����<p{��Ə��3����qU��vӎ�p���x*��rW�g&��r��j�V����A���r7�{vN�;v~��w.��w4��r���q>J�h���
�q`:�j��v�@t>h� �Ě9S� ��3l?��Þ--���>���Þ�rÞ�Þ�r��rÞ�hÞ�r3��$��s�j:-Þ�rß�r�.�mÞ�r�J�$��r�j:-Þ�rÞ�rÞ�r���r��l#��r��l#��r���n#��r�$#��r�j:-ß�rß�r�.m�Δm�"�rÞ�`Þ�r��l��l�V�l�R�l��lÊ�l��o�r�o��o�2�o�"�o�ґo��oÎ�o�
�r|��3�)����rÞ�,���q4^�f���q�Ґu&��f���q>��h���
r'6��i?���?���������n�����5lW^��#��n��i�
�qɟ�rê�]=
�q���râ��'��ns��n���q78�n��vV�is�$i��v�̡;��L��<p��;�����=?�e��<p{���O���
�q�Tv'��R�gd��r��j�⓵�R���Þ�n7�����n7�)�$KvǏ{vV�+���BN�)�$vǏ;v>.�>?��j���r?��n�
�q>.�*?��n�$+vǏ�wH"�(��B.����<p��������=�����<p{��Ə��3����qU��vӎ�p���x*��rW�g&��r��j�V����A���r7�{vN�;v~��w.��w4��r���q>J�h���
�q`:�j��v�@t>h� �Ě9S� ��3l?��Þ--���>���Þ�rÞ�Þ�r��rÞ�hÞ�r3��$��s�j:-Þ�rÞ�rÞ�rÞ�r�J�$��s�j:-Þ�rÞ�rÞ�rÞ�r��l#��s��l#��s���n#��s�$#��s�j:-Þ�rÞ�rÞ�rÞ�r�"�rÞ�`Þ�r��l��l�V�l�R�l��lÊ�l��o�r�o��o�2�o�"�o�ґo��oÎ�oÞ��7�)����'���a6�r�r
rǜ�����yÞ�r49�n��r�ěr��S����� ��
rr�6m7���c�����7c��-���r�
r';�y�r���lÞ��	�s���r��rq.�e��s4��b���sb�r�����m(��rÞ���8m�ᐦ��s���dΞ�r�#r�� ��8mi�r'C�r/
rH3�-����S��0')�r3
rV��l�/p���r`�0m$:�>�f��(#����'m?�����e��<r`��Bʜ��$/rǏ�s���Û����Tsf��B��<[������r#��s:��sڜ�s���l�� ��
r�r�*�nÞ�n�����n�)�$?rǏ�sV�+��B:��s���Þ��O��s>�g&��r����B�;9��s"��s���k5��rÞ�nO��M�r0r�r7� ������dW��;��r�{e���g��c�����Ɏ��3m$�s>��gz��r?��v���7s�mď�sV�+��Bڜ�Z�?�wӦ�7��3mďGsb��e���<?�r���`���=���u����F�m=���;��rW�Ƈ�r;��r/�--���Z�2�>Þ�rÞ�Þ�r���rÞ�nÞ�r�
�l��l��l��l���rÞ�eÞ�r�>�l�B�l���o���o���oÖ�oÆ�oæ�o�F�oÞ�r>+�r�̛mÞ�n[�����m��c#�����r1&��	r��r�7r���?2��[��h��ȧ���o*�e_��2ê�jo��y��rÞ�n������no������¡m0��_�����,m��?��;?r9*�v��b�,�?�rr��d?��k��r�̛mÞ�n[�����m��c'�����r1&��	r��r�'r��?2��[��h��ȧ���o*�e_��2ê�jo��y��rÞ�n������no������¡m0��_�����,m��?��;?r9*�v��b�,�?�rr��d?��{��m�̛mÞ�n[�����m��c+�����r1&��	r��r�/r���?2��[��h��ȧ���o*�e_��2ê�jo��y��rÞ�n������no������¡m0��_�����,m��?��;?r9*�v��b�,�?�rr��d?���l�̛mÞ�n[�����m��c/�����r1&��	r��r��sK��?2��[��h��ȧ���o*�e_��2ê�jo��y��rÞ�n������no������¡m0��_�����,m��?��;?r9*�v��b�,�?�rr��d?����l��xeÞ�dJ��r��q���rÞ--���.�j�
Þ�rÞ�Þ�r���rÞ�mÞ�r�
�o���rÞ�oÞ�r��n�2�n�.�nÞ�r>+�r�������r?���K������{�f��ol�8r�����-r:�����r3�$m���
��0' �r'�nlIc�y6����Þ��̞�r6�m=��{�f���r����Þ������*����|�6�r�v�m�����r�$m9
�g���r*�x�r*�s�����dl5i�b���rs�#r�� ��
rޒ�sa��r0�flW�I��al7��$j�����s�����&�
rޟ�����<?�<rv��$l�����s������&�
rޟ�����<?�<rv��$n��7��s������&�
rޟ�����<?�<rv��c$q��K��r0k�fÞ��� ����c���r������r�<r'w�*��K��r0k�f���rs�#r������r�<r's�*��K��r0k�f���rs�#r����
rޟ�����r;
rޝ�r6�4r4u�n��4r��mÞ�����%���r8��rÞ�Ξ�r��8rq�e��m;�)���y�r?��i���¡m0����6��$m��7���6��=��r��sV��I9�����<��s:��`��m;��s�$�rÞ�?��s��d?�����l����4�m�z�s9*�v��b�,���nǦ�r/�--���"�f�
Þ�rÞ�Þ�r���rÞ�mÞ�r�2�l���rÞ�iÞ�r�.�l�*�l���n���n�6�oÞ�r>+�r���6���m?��6��/{�f�
�rĜ�:���>���s4��nÓ�n�S�Kǟ�������m�r��:���=���8��c?� w��25��nÞ������KM�8��cW��_��yÜ2eÞ�y�r?:��3��lǫ���%o�� ���r��m���4=��{�f��
�rĜ�:���m;��:��>
�)���:�
3rǜ�>����+m��sB��~=��v���s��s���r�
�rĜ����r7��`���9���������m8��rÞ�&��+�����:�
3rǜ�>������m��s��:���=���y�r?�� w��24��j���s'�w��s&�r0��sq*�e��m?��?��n+���
�sV:��3�ri��=���9��k5��rÞ������KM>�8��cW���c��yÜ2��c�����r?��g2��r?�����8��W>�I���r���sɞ�rÚm;
rޝ�r0��sq*�e��m?��=W��������r���>��m��sV�I���m7��h���9���m=��ng�	�{�r;
rޝ�r5
r4��nÞ �)���:�
r��sH"����[����w���s��s���r�
�rĜ����r7��f���9���������q���rÞ--�����J�>Þ�rÞ�Þ�r���rÞ�nÞ�r�
�o���l��l���l���rÞ�jÞ�r���l���l���l���l���l���l���l���o�بs��"���Xs>B�g���r�:�r��xs4��jÕmÞ�����r;���Þ�no�����yO��r?Ғg$��r��r���p4��jÕ
mÞ�~���r;���Þ�n�����y��r?R�g$��r���r��xp4��jÕ3mÞ�����r;���Þ�no�����yU��r?ғg$��r��r���q4��jÕ�rÞ�~���r;���Þ�n�����yS��r?R�g$��r��r��xq4��jÕ�rÞ�T��Hs>r�v�b�iO��B^������)���pǏ�p>�v��iϝ�Bޝ�^������XpǏKp>r�v�b�iO��B^���ƛ�)���qǏ�q>�v��iϚ�Bޚ�^ƛ����XqǏKq>r�v�b�p��iG���G�!����K���K�Y���rC�q&�^Ƣ���B���b���B��b������"�9���y���Y�����B���b������"�9���yƂ���'��nW�����rV��gv��r��rÞ�T��r?�9W��w��rR�1W��7���W������
�s�0�0=�r>�iO�Y��:l3�����b���6/�--���n<&�Þ�rÞ�Þ�r���rÞ�rÞ�r�B�rÞ�Þ�r��l��l�R�o�B�o�r�o�b�o��o��o�2�o�"�o�Ғo�o��o��oÒ�oÂ�oò�oâ�o�R�o�B�o�r�o�b�o��o��o�2�o�"�o�ғo�o��o��oÒ�oÂ�oò�oâ�o�R�o�B�o�r�o�b�oÞ��3�)��
�r|�m>+�r���"��8r9*�v���,�jo�������+���s�XEM:�o��?.�io��&��#m6�� ��8r1f���r�?r�����8r���*�h�r���rç��Þ�i��ȧ��Xo$��W:�A�m��a���m�� ����i��ȧ��`m$��*?2�
ß�3��#�����[�%-���&��#m6"� �1;rg��h��ȧ���o*��e˜�����?��sʜ�?.�h��ȧ��m$�iÞ��s�����6�q�"��m��a��m?��h��ȧ���o*2�eo��R���nӜ��¡m0��ǜ�v��lm��F��m��c;��z��s1f��r��A��}���mÞ�y�rW���k�����rÞ�mÞ��s�����6������u���d��r��"��m��aC��m?��io��&��#m6�� ��8r1���s9���������nל�v�� m-�a+�"m;��`���m?���ӜA�T��s�y�T�ic�����r#��n�2�q��'is������m6����s9�����Z���y"��mΞ�rÕ�rÞ y�
7rV:�x�rΞ�r�
?r4�����&����lÞ�'O�r-�|j����¡m6b��i�:>���������r.��s�,r�m��a���m���C���_���������m7�����h�u�rÞ��3���<�--���ö�>Þ�rÞ�Þ�r���rÞ�nÞ�r�
�o��l�>�n��l���rÞ�oÞ�r�2�nÚ�nÖ�nÞ��+�)����'���gΞ�rÝ�fÞ�y>��rΞ�r��r?��9W���(��rR��1W���7���W���W��b���y�rR6�m�4r>>�i_��mÞ�~��rC���W�����7���7�����_��y�Uy=�@EM2�m&��rÞ ����rÞBi[����r��r�� ����rÞ^�g��dΞ�r�7r������r>��g��mÞ��[��j��l��rW
��+��rR��1���7����ߜ����KM�8ߜ�dΞ�r�#�s���mÞ�n?�����rÞBs^��"=���?���!am���r?���3�a��Xs4��f��Xs>��5��b�����i�
r}h�r4��n���s$Ks���r��s4��j��sǏ{sV���[�.�?�����(���BN��hÞ�n_�����n_��Bn�i�
r}h�r�	�sǏ+s���r���p4��j���pǏ�pV��pU�v��x9��r?��g$��r?��vӂ�������(B���oÞ�n������n���B��<��b���r���s��ksN�sn�+s��p>��pޝ�p��[p���d?�����m�� ����r?��r8���E��W��x#��rW�g&��rÞ�rÞ--���Z=��Þ�rÞ�Þ�r� �rÞ�iÞ�r3�lþ�l����#��s�J-Þ�rÞ�rÞ�rÞ�r���l#��s��h"��s����<6�rÞ�Þ�r���k���lÂ�o�B�o�r�o�b�o��o��o�2�o�"�o�Ғo�o��oÒ�oÂ�oò�oâ�o�R�o�B�o�
�r|��O�;e�"�y6��rR��yÇ���KM��x�r?��j;�m8����<�m3��� �y�r[�xe��y�r��8m/��rÞ����rC��j�����rR��1W��;�m����Õ�rÞ����y�rj��x�rj��x=��rj��;� ma��b��s
�s�����r�r[��mÞ�'���"�r��s���r�3rΞ��r�rS���r�rS���r�rG�����s>��x�rΞ�rÕ�rÞ�lÞ�n/���r�r��r�� m���rÞ2c����3���ß�j�"�vj
�s�������s����Õ�rÞ�q����ve���y<��r?��g$��r?����*M���]�r�rS��ă��B��)�$OsǏs����Ý������+my>�v�.�;��r�	/sǏ�p���p���r��rĝ�r���r7��nÞ����rӜ�s��sR�?s��=Þ�y ��r5��n�ڛmÞ�k;�mα�r�r�rK��r�� m�r�rW�2
����3���ß���7��{e��+Þ �y�r[��nÞ��r�r[��mÞ�'o�;�m�����#�s>�� ��2?��g/��rW��;�mx��nӜ�s��Þ��3��pʒg&��r��r�ʒ�՜s���6Õ�rÞ��� ���r?�����b���6�������r?�О;�m5��n��xe��d3��rr�rC��b���6���*�#r.�--�����Þ�rÞ�Þ�r���rÞ�lÞ�r��l��l���rÞ�dÞ�rÞ�l�ʒl�ƒlÎ�oî�o�N�o�n�o��o�.�o�ΒoÕ�rÞ�mÞ�k;��r�l�r<��rC��mÞ�y�r8��jÜ}l���m��y�r���n��r�ᐦΟ�rç��Ò��Y����+�rɞ�r��r�ᐦ?�s���g������r�� I>��/��lǫ�s_ ����M���[�I�M���/�����2l����k����
7r���rç���rÞ�������|l���nÞ�y�r��r�r��r:�-?&�g<��r:�i{��mÞ�n��n���n��B������r�
r}��r���h�&�5���x�rT�JV
�#�.�Þ����2h����k������sV6�pU���M���/�>y�r�
r��r^ ����r?��9W���9��rR6�1W���7���W6��O��f�
rɞ�rç��Ǡs��
��Þ�43��rq&�i{��j���8;�$r
��s����3��f�� a�
r`��j�7r
�sV��vj
7r���n���s���nÕ�rÞ��� ����r?��Ξ�r��r�ᐦ���r�H�jÞ�p���o����Ò�nM�{eÞ�~=��I��si�������r�t�+T�J���r�C����s	�2fÞ�����mÞ�y�rΞ�rÕ�rÞ ��<�r/���� ��rV�g5��rr&s�C��~=*�iM�oÒ�v���΃��oT�JV�'��y�r���r�r�
r:�,9��!3���?&�g<��r:�i{� ���o�0�*��r^^�=��r�Z�2���Ö�"Þ�rÞ�Þ�r���rÞ�lÞ�r��h�rÞ�����rÞ�Þ�ҿ��rÞ�rÞ�rÞ�rÞ�r���rÞ�jÞ�r�:�k���k���l�&�o���o���oê�o���h�rÞ�rÞ�r>+�r���*��r"��o**�ew��2���j{�5���mC>�>�.����s��&�&�8��W��k�/���lÞ�'5�r<��?�p��,i{�la���<� r:*�`��r;&�s�"�r���?� rz��W��k�/�3� ��(��W��k�/�3��W��k�/�3� ��7mm�r���m�"��7mm�rW��k�/�3� ��(���� 5���rÞ���-�s:��n���r3��n�>�����r��s�� ��7mm�rW��k�/�3��l�̛mÞ�yB��r?� ��2?��gd��r?��qb��iϜ�r���9��eW�'R��m1
�sɞ�rû��y�r?���ǜ�mÞ��ß�B�� ��7mh�ra:���s͜sV���s��W��k�/�3� ��7mm�r���o��oÞ��S���!|Þ��S���!a��7m?��r2��rÞ ��7mo�r���Þ�r|
rH6�-���������7mh�rÈs���r�
rH6�-���w�Äs4��f���r��sޜ�W��k�/�?���ÛmD��W��k�/�?� ��7mh�r$<���v���s�� ��7mh�r$<�Ƨ�s4?�n���s���Ξ�r��4rH.�~=��s^��o<��
���r?���k���!amÒ�v��������r
rH6�-9��q��,�S���!�nÝxe�s�� ��?mh�r6�r�vm=��g?��s@z�=��nk���r�r=����2���R����Þ�rÞ�Þ�r���rÞ�jÞ�r�J�o�z�oÞ�h�rÞ�����rÞ�m��lò�o��h�rÞ�����r���rÞ�eÞ�rÎ�k���lÆ�lÂ�l�*�n�&�n���o���oÒ�h�rÞ�r�
�r|�&q�mÞ�nO�"���,f��rR�^��=R��� <��rÞ�\�
r>R�9WR��w��rRN�1WR�iO���WN����ܾ�
�s�0����r>:�iW����#l3��K�� <�rOF��+���c�rOv�i�����DsqV�j�s4,�j��sivks8�����DsqV�j�s4/�j��sivks<�����DsqV�j�s4.�j��sivks����DsqV�j�s41�j��s�iÛs��5w����9O���-Ws;�����>l;����5w����9O���-Ws;�����9l;����5w����9O��mÞ��������ds42�j�����?s>~� ���2?�gq��r?�ث.�k��s>~� ���2?�gp��r?�ث.�o��s>~� ���2?�gs��r?�ث.�m��s>~� ���2?�gr��r?�_��r�z;siv?s:�����LsqV�j�s40�j��siv?s4�����LsqV�j�s43�j��siv?s6������rÞ���r>f�go��r�dsM*�i��"���,iO�� ���nO�:�w��r�i��"���,iO��#���nO�:�w��r�i��"���,iO��"���nO�:�w��r�i��"���,iO������nO������w�2�ث*�e��s>v� ���2?�gm��r?�ث*�g��s>v� ���2?�gl��r?�ث*�a��sɞ�r�#s>:�i�������6?
�iW���������Ɠ����0r>:��n��rRN�1WN��������r`5�j�_s
_sM��i_����� rV��gi��r
�s4��n�ڛlÞ��K��y�rR�Þ--����6�
Þ�rÞ�Þ�r���rÞ�mÞ�r��l���rÞ�oÞ�r�R�l��o�2�oÞ��7�)��
�r|�m>+�r�� ��(�mÞ�W�'Ξ�rç���o/���S�!x���r��km�#�m��S��h���=Ӝ�mÞ�yB��r��+;��z���r3��z��y��s>��r=Ϝs��j������l�̛mÞ�yB��r?� ��2?��g8��r?��qb��iϜ����9;��l��Ĳ���n�Ǣ���pZ~�K�n�:i��?6����.��m����r4ƌs�{~��g��mÚ�9���
��rǔ�s��Ĳ���n�Ǣ���pZ�<i��.���nk�r)㜐�;��.�
rt�]��Ku����#�����s�rs>�mK���,s9�����{��n�������n��?6���}$��?��q�4r��(r�����@�Ǿ�s���>���nk�Im4�(r�os&��g��mÚ�)���
��rǔ�s���R���v���m��rÞ��Þ�nO�"M��,i;��k���n;���Ϝ�~���s���j���
���r?"��O�!pU��sZ�H<��n��R���w�����r�B�sƔ�s	��m��s>��q�4r���mÞ�rÚ,��"�s�r�s��nÛsu�Ƭs�ᑉS��{��j���n��?6���}$��?��q�4r���s�����@�Ǿ�s������nk�Im�(r�� ��q.��s�����}����nk�r�̷���4r���v1�(r�� ��Om4�(r��p.��Ξ�rÕ/mÞ��-�s->�j���r3��j�>�����s�s���2�������Þ�rÞ�Þ�r��r���cÞ�r��l�N�o�~�o�n�o��o���o��o���h���sÞ����s�om��l�"�o��l���o���o�6�h�.�rÞ�����s������rÞ�rÞ�rÞ�rÞ�r���r���rÞ�kÞ�rÎ�l���oÖ�o��o�.�o�ΒoÒ�h���sÞ�rÞ��3�)����'���a��g��r��mb�$m����#��s����
������まĄ�r����
/�����2ǁ�Ą�r������=c��f���5������e���r��s���z��s9*�v���,�jǜ������/���˜XEM��ǜ�?��iǜ�&��#m6�� ��s1f��
�r��s��m���s���*�h�r���rç�A�i��ȧ��Xo$��W��A�m��a���m�� m���i��ȧ��`m$��*?��
�����ۜ����[�%����&��#m6"� �1�sg��h��ȧ���o*^�e�������?��s���?��h��ȧ��m$�iÞ��˜����6�q�z��m��a��m?Z�h��ȧ���o*��eǜ�R���n����¡m0�������lm����m��c;�����s1f��r���������mÞ�y�rWZ��ßi���rÞ�mÞ��˜����6��v������d��r��z��m��aC��m?Z�iǜ�&��#m6�� ��s1���Ts9���������n����� m-�a+�"m;��`���m?P�Ë���T��˜��T�i_�����r#��nÚ���'i˜�����m6����Ps9�����Z���y"��mΞ�rÕ�rÞ ��
�sV��x�rΞ�r�
�s4�����&����lÞ�'��r-�|j����¡m6b��i�:>���������r.��s�<r�m��a���m���W���c���������m7����h�u�r�� ��+m��sV>��-��rĜ�:���b���rÞ Û������<;��s
��s2��r�u�rÞ--�����>Þ�rÞ�Þ�r���rÞ�nÞ�r�
�o��l��n�>�l���rÞ�gÞ�r���l���l���l���l���l���lÚ�nâ�n�^�n���o���oÞ�r>+�r���mÞ����"��m7��"���v��8s��W�{�fm���&�+m�r*�m
r���,?r>.�f���r*������=K��n�*�5��<r�� ����s��"���<r7��n�� r��sH"��??� r
��"����K�%���s���jO��s��m�B:�)�$�sǏ�sb�r��"���E���k;��r5��n����W�++��lÞ�y=��r��4�,�s>��;��rג�G��v�T��s��J��m/��J���U�+my��vӦ���;5�<r:��sꜧs�ٛ�Þ��S��&�� !���bÞ�mÞ�d���r
#r>��qj
�sV�*Þ�n�*�5����K���##rV*�f��r���w���'�rW�������=K��h�*�5���m)
r'��*����=K��&��$�K�����i��ȧ���o*^�e���2ê�j������r�>�&���:�+m�r��&���?��s���"����K�%���s��jO��s��m�B:�)�$�sǏ�sb�r��"���E���y���rRF�m�Dp>���b�<�m?�a���b��Dp"���7��s
�m5
Cpǜ�����Ƌ��s�m5
_pǜ������_��>����'F�r)
r'��*��c��=���&�����(eƞ��;��Û����j$��/���<���;��\����j$��/���<���;��^����j$��/���<���;��X�3��j$��/���<��r;��m|B�m=���K���������Þ--����=��Þ�rÞ�Þ�r�d�r���gÞ�r2�l��l��$��s�n;-��#�6�oÞ�rÞ�r�F�$#��s�n;-Þ�mÞ�r��g�<:�o�
�l#��s��n#��s��l#��s��l#��s��i#��sØ�����rß����rß�m���rÞ�dÞ�r�*�l���lâ�l�^�n�Z�n�.�o���oÆ�oö�oæ�o�s�r?���rΞ�%��p�#r c��U��l���r$��/W����r����r�#r c��U��n��<m$��/W����r��]��l�#r c��U��h��m$��/W����r�����n�#r���l�rW�y=�����m|�c�����'O�9�)���lT�y?�����m|�c�����'��;�)���lT�y9��I���m|�c�����'��5�)���lT�y;��e���m|�c�����'��7�)���lT�y5�����m|�c�����'��1�)���lT�y7������m|�c�����'>�3�)��s�r9���
r'����S��c��P�����rǝ���������m�<r���jÒ�ĝ�&���*��im�(r���dÛ���������:�s�r7��p���?%�rb�3rj�;rr�#rz�+r��s
��s.s�r;��h�s�r;�����=s�r;��h���'��-�ya���w��r�r'��y��q���??�rb���=s�r;��h���_��������s�r5��p:�6�/��(/��{��j����:�����o���jÒ�T���jÒ����Ro���jÒ��ĝ����im�r���dÛ�g��k����*���	���r_�rf�7r ��7��rϞ��7��r�伩'��7��r��Gy6��h<��m���dÛ�_��c����*���	���r_�r ��7��r��Gv��r'c�>�7��rĝ���������m$�sƔ�s����>���6��W��P�����
r�r'��:��I��p6�2�2��(/�����i�>�����r_�rf�7rn��n���i���rÞ--�����j�>Þ�rÞ�Þ�r���rÞ�nÞ�r��l���o�
�l��l�&�rÞ�cÞ�r��l�>�l�:�l�6�l�2�l�.�l�*�l�&�l�"�l���l���l���l���l���o���oÞ�r>+�r������xe�0rC��0��c�����,m�����O)Þ�m���rc�3r�i�hÞ�nK�"!��,i������n��nÞ�n��2���n��mÞ�n'��2���n'��B6��lÞ�nǜ�2���nǜ�B֜�dÞ�n��2���n眐B��Ѷ�5�w�J�v��r��s6��s֜�s���s����=���7���i�r�K����laÇ���ݚ��fx=��r@��KH4�yZ�x?��r?��g��r?��x�r?��g��r?��v���x=��r?��g��r?��vӚ�x5��r?��g��r?��vӺ�7w�:mď�sɞ�rÜ����8-��s��s6��s֜�s��Cs&�r���rÞ�6��,m;��mÞ�n��2���y=��r?��g��r���r��s4��jÕ�rÞ�rß�i��������sǏ�s>��vӺ�7w�:mď�sC��KH4�?J�g%��r?J�r��կ������8-��s��s6��s֜�s��Cs�������n_�����v���rÞBpUZ�sZ�"=��n_��W�$��w�.o��ma��r�� ��|�����r=��n_���_��l�� ����v�
r��r�5m��r<��l��maÇ��|�Û����@��KH4�W��m6��r@��KH4�7�������r���s4��jÕ�rÞ���,m;��lÞ�n7��2���y5��r?��g��rΞ�rÕ�rß�6���sǏ�s>��vӚ�iל�B��&�5�wӪ��K�����r/�����j#9{s>�r<��r��s&��sƜ�s朣s���b�m��rV�y=��pUZ�sZ"��<��n_��W�$��w�n��ma��r�� ��|�����r=��n_����'nÞ�r��2���:��*Þ�rÞ�Þ�r���rÞ�kÞ�r��o��o�2�o�"�o��h�r�����������r���rÞ�aÞ�r�v�l�>�n�:�n���o���o���o���oÚ�oÊ�oú�oê�o�J�o�z�oÞ�r>+�r���k�h'm���rçoÕ�rÞ��'��r6�r4��n��r�������r?��rx�0r��o*>�ec�������g�����k��g�����
rǜ�"���&���<5�4rn�?rf�#r$>����jϞ��7��4W�v��0r'��6��K��s2�.�0��c�����m5��j�:���2����r ��r=���7��l�KmaÞ�r��r9
�g6��r6�
��0k������r$��g3��r&�??�0rj��W&�'���r�*��⁾ց�k�m#mϞ�����m���r7
'rH��&�m
'rt��k�m#m̞�G���8�c!Ò�G����8�c!Ó�n�S��_��lÞ�n{�"5��,i+�����n+�<{��n�����r��r9
�g6��r6��{�-���0r'��0�����<?�0rj��gΞ�rÝ�Þ�8�g��]n�����r$r��rk��p���������;?�r*��aW��+��='P�r6�r4��n��r�ۛmÞ�yß�r��f�,r>�8�fa���s4�����s���j��i7��o	������m�r4��n�
�s�ᐦ���r�H�F���EM��8_��b���7��Û����aW���7�Mp������e$��q���r6�r$��w�^o��mÞ��7�Mp���r=��+�)���&���*�����6�r�x�s+��rc��s������m6
�s'��w�Mn�������r?������y�rΟ�r���s7�"���r���3�����r/�����j#9�s>��r<��r_��s�������r?� a���v���rÞFI�S�K��s	�m3��r���'��0'�r6
�sV��ơ�r!c�r:��rơ�r�����r���<��y�rW��ơ�r���k5��rÞ�d#��r���r,�2�����R�:Þ�rÞ�Þ�r���rÞ�oÞ�r���h�r���*������r���rÞ�jÞ�r�:�l�6�l�2�l�.�l�*�l�>�n��o���o�
�r|�x��rΞ�r��r��-?��g��r͸qW��J�-1mê�:Ò�w��r.��mÞ ���r��-?ڒg��r͸qVڒxr%�r��mϞ�p��"�r�Wp>��i���mÞ�y�r���rÒ�Kɞ�rÕ�rÞ ���q
�qɞ�r�<�r���� ]��r�6�Ǖ�rÞ���Ò�w��r.��rA��qV�����rR��1W��x�r���m!��y�rj��x>��r?������eÞ�W��g��r
�qɞ�rç����oW���ǝ1������������'�����iÞ�y���rWj��S�q�<�r/���� ���qV��x�r��l!��nߚ����rÞl�̸q
�qV��g��r͸qV�xʞ�r��qɞ�r��qW �y=M�s^��?=��rÞ U�
�q���r�PA�3��^���f��pq#��n������6?z�i7��3�͸q>������r��-W���#�A�ǝ�0���6����-�������V�
�qV���ۚ�Hq��/m/��n���J�nߚ�iÞ�nۚ�ƕ�rÞF�ǝ�0���6W���_�A����F�
�p4 �j�� m��)m?���?��s�������e��������)�����
�qǜ�������+m�lqV��v��q�qH"���'��s��?+��q��{q��cq��kqB�qJ�qR���Ü�b���6W��g3��r��w��r.�--���f<��~�rÞ�Þ�rú�rÞ�eÞ�r2�l�z�$��sê;-������;?�,r���W��d#��rÖ�s���r�
rx.�x9��r?ڒd#��s����ߘ%����=���rÞ�r��l#��sÊ�d#��sÞ�sJ��b������s��4s�V�d#��rÞ�M��}���dÂ��$rɚ�d#�,r���j��,rǏ�sV��+s��B��$#��sê;-���n����<u�<��r��rÞ�aÞ�rò�kî�l�v�l�r�l�n�l�j�l�f�l�b�l��l��l��l��l��lÞ��3�)��
�r|��+�)����'���?*�is��&��#m6�� ��<r1��
r��!�S��k��"���nw��"�� m-�a+�"m;.�`���mW�q#r����������ZEM2�s��&����lÞ�'w�r6�m��a���m�� ����i��ȧ��hm$��W2�A�m��a���m���&��m��a��m���r�
#r4��j����?*�h��ȧ��m$�mÞ��&��rR&�1?"�is��&��#m6�� ��<r1v����s>��hw��!���rq��2��<m%�ê�������x�rΞ�r�
'rV2��k��mÞ�y�rW*�g!��r��rs�/r���=Þ�rN� r9���������n{��"�� m-�a+�"m;.�`C��m?"�h��ȧ��dm$��6��,r9*�v���,�j������n�)��s��!�'r�������m6�����rs�/r�)�&��0r��a��m?&�h��ȧ��m$�ê�y�rΞ�r�
'rV2��k��mÞ�y�rW*�g"��r��{�f5Õ�rÞ�M���o�G�m��a���m���>��i��ȧ��`m$������>�����=��r=��d��r���n���m?��n��${�f���s4��nÓ�n�S�Kǟ�r���F�ǜs4��nÓ�n�S�Kǟ�J������rß�sڜ�n���}���y�r?�� ��24��j���s'�w��s&��r0��sq��e��m?��W��W��ig��x#�����'��r9�zÞ�d��r�� �<�m?��mÞ���/n�䓘3��k5��rÞ�?�����KM��8?��cW���㜋yÜ2��㜋���r?��g2��r?�����8?��W��I���r��sɞ�rÚm;
�sޝ�r0��sq��e��m?��W��x ��rW>�g&��r�����#�s��3��rÞ--���ò�2Þ�rÞ�Þ�r���rÞ�kÞ�r�
�o�>�l���l�:�n��lÂ�l��l���rÞ�kÞ�rÞ�lÊ�lÆ�l�.�n���n���oÎ�oÞ�r>+�r������m?���K������y�r$%�nk��(���9k��Ξ�r���r?6�gy��r6�m.��rÞ���4r4$�f��4r���mÞ�x�����*m7������y�r$��nk��(���9k��Ξ�r���m?6�gy��r6�m.��rÞ���4r4$�f��4r���mÞ������*m7������Þfa��m���F����*�����6�r�v�m�����r3��r���J��0'��r'��mI��y6����Þ����r6�m=��
+��r?&�����lǫ�����˜`l������n��*������/�Þ�lǫ������ol����?��q�$r����!am�!��Þ�g?��s@����n{���˜�m����6���r�� m4��n�Ѽsɞ�r�ܼs����	��nm3��nò�]���4[��mq6�ik����������*���m?��^���rk��s������� k�����m?��^���müsV�IΟ��;��nò�]��4r����
rޟ�E���r��mI ���7�������cڞ�r��^���m��mI ����������cڞ�r��^���m��m���+����>��ɢ�
rޟ�E���<?��s��$��Þf���^���müsV�I��m7��nò�]���	� ����cڞ�r�� ����0������/m?������y�r���+��r�h�røs4��j�ϸs���kÞ�r&��rÞ/���mΞ�rÜ�x�r��xn������ k�����m?�߂��s��4���
��	>��+��:���n���͋����\s��מ��/��ɶ��cm;�߾��Tsd��rs��[s���n�6����4[��mq6�ik������=�mÞ�0��^���m$�s4#�j�Gs��^���;?�4r�����m��$r>@�h;��e���o*B�e���*���ǝ�+��Hs�os��?�i{�:h;��e���o*B�e���2���jG��y��rÞ�n�B�����n{���C��n���j�4�r�zKs9��+��b������nǦ�r/��2���r�:�.Þ�rÞ�Þ�r���rÞ�jÞ�r���oÖ�oÆ�oö�o�n�o��o�&�o���o���rÞ�dÞ�rò�lî�l�Z�l�R�l�N�l�B�n��n�6�o�^�o�V�h�2���rÞ��7�)��
�r|�m>+�r������ m-�a'�"m;>�`s��m%>�m��a��mÞ�y��r�����.����k���k�����~��2rɞ�rÕ�nÞxe�:�"a��b�7r
7rM�mm�(r&�?>�hw��!���rq�����8m��.��s�r���mÞ�W�x�r������rÞ������"�8��M�
��Þ��O�����r<��l� �.��$r�r9*�v���,�jc��������0=��m��c;�����s1����rc��s��!?6�h��ȧ���o*>�ec��j���n���¡m0����.���m�����s�7r�� r��a��m����"�m��4r>
�	 ��6���n���¡m0��c������m����m��c;��.��(r1�����s9�����j<��s:��`��m���Õ�rÞ�mÞ��#�	�����mÞ�y�rW6�g"��r��rc�+r��a��g��r��m{�$m���������まĄ�r����
˜�����まĄ�r����?9��sΜ�s��>���m$
rr
�s>
�p���g��rϞ�S��o/���'����y�r��jo���rt
�s`��nÛ�+��P��*9���.�
r����¡m0��c�����,m���.��O.Þ�m���s����"�8��.Ξ�rÕomÞ�iÞ�y�r���rÕ�r����s
�s`���7r
�s>��qj
7rM��+��dΆ�r��s�� �<�r?�A���y�rΞ�r��s�l�r2��rC��Ξ�r�
�s>��s�������Þ�y�rR��m6
�sV��M��ii�� A���rÞ����i!c�r)
�sV�����r�LE���<��y�rW����]x=��r��s�l�r2��rC��fW����]���X?��r;
�sM��m=��y�rW����/�"��rR6� ���mÞ�n��Q���v���rÞF�k�I���m/��r8��rÞ��Ξ�rÕ/mÞ�V�-'r->�>���r3��@��.�
r����¡m0��c�����,m���.��O.Þ�m���rc�+r	��m7
�sV��R��m;
�sM��m>�
n�� I���r?��r0��sq&�e��m?��o/��Þ--����B�&Þ�rÞ�Þ�r���rÞ�kÞ�r��lþ�h�rÞ����������������V���rÞ�r���rÞ�dÞ�râ�k���lÒ�lÎ�l�>�n�"�n���n���n���oÖ�o�
�r|��3�)��
�r|��+�)��
�r|��#�)��
�r|>�x�r$ �nϚ����nϚ�9ǖ�q	��i3����5l?J��K������B��q
�q`9�j�Gv�@v>�h� ���q��BƊ�y�v�rs� aƕ�rß�A� ƕ�rÞ�ql��m?ړ>?��B��6l?���
�q>ړ*?��ĒݧW
���=�Ϝq&��n��n�Üq7��n�рqV��i�$i�
rV��[���
rV��K�A��ɒ���r�pv4<����rӚ�q��sv .�y�rΟ�r��v��"y��qV�iW�����nW��{���~ƕ�rÞ����`v��'y=��s^>��?�v�s�2?j�s���l��<vY�3v՘q&&�n��n�Üq7��n�рqV��i�$i�܀qx��iW�����nW���ĝxn�`v��/v��r?ʑg!��rڑi���'����;;��q�v��*?��q��Ӛ����=ך}���q{���ך��Û�<?��q֚�*?���%����sm����=
r>ړ>?��B���r?��F�
�q>ړ*?� A��ɒ�<�r?���_��>���rӚ�q����=���%��s<
r'}�w�YoW�i��n�Üq7��n�рqV��i�$i�
�q�Lv`��nÊ����V��BƊ����YoϞ���oW���=W�i��n�Üq7��n�рqV��i�$i�
�q�Lv`��nÕ�rÞ����BƊ�����oϞ���oT��{� ����q��Ӛ����=ך}���q{���ך�(Ϛ�j;��W�l�9ǖ�q��BƊ�;?��qV���+m�Lv>ړ>?��B���r?��F�
�q>ړ*?� A��ɖ�+m��wV�i��n���w7��n���wV�i�$i�
�w��w`��nÛ�?��Û)���F�
r>ړ>?��v���r?��z�
�w>ړ*?� u���~��w
�w`��n�Gv
Gvǜ�J���N�+m$�q:��W�lď/v���w���r�
r4��f���rӚOv֚sv.��w6��w>��wƘ�wΘ�w֘�wޘ�w��~�
�-��vX>�����rÞ�b��Lt#7�n��a�<3l;��������q"7�ƛ���&u��7������6Ϟte�.�Þ--���V9n�Þ�rÞ�Þ�r�N�rÞ�aÞ�r3J�$��s�j:-Þ�rÞ�rÞ�rÞ�r�~�$��s�j:-Þ�rÞ�rÞ�rÞ�r��l#��s��l#��s��l#��s�>�l#��s�
�l#��s��l#��s��n#��s�j�o#��s��l#��s��n#��s��$#��s�j:-Þ�rÞ�rÞ�rÞ�r�
�rÞ�Þ�r�ڑkÎ�lÊ�l�~�l�z�l��l��l��l��l��lÞ�lÚ�lÖ�lÒ�lÎ�lÊ�lÆ�lÂ�lþ�lÒ�o�
�o�ޑo�ʑo���o�
�r|��3�)��
�r|��+�)��
�r|��#�)��
�r|>�{�f��
r4��jÕ�rÞ�,��q4^�f��q�Ґu:��~���q>J�h���
r'6���iך��ך��������n���b��5lWF��7��nÎ�A�
�qɟ�rê��?
�q���râ��'��n��n�Üq78�n�EvV��i�$i�Ev�̡�W��:Û߮����6���m��f��r���Ӛ�6�'�mW>��_���
rV��O���
�q�Lv'��z�ga��r��BƊ���z�h�mÞ�yß�r���,�q>���O������r/���Ě���՘qɞ�r��v>j�q	)�lǫ��c�4i?�p��,i���Ϛ�r.���=�-��p��6���m��f��r���Ӛ�6�'�m��+Ϛ�����r;�����v�s�2?j�s�ޑ1���n�������ěğ�Ӛ�jÒ�-�
���=i?ړ>?��B���r?��F�
�q>ړ*?� A��m���nÎ�A��=iϟ�
r'}�w�oW�i��n�Üq7��n�рqV��i�$i�
�q�Lv`��nÊ����\��BƊ����oϞ���oW>����0'X��K��6���m��f��r���Ӛ�6�'�mW��~��-��r�
r�Ӱ?9��q֚Ov&X�~��w ���[��:Û��K��6���m��f��r���Ӛ�6�'�mW��~��-��rΞ�rç�?9��q֚Ov&��~��w ���%��#?
r>ړ>?��B���r?��F�
�q>ړ*?� A��*y���jƜq��?�mÚ�v��??��q֚�nÒ���
rH"�~�i��n�Üq7��n�рqV��i�$i�
�q�pvH"���K��6���m�f��r��/��6�'�mW���-��rĜ�n���r�+mÀwV�i��n�Ðw7��n�єwV��i�$i�
�wØw>��9W�����rRF�1WF�v�ÄwÈwH"�y��e?�4��>�w�ޑp���x'��rW�g&��r��B�~�A�z���a��iĞ�qĖ�yĎ�AĆ�Iľ�;9��qV�/v>��c� l5��r���q>~�h���
�q`:�j�Gv�Lt>�h� �Ě9�� a��3l?��Þ--���V9n�Þ�rÞ�Þ�r�N�rÞ�aÞ�r3J�$��s�j:-Þ�rÞ�rÞ�rÞ�r�~�$��s�j:-Þ�rÞ�rÞ�rÞ�r��l#��s��l#��s��l#��s�>�l#��s�
�l#��s��l#��s��n#��s�j�o#��s��l#��s��n#��s��$#��s�j:-Þ�rÞ�rÞ�rÞ�r�
�rÞ�Þ�r�ڑkÎ�lÊ�l�~�l�z�l��l��l��l��l��lÞ�lÚ�lÖ�lÒ�lÎ�lÊ�lÆ�lÂ�lþ�lÒ�o�
�o�ޑo�ʑo���oÞ��3�)��
�r|��+�)����'���?*�is��&��#m6�� ��<r1v��#r���W�qS��k��"���nw��"�� m-�a+�"m;.�`s��mQ*�y^�U�_��>�����<r���*�h�r���rç�Þ�i��ȧ��Xo$��W6�A�m��a���m�� ����i��ȧ��`m$��?*�h��ȧ��m$�iÞ��w�����6�h�&��m��a��mΞ�r�<�m?�%���.��<r9*�v���,�js�����n��2�� m-�a+�"m;��`s��m�����s�+rڕ�rÞ�mÞ��{���
7rɞ�rÕ�rÞ !���m��?�<r��k5��rÞiw���¡m6���$r>.�hw��!���rq��"��lm%��.��m��a���m?��i��&��#m6�� ��,r1f����sP"���UEP*��{�UE>:�	 �����?�<r��%?*�ig�����r#��*��m��a��m���Õ�rÞ�mÞ��{���
7rɞ�rÕ�rÞ !���m��r2�$m���y=��r��o���8��i��ȧ��hm$���5�G�m��a���m������
����¡m6N��r8��rÞ�a��g��r��m{�$m���?������まĄ�r����
Ӝ�����まĄ�r����?9��s֜�s��n���m��rÞ��-�s:��>���ß��Û�ß�s<��n/�"��,g+��r�� ��.��0r���m4��fã�<��b��k5��rÞ��/����y�r���1<��b��k5��rÞ!�/����w���s'��y��?���c��>�����<�<r:.�`��m;��s�#�r���ß�n�.�-���s�"�mÞ�yB��r���rÕ�rÞ�lÞ�y��W��iß��ß����w���ß���7�w�Q���s��E?�����aW���-��rR��m*��rÞ�mÞ�n����rlm���mÞ����^��}l���m��r5��rÞ�������I�����`W��x�r��(i���->���ߜ��L�lÞ�W��\&h�r"��rÞ I�
�s���rÞBi����rlm�� I�
�s��s r�r=��������r��rÞ Y��Ps<�r?�!��Psɞ�r��sV��y=��x=��r�
#rV��g��r��d��r�1�mÞ�y��r?�� ���?��g��rǍ�s>���c��>�����<�<r:.�`��m;��s�#�r���?�<r��n��������H�������������gW��g3��r��n/�"��,g+��r�䓘3��r�u�rÞ--�����"Þ�rÞ�Þ�r���rÞ�jÞ�r�
�oö�h�r��������������������^���pß�m���rÞ�jÞ�r�Z�kÞ�lÊ�lÆ�l�.�n���n���oÎ�o��<rM��x=��r���iÒ���rΞ�rÕ�rÞ����s8��m�o�r;���w��mÞ�k��r���r}mÕ�rÞ�lÞ�k��r���r}i���s2��o�
�s���r���s2��k1��r���j;�f-�y�s6��mÞ������<�r?����"�<�r?����rÞ �9�sV��g2��r��sM��x=��r���iÒ�'��rΞ�rÕ�rÞ����s8��m�o�r?��%7��������mÞ�k'��r���r}mÕ�rÞ�lÞ�k'��r���r}i���sz��a��rW��x=��r8��ß�`����Þ�
�&�r6"�o�
�s���aÕ�rÞ��r`��n��s��s`��n��s���r�
�se��������6?��%7�����n��������lÞ��
�s�T���sz��a��r?����rW��x=��r��	��U�/��
�&�r6��o�
�s���r�Le���rÞ�f���sz��a��rW��x=��r������7���/�X�ǜq���EM���ǜu��\�ל�mÞ�n3�e������3���+�X�ßm���EM���ßy��\�Ӝy���rÞ^�Ϝy�
�sV�=���Þ����y���rÞF�˜��G�r��r��sV��x<��r�
�sV�=���Þ��ߜy���rÞF�˜��G�r��r�WsV��x>��r�
�sV�=���Þ����y���rÞF�˜��G�r��r��sV���˜�lÞ�W�=���Þ����y���rÞF�˜�lÞ�W�=���Þ����y���rÞF�˜�lÞ�W�=���Þ���y���rÞF�˜�lÞ�W�=���Þ����y���rÞF�˜�lÞ�W�=���Þ����y���rÞF�˜�lÞ�W�=���Þ���I���GP�킌�sP������s���ל\�Q���לX��GsPZ�y=�A�OXÏ�A�S@EMB��㜛l��s�SU��s�K��������GP�킌�sP�����Ws���ל\�QN��לX��wsVJ�A���Ӝ\�W~�AP���E�
Gs֒�GP�킌
ss��s�K�������l��s�S���}�S@EM^��ۜ�mÞ�]&@�y�rR���ۜ�r�W&T�yÞ�rR���mÞ�]&��y�rR���r�W&��yÞ�rR������mÞ�]&��y�rR^�����r�W&��yÞ�rR^��3��nÞ�R������cW���7���G�r��rW��q0
�s���r�Ha�
r���qB���ۜ�cW��x<��r�
�sV�=���Þ�b�gs ��f�s0����<�r?��ڛiÞ�y�rj��������6?��0��rR��1���rÕ�rÞ7	�
�s4��f���3��r���2���~�V�:Þ�rÞ�Þ�r���rÞ�lÞ�r��h�rÞ�����rÞ�r���rÞ�rÞ�r�
�r|�pΌ�K���(��'3�nS�����y�rW�i'���'�a�<�m/��� ��r�6��9'��!�� ���r���r�r'�/k����7m?������bÞ����rÞ ����rÞBi/����rlm?2�x�rW��3�/i[��mÞ�nc�����s
�sV
��7�2x����+���'�����7 3���s�����G�'"�y�rW2�x=��r���s�l�r2��rC������rÞ ���s�rɞ�r��rV�i'���'���
�ra����s
�s>�qj��sV������
�s�0�#��>hW>��_�����(ß�mÞ�n�98ß���sV��x>��r���l���rÕ�rÞ ���s�0r4��f���b�؀sD�mÞ�nß����nß�B������������rÞ�6�0�hÞ�Q�Z�%� q���rÞ��� ����rÞ�^� ����rÞBfj��r6��o��lÞ�Ξ�r�
�s��-W6�i'���'�����6W��ik�����'��F��y�r?��g$��r?��vӺ��k�%��������rÞ�6�0�hÞ�Q�Z����F��y�r?��g$��r?��vӺ�7��
mďSs���r���sl��rß�s���>
�s���rç�<
;rɞ�rê��<
;r���r�L�����=k�����rÞBx�rW��3�/�k���� ���r7���'�����7 3���
7rt
7r>V�9WV��k���� �<l7��� ��4r�6���4r�6�;r���V�7לlΞ�r���s4��j���sǏ�sV6�f��ryZ�v�F�x=��r?���	��r����F����F��y�r?��g$��r?��vӺ�7��
mďSs���r���sl��rß�s���>
�s���rç��?
;rV��y=��x=��r���K?��rÞ ����rÞBi/����rlmΞ�rÕ/mÞ��-�s->�r���r3��r�>�����sɞ�rÕ�rß�lÞ�����
7r7����4r����rÞ�r���r;��r���Q��4rq��e�Ps4�j��PsǏGs���r���sl��rß�s��Gs ���ǜ�jÞ�'���o��oÞ�49�n��4rV2�x<��r���rÞ ���s
7r>��9W��g��r
�s>6�qj��s��x�rΟ�rÕ�rÞ����1mW6�f��r6�7לolΞ�r���s4��j���sǏ�sV6�+���B���lÞ�n�9;9��s�Ss ����r���rÞ�6���6�9�sq��ac�r1��}���rß�sV
�x=��r�r 3��S���'��S��g���6/�--���N���Þ�rÞ�Þ�r�4�r���kÞ�r��n��l��l���h�rÞ����6���rÞ�lÞ�rÞ�m�p�bÞ�rÞ�rÞ�lÞ�rÞ�fÞ�����r���rÞ�kÞ�r���k���l�V�lÞ�oú�o�Z�o�F�oÒ�;��r���dã����rÞ�k���r/��lÞ��{�����r7��mÞ�y�rΞ�r��xsV��n��h����{���{�����r|"�i������r;������� ���ue����9's>r�iw��j���Ƨ���;��r��6%��xs>�g;��r���r�� sVJ��:��rR&�1W&��O��d�#+s>"�iO��k���"���>��rÞ���
Cs`��f�'s
'sM�4�))��(s>�f8��r��(s&����oÞ��{������r;��oÞ��{������r;��	Þ�nw���<�r7�%�� %�r'��/��.��r7��jã�.��2l!z�y��r?����`����{���{�����r|"�i������r;������ph���r�9's>:�g7��r���r�9's>�g7��r8�����r3������r7��iÞ�y�rΞ�rÕ�rÞ����xsɞ�r��r`���'s
'sM�2�))��(s>�g8��r"�iS��n��r4��f�� s>N�iS�����y�r?���S�����{���{�����r|"�i������r;��.���rÞ��
r`��f�'s
'sM�.�))��(s>�g8��r"�x�rj&�i������y�rj&�i;�����Ɨ�����{���{�����r|"�i������r;����=�ph���r�9's>:�g7��r���r��\sV��*��rR&�1W&��O���#+s>"�iO��k���"�/��>�\s`��n�r���nã�<��n���r�� sVJ��6��rR&�1W&��O��`�#+s>"�iO��k���"�c��>��rÞ7%��ls4��jÕ�rÞ�n�
r`��f�'s
'sM�'�))��(s>�f8��r��(s&E����n�<�r?���s�r?�����p?��rÞ���
Cs`��f�'s
'sM�0�))��(s>�f8��r��(s&�����nÞ�;��r&��y�r?N��S�����{���{�����r|"�i������r;��.���rÞ�n�
r`��f�'s
'sM� �))��(s>�g8��r"�i������n?�����y�rW��"��rR&�1W&��O���#+s>"�iO��k�����lÞ��{������r;��lÞ��{������r;� ��<�r?�%�� %�r'��/��.��r7��jã�.���i!z�y��r?��������{���{�����r|"�i������r;����>�ph���r�� sVJ����rR&�1W&��O���#+s>"�iO��k���"�w��>
Cs`��n�'s
'sM��))��(s>�f8��r��(s&�?�f��r�r>*�f��r�rΟ����;��r.��rÞ�n�
r`��f�'s
'sM�x�r?N��S�����{���{�����s4��n��\s4��nÕ�rÞ ��<�r;�%�� %�rVJ����rR&�1W&��O���<�r?�%�� %�r���r��sVJ����rR&�1W&��O��	Þ�nw���<�r7�%�� %�rVJ����rR&�1W&��O������r?���O��&���r?���O��r���h���rÊ�2���:�b�Þ�rÞ�Þ�r���rÞ�rÞ�r���rÞ�mÞ�r�"�lÞ�r>+�r���k�iqmƖ�s>>�g"��r?>����vr�2v_��v��r'��rc��s&��r<��Ξ�r��rH��~=��s^���8���O��|�Û���6Ξ�rÕ�rß�"��� c����
rH��?��g%��r?��r���/������8?�r��kϟ����y�rW�$��w��n�͛lÞ����lÞ��K�M��3��mÞ�p���rÞ�3��j�y<��rW��ӘhԦ�o�~�r���q?��r ��rÞ ��|��#�s>��f��r�����r���r�
r�#�s�� a���w���s���b��Kl�ћlÞ��K��n����#�s>�����rR�� ?����rÞ�3������lÞ��K�M����q���3��kϞ�������W��y=��3��=��,��=���r�
r��-$��/3��b�<�r;����sV��x�r���s&��r&�r���r�
r���b���r�T���s��mS�m=�yn�� a���w���s���b��Xo�ћlÞ��K��n����#�s>�����rR�� ?����rÞ�3��=��y=��rW�?�/+�)���s`��j��s���/��mÞ������I��y=��rW���s'���W�r��m8���S��l���<���7��nĝ�b���3���<��y�r?��i5��c#��v��s1&���s���s��s��?���ß�0��ǜ�v��,m��B��O+Þ�r���rǜ�s���r��s���a?>�g�r>�m8��rÞ�>������ǜ� ���r6�����s�␥!s�r/
�s��p��v��s&�r8��rÞ�<���7��hĝ�b���3��<��~�r���g��忞�w?�17��rq��i����� c����rΟ�p�.�i#��<���y<��rW�s��s���mÞ��K�Mx=��rW�3��?���rs�r��s���78��y�rW�$��w��k���lÞ��K�M��3�8������b����眚mÞ�'��r��rÞ�
�sǜ�b���røsɞ�rÜ�x�r���r3��s&l�r/��rÞ ��|�>�健'i�r8���M��i!��r=���� Q���3�����ȓ���n���Y���n��8���=��m���r�
r�#�s�� ]���w���s���b���i�� Q���rÞ�r3�����rR��1Ξ�r�
�s`��j��s
�sɞ�rç�>��~�r P�r/
�s��p��v��s&=�r7�����5���r.����4���y�r��6h��mS����W��y<��3��=�����fϟQ���r;��ϟQ�<�r;��mÞ�'��r
�sɞ�rÕ�b �2:����/��y�rW�����rR��1W��x�r���h��mS�m=�^k�� ]���w���s���b��k�ɛmÞ�nß�d���<��s:��`{��rT��J$��s^��)9��nӜm���c#��v��s1����s�~%mÞ�r��v���m5��sX��9��nc��m���9c��k5��rÞ�i�: Ýsq���r��a3��r%��m?�����W��y>��3��=�����k5��r��^k�� ]���w���s���b��^k��rR�m=��8�g����k��R��� ��2���s�"���rW�yä�ur�����r3��oÞ��K�M�?��q��rÞ ��|U���r��sV��v�øsìs'��Z�7��r��b����Z�;;�<rb�/r"��l���l���Þ�r5�rX���Þ��M��8��y�r?�i5��c#��v��s1&���s���s�[s���?���O��0��ǜ�v��,m��B��O+Þ�r���rǜ�s�����[s���kϟ1���e���jN��7��kϞ1Þ�y�r?�i5��c#��v��s1&���s���s�Cs6��?���O��0��ǜ�v��,m��B��O+Þ�r���rǜ�s��k�im?���O��0��ǜ�v��,m��B�r>��rc��s'��w���
r���<�Ds:F�`��r;B����rÞ��1Û߮��b���;��sҜGs���n�>�-��Le���l:��8�g�Ý�=��r4��n��rE��q�.���/r���s���n�>�=���e���l:��nӜ����c#��v��s1����s�~/mÞ�r��v���m5�rXJ�t;��r=����2���Z���6Þ�r��Þ�r���rÞ�nÞ�r���lî�lö�l��h���rc��r���rÞ�fÞ�r���k���lò�l�^�l�Z�lÚ�nÎ�n�F�n�B�n�>�o���o���o����=��rÕ�rÞ�mÞ�ng����r3�le��#r2��rΞ�r�
3rl�0r'>�/c�����?m|�i_������{����8%�r����>��3��7Þ�RB��yd��r����r?��g$��r?��i�������3�����r;�����s4��j���s>���[��mÞ�Ɩ#r>��g]��r?��q�
�;5��s*�#r��s ��3���Þ�RB��yU��r��w��r���r�L�:���r;��:������lgC��yR��r��r��rô������r��r�L�s�>�_��(��{V��n�����lgC��y���r��<l*��Ý����r�A�rç���� rX��mW�oÕ�rÞ�E��&��q�
��3��Þ�'o�4w�mƞ rB��y��r��Hl*��Ý����r���rç��� rT��mW�oÕ�rÞ���dÞ�n�����n��{V�oÕ�rÞ����&��q�
��3��Þ�'��4w�mƞ rB��y��r���l*��Ý����r���rç�=� rP��mW�oÕ�rÞ�}��&��q�
��3��Þ�'7�4w�mƞ rB��y��r�� o*��Ý����r�n�rç��=� rL��mW�oÕmÞ����&��q�
��3���Þ�'K�4w�mƞ rB��yQ��r���o*��Ý����r��rç�Y<� rH��mW�oÕ�rÞ����eÞ�n�����n��{V�oÕ�rÞ�5��&��q�
��3��P�'��4w�mƞ rB��y5��r���o*��Ý����r���rç�%<� rD��mW�oÕImÞ�a��&��q�
��3���Þ�'�4w�mƞ rB��yg��r��dn*��Ý����r�B�rç�<� r@��mW�oÕJmÞ����&��q�
��3���Þ�'��4w�omƞ rB��y���r���n����,�s>��7ۜimq��i�����rÞ�p�*�i+������n+��{V��h�*�5����3���Þ�'5�4��rq��i��J�c� ��:�
rɞ�rê�uv����m3���������rw��s�oÕRmÞ����Z�b� ��
�؄s��"5���sV�x�r���!���s4 �b���sƔr��&�����r�_�rç�O>شs��"���s����,�s>���[��mÞ�Ɩ#r>��g]��r?��q�
�;9� r
��sB��y���r���i����,�s>��7ۜfmq��i�����rÞ�p�*�i+������n+��{V��h�*�5����3���Þ�'�4�amq��i��J�k� ��:�
rɞ�rê�uv����m3���������rw��s�oÕ�mÞ����Z�j� ��
�؄s��"5���sV�x�r���!���s4 �b���sƔr��&�����rμ�rç�s9شs��"���s����,�s>���[��mÞ�Ɩ#r>��g]��r?��q�
�;9� r
��sB��y��r��*k���,�s>��7ۜ~mq��i�����rÞ�p�*�i+������n+��{V��h�*�5����3��Q�'m�4�ymq��i��J�s� ��:�
rɞ�rê�uv����m3���������rw��s�oÕ�rÞ����Z��� ��
�؄s��"5���sV�x�r���!���s4 �b���sƔr��&�����r���rç�8شs
�"���s���,�s>���[��mÞ�Ɩ#r>��g]��r?��q�
�;9� r
��sB��y��r��j���,�s>��7ۜtmq��i�����rÞ�p�*�i+������n+��{V��h�*�5����3��>Þ�'I�4�wmq��i��J�y� ��:�
rɞ�rê�uv����m3���������rw��s�oÕ�rÞ����Z�x� ��
�؄s��"5���sV�x�r���!���s4 �b���sƔr��&�����r���rç�;;شs��"���s���,�s>���[��mÞ�Ɩ#r>��g]��r?��q�
�;9� r
��sB��y��r��e���,�s>��7ۜLmq��i�����rÞ�p�*�i+������n+��{V��h�*�5����3��:Þ�'��4�Omq��i��J��� ��:�
rɞ�rê�uv����m3���������rw��s�oÕ�rÞ�7��Z�A� ��
�؄s��"5���sV�x�r���!���s4 �b���sƔr��&�����r���rç��:شs��"���s���,�s>���[��mÞ�Ɩ#r>��g]��r?��q�
�;9� r
��sB��y���r��d*�Ý����r���rç��:� r���mW�oÕ�rÞ����&�G�q�
��3���Þ�'G�4w�Gmƞ rB��y���r��Pd*�Ý����r�L�rç�]5� r���mW�oÕBmÞ����&�K�q�
��3���Þ�'��4w�Cmƞ rB��y���r���d*�Ý����r�N�rç�	5� r���mW�oÕ[mÞ���&�O�q�
��3���Þ�'/�4w�_mƞ r>
�7w�
mf��:��r�~�rê�uڜ�
����C�lÝ!������zÞ--����b�
Þ�rÞ�Þ�r���rÞ�mÞ�r�
�o���rÞ�jÞ�r��l�>�l���o���o���o���oÖ�o�:�h�r���rÞ�r>+�r���m?�hÞ�m���r=�����m<������g?��rƇ�r������r���r��#���,io��i���no��.����������{m��xeê�$���r�L��o��oÞ�k;��mv�e��s4��b���sb��eê�8?�8r��c������r���Þ�g:��rƇ�r���2�f5��r��s	2�m2r�r�� =���r�=�r�� =���la��nÕ�rÞBvĞ����iO��iÞ�vI���O��y<�UEM�m2
�s�
r���r�H�w�� =���j���s��s(��r;
�sޝ�r5��rÞ�"�no��c���9o��nǦ�o/��r%s�rK���3��rR��1W���0���v���r��rÞ7��s��Ϝ�B�� }���r;���Ӝ�F��7�ל�t�'�r��~���A���nŜ��Øs7��n�ќsV��iŜ$�ܜs>��s3��Ϝ��?��>*��~���r�Γu��t���rƧ�sq�e�8r4��j�
�s>��**�����(r.�3v��v#��r'��rϜ�s��������kϟu���l��mS��m1s�rI�u����=��no��c���9o��nǦ�l����<�r?���<�r?��ql�oo��rR�����kϞu���;�mT��'G�r6�8r4��n��8r�␥���c$���)��r�0�=��~��s ��r8���˜�`������s���o�������r?������v���r+��ra��n���ra��nå��'��r8���˜�<��~��s��ye���˜���a?2�g0��r2�m?��m=�Ɵ;�m$��nϜ��Ϝ���������mÞ��Ϙs&�r6�8r4��n��8r�␥���b�������rÞ����a?2�g0��r2�m?��m=��y�r$��no�����no��9Ɔ�rϞ�����y?��r?2�g#��r?2�x9��r?��g#��r?��vӪ��Ƈ�r���h�2�9���m(�8r4��n��8rb��e�N�9o��r����#�s�� ����w�Øs���~��#i������� o������r?��~���rÜsn�����rϜ�s	2�a��W��y<��Ϝ�=�������,;r>2�f��r����Ӝ;e���<?��sҜ����2k�� ����w�Øs���~���i������� o������r?��~���rÜsn�����rϜ�s	2�a��W��y>��Ϝ�=����.��,;r>2�f��r��x?��r��+�����r7���>�~�2�r'��nÒ�}���ro��s����9������hĝ�~���Ϝ��>��4_��rq2�io��>���r;��>��(r��B��Ϝ;e���Ϝ�h�2�9���a��W��y8��Ϝ�=�����eϟwe�^�r�r�"���8r7��n�Øs'�����;��r��~���8o��Ξ�rÕ�rß�lÞ�;���r�r�����Ϝ;e���Ϝ��9��r��rÞ�rß�x=��r$���xe���g��r���;��r��m��rÞ�j���!_��2?2�g��r?2�7��rf�/8o���9���;��r$�����;��r��m=��;��m��k��xe���d��r��mÞ�4_��rq2�io�����Ϝ���*9���r;��B���r�ΛmÞ����.��� ������r?��F���r������r;�����~���A�V�;9�8r��s&�r�8r"�?������	>���:���no��͏����s�������o��d���������4_��rq2�io�����Ϝ����B��sΟ��#��nÒ�}��8r�����s���r������r8��rÞ�l������ o������r?�߂��(r�"���s7��n��@sɞ�r��\s����(�����Ӝ�jÛ�yG�rj��3���F���r������r;�����~���A�V��J�;9�8r��s&��r�8r"�?������	>���:���no��͏����s�������o��d���������4_��rq2�io�����Ϝ�9���B��sΟ��#��nÒ�}��8r��=���������r;��fT\�i�����kT\�p��d��r�/����� o������r?�ߺ���rÞ�;��Ts������ל�h��*9���r;�����rϜ�s֜Ws������m8��rÞ�l������ o������r?�߂��(r�"���s7��n��@sɞ�r��\s��
��(�����Ӝ�jÛ�yª�rj��3���F���r������r;�����~���A�V��J�;9�8r��s&��r�8r"�?������	>���:���no��͏����s�������o��d���������4_��rq2�io�����Ϝ�5���B��sΟ��#��nÒ�}��8r��m���������r;��fT\�i�����kT\�p��r8����ޯ�����r?��B���rÞxeê�g��r����mÞ�p���rÞB3Ӝ%����s4��f���sb�ps��~���;?�8r�����r�
ss'��y�r����'y�r
sst��rÞ ����rΞ�rÜ��?z� _��2?2�g��r?2��z�8o��l�؛mÞ�yß�r�1�,;r>2�;��r?��g��r?��r��������8?�8r����m��dsVv�y=��pU"�sZ�4��Ƨ������ƫ�Mv��g��rR@�m>��g������m����r��r�"���s>6�g��r?6�p���f��rV�;��m4��n�$;r>��g,��r?��x�rΟ�rÕ�rÞ�j��Ts����ל{e���g��ry&�i�����n����Þ�k;��mv"�e��p4��f���p��2�=�1;��
˝ ����E���Z���<;��sҜ�s���b�2��6�%���5���E���f��xeê�g��r���;��r����l�؛mÞ�yß�r�1�,;r>2�;��r?��g��r?��r��������8?�8r��a2�g��r2�m�8r4!�n�
ws�ᐦ���r�H�F���EM��8o��`W�����M�;��r��xe���;��='x�r3��rÞ ��|;e���r6�8r4��n��8r�؛mÞ�yß�r�1�,;r>2�;��r?��g��r?��r�����^���8?�8r��2�g��rW��y=��x=��r����Ą������������Y�|(�ƞ�����jÛ���`Ξ�r�
�p�#�p��xe�������Ϝ;e���Ϝ�l������ o������s4��j���s���s7��n��\s���Õ�rÞ�rß�x=��r$��0���B���rÀs������r+�ɺ�ȓJ:�Pm��~���A�V����ro��s��xe��;��='��r5�.mo���Þ��;� m$��w��`��xe���;� m��xe�>�y.��r���`��Þ�;�m�B����� �����4s4��j��4s���s7��n��Ts������r?�*����s4��j���sɞ�rÕ�rß�lÞ�;�Һ�Üs'����;��r4���$'s>֒g,��r?֒vƒƝ��p�"�v#��r'��rϜ�s֜Ws��������&�9�֒)��y���mÞ�|�����(m7������y�r$%�no��.���9o��Ξ�r��*m?2�g��r2�m.��rÞ�+��8r4"�f��8r���mÞ�{�����(m7������y�r$)�no��.���9o��Ξ�r��&m?2�g��r2�m.��rÞ�'��8r4"�f��8r��mÞ�;�Pm5*�jÞ�d��r���j�Z�!_��25-�nÞ�d��r��xe�Z�;��m5,�jÞ�
��r?f�;��r�ᐦ�	+r�KpM��?f�qr�r�/�?�)�ƞ�����jÛ�_��,��,;r>2�f��r��x�rΟ�rÕ�rÞ�B�Øs'/��������=���nÒ�}��8r�+����� o������r?��F���rÞ�rß�x=��r��Ϝ�"���B��?mW��f��r��?9��sҜ�s	2�m}�rl�"���8r7��n�ќsɞ�rÕ�rß�lÞ�0Ӝ�~��9mW��f��r��??��sҜ����.7_��rq2�io�����=Ӝ�mÞ�yß�r���r�ܜs��o� ����r+�߮���rϜ�s	2�m2�8r7��nÇ=��8r����-r:��!���r0
�pV��IΟ��#��W��I>f�qr�r�/kÞ���jW��I���?f�qr�r�/pR��v.��' �r,�ds��xe���-���������s_2�i�������!��;����p��i�������n����W����Ϝ����ɞ;��rh�r��}��:m;��nÒ�}���r_�;r��s >�r=�L��r2�l��ds��xe���-��r��l������s45�b��s���j��Ts
Ws>f�qr�r�/�7��F�� A�
�p>��9W��h��~�� y���rÞ�����6W��i����W��i�������!�fÚ7?;��sҜ�s���j���������r=��r4�ds�Kp���c�������r���],�?x=��r$��n���Ƌ��j��s
�s������s
�s'7�nϜ��Ϝ�mÞ�dk��r
�s;���Ú7?;��sҜ�s���c�������r���=,�?x=��r$��n���Ƌ��j��s
�s������s
�s'7�nϜ��Ϝ�mÞ�dk��r
�s;���Ú7?;��sҜ�s���d�������F�����r?�xe�B�w�Øs'����;�DmĜ�F��ɺ���r�\s���Û���������7m;��lÞ�y=��r&�io�{e�~�qU�v���i����k��:��6m/��:�����&m?ƒg��r��~���A�V��J��z�;1�8r��sj�'s
��p ��r=��y�r$(�no��.���9o��l��ye���%�����r�r�r���&���r5s�rk��/��k;�Pm5;�nÞ�no��c���9o��k5��rÞ�;��r'	�r2�8r7��nÇ=��8r������� o������r?��~��0m$�s4-�n�Ϙs������m�r�"���8r7��n�Øs':������yÜ2e���rϜ�s	2�m0�3mW��I��2m7��$?�;��mØs'�������r0<�f���rϜ�s�����r�r���Ϝ�����B�
�sޟ�����<?��sҜ�c$ ����r0<�fÞ����p��4_��rq2�io�����=Ӝ�mÞ�0Ӝ�~��0m$�s4��j�Ks��~���;?�8r��l��ye���'o�r*��rÞ�j�Z�!_��25��j�Ks�␥������,;r>2�i��
���n��sΜ�4���=���mÞ�yß�r���r���rN�Ӝ����F�r�r'�������;e���<5��sҜ�s��_s������m8�	mÞ�a2�g��r2�m��rÞ�rß�7_��rq2�io�{e���n��1���n��;;�7��xp���n�2�9���o��-���Ư��lǫ�lÞ�ߋXv؆���8r��xe���_��0'o�r1
wpVr��o��R��w�����2�r��c���R���r���)��y�rWr��o��R�o��2���9o��4Ξ�rÕ�rß����� o����r�r/��>���r/��>���j#9�s>r�r<��ro��s������/m?� �ƒ�v���rÞFI�S�K�wp	2�m0r�r/���Û�}��`Wv����M�;��m!*�r5�mo��V��;��m$��w���mÞ�Ư�M�;��m����Þ�r6�%m4�n��|p�� �ƕ�rÞ�0'v�r5
pn��jÞ�|������=���cWn�x�r���(��Ƴ�;e���r6�m4�n��|p�� �ƕ�rÞ�0'��r4
pry�rw��a$&�gY��rn�m0
pɞ�rÛ�4��dWn��;�hm���%��
m?���ƞ�Ƴ��mÞ�w���� �ƚ4�;�dm���'��
m?���ƞ�Ƴ��mÞ�w�1�� �ƚؖ;�<m���$��
m?��~����;��m��m4s�r������?2�g"��r?2�qsz�r�����/x<��r?2�g#��rΞ�rÕ�rß���r�r���>���r/��>���j#9�s;��z�8?�8r��dƒm�_m�����6�r�vmÞ�Ξ�rÕ�rÞ�j�V�p���j�����y�rΞ�r���rÞ��m7��r���mÞ�y�r>�p�������rÞ�y�rΞ�r���r랒�m?��r�mÞ�y�rΞ�r�r�r�/kÞ��m7��r�{e���S��Ϝ���� o������r?��B���F��m�Ts"���,�s>��f��rN�J�O����;e���<1��sҜ�s��_s��Op������mr�r[�xe���gN��rƧ�s7�n�Üsn��f���rϜ�s��xe�R�;�Xm$�sɞ�r��8r4��j��8rǏ�sb��eâ�89��sn��s���6�2�r���4Ξ�rÕ�rß����� o����r�r;��>���r/��>���j#9�s>j�r<��ro��s���V���nG��ƒ�v��)�����r,�p�� ��|�jÛ�Z��f>��K��uj��?��ek��<�r:�`{�mT��y=I��o������ns��Ƃ�����o*�eK��2���s�0!���r��a7��r����*�m�<pV2�I:6�b3�����r1����1?pg*�hÞ�m���r=��n��!ƞ�ns��Ƃ�����o*�eK��2���s�0!���r��a7��r����*�m�<pV2�I:6�b'�����r1����1?pg*�hÞ�m���r=��n��!ƞ�ns��Ƃ�����o*�eK��2���s�0!���r��a7��r����*�m*��rÞ ����r�����r?�ll���mÞ��o��jÞ�p�������rÞ�y�rW2�j;��m�o�rQ��rÞ�Ξ�rÕ�rÞ ��r�r�/kÞ��m7��r��mW2��;��rl�r���"�
;p��4p3��K�����,mJ��"ƜO+Þ�r���rK�?p��.���	Ξ�rÕ�rß����� o�����p�� ��|�>���r/��>��]�����y6�?.��o��ek��<�r:�`�m;.�5��r����.�;;�8r��sj���"�l�śmÞ�yß�r��,;r>2�iG��Wj��?��g��r?��s���lÚ�qU��?.��o��ek��<�r:�`�m;.��r����.�;9�8r��s��xe��y���r�
;pǜ�~��m;��~���;�xm?.��o��ek��<�r:�`�m;.��o��rÞϜ��ÛҮ?֓�o��ek��<� p:*�`�m;֓���rÞӜ��Û߮��~���;�rr�#p
��n�2�9�������!�؟;�rmƖ+r>2�g"��r?2�;��mƛra�9��Ħ���8?�8r~��9!��b��?.��o��ek��<�r:�`�m;.�s���rÞ�?�rr��j��uj��l����Ɯm��|�r5��G���N�~�v�rמ�gΞ�rÝ��Þ��;� m���rç�!��no������9o��k5��rÞ�iH�:�Ýs����r��a7��r%�m3r�r��lÞ�'��r.�(r�r�m�a��m�����m�ak�m���rÕ�rÞ�mÞ�y�rΞ�rÕ�rß��mm'����l������m6R��Þ�r8��rÞ�a?2�gC��r2�m���r�*�2���.=:��Þ�r���Þ�r��rÞ�Þ�ræ�l�6�n��o��o�R�o�B�o�
�o�:�o�j�h�r����������rÞ�m�r�h�r����������������^���rÞ�m�^�h�rÞ�����r��rÞ�Þ�rÒ�lÎ�lÊ�l�V�l�N�l�J�l�~�l�z�l��n�.�n�*�n�֓n�2�o���oê�o�6�o�&�o�֒o�ƒo���o��oÖ�oö�o�R�h�rÞ�m�=�rÞ��7�)����'������;� ����r;��������oÞ�nO�"���,i��l���n�<O��n���=���y=��r?� c��2?��g<��r?��p���f?��r��}����,r��2���rÞ���-r:�����r3��mÞ�yß�r9��!Ӝ�2?���>�*���m�� #��R���r/��R���j#9�s>��r<��s��2���m���M���v���qҸ�m1��W���v1��?��d8��r��mÞ���Mq'�s��U���+��n�� ���r��c/�����s1��d��s��mC��r���s	��m�sǝ%-�����r>��:��<��s:��`��r;��4��������8��;T��v�$/r�sW��i;��e���o*��e���2���j���g��l?��s���2���n�� ���r��c/�����s1��d��s�~%mÞ�r�����m�sW��i;��e���o*��e���2���j���y��rÞ�næ����n�� ���r��c+�����s1��d��s�~%mÞ�r�����m��rÞɲ����� Û�#��f���<?��s���k5��rÞyi�� ���r��c#�����s1��d��s]��iÞ��y��?V��3��j���r0�������,m5����s=��r����s��n�� ���r��c/�����Xs1��d��\s�~/mÞ�r������V��N�;9�,r��s�s���r>��:��<��s:��`��r;�����rÞ+ß�n�� ���r��c#�����Ps1��d��Ts]��lÞ�v�������r>��:��<�Xs:R�`��r;N�s���r���7��s��Ss��[s���h���=���m��sW��i;��e���o*��e���2���j��-���r�>%m�����r>��:��<�Ps:Z�`��r;V����rÞ��	?r�\sW��i;��e���o*R�e���2���j�����r=��fæ��Z��R����r��s�#E��v��y=��'��r!��r�:�y���r��rĝ����r;�����i1��c���6�aÚ�#�h��ɲ���rk�����r�%�pJ�F��>�����`�h�rĜȒ��ɖ��r�ts���7��sr�j�q���JW��w��|s4��f���r#��s��Gs��Os��ws��s���2��=���M䜛o��T��Ξ�rÚ��� Û�#��f���#��k5��rÞ�,�����#��Û�#���>�.,�����#�h��ɲ���r4��n��@s�Hs���r��rĝȊ���r7��d����J��B�m=�=���M䜛n�����?��h(�����r*���/r&��rc�ds$��8��r��hW�����=?��gÞ�#�h��ɲ���rÞɆ��Ɋ��r�Hs7��r��Ls�psH��y��i�����n��Bh�$rǏ�sH��(s��BJ�h�$�sǏs7��r�$7sǏ'sH��(Ӝ�B
�h�$�pǏ�pɞ�rÕ�rß�lÞ�#�����r���g��ry�vӖ��>�*E���U���r���(���B���r�h�ryF�v�v��>�*�ƛ�����rÞ*�ƛ����ry&�v�֓Þf=�$�qǏ�qH��(;��Bʚ�r�hm�	�qǏ�qH��(���B���r�h'm�	GqǏwqH��(���BJ������n��ts'���������!pU6�v�&�7��rď�v���w���+��B:�h�$�vǏ�v���W�*UǛ����ryV�v�F����%�ě����ry�v����*�ě�%��ry֑v�Ƒ��*ě�eĝ������� Û����f���<+��s��Cs��Ks��ss��{s��cs>��*�F����%�Ƒe���-���M����6�%�֒��u�����v������֓Ɩ�U�V����%�Ɛeǆ����=���M䜛i����Ξ�r�
�s���r���}5����oÞlf��r*��m1
�w>��sL��Y5����BĚ #����� ���Z���r#��s�� U���r$/r��rk��p���<������;?�,r���W����0Ɩ�s���r�
rx.�x9��r?��g��r?���ߘ%����=���rÞ�r���r;��r���M���rÞ�sJ��b������s��4s���f���=���M��}���dÂ��$r���r��,r4��j��,rǏ�sV��+s��B�oÞ�n��<���n㜐BJ�U���r$s��rk��p�6�<���w�&�x<��r?֒g��r?֒v������>��*e����6�r�x�p��rď�p���r��Tp4��j��TpǏwpV����(K���4mÜq����mÛ���>�����r��s�sZ�sj�'s
��p*��p�WpJ�wpZ�7p���g?��sO��;���S��M���3��p��g7��r��
��l�$�mÞ���M�	��rĜ���rìsɞ�r�
�s��Ɋ����� Û����f���<;��s��Cs���l!/m1��W���v1��l6��y�r���r�<�r;�Q�� Q�Ku�������?F�i'��:���VB�g
��r��>F���l�� �˕�rÞ2:���������˞�����'�m��?���W��?
�iˎ�4��}Vr�g��r�}>
���`WN�x�r���g���6���r��s>h�*?�����n������r;����(y
��l�
Oux>�x9��r?��g��r?��v���i���n���s7��n�ѬsV��i��$i�ܬsx��vӾ�x<��r?�g��r?�v��i���n��@s7��n��DsVJ�i��$i��Dsx6�v�&�x<��r?֒g��r?֒v��������s��B:��oÞ�n˝�<���n˝�B��ϛ����0���(���B���oÞ�nK��<���nK��BZ��ϛ����0���(k��B
��oÞ�n+��<���n+��Bʚ�˝���Uƕ�rÞ����r;��Ǜ���
?y�	�sǏq���r��$q4��j��$qǏ�v>N�f ��ry�vӆ��~�?;��s��Ks���4���=���M����6�%�֒��u�����v������֓Ɩ�U�V����%�Ɛeǆ�m�Du>F����
Ku`��j��s�DB>F�� Q�su�� �˕�rÞ����W~�q���JW��w���s4��f���s /m1��W���v1��6��y�r?��i���j���r0�������$m5��Ї������r�sV��I9��:��<��s:��`��r;��s�$�rÞ�?��s���d?��˧�-`���2��/m?��2���d8��r���j�4�r�z�s9��+��b������nǦ�#E��v��y;��'�r6�,r4!�n��,r���kÞ�r(��rÞ�,�-r:��/������� Ξ�r���s>D�h;��e���o*��e���*���Ǚ�����ɷ�#c����
�s���r��c#�����s1��d��s�~%mÞ�r�����m5��sXj�1��i;�:dÝs����r��a3��r%��m?��p�`Ǿ�s��`��kc���.Þ�p�`Ǿ�s��`���c���mÞ���M~��2��*m7��2���y�rǾ�s��rĝ����r7����=���M䜛g����Ξ�r�
�s���r���0��Þfi��r��s���Þ����M���3��p^�g7��r���^����p�`Ǿ�s��`��Ib���r�i-m'�r��w�ìsƾ�s��rĝ����r7��n���������Ξ�r�
�s��%m?��gy��r��m��w�ìsƾ�s��rĝ����r7��n�����=���M䜛a�����lΞ�r�
�s�#gB�� ���$m����3�wx=��rW��s��rÞ�r3���z��rR��1Ξ�r�
�s��r��sɞ�r�
�s`(�j�kB
kBǜȲ��Ɇ��r�Ds���r�
�s��Ɏ��r�Ls���r�
�s��ɚ���rÞÛ����f���<3��s��Cs��Ks��ss��͝2��ƻ��'Û����ϟ�lÞ���M�5*�jÞx=��rW��I����t����h��Ɇ���x=��rW��s<#m;��sF�B��>�����oÞ���Mv�x6��rT��w��ps4��f���r#��s��Gs��Os��ws q�r6
gB'-�w���m���r�
�s�.�&���rL��rÞ �|h�����#mìsH��J�y�rÞ �|?�w��rĜȊ��Ɏ��r�Ls���r�
�s��ɚ���rÞÛ����f���<3��s��Cs��Ks��ss���l!/m1��W���v1��(��y�rW��|�m6
oB'��w��ܛoÞ���Mi#���#��lÞ���M�a,�j��s
�s���r�
�s�7�眐s�#���Ξ�r�
�s��r��sV�^��>�����lÞ���MF��>�����oÞ���Mz�q���JW��w��Ls4��f���r#��s��Gs��Os���o/�:�� ���=m���,��~��JBɞ�rÕ�rÞ�lÞ���M�a.�b��s
�sǜ�����.�)����nG��lÞ���M�a1�j��s
�sǜ���� x�rW��I�����S����h��Ɇ���rÞ �|����M���3��pF�g7��r���^��F����!4�r6
oB'0�w� ���nÞ�y=��rW��s<8m;�Q�� Q���<S���(���C���Û�A�����rÕ�rÞ �|?�l��rR��1W��v��r 4�r6
oB'5�w�\���mÞ�y=��rW��s<8m;�Q�� Q���<S���(���C���Û�������rÕ�rÞ �|?�l��rR��1W��v��r 4�r6
oB'7�w�����dÞ�y=��rW��s<8m;�Q�� Q���<S���(���C���Û�`��7���rÕ�rÞ�mÞ�y�rΞ�rÕ�rß�lÞ���M�a9���s
�sǜ����:�� ���6m����/��y?��rΞ�rÕ�rÞ�mÞ�y�rΜ�rÕ�rÞ �|?�j��rR��1W��v��r 4�r6
oB';�w�����mÞ�y=��rW��s<3m;�Q�� Q���<S���(���C���Û�1�����rÕ�rÞ �|?�g��rR��1W��v��r 4�r6
oB'<�w�����V��s9��+�����j���"�?����j���r6�����s���V��s9��+�����j����?����j���r6�����s��l>��:����>�r.�<r�r��r��a��m���j���r6F��Þ�n��j���r66��Õ�rÞ Q��m;��r8��rÞ����rÕ�rÞ �|?gb��r��d8��r�񖗪yv��Y,:5 �nÞ���oÞ���Mg\��r��m8��rÞ�a>��:��=>�r;��r|�i��l���V���r��ak�mΞ�r�
�s`�j�kB
kBM�m=���G������=O��aW���0'E�r
Bx>�x<��r?��g��r?��v����O�%����m�>�����r��s����r�
B`�j��s
�sM�m8��rÞ�`W�x�r��4��2�Þ�������О�yÞ�r4�n��B�śr��O���� �
B4�f�� ��B�6�����O��0���=O�� W��>��#����Ɇ����� Û����f���<9��s��Cs���r=� x�rW��I����x=��rW��ìsH��J��S�����M���3��pF�g7��r���^��F���=���M䜛c�����T��w���s���r�
�s���rÞ �|�2��m3����,r /m1��W���v1��!+��y=��rW��s��rÞ �|?gU��r��d8��r�񖗪yv��Y,:5 �nÞ�y�rΞ�rÕ�rÞ�mÞ�y<��rW��s�m/��p�`Ǿ�s��`�����2���rÞ �|�����9��#E��v��y-��'�l?��rÞ �|(�О��S��mÞ�n��<���n�#��=��8��*���W��mÞ�'��r6mT��K����ЛlÞ�n��<���n��s���M���3��p��g7��r���^�8��l!_�r=���3���V��<>���,/r>��fP��rJ��3�҆���s7�j�Ѭs���^���,r���Õ�rÞ�r3���z��rR��1Ξ�r�
�s4(�j���dΞ�r�m���Õ�rÞ����<���r��,r4��j��,r���sƾ�s��rĝ����r7��n�����,r��mÞ��V��l����%���S��lÞ�n��<���n�#��=��8���%���V�Ç�b��I
�y�rΟ��<&m7�Q�ڛmÞ����$���6��mÞ��W��<���r��,r4��j��,r���sƾ�s��rĝ����r7��n�����,r��mÞ��V��l!�r=��y�rW��5�nÞ�p�`Ǿ�s��`���=�mÞ���M.W��W
�x4��r?��g��r?�����v��s	�����Ξ�r�9�sɞ�rÕ�rÞ�Þ�dM��r��y�r5�n���&���W��eÞ�n��<���n�#��=��8��$��dO��r��mÞ�y=��r5�j���&���W��kÞ�n��<���n�#��=��8���$��dO��r��mÞ�y�r5�j���&���W��dÞ�n��<���n�#��=��8��$��dO��r��mÞ�y6��r5�j���&���W��fÞ�n��<���n�#��=��8��F'��dO��r��mÞ�y<��r5�j���&���W��hÞ�n��<���n�#��=��8���'��y=��rW��$��w����2��m?���;��r��m�rK�"-��,r7�n���s'�^�;��rߒ�sa��<?��s���2��i���d���rÂ�0��mÞ�;��r���&���W��nÞ�n��<���n�#��=��8��y&��y=��rW��$�w����mÞ�dE��r��~�v�r?��B&��r:��;��r��lÞ�dE��r�����W
�x>��r?��g��r?�����v��s	��������r�
�s���r����&��n��j���r66��Õ�rÞ��Ҟ�y,��rW��gs��r��~�v�r9��&��r�s9��:����>�yß�r��mÕ�mÞ Q��<m3��r:��;��r���&���W��jÞ�n��<���n�#��=��8��&��n������6��m=��y�rW��I��y��73�mq��i��"��� ��2�s�r9��r�������s4�b���sǏsH��(Ӝ�BZ�Ѫ�� {��*�؄p)�"���4s���nÒ�Ɩ�p>֒gG��r?֒v����>�*�ƛ�e���q)�"U��p&���,�p>���;��rΞ�rç�u�����m3��ƛ��Ɲ������ Û�#��f���<?��s����>�-���M�����ƒ��&���֒�f�u���e�V����=���M䜛����kΞ�r�
�s�#B�� �Е�rÞ�2���r;��2�>����#��2��<�ܛmÞ���M�>��#��r�h'mĜȲ��Ɋ����� Û����f���<;��s��Cs���7���[��lÞ�n��<���n�#��=��8��#��y=��rW��s��r�&�r!��r�&�w���s'�n��(���#��2���y�rW��I����Þf%Û�������M���3��pJ�g7��r���^��F�m2��r�&�y�r������2��m?��2������2��mm?��2����� �Е�rÞ�2���r;��2�>����#��2�����lÞ���M.��='W�r,��rÞÇ��!��Þ�cϟ Ç��!}eÞ�n������9��7Ξ�r�
�s��r��sHa�w�ìs�Dsƾ�s��rĝȆ���r7��j����J�������cϞÇ��!}eÞ�y�rW��I����y�������M���3��pJ�g7��r���^��F�m6�,r4�n��,r���7���[��iÞ�n��<���n�#��=��8���"��Þ�����r?�߲���rÞҲ���s'��������<?��s���Ξ�r�
�s����� Û�#��f���#��7���[��hÞ�n��<���n�#��=��8���Þ�����r?�ߖ���rÞ �|h��Ɇ��r�ps����	���r'�ɲ�(�sF�~�q���JW��w��Hs4��f���r#��s��Gs��Os���7���[��kÞ�n��<���n�#��=��8��7��Þ�����r?�߲��rܬs����	���r'������r#��s���lÞ�n���(�y=��pV:�o��Þf���rĝ����r;����7x�rW��I��y����lW��i_�"���,i��l���n��B✒s���M���3��p��g7��r���^�;;�,r�s��k5��rÞ�n����r8��rÞ�<���r��,r4��j��,r���sƾ�s��rĝ����r7��n�����,r���#E��v��y.��'7�r��rÞ �|h�����im�@sƾ�s��rĝȲ���r7��h����J�m8��rÞ����r�
�s���s
�s4b�n�� ���rÞ �ސ���m8��rÞ�Ξ�rÕ�rÞ��М}lÞ�b��
c��rΞ�r�
7Bl��rÞ ��#���,q�6�lÕ�rÞ ��#��,q�6�o�Ɯs�nÞ��k�9��r���r�
7Bl�4B'e�/�����jm|��i#����������8Q���<S��n������y�rW��I�����S�����M���3��p^�g7��r���^����d8��r�� ����~�m�����r�
�s���r���"�i��j���r66��Õ�rÞ���Ds
Gs'��n���Ɨ��oÞ���Mi���ƃ������s
�sV��g���r
�s���r�
�s�7?;��s��Cs���k5��rÞ�y�rW��I����t�����M���3��p^�g7��r���^����r=�=���M䜛������?��h;��e��4mc��lÞ����� ����r?J�9WJ�x�rW��?^�9W^������ �
�s4i��� ����rÞ �ސ����^��F�m#��rÞ �|�M���3��p��g7��r��p�`Ǿ�s���`��������� ��2��m?�ɲ����� Û�#��f���<?��s���2��=���M䜛�������fI��r�?B	��m.��rÞ �|�Ђ�r�=�m�� �Ђ����n������n���w��&��8B���2����s��x=��r?2�r+j�r;
?Bޝ�r�8Bɞ�r�
�s��cm;�ɲ����� Û�#��f���<?��s���#E��v��y*��'��l:��rÞ �|(%О��{��mÞ�n��<���n�#��=��8��(��y�r4l�n�$/rɟ�r��}m;�����,r�� ����s
�sɟ�r��|m;���#�����7#��
Ξ�rÕ�rß� �
r`q�bÕ�rÞF�S������=S��:Ξ�rÕ�rß����� ��2�
r>��g9��r?��r�����>П�8?�,r��dΞ�r�#r���mÞ�n�9В�v�����r2
�sVҝ�$��w���� 	�
�C��ym�����n��6��,B>"���9�|��� ��xm/���#�	�
�C�7#��TV���9�|�(��hÞ�n��<���n��B	�
�C���s
�s`u�n��s
�sV����/qj
�s�	rǏ�s���r��s4��j��sǏsV֝}V"�}�
/B�R,��������rÞ�*���r;��*���5�
�C�
+B�R-Ў[23��B*��oÞ�n;��<���n;��Bʝ<S�����r�/r�sJ�sj�'s
��p:��p���d?�����
�қmÞ���M�>��#����Ɇ����� Û����f���<9��s��Cs ��r
'B���r��,r4��j��,rb��s�����,r&��r$��rÞ ����C���r�
�s��zm3��Ξ�r���sVƝy=��s^��������|�Û�F���W����|�(��hÞ�n��<���n��B	�
�C���s
�s`w�n��s
�sV����/qj
�s�	rǏ�s���r��s4��j��sǏsb�r��;7��s��s�sZ��cW�'���rû����y�rW��I�����S�����M���3��p^�g7��r���^����d8��r����#r���l�����C���aW���0'��r��rÞ �|h����
r�@sƾ�s��rĝȲ���r7��h����J�mm��rÞ�2���r;��2��ry>�v���x=��rW��y.�vӞ�p�^�q���JW��w���s4��f���r#��s��2���m���5�� %Е�rÞ�2���r;��2�>����#��2��c ���mÞ����2��wm7��2���v���8��Ξ�r�
?B>Ɲx=��rW��5t�bÞ�y�r?�����lǫ��3���� 	�
�C���r���G�����ޓ�;��Мq-�x�mÚ�v���8��\V����|�(��hÞ�n��<���n��B	�
�C���s
�s`w�n��s
�sV����/qj
�s�	rǏ�s���r��s4��j��sǏsV����MӤ��r�	?rǏ7s���r��$s4��j��$sǏ�p:���+�smď�p���r��p4��j��pǏ�pb�r��;%��s��s�sZ�7sz��p*��pʝ�p�� ��(�<��W&��r��rÞ �|h����
r�@sƾ�s��rĝȲ���r7��h����J�m8��rÞ�j$��/S��l���d?���3�x�� ����r���:��y�rW��I�����S�����M���3��p^�g7��r���^���>x>��r?��g��r?���>�*����=���rÞ �|%����m�������� Û�#��f���<?��s���h���=������W&�x9��r?��g��r?�����v��s	��"���Ξ�r�
�s��r��s���r�
�s��ɲ��r�Ds���r�
�s���rÞ �|�������w��Hs�psƾ�s��rĝȒ���r7��`����J��B��z����W&�x8��r?��g��r?�����v��s	�����Ξ�r�
�s��r��s���r�
�s��ɲ��r�@s���r�
�s��Ɋ��r�Hs���r�
�s���rÞ �|�lÞ���Mӡ��rĜȒ��ɖ��r�ts���r�
�s��������� Û����f���</��s��Cs��Ks��ss��{s���G
���{��jÞ�n��<���n�#��=��8�����y�r$v�n�����n��9ǖ�C	��m,��rÞ �|�Û�\�����r�
�s�xe��C�x/r���r�Ґu*��2��d������r�
�s�xe��C�x/r���r�Ґu*��2���rѕ�rÞ �|h������rÞ �|���h��Ɇ���rÞ �|���h��*-���Ck��Û�m��ry>�vӾ�e+�4��z�w���>�*��������Ck&�Û�5��ry��v���x=��rW��?B�9WB�Ө��rR��1WB�x=��rW��-�6Q��}���e�������� Û����f���<1��s��Cs��Ks��ss��2���m��������&�5���e���5�� %Е�rÞ�2���r;��2�>����#��2���=��mÞ���M�>��#��oÞ���M^��>�����lÞ���Mx<��rW���@s`@�nÛ�������M���3��p~�g7��r���^��F��~����5�� %Е�rÞ�2���r;��2�>����#��2��M<�	�mÞ���M�>��#��lÞ���M^��>�����nÞ���Mq'��rÞ �|����w��Ds�Lsƾ�s��rĝȎ���r7��f����J��B����5�� %Е�rÞ�2���r;��2�>����#��2��z>=�lÞ���M.7��aW�J��='��rm��rÞ �|h�����rK�"-��,r7�n�ìs�@s'��B�q���JW��w��Ds4��f���r#��s��Gs���2��>�� a���r����>x�rW��I����7c�mq��i���������������Ɏ����� Û����f���<5��s��Cs��Ks	�����aW�p��='��r��rÞ �|h������r���J�q���JW��w�ìs4��f���r#��s��͝���7���Û���&Ξ�r�
�s��r��s���r�9�s7E�n�ìs�@s'��B�q���JW��w��Ds4��f���r#��s��Gs��͝���7���Û����&Ξ�r�
�s��r��s���r�9�s7E�n�ìs�@s'��B�q���JW��w��Ds4��f���r#��s��Gs���l!��r
'B���r��,r4��j��,rb��s�����,r&%�r���rÞ �|h������rÞ �|���h��Ɇ���rÞ �|�Ʃ�C���r�
�s���p�r�x<��rW�����y=��rW��aD�Û�������M���3��pB�g7��r���^��F��~����W&�x6��r?��g��r?�����v��s	��:��Ξ�r�
�s��r��s���r�
�s��ɲ��r�@s���r�
�s��Ɋ��r�ps���r�
�s���rÞ �|����lÞ���Mx<��rW���Hs`G�jÛ�������M���3��pr�g7��r���^��F��~��v��n����W&�x1��r?��g��r?�����v��s	�����Ξ�r�
�s��r��s���r�
�s��ɲ��r�@s���r�
�s��Ɋ��r�ps���r�
�s���rÞ �|����lÞ���Mx<��rW���Hs`F�jÛ�������M���3��pr�g7��r���^��F��~��v��n����W&�x0��r?��g��r?�����v��s	��G���Ξ�r�
�s��r��s���r�
�s��ɲ��r�@s���r�
�s��Ɋ��r�Hs���r�
�s���rÞ �|�lÞ���MӚ��rĜȒ��ɚ����� Û����f���<3��s��Cs��Ks��ss���G
���{��bÞ�n��<���n�#��=��8���dx�rW��I����x=��rW��ìsH��J�x<��rW���DsH��B�x?��rW�����r�
�s���rÞ �|����w��Ls�tsƾ�s��rĝȖ���r7��b����J��B��z����5�� %Е�rÞ�2���r;��2�>����#��2���:�U�mÞ���M�>�����mÞ�y?��r?6�s���r����;�r.��mÞ��k�9s��r���r�
7Bl��rÞ ��#��,q�6�o�Ɯs=��nÞ��k�9ik����#�s>^���)���s`g�f��s>6��W��v��Ds�Lsƾ�s��rĝȎ���r7��f����J��B����5�� %Е�rÞ�2���r;��2�>����#��2���5�#�oÞ�n��<���y�rΟ�r��,r���r�
�s���s4�����s���j��iÏ�o	��2���m(��rÞ��
�C�ᐦ��C���W���ÏM��0'O�r*�rĝ��
�sV���5M�j���s�����C���<���r��,r4��j��,r���sƾ�s��rĝ����r7��n�����,r���#E��v��y%��'��r-]m�ᐦ���r�HyО�d���r���mÞ��ό�Ü|l�N�:Þ�rh��rÞ��Þ�y?��rΞ�rÕ�rÞ�mÞlx=��rW��?��9W��Ӓ��rR��1W��x=��rW��-�6Q�
�CHL�-���#��Ξ�r�
�CHL�-���r.
�CHL�-���yß�r���4��mÞ��ό��!|Þ�y=��rW�����r��rĝ����r7��������Ξ�r���sHP�~=��s^�����
3��r?������!amÒ�v�������2�r��r�s�2���r�
�s�xe�C�� 	�Ymh�r6�r�vXm=��g?��s@Z���n�QЖ�rp��rÞ �|����w���s'��y��?���3��j���r0�������,m5����O.Þ�m���s�����8��k5��rÞ�~�
�CHL�-���r��rÞ�mÞ��眚mÞ���M�W�����/�+�����6�ǛlÞ���MӤ��rו�rÞ �|�>�
�CHL�-���r
�Cǜ%-�����r>��:��<��s:��`��r;��4��������8��jW���������r�
WCHL�-���r8��rÞ�d�~�r�[C���mÞ�Ə��ќ}l���m��r.
KC�
WCHL�-���M���1�� ��]mm�rWB�A���G���ъ����
Ξ�r�
WCHL�-���Ɵ����၂��@C�l�r2��rC��-Ξ�r�
CCz�-aU�n��sz�x�r?~�����lǫ�lÞ�W�������!a��Zm/��r5�@C>F�r<��Þf)Â����DC4W�jÞ�ƛ��lǫ�����y^�UÞf�ÊX��
CC�ᐦׁ����n���џ�r5��rÞ�Þ�rHWmĜ��Vm$�sɞ�rÕ/mÞ��-r->�2��Vm3��2���m�Pmy.�vӾ�?���3��j���r0�������,m5����O.Þ�m���s�����;;��s��s��k5��rÞ�Ɵ���H�ў����k5��rÞ�Ƌ���!a��Pm?��r2��rÞ ��]mo�r�ћlÞ���M�������r�
�s��Rm��x=��rW��$_�w@�����y=��rW����/ c��25^�n��pC���mÞ�y�r?J�s�������Þ�y�r?������lǫ�ɯ��0���b���nߌ	�Ymh�r�ᐦ�	?r�C/��?��q��,x=��rW��-�s�2?��q
�sHP�-���-k��p���lÞ�nߌ��O��0����{C���#E��v��y$��'z/m-]m�ᐦ���r�HyО�y�rW��h����\m��r��lÞ��ό��!|Þ�~�
�CHL�-���r3�r�
�CHL�-���r(��rÞ �|�>W�����/�;��Ξ�r�
�s�
�CHL�-�q�r���oÞ���M�ό��!��Þ�;W��v�$/r�sW��i;��e���o*��e���2���j���g��l?��s���2���d���r�ћmÞ�y�rW����/ c��24��j���sz��#��Û�#��� ��y�rW����/ c��25^�n��pC���kÞ�rh��rÞ��Þ�y>��rΞ�rÕ�rÞ�mÞ,x�rW��?��9W��Ӓ��rR��1W��x�rW��-�6Q�
�CHL�-���#��W�����/�+��rß�'�,m2��rÞ y�]mo�r���mÞ���Mx��rT��w���s4��f���s���r=��y�r?������lǫ��[�-���b���nߌ	�Ymh�r�ᐦ�	?r�'CS��?��q��,x�rW��-�s�2?��q
�sHP�-���-k��p���lÞ�nߌ��{��2����C/��Ξ�r�
�s����� Û�#��f���#��#E��v��y'��'�.m;�m'�/m%�mǾ�s��rĝ����r7��������$��v���JW��w���s4��f���s���kÞ�r���s��"-��,r���r�
�sz�-v.�e��rÞ �|�Û�q�>�i���������J��� ß�r���rÞ ��(C-�p:ޛkÞ���M.��=Ɩ�s>��gG��r"�i㜒s���������rÞ �|�oÞ���M�3��p��x=��rW��Ξ�r�
�s��m'��h����J�;7�r��s�s��k5��rÞ�p��M���3��p��g7��r��p�`Ǿ�s���`��/�#�hÞ�n��<���y�rΟ�r��,rɞ�r�
�s���s4�����s���j��i��o	��2���m�rؕ�rÞ �|?x<��rW��s��rÞ �|?i��2��m+��2��=���M䜛��S"�k5��rÞ�d���r���Þ�r.��rÞ��<�mÞ���8)=� ��$r���r��,r4��j��,rǏ�sV��h��/�;��0���(ß�B✚hÞ�nK��<���nK��BZ�	��mh�rĜ����r?�*����%���rÞ�:���r;��:����
�s9��-9��g���r^�f��ry�vӖ�x9��r?��g��r?��v�V�����!aa�<�m?��sJ�f��ryv�v��x9��r?�g��r?�v�6�����!���m?�Ɋ���r?�*5ƛ�ƕ�rÞ�z���r;��zƛ�U�
�s9��-������rĜȎ���r?�*�Ǜ��Ǖ�rÞ�����r;���Ǜ�%�
�s9��-���w��Ls7��n�$�vǏ�vb�r���^��F��~�;�,r��s�sZ�7sz��p*��pʝ�p��wpJ�pj��q*��q�Wq��qz��v:��d?����L/�� ������ Û�#��f���#��#E��v��y ��'K+m�rĝ����rÞ �|�mÞ���Mi�����#��2��=���M䜛���"�T��w�ìs���r�9kB���r�9�s'��/#����m3��n�����=���M䜛���$�gΞ�r�
�s�#�@�� 9��=m���.~��y=��rW����/�)���s`��j��sz��眐s�#��y������Û�B%����r�
�sz�-$��/#���<�m;�Q��pCV��v��r��$�aW҂o��='\*m��rÞ ��pC��r|��i#�^������
�sǜ�����s �*m6
�@'5�w��(�͛lÞ���ݖ����#�s>�����rR�� ��Q���<S�����(�� 9��:m���y��y<��rW�����r�
�s�<�m;��s�m=�Jx�rW��I����x=��rW��ìsH��J��S����h��*m���s�"-��,r���r�
�sz�-v.�e��rÞ �|��Û�q�>�i������������M�������� Û����f���<7��s��Cs��Ks���d�>�-���=���p�`Ǿ�s���`���+��Ç�nÞ���M����r�
�s�.�lÞ���M�Ξ�r�
�s��,r4����,r /m1��W���v1��9z�)x<��r?��g��rΞ�rÕ�rß�2���rÞ �|����r/�����j#9�s>ނr<��r��s���mÞ���2��wm7��2���q���9��Ξ�r���sVނy=��s^ʂz����-�|�Û�7)�j$��/������r��,r4��j��r=��y�rΟ�r��,rV����Mi��h���n��ß�r�s�2���Þ����r<��j���=���M������Û�7)�G���r��,r4��jÕ�rÞ�����r;� ��$�s>�m�śmÞ�yß�r>����-�|����r/����]m���wӾ�x9��r?�g��r?�v��Ӝ�r��rÞ�rß�ik�	�
/C��$s4����$s�L�p=��B*��hÞ�n;��<���n;��Bʝ�$�pǏ�p���r��Tp4��j��TpǏwpb�r��2���m�����6�%��5���e���U�V��ƞ�r5��sXʂ�x���S��M���3��p��g7��r��p�`Ǿ�s�Ð`��d$� ����r?����rìs'��g/��rJ�B�q���JW��w��Ds4��f���r#��s��Gs���#E��v��y��'�&m*��rÞ �|���,r4$�f��,r���lÞ���M,��2��*m7��2���y�rǾ�s��rĝ����r7����=���M䜛��S*�cI��y�r���u��~����M���3��p��g7��r���^�T*�l��ÇU�y=��rW��ơ�m���T�4�m�z�s9��+��f������a>����=��r�s9�����ú�y?��rΞ�rÕ�rÞ�mÞ�y�rΟ�r�
�s49����0?��i������r6����s1v����s������r�
�s���G���T�±m6b�V���s���V��s9��+�����j���"�?��眛��T�oÞ���Mq'�X:>�����ú����+?b�h��W��dm��V��s9��+�����j���"�?��眛o�T�В�G�O�i��W��m�����%i���T�±m6�V��s>��h(�����r*����tm`�Q���G�kB�������T�±m6�V���s���mÞ���Mh��W��8m�����r�
�s��m��c������s1�Q���s�1�����n��S���n��B��"���wӞ�73��mď�s���s9����n<��s:��`���m�����j���=���M���s��c��i��W��\o����p^�q���JW��w���s4��f���r#��s���#E��v��y��'�#m6�mT��K���!���T�4�m�z�s9��+��b������dΞ�r��m���mÞ�v���JW��w���s4��f���s���#E��v��y��'r"m6�mT��K�� �D���m��c?�����s1~�L�
�s'��y��i��S���n��B�����wӾ�x=��rW��y.�v��73��mďsɞ�r�
�s�$�sǏ7sƒL�%�����m��c?�����s1B�L���r#��s�����;3��s��s�sZ�7sz��#E��v��y��'k<m(��rÞ �|?i#�H���������r���sVs^���p�=���!�=��m��f��r^��#�	�
�@}��lx��y�r^�+��������Û�<?��s���2��� ��mĝ���#�� 	�
�@}��l��#��0���=���
�sV��,9��+?� ��<pm?��s�??��s���IV�+c��oÞ�n��<���n��B�	�
�@}��l��#��0���=���
�sV��,9��+?� ����r?�*m���M���rÞ�����r;��������
�sV��,���qU.�v�6�x9��r?&�g��r?&�v�֒���!aÝ������rÞ�j���r;��j���u�
�@x��vӶ���??��s������=���M����6�%�֒��u���m5��sX���v��y�rW��I�����S�����M���3��p^�g7��r���^���=���M䜛���3�?��h(�����r*�?��;�@>�s��K��<m��@]��������x:��rW�������,r&�<m(
�@�z�s9��+��������jƭ�@6.�l���bќ`eф�p�,x=��rW��y>�?��h(�����r*���/r��rƓ�m*��e���rÞ�?��s���2���y<��rW���˓�c��n������r6����s��m���s�țnÞ���Mq'"r�s9��+�����j������������s_��x>��rW��$��w������s4�b���s�4�uҜ�n������r6����s��m���s������=���}��9qX�����hÞ���M.��=Ɩr>��gG��r?��qh��}������r��a#��r;��;��r%��;5�r��s�s�3���-���rÞ �|�Û�q�>�iß�����nß��Ɩ�s�s9��+�����j���h������d�>�-���m���ml�=�/r���r�
�s���r�Γub��r��m3��r��5pʎ�?��h(�����r*�����r�����rc�/r��sҜ�	���rÂ+�������r��a#��r;�� ��r%��m��rÞ�)c��n������r6����s��m���s�������	��m���
���	��m����ƞ�	?��h(�����r*����Oj���i���s�?����r��a#��r���r��,r4k�jÕ�rÞ�R��am;��2��rݞ�B��"���wӞ�i㜐BJ�����J������d���=���M��m��rÞ�rß�7c��mq��i��mÞ���Mi��h���n��;;�7Q���@���n���=���y�r?���?��lǫ��Ǎl���>���c��n������r6����s��m���s������r��a#��rW���?�M����`ڞ�r%��m8��rÞ�d?���Ǎ��������r��a#��r;��s���lÞ����k5��rÞ�n������r6����s]������^�q���JW��w���s4��f���r#��s$��8��#E��v��y��'t;m2�,r7�nÇ���,r������ ��2��m?�����mìsV.�IΟ��#��n�����,r�� �Ђ����n������n�<ˍ�2����s��x=��r?��x�r��jW.�I���fW����=ˍ�W��q���JW��w���s4��f���s /m1��W���v1��&n��4c�mq��i������#��D��*=��m?�����r��s���2��m?���s��2���4c�mq��i������#��D��ɲ�
?Bޒ�sa��<?��s���2���y�rW��W.�I��m7��jW.�I���Ξ�rÚ��� Û�#��f���#��#E��v��y��'[5m5��rÞyў�rb�mÞ E��@s
Cs��r�
�@>��9W���ύ�fԞ�rSD�1W��i����W^��׍$m�
Cs>F�qj
GsV��*Þ�Ї}���r#��s��Gs�� }њ9�4�W��ύ�s��y��x<��r?��g��r?��vӞ��׍(��
�s7��n��@sV^��׍$m��@sx��v��7c��mďsV��.������r?�ߎ�
GsV��*ÞҎ�$7sǏ's���r���p4��j���pǏ�pb�r���^����r�/r�sJ�sj�'s
��p�� yѕ�rÞF�ύ͛i��r>�r����i!:m%
rƾ�s��rĝ����r7����=���M䜛 ��'6�I���3���I��y�r���qh��ў�M���3��p��g7��r��m<��l��@��rا@�rÞ��'�4m0�mΞ�rÛ�7�Ϟ��Е�rÞ�f?���О<gs��r�<i��j���r66��Õ�rÞ Q���mÞ���y�rΞ�rÕ�rÞ�B���s
�s`���kB
kBǜ��О����~��JBɞ�r�
�s���K���r��ms<?m3�Q�� Q��9�7�Ϟ��Е�rÞ�??���О<gs��r���3���֞�wk��r5��rÞ@�y�rơ�m���l��B��� Û�#��f���#��#E��v��y��'f7m6�mT��K��i����mD�x�r���r��ms�<m3��r4��rÞ��О�dΞ�r��m���mÞ�v���JW��w���s4��f���s���#E��v��y��'�7m6�mT��K�������mÞ���M�3��p��f͞�r^�??��s���l!/m1��W���v1��*j�Þf���r$�s����,�s>��7s��rq��i��r�ikmϟ�p�>�iß�����nß�BJ��s���M���3��p��g7��r���^�;7�r��s��sJ��#E��v��y��'�6m-��rÞ �|�rÝ~�Þ�y=��rW���7�r�lkm�ޛoÞ�n��<���y�rΟ�r��,r���C�����r/�����j#9�s9��s<��r��s���mÞ���MϞ�2��*m7��2���y=��rW��$��n��(���9��Ξ�rÚ��� Û�#��f���#��#E��v��y��'�6m�mÞɲ����� Û�#��f���<?��s���#E��v��y��'�1m6�m$��w�����Û�p���r0��rÞ �|?�ߍ�c���r�
�s�.Mў�y=��rW��|��m3
�@����ߍ�z���r6�mW��g˞�r��rD��r8���Ğ�$��v���JW��w���s4��f���s���V���r��ak�mW�����v���2;�l����Ú��� Û�#��f���#��l!/m1��W���v1���d���Ȟ�>T��G�����mE��r:��rơ�m���mÞ�v���JW��w���s4��f���s���#E��v��y��'�2m��rÞ�rß�7c��rq��i��mÞ���Mi��h���n��;;�7Q���@���n���=���y�r?���?��lǫ���W��� 	�
�@���r����f�ux<��r?��g��r>�m�śmÞ�yß�r>����i�|����r/����]����v���rÞ�r���r;��b���	Ξ�rÕ�rß�r�
�sVₓ?��g9��r?��s��lÝ���s���q��������r��s�sJ�s�� ]��@�S@�=�f���r��,r4��jÕ�rÞ�����r;��oÞ�n;��<����S�%��r�y�rΟ�r��,rV���?�Mi��h���n��ß�rď�s��Û�����p=��y�rΟ�r��sV���?�Mik��h���nk��{��rď�p��Û���Dp<��y�rΟ�r���pV���?�Mi˝�h���n˝���rďWp&�Û����@�+%�ƛ��ƕ�rÞ�����r;���ƛ�5�>�����r��s�sZ�7sJ�'s
��pʝ�p�Wp��pZ�7p
��g?^�sOZ��g��r5��sX���d���S��M���3��p��g7��r��p�`Ǿ�s�֐`��9���mÞ���M�>�����lÞ���Mx�rW����s`��nÛ������h��Ɏ���rÞ �|����M���3��p~�g7��r���^��F��~���=���M䜛4���<�;���r�
�s���rÞ �|r���w�ìsƾ�s��rĝ����r7��n�����=���M䜛7���	�`Ξ�r�
�s�#W@�� �֕�rÞ�2���r;��2�>����#��2�������oÞ���Mx=��rW��s��r;��rĞ��Û�BĜ��um
rx>�iӘ�B��oÞ�n��<���n��B<S��h���=���m0
rt��oÞ��?�>Ξ�r�
�s��r��sV�J�q���JW��w�ìs4��f���r#��s���k5��rÞ��)����r4�w�[@8?�aW���0'�m��rÞ �|h����
r�@sƾ�s��rĝȲ���r7��h����J�m��rÞ�2���r;��2�������� Û�#��f���<?��s���2��C��� �֕�rÞ�2���r;��2�>����#��2��\����oÞ���Mx=��rW��s��m;��rĞ��Û�BĜ���m+�r�nӘ���rcрw	��m+�r=��nӘ���rc�\@	��mr
rV��y��x�r?��g��r?��vӞ����%����M���rÞ�����r;��������>�����r�/r�sJ�s�� ��(�<��W&�m��rÞ �|h����
r�@sƾ�s��rĝȲ���r7��h����J�m8��rÞ�j$��/S��l���BĜ��8m6
r'��w���қmÞ���M�>��#����Ɇ����� Û����f���<9��s��Cs�ЛiÞ�n��<���n��s���M���3��p��g7��r���^�8�́Z��Ƌ��hÞ�n��<���n�#��=��8���]�Ax�rW��I��F�i��"��L@���cÕ�rÞ���@s
Csɞ�rÕ�rÞ �|�nÞ���M��i���ƃ��lÞ���M�a����s
�sǜȎ��ɒ��r�ps���r�
�s��ɞ����� Û����f���<-��s��Cs��Ks��ss��{s Mm
W@���r��,r4��j��,rb��s�����,r&�	m���rÞ �|h��Ɇ���rÞ �|�nÞ���M��i���ƃ��lÞ���M�a��j��s
�sǜȊ��Ɏ��r�Ls���r�
�s��ɚ����� Û����f���<3��s��Cs��Ks��ss��́Z��Ƌ��jÞ�n��<���n�#��=��8��Y��y<��rW��|z�m�t@���lÕ�rÞ ����s
�s���r�
�s�.n�������#��֚7������s�� �֕�rÞ���7Ξ�r�
�s��r��sVr�v�ìs�Dsƾ�s��rĝȆ���r7��j����J������hÞ���M.���a���r�
�s�#c@�� ����m����_� x>��rWn�q'�JB���rÕ�rÞ�iÞ���Mi#���#���<�m+�Q�� ���rÞ �ސ�W��������(��� ����m���_�7���!������ ����rÞ�mÞ�y>��rW��?��9W�����h�������#��iÞ���/qj
�s>n�qj
�sMr�??��s���.Y��Ʒ��k�N� Ξ�rÕomÞ���-r:��2��Vm3��2��!�� B>f�r=�,r�� �֒�v�
g@�� ����r�H�֞>����֒�&Wf���/x?��rΞ�rÕ�rÞ �|��� �
w@`����s
�s���r�
�s�7 ��Q�{@���aWj�;�='�
mj
@t
@>^�9W^�x<��rΞ�rÕ�rÞ �|��� �
w@`����s
�s���r�
�s�7�����֚7������r#��s "m6
c@'��w�(��9��(���s
�s���rÕ�rÞ�iÞ���Mi#���#���<�m+�Q�� ���rÞ �ސ�W^�i����W������n������r���rÞ �|h����
{@ǜȲ��Ɇ��r�Ds���r�
�s��Ɏ��r�Ls���r�
�s��ɖ��r�ts���r�
�s��������� Û����f���</��s��Cs��Ks��ss��{s��́Z��Ƌ��eÞ�n��<���n�#��=��8��e[��y<��rW��|z�m�t@���cÕ�rÞ ����s
�s���r�
�s�.n�������#��֚7������s�� �֕�rÞ���7Ξ�r�
�s��r��sVr�v�ìs�Dsƾ�s��rĝȆ���r7��j����J������mÞ���M�>�����nÞ���Mi#���#���<�m;�Q�� ���rÞ �ސ�W��v��@s�DsH��B�x?��rW���psƾ�s��rĝȒ���r7��`����J��B��z��	�WV�x5��r?��g��r?�����v��s	��Q	�a��g4��r��me��m���+��#��2���m?���Xv؛����������m?��E?�Xv؛�������`�������r#��s��Gs���n���=��,x�r$���C��#��b��ɲ���rÞ �|����f��*-��)m;�����r#��s���2���d8��r�n�mÞ���M�>�����mÞ�yß�r���r���r$���C�����#�����w��@s�DsH��B�x�rΟ�rÕ�rÞ����mW�f��r~�v�q���JW��w��ps4��f���r#��s��Gs��Os��ws Mm
W@���r��,r4��j��,rb��s�����,r&Mm$��rÞ ��pC-r:��������l!/m1��W���v1���T� 7c�mq��i�����m;��������m?�ߎ���rÞ�rß�x=��r$��0��Ȳ���m�@s���+���������������r#��s��Gs���n���=���nG�"���,g���r�ɛmÞ���Mi#���#������6W��x�rW��-�6����d8��r�u�mÞ�y>��r?6�s���r����;�r�mÞ��k�9x�rW��-v.�e�|����nG�"��,q�6�o�Ɯs�nÞ��k�9��r���r�
7Bl�4B'e�/�����jm|��i#����������8Q���<S��n������d8��r����� ��2���s4��j���s���s7��n��Lsɞ�rÕ�rß�lÞ��Ғ�ìs'��J�Þf���r+�Ɋ���m������m?��f����J��B����r��s /m%��W���v1��T��W��+q1��W�7c�mq��i�����m;��������m?�ߚ���rÞ�rß�x=��r$��0��Ȳ���m�@s���+�������h��Ɏ���rÞ �|����M���3��p~�g7��r���^��F��~��v�;?�,r��#E��v��y ��'Omi�r(�"-��,r>��g2��rΞ�r���s.��m���rÞ �|%���M�؜s6�BJ��/���v��@��2���m�������y�rǾ�s��rĝ����r7����=����M䜛2���
�M䜛(����`���r�
�s�#@�ɛmÞ���Mi#���#������6W��x�rW��-�6����d8��r�{�mÞ�y>��r?6�s���r����;�r�mÞ��k�9x�rW��-v.�e�|����y=��rW��-v��e�|����
Ӝ�r���r�
7Bl��p�iÞ��k�9ik����#�s>^���)���s`g�f��s>6��W��v��r���^�m8��rÞ�`W�q��G��v���oÞ���M.��='�mV�s9��:����>�y=��r$��n���ƛ��nÞ���Mi���Ɨ����s
�s'f�n#���#�Q��gm+��ƃ���֚7����nÞ���/qj��r#��s��Gs��oÞ���Mp��='WmV�s9��:����>�y�r$��n���ƛ��nÞ���Mi���Ɨ����s
�s'f�n#���#�Q��gm+��ƃ���֚7����nÞ���/qj��r#��s��Gs�� ����m���S��y�r$���G��#��f��*-��)m;�����s	��m8��rÞ�T��KHP�-���~=��x=��r�@���mÞ��K� Ç��!�rÜ|l���fÞ�r��rÞ�rß�7c��rq��i�����s4�����s���j��iO��o	��2���m3
@�ᐦW��|�m[
@t��rÞBpU��x=��r?� c��2?��g=��rΞ�r���s���m�����s4y�f��s�� ���r�Ymh�r�gm���s��2���m���mz
@t��rÞBpU��x=��r?� c��2?��g=��r?������K� Ç��!am�!��?�����r��s���j�4�rǖ�s>��p��,�3�(��� ���r�Ymh�r6�r�v�m=� ����m�_�r%��m)���K� Ç��!am�!}eÞ�r#��rÞ �|�M���3��p��g7��r��m=�=���M䜛-���7Ξ�r���r���y�rW����s'��y��f���r^���=���^�8��>R�'J�h������rÞ �|���h��Ɇ���r���B�q���JW��w��Ds4��f���r#��s��Gs���o/��r��rÞ����r�����x�rW��ìs'��y��g|��rOr�??��s���2���d8��r�̛mÞ�y�rW��$����i�����n��9ǖ@��8��;����m�4���,r���֣��M��v_���֞�d"��r��y<��r$��Þf������rÞ �|������*-��)m;�����r#��s	��m8��rÞ����+��mÞ���M��!��(�����#��2��'J�h������rÞ �|���h��Ɇ���r���B�q���JW��w��Ds4��f���r#��s��Gs���o/��r �@k���rÞ �|%��=�-����Ξ�r���sW��KHP�-���~=��s^�L���� Ç��!am�!aiÕ�rÞ �|�='�m%��rÞ 	��r�Ymh�r�~iÞ�v_
�sW��KHP�-���-�f�r���d?���_������ǖ@����6�؛oÞ���r�h�r��sɞ�r�
�s��ɲ���m$/r4#�j�{B���^�8��k5��rÞ�ÞfÕ�rÞ �|�#����*-��m?����,r�)����r��sɞ�r�
�s��ɲ��r�@s���+�����M���3��pF�g7��r���^��F�������T��KHP�-���~=���c��`W>�x�r�������lÞ�n� Ç��!amÒ�v���֨m
�sW��KHP�-���-���y�rW�����O���� Ç��!am�!feã�O�-h;�:dÚ����s�s�2?��q��,�� Ç��!am�!7mÜw��������e���s���rV���3�����/�Þ/�;��i!�m=��n����m=��v_���֞��c��lÞ�R�m ��rÞ ���r�Ym��r�o�r%��rÞ�1Ξ�rÕ�rÞ �|������,r4y�f��,r�� ���r�Ymh�r�gm���s	��m!��rÞ �|���r�Ymh�r�~iÞ��K� Ç��!am�!feã�N�-h;�:dÚ����s�s�2T��.s���K� Ç��!am�!7mÜw��������e���s���"r
@W��KHP�-���-k��p���mÞ�~�
@W��KHP�-���-���rv��rI����x�rW��ìsH��J��K��sF�~�q���JW��w��Hs4��f���r#��s��Gs��Os /m1��W��.q1��I��y�r?���3�����/�Þ�lǫ��s����� 	��r�Ymh�rh�rΞ�r�
�s����� T��.c��y=��rW��-�s�2W���3�����/�Þ/�Þ����r���I��r5��sX.��I�=���M䜛/����bT��i;��e���k&��#E��v��y��'Bm ��rÞ���r�Ymh�r�ᐦ�'@��W���3�����/�Þ/�?��mÞ���Mv�{��� 	��r�Ymh�r6�r�v�mÞ�7W��v���sH��^�x�rW���Dsƾ�s��rĝȆ���r7��j����J������l����'@%�#E��v��yx��'~m4��r�����Ϟ�p^�q���JW��w���s4��f���r#��s���r=��y<��rW��$��w�)��)�r�h�r$����x�rW��ìs'��J�x=��rW���Ds''�n��(���<;��s��Cs���2������>Ξ�r�
�s���m��s���r�
�s��ɲ��%m?��gy��r���^�8��l���lĝȲ����� Û�#��f���<?��s���#E��v��y{��'�m��r�*�v�ìsƾ�s��rĝ����r7��n�����=���M䜛%���Ξ�r�
�s���Þ~!Þ�y�rW��$��n��(���9��Ξ�r�
�s����� Û�#��f���#��#E��v��yu��'�m��rÞ���s9��+�����j��4-���
c��r�z�s������,r�/@���W�+s����xn�s9��+�����j�����rÞ�r�!�s�B�oÞ�n��<���n㜐BJ�<S�����r��s�sJ��d?������/���r��s>��h(�����r*���/r&��rcìs�Dsƾ�s��rĝȆ���r7��j����J����s	��p�l���mÞ�yÞ�rT��w���s4��f���s���r/��2���6-2m<��rÞ�rÞ�rÄ�r���&Þ�r3f�l��l��l�
�l��l�&�l��l�҂l�V�l�j�lò�n��n��n�Z�n�R�n�J�nê�o�Z�o�b�o��o�6�o�&�o���$��s��8-Þ�rÞ�rÞ�rÞ�rÖ�$��s�;-Þ�rÞ�rÞ�rÞ�rî�d#��sÞ�rÞ�rÞ�rÞ�rÞ�r�F�$��s��8-Þ�rÞ�rÞ�rÞ�r��n#��s�ނh"��s���>���rß�l#n�l#��s���h"��s�)�r�;-Þ�rÞ�rÞ�rÞ�rÎ�o#��sÞ�n#��s�N�l#��sÆ�i#��sß����rß�����rß�E���rß�����rß�m�~�d#��sÞ�rÞ�rÞ�rÞ�rÞ�r�2�h"��sÞ�����rß�l#��i#��sß�r���r�l#Ɲh"��s�������rß�����rß����rß�u���rß����rß�l#^�o#��sî�n#��s��h"��s��̊���rß�m�J�h"��sÞ�N���rß����rß�����rß�����rß���)�rß��o��rÞ�rÞ�rÞ�rÞ�V���rß�U���rß�)���rß�mÞ�rÞ�rÞ�rÞ�rÞ����rß����rß�I���rß����rß��)�rß�o��rÞ�rÞ�rÞ�rÞ�V���rß�����rß����rß�M���rß�A���rß�����rß�����rß�����rß�mÞ�rÞ�4Þ�r�z�k�"�k���l�^�l�J�l�F�l�B�l�~�l�z�l�v�l�r�l�n�l�j�l��læ�nâ�n�Z�n�V�n�R�n�N�n���o���oÞ�oþ�o��o��o�6�o�&�o�֒o���o��oÖ�oö�o�V�o�v�o��o��o�6�o�֓o���oÖ�oö�o�V�o�v�o��o�&�o�Ɛo��oÆ�oæ�o�F�o�f�o��o�&�o�Ƒo��o�6�h�r���&���rÞ�r���'=r�R=P�x=��r�<���������+�n4mÉ�Dժ�����������|M����J;��J;��J;��J;��J;��rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�r���J;��rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�rÞ�r�    �G        ��  �   `  �   H  �   0  �    �G          �  �    �G          �  �    �G       1u   �2u    �3u  �  �    �G       e   x �f   ` �g   H �h   0 �    �G         �      �G           �      �G           �      �G           �      �G           �      �G         �      �G         �      �G                �G           0� �  �      � 0   �      8� (  �      `� �  �      H� 0  �      x� �  �      <� �  �      Tp ��  �      @E  n  �       C U S T O M   �4   V S _ V E R S I O N _ I N F O     ���                                         D     V a r F i l e I n f o     $    T r a n s l a t i o n     �8   S t r i n g F i l e I n f o      0 4 0 7 0 4 B 0   $   P r o d u c t N a m e     s   4   F i l e V e r s i o n     3 . 0 0 . 0 0 0 1   8   P r o d u c t V e r s i o n   3 . 0 0 . 0 0 0 1   , 
  I n t e r n a l N a m e   s t u b     @   O r i g i n a l F i l e n a m e   s t u b . s h a r k              0  1u     �  2u   (  3u(                �                         �  �   �� �   � � ��  ��� ���   �  �   �� �   � � ��  ���                             �w   ���wp ����p  ����   ����   ���    � �    ��    �                                     ��  ��  ��  �  �  �  �  �  �  �  �  �  ��  ��  ��  ��  (       @         �                        �  �   �� �   � � ��  ��� ���   �  �   �� �   � � ��  ���                                                                                                          ��p          ����wp      ������wwp    ��������wp     ��������p      ��������        ��������        ��������        ��������        ��������        ��������        ��������        ��������        ������          ����  ��        ��  ��            ��            ��                                                                                                                                           �������������������������� �� �  �  �  � �� �� �� �� �� �� �� �� �� �� �� ?�����?������������������������������(       @                                ��� ��������������������������<����?���������������������������������������������=������<?������?�������������������������������������������������������� �� �  �  �  � �� �� �� �� �� �� �� �� �� �� �� ?�����?������������������������������MZ�       PE  L             �                      @                     �                                       T  (                                                                                                                 .text   �      �                     �    T  (                                                                                                                 .text   �                           �                                                �  �  �      �3   �@�8 u���8 u�FVV�   ^��uÃ�u�jd�   ���%@ �% @ �%@ |          �                         �  �  �      S DeleteFileA � GetCommandLineA `Sleep kernel32.dll    x��gP���7�N � @� �E 4��R�.�H$� !���XP�����^��������g�g�3�ә9ΚY�e��Z+{�u]��ׇ8� �   ��[[ @�?B�?�p[%T�$ ��ݪ5@�nU���c�XVL(+0
80::&(�bG�ã�V.��Q1A�:��b����?�FU Nd�w}�����6�I�del�[������0� G ��h�_�	��*�l��* �  �: ������� ������?	���#q ��m�:��k��;����a� H����]�����K�w)�K�]��o��~����O- �6���F��/�_=}�������dt⥏�ۂ ���������Y ���ަq;�9����bsh6כ���C��M���CL|[x��ߐ����P�gR�JW�	 ��8���9��G7^�M�3� ��\�a��"�KtVc:2Y��B����<��w��sS�6i�)���؃��������6�ߘ��v<S����EK!�<}��E' ~IQ׳����iM{��^K���ǠHm�h�'����C"�`.� ��[�o�ny�e<�$`�{�KkbaP��*�+�U4�q��<E?k���:�8�a��"����?[ht��U6��4�=���^�[\�qZ��3�:�ל̔/�?�1u�б0g8�:s�'Wh3:@��-�7�No�<^���̙{{7��u'��������S�q�f[rq0n�!��u��k4�H��}�I��{�Fڐb�K�W���6���yiC�0�-��Z�A���ΆPM��ƣ�#���v�Om�-]?��>�c���7�rV������ͦ	p�G�|�:y�Ǧ/�6s�56eku���
�W&oMZ��Z��ͭ}�ל�zܖ5*?����pj.�F���䈙��e������m�fQ�Hd��2� ��X�"u���Z�ҥ���?1���
L�=�y��q,����a�C�l"k�3��"��na<�����T���}l0�X����� 1ym~`�}m����BiI9m��ī_w(a�%�~��!:�O�Bs�l`20�sp����V�ʺss ��|���2$h~��'q,�^N��	߀�2SFC��)�t��7���N�zx��T��l|kxɄsp�6A��V�֌hB/.Z����db��ޟၷˆ�g,�D�fo�w��2#�`�j�/�{�*�3�?�Ywhl)	t��h�XO/%�Wĺ�!$�X?���E��B�aE[v
�q�m�qt���a��.Ҫ+w��]�b��$>n�%lr��rs1��2)`���|}��"6��Ҭ4�]���L��&7v�a�������3� 
A:���^�{^^����ҽ|�(��V�Ƿ�|D��ʰ�LA>3�m��"�}�,�K�1זɧN�V�t��|G���?:���守��s�����b�7�^i�������L��l�,ӂ{n�",�]�ł��ē�᭠W60��Μ^V���Zv̦�ü U0&�7`$�m�g�ڭL�_h�6�g��D~���Q��� ;[�F	�k�p��Uܞl�L��+�*b<�f�	��l����hL��O���Xa0&t�n����ܢ�p�D#�ý�"����m�Nn΢	hٓP�.V��W{jR��ܬ _�te7o�4T��� �Z�	
��!����]�I��-x*C�ʐ�2$��7ƌQ$�B�1���k�pL"��SK�K=��z����T�Q]`�Y���k��E���2`p�������]*���Z����';��j�q���τ'�%]]��_�g�)�II��(�	;,���c��&���(�R����[�ܸ;�S��+��sK�}z�k"�h1Q�A���8d�&[=�3ǝ��3�<'����VѤ�\��x�5W�V]���X%���|��f��27�,�E�X�����I�*��DS�+G�ӛ�c���F����������ܺ5������-�|���
�'+	��,�:�PuC(֋4�;S%!�F�ؒ�%ڛ���J�ۃ���+f������<N��
�"v�O���F�����Ϡ *Kӳ�������H�,�A{���Œ�ӳ�<��y��	�^��k}A��z �q{�.,�������q�N/�m��K+�tw���ab?7���J7��x��Z�@��jtmm��{[�\��Y�OC�G�d]��WϞEU`XK��	��F����k�hT`�رU<$s��膸��æi��l��[�����,a�,~Qqc|)�-3�5<+�p9�(m�U���DT�ƻ����7=�U�_���=��k���ZlgJĺD�G8�d��ȅ�8�������:����/0-g���rꪱ��)6f�j����U���A�԰y��͠S{whZ?�B_F/
B���+?�q���E�j"�)�\6]@Gsb���Gv�m�DI�c�� ް����
sƼ]�?'�(�h.YJ�®;�#"�������f5����L��b\c�d���cI�3~i� �TU/_��e�~���y7n]!>uԼLw&<�d�wZ����@�My����Pj��i����I��x=�й�~���;�t�1s���x�Yɘ�#�K�o���|�~�{[���|Lt��Z)jXǷL���I�;�Н���fd���{Q��jυ�_�5-��J��\5�4��S9��,*�<?,˪������]g}F���~D�DU-d!�-�>ҼE���K��zn��~ �5\5�#�/����y5�}	�1����Ѷ���(Л y�jPeТ"�7�Uq��t�}}�-�P7��P�r�`��J?F�JK�בJ���e����o������Wy��*� i�ۄ�`e��X9�8VY��"��䟛[G���W_��W��m�bZu����ci���]�kw&�o��«B�>���[��Tt{�yW���Y
�U3h�5Rku�^o�'���Z[���!�cƎ�fаG�ێ���O����X9գv��T��I�勦oЦ�f��bh�yE�;��/�SmT�ҩ\��~����ˊ?��� }k�F��d�^����,]^�g�w�Q�������I��m��ؠ^]��7��TuZ1��{9�/:T�S�.* 0�澯�;�.)j���l/�	Z�Qs)������p"��Y��Kx�� {З'3�xk�Gz�?��~�~a
�ڢ�2�H6.�,N�AQ��ϣː���gw���*M�����8ʤ�NE�貶$VL��h�
lW�+ŵ�Q�6��mv��C��%�oD�>���.�
3�l��h-&3q�I�a�8%�����l���~�a 9�6��pk�H�#���XXw��a*�9�1'�f��������dQ*0�"Ctơ&d�3�oẂn��"���+����K�w�-���Ϩw�zu��)?����D��+�s�P�$h�[�yy����A�6�La���=V��$:�b��Å|��^%q�S�&�4'SEŻ��g(�{�Ԃ�L��)��ߎ�j��H����X_7^S����� �<���@2'�j�� _�Q.‥'|kn^���5�!���{`��������p_{���F~�uGT��)�oQ�-&,��>�z�F���Ue	�A��x��G_��I3������8����]��[�남�я�L�x�i��3�'=嫝�\j���"�:���"󭠦r���ph��jQ�d�����!񒞨�x�o!hhA��_�A�-�:t��{c6�5u!�hb]�HO֪������7)�#���1�D�\	?�<�XQ=�1׌��E�!%��3H\�v������.�Ꟈ��xbZ$<�ޓ�pj[rp�1('��7�����E-5(��"N���-�����J\m`G�m�6%�k��BL^,����,B6
'`�e21��;"c�i���6��L��$OgxS42:��ͼ��f���S�t	<C�-3?E�Q%aAj �i5���U�K<N�K*��:h���dc_T�[��r5 <L[�p��|�������'�g>�Y��>�X���J)�i�x#�0�X����
��f�Z�g���|7�9z�vI�����O���M����C@�A��5F�cJu�9�C�_ iz5�@�=�V�f� � �q�]��8;�xN�1WAjmW{xY'�p�9���ܫ��?vs��"����.�P�ę��"��9ZK��*\�MW+8��p���E��#D���0���*1As4����M{�����V���S�s�N%;U�V�����*�\����X�Ӧ�y��hv����/*z�'��֤-��j:m[\��
FR�g�	��p<��}U��?�{J�H��'ׂ5M2\�u���;�b$��%B�L�(H؛�.
h�M�_bD�V��^�8O�lL�~������8����懇��yP��9����-��)�8���H���9(��w�c!p�_�Vڭ���|�\|�X�y�<&�����{vT}֡Q��a��_lH�c��!���W�X�,*����?2l�Y��[��֯ni�:t�ː���/�#���8$:���Ct��.��3WĚ��^�0��\�>�'���l�l���*�[2~q�I�O֡pnl"�������ް�x�Tab~���
��J��땣k��D�_��6���t`���}�\/qX"A��5�T��NT:\���q����(x0%-�#�s�l�t����W�_c�6���rj�ڡ΢�$\ħ�]�	E!IZf��:a
Γ�O9CX�u������-�`ɎS&>�[=�����(Gg����ⷅ�K��9�Eߕ�n'�pHN|�"s��F�kB�1XF.�`H�`�;&�ӹ(�5v�C�����9&&�͐:{Z�H&D��fz	��hn:`��.܁5:���UVĻ�  1�O��������᥹y�,��X^݋�~��C�w�� z�<���y;l�5��]K[�"	X3x�l
͕��X�,bH���h�U77V9 ��=&or���,!���$}��(��Ƿ���S�D�������=��f^"���}>�)����ncl��b�t	�|�*������|u�O��D�/�Oӱ��Ty�&��GJ�Lz��p����D�8���+ǣ�ֆc� y�����x����ɪ�MR��[@��C'�ƣ��r�0޻ف��c�Æ�ֽ58{�fk\o6�o�Iڤ-Z�Wīyv�߯�����h�d)�����w^m!�K������[���G���n�K��e��ǣb>"�%0���ې��}�S+��X�Z�3>�t��d1���:�p�hGl��];��I��J���'0l���^n�$������'�w���;������@��/�T�FR����ޏU�)�k2P�!�k�]��	�Av��gߝx0(�t�*�}��5�af�s�!��uC�ŷ��/4��Ο
��^��*H$k\�{���������l� ���c14���vvЩ 8��vHNU}��x��?�C�?���aeUKU0-1��ê���\}���(/(B\�3���S�͹��:�~;>��$
� �teբ^���$�f8�����M-N��@����Ӏ7�YH�Zqh���p30�Nk�䗀a�65 �Ų���AK��;%� 5G�R�+�����+��'K������`�q@|�6�;#r=n�fI�DZ�:t�\�n�r�6%�:G��h���ɄQ�r�CW�H�0���#$��|`�����2����CՔЕ���i���>��PtO\!��C
���8%���x6�/��AG*��x�ym�u.E9�:��zpGE|�b�:����1��+�rX�8�iJ��|�2}νd0l�@�[aI4f�zfo���`ks�}�"*��j����4	�0N*}��T�HOSFy�g�{����?�8n�F����\�I��H���+���4ʳ�]�Dؙ��"�ܕ������Y��-{P#Իu�6&��8c�q�-�m}�x���EJ� ����G�RUa�\���696���)���v��D�������_x��q۔x-S,���҉������I���7��U�!��ы��Qp���g����2��%���>�:�uu�����
U���������	����_izg��_
�!�k@��֟�6|�5,B�>�1+&p��h툯6�����%\�u{̓��W��I�ݎ)���[����y(2��'����Xh�����ky��΀~>�u���`����y�x'���ȞZ��^���Ɛc(� -��9���m�5��������;�˦��_GWd��h�D�OL/^���`��bmZf*�%�ѼJ{�]�R6�o�8�V�А���C��竏Ź)"�h�,6G$�w~q�v4�	࿳>H��4YJ��Q���)�V�A��^��-}WN��8�ݚﲃ���dPlh�9���Z}3�/�.�u��G,$��L�Y�I�ι�J>D��e�%ME(����eHZ9{�NDJ�����ӹ�>�O��DJ��OLM:a�e}C�2��$k� }���$WO$����ã5��Oʻ>r��e������ϙ�sAN0ˤ��bg��@�1ӵ���piQ��ư�Ɔ��m +�=����K�L0�6ά�G�MvP�hE,�,�;ҿ0.�XQ��N�NM~!VpT*~��U�Qo����v�>s����!O�$g���U�i��k���;:v� SAS�q.�Gl����]6�oo��zvT�R��G#i�<�nn	,I	Lso�T��賙���^'��D��(��W/��T���d~WrM��g����* Y"��>=�
/��Q٭;cbc�Z� YѺ_�"�%���o�~/��:6@k�H��~96���x�;^�؅�	�8��r9��U���⽑���y��-��"�uЖ����=#��aM��<>��I{[�V��Wn���T�7��(��>c��zx����ω��F�Rh��#�Vޖ_O6��#�@����[s��xx�w�)�<ɗM��W@9�J�u9#M�ؘ�`���jw֣ܣ�c���2P`Gk�nP)���S���g��l)�=�v�ˬ�5�m�0�t���Zw�ε,c�:�SB�Y�7���eʀ�V�'��ߜ�t+�L/N�(�av������kۖGH3G�W��|[r�Ҹo���ֽph����,N�2�E��:U����z=p���|A�;w��s˵��XuS�M ����q��O����2e�O�s���ǹ�f�6O�P�L��BPU�~�S��r�Cb� ��|L��R$�H�I���\��v�q���?�)bm�Dg%��΀)�/jqP�JX-0��� 6}����/Ueb�A�!1�갨�b���uJz��I��-fr��"��b���y�w�I��7�,���U��+}�4��4?X
��5۫��˫Ȯ��r�{���V������y�Q��y����r�i�i�lȚ���w��5�I�(.�\e�H8jsQ��_p0����V,�M��^�u=V�0��+R�y�5��E�C����m�鱜��Â�'jA�5K���QOo�[/�ck�R*�
�!�����V���#���4\��_6W{�+B�~K���
aU�<)	�Xd���oL�1.��ض�6�v"���Пo�����@/�����fx�A��Ux�g�R���d����(�1{$Q��x���b��3<�i?��y�s�4Y�}N�.�C�Dmu�����_P"un�D4o�ʫ����g&J�q�6��{A����No�7H=C76����)����ο#��g̞�-���HV�����	���ʹ�5��|	��0kb{���iٌg�q.S��c��;����o�n{�=�y�h��I;�)Uh��z�F���7�u2�oh��D	(~��L��a�"kL���o�\�WI�K�ꁁ���8k�vO|�4�q���ZE�D$o0��7�i�mi97`A"8�B�����͹H΋C.���L���� �5��^��x.�f)�[5!k������^�T����1��s�.����<�z�WK[ى(�UB)���:v���5p��{����.z�p��C��/�x͍������&<
4�Af]F�a�?
���a���M� b/��'#>�z��}2!�BɞU����}'�zf79�p�k�����"p�@fq����	��ß�U�z<�zL���\m:"�J�Ux�#o�{^�b X��ʵe^���͆P�ŧ�|����k��W8�1Њ�S`����J�s�Os{������$�����G�!0ޔ2��]!"g�Z�b��{������uk��ln�(��$+��C��6��ɿ�CNg��lUgi�;59>G�8�&�}ZJ�5�q|��$��䶦�я��E�?�ӵ(��?�e�.eM@m�;ߢ��[�o߳���q p�3���E����M���� �-O�K�����^x��������>ܬ�pI\�J��AR���l�����I��4{;n0;���ʾ˦ɞ�O�)F����ή��?����n�^��i��΁�#W�"&'-�I��gO�o5Z����9%�t�Zk��#���y�G@l�[(�>�WI[�s��7�˽L��ȕ��rPKO�`q}J~h��V����D?���]��^CXl�|g�9���7�]e����K���MYA��������^�����t�J<����b���o \Z�s���n�jw����=�'�um���/u���WtTA�%5�({�%���F4�.��r�0�il�W�Q��ДOŘQ	Y�ѕWZ�LBi?T���o���V8e�a�����N�M;ג���I���yyf�]U���Y��h�s�s��T��#���a~�Lқ��Bo%��&y�����QB�ݴ��k#���.#�)�ՆV�c�M,b�[�CV>>��d��&\�8��序ܸ(����:�
bO���L���3JB�(0��z���*�ӞD�C�CɜNK7��S`z�Ԋ1��m�<�(о5��6AQCA؊���w�#Z��͉���>TU��6m�dS�Ŋ6��u��K��6�Վ�^y�1}�4����ݦiW��P����?/J��k�ج�9��|5$q�"�@���N�8\���g{��Ȼ�( ��Hg��5!y7��h��|>支��~
��M �b�����T�(�4����w���4zC��|��tk?G�W����b��Ƹ��e����ad��75�p�+�u-&��{�Ը����q����af�e��E4�w��r5�P-�o���Z��X�@����2T%�3�Ne�a�-���\(ְ!K��e1j#Y!}��챇��5���'C�Kl��(9�#S��я��������?���_���o.�S���wwG)x���>���`��#��_��i�h���B������.���C��o�� �����c�V�oyqF�髽���/�؆���']�-h���o�^7<{�q_Xt��k�\1'2�5� 9�����g��)l��>N���p����-3���a4qHUq`��.�^�V�t��A�0~�rCL�MKsd�9�>�@��L�E�g�	��1�Mp�d�����jTy�)zJ���'�M�ՒqM}�ԁ`��Du.Y�hhx�R(45�z�?sr��;̉&��0r���T1�q
�����z��7����W�~"D����h�?�p�[�w��`�E^�J��B�Q)1�t��/XS6���nCj�	-X"�V��7߸a��J_��D&��4�����g̃N�A_�����s}�FI����Q��%�
��E���.x"��i^�t�q�$�`&��z�o�Kh��t��H�F^Y��Bz�����"������Æ�u'�r��*�z�Q���{�������ʿ�D@�;<���kP�h��Y.��G���LV��A��F�.	z:(�e~�CJ�����_Ε<9ǀ�����=[P	α	78}���</`\��;e>}{!tG�+�� �|���E�]}�؈f��1#���v�
��T�1y�@�����7?��{/)��й��d�
9t�|������}<[��w��4�D�����T����������ڗ�f��Z�Ҿ	:n����_}'���,�w��m�z�z����TQ��P{����7���j����@�*{�#*��'F���b9��4o���Y�[ny��7�$��Y-����6���U�;���/��r�5����N�<��C�T��(����Y�9�[M1 ���Ј(��٧�+��3��뢡ְp�G�}�<��y���s�r�2����s#k3-��Il%�(����q���>��I����}��� �d���~��8a�ppS�>,�U�R�|^��[���l����-!�YƳ�y��9k���z5�����x;���8&�����]����!���c\�O�5W�%^驵G�\���z�r�4�4��K�zVZwMD;���=�<돪u���[�^��@<J��;��M��~�{J��y�=��C����=����jtɜQ	��Ycm�`O&1W���L|v�8��Юm|��>Ϩ�I|�{���l�Tj���7�h %l���8��r�^��؉�y��\��|H.��7A_�_۳�3z�NT�j�nWmd����	�ߤ������e�Z9��"h�_W��->}'�>f1��%�����p�ܖ���~$ 7��G�����К������iҟ*�!���b�r�,�|	���������g_3�!� ��Yb�힨*"�ZLdۮ���{e�'��K�&��{��w��({>N������c�wMds�Vuu�n�-}S� {�]q�U��BրI
����+/ĕC���4w���=��6��R&�h�8���� �V�ŤW��W���*iiODs���ٲ~�R61;% %c�I��?���F�q~PZ�Hc��������[ڭ�=�W7��{�m杸��Ip�U�fl�ݫ�6FW�H9�����W�������ĳ���˒Si�CO0'EM�_Y�����]��)6���/�=P\�MA��,���Kd��D����F�QS��m����@�q�);c/����C��{�H��u�,�=�
��ĝ��5��N������fMw�O%_����3���yp�r,C���0��r(�.cB���{���=�y��ON!m����ܫI������GD�Է�=�b2�^׹�s��p�W��1��]9������w��]ؙ�/�������{ݔo<'�W`"J!�� !jd�-�Y�g��}����$�����&�
Z0�~�~w��-9�jJ��u���2w�}��9�Z��Ja+�U��Z��\��>�N�W�
#���b���;0M����P��?�;�_.��>� l��7��%.�6�x�iy
|�Ʃ�IhZ���4�V��S[RdĕI��o=lU��ԩ��s�ׯ�� ;���yz���w,�������v�1J�P1�;�g�s��Qb�������R݁Z�����Rv#��\l�Eg��[��DV�;�ے�g�X��9����h3~�G�0ME��9��>@68H��|m]�^�ICΊ�ꐣ�o�՝�m�R�Ԣ��0z���}A_z����*s.*P����#��k-;�i��z�[���.x�o������ ����	����#0[Ŷ��O5��"WE�T���-�3%����`���%h�\z�b��_7����qJ��	i ��Q�V +wȉ޳��A��|rmw�h���������"1��<�*�!��C�<�:JI�I\\�X��~<�&����ۻpN#������x�/�x��eG�hH�3	��?n���[�4�)������f�X*��"K�o���\����;�j~j�FE������{���C=�b�È����\g2�co��z?xdJ�G"E�(�J�����z
�5&�hS���_���`T����O�JHX�Q�o������܆�܁O�
�=9�x~ͤ��8'NK ~<��<,���Ԙk�����U��Ҳ[�\�ω7�V�q=U��)ސ� ����H��"��V��@y����_���w\�(T�ޯӚ��m�l$�>��i�V��� v'�����f�Ź�hSPjn��a^��䐝������G�
T�͓�K�G,��#~���y0���H�+�rm��$�!�-E>[�LO_��kr=����0q���q��D�)��hӼ�'_F���~���jo�y��VС��h<��Н�dr�S}�Q���=9^��Vy��r�8`�ϵ"���Me�g𤠂Fȕd��$)'9_ތ4�(o���4�`�����iVT���܄a����'�Nۣ��`C��wU���2���M%Yj�!��3\�����N�����x����w���Q�'�{nC����u^:�'
�Hj�R���}�Gts4�����݀���^�;I�4����Q�&6��G~r�����	KF��#�����^�K˙��5-��P���0-�7���Ϝ`�Vzyc`�}A9��!����/�:�D�s��jU[n �p�$Q@�jM.�GB�u
/G����"2#�,O��D��Tu��R}g���)b� 9�;NsϤ���U�s
s�%q��������7-_�[DeeO+O�����%nz�[��kK�!�kpS�fIQ���vSIk���Gv%#p�	M3��A���N��J+9��K��N˹��/y�Ǒ��go���]�Y�lD.�FNg��C l�(�Fv2[�J7[����;rR�4g	���؁�aO%dS+�*!��nj1�j�ڷ�7��e��y�7z�g=uۛ�@�Ԓ8neI�!=[�@����_�X:`}���|�����9o���q�<�H1r�&��;ԛ��8>3��̅&�s��l�5��� ��sU�#h��ck���ȯ���Xq��pֶG���O����W<(�0�nb��7к��#$����:ȼ]�Ȉ���e��*���z7�'�h8m\ؚ6����[eDa+�f���������<06�ǲL��NBU���4MG�"2YN#���G�Tx��߻D{�Tr��E�f(X+:�ܝ�1_�嘏��i3sL��$+�T�S/�2����z�DzCl�È_�R��;e�.���
,/$�h7���ŕ(=5�4i�g�j����2��?��v��]�i�wS��f������-a	�dur�hoAշl��us����=e4h�t8z �{�������0pį�
�zb*��a;�º�1c�\ͺx�>U��� �ed������I��=�#�rӆ�҃�ʎ�j�O�y����?k������������Y���[iONs`'�k~sA�9GB���s�N�F7��Q����AC :gv�@kΐ.����,2$F���D��i1��M� �j�I�		�mR�͡%��m�_j}���FB�M�Ȧ�D4�fd��2
Ϥ���@p`�l9��K��!W����M�xϤ�ʃ	ϻ7*.�]�'�Q�̗"_;�^G���SS��#�D�rn�|��d0O�jo�BsT�V�w�tCj��`�q����BZw(t/ ���j	ƃ���4W%Ne�4?���}7��Q3�N)�=>uٻ��2H7�^��=;�o���u.��83�f��wZr}H*,,�2��,��zJ�����|Ga{��z��
?��!)M�:3.x���4:��V/�tz<_	��ёW��/��UJޮ���� Y��f�H_�H�.&6�Qc��_�9s�l
�\ �~��B�<��dؕ�H8�e���9F�s�n���3}p�X�M\���:�	HN~Iy��<�����Z���f|)�5/�T���>F�?��UO���������N�KP�UIC�򋖦S��ե����1߷�g����$C�B��u�uYp�d�d��c��44^X�l�l��r���"��B(�Gy̙����p �����K�2YЮ	�e�L�D�6�3�&��@j֬�4��`g̙ˢ��@�LY	g���Se~�E! we��Y���4G��ӧY�2�;ue�Eb��2d2��@����h��$w�!6� )^.z���gjN�>Wk��DcTYr��G*�*t�siii�M��\X:�� B���'x��A�Cd�e�Ȯ"q�
����ԝ{�ߞ�V-�K�?�� w�.�}�Ů�h*ؒ�[�g�S0W�wy'���N��Tܚ��ѽW�����A�;�us�kL:U��	K�%���x�Fk'�$'ة{�!(�'/��ln.�e������g@��[�N(��œNpU�E�/D�^x��,�+�t�nZ>������w�n�l��7 �����o�oM�tغ� '��a9� �~-�N�����Ax-�vj�@�ug������ۣ��aS*@xO�n׽y�0�N�)ú���p�I90m��8.���Ԭ�J�������c*K�k��j��5��DZ*벾~%�sf�M�4�p�.���5�Vތ�Wv5��DpEه���(4���Ҡ��ieeGM�OS����KGO��a�Hz�L?t���<tv��Q�� \�>X7j���-�d�R��fQ��_���%>l?nj�|���U���S��ľ�y��z]MC`���T4%6X�������t�������o� ��I������F�����8�Í0d�����L�&Οy�}hop��F#(2g�Yq��ʦ����;��Gmi�����me�5K��2�JT�����bC�܄���>�	���@� �&�Gʜ���%�"#��!�z}�\����C�Hpş���� ��:���J��JS��x�i�L��<rǍ�/�-�˵���_�I�]Ey��&�i坡���A1�"Sn�V�t��׺����60�S�,B۵��4lV��m�bCdY�hN�,k�O�Xڧ/<��۳����¬"?�1!F_��!����(?�:ރ�v)Z��P���II�A��12~�B����o�Į������%pJ��xe���5�l��4�7ͫro�0i�@ ��֙r|���k��6%��Ԓ>e_߀�A�r�o�o�UV���7���ij�:15M���ML`nX��C�T�����[����g�0@&j�*$�����!�������� |��􀉧cz%����a��Mb�O Ԋ@$W�[���j7𩞎�P��&��-��q��+�����8Q:�"��TƸwk-�$t&-ծ`s����U���\z�+�Q $��C0HuЋ��X��lL��$]�V�4��.�M�Ċ+xg��0-���F�!�P���R�9�Ɠ��.�+2�GUǭZ�>`E�@9�����w]=挭��6�X#��!�^�o�Pˁy��*,8��,��H����,�,z�OUsD�VD���]������K���HpF�&)Qk�<!���H�a��v��VY�|���lG��n-��ok��@V��Nu_����G`l��
b'� �n��0�`�M�$_,��N�= �L;�J�
�,���#�d�L!\�\е�J��������3j5]_)g���d��dMi��B����"��ABxd�n�eI��f��؁%2�܈S ��C`j�կK�k�K-��j���+
3��|��u�%���}���u�2P�h��h����;�p���E���vaV =6Nh �'pb	\�~\��)����	 )�I4��|�*d���ZB�X6�Ȓ��� ؾ�T�wbsX"̔b(�	LL-�jT�Yu��E�x⺖�Zv�pwhw�Q�D��6ڥ{�^BlX�F`K��b7�Y���}Ϸ/j�!\��L�|�*�I�M#�R�\��i�{.4��UnY4�5M0mQ%�%`� ��{b�1�_/-oK`���"ӥ�mq�����OZ�~%�*�L�ڃ�G�%�����H�;�˝[9������a ��H�<�y��Pm �D��ދg�{��[�W��߼���s�QRgoF�S���%����s��	ke�����s����&aZ2�
lF��U	AeW+�j1�kc�;��9t?�4 �~p�a�d���	'��WՃ�#�����ʒ��Y8N���~8_�Y���X��r`�!�x�tKG�3�P�`*@ ��d_0��b�w��݌);oTtP�Z6IK�O�x� /��Mn�x��ǉ]R���d�5c�Nz�O__3���(��U���g7̘�0�-ˠɾ���}�{�d�R�}c-)*m�$$���-F�%a�J���f���<�s���}��<�9����D�4��8w�o3��<�ߢ\Y��Wa1^��R��h��W���>��������,��J�0N�">�%���H�+�@n�
U������:x�p�
y��p�p ؽMk,V'�Fڂ�2�m��;������ܦXƳ���w���_p2���Q�F�t���?&�M)5�:�� �C}�,�:��r<�3�;$Ln�@%�S��1c`�*:ϣ�����@�W�B.� d��=�[c����h��}��X�<^!3*!���0H�eH�Qw&xП��� 84㔾�tV��V&�J\���i�!�Y�@h��5J�ܺ�ft��tt~���pV�n��3��t>�bt��h��{�*Y�jn��^�3Uѽ�u��s��ҷ����)������z��YY�&�CJ9Tge�)����w������6.�|3���}�*�-k-�嚂��N��<\��ϿVt[�E<+���*[ax�p�B��{���7�Ș��s������$~�J�T�;�����*�4���\��R�KyL�e��ZWU6ռ�k�t<b�F'Y�y�QPT#�\	�gI؁J0NkN�8�.���̗�Ż<
��r%P�Չ�y�t7�K�S	ٶ �\��Z�6<V����&��qlA� ƍ�_�����eB*��-��Vd#Z����VZh�s����D�Q�����kFl3jZ+K��i�l�m���@�(�S��bͅ�ဗ..ܓE�5����"1n�{ZZA
(^��#8>"�c��d,��U�n�:����u�����7�z'�|?���ޢ��z�����z������z�2(�Z��o�^����hb��k�9p�'p#��m�W�iڋ�����;Kb3� �毹9BFل5����$���n��:MNV�'��0�4f�XR�����u��� Z�fp���n!B@����J���yG�`�,�E��<({e�RHbA�T%��g'x��ú(Y�A�6����9-1��zF�W.{�j��U�_&\�4�z-).���D`��y�m��K@v�v���"������7�I�9�[s�I�������B�3
� pQ�X�4�=^(G����^[�k'^���d�Q�VF�%�e��H��-��ʘY�F�������d�/�՟�THS7%ȯv}ijИ��+*��?Q�j�� ����ĳ�G) `��o�xA_Y�Ix,s��T�: 1T(��!-_v���?�TU���{z��W�ǁ�B,���i<
�����f�-�	%�W�K��
O�Kz*|.��W{�PX%5�g�A�|�t̼\D�Ԯ�9U䁿���(ڠ�n���JE�-(n�`	�"�C��4g�Z�X����+�d�G
�P%n���-������dm����/r��u��"�t�Ŀȵ���q�����Pf�;�p���[T�^A!���M��B���PU�]i���]\�I�Ձ��0a��Z�ֱ]�t������6�[`˃G�%�j���]���e����=9h��_KP�!}ee%��q��p���;s����*ƾ؟w�j	!�L\���f�|mD��M�}=�A��?Wt���ƂF9�Q��E����=�V���q��<��s�c?q|���=Z�J���8�����P=��WV����r��q��+��q�`����@L͂_���U��c-<(�bp��0j+B��u�z:~�ղ�W���_���4�)*�
��������waf�nm�mCi5a��Q����VQ�����Q�� K��Wt�U,%J�3��]+c���A&( � ��+ZcyOں ��y�P�_���ʙ��M���i=�x5#:fC!M��~�
�fD�I���Ƒ2~Y�l_��g�xv+Y�f��+-$�:��L��ֿ��Y~~ ��M�� &�e����������\G8�𿅒C H@Я ���5��z{���t�HXgX���ض�?�y�x�:pWqdO��<ުl�X �d�lS�F���m��L�5,�5b�Qq_�7~�d[���7e��@��̵�Н��������B.A���� j#�Jm�g�M�����8���a|��*P�����6�Q��r�����4h2�D�;�u0�
��<\��v/G�#|,�X)�����u�8N<b��h�^7�F�)]��w�r�1��w�U��5s��_j�}�>Y�j�����ҧ��g�O%'/�	lT�n�������[�d�����ވ���C�;���|���D�G_�eJ\d��w�IE\L��F
w�(2��c��~�|F�n��'s�4�-���̓Z������n����4�i�χ��Rb#�b�i6g�J�������Ӕ���2s��r�� (�J��fT�W�Sz�}W]�/8�T���*i��޹��?���,��`���9J$v-Őmقd�	I��jF.�� ����T̎ ��X~xN����֖]�"����-��c�N����`���f�FpA�X���V�*�tׁ���(��u8E��������f��#�ǟ������<˫�T��	X�4��Ř�����P�G�����1u �G�gNIT�0g��+&n�.�Mn�F�(�G}�Ŗ�3N.DI��"�y�����s���*�ok�A��7�%�j��L�yұ)���[�����-�+R�J�|�S$?����-���ϴ���wuT�S�h���o�`�2��%�K�B~/��0�1���ի	�c 7^4lj\ �'IL2�>~���+O&·vpK"s�N�Jk7����(K�ҫ��N��
��U>�h�>;T��&�E�+���*r�N�Q�V���� 2�)�D���z���W�J��~q̩꫇�q��T<��B�����I�U�N��1ja�*��U%[[��,B>�/2-�p#8����l��bK��*���f~G�7��
?�`�Z����w��-����E���A�ٖ�.��6f��S� �����jè�kv�'�BO��]�>��{{A0p���rԲ�R|�fVj筻7���43��⛱�h�[d�T���M�O>^�})�Al��$��~ ��%�ԅ�AYy7nJK]����� *u���Ε�)�h��*tc]`�+	P7WNx���3�G�\D�kW3��H7tQ6%�}ٹ覅�'��a�?7�I��M3�Q�4�V�*��j �x�.X��L~��E|����-�҆F��K��u�*H�_%e\B8HZnYm��Q\�[�[�H1���^i�"�(�" ��|7x`�X�� ����y��!PsŃ�_zɅ������8]~�?1���+����EP��Kɰw~ ��s�x/���0=���X�Jh�Kf��W������W�L�F'�kf��2��U�G�ԭ���� CXPH�(���)O\�!~�8{^wW>_���+��]�`�Bp%�۾3�s��u���5/D�J��/��<\/�s g�Z�9*�!.��k+���O�bY]Em�[�Ug�c���%��=ZU�Q��i���ȡ��S?g
���
�*���y5�^��5���ܜJZ²wP\���9�@���*o�H�������X\�G��/�� � �R��v0�C�u�-�!P�� ǃ���T���(.
%㞿�r㡜���jX�G�h����x��ߟH������/Q��e��6�R;]�*`VD�aH_�q:	H{�3e�O%��3��9�}jہz7A�d�4���e)f&%��7�/`��^o ,����� 9��Ѐ�7���mu}�ˑ����e��w�B�*��� �63G�޼������.8c���3�tV��%�d���!-��L?��3�	�I47��Z%��jn�?X��a*OM8�w����A(��l�qh�{NMA�m?�����m�I:������żP�n 	�[tA��c.�|�w�w�psd�� �A<����&ª����6�4+�{�V�M��&� ����G|�tk���f!�6o�W�L�	�Yv�`rkz��f8N'�
��\�/��`�Ƀίy�O_ۑ`����6w�IS�^��~ߑ�)]��j7%��}�CQ�
B�(?�zx��ߓ��ݘL�	�֤�P�Ϡ��Ȑ���xaս �rf�'io�<�i����}���g��fпb�U��;#���@��q��1��ʣ@���'��qr)Ѯɉ�����׊�!4�o�e!�"7F����+��]4�N�"�#c>Y,_{Sdټ�ۻ�II�D��ط��?ީ��tDl��ȳ�3�f� K3n5k/����3C=<�J�1UBmf�x�o}k�BR��}0�+N)�/��x��D�*�L�U�pN2�bpc�E.����V��|�ȃ<��R���$F�U��1gq�N���xA�[�X�><���}�S� ��c�PJi�5'͟i�>�ϙZp����;�31�F�N)�1*y���P�^c�Bg;�q�l�?�v��=�B� ��*}zm����u�;�rF�?Oq���N�:i���N�����Q�K*e�o�#��!�gZ*�0�a��|���+e5�:O#b���ʛ�8_f��4磀�T�Xk�R[ڒ���7�����@`ر���h�	\�n�s��z��v~���q 8�t�+
�M~�+�P\Ft�u�����Bl4�= �?�3ZSN�k���|�|I�j����'��o��俑�Ug��&6Q�ME�4a�F�E=��J��Ů�vp�nff�{���uI[JX�G,x�w�9�����#zAy�i�
K���z��͉h���\�t �59y��X.*��v҇�a�x����<�����9<y:�=Z�A�'������3�c�������r�q?��J�`:��ժE�/1+�܌����d���(�?4S� ��YV���*StƗF1o�v"I���C.}d7=C_�]K3�J�FQji�޹}�y���>�G��F�G��������e|���Z�����@	w�b��Rs���\u�6�w`J;!JHN���汖q�Ȍ��T�&�q\�A���`���I}R$>����W��:r}�X5ʡ���Z�$���S�" 9�紗ܲ`��(��������� �����9h8"��$�/A��J�I�����	E�'��';}����ʟ���al��d紇���j��N�)���	7����kh��2���rmrI8��D�U�`������Oh2e��;mЄȄ��"����6%�vj��8�e]Lb>Dm�����H��Ec��m�}H��%�@�kq�#ۧχ��&M�GB�)󠠣�����S�`�<�^ 1�=�ۮٔ}I]�Ǟ驇|���g�8���$-����r"}���Q�ʇTF�}�9 q��WA�`�3���1L���=���Ύ͍���L�]�S����s_��ȞOw�dٜ��`�P2��Xx����C66u�i(�3��P���ſ�m�H�j�ySw�rލ����G(�8�@O���(�I�J���!Ԏ&E&��&)1�D59�=Gv>�-đv��������p���9��6'�"h�GH�궙�z��ӓ����K�������Y_��N����0��y��g�(��giȒ���O)Y��%3N�)'A:'��G�?�z6i�51�0�u#�}.�Y�g�(�d#����
B*,e#��Iz�NA6R��?..m�2���X�SB��q���۷�����*q��4ćLG���ߠ�F�O���=ع�����ӭ�2�3�*��N�f��� �:�{��=ȸ�&��E��ռl��DDP�\2�������>�6qW(�+�)gJ�TS�:����1����e�`߹u��F6ս
㺠�<l�>�0���e�"��[�< M�Q� �**����u��{l��{M����5�gl��Xᰠ~n��Ҥ{SX�w�Ĭ��@�l���!o���e��o��~Ӳ~�'��jY{:���1 ��p𬥌{�m���,_�r�>��˵X����)ug���z%l���OPO��M���H/������)2{�)Tr?�u���>5欹3�s�S�h�������1=�L�>#���|��9�3�ǿi��u�/��$>��U��[Vl��-�'�栃|p r��GDĽh�o���|r��tu�x�5�~���i04�s�`�b��fZg_2�s���ׅ�Z��?	j����쉦�)*[۴����06��f�Ùu�ɽ�^  ����+�c�j����>=��Z>�4���*�e&����8��ɎJ�<~�<rߝ_��g���E#W��D��!ge��?N�<��Sd�̎CA3�Ѯ�*}-<�a�����UT�/͙`�ύ�]���T��qY�3N���%�����oj�F��^O>�|���th��/� n�E~���%�ir�IS�@է{�`b*{od��q9ǷӠ]��d�g3�_�K���������zzr;E@���Α?��`�W�����ӋB�o�k<����d9G��yp���m�c7,o�|�Y�߿}�7�@�Ȉ��u��5;<��.����ܟ�s;�}7.�,�-��)���b���S��E}�������W��/�����/���G���06�V�X\|)�߽x}5�yp���z0�����;n�-��]�����k=e��!ϲ��1\K&�>?�h��-zlL�S�<�/[�OF�TZ�L��C	���#k�g	;�>N��HA���x���To}�8�#�z�Pf��{�Oz�צ��	0���rLK�j��j�l�����a�Ȩ�ĵ���_wD*N=z���#}0E������@ug3"������έ��bx�|����8����slBf�^�����*�i����7�������(5{X�W4yb�E�r�7����HM�o->�v���|f/`|�������o�� ���]�����v~m�K�2	�{l*�K����n"e
�g�&�0�m�g�l���I���i����څr��Lwc���Ǌ&�4�Od�ʚ��8kPm �y���p#T�t-��Af�0�=ֱ�[5�H	T��Q�7U���p���L��0O�2��9�x���N]��-�k*�Gw�ȶc�~�~�h&��WCIt�_|w���j(�<��:��Txƛ���}әHl9w R�Q�|�9��Lx���&+��5��������}��
���$��?����(.����d���OU�:�W����.�QV�,�8C��V�R�)�+�y �H�ʣ-��pߘ����A�a��b;��'�8�ʌv~NP
���h�T�.�G�+JT��ߝ#�en��$N۴؃��e,-.i�(S)-�.S�?�|�Ț,/��x~�ϔ�m<u��7H�ڶz��A�ڛ��2�Mhb=�[X�l�1���H.<�5q�rz�s����2բ����T�V�u� �5�/L���w_�Jb=��q��G��  Ky'
�[����#�щ��]뷏�6|���kL���j�!��c�`l���ю���h��G�*7�&�z��_M-ߘK}�y!Ь8���76d��,����2c�u��JQk1��O��s�7D�e���<���Z��"�n����w�Yj�:=	)�f| �Hr�?�3!g��3����	Ǯ����S��SXy@}���W�\�Rf�H9.u�+1�B%�w��|�9��b,5����$��}!x�g8���s!�C��4��9Nd���|��i�n�zvN�	.k��{�/���wrkO���H�42��~(�8��j	�OI��y)�}�����z��|����?����{-�cmM�*�����7��^L<Z@M�c��;�8�5�["��ӭ ��@Ķ��N�}�Fr��=L� W���"s���j�0;�Q��=��b���;���ˋSzR/ �����s�����E����J�W˫n�>{7�`�	�F<���s��~@�c��[�4;gg5]����j	b�#�͕G#5�����N��L����x���э����tt��n�h!�8A���)11B�8�[��݌yߧW����u�Bq�o��쑕�>�Ľ�̕063�g���9��"��թӘKS����[�G7
�w<��;�������Ņ���߃
I#i�5+�9U1� RCb�O�8y�����w���_�s/�����WPX}6"=����t�E��UV��ڑ1*..��=0#�����Q����+ۓ fO����g%7z�Z"юW/B�)~:TN:V��Ǿ2-$;_����͜�\�@t�� ���E�����%DϺr�?�G	Ǣ��sH��>�*��d�ʑ�_0ql�O4w�F͑�BFg�I
��C>W�㙙�nѢ�.*b�^�D�
n?nUQ	�7�
�x�d��d�����*nG��o�ƾ�nW�?0S鲛1�<o����o!��[j���kc�+�N���]y��V����m�/5V�7��sj2b��T�Mei��S�o��եt��V�Q�X�@����KB"s�{�g�p{ |n>3e�u����D~��[O�F�S�Κν�����E��3���9�N�␙�غ��U���&u���/ʂF�x}�P�`!1s?��݇ƪ6tn��$%JP�Q�Y�(
��t�;&������k�l-�����V��h]���آ߉"��#X�쉬������Tp	k&�¦�5	��D{�<)5�͛d���KY��Qt�vr����L�y��gd�5hՋ�BI�X�F��c�'��������zz2ҝ���S-�a���-����`M��a������Q ���\��c�\���x��yt�[P���W��i��5�+��
{�4��>��/�0Z�bN���S�U�H��ϰ�&�����[h��Q�S�q�ޘ��eH�kF��i���O�F��萑y?p�w,9ݦ�O��-�Wy�//���E�k�m��y���m:��'���<�Pڟ�H��]��q�Ÿl{GA{-�ô�SY�~z�n-�d#	���z|w���f�j�}~�#��?�/Y,�Pb��/%u9j��aM�ȭ9��=��Z�ҙ�Z��D��H?F������v��/��V�ʣH��<]p������Ĥ��Fꘕ��n�֞=o���E��I~�����`��q�O�Ҕ\.u}����<�񃙵��&�1^�o�)�RbX�㹁&`Y��i�ɿ���'Mk#
0��ؑ·h���}�خ����ﲞK����Ԯ�������hq���K�R٣���㝡u��nK}k�{�T�d:v4y�jZj���D��oz�=)���<-X=�mã���,���]��^#D�22^�?k͞�Q����q�����_F�\C��T��:9����b�iĔ5G�w�C"�e2��� ׭c&6)�ɴ��	I�̲N���߱� �
�O���q���UOa�P٪����p�X��q^��(�ߌ呬jQ䧜�XXG*N����@��(������6 <�4,GƸ��G�\��j��T�����yq�'��<��1H+�k��W ����s~ q�
w�\
�B�^\��y�z}�'}X�441���a{��iuQO�}w�޺H�Z���*�g\����`$�\>A�<뜻t�P�<a�<�i���F�K���pj�&_��̌㌎V5�/����c5v�o.z0�_��MM��%����m�պe��L�g},�/�������0|�#{l�d�!ѰB֌M;.!gZ��O���9��>ֵ�����0B�}.z�4��-_��0��;Y*,c�c"�`0��!m��6��UoE�w��_b���^����4��/;ʥt�pY�n��5^�z�5����Ӹ�A��#�a�e)G�k�%�2��k���̠��J�b�]�|U=�@�+I��{D�Ò�/��K��1B���`�S��W9s�S;�u:x���(��˃��e/t�^$j�B/��OT'	����*~^Ps��#�@�a&S�rF�].^��+���#�NZ�2X��D6��sYq��ZZ���	�f;���>�4W�K�<x��N���B�������fN��'"�KQ��;���)4Dy������~�aSF�������G����Z<'"6�;��}~l�"�p��;��SEd�z��k�p��j��Fj���U����+�-ՑV����h��wѻ��)���_����6mwg����F��2u1:�����I���S4�K�}Q�w1�_���Y�
��cm�{+�79�a�h܆��QJӥ�R]�H�_����+�T���{���09�}u_7�\h�� ����Ys1���fSK9�����U]2=��9�?�~v���{�l��YC M�O�Ġ�7�ݬ��L�z̷�����z�v	*�=#�}��
�C��1~/�7�ݑ�6*�M�U��P[{��Є/�/�T߻�[baR�lr�4�Hw�-ę�B�l���0q��d(  �V�i����V;j���xǑz_#���rs���EJ�+WUVVE1�˥��˗˹�z,���Ih��kI,�����9��;����=������@׸!,wIߥ�o>�i�.�+�Ю�t$�&�I`J��q�4ZyNR2��J���6�V\B�!a� �۔����j,�41A��B��x������h:�Z��q����#.��}�|��SR�����J~��t�g��ǫ�����V 	���r(�+U�-Sc�a��ڶk9Ѷ�� 9#'к1O� ��^��`�i�˄�ւ�O? �s7���(wh��{��5�k@P{`kd+U���2)���,��R�6�`��{�=�w�Nv;�-������~�~�~�~¾-���]�Cii���ᕶ}�&�x�}��zi�RM���8��!y+Ϳ�(��Z�爹������9���j��P���]�-9g���I�
7�Z�O�
:���b����d�$�ҏ��
93F��#��Lh�>:!5u��%�>�u������zc8����\�� F{�ic��>܂�)8�k�;�	gQx�f튟!��{`����,��3�.�W� \ꥷ�s<�[χĦ�-z8Nzf�K2ύ"�F2��-I+Ϯ�����Y�*�NI�����q'�ss#]�Q�+�R�y:e<s+9��U������4�*�X�ӊx$�
���+ca��艹w�.�Uvj~�I���R@Ե��"�<te��YBjDn�dEUش��i���Z|`M�l�d�����tGTyR��6	��|�#ɓ.��4w~�I�w	3@�\(:gl(e3&b�����M��$݌��'����H-��c��
�tmH�t�А�ѼI�A��'���,!�H���suf�%�\�fo�i&��+�Yh���{��B�^��>�m�~n^2�}�����˒w|~�v���O�Nyj݀�Lj�eJ��nTF�9;�Ntҵ)��^�ud`���v�̳��� I#t�U@�֜�<���l�T�A0Aɦi��Nxث��@�_`��2%i�Ś�3����Zt/��3��^}4�8	���y�sߟ�oh���	氦��i�ɰH_���nI���y��~�����]`jފ�Ew�tj@R��������/����xh����g�j1�����Ԧ�"G�s����Ox�߯�Q�c~�鯋��=gݘ`���m�����>�������Ev�B��\���/�-��_�Ҏ[��']�!���.�X���w�Pc�&2,��cbS������qp0O���_Y�B�=��xFƅ����� ���DHj&�i
yjW���q�#�90��=��m9~��\�\�G	�����[�dT<��!o��LHK�7��s��k/���� J������q7d���z9��A��ӡC`<@2	�! <�t��^�xN��O�
u�B���ȣ{_}<�	<z��z�=���2�3/&.�~^͡N�1Ϟ,X�X��h�%��5H��Awũ��Up�d���$��-��f�B�Ŋ��R/���|���Xѱ|��0�m��%��[.ZQ���C��T��~��T-�qr� ���9�VI�-��-�cR@8 4�Gʞ�֖��]d�7?3�5��ᒚ�I�l|U�9��byh�q^���*�Ѵ�����"�^'����`.�{Q��D{�T�	���S,1������:��(���_aOJ	~|�J��i �NJ���[
�Ut�*Ũ����JA[p��,���(��� �!^�k�Ey�����5�9�I�>+RE����8֪��S����'W��_�=h8���*:x�b���?)��/Y<T,`x�!I�w�0�tN��<��~'D%ÿ���ʥ�]46;x�*�$�ީ��$�3u̒B����0� ��$����~]a������n�l���z�u�n la������"�yv3lҶb-*f)q[�B�lJ���̾cLu����>�L@j���ѣ����y���a#�W��9�_���l�l�-%#@��X�!�i��.��A"���B�R���p���0�J�$S�aD+���	�5ɲD?�<�����U���F�<����-���L�����R��6`��vz�VA ��8 >�4:9@��� �h����а�����_G��m�
�.���SQ6LxX�<М��:=i��xb�y��֋���c�ۿ�i�}�ޗ��蔝D�+h�~�Et�??(��[��� ��|R�)~n1*��z�m��O������0���H8��Ҁ�p��>�kj�:�pљa�C�mE��w��G�+S�K���a�\Z���~E�O7"y����S����o"��	@�87n܃lx�޴S.'�O�u��_���{N�=)�v��H�j�΢���B����9&��@����,Jx9�t���������)�w�r��=n��وJ�	�NJ��ړ�_4�~B�'�\/7�{'�G��P�?�gHK�:�n*tj��/q<���P�[ժڋe��΢���Kn�!��zpY��?��ԛ�L4C;u��n������(«v0�Jc�w�����x9�j�OQ��S)�yB�aL7���2"nGS!E�jy���oZ�v,�22!���$i�O�yr�}�D��~�ӳ��!���Q��%E���~�Y���!�N��R3#:s���b����wu0P\��y������$q���?g{4Y̐���;�"{��+�c#�Rkǅ&'�#
XV��?�����wG+��������� �����!`M�b��U���1��j���>�1?���;1�-I�׉'у����e�䒁�GLl4���i�(��hU��,���NpG;���МsO��֙v�$ԢАoX���T%��"�&pm�����5�D�8�έϏ��>����ı����@���DⳲ�MF���t:�KoX������cx���\1(1��qi�{�x{>YL�]+���qKSy h $|�5�`e�gIpX��_�Մ���Â't�H!�S")��yJJ�[4�싃kp3X�1{�~�x-�ͫ��wm`���6��9�#���C'3 �!a;�����s7���@��p�Pl��G_bN0(����d�j�޳�lk�:���_�|)ICt�Ev�������i��(�A�Ӧ���ha��w&��x_^��	��Ə���˭�K��yY�=%'}��6�{�&��W�t��ҳ#�+��;͆EƬ��/�L����sR�BK�E�A����eϪ�dZ�4r�>���,I/��h�@����d�����_GG���G���B}y�"�YZ5��ߩ��[��k��W���3���`|q�j�t���X��a}v�ZR�(S5�$�X�ya�It�Ɋ$W �q�jǧ#杽a�n�r���E5����_���9I�����Q��%�6Y4Fs��l�A�D����@��>2䎂<�� u�+7��q�����v�k�F% �/#�6�K_�z���F�:�[
x"��b��6xzُ��)���+�L�M��A��~�)�*m�	�ƴ��P\��z[�.�&��	
;C�3��mS�O�񰣬�z�8��&�pvL�����������& �p�x<kc��5	HY���}����4=��r�Z0PD�?ZwV��rU����8�5��%Y�WE	�b�hX��p�8K�~t�t����ԓ�ܪ�����b=�5)�nwi>���X���x>!$K��-橍�m���������*�0|3_��{#�*��`T���ۿ�&�O9��4E��e^0�P�:�)FS+_Z�7<�a �G��d$����<��+�y�8s4L��}��>I?Wk+_G��oZ����K��eͻ����I���֮9W�~�T��h���WE�xm�v�Q�
�x���M��� �����#7�����v���3�W)E�����I�<����DX���#�|�%z6�ΏվH?t���GϷKR~�*8  0ef��8��.ɍi�7�@�?ֻӦ�����B�,�3��m*�����//��|��a� �݉��ʉ�!�-	B�:�2�H���U��k
_�ɚ�8&�C0`j�1��|�^XX����J�
`�J���� ��}�U!��-��t�Bw�_�	SX�"���]z�[݉�<��b �b����%gxE�q�h����n���}�ȗi�����K�����˱��Y�A�<TNnF!��Ժ6���-���/u��g�-0Y�y���q�5G"�7�Ϛ�ra�Ӱ����¶��w�mW@b������wVJ�S�n� _�]�;g�~`�s���P�O���=;GB���-P\�'5ƈ��c���Y�<ݧ���nq��}�7�o]U�wio�������,9Rv���bѤ?98yn������M�˕���Ծ��{v)��G�#;���{��=(���~��������6s��cD�&�}=?}���7��{� ��	��������:����Y1��JK�(��;�N�K�bnE9˿�^E��>�	����"1qw3�W��/�V�Ԯ��V~����9h�K�p}�p��'��_UPiGF����mZV=oB7�'a�A���m�{�k�2�z�U���;����9���&�١�i�D�?��ͯO0i�OOv���*�U�)^��4_�(
j�b���n��^/�R����q±�lp�֭�
��#B�H.�F�\�������G�&7g1<{����Y�>��tz̼S�ӓl�r��w��|!�m���gN���Z$~��|��!.o��i�0�$�����~����M�i:�N�����>�������i.�����}hcp���6�Bl�ɑOAJ����ÄE��m(_�#���Z"�� 	�����u0		K�����W�[H ��̸f����P�N
�������9��0��u��ǡ�3G1���6�!����4���D�:�ӎ�sx'��D��֝t���t�c]o��w���|Y9�cb(���;�s��˧F��k��A�u�>$&V�jF_c�}/~///L���Cp.O7��\�ĄW��y)�B_�,�I�Q���+�5�U	��t�,�����UA���V�V�b$m�zֽ�,�"KE(��u-�$�T4]��.�ﾉ�F�5W,iNS\7,�-�XM�шH�hP\Bs�7�W���e�YI�����_ 
{���+.�H�m��/`?����[\	����܏;�L��q4�U<	��P��s��%W�9�2�\H��j;��#�9L�,vǒ�M����PhumóN~�붮������]��Y�¼��7�_z�ݏ���ր2����얧�2R�����)��QY��4�>�X͹�'BU����C�V3�V�4����o��]iȏÔ��ُX.���I�[m��u�oՋ�y��	&޺:�?��))-�#D��^�|�[�c�C��kj��G��U1�/V�ws]9���4PE3���3C�kX�d�`R�q$��0*G	����V�M�ɀ.��i�Ӂ�����?�Y4�����G0���x'q�Wﯩ�&��3ވ��[>�7^�o��x��=cB��X��X��%�D?OEgb����5T҇����f�PD�N&9���_���?�n��`0��!Y�����}�-fP�}7�J�$�RQB���,I(�eI�P�P�|{����׹��<��uϽ�s���<�z��<6얐T�t���a%v��_�oG=�w',����㾀,���'�Y��������a�AY�����bbY�8���!����:(�R%��Wd1,Q$���qb	���°�p9&@�)k-�9�Z �a��G_vC����n8G�����P��U�\��w����������/�'�j��'
���>�X�c^׺�
�=�����W�=���y�l��#�<հ������Jػ=D-*e։ͤnpl�����&Ed*_�;!b�������{��0�?|])_��Ͼ���v����KC�i�s��YR������m�Q��n�:�-cS�3�~�'w���l�z��E=c��hY?�7�3U��Q�)�tcښ]�&�����ԹHL��YXl�v����΋R�$؄$x� �Wkl	��Hx=7?ץa�|+�y�R��fE�B�k�9>��m�󊭟׼iD�j��1\;~���͗$~�П�
�`ւ�V,�M:����X�T���	;��e�M���#��oXH�!�_��<�δ����HQ��B��0�뎣����u?>��ֺCRo�T�W�n�t@T>Od|�*jS/?>'� �;/�;O>�F茖�:���ٲ� qiJ�5�1{_b����[T =o���|�aK�x�_�����0�W�|��~I�_�Hp"g߰	�Qn������v:.��|�]�^�?�нo�������&g n��E� �u0��]݁ʽK���0|Y��P�������W=��*���S���N�Fnd-Lv������Z��w';���.A�VW&�خY�A��.�V͉z����[ˊE`͵N�	�7"mؚ�b�6�u��[������X�#�g�ͩ�	C��������wd*�}�ݕŸ��S�t��)�>dK���nB3@3�9�xZ��� ;ct�#��*)5{����!��I�\
 gV���k���ĩ)��'&�]nv�Z�3s�	��G��$;WhZ$x2М��,�]8[�7�ަԲ�]F� �IA�کm��� �h�4�Ή�3�n�Ń=�������{��@���z�=�w�$��P	�g�oQ��HW�0�!>��H#ߡ�v(C7�����_]�g��fas�#�<�И��mt��KP[T}��H;�]��YG�>�d�e2-L���vV��;���[S4����+~�ۭ�nov�+�{��8��K�[�Za���Ѐѕb����\+]聩9T)I�4�)�|�G����`�l)�<+��T��g������J�������"���v����v�z��n%�܇_
�	����
� D�~}ۢ��������|Ԯ�d��>}tw���2M����
�i �@�nÊ'O�G�#$���h�*�!(}ܶ8(��8����V�4���c�U�$��5���@�3�� �@
6*-�6��w�����2�6Ԩ0d �!�$=�a~�4do�B�:Snp���x��ŀ�#_3w�� ��C=��.��xSۉr_��p�����������$�E^����T���GL4ޟ~`w�̧3
Ɋ�U��Ћ�^�lLK�<2� {㑈m	5�<^��t�Z�l w�u=o}?D��G���>�1À�hmw���Bٹ�|���{���=�Z+%�
�����@���Y�5O/Oc���� >�@}�����4�4�Ror��Ch�ٮ�������|�o���{�� ���S{���0?�Ĭ�G5��ej����y��C��xm�u��s)*����2��T����ц$�'#��:�y�~�Ǒ�E+���2Z�ŀ��u,�\��#�r�D�˚�k22Us�7�r�r�4�M��Y��d�CkL#Ռ	�D'��Ee?ap���n�}���t����"�_GC���dЩ�9��u�)�����3�=��wӕ}��c~mt�|H�^|B/k��	$Uh=�����⵱�VU�A��a�?��Ћx��8�������Ĕ8��C�20�O����d��������gM��t
�� 偌'Or��ը���A˃��RF[��@{���)q��L��`�1��C��o�3�?��y��M똦^q�4P	��q�Y���ڬ���:t<]���y?U;*�+��������I�hGa�s�h&��Ȝ�dE��Bj�r����V��9����0���m�52���}�'ޙvJO��3� �Wo(�(������d/��v�OKb~�KԺ4yԐ[��|s�)�cUs��������S�)�P��o�D� �N#�H^Z�C�wG>��=�^:�g<��uG��Ӄ�s��F��2?m� �m{�=-(�������Wp`|~~tF�@e�r�q:@������Ѳ0��%�ρ`�&Mhe���Y.1�͍>���i��8/��2xFV�%,�^�{���������?�4�&�JD���Ǘ��ϝ�q�z^ZRl�����������ϔe�ɸW������/l_��.L���m%��x�| X�sGuAPE<޵;X��/@$�)B�"TQ1�A�������mߒ����G�̎h]��`,ᰵD�WE�ޓol���9��h�B����k�5Fv��* ����� h�:H!�5_��C�8_;s�nz����r����^zA�l�ӕ
K�}��=&�����I?�޼@I=A�jP4���]h������:"�Ī3
��U[i�c2�6F6>�i��#Q�\5g"��s����wU��Ϥ02�Ts_˿���?��>4��.?tl�c��w���`��gV��S��";�#��k�3����]���*=E��X�l˅4�[�� ����Fj��9�e���.��}h,�K��:D�<�G`o�b�jb1�:,��}��(�BD�+�7�#��P5��	]�B�o����+ތvs�?y�V�h��]�N���4 �S�wF�ƶ{Ф��#,�T�>\��M4��b �u����_;7\� �j8���L'�Q�'MF�on:!�6��>��O�IGR��2�~}ƣ4�S�~?�� H܏���X�Ĥz�����l�����vs��8�y&Y��F1���c�%�ް�c�b�@T�UCw�7;.�����K`��3����(�qB�H��+�^��]�>S�*w�F��q�*`�i��?�V�wg*|+<�Bǭ~�Mle�XP��"�n�/KR&��ǆ2��t\��omno:. Y��âF�?�-..�M�"�5�o��>�l��:S	Ѳ�r�������H���5@���pr{���!dL.��K��r����hFK���鍇�!��﷈�Ⱥ��+,-�����������D��{!�C�9nw���/�%c-�쿅h�q��GC��=>s$��a(�<�~�2ݟk�&>��i��Fzk�q�?��a�2����0�=��ј�d�|�Ly\]85��! ��T��k�L1�x
��
K&���L;��������A�7M�6A?c�ϖ����>�-�r �0����ԥ;�{�Py1^@�O�ð�i�=�E*��>\=�0�n���r�TZM��慕�"��I��&��s���x�b_�4���;�Xw�aO���?I>�WA�8 fT�RE�[pZ쁳��8(��iw����˄b�bJ՘6�@s�S�E��(�B��ڣ]����NV�QԚ��w��۷�VAי�K*[�A?c!cT���eĠ�1�	�O4B
�6>��!60]���Ɓlڑ���g7�r�������k�k�*n�i*�;W�5�Ŧ�+q�x�=��2����B�������7X�i	�LE�ƴ�R-?���~䗫��a����6�ϗѰ��G1e�}J�_�8�>W���V�͉8�rw��."��/$t�4};_���Z�Q�H	��8���A��Fe������ʦ���� ��c0C�X��ŏŘL����(DY����'�wG	n�	dp^~��!(T�~̠m,6��NGQ�����\���E�������2�1?�6��S����� ���qU�S¤^�t�yb	�7����������xE��Q��,�wW%�
�68��x�Q�ێ���q��wKI{L�R�J݁w�"�
����o ]!�x�2����߮b[��*j\_�"���t:��ig|(��1:ߎdt���@��]O.��M7S��M�����X]�\f,HN�����nO[53�۟�y��UmwI��nZ]7<�k���H��~�hR/s*�.!tu�G�cF�A�� �J�����h�_�q>>�Z�ĖO�,�[Vȏu��))�6z'\�
�έk���h�ڻcm�	�n��Έ��/蕢��fs���-k���u+K�K�t�֘V�Y*+S�G풷-�aݵveT��RF��eaC/�7��g�z���ɩ�Wo�����0���+�ٲ��=\�~qteR��/�D�l�SO
���b빿�ɬ�$��70?ӴO�xw>t����� ���r-zT75l޷J������!��8J�T�/h�I��|�)�oǦ},�r$4fB�>x�})Q�Ƃ_�ܼ*����~yF%?(��T9@�b�1�Ds�O~�=;��A��ih��Q�j��ֵ�Ԩ�A6�����3�w���,�l�9��$N|�z��V���{Pl�l���N	p�<9��΂�y�v����t�%�����¢}�*��$x�a'�N.��/G��B�[�yPu�.�":+����A���_���\S��*D5���B
n�I?�X��z�4�����މJ��;"�=�+f����|?����G�u+]��%q_~�A;�f��bv�ҧ#��Բ�}ԩY�C3;ZGC��b���H�̴'����ɸ�}'���E��Mٜ�n�ҝ���3��Zُ�Z����7�I��d�G(U�n�Q��ۣB��f�c{�}Ҍ�w���"���*�j�C���j#D���Gm��c��.Ѣ{���([�.�,��\�c;S���{�b	�C�$5������A~����}qI��E��߽�89O�}�y9]�� @;=l+��8r3o�Zw,�j$U���?�����K�'>�	��,.�_=Tl�С�v����d�0�����0��dh�Iw	b�?�(����a"h�u���Rv��p�����a�1�T�\�+J��uCy���E���Z5�e��������u̩N7�n�zȍ��Ld9�P���*�J�z��1T�C9)Y���h����7�& ��ٴ!���3�i�<^ �9� �)y"�w��s����c�3C:]L�:S
����y����IB��)�P\p�z����}�9�"�Ú֟#S�؂��<���sxcԅ�C�<
ٝ�$H���U������]�Ş}�OM��1�}OȮ��3��;q��H0����vI�q�l3��=O둟,�+c��P�<c�������������H~�X�.��j#Z׉$y���|Y�V�_ʏ�o�J�!�N�Y��G��9��� ���#&"�K�H�m�~��ke<e_Cc��g�r3l���ND�ٯ�/���^vv0Ė��BH�B~�<�*���]�oV�[:�ۄ��%�٤׋-�1	 !`�h�uщ���}=g�a]ʠ�|���EܹA���V�H���-?��G�[���'JX|>e� j��l��H�rz�I�l9�A�X֧��׽�X'��/��Y�����e��9�~��[�J�]�)f��Dw��̸�+�ggap�x�#��;?;Av�zX�/�H�2�.����`�B�o�}����r�j|�_�������yG�R��;\L��p�[al���i�_�D
>�
���<c�4����'٥��܅p�%���'��@)���=�=i.�Q���s�cK��]�޸R�S���O�8D�<[YC����m�mN�W5FZ#��~��1���ZwZ`��E�?N�����J}}B�y�������t�Q�_��G/��td���z^o`�?lu���{�-ʬ�S�O`iC:��8nx��V�V\�T[#��(��%'I�	3��b��{���g�K���k�K9׶	d>[$�k	�i~L�|�r�#�]P��+��� /��A�� �歜U6X�~_�˫F�Q�&���4(z���(M䰆Ĕ�`�~��W�b{��{t�
��q�P� ��c��U���{
A<�h0�n2�\Z�A9,��s�Q���&���1�k��^;�Cឺw3��D<��FA�	d�1�������b�����]U�6�fB��s���}��Q���y�� �7�u c�`Y�n__~��%�8K�.�5i@/�D���|��/���8�"%�Ìv�W&3\rwh��Z<:���3�v�\R� ��9�>j����� x�b�`�P�8J9)��b{E�R�
6�e�_�w�Q��������)T8%;����f�[�t�m'@ǊG���"�E)��[��m"�1�~���!x-D����Rr6XAj��K_�M�_���@߾�_����Wt6��Υ;ie%�A�?�ݍ
*7W�0ك,4&�褂�x"��l���w�(��/�|i�V����}��M4���zo�<m��~s���J��M�r��,��lkI��L���î\�X,���W����� Ór����s�S�Q��S�Ov���� ���|�W�?� ��?�Ba�QΧN�9�=�)u#k�߮��M��j'\�����Wb��`�Q�C$'�y򯖓g"��`A5�l�]i�ͅ.�Ð�o����yE�W��WM��vƅC�LyU�K�%�m��^��P/X�i���y��~Aֆ������o|M�f���	~���Ô��bvb���Ց��.Z��t1Р�Bi"���!��`�:�r`�,�N{����� �"�|��)�K���ꄎ�?�����3��dfa��^��$X�*�9_�M-�ϋ89ނq7�+��j��͠K���j߽U�O����m�~�n�HEU+v��!_��X�Y�d�T��4r`H�{��c�ݡ\��/葚�'|�<���AP���Y�n�R���hi�EA��F4������
:X��,�,����]�i9I4����Ŵ�JԈ|��D�ӧ���a�f��_���8��^����,᪔Ԣ�YiT`��a����:�o?{��ﵸ9~�?�\l��	����ġ��h�RD���g���{�.��!?����5�N@���/qf�l�~C���
������q��K��Q<�����p&p"/|n�ʥ��}@�&B���b�/�/����j;Ѧ}���4Ku/��F�eAT� �E ;�<C'G�y�����Mc⅗nm$F�x^�UvP���w�I:Y�A�[�<�?�~y��!����yw��K�H���8��#4�oݖ��a���{=�B٦u\�r�@�ƹ��}3��#x��฼k��wn}� ��.#�^?dSһ��1�r�?0଩�hpG*ZᯓϹo��g)�=�z~��̼>�Z�{a�Ϟ~��m;�f�ĩ�����t�(r���^S!�e�d�@�0~YQ�����k��²�'ůD�IbZQ�'�`�Թ��y:�8�tu�:g�\K��u��y
%x9��T�,�́l��y$�¹��o�ڀ=ܗ��LV�4��lQ����sk��`/�l��.:Ue�����ua��1�Z�խ)(��ވoЎ����:-�L<�0>�Rb�l�~O�\�}����0�뮭����^H�${�:���������j��uMp�,����fb G�?�Ձ��\�	d��7���H:��b	�'�5��|=]o���mv�jt6���K)�pe3&4�$��1�������aB�j"�)'1[05�5�y���y��H�3�$= :��3VP��`e�l�x�ne�w�"���h���vRrN������\�ɻ���&�#���5v�z�_I�S�HjA�����.��{����|+���_�z���g,��~���gO߃�����Y��W�t���]M^zh�.��0�Y��-g��Vw__��6�.��RŒI�����~+�c_�K��yp"� ��6�n�aXģl���r�E��ƚ��U�ě�lװ������r9�Y:��˕���	���*�����vOd��/��	��ǹa�����LP�'�
\K�*mC�#5�<�>��X/2���^�Փ2R7�?�-9S�e 9 ��K�@l_�*?�M>}2(���a�4��(F�ؑ�I�����y�ST@u���`0�h7�T���(6�|��(�ܑ�H �d��� �8�S(�F�/����)P��"�1����;7˨xг��y��˚";@)\�H����@j��|�n�sNE�U�TϘ|Wz,�M�~߹6��Y>3��7�
}�z'S�ٟ(zU��#�g�?ug}���^1�^�2L��<������ӌ$��z��}����5���#��*r�O�{��{!�������O��Y�> �*H�螪a�*�QR��x<����뱯\L��]��Y	[ِ�X˔��C��]?SЎ&Q4������.61�,�<D,X����R�߸'�2,�ՄPu,��hXT����)��
���/�6���!t����F���-�ot�:���ꗣn�`�b(�G�4�RK���ա4�r�VI�H}�TM��q��@�J#�A�j���]t'�Gɉ�cW��U4��l�b�n�[<�McӉ��,�r9�o�_S��I�3�ч�+.���\d�l���U
�`t�A�w����nt��ї7��:RS}�z�j9;o�j���e�ٷɏi�m#n��:Tc���3�WI�\��l�O�����J�d<��J���կ�;p�6����I,��ۇ|l R
���J����Z�W���ޡ�Iv
�����Jyj�嫶6�Z�qۀ5 ������1�D����T��-G,崁��N�������x�ݷr�W �.�x�@S���c�����r���4|��ӗB�o�J<*�Z"� ��A�_}��;�y����;k9Q�k�@I$SN��� �)$���)���\cU��'�E�jL�Tp����B��>e�.6=8C���箅�żd�{�-?�V�13b=�j�6]�&=�l�qXi����o�9��*�݋�5Tg��՝�m��֭��M�E�M��j�e��[xlk�v�\Y��(6��U��6�xUt���.�{�:�P�$�Z�g8�4a�f�:C�4y�۟�Z����<jT�b@�`(*̉Y�Dq��$�0uzR���`�Ws�6�%�_<���m�<����!���;�[��	�G�?0�w�hd�(	���[�d��_j*r��M��5�=�]]�@�B����Ǚmª�����MW�d���s��"!k�du�"GU��!�����������}�/�����?3��ߠ�va����a$?s'מ�%4�A��V] mp�mP�7+�����
N�K�+�zEa=�SF��F�w~���բ9�*���ɲ����K-��/��t.ge?���w��d���|R��=>a/�J��K\lNC>4F4S9�9����kBz��&�aaK-,T�r奋HQ�J���}Xq��ǒ�N�@K(xy��A�pB��^����L�$��d���#u�;�7��&��R\$h��d;�❵����	�LOo�J��h����j'(.� �T��z���m��.%v�Q�6�V�n�±�83{���7lIƄO�>�E��i�d��ٲ"��E� �U-x`�-`�MKߺ�N�����ML �{��T)����WG�t۫ǂ�/�}���r����{
Y��,1m�3^p5�%����:c�8��@��J��,з�?�$��ܬ���kwm���S;l�-�6�#/��1����x\YT��=c��r@G��8�i�%}\9v.ggŒ-纏��ߧP�!C���
qcv?g��DpQ�hT����2�3���I㥗'p�Ƭ��wE?�x���%�F�aY���TT�bfN�z�д�?��&#|I����84���R�Nwt�[�x]����j7h��tb�2�l���[m�Y��ڌ_��SF�{�H��\��<XԎ5��#[��܏��"̣[��o^{��)��q�"���R��kr*ÄZ|�2w�Ŭ%����Ώ��33错�=jW��n'_������ ���+��zQM���U�=NU������Ⱥ�����@�3w��\����O��,2<���w��Ֆf|�}�W�A�Q�N��ZG�#�N��xk���?L��6e������7���*�ck�B,�Y�}ݞ��^�Qdn�o�8�Cv���y��*��ي}��wa��Sg&E۷�c���
&��C]���Ǵ���o��ST]3�������l��}��v`���_���)�}�����4��Q(5*3�bg{M����Q�����Gf�K9x��L3����<^(�U������#I���
��A�Eԇ��E/fo�����|� �g���-��g���v���@�� aF��#с�;/׹�e�H���C���w�,�.�՞����-��x�p��N���uu��4�l�r���_Xc��尉�	>����Qx��7�o����F�Ճ���Y]�[��U��TwVWCkx>���_��Q�A�o�_M�A/�ǌ{�j�/����!�1��_��r����t�j�+l �D.�r��jo�ݺ����[��\��؛�Y���q4+\���w����7��x�,���ET'�.�L�$���x��W�����$ۢW����D���?T=)&w�j������CSi��"����,��S�=��/�Y���̉;��Ke�@X,��o��a���흨���4���Ԗ�ᜬ�q溹�
~agW�K�R�#�xAY�צ�e!� \_h+�w����S��i�_W��Q*q�c�R����>9�����<6fփ������I�>�,�?�V�s|�Y}�l斚Y�R���.���:���ndx;2��MV�Un�=W U���s?��<X��������V���Xy�Rm�{9yB�E,L*�m���h�18���J��kݤ�E��%�RX�Y����HwE���z�(5,��2�9��>�d鏆J��
�ɿ��n*�s���m�茤T|�x�}���E���r����u�dũnHK��2�I�7����VJ�����kq��=>
�,�0�Nt��ߺ�J�+~fy�퉗�� ��!�o���-Q�@GU���\EՌ��%U���I�%�ԙ)3��Z�/�0��A)?�N��}na|cs�8��LH�d��L�s��'8&)�F2oA4i�6á�2���P~k�&(��w�Zw�-CX!���3|R"���,[h���-4=�*T�лx�=3?��Y�u���d��Fv*~}�hs�̵Cg��;�KI�
kb�|����<q���\������"�Ґ}rga�������o1�+�|���1����q��|��5<}g��6--su���{ϴ*6~J�����< +�w�Q���͍��o}~��I�.mP\�&��Ѧp��Ƅ���7.N)�$!v��g�JZ�K��o��k��5�v�Z���3Zيh�ܖm�bn�'������p7�)p,��fD�i�Z��q���Eo�"��\���W��b��@��G��G"��0�y�0����Q�)&ȋO7�%;�S�ss�ʯNֆ�͒���c/l���e�YOn��ug�T��-_�Զbk?�O=������wy!M��]2S�A_�ތ�S\T�Wp�E�c�2n\�����W;6j�0Dɞ�g�x?��2D�O\D;\1��y�ȓ��p}~��g\�R�'y�Ú�W[����<.g��f����g9��r��׮7(�a����Ta>�Zܧ�{qU�;�\�o^ϩI^?�f���I'f�u���@��(r��pj�W?���G�»��Lƙ)�2���Φ�u��nle���$5o�� e~�c����z�"��v�,շ���{��츛.YǞ��*�3Ut���N�.�T��mЄY��#7���r� ^//9:�:��Z�}Y�a;b!����q�p	�(�uq�u��3��E��: �]���_4ڜ�r1�|z�:�ݜC�Utd@���_���J?��:��2<d�\0gޗ�#=���eg���s䱛��fk��a��W��BR���Q3�ف�eG��[��o�ի���^��̑Ϧ^��{�z�9�^�w�8z7�[,��h�����u������aFJ�_�:��>*)h�ƽ��-M��V:��V��A$���^�y|~I9��A��SWdj���k��Μ�YGkP�o9sj��������&�Hs2Bh�=20�d���߻%����8�sk�8��W��ckOB�Dj�����g����JI��-��8�:�������/a#�x��|��C�IwN	*�:Y" !�rv���U�GUW�A����jE�"�USN	�g<�a�����XP��؇�h<i�x�,b'g͡4�����+B��%�����P�)D�K�Q*�bgK	��9X��t��LWIsk�y��ĳ��*!IB�i�x��ut��x�4��\�k���3�B�㠊9�rϾߞO�8�n����6����"�⣋�.s߈.�����d��׸u,rli��kmR�uU�KΘ�:|�|D����қ���f�����~#8o�<��eUogC�3ӟ�o+F;kƯD+B���� �	�ODv��0�%K����#"$��T��<�u�r�ֽmZ��~�����1��ξL���A��)<]�vMŻJT׆���Է�`B U�pН/ x@Je��N�#
C݀�qRz��c��@���>������半�_�ח��j�%%�JN�諬�;��	�&qBb��2.7#]lIuD�z�nƝ�O��P7W�X64�6�W�E��flv�kqW٘��}����d���lIM���m~������~�#��d��_�� @[���	^ij�LП�
p����q�M�i��N����EB�07��R�V�i�&��<`@X<�����D_�vj-�n��gykB�iঃ�t �{ �	�}Q�-�6�uvi��Yq7��>�F� /���zN0�5��Z���[�
?�R��Y)�X������X�N���i�����<�(w�}P@~���&}�&�x���G������eZ>O�������o�������R[�E����K@�t����U�M��m��W��=��W�X�9��Y��1��w>�=�Ux|�7��N���x=(�7�~����QY٧��C6;��5�܏W.[��?}�v��B�����a�`?�O�Y��2Z��v����3�`��)�� N�!�p��a#Ϡїp�(�0�^M&,��8|�ɜ���z��s0�!��"l�d���~�4z�\\>�1mW%�}�C+v��1������)�j�I{'�K��p��O�3)��;>�[�0�pi�����v��ߕ��e���.�������tHR'&=��>)�b�g����ň?B$���1O�W��'l�Un��+��������Ll-��O��:u����?Uc�����[롍����?ј��ߧ���_lɲ�S��	�;���%dA��	'n���p��6���O��M���%}S����q;��0[�[��g����g��`GCȁ�tSϕ�3�N O�����o��߁�,V �(s��
�{М	�F(FLޏp�k�p�u:9H0	��>�c+������]��z�{ �3-8����� �$M�|�I��Iv��/��	��^?.!��)}# 6 Kɼ��vn�j�:�bq��XB�Zh�3�^���`0�2�n��O�\���D��f�M|���������4���tz�?]?죒�+ ��O�q�@�	��g��@1��K0T�$���*>� +.H����n����<=�R!J"����'�����qQ]QF���耮��2q��!}u�$w�?�__�^�ھ�� �ݳz�n���ؕ.�Q���I�m�1�Bi4-�~- ����%��}nP�Hz;��#b��"�B,cBc��w�T�U��F*���0J@���§����yf|� �k��_������Yy���1�I14~�ǭ[� qǐlbHp�s���vt��-< ��Dw�&���au�YP�K�Ύ���i���!�G���Y�
���C�Sh;�����<�� V ٖŊ��:J���#��"�� �c*��{�2�������uv� �W&v6����ߜ�͌�m�Y4+�������ct;.���f��ԟ�$b6�qL�=��(� �9u�� �u�c:���-M���3D�m�6�܆ېh��|WH3g���B��Dhq�9��!Q���������<ӘWf�ɤY�����d>����1�=�%!���`K�� @�3+	�8�A�TT�}hjQG�u�MD ��T��e*A��V��P���t��~�m@�iJ�Ƣl'5'�\*
Ÿ>��M�cJ�]d�	Vu4 �=�Ƃ�y�]E�X
�������Җ!L!�(���E�jz�Zj�,��L�Lj2���q�;d{�h\p�wHX���"HQV2�4

^q
  �P  ����y  ���o,���A�P(BM��K�^�/��&� �<BT�8U��2��-�8�IWs��;Gg�|���e��S?��/�;��mlbjfnaiu�ך�����?�SDd����|���������/(<}��lٹ�.V_��v�F��[�M��[Z��i{�����i_��೗��_OLNM�,-�]y�����O_��x߾��w~��k��Y�i턷��&	S-0~C�!��_��#��ѩ*�����X��7����K�_��e�s|2`T���Z������3 ��D> ��
�2��Z�y�6Y�?>Xx�p9�,�sgw=��r
a!��a�z����C���2ě�YCYs�ӭX�{6+dr�4�?%k̎�m���r��J���1�d�<cx���=��~! ��k�j��������!������/:���_L��dsu4*���;�}`�c��/48"�/������3aDW':9��1{w������zU��^R�DWlU��;l��H�m}F�&�:9�5�/*��o���/m�>lL�u8E�'�uK{y���c:n��i0x����zʇ7m���£B�4A�_/LNJ���@E��E��$��[v}>���@�s�h8�ϥ�(8ڎh_ ��Hp	��_���8H�	ެ�_K�i�~'�%�F��4-�M4H�L���4��Gg��q�"E_�����q	g��tUS��v�g�ȣ�^wP�hP7%LH�fÿ,+����Ma������N�h���O��A
��MjM�闣>g�(��e5��T����=�ͫc�T�4�}��f
��)��C�m�@�0isiC@��!<�T�MP�J7A���Ynd<aSy�7����D)�I��!�g6�)7Swy����W���l&�k�ڧ�t�?��v`���?���0pSjl~��[��^�v��nv3
�%�/�e��lv����7oC!�����=��� T")A�PD��k�-��`��?	U�x�QV�}G����-��Ѓ�ؕ��C ��7�)�i��P)|Zd�*��=b��
#��Ԇ�XE!���~3`�8{�t h�����h)�\fPLg�p�7��:p	#|���l�� �ah>� �@%5(�	b���>ʿ�_��wn����F��0 �٥��c+o��@� ��A��i�� ��C� 4
"6��g�dŶ��UppX%Ut�xv�^#U����	� �3�3�-C)=�5�Ѡ<�����}p7�kW�֐�۝T>�����d��th�"eP�|�h�}BzM�Ic�{F� ���®�*MV��c9#��� ��a4  hx X  <��V:�� �rR� ��#@%п� �/�-k���WRRR3ˇ�g�p�X��=�l�F�?[��'!tg�����MX�?��
���^D�_�U�D�g�C<4��&[Ń		(P,?�P.\�-K�,[NbJ��!8���&�xԃ����MH<�p �& ~�@[ѐ���ٙ737��}�������t����Şe� �͉wvi�a��blwg�pB�AR���jv驄����ؒ[��߄��.����/��	sCY�R�n�V�F6��7�ʛK�/^�>��6�ܜ�ǕO(}H��ze�G��~��&��[�ۛiTD�\^R���ٸ9۱7���)� �}�m��B*��;�$�a;W�-��EMk+��s�E�B�k+��ўђ�*��ښ�g=��ϗ��@]a�,7�l\�K���AnHNj���x�Cf�+i�'��#�WXn1+Ӕȼ<��F~
R?�� �A�Q>���J�������J���� n�:A��
�Y�P�!�H. �"��_�>��6m8â�����u �`%`�r�Q�%��u��(7�Ҁx�c�r�^NW����>@��e�:��1�8.x�sVkVE?����S�a7�����
ƃ<�-��J:�V�o�}Ps�0?@c��*��Yx�6>w�wB�����0{�z����_+�C&Nv7�{���k����+Jϫ�۽��7���/�+D�@�[F�>�K��M@�Q���F0n�ҍaܕ���������b�^���������p]�T�΄�o���\	���pC�D���q��p�\!Y��D��;Q���@�gWM���T�&:�yR���N�j�#�6�վ���e�:"�&� 	㳠
��3�,�ژh�!�@S�5��u�B�(�6(��F��������Ӆ�д��.��Yz�H5 5v�e
gЯ3�Ve��N���a�T �f+����@��x��xSU�8~Ҧ��BK�V����b[C��&�GKJ��j�'�ږ�4�a����2������*���t�8�zbP�v H���Z�$}���߽�����[9g�_k����k�Sp�!Z=��
B��9¿�U��������_U����U7�߾,u��ŷ-����y�,Z�XJ�uA�RϢ����Mu�޹x��a�zŧiy8l�0E�8��n���BT����(A�	B-����L ��'�-���-O�^G��UQ��:?���\��S'��g�N�Z��6�C:!5^6넅Xv�NH~�
�G�|�0i�J	�W��x����]�
��a�o�n���8��"v��K<��aK�-��'�x[h���b�,\�M�6�XuA������_�K�]��f~u/  ���� K � <�� d�: Hk5���$  W�1 @�d  ͭ^ `X 4��'�m @��G � � R_ݗ/#B�Q'<g�	�� ��mHp#�`@)�"�' �xn�	p�s�6 =�]
���, 	�>��	:�j����w����`�$��� �$p�xu_����G'\��}q]�4 S ~��J�� ����>Q'�HX�n��2�� ���|�x��x�� g ����\�Q /û�f�|�Q W��zp�m�� [6C�Hw<7a��L�ї�3�0\`O�~��lò�x�)� U K��Q�qd��'^؁�:��)ג��ث�ӣ���p����h8(j83ַI K 6�HH�x�`��N�zh�� H����q:;�l����ڕvA�cO|�
�����1�'Q��T�A��j���e�n�����b�)���62SIo��� Cj�E�0�#�٭[�^6�k�R���I�Psn�y$ƻ�>g�x�'ß��0d�d:���=F5i38}�[�CJ�2[D��
�kդ�>[�Rހi����6ZV
DQ�Rނ�'���F��%�5�1�&@u�̤���p�f_��)RG΢l�B
��ݡ&�o���u(	�\-F=��ڛ�l�U�%��N�@A �Xa"��@��z�ohx�n�7cN��ݢ�Q<�nJӳ�5�;*4(b���g�Jf�w�b&��j������<|g��l��L�2�@_x+�D��t�TO5I�~ɨ��դT/�}F}�8����F���>���wCҩ	!N㝗�-�������vݾh���oY�L�l����ٲ`���5[,C:`�xS�=��O��q ��o
�M_�������n�G����e��ݑ:a��KoY��X�xɂ��ݩ�[n�*8]���]���q�B���a���$���.^��LJ�ܜ�[��E�����._�t�����.ZY4���l�t���B��b�3[���Ǐf�T������Wq��'_��ʊ�N6>R�H�ݤ3�3[x77��d��CU���c0�������y3�<�a˼+����A��!�f��z�?��r������ǜ�F��擩Z���Y���Fe�*K�WEu��AW� �|�R,ӹu���X��GUe��3��5��N� (5�&1�yH�7�⬅O��K��;��W�"��X�[���&�j��z����\�U3�0����l�g�)ؔ�q8?�}�F_�8�\��R�Z�ru�\��I���N�2�*�C����������S;������z�7֬0ŭ�9�5���#�ҳ"Q6��D�L����y3�3z�Ia��eyBi#�(��*����$3w� H]�"��bӓ�,��b����VЖ�Q ���쀲A�I�������KҙX^S�r���xe��k��yM�9If��:���0M�A�F��W��'C4eflO�1:���[��S(U���g�*M���5��a�|G�R޴�B��4����9���y��w�������:r.�$����I�ܤ ��n-RU��u��h�qh,�qܩ�$q��cm�R���W)��,ʝ��T[���S��%��c�:I��:�)��Pϒ�F����c o8E��Lj�&��[p����B+���YS��(�[7c�u� ��d�gN)�<�h��^��S��x��g��x��+�@�-"�A���YC)�jm�3���Wǡ�V$�AH|�Һ5ҳQ��ȶ��lk�mm�-䷵8�^��vL����Q (M�v>N�a��;�1ךSpq)�9DZ��#2�Ҭ�S����-�IU��e
06"�d�~tF_8����hp+h\�u^��|��CC�B;k����gV�����CV�u�=܍޸��w��,(���i^��)�g�G1��0@�Ki�8�\z�R���B�Ю���]�O.c��/�|��< W�}
�j#k�΅A�������g\�|�s��W^=�̧�8/�u�<!O��*��l��g� �0�pک�t[&`×QL����k4��Wa_MIK�g��|y	C��OY���S8-�V��'�ź�/���z}7�d���Ð�7���vD��;է�v���U��ѽ�O�~Tqڛ*�av��r�H� �a�}`�A�D�W��	z��۠����\�b�W�e<Y"���bՄ�D��Y�d֜��Mc�l��z;vg<��A�KLJ��$�����	����"�h���0r>Mv=���� k%�2e��#eZc6������Py�.t���x澉��b��CE$��������#��.x����Y�ʡɄL��xg:�	�"i2�B���ڥ�(du:]��ڭ;�jR�'O�2��fW��V)���&��Ȁr3�i	4��+��������D�������Og?�~���.P��
	X�TA#BT����wA;#Mi9�r�!Gy5��ͪ�#�r�όs��� P�j���}�0��C�e����E��i�>���N���A�!�9hj�7�C���}���7s����DN[(&�#�.�3D'HjC�n=�����a���" �Ό�ř������3>�R�y�1Mb?Y-�FMZ7!ض���+�-xR�%�t���b&d^�9?�z`٥���Cku���N}���>�z`�l��q��ۿ,v�$�K�V���w��KΞI�z�-ֳ+�k{Wf�zw���w�9}��؃'�IƁ�B��;��z��I���:�rLH�	�S���Qc�"d+a��-����	ө�E;q:!��n���$թ��t���|=���k�����dbf؞�-�'�!��������d�]~#L��(�9�mW�Ht���R
��M�7���HXW#��ࡼ�Du}r�����o����}�g���m�<�<A���)J�;St����M��Y8�S��)�c�����:z�m�G��S����q���1� =f��c�6z��@��j|D7�۫�
7�eT��u�m�<
�
��A �+� o)�~Z"�s�7[�״8��%���w���_����g��i:���:S�����T��3�o�yyo��yMq�#���Wc?y�Su�?p�S?�����(�j���a���b�()�����ɫ!L�H^�O���5H-��X�N�d�]D�O�?�2ÞC��B��m�ȫ�G~=����ʦ�?H�����"=�n���jxd4�,���D+�i��#s	=F;葓J����J��ǔ��p,��M����I�Y��1�D���i�xȅ��%r�$��)����c>�a\�������7��V��N���������p���Ӌ�<X��Us��:Xgi��z�e4�V�Xjﶱ��=uM� �0�L.�V��c����5�)v	�9c,g�;�gP�Xn^���,�Ѧ��h�^���iO��n������V���?9'��bb`M�A�YC�4�밚��|<]uw�����n���u�k ~�5�^��,���ՆX"���E+��K,.gS�J��/ j���.�g4���{��J_���e�>��Q_�1�n�	},��"�'ҿ��M��7:����]�ɳɱ���~�����Qo��d�Ȳ7����|O�C&d�L.R*�4��b7� �8B�g��Ѳ='�df� 2:�A��6U��Ւ&{"�������m�&���*2R�{�ݤ��2%�D��n�ٞ,W��U�*��T��I`dQ��e˫� ���KTM��J�},���x�,A�f��q�C�/�8,�QfY�	XY�Q<J�ȯސN�I��)fos��ڀ�"�Wu��ez@Idq |PM�Q?���#�₥�5��fc�ґ�`���b���~��I���5���ŕj$�gC� +`waBb��w5���#���;���������	;�b��x,_��^qj�quOpd�n�w7W�ivu���2����k^~�%���p���8��d�C�����FAx�6w�_F=����w�X��l�h����&�Ezd,��T���[����30f^�������Ѽ���HM���8Xl���H)�"�,�J�A�d��gv+�^J<:�xc$� -�e�8�?>�[bc���w}�~	���:���s��� ]!`W��<��ìp9k"��g�r����L�ҭϸ������`$���,*�,�P�xG����s�t�)����Q��{&���ٻʴX���Q�i�h����hM�(ߍ��H�3"�Z��c�������V�wa�>?��T$���,�`N�qz!22_(�T�����f���«wl��>\���d�}c�T= ��Y�ˊ?��?,r��&q�_�	X5D�j[޴I7a��l �Z��0<t��LH̑����l���rV�)���w���o�+L�XR�f0�{�*��~�o?Q�nj�⫯���_�;�i�0'�?B���h.���r2��Df�d|�A��nRKh���Ӥ�� "�ɲ	�$�_
ү���k^���|��1�V6��}�t#!XY8���f?�U�L�(����w������9�@"a���@	_O�+mH*�ܗQ�CD�R]L�P]�
9��㦶1 <����Ӡ_�Y��aZȶ8(+�8~ ��X��-�e�0޸���~�UeN��Mq�j��Ōz$δWf��v_ˉ�z��6�b����/{6�v�ٗ�{o	�*�s�H��Α��m��7��T��$Й mz!vJ�Yq����t�K���i�DZ�� ��|͞o������ҫF���6���]��b#`�r�����΀��Ʃ$�7���3��?Ϊ���q����&��<AO���N���ٛqo\���8=�х�I�ȫd���n�{F10�7o��Տ |�&�!�tO栛|��?��#�|9H�ױ��\����|��1��;ێ�Vg��(ߡ=Yd��N2���U�5 ���G�^�|z͉������)�� d��L���0��|�DP�'+"�K��'�ثd���U�l�!�ФC��I�<m"�h`�W����[�~���o����:�q�U`�ޑ��������Kx��Mg�Q)���HT�U'�h0�D�X#;�D\pd$�A�(�>�x�Ш����Cnn��}��C�#{/�~d/����¹��t���SC�esi:q��x��x�3�.k�����!�i�4%�o�� ;�A����Sζ��݀��C��� ��!p롸k��Z�p�ɓ��Hw�C�1�-���e�����p���"z�p�*�<�x�M��P�T�LFן�(�X�F���!�ZK��3��a�M���d����O#�Xɵ��3��q��>u�^�=1�t

<� 6+�dܕ��N4�B�eֽz��~�ڼ� K�����.�|�M��\E�������ۚ��-%�`(�&��A����fm������9n����΃�[v7"�6g�^]Л�?E���q@��7��H���&�mR<P�9��1J=��ӼB��}��Ү���}���:���i��nN�s���2��D�1�虷l49w��V��e#e�q���+�|a�~`8v�������#NɷS۷Ӱ�o�!}��l�b߮��%�R��ʎ׊���jGerm�\��U���.���\��zNsU�":����!]6	HW�_�����)a��*c�xX� N����p�U��:����چ r�6�v�z���M{�FR��t�����~��w��"��zN�EA ����"�i<W4�s�������W7	�#.�kh��=��u�0�e�d����fˑE If�d�� w �� a1�a����8�}�w��l�{��2�g�e�Lx�&��������eXP��-/|0|��r�� �|a��[k�\�}�l��$���?7��6�
�����P��+͖� �2[~�
���l����}1ϛ-} �h|�l9�,���_ @�j�� ��I�#�?����$�̖" �D��8͖���̖;!�`"���qx/���?
}  <f���a #��
`+������@���?�-_ L�l�|���r��%=�lY�g��$�=�l�
� ��9n���9�ZC�w<���` ��lw=�; =���r�a�B�<g��@��u�� { |�D���<�� SN�q���a3[n�7[���1 ܋�Ä��b�_+�}3,�� <�_���yf�wN��^c Aޟc�=���!�x_��g �m� ����Q� � ���o ? ���[�~������x���On�i����c��x�?CA�~���ْ���߃��u��f0�-�=�(��s|A���~��� � m f��P�U��=��C�ӡ��!�t^n�[	������'���X,����}S`;̖���-u������c��Mf�s��s/�3}���>���v�끐��pW�Yze[W�0`�.��k�k��IXc�����yVϥ �u�g� n(���<0
 �3>�z�3���g��� ��~y��8� �8���l;���{���l��	�/��k�ҭx��/ϳ�������g7A�R�ǻγvR��Z�������u�w����і�y&��졳f�W0��y���γ_©���������o������M����k ��(�S�lW<<���k|�E����x�s�E�-�w>�� ��}�9��6�Nx��Sy�s}y��ߑ������rw�ף���c�|��#��^�%�3������'���?���[���[����wA�K����� }�v�~\�i��l��R������B���������Ð��k]���kC��b�^�������/t�7L�q���OxQ�Hy�ɚc3�5<t �T�zΐ�����l���j���Ú���O�HصZ���?jM7y�4�
/3=?���c�}��'Ԍ���uE�t]����]x�s͖�@�_x�?H �3�@�tQq�������g��w�ύS�_���Tۭ��������I<趽&�u�^C���E��pW�初6�>�'���+��T&
���C����7;����5�Qo� �ˮ}�?�䷉x=b��{�W�
�m*��ʷ�����F0�@�
 E1�2-َ���$��+�Y,x��:/ ��g��=�yę��N	,vđ��'��mE�-PW�2T�d;-�:�v%?���4���b�ʫ1�gؕ\��b���wp�mme���%%sJ3�g6�cb�Ax�(�!̛-Z�Gf;�H�7�w�m�.	��e������e�ta`=�����2ڿ,�rۼ���73q+�54�����~��Vｭ��yif)��woTcu'�;pJ�`����z*������Ĝf�׀�uQ9B�v7"P}�N���x�_�"tu����C*��������αX7�W�-�~�Ȯ�]�;��їp*`��F_�xz�[;"&�4a���V�C���t���*x���<Te`���v���Z�밑,��/0t�<�ǩ��x���KMB���}����h(>�����ª����T^�O���%5C�J����
T��m���#Tyu8P���u��\C�|���O ���܈��ߣ8=c3�B5��Հl���J�M{@��Z����5'h��Є�?`����}$�Ж����feq�4�������� �yY=�f����Uº�j:���I�*�Oe���걂Ǭ�R��M�9��A ����#�	'�8A(�6V&A�[!�qWcI�C ���.�(����q�4��v|�©�w�Е�dhE�$��i��F�6H�K#)�>"��'�ɂ���.�);�Q�Ugh���)����q����V�l�h���څ�,˺T���e�W��e�f�wY��鑛�S��<��2�*l�+;��e��X�v�@Q�)p�g���z~�L��@[:�#MC�7v ���Zc�p���e�x��~���e��a:�O2Q�(�Օ�1P�TO�AI��Ǹ�wMgu*R�¾ 2LSo�g.�:�������I$ͥKiG����l��Fv-W�K�H��=X���j���K!�	fA{Q�O)c9�n�ȡ�|Ic�D���u=�P[;��9�!,�o�_�4[ɐ���Ԋ?B����in�(h*� ga.=
٠R,xg�w8�q]��ze��d]x?6'=0V��Dc6��nc6H����ԟ�4m�L�����/�R���SQ��#�Y�lm��p�\��x>�� �4�Hyu96f����R�EH�Ya:�)�@�y00{j�"y`����H�^	\Sݿ>ZOM��<��W1 ?��»�t�(�y5�(e�,P	�PW��y��:��G�A�����(>󽌭�H�.�ךfA��.b�UGz���v;m���R����#?-@U��*��
-���x�] �P����&b�˼�ո�K������i�}�R4L�ά�|��.e+��q!y��T�d=.��3#�}UJ���7�z�A"r9n�}Z���'H>y�.L��1w4.'G�l��Q�����N����Q�F�7������Y�r�H�h��c������U��M~�r3�݀���~��w�Ń�w�@�Z�<i2��^�F�CQUS�Y���[�[�~��P��"�E@?P�P�������Ԩ����S��1�nɿ�){ڱ���إNЩ�/��jy���$v�'���4��<O�QI�^��������~�B�M�\l�}��K̑�BzHh�d�o�+8HQ����z� {D��b٣���cfI�b�#�
��s�����ހH����o�]4�R��Ez�4\����v�V_x�@Џģ�U�[@�Zk����1g%�����O�u0�~[;�Tȫ��"/��DW��*N�Aڈ���Qn�3⨯��ecqZ|ࣖr:��ŉ̇�ȍ�ڵ5 ������b��&�U�A[��ij
�� ��)�n��D�OB4�nq@`��SO�²�ƘF��D�PhZ����A�N}UO���4�)��pxI�����f���e&�:M��5�Q����#EƋH�U1٫�V�Qͫ3e�EU�t5'�rU���'�۪sG��/Dr}��D� �β�{ڂ ��~M�������ؿ?��9�0���"@������J/b�P׀j��:�w�%%_��n��Wܤ)�3�,5� ��XU�:�Թe}�n�	�	"-f~om��4�!'.�ը�!SP��ۥ!u;�ʐ�*����p���0Ny~R�/�"E�:U[��aiS*��=�:|��) ����F1'<�o���y]�Ѻ�ȩ��q��j����w!j��c�x+�?���*)}hcm`9
=�=�|O�Ӱ2��������@�V�؝n������J\5�x��#�97�=�$����$�"eɣ!@�}cK�
��nE��\�6A�I8�
�RT��P��X(�4�����!��{{=���!z��=�zm��C?���R��yL�b�?դ�4���l�V���t�Uk��d�	� j5',��D�<����u@�g�E֓���6eȿ��El繃�����[�a�=A�Gi��&�4��7�/��DK�BI�-��[>�w���\G1|�A�,��$���x&j*2����r84%�&[;�����
�Q�Hc�T~���%%�$wSd�**�P:��P�����r>��!.ɢ�%�X�[υ��hu�W1�
%�ƒ�kI1V?�i⢱K��,���R����P�]��q���������Q+mn��v3`�e[{� ������_�]uH����RT9p~��*u[��n��p `���@�� �g���@^,)��ާ ��0u:Lo"i����߆nv�z�/}�Ry�e��Da��C�����Ra�p��XXI_^>OZ�p��y+�;w�sbެ{����L7jh^��>t��\�Ь�n��>n\zz���^9k�%K�s.X�|�Ҍ�)�r�QU<x�I�Q�_�fG$�v;l@ڥ��?�>
_E�\�W��	D<p]=x��[+�Rv�	��p]L|'���[��\��D_U��J��C�|�u��	�Eb�w����P0�� �3�R��^x!8_���" @m�]�n��g���X�dS૝@H�Y�`�+����o_�c�+��F��<OM��� Lw�D>&���@s�ې� */�L	ܼ�XV4�����-�����z!=5��(GN3��^���Q���]C��j���(�FG��g�F���c�	+��E��ض<�n�@Ah�;9�(9�U�� %]��R�����g>G���,������|�+{R=��}JfRA5�,]&�F�+��(-�cM�^l
�{Z<��"�O���@tvƙ�����zI�K`[İ���[�]��Af��8�&yE�G�x(�@���-`$+	ҡ2g�'y���T��a��-8�埩8x��ʟ�GE`���^�^E.x{}� �`]\p=&u���O�8IA�(ԫ3�P�:T��kQ�ڟ���_�@��pi��ynf�-�1Dr�-�JA��p3�	�u��7���
���<܈T�?D9��ٙ�L<��5� m��B��W���58�bBu��`d?��O�����.9�x�WE�X�.(	�K���{�$�Ԟn&�*����*q��-��|��W�8��_�|��?�lRF}�?�� ��{��_�L��C�����\>���  ��mڅׯ�k��B��jv�fQ�Mt��U���*�o�T��.3C������਋����z�m!00��13�x�p����H��^cvp"�GD&Tb|�5$�"x#_�"�(c ��&d��ч�[�=�Q�U�mSG7Q��)�.��5�]c�u�NF�j�XG�����CuA�y0U�h�J�ƫc^�G/�w@&5�pj�K�ԏ=�"ԓ{{���<�?�S�����7���z 
�v�|?P�H$	|�\B\u� �u	:}u�ٝDk|���~o��bNY�=�*p��нW���c�#�ZF����|��NF���fm��8,�q��.������N�!��w(^���ǿ��h����.�[`������4�ߖ(G���꼍S�P�u#ߡJ�u�ѷ"Ӷ��(I-C�]��.p۷��f]C�A[�n�0�i��ׅ��;^�v�z:^W~��|'�~�:�n>މ�W�����M��7]p?O�ě"��H�5Z�{)q�|��C1�Hbt�ē��c(q�|��Jl�$V"�{k�u?����ԅ�D���o�~��5�{!2]�m�d�7��-��g�%�d;�0[���y�Џg0U�`<eP�_~AuP���Y"�u�_�@��������馨�3!r/3���� ���4a#D�K�F��H#��2XE����{Ak 2�t���.\j�=N�ai�4�?~��VB$� ��]�'�%�I3��gtK�Qnf��� ��FѼW���ks5P	�g�;�|�D�ﺗk�����7^��l��ޟk��u�+��{���D�,_e`qxK�ͫ�aB>�;�����^���Awjw�{1[�r@14�ĝ�4��<҄����i,)���ؙ��\��EI�G$�r<܀�����㘫��_X�:Fւ��'.x�ĥ����'��P�λ��r��B�,�X$���fcm6~��)���Qm�]N2UH�j�|\�W���C?c�hȚ�Yk�?���eq��ñ�أ#�������??^�n��]�U�#&J���z�(�5	�6<���Vb0jWmMZ	C까�%�Z�QDOO��d
�
Q��?p�>.���3�1�K� �ݳ��)<+�h�(x|�t㙆8O�_�K8[��6=H��v�qWq<��4laVv}0�N������E�F�R����H����K�o�T�q�W_ed��YY�8�۠��h��*����P��^���~���5�1����,��n`/rU�zo��1��3�z@ꑵR�n=โ-у�qu7km�2}`�_�|oğ=��t�H���
ʲu��7[����b����/�:_mf�:�~�T4��O��*���i4������r�([�'�܌��ԋ��#jb�r4�����R:^�	n��;�Z�y�PN�n����)p���w�V	�����rI3#o[a
�Mja&ހ?��x�.�A�'�;�I����p}�f�8#'�0���-�#Y.�|�����Q�#�=�(p��/�f����&�A���~�0�r����)�/��<@���r��n����h�}�2�M͝!�M�2a���x����$�m#�-\�{ˢ�.�e~���8dMs���$����ۗI��M���hiW?�=�m_��n�[��-׏9�P���fK�j�L���f�)�1̖� ���2[, s � �8���w��ݼ�COs�~�G�g�5,=}X��QY��s�>>�J'k���+-�/�����K�3mA�Bhw�kHx#C�EQ��G�����}����ߡ�4��>ۏ���Ջ��u��-(��~��h�?�v�$a�/���c���w0�_����#�u�}��'�g�[w�֫�'$G����#�_�K��8 ~��r�=��7&l�
�����ts�wsOs+��| �k�^�˦9��]��.j��L;���(�:= �o��1ǻ����^`?�{.�C��M��u�s��F�^��S�� O���� ����!��Vz�����5���ws������vs��u�K_$^fz��K7<��^��!��F@}���^�-|�_���sxԛ�?���?���n�_��}77^,�[��������W��ָ&���χw���D���s��� ���﷉.�Pl��\gBcW�E�MDb����\j��~7�(�2���֫�Ժ(r���g�6)G�����chGȞ	�
�������poU�-%A��Nn#z��u���Ȫ�C�B=,*�O����Q�,��{ϫ�Ց����a��������u�8�P~����'�z��"M_U��.��x�7��OoD4�` Q b����9\�%ѭ�cg?%uL�.��.�oƾ|��5�Щ2��}g*��l�h޽�v�l���(nsyD��&�Vf���l��A1����0����!ݫ���S�,��,-y�X%�5�zHgk׶4�aaZ�&���(��&�<[��f
� �4��/)��e��y��;�o3�I�ez��F�z�3x�	xH��z����x9����y��Y+���声�/b�=�<����������9��#�����'`�=,��+A��%���k�0�(�[��çP��>�%�Z����N*N{���RW苝|�j�k���~T�TڕJT0;�� R�N�C9�Xx��:m�����U��IW]�b�xX�c�5�X,�L���$[[��w��(}�)vM��4��5[�.ǳZ��A&� ���Y<��*̈́�-���()ERK�>�]�U0�+p����v܁.xMV{U��	�V��xz՜�fJ�B��� 7�� ��l�.ŗk;"����W��{�;�4nd=�l.���
G�ꢱ���X��Ec�#�`�l@%����(v�~���6a�S�l���=(�z�qR��~�r�eh�M��ź@�گuf�#1�X�#_܏*->�k�t躁��O�y�Fx"�l$��t�O�P�0��T��d�4�Z��S�oku(�q*��d��U��0�f����G��5 $��!�B��vU�Ķ0gpe�� ��F_OrMe��ֈ�o��<9Z��hZ֛Ţe"D�m�;͍lb�Oe��F<�8�ܥ7��-||��ؓ��Q��(
���{i��dap<Y��lE{3�,��Q~�P�7��F%�2���%�[Ofޠ�%����6MCl����H�]ʈ��	.��@��0�yx1ůS�:�Ǆ�Z�\��W��Cۃҥ̄�i���;��gX{J3Πr�i���k+L�T�D�Y!Z��!�d��Y�d�`d	9��]��qbgW^Fs˼�Q݇,��f��B
�s�'������k(;�v�l$��Ъ�=��cP��)���%��x���Ɏf}s*�X�la@~���*=ϐPf<��^�xuy:�ӹ���TU�<=.`Y�hU�X�6�HB9ֽ+z�a��{�����M�#�g���8���%Rw�`:5�w0����>��?�񊏡�E�+��o�Od��I��U�X���������3<��,��3��ӬM�k�����#\��2]�i3TŁ�B�����?��lk�'�aO�%�"��\3���C�/��6�?3{��w��t���"��5E�[sG�E4n2�dɶ�w���G[�N	x�u�������^k��7��N�.7�MN�&w�.7]��H�ie��V��Q���y���l�vvpk�a�G�(gO������l;��Gt�x�K�"�mI��k��f芡@��eC�G3֢�	+��v�-�Ϫl�uK���lRؾ�:�d�r��hhJ�5���*SC5<Jt$�ǰ|2�\�i8&�AMW���C�6��h<W�b����n����b�t.���~���e����@��+����'�A�X��L+۬qX?��v�\�ru;��~y�A���^ϥ,7�����.[Me?Q͂'Pu2��}�W��6��D�:*�mO��F?�T=m������F7�dO��Gxz`W��>GGcCU��k'�İ����5D�.*w�{�IO@�h q�>b0�僀U�b{�)�.�E��h[{������<"/;x��|��m��!��\8�8��[���@I��c!% Q�M��!w���J�h���өui����k��65�@	�EL�N@�`���ۦHߠl�R�����S.��&fO�!�J�\����?��=���*{*�T�����qXHj�K��gt�)���rB���*5B���7���%�l��A��۠G��΍�k��I$D���F����ͪZ�K��Wy����yø�ؑs����rN����ٜӔ�Z�݌�J@���c��l����ӕc��b:�H�˺��J#�ִ���y��6K}�:t�(�y�rr���f����@5Fi��e��5��o���@�[2`��|
,*4h�j�R��6<����5hEw�BX����J��c�P#�=''\�R�J�Z�����w鍵���9�QV�ƍW.-_��/��K��K�����5iT_E�����X<�QYjVK<�Q�k)'�bi#����pEz�#��Ņ���@A�tU�4!_�!_�$߶����U��#�l���N��������j�'����N1�z�4~M��2�<��'PHǇ \��X����H��jOa�zʪذw4�z"��Y�*5(���'�N���0�f��n�#����i�=d y�b�m�Q�1�ik�ݏ��� �\s���]e,ڿL<�v�4�,[���(�Ε3�pը4�����ސ�j�I�h5���o(��Zf3yE���e�	s=���+���:P7��+g��'h>���!�<�ڀ
 ��5�OwB��aUo���P|ų�PϪ����q9�����(x��!;�3cq8��)!�[W�&=��E �[����< Cs�1���3X�_���	�U�0�
���Ld�.�%�-��x_������
F�iFTM$��!�e5c9�h�\,VPϻ�� V���Ŗ�:�S�Hwa���M�6�J �x�V�UA?�г��R~����j$�����l oY*�̳?�����@��M���C��t<�rwqG�cȃ��dR�s�2f*��!!�cd��ϋ�5}�Y?�h� 
�#�E��[4���=�0cUc-~xf��\���-8���;�3[�墚��z67���k}w����p%Tg��N��^�%x�?'u�ȹ��bع�7`��='�����RZMÏ�`�ܻ�j(�+(�5#x�[<Ũ�ex6��p�4IDE�8ļ�<q�kL����P�����O�Mģ�>�; �J(9�@�k:`�m����)��k�l1Z��D���CJQ�_a�G�U�%J}�@ox�6�ك��E82,)�c�$5>��W��V����@CV19��) ���������j�(�'���->�́����5��Wo���JF�n� �F{�3��ڐ��RLP������)�#z�<�~��,ޤ��aI�j$��}Ũ�G��B��@k���T�t������
oiBC-5a|�	��(^�ɭw(_�j���ojǋJ���A�&C��%�`cV�v4�X�g�Ԡ��?۠ɸ��+�Z���5?������3砵�P��bH��9j4Z`%{��/�s���������hZi��I�4h��#6�=WC��rI�{3��r�ȗ7mg=OI{X�Y7j�=����Xx�|Z�0���՛�;��o�'V���6���v�a�b9����� �Gϋ��k%E�0y�@�B�P4�¯.�G�w9���h?�7�����*���۬}�'i�m���#��rOeG]d�m�E��|��#t�G�$7t�Z���Z2�n��Z�������(�?V�W{���b@Y�WL!��SA>7�O&��]^>�|��O��-`(٧�����R�ރ7�K��À��@c�s��(yL$��ߖ�ɷN�;_Pi���HWwL��t�OEG�'9V�
�g:�p,���#��<�ɞC�p�����^W3"���ux=u8tC�.�>�N''�2P�f�t��Z3}�d=$]^�X�F\e(��=�xP$�	�j
��O{���Jw8�Nw��P,�ǤK�a(/�^	D��W�ThG�ڡ��C�J����+C�8�Ui�\�.��#@d'"�}dt~�
���D׊;��.W1���1�Mp���UY���V����I&���2KK�۰0�(*�~�4�I�PY��I�V���4��I���B�ƨrp^�i���k��V�q�P�����߯TĖq3�@҉�}SE$}�� �vW\��x@�%]�7�C�*~:�1��V�`nX^���ɪ4H��JC]�����
n���\e��ޝ((��76q�w�+��V�;�MF#N�P<��i	qR����M��T�ltЫ� MU�Ȩ�lb{IA_y����zeeU��s>����kc�w|����W�iO.)�$ѷ8�w�w�_(Ϭ��(_�\ ����N�K�R*T��.�\%u�'��]�+��Jf+17�^��}��J��O<	�m!$a��E�2z�(.�s���p�[��G!���=~�<xˋ��1�����Y�H]�l���a�/$b�	�"���OgϪ������9��O7ш>,B0�k@�6~��-ëҐ��7� O.�r9Q�M����\�_.�5?ё���}er�ȢU��benE'*n!�?A�v<����@��б�M���#Y��T���S����! V��B��E+�Jb��n��ص�ߋ���:<8�d�e�	������N\_�K���ī
�x2������y�q�C��
+hg6�:N/%�D2�@�
`��P޷`|-v�[G'��S��6�]+v����?R(]�*HF����ÍX��v�����:废O��s
$$u>"&�@e�=�]�����A��_�!BP�L$Ý���U��YyV�{�C�b����t_�O�z��L���:	#�\���]H�{ʑ"�ҥ�����O�����H���H:�/�%��?�i����5��3��rO7��QNt!��j�������N9����!���9�=�??�-���RJf��ϱ���-�q��� e]5	���"�"՞~�j��]��oXC�W�y�,vц���8Z*��"�9�ǐ�i�:H����j�//���Li�q]��<ւ��~�O��\��u�C�wb����ph��+;��Z��T=��ҕxT��f'w����:O,���nt�B��Q��c={�Äg��ge��)���"��c���ʘ�tN�M��B���j*va>Ϣ�FD.h����^��(Xī���
2ǥܺ�S�9�lmU���A]6O/��<�9�7+/-E2{'���k|�2�RS%�j0_.�o#�1�0���S��Vt��a5���ho*ɞԃ�,�MjN%�$E�xd�&�i��vN�������h=���f�X~��+�)��1����$�������ze�r��Zv��g�������E|�l���_�^�i�2	n�P	.g���}�U�ۥ��P���l�EJ1�-f])%B �r���y�4sN�I��j�TH�ުdA���k#�Yq��� b����~��)������UV-�E%��(���U�z�ܻ۠Ie�qG^���#c*��"����~�{�2�F��在ĲQ;H�,��Sv�RU4!"�̚�,�#�P���V���@4����O��RQ��� ��Q��c2��}�Y���$o��'��֟4�߯|M_��jnP��t-P��U���5e�H�'�]�W�p^3��.��=�X^��n/�-�<;]b�G�$(�WU���.ͅ ��?�К5�]r`3b3-��e�]o��K�����+Bݥ
��$l�T>�S)y���[X�:5�s��"�gǘ-T�t���np����RE�UU��~GQU��02jV�(e�]�	B	��HnF�j�i7[��JI����	�Fڠ����������+�R�fUD�ut��;5�*�I��y�]�����O��S�����܆$�L�Kt�OG=�ٍ7Q�hO2��gNR�k�5x�e8��WaJ�uT����o��\��)xb�<�*[+c�?(LV�SQa_�����A�C���+j�ݧ��E��3������2OKg^�6.ǈ�tƿ)�����A6-R��J�6x8����Wh	D�P.9��%a�!���Tpw
�P��a"��B/2B�W:�!���M��_�k{���/���v�͍0������Hv\�6��N;P&���j�7��ѧ�f�*�?jm�D�g+ �4�~j�� ��j��1>S,�ZE���X&r� ��ڍ���.�9  ,>;��r�!$*'}(`��F�B���xH6pZ� b���R�}�t�=��xk����Ύ�iUT��B����ץ��S�Z����U�z�~.�w�sXK��U��9���é�M�7
�*�+moL�D*�N����;:������Ǡ��T�KN.c��|ڦ�j>��� *{�c��ﰑ�<l���H9�{�g ]�̗0�M4��g�/��mH[_�?[jk/���W���Cـ1Y�����RCΖ�l���!��������Hj�"�ETN+��<����^ǐ�OIJ�M#h�H��P� �q�G4�O�x�@ yg:�r6� ���xE��b�z���MW���(�pE��i�֚��t�t��Rm�����|ڿ��^�)��S�̐F�<(� �T�~x���f�� J��,9UT��d~���V��zTh,�[�sm�kg^̞��7�{ư�t��X���=ݭ�����T��3�T"�����%�³���]�tI�'���ld;]�C�ނ(�&�dm�<Ux-!.�6�$0�I!4���J:H�������D23���.׫� ��J�5�2^�\/�Z��2�`�z��;�����h���F$�qod�R�Vx��%(ܴ����t��-4�Zz��������EM��]_[�h���F&Ps����|���F�n"��/��a�G�q#f�$�/X tMÏz(.�)��h38����U�\�P�>�[�W�'QcE�A]"��Ÿ[�nŭ~[�CyLK6\�#��1Y%��\W9��P֊�F�R�'0��VB�Pi��dm�!0�j��?����[�y�Oq�;�k����������>�,���ԩ̬FJ���ԭB�0f>���ګ.�A;J�7P�'��l����>W��ZS�I{:i@��i�� y,��3������2�=�.��f��a�޴tN�Y��?'���X{�.�^@��������+�O��f�
{���2oV��a�V&��"oU�/�v;���a!M��}}�[g�
Ag�(n��ވH@�Y�ΊYU��K���`u�UFޭRT��-�2��L�7����X:������x:����ʳDhZ|���@��fN��A���V�Q�<�J��i�����/�*�"j���=��f�h3��P�g|������'����c3�j�J9]��_�РL�J�����^�<;�w ��B;�K�i�Q���_��4T��vh?q�u���'H�>=g|�>�Q�ۿ�nyv;k{��ƪxxwE���5�f�-��P_%S�V`ޝP֕d�X�FOz��D�Bv�c־�I�r8A�P�ߨm�0��0x���鈢u:�!@���T�O���{h���Ѩ<��2E�d� �A�>A)���?7���{�����.����J�l���R����`$���4GA��입�d���4�(%��Y���,��7���0�5��Q^OrŲb2�M��{�sKqX�o֕�P@>�P~;A7�ܴ47�ZLW�N;���Pl���N`��J�+�rx �b�CY��s`�P$n!Q�!�\Z6� Nc�hgr�2�v?��o}:9�>�v?qۓ�V͘0�*m�-S���j�B�o*��"W������5H����\h�3�.��SP���[��v{+tx�|,��w J稞o���8��e/6��L3#fV�j�0]h���5u��@w�6q�Hd�"ԑ����]B�&�"��}��%��c�:H�·�P/�e,8ɂ�2_e�=��ﱕy+���[#<a+$e�����!Y&�h Z�O��ہ��,�{�?�x=������p����1�G�Te��Gj����9��l�\i«HNeG�FY���EN坿��	�AY��5��=]��`���D+-���	X��r4�Yr6֧��c�&~�*M��*uu`<+��Z��K��\(��=�!��u3�8^�;�1� gv��q�h�H亘Wנ�]�e�ȁL�9��ㅏ��{�Uq-��&�d��]p� QWq5��ݐl�@�l�B�WL6l��w!�&�DY/[m�}���i�{����*m-&��P[Q+�B+myu��6j��1�=��ܻw���}������w�=3s����3��ބ����$��ocM��VV�ꢽ���l�㊛ai��Tl�.[K��UM[~A�$:`�\*����'w�1w�,�t������R�]r�K�������R�D�#��H�t�9G�N�$~��%X���it���@�!����#Y�`���d�d��FS�,7���<���]5���������Vd�B��y�h�fe�"vZ���T ��u����t���i����A+���k� �� q�r{{-�f��o�`H�*vw�:�7�]*�s��J���2	�$\ve�����K����3��]���|�{�<ZJ�qţ��w&^�.�?JKF�B��x�iXO,�aM]:�9��]�9��jX��>K]U�SV����^/P�+�͠�����iǝ���=��4�E�6����@����?c��x���M��:n,|�A0䧉!o�:)^���4�����k�-@1	١k_�q�a��_��<���u+�%"�'q���Ļ�t���c:��t[��"��0���t��M�/�x�I���?�
Τ�I 4C���n��H���H=N�p?]2�� HG����ɷ�,w�ě�ỂG�����=n9(���[`��������^���V�Cy[ �ꑵ�������E����L��7�)��ͻ�G�Ϫc��2P�0A���Q�h���)֌V���}��i�⚳e�Q�>�-���z����o��/��n�������?S��׾����i������ԓiQ_S��V!��>��-�P�扯�}�>��]ߡ���Wg���׊�6�-�CyÝ�ބ:@M^F���?̑H��MOr��웭���]�OD|T��jĨ|��O�8y��KG;�}/��x��5�k����e-*���]�;�����G8e�n����#|�Y�np˯G;��o�ڣ^���U�nDG�u�q3v'��u;�ۯ��|��&� ��_�%�1����Dym]��*�yX�?�M�(�� �-��bn��׺_'��L��Z����IYF=������_��G��%}�g��+��A�F�yp���7 �����v�b�(�O�e�F�-��gc>Ay��k��V��:���j�v�����(^"�[S�d5(���6�q��a@��0
S1�.M��W�#�kzn�Q�4����I�eҒeˤ�ȟ��U�?�K"6����1^)�"�rq=1@�8���7��������G0���N�{��%���*O쫮��@��@���Zx��%�]���V�{�@��x �q�׵�)��^~y�:R�М�oB^	ރ��5G����[���%\����xddzY9V]��_'��-n�̐��a ��ף�!���z��瀄v  D����o�C�4|�v�o�﫮���FRY����~�O/���\W���B����!��奾ZG�ͩ�� ���rH��l��F�Uv�!)�*��$��<Z ix�u���i�L�������F���=�A`��|9I��剟{g���S�H���XĲ���2�?H���ʡ�nZ��.`ą�+��J��<:�ާ���w>���-���=��������Pm$}RK<�W��?u�"|��j�V���&㪍/�����c//�e΄��h�JB��NҶ���^(z�#���o� �-��g|@�!Lxн����E�IW ����t>��"tT� 9sg��U�k��
��x1)��_����fA����c�rރ`����]�8r��_��ۉ��ÑF�H����{�l0��q��P�]�`�#GC���Z�!UR�-�ˮ=hG]�W�W���0?f����d�
/��'�\�d�`I ��z���7�xCD)D,�
�Vɕ���G	�*!NUkD��ҕ�1E�!��z�Ϙ҅m�C�\��%��jNU�~(��4����\�LD*�	:��?Y���E;�Cx��㌴)�u��g�"3)��t:�:�&V9� ��E�M{� ^F#yg�:�2=�̎V���he\�0(hkܹx�N�v�Og��=H|Lfa�i�����S�1��:��ťK���5:�*2n�4��x����b�!q������]�w�we��
��
�78�VO�>�G]>n��,�!�|"�=@B�\��؜#�]�$L��o�{�Ä�a�a4�9lh�Y��tQЂ�T^��4��-�TC�)z�3�8�y5fϏS7���{0ҎK�S�tx<��ɋη��CL~�0�K@"���V�^t�qf�D��N�-+h&�rǙ��0�{c��W%���!�1�@N"��f�z� �������}W��$�=`�}0�Ħ��t�����H��,jmu�T[E�'�n0�nHZ��Ic�88@��a�Ɇ�W%���s�2��e�]z����c�������`L=RxRjڅ�Z�+0Ʃm@�BSR�������Z��k�lN�pu�h���881ՏUv�݆lՠ�	 �Bv@Y��/M�h�-i��a�ٜh6�c��,\7(!V(h:�`^��5�aQ�UT���Cx)D���g�����>/sU����=��"��;f�A�9G�K��ܘ~���u�i <�6����%P3ʽ��I^g��c�;%��h{hD>$D!p;�6,u|�g��,��oi�J��"�s���ۚ5��Y��
~&��D�1����?���PM&��6��*�tX����χ�:��`�1K���N?9����=㰨b��\��H�A��ɋ1.��:��i�������/[4e.�I�������С9j�ˇ�H�-TR�j8
�FS�q��$b$c#�h�vy��"�@<��+�N��p�+�V4B���v�;�@b�"��{�a)ߞ�0EzYa�"�h�����^��>J����-.z���0<�oè�F!�DA>�D�g��"���)Br��$0�����z�x���A<N�/!��xIg	�<�fÔ�ޒ?�z}xaj�y'��K���3kk��t�!���t2�+"}�*�!5#�b����e�'��p:n"�ԕ��ꨨ+5�e���/7>2�4��
&1|*F�O'"�pK�:hj2ٔ�����1�.�pb����W�=K2c�[	%��4M�u2�d�]�ui����i��LJ�E�(���.,W+ex`t�?�}A	���xfx5l�L����Z�Ri��ܱ���]Hwѭ�E�-:M�`-YsS��}a-�/hs)ż�)�Fɨ�a����=_���]�M���5n�T��,��¶�D{3A��)��ԼH�0\I��@��V�:`���Vj�� ����(�(����U��#�����ú��W ��T��>�_~ K�h� ��=@�G���_��"O&��놁H5ͪ����∙�g�q�8/��1x`���6���&�{��U�?���[@���%ʬp]��0�R�kݾ(~�o#�(�CQ�|S�R�8kC-�P����L<��g��4(T��0���~�X���S���3��N1K�b�������"�m��'�2�"��i���B4�u�f�e�3�z�)�_8��c���G�q��6Mb�B*���H!�US�8��j�(�5�%��]MS<dڃ���M��Q
A��v\{p.��S������o�4�F��}	�-ң߷/��a����2'���BD1O�\���<v����Pd��Xd����%��b��U�{}�Jg�y��o�碣���Oc�9)�H���j��
�����
<)�1����Ec*j������������@�4�}��OH)=r5�`w�P�s`�n��R����v���z\xH�Le4���~�����:#t/�����)J��D�.O|�NP�R 2y�X� ����1�?n����%B3�A\�S�]�1��!.�n��X�UI�N����_��d�'"6��FD��	���i1�q|�R��~|T�5�,o�d� %2�\`��7�U/Q�N#õ��s|�P�4�l�+�ţPL�n�qQ/��|���S3��|�.�\��5�#�G;���0W��*N,;,��-:�Ңٲ#F��#$�$/(��m��=n_�բM�����1��z{�:�����b�>�:QÌ����~�Y�ly�ɻA�t�������u���q�����R�����f�����s�R6�F)Z� '�V�Y�t��/E+T�+F�k�%#4a���}<\�j��."�ܮDz���2ڪ���U�T(���mJ��r����dG<���q���Թ�\A�����x-5$jxE�����b�S�e�f\ئ�kḚ���d@y<S�}�V�T�Jq��!Pm�m�s���
/UC�Л_���>�`�Ji��w��S	�Q��P����FRم�,��t"a���s<,��z�u�k�NV#;L�Ic��Each"���t��5�Ȋ��ㄣʤ1*K)F�}�٩��IpB+���j*D�Ơa�Q�$6e|7�Ξ��). �EȽ�+Nb�#_�~��"�Fi��E�Q��a����G�#��O鐭Vl1��E��:�I���A;��[ϗ�~�b�i�c]�a�E�=�����]���.匴!���o���+dǣr�{��>sc�Qq���fv�����Ge�E��O(r�B���
����3�E�4RF�O�T=r��yb~7~�>���AHƧ8ު����iC�[��Ŏ���Z����@;j���+z|}P�na"]|�.W��H6U%Dgr���q�k�Zk���Ⱦ����
��}��[�a*����*M�9yݞ���h�kDX�Wߧ�' �&�;:��I�D�E������K�::�΋$�'%)��O�JI���=R�6GS)��Ye���˔lfq����p{,����Fٹ�1:IF��2�k��p�q�Kn|L�����Z#�yC�2k>��݌���e9Ѳ�Ѳ�#���[3W�A�}�+�g�̶##;Y�zt�����(���d���D�h��aŪ14�J��p6�f���L��qx��அiWN+���0Z967��O�D?�3��3V�{���{[Vf�2Z�j�L��!ʨM����ޕ���)0����c}�B��h�G��za�G�U�s)�؎�����;��^_7��se]x2�� �\�l}Zt$�V{r�3胋kzY�(�0�0�l��m��;D}����gR�&MP�5X����h�@݁��g��������5���H����%F!�(�/uſևZH� ^#�k�u�)��D�̩�k�t���Ě�zy�1Zf����c����lia��tc��z�vC�{�e8d�S����9���������
AUh��馞��J��a��,����z�dH��eڥ'�2����|Kxnl��h�!���w�O}&��CU�"8eԅ�W�9��c��Jl�	}T^a��{���)�_R�^��;����@���B"�OЭ;V������(�����Z��ay���S/��6#��ɜ=���fටV(-C	�1��!ie?x�(E��0y{Iݚ��\�#}��\�N����k+��2�ׇ�`.Z��'7H���"^�R.3�E���A3����Ѵ�B{�FH��0�� �6�eFy1�YUCƺ$e����/��K��:Z3����鑞�u�����f�Q+ئ�P�
�q���1)H��J���7z}�rj�T$�m�&J��<���G����0G�qTۅq�7�9�z:h��N������ͷߠ�¿If�]ɔ'�n9���w�Õ�j����$p��G�!�À#M��6�E�.Ԫ��4������>3�w��e����4y���'|��1D>�(��̰�d�%�/g:�\y�Kt���=$Fb�^���fLl3�Ґ����?9�d	0/�o�ݎJ'D�V����F`��뿐;��0�����P]�ǈ''�F{h{�MZ�(7��\����m����Qd�v~���kz��@~�w�E��*1u#�[7�Y��9O�lNL��az�WQz�3q�,M�S�$��!�@�Ux�λ�tTvCx�*��brX���<�^���Fo���I\m�n�9�0�z�[��|*QC����u��J)r������2���Z�Б�>�*��F��Փ�
�����<���g3��^?f4Mn�����ĭ#-�8,�$�ch�.W}�X܁�<vL�����a��G��ʬ��5���g�⧹�����(�K��Jx�L,����<��C9�w���f->5B��u��5g���<Α�1�'h?1�O&2�P��o�{Ε��K��,~;�ڤp�P�eA~��{�4T�5ﷴh����[sS�)�7i��6�_�>������1���A��1=A١��]=��h ��
3�-"�6Qm�'0Od����;�rM�YE�C��T�����S�����(b��_x�ߥ��;���?��%.��l��%�y��b��%Oޚ�Xa�I�ּ��4�8O.��:&&]sz|?�Y��΍��t�v��C��9�>��S@} �4�gr�"�*����H~�)5���%`��yٛo�R��8�$�<��H2H����ABc� ��_�L��Nf�i�8�Gb�ry����E�!S�٢(,ɪ*������+��>}(�0�3=Wiܷ���}�'�2�γ������G��=m!�L.�+\����g.�YW�iP�؝j�ș�X �*�M"翊���}�#N�VC����2QZ��x�(<!�v.ަz�.1���6�=�L�p�j�.�:�ȅ�,�8w7�(����9�W��	�[?O$�����l,\w.�y�F"_'\D^��a�(ĳ�|<}W���h�������-���V]w ���%}���E����f��}G>Δ�Nw���ஂ^�,J(�w�ĳH��7��4�$^u��Uh�+��B���G;�(���zד���<Q���e�/��}��k�:k�:��x�Q*O���/ ͗�	FN�K]n�S�/��o����c;1�f�5�;�9����&�T��DY�p��~1�G�ҿf�Z�M-}Ų��89�z��N����Uò��/v�I�p����i5:�\�(�h�B}��:3L}c��p{ݸM�N�d��t��l3�r� �t��� �ܚVd(ô���P��ّ!��;[�\z
�#Ob��ȓH=S��#N ZE���%���F��Ə
]Q��o;�Bwc-�IO�e���dC���c�������1�a��1ͧ��H����r{S���S�n���T��S"0`3iB�p�}-.[�g�bB0W:�U��T��%<�U2��~C�J��E毛�ڰ �#=���A�2u� z��h���T�h;�#װ�H�)�#22'��ak�g�"#+$�Α�x�1o��A���;G�ek�Α����\�j�9�[�ᗛ���;>�?���0��iNm�i���"�o/W���{�H<C�:�a�:_B�:�h��#\��̴�r�כu��U��{���ADC$�dqyx����c]�!��!;,��(De=A��&cW^�#|]�V#��C�8]g����W�	����'W%�򴢷$'��8�}7�����*�W5�}��Û@P ߗӪ�X֡vT�	�g���	�7�:.��4������U�0��qӳ�����lr��鮏��!p��U������͂cñi4N��up]���44ò3��zNgN�1�R����{��u=�BC��H�ި.�͏#����+9}��k,9\���~�q�&h@k_H�������������c��淍J<��_�c?�-4G����?��w�.	)��6%��`B�O�qPy+Wa5	��;A�m�
[�P��4��MTa�	�:�w����F��OG��@A��vjD�"�!����
;8�\**o��GGhQh�zF�e/b�ǂ?٪R�H��Q"�`�F�L��PC���S�u�N#E����1�K�#�t{�tc��.��l]�	������g;GnSa3�܎[a�f����җb+_�A���8u7������إ�2*�u�hoh���+#	Im|,��GZ�z���8��*�n���L����;���(G[B�W��N��#C�x�;"C��ȍ��>Ey�>7��`��q	�D�f��]�;��U��h�Σxi��:��6�b��d�=w�oG�5�l���Q0��Ӆ�O+���\s8����KN�������(
�Y@���m#�?݂��N���М \U��Kl
 Zr���aO�9��w���9��hB��]�-(�&��	JY�ҹ����^!��O�����G^4���-��(��C�F�R��S8������pZ�k��G�AT�x �9�М�O�1+C|}O�֨��lF�u��*����&pI�{I_&'��!��R�L�;@'`��[�������m�'�����t[��x���4xV�<��l}f.���Td��d#���Ͻ���ν�W���w��u��U���sk\�_<�^t�p�183����`�[4�?ؓ�N�+P�����u*J�u��$;��2/��6`�E�%�����6������b�(��k�`�f���6�yH�4l���}���2p_���^/W�B�i��m��Ur�F=���狃�|_�sܩ>���!_����g0sZȰ7��ě�ut:��^���h���w�hUZ�n?�Q�-����������0�/P���[>�0�~`���:��ӽ�=}YȄ%�;����e��k��_u��������b��cQ��GK�eGKj���B3f�E%5�>��MW�\
�*����[��'�b�ձ��X��tz�+�C"�3Q�Y�D�q"].Y���O#�Zp��--<Q.I|V�:GJ�J�%CJ���ei���$B��*�����V�������/#�,��S�n�+�ޏ��k�HQl�G�,�|��l:n�w��/�����>�Q�����D`��#��ph��7�U�h����.�#fc��a��i0I�}c�t(��X�v]��6���
�c���hǠi�+i�	!W�קH�_�6�L�G�v��v+�n�o�E�r�?V+U�V��_1�R:���8��|ƹ��i�a���uP�j�߈o����i�	�����D%b��PG�H~%��j���T���O9��E�C�<�'HAm�����[t��li����bf��c���#Ӯ�%��l(�F�j�鑨ZD���/���G�XpT9)��Y&a��v)g�߀3��ma��tQ�S�.�b�����Qp��75i4���.�:N�*�s����@s�s��odB�CM��#��O�g�w�n Z�]u4Vf�!��g�X��o�Q	��-$���S�po�ڿ��][q(󫥖͋p<n��b��==)��U����F6�4����7�덆(_�i�KQ�P��>�������V����Od��C%P�^tH2$�mnqmk{�GR����|N����M)���N8؟��#��'��_��Q6����I�F��eQ1���8M��@��33t�xXB����ܵ@��"�� 0��YPaP��= �XțG����)�P���aL/q�����W]4C}u#3����vy�@b�_3"��.��ŝ�t�?�a��\N�3T�����߂��N��ο{���ſ=����� P�P<f��	<A,o�柃yu�:>oĝ��o��RȜ3�3��pn�~%z�-���Y���^�9���+}��q������Uq0+�9��,�NCh�0́.�aѯ��	���9N����E����J�N^.u�Ԗo$Ŋ�c�qN��V^�3�b�$Y_uy.B�G)���o�(͂��^	��G��Bi,_�l����J^�z������	~�Gj���jK���$��WF�m9��i�4�̆�vis&�����NYwlE7^$\re���8��ru���y�sb+�O�|��H�����rA�g�3��Mf�[�&<9t�ߋ��9�� Mኳ'��UI=MY�(�>�\`%��!Vi���0=79W1}T5�Μ�q��ڨ� �T���kd�\��
��ƛ-�tI׹�qtrW��1Yb<�wǮ��tXe�K����
���+s"oMs�	1:L���ds���#�,�{]���&�5�}J�������fܹ����xp�Ҭ�D�r�;-%�¦O�紧��0�}t����W<�h&�Ur1Nf��\�����݋t���I��2BK�L���/o�t:K [��*F��Ņ�dʇ�f���o���q��ћQ?~�V<��/`���H��n�Ky��tƄ�h��d�G�oX'l���k��=�8��N��;oy�=�uU4L+�
pKƆNo�,��iZ$n�&G�f�HM�s�;�6��j�yܨ�_��a�	����FW�s;Ft���&E
�q�]�8���A��!�q4p�ȉ�ІH��h��@X,�y^��B9ù����H��Z�� ؂I�2���w&>�8��<
�3$�h������1�P�=�늕����x�@rL]h�/�8ڌbSO��(�Q	�y�sю�k/��Fe"���J	�(�<a��9�\k�y e������w���3Mt��?�����he�wm����+RZ�^��0W�+$vz��_��7(��G{��w�"�Gi�(���D;�ɽ�	1+L�%ҭ�R�r*�.�T5(�����><��r��Ipn�u�_܈�)֐hw��6rV}=�����T�ֹs�ɨAm�FX�P�렌�~�tO}��J+?�H��V�7k�{1�nT9 ��f��m�S�$s��I(��z�q4���Oа	����G�2�4j�B�<|���� 9�AE�0����^5u�m��3��X�s}�Qy1�eD+�� hH?J�����'$O�"��k���P�'t2���� �	Y�����Пے�B�c��syb`K!���GP,��Z!������a�  )���q�B�w��8
�Z]�	b5��m�����?�׸�'D$@��5���Hz�ĝ��D���/� :a�>����b]��4f��TA*�x�[�U��텏 A|�D�>���G4{$�%6P��c"�#�F͹���60��x�����Q��0�J�\�&�̼��G����bO�nG�'����O%�c������z��r��68��/�Bǰd�[I�u�Y�1��s����aH[��u�d���Z�%,x�w��n�ߜ�>��2v=���lV���6+�NnXoz��l\ŗ@z�F�ՏަGz�]�%,^7Rw�H-�j$�CcN������h�>��b��6������4�n\���fi7~hw&�3*Q�vE�7(���FZZQ�^�EI_��5�\��(#{	�� �/GQ�lzQc�+���X�4�yiz:�,<Y�*���2�q�)n�5k4�);�:��K��:���c��#=�9=0�"30Y�67z��r��FR��Bw���Q���_O(h�p�\��fE���=��(��+��bP��fC�o?/�O2R��Ey��"E�y6 ��ս�r�^~]��"/꣺h�>�cX.������7�N	�k�YD�,�GުG�\V<���/)w.."y��'}�G���#�����E���B����ގW�O�(��7$p	s�e�^~�����7cO�����V�f�-7Da^5$�n�oj���ˡ�ɟ��]�pZ���3'*��'�Ǻ����d�,��丘Bɦ�cNk��VK�����͗.i�%�iZxz�l�t�����gz���o�\��ȧ���Ƣ���-5�����{3:��hu22�!e�o�4��d�5�������e ����=�xE��8i�]��r�>jF=WL�~��Ky'�C�.��2Ӂ��(��0##�T��#~Rz�?����	���/��+;����p�-�>|�z7#��ݬ\��=�I��W�
i�VY�h�� ka�D(ly"z�nZw���}6ˣ�&���)s~��m��ʰ��;�h�6:�\ӎ��bm��Bd��H2�?�s����f=J�j�T�V�e�Dˇ��}߁d�,�|��CQ��\UbLd�1�r�2��h1�ƈ�/ֱb�,�#�q���x�S�<z���P"Pr��l�i�X�d.G(���S�w�xOL_�/%\���ksQVj@�X=�X�ߌ�-ѯᣣ�d�9Q�����̟3�
a{30�kb����ǩ�ߑ�����U "j��M�g`4:xLvdWq4ΆG[x��|/0�3q�?e1&�O���]�%u��PHg�q��pA6��,�d�}�S�Mr�$��	�^R�R+��rbj�.Z��zgS�bҏc�T�1|W�]T񫨚��w�NE�"�I3K�*��Z��z1%��w8h�]�P���X��A��q��ىđ̽xv6ľ�K�}��%h]8Roc��޹�F��̇�ϢG�7B�#%���dl�v���\Vp$?�%�(]&;-x�r����O�T�������G��������o����R1s߄������-���˯rc(�P����R��7b�v�p�veי�٦��I�a��a[g�e9Ee���[������e���C����cj��a���+��:����)��>�{L�ϐ���9��.K�+;�5뢮��@C�	�y~
٘��Pb3֊�>?-����l��Rn6�ڕf$���V�[�@Rb��
���G���	�;Vv�6�� 2]j��0�#���h����<q-��:./�� ��bq;;~'ݶeBZ��}�q������8;� k��f>6��j�T�^�BXx�L�s��/h�����%
�¢�./���!��;���FU��)Mn>�n���ͺ��mch�Ǹ9���42Xt��&��K+^��콣F��������h�c>g���!�X���'�GU����A�>H��b]���b24�K�!Xd��+�g>����*�X�<������f;d|;D?X����>�:�޽}�_ w,�m����1F�YQ�<�qs;H���$�C4k�uC\7�	ʜ2��PD�+��g� �ܙ��%M�M��9�6e�՜厛����嗆��R'�9���r[�I���8���Y,��*��r�P�c�C=�?���n6=W6�s�0�c�b����d�uͽdTc�A>����%v��w�%/p�A�Z�r�Fj����*���p������°Yv��q�ޜWXiޑez�>x�BT�e4}�c�!�Mb�l���w�=�;�1tΞc7u�=��Z`nj�Q���CJ̆��3�I��P�?��4�%���֭�_��&sC&���0D������_%��h3K�[M�O.T�V��q02V�p�R�ٴg����C�,�j?t�Z����D��h�0���k�F��V�43G��[��c��-�����f<Y��B��(�����ME/�Q�ߦ#}<�+zon�+z�}�Y�@�<�-�e�48^��ɕ]�><^��*z/�aٱPݘK%g����8�s�YZ	Y��������B[+�"���H�,�Nu٘��E;�'uq�P����׎8�غ�0����H?b�U�FE��4a~Iٙ:��_rp�Җp��7�lK@4'�W��йz���i�X���'@��V'����F�� �Zk��E�����~������������~K6��d-�Lc�࣑���;����������J���o!�]��g47F��r�Xx�d���P�X@c���s.��H6ڎ����s�݇�-ؓf���@�F��_�~�鷍~}��_?�VЯ�~�w5��Я�~���跔~����~�w>���w.���o.�Z�7�~���-,�
Xi��w��7���-�i���oxUŜÿtޓ�Ɗ����������oYx)�Rę�O�f���[ŷ`�7ffl�H���z�w��:��QԬ	�wk`Ol7�r'&a?X�d:)	;0�Ƭ�q�YV���` {^;��\�<�{e�����5��l��z��Bx�*��Zyo�{�kqim��\���p��Q|KK��2�V�d��\ ����ঁ3����,wB�vB�tN�יj������n:�8	�p��5��n�Bp��]�@ͲOAC����fp9�恻\�jp�����W�����w����÷K���3���$p_�w��]�Ex��{�}�[�-�p���i2���/�1�4p�St�&x6��\�o��.�6p��	�w�>��9s
�pw����j�\������?��yp��;�O�΁K�
���Mpׁ!��{3���s�[�jp��?�;�%pπ{ܣ��~�O�|ㄧ��Kx>����M�ʦr�zxb����"���.���� �i�)m$����3p�Ỏu~W��lp����hO��m�h���i�h��f6N�� �0���r�Y�e��������x�y:�8��2��ݢsz�eA/4\�����,[��+�����P���k�?$��[��w��b��w���^'��ݺ�В�O�I� kI�45xK|u���ʰ_jZ�]��*�=�ݧ���m��@���:��[/5��0v�-%�`��"���޺���V3G��^��/��V�S����Z�[�J�E�&/P��|�4�o.i�@��N���U!�]���Ju!��F
*[�~oY�߻�nƵ]W��������+X���.��eHXE����vV�J�Buw��<[\R���XRZ��(Wq� �.��`�a�
�����к-T��4Z�X'�C�с���b�4�d�R��A(�v@n�<��7{�[��-^,��j�^�����@S1�����8���jo�5���� ѓ�GY���ٝ�򪽼�=��t�H�ji��:�׻9�?���nj
aC�ׅ�L*�V�G��a}�4m�m[t˛�~p^~�-� s+�����h+f�BM9��9�ݒ,s�09�J�����ޖ�$��_*�o*��[�4yyi���/ j�5�j�mЩ>ք�����2isoQ, ��zƒ&i�m�	��V���_1�̭"����"����೫.X���=���٣�4X��Ѱ	�0H�B���YCڶP ����/�N�޺������(.aW2�X+����ܾ�m"A��u ia�Z�,�jh̼��m����1����c���'+Y�7'ó���	By��݁E#\yH�lv����D[�K|M����˽��4v�N�S��vyK�;QX�YM��)�I�g��\uM�g��H�o�x(��h�-���X�e��a��#��V�R�B�մ���ya<ا[����h�1�3\�'O�!x'��2��!�sI�-<�jk�z��JZk�Bл���Y���Ɍ �/o	Iu-ؗkEy����akS��l�7@߲b��`m�?�3!%�֐
��H���Ѡ��;E����o��_�� ��*�;Z�[����
{�ۓ�^����-Hŀ��:YyG3��ĸ���?4a6�A/Z��2�)?|W��ePҺ%P'a�#�j[ޭM�ޒ�@�-XX�PJ�a�h�o�n�%G�glr�%�4]�Kj-u1V��. ����Q��t�Q��Z���M۞��ҶK�������[=��5w�S?m��S�D�딕ÕՐ�m�^�����4u}�� }�1�5{���٫	{���S������2h=���<N��\>nb�l>+d�������࿉5���ٍ��\�� ��1�����p�M�������}�hc�Z���V&��	�������
x�*�)PX7�;b��V�\	\�=�(�ӄ�e�|b-�0��t��a�b`tm#J[�w�E`k�L�5;4;4������Z�$װ_6N�����K$������7o��m3���e_�m+�~�m��s�jt��h��J*��@6ϋU0YyK X%�7��̿���@]P�%��0$���B��QqQ�k�ÃB������44	�b/L@ �p��ǃ�F@���l ��g �/ڸKZ[�o��ʦP=�8�߈�Bs���#Դ���hm���B��Q��'N=�*�f����;�QeQ�%�'���`-�Y`Sk�	{'$��Z����]�r5M�2Q����+�⿃��>���%�JJ�	T��֊��M��F�����(^3F;ec¡��[E[Լ����ڗ�0�2�G���tu��`�{��'���lu��-#�f�R�������
�2Fё�>� nh��Y���S��?�o�ث�A)�e�N'��c�������vڣa�9	�j���:��ă1a9>:���4���t���=:q[:;m�w���ўs�s��K�~xކm��4���:C�솧�^x��9 O��dHg���i�'�e�|-��3
�O}:Ng<��3�O�²��|yc��y�C���iֳ���<����~�8h̫�����}c��ƀ��w��1�ƀ�;<>|h�!����1�yc�ƀ;ǀ���6|��c���?0����1��1�Cc��c�?��E�~mK�1��:��9Djجcq�ߵ5�:�cF����cwh皻u���t��m����4~0�����]��AlP���`孡_ֱ��L$g��1͑��[:���?'t�3��Q��>�c�4�WlױY�����]����t�)My<ѥc?�� �e^��g��r���dz-:f��lO�o��>M�Y�8ip���-I�.G8����ǜD;��}g'�?x���'B��S@�� �ٖ�����̩�M�g��ݝ�����R��ol�\h����"�ϰ���ݗ٘�Cd�M��!�� �$>�$�����ݻwߣ���-���ߤQ~�R�"2��&"�_,Ϥ��hKW�Z4 �4\�6�3����
�f��!f�j� W�M���B��ط�������	(���K����k��>*��@c��mR�I����޶���y�s�>+���hmje�Sb>�c�w}!�h�oA�oH]J<<dj�Կ5�cy�u��	���1�\!Bj����C��6´�{+�l"�Bq=�yTr��r�И"D�]�F���E�%�K���&M���J�?��Xm��4�>�g��#���F�/�*s84�5W��C�����V��p&�#wx��E|lS����?���R�8�j��+h�_����%��Ɍ�2&��/�84�b?��o��S7��"��5���6���r%:%^�&%�����{9V �%+�ƌ��[���y�i^�2��D��3����4rg�1�l��YAZ2������z33�;s%���b5����c6�"��$��_0��Z��´]��J����"����Q[��)��]\i�c�i�)�������_�w��
�Eŵ|�6S����P�~J<_���W��4���Q��o��E��}��N�hC���r?}�<�:���\lD�{p\�������Q���QpC��(����Q�A��y?��䗥)e9
������,ƯtM��t%�~MO�����V���y����%���a�"���g�.,wl�8�����f�]���Ÿ�����%=9�Q��ڜ�!\;�w
��!-�'��Eڸ���t��@�v�km�g�B��<񤵫���]��`��F����=��ݘ�����+æ���R��+hƛmͷ�EG�0��q�O��ѐ���T���6B~7��q|����*��h��Ȥ�*ݞ��Pk�fܼ�0��m�+�*�ַ�KZ�`S
A�iP�?�l�P���w�L/��W:��c�cQ�JV����G�'�
M��eM��귲�H�B�M�w����o�)q)T�oH|+�o�J5ߔ|؛�������%a뾦`*0#����[Z%��5$���DV�OB$FMe�?��o�.O2���QlDrֵ4�i;�O`��ސL@���Ԁ5��vw�5�q�/7S���3�'�T��D��t�	U{�M[�)��=���OҒɺ�T�I�G����zo@J�)�؏G��;�^(�R���g=F2uR���g�E�O��ׅ'� �$q���=���C��;[��*�t��Q
�TW�~�khг��]��Ҁ�5�f�E'�Mi��L���+�[����	젵��6PfI�g��7��[�)�>�&)�$��^�B!��O�y�J�a��I*�D��9%(H�/m
�u�E�ڭ�uҶ��<�M[��j���X�X�5��	�Q��̞i�dW�Z��S#+���sP�	a��U�|9�%M�&��G��mfK]SKS�&m\_�ƅ'�(���q�;���QU`C�ƽ,� ���o��~&�#63�]�[l�؇�YqAB�;n�m����o8�%�ɖ��Ŀʷ��7�h���з 8��ԗ��m@�qp�m[��P�2�&=pjNʘ5������&,�7(�u\�b���AќV��8T��^���w<��d��o,ǰ���Ƅ��d�	���m	�Ca�G8,��D�M����8��V��U���Qґó���d����P*��k�e$�[{>m��ڪ�Z6y5�ms���lm٤���j������$����)���P#M�=�u��5�oX�2z"�3������*>%�_n�o�~<Zݮ���w���k�+�Fp���������Ц���%M��Kl���p$N�8�����v�4�ǥ�[V��mb��\������5�Q>+I�[�{H�W����#DRne����9N�tI<�����x� ?0������WRӘl{�0�`��ծ)��M�<����>�2[nl�݁�zo�|�Ж��f/�l���;��ko5�Q��/��A׮��oZ�h��m�ٝ����ز�G���a)￿��Lʱ*�}"ir?(��)k�p����f^;�[Mp{�&'	�i�'���?C�Y�Vo�AL@�c��^�͂�e���>�jm���_�
�ʺp��cd�h��7�[Y��������}[<�)L�]V�s��)1m�J�ֆ����4���1<�c�xL����o41�d
�Ȁ]�T��ȀE�����+��-�`�Y%�������Rp�s�8"�j�Z����sy
��#��M-^k�l�_�=�Y�'H���BZ��[�V�^k��~��ڢ���������6F�>�P��d��Ri�rom�X�6��Sp[��Ad�ρ��B��@��Lt��Eȿ��)�����`�5QXC��>�q����zrrVd1�
�Z�O�	�$�	Aӄ�\�tYEk�fk��L��lk����k�dm�n�H�1˓͈u��sq�����!7R
���M�M���W�5���[.�_l~�~!d��45^4�D�i�'*��J|Y����)+���5oK�&Ռ\��f+�Ef�Ș�Q�S���3?%�:5&�E�:	�� rN��Km8�AS�*�����4�Qd{72�4C�ˣz�(xu��	+Ux��p�6I��s)���ם�H3���Z��q'�ͯ0�԰��8G��D�A��t=y�8�
S:���5�WPp�c�^��[eZ/�=���`4CЅ�7h�匭��.�
m�^�Va���_{Śjl�*�֭��Nc
/�)n�1׷���OM�#c@`�D,$��-��]ΈmTg+Ԏ�^>b���O��yֵ��8N�>��5��/iԅD���6�[x�m�͖VAD���2�������G �C�x�3�J7��3��}��6�dh��m�2���m"V��S6S�],�V^&<�ͣ������ �p�f��:��^�i/-�-�߁|66�R!�&��J�З��j�m��HI
3��ы/B����YW�&#+�y0�ab����N��<j6��W����L{�%46aՋ�O�[�B��Q�*�#�y�D:�e�g�=��I� J����x
gqd3��Ĉ��6
濐�hߡ*1�;�)@��� ��͌<�˞YI�X��jl4��WnX�p��+�kH.2��apZ�+ҩ�0j�0�AV�Dg8��\Mt֧��'r1�`b�aXǼ�C���D�k����X��!�jzJ{�R��Ўc4/�`Aa����|���p�2�x��w�v�����1�<�Y
���
�צ����XM���ˊ����XX����q��y��XqAAD7�r�X>\��p�n0���#sh.�����\�Y�6А�2`l�5?%������`70C'��Y:<��i,�F;�H��M�O`:]B&d�����c�e�碴o�<�K���Оb��5x�ǣG�B�}�3��{ʦs��v�A���/��NgŬ�M.�ʷA|C�Θ���_?�¦�asY)�R��°ʞ��¦�a�(�t
[x9��
�g:yj�z5�\
���� ��s�[DX�6Ck����6�
[$®U�f�a�S�L
��v�
�0,��˲��/��
k��Ǡ�,�������r��`�x��\H�Q4�4P���-���}aXl��t'�a�����^��pT��E���t�j�
Jw��MMw��E�N��󰝤��E�U���t'�ak(�$
{�9G��A�<,�:�I�B�ӛH�x�F�E�m������x�A+�~g�~p#���x�B)�����'�7����oe�������a(���㨰���N��]���1?�����%}�y�I|9]�����^�,j�~��Bq.���\�%㴱�j�*ϩT�!|�8愑S����Q=���ã�]�L�k�q�x_Ħ��Q[ʦr�a���g�7U�a������/����3]s_(�%e���<t��H.RBr(x7�K��3��CspK���x�E8c�b�Ǯ���p�ǆ��9��q<��3k<�Ƴ�S\N���Q]R>�F�$��t��)p����E\���g�̷���8+�$�Q�����׸�����)>Ìz^VN(W�>���t�-��"=h�IW�Wt�ӕ;]��ͻO�Ӟ���y =9�*4�ԍb^,��,�h(}��O�� ��(��^ͨ��h�HW��G�÷�Q��5�OK��5SZ�)� �gF�������[�&�z~?����_)���'�ʦʟe��dS�\Zm��Qg��Դ�4���s�>�C�u8%�*DZ���ǀ�g[+��M]���e�44\9�5�C�7���R���=W<������S���=� @��Kx�<�Ҟ�X7�ل�����\�u�����2S�\�\�c�F����J����'�E��Gx�<w�\�޵�7.Ʀ=�|��:���ż�k�Q�%����!��;�m�/�Z�8pF�(��� I��%d�r���8���(�?�-���p�y���fR�½�.E��^�Kmw8vV�w�_P�8^�5rFY��ԶP�0��Y4x��V 8֠�[Ax�m�
���n^᥶�j��^��U^j[�<p,���!�Զ�
��1�F�g�O��
�}�<�_�ų\���c<����Ż�����r���x���|��7���_k���)o��cz�l��3��-<p̩�[Hx�S�
 �i�
oJ
^��Seji}Cx�����,���"<K
^1��cg4xń75o	��c��xKoZ
^	��c�5x%�7=��������S���=��sތ�~x��)^�]����b�MH�-%��)xN��r5xN��I�+<p�T�WNx���-<pl�o�]��Wx�X����H��<p�Q^%�YS� 8��o�]����ul8��?��J����1�1��)�]�����c�4x�^n
�0��c5<��9��$�!�}"�I�L����o��pp�°O7�-��.7\���]�
p���_	n����C�C<{�sr���y�3Q�eEQ��Q��D�;����Q�e Q�e Q&eLQveQQ6��1c(�r�(7�g�(c��(/���(o�2�(��e�����!���=�N~?�֤C�(s��{��\<��n���Fq��i�^c�g�����s�U�[�;R�i��w��g���ݿ�������
>��C{y������:U��v�z����3`tfcc�/�&���5~�I㧔��W�OI'������ӗ��ާ
��������}K��?�{��_�!m��_�1?-�4~J:�)��ɢ����"h=�LPGY�*�F�Τ8��ӣ����Xn��v�l7��l�����iƧ��G-s���`��V�V���{^e�����mD�
�`U��6�7=��epm�����T� *���y�.�EbtGS+���
��Q��:V8[�6T����)������fW\#�g*�M��S�H�����v)�ƪ'�����!�Ct{l�H��r���/;^�F-�Yi�^�摮�y����B�7f��XN�!~�K��N�mWCؕ�\-�����6Q��)��r����م0+�wp7B��f҈SH��/,O�e2ENI��ʸ�������,4F�@��W'n�m"?ϳ��66+����<�(�� �m"�naצP�?��۽ʄ�Rl`a�c�����'ܣA��[����|6I�/�=B��etc�K�^���/��y4߭�Zu@�B����H[?L���
,�{0��4�����އ�ό�跛���o��N�bv��?�]	XUe�>�"�b`R�np�� 
���J�%��d��i
�9DIjE��T��ԯEef�JeFFEj�9d�d�w���̿����Ͻ?�q��{}�[߻�z�>g�O��߱���;��5B��jO5j�n��'�<�Z���r9�[��/t��9���
���nG�0�s�sa��.t��}���[y)^|�i/�eǂ�&!U�?35�DkO��Z��h�C�h8�y�pc{X{�B�`�Cul�u�*â[��S03U�nXd�mu�մ���8�˿��^Z.���:�zf�ٟ��K�~bf�c������JefYw�,o������Q��R���u���F�6�R��a~���ɒ4Y�v���u��u�r]g�=���q�n�9����싴��瘟�W���z����������Uz��<-�u�"ǚ���L�֝�c��"C���ls��T��@�Ǝ,2:^��؅�Q�s;\g�cz����1sD�$*	�F{���'qx7���A�R�pk�ûѰ�D�>��7��tLX4�����ԍ��Z���؞=�N�$gjxS��k9Ȥ!PE�h-��4�[#pV�F�7�i:gi���ѽ��m�Z`�a��Ҭ��^��}+n=>�/�o�u�1r����#F��a�(���#�+�&�n��i�B��ޡ�M�1i���{~d��hǹt�3:�g����xعK��'���@s,ͳ��W���l8�[Գ�;���M�qq���U�h�����h���욡�n�m���j�U�j��$Y;�����iL0_[�Tk�����Q�r-��E�-�ͽb
5	6-���,����kk�s��k��7��ݝ��j��֪�"�*fhn���ҭ�t�c��˫�N�&K���"@owR��@���'[��>v������[D�L��"G;�w����f�k��#�X�6;Co;j�إ�ې��wyd2�����ކHk�C�3l�0P�Z�)�|"�el~bɬj�ʹƀ�1�����S�9���-q6�.�آ�*)G��::��R��#G�7yv�Dä�UЉ3u�kd�#����3;[О;�"C��ءkW��,�ȁ�ZVk���T�znL���k�s��6���=���Y]����滎E�p�۳cW��l��R�����������W�����o���n�}Y����;�{�uש�X[QUG�^m������0��VJ_��N]���ԫ�{�|�}�r RN֬0η�W�ӹڽK��:��c�Y֐N���H�9�u�s6n��б��ь\{���R�4�E/���p�����Fzf��������-����B��{tZK�/����v����Y:��*>�j�'S�ތN2¬2�үcƵ�� M��z<]��Ng���Ιr4nl�`��W�E�N��������Z�"-�\�ehc;��8��9���S���̴vf4ZWU�=hc��d���գ��V��wd8|��o�ȅ�^���F�Ni�5�����1cW�n�,5�oލ�����4�hz�G-y��o��+,k3����"s`�b�b.�=�u��=o�ue�n�+3Z�v�?�K��UB�%Zt�j�q���?���G�hە?Z<�hfqav��<`��}��
�V!�
�1OGt���1j~��M�cC�E^��g�ٞ�U��0b���ܷ�.��b���Y���B��4�ÿ�V?��e�/ii�Z�rP?����5���W;�n��fF���z�����eL���:�Z�-#�7��yV݊�u����L�=]�={�n5�A�ǎ���ʿ��Z��u�}��~��.�v��cd�>���7X��4ˬc�;Ϝ9r��0�s,gEU�Õz6��Lk��t�ε�>[E�j�W��s�Z���)9rx�yv��V�$�=d��u$�t��+[��b�8uT7cXЛ���Le�"��6֧ן���,8G�ȽV��bL}�3��u���wf���>�iߠI�˧��2�K�Sqb�<�˻��o鯝Ͽ���׶Qe���2��M����+پj�^�
�o��:�U-�W9V?l��^-EY1j4׭�����f��Ǵ�����+�*4�����.���ʷ��ܖ������1���8�w��oD!�=�����AC�*Ek�q���e�ؕc�!FmS7��c�_�W����h 护Xӓ�׶���7�ʴ���U����;���J�f��,k��F�2��q|�]�`�d��Vi�f�gu[��y��C~o������V:�#L��{0�����u2D�"��&�Ok�jb��x�x��K4�?���D;�N�%��P�%erO����_�^�/�O�I��H��"�(*���|h?ڟ�:���i��'����A:�Χ���z�c� �}��@�F#LC13���le��P�d#��F� ���Ď��q�\"w?7�[­���6p۸�\3�=w�;������e>�O���_���O�?��NB��^xA�$lv	{�S��8B/&��b��+>*�,^�H/IG�f�;��,��9]�%��]�^�`e���~�E}�t	���Q�E`��C�N�]�l?v;�}����a���1��������8����x>�4��
���_�È("��BL'2�YD!1�(%���u�&���I�K|@�'�ǈo�S�9�2�;a {�O�����>�ه���E%QY�<jUA�H�S�%��[�ڇ	e���;���L�žξ��f��ٞ�tn6W��q���?Ο�O�����I�^�WJ��һR�t@:&�H�J��&��%�B�I�#y���
���V刢?8����������`�S��߉�$.�c���T�A<����G�2�l�"�߉�����?&g�K�5�O�&}ɻ�����$MJdy �X ���pjX!�*����~��j��R�T�J���P�K���j��+�A{ӎ(Ei�fi�CG�Qt�5�N�S�t�6�.�M`�t)����Wҕt���,o�k����t���O7�Mt3�B�ҧ�3�y��Dm`\ƛ�a�&�A�@&�	fP�dXFd�0L��3IL2���`2�l&�)`LL	��)e3�J���b�ê�0aekam�zX�f/��id���L3�´2��3�y�s�ic���z�ެ����,��A,
�Ʋ";��`��x6�MfS�l�����-a���b���d���l5[~���ew�ul=������L5�G�f�<�{���^a��v��ypޜ���s�rA\0�r$�r"7��ࢸ.�KⒹ��.���
8Wr��
n%W�Uq�j@�Fn+W�� ��s��n/��k䚸�Z�V�g���%�
�Ƶsޕ��yޏ��>��y�'y��G�Q1��$>�O�g��|_���~_�/�+��|%_ů��~#����w�u|=��o�����F�	<��o�[�S��<��·��Ap<o�G��� � !X@R`Q#DQB�/$	�B�0C����@0	%��TX,T+�J�_�B��Q�*�
;�za�� ����G�f�Eh��vF8/\ڄv� �����#���b����b�,�")��(�#�(1^L��q��!f��I,���b�B\)V�U�z�Z�7�[�Zq�X'֋��q��_l�ģb��"��g��A��mb�h�\%�[��$)@B�@)H
�P��XI��HR�#�KIR��"͐2�l�@2I%��TZ,UH+�J�JZ/UK5�Fi�T+��zi7D���~�Qj��B�n�Z�S��tI�"�I�Av�=do�G���eD���`�I����r�#��Ir��"ϐ3�l9G.�M�J��r��R�����r�\#o��ʵ��N��w��^y��(7��r��*������Kr��.W�C�V|?�_	P��AJ0�DRa!*�Q"�(%F�W��d%E��d(�J�bRJ�J��X�PV*�J��^�Vj ��*;�:�^iP�*��F�I9�4+-J�rJ9��W.)W�6�]ѿl�=N����7���(��A(��(�F�1h<��&�)�4�Fs��]�����
�e�h��FkЍ�V��;�:�ݍ6�{��h#ڄE������<z	�����s�<0o����� �� ,C1c1�1
���$,K�f`X6��`&�[��b��
l%V�Ua�j�ۈm�j�XV������S�&�(֌�`���<v	���a�]]q����!�6�{��x#ބ���v�@��7�C��D ��DL�I��H�!" ���D�L�3 g9Da"J����}[�A�d0d�4���A�����I9_���h�������=�G�av>D�>|?~p�>�7B9ųB��/�!���+����G!��(����?8��>,]�z�!��B��^��|C��W)Ô0%Z����&~S��ԽQ������+~�}�a�]k���d)�,�y��Hzs����!l_������B���%@$���P��Oa�8\�0q�$��.��A�# �bd	<*��@.��ɫ�5�7��W��e���(%_y�ܠT�QN*�f)�ڳ P��=����bC#3�U��0v�v��?�o�?�O�=��D"��ð��*�u�k�,�G�?�*��Rk�j�u���j=����D_����Lc�@v��9�0�߲�"���=C�]����#lQ�V1�	�U����~W}��뇝�3���0z��~�&�y
r�;�����ǐ�.q������qq��S,�2�\`�o+�)��U\�X���:{[�}Ն9���#�r|��:��!�?��Ï�߁���/◁�^��ĝ	w ~D`=���_�]��[ʗA7z�^CW��hfp�?�Tv� Nᢁ���� ������x�A���J��6PQ���6Z��L��\H�������� m#s�0��m�b�s�������Z�E������k�^N/8����q��	�U���x�S�<S���S	�YHT}^�]���M��fB��b���`������/��D}o���5�=�0Tw`�d �UH����ɛd 5�ʠ��j+�.0��`��?��?�N�=��n�0�O������l0;�|�x�7�ø4��\o�`/?�_�/�_�ῄ*�E�'H0�x�~�u^���pQ���1D�9�(�*~ ~y����8D%)R�4�[?�~�zdL<�a��y�S�3��Z��9�?�I��L��U�5e���rSћ�d8����H�6	��#�-N�=��XFc��X:D�ǰ]�l�=�v����M��B�ax�6��V�ܝ`����k�����P��}�2r-y�18��M-���X��G�7�w��M��E��{�eC�&��V��>�(v,0�r��kl?n4'pqPI��6q�p��cPG���M��O�W�O�2�<�%��z�}�c�p��I�g�W��n��8@�
9��8q"��I-����5�s��^� ����O��W$-�8�,��ZMu��u���]2eTU��|��w+��Rvާ��ڸ	b����Pt<��w�;��ؓ������E�a��^��?n�=!�
�	�l!T�k�W��<B�K���]d�-T���0��S���Z���s�'�^�|�����r�p��/��������P��P�d2yL�+�A�>���N�ZaT���u��*۟{ ��vD��u�B����h���- �����"U�(�l�8�iy00����F��z��71�z|�L�M|��5��P���r��\C>C~L6���30Ooj&T�ǡ�s���<G�B-w�����x:�U�F�8w�8Z�\�(ބlGHE�#��&�C�W�dF�$*ӔY�le>�5��ruM��I���*F�ax>���ş���kq��!'����WP��,�u'JO�s���Q��^PFAX5�/{;��1`יPs���b��]{qwA����pk�mܛG��h>�~�
������ *CDIL��9���%�l|�<-	�$`�J���H��� y�<B�/O����K��&�?�����x���W��PB
"v������,D���P/t�U LE�C�Y��� x���5�k޸/�����x*T�K�Րw����<`[/[��������},�DN'ׁ��C\
~^~~rM�'5�N�,�(�*pW�?��'�o{�����&v;{�����Fq�PWN��2�X�B@��� �B�	��k��ޅܿ2��W��
�gȮW��Ȋ��X6pf��R3[�~���V`����Vbx �B<��@���j���=o�i��M�'r��Ƽ�B3�f������:;�r�;�{�\��Z/��5�~.h��Mg''�7���qvs3�3�=G�;�:�3�N�5��	�w���\�5�KK��'N�$���	Y��Z��>Ƒ���ӊߋ�M	��M��5�}�ܹ��p��]^���g���C}�ܪ��$Ny�eU��4+{����2�����)���D��<$�pN�	1�������|{[NF���C�`t�~`��Jcn&�hJ�-P/'f�5�g"	��&�Dq��Q�qHLt������������Ȉ`$(}� �@���1(��(�*:^rN`���({���Nn��U`���ee�/B�K��CB��ps�׮���Ol�s�Sb�G��|���l�=���0�C��V��|òa�M�)z����~7�%_�=����7B��&��]����_6��-�߭z�nℳ�!�Nyf��ꜥƯ{�n3�e{ϐ/��wN�p����K���ϖ�1��mWj絻�?-��mT��+}3�����iϦ軥�ʮ��v}6�Yi��^�t�Z�6��ץn[��s�_��kwN<�c�s>9�zR�,�{ׂꑏ�������g�~��6Vz�j�~��ǯgx�����C�v�g�������1.y���**�]���ĵ�pt�.x�հ�ԫۙ�--���d��h�@_�h��^�	-{��W�*,S!�=�Bݫ�*�W���}���(��;t�fœ㾊��uW����i�oO�����Cy�����_�o�5i���pR\Ӯ��^M����vi�ɵu��D����b��)/t$�E�ʢ�ɛ������%ջ�?6���Go������sg���C�;��_0*m��d��C�}br�=���Sj�Φ<F]}�ַ֞Y�従E��z>�������:��c�aS�O�n�鳩㎲S�9��G�
!���ϝx����s����}�O��E��ߟ���w}�߅ow��V0.$x!Z�s3��S������3/km�c;��v�#�������;�S��z�+D����#������,L7�� ��Y����L$~NZ��(;��	� ɢ$F����K��8����;M�W�F�I��šs��"�04=?wtafA~�є_8otx|�:F~aA��>!3+4X�uhLR��e�QQ�CEgM0`t��ZT�HbۗȪ���\�`.�y�=���}�''b�h_������Ԣlp=S~���M�#!3#7?/����������,ǽ�9F��ܩ�
'�r''C]���n���\��n�����=��á���q��h�ԍ�;�׶gI�C�s���~Z�[u�q��#�g��oo�5l�3'�v��k���u�����'��S����x��2[��!g��k������#i��}:�����k��Y���,�Ͽؓ��Vv��ȗ��?���c�'�[_�hD��+k.���k?~[�+��]Z�[�~}2�w��c���ܡ�f�^֛��󚹠mټ�Y��L�~�pp�����L�}>9u�Ħ7��V�ܿ$7��ץ��/��}���}���=��Ψ�R������V��U���\�Jх�>�מ�,�F�����<�W����G*ws���V5qur����CUh#xw�8�(5�j�)���((�>-w����T/-w
o�Q:<�d*(�G����P�R_V�R��mϔYhR�R7:1j��-�H�8!+�03/=3Xߡ�T��1���`*4��r�y�I{X��)X�\�f�\�_���Bҵ�d���	MFx��E�	X(l�Y�y�4��T���DU�Ȑ\��E#�X�����BO8�rb�5Fp�#`S!C��̈́7&��Ҥ�VS������G�$�991�+�Wh��mR�$�q��8	��A�3�u_�¹�f#�	Iaѱ�S��b��#�����艑HXl�]���i8�S=;6:v<�$EE"�#��q�kt�&.z\txXR$/��Ób�G'����$ũ�xN�L�N�kw~t\,��	ׁ����I��:Dtb�d	��� �xZ�L�� ��m�929>!21��
�39B�b{����/-��K@�E'Ū����Ð�0�1|rLX?9!>.12XdjtL��96R3RL�vAx\lb�ɠ|tXL0\�=�|�E�8�U61l|db(���S����H8+&,�m��ncg���3�ݜ�����TX�[�$�f�H��Y�k�ֶ*B��S�T�����H�m���TuC*��m��*Ϲz��3̛�E��z�L������s�g��4f�e���q-ۂ����^3�F9-m�t���o�{@Tqs�zg@���Hh��Lgt
��N�x�Yq�[��9�H��і��1�1���"9&��������N�H7��u�h�9���=�Ҽ��M)+�}���S�s���/��Ȼ�ݣ�ݑ�8}D�$a��7���%ǟxͫ�����c�������s��kQ1����}��FD��'>{�œUN�4|�����]��� }>^!����?/e�BOof����ʇb�"�`����_�]��E~M�>�.��z�`���8���v�A�]�;\}����=9;�Fā?����ko�۝��j�R���&v���!���43�r-�GC�ܴ�"c�#�q-w2x+� D>�4���|�1+.oU~���}jl=��}ob^+�����l:u���+L��įى���o�A��\�#x�����#�?o��|���k]h�]��/>�����P�����ʯ��m�vˆ�)��oպ�_;{(���b�O;�b1��u�G����~<|����^��<_��:Q�<>�{������?�[����A{�;=?���{��K�AK�ܛ�o������!sn���������+[�b��9�2uȇ��
.�>6ְ���c��"�l(wj��h[%w��i���
����ʶ��#��G���e�k� �q��hE	���b$3��kS�?�W\�V9n��FGP��V�|nP���6��߾e�S�k����|��^��gG��}w��ל^�_�����[�p��h?"N�sb����\w9�O��#�WoM)~����;^7�T���K��.�3M���u�G����O]��v*̋��mc�A�~^g0��J��MZ�       ��  �       @                                   �   � �	�!�L�!This program cannot be run in DOS mode.
$       [��O:��O:��O:��O:��U:��O:��K:��-%��M:���&��N:����^:�͈<��N:�Ͱ��N:��RichO:��                        PE  L ��9        � !  `      �  �+  �   0                       @                               04 �  h3 �    0 h                  :                                                                                    UPX0     �                        �  �UPX1     `   �   ^                 @  �.rsrc       0     b              @  �                                                                                                                                                                                                                                                                                                                                                                                                   3.00 UPX!	ta�>-���� �[   �  & �_����T$UWVS��4��Ut�]p9�� w������B����$0�El;�s���\$(�uۻ�oMd�t$$�|$�	f�\}{��3���3f�4$)$���n��+�w3ɉL$,e8 h7�}�/l$�D$L�-�߾��|]M OX�N��0������R98t%�
�F;���w��[�R0u��bxf;,u�
��/�	s>*��lv���r{HR�!mc�I7�RT�Lr$7(�!9���!�d���r$��u�2ɑLF���$Gz� _�L�At}Hz�2!1s!r�l?��e���Y�(of���� ��y��l�	�ŀ�\�\��dK�\�S����2 ���=Ȁ	R
�t�Ƀ�&�c���9��R��A9y���0v��x��J��$o*��8:6��|���V3Wt-
�t�e �Qf�O��E��� 6�/K�v������?�c��W�����3CuF=u
F7v����F+e;(w��ϷuL��ԉ��B�Ows"��N�Z+6�Y�3/-+���H7]ha�w�������4[^_]�
GVMat32 optimised as��ombly code writDn 1996���-98 bGilles VoantB�ۭ�S�X��5m�P�
3�tQۍt�Ye ����
� �[ø����N��$�8�<�Bp��o�;�
�Zt|%ځ���K��؉&�-�7�)�|��r0���վ�jd�|q����؃���5(C$-���Ös\4�,�>��[\8�Iz�$�[���#�O;���j��?���߈Լ�D1��u݋��m7�;�ω5��y���������8x��w��023:u�D23D:����u��u��q�� ����	��,��4*M+�=w�"�;}L�{j͆�^��x���n׉Jh!}-��۹n �,�K�,�a�Y0Z�oY��$m68��6 h m,h�#�)from B.;0�� Ra3er,<8Oo��l� VEWߒρ�?�������_!^� S�o~хہ�U���A�����r�+������_����w�������3Ҋc9y�D+�V����C����C9���C9����9��������vM8g���t���޶FHu������w��.ǿ�5����hb�1][��_������ ,(�ò�H�<�D+DV�����
T�j�Dh�yklW�JQR(��A:�8  <@�oou
�u@�jPl{�n�����t�RQ ����.��t��^[#8��a�b3P�"��nVw���^�PC��k�eL�,��"l�]	<����?VW�}��3����h��+ʺ���(���@
r�M5��[��¾����3�5�~��Nu8P�B��ؐ|�1�}�_�n�^e�vhdl����洼��S����89�������3ۊ�w���3ˊ����������3�F^����r����%�ef�l:����6肹*4O�m�ٻ_��ˣ�z�&Ju�.���0��@j��� j���0SUÞV�X�;�W'�.��� &��:ͳ|������
;�u_^]���[� y��~G �W=C�G ����
|(9W$d$���̎����4�ݏ�7 ;�}�L�ۆ$M���|�	�p����|��m���;�|�B�'(i�[��|�&�w��kh�Bj2�h�R�W 8�M�����w�nh����^(���r|�>j�K�NH$�E��6��U�F,���D���~FL��� ����VLO(Qb�ж�V:F0�(>Qm{��ND8�WQ�<V��J�I�K����P/}�ޘ,��0%����m;YR0�L8�fiE<>�����Wz�F+P�Hȉ��|op?�,���	Lw����FN|���G�X��W�GXN���Vkn�>r��� X�,�m�
П��ƛă{*�@09�+�GP�n��A0s	;�Yr\�[�C$� ;�/��v'+���{4�/�Fk���r�������sK�kdT��C@���/03ɊN�u��L#�5g�M&{@�kL�L�j;CA4��f[�R�<#�!fG,�#��uw8f�K6<	HB;�v���d����ĿH;�Vtc�p��t\9H tW�e��$t�H�@,�7���VN���}�o�	��҃�G�Rm�A**�����f [lV\��%�X�qy6�TU�Wz�l�myz�
���]j�8�����a����	���l���|{��v�|V�X�I��>��"��;�t�JTÏ���t_R9_|t9Y�-47�!��W�Q��x-���١洗���Ot��\<p�NM��DK O��~lvΥs=����ܶ����˅C�lK��q�;������aF=7u	5�P�lNK���#�B���}�q�Uhq�������ux(A|������y�H��vś��x3��dd��}��� ���rq�o�����Q�<&�ٿ3�)�S0��R����%>P"�C����, S%loF���u7Z �����n|�ul��t�@�v�K�������%�2S�lm1��X���2
���*��|�?@�����>b���Z�(��*W����ui;��~���\���:I�\\t��f�?&��f����J�h~�L ���S����#���7�!�<���7���P�`�-0�k0��]��-NYH7�F�=���=u2|IJ��Hf ��?�]��!pxx����`�>�PB�_��)�5�uA^.�/VI7�.]%v1�X�v�-m��Fx�}k��*��q�-�.=�|��l��+�qf+�[*`�@Z�VJ��^�OD�W���m/��
�x�*tq|�1n��PvM�p40�F�lk�VE_A<�R�2rF@8NQ��u5V�0>7Q�sM�m�<����H_$��_�{����0�`��m��<}���%�!�:E�uU���@�������ݻ/��]2K�+�Uv�('�UN��M�m;��CSD8W���w���<2&D����|ݶ�� �8
�I���<� H�p	n�T�� ��s�����r8�ɲ�D<<ٲ\J�ֿmzs+��_5���o3�/����N񉃜ǋ+7o
@;��	�t
�=7��(Y�U6�R"�V3�v�[	�D��B4
��^�<WwtH��<Q;�ض	����"X��`|W��|�~6���Jx���@�����A;q���.�rd-߶eTlrpX�r`@g$iٷ \[_зx���O���;õk{,��gl�w �c��E\�����˫Nd�l�-́�Td�t;��K8�r?+ЉH%Vl|�Zm���M+�,_�(=X_BQ�\gm$T���\!�^�M!$+�+���;�c��NF7ȭY��LRP�h��ZR�L��:g�M8k�'Z�;��Rc`D��ّ�1/�PX0�F��^��.��]��$�=�<BCb	^��$�C�S�Klt?�njuN��ՙ�G��ȺB���1���)�rq�9�-�/�hsk�VPCT+�+͉D�ޢ�%i+�T�q���k���;�r�Nudk�A����h\��#Ջ2`�Ka��VM���.��Q��P�?r���	�r$���<=�vE��O����.���s��B$pʍ��݌��h ��}]ܸ�E�;� ٽ�@�V+ÉE�E~�V�hU0SQR������iu���%�-)E˟c�ek
�^��{Q��:J0��=�'�`60���,�����}6�A%@�P~0��TwY~L�Ny�U/]S�D{<&,8#��b�
aV2Fhʧ�P1t'�m2�wp�B�u�-�W� �Hl�V#s�L��/ۯ��ˮ���LF+FhHw3����WDU!�`K��'އ*5�J�"�
5n�}Ҋ�˫�f����= \��5�
s����\��Z�m@�l�5���7����6��dH5h���б�x_���o~+�;w2�9YH3��{���~@BF̳U�N>r \�HCN�,7�F�P�NVF�~nJfMu�IkX�j5�g�0k�Px��X���v;�JN�n��F|@����D�	��Z��[Վ��Lp�tU����E��:��,�f�#I;���aI�����=���D��	����r���ȅ���ztq�>k)�΋��rwź�_��]Y��-�t��^]�&�J�'�Q��40��5�$��9ɓ&'�5^��\L
0�\l	���5X��v�hmVp+\�X#�ˎAFx;�sOM�H�>9�Lw!j1�ju^�;�-E�hݑvYo�Ȓup�94�|���N~cl�Np��,�l���4�i\'�H ��щ�S���L2���=Ѫl���P*����È
�5������\Y
�(;�*����bHQu���YAy`Hd��pb��V��06
��n�Q���ZP�t��A�Br�p`�W���IzD���Bi��B���B���u2�J�K�BI�h�;��h�� N�C~8AH��3]V�t@@Җ5�,'�Q��d��Ҏ
���Ru�@�Q1��@���`���L<��_#ź,��:�*[+��x�, �d :FA=�w���uXU�`Scm��^�_�����4n�u��%����.� ��AGA���n, ܏n�Ь�~$xt��T_nk(=��m=��j<�vЮ�n:��;����C4� ������{T)�	�L��r�lQn��n�v�,B��:>fy�f9D*��o�~utABA¶KUP_f;1�B.�"2m�^�rn:	�K����+ӻ��~�n��~h��}/�
Si$VG��̓��@P�9�СH�L7D��A��吠����U�+z"L����oX2k��d`l��_h�����[����h؃pH��;x��@jdL���8;����l,V �u $(,˲,D HC-˲@8<	ւ�P�ш���9��PX���QP�։UT��^�S� �("+����l���(�E\ �r8�V�uHM\�<w�<am���uw0|<9�V�0K2����'��h7=g��<h�p��B��C���-ڨp�h��Q�Yt�>`uM��EOUP��n{Q���@�m{s�����H������T"',tm��nX�/-D 2�ׂWT.KM���Yl��E.�Mw���  �t}�l�C�P����Q�����@E@?��}\�=�
l�z�طP�UQ{8�wk�� q`
fV���ܯ�%sU@R"̶ꖨ^+�'_$t`U�#_�A��4}	3}�g�fV�g4��\��a�!�}��)�_��tP�~�9�/u��GNFH�@5�-ŷ�G��=t*B3K8/S=��w1��Sp�S�%b P��JK|.&��h}x���C��#r�uEl�1����v�-l�'��������A�)FOu���^�t2:���� ��n�O�-��v[@�ˋ��u�6t�kH�u�
�l#��t��_$-ZP���o�D��V[�J7CoGmAӂ3M�����V���7����y�
?k7E���p����F��DP�kQ���(�����j<>�B t�ѢֺGD�찢�s�@�?b��D��u��:P�	P���m6��
������
<rK��v�H�1Y�d�=�8q�����ׅ)D[H��M�TV�_�QV	P�z��\����rNR�h2E8����F��������#H��шj��M~]��}���9Xz��N�G��ME<�C�r EMEv�,?�UE�G���>U�bM,�oۛ8umD,L+�܆�R�(U�H��W.�LS	Y��hP/�6U^�.*��O����F��}L���pJVU-F��.���<
�h˭{\�r)�o�,�-��Vv; �j �RdѾ2��~U�?=��F��� ��U"q�XWv���E&P_)(����C�M+��˄�͆��=�;��_ͩ��h�	.K�_%�a�\�+���
���1��<�,aM�'�
5(R�2�&Ē�6�>�7ė��t@u��~8O ����FVS���+-y
��[�������x�fB�9�~x�W��g�.���j;�$u��R�߅\S[C�X���L0�
�WU0�FLC0!`/ݸ:�m�c���Z�`W_WPo��C�-eh����I_���;�Q8P�#Sc*����`/��ۄXSM0R�#�3�99�u,
������n�3_D8@�S��g8�,,=��B�~�<�H�#��A��A��j�ྐ�����>��y^��m+�$��#�HPWŉ;�u�%�HE�w���H����R��}�~�+�=a8�
�	�r�e�z��?8��g�p�_a�v8Gg4��Ʒ�L����s3.�!({�&��Y��fwf�p��q+^Ќ�H5"�Vo���ɇ~D�)���Vq�;���P1�0<����ݺ,�#��k��=�ך�[{~m����X-U76��WR������H�c�n��|ko�GT�F���u�Vt�o.<"Hh;naԈ=�#�i�L����HsM�r'�~F��S\Br�68��fc�]�U�d;ۥ8<���)�\YF`vD,�N��c!�!�`>u�3���\!�zϫL0�G���n,�x��@<"�I,ki'�=r�)V
fa��s���I�b_�Ru	�@,j���o�L��}cf;/���/fVV�lH��ơP�S�!�W(T]��Ku�MɢC.f���G�[���x� ��8(���p����V�W���k7��B@t.A�Sd���8%����+(>���5��{T�
��b���
Pn?^\�%xSPN�� �:)x��.<@!H,lPP[OcUK�M�%�͘@�paa#Q艋]�]��u��
Z���$���>u�WG�+8��(��F4�k���QJu�g t�
�e�`G06�� ��j�.�I��Th��P �
�!6@$�O�f%ڐ0(�t��@S�(t�ۚ(�$+Q�V���3s ����
Dۄ8���v�0�@Y#��0"�V�8F8|�P戛��C�k�K4��e0�V;�W�K�Ds2H�,� >�����.�n��0��>�cx.s<����H�>k��L:ы�����%7���G1pr��Zn��7���2���n�w�c? ���.�*u7�+�?n���2^5H$R�H�e)P4Q<��U4�Z�\y���S?DRLP�?3|
6�(����/Y,fƞUn^xC��s�7�� s,3�;���粭܉`qO�|��?�@'arԋ֋��Ґ�+]8���8�;���v;��Kl*n6P�rE��5,�*�_��W��|,D;�u�Vo�%�s(;Ʈb;ZX�5�s�HT�]X�ʵ5uqXj�K�S�4Ǯz#<�s0&ak3W\8�3I�p�К^�<S��ڍIu"d��;�l�n�N.�� ,���!�Q#`&ev0��vi" ս�DgH�2���Qmh��%Do�L�L�n���������b�C,B.Dpw,�s6A���_%?�N��i�t��ҥ6G�@�?��ǿ�%����Ё���v6w���l;Hm����}A�ӌ��:�_o|��F�C�C�xM��h���A��
��%�;�snT8M���!ONѾ�JlXs��˾�Ead�,?�E���z�(
ڭW~�g�a�V���pmr�0do�ܸDs!<4s����1\5�7 p�vr�$V�K"CN��n�QP� lR\��]��X��A�,4�WQa�-3����5�;��þV;�s;��J�L�o���
�?�fx*�A6(r��|t�=��\�[�ҊT���6~@vo��5�4s�+����Ѱ���{@88* �w��/�H�����?Z�$���;�sC��[��"�s�>r�!�|]�޷��#��j��Z�B��tB�-�
���+�x���o�P�4|�I��L�^�����?ޭk��@K��w>u�l�횊Y�
\����u]l�f�"VQT@�;���	,0��h�?[8�AR�<	���D	Q(�X|3��=�VZ#.,*^�dr�j8r�A�s%Q�O�B�焅#ZX���{_k,>ma��V)�ʵ��L8 ��e��?�)���s���T 9W��IG���Q�Y2����%��|�) oێ�H�s�ϋ�h�ʋ�j�Z��L.@L �n�8��n{GQ0�>�B&��6�F�Ej�P;ơ��L���������o��NC�]�H�j�+��+9l�NKLɰlp{1�i$Q +5���7U�!k��:C�2jZ�w�A��KF@a��HHQ�yFD�}�#MK S;0�!��\�ƄQ��R��Z�a8@��9�j��/�wO8���Wp� MKR�c�#Tm�%��,�5Սe������
����V%���S�PӰ�iHK@\��g��� P�LS�vMr��N+��p��2D��V�����TH� j��&��=X��ɾ63�@Z�e0�m_]LV�s`S�-�!1��uGVH+�����VqĽV5@j'LJ�f�ǳ�0�|N�ep����KsYS�t7�dI���o q�.i�>+Ջn4�+�58f�G��C.�ǐ�v~�j�WxK^!�;|�
��~u0�0\ƻˬ;������HC��2t3j˥�4�5�6�8�k.��=�>W'�Z\��'U:� [1�<W �G�0[2Z$uWI(�]$��HP�@=���@���(H(_���<40[%0P�O���+�9j|��\5,P����"�5��Pp@����H"��Y!*��W��F� ��ol�LPA��^6W9����V����N�����N,�N���s���Gp��%^�\��3U'm�U

�2$�,<�F�^��1OH����/��l�ֶ�h��W��KQRt{����h�lG�����ʜ@<ү0����,�
�,tR�t�H�{M�]&�c@-H#*<H��uh���7�?6�#=(8}y��a�E��HS�R6�W$:,,�s��E7rȐ�j@���#�:���6A�mVq����=k��+�>"ж�V��T��抙���}z?�|-��RI6��#@u:{o���PH�K�l�%% ќ]�G憟��l�����9d9at�+ُ>��Y �<��-Ur 9A�[^�2����\�Xo���Xdx(9G�J��+A�B�:�9%�)�سz��?m��Kٖ:�,��#D0�
,�)?4���=�H�>D�lq�uc��,V��h�
�_�
�2q|�p���nZ�4��X8���p�MB,�	�J�\��AʻIZBst��^uX�I���x&`�8����� �ةx��
�����
�G0����L5;,�8G��+��!��j:/���LkM�4��o�DNͶ�m?TR}MW	���L/VOH����9,QW:n|��v;��AMXF�HU�Nʯ�6kL�2hfB����P��_ٟ_�L������ j�7OAr��o��涋�@CA�Bz�ri.C'�D�FX }��a�I<���x� a"�$���YPq�Q�ԙ~<;މ\>�/�AmkW�s	+�N��	�,��Y�N�:Jv�E-,/s	:�xl��D�/qi����S�Er����T0#����΍4���׀����U`h7Hu9R*�ݎ,
�^6�8���etǃ��4� 1���#�H�� #S��4�1#̔����zfX�'iuO��}מ,�zx���Er�<\�L'v#�����s�+�Z�໎����+�?���;�r��+��A�F�Y�Zsk��a7�-\��۪.�S�v,-�7�[5v+߉+�AFOu��=7I=u�M��v� Ҋ��f���FG��? ����r,3r��
r'�� X�����B;�c��g=���K!*�ۊK΍|��Ǎ��Z�I�Jpm�M<�۬/O}N4y{�Etl tRq�J�S-V��.���X�H1WX��]]��t��-V����P��R���P��B�Em�1�QmS-�
��+���:T-�3��,���=D
b��Y�?�{ fT�T�#�J�;�LD;�l�w�f���_��8
��;�hg��@%~�h:�F~(9~5��4F�j��m�'7>�6*"Vhq�ωz}�����������|YTl�>h�J0Q�u BP��"w��`1| ��k*AOV9z��Xv\nI_۲�V��	��ʪ ���	��jRQ�2����&/A����vA�> �wU�j�:����ô��K����1��|C��Q8#�F�eI>	��YA��R�2�#�5��B�s�*�d'U��/}����j�I�qk�P�(�~v$6�!(�Mnq�>ݽ����UF@v�wN����%
�]D��U���1��K�!�V�����g_�hr�%����&�h���2?`�h�W��u�U��M�,��u�Ũ�"zF�zmɠS���ִ9g>DT؝K��9�
���c���Jܶ�\���h�I4	`C�K�;�HBu��:��H���7��H9
!�H.���te52;,s�15H02�"���P��!/���[�duǜk�&�grjLf�_�Pcx��n�B9H��[BK7�
P�9[�>VB�Lr�)a��(�!n$�_ �0^�+	O��;f���e,�l��@����|	�Gc �.݆��M��O�.M�\P*i��Nu\��k�Q�QG ��+?W��ޠ��G�^�8uY��
l�VUA�;G0tK��t�WhU-`A���;�r�X���B�`Z�\��Ss1O9�{+뭤� ϙ�9ɭ � 8t^�]x!��n��u���
W�-��a�B� 3s"�:Ԉֿ�tu@��+�ŭ�mq�<+Ћ�u�x!*�c�~ʵ�V�N�76����UXe3�
���E,h �#��e��8���^'%�D�c]z8QS� /j�	A̷���$7	Q`�O��TdU��
��SQ]Ryy�W{��S���(����R[�W�R]҄�mG��ƴ_L�YS��t�W`����b0)��p[ā�B:*�x��G	�֦i���TX\`��i�dhlptx�sPo|��$�����䈌���7G��T�DEJ�����u�9tau}(��{B7E%9�:��ě=���&�l�[��:��+�98I6��A�v�z�.ص�s�?��d@+�v9>uJy)�[�;�u�;�I,v�J����+��s�wo��\�T+3x%S��r���m�z��\�L��M@�yX�����,�7�%&�LXI�l�z*�X�m���:t#�m܌�u8������rs�!��X}WC;�r�{���6A����jLCl�;O�+�8��R�"(� _�ލ@<���ƍ����ُa5x� T��J�t���'�X8PL+�#:"w�`�P)aC����B+���aSK�i!�H;�d�PB��˃�6�+7��h���6l{�~A]}���}#+�r틬��'@�8�E ��6����7�G���$0U(�ǋ�؟�ҍ���D��^�{t>��@�@�M�%�
C��+1x)����X�ߣ0+���+��Vt��碇a�\(�׆�����L(���*ӈ?��k�,6�m�,0�ؕyxI�u�w�����4Ҁ⠀�`0� v{��t $V��]h� D4!!

��cRWh [��ȵ;�nkP!8�q���_�0�)�,��q�<�_ r�B���t������u�:Gh�I���u���?bOM#��t �Ju%*�+�*�+�C�u�� ,�,��H�$�i��:�^ @<���(B�"}ҕ�mY�$�M������=�
��<��r��C`@��=,pW,�C(W�h:PԨ�2���%�:z>��<0�4��W4Rp�+��Pm�$��hK`\UR�j0�.ͅӖ�Lv����L(H8�~�(r0L�Q�V�{`/��RQKu$'�:���*��jw[�P�gp�&� K�5�Q�C�0���C�u�Y#�t"C�|#�E/#fS�v�R(�B�$���*#��:�XY��G���
\%���]?6���`�e�`ÿ�Yԋk4W�#��F��t�nQ�bvBn+�(�6q�]�Mib�% �o V+�ThK�՟�	C�[��<U�Є#�5b���@4����P��>K,�v���
u~A����(�Fs4!W؅��+$G�WɁ,'GWV ܡrѡ����Z;{�䌊��`�x(����Q�5EW��^���o>>ԍ�o����)>w�t
(ǀN6�	Ә��$���=�	0�f,�2� �}�ܬ�d�s���O�V�nb{�����C0�Iu�慵��t
��>����g�Ծ�Ȩs�O2fU3�Z�O8܀؞�~b7Ub�ßWf	��￰��p���1�x�ۮ�F��7+�����CA�	f�j+�_f�X�����^[��x��A�a`Y�RĄ��⁎v\��jX���. �a�]���{�G��A���N}�����-A۠@���@{[�D��RF��|�����f��YV��y����fJ�޸N wx;ȡ�~^��c7w�瑾3~��<�'9�~^�G�~r��;��3NύT9k��臎���f'ʍtu�Em����+�<���	 D���$2):lH ǆ&����y <�z�;W�B�|�~{6U�.t��t���qaL��Q�q�gO��#���pv�
5
�����P+prw��MQ|���;�wqW�b���WUS�u���O/.��,1�"ȍ|�(�G~Z��]�ϓ�V�VB�q�.�=����_��[��&B�^�Q�,�ݩ\�ܝpl���7Wڋn���E�^��9�DnC����)Y�.��}Þm!���}�ᷴP�P� AP}^h|��k=#5��[�9B)2Q�u�h��ˏ<(�8`#��9��p�3�l/�l���m�ɲ�L=I~^k.n��fM4���ZA����T��6�Ƅ0P�jBh�W�M@��|�5P����}]��E�����A@6�F�E�VJM֮�F2BL��,֢ǆh�X��|��]��oDc�������|SW��5�c�K}�؋h��s�1
���X����؄�~�HV�@�����L(�LJ��s�X��1�o���������f��!��X���⊌.J�:��B�E x f<:^�w������"7$L�������V{3�M⚥�vhG��*H�=��s�J��#R��ݬ9�8dl��4jr��VPWff��A��ot.�N�m)���j(m�6����ۻœ�}ڴ�y"���0�;�ru�^9�(�wA����3,��/u8���(v+���}��ቴ�1��~��ŋ���u���=*���]�J*��$(�#8��[��mW h���*D3m�Weع�G�፺@A�[�%'���(���N[���F��Q����̈́��]w��0�+��F4�0�څhV9	f�=u�~��|�@;�~U�G�O�|R;�`�[ 08[B��Lu���|)�+��<��O|k@Rǁ������V�z����lh�c�X)�5ʙM'N��<��,sH��=x��Si�����#���V+���m�&�H9�ڬ-����6�V��jE�6 ����H��Q�=�E�C+�)tb6���ϒM�N��0���?u8�o3;���+��έp�����׵���VH[Z[�ɩVsOW0:��}u��..m� �V���t$+�W��<~[�`
����NcA�u�ѯ7�a|6,�x�N��mTLQ�J�Dm�BP-�uh5��[۴у ï��� ����g�,�ě��	�(��[J����.��ȱ�v!uHt����}��@G=�J.8Q�n)n[S�V�H��Ћ�ú]�ޅS�뺊��۲��f&��Q�.1�CUf=� >��h�M&�-}+��n;�}
f����̱#�'t�O��[����
	� <v�
�k/۲��W!,�
�� ���cH�o] �-�W�P,��,���p˓Ѡ�d�ŉa��9-f��E�X����@�b\�a_@�~_<B����H���?�l�E���)i(�~9ùB��� �����16�vlZۗ�-�ȋ��(��\#i��J�y��f���ǭ��]E#��!�tH�j쎎h�tJ�$�!42��9�*6@mX�%�!c�a�n����0��E���G�۶����LBK���;�w�};�`��vI;ֆ�D�b�<��۴�������R~g���z��C�`YH�x����9�G�x8��f����~	�T7�	P��E���d�!�`�	�J͂8F��Y�p6C�����	�^� ½^���]f\�*f+[��`A�~^��.��Y��>"_@������]����]��
,�2���2�@�r�L��!��'�H�	~�#@�[��B3��Zh�`z��;�%L���jɀ��m�4��O�jr	�����f�U��߃���`3SK��[4Ws�pX�[Cb�Q�J�*KZ�A*M=r��W���4�%�����mJ��t�B��/$�P�Pr�,XP���i1���e;��:�B�s�\TY���f2����)⊚����v����f{'��;�~qأXtP�������X��CԞk��^�@�馘�B���T��ʬ;�{�$pn���L��k�4MYĮ꣐� �-b6��Ի��1���܍ˉ�ڱ����%3� .�S�O�BtP<
ߟt_*W��������xE�q���:lx���z���j�T�b�,�0*D���;i�g"�Y�,�Y��҄t���H����$�Y���X����N�d��XʉL2MAw\��8��O����LCb+E�� �����_9Q_��l�΍��E*z,�bEztҰ�g�]����Iu�U�̳<�y���(�'�G �]}� ��4��D+�A1��H��;׈XF�_���C^>ߠ��TV
��(�������J�������B@�d9�V�pRД �m T�{l��54DC'B�&uH1t���Ɉa:OV߭�V�&~?K�QK���~5��$[Dp2A^+hI!_< ^%��u"C1�tGVG�IU����nV���A��e��E����G�ձ�����H�o��H�N�7h{��:5C@Iu��4u�[� ����q pH�y)�}+�j8�>(p�Q&#ϓ��48MT��5R,��G�{]��f8�(~#3R��A�(�� �F�D?�P��O���:�u!��t�P%6�
7��#-�n^��� ��V�?�LA��UuxSM��������
�BF��a|z���<<
��R��t�^:�8Dt�|
����eÏw]��`�����)�En< Wt@�W��,"v���$$��J4�l��Z� e&6�/�{,����jQW�7It�~��z�B���BR���Uu> (%r�ି ����Q�����){�t�<@R`RP_<7��;�r W�@8M(T)�h�e�� S��<3�h��U�[`�I�8��C�S��2Ā�L��'��WCz\l��ٗu$
Q(^����.`�0������ ��OVjR��hT��g-T$:�
iƣ�?F^�OB�&�i#�Lk~��(V��ы�4�@&���W�P��@/����j�K#p��1`�	��O��V�́�4�� L&�ls�h�L8��Y�
��86S�;�#����@�����;�w+P�ߩ���+��E��L ��]�+|��ďuX�Q��G�B�B�E�6~.ۼ���<0Pu�|0Kuu�]�@q!����;��E%
;��hA�"�sD��[���&G�m���54����B�a@/�T�N\>�3����P�9A.$o���'�P��Rf
!}FE$�$���Xdk_�Wvw�����G�Oo=���������(+�ْF�P��|9>[wK��|�K�U����7���QU\ ��D ҹ���FHd9;�\<,�'�J(�,��6$0�4�] 8<D�r@D���#;�0U)�6�b��$x,tl:	|+��>Z�8s�-.m�v.vvbPVQ��X@K+�ru�@g:��_j����:�Br�S�
S�l_؍�t�Rv�����F7<g*Vv&l��N荤{�QrR-8[�ݕ��~ě����Bto@���6����s�8%�ɝ��D����@0Ȍv%9�o3��W�%������!pv�BP���tɲ �=.��#53�V����]���r	����V
6��BL`smC��+%�j����N?�r&�lO$�{�*p�Nx"JAaV�ɹh �#�AԮ��W��^7�f^"I��N@�
Z���;HuL.
�x�9G�2��P �V�����%��+��x�E��UP��ں�4�I�`&�,�\B2�:V]$��%;R ��(�@��[whXQ,|�W�6��SRw��!��L��	��Ow�Z�je �`���@��!�u���9��9_Dd�+|,WE z���P�^������4�jl���$P;�R��c�"�����Zv�+ÿ��K�^LuGK-X�8?:tWl�m�4<�;�7TPe�)����@[��`Dh�&���Ixj�P$(�&-,����h5@�O@8XD�h6�GxU^��.��V�w|~�oV!�Ń��S��5wGN0�1~NB�t�AR(�
A$��N&�����9�]�� ��!�i@N>U [W���4,�B�H��ac�5]Hb KL�[��IP<L��D��`�J3@�@HD�d��7&��.GH�M^BFh��V���[x�!M�:RB���<M?�\/o0EW�.Y��uf쑹O�p|��>)�-�|�ez�I���2pa��8\vRS���BÆ�
9���h�va�`�A�!Q�	��'�!�$JDm`���R�;�)��kW����<R���}<�\QiX$ndګp����&Z�L�gs����@r�%SšT��ʹ֪�Un�FV����+Y��n�M�߿lp)�p��v�G83�c����~����PqEB�=�.^\ZT^n�:7+LΉt� ��.7���hV��/y�$$�yS�JI�v�@|Y��+�/P\���� ��_\%cF�6I�-���~H�����!ퟠv5�K��w`U���{��ah��S���8`U�!����Dgc{�X,$�]�w���	����s��Tͣ��HBN@�C4��Q�臙�x@%�G| ��7+�YO�($$,��m;��v�!�Wߠ��J	�7E�v!�iR��SW�����vY�v�>"�t@���5t�|0Wh�h/��#B���P�{q,�:����^��ٯ>��h�-	g��Q^�o�Vb��htX���F�MR�_�,�OW�G�m��I_	�E=j� z�w�0_(74h���[�~��O� ΐ�}[�Pt�,!��耣:k0?�����!v8���3C�m��I;b�=��d@�r��E��l�zu��]�\Ol1�	�\_��L��
_��׀z�Qض�lVh`<HLw=Dx��d�E0�38.Pi�9�4]T�A-�Lܩ�c�ϙV�jRps��"zFV`�{v`�
23����D3Qm:�)�df��k-+�%�/��6�VSW1/w��-׀H" !�X�"wk��\u\6ǰ� $Rjc&!�o�pm� �E�$��� "��P�*X��*p,��Mid6��T.@c���`s�s�(�`ډpp.dϚ۵o4N�09� ��e�9陡�!g���b�U��y��ڳl;��G�`�� ѹ�C �.�P�q��.�q������v5U�	�N�hu}CU}4!�uiuSu�$54�?V;\inġC^}SR��Pk8@3kQ�g�d � �Vd� A�q4BKo��$u?�`�䤢�2f8Uٶ�@��!04�کh8D���v�oH�G� Õ�V���~��L�w�����|�� ��"IRe�?�z��X�b�0C�UdJ 
8�����v#�&{�=�Pv�B@���B3ri�޽�Ƌ2��r��{1���	�^���[)��^�+aM�D���U�n�ՀJ`�f�b'd�%��E�Zo�����Q�~d�W(
K���I�!���~���%0��Uф���$m�SY&X��v *��*C��136*j
�A"�R��� +ȵ����К�~�+����V$a���qL����C�]�<���;�.vT^u�:��U�WT�L�-��1˟o^``��QS���F���nw�"��+��ʨ]��t�	u}D}�a*�v;�#�б��QOPR�s�>#SQ�J����H�hp�]��$gi�"�<Va��$���M��/k���KTR��w��,�AR�%.�E�~�`Qj�CU�U���`��Dth<��e*t�ej���QCF�lyUWP����pon@_�
m^�1��+VFTJ�W�je�D�Q_�Q	s4�-p�vu+�\���.t���k@��N�h��U����7�����ރ-��L�U�U��Ym���ؼ��+Y3�u��"��%�hzܟm1��M��_L 4�@�[:,�Y+�{��E6S���<X��n�F��v�B<���{�0ajt
!��u�J���W�OB�ٽ�?�_Ћ�f�:�P�LW�M��Q{��{���Taϙ��/B��3���5Q'̍}uy��9gu_��Bv-UK󗸐o�+3YW<�U�	���Hg4%�S�ä*9����ov0X
��%`.u�t!T����@T����tR���B&Z/#@�dT�##c�%C�0######## $(,h���Q��!=�}k|�5��	 -����mU��ċ�@f��3 48<-@�u{���[Ԍ�=��;���/�P<u+��%��"~�c��%� ~���pcO4�,��N7;��)�L|/�xI�}o�t��ؘ�0J�b2u %� �6V�L(�l��}h`\�u�_)����X�To�`��	�uB* t9�6ދ5.�9�w`'�~��v�>��X��_P�Tŷ�|��VW��}��u�dRfG��-�����V`�v���(m��y(��b'�j�Dz
 � �#
�
�� deflate 1.3 Copyw*�right�5-8 JZ���ean-loup Ga�yZ�� ���m�3�_0y��� � ����		T�}�A}i�i��	
��i����i=�� in�7��(Mark Adler KW�{�co{�{]��wk_��4M�4#+3;�4M�CScs�`�4M��� C2dC$C2$Y�I3 pO���-aw��?!i��i1Aa���iv�@���i� ���i0@`�K8������0!	����A�"�%k�0l���K���g	
	M�ty�L�,�4M�4l��\�4M��<�|�M�4M�B�"�4M�4b��R�4M��2�r�M�4M
�J�*�4M�4j��Z�4M��:�z�M�4M�F�&�4M�4f��V�4M��6�v�M�4M�N�.�4M�4n��^�4M��>�~�M�4M�A�!�4M�4a��Q�4M��1�q�M�4M	�I�)�4M�4i��Y�4M��9�y�M�4M�E�%�4M�4e��U�4M��5�u�M�4M�M�-�4M�4m��]�4M��=�}��t�r 	��SM�4MS��33�4M�4�ss���4M���KM�4MK��++�4M�4�kk���4M���[M�4M[��;;�4M�4�{{���4M���GM�4MG��''�4M�4�gg���4M���WM�4MW��77�4M�4�ww���4M���OM�4MO��//�4M�4�oo���4M���_M�4M_��??�4M�4���i���@ `�i��P0pH��i�(hX8xi��iD$d�k��T4tA���i�C�#�c�i����i����i�
i��i	�i����i�Mw��m C2� 	
�P2$%C%C�}B �2H2���P�P�B�P���a�ݳ[d�� �dHJ�dHTB(*�Q)Z7�i�@7
���i� (i��i08@P`�i��p����ａ�sokg���{c_[WSO�}�KG<�@ un.���zip 0E5D8�-�"	7 )"�a*�AV�7(HP1#@~�.g �/�%c���%<fd:%d> :����(invalid bit length repeat�.T�too�ny����or distce symbols?���eFlock/��2�_tyZPE�eL�*��+l��>�m	/Fnee0ctio��6�nary+rq-{۶�a#h
ko�ٶa7r[w����dow�izSunknn`mp���n2ssZ�eqo ���s`\��b�CT;�}�R p0�4]w@�P
`0�  ���A?�@Ad�X�CA��;d�Ax8�d��Qh(d�A���AH���lTU�Ad+t4d��d$d�A��d�AD��2�\�T�2HS|<؃6��l,2� ��2� �L�� �R� �2#r2�2��b"2� ��2� �B�� �Z� �2Cz:�2��j*2� �
�2� �J��4�V� � �3v6 �2�f�2�&��2� F�	2� �^�� �c~> �2�n�6�.���4� N��I��Q���� �q1�� �a!� �2�A ���Y �ɒy9 ���i)�2Ȳ	�I�� �Uȅlz�uȐ25�e �2%��2ȅE�2�]��2�}=ڃ2�m-�2� �M�2ȐS�2Ȑs3�2Ȑc#�2� ��C2Ȑ�[2Ȑ�{;2Ȑ�k+� ���Ȑ2K�W2�2w72Ȑ�g'� ���Ȑ2G�_Ȑ2�ؐ2?�o&�2/���Jb��O��(J������d��d(J��d�ɩ(J�陆��dٹ�J�Jť��d(�(J�յ�d�d��J���흒�d(ݽJ�J��ád(��J���ӳd�d(��J�����d(�ۆJ�����d(J��J����רd(�����dϯ�d(J��񆒡���q:�W�4�{�[�Y�4��UA]@?�NDsX֯��=M!\ �	Z{�fyV��`�A9�99��a�CN`9��10�C,9�Ompleˈ�dynamic*��_�s tre�oversubscribed'��VK�	ld�G#���e@ty9%�xCs){˖�(=c�(e��i��?���i�?z�#jE��#�a�37����\� ��@3�{��lrbawb�5�����xؐl�5M�\P<,�k۳�at�l��R�k�=buffro�r's�i:t���moW�`�M!s�/萹�*OndتP ��P9
�\����L�GlobalAllocetVU6��F����-fflushκ��printf_fdope.f_;�]*�nomaQs(���fve7y�T�dclos�kmYv&#8s�	��kwnuU���tLcT_;D�r��~���7�"	 = '_:�y�"��&����<���;"�S�H������X_h��n
i��d�D5���l��L������ �+I� ��e����&N��qd5eM���� 6f�?ao�D%`s)-9@�� w����JHI))�g
{����}����j��������m�})��%��V��M��e 4		�	��ݷe	  [��'������ � PE���o~ ��9�� !��T98�:�ׅk�'�q��fg'47�`� "x��u*<���Bu�����dH _�͍.Oxt*����na#�`.r�B�An�u'�in��@.&'���mJ��Osr� l���s�O��R���7%c'�B�C
�T�l      	 ��|$��  `� � �� @��W��������F�G�u�����r�   �u�������s�u	�����s�1Ƀ�r���F���tt���u�������u������u A�u�������s�u	�����s���� ������/���v�B�GIu��c������������w���L���^����  �G,�<w��?u��_f������)�����������ٍ�   �	�t<�_��0h# �P�����# ��G�t܉�WH�U���# 	�t�����a1�� ���^�1��G	�t"<�wË����������$��f����⋮�# �� ����   PTjSW�Ս�  � �`(XPTPSW��Xa�D$�j 9�u����gz��                                                                                                                                                                                                           �                  0  �                 H   \0           `�  4   V S _ V E R S I O N _ I N F O     ���           ?                        l   S t r i n g F i l e I n f o   H   0 4 0 9 0 4 E 4   d   F i l e D e s c r i p t i o n     z l i b   d a t a   c o m p r e s s i o n   l i b r a r y   0   F i l e V e r s i o n     1 . 1 . 3 . 1   *   I n t e r n a l N a m e   z l i b     : 	  O r i g i n a l F i l e n a m e   z l i b . d l l     2 	  P r o d u c t N a m e     Z L i b . D L L     � 5  C o m m e n t s   D L L   s u p p o r t   b y   A l e s s a n d r o   I a c o p e t t i   &   G i l l e s   V o l l a n t     | ,  L e g a l C o p y r i g h t   ( C )   1 9 9 5 - 1 9 9 8   J e a n - l o u p   G a i l l y   &   M a r k   A d l e r   D    V a r F i l e I n f o     $    T r a n s l a t i o n     	�            �3 �3             �3 �3                     �3 �3 �3 
4 4     &4     KERNEL32.DLL CRTDLL.dll   LoadLibraryA  GetProcAddress  VirtualProtect  VirtualAlloc  VirtualFree   free        ��9    7    T   =   X4 �5 �6      �  p  �#  �"     �  �        P?  �4  �?  �;  02  �7  �:  0]  �[  �[  ]  P[  pa   b   �  p�  0;  �;  :  �<  @>  �>  �>  �4  ��  �b     P  �;  @:                                                                              `�  `�  ��  Ќ  ��   �  p�  ��      ��  ��  ��  P�  ��  ��  �              ��  ��  ��  �  ��  7 '7 07 :7 @7 H7 T7 _7 m7 z7 �7 �7 �7 �7 �7 �7 �7 �7 �7 �7 �7 �7 �7 8 
8 8 8 !8 -8 48 <8 D8 O8 ]8 j8 w8 �8 �8 �8 �8 �8 �8 �8 �8 9 "9 39 C9 Q9 Y9 l9 9 �9 �9 �9 �9 �9 �9 �9 �9 �9    &        	 
 %   !    (    '    "           $  = G ? H > K @ A J < B C I F E # S R O P Q  zlib.dll adler32 compress compress2 crc32 deflate deflateCopy deflateEnd deflateInit2_ deflateInit_ deflateParams deflateReset deflateSetDictionary get_crc_table gzclose gzdopen gzeof gzerror gzflush gzgetc gzgets gzopen gzprintf gzputc gzputs gzread gzrewind gzseek gzsetparams gztell gzwrite inflate inflateEnd inflateInit2_ inflateInit_ inflateReset inflateSetDictionary inflateSync inflateSyncPoint uncompress unzClose unzCloseCurrentFile unzGetCurrentFileInfo unzGetGlobalComment unzGetGlobalInfo unzGetLocalExtrafield unzGoToFirstFile unzGoToNextFile unzLocateFile unzOpen unzOpenCurrentFile unzReadCurrentFile unzStringFileNameCompare unzeof unztell zError zipClose zipCloseFileInZip zipOpen zipOpenNewFileInZip zipWriteInFileInZip zlibVersion          �;                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              ]� k�     ��                 P�  �             y� �                     KERNEL32.dll   CreateFileA   ExitProcess COMCTL32.dll   InitCommonControls                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                      �b
s~g r r     �$4                                                              ����                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                  RestartApp.exe                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              Themida                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                               $$$$                                                                                                                                                                                                                                                                                                                                                                                                                           333333333333                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                ����                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    !!!!                                                                                                                                                                                                                                                                                                                                6666                                                                                5555                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                        04-1                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                         �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                   """"""""                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                        qqqq                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                        �ŋ�`�    ]��34��	��U���"�� t���   � �D$$���jE�   h�t���   h%K�
��   �                                                                                                                                            U����`�    Z��!5���E�    �E�@�E؁}؀   t�E���4�EC��E�a�E��� U���|���`�    Z��j5�E��]ǅ|���    ��|����ÈA��|�����|����   u�ǅ|���    ���4�u����  ��7Tx�Њ��Ku���GF��|���A��|������   u�a�� U�����u�E�    ��E�F�> u��    �u�}��E�    �m�E�    �E�    �J�e��E����E�3ۊ0��0r
��9w��0�"��ar��fw��a��
���Ar��Fw��A��
]��E�}�r��}� v�E��E��}�r���;U��x���� ��E��� � p  ���6�GIu��""jI����񎆭8Qe 6e�&�YW��\�i�J/�Z�ļ�>7��\,�����
[?l�(s��\&�  ����4 g�9N[v�Q=т;QFu	.H��e������8Se 6e�&�.�q��  ���w�q4���3u g�?N[u
��A��=��@QFuE��e���b�R�M%���Z4��R�M%V�^���8���8���^Z4�ėe�����&m9���\+�݃u��J�� \��g�ڼ&|HWR����^\����1��	���\�l�Ȇj+���y�6�ag�6��bȆj+��͊�r���%��n�ʌ�`�؂��g��ei�o��c\g�� 5<�l`�j�iX\\�)q��?Z���˯if��$��P�YI��[*�?�x��ebYg��ܱ�Y� a��ɸh(b���i`�������|��;�r�ς��W�ᦊ9|���W����  ��Z�f��oF�hE&�c1g���K   �U���o+Q�nx�@J8�[#2�S73k4�"��k�|��"Դ��(Ս�|�p�x��փ�~g���q��x0}7�9��l�.5�[63nq�!}q~[63k����"9��7=��[63k<��"�`묈�"9��7���Y8�@@3�[@�%5|�gɐ|�77��*8m���[63W��Ţ�3v7 1X63�P���X�P�.5󑞼܍.5z78�x����
8�s���98m˯�[63�ˏ®m�u��`�3=��[633U
�V��6F7 l&63�@=3�[�(^佐-���{�n�8�"=�[63�93�[���>3�[=��[63���~
8�������.5dWx��^t��lH�.5zo��{pt�ɱ	��`�%63� IW�6v7�^0 �k�kTG�m��|�7=|�[63�83�[#�[63���a�襰�|�r��{_�[6i}0��C<�^�@q�r��4�qմ!G"�o��"=��[63�����.5zo�4�x��f��V���d��.5\�}���
8�����"�p��
8��xv7
3�[6~>��ZU�V����Rm�P�"�qFW�7G_����0�~*ľ���m��r����|{̡Eh��H��N�����Ÿ&�g-@H>�:��Ũ'RI+$�yt�+�~�q�BG*̶�W-�7Y8��63�}��[63�"63����U:��?3�[=z�[63�x��7Y8�r/��#63�J��+
 ixHR�V��.5�^�@�73�[�7%63�����.5zX;�x�|� <�Ŝ�k�H�"_9�[6Y��7�W4�V���.5�[63}Ö�Y�Q�Gi�@�m�;ڏ��[63��#BY�k݌��b{���3)�*�7�[6�f�����@3�[&�p�%4*6����5J?<G��39��7��[8k�����[63n�n�!'���nè	�?�k�D�"�]�(63�x:����qHu��I-�9��z~g�8�x`��[6����X���0B#*�Z�[6*#��`[63��F4�73����.5C#*�z�[6Ә�x�[63:��iE�}~�s�/,*�m�Z6�[63p+��;��1�����5]��j5/*�/�[63�T�i�[63�*63�I�Rw��S�n|�Cp����"=��[63�3�[_�[6�J���G�j�*�0Ou�&8�@43�[�r��<��'63�C��>&�fX����ǧ6ݴ#�)?3�%63���3��@Ò{�D�+63�JJ�bA�[�ז�]vNx�Ø���Μs�|�7_�[6���Z�Frk��
1_?��dr.5Ӓ	0��53�[��
8����q.5Ӄ��"_�[6�h�3���x���c�y�ʓ�d�.5 5&63�@=3�[�;��K��֠�=�P�o�䰝[_�[6e�e�Y|�'$hd&i/�\��a�2#*���[6�m�p1�"��
8�}�|���j"0x`�[6��9k�}���|Χd�}G$8m��"=��[63�@<3�[��,�&o�kd9��{,x����
8����"��m���"Դò���53�[��#�
8�~w(n��#�
8��73��d�.5��{�I�	9z_( �@�2�[_8�[6m� �E�y,��53�[�o�
8���l�d��.5}.����.5D+*�4�[6/��?B[ �L�.51-{$�p�^�xAE�n2�Z�4<�x��fL�e0)���1Z63�53�[�~�P���/2�{մɿ\mX63�P�1���h�.5+�[*2���4�.5zg�����{.5zx���H�.5/p���"=��[63Ǡ�0�.5�[63٘oC;�`�h�c8kص.5��'63�$�`&��S:�O�>��).��wnN[6�)oj؆J}�:��;k�@5�"�)`��1���a�k���X8��(���[63(�-�рf!�'0�\D�.�h�[8��;mKױ&� ��-8��Z�j��4;��r�j���3���3N?��Z�kZ63�%63�p�q�����lGÚlGÚlGÚlG�NkG���e�P��T�7s�eG�JÚ.�܋�H]� �9��t���ͧ?8�e�P��TΧ\�PīT����e+*S'��c�;&���P���*u�H���ñ]�H���N��ʿn�BIJ���]�HОkG��LJ�J#ç;�e�Pl�T��S���m��{Q�鉆{Q�C�Úl�Hp�TΚ��ĚlG�?��]�Hj�v�eCf����]�H×�GÚl�#w�eCJ	�
��1����(�lG+��	�cu�G��m<��
�ˌ��lGÂ/����D�p��l���_�e�8l�TΎC���m���jG�:�4�o�,��x�C�mK���КlG�ȝ�КlG����񪆧mI��CÚl�\�Y�GÚ���ȝ�КlG�����bÚlI��CÚl�\�Y�jYoGÚ�V�Z��ZAP�lG���!ȡ��ȝ�КlG����,AO�lG�?��I�Ϳ�O8KÚl��m�;�lGØZAP�lG���!ȡ��ȝ�КlG����ꎆ�md��jGÚ�ƿ�lG<�lGØZAP�lG���!ȡ��ȝ�КlG����ꎆ�mJ���r�բ˧m��L@���ī�jGÚjYoGÚ�V�Z��ZAP�lG���!ȝ��m�Ț�H×�jlnlGfGÚ�J���r�բ?�m�B��=N�lG�+J]�tdr��v���m��,�ė�UÚl�Ԙ�]�tdr�:�lG������+���,�ˉ˚2`˚l��elG��UUi)�(/�:�U�^�|0�
�?��wK���͠VVTg� ��L��#�$y9���-���{����ϙVV
g�6��L� A ,�;+�����8M�� ЕVAX*�61�FHÚlGÚlGÚlGÚlGÚlGÚlGÚlGÚlGÚlGÚlGÚlGÚlGÚlGÚlGÚlGÚlGÚlGÚlGÚlGÚlGÚlGÚlGÚlGÚlGÚlGÚlGÚlGÚlGÚlGÚlGÚlGÚlGÚlGÚlGÚlGÚlGÚlGÚlGÚlGÚlGÚlGÚlGÚlGÚlGÚlGÚlGÚlGÚlGÚlGÚlGÚlGÚlGÚlGÚlGÚlGÚlGÚlGÚlGÚlGÚlGÚlGÚlGÚlGÚlGÚlGÚlGÚlGÚlGÚlGÚlGÚlGÚlGÚlGÚlGÚlGÚlGÚlGÚlGÚlGÚlGÚlGÚlGÚlGÚlGÚlGÚlGÚlGÚlGÚlGÚlGÚlGÚlGÚlGÚlGÚlGÚlGÚlGÚlGÚlG��US-����L��?�,������r��A���Ѧ��BT-�"/��S] 1�;a��-�[�[n���å�VBT+�%.��ST�'y;'����]�AC�E�Ö�A&<����;�&G�y9kGÚlGÚlGÚlGÚlGÚlGÚlGÚlGÚlGÚlGÚlGÚlGÚlGÚlGÚlGÚlGÚlGÚlGÚlGÚlGÚlGÚlGÚlGÚlGÚlGÚlGÚlGÚlGÚlGÚlGÚlGÚlGÚlGÚlGÚlGÚlGÚlGÚlGÚlGÚlGÚlGÚlGÚlGÚlGÚlGÚlGÚlGÚlGÚlGÚlGÚlGÚlGÚlGÚlGÚlGÚlGÚlGÚlGÚlGÚlGÚlGÚlGÚlGÚlGÚlGÚlGÚlGÚlGÚlGÚlGÚlGÚlGÚlG��ULX4�-�E�SV '�;"��3��w?�D���WT,�'���?�+njT�&�5���J������WR*�)�@�  )n�0���|�3���˙�*�3�:� �)l�lGÚlGÚlGÚlGÚlGÚlGÚlGÚlGÚlGÚlGÚlGÚlGÚlGÚlGÚlGÚlGÚlGÚlGÚlGÚlGÚlGÚlGÚlGÚlGÚlGÚlGÚlGÚlGÚlGÚlGÚlGÚlGÚlGÚlGÚlGÚlGÚlGÚlGÚlGÚlGÚlGÚlGÚlGÚlGÚlGÚlGÚlGÚlGÚlGÚlGÚlGÚlGÚlGÚlGÚlGÚlGÚlGÚlGÚlGÚlGÚlGÚlGÚlGÚlGÚlGÚlGÚlGÚlGÚlGÚlGÚlGÚlGÚlGÚlGÚlGÚlGÚlGÚlGÚlGÚlGÚlGÚlGÚlGÚlGÚlGÚlGÚlGÚlGÚlGÚlGÚlGÚlGÚlGÚlGÚlGÚlGÚlGÚlG��ig���?��I�]k;~���r�Ͼ2M��&Ι�UOi0�h����Y�r|/���6�=��Lі��]-�)#��SP�]�;t�(�|�w>���˥\*�3�� ��*�.^�&��]�AV�����lGÚlGÚlGÚlGÚlGÚlGÚlGÚlGÚlGÚlGÚlGÚlGÚlGÚlGÚlGÚlGÚlGÚlGÚlGÚlGÚlGÚlGÚlGÚlGÚlGÚlGÚlGÚlGÚlGÚlGÚlGÚlGÚlGÚlGÚlGÚlGÚlGÚlGÚlGÚlGÚlGÚlGÚlGÚlGÚlGÚlGÚlGÚlGÚlGÚlGÚlGÚlGÚlGÚlGÚlGÚlGÚlGÚlGÚlGÚlGÚlGÚlGÚlGÚlGÚlGÚlGÚlGÚlGÚlGÚlGÚlGÚlGÚlGÚlGÚlGÚlGÚlGÚlGÚlGÚlGÚlGÚlGÚlGÚlGÚlGÚlGÚlGÚlGÚlGÚlGÚlGÚlGÚlGÚlGÚlGÚlGÚlGÚlGÚlGÚlGÚlGÚlGÚlGÚlGÚlGÚlGÚlGÚlGÚlGÚlGÚlGÚlGÚlGÚlGÚlGÚlGÚlGÚlGÚlGÚlGÚlGÚlGÚlGÚlGÚlGÚlGÚlGÚlGÚlGÚlGÚlGÚlGÚlGÚlGÚlGÚlGÚlGÚlGÚlGÚlGÚlGÚlGÚlGÚlGÚlGÚlGÚlGÚlGÚlGÚlGÚlGÚlGÚlGÚlGÚlGÚlGÚlGÚlGÚlGÚlGÚlGÚlGÚlGÚlGÚlGÚlGÚlGÚlGÚlGÚlGÚlGÚlGÚlGÚlGÚlGÚlGÚlGÚlGÚlGÚlGÚlGÚlGÚlGÚlGÚlGÚlGÚlGÚlGÚlGÚlGÚlGÚlGÚlGÚlGÚlGÚlGÚlGÚlGÚlGÚlGÚlGÚlGÚlGÚlGÚlGÚlGÚlGÚlGÚlGÚlGÚlGÚlGÚlGÚlGÚlGÚlGÚlGÚlGÚlGÚlGÚlGÚlGÚlGÚlGÚlG^V�6�N���J���GÚlGÚlGÚlGÚlGÚlGÚlGÚlGÚlGÚ�/,���=�3�z�g�/kGÚlGÚl��lG#eGÚ�[|G�����eS�<�e$���P�cI���Wd�H�!b�H�oTΚ SK�;�lG�<;qe��S��H�oTΚ WSK3HÚl���=dͧa[oGÚ_$n�]A��lG��ZŃ�l٪�lG�zҌY��c��cΉlG�X�������=+�망�H×��Ěl�f<8n7��eG�GÚ�G`qGÚ��I���GÚ��s$��GÚ�=p���v��G��ϗ����D�:���T�:����S�P�T�����eF��lGL�B�⌓�S��l��lG�z͌f��d��cΌlG�OԌ�k��P�TΡ�КlG+0c�=9ҤS�'nGÚ��ÚlG-�`#
�G^qGÚ��G�,��GÚ���+�<��ҾP��T�<8�J͚ۢlG���4�D���n�2Bm֤ęH��I���6@Гe�P��T΀lܪ�lG�zٌZ��c��cΉlG�[��>������(�lG�L�Q<�YZJ���
쪖�jĠqjT�����e��� ����e*:�N�ȗ�CÚl%D�<T�x��kGÚ�GRqGÚ��S���GÚ�܁�h�I���,�L�J@�L^����>�W�e ��T�7 ��eJ�GÚ�˜o�HB�o@PxlG��GÚʘ�*sy���/;���6�;�lG��ŷ���H=�TΚ�û�lGjGÚ�-�[�lG��۟lG�R0LV�CDN�C)�lGM0�I{����H#�{7��d��H�nGÚ96襶%D��A�jd��nTΗ�IÚl%J���pY�H��ܟlG�S0LN�CDN�C'�lGJ0�u܀�/DyrI	3a�.H�*>���PաT�K��͚lG#��]=w�ϚlG�":�1���np�\vuJJ��٫�lG�T���&?�3�/���^�0-A��t�2�LN�CSH��җ�a�GÚA\�!��<�"�)n0u3�w˗�'$P�[R��<řH��lG��y\��>�^
V����?��el�ՒT�|e@F�m�)�՟lG�T0L&�CDN�C�lG?0<�V�ꈶ#��e7��e�P��TΗ�IÚl%J̝��7,��eJvGÚ�GTqGÚ��U����GÚ�ځ��O�/-J����Sѓe*�S��!�JCMÚlgZ���np�npRÚlS���7���*j�DDÚl��:Y&I�_JN�CI�:���k���c��R��ߟlG�F0L6�CDN�C�lGA0����#Uذ@ՐT�m7D�e�P�)f�fGÚ���k�2���H���G]qGÚ��T�4��GÚ��4Ɓ���g��G#�l��e*��cִ|�HB�2F�k@PlG���_�e�P��T��]�h�lGJ	/��@P�lG��[��n��[e�H�~�� w�H��s�kƘH[�l��lG�z׌h��c��cΆlG�QތM�,���k�T��eĠ̓T��G����f<�F%Hė�Úl�͚lGlnii����IZ=�����HB�X�l@O!kG����b�(�m�͚lG�Qɴp�CÚl\���;�n�Z�<�3�R�Kl� ^�H��۟lG�R0LV�CDN�C�lGM0�}��E���elG�S֐��������-ZPBֆ�m%J�%���HĚlG-�L;���GRqGÚ��S���GÚ�܁$��J5.�HCGÚl��A��I	7b��#?~�mGÚc�$o�H���G^qGÚ��G�,��GÚ���/�G��#����ʚlG#�-zD��or���-��S<藓�l��lG�zԌ[�c��cΐlG�ZیA<6�Nձ'-�q'D�,�i��Ӝ��H$=��<Y�H�mGÚ��q�H�<9��J��#�JCMÚlgZ���np�npXÚlS�N�\p�ΰo�H��f��� ��H�6���ڗ�CÚl%D�p��� W�#��ܰ���X�e����X�e���m%:�!�MCMÚlg[���Wnp�npRÚl
Tۚ-��]��lG��-FW��*?���e*��ܟlG�S0LN�CDN�C�lGJ0Z�� A�S��B���T�pGÚ7��BÚl���p�&BmN��)�uR�[�np']J�@�Q���lGØ�G���"1d=����m�f=�HA���2C���oGÚ����l��d�H�`lG��)ϴ@�����P�)f���0�:l�)��lG�P0LF�CDN�C'�lGK0њo���DN>���X��HI��6����e��۟lG�R0LV�CDN�C�lGM0�/p�&J�DDÚl",(��lG�yZ���d�a{mv2��i�S��@Úla��'$P��np'SH�����:SH�:iR�SH��ÚlGm@iR����_�np��RԼP�D���T��`+��Rd���ϚlG-���)���� c�H����|�HL�X�CEÚl�+G�Ш$�9����:,��d�*-S"�LCMÚlgd����np�npXÚl]�N�DLu�ϗ�\Кl@F�C�ÚlJ�}oT��>� �e@L�lG��>D��eʍ�G�7TeG�GÚ��CÚlĨ�T��G�GÚ�GRqGÚ��S���GÚ�܁��㪭��<�C�U(#��Y3��lG-�y*�~k�[��H��s���x��H$��e���m�C�
�͝lGÀl٪�lG�zҌY��c��cΆlG�X���n�x��_eGÚtӀV笴d�IÚl%J���3Y�HЗ�pÚl!�JCMÚlgZ���np�npUÚlS�╚:�~��eh��w���@U�T΀l��lG�z֌e��d��c�lG�\Ռ�ݬ�<.kGÀl��lG�z͌f��d��cΌlG�OԌ�h>j�M�T����GÚi�L�H�IkGÀl��lG�z֌e��d��cΉlG�\Ռ+k��4ÐJ��\j�HJ	�J��.�؝�ƚlG�~lG�}��a����W�J�-�j�b��L��̗�HiP�%:�L񭆧㻀��H�llG���e�@��T΀l٪�lG�zҌY��c��cΌlG�Xጔ���@q�T�e�˓e���lG�P0LF�CDN�C(�lGK0d�J���Ǉ����㳐e�H�jTΚ��E�lG-)y:����lGJ�.�܋�H_�L�ϚlG���J��%:H�np�̚lG�T��_��5�k�np@B�lG��Q��fW�m��n�HJ	�l��Ê��HJ	G?�m�)��lG�P0LF�CDN�C�lGK0�{_u��blG�@ڶ9R3�S�GC�l�@�jT��U��� �e*nGÚ멵*J�c�%Ǹ��HĚlGAW���vv�P�A�t�`�l٪�lG�zҌY��c��cΆlG�X���L����X���e!�����e��!�T�oGÚBh�*J�����oc�R�PыTΗ�;Úl�˚lG�X�9ʱ�ڝü�lG��ߟlG�F0L6�CDN�C�lGA0FR*�L��䶐eS�x�eZ���e����﶐eJÚl%Dː�B�Nj�l@OylGÀl٪�lG�zҌY��c��c�~lG�Xጯ���e@D�lG�<�y�H���w�H×�PÚl@Q�lG����e���T��<�e�H͟TΚ�ú�lG�+k���řH×�`l��lG���aC�oyK��t���#���Sٰ�1�T��H�e�H͇TΚ�ü�lG��E�����H�ZkG�`lG�r �ytB��3�˚lGG	gT��Y���eL�l�җ�ʢnz��f�e�Āl٪�lG�zҌY��c��cΒlG�XጃndD��=Úl�ɚlG�
ah�wIMbCBÚl賹-��fk*��lG|��G�$$+��IL]o%I*¨MnTΗ�Ġ�oT��g�e�u�G��lG�+�T4'y�椝Ark*��lG�Cڻɨ�����֖�K]o 5jT�7%�eGcGÚm�PÙHC�M�H�TΝ���lG��W�k�癙H�_lG�cGÚ���Ih %C��nT��>�h�e�͚lG��>Dg�e�͚lG��5�#�췐e*B�2]�l@O]jG���{r���v�Hė�yÚl�����W�eBH��TΡ.KÀlܪ�lG�zٌZ��c��c�lG�[���칛�B��ƴ`�H#��eJH��T΂�d�YD^�N�]��4�w��CÚl�H�΃���xw4nI���\����lG#�6,�e@B�lG�=ʢ̚lG�	�8�r�V�P�e�����W�e!�ACMÚlgg����np�npUÚl`��+�;�gvJ���lG�P0LF�CDN�C�lGK0!��e����o�Hė�]l!�MCMÚlg[���Wnp�npRÚl
T۫O_���"����eBH��T�=�)�۟lG�R0LV�CDN�C�lGM0Du����&�7��eG e��ۑ�H��R�+�P��T���C�e���3dͧa[7�ГeG����IoX�����H�	���m\ZR��VS:��P��+E���T�7�eG�GÚ�GTqGÚ��U����GÚ�ځ��}�L��oGÚ���%�H�nTΚ��͚lG�+@���;v�H×�Úl¨e�T��뤁7��S��H×�nl!�JCMÚlgZ���np�npKÚlSۼ���>��^�HQnTΗ�@Úl@��lG��[K��pT�7�eG�GÚ�GTqGÚ��U����GÚ�ځ3d6B��E�l@O`lG�<9�����e�H��TΚ��Y�lG��ߟlG�F0L6�CDN�C(�lGA0�V�p�����7 ʓe�HQ�TΚ���lG��՟lG�T0L&�CDN�C)�lG?0�Yy(6,���;v�H×�jl�@��T�7�eG�GÚ��^�H�wS����+��2��7��eG e��ۑ�H��R�+�P��T�����e���3dͧa[7�ГeG����Ig���8|�H�	��m\ZR@kH����+�ʚlG	����q�C5�H��TΚ����lG��b]���w�Hї�rl�T*8B�BA�k@P�lGÀl��lG�zԌ[�c��cΐlG�Zی� �q1�t=�T�7(ѓeGIÚ�_�G{:�ˀ��HJ�����lG��lG��s!�>1`D3�k�Q�#J��lGQ�B>ls݁%��r�@��U�"�$pch��vS<����!�<�|Rl� v�H��՟lG�T0L&�CDN�C(�lG?0(���1uK�E��¨jT�:�G`qGÚ��I���GÚ��@ٴ__�%S:�L�~_��J����H������HL	Wk���Q�9wzpc"��v�B�CÚl��@ڶ9R3�ՅC�+��w�m!�ACMÚlgg����np�npOÚl`�,H��lG�J:��&���<qӨY�]��!�T�H�YY=⻴��H���>��GaqGÚ��P���GÚ�فȝ�lGC ��V��ʩ\�!ĝ��e�bGÚ�@Q�lG��*SoGÚn� �ϚnGÚ��T��H������8l����g�	#X��L�3A�':����ȉ4�1��|e�@��T�<荆��GRqGÚ��S���GÚ�܁(�Z!<�W����r�HfT��GÚARp��d��e�x5�V�Ĩ�T�P��&�lڪ�lG�zӌ\�c��cΒlG�]ڌ��P�𰈗R�J�dlG�0�m�ߓ�i��,���=W�<�Kˢ�lG�%ѯ�m.�?�J��6��e*i�|e }gTΧ\"�?CMÚlge���np�npOÚl^�?��;�¨��T���gI��zـq!�HCMÚlgh���_np�npUÚl	a�wQnGÚn0��QRS����gc,����휝�ΚlGS<�.'ٰӀlڪ�lG�zӌ\�c��cΐlG�]ڌ�!NS�3x?݉T�iGÚ���F���Q��gGÚ,��yW�ꗱ�#�Ę�T��íė�FÚlĨqqT����W�eĨ��Tδl!�ACMÚlgg����np�npSÚl`�7��e�T΀k�O�`�;�՟�lG�P�m�AM᥆��2H�ipc�b�I6����&|e!�JCMÚlgZ���np�npVÚlSۏ$��j�m���b���;��H×�{Úl!�MCMÚlg[���Wnp�npNÚl
T�"�ُ�H�s��b��������HB��a�k@P�kGÀlڪ�lG�zӌ\�c��c΁lG�]ڌ��9T���CXÚl���X��%f�:�L��P"��GÚ~�u�԰�h�6��1�k�˚lGS�~0l�����I�mZL	=��JC��!ė5����~e��i���H�z���mU�TΧ4��e@��lG��<�x4IÚlĠqT�c,AO�lG��0��eĨq�T�7��eG�GÚC?Úly�bRv�!��'��S=��GRqGÚ��S���GÚ�܁�p�Y���A�)C�"AM�lG�?�*J	�c���d��HC���,���lʂ:�۱S�E6?&-S"�LCMÚlgd����np�npUÚl]�6տ���e�����V�lG]��{�e�XkGÀl٪�lG�zҌY��c��cΉlG�X�ccv�!Wʃ�ut�@�T�Z�M]�ʍ�G��nGÚl���Z#���͚lG��L���{����`lG��ߟlG�F0L6�CDN�C�lGA0�#�V��Γe%D�2vA�k@P$jG�Js!��lG-�TE����Úl%J��ė�Úl:PA�T�tL�GÚ��q��lG��ߟlG�F0L6�CDN�C �lGA0��<�[莘��/Z��G^qGÚ��G�,��GÚ����?@��T�hGÚ���Z�^�x���bm�C�,�ÚlG��f����5�G��ߟlG�F0L6�CDN�C�lGA0$L��P�m���>����7x�e!�ACMÚlgg����np�npTÚl`��u�O<�F�B}Ěl��lG�cd���,����5[u��HU�eFÚl�&ZF��ϚlGnGÚ�Ƽ��H��eG���g��e�{��Ǝ�lG:%���kGÚ�ˤ��H�ڝ�K�lG�pGÚ���tJ���CFÚl.�F=
�tLc����G]qGÚ��T�4��GÚ��6�T���� X�s��lG��lG�j��Up�w�JZ�75�Sk@Q�lG×GÚl@O�lGçE�`�����YUv���lG�J���lG�elGØV�u_����{����lGL�L���GO�HC����lG-�T�B�o@PllG�:����HC�6+Lkh�C�͚l!�?CMÚlge���np�npOÚl^ۯ����{���ȚlG��> ���lGC�-�!�lG���lG�P0LF�CDN�C'�lGK0�'HV�P--)��tH�GÚ���m�HJ	S^�C�Úl��tA�GÚ��٩#�H��T��t���lG2��!�JCMÚlgZ���np�npOÚlS�����¨�T��>�ēe�@udT��xLN,�˄��HBgl@OFkG����e�˚lG1�z�(�J��w�l��lG�z֌e��d��cΕlG�\Ռ�:�p����#�˚lG6�X��$��L�e�c�m�:ƞ�G����6�W�e�@I�T��3͓eJ�UjTΧ?�e�˚lGś#`��o	���ܾH�T�����e�F��ꤼHӢ� ���,6�H�%���r���;�lG�c,47��eG��m��k�HJ�����C�H����X�H��%���HĚlGJ�b>���_��HJ�>k�����l:@�oT�:j����H-��:��7��H×�=Úl%J�m�t��H�	�A�����H×�Ěl�͚lG.���e��+��Hė�Ěl%D tA�`�l@O�kG�oGÚ䶂�'J���Y�H×��Úl!�LCMÚlgd����np�npQÚl]�C�^�{e�K�e�P:d���e�@E�T����e��Z�ASօPաT�>�G]qGÚ��T�4��GÚ��(˓I��K>��˄��H��lGÞ6��<�S<�JN�CSH�ymD@Úl1e%���a��[P�J�����cΗEÚl�I����՟lG�T0L&�CDN�C�lG?0�[�a���]�S�@-�T΀l٪�lG�zҌY��c��cΒlG�X�Ei�]�dGÚ��c"���*u�H-�Қ����d{�H���~��m�@��TΧ\"�?CMÚlge���np�npQÚl^۹x�ul7��AÚl@P�lG��Fn�@L�lG���:�y��r(��Fe���,j�H��X��G]qGÚ��T�4��GÚ�������Z��>�W�e@F�1"�JCMÚlgZ���np�npVÚlS�:3J3S�A�J�
W��ʬ�ý�lG��ڟlG�Q0L>�CDN�C �lGH0����IÚlǊ�!dT�=%F��_~g��4Y�HC���{���H�lG��ޟlG�U0L�CDN�C�lGL0;�f��>�̚lG��/�H0�$�e�lG#��[�e%: M+:���tG8IÚ�GRqGÚ��S���GÚ�܁������l!�ACMÚlgg����np�npVÚl`��L	<��÷O�H-�/��cG�<�S�E��nc�`��H�:��ߚ�H]<�e=3IÚl@��lG�{H��e��|C�Ěl!�LCMÚlgd����np�npTÚl]�䍟d���͚lGJ	C?�4HÚld��T�Js�������HSnGÚ��մ�i4IÚ��ÙHB�j@PflGÀl��lG�z͌f��d��cΌlG�OԌ�t��HŮT�dGÚ@#@�[/<B�lĠ�cT�tL�GÚ�U7r��6�9]���U�lG��`��З�ml!�JCMÚlgZ���np�npQÚlS�ߔXU�&��<Úl@O�lG��x��e��lG��zd��ʁ޾���xLN,��x�HBgl@OnlGæ���řH�di� |�Hԥ�(O5w��m������e��tF�HÚ㻐b�H-S&I������	�lG�`lGê�,+��!OV˩����P3IÚl¨��T��GÚ�GaqGÚ��P���GÚ�ف�-�s% ����dřH��@�m�J�CBÚl���yL�T�7�eG;IÚ��̚lG�pGÚ���JA�L��2���Epl����e-I�т��5�D��\F�e�КlGs�9�Χ?8�e!�KCMÚlgY���gnp�npQÚlR��%�;柾�t �e�P��T�<�y�Hl��X�PU�T�]�[�lܪ�lG�zٌZ��c��cΒlG�[���a�P���̓e�H��TΚ�û�lG���lG�P0LF�CDN�C�lGK0�tkA���Fe��� }�H��X��Ӝ��HB�l@P�lGÀlܪ�lG�zٌZ��c��c�lG�[���m-��dlGÒ(����G��=`�J@�pT�P��#��H×�ilL�ͼTΧ?(�eĨ)�T��jGÚ�y��i��jGòm�wÙH�	sU��uw����Fe�2�a�Ͱ@U�T΀l��lG�zԌ[�c��c�lG�Zی�!��L�v����d�H��jGÀl��lG�zԌ[�c��cΒlG�ZیO�������eJ�㻸řHB��l@PdkG×�PÚl@��lG�gGÚ�L�4%����Z�+�PաT�YBÚlIt/�m([&m"�h�n�pGÚ7��CÚl�@�9�Y	���}�����ԙ��,�Ҷm2��8�[S�a<�m9�{n[�c���g
{�H��lG�Py�Tl�T�����+D����rPӢ�lGv^%���'��?�7��iư@5�T����e�@E�T��!��e@J�lG���%�e�Ӏl٪�lG�zҌY��c��cΌlG�Xጾ��L��9S7��lG�~lG��H�\��C�R%~��Xe�l�eJ	^���kY�HJSV�i��GÚ�GaqGÚ��P���GÚ�ف�BÚl!�HCMÚlgh���_np�npSÚl	aې��)���X�CCÚl�4"�ͻDL�P���C�H]<ꡨ<��GÚ̢ʚlG�]�1xl�0�*C($=�D���e]7�_�e���Q��7jA����\�%��eR��#��H�eĘqT�k#�lG�ڝÜ�lGB�T�l3ͧ���e�lG���?B�:��k3�7�W�eI d��kY�H���m���	�m�B��]�j6��@�e�P=�T��oc��H�kGÚ��7Y�HJ�>k�4HÚl��IH��H�kGÚ��˙�HJ�����?x�H��*<�7� �eG����s��H�e����T��>�W�e�)��lG�P0LF�CDN�C)�lGK0N�|�������:��Jb�He=9IÚlĠɕTΗ5�`�G�]H��b�����Cgl6|k#�bIm���UC ��s$�āK8CÚl�Q�A�l8{Sp[O�D�!RńT�\�*D×�FÚlBPE�T��GÚ�Ս6����*���׺)H�C�^J�C�ÚlGÚl�#lGÚ��x��Q��>`�e��n�Ƨ�lGJN�CL IÚ��c��o�lGJN�;B�d�M�kG��c�+JN�SL�HÚ����O�lGJN�KL\��n��*Ż�<�Ư�lG-T&LNHÚλ�<�ƫ�lG-\&LBHÚ%��lGs�>`�e���E���W��CL\��n������qGÚ�un@P�m���C�����z�HL����3�HD�xPÚm([���e+H3ᦧ?8�e�P��TΧ\�P!�T΀�ÊlG+��GÀl��!�T���h��e����T��d��e�P�T�7G��e����Q�������j:��$͎��@P�m��?G��e����Q��]ͬ���I�C:(`lGÚlGÚlGÚlGÚl�Úl�dl( `lhÚlGÍ�GÚ�I_�bG}�lG��k��cl��l���O˚qQÚkC�t�;��Gç�J��gG�lG��j���l�l� ��ʚ�RÚmu��`E��Gç�I��iG�~lG�{k�R�l�l�䙇КTÚmr�`�L��GçdI��qG��lG��l�al�l��v˚yVÚm:��NC��GÛ�J��cG~~lG�uk��l&�l�Θ�QϚ�SÚp�P�D�?�Gç�I�	jG�lGІk�vel8 �l�����KPÚn;�du>×�GçnI�nG��lG�fl|�l��l�왆�QÚdT�z�B�ęGç�G8TiG�lG��l��ly�l�Ϙ4�˚SÚca�)S<�,�GçcJ�)qG��lG�l0}�l��l�Ν�̚bTÚiD���A�S�Gç�I$BkG��lG�l�ܑl�'�l���К�RÚmg��qL�e�Gç�J6�qGܐlG��l�Ccl7'�l�&�N���QÚmB�3�I�O�GÙ�GEGoG�lG��l�cl��l=���Ϛ�TÚmW�0�E���G×�I�,kG�~lG�ckeE�lQ�lW��{���SÚmj���F��GÍ�G��iGI�lG�al���l��l��xϚQÚm]ß�A�Q�GË�ISfeG��lG�lj�kcl��lS��v�Ú�OÚmA�^2<���GÁ�G4fGslG�_j�?�l��lU�	)К�OÚm=ý�J��G��J�OcG�lG�rk�ؖl(�lO���OÚmk�.C�)�GÕgGU.dGQ�lG�^lTk�l��lQ���R��OÚmQ���I��GÓ�J7siGF�lG�}l�Y�l2�lKŘ����4TÚm9�d�H�ȞGÉ�JckG��lG��j�b�lh�lM��D(ʚ%WÚm`�#<å�GÇ�J�]cGg�lG�xju�`ly �lg���FϚTÚmaМ�I�9fG�}�I�8qG�dlG�tk���l��liȘT�̚;<Úmc��OG�ɞG�{�I)ylG�lG��k$��l��lc�>a�>Úmx�00C��fG�q�G��iG��lG��l⥘lZ�le���˚�=ÚmJѬ�?ô�G�o�G,�hGόlG�^j�J�l��l_���̚�UÚmSѻpI�J�G�śJ�xnG9�lG��j���l� �laĚ�К�VÚml�HD�˙G�ÞGF1nG��lG��k��`l��l['�q�Κ�OÚm`«gC�ΕG�y�G�5qG�lG�j%ӛl�l]̝��ɚ�QÚmdЃ�H�z�G�w�J��eGO�lG�jj$��l��lw%�z>Ě�XÚmOérI�F�G�m�G�dqGO�lG��l�ޏl��l9�HqʚWÚmIĽK�2�G�k�JzkG/�lG�vl<��l��ls�P�ʚ`TÚmt�+PI�
�G�a�G�lpG��lG�kj�xcl�'�l���T̚�KÚ��oqG�z�Gç�I�zhG��lG�yk�K�l�(�l���ΚNLÚm:��EÚ�Gç�J׫pGJ�lG��k.j�l(�l�����͚�KÚmx�<F�k�Gç�IxdgG��lG�^k�<�l��l�˝�̚kTÚ�d�QD�s�Gç�G��pG�lGɑl'6�l�&�l��_���KÚ�G��Eê�Gç�J5}jG�lGǆj�el� �l����͚wVÚm`�6}?á�G�ijI��jGρlG��lxQ�j�I�Jgnp��	g�B�|�^x�νq��fHL�1�ϳ��/�;��E�	��oIr�¡��ѝRD��?��G؆t[��1xЋ�L�0�RBr־�%F�'Y�D�m\c��|GZU���Be���\S�o.p}wx�I[�T�.8Y�Yx�a��o��Nz��]p�<��I��9̺�ML��Cs�l��j����P�cY�d��f�&k��+���#��ft�O��Qiǲ(���d�A��^�qܽ,�l���jT�abĺ�]~m5�Mj��W�P�W��[�J�!�7Шd��;p=�։�\�p�Z�<H��ﲞ~WQ[rJ3	��nĀ���yeF�b������.�W��kí���n�O��&I=~�Cj�������v���nY��}BᛚJ���	"0$�J�Б�F�nbzG�h�F	�ܫ��Cx�f߈ h�j�k�-U�J�u5i�%��\�?.eR7v�y��jS�H�Dۢ_� ��������<�a��i�G�.@V��B�m���C:izCk&�7z�|��xa�N�����6�� hm�G툪��k��k� o��i3�q�\אuhҢ�b�C��QR��ɏ�����8QwǙoC>Yk�BW�I��:r�G:L
��e6!��k���{k8+n�I��}jW�t6y/�d� �ǟ���S�;PC���ajY��,iI^�������s�)S-M>=�q�솭p�����]�K��bqT��{iJ-�������@�~���7|Y���F��F��[�)��ʫ�l �`2~��h���Vg���"�)��'KBV�j*�8�e+~I<�P�PV�����^P�qNn��9K�v�?��t�Tg��QʭBOa�_A6H����������QR��dFam�&��h#\�AiZh>Dݯc p@��[#�������E�OL�%�c�����9���k���ƨ:�㵀�f��\��nqFP��+E���dz�I9G��lI�����\���&x����BR���A�h��n���ϑ�����ʛ
p,��Or�;��<\6@��ߡ?m=�c����M��X��9LC ϥ�J��>o��d��A���Ӹ��X���t�7��B����J@�^M�.{�٭IK�ւ�8��x&P)��:����6q�{�K�@�Yl�S�A���|U�0鈘�Κ�(��1}�ѝ�eY�Ytu�g���o���0LK4vQzprà"�͚�#����vN��k���D����n��
ڭ�͋�_�5���{bZ�ZCh(�m/�<�3)�ɂ˫��Ta�A6��_�̪�S�%�^�31<I��ܡG;��k�obly�ĎV֚"�y>�ETCW��rjJn��c�����y�oǣD�E�ӡQM6�C3b�kr��O�}����v�,L�M�m�{x�!�N��/���ak���j܃d>�?sǖB��p̺��Sma�h�W�*�F1Β�Ry#�ڈ�+	��F��IW
A_�eo�k�h���j6�cU#4H��\��eW��X�D%��iH���␈l�鄀��HQ���](U����lk��k���'�X�T6;{�kDc��b��q�I�S�'��UgH� �4�ʴj p0ex���jyl" sJ�d|��FC�s�2���Nic�"�hX�/Ӏ���ԪK��fqf=�p�o��nVf6�2!Ӹ���Y��7��~\@���NI��ګU�H�iwLk���~maM����b��.��b�#������V����.��[���[�B���cF��E�����g�f�AEqj���3����ĝ�F;3�P\�Ąx"�"����Y�o�ŧ��HeH<��x1,L�mz���~�Ù�G\jQ�;sV�W�1���QǼ��6��*n�-�+̎k�@�!�.'uN+�e��H����ݱƙj�x��텛oG*Y!	ĪCJS�ɪ��t�xt%4�.nk��~���+���:~&T�7#�8nZa'�.9��`�J��h�̎j�x�W���W�Q���C1`۞�F��bUt�����A�C��OwO�,�d|��e���kH�4VW� �O���d�*>�m�/���5�8��̥��[�n���~��Da/YD+q�~�^Ku��T��]�bJař����*nz�oz�.;r�k���B� �i�ڦ��o�+$6>ҝ��0�hrA��Ud�}@��Mі�7h��b��M�����)a�����GU��wK�]�/��ELҼv���L�^#�}x`�'L
�c��;��I��5׹㡓h[1�3NT�K��8B5��G\!f1� 3O��I�ɸ��k�;���6ʚ��q�T5DN���,��,H�;�T�Pic��9����~=tk��R3�l*{w�?m��:�K@�������l���0vn-�6�7� W���j����_p2�k�-Rþ�w]�9"�򝒗�e�O����l/7'�s���o���gI��q:x��E/M�s�]șCH3J�����uW�aq��A/;3�8n�Z���3V��
o�'�_ó�IkS��yЏl��r���:@B8�����u������^.}�_���i2Ӌ�>����'�S�������|09��[v�x�L��U�X�9ۈ�m���j�[NC���g�I��poۗ����Z(X:�$:�b��Ľ��Ӌ>�[WPu�>n��\y�Ms���+W�&�~}�@k���0l�H+NWvP!9[��b`t�qH�kN|9�g�k�a������(K�xS�t"����2ݔ ȅm�w���|!�-P�xm
�����`�n;�ל4[o% ���Q��B�8�R?Elܦ��:��}z���õ�)���-ϊ�~���RJ~�C��~�V|�����0ӏ�P7���������"y�@^VRpo�̝M�7~����2��Q+��=t����[zQ�[��b�w�Ub���B����j��b��n��4�}��FEop`B�8B�i=�����8�@�v�l�W<��}ix$�VǇ��M�O��n���D6�j_��Ӝ6a�&H�䬺eK�iX_ESse��k|�f�E�$Te\Ih]X1�b�A8�c������TЅK�ˢ�
9M�r�|K+��`k
�MG��/���*J"�����w��N�)ɗj�5ȃxx	?o��� ���s�/�D��<�ˢEtkiy�D�T,p� oTDa�hG�r�g^!c8[H���5��\��:�z
��f���9C�Wi�*�+���)O@��$Њ�i̎di���6��&�%o�Q$r�BX��28�:*���lf���t6�E՞c�؜��"�J���=�[�a�K�]�Ȩډ<��H5��I�C���)�̧��RF����gE4�<�;F`�b�:�.�_�� h�0��7u�<�����\��M��7S��܁�k�$?�d���R@1�k�{��$Y� 1�F�1��4�Jϥ�1�������bcC6"!�jx�hV���u|�p�+M�̇�kbJiS8��5�7���<����c�[��h�grV�IB�/��c��wjÎ#�g#L��_�j�Xj�m��м>��f4Od��:؟�Rs9���c�wT���(fQ�cG����8ϔ�yf�#�R
�����i�T��/�b�Z��t���킝s9U5/��Fޤ�f:��F%m������e��L����uhjS�9�g��v�e瘙g/yL�h	��O�)P:h�	~g�j�� _z��@�m4��"�-:��n�(��.�����GF�OL�sFM��c�\����Yا�c�T���3TB�.n��:^����F�/q1;�&._ �o�%���S�9�I�/�AC��T	J��\�A���E��:U���Zn�)�/u�?�ŷH	A�X)�Rj�K�x�Փf㇧�ˢ�o�
����~�a��d�L���^`��s��:�x�mj�u�C�)`�)ߨJ�;�Y��:bѷ�K�W�:�U���_
�H�4M�uC�I��a��̈́���%0��;��:?����>Z	���^��w�_�tס�g���i�&�/�}����O~�z��������ʀBc�򪛿V�{�Z�-�܍�J��ږ�f�q��� n'�����U�0��c6����nD���GT��3�[��bf��Z�c˦6�k�I����C�he��Li��8C�����J��C��o�|��o�t]�ꄺy<�n�Ju�=��U��5R�)&׻�*b�+O�*x������v[�jb�.@�7�GF|dC��aV���T(G=��JJ�j|�C��J���Ё	�A9�c޵����z��:�jj�b�L���/\�E��%��:��g�ne�z�؏��R(<�2��zz\i	���(+zص&���:�q�U�*)[(��[�=q����yɤ�GI�ڂ��_nX���@����w
7J�j�Zp�'�m9�M�^kq�C�'��r�O»�\�e��/��3g͎�ZYD�ycv��"���c�\0�Cc�� S;�Vk0R�_�i�#h��Z�I�'a�k�g�NMi���}�F��=���@�n�%��4���\C�nJ3�
3[Z��v��:޹Z�;5�|T5P�`ҔC����^l����yD��+]�\c;C~�:<�u��B!_�.���cj	H��e�:NxQ|��ӛpkL���f�mBO;fF�l���)>`�B8~���Q�(hЫ�im�9E�v�C��	�˰��˻nXw�$��C )�
G__өl"%O��ѨJY���ĺb����%��G6c9B�B��Y1��x��z���g��;7<���xq<�ϗ��~���&>��T���yׇĀJ�� �p�l\�S��:qѴ��I��f�4��q{��w�*gm��;}�fs�PY���Gb��gM9D�kg�t�v��$�ky$�?��m��}�`e��*Ge9`��`3�d��1?�~�Y��Z��}�FWʚ������S�r��0Sd��GB��z_z����QM}����rRbXBj!{�zJ�7��%ex���C �F�?��/C`�Dį��e��BTefv�a���������W<�J�u�k�G�1\�h�s�G��ۢ�6n�:�
�Qzw�UC[����Z�H�IWu�=�z�eC
�R+��������KhOYY�{������J�w;&���x�ɷ�jٵ���X^�?Z�q�> GcK���h��B���&o�I�J�R ���Si�@� ���}Y��G��"~�MI�qy\�B2� u�o6�1�kKfmy��bu�����Y��9W�_=��m�τBټ�"Z�9n�jw�*��M�c�dh�n[o�!��2�Q-{J��v����Hö�]d�fzǊ	����˳�Cz����sw)~����*}�'.�O^��j�ek�̹j��T���㓩�Tk'�K�3[�+��p"�4'���3��UI�.�od �G`�h���^Z�-l�+	�>u*ߎ�uUAܜ�Q����o�Q�g��EA��M�T,����c�~ޯ�J����)��Zv��|U�lR�J�)UĔ H�A�`Psi�\^h��߆�Jcc��q�'G��>6(��C�Wu��B(�s`gC�# �&���=�l���RYfc�JF:Z�V�-kv�TP�|Rk,�-
�t7�����,�&r�kv��%��4]tS�ǂjzR6���9��F)�կO
�O���H��[ê��4�W�ُ��D�J�c�쾬2��ILHj�0B+�+���I���u *J���M��.�}&jc�OF[�n~?f�$|O{��V@F���
NZ��rU�q�[��?��oAF��*qHKlE�%���'xN��� �m�u���]�� �)�����[#�^shi$��D+���Z�2(j�˵��?���I�r�ÒF�����߉0�7[��Lz�R�?#r0��B{�����A.)���AT�K�oU2��)��C��y{b$�.W���Y����a���sR�1| kDҩGc9�ڍO�'��'�J���3��fF�e΋�8S��Rx���w��N�u����vs�i���ed�*��+Z�,Q�P��E*�\��Um\0����7���,;`�v�I�/�u&Z�����d������g��j�hQB��UvT�0���C�A�p�r�C��jl����Sh��)�=�����y�ȶ(�������*������-2L�=�Ju_ט@�>"띄�E��0�wݡr[�}� �ikE���:���s��gB�GIV�j����w��D�.Ѱ��N�)�}�"	|�%�d/�c.�B��&[�F���%E؃�[F/ ��um;�"cfo�Re��<ou+��R��AE�q����b�IIZ�MLѪ2�#�`[5�G~_�}���v$��f�z�^��sOZ�Pq�kS��*��.�Dc���~� ��=sز�'�u��UȺd#cim��w-�	hͨ���i�jiIR�d���U8D����>�K۳;f]U��J��fC�����_��M�iOx����~�z}_��l%u_E:۟nk�9�7�nF�yk��5¢7�@�v��Pj�1�v����:�;.�B@J;{�C�P��<LI�!��4I��u���"i���������=n�c�JgGA�m��}f[Ɗ�K�cp�e��H��A�cl3���'�$�h��k��]�C�s��EK[�'8:w�WRߦ�ƥ���
�Kma���Q�:f�����S�����������
��^Px�˩36�@t?�C�plj�b��+��^���h���(m�����:7�OZ�_�6��kB�9�,c]�1��޺ue|�fYT��MQUB�,�z��:�p%������iE��^�Њ�t�}$r|��v�Qy�U{�k�C�u�/I��poA䝰H�p��<�pGm3c�e��X�)���wS�i�Yh�yd�	d�����g���;Y�JѰ�R��,Zb�u�k�,ksT�O�F{��*:��M�b�(�T��owӻ�k#|��)3(�)���܃
�LF�[�B�s��`S+��<J�o�=7�Q�DFG���J��йOOd٫�x"Ԯ]�qZq-�����b���)�e9?�/����fɒq���j���o��H��"@������=��_Uw�l�Lb��1\I�w"�]�˰�f̬��jq����dW����Ī���:��/Y�}�JoM��*%B�x"�IU�� ��5і~�v'��Jb�㯏C]�}���bZ�3�g�3�&]4��
�,y� 5�:����38k^����|F�v�X#�\�PMB��]�x4�C��M,,�a�~��Pp�u|�fҞC�d����>�hv9�k��zI=� �_��g�c�,�x3�R��4l��bs� ��B�A|��R�˜��`C �K=Iv�����U��x�Bf�B���ڭe�:A�,�׬q��ڲY�ı�>)��8��ZbnQ��W�+�x�h�E�5�pH�\Â�b�U�@�f�R�ϐi;Д��f<<�G��?k<���)����m&�+��7�#P��xd��m9D���Q~�М�ba����C�Q�0t��&�`?9�:�*��� �B�<��Ap����^r�c��Q��'�����е5h �=ycD\E��Z�t�i�9�EX�Jg𙱗>�9�e�7��JG�o��G��������%��;�eQ��k��jJ� Va(e�d����r�H`e^�[��"�{����2�?Ô�<�WQyHX.�?#��a敁�v��ϴ�lp����:������ �ҊxƄɍ.`N�f"�C*KA�����Ɓ&=Kٿ	��,���+-㧆pЌ��cW�p�Ao E�����fH��d@c��~ˑl�( �G���Ia�����Ů^��w|�m�0��L!����.�)��W@m$w�l� ��+Q/}�.�h��i�-De�������m�0���q6�s��vQ����7=�ϧ���pd��&q�Ul���������gBGͪ���n;��n)��V��Q�3�a�.p�f+<���+�\Y׮���J�RtS��֓*�~���k�ō�����αP-g��Jt��P8>���P1��������+W@���L�>����C� �.�J%q���.���2;.&�&h�s��Z�r��X<Ҟ�Jd�w$i���q�Yq�� _=��O�4M#NV����'3�U��	��
NӸ@VT̙p- w��%E?q)�V �B�#�]��R<"�`���ZO�O�ID�B�o�A��ݏܗ��(�0=�:W0�ȩڀ����6�"P�*������d��W�Y�f$��,em��(2�*x����\���)b����^N"�V+�� q�?�nM�O��Gg�'�@�"�YDr}��J�&Lܯb@���GA��	��8d�>?3��p����i�'r�)7L�Y��f�|?J����~R9PHc��ߒ\�᥷�����u3X[�97���w����r?�$Ϯ�A� 1�<r�'za�!	@@�yt�$��p��@� 
!7�x���k����@�*y8��DZ�E�l����0f���˖��L���@���I�V�O�`7첚 C5�0�~�j"p��0��r\R_���(@B�X_A������r�|;�i7�t�0I��j��P�qH����g�PZK���Y��`g"g��\�keL�&b�A�>[�J��av�8��P=��-�G�$@��Ɓ�t���\�wB�g�e��Di}��<�ϲ���m2�DZb���#�<o�����v!�<ξd�`��C���H]؉g���Xp,�]Qu33��3p�2x�G��mB�B�<��Աi�"V��a_�&�2�I)I|�/�zr�Е�W´/I�:��Y��~f��/�j���JdW6��V�_�< lS�e[�ސ�{fЭG�f���'��v�o�h��g���ԹQҌ��S��8���~{p���o���B�%~O���ɎK�sJ�rڨb	S�K����!��21���BU��`�D��^F`xE��^͇��'F���L��_����G������sڂ�%��m�G4Bj�����%.8E���!��R:��/V`�;͖�Fy���QH�l�_w�f���fZ2@��S�'��{�wx_N��v�k%���W�D���^[5]�9�M��@��l�S>��	js����
fp8_��:�����׻����h��(4���@��2O��wKb��-�/W���
]���i�JPB��M���GSwSj�^��*������md�e�c�J0��"W��2�uA0
��������[�<����,�f� �,��me�ݖ����S���Q1�Nxc��V"���+ϰ2�Հ�am@� gn�
FՁ��}�l[����߆�A�o!�܄k�<A½J��X�U7|\�Qm�h+qD٫r��s2_��� DwWi�ڟ���k1�5>�����B_K�����?�c�F7��G�[���E�$w1A��O�˞W�=��Bf�d��+��;]��l���ɭI��%��i�Gκ^>�@�J��,g��W�+��!I�CT��;�����BB4��/�3Q��)��E������fr���I�M�C�ӱ<���Lv�c�� �	��;�(d�I2��]�F����^Z�զ���iᏇ(L���ޏz?I!�0ɛ��OO��)?�oR;�ه���/_h��;�R���,����tp	�G���������eyMI��{���v�3�K�����&{U�H-�(mЭ�r�Ok�a5e#vD�����B�z���ӳ�%�p���

�{�f��y�a�~[���!8vE0�˛�Bs�rC�O��3)����$H�nQ��5��n�;����羷(
j��0e^ڼ��I�o�Q,����ap�w��H+b����z<t-w$��t�*� ����4�p��f�A�ߦo��O��XF�o��s��ea�I6'�P��p�iכ�U:��nh^����l쀇(z�䘹�0�,��y�g@[\"�3�F3�@������㺞Zک��9z=!����`�0/ �Ac!��3��� �O�'r���I�ä�����>�˔�u�q�������Ԃ��.]R��5����G�RP����j��v��?�V>�]0�-����3�E�q(�����4�{��r��i:��(�Ե�M��p���j6w3z�I|n׉z�2u���N���I�G�V��,`��7�ʸ��{'�ǿ�1���:v�
h�������Ⱥ%�p��/�F�A�x���s�33r	DfS�'�	�"I��[����%ř��bf՘���Y "�4dA���4�><�I&�
�R���6��2��Ƕ�W�Ʀ�6R�9���R���/�5��'|��N(8iP��k��ï�@����7�i��A^����KE�_�x;�I��pUo�6�#v�8%��u�����H��@p���M�_4�����L�N�1V�ɣ^�1�%��W�s���x��f���~�x�����p�yb�]:��q�E�V>���Q�;_4\�A`�b{�ν�u^�F0�{gA�=T��>�'J22W�e�n��uj�ջQ���I�����Hd���Ui�͂I�VKZ�n�V���r*?�م��	~&WG�} 1��p�b�o������؅��;v�&f���?��!�t����b%�>�-��@��*�`G�O�%�w������گ�>z�B���r�:���`����ڄw;��vz;�h��o:J_l�B0W_��ֶ�i���S�r�/»�&�'�/�0EL!1��XD��(ڏ��>_eS�2ѶmAl���\O�^��v���6��Ҟ�P���-������I^�v������^���D$�7�wr�-�,Q�r�W*	֤7�?��;�����ҝs$�z����ӼUn�(Ճ ���+�n�q���(��Ä�P��ꭰQr	nʇ���5�����Zӝ�H2ѭ�&%�O����_�9H�A�@� �6��c�6nvj����/��-����v�r���Nc�%F�G yt�!�}��g�(�o+-�5J��[��ﵿ&��Μ��&3B��W���W�@��4��V����������{ṓHto� �k�0G
�^����n����א�X��&:��;���M�;�{?H8,���D�/O]b�g����A�P�b빂0f+�]^��7G���<�X�#J	������T�PC=L�Y@�_�@KH��.���y�ظH�\�xZ`CS�oV���x^����ϸ�	.wB�0o���'EL��ω:+��I�,<^W#�&��f��r�I�c�!Q��r�`���nx�+���n����=���WN�6-�O׼����y�ziAlvPh�
��Ь��^�x�	Zh\F�l���R��R5�/�`��-f�b��������q� �2�8Z�d�����o/�6��K�T�&j��A����Mx��m�+�m�;�zy��}j	��ٚPS����]�`���ѰPڼQ���>`�(V�� UVhX?uw^3�s�?&`�Y�6_����%$�Ky� Z�)����/�L���Z�ظh,�+���Q���k�_\fb���d����a��
y�V!F}��%��c��sC��^\��0�[�����0QS�w 
����N����,�ö��	'	�)�T�P�A~Vb. 4��a�o��ZEH{X���<�L�N�i������C=q�8�����O��(X����ݡ�h?��Ʒ�)�-�FG�9������^Fb�.��|p���p�H��}���e'j�0���#�[s�;��Z0�V�� <	��� A͌�\^j��F1s�3��ט���F5��T
��2f�.���؈���a$Odwe^E0	�<1� ko )ݱP۰�ɀ�������;4�����]W�@ہ'	j)�+��-�e�=[�+��	��O4��qs!���Yê$���֘ d��ieA-Gw�g`��|?	Rډ�)���_���!�O?o>h�DHAء�{AJ�T�'$a¢������������X��� �nWI����r1���
��ȽI��@�WT5�b�:�Z���Np�p��zC�� %³Gq���鎞���Dq�	b� �17�@5
��H��R�h�d�]Ό~`A�ɥ!&��/wq�`HvK()��5���'�lT��x[*�s��.��Hx�-K�1�o�t�	�vt�X�/���rbVL��	�#e���ݽ.@Nfm��%����k�����g��M�]�Y�T�����7Z`;-�	�n��i�cK/	cF��S�+):�"K�����R��Ū�!^���5����6@��n���f0�Thh3�TOl�+�lQ;��s9���G��Sq�`��e��>YC<"���q��<QP�)(���%�X���^j���&?�?&��Ű^A�������K1�|Ĥt9
� ������y4LX'2@v��)��V��)�ra�����'d�/�G2+T�`-n
M)�	�����t�����]d|`T�Io�髨�	� ��pb7��
G����%0q�D�z6'~"	p��&@
���<��,�d�M\�]h�I��E;Y=$j,BՁFW��>O`�b�3pb��6�4���n�	�y2L)�I*��6Q��8�[��)�2H���ѢR*�B[���!�������~ �KoJ^�	G[#,~5>Ch�d�+<�y4�5��a-�pJ�&E�.�~�.V�L��l_,>)�> �'-�3zl����I���n���`�Z1�^P��I�ORh'%F�EX�E�@/!p�\��H+A�~5a��Oa�
�+A S�ilZ���߾�|-�`h�~p,����ʿ �A�������#��$6ש��$�Nj��ǣ[�W�}%�<P+�7
�"�ժoO��� D	ke)��&3��錠� {���kT�P���
߼^�T!ڐ�/�x�^��H[��5�(ᢔ['[��P� ��(�X��0��Q��*��'�2������1��1�iM��PT���I�M�� ,�	i��� �ohn��wn`�h(��`0�?&���FX�,%br? ;l��!�����������Y��"ɟ�5�bN�t�^Np��g�/�?����6"�:����w)`�ъ	`^�AQ��\m���K����3����)ۨ���,�_<W"�/���eV�U`^��7�'�jC���L~�:�_h� �a�͋��WO�Bsb#Z�0DÕ��g D��~��� %l21�5�+��@����)A娠��k2�[@�)���Z {�1�h;[m0]�@��*�UY��g�,�E��9���灐?�` +\��-����؏J���z�!�kN8�͛mXa{�O[�Ì"�}Z�C7�	���&;�{��*�O
&��(`cB9��hS"�Ŷ �4(n�1�\���A������P� ��&?e��S�/`��5�U8z$i<�������ְ�D��5�0�q�*0���U?4}�{�Ai�~*�� �ؖ���NN�I�[Ԥ�Y�hv�S䨖�1��3e��К�T�|�9��,��)��%�ځ�f6(pXqQ��?'9����(Ͽ��#���=��(&��P4� '/"r�䗙6a�C0 ��e�lX�т����:��9�m�
Z�����YQ~�h#<��I� ,3QZh�[U"���K P��d0i��	�}� u1+�*�~".�;�1�4�0��c,�G �t_��R�@�h!�V |^%�A�]K�[�:(-����.�BӘ���3Mza�,�]dC0Vƀ�l����=�gfQ�)0��Y�!K��T�k�)�^&��\�㠝%nI�u�"me�5��=_ː��R� �k���DzQ_1��9U�yX�k<�_�� �^I�>�|E�z ��Dw_)O� �U�n<&m	�M�"��Z|'�b�GM{�����xP1~�./�Z�g�H�ڝ���0��
��(�Q~���3�\���x��P)�ib���j�� [����%���R��K�.�|�ph�La��o�`��Z�I�.1�D$�� :	-��=(��@��/m���8y��^)ÂJ�l'}���j-TYG'j7 MI�U�~O°�x�&�[fP@�-Q���^A��/S��pb`H�!�����hDKE�Ȯ�-:]T�|Y �G�P%4t�jH�y�Ё
�?�ȸ��R%Y��[�~q��0�ZR�2�հn�0�8�P5.2>-E�	S�����P('1^冻 Ɗ6CNޠ�� 
5&\�r�8��)�!���dZ�{�hBV�X�!�G^�l �,�|f�b�@��Oܩx;8�w �S�(�Im,u�2?<x'�
����������xA� J0�0�:4�[�ݤ�0�v��fHB^R^�xJ�v�8�J��	��T�Z�*�>\Ex���9�`F=o�{e��S��iz]��1K:3v��9}	٦8�e
�*�(�� �Q��ze��(-�(�)��V	�f,ON��<.��%H@B�!d%Nr���0��B� ȵN|'�>|�[-BY|��[�ky�Aa&?ig�+���,���m��q������9�$�40]�N	������Ϣ &��^	1�I ��S7�Ѹ	�X�Rp?^@��0�!�ܽ{�c51n�Kp�|ӊ�=��P��@��x�E��#���A��P+("���}�<��q/��l1/{(�j�8,2�f������ ���ҹ{)s���/?��Bp	�v(�E�|#��R�����Y��DH�=�B����_UKv���r/�] ڤ!��>�|����a����x�V�B�� ���� QVY^��O�R�+�D���oZ���R2�U�v�� �X�h�YY �V2W \��3���ʏS�\ _�[�����#%&�h��	Ԫ NR�FS�bQ�{�U� �o�6X�3:>���,d�x[S���*>e@�3u���U]H��P@*�%��<��7)�b�_�3�A�.����9�[PpR	��i����;����0��=�PZ�~ԫ1w�{�YS,�Fo�j~wͼ�L�H�-&������RgC �L:�c�J|p�4�1/�)ýSz6JV�[N �f@�8���y
ۗh1܀X)JT���}�Z�tk0h�a�?(��]TƉ�㐡WeNR�>a���/0��#���-O!K�@>��|���΂܊(qV�\��ͅLh'�>��ܼ�UגN��s*�^ް�1�5�.Z-xO�!Ў�Bv(h���L�J�5'[�X��5(]5qƊ �
���2�6|T����S��G�[�(�h"�;�@ML�� Ȯ
�Y������%m���C�|���L�%�$X�w5�S�)�!�_"�:5�:#���aZ�	.:����v��� ��&��U	/� C�� �q4޸��t�?C����$w�J���}U )�錟�h
��rtJ9�*RL�L�:�Z`���KI��B����Ņ
�p�R�]&f��\�`�J�� SWh>MiD_���y��Y�kS�2�~$[���_��'�e/�%�@�2"�`T�G/��Р �ݷE���`t���� h�	�D逹������
y�<��8@C}�(�F
�B!ڬ�ht>�=�b����K�V�*+�R�-gk4t��\	����	��F������GkH�7Cv��9��*��I	�U������Z���!����L�K����$ `)ѸEGP]�n�kڥ-s���q�k��y��=��η��ީ����'�Y,z0/��&(W��2#J�I���v�x\��%�d�Z �<�\8oH�@�(SXꗚ�޾A�9v�G���gG�a��huZh�.v�dúU��=���6Y�IX�ݺ�@�[�Ǹ(s==0�5�GA'�`��p�V�*�a��)ӝ�Ih�t�9��H��&Z�/q�i�z�[��@�^�X`�N\h�D�W*��	�/	�3�82�,��Y��J�I��|Ha��AY�k;Nu��2{^��[�X��du�ǹ�h�%)���k`U��1ت�hQ���2)��Y"�<|� 8��\���SR�u��(�Wa����[�Pˬю.���H`{v�i�10K��즔�	ּ�w�vY�����`�X,I)��_jр�6�{��O���>�G�U��ӹ�	I�.�A�$��	��h)�Y
�nXP�;�5�=h
hP�o!�*����`�hdJ�&/f�	�wC
R�§�A����{�B%�W�����_ء�Ą1) ��uq�p�.-����Y�P@�v��>�dLyZ����&�7�k!J袳N���sLh&�R�9P�c���D@��k[L ��p�J��ݴ�Zݘ�5P���z�2�����)���>�#���a��b�Q�!�B1wf�����]/Í뭻$v��C';h%� ��o�f�:j1��pH�r��vU���g����`n����<�t�Pi���J�2P:�c_��G�@���xY�n�m��(v���Հ�~}�S������y�[5?�DP��1e]
�%�iX��Ee<X�%(Y�AY9�p�a>�h
B<5�p��<�G)ؽ�	K�qE��wo6�@J��wV�/�j*A�E@h�2�>a��G��`l�8<^G?虠��`5��v��w-qF�\T�S`V)�` �/"<g�?�/�$鶰�"@v5�o��"�	ר��rZ�C{�ͼ'�st��w	ݐ��O��)'�^��P���É�Q�`�	�-���{t��i��q�.R�N�ZF��@p8S�u^x� 4��"!ʽ%U�]dh	�+�)��5� ���PI��u�%,#����*�r���0�y�;H�XO"P�E�b# �[	Yh�g�SQ9��?��<�[��(�-�f9O�����kͰK��L%|��� (O�)��*��9�� r�GHR-^�5��y�n��zi���S�%X^GN��*�*(�q�9dWR��@��#l^F�Rt�-�l��_�)�����p	�O׌��(��������ݬB�w +�dPFZb�,$���@���ї� ��#���#��A��&;�e�p�T0��%+v���x2��\���+м�	�ai��:p�Y�FDx@���-1��� <�����qH��� iv��uԈ�\ �;�P[��P7�]�{o�s� �CW���h�r�fH��1����$^y �gBHX�Q�)�]�g�FCb�v�� 
Uօ7f8r�T`>|d��V_Qm
n����s�R���4���X	AY��-�z��@1O�	�U��Ff%:%D��G��k�� �3��0�f[.�.U,�(���Á�.�&X`t2�Q�<��X"'�'�D��7S�2��ԑ���x�l/	}0�q�����	�5E� X-�O85���!=�;��	�E?�� .�2Z�ى�����i����b�VG}�d	�UP	~a�_E�;(�)��Ծ^	�dpX�p���fRe �j��g��Ll�B� f���.^FZ�>W�/7�Z\�04Df��d�v<Kʼ%%��'�z�8���"p��wW~�j�^���Z�� �pݧB�ULT:�@X��� �ln�W�{	7���wbev��k4	Z�E�@#h�~� 1��ހ��=�*�1�^)��5v�T�S�&�I�ueF%I�ҧ'~�֛�'~�P�N��S�Y�ݗ?�	X�=,S}+�&c��r���	*[Y�aO�%U!�]�ED�j�׸��XS�L�Y ��~��	1^�4��K$��Ņ��\��	����X��P��X��8�;���(;I`K�<)��KԬ ��A^����ì�)�Y��U����1�B������p�T�N��D�hS��<=D�Dy+�dK��"���a3�fY�!�6�h��uՄ;���ĂRVPl�H��s.Zh�6q��h�X_E9;Nv��1�0��Z��p0# �?�Q�rN�T�2��
;*�M���j&�I)�Y��(��R��� �Z ��w�Sp(6� �������Z���|V��]�����}����̥k�0/'Z�	�����=���A@6�i-�J{oT��>����A�-<��2PZ���* �5|�3)��b?1 *Z[�zp�MK��������W?�O�9�Pe�c���� ��k����7���7���k�I���'?T@�B��p��X���~�!���8��08VW���X��,0�S���vL�H��!������8T6A��`�h-�0��8�r� ����u�)��kK��fK�Y��ޘ�[򢅔`!�1���ky�\�	dP!�Bn����F�$������)�Z�� �>l�u��M�z���h�H� �a�G�6�,��9���E��'m:
�Z�U��P_V�8'�j�,A�݁�w|��Jy��,)�c�r:D���~F���,�iҘ��WH�b�h�2��]�') ��X��F-�`�8
��?(���	�.6iy��* ����Dy�]xm���5>D/	B郬 컇qO\s�:ā��1߉�`?⽂��;HV�f�� �m%��P�xI��pN�z#q;��!�W���])�	G�4$�_e��b@\^h%Zd�q��
2y�1�<<�%k�fJ��	!��g����Ky)G0���x�f0n [Lc;��0SP^��j$}/e�)X,�o��P�*\�	��z ��'�G�C
�� xM�d#����ٍ����wfh�}�E���������3\ؘo�J����3Eqt��4[20h�0^r�p0�·�$^IQMt#�K�P��#8��>�Z����zv<��=2)� ǇJ_hO�r��E�P��8�0R��J�Z
��o�D
�iN<_Oz͞`��8H8�� �X��k�`5��U&xOE����!q91���)L��K�* �+.�J�v�x�3��hRP�m]n�jn���A�~ |���YL'������@��Y�-O�W�B�M �`^�)�,�h,uc�j=�i�R*|s�Z'��&b�t��W��>�f ��8�J�g��H:��U�N��
&���%�0I׹K&���8[@;�Q �3g3�j��5����`*R��	�Z4�NLB9C;n���X{������Uh	�B3��[A�����i�XO5�^	31�p��h&�(H�Gap��Q��Ӱ�v���!uȲ$Z� h.n��9-�cD�Ҋ�w@h�Q*��~��&�N&_��w�W&�8�k�_�T]ņ�h�j�I6��ngj��i�(�L��^��Y���z0k��-�+����R85LwS^���%��Y��`��[ h�Mx{_\���[�5�,���NEPa��J�)����Cd�v�i��-��!˭ֆ�IZ�<S��o�y�A%Q4�*ϙ�{4�'���ǀ����(>��ŕ#�*��b2/^A�)X%�烱U 4Y������������� �h�YvK.9w�g�5�>C\P�@�8�cC�����0��������IU�?6�L/��{��31�\�p�yE b���sX���a=Cׄ����nݲ,5[dZ���D(�S)� �g���Q^Z@2�
�JX	�x}� Q�!3�~��̺	w�	m��-\�gz�=�lQC�@	e�	�qр��=�_U�s�t�m�f�L$H�*�m�$)�P-Z�a��~Q��!����94�	�v�"�	��6�yydA��"�H1�KЖ'�O��NQ31i�"�X���J�]h} ZS�>6�nA��NMQMn��[Y}�'\[S��8�Q�9�K��_��X�M.-t�a�u�3@J��q2 �/�"Q�	��Q��2%N�#Z�J���P�-[��^�&A�p	��o`�-�`C|xF0�JL�#���$�)�-� �G�4P��� ��
�o��%�����>~$�Й$:�(�(�����l����\��_�H�b7�D���hDl`NŁ�f'�p^�d[�'[�>	<{Pɀ�ҟ`
�l��`��)ى˽2$��\� ��~\)r��0!�%V����0J)�`i�xo&��}E	�˖�i�P]*�����,U�+G)��`���֝SHy��PW����_��%������H����������1Sf��p�b���*uC�׷5����3���k��K�ވ(М-�Fw����P鰕J����R��N�낕� ő{����C���i%$+
��� ��3?q(�R�z��MN���/�V �C�D�^���*3H~jk�x���r`]�a-����?�.N�N=*H9��ʢݍ%x��l�eX�g@�@��p�Lk^pxiv�8�"0	�����`'r
���6{���J�,��-�TdD��À<0��-3`�P�9�Q�ſ�7+� YZfh:�`��<��(̀�j ��kH���y�+���Z&�Y�kb�A�!xj���%�!`��gh�.���` �e�U}�s�'��\-h=HҠ�h�KY� �ǚhEց��.B�_wOhvTz%���#)���(��h'�@�G�K2�@��^�ԛ X��1�r)��Q����W��~n�����Y���g;�AC��q	��
s>�Z����7jĜ�. �_����(t��(}��Z(��?@�5l�7N���e-�C�k ?��va�el$��E�Q��6�W�@)�_�:�m��#�"�JL��ޥ�L����-�B�:��ĒV�&�c���!�����ZV�H��;� �.�?��O,}���Ne��{`3aLo�$����)	�h�!�9�<�U���͉����� �.b)ڽ�f��A�TѸ���r��n�	g}� Ļ�FT>��:$!t�Q�N4�ME�ݞX ������	������T_��-�.	�-���. �@�	���V��)�hL�iR]e����Q��4Z]E��-3�IӐ��XG'�[��4ꎽ����?l�Lh2^�x ��ؔB!�s����%ޫ��M���O����{(���bu��X�0'�[��06�fO�����?>r����9&)�tr@k&"#�x=*/��5�$Fh��1�n���2-4tr��^�I��v	�$1�GWb��������!��}&w��T�Z[x���DJ����QWx��9	+�p�,.��H�㼿8�_4S�Je��WJx����
�v�ӎu4����oC���S���	V$	\PW�T��N�ˈ��u(ņ�(�,�R��M�f�U��9�2n�"����92�s�K�чڝ��2K��ϯ��f�6��U�20ʀ�f*��'�rz��[N�L���*���fsy\�F@_���ЕN�*�1�2J��^k��#�V�`���[5���cE�e�Z�Kn��hB��55���]��yX�s��l;
>�<À�����_�	(�fPD%������1��*�!Ok���_��U�v��h�y�MQ��P����X	Y0w w��C�4�ց�h;5�`t�*c|_�T3X8�r�%�V(ZY2���9��C_�\$Aj����t3H�<W�r]�d�/��Dfr[��$1r�/X&��!q��MHO,��@Y����U[�>��v������$1��p5:Y?ʸ0�
-�%Y����O)h�@��_ $'=%!^ ��9��ٞHN�71�29��Ӵ�_���DF0��lAN� f��*��y��$ ��	,���	זB�8�~��ї9w�U{ŏ�	�S�)-�9�} �>n�x4�g���Xs��?��K톤�^ZDe��$�A�S{~��Qh�/Y`X 	�k,- �U����t$]���3n�8�J�2�[N4�@���'�P,�-^�ʹ�K��1팖@^����dOJiXi�/�<��*)�j�z�� YpE�5��(�h�=������b�@'� �V�Uu%k+�P�^�ڗH�_,d(ȑ�hc�%7���Ef��yܼ����?�_JVo�Z2U*�����NU"�4S<��@�n'-f�� ��!���SX@�=�N�a-k��ȾK �m�J��i�V �� M���f��!D�~�5��E K�pC�������YhS=��2Њo��r�1���!x1�����	<iZof�@J��Е��l�aW��h�š�Q�VD�E^�=PTڬ��A\d��3��*�w	Xhs0;
'��^:q����\�?����S����^6Ϙ�i�?�[�f�����+� �
gN�L��X�?0M6�K魲Dv](i��9��-�)j�SrWG��� ����_La��`�xYHSD�UXy���,v������lX�@
q�q���� �M�kK1��>](��J���yS�#J�E-d:�c��ֆ�D�,���!�Ŀ��1�E0��}����t1o�(� |x`�6Sh=$�;%$����0��i^##��s�P�0[h��b`K~�#�@0�<�����^�$rFL�"�h	 :K�h��,�V[� �����F���r��t["v��
#Mߵ�������zRa:'�_.�"���`պ)�y���~�`�(���M�+ k�KNXm��	1_Z`�iiV)`�%Z�����1T�R]�s`SR
ȿ	�"�l����T�Q�>�&]G'��P�b����r��ѩ�\.sI���g�)�II ��VH[��A��D
�m��ၽ��#/ī�| ����'�����@�!0h�n�HT�+f;ٽ�b!�\��S0����grEa��.3�B����UJaȖ^��xQ� �H67��hH.�`db3o���騶�]t�O�I-�
�Ȁ{�yT��_���C!h�{W,�!��";Ѻz�)�T���"��d���\�;_ȝP���;H���|a��t���B6`{�b;�x��'*;_&��r����}_R���~4���J��j	��M��piP��e)л��l��C�v#�?2u��i������Aˮ��C~�l��=��O�n72;�<h5�F2�3w�A��,���R�z#8X�[�G�\�B��15��Kt�N��b	U[Q��� �M�V1�)� ~�,��Zh�٭C����oK�fZ�h�+�a�։�1����� ���^^�=��=�׬�QS��3� ��[��(�<\���]/X��12V+�A)!x�!��t���")�'���umc!_>�B)ú
VfC6�I4[B�-��>���+fX�/�I�r '�)1Xs�u�e1�^��hu�G�E�XK[��R̀Z�x���Ƭ�5����1�ֲ�����Xh�)�E�8���}�vP��/,���BdN?�I��[��z�vzK���gi1�]`m��	��� ��5� K��+ �j�׎�T�w�6�Z��Q)x�^�"�����=�Lu_�q���Xhn�
�#��OT�2	H@5�b�?��p���j� Ɨ)�|.�`]_�[�����9`�\�n�PvU�������'���/��$6��"'E��Ybbr~GcH5һ_�}Y0Ư70W N(�<�إ���$���ݎ9���b�Z�S.Z]�y��U&�\w-�MQ����_$[[����}r�'��hHx0������Q���dU�]� ��]�\��7f�g�Ӥ�vƗƴ�{��x�j �Wt�aը�/T�ޢ�^آ�X<�K���T�𡉰Y��%D`�z��~�H g�z�+�[N�?�� Z�k�M�o�#�d(/kr鑟�Әs�Z����b�^` ��3/g���1	o5����$CB^���N��"�GX0��yJJ[�^b�����ѫkRϘ�E8 طxP��&��D�hX":��e�%���*-��r'"u�f��d��������#��h�t$�i!�\_ZT8	����Ս�px�wX�KO�-�p�K��sb;�V�^dB�!D,E^~��OE��\�n�H�{Lz.�e�;���o!��c��Q�=��!��*�n	'���b��D��ָZz>�_��2?�0%� �l�V)��XN3�*�D�ea�:4T���hTF�d@E���3;^mǉ�����}�(7��(�������`�� �X����@ֻ �+�\�6[��)��6���D�^ �r�b�@igYܾ`�Ӹk,)�]5]��# �I~=�?SЖ�AM]A��C1�`R�P���� �BQ�A�����"�~.��R��
�q�����{������(�0�P�)S�3���߀�;����h�V"Ök�U��&(MP�m�h���8�!}�YG1F*�;B���t/��v��a'j.�IV12#�9��۽p��1�.�w ���.�(��c�n2�͝�P��f\8P�)r��-��n��$_P����������^����	G/�ո Xi����m����&�8�KHIB_������q7VH�r'��|Y )9V�(,!0��1��'��I��p�Ʉ0QBB�����zT����\� �';/-�Y��;�MV�ٞ�P�n�`��Cc�j�	�W���� +��h�(Ԙ��P#6�^���})z?1���nF+���?�|�{���-�-n�t���o��%]Ll�/�T�T� Yk,ZM'�{�?2 ���qͽ�����F	p!Љ�Wܦ��d���,,�S�1�Tk�����;E���4�K�>t� �c@�f�J��)�v��W�z���XL��uN����ZU��"�Ph�*w���(�
ЏJRW[�q��� ���9 պ�[�A)�Z�O,m�p���*
��G�CX�$��2aO��u %2�J���S� A���J�U(�-}[�٨��GZ	V��>�h':$d�\]����2
�w Z�9�X1�QhU$J3+����dK-�B�YЈ���kǀ������	�0}�T����x�#��qDw­q���ٸpe}T%�Ak{������D����2�y1xq����JjԈ�hVf^+d@GX��V�, %�0����9NK`�},Q�8Lk�?�r�@�$�1���`9�=?���[(�QB�
��?��:C���]�|��d
U,*���+��h��,̂�	4Ct���b0xF��#=�-�良����I �Yo��|2�tB�|����*��Uo�D�&=M�I����p�O�G	�K����㔓�Y��䪰Ƌ�n�r�R���80�ۀ�� ��'v-^��(��h�wjtZH@����"/�a0P��5$�$�(�p嗴G�_�&���'��.��ɰ���%aQ/D�te]�/���a�7���t�6�Z	 ���%xt�8�1^��X�� [fY��k�h������e�� � �4t0x���
f�x'ö��С=��t ��~T!�Z���S��ʀ�%�T W 5�^r `p�b�k�U-������;�-��~�S�>X���ҷ���L��EN ��?����`P�+(�0Z���⺑|jG@�R�>(=7�`p'�!�:H�Ԉ����a
�X55.���w.������Cb�H�GH�.aK�1):�lDUm�6�"8>�z_�)��e�?�T
�P�0"�XGs�L�(����|e7�w�v��ZA�]�a*�a
c#h��yo[��,�4~ 8����	Hr����r�<� "/O��n$s�R�@-H(x���<����>rO��W�Z���5_6�d����X��Y�@
��h�=�ռ�rF���ŀ	��)핈�S4��R��i����s�8��hR��Ft{��4����6R��өk� A��9�ֱ)_�>)��h�j/�T&���`���`��ne�1Y��~h.�Z���f�K1���^q�-xTkRB�b���X�fN>��P�.��1������V�S��5����>O��>	��4���~��4a���}��8B��>��� BY�H:�I~���B��|�]��L8(`d����4�����o��`ݷ�=�{ja��0h��jZ�ph	VqTz x*������r?Z��ex s���ZA����aK��Sh���L��}Y霕�)ݢ�U��?��<��i8V��6�B)���0���}[��ϟx[%�X�\;7�p��"�����1j�s&h72����`�V �t�W��zN�B�|`��-t���*����[7|�ՌZ�лK�����n�w:�XxP�`@a2i5�K�{��~P:;pL��T�}l�_��F@͸�,Qc�

;j�]8/ Z����p
%��W��r0:	$Z�+�_N�d�r@o�������~�Q�~��K�1@C�/�#}I��/Wn�%,E�������B�^�2�'�0U�V�1�(�[�/�(��|ʄJ�h'�}�c�:	ms��t ;O(�-��QF%
�$	�5]��(W�(��z��!S�e����S1#�(���FH���R ��8v����
��yCG�,=��~����F�$��������� �X�dpZ(� D/#�3��h!I� ��v.�T�	s*�,^3�i�N�l�	�2iS�'��& �3Z�,�_z"Hs �U�,��V����Xq��U'���
�H��O6?*<R��8(j(Fyfb��D~��W=MG���R�t���f����{���?	�YT��m�$�>���Y��,�8���=ܘ�]?
P���/8k`)o29CWZA��xT{0�aJ 7�a:��+g$�h.�B6k��9%���RO��8,� �V�i�jg��R��|HH�)� úU%Jw@Z�d�0<��#��"[IM��r	Γ����A0~V��K1�F��*�KG~���-Tu��s�L��f)�Oh�>�F%�a� r%}_(��V���; �5�}:��9�1X_ �/y+���n3y�\�n��!*hE�\�P[V�A�j(��&�D[ـ�j~����-�x�_�������y�J-[RUf��#>O8pP��b�Zޞ�]O!�* �ZY�o����`��X��)�V �Y �Jf�)3N@;����:B�,#3V�*h�/UQ�@�B:�PnÝ_�x��B�B/�'����	tS��(�m�5���Z��	�_�XYh�t`X�.yCH,u� ��P\�PW�X�*�!!���oM��pB�ԍRVJ?�~Dr4q���e+r���K�:��n;��G ��]B?��.,���L�����![�3�������)�Ad�C�������҅<ޙ����6���&]�Z���S�dRD�5�yJ�63sI��GW>��)7͉����n˿��D�\b���Y1K�� m"�6����=!��1�S��L�1����+
`	�-������T���D�!�}� �
}�g-h k]d�t��q�X�AN+9wԐ�KG�l1�>��P��f3
�$P���چ* �JQ��!� ��]�����\[o0a �s�U5�w��$�)��Vh}s�JH��	>C��9&��]`��^��M0u�^A2��+����ڀ�K%^��ԣ�j���mVԖ�Z!��l	z3�טƥ�R�[z�gYL�
�fĂ�w��W1�)��v��)��_2��ϗ����8*�����EC���
�� �}�d >�1�)ٻF@���t�4B�����ӣ�5�
i&�vݾ��t�`QTR(����3^j�e�)���<��e>�	VIBɢ��c��YvH�n�e���kEV�/@���j( ��J�g�X�!+E���*��-�~,/d��/~��&�U���B�	0���ٜj!*�$"�$��\r��+;�#�nJQ���=�PJ9�%�v�P�p�)��U�GnZ
�5J���W�7!N!(�E8 >\%o�v�.=��@ ��i?5��@sj���Q��A'@	�K� ��E�K��Hi �G�Y�c.K����Z�A�u1���/�����Y}����羚�� �Q��~����fV�����j�5�k�d{��	�[��]2ʴ3kt-SG�%�l�C��-����6xE)i�0*���&�;�_ ����حȤ ������pn�E� ��H�W�^,�~�����0�A���]������A�3�X�J0��J�4��kR����n-�LBf	[��[�����9����+�W�l��)ლ(Ӏ�A`�R��$0�u�*.�[!�l�mB�GA�_��4�`%(�`��h-7�v�, �]�-0�2)����^�����	QP�>���H���R)��=:'n1�s�w)�C��o�Ȏx�l_h-P����n	"���v�;�h��c*�	B`b�]N��=e�U߳x�B) ɹ���(}��-,�P�;�4ޭu��0�gm#q��-:~Vu�8��/�ni⻧h�2��N]�T;���_P��!�;�6�mH&Ʌ�J�~��	GW	a��%t<D=؜o�sc���-͚��XW�Z�?�2i����W �TF�o�m��Q��j�[ӪqW�����S/�m@�T�. & W��x	I�����ԉ��ˀwH��|
 ��~�����PW<1�+�e�D�ԧ������s��^G(�@�鄂�>��LI.YȆ鑳 &��D�,'a(��1P�@@5	��	�����1%���X:?�i{�t���Q�a�� ��Ғ����ӘQ� �
�x }p��q_���k�61`����`Liҿ����g���B `#Yx-<�h�I��>�cC�r���l�dC������
VTd��8]ǩ��B��2>Tj8C�bN�.!:g���a""
?��qH0B[�  QhdNZW���J��[dV<��('�
Xh����<�`EKL(��������،O ��. c+��)��G�C�O�0��-���zeL���lꠞ� ��-��5�Oz�Pz�y�ʹ��8%�!n��!���P�O^���ƛ�P|�z��ue�%�.E�L��F4_�})�h)E政_��P`Tu�y�
�*��Q?��O�s�1%�B�7s��cɉ�P��UD_	�v���	�{�n�vc�63�Cc�����|^F0�_!e��s<)Jع���=�K��! �^��f`�r���2
ZvhN\�}���njQ�.��x�Ʉ��@X���O��¹r����*�tJ�tԨT�����\*�TO���l�!˘�h�;`@��I �1�J���	�R��@jh^֡L����Ӊ�w)�W��I9�Y��쬕���l��2���]]Y��	h4��$��xî$N�b�(�v^2w�]B�ü�?⚠�P`�u�3dIS���8g �GUo
*�4#@j���-l��=n-X�����r�$���>8	h8H�R��2�}��w [Q�>Z�.�=t
K��נ�G�~'!�Ye6�@�h���8�r�T�L����O ϸ.�Ok�Z��6�7 4�Ã��V�Z�l�0w�x��L�&�%h{�gFz����&�ػ!6b�@�����	�	w�� &T\�1�_�~��p��!��;	P�8J
O��Q��&dD�	��g])`}hE"q���vB)�p��圄h&�:,aPhd8Fs�LQ�6�L�@,O��R�~=X1ռ�5I���]�E_]��ǥͯ���<�!$�&߁�
k8ap`�	i	t  ���/0���c�}����.��[����/�$�G���-��JB��;���f]5��~!� )	��ܐāF�>����f�b��(�!���Z>�s1�H&
��f����l�3>n���g�h-�-ff��aB� �W�
��|,;�h�s�_��lAe�1�4�����h���N��B1�5S�}��[����"���0���8��_k�@���^O陲
T��@��H�Y1��B��$ hͺ�},�g[�F�n��V�/`QG��i�)��3\������[1=Ի	`g#��Qj�?��-n �p^��cr1V�~�Cջ�������y�.*G_�F��Y�b< U1�!"�A#�E	�@ ���-��V숋Q�Ȭv��-DP��%�l��_K;����-&/[B�mu �a������"�/�=�C��n6Z��q���s@���xW&;�	P�:]���A�(����[�����Pk��x@�x=��z,�?����E�@��3G�O 1�Q�f4$A�,�=�wZ���~�k��/(�I�KaԲ�IHP:��dyX����z���-,_>v�)�Չ�vw�����!u��c�<���W�	W��A.��(�ò����HO�DӰ��,IP�(_r� ���X���B��x��~ ���մ����o�1X�E!9|��[*��?>�Й�2N VoP�n���'�"rNvF �>z;Z�>�F�
�d�UD����Bt���ŋP���8��F87���]�?�n{+�(XR�N�h&)
������	؝
q,J"�f��6�ц��찅�@`X��(�`�
+0�f��K��3��Q� K�{����40
ʽ�e§>�I��":0�QS4G�ѹ�1/�6��J�X�W�fD7UR5�� ��jo��KC��`6G\7�H)�(v��Q�k�$��IX@�M&����h�0���V��ėօO�N�9�:�,��]��Ht�P���H�"	4�y���$��N�������P4�C���
0nK��h}�1�u�yV��Vo�۬�]u<\��%��%J��.@�!G(�P�hN��y���3鯲�r��VZ��[h�o�6��7;;��8��=��F�6�@�
)�P-W��V�����k���Y?�Y��(8z<Kο <�~��j�����9�՗���	���!KX��
l�43.h�!���eU%���>/5T,��Q6�9��nE)?�`>��DU�7�F��N� �f�	^�	8[h,�Y,����#����'��#�V��Ab>��]�,���j+���4M�����&�I�e�c��X �"�j	��Z��iZ`�Y�[i��uTX;�	_��{�w �ͻ�`0�+>�w����&�
Q��>�L�$���Y��#.%,)����%
�P�����V	)�Ti e�'�L�I|I�/�İ�����@�ƿNP_O`L5�r���������	G!���	�l��]:(-��F�N"> �J�H1WH��h6E�̚K%�}w����IO�U`GQX�����:�4� �1~����RCD���>���Y%P���<�W�df����wK�P?�',�I^�T�e���1z�ų�iz	$��T�Y�m�������)ߠĊ
'�2T�Ļ�0D"#�?�]�aO;�
���� K�U�`[�~��I�	��ݾ���\��Z$�Ӳ5��Q��u��O߬6�ဆ!Qa� � ~�2���:�Çn�X�3F�����ь����R���Ki�K�.N�������a�m�XUh�Gv,��:�z�C ��/�ڛ�]�$p@�ﶰzh/�R�4�ӟ�Ph�J�M��H�_�^���zl�q�f��8���w(|�V����_�QN���z�������1�+��N��f�!��$B ����9h!sbA]p����3��U[��쵤���9�d����3$\P	��C�"ߖ (���h�c�`��{p�r������f#үǿ�f��(�%��.à8J�As+^p%�;_��?[O��Xc�? <�^���,_)W����!+�`h%g@�x0����7��ΰ�^%S^`�����i��Q�6��3F�Qv��<K��7It![@\��!GeU�%���a��H��i?��<�?��SȊ�K\A�;^�����>n���r��w�q R�Nfe�2�����$p�-$ �60cdPѮZh�2��	���Yl�{!��`
Z�%h��V�o�J�.����ߘ��(w�AbF���|1��S�Ȗ���S�!�0�h�^a�@	"���eU����
��r)�@����	^`��sQu�P�v^��I��z9�� ��7�?Zw�E��z�/�| )o@��O�
�rZ�t�%u���0����\1�V�`WKOZ�XBJ�!�����Nvo9h@�3XJ
(M�P �ж�D��ϓ��Ub���P��XNE�����������(�j�_�����:�,Z�/8�b��b��l1��('��L2��9h�����s�
+�o@�`u~A� ��)�+�s3���O'�W�1b[��&`��+��s�$���G
�AO��
��j_��:ߓ^��FZ+�\�>��P�J_�n�E�U��N�p�\���,�*v)Ub��	�|��ho83Wx8�&�k��:>I`��o�/��^�՘�������PAv�Y��b�UY.@����s�%����*�W���;/�^�X�P��X�x���'V�6uyE���"�͉j��V��b!���jV��F@��h�W�p�쉐���8=
O�����^/C3ص�c��� �M=9ŜU�X�	4�V]t�If�")���h�J[��S�M�]!��BV�A�c	+�l/Yύ�0�; ���H��ib�@���	-�v N�}	��1N������p��$JAW�D���V$�2�eO��2�,�Y�0�m�O��B��+O`h�m0��
M��@�"�_\'f)�.�f<	Q@{�2��}O7!v�k���.w��r�	�*P
T�)�C�|Ws� c�B��
``.�9�0��	�t���='@�Vh#ud;�}d y{<4�a�s1�d�)�;�ڒ�\�*� 3�Nru+$�ٷ���!����}̨	�.юꖻF�)�v$1��4r�!��Q$LHO9��Y�� ��h&��;6����ӏ�1�h�#�h��_��K�b���[�9q s}_ ef�	�U�+��B��6��u���6�v�a���g���7�{'���#�P�}W�~�3�$�����\�m2N��h�n�G��_�ϯ@}��SP���)��@��r_Z��D}���.�nQ��	Z�{�u�(����Hz(l4�q�^P���X�G		���$��Qce9�>F2�T?��^�Ɖ����k���ހ�5�P(L͠�����X�t(3������	�&9~ ��1K(��u8�k�M	�	�C�G�#@	�m�:#L�]	�%�]䠐l	�L~p��nN)�<ow*�Bc�A�1�5Z*�y��rS���D Q�fuN5�~��w�hqX>�cPO�A�l;��%^�g��c��_Dg̺t;�}�w0K4k#�i���C=���3��_�[��� `g>Z�	~K},?{�P��Y�r�%���/�v(�Dz}7U�s1�u��\Hڮ�Yv
?��xۮ�t�iZ���H5Po�9�P3BZ��.O�pvM<]���:�IR�Ѐ^�$��3 A��9 �V�e[-j�o���¹w��!��5m�gk��P/�5}J�1
 X�T�(P?����o@��Y��a�%sCo�~�@�i�g	��|�b�b<��������-�����������E%�R<��H��^�O����Oؼ,��'{i(��U�Da,����8�9±)h��0��M��N4A�@���W�4�I��Q"0V�O.�@�v	R)��^��+[L1�����S��"KU��,�	%R��������X)�����a8{
-Z~_��t��U�C�H_�Ɛ\@�\�1�|{�HT^�<Ԃ�ݴ���]w���>��C��%U��S��, P]�i����=YϮH�;�1����`��6�\��t[�@a�XAJ�(�x���- R�W}��1��?3��&o�
W��EW�Ŋ�U�½�b�_�� �`�N�?T�9� �	01S����U@y�KH%�-�(걷|��p~h�X��
�T���N�
y�<ŸrZ���!����PI��0���%�jа2�t�AS����w�l�U0�F�9;�gB	K�E��Ά��MNۤ���.\F~�b�-&�V-�[��	�$@('T2��/����OY/�>zf���L�)���Ro�%a� y-Ms�;�'�}��A3�?�%nRUZ\�PUh��1]���t�f�
�@&O/T�R���8�a�(��w�h�3c ��m`�}'J�0 �Y*9��fQ�M�����τ���w��0��C[3�\�d��IM�k��}ݱ��ܭO1�`�/����)ʇ�Z�^} 3���|�/	^=�Z�G(��?�p�%)ؽjso5�x�����D	Z�e��+L�A���H��m;D���&���[	��/P ��W�.�M,� ���N�w�q�91����DȾ̰R$\HoA�]�I��
�Gxq��\#\n?s�%���-����5b���8<�
+^�f�g�����PQR�޼��G�XZ��Y�⼾�nA�S�I��\҆������j[�F� ���v�p���:��z���!ʃ�g9��>)W��_�Q; ��*�P�]��?2�PW!��u�
��������v�<���xN�B�B�^���,�4\���#�*���V��G!�ķ��ף�i�4�ht�W��#9�C�h��A�q�k��H }���^uX�vO
���Ҽ0�n���������-�m�uY�_Ryx���z�@�XH� �u@5�P[X�~X�y�N�X-^@���%���؂�1@0�D�H�p���N�[�I��u��k���	���;ͽ�=�O�od����п�,c�]��i�
��ú8�����o�zw�j-�K/��) X[�g6x�`���HN��p�L(����r  %
w��b�!YW ��Xbx��hE���o��*��dй� �~�Nf��1����F�j�?�ְ��-o\T��Yye?rX�
�,�%]	���t�h�p�ý�?��O��+�	�
D$]�N���-u;��̐Y��{I�鈭�`R���^T]��9���$	�T��.t/�=ҩu-H�6�pFJg&�bϥ�Z_S1� ��g�^�7Z!���.hOp�� ��w�O��	b�.u�)�Sz4K�R@�5vMn��9HO6��;#6`I�],�4�����0�!�:8�7M�&� �q
�{�(�5�,�+��,��e	:�� ���sZ�t���[��n���� Q���t(��p"'\�ҙg��а%�V'�_0�n�_Ь�@� [�a^�E �
g'%�"�\M����"m�T]Fz�g~�Ue��V�J��!�
a	�Ai�j 5G��+��@0\�(�5�d4�H)`h~�56���z���1�($/� ��9��U��}%@n�:^����#<`Ք�'Z����I �
J?&��<D�`��v{�Г�0�rU�|�`��Ow��h �`+X�o3`h�Vd�H+(z�%Y��ssG:���W��g�� �Y��v[���=�h�殼��?k(�fh@j�>�p�X& �Y@{@Q�5�nV�
�T�w ��Z�YR �b�)L�"����	1N�#C2(e��B�>~M��Z)����Q{�L?�5%�.V����v�%�,ӓ�1���$)�T�(����Rp��+��P��R�YX�ZS������Sꍣ����/�o��=P�-i�FH�� T\�� �Ъ1�5�P%�J^x�~��Aa�bvb����)u�CA�9A�rW�E�p]�(��%IB�v[p`����ܨV�#[�]¯W������[����4�]��r�(b����OvT��J>��'��t�F5o��2n�5D�
��i!�����A�3[��1iOW��Y�&�C�S�[��v0�آ��í}8V)��$lac-[�h'�I�<�Z�tޠ���@���@@#�3����)��z^�R<�� aQ ۉ���\�)\T���u����d��r'iG�`7 �E4j��8�r�o���j���B��ug �u�֋3�6���	�p
����I����>Ta��@�� �� 5�DN,铴\��<�b^W�.u�I��|�6.�TQ��
e��N@�Qh	z8{U� 2�s�_��	c�a�?�)�u�-D�H}�&rܝ���:�r⢻������Q��u���&�8,#0;��|L�Խ�n�y{��FJULD��zJ�N��<����W���.�%1�F`9��/���`!_X�@1$�]��BVWD�@ӹn!c[��	5FE��)�gɺ)�u��,�	���R�Q ��@�#���vQ�dq��c���b;|��`x���_8h'�kt���-ݾS7�!�y#!�9�+d��}1����;�Q>J�LnCx�w�A
�q/�X�+�"��p�̉���n�O��!����drY`��⢝�	�V&��]@�G�4����_@ ��:������)�1��$��� �r{o��R��?]Q�2!a� @� u3>RY�[��V����§�X�l��h��jW0�\A�"PN��-Y��
.J����r�q��
Z[�Uw�ѷA80���� �&�I����
��%�9Ӥ��-�O+nW���<^��Z\L��|��}���\�n��^���v7���0n>����V~V���qc�O싁�W,�n����o��c\t�+.�e ́�,_Ӵ�	 酂<SXw�����h�wb�������yK7 �t �[J���/��o��̧���Rh��%J[�" �kY2���0K��7=Lx}M��K�.���`2��Q �d?�>�4_( �V֐�q]	)�Z]���fh�N�A������ |�N[0�h����'z�Z�J0��[�����K�[��/�p0p��(`�*5�DEC�tAKf��ƏZuѽ�*�J@�x�v-T[���4&y�$GfY����
�"�X��-��!�x�k̇���ɼ�8QT�%	ER�r�;����q1J�G�A���NIZ;�L�v�F� *�@�1`�:kh�oS¯�kT�@�M1^�e��y v2����0�v��P��4	�,����K��w0�cm�`H�%ۧÐK]�h��- ��@$��`e�EaX�C�".a���RGqms1�h[-�pF�qp<��7��#	��n�����=?-������N��y�%�"WۡI��K3���`��Z�~�mi�+�m	5y���f'�-/�����W�n���w������ {�@	�	���IY�����ydaӮ}%R�(W����k��_�αo?u�׹�LNX���ZػE���z�w�)C0 �\�z�&k����T��Z��]��|g�
�$�_`Z"���Ng���+���L���1ݧX`-�>J�VD�1w#��R��W�����`C�1���."D��p�� S�X.��I�D��k)
1�_�Z�9�?sB}D@JY�o1'����)܃��0Q>h�>yK5PP�1��^�ֺ�^RqZR��I��L�S�s���P�/�2�C(����ؖ�i�������X���h@J�f4(�cӊ��8X��{���aP�~#)\ �.�5�MZ!�WW�[OR�@��
\��:b����¹`
�g�R�1h%>1�Aso�HKr��0��	Y\�����wO����L�	�]�j'V��(0 GF|JQ��1)Y��X�1�!�Y��P��Q�[��~ /�p��}��P	��1���� �)���D�lL1���/��N��L��P./H��ϊ'אޗF0��r@%R|�7� ����!�����ۿ���_#7Շ i)F)\���Mb~�`�]!<=@��_p��q!�ɷ,��<�Г�i7|@V0�-LY 㙋@�@�p?$~4�Xq�sz���wi<��Y�ǽ�%��c��ܷyVɼ	=�^8�Z+E�Q��;W-T_>�S��	8��}��鬠	0\���]�ŭ���[H��X�5��`��(WǱP0��{���s��`��[u�a����k�V`V���}�>���B �DH��(V�J
wnó�zXZ6	`���>����G'n_j�ƠZ�0�`�\%�C����.�Qe!�`%�I�鳰'({��0��K��v��	ň��H(�SZ��K]J}K����Rf�y@�HL�v6	zb-4xA���:���ȓ��0$8�qZ�R�)�w<�����C`�9�;:)Q� 鶈�]�`�6�VO�{��3���R�`�� � ��0�$ h!>XH��Z���V:� z��y%���)]:�p�u%!�|{h�lԍ�/7^Ն�	���~���QC�?(׸�~-<5\_$�<�YW��`>@�)�㟉P��L��'�.�7��-__ܐ��	��]�	�( ��� �1�ͱ�`-�N�E�&�j�5��S�-y,b��w4"�Q�&�\���E�KUe�-^6��[��mF�k�����(�������M�k*Gt��f�Kf�ٱ������Bp�[%#}�ݓ�-	��<H��PF�*�	�OP�dt�s�.m�X�,�U�SOi�"��p��>yc5�e�ꄛ��~��ZS�����7^���	�JHuޡ5Dp^��pX�
��zʔ��ac3�*��K�T
p�0�1����o�4�'@��{l=��⁺A/<j@����L��`_.�`�d�
�^�|2��,���1Ԧ�mq��$�^&�^1��+�	~u��ih�d���*(�1���D.)�ġtz�=�!nG��p��nf��f���RTZ�Ո�)v�@3��;L4dO�,~�JF"�U�I�� ����B7J���sL��hǭ���v��H>�b�Q��NE�c1Ր�	�.0X!�$r�D��1/���]�)j0��bx�1��c_*�h	���l�R[v
Sa����f.�r�SDXRU��Gj|�g	Tp!:�v;s>^2Ev`|9n0�c?�
�u��$K��}�P:�?!��.�������iA�g��Av�\�.0��-�O5��3NI�����BAx�ִK0�0Fb�>_����U_�C�w@�x����f"[Gp}�qL��$X!	��nĵvy�w]^ò���y]�j;�WJ�`���h]}�gYE��^qj��G�����*h���<��[tק R��f\!�	$����)�����
}�<-�3��S��Y� �� �ӊ[{Z{��br�W��kCנo�?'�x	����J	��e�d���a���S�9&ρH@-4�>�rX�Ǯ���;�ʶ'��b����7���u�؃�	�)�^�K'��l�u�~�)2#$�sZ�����ц��;�l?������D��g���>�Q��(f%�(���(�,sy�y� �X��J��+�:����
םt~W3c1��Y!�(A�/OR#�J]�]����L�&X�930I �7@~��I��� �����h�H��T|簸.w�Rh4%��0�3��!OӓZ�����]�@
�&�/c07n��C*U?�0\|��G��ʐ����I��B��0Y�@p)��V1$�E�OL�G�`��l=�%�x��b�䆼F8���E�6��$�y�r������_z����J<�@�&�FW�
�V/�	��	�~�-��I���m�&�N
 j�UF2%nok�׆�$��{�ĝT*x�V_��w8�u���ݸ��oH1�7zԱ �P�A24�\(kyB�/��(Ӱ�/�Z���v������]�3���[w���kȥ��<� �U{Z�p/�M��d��`_-{0�8�\�X�?7`����.H_d@��6o�O���!,+��?�\hka�Y]E�>�0�������'[�P�1 >�����1	�s���ŋ��'�Z��~Ow葰�-��SR������+��'�Zϝ�W�^�F- �~�v5��oq�dr�@��hRN%�l�)����$�6X�zu.`�@���ࡏ
�gN8�1��i%S��	.1��u��F5	�n��#6��BX*U�.���?9vOs�h�{����_�z����N�|Q�0٩���%�	��8m�L��sUA_O���. �����{�f�j?:'��U5��!��.���9]����P�}%�z��S&J �Xj:��9�!�]�a��@ 0���4�C~}1oHtR�� ��4��0����`;�Z$e�PY�W�
_䴐Zrn�7���d��<�vJ����Q5P��T�b�a�p� z���\�H�[���1��,�Wh�u��F�i�n��LK3!o�qU��&/���N�����7Q6��
�f:�)�������^�.	��!F�
=�����W�R;GD/)�ှU8\+��~lZ��/��)�U']_�P�`�a�:�U�-t&����!;�� V��$xf�D��miHtU�^���-#�3P��S��s�9W��=�_\!x S�Z4�n锔�	����R�� ZfP�"�ꢈ� �ܫ��#�:B����+�=�?���joc��À������
��[����a!_$(��|�,	����z[�X��"\$I:�R [�{b�-�� �w='�%+�fj0�]/D	��P8Ah�eW���u1઄)���hp�^�X�yO��@�/[b"{4l?6�:(Y����xuK�[��O���[����JԤ���o�$`��U]��|zW�DEP2')Lf%��w�����?&�v�>���`�>��(��4�<�q���_�A|
Q�L�)����Љ]�ڳ Xp�v1�A�K�OFl�Nj�`��(;O �C��y�.�K�%���:��� ��[�� <g��a�ڻ��)Ε��x}�p�`�T^jh/���Z��|���V��- #4_&���*i� ��#�%���q�
��V'8 	�5�B})w��.�9	2w o��ש}�2Ŕ�U�V�J�`C���ʀ�
�z�,q��-�K�U�C�-�*g|�X36*1�|��;Ӛ��z� ��n����DـL���ǀ�G}G�(�%��>9L�) ��BE1T�p�:�4��:�LgA�e�տ��
*�'"���D��/��i�Bz ��#Nr��������8&Y~�Tt�K<��!co����r��]5�1��X���;Y[�/�����ҥ݉ ��.���y��#'2�u��=�M�o{���5@�d�h�S�1Z�M8��o?*�WX-_�7�gPf%2ґ��K�]��b�θ���-��� :�p��5�as�)��g��X��*��v�%�[�e{B4o���+;�.��=��ђ�D~Z/��
R鐻� h|A�_^N�ޯ �x-f�L��~)�5CX��b@:����Z�	�{�{��E���:�Z�`��)]K�W_o�!���LQ8[	Y��	�*��_䩄d<�>2M7��L�6Xrh�)7���L��]A`�h^�����դ�j_X�f��aUs0{p'_iЈP{	�1i �!�?)��'��PA0j��hK�>�����4���R;\sl��@� �Q��te��C�Ӣ��	[�Bu�v(��m&SVIiS��hh3\C�<��7В'�r�����E�>�%\�*����Hl*�[�k ��8���W͘�ֽ�k#p[�jE��C��H7��_�s[S���[�����;��x���p�˸��][�D�����*  ��Mb<��HӠ�!�,1ҧ �Ė)���?M	s��| ���Y�h�o1���h)R,bKBa��{���[.d�#@�/I� ��hvV��Uq�I�9�3o�)u��1�kV󩟊R��-/);�^��Be~��k�E)��LW�TF%��K�6�}o�hF2�[q�XB�pN.�z`Po5���LZ��v�1fY��6��/0�{ZS���a͉(� �)bK	���r�p�d%���>	`��2��_��`�\�_}�(�H�H'����tD������Ⓟ�_�(��b3�U�&�s?=��_��+5sW1�V�����9�	�}�-b�UNi�IH�er/�e��j&:�j,		�e/��������k}Q��(�H��(SY��b ����1&��Hx���F
)� IaWV���PW�v�cA��_��-d3�uXa}G��u=M���gm,��	�5N Eq8�h`M�R4������Y1���V ��l���0[�V�&!�
�7T`6F�C���ʖ�5o�^J# ��s*A��Z�iUX�I8��O^o�h{��`�����X$�|Wy��R��P�;�Yn�?Z�H �s�/�v6(W���1�_�O{	���Ɓ��;Zn��	�,�m�ц *{���������X�vP!��\[�_��PS�9������L���H��<1
�*rO�-B�ʝ�0RҽB>���Y��cn H�-+�r����1��_�Sx�G,���C������OD�tp�MF_�M� �V��;�j	zV�?�@���G�-�%vC�"(j��� >�U)�����70%�N�������-:�uO�ߟ�(����V�Si0B���������n�N�E���[��{�-_�^�)�1���Wh;F�.Z`�S�p".BH�[��0/a7��$ɦ]��Q��%}����mH �侉�5:uj�D�� D�Z������^����=�B�B�Th 	�iU�2	���i����k�K��*�����w��P`[�8�~���Z��yW�x� w�y��������Zh?�X��{9)�<h�/��Ǵ�Y��*���f��3�>���,ӽ	�=3F|	@�l��:@����S`&�|�/U��.�<�T5\V��D���}|-�T�b;� �n��߉O�"Tg
�oC%cfB�t���<]�vN�-�(+����`Y��+�φP�icԨ/\!t��_��s^�ؼ����!��Ip��Du����9N���GD��h vA�:�Q���%�zH�B=gm�X �0�(�f�����z�OM�TE�T� �f�B1��܌l�z��T��-��ۙ[()��|w�ň�Ph�&�WY��nQ7g��H|���h�#�s��yY���(+U��A*l8/��q	�	�L}�QW��g?���5�j���{P�rm�@
&�Y�/��O�(�Y��'y���؛B�XWHx�,j�^u�:��I+�=�EAy�<�J�p�t�0���\qǳ.�H��!kujP鸍`^�J'�l��SUh�j]��%q�e�hʪ��ǽ
��IW�_�2��� RVh9D"^^
f�	��fMz	*T�_U�� �Z��hк4;	�4|��X�	z���5C�������~��T�	�2Z]�J�=;
��ʾ@/�C-jUQst J��EV�ٵz5��l��v3 �N���!���2�e�3(�~��{0�b���~����[)��H��Av�N�Ekh��tAӭ���1��o)���!��6��U	~_W����UMh����y^�@�V��1v� �� x~��������!�Ju>�!����Tqp�v��R��@ �w0�f�; �xP��̀9����Y���Q���X����	�� ӵ�:���
�����C	��joR�$���|rD�0-�>X�z
��0M�c|Z����}<�(���7�n&�P	��%wЯ �bz�e��%*i�U�ڄ��R�V^��d�"�vYI��+���#$�^�y��`d����q'��"�Y]N�	���m 
@R�ÿ��
)wXU� ��	|�3g��^G
�*�� PS��:-�(W�{�8����
4����'r��/�GY��r
Y�hC�;����=¼4�k�~�㯶4��i��O���_��	����/0]5x!y��
������8I �5v
	�ӽ	F� ^��l%�i|�G~j:)� ��A�p��d0�����������{fh�?���	��Vq!�>�mÛ�#���(_��1���ֈ�.T_���ո�v��@ZJ<0�Phk�j�:-�-Ki���+�W���I���i�K� h���q]1�ջ"'�X��gH�H��[d�������0XY�_���-xG��|��8�M���a~h48�N�h��'���t�t�J`J�zh�6I&Dr1��ǎ�����kA8�Գ ��b{^���e"�a|�z��%=R�8D_'g��j	X]h1(U#����������`
YԪXgN�J�R��u�3Q3�
Bu�	�S�j��J��ݢu6n)��Ҹ��;,��68��kd�<�!:	ɼu�_��W^�ȉW<�l�d� ��W���d]VV��*Go�JQ�$��%(3�ZT`N�J������!��
h�^�,��	�bH�9C���XP��I�B-�M�[��I];�}���9��)�v���^
��{N8<.|tV9� ֫�ZJ�1��j�2�!��d���{%ziru��,Q��[�GJ$c��� Qh�N	��]����KOiP-S�-�5�>��?Ӿ#'#R_�KYv��D�^��}�ѐY��&:�BZ��D�	����hcmXU�챗|!��^�(P��X??�����3`Fh,�E��ZO�bG�\����oF]M�Ug9Js� I�t7p���$��I%���+L X���t#4cY�6��:%w�P��/�%���G�@2�T\ɒ�O��Y�1료�I_��Mr�J�mw`�q���|�Z�7��EI%�1�y)��z������饠�`�"0����1��������W�oI�"�z��nJ!`��>�;�W��
g�{'���UL4��_������QI��o)��+�S���XRh��V��
Qt��$�/@~�Y4�F��Ag])���5�vS�bq��������t#�~XZh���YMp��lf3�$��$��2�"=,��X_R�-0)U���4�!�h�:�!������k��b/P+��o�h�@]K1��Q#��.{>h�pQ�Tք��P��-I&N6�!ؾ��?�='��h�Nb̏8�9J�[�-Ċ�h0C�I}�/�R�E��G Mt*J�g��}y�o�P�eV	*F�5���[Y��_W��fw�7(p�y�t�x�`Y �[[��x�b�m�΢6&X�gZv��-*�kX?��+��}�vDث� z)X�-�J`��{������я(q8��"0XJ�le�ԛ�U����2Q=�>��%PҽZ�^�t�п/Z엒���TR
� �G�@�A%�z�I�_���A@0nd	l� ��6�v�w.���%�>�4�A�T鵚�XP����b���H>hbYj)�F\]����)S����������[��^�mf���5�B�e?�# �W�U��`��.���; ��py-�n'�.]���#	�u:X0�T�I�E�
!~��/Y*�@��G��h��d$5��� �SP[XC�_�ۋ��:�Ҫ	��`T��54�� t |��!�Y��hc�����Pun$���Sk6?���FK�AH&���P����CH�����SZ)����<��BN0����;��p�-���aUh�,�Br(�CiE��Z� �`���Sh,go�N�ˀb4�{�]�|�d�X�\h����@��,7i��� _^��W�L���Ҁ�w!%���(L|V'frN�@��CY HV+�>��H @^���-��	|�]u��X����	~��_taW>hK0o8��c�
	ҹKE/��/��W�G'�0}�v��!���,r����nT��]���AW�;,+��<!ш�eC��BlG6��5��G`�F]e$��9k��W��d��SkE��'���!�����K,����l���)S>x�@�	�h�(v�X��%�"��A�Qk�YO�	�w2��YX�
��V.��(T��8c	��$s�*H6�v��5\D$@v~�	�����b! �l�O���[1�qQ�%@�Q��4�!
m�%H���M��v��3=+�-[Qh�F8�;��;@v��t�%P��00R�dD�����_��Z͗�(2�� ����q��Ͻ�>�!�
yK:�nuHռ8W�@ۀɫ���G�v��7�~��i�I��P8�	�J�^p�	�0�^%e�&\��(v��9�U�B@}0QW�ح.-p	(�2��x�D!��g@�e�6Uv�
�t܅#��� k�i]V�����a��c���xT�$-5JH �}�c%Y0�e*P�)Š�{/Qn~f���e@��%�^=T4���v�~0y��{���Q�yƺ�����h7-AX]��K�Xm���M9�G���5 �^y��1�Ԋ[�V��xuq���+�eb�V)��0ѷ�gNQ졋RUe>�3� ��o�f&��1 �)ʃ����P��ho\V�_�0���%��$J�f&�T���&!��m���9�hRD�5%�Olu��@�-�Dy�<�.)�[^�^[�*Nڅ�Ȱ۰�ZM�e�A���ɒ��)����l�k�1��J���r`:��afgR��VI;S�A�������{�����������Q�_+U� m�`.,	�O]��Zh��.W���)�T����A����aD�y�-&N_�`I�*�O3����51 ��{&�p�0�V�9HB�;��yHȒ�����-l[t2eh _�K
��!CzX�cu���Ձ�Bo��f#a�N� ��������XnV	1�?#:�����s
��2M��
����E�	uX�^� �G}
.�{�;�Z����Q�!d0��zFh@I���X�L��t=UH�w �W5�:�(ș�J����zpg'��2,@�C&�� ^'	.)٘΂H>�J<b6�nd�y�.^.ߺ̮8�Vy�1�k��0wV�iMSQ�Z��O�۬8j@�K��u�����?
��~8X����I^�`��|��&����ל�¡@��
���r� R��щ�1t��[!�_��pz�[!K�eO�@�S+w6�r45�	�;*�w@�h&YZ�`��t�_#���e+?�$I.0�c��ỳG4�Jh��"�X�p����z�}���^�A��]��.��C�,�$E ��Y;_���~��J�������v�z�n�tk`�����u@+�	�B1���o-y^@�sq�*h+���zN4���Fh�ù��X���.KY�+��pJ雨�����Ҡt�"F�[M�z&��48��׏yl�9�I'q)(�ƴx%T��~E�����4�.��,�	6>�U�A�x�`�î6ph|��Wʋ�_����$'�,����ad?�����v�8��)`/�l�gO��_�|1��X��*�i��
y�v���"�Jݱ�#��,+�xj��,����h�M
�i�
�� �'��h%� Y}�̫���W;7"�A��/[B(�Txq�(�[G�*�{��|]E{����ل�)��A��Qla��n���� 6�<=}�Sh?zV�\/���i;����SJ=�+��^�=���^p\;�w[�/(��Y�Q`�k���%[�*i�m�a5I�q�x;��R��f�@3��8`Z��:��&=EƢ���k"��/��'�º܈CܛN:�,��*�����i��f�if�0�>O<
�H�����%�I0�i�5��,W�x V�T�K�l�	Z�AȜ�n'�^Me=�Mh<탟�N��vb�?^�>���*aHW$��(�v�#�R��H�� @ 5�\�JgH���F���xHo�
�I��\��`�Kj�6�%��E�N�!�o t��.��/b~R_>eM\0&hp.�KuN��ȕ���	�RY�h!O����l��X�s��.)ŕ�׀�g�_� (���@'ZB��������l5��1FĀ���fY�u��@�h1-�Qr��\@�O 7h>$�[�3 �5@-�$�
��i�o�9��P4��>L��V�2Z�=㦠!#E9`8�=]��~+V�J�fO�^�z�]r$_>�CaC#���<���0��09<L�I�/� ��� H&2-�du R}_.����8�r�1@qh'O0�XM_"H��P��=N�ЋDV��-pَ'���R{���-J�C�[N�) �tEe���[��[�}�~逄�]���Hga
h�3拌��4VN�<Z(��f�@��
�B�l<~�0�L|���g�[�нD�(9w	���-\�7i`t"�/_U�B��Q�=F@��(�6�s�`�<�i����8o[�hE�-*Y1P6q�����5e!��)�v,��0��Ѱw�k�&���
_���HR�)���GHVPl�A%��; �s�h\����
���o�����`:�"�(+2* ��d�l	-�=��a�A�_�(��Y���"(��$��A��W���h%z>���]��_�9~���> rw�<=&X&� �J�H����:HzY����0!Q|a-��Q�|�?e)x�x�rK��F��J�?�uhoA-X~$-�ZW��iej���*`��?T ^M�f=.��#A,bK�s�v���5�MU���	RP��ّ[��t]��}���+���e���w�p6e�{K>hJ��/RX� ���۵�����6��	���/e���@ ���<q��.'gޅRc��	��V��� 
�P$��W��!��V-���A��4��|�-�ٷs+Shz��Y�AB���nS�@��Ac.�B�тah�1j-�`�Pt���z��:
��R��3�,����i�����ӄ��{%4q~�c8ah e/��#�#	[L')�h+�uZ��$&R�Kc_w�YVQ� ^�S �.�x�G$@���4�A����N����k�e��P�R831��#i�T�
��	�Pd�L}Uh�W��CAȽ�F+1����l�9v?)�Yg@�K���@d�w��$A<��[��R���ʦ&W�8�k[$�C�Z���-L((�<�Jg ���6�J5/��B���_|;�M	y�~ŋk�S� � �Gd\�0]%��%�	�{Aֈ|�d�!F�~��Jh���~���P1� ��uF�$=Ry��`�( �J����w�b�B�=�����Z
�[)Oj�?��csu`5'_������r1cJ��*�\�`B�n	���/H�z��.����+�D�[J4�%J� �=����kw�#�+��,oad�h�w*����u����.�fp�.p�'��D5�ٽ��%@���@h�U�U�C��o�-�>/���1wō�-�� ƽ,�=�����k_��FsA_ t� �pX�J��2� ���3 YX��H�
��|7����<ym���0H-��
�1Ÿ� �"W�=$�RN�.��xqs��N��v��	����r�a���� ��Z��'/��A��|��p�<e�itݞv$ m�a�_k�m��8���H��v��@���z�v�!�cU>���Y$�w(�>�3W^�¦}t�)�Z�%Y�]��k(�zb�`��X�i�l�tHC	R[��Nb�e�K���Z^�#!Jo؁�bQ��"
v\qХWg��rxU H��-�Jv@��f��5�l[XP�=�|�%,h 5H��0)�+QO��t�󆂎zS|3��\ڐhMŪ���5'�'�*no	F?�	�P5�[��&sv��|�(Z�p3��?�0ߠ���0$D��1�C�L��y0f�D��%�(�����1��ܞ8�(�]�y������Ĉ�,XNR��e0�(R�ZY)�!յ�b	o$�n}^��mz�$�i.�巯��{S��D�K���W��Qh	�Zb�pz�%%���CK���!_���Xh�zQ�E3�S����~�?��-;+́��iM��a��������
3����M����]�P,�e�'tX�̤�0�����靆�Z�xd�O.�?�9�L`���
'{/�鹀n������Ƈ-W��=�0>t�n�����J_���	�x���>Hh	�o	�ǒ,s�M��	>v��ҼUԢ�8���̸�Xn��U�F?�zkJX%C���ԕ��[_��`}� ����<%�⑀@�.>d�⍁"�P��H�����KW�xG<h0����2�[ր�շ�%Q����X�@�<�������Ü��L�	�Q7$�A�+zm�_���L������Z<���x{ZQR�3����v��N�,Q���ab"�U`����z�nhd�R�\7�)�]ҝrF魯�6�.k�"J�>	kf���s	��f��X��P��w2%���Pc�H�^0XV>�JwƉh�j$U�~�����YF�4��-�o����Y�5���zI��+%�w�Y����g���x	;�5g(B騣.���|�Z��ܗV�x�8�K�*�_aލI?������]�P7�}w$pB��$S��">�]�`�:�Z���*t�����сV_��/�%���\(��������ԺZ�L(�݌0�	�2}�_^���>ƅ�C��(N�"�6���	�ܴ�A(�X�ba�# �ȝ����f�s�htCRݑ������aB�@��_h�O!hBh%�iQ�a�� ,iK�C.�sU@��kEIl�����0K$<E��� 1B$(��Q�;�$���.��01ˮ�0i!)��L���/�"��ꀰL�7�;h([׏��)O��8�O�9� .�'A���f,Yu��Z�c1�Ѐ�o!P{�>hCH���,��Q0�gB *�R��y%r�X0A��P�c3l}�٨��Q���ǼaX��@�5d
�RT�\�]���3@f \�����b���X(��F]c;�@|�Vo钏�r�=a�� @1��TK?�83<�3/��v	h�#�����_!�����=@�Enk������T�PQ�HH�X�A`脾�c��H47�XQ�햑ʭA�PQ�%�@���ȕ L��&C� (�Y�KBEWf)sΐ�/�M�����l�^�v[=�޳� ���@��;��c(0���L�k@��3Rh)^�LX 0� 
�~V��� y��˱��x���e�(�)�^�M��ӡ�V4���v^����0��fŁ@�\A'!,�S}��p#XM�p�~��	��Tq�_�\�)�]C=�L"�d��wP��-	�Fx^���߄�����k�T	˭�h'yQ�	T]_Q���p^ �J�Y�IQP� �VR)�-�iCr��.�;�>K��1�0�~�&RA�:9b�w�+�s�hj�f@�a���X��8�-�dc-��`H�8	b�
��Q��-lA��hC�抉�}��̭]+��[B�!Ȕ�5>�h��߰�S�-q�#0eM��%H@���j�C��!��
^	��,\hO6̱� ]LZ�"_V_b��!ws�0�K7Hp� H�1ꉕ��D[�(�io�|�$�~!�b�_��YXI>���0h;}�u��o0E�
L�/��@ʑ)�J��=�3�L�͐YU�P�$h)�H��V[��*a��8�z!�;��b�VV�?&+�1����$YŴ���;Z��`����G�xN$��SKz ,�3kf2�����	D!n�#r���T�I���I��D�x} N�<:��]Q~�rc��>R�G�mhI���&U��+�\	�3+[W�2A�J����Pa���+G`ht�����e�ӳ��V���	���__�V��#.�"y�o�gW��8nWp��k.�CC�h�5vX7-��Y�]et2�͔bGr8����( p���wA��j��6���\I��Qm&}z u��)����ęiY���sP���w0?P��rY���fh E�d����u%\F<z�ƥ�W���,�T�]!��'����;�ˑ;�vi�@|rP`ʫ4���0�#��@�H��2����/�G)�X1�"�%Mk�!�u`��8Xr�{P#1�_�_��	�8Kt>O0N)� �&?N�ڤm���tY3���}��.��Z��^[�`�q�^Q(��ڒ��*? �=Vc��Ĥ �<�Z=,�Pt�P?,��x]�?�)0R�h
H6��L�����{Y8���'F���7������P����G����7#�k�m'uv�aX���kNU�iPVh�4� �A:���,߉��L1g��P��Q����~����.�@��S%�Fjh��4(.�\�
齗�-u0��~:�|����E �TMJV���[��0 ;��Vd�Wރ?]� fS�9���,�� �dM[HS�+�L@���H)'�[߈�|�	��ϳ�'�]%�	u�_qW!�^+F͉m��EYh� �*s!�XM���V)��$�p��(�R���]>l1��J�\��&�Ђ��<�+e��A
�r�y\t��q�Z.���k �Ʌ`��@�/����"J���d���e���l�T��,�ߨa��?����*�Q�S�d�LUQiHu�A	� ��0'p[\T��	]gÏ�[P �V|�ߡF22�U�Y�DجT��Guk���Y�!����<j�'y�����^��S��I�_�f߈�(Ư��o�p�qs,�]�?69M �J1��}����ZD�"�i�E������X��FgN4L�z
�
�Y�|P�Wi���� %B0N-�?�����B�x}� �o"�ش	_\�v �Ř&��i���:4���CO��ШX�TLgq�B<#��;4�Jj���O��1@��*J%}t��@\�CJ=�-�X�܁�X���1?�k�2[��Z��~(K��)�鈻	�k��:�����mj~}����Oz�T�X�!���| ��u0�˲x�(`�
���${1e�O/�w�	�� ���ϟx�N!�c%*�z�)����J�����0�T�j0yY,�`Th�2O+��J����
U5İ%N�x�	jkG׀z������_K(�a�\���p��ٻ�@�n*��&h�K��e�RXn��#�pXX��fh`W��� ��-8��	���E��έ}�[�s�|Jt8�B	������J���?�����U
���Z�2�����g�M$� ��Bܰp��0fT�^��o�
�Z�JB�hk��"X�a�(�o>+�K���1lCټ|�i�U�Fn$ �\o0~]��^�#�ǅ��v�- �hm��J�^i���j����~/�K�>N�/X�~8nN�p��d���-;�)��P3��K~a��   �X�h�����Uyr\�t���r�}fSV����p�b�c�S	����=��M�p�@��g(�Z|�s��v �Y�H"	�F~-��*a��
1�U��E�_���Ճ%��p�.O�fZ�� Vh	!<�_����=�[c��X-����w�'�\	/�8|'N�0\�}��b�zB'�R��u��@��~�BM�e;�<W `k�JǴ���o���b��Q�Q�Ǥ��0��|�����u��%���J؂�6%ݞ^�P�m���;�z�Tq�N�R�x8P�3��k�Ȁ��1�(x]Q� �8ݜQ�� �tP�e��A�d�\hAL�1X�a�cP�\�J 5�}�{�G���[Y ��y�y�`��JXH!z7C��]1��n��evB_�( ��c�]Kvh�w6gz�1Q���	�h9](%�0��e['���6Y���� �*P����4���:�5r��yU h}t"]�1zb�X-�8�v����
f�ʩ16�S"K�1@��PE��z�ݪ�0�;s�`F�Rh�y��.?S5��~�^����	�	3�	� �*y[ �7�`؅�����'�r�G)�I��@���v|���a]3#��j��=�Z�M`�-���'�+U����ϰ���X���,E)P��A�!e(9�����*���i��x��mA�;lX2.Cǋau��?�� ��&����RJv��h �`��L��3�*[��zF?��� �ft�^�sE�)��Y�>z
��� ������*<��m^= ��op��$&u���_(�B�G���Ϭ�Z�$�,�� �w �)
^k�ɷ{U�N$F4I�(��`��7�/�W	 �V5'ߐ|�`H�
 �Z�W"�T�Q��I�k�^�P����`�)ܴ�*�%	�~��&����hܷ��L���-ޞ�p�p���%���S�T�@Lq�)��-hd�,*#^o�X�z)n�@�Z���"߉�|�ke��Ě ����j�__m_'�&K�^���9�/�^�V��W��&x(W����6� ��z�`d���<E�{��`>�/M�S!�;o &t�g��G�o�+�35��[��/��|�ժ�93(�u�������8�#	�Ͼ]��g�������j�4�
j��%uDc-58A���<Oh�nl^6��<���g/ g(�Y �/h
��9��!�: 8G�m���UtP��ןS�4<��y�.�w��0}���`$�Tu�vj �&�%��SO~���5�]���J�D%�(0��)���
c���_h�j����w� ���W�_� �ʇ=Y��	B���	��!�_��-Œ|k�P�{ 
���-fzD�L�~a�;�{�q���<@�4#�Ar�
4f��i�\*�5���@ðP��(�0����ܶp�������<Æ����g�?���f[ �U.ʷ���l0����ƽ�M�1��a��Y�D���
w���8��w���P hQ(RX��:>�u)�(�؆'��`p�F0`f��߿��k׫a,jC|P��qS��2��_��+�`�ӟ�8���n+;�X�G��ԭ�))˽�p�����gE�m�޾��TtW-��oK�ͫ?�E�#����t_��rOx�]�:�8ɞ�VM�n����`okK���LA���/�^[��J_�R��ȵ�jp=�3#^[�ԟ�n�d�(�RP�\q�険@���&V�/�ӹg�L�v�n��t��tP8,S(��+[Ye}�&� 5�<X7� 4��cO^�����$ �ItK�x�����0�G�7��/}B��+���@�L-]fՕ���o��w�@�b	���Pa.3��<�8z�JAa�����}cq���*I���/��s9BQ��Ap.�~p	�[h�\�O�/!p�A/�"h@��~�N�[]���b2	MF L��X��L�/G�����L��y��Up��ء�dQ�x��\���m3 ʽ�n��p�6Ϛ��wH}��Yh�aHס�Ŧ1ݺ^B��2r�̜�Q��y�$,�����v��4���+�K�͉b� ���0���if?Т�O�z��b\UY�܅�$>��X_�죂�B�}�pDY�|����ո_�8}�����r���9@��UAR5�A;��1�U��ۄ��W�L��h�tX5Y�ɦ@K[�Q�P�$�P�Q]��Z�̡���LЀ�7&u�H/�Y��E���N�Z�(_#��J���� �0�T{� �N�򅚉D��)������cN������5*g�Lp��0V1�;fzq_B
-�0�x%&m!��h8�_?Ԕ�lk�~7fW��g�K�n*�ª�0���X�����*�][�C"�9o�B �UJO1�DW�Y��R�.S�t��ݻ>!���	k��"��W����M�:�0�}��G:�),�y��E��fPW��O4�A{��8�Npon�_	��D:9�#�5�`+��u5i4<�Z�d ^6�{)�Y'[^�T�Јп�h�,�%�S�AB�Yw���n��%�?�' ߿�#�8�GE8k>W*������Z�,��[ZB��=U~�e�-s�VV< ��ì��k�e�)s+@R��	�[�U_-D7'N�^��L<�y��U��W�ZK)�J��/���|�X���Ԗ���3XZ�*1�8��	�+
_��`h J�q7 ��a3C���T:!�U<�K�+t ��1��4�"0�(�ˁ������4gc����l{��K��i�n���wr�&�ֻ�˜`nh�Z#ɻ�G��9�P�<�J�r����&��88#F�"�+��v��jE
�J)f� �Jt=W��vW�	f�(�h��X�jc�<�2�p��������:�N럍J�4x��L}�E�1�Oh��ՌэU&����<Ȁ�h�4@Z[�s'K	���Th�L8:.|��*L�<fX��F����,S��E.���mO�Mu�$�U"�p"��}�iY��br̠�h�s�_W�7�F�/��J�sA�p�w��"Y|XP����&�"�X(/d�Z�\��]w�v��l����謣�K6�oo�I^.C�c��+صW;��+�|,�������w�Xe�y@����R�#Ȇ?L��'POT��@<�h���D�R	k�5����<c�!иU%?�D�ØV�0*� >��]!ڸnD-@H`k%~���L�a�W�����x���
�Ҭ,r�3Qe6Z� t)\GE�BM,Il�ʇ�  2s����v	)_�h;��y�@vY��_Xl��F% �H�3)�@"���tPۈ�<l��� ����1N)��Z��G�iHW!��r�>tp^L�%@�[2	���h��=P���X(��@p���L�/e
��SY��!� ����c0���dt�n����O�8�q^�3��?�b�{
�C)%���`�!��[��Gx�(����Q}'�M�}"� �xYRS��*��+���Z�7�D{t�q(���e`���nE�pR�X���?�3S��vD�7��P&�!˝`��� 2W�3&By��1����8H�XA��/�=�%�k@ ����p�log�xi���eJ<����bl��fS��ǣ�tI��=�򼾁Y�A��H��N��́;c�n+��(�����n��k�%H��L�������ս�O\ \��'�/�ʗ���ί�	�-�؝q���(1%	�D/��������;�g��揈���رy�	�#y�T`;hN�gQmہ�+�`���;���K?�z����H
�S	��;�h�*7'`���J���ي�C;̍1i��܍�&�~�T��K �l����;8�p�\��z0%f$ }����()����7O�sGy���	�'��l�'$P(�dMu1*���)N�Є?G�^M���[���`�Q�df}��c!�'�o��	��
y��!�W,�\e���P��X��V�K	�}%pҌ` )�!ݷ�J%��~���:2���z�)ռ퉄�U�]�����"1�
�#�	����]vC�@��^��L�P��=3.�σ�靌`��z�H+���7�-�]T�����jv/�c�v���1�Ȉ�$0��|�x )�
�k	�w�ِ^�J>>�X,�+�!}M1�/�F������,�sz�j �|�5�����Z�~����?��Xd�Ӱ���[��P�zoTx���=�V��FlNW;�h>�.D�v/5Y4b�,"�O��!�u����KX�-���AM���c�H�QqJ&X� �uA�� ���X �Z�����'����[g�Ϡ>#��D� ��`7��n���6��R�
��U�h*�{G�
���%�-c^��J -��ó�%ߪ�[�����w�[U.P�'?W�7ؽ�4�Y�Ȣ}ow')�D��t:[ ���)�p����ΜZ[����"��%=��O�=�� %�쫂 �U��Il�$�0�	R�����%���"B!`�e��?ǹ���n��].N����ނFg�|�/�:��pUPCݺ�t]��+ ��;qx��lJo �/p�V�	��q]~q�	��TP��n	����0񒕒R�ٸk�]'[a�����|���N
�-��晆�o��2+�Ψ�v��g������^���]��TmAS���4,���]� �c�ҿ[�P�[�B���.��b�RA����X�34�0y��W/khE�,�!u�
h�k_�K��#�2"���@!�%f^v�i����\�кj?�c	�HaH���ן��ύ}��U[ �'����U������D���y� 4W:��1�t����2e J�|����y=HiUT�e�m^��hz����b[�Ԑ网AgB.����FD����-����S���-�g`2)�P���!�
1�Qhcj1yz.�-���rKV�"I�1
��ޖ�HPyc&3E���CT�n~gh���Y4�F,�.�1qZ���>�p�:x0
�gdb`�/�0�p���;�J,�"��ΐ�":��%Ȱ�R/�v�������N�H�����u6���Z��P�-�%]�T�BL���ǤTW�G���P��b.F��@��W�M���Ä0 �[(g �^�����p	}s�BO����B�S@��9E"��s\��[�p �E�ˢxm���@�OA q���>�M�%�{���Iy=O��j����顆���� �_�������Z��(콰\Er��
�j0�nXw�v��^�)��0(%U	&LS�-^@'_���CD�%
}of�/>��_�W���N�p~d�VU�-��S.�g��+C�	� �^-�b)�L�( �h�����M���$
hL�&@� �Q�4KK���[ڸ�J��+^�1 ���GR=x�P�^�E��@8`;c2~	GiT�P�>��H= �by��`�Ks]'vv�z�%��Wt�z����p^�V�gMT�PJ�<��v[C:��>%��@���^��:�+_������(G>��1�{ �j��~ON"�־]Y�=�}mH�-���� PA�&D�q5Z�^��Cn�E��� 1Z����[�¿_� ʯ嬥'1�����W�B����Z~�V��k�bn�{�	'�Hn�$r4��c@��Y[���7��(�	(�3TY �Z���)(��ς�������:���IJ蛵���C�;Q�`"f�X	ζ@'!qB0�Fz ��0�xR�"l��� �-%M�s��y��8�b_�s/�����ZAb����	Z�-P�R�B!g�*�d��tGy3��xKz�p>�p�E>�Е��� g�F�|�w_��oS?�ﰁ3�(��a]?e����&l� P�8O0i�,%a����4`1��^�PQ�W�IN]�V�(f�J{Ѵ'g���!���]z�XY7�@7�O=�w�Ó����ֲrԼ���l�%�Y]F�5�k�bO��nx&^�By]J�K=�7Xr	g�����8�	��B�WT�K�A.�t���
	�?gA��oZ�`h�Y;��^0
~���S��K�PJ��{�p����,�/e�^������$�5%P�#�d�hQ��@�U���
V�3	ܙ���2�x�d�<�q(㔟��3
1�����<��xKr��W�0��GNͻ/�^��!���}��ш ��O։����' ��tNfs�L%nTUK�6
 mh@A�YZqB�� ==-��^1ۜh�4������m��fS���"�U�F?}�r/�`-~���`u�F^
Ijw�fArGx�-K�&	��)�Ulҝ\o(c�udy���
��^"-}���	�	w�{����~�`�|(J�?+d��H���]�!O��S�?{c�<h�p*̽�PZ�!%�]}��[���i�
]!N ���͉Wa��!�1l�� \A
'���:/Z�m��1U��B�����KK�a���.����]chdS�+ٔ	�v�zW>?�G1i�O�|�ۯ�8��ыh���k�e.iPS0���(�[�΀�VI&� �Ux/[_ɥz��K�`��Q>BYAj�PJ�k��� #K
Y]��G��pےf��~�+�x��e�j鉁��
*����� �\�G8�n��
/ՉA����[�59�X�%,"��x+���0n��ug��E�~�91�K�9�K�y��p;���Ks(f�  �_@-�$��W;�CQ~�}�%�u�ζ�������Z5@i%g
�d��v�3u܍*n�4��O�������T�����J����T�J���lP و[���kaǾ���Ԁĳ�K�����$Z�������h`_'����C�4Kk���37�_��pBir.��� g7���C�ʨ�K�j�鐜����N� �R�K�`�X��}�	qP�p�6������U�xg�k�D	��B�T.�[��c���
����4������7˹�I��F��U�h�����[�_!�b~Z6������a5�C�LW-�zc� ��$7$:fZQ�� 3���Xo!-�	} 1%�]���*��҉
�{�t!S{�� �&U��h_���		OAu��S���^�JG|��2�3�fR�9^_Y��<\?�5HJJxŬB���v����qT9��p���v~�j81�Ӈځ�f<�U��ޭ�[�����ݯ)C�o"�Q�r��|�`�JQϿ���0���Fr������wJZ#��<�N$��*	1�s�P���Z/�|�R-�{R#o�(Z�t���Q�f�o�{�uY��ޔ��"-;�)л5fD��b�|�'!�aB��؋�"�KK Վ\��vIb�-b��*�������v(W���(Z���x1��)_�[G����m���f"��1A+�
�q�O�o��AC�uw.���8	�I���z���-�'z5�#;S�@��Qր�X��M�����������"YZ��<U^\�mx�^D	�H�:�{<Y��h�X	:���1�W�C�����`o�LҾ̠��{ �[�AU���K�Ȓ����O�e'p6�bp2�t�c{eKΊ��R��m�.2�E�J�B0I���@wQ�}��1.Y�������5�.�a�� ��	��<Bnע31������� Ֆ�:�wo�NH7�^���� Ũpb>1�H)�D�:b�¶��Vs�m�Wʠl��|'>�&�#�2�$uv@������*N�] �z���Y��6!�ܟiՑ�5@��eKǐQD"Ē���_-h^�_�Z������Ա[z1� �?�~���]��˱�������Eiz� ��4hLXpAa৶]hC�^-Lit� ��� 
 2p�8�J��V$d�\~�A�57�`)���P��-�E�*N;��ޞ�+��k����4E.�$A0��Nl��s R���ʀ�"w(Z ��	~��sW�i_ ?�����\6Qp2��xp��X��G'p��k}�#�/������U��K�@X���V4zŸ����m�$7��`~���L\�5�H	܎ ���������.�OZ��s#,z!�^�"ޡޚ�?cFC	���b���/��7��P�fe `]?&��i���m��_D�}������,|��dS��l��^'��}&cw�%^��U�yV� ��L!�%��}��<5�NgP�1)��v���� �nV�(�&ڝ!D��o�#��|�� ��&m��d7�+�Z 3)YVR�	�:�3s�wK����A�z��ӫ"����\h�1�2�^?,� HD�p�谯4��0��i���|�O��a��̯�q*�PT�!�o1�	����E�i߮�TE�s�P��iq0��D/j !��[P��w�1�o�����{ ��z�|���S�7链qA�x�o�a��	��Q,U��dUA�R�}���\����-����h
'v2%U��?�H=^@�T��ޗ��x����u�N�%)��v2	3_�H U��*5�����`��m�-o1���(���.Ke�؃fQ��(o�D���~��"h�}�����5��Y��	F�w~Z�|�8�l1Vc'��	_ۊB��A\� ��b=��Z0�<�+Df���{/h���/mK]`~��!ؼ�`��	G�F3���hC|M�����Z��{η�KcWlU(��$,Υ���v�<�F�rZ�	�v��e��a SP��y`XY<I��Ɯ�e�4[�|��}B�8\@���7��Ѱ�Y���)�w5��dNa-��OW~�_(��-n	=N��>�Q��-V�[�=)`F/U_�͜>PS�	GKBV=�e���鈤y��Rh�p�?BZL�%�.c�<��.iA��ᙴA�1���!���8��_�V���8d#>	fcq�hu0��/��xL�W3��aR��u��1�p�gZ��1wgd��X.����0�i
I��)K�u	�_ZC�;�O��(5h1�+�[���N[������{F0��G^nz�U�^� !Ä>�.$߅	)�_[�
[-� ��Y�T0�pK6�ظ�8�O����'h �I�(XH��iF�u
�3��Q�V�_ܼ��Df]PĂ��Ch��5~����'��Hs��\�[;��F~6�8�s�7�%)���@�^h>|�ZE��͠��/#	ԁU�28?G�
�B]؊��}Yvc�Sh���ȯ�t�u�$@vI��"ľ֕X��o���@{ �h
C���<њ�%�a Z;�`I��R����-�[����	�R@KYX��� 1[��)GX��	�������e���z��L-�tob�`DX�w�N�����D(ޮƿ�[����L�`�*u8��U{$\� ]N^0�1'J���� �N	�o�U�wE[!�G�����_���d����Nk�]�$�Y�:��4#�o����{[���[����W�������88��λ�#X$Q�����1٤:M��,���6ayFk�"z���VOH���B_Z)�:�e�	
�~W (�X��f��.EҀ�m!	B)�[ �̰�,�WPd)�@��1�> u��~`@�;�?�ځIA�� ��b=�Bc}.Hx�w'���|���V�d|%S]u�y� 2���	�KW�������nJ��{�H�!�0� ��~�{�=M��5ΓÙ�
/��1�DH�Ox�!�(��\�-|ݼ%��'г�\���p6x醾 ��� ��A
`v��P��?��I�eiva	񮦻��Mz���iZ{�b���"¬z�}wdz���(��XM��Nݩ"��G	�Yu�J1��U'*�6L7i�9;�vœϞ���F>�ˢ��������H��ZVh";}d�J���)��=�>��X_� ybs*��(�^��{R�^q�8� 0MaA�L �*�0��%�h~��^���/��u����� ��2�8���kT#���*F�r.�j�m�o]��_�b P���}�ȃ�@5��v�Ydت \[��j��?Qi7@�/)�(C�-U��	���	W�S���>�|��.�<�.4�/� x�^PW(�A6��=L��q!���?�J,k�-(`|����!+��L�M;_
�j�I�7�quP_��^�[��s��D�^1��
�*�i�<e�~J����S��Q]�Vz`&G/���@w�~^���E
�:��T��,(1�O��,0��.x7]餁�,S�lp�	���7���)���K}�X9(�zh����791�%�V�P�kC�� ADPKe��%��S��z&�65�8Ue����"h ���a\vD�Ge�qH�s	��`W䇁�^:�ؓ:�[z����ihz-_��"�<���;�`�h`�� �[7������5��c�f���UӑF��L]���?�H�'Y�*!��xᠻwGQ�����`n!�|�о9:'U��k��ت�����^r�{��X���l��������3| �����*@o�L"�.�� )㝽�+(@��d^�y1��,��;���~�Z?���+�w�z3+�12�]TV6Wږ�l��;~����'h�bv�/���i���o������w�C��נ�EV���ZP���X�x��@�D�l�>0�`��[��A�P*�9�>����:������yҨ�`t.%XV�	!�w�+;d��N������k�ҁA�zA�p%�GzA"C�j́8� <a8��_�����Dh#̐�}[3��:��T�-�G����U��[���	"o Ҵva����N����q�'�y�-�. �>Q� 1X�p6',+wF�������}�rw�!�~TUB�PC`gVW���@�651LL7�y\,�?�4���Zτ��Y�sT�C�LY�f}{V�)����	.Z�N2�a}H����+o_#	-B!��0�p�� �qU$���%���RG�F0Bh
-.�^L!��K�' ��n-JB�%�M@��{�3��)����jfb�2���%�h�X��ɑOo�W8#��PY<&����+}�Y9	"#�A���@	��/:S�����	��oc��8�#\������@T�'b�}>��yy1����f�����h8�k	�v�y/��<` er�l!�Ю���r��{C{[�1��I V��6/O-� �]h$OTi�����,�aRL�-;m�K�(ذ�-Ősy�J6��?td3&�����F@m��=8����\1��=_b��u�p�JP~Iu9"wO�A�PK�!{�,BgC64���ufN���:�Z����^�E�/�Fp-r@�Vh������RUѾ�z��2N�AJ�t	C�ZK��z�C��7?�x��|�R��>������_ ��2�a@�7�rI�W�4p�/rx���/q	�҆(�P��� w5�l�OO��:���긻;VG�7g�O�1|u���4�{X�=s�v�ԳB�g�#t'gh_Y�f��#h����^T��`w�b]_��
�6y	LF_�� Y��@K��d1&�Z�&a�l,���Jh�2)�! _��96J�C������g%jK>���V6n�X�A�W俹A@h/�>�^�M	6黃;�CQ!�� =
^DXV� ��[���%1T>�It5b�`�^h8CK�p�-F?�XV�K/�=�ׄ��F�/U�v-6�*D��^��N B�]Rh�L�4�V X�Eى�)�[Z`�3Zi�V �5:0j�GYq�:�~�?����l�Mr���`���ȃ_��j�,�n���-h0�j0�r>�sf宵o��8�~>�!A{�.��u�y�,q�`h�i� } j�,��Y9�1d	�i&�z�M�I�o�t2=�@��}��- �Emu5�`		��\�̸���,A<N+�w�(ttiOv�_Cǜ������¶_N�ktȎ��J	�5<����i P}���cp�WQ�3�7�rc�A�3�adU`�rnäS�ʦ��'��Q���U��|u{�>6)w�3_j�ԎK�3�z[�������3����Joxޗz������%,3���g5w��.���Q��L��||	W�\� ��KD�H0?a��!���)Kɯ�CM��[�⩃�AuhF-�Zx{/�Ւ��|5	����Lc
�9��}���-Ԧah+]8Y�F["K�q�
S�qzh��^gaw�
{�롰��nz	�x�ɼA_����W�`K���cK{|���R���f�=��|gVD���<R]N,��8U�P�-!������T�cPs�t;	�A*�4��@�Z[�k1�j���� ��Nǫ�UP�(C�J��
0U�v}KC�	�#	U��$�_o�����<�9�eͶy�!�S���%���]@6�(+[�v^%վ���S�����k#/
�֗\^`U��'�o)�PkP�~�:�4��Q�����:\0�%����s�6�Zi�X�,�Exe�0��aP�{8�[,L���P�Ьh[qX����z�E��U�]{��]E�%�TR�j0�PW0=�@&U��W�g��ʟ!�2X�%>��bC:�`7)�`���!#����]}B�����:<=�Ћ]O�f 1�!��uoP�p�^���	=5_�	��0���^:(ں��Q���i�!����R����\�C��&=$�I� q�
��pY�/	=)چ�V�]<Q������UWh6i�Q_��#,81�A���o_!D;h��s�#<�z*���!5i��	_h�GD޾98D|#險4��oK��F_V�S�� �y�dY���_�=S]�H���G>�Shx�B�r�	�x��R;L�@(_ؑs����f�K� L1��R�4%��0驶�%�B<&5�0Z�$����sM)�+����œ���:Ż�˽گы�}�&!�_�N��'���3T$WSR��4��[�Qy�`<N�H��PgWZx���@ֵk%"2����-�
��b�KN �����o`$�鶮��7��p_��� �fQ���L0ဴ]�à���pə!< $5�L�`;!��CZAc� |O�@�	%BG������w�
��M�����GP{�^h�2��[��HH�B�����t�Ýx�cf<r[*�4��5�/\�PrF-��(^X�p�h�[�z���b)��J��W�d�R�ـ����\��O�į�c=��uvt�d�pH0�5_�B('����]���R���_	�d��v�U��^j
�o�e�ǳ�/��-�`}��Z
�U ki�~eL	���"_/	�A�@|oX5Pód��	f�]q�I���7��$��"0� �,� XPY�dP�	o/hW%��3y�c���\j���@X�ёhgk̯�+�gj�բ�n`ẁA�n����]�(���?�v����61\�
�AR���&P=*�d�QSh�}mL�4wuZ|�Í>@Tn'�Q0�Lx�h<;8N���u؂]��h%V"� ��4(���I�z��;��*L�Ą -|
�F���F� �NR��*@n`/�����9�%�|��B4��_��D������:���1��,�0	&�\��t\�"�V�G����z��˿ަH�䓌Z)��k��f�о�I�i[8W[sO�")w�&nh;�F%}0�"W�� �K�#- �?o���� �;V�HM O1P�0�X���RÔ��{�� ���s�~uQ�>��t#�B@�v[/G+�Z�]���@1N��� U��{�C�2L
+ޔ,�O�1hez�����%gryQ�b����f� V�<_�N7m��A�Ë�NX��3����"@��'�+�����xջ�~Z= ��	7靉U�<IL�7�;�\��S� �A������i*P��BI�.)���A�n�F��P7�]!���5�h��V��^&r�|�!�3ʀ��'�W�:��ŕё�F�3�J\�g�x~�Y�'
#u��1�ʏ.V�^
TVAg6�H➖���5�8,yP�)�Z+�	:�-	_�u&i�����>7�۱� �X����j�� W�<��x	;�m�2NU�Ӫ���@z�(�t�r�CW�a	��ߎ�0P���;Vp�ry S�K�����������ZQ�4;O��D+��G5�.j�$o���q�+ ��y�1�)�R1�ڋZ�2e|&�c�
���O�m�{-i;���I���A`���O`�� [1�h�J%$����J�JK�o�HY�!���� (��*2�};�7G%H{�U܊=']VT�1����δ�y���`Z� ���_
=�/�Wӹ]	����.�� .����1{�@	����/��^�1>^[*�W�Kb�g�ݿ��j�^R)q�x�d��q� s��1&�_����`�!K�ʭ����6���I����΀)џ�Q�q}���0�:�!>`k*_�H��'�QVfbY_�u��ϓ	DW���BPV�i��? ���>�f!�[a5�>� )y��G�0�qB�_n�cW�+���N�3|�j�����$� �,xfh�*��H�R�h��q(����)�J��i�^���SE�결Ga�20�ӈ﷓M�~!�V�`g�:�T1`��s�Q��=$���B|�az����#>��	�c�9 Y�;,j�0)/�1 ]�Rw5�0�^3 "\�~鰱�>�`�r;�Ok���L �gQ:��zA�/3y���|%9Sw�J�*4F��5t0>���N��#=�'�GP��4�E�8
8X[���hiL$���^�h��2h�3�^Q��'�{�;���|�[g��ON�0Ȍ��`�SR8&5�Um���g�<���By;K
U�m���$F�����}N����/�&��]��RDdX�W���$�?#�%kA:h�&{0���}��[���}����EF�^�W���fOLn7� vQ�[P`�;\����%�v� 6�����0)�@:K_��8�IO�k���Q4~[^�ޟ��,(�Y����,)몐5-%:hb������a��Z:q�u�
�+�c�s�l8�T:���$8�	Ѽ֊���%}t\��QLE��z�����ª"��͂A������	����Eվ���b�l �-hz�G����QX(J�(��6 Dypm�{�ik������q��u ��L1*E�M�?'B�;��ZgIo鑗xJ���$�H"[UHQ�eY����!��J��W��A�Ť��*��;?�_-�>�L �)zR�]8%�t�D�}�����J/`�P� -�r`>Ⱥ��^�Q�%���F�RH�Z� t�a)��*	���8b�m`�������f3K8T$����i�*��	���U�9H�%���B�\���%
�T
�e�h^-37+�O0�4�w'0X ~V�JYUhZ�ǎ���YsiG��<�V�ԗO(��y�hV�aY"=�	���X	��'w��T�h�dsH�C�d��K��}�������
�-aG��B_���x.�-n/�R�\*u ��&�O/)�̬�#Z�U�UZ��!G�n��3�_I�Nt��B	6>	��O�_<#�	�NS0%�D�&����5� �@��!ؿ�/'�QH`�S7�����
U����)=(2�U��	�Z�|�����ꑎ��H :��.qN��)5B!՘�P�	����_|C?�y{���.j�RW.�̸|t0A�h�1j��)ڗ���L��ْʢ��X��L^,�hݸ=��(�&��O,�?G��1���~t0-�fpPQ�U3g��b����-ޘ�q��N-8e]F%��:�DUȱRq-�m�	<DFLAc��P	�e� ����p��wYUX�sZTТL% .ӹ���������Ы>� ¶{��
���l��J)�}�]����t�P�V�
&X:�^L�@�O찰W���	�x���̕B�'� C�0�ww�D�hd��"���u�dG�G�4��U�V�OA��%�# o#��)W1{���LH5�/��d-�N���
�ʠ���-��\R�����s�0���z�j�����z��
�צ�$T� �C�?���J*,A�ufL|D��'![W �W:h(�����fP�/��VwQ����[�Q`�A��UQ�@��Y-'$/Vº��UlG�0>(�c�'��Oh�_���.3gJ$I�uh &����p�A!��Q�
��ѕ��h_s^��h2� ��$�@�'�.lXj�|�r����G�N9�Įp��Nƹ?�Z�,w�~�@��@�f!�1ɵ��i�{h3|���������D!!! �vq���VH�^�?��Z1ݒ? Qh��%Y�y��e�o��&s.��X�O�5!dh "Q�MYW������Dȭ�ِjL�p�<���N��Ru�(� %�G���̀������X����6U3��{v���.�@3�Iif�G �Gm-5�I�D�E�c��)`�z-d
v��M�@	ɀ��C��ߡF�2�uT��C2�PB$ ��t�K�^W�C%אcU�=)T�#^��K��Ao���7T�a���kM�>Z`�Q,�����%O1�����$0�B;��D��:P���v|ݯRB��~��f�rN�;���j��Xc=�)V`C5/�_�!�h�J<�7�Od�f�GxD
Z��{P�PXѺ	�3��-�.JnT��	B�U��01y��eW�G'歝���e]��fR$�N�)3_?V��M,ftH��G!y)�0d�?͌T�`@��1���x7�TDQ��(5J`��1Qb�i���	�uW.k ^�ʀdQ������W"
<�AG� 	W�D2���S��������T�XS���v��`�����2'!�9�X{XD���'b's�zJ =}�t�입���	���VTMj:˸$�
 �K1��kfp@��=Z9��;�ܾ��gb���$���4<�jTl���ς`׸Z5yHa,i;#�}u�(�1��"�HE D��V�Ofa��[A1��+<k��2�_I9��"��a?�ۿ	� d
 _-\'0}��^U��c�QR����d!.N��to�L�X���?WF/�b��-�/��!���=�0$�d� ������� L�
!�G��j�U=sQ���-s�?�%�A� z�� ���r��L�k"ז�1Ywu0�M�4=_Q3�����+���
�T�!�9����-Ϝ!TkIݦ�
h�K���Z�'yׄH���S�9E駑����w�H-�L�9
���Ԏ%#��(�%�-����	�%	&E
B�q�-�h	_M$Y�5Y~��z���FH��x���wsu0�9�\S��h����g\� �\P�Q�#5BǛ���%�,}|�w�$A��	�ӏiԈp������(��ǭ h�E�t0�[�_����=���1J�ܻi,"	�u��i�ǁ���+���H)�{���lg�	L_>Q�\Ԏ����
�X���BfK�(��-��Py0e��U�&}D�%_(�]SWfa�m�)�BI:��A����1����p�:�ɔ{��i2�J�.!e�%�o�Uˀ߸�p8�(�S�mZ�k[0����a~)����B�U@�r p"��K�&BQ`��!)�YP!���T�H��W�[)��
� �}<K%6 3;.518
�0N��u� ���Ȯ���}Rl�Zé���;� gƻavH����_P���Y+�j0��_��
���;'p����r�_�#씉
��!KHj�3�x	;�x}k6:�肤�?b�W���u&�P'��k&�2����(��}�n���� +�q���j�Xِ��e�>P����k�����h�M>��5Dl`�2��`K���>8���U y<!_[�g��Q��r8�Lj!�$�-V�/]��pH�Z
����o�U零���S��T!ˣg���@����IPL%��f#bHW�"�w�2��r1��X�� ��:+ �V�u/�|0<5;LUp�����Ș��L��^��$9����@͂�@ ��� �.�;ioBg�=hf����T���?&�P7��/H�X|	�</ cՕ���nW2[������:S�AS����P�6H��%Qxs\׀X|J1.��?$X���e3ZC<	 �Y����3�����(�|��k;�h�%�-rX��Ii/,W�� ����x�p�X�00������������ұX?���6 ٽ	�|�qy��/�a�j,�n��-�@I��]bRqd�8� �r&y`�(qaD�����p���2��������wf��GI�3��h�6�]~O�t��z*٤}�u�%�?�~ ���\�۰�W 1�	���z���t�I�z���� >�4;4��`�G��y��H�q+��Q�gߍ*�.�k_z�jR_�J`�D�)���'v@��;�?�OQr� �$,c�7f�d.�-4��c�7��.��A��A+�z�ժz��"����7�%�����L+���-[�=���+ �D��V��	�F4q����'.!鯞�^)�\Zp��w�A �����0� W�wW��Kˀ��Q8i)�_�h,M���o���(ʝ�P[��/�
�#	S qU�\���fR�z9��H�q(�,�Pg
�~SA�$���_`�S����a��*������-[	�
�:����)	�\��¿֡W/�1�6l2N���!rt)�J@��\���5�Z;�?@]���Qi9&7��nAذ頨^
�2ĵ����O�I*�5<�j�D^A�e�l�]isy�砬��0���h�xW�\���z��ab̄82+�r'�|�Q,�Ph X��^��>�5�1YhHm��h�%!�Yw3�W�	E�����K=��鍢n�ꨲZ/�J=��b8��J���J��7g��u��G��W��Ɠ��F��;�F<���*/�ڪp��p�'�b�rft^ToH��X������4�p����p��7!�)��hK�:�ۓ��|j���h�D��J�� �R(K��m�)��Xc��=�	�,.*	Y_����o깉Q�.�u#��ʅ�ʥm34�������8���>���,	�?
Q�q�����0��	��!K�����h��7�vb��������חV�A� �E��':���)D��9,�����!�8XB�z(�Q�0�f�: �˔���p�F��Z��|Xc1 �-L">:H�)P��@蔃�glX�A �KF+	�X�@���XW^��z@ZH�;!�v���mWrђ�Q�=B��=��&�0�Ҝ��C�,�G �N�h%M9U@���rLP����0˳	zh�KQ���Cy ��uiV���|J���8�r�X��=�@nB�n����9Gl�~���Pb`�o)_���p��a��S0L̐�UY]�r��/��>�3*k�V�6��Q��1�v���T'	�@�";��ѵh�js^��yA~'�Aj�n1�p;�g��j����.���^��c5�c�k�J}���?/*֫	��U��قp����Q��@�Y��� p��(�h�th ݹ�SOh���c�3��G�ľ�~0sgH�^�v!]1�ob����
��/F�5�	ggWf��J�S	#:O�&��ĸ��I�S�Ix�$>Nv�jYa\<���,Yp�/���v.?�ˊ�(�e)�%'�o��H{W��ŏ�����*���u���	v��k�/���eg�I�W�O{��/0o�L�1~��w�=�_����w���|�'�$-D�3׸����� ��Fv	h*{iS�,m]+@�&؜?�`(���P��-�ri����w�>���.
�,@�8���񀜽��1?�]1⼧g �[hzf-W�9��2%�x/G�Z��mS=����\�=ɺ�<�I�z@#��u�yda�w�[<;X�&�l�����P�Q����)����Q{�H�K�(�k�
�f��-�rH<���݅�Z����O��B�l��(	�؆^�p P��}�\���-UE�t�9Phyr%_Z���A0�������R�A��zS&�'�o��@����eƁ�o�A��*
:����!(��G^O1���*��;�3	iU�~'��˃ͪ���
W�NG��Q���������p�3� ������<\� ��٘5[u���I�m�Ë���OB%:�m	�	u��^���������� �/��UR�B���xd<S�UӀXl?9��ZR��'Q��i�[���(����mO�P���t��*����O����Y�Q,� �5�W�	�n@|!/�F-����Ա��z�����h�'�-�f�Ϣ)�%*��Z��2�2bM_^�`Q�:�ǽ�Z0� ��}5%M;S@s���m����x�%��zY_�bh�A+�T}8�
P_!N��`'[�c�����(m���r_I���;�+
L6L��rB��PSG�j�<�G�FC�N祾FH��NQ+崲,	`w	~�B�ga*Nd1%,�RA�O렢M}�Ԁ�w(�|���I��u��B%`qV ��۽�w�T�,5�-.�-� �!�0+P	�H*	}u��.
��jb���@�'��u	���Ҡ $AN[%@��v�[��:] _3"�Nݵa ��a�hh�r3�V��"@4pݿ�����}�Sa:J龵Y:�C�	uNNh�!D������ �E�/r
��Є�%c�[���!�+	�̿Q�T!���k����]��0pC��x+���S�g�U\Mu�W��Rz�P჆0} �-�,^C�Z��qË3iG܈��O�.1�,o�^��/���ޭ�i��\e<�Xhja�	̜+���0W;&(���w΁
h�l�9$R)�^ʁ��oY!R���[�/_x ��@�W� �G)�5�Hw
��a�K��%Bz$ V���	�)ʟ`[�	[1�X�ݖ��p	b7�!�kY�8��A'�rp��1:�(>S��XQ(��a^{�f�~A���V��XOV��O�!>i�����v]�2��r��\Z|]��OR
�6��-xH�'8�������\�.�"?�w�H�Xu@1�;��@�w�;���������t�������#�-9J�p\^=�O>�!r�K��Q��% �3?���KR_z ���~Y��
�d��+�l�ųH4�����}[�|�H�B�X��{6^�__��U�%�H3�)GN]�A�z���r���o���)�.�I��)���`�Z(�,�� �E����%�j��VP�!/�	W2�����n��H�VO���w^����r�U"loSJB� ���4h	�	'�����z;�u"i_��_����qJW
�Lw�eA�c��>DY,NSz����=�j?m�90�?�i���^�^����2�����@� )�R�P9�C[��-|��V�ˣ��!I$��n�ܡ��:�[�>���(v��x�^6o6J'c�#<B����1��ڄ�x�픬�E	)�]VPG,L���x���0\�f:�����c-�� ����<HH7�e��
��ӹ	��]!�w�dR�Y�|�@��`�B�� <C J�ҹS4��%��`OI����h�9�7�1 �k[��} ���1�������<Ќ��&2Z�s"p���Ue��I�[3l*�'����f��oZ8�aU���w! eW��"
�'�����F�^��D�4��S�g�F����h�݁���b"|����!� �]�/w�OC��?���_�bEo�����逛�����X�>K<�-�֞�'��v�N�N�ʸ!~�r�t�%_}0��2'YZ�A��b�H�12�-�P�@���Qp������*4��C�̃W"���\���`cS�R�^c�� i�u�\L<P�gB��_�	!T�~w��g&�d��<��-Gy�E�=bN��֮��G���=��;O�5L����`Ӑ�T3�zF1Ld:�n�2P���8%jTp�#����5+�� M$��	�_�$B���ktB�,���'@L:W �Y�&陲Š[WѾ�5�>+b�ՋOU�FO�Yr�#�e飻�Tv9�p0�h*q�/�d2=U�K�T�x�2�xH Q�oR��P�	��rU��`%� CL'f����^��u4����p�\�?a�[�������f��4ʨ�����B�S��X-\Y�ApN��şq�X顷`�f1[�qs�����h:Q+�� ��p`�־��D������5fn1���s��l�~��-�!��Jy�α��,$�E{���F�I�ZT�k��:��ʄ��(A?SY�ޒw!�>�y#�w1���U��<!��l7�W8��s_���@t��P_�&�ZɆ���X���,S�{	=��M���b�݀rhs:'H]��^J�r#o0�	�����loz��ٜ�9!�9��]�"��Ȕ�#��U�ԕ��)o��a����<���7�
���`#�HTt���sJ��F{^��1��a�o �P/wyA3i�<́2IQ�#Z�p^�\�0!Qh	�m�2���H�oRv�|���Ȯ�0�u��@�S�#Q5�����0�5{�Q�� �dS	����|D��_	�B�U�V���hW#UYI�?�8���1��)�ps?S�@#��3�ҐG�N"���BSTЅ����X�{���h_z2$�Q�
�޺Yh�iH�?y�D�����H	�b Q�%��
�����f��h�8��u`��.(���p����c�j�<
%�`�)Ǖ��U�	��������B<�|<kpL�v<��C��\��Ơ9BQU�M)��<	7Օ�CL�8Z��T�F1yN/1��|z����}��M}�OI�`�"�Ț�37[���J+��em���_� U�?��<�8���m� ��(J�M�S�Q�t�O��u~jTq.˓-'������P�2�n��i]x�Y��N�C�HW]y��!آn%]�M�2�
���X�� d�!�1�-yH+rR�H��{�~s�+��6S��c(T}c�L:b ��] �!O�KF\w"��$ hF#�A�i%4w�/\��PK����7��/����B�[B��%�`���,�⌓<���k^�a�U:�v��f`Z�?EB�ם��/ ��l� Z��1�̄F0�?�j�`L�k�� ���&ZO)Һ����U�~���%k!��L*O�Nǜ�����}���k�#:F= me�)�~��@\�U?jA�ks!�`fy_6���9�`G��s0��*������������w�-Ҳ��RT���ykq6C!�f�m��d�>��k�ZVO�����I�! +�^���-���ؗ��8j�gd��~ߎV��Q�m5���6��=�A���`rM��	��}}�¦hXYz�p'@��Jdz_��:�����O����2&�<F�q3�J�`�k��/��V�I�/��T4���#���$4q[��h	�$@�oZ�xkN��CxB�N&���&DC�����!l���D��,,��ص�M,K��e�`P陧��5�
����.�:���]�-�hO���K��EI�-~YXQ�aj�B���?ӻ#{�H���f��e`t��	E��c�'�����'�q�iy��P��bC$e�x�%>���V�Pp�f��0�C�z��|��5:�*�ܷO	%q��]���[�Ұ�>��wY?���S����{�2[��~(�ć��˱�j���`�H�y[��q����K������-�L=�LfH#~PZ��GL�f�a61hcp���.-ә���ҁ��A�f`.@�x_ �)���[@��&�~(�w(����P�	�b r�Q���*���='�,�@�Ԁ[�^����G��tZA�.���-;��9�XRZ��b_��FQ����X� _��S�v�X�O�[�Z�	�l�q��s��n	��<A�*�*0�R� �̗��n��f���(��aZ���^���ʛ�T�(�Ó��Խ�r �z-�чP��fQ\�B�(d@��UZ�l��&K۠^��<��[-�N�U��*�M��]��G2��)��!�[1\�1
��@�(�	Wg!`U� ��o��9��du��Nl>Z�[q�K_�,�h�=Y^�-�A�Zݒz������ �a��B���N(R�-r�t=���Yu�����- ��Iz�s�IVF~r��^U��fhM7{�=����k�c���
�O���zr ����զ�~C¢�/��u n�`}NK��;�	�"n5����4K���z�>�T��E�r#�r
8� �h��qO�0���!jOxbLy#�<�=�c���.�!N.f(���q	N��� h�D�0[���vM��E~jSѶ�a4H�����2	�W�U��m�a�+30)���y���*�m�190Ts�B�A��!�'���	xt�/�w��5�����%�'_ECb"z�,%@��80�PACJT��U|��d3eJ`ʲ�r��;����	��_a�[�P�S�
�����N���"�4�-a�R�Q���MQ�y<q/ �=�� JA�AD�]��^��8��L���y	ȃ�/[��m��	<h�Y_e��J��{�W]VƂy7W����!�@d~���3x���,vM���G�k�v�������0 ���İ�N����)Z�����/[R�T�]��b�X���n��X��,1Ws�� ���gc~�Q�F4�ʾ��A?�=#4l����~׺9PS1�B!�1�h��XBv]�|Ўpl+5x	s����Q�F)^��haK���cz\��~ �0*�W_�����W���9����EJU�+	W��D�J�g$$+�u ��{�°�����p�
��֣�%F+�Z���]���!P-\��j�1q��t����ѿx*���+�Ǣ���Yhx��	����ʜ��Xi�}�w��@}-�96�'�)���R�SN?�2�5�h�A'Eu��¬a�P�줝}�R]:���g>�E�X-\�:������LN3'0�z�%~X��òYXW��bA�1(�u����'̥W $)�ob��<}g�&ٯ�Y��H-	�zC���C(>�r�_:Wg��0H.
(-H�W^������{�r���8(WFl��5a�f,XsIw��<��n���A+puR�L_�%~�a�
�[;�/�A�~_\6R,TZYى�h�d'En�И�V�vI��[�)�?��R{}T�x�)����G���>@������7(�튇�(!��ou��Z�CM��Ŝ����0{�����Q��Qū=qc^�U!د�0\�xt��_��|�"���b|��J��$Ҧ������x>����G;���Z��`�r,u źS}����+&P������_�j-0/Z3�z>�B��������w&o9���E�����^G��͍�3�8�x�/��#k]��	����kb��W��3�9h�d��-�+��k�����tc�8��SR�^e�,���]�	�1�)N��
_��8&=W��]
�����۸.��pտ�oA��O� Rd{6{mS���yWa��(�@�	
5���t;r8z	d%�'U��蚢�W��Gx�����/�yWrU���?	�_u�,�z����[�+ J�ם��b�%����Ɲ�4]T*V$#^	]yC�S�yƂ�	w���Hl����\d/Ró�w��F��0��dv�z�-:iV���nެ�M�6�4�ئF��~@v`��M �F�Z���G��
J�u�%��)� 1�$|+@�U�,K����T��~� t�C��D
HV *b�'O��0E�����2���yXm�j(kr1�$��Yv.P�G]�f�{�m��v������2���F���bO_������׋?�o?��;	lP߱�X*�k��T�� V�YSDs���b�I0�ھ>�'V�{ uTS�<1��0/@�pZ`NRq:}�]��N�7��+�� üP��1˿�X�Þ^�VM�1H�Ĝ1�)��M�I���o��Woe�Y�j͹�i��qG�.�b}B������P�S9��1 �����!��3W@]�؜�>�V�-�
!�F��u�Y�H%�)ny�J��@����#�>�ʧ�^�^S���HA@�C�$����X�4?��3N�x�nW\�w�vg&��Rq�40̪��0\���P����9*���<�0��i�݀�5*�d���~%�G�Ӟ �������%MyD��`���	�N���J�X#n�x�p�����]���U�R�0?Z�[���  �^+���]L�À�?}@q �f����U�Ԗ5B)�]��b�?���
�	��_�l�=}��	�I�ۋS_����`���0?�p_�԰YW�-I	������V���0�`��,6^f��qs?~�p{�"^��E���h�^U����Ż�S�u��`���-N�^��na]	�~�|<	��X��	&���e�>N�e���!'��`M�0�(-�%�X���6'�ۅ����B'g^���]R�����Z�l�D@��bŘ�Aa���Hz�U ���%Չ���`S]/rP3�|(qC�����-	E����D�Y���]s֪��$������]�k��={��4;򑗫/EJ0U[U��a܋F�|��g���+[8��8�;c>�^�b����h`up������>�y$_m�Nh�:�G����A������p��A�2\x1�DuW��@R	h�3�(B'��@��_ 	D5��o���%�:�ۅr����o�1��4Ԅhw!�
fk��������\���E?���z�y�wu\}�͈�Y��Zs����R|��S�h�Ӑ�_�������RB6�+�>[�{��d��;�T~"���̙��W�S�!���*S	�+�)�}}5	���Y��ƽ����R%A�V/�EX-�u' `C�vX颧�ؘ�	��wuF����,fZZś}TN��4��Δ�=t�/�� {
��z�CHP�h���z����C7����hM/v8`���Xq��2A)�� @!�	D8=�dJ( 2�]�߀P����
���}{s�iz����b�.�0����]:� ���6�1�M�VLJ��[H��e[���hws�V�0Sb�(G��h|WF\�F�H'_U�ag<h%}T�d4OX!����S��p��2 ���1��(���x?B)�R�2tʼ�Uw]}X_dK��qN-l��ѐ5]XEtA�@�"��;d|v����`sL�+��/�p|��> z�y[�~o%�8B9uQc���o���K��W	0O��{�(�� �(-�"ߨ�.)��Ք�*z@�����vf�d`Ǐ�'� �? V�`4m)�^��k"I�p�P�ژ/��}c,V[`��0�:%�X{��w��S�a-4Y��M�
��OC�
_:,��d��H�����r��E�X������J p3+q^
o"�P�a�����ׇ��(n��Һp��3��D1��d���W�A���+x�ٲ�9����n�q��@796~U1J�Дt��
 �w:o��4u���{��w���N~�8X��]S��#i�g�xm�U��Y��]/����U��-� _H�Z)�-r�k �Wh�v��l_&�J�z<��2�:y0|� 1��׀<>Y�}��Q��i���o	��w��\�>�/��]�a��K?��A�#	�GH@����0��w�$��)@�)1(����h�h?�>mʤ�60�v�5)��L��WUF +�x	AY�)
K%�X�A+Q~h-�7|�P��0e>1DJ�(�^��P/��<eW�������A1�T
��f�K�h���|$�AM���LP�/�X��p]� ��������t�W(�O ������/�N 2^ZY��B@)����_!�]Y?l�y
)o Jb�C^h�Dm(ZS��&�k�m�{�|��L}�w��NN�����&�K@�Rh�� 0]W�sTJ.!�_C2
 ���U���e���������&�^|u	"0�߹�X�vRsVA�/�h�ł"+yWQ���j�ޓ�788m#u�����"��j�Θj�p�|�o��*�AS�9�2;ԡ �3[S���&-z������J���S�y_반�Z��L�6j���*�<Q]����9E���H��D3�$h����&(�D|�q<�xX]��UD_hQ��6�	���
�R)�Y��n���l �[h��ST��v���������r���_x�bE����Q�?�p�UO�,����i� }�#��"�_�(tL��AX`9��GE4�@%�d�b i�15�;�<��!��4I�Î&6��Rw�cv�0=�K9�d�N�Z�;d�HlH�8�$��<]'4	]M��_,��a�%*Z��8ڇO��0#�F������rRQ�h�)�^�;�1QL�$YO���;�����z�<��-��dF%�'~õ�����x��j�.s=���Pv~��i��k)��è�ф��,���`b�9j�^ �YhCcw���%`_��T3h�s�X0$�������n�W����|E
�VO�v� ��!f2 -����%�`go�	F}������Gj�'�nK\a�p�p��L]j��$1��Azű����h>> 3��b.0�|R�6�i����>p��O���V�.q�0Z^�҂��d�� �T:��Pq;�]06��B͕*���%��d^�(.�;^Rq�c{��+o�v�K��X{�ā:0$t*�?��@ b����}`R��P������Ӟn��(���n
��K�T�	�)�L-���T�}��(�_d�K4���;�ª5w���]��b��@��h���H�oc�W�M-O2E�T�#�]���e���	�A1��-DR�n{'%)�_������l~H1������X��r+�k 
�X�X0"���`�!�01۪�OԘw�J�¶S�q���|Ix�'����B�^�-�5q;���@��[�}��s �fV��
���b2���M/Ɯ< |�Z[�б�M+A���b�;�]���>",73,t9\O-�@N-�W:�҅@����ۨ!��6>��
�9zԜȒ��sC��n���\��r���[
��{B��+�x*�\�i�+b��< -975x�-�I��_��š�쇦��`IH�kY%cyu�����~���0;3K#���5	�\]�I�X�{�h)H;\�鵔f��W`�f�Ǝ��8ʇ�D��Rx2sv�zc�ݡ1����O�D��Ll��؂�)ˀ�4^@����w�K>��P�`��e
��z?f�pPW�~�_tZ@|�����{Z�D��{`<-1sf_)�'K��S������a0����R�xֽ�s���z�&k������aO0���0��b���{
��dR����M�&�� Z��z:,��})�W�bu[� ��I<	����JH��@�Io+	����2��T| �]LleaB*�S����^P�w`'���z2�P�B�ǃ ��d�Hh'�M�O�Y;�bI��
uVH��@��2`AUB�[@��5/�{Z���_	�*�x�������<���A#��§����9���H�!�%��Z�?/�\��w�
��j�~O.X�%~�m  CU}�`XT=�~�%K��Pܗ��b3U�@��7��1�9Y�8���g��h��PˉJ;�N�
�P06B'(8�\ϙ���H�,�@1��,`�.���A:��P�x9���r� [Ĥ(����f Z�E����N$��U郁	l�|[OW�C@��`������Ŧ.�s�6?uTW@��nI�E��X��=>�=�b��b�	(�%��3R�v5�-����<�3j��ɀ����x�,����hv��5�K��у�1v؟JL����	 
Q����.����V���A�'ׂ�^����.1N*/]�9�{��@�1M:P�q�y�'u�I2}�h���Q� QO�G�<P�Q�@E
����7�#1��_�ޯ��G���ZY��&�@~P�X)l� �1�_o{>~K�(��L*vr��2;~Y�t�\,̘�*TE�a@����R+�}n��0')ч溠k�-B�T�M�F!��N�j��St�ZH_�C^1�	�@�u|M'骄�!�dT����o��ב��j�T*���Y 2X���������Q�� [��Rxt���A�k��äN�8C������1���K�+.�(6O�a�^��/Վ�����D�6"�w���0��K�������<�0)�x �Z�Yhvw��"o��C��_+̪�-�:Wx�l�A��2X�'���y����W؍l_<f�H���h
_F��f����Q��:�m/f���稞�
���W����H��L�+��	ԍ䓅���nɓ���������D�G+Q)(�[�3�2�@�fSP�<$����㿘�4È�X(�ܻ[���ج[�Z�}	��M�h�Z����q�Zhо>��u�<
Xh�B�+�*z\Q%Z^F@��}����7�RA���H-$�E���
����_aL!�:h*�Uf ����R�# (�Z�݀�s���	���YݣJ7PV��R�	�:�(��� ^�T]����yA�����ݸ���d���������� �P�(ȝ"�NbCh��ݝ^���@�"����"�����g7c�� 8XZfQ�� v˾r`�A�}�-t^'�6iӱ�RT!^�0+��	�`���_&J1��>7u�Nθ�x�y'�(@�WYr�4bJ�堊�#1�[��Lr �p�b�F=����y 5��o��(!��'�}�,vDcN���������myk1�鈥 �R�-S�
!���qh�}��`�d�[�IY+/�h;]`����v��e�z��)�o�.�8%�u�P�ԓ�Fy"� �c��
�� ��6��p��ۋ/~��(A��`�h�
;^���O��^Ĥ�����E��f�XnYh4	R]Ct�($�M�͍r`�~�s�QbDÿI�a��SE�	��~��I04O��jO'g���/)���E15!^�XLK�O�o�0J�M)݄��	�loJ��H1�t-���� �[�CZ��q=.�UA��:��b5�`6M������鯥r&��ɗ3~�)�&�K�Vq���*��d0�4Cl	����
�b�c�/Y3j�V�r�_�OrS�,��1��G�Yߠ���-�ߖ���Wa�lf�A�u�EI5��A`Lf�D@�z�� �0�P�"�X�Wm�Ph=)�w�Q-�w�RIp5��q@��SR'[Zp�5h�r�Q+TS���j뤀T/`'TCb����b�Oh�$����(����)y�vT���0pX1�[�Uդ�F@m<_;[1`N.un��,\@�X
rP��v��!��)@R��{@`0����o�����$�O��Fo��1Z��qfp�TP>��$/AYW l�Hb���8*T3��+_
����u�� 6Q��/�Zo��~{(ب�wTP4��9*V�j��_����r#)-���y%հ��%�vG���3�%��:]|��\ƀ�#?�51�]�j�'hRo�ܪ��^�����ź��8� h�P-��)�/_�8��6=���ӯ��O4&��o�a��B�R@Ј�F�[��eI��?S��������fP�(��XQ��鄼N�\+�yV�̆���`�V5p��N�B�ݽ�Y- ���j����
�"���/VNR�{����5Z��7ZJ\s:��*�Z߸)���"o�3���M��)J���_!�^����1nq��p�-(;���O)]%UPFZr��
1���s9�X��g�^Q;i���A-9�)й2I�<V� |g�e�@J��h.NQ����r9o"B�tU�������G,HJ��h���Be^��~=�.�J�;�,O��0	�mX�[T�0�-Zu�Jq+���"�X@�6� �-�#��*�Q(�<����X��5 �f�a��UeL-� �'mK��|�����RY���!^%W��<V]1�w)ᐚ�x'(hRK����"�8.�胋2�`�
v�Z���؟83�D9��C�54$��F�Cp�b9^؀��^�L\���-��5W�����Z]�5��O��4�+��c��5��#� 9� �r1w^Q�5d���<J�݊06�K��GJ��R9�^��ov-�,j�}�hJQ���$�U�9B)TZ�48��a�Z ���� �,v(��h-TG���(1���Q��;�"���E=p�F	5��F,�%��.������o;ʒX�A��zM��w������̎��0�Z����!��	�uَA��*�{hO��U[Z��hs��-dM'�_�@����j�h*	�NJ��t,.up�Z�	�Y�)h
0Q�[��/>�-��A��ipn�9�����	�  ��pv0�������ꦉ�o>�ڹ�)��A	�{�ã��BK�&y�o
���_G7��/�{ �~`U�R�W|�`�s�\^1���Y?!pK^_
������?����!�R�2����u������Y�Q(���ǘ�+0�� ������!��M�%��ܔ��a��
`��4����V�p"����X�\�\�t�$�l��*3r�Xu�4jAn._5h~��9o�
^�|��	�=����w¿��0���O����g�#2X�Mw�P,z1'a\�
 ������t����X��Z \��;e�T�pL҈���j`g9(� �.�p��0ü��]��n��h,�OHc�'r��,��r�5�IN�ؽ���k����@�W��P_�!�^�g˞�
�
�͉Rޯ��2p
�vI�����m��1�p��9�G"%��V$/ݗC-@)7�aR8��Q.¢	*�l�ح�^_�ݜ���Iu��3Y�`���l}����P��[CJ0�����9jA�����������żi����?�W;�� b1��Yb�x,w�X_����j�#�a�&PK���G��H,D\�{�y�(��Q�18� .bG~P��fm^���\�`*�E�$��'�����B���XL�	�{�Ƚ��mW��OdI1 ���N��t	�i�X%(ڳ�OY�*��E�]Q���V@T������fY�4BKq�@��!�N��1�	�f��l@��o/��e""Y���|fh���#�,J���
K������ �YJ�i�	 ���-�TJ�b������V��v�DE�r�Q_VH`>K�y���h�,@K��)r�c��(�a1k,X�B�/�½���i�Iѫ FO:�UX1��%�
h�?w<('L�~?Q��C���l�`*�U�+!�^�Mdz|�!�\����>=��s��V.��/�Y�6}��!oA��E{��<o
]�z\)C��(�a�Џ'�^B��~�k�`����ZlvA��cPI G�f �)�%Td��SU�MXf;/�Z[�m(-���a:C�:���+)�@��nz#��A�}�x���p����>�Lk	gT`������C�Y��MK�YT@�t3���
��9�251nz�%�jh~�fz�v��j�������f_�\��[�,u���A���P&N�ʁ�]T�ܶȐ��&̤M��a�u�����t~1ɽ�c&i�0���fBIr�29A��Ď�(6JX�YZ�ct�<� \�)�n�|�\��iu��X� �\1����HY��<�s�h�������1X,콠��i��_�E�^AT8��O<VL��PZ�	�aYFR|&���[�z�e6Pl`�o�$m�1��<�=�T��xʙ�	(+�eLƇ&��+-�α@�1���({�` ��
0@!_���TQ��?~R�XTۄ~Ä�4�`B#���M/h|�b�Ğ`y���9�J�8f�<��A)B2�]��@(��B	���P�+Q��;�*,li�{�A��*��BY� ��!�S���E$��
�藥�|O�2V�<_B�b`y�ZQP#�ݐ���/�^�c}�cx[�*_!�fN�$x/�,7�ˈiV� 7�۸mk"�A�@��l- �|	�5P
+��B�WJA`�ϕX�3)�`��Q H ���PRY)»�(0[��:/�ZÑ�NQ�>��~�ց���n!�(r�B��؂�ཋ}�����<֟�?K���_t=']輡z-&syu�Q�v{�i��=p%�l�R���t?�Z��;_�(� �[��ku�ߖFN��Q�
���yv��
�4+MZ>��C��Y��7�mV:�5�$��U�s�)@oY�A��?���ª;��%�	3hX�.[Δ��VK�/K��
3��K}!��$*�XY��'.X�=^�༉���(V��Z��(y�'ڑ/_�E�Q�g��i� ��0<s����o�^���� `����1�?�l���Ĕ�y7W�����R�)Oc"A����H��0�d���p�
@�hRBc�=�ټ��@Gw�#�ՠ`	�P�|Z&��,�Hs�W1 ���`~��o����c�X��
�!p��O�$|��~h�I�z4��Nޏ&����_5D)ى}�TY�k���Fc\�qޛ �,x�b�(G4�a[t0J&ˍ��q_`�%�u�b	��z�%��IR;�/�p�X�]6%}޳/�}(Ђ��m|�-�@�is�Z��	4)	�5�h��Q�o;�RV��c{�:��I�A�hE_4��xp6�}�8���X�}-T�����U�8~	[�hɰ8�J��:��25�9w+ �[{��%�V��H0�U�K�Sw3�f	�j��rKQ�Y	���P��p�,U�y R.�#�bX$[Pٱ ���lGh@G�HRlZ����o>�ۘ�\~'�v �|Lי����B�?}�7�#l���n	3o^}�7.�l���N���G�>��H\��7<�����]-U9y�|���� mBr������?.�`��0Y������Ҁ�!�)R�Ԗ�D�Z�
�!��)��v��@,\_yAi%���,�1/�H*�:ej
�P-�#i�%ߗ�;,�#		��̝��	.�a�� C�/LzW�odG��a��;,$p9F�1(��Œ���e��I����$�c3|�п0tW$��/q<osrNJ��#R�r(�Y,?�}�?�k�'5�C��5G��`�gQ5�n�liX �
Zh�[x�I}衠\�_,!�^��PZ�1� ��@\�E��V��Kp�ut�A`�s�f!hÉ0�a3�A��hEʾ���-���)���_����fFj1y�bk�:] LƏ*��[����Miv���	�y��~�bYwQ�Z�	��TΥ
����4�!��;�^�-T0PW�]��HAU �ͮo�M��9�� ��8�B5�V�a�L詘ME�9^� ���-`�顨���EF�#�
���~�r��	�J��q�~�=�Z�����L]����#��'r!| l	*�p������wǫ0�t����qY��,M�6�*b�2�*�h+ʈ���@����H�[��/�N�
����bK������Ph&[�Q�0J��O�!��DQ����Y(�X�р���;s�(�(%=J�"1�-/�t�VU�F8�xa�>��'��R��n1�a����}����!�����/�I�x�R��ʍ������P+a���
1͚���~f2[^¢F�0J�����ʹbC*��Q	e�U�u�'�����t��SNY���g�,�L�,R�l[��-�OϽ�ǒ�=6�p�	I{~[�����Ju@�e���p���^OJ�ן�)W�	cK�'���p IF
/h��T�M�
�V�����1����`i@�����ї����ը0&V(�n"`.��/�I�v
O{��h'wF���8� } E�@V�Zc���_��-I���������V�Q�;^�<�����(ث�~[��_9ƭ�]�D�^��S�vV�c����Zy;^ ����"���W��W) �2&�����C�7�����$���ݹ{8+�K,��<��o8U~]s 2.yZ)߽	7d�%p�}�X^A��7�G#`!��g�=�w�������OoBlCa�����X�e 3
Z� P�EV���	h��)A�I�2T�f�aO]�x�� 
gXH� 
�sU��\L��Q%8X�g !8b%F1]�.�3R=k,>hGc�5�Ja�Ժ�w)*4��Եx"�Pʙ�;0���v�\R�5�K��`"h8ba�*��'sO�FL�[�(zz���4�X����.��	PUk�������-T�h6�W��p~��O\�=w�:�D��O~��ą�(�YV�$ګ�w<���	u�Xv�k�/�hE�T{6�}�u��PPHZ�� �)8c"���W���x������p�\F	7�GLA��O-����?	�F���5D4u���p#Y/�Hh�O."⸏R�!���O:�R�=���-P��YS&�@�sz"`B2�:���`?��,`J,<I&U��n6�1%)���$�I���D˽�SV��*	(9����I�ƙP�R� !=�J�s�]V	��kB1�`�3Z�/�@��_
�v��A�*�I+T���b�A��KsՒ uƿ5F��W��df�쉂���Ʌ�>Rr�*v�[�P��[�g���3�;@�)����,X9.,�}\�{����,�Xҹ��0�]�MU;h�F�")_!�W��;O�+�N�����ܻ��0
� ��)ݾ�X��	��T��AI����,N<��q���|3�N���3(J��������U2,!�<+����h���@���FRh@	Z1V���Oa�#�N���%Ձ��]D��g~0ν��n\p���A�}`:�r0I�V�b|J&B����_^ �K	|1�T�d["�]��Ij�/
i��'�I�b�����Z)�_s��v�k	0��1���ِ�G�-�Dq.|��Q�R��� �iY?�O���x�݌�Q)H�p�R�t�7:0����b���<�
��yN���k�,�U�U�
!Х�@���,f�$&|S�k��+�,K)�hTx|�I�懿TR��-Y>��dl��X����J��X��	�.��1�`�~�`,���5��>\�%�<%��V&�d�(\�o/�co �5~|UX��h�xK��E@�rj��y	 &3Pɀ�y�q�tfH�����W���(:�=* [9��J͸���&���
Z𸹒�l��%�'��OV�����h;�!K����2h)���l���G�8��k�(ߘ:�&i��1�x�<�A��1
Zܹ����h�J]@Y_I�$��$�I�W!F���\I��L'�]RW�
\��]d׬�X� ��T��)Z��2`�LP�I	�w�	Q�r=}����Xp�1�<�#CHv#>�G�O�}�IW����������0�������U���3�N���e�<���2�h�� ��V���I%�Y�� E�[�m.�1��W��2�%�q/�8C��
���՟����og
1h�	D��	QT܆�Jz���,��Hվ`-:X�3	_a�� ���J� �;/)�-�Zj�9�p��[&M�G�{�_ȣ>�|����311�>l�KC#�Y�����D�¤���e}�Y�6Z �E=� @-�W%�N�15"If{@�-`)���Ȋ
[hD;̚%����@�R)bf�-fݟ���PCS���J0�mc5!K&����'�|���%~ޞ�h6	+4�������f�-�
��P�(!� 40e��Y3�ל�?PS�@X�+��#����Á�YX�\�E�kh�_Y|�' �m��X6�0����?v���1�!���A�s4�D�/�]�E��"}d���1	�H�zx���a��
	)MZ�~N�l�8I�Z����I I��"�x�g���C���Xoj 'e)�]�A�������L 5�<��)72�����4�R`��	�'��Q�������>�R⩁�m�!;�$�aF���IA���N�(b�F/�ˊ7.j1o��)�������K��0z
T�y�W���	�#!)� 1�����\�5�.�l7}��`�d�z Y��-_\��%�cd�=���-$|Ϙ"?�/��)�b�L@+?��I��<��`l�`G)ME�I�Z��C��؍ p�I�	hfW��sSJ��0���A�u~�	��m�z bv�T��� ��@$5��uO|E���Ȥ���ՀPhzF +X5A.#;�/Y+xY=L��jx@uB<w�x�����YJrFP���}8@)��]*���&hX-yQ ��n{O�	:����'?0fQ�r�R
�U	�t'��Y��j�
�Bk��EEZI$�P��)�u�o�h�L���(�	��]d�HT�d�/x�EQ����fWB��4� P��D�h��C!1�)���`Z��z�9g�r�D�������%���d�Ld:-&��
�� I��Z�����B�[��q��i8�'�O	�31��Fh��|C`�@��m`K�5&_}wu0��B�?e�����?P�(Np�QP ��k	!�� wf�5�q����ls(���0	��Y S�G�K}�K����{&Bw�7�����ȗ[�' 8��;'^k��H��)_���eD� 
M���* ��|�y%Y��Rw��T���k�gV���P��[�@z���s�qV�R� ��P?��Ýk�>ޗ���S��ضc(���[�ހ� �_��]p���|����U%N~(w4�1;�q׻r�u1df���^k(��Ҕ�_��U�3��C��\�E [h��`���Ʒ0�
FQ������<��o�c�~}X�,���YF<8�rV��X/_]�� �]
[��Y��&�+�3�Z��vY���&C�J����,�[w���Hh�>��!���/ݑ��o��%�vv�Ws�\n� d&zD��M�E��V1�n:�	X{�.K� 1v�h�K�v�bO1�ي�%Kɂ�V������}L:v)�R�H�QR���_�^�������B�(��i�4���d,^U����e'RT���G#
�E-���Q�����i�I��Q�8�Wԣh�o�T^�=-CݪZ�����N� g��;��Œ���iv�Q{�W�� ��$��8\K�^� �%��WiYA�=_q���0�m���q(��<�ʽ�Z�/����B@fh� ���m�b�G!�d������f*I\g��[Rh�Ta�˕XD(�f6����A(�ȕZ:�z||:�x���1��g]�I�V�.S�r��wY1�dg
^��2<�Q좝@b�r��,�F�v��ؘ�	� X�gf+q�(��A�����*VN�*��Τ��<�{���7�#]4������e?/1Fb�@����]\��:+���\�c��a��(�;���_�[��Bp��Q]�%��^H.��Tfn��;�ۚ,��6�y.c/��%��^PJJ�ι�A�"�{��?Ԗ�J�@���<�)�h�t��rJ�������w/Fޕ`B�g��-�籦N� �4*�����f��q�R�;2r���G�q��)͠�R�VeP��&6Zb��`H��&j�ܖ� RsU�rq'�]�鄿 �R�@(��p��
U�^�a��5��~�}wX��f��."�-We��֓h��^�ߨ�h�`��s�*A��qL6+�e¹HhT R�C#j���@��}@���;�N� 7Dl_G�l��c-u�
�G)�ZS��#�N:V�?��q]���D�e������-��>ʓb \���s}�����5�%L{.�c�U�Bf? �Y���� �#Vh`���LU9Lw�k��R�Q����kE��r���� �<T��Z��C���������'�z{�:�؞z�@T�O�d?̚��_���\rO Z�P�^0!�"��L~"$S
2}� ��t�1�]�w,���/ ��'�NI��E��/w�?X�Ŗ@W<˘<��+�����qK;�n~lf�8d�L�7Y
Fj_�	��>� &�En��<�w�w��{)���S�1� _l:�a�Ɲ�	@��@5(�%�Y9
궖}��m\-��1�����YV� ]�#/��z����o���?�Y-�8�B@�ė/�V��|\i@Z]��'����,p�W� L*N[X  hFYZƈ	A�;�:�/VV2i�?�5��D�#@|�;�������Q�@ �Y�(HD�y�dJk�&I�) |�0cH8b�m[U\ee���Ã�>��z��>q~-7�	
y )��̳���+&�/<SY1�`LG��Z	 i،�\C&pl���������� �Z�"�DK�ɬ���KV�Þ�4��f�9H�P�1�)��=��x��0�Q�z�Nݴ%j1��5]�/�bo�&�R}�2l�h���$w�,� 1��x�-I)U�'�RhDL�3�����꘸	F�y�[鈧P��>C%��� BƗ����B{_�e�(V����h)��1�No��0�n�Jy�;�	k>gu�x����1u!����~a�Lh�Y����Bj# H5-9-7��_�r-�����S�<���:���
�`*�ړ���"r2'������
�\@uf��vQ(��)��j���v�!��'A����qW��	�j��
_�\��m��\�v�K !�m2;�Jts��J}\�Xx�ky����0%�(�T�0��Xu���%	���25,8��B��N���0��@�b;�M������hk��k_6�aD�	���|ؒ�@� �������#�������~�.eEd@z�՟r���}>\K��<q�V�Hp�������dp��r3�\-P���@,�w�׈"%�!a:�kh"��L.<!)�f�^'u���otJ��`�z��m�K)��lBp�{����� D�^f�ȸ?@~}�Q���.Z�ͨ2/U�[�\ ��� i����ʍ��e�4�&��o)��T'���d"iw^�s�򸥥,�k �cVP��v� �T"@ wZ!�`閔���C�4��pх�o��� �I!p�3Z���tA�����7B���W����Z�� ��L�KFI.���șw�4I���SX��W_	] ���n�}1��5�^Ҡ[R�j�%WU]�R��x�����������ȥ��fX]����"��b�i�ݠ�a�tPZ���<����U�'��ơ�u���)��EaR! wV� �+��^����B��u�P&M9�&O	��y����}�q[���h�IU �B@�FC��>oJw�k& : 5LS#�k�u-�+��1���r�]5�L~RZ��fYXx?_�P1�L����)�}Xe{�)Yf�Y�i�Z�ٍAU���L��e/���SC�J[���g&�0�e �v1HO�^�a��6T�[�J�2�Y�\~��Y�v� ��8Xl����.��}1�]
1�`@����<MV��-���R3/Ѽ�/�f�At@fiG�N�4@��\'�V��������U O�0�R��&n
Ѽ��� �)��6��顔U�}Q�z�H���A�Yq+L`�a�X iD����)r�A�Ph:�12u��<�귑!��8NdQ�k�ד��7��<P��~�,���;kqU��0]�Ȧ	��co;~@tN����M^�-��R�O0��j�k�{
�o�
�ڦ6���"�?	�I�	�<���
1���@!�[�:�aXşD��	�q}��/[0S�����{����.�<e�8)����HV��5�	�*K��
2WZ�)�݁���I ��^U�ci���m
��/���d31�Yӆ��:c����p��i� �}VtH��5���`�3b|7��5sq6W�h�9ݎQa�1�)�S�	����xV���?fB!Ÿ1��б��¶7
 �!C{L�����X��h����yj�Q�iWю�����ϴ6ʆ�������K�B�Ƶ\�B��W^��dΫ�-~�ƾ��0�-��\��#4o�oA�/F�J�)�X!�U�Bx�ܡ���g���Θ��[Lt��?Nԩ����A.���^����������Rs't����o ���Yc�`L&j,?p� )PhW��`s��dk
)���p�����=� G�vhѵҥl�691���BH���o�.��	��/����c�WqQPbZ�?MEkfk���W�
S�BK�L��a�߅�z݃�MI���gź�jPF��/���6.4�!X⤐�A�6�L�y�E	Q�>�L�8��ea��}=(��_���eC�� }Q@��S0�.��`c�0�H#@
K6���rm1Q*iT�I>��W+�B�_!�B�w>x���K��tĚX�pq/5���ǘI\xI�� /�-wWS�_�mIyu������W}�"^��d:���YQT�9s�w�ȯ9�a�@>�;�LClb�'i�^	�HBDӅ����	A�ڌ�d��Q�(_�BMXE=o˻���'1#��[�ji�Ҭ���'!�h��ָgM-7%�� >���H<!ntk� ��fdXy�	`~ >�!���:�)�Zt'���z�<�M�Uݎ�
�dI����,�U�WB��eX�_.�61sBf�;���̻p'�P�	���]��w��'j�\&���@$H�B)h� 0_7�HJ�2閐���\dM�McQ�~�饫Ŭg��kj�A���6�cǤ����:-Y?jO��U2%�bZ_K,���ɤ����~<�c��>H��q
�G.�;$j ։�)��
���hT�7�����2ua�]��x
����;��u8���2�p3 �fZ�h<p�<|f�V7�NK�I^�M7Q��>����_��.��~����	R'�G%���X��=�\��BH�z�>�-	C�å$)�_0J�,�}R��O�W�H8���mj>��!
V���
u���S�/��,���%�-���Hl�x`iIS������>�YpH��F<�h�E
^^� �!�Z���OK�Gh{�]l��0�_������z%�MZ�fP�ƈ˲X�/g(����?k-�]��C���U��pU���֖��IZ�)�k���1�1����3]��(b�ZY�g^F����Bib�]�X��o����	�e��
�Y���CC�n~3���X�r�^��$]�}$�J7>~��.�RȾ����c���Y@UTL5G"����zJ�@eUR�A 0$�'M&,)b�N�	�f�KZ��[p��J���@���S��M��G!�)�;���d�$�}+�#��O�8[��i����	Ih�D_ ��<1*,�%���	@�z9%Uk��/x��s�3Tv���qG U[�yQ���9	D	��P���V��0�� b��n%B�)P# �N�4@-lU�s[��)���oCN�(���xN<�_���;���ɮ�Zh�%$�^ɀn��T��F#���D��$�����6���s?A����q�|Hv� �"�a/!�*���	�L�|�Z��=%���y�L��+ ��AsM��Hs%Z�1$C�`-�3+ח�@$H0FQZ˞_�a��z��b�ov��P����=wy`��r�RIK��� �[$J�������w�r� 6U��C�s)���F^H�A�F��*k.f�A!���_�,��B��}�܃�[!�R����^�FN�xX')ez��c]Q@�1	�tu����T�����u2ˍL�n�^;ܘ�BV�h�@c`x^9IZBPz*HA �c�XB$hkgH��*��!�X�X��%Bl�1��z�ӯ�CE8Ole���'p(-����P��rcF�̐���� �O�^��m�\��Q��~]�d�}�jL+7�g��=ik�0~怙Q�<��:G�"CL�=�P �h��H)�|r_m��V�@��c���2��/}!���{�x����YxA��	m__�/ �<n�&X �5�r8}	1���P雜_1�?&�h�,�o���y�z0�@�?�@+�x�
� �������(�>��`J��ڰ|���ށ�cm%o���M�7"����-p
�}^��;�2/�'~d�1��O_�R���<�z�5���,���r�Mq�SZU�R.��2:���z�6GC�A�:�_��t1HXLU��L��ϓ��P �b}H.�6�J��%a�.o���h1yf1q��QQZ��J�[l�1�v�K�` X��h<! 7Y^�*f(�d��P.9/�-x��@�Q��]J�L��X^�+�ӄ��q)�@�z2�&ǹ�{7Gn1��%�;�;T^��m�Pv��`�	�T�c�y�@6S�� eIQ�8�+��ܽv�k���3�v[-D!%{; ���=)Vء��ԺS2���>��a^��0�%O��[�}F+��-�=6n}�{���������:ţ��{�y�X9���;���6���<GE=�*W��a*��Ci��L�;���8ol&�4��^�v�YO	�y��.���3u����M%su�֮�f�)��,O6�pR*���¨!����� �) !����HR�1���H/� Y�������#��N�S�N)����`y3�#����g��{Zt��d���ٻ4>$RM�6:�b��w,)4dP$��1�?�X�w.		~'�tbs�R����8��nz��_k�.q,�� h���M=�=,5��~E��jirn���@�$��\�\ ��)�gE�@��M!�6-)�v��2���$�a���@�4V%g�0��w��$1ŭ_lPb��>ZX/��ڒ��� ~D�8��eLGOE�lb�ʯA9_`��4�7�Z0$a�e�ܮ+'�(g��F`GgWG}�c��Ś<���XS��%3Ji���C*��4�?9�'�ײ�u�����P\��Faw���O.�(hX'�t�'��Ʃ_V�Cv����Z�w�w}�fX�����`Wn�h�zHX0��&����� �t��R*�t���*I�@Ap'����!Pv���p�	�&LkF� ���V��h1Q��@��nE'�b@��L
g A�Q�KR��Xzn���HJ��U�7��<�ʯ���X�XI|���h8�[O�p��M��K��P�QP{���7��
Zlq�}��V?`f��{�rX!�����ZW0��|� ��8]�� 'P>o�Uh�]`��';)�X�ʂ]�_�/_Eԁ��a(����'.�	�BF���i{)�^1���(���./�=@�	&�E3�X��4]2�A	��1�4�s.�:���+�e�r��D�!�+�0	�;��K�x���>$v>	��f�-V.}3�r�{��1YX���U��r3Jd����j��hzbr)}�MX��z�ӿt�������{P��0��}�&'%F�=�20G�tg�_@�[�P�a.�9!�M��z�JW*Q�Z���0[�y	��H\���\��#~	`Dנ��x�9���{.����6*��	hJuk���<�S�R��h�Ť�������@<[�6�F�놹_]OӲ6Ҿ��	�7Wʊׄ/�z�EH{C|�W��<�e��Wh*�r6����e�T�2w*���HY�W�A{�����1����ﷁ���8��_�	�����N���fS�J�����7P8��,���U��B�C��@��~%6V��*0Xr)���$p�X���,�̀P
�%��=��.4O� �����$��c�
w^\ra���퉈9�{*�h�S�U1
 ��F(؀,�,Z���HZ
��OHe�0I�5dH���@��Tu^y�H��P`VŮ2Kw�Y$
N�O��ð�HLJK�y�O�P�
-D4?�	�"	�W�!OWā��!�n�B{9��[�Zs�K<�w���
qh�@���7բ���``h�r{oY�)�9	l��Pq� N}R��a��1��7�ir	.(F|2F���Y�~��?_��Z&���|�{m-lM����0h�b�(=6Q�y�r`%O�n��K)32�L$5E�@�m��1'|�����^�����m[�C���c�_]�I��ҿ��B�+H1�0�=�eC�ث� !�ZRh��_^� �i�ۘ7��Z��u0e�Ds@�n���8�݋]X��b�N�<��kBZ�����w�� �n%U��B��\�nh������*�D� �Yt�l�� ���JN	q�۰�1�.t����I��\xѠ��2�R�`��tfh��J\^K
��s8�s>9\k,�0ʝ׼�����hn΅�bw�M���L
����iϩǵ:"�4�+�ܼ�~����Nj�Io���'U[���9$�E}r� 4նۃ
��pQ!w�%���>xZ���3'��A�-j�ixK�{�	�_fVVN��zHSX��F7];��ٯ��*�0��`K����Y���PX����X�lJ��7�?�� ډ���%΂2g��/'�9�M��J�H��M�WO��~J�!���=����(����!��hp�\d���/�����=�sm=�m|O�]ѭ���"\>J}�ڠ@ �	H1hZ���u���Gaht>�MX]1�(�|��^D�����W�a� �Ũׁh%84��,H��u�C��DU�4�Ƃ����	WӁ���i=� Y�!��^Ivj�P��������Ɋ��8d1���X@c+i�$)�h(|L����e��K�����s��� ~���F�w�2���^�xd�J� ��*p�[���Vu ��:fY�hw��~��w	���4�7��I!���h�Vӿ862�Q������r\P_�����ԅ�C�l5Bp�e�]9��C	�n91�0���F�	h�o�Q,�J�w.0"?[1�t�����G-aV�	0��jj� dT�*�OW�*�^���'^����a'��ɺ,!5�1 ��B��}�-PYx"�`��rc������]����e(ڈ$)���A�6����i@Cȕ\}���H�pXR�
�h.8�oO��[$����3��:��!ј7	&l��b'�{%�F	��@P��E�vr��ۉf �87�X)\�k� ��{f�S�"LՃ�.9��'�\���}�K;�~W�j�q���h�B#;YT�`��\%`/��!E �劀-B	�[[�B/�PK`
D��^���!��	馗-�q�׃~)��R�r�P�_�9y�71_�h�z/�`�kp��W��
��1Lz�:�qn��G	'�V�EZP��II��$MB�fRP�Eжb>��\���u0��8��F2�\Wxy}�߂n�6���k�PbºaoB����0X��F�G�78�	'�hN�AI]���d��j�ib�W����Rk-hWc�p��'���_jʘ�hR�	$��@�J}�bN&P�$k9��a1A4z�������K�[W �Z������n�rޝ����Ka��P��p�~�K��V��Z*W�o�c�J��G��sM���"�2�k -��ȹK'�)^D�n� ˮҡ�nAhtV1�opG�P�w��O��h�H���6�����Mr���v�V��4�� �۾V��Qh�Kl��-���~�p�G5-��%}�q[e��(��6n��V��0u�+��-�xc9��:�=Ȓ�M/�f�Мat�@��V$"bg5�F`-�Y1L�m3��Z�u?�c)���s�Œs�<���3F'D�����"5h4�%���M���I}�G���z�K�;��i�
�T �"V�	1��ra�(Z�*��wP�Y������m�����Zi7� ��s����mbi_���nC��O�w��g��� {�c��_���dEN	��]/�IK���������	�	w�A�:2�ğK\��˯̭ y�RY�	�ph�4<`@��J�i����l�	/�	�t�-|�zuHYZ� O
k�i}��
�z�6���	�1�r�/�
[ث?�z����pF8�)�s�#/sf lm��N�­�}Bw��&��r%�H�z�k��Q�����3t[>��xÐk�?&�`�w��d�2c��1�P��2�5��}�]v��t��5Orh���\/�?^��SV�b�s1>�u�
���A�)e�̽y/7�pa���}O�:�B�v!Pth鈹���T���q�0�[��S�ĳ��,�^�3���Z^UrVbPP�^ܾ�����ЁQ�����+�9E%�bp) :}��af�XA�[��x���1	rLݳ�(�Y��X@U�5I�	� ;-:
zH��M�;�y���5�X�9���S��B���c5P��W ?t��P��{'31�Ƶ�}N0�<N�`�kVze�GW�L�O�PN���)�>�Cz	:𗉂%w���A��ӭ�*`��ҏ���Ul��}��n��H�(.�;]V�i��}�T��!�]��"6(p@�XM�L�+37/�1cN_�����t���|�"-���B@��e�O����W���tO������	��W	e���\�d�(��I_G���W\��
B�N���A,���\gy??�^�?��
pB�F	V�� �.�S1�ʀ!4E�� �@�Y�����ufG�Q��РXGmZ�E�Ќ�#�^ŮZH�]��	&`��Lc��D�
��A��E@f͖K����d�>�!�T.��eո4>(�qq�V��dI�(��-�i���=(��������Ƃ���h k���R?���e��`�BKΩ�&����K]�;�C<N������t�:��h/��%;� �H �S�o���O���!�����_����0QZ��x�8�p,ϩ�p�<8'W\�h�t@$��Q+��gz���A�,7[źbX�`ZH����nz�	x$NzՒ�u�P`r�;�M���A^�)iң�=я���gv�x�R�#N ���Z�)�&��!řV��*m�Gq����>F�~Q2n�ʉ��$?���b7������{�r�RAJ�^�;��������Pv
�X^VN���?�	O>��S�0W�q`X��*�]������l
�Q�g#f%��K�nj-1���B>�!����6	��H��z��o���Q,W �k.�>����i_��t� 
>2&n]��W���b<@�0�P�y���ɀ�5 �\�9��0���?�V\�b�F�"¨�o� ��¯��-WTk`�0�Y頰7]�OW��U�@
链��)rt@�`��o(�1��,3>Y_S�/����_�A'~��Eꮡ):�j�'����v�	��r@B���	�u6�';Kj�_�������8����m�5Z���^�Y� ��{=O����&�7�9��M6���_iD�pn\��|�/	�A�/4av;T�/ �a�OM��-r�~�G��"_����@���7�ֿ^!R����|{�ep%Yt�6X)k0%cP�=��Ф�PzN-����{!�y��a��+u�����`����$,Z��ړ;��%�a�E��QK:�w��B�󃓴	�!&�
 $�}pP��&�W����Q�b��Q"tbfo��"�\��ʠ�`FQ���
b��	<h1�D�kE�����^p��W]0�����x��/T62��d/S#�1��Oo0�!{�y�%�����}^���<x�.���f�12.�ч2X���@F��.`���[p'�xV�<Y��H9y�Z�$
�ao�?��>��)4QQ�|qՈ�	ɀ�9�P�q����	�=!����:pxى`�-�e	�b 	�q���dS����6�v�'^Еa��U?�~����F�`vI��2��;i
JVX5Z[�
Ts�d����g�oV�*��-s	���������5-���v�2����-�	1�`���I>v$ �2Z��%�`�����?0�K_���8Q�`hV"U��	�²Ur�2�k��UX���O���PBq'cS��h�p���Q�L���p�s���Q�T#�U�,���)�Y�	XQw��%a�6E�+�/�������pЫ�B͟+�'�_]�s�� &�+�1��C�ޕ��}F�%wY]��YC{L1d�?jm�꫐f��}{�i�a�����ն�5���������Y��X*�oQ�_���&f����^;kFz��I���YS��W
�#-�Z�l�]�Ӈa��/��b�hN��ꬄ��Ԯ-�`�SO
����z���Je�� ?�ÏՑO���!e��1Ӑ�Vzi{	��I�ā�!%z�j~T����\'���U��B<��]!ˬq��1K�ȥH�Jt�h�^5����W bx&R���k��,	���y0B�r/Y�Z�	���c��GP4����:�<��Ǒ_�L�r�t�QȠ�`~�i݃���L:9Ki�z �?X�/)��ţ�~Zc���ߟQ��$�GZ��9Pk�PN�C[�q)
���\�
�T���sF��w���1/��Ur��>�&�㹤�	� H5�X0;	��|Q��3�R�����_Z��)`���f5X(�,��b����3����y~�	HuF��mp���`��
�����@o.�U�[�u��������[��-&�e�#H�!v(P��(�U�p��_��PPɈ�o��e}�tE�M4Ɂ���\`�R��J���A�R�ۅuM\X��G�h�qP@E��R�����0�N���o�� W8�R��>�s�a� ��f(��K�&>by5:" 0G@2N����'p� ��n�FM�A�j���Ako}e/�8�[Q^/�T��O�HW/����{Sh�5&�M�[A�@���{-/H`��>x��Pch62�^�� C�K��n�)R�u���B�A�	'e\�X�<�CA�鲇/	�Q;�_�n�1���W�k��4��J����18��v
?J
� �)�h^"MG�h8Rfp���ß]�%�XR�vS�PE9�
_���"���4����B/׀�!?\�AN���2��"Y�'r}֗��ph���Y}�E�Zp�A�)�;r�SR� K���	2{~9|���֡{�V}Z�<52�_X-'H��G�Q�x�1�wr�j��fpZP��S�Ȉ�a[��Ν8��|��?D�j(��7hIdB�vܗky��N�G:��[}ր%�����z�(N�C��]OC��2V�w^�q���,����ܳ�_G�a��1�$��l$U!?8��	�܃ v�P�iY�p��Y_�,�� �5L�uxi�~�r�_��' "�F{�
����A�/�!�>��Z����$_�-����8�;끋�MoP�(��J	������^�Tl%��(	�U`��	6�S!v�]v 5#���U/u��>}�3� ��s(L�*������tP�S��m"!�G����hAø/F��??x��^8<x� �[�"b��Uhݞd�i]Zԑc!�J\S��0Ҡ|�{�F�~�AUTp��Nº+n-h�,�	��������ic����	�HE�ʴgR_b7��!�G�B�c��D��K|�1��X6�F�/��f�nH�r����;�������j�	�EތJ�E�/�\]U�xNG�`���Z'7�*�GZ���YF K�Q�F.j۫�pAuڈ��E]"��dQK���>����@�Y�?e�+)+����RJ�-Q�^��E��� �C���Q����"7N �]#�y�%a��E����fvG�%�w7��B��<�P�t���g҈4vI��
��̬� �
)�-� ��r61�! P{e���c�������.a3�} {�o<;B����u|�_�K��M/��Y��gͭ4h/�Zs/�N7�a���G�.�	��Sb/�y�Z��[�v�/� +L�����A�/���0Uv"P��� ~�vX4W_(������[�����&�`M
^�к�m��
�N^nh �w9U:�X5 �� ��!-�Y�Lrx��`^B:d���1��h�b�q����L~]%��W�����!ջ�e.��� 2c�m�h1_@xnD	�v鉠͹3T�8#I�pnC��O� �.�|HI�n�pĲ��5��N#��(��
	�,��t�quN���N���2q~�b��Af��-��1�R�d%�Q^T!�N�ֳ�������*��9Q�]�%�ku�!x�"�6��L�e}&I�׏����*�ǐx;�?21Y�=�y�i�R�x<%CTuG�gZn����W����R��L�鞇�^)]���'n9�:GM0�&��<���a�� ���_;7��U  ~�H�)r�$[e%MKd]��i��	Ku�^�_E2'�Q� >�2�s�X�?���Z��߀�^�!�.6����yq5`��K�������)�����--g�I�K������?HaW��M� 3-��y���m�i��u����]�h[L���3�H%��2t�n�>_BJ+�A��P����h	�W9M�;�1��쭴��\�WqZY�3��Am.�ަ �WE��?X� �6Uw�9/�g-mV��@��	� L7{�S�$������B��pŮ���G oSg���BG�QN�����9!Ë�aK�$O��v|!��56T( 5�%�O���z+�~/�\v%|�T-A����z�p^�fШMP�u�h��q H����X �ڷ��R@��}��v?��B�!����t�<���aߘh�}�_��)���_Z�!.�����$����>���(�� 0�������L7�G��H,�(y�I�J�ș�����vw~N)�b6��BY�o�<���l* W��G�A� _��\�b�eR����Q��'.t1�\SˢC���՚��~��Zk��}�]�t���cT�V��:`�5�0v��L&�o(�6�c�0Zd0�P��&�tO����@�1�m�
�i�ܢz싱��j�Y��C4X	�J�q	V� ?R�p�0�E���e]�iLxU��-���F�Ј�~�ٽD�m~��f�)�b�E! 5U����g����9h1�4���=�k8 7Nk��� �ҹ�� ����ҵ�+�,���N�T��	�t�m F,�oM���h%�eyƄ�����	|w{"��'���A�P��K۝���p�K\��VPh�#]�(��j����Av\�X�L$�#P��fSz����Wt	�nG�aG�"AH����D�Gd�Z�tQ�D�� ��lYZ��A�h.�+mgW�qb5�_�5�uZ��	\h'��,:�as�΋�q	i}�q��>i������U���P�����hzn�I���Nk]�ߢZsX�L2�y����֦C/	J��̖�pD�P�BTA{��s�-.�t�I�-W�_���@7A��*H6`+9E�-��f?K���(��)��/Aj~7^.ae�G"�p�В��]�/J�X�B��CM�Z��'Tp�7@h�QK|��F���v��_�����;V��
)��<�"�-!�WJ�lKg�S�S��<@��8lC��i��s�Ŵ.[�,�{h��u�F����20BpI�P���o�~�A���7��l�a���!,�O� �%r}n��V�Mc������8�uHE��LAeRw)��|	���DS���Ӑ �6�~��&
������@�ƛ�h��#
�)���`^F=_��IR@E����[�h�S��h�)��K�)�[�;cdXP�|I7@��S�&4��ƀavQ �ջ�0*q��۹L�;[������2X%�Y�d�	��� P]��n�J��~��7Y�z2Xd'|1�AϨ�O�3*ž��������_!S�?f��Zg����� �'i{�߽q/ZP�8�+��1�K�y%VD>	�3�ER�#�C�����y%�U�/H-�m�c��3�É��*�
0�����`�h�~�qa�_����Ub�]\�'h�SX�;x����X���a�1�K9�kR��h�u<���t+�/$��:��� �)H؂	D�#��G,�a�Q ã]$���H�&t��$d3��^�7��>|	��蔠0�d�')��l��O\
��$<y	������z\'��T���M�(�� ��uH����31�pR&���[Y��X�u�B/�"���Y$	*��]-B/�
w�BJ�e��~9�Ѕt�k4�<� �>nӽE���sl�P�P�h-��1�+XY�G�i��i]��
�H~ɜh�"�^р�%�k� ���
���-]����.U�L�&�5@g� h�Y^]��b��P�N�4:��n�q���HV���u��� 0�-(��Y �),�vm��B@�!k}QX	]0q� :O�t�} d��A�q��;�Ri��g�:T h�sQ�-HP�'�
��v�XK�]F�l�?�O��Q�)K���)�	���P�.@����d>:��	邢�] �(�x^��*�oH7�d�� s�~�Y`�;,�U�)X��-�������c��[hRc��1�?�d'�	Ŏ �L �W]UY�k6V|C$�>�ٟW4���ڔ�L;�ϡ��
�����]4���[�=��`
�G�{��p�������q�W���s)�!E�/|�6���+_)r��h�
� k��K'(�-���h���P���T1'XM�;�K���@^�GJ%XF�~�8 �BQ	�)=�1x�0������͝*|wd�(^�[�ZV�S�c
�v)�	P]��輀Vho�5`[<�c/;�X2W{�J���i4��� l�"��h7��@�%�	g�a��܅��7��F0�NZ0~��桏(p��Za���;-R��.��Y�T��h�O\퀴�*Z(�����0�4`tZ/�0��R�{��YEM g�ϳ1莳	h�Q$X��߻E �~��d��Z���bkƀ������|l��Z�1hq�*X %T5�L:=��hb ��-l%H'���; 5P���h8u^�u�*�69&"�@鐽��R���z�r�J����"���Az�Bn�&���$�z�٠�M�Q�_�/�0����`��g :Qh��j�de`�\�x������+S�����{v����w
�d�����@���>B��K]��O��2�ZY� /�t ��@r�)�4��"!�y��\�A�$���
&H�%�h7y��T��}����F:�O� �.�,^���r�ً��k%�+0<b(W hTȴ���һ��t��hVX���4z*��e�o�d��RHr4��jnL*�(����us1bR	�u�J��
e��9�T�::��_���	+��eY!�p�g��\P�O�q��8�3*U��].��C"���1�k�k�������W��o�E���o�.��c���z���)��˜�h+B�p��;G����Q���0�ۙ� �}^8�ܺ=�.uV t�k�p2% l��>�^�4n�*���x��L�Z�o�dU���'���L��T��}��. � �Q�B�5T8x�,Ñ~�M�%���1�!`�E+��S�rh,H,�o -/TaZ�I�����\=Äp���M@�0��V��Y$���ǧ�ða��� p�7A�NCsPh�]G&gM釄.���W�o�n���W��S� ��>S�)��L�P	h�Z9 ø�u'H*��vQ��r%�za� �ݴ-^�� �7h��Pvz-�C���A�g!��,�� 
��`�M�vۄ�m��U��9)/	��'�&�Qo@}S?]����$�)�!=�_�e��^�u�	f�h �R���[Z�ؼ�g_I���נ<��ֆ^)A(/mHDqM��_W�C�8h}���x~t4������LӤ� &	E�� ��[0�M��0Y1ӗ��TK���)zQBq�B;�B����	UO�X� �S<�Yv	P��}2��u!L�Qm 3���_�I;O �l�`)PU��D���%w#I�L�\
!��@�Y��,=���5�e>���k/,\�aw�r� ���{�-�[�H�|.��� ���~; ��I�%���	C���,��c�I��\L���������'�`���Z`���Ah<F�$�I�b�\nx��s��ϵH�-��r�����z �\R��S�2�%gk�j�v$@\m4o�����zSO�	�`n���No�aK>F��[��?��HJ��=�/0D\Z���lO� JygPw�����>#A����3���/�.���^�rA=5&�bD@V)��Mw�X��l��z4RdV��v �Ŏ�l�����+N	�NO�o.xC� �-V��w �21�^5DZ<�"���t���߀��?)�~�(t����ea�Ȣ�0�b�t@�Z��qh^X�'=[_7��t�0�M�K�&���-�pyP�Ԃ�h����j��4�0'wE��1��Pýϒ���rK�RaӐ�K�����o)�q����%�D+��X�5�Q(�1�8^���� �A�~�/g�H-�dV�H���\�55�����ai~��o�S�q��,?�P�%)�{w8��F�j�`-�l@�1EsOП�Fu�	p�O| Ph�;�]���t��p	K)0����C`W�(�ʅ�;�Z�z�P�3`�_\65B��
�y����^f�z�����, 1��@����xfP��?��e�X��1Ag7x��yT+�D��e`K�J��W m#�~�ڽ�[hr&JordR���:�"#4{p*~� ��L�$-��vP���h�6" A����W�����i�*Q�e�� uh�X�j��ï~ ���3Y�E��A��Eg��Zlp �1�q3��)^Űk�$E��9j�Ԝ`�2Y�4Z@#S�*9�[A�<�	+bHV �U���c�"hPK`�����;��!y|�Ϟɯ
��i�$����U�@J�T�f�-�\l�0o���,z�L0?v\n�A��e<\(A�����(���Q�!Q%������������F���P�|	uQ�Ph�IQT-�.�%E8D�~p�� q�4���˸E[P��¬z�����>�j-vFq��@k �C5!z��|������d򀤸o���:$l�	�L ��� ��oh]K>�=���f2i���T��"o5�^s�����?E�����T
T�{���<.$W�4�h��	'b_�ʽ~Hb3�S*�����.���q-�@"��0Eb�g��(ꀘQ���8 ���,[
�	�B�Wfo���I՚�`�W&	�)�W��	}����A��l@�KX��#�]�������Rt�<ǻ�J~Y@�V�J�ZW�/P��f��j%pW��aQ)oū����ɶh>ˍO����[�/��p� ���fX��~sb�����.��f���{�S �0�O�@��&\Q��] ��YuKW�39x�/!�����P�Th�&z��O�
@�ķ"����%|I�B��v`�B�7 V��k1�X��� ���)��%n ��5D���h%�FB�GN�˯������2�*$؏�)��1���ؔ	R��e�b��\��of�p(k���D�>n���� �TP�H,��>�0���-��h�8��[�4�R�@���X[EJ�Q�Q��w�	w bH_@�+��&���{>-�����Y!�k���aƭ���|_!n�41v	
h�pw��۳@�?eg�1��U1�.� �Ph	�JY0x/pU�F�ڻ	��I�l��F{�p�'�0�NYHA[,CVO	AZPn���j*낊���e�Ǔ����>K��-� !�ZR�d(0�=��,��9�Ѭȗ
�����,� �(�J6��	F�x�-|��"P��w>���h�]a�� U�8�#k��(0 �E�iD?^���J�J,�:��|��F�W^���pv^.����JM��xF<Yh
鎕�-�R�.��2Uk�0�LB'�����G���1-~��T^u�zX�	��{�	�h9[��$SK�}��)��
�K���*��V�T�ю]��}
�F�K1F�[)֯�E�CD� U���?�7��� Ɓ�r�}%��h����$���D�����7��� =�Y�1Gx �z�9�<���ļ�K��%�b�u������C>H����p�O���6���N�fi����y���K��P?ȓ�`=V� e�O_���x��XT�iL��O�	5�N���"T.��W R�O�`@�]��3%�V� nk�s%r�5U��[��6����#!	��.� �RQh%$l.������F�s&�@�(c�h����{�dP�A�
gJ&5�r�Z p��M���q����>o.��|��n�B��	_��y�~�~x�z ʸA<�IP�`�v��������A���}�Uc.�{�����ԧ)��a.�扌� B�DzM|���Y�@��h�kF/�y�a�+�)����4����N=�
G�#���c�!������6r�͙�u`�%O��4�_�#<`Q�w�B\A0�1I�9�(���J�\w�ne��'�E�$>ހ럷?��� л�o�BfD	٪,E/[���0�c8�%)ݴ+T{�>�d���`s��Z�'�.&i
r��C�����pe���)D�'1`gm�;H�7�0R�-�=�;R��T�vx_���9	�Ⲣ��ү���������0� Ӏ�B��o��\�<�����Ͽ����F�ئ�h醸�z���U� ��9�p��l%WLWN*���_�8 ��5�z�w-
m���wHrT�hb,�r��QQ���Љ�j����f���H�o}�@�D@�%���`hSy1�*�bP��xc-�F��D^��y�<bM���$���L�ħ��m�h��[��ǯ��.Cs�"�]r�ז %>7 ��A[~Kr�/*Z\��u�:�xO�B{�v��f] ��n���Y��\��Y�wNSh�z�IX%� @5U�>�	�)��G���)�F�?YU�ښ|`cXCH���+|K�����E<��3 Ͳ�N��U�}���Z�����-��{I�A�7�p��{����C�-�%a� V ��b#D�K�0u���'A)� ���c�$1�l^�5Rah��h�7k���gHp�Z4��$ Ng=^�W��0�q:3{���߄�k� y�t鞫�<��Y�|z=�6J���%%՘��X~R'P8�͜%E^�۽���W'�*yQ.+ ���K���!�4��̰Xf\Q���*���$YX~����J�~��Z�*��sxSxY$̌0���&a������I,��'GA<"�/�4����'C��skA4Q�[l�hH��J� кB,7Z!� 	J�6�a��(�e�a:z��)��[�@+�_Ҁ�Ta�����0m��j�u�W��gH����*g�5������s��T����Ćh.:P0��Q��n���]"��*�J|���9�/� WT_�u��=���[�R>0rh��7����/���Q���-ރe^��zPؾ�j&�{&`Y��Ȑ�%CS�R��;XP�O�)o��vP@�$ �4��;��G���#��	\V�A邞b����uG�)Vq� �������[������O�P���w� ��Ha�~�G�v�E9�t뚢U>�i�@�r"좟����@�ﵥuM�@����F��hT늀�K�C~�%[a�ňz���K��'����]��?JU�,KW�[!�1�/��L�Q�GX|g������FSV�^h�YF��9T�*)�����~)��3v��+i��Bt�OS�A�K�bk����$��~ �_��Z�{��Ǘ� �=(�0��o`��'��E��cΘ)���wL��I`��r��颿�MJY�8
h�=�c�1(��Oe��Ψ)
���|�~[���-�`�\^{��\O�x�b���k �T�����}�XDI h�6Y�N��0��9�K����vQ�Ĺ�9C}�[�s��{��Є/�+} q8X�Y!�P�P�L�7��������0���?-�#)�	^T��BBW^���mTr�/��� �խ��q��� AEj	�Wh�\r��z¬��CM�����v|1�J[
��hgQX~	����ъ���O����k�HN4pZ.�IE�L��ɺ=�2��ܬ��+z���J�ځ�a�B�2$;�w�/�Q�X������X ��?�hph���`�A#qE��'�;��pB!���O,��'��E�"\Cd7��;*�=``ɽ�_.�c_\���%��3�`a~��X}�ZA�hΠG	�d�\Qh�tC]�kbJV�X�1ʷ���EBr��ǎӢƽ	w蛠\/KT0.!�^8�����ಽ�+����*@1[����3�nQ	�����>�r���X\��_â�^�-��t���$!]`"�8�U�E)�-
��XSa��J�^,B=�ϟu�$%�F�m>'�t3_1���%��w�WNR���\yl���	1�Q�-����7e�_��``���-u�dkfZ!����u9@��Q�nb�=I-���C��2��&��?��{�G�x�t�*���"��"@H0��f~S�@���I:XMe�fq�YbhZr�
�����w�X�M�bRsG�7< .-����1�)�
��E�­!�W�`�C��=.@U�3	����jH%0�q���Ȫ`�eZU����x5��b��HT�[%-+ڷ�>/�N��h0	��>�@�Z��?1iuڅhV@���O�bi�y�n��%����4S^'��^ɾ�d�O]�o�٠຾� F��������'1�mN�1wTm�����1�鰼W��u� 0���h"��.�0���0b��(=�ټWæh@��]G}UB��¥QRA��O�
8�ADӪ����c��2��ru����?�s��x�-W8�3�y�h��/c��I�<-�TV&iqB�K���_��!L,��9s�Wh�"���ܠ�,o�a��0�O�Z�14%P �ɝp�`c
�E����0�b���:��`z��ߵR������Z���LU>�5��Sa�wſT�R ��eAihv��[`���RJTl������	�'���!�R��� ��	�(O]yĠ��_C�+��Զ�p�Zw�O�ՀXt��Y�O�u;!�*� L��;
`���xX_|�sŻ���pe>/}-��CN��Y�)ݹ�,A�Sgf0:I�}�@e�	X$CVC�	 @5�[��` ^�`&�J�2�U[��i�G���{f�X<�(oV
d�%0̕m$@N� �1#�/&�;jX"����O����	-Q~!p�z4��^)荚)��A���:1��6�U1�1� ��ڷNϸQ ��j!�1��ǘ�r�Mz�P����[�>��s��G��J�k�{3+/�I[z�m��д�ٕ�}ٽI�e06rQh@n
UJ������A��nj��~.��<��N��)�i@�h�2��2�W�5�4��c:WT	���}�8�=Uj�?�g��1��4�����d�����T�e�w��0Kn�bO)sW��?�B&_��T@sz�y��[��;']�	�$��f�^.5-�c�1�"[Q>�W��9�@}���{��aN��>Pp`�H-�MG\&�(�0;��eՀ��Z��fU4����G��m	��_��ID���Z��A	f��8ǐ�-���~�P
�c���1��>i	 �=,�S�p�N��=(�,��U	R�Vz_�Q�h��_��XQ�X�;�����Y�ozĤ�b{�:�+�l���s�UZ��^0沂�.d�h�b� Y�p�)��Q$�x�~�3@1�!�	$���n�a��W;&�(���׼�)��aP�B"��
W~px1)���,A��͞��(z�$��Ec����ܠ���bi1��m��k�J�HV�u����̛;9�m˰��d:tZ� ~���5���æ���䅍>��NES���ٔ�t��W�1b�4J2[���Fn�	��2�J�N��8\�k�t�+�G�m~�Y�4 ����QPt�5u��
���o?J4������ĝ��?ɕ���:�9n�)�B@�&=�`'�3
�s�x&>��-�K���`$��&:`j�b]Ηa*�<tJ���r^����] ��V>V-�|�p�A�,r��Ik�~�PR{�痁=LGfp[�^���؀U��&�{��=���E����eMU�#U�>׾���G��h��`�*,@�-\�@��=����(���' ̎���	.�hK�i�i�z�����-�0q�/���� 2�X�{~��O��� �y?�!�cH킞X�7�`n\h0�5���IoD)c���b��fU0��,��<)�����e]��|�N���ǈ�%⺈�f0� �ͣÄ��Ê(���3@�Dԟ�2'�"B� 廒t�f�W�lH��'�<GH�;W�hձ����f�V����F|���TO�F��p��[�;B�ƉLM��95�X�Qw&֠��Z)�_=���8�N���"H- ���;���:�1_��;��) hXJZ0�,��en�z!dD`��r[^����*�Y��<�Z�-^k��k�NP/�̱�	Mb �Q��& 0W5wB/)��%bq)d��EU� ��~[���F��:!\�u��ڒALZ�a��M*'��5�K��Թ&�<
�a�i��,'�)�E-�XA�'d��#ao h��e:\O��C�o�� v�*Ԓ��K��9�7�ܩ�� �Q������.�#M#k[��T]���2��=��sG���& 2�hkZ}���O�E�.�(PƧ���~���,�a�2�����D�=@�X�� 5�h���9�T-rF�B�(:�K�/�=P��Y!�z+�@����Q���0⣔���'`����R�O2{w}J���9��8�܀�.K�5�Wh�8N��1��� ��S� ?�P��~} WHrh-X,y� w�{|+�,I~R%#`Z!°�cSP�VV�A��4��r��+�o����� �q	�+-�u�*�����A2;��V6Z;����}����{���?aj2h6L���I&CU�����P���8;q'�=��c�0;����>�T�P1�M#$�ZR��L�rpM����D@��W�D��m(��_T<��`%�#s�	��u��kz�2�T�cē���]	(ʜ����AJz�&��-�k�]~��ξNQ�"��_�J�%�0��ߡ�^�����	h	�X%܎8wg�Bv�O��W���(�&�g��]��l��m�@ �N�@�<א�1ʟ�"��a([^�*L�!�	o����?�1�KR�G�Q�CNd�ʒ�V��\���܍P�,��H=oHTHFZ� Y>���)i�F���G�2�� C-�h��y&X}�>��[<
��t,H0�p@L ����)ݽ	9HOF�:�9�s�.���?�x�nx�8��K�J�������_��yfn�nP�ߖF��J�ݦj�Շ�ȳ�0x,�s{�Z;.UV�T	�l�53.�{��U�I~��&R��)�	YhS[�� F?|j^hz$�`��g����2�t��"�M�;�W�v0�p*�oK'�­UvK�t�%�
u���I~�(X5�u����e����q�V�@�6�r �_ �T&)�L V�#v�Z%�� �d@=A��~ ��k�V��`&>Ǡ�0��gb���߅�(؋�:�x�B�)��<�Ўj�`�J%B$A�U����c@1�j0ֹ[eL��`1����:�%5Q�;���
��]�n�.�>O/���O�L	�$ּYL�9���I������R-��dO�Wq�� "{�"�Mi?c�Rk�ŷ0�DS1{0S���l{Ph@8\X- dC�?]�g2�}��TZ�|[�%�XV`� �f�FZ��a|��� G�۳�!����\�����9<z�G����X�w�0)S�*O�ZV���Y�zK�5�"Me��c%�CT��O����l�靜[�o��f�h !�.u�á��i(@��ո�0���fh�t"�z+N\�� ��OP��������L�	%~& %h�P�)^��\"��2�P��
ZS0�l�L�$����ؿ�!��
��d���4�Wb/@B�x�)w2��}nW#.5�&�2XPS^�.>��|;b�^޵�_t|����|lA����&����BKr�@|f�`�A�["���S!d*�	Y����u��.X���-�1��6h#QD�m�z��٣��8}S�P&�KfQ�"��(���,�yR_��l]�%�D�{����ΈݡD��z*����^[�Jh/����?,��� [Z�������x �X�h���6�%^dbJ9�����3Z��{�I ��c�6�mR��NR����p�hd�f�Ǌ�+z���G90x8G�L�k"o�
�t�h\���I )�_U��l�#���Һb�2�;��)H64������nu�D���!'����"J	�8���>�R̬�!	9<�ip�Y��?z��_o��[�����1�!Ő�@�h�"�(�˞���/��b��W�x*v'DH|'v������)�9�Y-��*��\8�����n�m(�,(���qϢ��+=n.�)�F��}+�� ����A�.%�x�O�;,Gi�o�n��n���$n�r�J��o R����b���)�NZga�JF�����h6�S��;��Tn���wPY-!$��ob�
+��Ob��G�{�(�4�PF�vHޔ��࠸ �r[:�l)�f1ŭ�4�y"�Dt���̠�hj�+XH�@zP�^5��	)� �'6���qe��E����Z�a�H��/�'�M� o-�N1�Q_�+���+�Ih N�[OC���A�(7v�B?$3R�����-]e�tyV%�}o;e��;H��m�E � 8aw��qPW�K(�#�D�zn����J/%W g�34{0dg^h�b��B��26Rk��-W�_2�J���M#�m����5��&��H4-[g�%!
k�K0���)k&���\!\
�B~ˎ�S�mj����lhU/� ���	��
{AP��Қ�A��0�1§�� �S�?��`�`%U�-��/�p���A�S��zD�d:a�hPCj��86�ޏ��$!��x	� �1]Pdت�vgS����8�@�!�[]�õ/�
�o��|�;��k�7�X"�	_W'o0V�\Zx��+�z�	4")�J]
��+Z�D����9��&_���*�-΋�p>��	����9	7�;EBp���ސ0 ��@-V!�x����`4M��:���AJ�8��(�[h�;`!�@n��}�>z���V-�~��B-�����"#��� S���0y^H�<� p�:0k�x@5g�B��z��Gs�@F1�_�)	��~�x�`!f_�P*T/�`��s��K[����J����H`�Q]Y��Ch/"�U�;�-W�� cU_�m6�
8,	�zXZ.�w-Ԯ�H��I3���%��e%�,D!Z��[	�H1X	'�Z�r�+t�	)	b��P��uQ��3i��hnH�n�������r	�!ue�G�<<�\ȦX�hoYtꬵ^�B�&��Uď	�|:���_�4�g�z��&�9�%@��y�M�#�����/� -*Qs�1�-
z@�����0%�`�7�y����7�t,W��
�"�y�L���4!��,�О� Z0�YQ�d�Hs�v��'0�0����'u���1�0r�nnU-o$�kN�� �!�-�j�;���')|��h�H�քr�@2	�}��/ û�mYhI&�K]E��tfB41�[��'/@�Őn8Uը�Q� �3�)�X����yc�@E���E,�%471���f��� �sN8�n:`!��iQr{��o'{`��KG�����of4K7�0V��3���F�.��3�k�=�z�u�I�Ph�?`|�w������j�*gF���nJ#�E�j:-�G��S��ePy�,�1�A��R��D��(9ڈM�'�����F2�P��a-{y� ��S_KV�l�Q	���^��\�	�~}��x�6��,O8��w�Yfh �h*����s�|}vw�/�p�҇	�h<."�P�Z����R�� &��^B�2�]3IS�r�?W�()Ŵ&�>:����p����S'_Q�e�sg-ns���o�:;��5*��ݺ�{oz��5k�}R�|��h�eugr����8 p�{,0�y�~o_[��uq�W ]�-�:H�C�X�����ЮF�F8� ��U�h�("%�4@�-TH��'Ap'�oz .:h[0�1�r��+�6�@�3r'%^�����oX�� �|I�CB�@��7H$1.1��`2�7B@� /yS;�Ih����V��Z�'�caCI%�g���kXd���[bz�o��<� �5���9}[i�ю,y?kA`����O�������;ې�/H�,娀��9��*�{�
2q�,��A��j~a�@xn'��4*�ҹظ$uqK{|&j�T'�.�2�e��0�ﮣ��G����;+�[~�Q�����	���_�)1�	
8�~�~��9�.H[��|c*�{��!�(������T���Ӟ�/*[_q+�nN`f��[�	�va��[Y�b�_�X;�0�$���]$$K�U�u���ܯ�h��[� �ZhWL��&,�A��ʤ���KƇ��ȡ^.X�I/{8�M�Q����2ͮ�Ο�̰��*^l��1[�������T�T|��	�����")��1�Q�!�9u{����G�Kb����(���1ZX��`�US%�P�#t��))�$ 	�	'*��X�nr�� fSh"��?��%��M���u��N��#�>�y0n0ޥ[���2q�8��Q����� �x@g)(t�$HYR�CA��\�I��٧ttX�'�OX	,d6�<��(u8��8�w5���$�O�p���4fT���A�8�����;�������׽�m�	u�졣����[+���P��0>J}��8�U��!0�s`�<� ���rj�=��`P��[������1��jө����z����S	�KR�lΎ�w����X=a��<����t���u�x'ÂwoB?D���}A�?�ۃ�Sſ��i��~	� &��AMx��io�o���
	�ɗ~k�����u�Y��nowU �9>`A��m�w��:��S%�+��6�~j��Ӫ�G ð�Xl��|185�:��g�Np�A��[����*%4���f{,L|��c#`&(}��1��ʽ+4�t��0 �R��@�Z����ؐ�(�Y��L����L��0]z���.�c�Ln0 hQ^�f���w]�|\�sg�K�|N��Z
,\��C���q;������ ���P���B���#59+����A�g%�upu}����a=�&bvhb�y��G4W��kS GW��e�=%&P1Z��P1]�y����C�؀�D$�Kq cb�RI�	�>Gg��x Y*�<+��^��E�f���0m�	Ά~� ���4Ҡܞu�,�L���c3[��R2@�S�])�ۗk�,���t�S]��O�I�>�e�)�M��N�J4(�(��%-��W^�XXh$lF������O���@�;�;� ���$�,� �A.eoC%h��b� 5�'�>-�%p��4�G�f�k� r-�^lac�k��g[@�^�e[/ho~3e�)Ù>e�`��.�\�{���{���<��J� 0�B�{���W@'����B
�
[��%d-�۹̥Ps���'u�	��F
(|	���#P�Q�t2_[� {Gn8щ^�΀Ll�9�H5����>)� �Ө�2�A��RBh�N!�%�wU��aM���| �}�X��v��T[�S��QY��N�ȆFnX�JԀzsI�	�t�h��X9��J��g,��L%�4��z�Q\���}�1��Z	�X���S��)(�-
��z6HF!)͸��R�ř��Y`<�	]~@��)ݾ��>������!}�
>�'*B[}eB�W����j�K&M]�ܢe���ܣO��[I��C>������8��q��$�oM_��H[<�h=u�][��.t��+�K\R�gB>��'v��}�p��;�~�x\3@�����
&7��HO����)t#}�0�_j�K AܾD�� ��	���� V��2�)`�.���,wdz��5�9%�<�������y?	�J���Z5�d��w� k^�X�c��۔�08w��R#J
�e�B�(4���s�L*�U�K��n^ߝ����3�1�^΂�XW�R�Ć��M�h*'�~�/�|tC���͟4Ȱ�H���1�=�	��,|&U���	�yɃ)WZ��d������AE�9�h�5*�����
a)�P,���u;�oYnN3��O�=�,�nǗ�������y�%��0��
X)����R�>O_F��05}�K��\��#�6�f��`�)~\1�� �7%��t�q�N�؄cX�1���輰��S���ٶZW �PR����6�x�P�Z������4 ü��e�d�+���1ۭ����VH����^�d��0\{�<�[ r�~ -@�B��nJ�x,R_��,�-X!���O�*�Im�/�PYh$y|w³V_���FAn�1M>�_�[]����}m $ŻV��� HzC 6b=U�0�'�7�p���Ē����j��>J(��j�3	�	]�1�^����L���)� ��|!(K��]�zu`����%�y�b�5�H\�L;�K�d�R#`?��:e��1����Ň�ђ9�Aq�GH����$}D
��p��J��0W�E?~�u�~�g`�O�]��Y~�s�3�Y�b1Ð����E�������1�Q_I���QEH���R�`S0�� V�&I�Iq�Z����"Zw���`���y�
�p��p�|�����TN�0��/���%_>�i#]F.>�*�f<7�}�͑ux��.�2���@��=��E!���g~8��C�CpM�g��K��d�]��s��\�����������4���A�Ws���~0N���Z����uE��D��-X��$��q�X-
wYbœ�d�<�R�1KS�z��a[h��wn�p
�jz� �굶�ﰐ%M,�E\4T�ȯ�&��fQ���5��V[�I�P�
��WqL���P@1N��a	h�VGd�P�
�v͒�PH�^���]%�Za@^F2!������3%�dE�b=;j\Q������-3��nf���5�)b���1xe'�ՀM˳oLOH��M<.�6�v-+9x�6)�E�L�^!��rs ��0�b��[�?�T,w��	Z����o/	)�R-��r�,pHx=���@�ͮ���]����p����w2����="1�SZK�ʢN�p�鮧J���|w.Q^vZn������-s��"�)΀��N?Wn�l��I�V�5L�@������!��eI{��Ǉ�D�K�sy!�	\�N8\JN�kR	fh<ZW�Yl�r�~�Y0����X�-#a�����Kiu��A��f��։Gx+��$��������߀�FN�8�i$����-[�AC�~�U�m9��(�0����&	s�>�.�׈�*��f��հ�{+�ф fR�Ɉ��S�b�u~�r�q}D�T��c�y�+�C|ւ�(��2�Q&Rh3�+�wH2�([�{��0/¬�5�#? �@;��U
'L���`��{:����j�w�Y�����h)C��yAw�A��t�J���GQm[L)�]���/AH���x)��C��5u�%�GF�S�(@����(Ϝk}uA�!�y�!���D��7���I�-�w����N��_��ݐ��A�O>���K���}|�HU[�y)~��A����P��-�4�$ W�<t�D/)��(�7U'H���Y��%L��H�H'p�����?^[���Зŧ�'{h�ێ�n���J�♞�e��9Bf{o��̏�t�XE�_	0�r��km\�/��0�s:ô ���ݲd��5����Y(��X Է���������C��! �������0��BrO&��	����]yf� ��e{�,a��k��R�XF|	$)�ZZƀ�8��Ϧ�q�@�b\%WZ��A���{��e=�M�. `^�h� V�v�s���>R��>��xO�X�لd�����A�B*a��ϭ��!PLZK ΅^��1�YE	��g��z._��1b7�{�	��>�&A�m��QT��8]wW��P�R�%�Lp5ܛ] N�Q��B[���� n;�/�#_���#�H|B<2
ZXS��Q��������*�^G'�����F�4��c�/	EP���`�B(���B Ӵ[�����@����B&cԝZ��:d�{���;[=J�?��j�hng/� ��)_cA��^7}�=	�	��U�'\�T���b��u�R�����p�N WZ0�1��O�`]ֶ�=�V�dbb�>HF &����c�Z���S�25P.���bu�	V�'e-����1'�@E˥	A�T8�h����b^Ut5Ωb +ŝh%<Q}���}�>�`�y���a�; ����		��l	�_L��aa�BR���� ��Ap��Ha�8��Yx��J��X��,r�0����ǿ�b/Y�qJ��1�S�
�})��t��p�wP^�C�Զ&1����8�Z=��8@2F�O	E�h���_�.������&��w���1��:��c k�@5s~��`0��3�n�[��s�
�u���U��w��Ph�[5^D-s���C� G�j�g�T�0�/�w6���>�Hk?	?O��9i;�P�7R\�JSL�����_�g���Ƴ fַ ��U�x:z��Q�K!��R��a@��oXB��Y&���Z�'	6_��i�������j��0\��>V Wh�m4[�L��� =�;�
&p.�(�R�X�:_di�3��`��=����Yc��N�1��X��Z���� C
����e�v�̦�Ŝ0�����Һ��6�uQ�
��+�Z��+�N�PӤDBjm�}�lz-GbZ�U�Ӱ�;3&������,����S^)����X�D���%r���	�]Z_�ydb��U�t 0/�Z+�Xy��}�	�Vz2�F[�h�-H�;1��^)��.�Yz�'0ٸ�&��"��fŬc
	��-����)�5�1z^��k�q���f�X��U��QN�	!���c
�8�"ku�0X����U)�H�iC�b�=��,Kü��h-� �R�V)���JY�������x��
��V�e�[�㡈@��)�2M�l~�(���K^����[J�,�L*;]nx%|��9��|/��^��ڠ�S����L�[,���A���`M�����CXA!�W�l����,h�bM�<�~L�f/V�ِCh��b�/�Y�43�M��=Z���������(�=0��^	�����h`��t;p:���Q<���.� r���<���8��@�PW	�>'��y1���hb�k_la�0t7��@��D&�-:i@�4Uwh|	>�/u9����!���	M�oJ����E,�	�W�T�%f$�sw��u p�):~L�
A���(t�ƕ��ӂ����Q��]$�A���h�I$�G���Q�.	 �ړ�0
8�B1; ]���"��Q�;�|��2��ՐP1hj��f�D:�0����N[%(E�	^	���X�-��퉉�]e�1�bTX�{���}n�ŕ'��P�zOf���h��(�諰��J}�ڄ�^��)Z%`U�rk� oR>��:�o4X<� r_�釽[�bX[���f���:��Zd�Y��JQR�]��2CV�`�1�I�Xd���? Ƚ<dk�"s/�c�&X��	�<}��pzM_:��+|0O ����_��
8�%ZVJ>�"W���B.����< �U!WZ�o�g�d�1�b�O}}w���TRė�P�[�dW��[H�d� �ɝ���Z�j1��ű,���x�x���\:P�%��C��Ā�	��$ �,^z' c�bh���!�l�2��-P�mO&-�h����]}Z����Z���3}�;�vZ���c���	3Y|X>j&~C2��p���&��:9H$Gf�^�[^Р��8�1��؟�J��-_ 	���	��<��|��;�!��xZ�9h�cU���1�g�*�f���BTXB��� :6
�%�AV+�~�m�NJ������B��8rBaU\��h�Q.�ѰV
�Bl@�K�:|�@�-�{��)��a!>*���������O�(�!N����-	�'>;�b �l�n-ckdW���5
 r1��(V%�x�'?s!خ��/k$� �#���/)��cZ�tYY�@�k��/�g�(�����BC�T���Y~����BH-G�r J9���[�������b��V�1���+�c��MD����P��!)r��,��`yhwD�]f
!FS�����g���~��Y�����h#�Z�%f)�����HMV�dI�W��1�W%,qB�*8k���W�bC[�;wEp��hJO��E��N �j��viL5:��nH%(/ho4�5�q�E��t�5kI��Z�Wk1�X8\Ɠ-����	�hX:U�q�̋pvQ�1��b�E��զ.�F��uS�:c2X��RX1>
g�QhY���� �w� ���/�w��eld��W���[;�Q^�L��j�q�v!�rA��pv)H�jL�L�Ӿ��o�b�cy	n�~ńП�����,w���v��0U	X���2����SW��lRj W�>�bM�^��?Vn c�\�P�-�
VJ�C?_~�T;u�c��p�e0������H��s�{�#p	��oe���'�.Xh}`<�:-"J&)�BYp\���gq��ix(|�`!Cq@��\u] C�$e�m�$��pJ�Y��7:�*��k�%�}�����so򆫈��SmVM�+�L>�@�h��0O��-���^���%hZ��	�/K���Y�1�����xxi�\�'Z"��}~C �@i�^FZ�$J��6K�𤾲�S�>
��ԣS� X���\�X�i!�D '��_JN�X�'�	�3(� �`�8"vv�ڂ]s(,�`��?�XC.��=��zXE�/?xQ� c�B�+[h�G���I��Nm�_@he$>]�͔6��ډ	�t��H\�]Q�����Fh�3/���Jk}J_�k	��H�_����ē�J�A�a�3�}�V�������9�����n%�H�$*��uo�4	�#�q� �N-
�����ES
h�u��/�z-/9*� ��p�pc$�M.���X�#�'��Q� ��a�X��F��%�m��	�/6����P&�B����ov��a�W��U� we)�H�-�$Lr�#��!}
��J�t�,�GQ�FW@|P(��S���/R�� $�*OW�m�	E�L�)!C�(�uύ��I�ԃ��q"�`�[N��!��a%�,Kt��[
���[��q�˨�7(Jّ9��+�(�P	�1]	3Ob�69��L�"��`S��'xb���,�^!�Ɵ�.J��1���0 P[����5&H1W �W��J6�=�z8��h
�,˽�~HM��|��֏����p	�H1�t{�eX|i��~�'��uw��Ղ�5�	)yY G6�`�/"A :7s��4��;�7�鲇U4i	�&O��S�W��0������B�u~�TZ��R�g �>�\!	�K�w0�\�X�x}�_Ay��;<�, �g�J�e�T��]$F̏/r�%q)|���8��W�FH!��1�^�4@�P�NvG�����W�-��z�%"8��1�0�x-�m����j*�8����ހ��!H͸/G]�m�,6p��3f�Z��qs��,�q�,�'PUn`��lO��l��廧�MD�1X�0?"[h�p'���j�+L�.O� ·b�_&�1%�1X+����) hRv�K�$� lC���nڠz��^�S���C�1$�]�'�	nh�_U���Z���[��S��R\�v�p�B̠��o�|�Í%\3�K���] ��sX�� ��3�ᩤ<�Vi��]BB�Y�o˪W��P�Dn�}̷�́Q5:���נ��*�<LZ6A>�Iz�J���
�8@)XV��w��U~\^gS��a]'X{�k� ���u}�����5B����U�~�%S@����I{d(�)9>uFc��	�������(�Kt�X���t�ebR&[1���0;ň�m�=��i�x\�2c���4��)�m[���}D��`ɹOS*I 8�s�)���<Bx��Ui�\�߅�	[���]�%w��J�����_B��.�}�,��#Zj�z�V��˸���X<�Zp��MȮ�%\�J)~�$��/�D"h	��FUS�b��ޥ ��_Lx-U�
I��}|����:����A����09"�2�lR��) #XQ�
�~�8������������+֜�U�����P�&��k}.�0���� ��[F�Ɲ�QR�#5_:�	~�δ4����ޗ��� R�^X��K1�M�n�5!@�}���$�8��%v�nć	 �CY� ��/Lq��l/�)T����P��B�e��8�16W
��	��Z[e���b�XvX���:�w���a �ZQUW�YT'R��XMJb��h:��JV��3�t�Q2j�XШ�G�<�B�:Y�6qH�S�pI$�\E@���P�k�*L��Nm�^��iY��r/���ф�݄���p'���~%ߥKb�� K�>҃�N	�>*Fp�' H8@(0B
�S0�
����0� `�#�R8�fecVV�3��d@"����Dc!aq1���>WI�h1R�*2�A q�h��Wg\z066��!��"~��D0�H*��x���N��N�8,��n_Hq��TP�3�Z�V\S�L-�	W�K������8�P��fMd�,�� �^���%
y\�-�{����"�|[^�����O������ح揰A,F4j�S�����)�
��O����Y�K��Ln8դ�f�p9U�~ 
��J�ga�hA4:-�z�à�"�E��>i'Ɠ�])V^�hMU��@�*Z;
�[����i����0w�@!�+�d��ׄ([#K�:!���o>/�/�T��0:������q
�0�%壏����|��^�m�`�~���+��kQF��-�����*�!Q)�𦳕r5�J�� ���:m$h}P�0A�^	�|YQ�: ������IP�џ�tT\�}	fM�A>�����?�)�I.��d����[�z�Ӂ�r��v7���B#�����~��>�X�(�,	���#�Sf|ok��P�b�?��s/-�P<B4�S���- O�N��P�X[�_h4U02��/��,�	�{�Yu �T]C�QSt:��=i�<x��)�I���E��_�AF��+�\r�D_=��
	�V	�X�X˖?�ը��h�Y��UVP3XWh(_91����vd��/�� ��AS�~q'1�.���3 �R6P���!�h*����n�|���'	��2Z�=Ԁ���	�]�*��A�W�q����$*�%�+���hpzܜq&�U��o1Qz�b�����	��)�D 0e�d_�Y�p{�,�K �A3UL](@�_��j����-��:z��J���h2�dK(��w?Z�d<�,�M��r�F
0y��%�)@�8w���s9�5D���`��>��ԣ
�I�����Ug֧��R�}�f R7|��Z]�� �y��^�����Q(YrM�����P*�<��N�����C��|#	D����[�Cfh?�0��AV�I�n
^f���[P��-2�]�)f�C(Ҽ��٭�U�R ���7i!��~�-����|^�$M���@v�x��3-1)�f^VV��4M��
[�Ϻ<�PB���U�C�f��b�WLMh�G3� �]�E%�[^7��lT߅S9DЯ�	E��J�Ey�\����~�ڠ��I(iXK�%��jh�b�7W� TTwன���e[	��?6-��u�����,,����`ѿx��ٲ���������R�������X���$0�A�ca+,_���v��e
j�s���HlFu��'�8p��P�>�]�<�8�yC�P.���F;� �L�If���-ae�$EX��8�Y�0r��h�/�:�9�BW���	��Sz����R�38%^M@�sP"\Ju,�g]��-3yW�����m���b|�Y ��se�cV��h��NZ��X�4a��n�!Lf��c5�
%JPU�}��!�j(X-�<b#��i@��d� �ݸ{P�0�n0Z�V*�C����A� �HE���a�4)χz�_`m��5��!\9�{�^���Ь��,t� Y��R�N��X�u��J�E�,���W �zg*)�'O�1���W�k�f%:^Y'n�k=�C���B(��'�Ib��`=�����ϭ|#�_�d���.@�Aj/�1_n騒��Y	�B&k/2	���)'բ���%�-F��7A�XA.V�Jڜ�)����{�U��xU6�8�-�@�/J�>�$:ދ�]�|�"�Y��N�"�(�f[yE���	sY��0?4Jh�;B�K� sq�ʜ�C'z����a L"��5K�`002_��'A)T��\�g]v�܏��[Đ[	�@q.%\b��n��-���<i��b�4ug;	��r��-����M���m�@SF>O1[ͪ�R0"B�
GwI4�y$	[�-�f�+��&³� ��(]�}8��K#��;> P� �u: @r*Q��������D������HX�������B��i1JF�`H`-.x7]��-��ސh�R�M�'q�^>�2� �S����s�2Ǻ�Hs��v_�㜖��a.��V[E%*�Rq8�>v-&�t�E�C`��N0�p*,#�[�@r��D�%��4c�fjd䩻��8	���|	��7����g�ϐ��|	f��~F�X��h'�V��C�N^�m58�\�A_���`���<��ҁ_��=����	��[��(�8
� -f�/�!��]y*ru徐1��S���c �2�,ѷ����.;���`;0�,V(�A�ß_�e0�A����;}9�C�N�
�̅�тuZ�	IB�$>8=_�h2&i0���x|lp	�aw�g:�4�D���OZ��`�-f(V|��,� ��b4
T��v��L�H�7�?����� 
򙩬�`�g�:�=Z$�ʡ�I��Y!xV*\�%�^r&���$���{I�	� �f��h	FQ��p�" !ڸ�w�G� �5�Efu'�� ��-�UXu?D�XC���Imd]�5h�b4��r��%�SL0Љ�>k+5o�1����|�/��_:�Y�L� ^�)^�;����#��.�[\ @$o�i�0<1�5y2�����_��*	s��&���X��p��X����o�0y���u�=H5Ke`91\W����@�3H*);ϸ�����B�6�������1����X/�O� ���Z�����zu	��{=U�Q&�� C�e
�	�W�
0�Ss�"������!Q��5�y �\`��IK���fjN�7���H�}8�cMY�T%�&�
�V)�q��_q��5�Z�����L�h��?o
EJO�㦎�ٗ��b�|(_d��Q0�	��|��hS_}嵄�����Q�x/KC��O��=��=_��Y�K�u�o�i����N�q�'y�7p�ݗ�Ó�р+1ZxA*�v1�V�My,Q�JH�j`Nq1/���'�֤��hK(�����O/�$���D-q	$XłR;52Q��X[�bX�a3h�a�1��W71`!�`� ��yE\@`4���^�@QKwO7��w�W0]�X�	�N�uzӂ���
Zu|��Y �1�f�ȉ�[v�)-т�Ih�WH]���-'�K��t_`�V�dR�X��o�)��@�l@5���.�O/#] ��bh��Da`���. Z=����?���hF/9S�6��.x]4>!�� �Z>��N�C#aOL)�����1`a��l�oX�Y���f�LO`���iHO�ܩ�o��&Cl�wͺ$����j����Wg�wC�{��5�[J(��9�=!��G���hR������d(��� ��N���]�q������",���źK��̀�&?� 5�ů!�]�1�焬l��[�	�O���ei�V��j�����y�l�#�Ɏһ��[S`W��hY��-�%�$��y�o�Lp�ˢ\�db<A>�~(��0�x~�y[1�z,)�;z-kq׀���ſ���� Sh�uPX�3��N\剴iڈ,ߑ��������Rh�3<��N���-V�)z�}���\\^����`�o
�]h�f�B]Oep���~�^U� �-+B�1`(�fX�w�� Ci�.�7@~_�༂���I�u�� ��u<�x���.qG�Һ`|�������1r��0�J�a߄���뉝{��]Q�L�f�ĺ�ņ���PS���<ZoCA_��HRJ�ǅ)�?i	�\�T�v�}H
����'h2P�} 3�m0�[(�Y�R��ۣ�]�8�K��c��>�O��Zhav!8�#�M�@ص��I�z��.N��7�H����Y�Mhte�_�RLEy��U��6�2T'fr�X�Z��G�|hq�z����UL�K��0��$K�8&Q��BO��/3!"׈_����hfy� �ΐ�铈����N��-�%!R��Q�`�ށ�@�K�N4���N��1X+�
Q�]��5�.+��lE@�1��"��V�;$PD]�6�i+�֭���xT-T�f4	�pr9�	�]����d>ʈ�����:�6[E	��.��N�hZlM�����&
��K���l����oO���8Q
�fw�p�k��G<�^�WAz4��xX�5.8����7�YK�(��>�#���E������:�/c\|!]I�'��%0� ���e���:/bW,�a>��J٩��.)Ib���1�.�BL��ܠ�!b �HYX-NQ?1V�Ɵ�N%޻�5o�!���3ߧJ�
cK�׫���bʴt^�`�hI?�%��K/"�mz� ���[�N�N���`&���Q�m~w��;j�9F���J���h�
)-.�S-ZR{3 �Vh?<yPd=�Y��ю,0cpC�D��O�*/�N�9Z�hv�$+Ư�t�)*�YY�M��TX㨇M*��rpD��c�l��&>��#Va��+[_h���	�X����-#K��	)��UL=JP���N�9��e����YK`|κ�O!0�y7\#^	��@��%��?xE����-� X1vz��E5�]&H��^N�<k����൸��:�:��Ã!��1z���L	%j^������(���%���� �������qO��3�lf[Q��]3m�U����KY����Q�{颠�h	d,
�����KT w��Y�y{C����^	��t���A�X�� � ���H��W�Q�';�9/�Z�ZW]g���4���%�ı��N���Z�/��/O�\��j�9-1��p�>�2�^�/�^���s|��lҀ��C�5=�4�!����鎠W�>�5-D���x��[�Dt�H��K���R�]鷙8}��a*a��B�)��5�8)1:�)
*���?"�i�;�[���	�o��S%�'��R+�� ��-eH%���4ˉ:�g�̥@���~?��z�T�C�P�ɥ4o� 0v^|_X��H��P�=`'�ÆQ����<�{@b�6!�;Za��pm�X�z|R4P����E�	 Z�ud�$�|�̹EIGp�0k�z�`�oI����J�BAj�����|���pd��ϸ�;�X�E�A` i��n
E�e���	��I�VL%�/^����O�QS����3!N(^���&��I�PT�yAz�7\�5�\�,��@B�ަ�<S����_�O?�2�`��i	B|�$�������u��� �p�O�-��x��0���=U#E{�1Y�,�:�q�l?��_]�� !ú�X��t-�	�@���w4�/�1Wӛ�;��q��kw2���\
��[Bt�� �1z�1�I�T1����!�@�8��B�i���$��h��֟L.5:�X�/
�X�`U�ɂW����ZYRF�'2��{�(�Q����1� �[씱��.�/��bW��]�Sa**�N	=���(���(бr�����
hM���
(����Hf�tL7 W�]2�k� �s�0h3[��6&`��X��YQ��A�O��Z�1wX+��0�8�	�́��D�0���;�5�I��-i���H+N���5Ig4(ɠhZ�#]�^.+_ޔq�[�쒺N���5�7��9Q(�Dx����Shc#VRJJG v�Z9H��27PV���E��|Sh�p4҇�7R��OcH[Y���U�=�j��(���p�1�`��x��/��|i�t�nN	7�+�	��	�'y	:��P^��Z QhJD��N��z]'IwSH-v�E��_�%U��^�I���A�v[n�1���鑔:^�6��>ʰ��^��Γ����
�J�9�_H�!?t���	W���U}J����|QE� �W��-��+��O�m���K\��Ӊ�T�x�� � �tKX�=%gcwȔ�p[ƃ������{%1�h�c`�F���j
&�,�� G1w�(9����/��r+`*�HnA.���×kK8~����ic�.@����w��u�E�����DYr�/�@e� d�u�q�w^)�_��f���W��	���wH��0q�h~//�P�������F�!��z��R�Uъ��0!1@X�hIR��:��?�o�Vֻ��� R$H�`͍X�L��|���4
���fBܬ��{��-w~�%pS�QحO���ڝQ�`��?�x� hT�S)�^��-�{!����)�nx�[�f:!�5�-�6@�Z�4K��V��D�	�Y�0������
�@�� �(�P[�� `� �la�8��>)�NY��PZp��.Z�N8����@�(�i�ò_ >�U���1��򣝐�~���R�<���M7�`E"�'�@����?u����>�02wW\7D�β���ȺKX�[\}���b��QX��;����U\8�s^����
p�aF�N���{^!���WqkW���$���,��H1
�S�4/�)~���5���T�')�����p�CaB���ځf]1�:�+����l8@��
2��WD�"�N0
�O@�-g�V�u���_��tM-IW&N�0()Ǿ������R/H[�QXP�D�+�xY[n"�&5^E''��~�b���������#p���;�-4Ǝyo�E�C�S��D�	���@B	����~�5>��`:�;&=����{��7rj�j����)��O��� 6�s7oLJA�A��!8#��I�zĿ�E{�˱�ؔ�y 5�D�A��W@B�`��)@��a���� NZD޾>��=�e�w�#�1���zBm�xӧ]�h^�F_�.v�t`�#(1�.	������#�b�ʬ�P!��X,,f��)ǀB׹k.*�V������
�=���/���[��������!0��5h�zO#](�[0h�<G� ��H9Ĳ�	��a�_ة��7�\ ��bL~+W�K���M@h�J	Hb�e��A�[fr�.�D�K�!��Jn�Q����v ��~-U1\:����"
�c���,!i��Y��0DL�	ØWZ��dKN8�&�ˋ�O\6t�o�ۍ��*�0�(��_Ro�"V�+�W�/��U�Z��{���h?d�i���c���3%5�`Sh �4�aY�?�r�uA�+�:�ffhj�4R��
iZ�����l�:�V��8�\$�\ch�.���H�?��°��
�*�xWB
ĞFq�M��(�����j�� �I��!���< (�8DO;���>m,~��*��KKi������\��K�������E�Pr%C�3���լ��N����[ͩ5�u�1 G���Y,���V	�.�|���-0B�1��3)=?9��\uK��!
D*��^�C���ì��(���ߏ��I*�ZK�0����� �Y�I`+U��<e]}9���"�~.�v��2M�p��z�P��S�I@O ����*��vm0�S���N� ��h�<�T0� ��_İ/�	�lC��}���u��C��h4O"����K�
X�3���޶����l��/�q���~��~�����5r�\�ף��^+{�{���W�\+X%΢�\+��v6��<�V�� _�=X	�2�3v6���<v(V�b;^)�l�1ڻD�e��L$֯��
�_��V>�wY��"'���:����(�X�/A��+#��X���i���}��y~k�tX�;��`I2�T� ZC�c��}nH(q|0�"�}��O �*	<����M���G�s)ú��-B� �w�$7��;�%'�����h��2��w�i�밃10�]��ÝU0Ѝ���ڽ�����ݰT�> 
��@6�^����*��"� ZP�%O�E��~���+��h�b|��Y�\W�w^��t�j-~�Wh}j�� �W�K���k�I�P���1Ų��R/x�F	&+:#���D��4�g���"z
wV��т���N!X����_�� y�$��IDAFI9�EoVG�1�x.��'���;P/	I9l3��]�O���&1�RH7w+��u*\�	)�W�}~*���~����_�Va7�9.��fxNR�ȋ����{)D�2�8�|�f9h� �k�<���(�
L��!�f]9*�5��,{K�8�]%���m(L�Y6	j��hn0���-B~�1)�E��u��Npd���\3: �#4�Q��8�)Ȑ���0���+vlJs�/ �5�Z�!ZӼ�$�~����YhRAVW�6
Yo���c� f��th�̜pN��<Q��;��%���Y���Wa�x����P	/��)�}�r�'���V����K�BTs/[ck@���V�A��'{M.l��-�(h%�K���,�&��	 b"A�`�NY�߀8�f�[�,����_���:���ň�D���8� [h�����.^�@f-��Mo��啀���D�����tfU韔���Y�uZ����e����1�i�Vp�0�}Ĉ'Q���H��	�^ȁJ�
<a�*����HZ�/�K���P�Ǽ��]��񷠕��s3-�}����0�"ԣ}O\���+-0B�w�\w],k���N
�ۇ���Y����Ts�
�kk��� ����P�:� 
M�
�E-z�� �'^"h=r�"1���
(�R��	�&�ǿ�%{wb�W��f�F�ZX��K]B�Ý�}�'D@�^E�� ��9��?BJ׭�3D�
[g���j���5;?1�Y�rf[\�&?p�߼�Z[������K�V��ͺ2[m��v5��ѝIU���z���m5yV�i�+)�^*�,��0	���O
�\�C^L� Z��z���&f���VP�GB�=��EV0&m�i8g6�g'�K����r߉<�s2�n�S��Ǻ=�|9t�K��X��hL�&`�B�!(S��;�P���	�Q�X%^�+�}��-�#����1�%��9	H��������)�&�-�.���>GM�]h�ųML�(y�;_�_�$x��Ԥ�;�L�'%i"j� �	��ń��>�~pI��D �'����vqP2�"�?ȰoY�!EV"�.{3��	s�g(���jT���e~�B��m|��^���uŮ�-!z���铋��ȸY�ph�!�i
�?f�	@ŀ�����@�z0\!�7���)�j���S�ʹv�JP��J��B	��S/�ܱw[�����AjW�ؤ��w@���׿`'���T9�'(U�*s
N,�˻e�}|W�h�;~ �Q��b���f��2�y�`�1mEN�N�w&q�R����x�~�G��,�Ȯ �T^�-K
U8��!�M�'Yݺ�s�O5E��`H��U<�� 1�-dD��@�����o�h��p�]EN���.�}=�.��p�Z�͊E �x��)'�XZ�hN?�D��o��]K͐D�rW�5v.�lH��� '�Z�P�h�2��WK��jkKX�ɕ
�����d��g�kn�������� $Y4��tO�!{7>�	}E-&U�$���;#K�T�B?�@.�A��4}��~|�!�kH�\e0,�� �!ʽCb�z���)��4��Uf!H[��%��+D.�-XV��Wś3�1�V��>�}.�y6�G��a�ɉ�0j|)<�X��z�h�JD��b}z�Uy;H)X�4��>Xs' h�#�/X% �$}|-�	���5 ? f1пT�QT��z��̎	�)���.kW���h�o-~��T���@u�?�[����?S>� jh(���AMH�r!.�� Uh9sNX5-8��[�e&�Β��8���(;�
����ˌL@HV�S\��2&^W �V���}���W���K��t Qˁ�e_\
@�MA@�f�O[�(�/�RT���8pZ���h�-�̇�!�2�_0�\�K	���=K��y�ZZ'�iД)���@˧tb���)@�^�|�������4�.]�RD+�@JGC=���sa���k�5��1����
�s����������ڛu �"(г���z�U0��
�0���P����=o<ꦤ	�j1�m��H����J��Qq�>�)�k��kE��� ���|�w�i�rj�hbK��-�[D<bY�3}���t��������`0ʗ�w��r��˽�;"}[��Ə��	0� �|�[�SH �����b�A	��>[Y�����9š��|0�
 ��\���f�����2�n�x���X��1�x2�J��AZ)>��˷��o�����g�a�����5>tB�ׄ�^�Q!2���-��G�����	=�f�L�Ak���jH�#��J����_��J�3n���m��`�6w<*��!.�2�S9+��Z'([�P��8�{�t.R?�@�~�-���&�W���O�U2�b)�(��o�A ��w�>_N�%��C����Ϭ�tZ%Wp��jF_A��!b�h��4 ��O���Rҷ_��-k.U�	6���)>�h���g�1˫Qp�h �V pY��$nO!�eo� ���A�|5n�-��~*%)2�B�|���_��.p��
TVi������s�u��җڮ {G�)/1^и��q,�չ<�aK~lCݩW�.T�4)�vB��}R�<�R!�°�}][r�dlB�k�Q�7%u6�����/S�P]��Xm4B�a�!VH4�@o`��ѐ��n�ڠ�9[�;�l�I�{$+�5�H��X�����;�p.�F�YӅ͜�hDYW��C@j��_$�3)��.��D�|l�\�� %�,LO@	-n+w{1����g�!b��/�Z 
��Ԥ��O�c� ����n"�1	�m)�hSuNP ?�&f�O_�y)-)Z7����Ơ��Z��<�`�p]K�����W�YayX6�ݿ��/W�,�Q���9k��З.Lm� �(��M�S�? +5yh�S�X�ؠ_�0���V�� m��]���YC�1o ��R^��0��c2�~/�����GP�1'
Z|�POI�ڹB]b��tN�@��f%?@�H;2Q�T]`n��pF=#�Bys-�a�;kH{�A���Bm)�����f���u�秨B*_��'F�"X��)ô|��� �_&���`����	/7b�U'e��h�u���>ı��0�z�R�W�C��O����,S���(H5���!�%jB���^{0�	���-o�v/ܠ��y�X���WS @t�5�zv�O9��t� ��A�/4f�0��`���b��4��;��ц�X-�	u%tN �sb��q&�1�^$ A�"��m��P`MI{O�oHLK�;�]�v
o��=���^��VZh��W�_�5�N�A�1����L�8(v. �6��L
�D���T�)B��%J-`�
�JE��H��Y ,5�
5{Cc��5		ԯ�T�K	�"�Nuu��}	��O�l� �W�~�>�J��nTM��xP>6?�O\8}
�{�'�X�g_��!���S h�R�8]��H1*'����H?Ό�?	��$�`ͅ����	�Z!VŎ�-����4MZ؇~
{n�{_YU�^yo-cn��D
��W��V�g�ϐ��Vf���ӗ�������T/�"V�b��wY���6q�����	b\\Q1��+��ِ�AWT:�`��O�<���I^�˗	-��Z�K ��u4�S���Q-y�^ �C<yR�ZH��K�����_1�}����idG|��\z%'���D��	H���L)�%X�|q������
������!_��}�,)] �LJ��X)�S]��ًZ�bE� ��N�\q/�=�`#��Z8�h)�}�D����!g錏.�	x��Qh{�jr�1���9ZA8,�h�'� Ͼ�PWh����M���/Pݰ�S�Ð��	�1�* E�Yg�3�I'lA;�cÎ�	Z1+������C ~S�f!�h�Z%׀���N�VءF���fB����i�@y�_�������r-?t4�2oZն$���9~xnP�P*F0�
)�HܺJe�iy����M��	A��	��'��� �L)�>�߀hI`�,YA%��@-�" �.H(q�˰���xp�< �4XI��f'RJx-��t���pa����u�V1�'�~��c�Ӱ� Sw�s=:_��x �]�D5�Eǯt-W�i���Q%�/���8�Kp��Y(�������_Iۤ�I"}��b7�=!���X'(/[_6�'�A_En���0��Xv)K�:/xS�VQDBGU|q��@���m��0��c	��Y�N���)�1яᦖ�Z��,�� ���V8[K����%w@�m��`'�a]�/�d[�_Q?���qK�>`�p��-�#X�Ĳ���A)��1{�_���T,0^���` ��%�8�{B������W����K_!B駰o�)
E0��>�N�G��v���H��y���;�=x:q��I{�':��ӽ��.C�$~����k���}���s�0����8�+=��M	�,+�_G0Ҳ)^#�����Ϧ
�?�*��1&�-�U28wq�k@�f%Az5�	���r�A'.b�!�f.�p�UhH��y[��K���Xw_%m�G��3�R�2��������B���1�ȋYfp�'L���ɸS��-�U�Z �[X�}MOx����9m �� H�1�X��yh�o��& mS-Q�>T�!J�ҏ/�`#R�|t�@���?�:�)P�EV�Y�
�Ṇ��[����(�;�@I��v5v�A��R�R��J�.%u2�|���	﨧��2`Yn  wM�2'��Dꁫ&��}�Mx}I�����6n�ͺ�@���k�T�ҝ�hK�-��1� }Lt@J%IQ$4��	����^o.��g��; �W��
�^[�Aa����.�'��*�(-`]�-�#ҳ
qnRm��C��; ��Xb,h�`{2[vX��������D� �5&�����1��'�#���8EWH[�J��%�'����p!cIL4���1���^ �����z�tH���.#�	C0)�P�9��%��ȉ9��v@������?���#����5�N)�J��!h�$���k:�=�Zף^���'yC`���#�]B_ ��5* _~-�X�8�Bn��EX�,�u%�
ٴɜ�;GH��:�	��}�!����'��m �Va!�]�CeQ�,���uh��2dF���s�+�'A[Wrd-!Ys�h+M�ە�(�>$	<��@�2 ��N!g%�j['�rƲ�]9L>f�g ���9�6a`�h"=�����5��t>
��C����d�X ���3-�0%	(Q Y1Ż
C Zy��@5�r}.�X�9��=�w`�/Y:SA��8�%�J{2;uN����nXiJ�B�*Z	u�H�>8@��p+���CP�8�#*	՟	o�q�D���<@A������pr�o��sQ}�'?�:�&���G�6(�-��@V-cK��Jk�l�O;3�Q�1c!�:����A�ȒA��S�1�Y�@�'�Nc���j��^����g\n���ApH�V?j���	��ܰ�X'� �2A��Bf����h��c?oX5�N��4@⺛>�Ϫt�z��y�TU�Z����B2Q{u栠��B�����:ǰ�sJ3�!�_��ѧy@P�6��CNN�*�Y$`M�`�^YX�ʬ�/����^���@�1{�/Y����
-8M�<��\[�P͝L�	��	�h]j,��`HBY�m^���\[t jѪPL֗�/?�θ��X��hO	鲜p�9����P�; z�|M��G�t ��b�}��ц���a�0��|�]�#�Ը�|t�WV�}�à�]y8��������	}qY;��_�}3�\K��V:�Bʰ�4�)�,�w�xZY�,2�^�����<������zĿ �:_~P�q� ��]�O�T�@X9�P�- �qp1�hPZ!̥SJ�~���A���k�p���~��Ů��%Pݟ�FP14�y*�Ez2���Dj�%G������fT<P$�cs�\�"1ѐW�mA �p`�x�׃��0w�4����\�$_�5h`HpMW�?'�,8��tz�����!��>�+	�S��Q�tj�Y�J�fS�����v�z�a[2(�;�dH�"�ZC��\RT�n�U�_�i��:�0�<K#�9X< �L���
}>(ʻ��닐�!v�>�~�.I���6+�x ؋��)9W �H�z�P;I�*.�/�f����,^]��vH��5=.��02�Ģ���N��#�
�4H^r�̎}l)Nՠ9� 9����h�;-wq��S�!n�a1plȵP�/<LQG	#
�P�����Q����Ѐ@?�	�h�f���S'__�4.��a��/0{O �+BF*�_�GM��6�h���ָ��e-1Yr{W'F����iM`<N�Gxh�7g_���c@�0-:���%�#-�B�P B�-��X��)�� o�(�<M�RC`-�q��VW�=��e�Oz�3d]��"����_���,X�3!�X �֧ݩ��J�Ly0C��2j.yL�Q��I��T}l/�T�-U>&���,&���P�^-����[��Q9��Z�G�y���f-�K	���1 �!�=7
#�w`83LyP�r'�A��O ڍ�)ݘ�	]M{��4���hbP�f��#�N����{�T�'�?9�� m�~1x�	�BLC����O�"���QH��@9�!��j���@* �:T@u�0
ދc�����HVL���
���>B�[\�A�p�S��Zp���!G��
Z�OB����)�+����[FP��@(R����t�l��=�-&
�?Ո({�\��b3��T����4�"[(�~���h>p�� ��m&'�/R���q+��w��S����_ �$�A���!k`���$���٘o��M��w)�� 1�r�l�	�Q{
�b�C@�_K��_[PR��NE�Z,F�!v$���d�P��4CR�:$�,$�]2�u�ʋ���9��D�2"Y��$�E�'��,C�Y���1�_��Q �'�������_T�z�����hb�½�yL��\�|^�q:P,J��S�[��ǣ�9�����Z%���]'z��Ik�v��VW$I��-�DKVH�n�bK�V�5�z���R=�u/B�%�[	*Z��s-�n��t3���� �[��Dc�溃�z4�`'�0�L;��j�'�1��@����� �B"�\��#3?%
����_!h�\�nJ�>��-�I�Y��[j����~���	�^�(�����������ݜ�V$���aQ����p����m�Aw&o�}޾��O1�¶���Yܣ���K@�������[��)�t-��t�at<>m{�Ѻ�����kT�^�J/�L����Î��?^����5X���3D�n|FD^�T1��dv)ɒ���3��Ò��r���8�F�	w�N��^�����p[�~�$�e*�+�		�F�v�RB�q�_�?���b$�Wz���ٔ�N�-�ֿ'}\h���[���l�-��ʄR��s-�!�DP�eCZ����=Ш�a�D�wA[�a.:�oPY�=9���e��(T\�
n��J�ěx��$b�x�*%�1
G-� �Bx� �5tv)�8� Yh,J>a��O��S�e��F���Z�32��܀ Rh��	X[�U���%�A�@O�p�J�d�&�,������i+{��e8:W�sP-Sh?6ddA*��1H)�!̐6��j�8whp)���i����5�'���q���$��X1ʇ�WV��5���]�����w��N��HN���{�x�Y�B	�M�!QJ�\yUT��^��1;{T�#��K�Z�;��2��W�	�8��W���
Y�"$��	�J��I�p�S�'�3c��0[Z�B��輥��X\J�k����X@��b�OX�I����N;�4�3\[$t��S��]�9'T�Z�M�'T�S�cHՔv�Y���<�G���)�C��RvJN�(�LfA�� � �[,\e�O�?>��+���\�k�n��b:�`PBO.�3_�ƱJ����u
��]����n���-Q���R����3�Ե8EKR�C@h/*��τJ����Z��R�3[����a�|hX �wq�b�1�S�B�]������ ��=��w�WU��h�a� AZ���Jc~�P67`����P�A�xb[�"@�	�-W�i	��O�YO�r'�]�	�0^�DZ0�� �P�]��_q��i,A$��V��@,%(:铱���Sj�3R���2�cܡ*ӆ0��'�^��:�	������V	jS ��)�e-�NP9q�" ��d�x���%�@�<-�E�����p~�a{b�1��ຸ O��m o	r鈉޸��E�
]��f� ����)���
R�xGf�(�p+8�oJ�ݸ>�f
�{aCr?1O�d��U_kdSбFk��[c��!�_�V�p*?Q� �v���) ��Y!�K_�	�="�O�YE���ӯ��c>��d�	�AI�eVi�1�Uu��'NyU��]�>Λ�V( �N�+U� �~_L�p�{5��7�] h�A?9)]9�ځ���W��`�r�Xwo܉�{}��IQ�I�_&�!���ڸD������^Zm
:V3���ش�9�@6�+������e�~7�����c��2op*)�O@dp
��.iW�X8]������������5�R�'�`|&*�`�h|)V��	<*�Qz����8�p��KbǪ��(�Z��PR���S0��X�{Ѭ!���݁D���a�Ҕ��Q=�H�TD�`��+_`$C��U&?���+_�L[;g���}�6t������� ׀�.��0���������M� K8���\[�NQh�<�4O���ƪ��㾅�h[q�pF� ��/'��5AH�4����fJ�O[-��0��z�uT��F�r�<P���G~�50�W:7ŔY�O�G�p!��E8���B-p���@N��	gw�B1L���� 
�M`�-��vE:��.D�o�~�ErƨI��r-�fG+w�qP��1{�������@VA��	�o��A|Ym��UX���~n�$+M-��S�mu�v�#i�b�/����n.�~$;2���L7?&:�U�>�塩d3;���-�]��|dL�`��0&z(6�X�\�T�"��C.�ïp-�A2"�[������m�* �J�w� R�׺�0���M�`	,E"l�tq9��ڇ@�ؠ��{1i�.t �vu/�Z��k�1�#���� �)�=E���jc'�ӹ�����\H���>!˸�w��ٚw (w�;�w_T�N�O������c��������zm\W A����U����e������`W����6_����|�t!���t�J	������������KS��n����M�ѴT?4<�h10��`Db�cN�|Z 빒>���'0{;Q%U`}�r�����8h�O?�@������<<-���:0�Y��"�g4�f��xmo>�iB�~���W��yy�c~_5�1�hGc,��륊Y���$EL3���U	1�*�5j�����c/&�O�@��v�1��$�H	�Ђ��[�����0U0i6��[���%�):N�P�fӂ:
�dʽ ��h�p|�U�b��9u�0��%2�s�ӈ��q�h�M`�R~�S��_	�i����,;��������\}�<�5E���*�5+�8���8}6%�����r��c�m)�1�Ikt,Z���Z��_謰X� ���߰1�n�P�UE@���`Y�i�L�s�b)˘� +VIf��>�[�,y��-ZQ{��@�i���}�sE��pO���Q	��~R�x8�z"av+��z� �K�HJTS.�F���<7/��Ж|��.�),Ȇ��Tr`�X��Օ��đF<0� ��(�Xh/k,yl�Rb�H�L��q��~����,����f�O�U!	<��[�V(�������K���� ?���X��f$�; x�A�+%9W������'�Z��!�S���s#�V0�ІB�1�He���`� G�/�]E���{��E���N�^|���ub@ ��z8`}��G!��D��C�ٺ}�ߪFp���bM�O����,�Ud���px�Y�68�j��U�^�NȰl	g���գ,v����n�J	j�$����x�AI
n^�'��Q���Ԭ@�hTj��H^K$e�
Cȯ(�]�;)�[��� ��Ԍ�>�O�|�m@4)�ԡ�����!n-�[^&���>1�zHG�c'.�o�~f'Uh�,�k�D`[3�>����Rb�n�w��ARh�twz.B	ZS�0)+kA�k�����ج����wQ�P��9���/����U:�{�'Xi�����2��we5A�٧w���/�ad0q�p ��/�ԼXLC��X�`P��?S�������	)�Р�חT��H�"�0�R�X��
�:@a/2�p�~$-ȸ �)���@U�Fڰv�'3(��Z�f#0���*���-0h!3���MN4�|*}	v�R���y����F^�>q��<Vo���qu��9
v�{�cv��F��R)ÁA	�v p��q�S�N���^��	�)���_ �C��x f���q�r^g�##/�hGXwA@��)~�P��b�����Q���6�
��� �Gſ�W�S3�^"�����U�P��=�2�ۇ��0���_$�H�:��Vw��4�^�;���zR����vB��}a+q,Q1��+n�`~�dy�F��|��(v\|�:�Ax_DG����!�+`�To�Huk����@�('C|Z@ZjV�4+r'0�ߔ�`-�B��'4 �2�]�"G�E0�o�
�ב��j�,)	�][';�D� Q�h�>9Z���%�
m�HK�;XQ��^_�-�?��;��X�п	Fp��,�3[�:)�-P�պk�F��$�=� a�4���a'��o$��W���>t+@�L\��fJ��q~�v�P)"��kUC)غn�F��D?`)�^ּpɚՉ�U�ؗE�ip
�~����Q!�.�9�?�ꗸɂhV��rk�;�@.Լ����d@��l0�(3�Z{�HFOG��A;���Zm�EHe�'	�kb���]�*��o+�E�-)�!�/�����^�B~�1��ť@\h��̪�$�`N�}��A^��[�1�V��]Z�^);�	�3�G�/vQ�o		�m���0�p�JG	�  ��I X`����	%��+���RM��Hγuy$2��{��S	HU�_�_�%�����9�f�-�%��rה��15�6\S�y+�� �W^�<��;#|&)�O�Q'>�s�Px!�K�~���! `	��Bx��zk��ټ?�+�d����}�) k�Nd"�v �pf��ʬ��%XH��KoN��Y[1��- d��5>V�9�L~��?K��.2���r_m���u&6��UX.^���hO*�&B�%l	WPt�B�j�:�F�8��B�AW�z�����S�V�4C���K�̐�%�tmV(<u���qy��S<�Q�|!(J�	(vC�l*�'���R>�Ut��Ex����4��7ty��̴��q=[�u�^�j�\^U&��0���`)�a�>�Aڽx8a��E�gH{/n"r�]j�bQhI���1�xA��d�	Վ��<��Ú�*�[D�J�@ϼ���U�;�� ��h�l���)pX]�$@��N�a��fB_h��֚�`�]S�T�@�J @p�[���R�m����%�'��cx&����XS�0�[o����@�Åp�b����V�J ��1�$�|%�t�EV�Ah�9|����L���%�n�:��!���91�^��a
�ޑ�fB��VU��"���(�#J��q�F*5�;��}>Ϲ��U^ʯ[�I�!'X]�κ��C�
��%|�5I9�@>���-\��:���P�$��	���A"�� h�yY�ݽ�ս^���Ƙ���AC�@ں�%e\y)/��U�pm* �:@
�'��j5�lUu��egA�+�*�/^@�}[���&���';'uRB�}�:'��Z4H��И:u�}/�a�H	��6\h!SU��Ui����!8�w�}|����I�g���^'}]����A1�1�+��z�1]Qd�������q=vl.И�d���z��d��h�����JY�7/HUt��y [BR�Eށ^�1> ��E1	�r!�ݐY~z)�s�q� \��	"��s�Q� W9Y��0� ������glGK����^-����G O0���s3�_�����.(n��R俘���Z!7�z�S�?��@�ل,[��uI�t��CO�+@��%BJC��l
 ҉)��A�Ē�N�/��ޘb��<!�Xe��P��W��"je����a1>h�Gk�`|����q%B!�`�h8K-��+�w�i�] ��e
2/�@Ïg n~�t�J�����L%�]�:�ƵhsV%WoxS
��kbWE��N�,B���\�y		��0߂���D�:ɛ�RɄYU��	3�w a�C�:��$M8�!ߡ;���=$+�pI��~�/�up�]F�>�=�L����P�Pg��p�_�!c�K�}f���!����ȳPF
k�
2��Z��Mj��^^ԁ��(.݀�i}���m��	�u�B�%�_�V����?� ]j�ؽv mM���p\%�\�Z��
z�6�L4	��4P,4C��0�Ҡ๺e�M�n�`�ɚf�@��4� ���^_����-3/�cS����/�m>'�iX�<�%)$�D�[>�l�?&\\ٙ*�����7-&@�� P�V#��_��6|f��O���O�A4c�����å�jU��:j��/�8����1Ҝh)G���W�	_�)�����C@Sq)\M�`���?0p4���X8�$w=-�W�c�������ͿX�F��0H�p��`��F�^;�w��d��r9�0�-l��	��! �;^%�~	1w����X���n�_����Pһ zw�}���:�E���P�@5�Hc� �Jk�Cb�w�]K��B8��
��qY3~ɹb��kE,VU2fEP����YX��t[�~�ŗf�Y%F�S�a��Y��Vz}��}��|\ P�Eq�|H-CZ�;���%�,X��x(P��Ц��F�Ӂ�	`���T�%fA{U\Z���,�oIE}����	>#)(~	�<�?�_,S'Cs�5�* -�C�I��	�~eؼ)����n��<�!�f�'��Qe���d�]�
�$��Y9);�]�%�U�J }k�| �-�(
'��G� j���ր/ƬB|�y���p�a:J��pX���_��t�G�on�S�	�ǅ��[ �Z�Ra+��?��O�eM�����sSgc��zb�_U~ty��|��u��mI.���e��&+�+�Z�]YNA�\*��^�@�a�ɜ!ٸ �45�+|Oj�^ހtDuz1�	�0�	E<\0��"����)�b���_��hS2B�x�,0�	p[���noU{��K
�����n!=�_��Y�����<��F�I��X�TXk�^�� �-�+�<���w��QR�*�e]����0�02%3�,S�- (�Odw�`٦)�� ^���q]p`7?t����%�c�Y-Kv��6NLMpb8��h>N~L�t^�s9��kOи��~M%ȩ��*�%9�tB�U �_�v=���!YA
)���:l�.T����p��1�^Ul���C�.1���O��;^�zjNW����qyޠ
gOV�&&LT�4��PmX��7�K�7��:���H{�W��L	�a���1'��� .���4�3�z:�`�h{��U�Q�����F]�b�@͠�$M~��
�1�h�.�2���:m}��(���z�/�	�C�/��e�����'�b���U�S��f�r���+^�QW�*�@(�5H�L�![���UF۵c���V��S8"~� 5g9���d�N��m&!�fX\��J��P�����*4r�J^�����J.��M[���д/ݠf�I-P��Ð�,�L�8�N{�}��%Qghz)b��A���	 a�oq�+�U���'Y�r?�#n�ܛ��s������3%��w��8%#dT`R_y��!��A�	��u? -yBX�Y>��>��������`��p 4W0�(ހ�%U t.�[+3�:�70�Lo�{�5A���UP�02�%R3�Y`��J6��T0�@LV�K�"EA�P�:����>�	����U��%����V,)�S���5�$/����圉oc ��5�E-N	נ���v����`�]�;����f�L�fA*H��I1z5y-�0j�P�4 �z�
5��'�!`�aH%�^P�[I%�w_aa4**��:A���4��/ �B`}�__ީg�a�S].�A����P���>�3�$�t\� ZRfSP����en�	�[}�K楠���=W�I	U{��«
q��-�f���j���x<(�@�hn=�f�VI�zTߺ���@�C� �|�A���bY ƴ� �6�S����BIkvL��� rw麰��!�ҙ�1Sͥ�ާݗ�-��+�w)"�:^�Y�|�$\�TA���{��BEU��`<��� ��.Q>1_ٮ$���PfT�`�kf�)_ٺ�[Z�d�!�(�O,ژ_�p��N����5�)KuA� ��1��%qj�5ꖄ�J�Ŕ�%]��`@R9qP�CP��!1󋏬�{�&� �o�h�l��}8Ny	uY:`U�6S��Fx	^?\[GC����F�0
 XQ��e#_����=� �"c>H��u�]���Z�b�s-	�!��O��R���k�U�M�ό���zr�n���-�����o]@�)��H������QSY���"��?��C;������n��
y�<Ċ{���� ����r,��i�/�0
�ǚ�!��3�`��-�vv�� �)���_��$�e���}K���י��P� V�KF?�X3(��:l�+Un�e��Aզ(�I�P:� �ˇ]�s�V� �OEh��I��&ZN0�����ɀ��k����1a`IC8�0�/��.BV:P�HUxK 0d<[O���[Wf��O��7�<cɎ�\0��YcP(y���qhVn��H������8eA��SZYUhe]?!薾9���C V���H @-j&�75�<3������Z}LZt�c����I��f��p���?%0rnO�*1��	��1>pF?Y����F?0јs$`S��(�[ �D�0�l.h�`%�{�\K����'P=�y�C������<B��=%)�$	�p�%{$:N�ZxW'�l�&h�7����~SJ��+!pm�\7�W����|K)�ۊ�%ގh��! �TF�c���@i�؅񙬬�5�#�A���U,9ꆗ��L��X�:� �^���PW�&p}�O`@+1��� #	`���F����Ѻ�����R�#�^26���1�����_M��W�D�)Ld���_!�`�Q�Yf���Z#�	U	wV�����Z�#��-|@
7X��Xh�KC"���J���*�<|/E���f�[`7~	k�^��a>Ŀ��T���Y�o1[�����/N @��@%�7vq*�H����I} �j#9��gf��x��� �1ؽ�AN���3�A�M����`�麽N	�@޺�ȱ�L>�-�F�<Ce�۽��lE��'Pr�k�
o�c�����S��Ey�Y?�S�uJT� g��+Hf~�`J�b}����C�E>V�.L�	�l���r]3x��`���$[Q�@�rG )t/�.�2v].[�	���.(j�{0��i\��c�S� �=��t0� `��s 5�d�o�����w8�"�'��ѭaJ&)��{�;�;�]��Qx��� |K���XX��`��(.J�+-
2Xn�fS�ǻ���锫�C	�,x#������v�/�E�f׮�Y�D�7�k���){�%C���Y��4���-��@�~Q�X�V$�w��3H#\N�x�ީ�Q���Q1k`.�)�T���[;�æW�V��o��9K�8*,�x��krzcَ�D��M�����bTF S��?�k�v@*�IR�A������`��)��ڕ������K^e�+��/c
��|�>I��6eC�^Z�n	��#Kc��)7:L/���X��%vC,n
�羣��X�G'��Z{(�_/�SS1�������VT^Aӏ�<R���y{g(�K�� 0��;��5�H(B�v��3��2�Iv����3���W�m�7]Cj�j�ԦI���$�� Z��6'�8,��/�~���>}) A��V���N�����)��^/���{|Mh�BT[��ne.�Á� �4*�ʿ)��<U���-'�5�(�S韃�;�	�d#�� ��j*��1.�Y��ܪ��/�	w�.�T��hI�]�O���_	P]�yJ�H�-ZT�RU<h�^�L�IK /�a��@�-�T@fh�>������h��Y�=���r��X!/,�펟�D+����QnNbDWF�&�%���3����Z6	h��v��ߞł��'����, *Y,��9>M�����镈�1����[.`�	�ݲ!ܑdZ·�R�G&�06YF���H�o��;{�N��Z{�X��t��gh Sq96�(Jp�|�� �S��/~/q�
X�!�>�,�faD)L�<*Z��9{�-3�ؿ�Tޥ�>�ڋZ[��J��}�!�X��Q��/��3�9�w��0K��	�BH	?�WzzO9f>�>�(%�mW��q�h�b�sV9pti��|̏Bb|��@�Y� !t`��-�;��#B�\43X�J�r���cN��|�`T�d,!�ܐ'�zjAX*	�a,K�b
�m�7H1&�l�������ܘq]���A��p+ U��AGO
�\8Q���	�$�<p�p�'؋@Ɇcj����_�E��0SRc6(��@��BK��|�ԗu��6i�H��	�ߔ�gJ��Q[��O��BJ�:�8Ì4�7���ɯ�΀��)h2���*:
X�?��:�+�qM~=HO���^��O�c{Д	�?_�#L�*`���Û�cX���Q�5Z�A)^�rk�,�
M��S+	�]� W+�Y��_�K�W�i�q�6�$�	�\���!����XYAr��-�m��e-h����-�2ZI�~�)f@� �C�6�㟀� \GB�e�,��8��4 �xH�72i�r�5aM�n����F�D��͂;�S�� ��!U[��NV� 3%X&'b�h�3��.��Zq�`Ä!8�oND��V�!�U��EPH" ��S�
`wOh���V5�&!��;�F���4�\����`�=Q������ʒ|~b�Y��פ"��O���#+ '��0�J �X۾����%$p�#��DJ�d_w��${]�w?�_ ����X^wZ��{I���si��T��� ��|�'H�?o�"ԑ�Pb���z��^���iD�1�/B�2ý&�# �>?1U�S�g�����J"�J��[v+���XbvQ�z�"��������4r��X[ fYh>�;�+��H��-:?�u	|��MHOaĪhP�� �[n�k)�h�*֍�+"��84��7s�`��k��
�hq�V8+fp��S��ʧ��9�?����;���?�1[h�F�G�1½�1�cU~zoE*����h�0�|0T���*�#�?����� �-h.:�	r .hep�({Z��=	��M�G�鴃����6.��
8D��<$f �=��џV��]�2p	��]�w����0��k�\����!C��a��S�Ő�ƿ�xZ��D��2{-�Zx��`�$�6�@>�.X�-�"��^� �1�-�5[GhC�0\gv������0*�2�.{�bV���,�	HW�c�w-�FG|{���	�0����N�_�}�_M/�RK�$�0h�\�k�!�)އ�~��h sG&�*�U��4�.O�ѻ?ڗ��v	]����jw\Kc	"['P%[�$ay�O�	�ſ	<��iT%b"��a���ө@�MZ=�˰�Ld8�U�f��_�`��WZ����h*�.�n%���2�����ά��8,K3 /1��<���n�����j�Q)��?��4�6�o�C�� Һ�{���Q�`L׺�W���#DN1��|�U�� 0{IX5�!N^-���Z�mbNY!��
/��/�i�n�b˽�Ť �OX@d�PȀ�9:�P�R}���`"z�	[ WJ�v���\<�}\�@U�R��1�}�y�M��HJ�t(����If�BRхX�oH~ ���_(���R%�.^�$�|�%��S�"!�K�N�����+�} R�Yz+�A�Xk�@��#'�):��g��u�R� �j�H(����N��E�|'�� Ӂ��it0�x/�0��d��
��}���1�}�"��Hq p���X�����=��yp���:�}ߍ�).-Y	��w{� Q�3l�
��xdZ����2���^� q��{|�����*[��L�RXHZ}����j�7^��P^������=v�ʠ�F.�B�+y�v�|���[r	�ލ���p��J�<yc z	�к��*�y����Q��2_?>{�	!�s�J	���ۻ�i�1u�J [�NLS�� �ʅ�v���#��TDO��p�f�X����qn�$1^�T�`w�y��V0t����w�	�N�MK�ނ@PhI~7�6��HE�A?��(;���^�sN��8l8��8gZ��Ҽ�$�8�JA��C���\�p[QU�9�F�S���X2> �$/��R�������������N[����$0����Y.�'8���X�0)���'Ϟ���H�>���,	\h>nD=|���Pp ),	Rw�%Q�.(k`�� �@/i�m	�H�W ���U��I&�yS [Fmo��&(
t}лN� amQ��#�������n%:U6W���a�TPཱི�H|�%���0R���`V �Z1��q;���(-8c(Y7�h�,�򤣬�t(��(�[�Ǿ��0��'�.�H �_,����.��M��0?�3h��>AQ�܃�8�v��|��)T{2�ZUO _f^�w:�# �cRKJ1�)�-�&��_����+�t��[DA9��Q���c-v^Kꪏã� Z����{]J�����sb�B	f3�%k}尿�+�2@���0�B����h�<F�М �e��K�������v��M�r�kH}�@ߒ�ubA�[��	SN���{���� Q��g������-�p=b�u&9�	ʘ���.� s��!C.�׺��X���p�����i��r~���o����? M��TN��I��:�!�	�f��h�pY���X|&�}R���L8@1*]Z��7^whF]t�c���)ø'���f6�H�%D>鄸	8jN�'Te:�ǒ?��b��]��(ڄ�kn���Y首��f�ȋ��Va���?��PǼ�K3�z�����S%rDZ��,ۍ�!�*�'V�atvh��ye���?�Z�3��)�@�����]�w��c� 52�)�vo��d-飿��.97����p�jld
*��	[S_����[,���I t�O)�˥����(����F�n݄�����]��D忧"�l�P ��@�V�jc�d; �mk!�JY���/Q� 9�P���I�W�q�*�	$��)�Z���x�3��"�AiR(`J���o�j��(AUT���=�0�� p.��' XbuL%�j1�:������4���J��aZ�`�����Q�m����ɸ� ��N|"��p��l�$��//|�1(��``��v�t��G����z��Y~ӂ�L�e�2h3pZ�;�*DK�qhT�;�����N%+}��Q���|�
�:�@���6V:,)�	�նh�;` ��e�!�K�i�߼���Q�nq ��fa�ŸN$S���-��zoԈ/ ��!?t�K+�)� ؄uh[�	��٧V 13�	��Zs�g����ܲ����N��% c����<X�����^O�z�;C�0~ A>��Ck��x��c|�Ȥ�����@FAҽ �� �f%��%��̽ ��k�w�V~P��)�k?|9���"�fq%,�#
���[��Z��W�tu
�rd�L�r����t��X�v�뽵�����Q���E��X[Z�r�QOY��D(�(ZMpA���~�w�Z{~d��-�1@��3�E�c)��58Q/��X�M'�|zgY�1�>y�'�L�q-F�u>�I�> ƴ�@Ӊ��Fiy]�����a����XZR����&	uD���J7���}^��4
H(��K^^X�ޱ�1j!��q5W	��	�~�
>�S��β8R%	ux]�ˏF�p���C����ړ��N
ߢ{�-��~��:B���G��_�`�\\u'x�_P�r�Oj2�)�h�>�s�b#xУ�aR: J�xh8 =O�v�&	�L�9��)�dYn�� ���B���j�x����[���uN��\��U���� ��i�)Ӻ gP�Q����|�	�h�(QZ�?�
�,N�Z���>8JB�2k�<�!J������ɽ�q"���d�@� '���\g%J)�� �} ��^?��BL^w��h]^5���|�� ŚF�ad�Hlh�:�VG�%rɥ�.����2��`�]U��T����;����M�fQ�p0�`Y(�,t��S����*�P1�=���[	���� =�	Xh8%�˖�o�RD�����]}̢ש��R��s�����A�b,� �RS�Q&�ۃ0��[��0���}�i�Y� �9}���E[�DO��%Bg�J-�M]Oa�8�)��T�	���� ��-r��3I����+F��f�X1�:ƙ��J�p1K�E����ߌ�!X��;G�?�¢buUg<�:J�G�͢�gJ+ ��h�e���`{��MB�ut�
nd���Z�&@��<�N�9���1�����[D�0�����U�R���(�W�Y�������h�|4��{ �zZ\r���SR	�q���CWZK�`G5^<o�bx\�&O	���lxLN`�,]�S�	�.��E�{ ��k,�$U-�T�S��m�9Q`
8�^�3L1�>7��'N0U�5��~ ]��Qݕ*��q��f�%q����	�/�_1qyh�6~O� �8=I`��g4@*�QAj��uV�}��:�`��!��6_�����Qb^��.z���Y�5A�w�x�&[H(�b�-1����:�3��[h�V*�f��W�T2�bb��{v�� ��=h10�PN�*�\��5�����)�����8zB�
T])������DJ��r��iC��0��$x\�$pLK�e���7>�~���`OA��9�������aZ@*�̉�(1˖��Oq`����q=G�+\Մ.싰�I/1�l��)���`���Ɉ �Q�n��@��\tE%�*X~J^��Aֈ�ø������1�q�&*���'������k��*�UDW��hǾ� �te�ِ8N��ʮ��-�)_�Y�f��-�S���-D� gdK鞚�b52[�%2��	�|�,���R�7z���9ǀ9���y��Z�!-��{V����Ȇ�&.�|�,�Y�=�Z���I�
��sD��-N{���DX/�	�v�J� �M^�@�Ze-uqv�%F!?�@�yRA��,�Hr�@X�N	�z�gU�`v]Mhjx���I+)�X��M�� �$�Z}b-	#�Ĩ	(_h�WF�-t>h4'K%�tN��%et9�_��ձ��%b��ݤq�t$%7x�(À�}�]~��h�!�Uy��U�� _e�g_�,GR��Q�:@�� �����G×��m�^K1�D������Zx��|,�4l�_���u)=����r���w����N ��Ʉo���GK�-�å�Q��*\���`��WPA�>_(���T�`�B��Z�������e�J��lx���Vf*�uI�PP���7b/�C9�c�T 6g�5�Ґ ����A��)L��J�J8Zh�����"o{P��NZ	�5� ��oh� p���������5�����+������{U�{�7uthx�B���_��,��Q���n/�k!oT�Áp���z�q�;t�?��\[ ���I�[�I��Há[B����[Ԁ�1-Ab�&���=���>Ǔ���R��'_	�Հ����i�}V%[�Ӯ��h,X|�/�I���>N��٘=��{-�%�X?�k��i�J�qu�G��1ߎ+P����Cl�Lnc�!ʮm�#��Yv��
�G��i�j �3|&!���GAN)� �J0�[��h�~ܖ4��^�w�z(�~ϱ�P����0��*_<I�F>���r����ANLPn�)Z���ɀYm�]1��З\�I@�Z/s������.�{�4X��3z��HU��	��%�D_\|��<���� ����sg ��>�C�H�}Z�[�W%'ܥ�*:%:]kF���Y�K��LX�'���%Y�R��x�S:�k�^<>��ʃ�"Q��zx<�]xM��&!��T ���vN����`57G	����;=��~ǭ-p}Yϊ���5�Acqx	�j�����q[X3�y!����鐧A���6�8D �fRH,r-kG���S[���	���5G�vKY�c�Bp�qK��i���[s�Iq���O�4PP�	'ڶ&��D�_h. PX-�#�X�,��yKؑ0�.R�h.�3���<,�����/%�ɉ�ڐSc �J
M�V8��y[��N/$$�J�A�,}�%0E��)�.-�;��=�b��h}$�;Cݗկ���Z1^��] \i��6-,�;D h �"�VJ��@^�~N��q����|�1���J�����UK�����T.T�R
xl�	W�$%�q0��S�3&)ye�KU���B�˭�H���IO��)8��[T�!��J�&4����vKӿ%f� y�bX��AqO6�;P����-�Su�K]��ƥLP�H�6�s]��4)h�>�:pL)��E��t���ѹ�L�(�J!�O�l;};4lRhH ���G	)�_c!��e×�a�sj���	�煴���]�Ǒ��Ōd2ˠtR%Yh�zl��G
	�~k���UP��Zo��Rĸ�"-8(�[S똝B{-n/-�q�~�@[�h������\ր*`ʽ	��I��|��t��`Y���T�J��Z����y���d.���?�X���W�8�+�B![����n�j�[��/	`�vC@�2�C�� �Uhn!^[W����01j!1opʽN�����L�[�lt,k|�P�
�� }=j_"C���d�7v�?�ݐXN%��
�Aa�o�	��F��*� �|Q�^�X��� �	Po+ C̐�迏��bkѺ;�dr��a��lM�0��F�Ǹh#�M�� X[�� s�4mo�@uK?Xy�,� E��4t5 ��qM���/�ѕl�LX���ƒ��<~����xp~���y
e~J��@��@x�
ӵ@����_�&�B�_�p��<�\�|����n*��`Gh�7Q�H:e5�|�� ��TJ��3ktP�?/�"���61����	] �P��iCrC0Ђu�_}���j`\ڇ�����Ś1���X8	_�[�IgU�h�N)%�����!�_Gц�f{��ZC�s �Je�gA�1�p�����;��ub5w�d� �s�!����)�_h $��Ld'�.��bK2�0�'�ά?�Q��\wX�	M<]����(&�'+h[������_W�����A�����S1ꐌt�` f/�z)�!�ʓ��_Y�������I�|2(+ݤ�����_:/�P� �:3?B)N�����P&7>�h2�u[�^��0��QI fQ�� ˷Ԙ�M��P�%e�x�'� ?�Vk���c�
��c��&YhMy�="m�Ӵ�Mf!��_緧�g�$.���y��8 ����	
<�S�`��ME�8�{�~ʨ��}�]�P��n���W��r��A�������[9Z�<v��*!���ۋ`,�l���u
2�L�,.H�E�~�u�>�I�z&��] ^ݜ����Ap}��4\/�8�Rs��U�{D^������`*�k���{p�uaS ���n��,o1�2"�~BO8T�5�n7��:��-^R� ��l$���0��^�/��9	2��_�Fhe�^�)�z�˱X�	��������x1>Љ�w3�)f:3�]�	[��Y�	�6�XN �ŀ�E ʴ��]��\�|�H���ta3jz���#�}@t^1�3+��@��Y�����k*Ո��ogȑ�ݳ�_��9����g�2W8��{���U��xnXF��_X�L��%jYH �A���L<
 �/C�`�2~r��P(L��,��[
\:�3��0������P�m���K�Ax P̢p��;�؅�0��D���Z��E��	̴�Zz�Y _�h�t?n�_��x!Cfu�~��\C��T���y@br��^?4���V�f����l�HR��fh�Y�/o�oZ��i���,�00X�%��@��� b-�!	�� ���5�1�;��a�(È�*�f2ju�	Y!_��%���G�( !9U���k��	���>��.й�C�ܰp��{���L�RIs�~�{��v�>���_~�/ټgR�c�E�׬���������v�1�!��V�# /�U�� �%N��үC���W�ם��������C
�=E`�=J�P�#.C� �U��\�M��]"c/�&Fd>�`���n:%�0g�w5p���!��x@�����/�N2O ������U�LB��!�4
���ZB֥�Hy7�"֐@���`
��ա���zJ�G����p��#����o�[	������;�RX�-R���H!�+.��4�3���d�n��	`F���x�P���`�Ĺ*���]K:`��L�%yI�'~[���v�XS,���!���t��}��2o�B<����2��p�Ǿ,��(W �BC�<�qiu>�"}�oP%]�XZ2��\_10�dX�, 5�]f��Z�B{�+��;���6�a�Ҩ��i�o,�� �~j�3��G)W����'#��$2M����;��W �,��1�_��Jb�sA�,OD���uC ��MT�U, �j1�V��/%�~|���pFD���wQ��%/�{�?��~�PC`9�h�z���	�]���Ϋl_.@|� ��skhJ��]����5�?�(G�%]��uv��h���I�=��%/�T��oEi�$)O[>��������x�P���w{[�~nC���0up� �R�s�[ѽ���U�(�э��N�4�e<�o��u��[��^L���\&�Q���MZ~\5Yc�g|���ĺ�7�H�@Sh�K-f��"�S�X-�=�{Q��o��7�?w_͚BmE�����������v{ax�{�ߍ��/�@��i�5�P���'��<)
���ɐ�48��?�*�# �X�	�Ht�\�8���~{q~G�����_N2��<�u�W(�'}����'VǴ�'q�T:iuN& ����^�j��]�c�P�+s��A�>�|�FB]P�0G���X�p�@-�k��Y%V�;i�k'!�Fڀ��^�h�P�X.�|���;�i�U�;����H�SXT�%�B�S��DXs�N)9F�%��Ab_W4/�(?����0���D�+���JP�c;�~bx�kFh�In"��� �-(�a�~�G����A1�I��I��=fX(��єx���{%[�YX�ء���h�s���	�d����\8���+�"�pӑ�
Bܴ�����������'ߔy,��%`�Ff�LS% Q7�"�w��u��Ua�.�Z�h�-����ݡ%x�	�i�z �I�.�� �[T�|���8h_#h�;�=�>���l�T~8�����x��)����:���_�A�t�P��?e�>��`�u�.����r'��;�s��  �{��[:�˽�K��'
u�0".?�7�[������^���� �`u�w��w����&�}p�!���.�BZW��� G��
k�&���! �25Z;K�$H �?8/����+2)Ѹ�H#9%Za3.C4-��sh���-q�a����1}K�L��ZP�:��"8bF"��7^��0hqO�il'�)��&]�U�R�鎟�(~c��/Q�,�{��R�	Ƀ.��hV�~�TFn�Gjh��6�pt3�@7�Ss!$	��k
')������1�Q:�a͈�*������\�aU��8�@8�P֠�Yhn&��7�>���ӘA��Z �-�*�p)����2f|3�/���~��s]�� �h�T�?��(v��1�X���44�,ݺ�7Oa�q� ��Dg��p�'�����\H����7�_�>W��l�ļ�(�	h�x夼��	�"�@v,`�rxnO*�e
���
�A������x�|o��T��#A,b <�f=.�T -�/
�VO�5�6~��p�p7��@���vV�	��JL���E����V�4�7����)�w1�h����d	�L�yc��&�n)� F�5�#�g� �]��|'a��%9[�q"�/Dd|����1Aq6�*��O�i�c��0�Y�_E�1�[t4h�����ϧ�3�1�Z��9)�W��^|e˱� L_��I��sj�g�K���_�ڸ]�}�OF� U�rdq�1��*b</��σ+p���tI�J�%��%w�� ������.�O�r,�:���q,�~�^��@C�!��_^'@�G}��q{`h4u;w鱯Z]� �SZ������3�*��^>T��/��Bpz�W�Tz��1P��)F`T�* 8����> !��K�N�-~�����3H�7�{�g֒[H�qL�pzA0�S-,/9Y:��9����Zad=�.�ၻ��?视���	���3�[\VOd���1�c��qMz�0�|	{�%U��S
�]����F	����>p(�u����h �=,x{�����U`�R�H�i��5	π���|��LV��9t�A�\��&u_j�D �BG7�)��k[Xx�	�#&�L��YXP-�N����R/�
���g�J��)��o��e�t!�XZ�6�YR�Rp��gj%���)�j3�K�8����0}��a^;
��X�Ò칳�;��oP4��g�x�q�WV�$>�����~w�Ⱥ>������M�e ��W�ftx��� ��ܱD퉂b^�CH�I�R)�JX��9GAZ��J�:�A��8��A�R�eX�a%G�Б�[%?�����b�B�She�  ]Z�A7������}��!���������-� Ӄ���	g�pI(Z�S��^���K��� ��Xԃ��4P�0�x^oI�K�t��I����Į����4|E��;�h�kqk��v<D8� K}X�-M�	 ��czY�c)_1�Q2~�����+/(nYh7Q�]��S��F-T��rX�,�N�ɕ->��ao���83_�yK;�%��z����&R� ����~�:�-�.�C�d2�MQb��H��@���1D>�m��ﰡ�u�C��8�-	�  �3c�x]z� %�q�R-���Bî؟�qR/�/	��N)t��""��X��)!S�R��YP{�CX��3�K��2�BS`��h��^��Bq�'�B �"b�3�X��^0� �70��N��}JQ����avkL<��X�@X%?pZb���@�&,�,;ŧ�ު)D�-a��	�0Z�y�<�oCzO�)|*�t&�-�h��8&`�+i8q���F�f�����_4[��
��g�A��e�d����Қ���kO\h	�trfTzZ�`���ku$	 �P2;��W#�]{�]b����fh
������xA�15 �f-`td�G�
B��&�%zf0����R$/\~'��hFE�eߐN��;/J �sV1����LO''l�C��ك�n�5 �t'���͑�%&n���r@�Ц�R3^�[&�Ʈ�Z��6��L�Do���G�W�J��`c�Q.9ï@C�ml�D��
hr  YgZQ��asA)�,�Rz���gԉ�w:���q'��0iCK���GoZC���b�`23������I&�\���^Q��\��;dF�++�*�7�PQ�=('*	ݨ!����y���X6>?%�fhz[] �1+3p�Ͷ�=��q�	����	�-Y%�a��_�%���KA{��'5�!J� �4uc=������2H���Wd��*Msb�]�n�^	hy\�� l��H�+�΍@1p-͔�'u�B���V�Q.�q�vH�j1$�^� ������a�*�;�\2�K���i�J�f��n��~��z�r+�$ 
�r�����;~8���Ggs�C��`4�*�|�TKӽD9���'|luwqrH-Lu`�"�*¡�q �l�q�_9�+�nj�%��Y-h@�	�X�M !��1%�<¾-�$��D麸���N#,��D��@�0�[ ^��.Yv�$�%2�	����@X��4x����~�0ݯ\ZZ讲0w|(H�bL�ur�_Y�-�\�Z����	�/�t$����t��~���`�5�/1�T�ͨ�>�#������^�DPZ���3�3y���i�x�(��vV0%�`ZhiO{��r���@l&xf*�X0jU�j����ߛv��!	�)� Nh�C���ݛ�&�3� �*�?� �P��������1S��3.z
D�>���o lű�)W��3�>��=�N$'�Ņ(*�'�.���u��y,Y�L&�a��>!�x$�\�^hA~=?�@�QTY���$�D���J,^�@�&�0�,xN��'\�hk(���x5\0�L� ��IB��ڇ�fS�4������R{��2����N%\�:-�ޫ����F��Y��U�B��W��W��#��;�O��E�Ho�eJ�D��>O��@�������G&�H1
|9�7Hd�,M��v8���sW=�뱍O��!o��X�Ym!��'�ښ0o�`�x|�"��y./���#�o����X�m�����2�!�s0�XҵՀ�gůa�(hu'�*�_/��BX<OY �Ȑ���EXu,�fNkGѻ�?�]��h_V��� �6��U��`�%)x^ـ�1=�!˝ձA?�꾨��3ȗ�AX'������	g�;��0�z�i��|��0>`��0:����	��ˀ��cw ��4e��$��(��8���)� ��4��;U�wi�T�i�Dims@��X 	8,��K@�_���JF,h*�*'����m�~�ڌN���n�Z��*�		,�aV�+��M�����ƀ��(w h�EQ8�0�a�j	j�}�Ӏ�1�')���+[ ZU�6{�D%��l�4�
�t/np���Qn�b�1��S�� P#�7{,��K!�!��$��\B`U,;L?;ˋt���u��Lf�J�}^l` >�V��S	��xO���� ��O�%[�U���BTR 8�_��ޗ1`Ƽz� -κPY%y�Zp�.�[T�#_b��p-��a�_���i{P�	�^�DP��]�hb(�Ӡ�0�r�&{eQ��a>�6}�j;�4��,a7!�F,�V��x�W�G�M���<Y~��age�O�*"�3P$�>F�{�a	��pq�5�'Mb�N?%R��O�z��%qU���h}�E]�a	1�ŎBV����>�h�͸x���\��� f�ꨀ-�(Ԁ�u��:����8�% $4���V�W�@ )�_$�P�`Xm%�	� ��'��_��V��5���7���^{ C��e�
��B_�"VOH�� �?h�]�_�A�E��}��n�� !'y�Uƛ`t���;���L�k4]$Z��!8�)�!#z���k W@-��)j��I���Rn�%��VPޣ^)�h��U��A�8|~��í .�2
Zv�,�ChrK5��&;�L����Xe�	f�y��n ] W�F��k�Bw�J�:�*�Z����Z��j��)����𱏕�&��Z�G��-�
��H�14 ��9P�+�*��zʰZ�YN��o�f6G�I�.�E��ɻ�pJk�h�q�m)��Xu�v�	���N�k���^�U�̷cX�7��n�B�o��"/� �` Y��d%�^W�.�hiU��%_�;%w������vW����R=Kȕ� oBlQ��5'���H�.�i2��@�@�}3\T7J���4p���K��̠#-�	d
�s�r_N�J��d)1�nVT�C���I���~�D;�h@9(P�8�09>�5�z6�T�;��CE�M�2Z`���b��q!�k(�P���������/�.�K+p�T�}�Bxq�m`!>-�Py�	ÄW	��[�0�j.�8�OC�M��zY�2�)�~�hĿ�@�A,GfD �9(�t����+���9v��kLP��C%����<I�b\�M �t�FBA/�X�B	�w��{�;���)إ�4M�^���0����P��Z����9B� �E
�~���)��wY�Ҧ�/N����:�?�Rl�
Da�&��O������8�6\ ���c���͵�p������	����ǭ�-�,�ҹ��Gt���b�H�-I_0jA8	�����¢�� ��2�|�t� �0�X �?[��t�vw�"@օl~�n�L��f���K�Jʧ%i�l+�$��J�����y?�@K_���"����W� ���|t=0A�7P��!�[���`rhL�=Ԗ�A.�8�Q�~qi�=J�.�Y#��	���Vbs�M+���什@_Z�H3�H=
��!��sQ.�~���&W��pZ�pO��U�d|���}{�>�h���`c��AOz�ٛe��;ހR��hl��0�� ����&{��LB%�y�F`RXHS~��y./�)1o��J���`D��-^��j_H�B�>\hKJ��N툦u'�n��`p>1W �PD�\Qh-t�y|��0<���R�1���+����({�����
l������a��B��rpNl��PLh�dAQ*�����X�q���( �K�N*����5��Z0G�rH��%�T�-�1%U5��w�Yߗտ�0�������;���Y�8R+���]���.陰@���}�?c+��W��W��H�~i]})�}T���o';�.�(���$Y��������g	a�K�������H��1���T��VB�<x��I�����b�K�u�����R�-A&)�Z{�p��"��k�q�$!T�w��d�O� ��u^E��a���'p+��N���<z4 u��n�HJ��B��d�}`�(�P?��O����vyi�}�9XO��@ø�?�]�sJ�������wN�BЉ���t���o�����@h,���ߑ!��/��9[�1w��6}Q�R�{4j	]|-	�� �[��#�)�!�a�n��.�_��7Y��@&�K��&v��sO��bCK
ȏB���V�0Yl��������!��bRh捝~r�`�x���*��=_���,A� �A�q)ښ������>������D�?�O�|���l ����N
%Y���'&Z� xQv_)т�wR},�ƈQ+�>�L0D��>U�Fg]��z��1��Ϭ�Te]ëo��Ӣ��^)V�(-"9����.0
��M�%J���ZG	�Z�	4��[b��ʹ���Vk�U�V�9�����_jh5wn�	���?�p?�x���wz�>�p��!!�*�5��hFn ܮ ^�����`5�ܡ���>��4������\OK�b�CE���T?�:ev3&�5)��3�V���� /��s���u$���bP��X��;���S��ׂl��'[����'�ZI�
�yJ b�ޓ����s{���1�yG�:\j7�g�uT%:��şQ/�����z�b\��s���P�~���>���0�[�n18��X��Lq(��_��"���N2W��F����/"��3���q�A(�I#�N��x%?�ʐ�0sN'����}[|�V������F�r ���.�v�-Y~�w��P��Rh/�-gD�3��XPh���Sbl`f��N��h�^'7#%i��.NxC�v��L�H̤%͊��<M@`��^sD�)o8!7l��\S�@)���@��Y���n!�E��i����ш�fhC�$L�	0�/V�z��\@
L7 ���(�,�/��S|�S�x��:
-.Q�1�i��ԅ(���UT7o��h�K'���Rl�(��v
�F*�O(Z�q;q`�u�n�{
�{r��@h�� �7���d�e���A�1�|-s� )��P��| �"���}( �n�dGO`��i�$)�H�c�Ոj�����c;p��,^��q�#q 00�Y����' �_���h)=iń�V��!�t#�ڞ�`�Ō��pc#��*��l�aaV�_��/�0��}�B�E`9��+���af�+�0�F�9���B�m�y%�[L�1O���_@<�S.P[|B���% �Zh�E�O4>���#')���A�f`�@Q�*�h�v��AP��e�0�C3	�)�ꍄ;�)y�^!�v��fR������aSC�Z��
�}��S���XHB:����-�B֧^0�4K9H	�[@��|�����o�{H?B=Zz����Bsꇆ|�(H� ����b;�O)w�<-yVI����~f8WC6a�	��h P�p�k�[	�$�W�-�K���'�	�5�jNP����U������)��J !Z�G$-N 9a�v
S�#[�L��$� �����H��LXe-{7>�y^��*�5f&�
<<�t��+%����� �TJ�*!�-�|NNض��'�	P��͟��>�t|/1vW����)k�J
鯩�	�҅��	x ^����(�Z��Q[�D���5*bHf/���c7O�i���W�5E�hO3��!'���X[����D�����)x���1� 3[X�M�w��@K"�FV�xI�r����u ���xqP������
�ո4�	�٪o�Ǘx&=g )�b�G���wݱ����� -��C�!���\�~/�\)U���1�h�WV�cC�/_"��պ?`ՖҪ��	htJ"�O��}	�f�PA�G�2�DO,��!='�?/Wh%?�(�j%�O�2!mL��9�Ъ]��8�N�˱�sx�h ��PQkid��E����!'^Q_	�s4��b���;U��B+�=�b&1��!� �����Q�`Hg�1�$�E��-�?�y���z��XTYK�V	m\p���z-,[8C�Gt��(w�E�
��O�~���]P����,L��
��U&�ϴ���F@��7	���;�(K���]n<�'��90�1����m�V`ςgE\AU�V	�]�Q�K�W=+9��nV+Ph%�J�]�˧H
;%�i}�}H��^��Bf�5���z5v]��[	0�)�#�R(�e�/��Y-� �[�1��`�#�p��&>�^N	� �o �,D6�P�$|�tTfi�N��9��8('w�����Z�f�);[�zSq8z���D�L��J� K�p5YPNh�f�1#\�01�	E&y<W	�y�f�#[�	��a%�X��`SfR�N�ЀZ��0��߀�}ڍ@���0VFZX�y�/��N�(�Tg"/V�̅�8�K@#/'�9��� +l�y�ԓ�L��;�d����`�jQ�X��A֋�Q P�:��zP�Z<c8e��T�p��	]�_T'H�p�Z��a�����ل鳆DDf�`kЋ�5��B�f`�~%�L�'I�ׯ`�2�R���7 ���*`%�M�^!�A��|
.� o�s	�k�W9>%�Ԗ%�/�=3��jN���j�v0#�c W��w$����Y
��5�uK����h��Y�`)
x����6�d���7?C�:�|��x�ڽ��q�����
V��%6�O�����w�Z��$˿��=�z�贉�Ҍ)_s��#�\�>Ĺ
#?w�Y	MvV���J;U"�1�]�FY6���1� H5�� ��B[C��Zh}K!���/���["�XZ�z�$|��+�
	�{�9s'u��J�4�1�C�VPh^.)��� ,��*�3��U?Q0�ԶT����M��]a?2j�D_�/�	�d���2���O�s��:+}��'BA{��1�U����$!~�9r��ҽ1�-�-�JO��`jYA��b�=�9Ab�:�D��!_��}Pi�>ӸAR��~EK�@��[f��W

_z� ���1ʐB�yL��Xb�`v0��o�f,��eL+�s].L-���[O0'�����0�quJ����0ǩ����h\�nSg���>�g�o��G����A��w�6�%!�ЉKvn�W�|j�T	nRvJ��H��c���T�&?J%��xԀ-!i�J/��4Jv�}/�����?�iӽ58̰�G��(�q�h�C�
Z��'�V�Z@�k`3}[nx	��Q-arbp�F��0<�m��4@p3�1Үʽy��}6\��5��DJ���g`(-�/�wU,]Nd�"�Ż}�l��
	����ӿV����鶕؋����O����鑩&$�U��/J��E?��*��*���g��;pt�q�v��dח'��d_��8��� 9s-�K��{M2`�~��W^���7�j��-1�^:~��!��b,�8���\!]�j;2h����c�HH�{��U^S�:7�K��"��`O��`)�{`a����G�����J�)}` �_Z̤��",���U�Oi 3c@kX���m';_�.�Y(v��;�<�hՈ�(x��$|�XQwJ���~�BN���y����䓢�þ#�^�>��������d{��Q���^�)N���Xh�7�/���=ѮƚAѪ�e(E�[Z�02ݪ%+ ��ͷC��w��j�K���1��^�O�=� �k�n�2h�Y�J���L��vr��!�U*�E�Ĳ�Ʈ�	O)lz�S�7�����_�)-�f �iy��50v�Á^X��/�.�g��[ �M�i���)�����D
!�VR�M�Z$�h'.�� ���J�����-� �y9j6-	P%4FpY�K|w�Y�,0�I�����
V3��Tg�%P�i�`�̊(�����CK��a�y:Q��̹F+�뱒���������%6c�}�%��t\�$Ah~L�� �u?K�,5%o!���P�1�!�2L��-|�y\k��N`��8�\�O髹N��G:�m+!e; K\i_b �Uh�Q�]��Q�Dt�& ��>�\�ڊ��׆8�-�Un�1�F��	/Utz��e8X��0\]� $GB>�r��}\Z#�ZF�W��1��	��4���Khj'�aK�qY�{A";�|`r׏T? ��.�	�=1�~pJ����pa��o.�w.zi	V��(�p��ߠ��C��� �I�K��Ò��r���Z[���QL�?�0ꋈ�
����v����f�o���B�>��*�4MafCK[�֞����S�W%)���}�;!z���&S����§��a(lF�>:E+ߍ�(���Ԇ��Հ\��3���Ō����_�Z(o �@��I��8�!B�ou���_�
@��w�HC�׳��b ���L�"�\V�
��w��
���$X���߻�T(�b�	�[����)�&،	C����D�1Gb�!n��)�;�ԑbRii���AYpŕGSz�7/�bU^w�n�w��[S�y`���r0u�>�u��6�����>Wb^�ιFk�W�h�$������t��0��,���t�O�~��>�	 UV��{�Z�@�qw��N4m�Z��� ���B�qC/_M���h_ƸA���Y6�tt���b��/�1���%&��,hy��sT34W��L��ؼ�/�����U�س"Z��"cg;�Y����˞���$����C�Z=:�G;l �=`�m��5zf��2 ��}jQ���hXF��)�K�ZM	>}�{w�,$'7�Ya1�)�p3�|.h~�t���VVA��;Z H����N:�s�q�C3���1ѿ�NX�i��Q�4�`:n+���f� $Hc~������0�Ɵ��&�#C��I ^`r�EcP'�Җ���<�^����}�;��yA` �"`�Gg�6�c`���$�eET�x�pP��>��Q���]_0%L׽Eo[g*��<�%�DT�pPW2��eB�Too|,�'�A
���h��`��Y@L/+H�P�h%��㈹�_p������+��h7K0۲���B��9��	��Q��Pz��鱼\j���o�H������̟��d�	 ���:�Q����00#��(���B�a�>;��pC��L�XM��Gb�Z�y�(X�u��@�Ik$�	BJ ˮ�;�	�1
޷~����>�v���2ӓ[-fKi�Wp�pȕز�=-���ɂ�,`R��_Ά^���.h�-�J(�ϟ`Ƽ}�����w�s�d,�*�����
� �Z����00�Y��Y)/��A�WX*b��X+`N�z�t/3��x@��	"Vaִb9׋j~`�qFr�Ek5���� P��^Uv��)�₮!W�XP#:b��1O�A�H?�t���ou?��R�N���\W.P)�a �:�Y�Ҁ�!�]h^9���߯�I���52Ҵ@Z�s,�1��q�J�qc!�/�W{09�H �f/[��,�#}Y;x�3����I�)t�5��Y~�#ֲ<ށ )�n��[��H���W�R��;S��n����;S���^�']��%~+ ��
�!�J[�j�`͸�vJ�/	��.�M/���{:� �`c�����5f��4x��!��V,���	U��%Zv�<���c�J�{d
���Vb�ĺ,a�ap/PL�;L�O�I��T#	�`q�`(�+�	�1�I`tp$@��镏������t���j9P0V-X�)���Z�*�mj:�>���K�<m�8�N��X!at��!��w������fW[�G��-
 -�M�~	�K�n%/����:��J�FYX�����aQg�d_P/hq��1/\�V�����K��]B'Q��@H�"��t[O��k;B�u��p��w�N_a��w'�h�F#�e� �WA	�}���&�fY �a�;�HЯ���3o����h���[6�����Q���*��f�HZ?�A|b�O����TBJF��xY�@��+��D?&J�{�mRL7�(�G��22��z>��N�G ���Z�ŀ`)2����Bh�E�O8�&.(��G��>A���S��]R���\�%�k&	a�@��
Z�TC�g��H\]X�
@	��J�� A_��4!o��^1]ws(��/��J"a[+�����)�p=v+��k�M�	:*	j��R
����T�"��� �B�N��h�#;
#KR�>�h\��)[T��H,�0�� K�	�ߨ� �.�2��� NX���E���hfT�+�i�+� ĺ����`��j�u��1*$�V=����,�CңY��&����X_��%�h�1;�)Hw�0�aM�\��Z��zU�m:i��IqgN��he�f	�~q��;�j�y���;�,���/�w�@��O�XZC��0�F1W�� +�)�S�bI��m�y�K]�5�}p璈J�� �� U%2AO\��(�;�`c�e	�[.1q�z �)�T����I�Na�b4^�`-�E��9�ZHTz�A�@QP0Yh_Z�3��t��|��PS�09� R��΀����/�y�W1R�/���C�m �o�?��P.�3�(�!x�. �O����v�o8�@%x<A� �l(��YQ����1�~J��J!B	�D}�u���f�$���<�W�	P�BK���ThS,���t.Bz|M0� ׽^��u)�XK��F7-�	�f��&nB��;�X�N�W^�Ǿ6��hI6	H8���)��҆� -�#�l�- Zg��p�'`�#h����	!HA��,����*�����Z�d����_��ȹ�҅R���J9�LhrטΜD&�[x�I��`�\)mL������8�C6�>���?f@�/�����-��U�Ju+�ӧ:.�^V�5��4���	&r]@��`���5��C�\<9)������-�qr��U&Z�
h0�z� ?_�Y������l�3$)�B��ٚ�â1������}�Ua���E��꥾�l��AI�+����)ȝt�R@�\(�L��|?� 5D���£W$�ۈ��Yr��op&J��p��1��_���!|��;��hUz�fT0x.SV�	Ry3x8�+��ga�����U�PZ�� p�v�)��� �͈A��%�v��ʝ*P �1�T�z������I�k�(	 n �!,J�SjU&|0B"�\��@��­���u,�ZOWxph�<�u� ��e��]$�|��=)2a��`F��~��:m���N6��Ӱ���G%;VΦ��8N�C��^�ڲ���S���1XZ[�P`�w_�L�A�%��[}����V�
��F��	�6ؒ����_��=�X!�H+A�(:-aх+l:�`̽&h|[P�P�h%������E`�����(�;�d����	_�	�U�?�f C�6��҅��3'w���$ꜗ؎�3
��� R��X�rQ�:�9�/!:�P��2Z��@5l-+pu=F��$4DW0ZE	�ܶ��:�����h�@]�^����X�N0���?3�Q���'U�(������z��������W��d����G� ��Y>������}�E�ʹ�R �����״��ۿ���& ُ���\C��T\� ��G�1�Y�J��,��m�v?��L:����!�U_��~B=�u|����RU�bk߶��G���������( ZVhxR�jS�	XTSp���]Ʊ�^/YWv)X�Li�.�u�V�觼+�x0bjLBd`��v[C�������9���A��|��R�0,]�g�X~	%aP�E �[�7;�\B��ɠh*a�$d�e%�W������^�,�r�M�ނJ�ru,�R	���@6���q�����0��(��	W��h.>��K�{h5`QE��������)�ʲCV�!���B%����0:�'�t�%�b�*�N+�y����D7J��S���axc'�yF���!�~pc���{����J�l0U��]Ԛ�I"Z~�hIu� l�'_d����`��?l�\�^�@"�p�E2�[b1����,�5^�6����*�3�U�%(�uo����_�w_� a�'J�2�]VP�)����&�5(,cM���8���F���qZu�n��K�;��Z�Q��� J<�KE��ַ����� �P��9���NO&H>��)_���-b�T�'|�`Z�O���5
9��1�g�Q*��BԷH��il>A�KJ�#+�4R����U��\��1"+���:y h�Z>]�p����К9�^�~)��e_p	�~�ک��6��qb�}	��Wq5��>�`󱝈�0g ��RG���qp�s�$��]�N�z`[�\� ��8�e �E �� Rh�&_)�ǧO����4�Z�a�Ձ���3�� _]�!��L
�U]��W.��"L�Z�1�]R���3Y������׳\�)뺙�+#?����J0f�j�%N1����_�-ur����Lƀ��`"�-VCz��qn���U�3+�!��D���V��4��[�q�⒋J��~IH�HX�w�,�!R<��HU� �50s��:�@��g"�O�F� ���ܮĿ�xD �?h ^3[V��t)x5Kk�	��f�7&1�g�ٟ@`��0�5�\he��J'}�t�wB�u\�P�!I .��Za� �S�����^�A��?�|��y��)Ⱦ�AeP����T',gc�>��%щ�(){z���&��|�N��n�F	K�����>���cI7)���%Y��^��&_Ӿ2?�G^h(i�`��ɗٱ�?/qz,]������c�W����UG�E1�3d)�0��Gz����L$ +}X�,[�L���hP�����[�0'��Z� Sh�T]���Vk�~� ��&l�=W���#PpIo ��Te1˿	���A��(g���$Z�^�lR�0!7���~v�W�_��l���1�}�Є h^b�PY��5���4�?:`WI[��J����a[a)k�w)�0<ԕ����x�,	L0I��7� �q�r�-�v�
���FO�O�Zop�g��N��H���x[�N)�:	_��'���+W�,�Y��T~�i����� <uL/qZ�(
����+�0��2^@	K�)0��K	�gE�M����&�ʚ'/Ȕ7`�X�y%O-���9՟�0�
��{� 	����xk�&̰�Xh���a��D�B� Jg��Z�ܴ�1�����Z�,��!�g�ϐ�͡.$�Qh[�Mw�>� �(L�c>	*@-�ݿH5=7� �	mYQ��S��
.0�*~p>)H��\w����9��BK��&\-3�`U�J�_:�K�7S�5D��7h��'O�C��4K
 ��? 5X-�8EA��H�� j�F��URLy} s���n��%
	u�s����� SU?y)O,ٍ[x�[��Z�Ag�/��N���h�q U��s�0ZY�H,����>��B��j���ZI��5��!��a{1����"Z
���!�`S�kLV���l�XQ�%���h3B^�[|4��ܐ��V�{�d��_-sE��C��~wX��[�u���z?ég/�|����e��c�~LZE!�|����C��R�d�QciV9�
���/H�|M���O�(݂C*]�v�[�1�h�����)ؿ,e�9x��.( aKW��e-1s�!�htf��{�-@�K��A:��ZXW�'����A�x�-}@X�� �(޽� /qxEhF�0' �Y@5+�Ɖ��]�C=��p��)���IP�	'[�"R/f	���ZLڣ��3Z[�0��<U�h��Y�C��	}���%T�Ȱe��6ix%wgq����(�+I�WJ>��\A�E/�Du�C�¯�4U�M��}��sרV2Sv@�p 阀�<�v���BC5�b�j[�CsOZ��ը!n��|	�DAx���-y���BѴ �ܖ�wHH�[�*����y w�)��B��h�A\%g5UdjK���+�}�>�Ĥ�ڣO�r�R|<�A�L1�.�=`�X&�m6� ��}�1IA �9&���<�B�B��A9e�nn����w����=,�/>��hv�%W��s�D�-;�-!�^�W��_�(�����3�[���(�$����Z�\m	�g�~���ط@�f��ԃ�;���	!طk��5�{��.;��kp.�l?��$� ��J-]<�MA�Ex�,C�
�.�-��	0� .����� �^Ӽ�\��N��B��B����v�L�5�]�= #gm���/\ ��<�D]q 
�Di�����Kſ�Ih%;qW�!0:�[�L0�I�y`�WX�]�Zǀ�^$�#;P&@U�^�R�~J��5l��o�r�Q�{�P�P����4˩H��&�o���M ��gN���LJuc��W~���pt|)
���b�J��w������	]@��iu�_>1H�R?���TLc�8�a�UT`����W�-h!�	VBX�H�@'U|4�����9���P��H�)1�L�7@=x*%B]@�u��^۸6^�E����`�9 U��>�1�i_��r� i<�\I�9?�|�]&F��ᔹ[� �Z��~�a�\H�
-d\�@U��*��_��@�@,�W�I�vZ=4�:��h�����_yLF2Wh�0'}���
T�2�ZY�1��N{˶����0�9s�y������ǆ�f�?��J������܇T�^,U?���ʱur,�HBzZhr�c�	�\1��+`^�\�p�sm�U�栖��%�S��O	�W	����W���->V\G1�^f	�`�~#�&�%.X)΁��I'j�jL��l`��h�[w�A�o{:?,=�Ak���hyw\Y�r��4ɧ���sYV�ށ����P�%O�Ud�{�%�)|���]C`2���+-��éx������)��ĸ�9x� �d�>���� -(���pk�\�Z��� &V��0�%^�o�_S �[�.5�!)-g@����_�G��~�י0~�'��BUō�w�S�S��
�_hMJ~1V���������ؐ��Ct�g�w �EI�H���-�h�)!�Y}�	a/�V�*7OW���������L5%;w���[�O�������h;͙�%�$u�1���X9�G��rs����5In�yD=HT�;h��K��J��f�=*Z%���,'~Q��(D�����H�W5�,Z?��^��,�$�1���/�Q�ǥ6�w��YC!��D� %/c�hџ���G P� _�8W�ۦG�TD���S�H)�����fY/����1��Q�Z`�R��.�k��u)�ud"�6O1쭅=���r�4ݘQ��đ��_��\5½�R3*�r��P�żz@v���9� l�8�UhD�� �
)�����,�	z;�BA8bQH���&(��+W7�������@Y1�9jfZwiK��?7��&�%�Grd��®���^�ɰ��f'4K|�8�����0��C�b���0�>q�.�������Z�:4!�5�1��[*�B��U�#�<
 c�7|�?�z ��%DBPp�_����h�p_�?� YRS���ڼN�=%�ӗ�Q3�Ź�7�"�%xa�� �����ދ �Љ�KٸN�"����Dh%�Z���&��)���}�z�N�-8�+��&O��O	��ax�0���T�r����:��?�����kj���g{�-�*��A[h�~�CY�OW�Y����<��l��:S�	�y�X���+<����;8Q��#��(�K�?oϐ��R�X+%]�lh��O��D�eB�}b�v��ath�7�'ߜ�u�7��b����&�PZ�CO��	E�u+o`h�$�Z�x��S`Yz��	��ȟZ�+[�d����m�騸��ړ��V `�O�D�b��	H�;� W�L_!����hN���:�@�Jw'�B���%�]�1�~%�X�:$��	[�_X>�������B'rU.�_#�=�ӦX�:��B���\� ���s�;�X��Y(5y�	-��.����\eH+7֕��R��Zk^�����0$�5f�v�j(�	pn}c�P�/3 S��.!h|��
[Ҧ�x�1��LJ���"��G�b���4Z��{����aB_+�|�����z�c�7̰�T[���.��_�V���al���
@;!�=���y_�w�7b��-RQ�����
��[���J>`T�cI�B<����G�RVpR��90���<׸�>�L� �Ea2U���]3����:��	��{	��RC�	K^[WRI!E���ŀ#�a��HU.���Q-�
�(��"��X9Fu��.��v�!�j4Ur���@{y�����\I	!�-M�}Kn�* �(�u �q���!Ϳ������E~�����o 'X�֒t�d�%��MU��l�!a`�ߗa��_.An	'�@%c?������-�uE��ݽ*�yG�'B�3!Rh%�Wr�Q���i(�A�}<��L��	h0{��q�+��a�2k�f�#U���J칲��2�����:�6�1�[	����L�!��!a�4q��Bٌ�l�$}--��2��b
�߸�QV���޹�*�Pp�O���[u�ciծ���0{B�����]��J���1�U�+~�i�I�� ƏE�dS�0�O�kӡߋ��ZY� ?��"%.�/CtLO*��J���!�[�����*�}���hJ�z�<t}���|�Q�X2$��Ou��l<[7�� �] ��qg�`B��s)�R�	�9{w��N�@��Er<�I"��)�z!�5?Rs~�[A���"��p�'L 7(,6+Z��O'��r��]�o��/�{���|�p}�#���EJG�������!���n�[�^8�����j��ɨ``�|�)�K;��f�>�*�����1�c	!��V�<w�[_�r��y��w���U��y%{ N@�"U��,(��^�$�
�4�뱽�7YAf6�� �h�4���S�������R_�F��/HP��[D<�+�ou����}9�~}��,���YÏ��Z�{:쳂�b]�P����[Y�C�Ö��-�������"-��$���R#?Z���!�.f��@	�R ��?��y����8��*u��e�A�o�hd+�I��k	�Fcr_H�(ǀC6�y��|����{���(�M���0�^Y�G/)#FId��C�ڦ�^�g����_�%����S�y��kNU�9�bpl��%5Q6���p@�E�'��H?�@=�o�,8��e����f�:"��з��א�j(<O �lb�ڀ_Ͽ71�|�ӕ8P)�]���ph�T�yG,�K2�	�}��?����@�o�~�V5�G=�G��\��5Cփiqa@��I��1͹9�7����܏`�y'�>>@���$�`Ɖ�^���%?��yhI�-����-p*�Z76�wF>ZS�����������Q�!���z$/3�q}m]�%_�G�-pI��%j�,��Yj�������Z�*�:�:U��(	#�|4���@�+zK0vU��ag�1[��*�����]��@E�s����8@����:�ee�u��*iP��]�;��1����:�vÐ4�ۀ�����9c���U�/K�$���8���'!�i[�xuP�pK
3�܁�_`������˕��!h�<q���N��%ۍ�\�ڄK��^�铆����Y'�F��Y�ѵX��L�9���A�ڀ>��ѐ����
�(R8��d����X�^�~�9���Fyi�4�2p�|�A��>�.:�{��3�� ~ 4��;(Z)��P]�z�@����1@�T*wQ�Ne"�$_�im{��6�r[��/�@��sG7�'[�}�N���PCo�W]���|�?�i��'��Y�����71���|^����]&C��v�-�����W��\�l�`pA��<ؽDO1����J$n�`$f�%T/�_z��O^�@1�XZ=�Y�{m�~�j�9�-�J�L�G��������CUhC�f:6���g�C�ﱧtj�}Y�3��)@��!� S�x�s�a'2h?h��>�	/��EA yX;�����,>|9@�7qP0��?2%	��.ߞ����tf�Zv��@��R�}b�^.��w����$�$��*S��Uz��W������������v��w���3�qO1s*	�'�|.)N���U{� �4�r�~K�V��_��%�c��H� ^���3�jQ�	���#<`{��YI�!}��]�NA�+��a�;�B#�w6�/<ԟe����B��W��hz3{�G�����1EX`^	I,9 ��4�^�� S��"��c����˖�	��s�tXBZ��M��A���l��9$)��14?(�pJ��(�$T�]:�Q�ϣ��E1z�=J�md<jY���\L��czSs��Q���-dT�R@��0� q��1�!�I ���ap��=�Â�%0������_���̓�T03�����Z��,�7���x(-��+N��/��KW�o-@r*�}��D���X�,�nP浝שoݫb��}���e8+!��
��,�0={����`��}��%�Y�bE�B��sE��e�"I��b�3��P��'�D勪Z��	����Չ.���]�����?�@F�Oo�*#ޯ,�4@ (�r
L��3|"��tM���97�m�W��y{U�r�Y �^� o�~�@01��RV�iqI6Ve,�����n��!d��vo����銯��(�N��S*� *[骳�m�Ղ��V��Hq\�4���5�a`U�-"�~,��J�.~ы�_��u�dO,��N@RQh��x�C�K��;�3�Ba��ߋ�h*��K�v)W��[	U�t�������'6[��!��m&')С�+A:�ӹ&,�#�.�re- 3j�@H54q�: +O?�U�Vp��{�O��Ĺ��*E�s�����9+�����wb�}SDd3�k8:�R��%#~�E�랕��O���y�-�[=��<bU	��f�܈]���	ζL��ԿL��[Ch����	s�Z�]���W����V��ɠ]��_�[���h`~<�֗�T���i�Gd(E2K��@���"�`�M7�h���W\�G0�_'fr�K�0)r�t�}�?W�uܿI��P�b��`�?�O���-���H�xҀN��&M$-��iBu�tf Wv_7Uߪ���K�`�Q�:0hJY�e�5A�[�o$O�9L���?N@��bh��U����9�����g]`�.4Q�,�S�x^-W�"V���c��9sO���4648K����BO��+�J~� ��;�����J��]��'	I��Q��J���@���涇�)�1��0@�A�n3oC�a\j������Z�5��W�~τh�_��P,AJ*��
�=
L�Gy��`�)ˇ&�[F��?�'!��`�[,�{hKv��ZI�����q���OF�'UI�޻b�M][�aD�.�� �s	��(�7�?'~D�,B��ݝ{���Y�:.s3�6E�h�ʁ�F�+ ��(D��w�k7�E��(!���w��I>
'��49h�5�NP��o^ �p��}�Q��h�d� ����Zs�	הp(Z�(l��)j�\J��� ���L�T�@%0�X:�f���7�o<&겈�wS5
�7u�U����J��Z� �S�:��9��k	�e-����H�X�$�)�����:þ����D{|��n|u]��f+�.D����c���@�&UA�|`�����vRŖJ7���TEX1C���Kt*%Y×pp����ԆP�z/p_Vށ��h�5p(>b��^�`[��ӻ�9Q;C��+�)�WA^W	��]k!���B)G@~/.���Ӫ�r}��J	��	����9KD����^LS�J����ނ@2v� ����JZ:��	X��R`�l�*�?�ԥ��v��]S�;�ƒ���z��~	C8U���k�ݗՠv[��`z����@)�-�s�[h��/V�|�zKC/��yp�K�����d��$,eN>�/3�
�Zoz@G�@�JZ\dOK�0[��vM�y��U���2�y��CS�B6A�/8��޾�g(����ʟ�]�Ziu�pLP�	��p�iAt7�� ��G�vh�*�}2�`ق����xH$��3'_¢L�c�a�?n+�|���Yh������3<W��� ��o�+�z<Z�n���ڸ�~�ޏkQ���=��J{Q�	�ȵ�_O��h(.q6��x����d�Dc�_� PPz4��@%pބ� %ĳ����Q�Aغ�p�$ 4n(ΗU"�;]SnR�C�h�K	�{���Y�!�E�����-|Ү"�t`�jҽ�F<���x>5vX���N>b�_�,ɋ\�8M�7�H9%0,)�}�a��%��M_&aKAZ����d�^�Q���>#�E�g'a��Rk2�T�;[)^��| KiJL 5��N�2G-z��S�|�\_`[G�%5'�U�)��oV�6�Ba�S�������k�x�6��4�m�?k���k�J�����̭�#G�����U��0ʜ8 �$#E�1�)҉�V)�}����	{�� R��>:5a��;�ʽy�AXZ0�oE�0�,q��X|8���*��P��(Z��m�(U�����
ٿ����A�1X.�ſ�\Q�3w��0�"h+5�y���}}8,�F��<i�V�J��b\z�8�c.x�&{�����I)����B�\� W]?h�d�<�Ysa`41w���IxN���BϾ����&(�<�H>�{}�9ZfhtV	��/E-�KP�<�&cz���Q�o2l�3`pR�i]�_UYs�^,	m~���DV3�x�j��d����T��f�k(����Q����as����x����\�jʔ�/Ԁ������ _�-��X���.l bB5D��J�?�)�T0�CF�?�_G��| y2���M��+xD%B����>xB�%|y�P?�N��¼��i�����]�8�w����>��`=sS2y����"%��$����̀����(��[���/�S���Z���6�f)�J0�MO0 	��7��JU�]ŻE���+��Y�����n��i)�����PhE_t��~[0�x�R���(��C����(�������\M���	�P)w��3�<¶����^��}<{{�@(�0N٧ P�w3�M�4��X��m��8P�Ed��@�'2�u�Hz༬%X�<=�E!�uтi��W����1Y��%�?��{DJ���<<ͭ ��!�D�Y
�YIM���ݞx�uM��Y�wNVHZ}(��;��VNX`�g��ƀ�Yw��S��A�[�镖w֌���社����j!�UO�ؓ!��G7`kI���P��R-��V�� ��,_ U?X"������͂N�m�)]A�R�u�`,�@�������]r�^Ւpj� ��W3�"�i�����UC��>�#���� �h"�0Y��u5�(�j
�&f -�u�l�f15h<�.�k�(��� )�!��J	���/�8��OV�d�����z	Q�w�x��z	3�^�G�[��>�\3�d#�Dի���4���03]X-{u�^��/�`�PWh�~�k�t0���Kj\ ء.�����4�`d������?3˯N˭q�*�q.�NH\�N�@y�W!Z ��>.铰��a:�5��,Llc8������� � 0�Rh�.�OZ[� ?�a�q ���@�X�1r� �)��h��yLk���Z�5{ �]��y��:�`aTo{���j*����{_Dt��ģ�_1w��%��|�=��Y֤/,��`JoQ%#x��D�?���2Tj�V�w����Do���p~AwC$~m@��])�A��4Ll�K�utJ��qfh�rJ؃�j��c}����	����b��	�k������b_@�S��Fnx���,b%��Jn�ѷ�����XVL	��ֶ�^�l����g��^�,R����4�]��3�f���u�m/W�R�X!����[��h%cQ���n	�}YliU����^�
u�c.��)w�PV�<r�b�1�@��R-Z}_�r���~	y*P���j��A.��x h鼒�b!���@���y�-�9���g%ԣx"�H�O:��G[�j�hgV��Y�NQ�*���g&:O3\}	0w8J�b�
4�鱗�ob�2�g`N��F�IK�~:����[�|��N(���P���֞�<x%��=Y��Z�]6�0}��9���
04���1�����ia�����%[eή�LN���'ܞ��-�v�r�vau\�_�o�1�!��9�7�߈��Y����%F�!ˠ������wDm\
-+�!�ל, �ň���R�D(��� �������L�xv'��lZ	�r��}X(XRT�:��VO�˧wJm���4� �\�T5�I�銹����}P�h2^0M�.�	���#0B�	�!bBUh�t	�	UX�}�0�f��O���ʍ� �G�}���EY�E�#�-U4�h�tQ0O"P NĘ�2��,��]P�[^r�0�>���b%�%W�+T�;�0�dmE�(1��'�r#	����W@�*7 y]h+!j[JK�������DY���|~��D�&������l�{���?��GD�x��eǑ��:�����~�S�K��H'��@f��Z)�%t��� ���]�P�[���ۀ�`�ܑ���D:חs����h�ywJn��f	X�%[�6�%���q�>��W�/D��@1^4о�����Bk�#��/����	�_��׎�ut�^\���D��0Y�:h�v�[�4T+�'�BL�O�4[�m����+O�e��54!*(�1[Y�j\�Q� Sh���O[�3鯺Z ��Pn�h����Uu4�8
�B�L�n`M�{����C��0���A�.+;����X��b20u�v 3��W�,��	�~����ZeP9�p����`)��'��z#h�S4L��� ��N����-�8�7=�X5�bDir�p����Yo4H�+�e�.OP��b�#L)W�ZD�^�VS�A���	{�q�*Zt�բ-�%YU��2O85�%�	����J��ǀ��n���uf"#�<!�^`}h�w�7͒VAlt��a�Y%��b�
��d�,��)��;љ`�l1��p��P�$
q.�"68vt�'��I(?A!&�"����h{� t`
�^ 1}(K�+4a	x�P�YU�� ��1�ܲ`h�~lYAD�U�5E�f�����J)��ч��fG$M���g<W����p�z�̢z� �U��J����Ӫ�	 5, T��YXP�h'p�W��O?R��Qrt,��L<_�J�{�͘_�,�E�$���0�Q ���4��j9kۗg@oF�2���
�f�p�$hȫi#6B�+��}��E5�Ka]�00�X�Ei�T_/����?�q!�ח_�%��f,����n���P�V��>�H<���B�k��@$G0P=ż?Vx	��XL��{lH"NK�-�V�KZ�1Z�0 R�cP��$	o��� 4(��,�S������G���+u�i���u����(���,v��}Ռh8�JO�V�3��>��f� ���CI?�Yզg��*G$�`S�J�`10���0��{�lG:�u�{��NL�Sːk��p�Op �B}�"S��pF�h�[)ÿ	���Yg ;ƈ��X��Z��=��:��K �v
�)��t,h�$��'�@i�K��@��4(n�X0s�g�)T�N�*��{ �a���T��c��C������n<@ҁ��4?z?��n�s��P],1�+%�ǽ!b�}��EH�h��	"��PZU0�=/�ĿX!�M��d�ݫ�� m{�E��X��/���-�p� Ъ7�R���x(-�2yC��B�%M��[�А&/p��8a��?�%�c��Hm�/���HYl'1���¸6�ۅ[x��S��f֘�(1��L}9B��_�!���	 �O[\!`�a�`���1\h��J����1ݺq�J��R�tp��.	�ny�i�z/�>��[���i�!�+�u1� 
n?�w��]��"l#`g]z}�.�fXW���x��G�w�
%h���KN��ܖK�D��"H]zс�/~!��+����h�'%UŅH�	�d!�FX8- m~�&e���K(>����؟b��%t�Z�E.%D ���+���d����qW�)�/�1����e���պݩ`�H}<�Pb/����S��u�Mv�~BX�QZZ�0oZ8�h��A�@��OvC�4�@����'����ؠ�#X�.)[�
��(&h�'Z]ף>���8$ULXk;OaH5�cOh��(���K�_�@�mSZ�#��{�}�ׄ*f���8�i�T{ƭ�M{�8W�ۨs�������7]/�~`�s��Z0 2Z^���QhB��Ѫo׬ʲ *BF�(D��2��O-*ـ��>-GJh?��˂��}t�G�;���fP�8;��HF-|�%�TZ�:��hGST���t0p���$,������i�0�M�����y"�NJ<���B�j�0��NWc~�z��WI�y0�-����g����	�tVY�eAP_!�,��)���[k�G��߀�MUl{YJ���;�F�]/>,�T�+C���Gg� `���L�8!^���yp�n�0��>�~
�P�{]s�%p��'�z�?�5��S90��("H#m ����	ٸ	�['\� o%�o� K-�����/���^�W����B=X��N��z��sU�hB���d�n��Ls	��~T�;)�o��	��.Մҽ� �=(m��{4n����b`��[lV>bA�h�8Z�o��m���{s�')���;�r�"w�]�1�v�P{�-T���
�Q���mc�h�&���QciS'��A�\.�!Z�	VT^~�����v-,a8WZ���b��0�ތ(�fY0�	��ܺ@�B�s����{�>�.\���ڽ�����J�ҁ;�Bl���U�''��t���YF�ݓ=���<V)��O�����_����seC�*�0�������ϟ!T��̭��%:���<�x�-�"�)K½�[�yzn��Y�\]��a���S�%#P���%��UG+'Н$�%Z$���ho|�]/�� ���i5@W�	��kت Y�7*Kw�j�M��hp0?����� V�yPHA�Z�� ���c�I^B8�� 1������r�?Ch�hw��xvG)�ɖ�``���0��$|����$��`��	���U�3��۱R�I����j���
N0��8�.�H8�& s�'!
j�����1ՅM���i�.�_5�,����Ҫ�&ʁ�� -�*ur�;kpkJ�B�������?{�i��Q'he|w/�&�G����1���h�[�/j�:�������V_o�,�V�cGn?���/���xH|Y�~�(�[B�6R�H�L+� �G��Mc��e�7�g��	��*�6� ���H��6j�ƢDS\�_82[���^R�d5P�A�N�����.h�*We�}D��J,!X�Y1��'���)���%_���h��:/8^�5h
$��q���D%(EkvS@���$c)ȎN!$�X�DH�pRhqG�K~ W�[�s�i�%���+��k�P� TrZ"�b��%,jkq�)3^�M��1��S*1�H}cC�@��bF�aAQ��~�z�����1̀HR�a��f/,!��LCD�P�LMO�P���߉���ѽ�⾒X"�jU\Dr�3᱘����~���^�rX3q�e�@�h�K-=����[SU�֋�U�������(�������iF����<�q�8�X!aFM�_��%�q��qV T������!s!�n �by���]k�J�^2pǸ�*�%5z-}o�U!�eA-0��Z�VnRw��_��̿�W��|�� �b&�?��ɒe��+�~I��k���1� ��h|�kŢP�^4
ܕ_[��D 1�^!�vQ)�\� �q�Q��	�� ���QS��e�t�^)ڀ�o��^���Y�����Z�����Urs��ׅ*X�6���@��sRuڢ�z�7�4��LE�`��J�� �H���~Xdf�	&�Jjp���B��)��������Y�hI�P��|K; ��fG�s���N�`Kl�Z.����e[���t,WÊP1,`z��/�a���%��!Jڭ_+� ��.Lh�KG��خ��%>��k+��I ���_�,�i� ��T-��A?�G[1<֟X��AE�lA��d�������5��V89����}8�B���%��g�v]�����l�=錗n��]�! ��52Yh�ah[�� S�0�[Q�v�H��1�.��N�C8�8��d�60`��349)<����w0>�2	�JXB�`�,^����_����Ly,e�Q����_9�E�ж�֥�I�)+���b��+�9�_�G�^��vt6��B�e|�J���"��h(�a��nhNel�&>�/ۣ��q����.	b��'��h�ї-ڮ\�����Xh��E��-�#9*����r��8�^��A|ML��5	�cD�2��J�S|hO������Y�y�����Z�"N|U���-S*�d_���/i��j�j"�^����(���^3v`��}�'����W�H��ZB#&_����%�?��3�)�J_e.�2;96I:t�[s�`^��∰a[S�9:� N�(����ߋ_Ո�O�,�R�f��z/U�Z�	Ee@Fh^�#XUF݉�[�����؜�5@�]"}����h�na,�`�|j�3rc�"���⃆E���cRz��fS���I�hd�*ٝ`�0a,�,�,b��U9�JB�	��� _h�b|������XTe�L�&;���2+	2�׌�DX�~%P_�������F��I�_P)/}�8iH�!�/�n�~0�,2��u��/��,�(3�����`��1�0�Mf�6R8&zp�l��>H��#SZRh
���jHqpN���T$ok)�$CM ��Z]ڔ!V�q��&�3W�%~����} �-G�o1ú`���(rH� )V�+-�Yx�Z�-x1�6�U���h�|�W��5�O_U�M9|D�4!������ݨ`��V��o�,�1Ѓ`�4���%
[�@�T�RW���V�W;�˵��׬�I(��X5�J�y�*�z�VA���Aj�O[8< �9N��W�"*�_��p� ��Ii���?K�!�1��S�0�Kh�e�x�N�p\�2�w U�*b 	1f�d�AT-�c$���K#O�~XbV����YRUZ����]�&P��S�:�=�+��́�"���j��'Z����U!`�����a���W,K^���l��������1sG	-��U¦�W���vU	R�ojrW�!�-]��(�!NR�'L�шhZ�o:qH6(&�)h}�M,5��G�/�"J)��6aM-�Qu
 &�%]gP�w<�+�PB�]Q�%AL�i(_ �Rm.v1�o��*�l_�n%uK��oȯ����ô��.�@���|��p%J�cPu���K��T����]pzZ<��}(/L��P�o�&T�-'!�ܴ�`,@6(V�/�ۄ�1��^��[�O�Ū��H#�� �A�.�d�ꩠ�\�.�R�q��T7%����3�RI �.71�|�)�p�	+j`8����0Z�iO���}5����馏��Ga(��#������ �Z$,��=[Ìݷ���0X0�Y
�%�Hǈ,��tC28	�BD2��ex�%!����w ź�*9W�B���S��\����-:o��r(޵)��, R�L!�P���d����RD��*��%4ܟ9[�85�*�'h�'&�Z��_�]�zH�(%WV�?�ؒI1g�S��NZ�|� \n!��o����羄��ŕ� /k� ��V�@��.f��#D	�-������^ �5�K |�)|� �*{B1��T���ZSȑ[�a}+ ��(!��&�(�~�0�����l�(�LZ",��'�j���bh<K9�*�,Vo^��dj7DXd_�̴��E8�!̛)N�)�z�v��n��>|������ �R�g���oğ�I�C�_h0�-�*(�h%R��[3
d�)����sM@}Oג�B���\ ��a^U��v'� p��U��\<��p	��j��17�(�,ʬW �ALi1�N_�m��<����5�	�Xw�j����q�Z w5���[�R6��^3��O�0�jH&>����{~`|�y������a�0<(9�X�����U�x2ZKW\�b�~�B41�I9�-�	�W함|\!_@���B�)�@��z�Hͼ�(
� D3�$�/)��NyR�y� ����F)���N및"c��fP��!���r�_ݖu'����4��SUv.nNҹR9��⻋���h�a3	�D���w�8��ۻ�w�rR��������*�V�A;��ۼè��v$B�l���S�uP��鎯�4��Z��fa�j�@��kIG�H/���8��hV{��g��쉷V�X����%ׂ�g`_�(u�u��X �09%�HUY��Vh�AyX
]���ݨi�I/x]́���	��a��� ��\#�N�}l��0�`J�,O#	0�$���@ȕF!�1��	�� M
����O�� ��Ti�p��FX���S8�+��>��3�@�1�I_GN�~K���[<��+�[�`���WY��#8�	�O�da��@1���RS�w	x[N��߀92%z1���f9xh�mX-�	`v��LJK�	"Z� 	z�6�CAk�G�!�ٓ�Ǯ*�T��rd��`c?J]�ӛW����B4M�'Y	ޘ4����
K�?�� 0V[#5�`�)�_�Q��T�C���	:�A^��,��N��4�'x~�|L�h�wO-N �k�|�H
4"R,!h/�m���N�(��%���C�O޸�(�	�c���܂�^19Oa�+�%ܫ��u���v�����Se�x���KL�/�&Rr��J�
׌;]�
R��rWh����^���в �n�	ҫpb�_	�Ѭɨ�F�8�4A^:����*�ְ�(S����Nx��=n��N�<�b�@���3��
���P��i/ آS�&hIX�<2��}�Av�e �j 
�)�Z��k����(@g�� #�� z�33C�[���$Xa� 6�W2��\PA�i����;���x��,��d�8AhUd�Y�8��[(�,d��!�	�`�Zx�+��A�#?��A���/n���[2����8	2
F0K[�P��X/y�3��	U��	�I�T�-K���k�\�@�9ow"J�xˊ�W�S~�DZ�?��Ҫ���%����g��HU����D�P�5�y���~K�D?�@���RuYʓ¿��h�d_�����y����d
2�E�Z�P�]xA ��cE��>�G�
�r�&��e��'������	�h~��m�F0h��W|����w1��y�)'7����-�@�G`W��~�Q�ķ�`.�S1�&PJ8`��� ���A�pl(*h�	�XE}��1Ò�b{��w���:H~�#���j��*���`v<��[�zx(�Y���|T-��� �Q
'�%?U�N��Kٰ(�`;`�Û�0�-)�1�.�B��]����P��>k	B}S�B�X6�b���o
=��� /���������F�<�A>��������Y���"���H��@|�e�b����n��=&9��?�H6�⁇\��E�%wt��Pƈb���[��0ZhE�T{���0�� "H �,m�`��V.��?�wY6DV`ʅq�	 h�,FJ殿���4E!��|�9h��N�l��� �5]�y��^�WjnW �~A�O.1�3 Ph�
F|��Ԃ�@�S`�m0��RBP=���9��l%�ݪ�3Ϥ��=��Z��`�j)�� �$	Sh�F Z+X)(_~�?CA%_d� �G ��<��hH_��	zS��}�������<���U?t���>Y�J��&KRI��2�'�q�M Qh�/�w鹕r�~�s�	��_�	ISO�)�� %V��5*�$�X�QetU��^.iH�	��V� �Z������n�6������L
�(��%�d�.)�Y�����c�N�4���-��v�K��e��l1��`�/	-i	��+������Y���x��h��0E��y�^�� �-��0�hK�b�ڹ�}ՉM��G&��fɨ�N�l`��H6�0pUo1V�@�^�~�n�{�"$T��\���	`(�7��~%A`��]�v錾�Q��r�/��P/���� }W�S��_�E�Z�Fgv3s)�_��*Վ��#
�Ƌu�(�/��@a�&�o5�<�0��;�2�\�)�(�$�X
�@4�J�
9��f�:Z�õ���#�d�oH�.&]�%0����ng�d	��BN��+mA�XY!{��Z���w 3��֮?�o ��������0�X�ꁜ�4��f����t�cH{� %b�*�����a�W)�?�~8�I^�_�1��{;��)Y_;�0i�j��q=���}:MÊ���~l-��UQ�'��h�Ot�����l�鰪^�<l �k<�\A�&
�nue�-I���M��_��Z0��T���Q{ h:0+�j�
|Sy���7'(RL����x7ޡ1�ik��Pg	o�f��l9N�<�V�#�����d_R��k��
���P� �1��,rU��j��3TPve^����w���������"�0̻!'�_u�(�Z0g\��MEJ t4�1�/[���5hVm�&���Z�jUıY�:i��oyV%Z�вJ���f&J�=5�n�Hk���B2]�ܗx�� �Z�ȕ�-��n�t�W�u>�[�!�PG�x5h^r�	"8�njOW_�.ZXC�6')1�5�I�$��J&i 	�	�\޳_B���q\���N6��ʡ����E��B����Π��*o$&^���΄��`K��ES���+]��@�!�ޘ�)������Ah/�y��	�]�p���4vm!���?:���Y[Ϥ 8/{���6�3����c�)��T;�zA�Z��'����pi;�}�'A��Y�I.�i�>�g���pľ����!=���4�^-����!ÿ�m�T)
��+a�,� 	.Q1���/w߿����z_�<��#�}|:7ۀ��%t,\1;ϸw)�x�
�r�N��t����<JA�g/�9�yU0˾���<®�������1��^���E�����ϠBT[j�F���낤"�&���1e!H�գ��)ƨ���j�|% �7���1 뺾M���I�t`�h��d�T�5�Mτwm���-<e��ĵK�UC^�ޙ�/�4��Q��|�0ݓ�'`3טn��$�����#�"� ~5u����x7��LY� X}afQ��� ��h�d��(OA�0�X�
2w�s���Զ�� E8l�,�� �"d�-	�7�!��W�<[۷�)� �d�_�Ko�lP�	��r[C�ع�C-UFܶ�h�NI�/Q����0!��->\&�5���J�v���hkȝ�%hs�r��W��W�qK�[z!�(��0z�r���Q{�s�wy4;]h�=s]	阕�W�B)�k^� ���x�.���J`(�|�G�ِ��>9��T�=�X��%�R���%f(�( |2�Ga��H)�Y�S?00�8Q;�W�m�L�O�(1��5p(���� �N���G�&��\_�铈�p$��Kip� �]�n_h<*�fՀ1�0[V3�rM
-�k� B��I,�֤��EXm@��=�`���^�_M�	O#S\R�hHF���
2f�X���`^\4�f��k4�a�S�� ���8��P��8I#�CJ����4Ї�k�9�^��RH���j��N�N�!�$����K��/�	i.�ٸ�8P:N�a�^)�-E
�����ڄ�)�~%������Z��.h��E� sQV��-��	����^�P�E��D���U� �h�xq9X5�zW"V� �^�4�	�'�&#�%�Ms��4�,���k6���
����3��f��[Zut��U@�V09_�����2w��5��w�&�� �b~�<1��X���,n�c�B{��yepܲ��!�-�|@����sJ��HE���x-��נK�fMd�'t�*h15�|�3(�ZȀ�T������
�:���/w��XH/|Wh�جA���uEe\�K��5%���Ʉ�:��>� ��~&E#, �irL�L������K��8���� �,Z(��C^K�O˅�ys����
0�4E@�P5�^���\fd�D*v� %^hqEaJn�w��!mZ�D/W~3 Uh�J]���(�ig�)O�!R�<�)x"����s��#n�[(t`H�a�H�޼%�4Ph %Xݎ���W�����R�����*	0�f[@��s��u��ԋ��]��������?[{�*��������#�����5xK�/W�~���hUp���@�
�Dc���)�;Nj'�[��s�`����z���x�M��&fZ�ٮ��=1�i�r��n�/P�� �p�qu�`�)(�-v_�8�h
�hR!��P��6V}	�̮���<p	wǬ���!�~�(ɕ�=S�Ne�XvP�J>B�'޻o~�O�d,3��&s@��`.�Hu%,!з�D�{}���UDﺅ���]������3�5dB�@�%(OF��Z
��B������/3VyK,��W`�_�|��XQb
4�Uj�v1X�r3A=M�l�	�u���^'J�I�/�1)o���:B��}ZK�c�}���HKO�x�a�h�,¢7��QAbI�j��\!��0f	A)/� E���3*��"��^��Q��-V����)��p_PE���œ�����_�l�;n�P`�tW>sh ��&%�q�ߕ�A�H%o�G>ү-~h~#���Py�O�!|ݽ���h��"�	H�f ��w�%)�~��W�����e0S���2��<��2#v�>�[@h76k1���N��E�����Q/	Z!u�4�t��K�` 1L���ʸ��CL
a9o6��� =���!�X	��3����荁����Njf�OJ�/?�	3�b���5'�&
�>�=`%�v,	�a�l��σ� �v
���{%}2�\�c�TK!|GLE�Γ ��!�4���7��.��j\E�^�<���2��_]��\�uU�[C�v�/�5.a$��鯦�^���<-��:ej��*�^�R�B�Us^�Y_���D��?*Ek�}�"{\ �n)0�[|�t�y�/�-pl��(��e�z>���B�cd�u���A�%�u�H�;�m�g@ �<��xv�~C���
`��騸���� �.����(?Rʨ��W�t����Qd�	ݹloe@��90!^`H.`1����i�)������!պ��)���0�h�p:�\�Z��t1d
9撁�wg{�)S�~�A� _�8:�2��v.��V�yZ듸� R��>.zG(�?ݺe�J�~���3�[��8v�Z�=��!��a����C�U�E�Y@:��ݡ��x�����/����Ŝ���B��2k���H�C�z@�ST��X .�%5�u�K��7���O�H�	��9��R��^���W��[��V�5�-|z������!�(U�H	z��{���-�=֒4��=�f-�^�o���[���\�E%Z�D�Q���� ���X��1�~Σě2��Q��/{�q���9�[f�W��G[�����m}�:+�0`��P ����C��.����8Zr[�d�K?���ua�Ƥ�%O��9$�� eaL�(���ː9�n/4�lٳ(z	>x#+� U:�̶t�XRv2d��1a���~�P"�2o�KM�͓@�m �CH%� ��j�W)�-�����Ul��{.iu�>�֒N�R�|$��}��F	���/L�"{j�d��y"qP*�+�K������J� �h.UD+_~h�?�F� [���x+-���PFZ���v��	'�;�'�S�c&� j�� ���-�7�>� b[Qhlw{N1�=���p��0�)iJ�%Sߚ���H������X����tRK�.a��Q�Y�&6� �qʋ�}�����ށ�	"jze%ѳKѾQ�l�1ʝ�<ʻ$O�꤭���;�X���P�=o�#�K
,�h)��\�	[vwN�t�@)��5��D���h%@�G�m�z����(#>	����!�9�q�u���*)|.��}`e`�J�>{�P��4Vf_#{�kؖ�[��cp�3���@�h�;^����*^	�<�� ��o��X�	>�O�N������jĪ�
�}�0��H��h%k�p{P}�:�X�>[V�T^\5R4�qk���I���h� �7��Z�U�̸;3&�T�Y �
Ug�xEt��$�����0p%���:��e|���\0%]Ә���|��L��(�Z� ���d*��A�˞�s��w$W0Nǀ����n�~y�PQ�e�,��>Uʨt�RW$fY��nL�v+�x�5�RB����W$�D�_AK�C� !%�t1�)\ТZã+��Hބ�@���. �|���G$	��d�_ٕ'_�i��9��d��h$�R)d��e���Z��4�M���X㤑��Sn���]�}��E ��?�cW_F�M�q�/ɋ�t�)�h$f�����)ǰ60x�h\h��G�`���2���G^���f	{~�̫�sW ��*�(@�ذ�	D�8�U����9�S̽>�!��v�Wq��א��e>"/)߈�
_S�9:�,��[�#bXԛ%�ͨ-�6��@��C�zf8\(U��Q�C�~)���O�ˑ�l�t�`��F���E�~��}�\a �e]������T���@�SP���o` i!M^� "B�>�6��\R�O0�dy#���/�h�Uk�)-4			�2X��y�f��0�Q�O�Q�V�@����o���&x���������^�*��/�;</�`j��y*����U��h^��R���0�6�b�xɀ@�z[[}Q��1��8�x� �wIMl Z��'�c���:yE��p�*0�5� Z�v1��l���R�L <��[�ᵼ3.Q��^/u��̇�8Z8z	C����UN����&
�n��	�q� �hVN/%QZ 3�ʡe$�� ���1ְj�Mj\��S���a�B��a2���vi=��xO1�� ��5κ
oJj�⿀��=Ka����Z�)�����Q}����]4����R�施 �%�L��^l�ON� ӣ�w�u�;��Q��'�u?��r�8v�C��@tXG�:U�)W �J�Ƀ��_�w%�4�'h�)=��Q����h}�5Ik�;�0JѮ)�<Ɉ�VAh
�D}�u:	v�)ʅi���W<�(��*w r}�ĸJhWA�?��V�O�-�A��:��MV��WG�H���)��^��h?tdo�Z��'XY��8@A���>�`^��mF�����!H˜JB�bU�iV�A1���Smu �-���;�}j��l���� �����A��U1���E�F�P툃]m��>���k	w�w
O�cz�A�a��}�h��-'������ø�ֆ�J���,_A7��8v~ L��yMS�3�b��^
��)���w<	�1�X��#Z3)�1x ��~$Kk�? ��hg�w�=�����8�ԓ ��g�S�x'O\�@~.J ]�:e��×V���yw�	�Zנ��h����� v�p��1��r����-�4��a9
"�w- �tR���O��T��C�Xr���ZBh�}p?)+*�d4��~V��M�/ɼ?/�b��1w��_��P�^�?����vJ�o�*�h-��@�6V�!�P$Lk���h�Z8�ٹ> ,�Ow���HU��$�Ϯ��	]hm3w����
u؜Z����58L�?[l�AYB-�f�	�Po�te�[;AWP�45aJ� w ��->
%��[�V%���낐�p����w����Ȋ^�\�D(.��|�-Y�������h�!Y�	�(g{	 ����0�haTQ��'�]Nd�ڰ�JH��t�_P0h~%�'��<Ï�d�h�MY�%s;wf,��Sp
0�fQ��(��#.�[Se%�`��opHM��}<�h70�G	P��s�|�Lj�y��c�V5����- HV�2b3.�Y	h�y	���Vq
!C ��@W��bW�U[�����_�p�jT$�~�A��q^7��kV'0)��n�^m��&~5E��!���̷0����	��S��B��G�`G�T �P��I@�pIS`l?�[�X*�T'F� |V!)�_L�Aj��$c�x����f�V�o �(�����h���?�J�%��7�?ߪ1�n WR��TK<�@�B�É�� =����T�J��鋞���Bf���Jk��(�JH�)�/�X��HI�jū��q0	|�a�_�X5�]�_m���XN*`��L���)�����������LKG�Һ�}� ���tQ���9�p�$/3���`�
�~A��Lj���JL|-_bV阳1Rk��Ɋ�s� �Z���f��WF�<p;��X=TE�ݠ���1͘� �
��"\/MU[1��;@��	r��
d�A��8�#�Hs K���1�-�s�7��B/�E�� ��u�c���T�^s�:|�d5,����ܐ�[ �܎k����m<W��h���k�YH�O4��R��0�E�Ș&3Zx��D@U�����#�^jԵ���B�7-`o]���9�z�����K/�;6�(�(VFTJ���3q7Y\.6$��%���{/����Tt;!cA��c@�,Z\��5(�}E��\+X���%���	�����-x�8o��l̰�(p4KY�v��R�����u�+
a'gW��.���'����B��2;0oa�g����^�Ё^b�A�=򀾜 @k�Ο���a�1��r�	bUsJy��h�02ａ�4�\��7&`[��	
�N� �y$d1�颻�;-9�����ϡ?��:f=� �6k���(申 �g��B+_2���� �EG���n!�X��i�i���0�d�(�|d'��o�W�q�|e�XKW�eCf�gP��Vt$�a���	�D��B0w7���d)@��pv!5�#4'�/�	�f�@� ��)`�,L��=��\��4��������?�S�Q�6 �*f.hJ��%��S�˓��Oˮ��%Y�f�T�?�܄W!rӗ�p&�{����_F?�r�Ox��.�d~�������h�T�Y-yn��g_a��>� 0�������u��)�0&V��O��o�_��{se���y�1��1�Ut"�y0�}d2N[�!��Xc�I? -M?d_�5J ^���1b�\+�����{vaH����P����0& S����UӐ�Eu���%��\њ �=)�cˠO%���E#MW�Q��cp|h�~qW��=�1ٛZ,<��n N5�~�ԃz�TzG�^"�1�*���G�z���=�	-c�;�0J|��'{�\:������.�Q��'+U���VMy�ZNIc@�������>|z-V+�f������:�纉̀�g[�нnA�_� ámx{"�J̰_�KN}�f	Lj��1!�	�p�p^v��6�>!��8����qFA��nv�\Vr~����#�wO=W̹j�8�� �n�D��ܲ� Ycaq3C��@�U}�T�J� ��f1ʕ��@h:�O���O߮`���I�.E��1��L�,��Q��ş��hS9���e'�|�/YY|J��3��6�엵H3eH���PL5	�/[�� j�=����a;/��U��K��z���7p�,���hNe���1��^ ��-xt������ַ�W�R�I�F��P; ����@�1.�PGri o�U@�z2_�fYߠ��3���*_s1�h�+�L���%�)Vl��kW�i5=$G� ��g����rw�.���#-N���o>J��jյgu2�\愞�h������jȆQ���ɀ��	���:Us%|#aU�DiP��¶^��)�@��?n1R�4A(u	 ��ڜ%H������^_T/h�V�Zb�\<�	�D%�<�*�[p���W�o�c,�������2Hp����`�G8�:FΊ�B)�!�10A��Q�=5�hY	�x�LW�wC[�i�������S��pĉ�ã1���A5 h�9^G)� �	��+�=uS�r\��Lw�I��_��@>e3�"P�[�hˉT��ס��m:����ӰZ ��<ނ����(��_3z�;k�1�<,&���ņ�Ӊ���yW%ZQ��/��Sw>{,£���d�����J�^�pj�U7������W�E]fm �F����?1ڧ�T�%E6J:�k�k�\P0�3�\Q%	r�ol��p 2�SqH{.ʸ{5��Z�4��H�b7_R�F����Q�⨖���������V=�C���3�^�i�YX�r&� �Z1��`p��]t`n�֌R\��j�^�F�2��>%]ua-د���]��b'U0�E�u%�˺���h9j�����h�Y�W�W�Q��=��"?�7LQhQa)В@ܴ5�`F�*�m���Y�>/j]T$1�ṷi�{�-�׾��,�s�I�,A��n%��R0�a��TO��e4����#�X�{� �	/�P�y���p�Z���2?;��S�{�����U�ex������눢�v�&5��d�e/�-�*��(�
��eg]�˿��J�!��W�1�MT*򥥮�*�w녗�O(CW`�q��1 Z��p=j��kO��E'TERZ��EA�����N1�3޲���/��8�	�h�g�;)I\�%�:�����!��$+n/m�ִ�,wp���M�Ln--R�@tM	�!��w�^��0����R `�����78bM�IX� ��1�*���{�l��uF�<V��\A)�^�q� �R��` 1ː��{ɯ��u�}:P�K�"K��F�m	�j=�s��4P�M���c.1Fy4Y^�@���>�`��}�τ��,���q8e�����Qոp��[sa�%$ު�Jm(��X��Z��P�FbJ�8��_��o�`3�A��sz0�dT� *)XZ��C��� �;�6�R�@Z�@��l-^Y�}�*����h��V}.�x�!H��_�7�5�w��_8	���$�oB�B�ȀGz$){��L�ݱ�����9(��7x#h�XX��� ���G�:�)9.4���B��#!?�R)��i�!]I	�����1�P9-!�s��V]L쀹�?D��c"5<2�S�4�� k���ɐ<�[@^����-0/0f�mq7��W���x'�Y�V�4�aaU�Ő��T�S���Æ�+�}��x@`EZ��&�� jD�����+��z,;P�D��w��S�Qg�|ׄ����d &�N7��W�|]Q�F�uYZՈ����K����xXr�J2��h��?�C�j'~!����N�\�DZ���RO�S�У���d����?M.[�
�YV� f'x1���S]R��J��5kgI��Z��7�'lec�@R��s	��W�I�u"x��F(��d]u�������)�7�a���`c�� J'�
A����]-eq�l������dQ\J뢈���-��5���$�N� �������Y�X��PlsU	�lqZb�?h/��`m%k�T]gݔ�
�8� R�G?�q��j;9�)Ep��AS��h�K5~e0�«��ȮV95�q4�ӝ�oF����	�, \�EO���2��*A���E3H`h�V����%���0�J� ���#��&�$���
�X�1����-*����Y���Cd'�����ǅ�h􂨎��W�B��ڌ�[�$��V��.�]�Df���e N�F��Dh	hU,0�zy�2��bA����XǬ�4�Yv���f�|p
��	�Y	q��> �yi��'^�m�ԟ�1����8{��v���4UG��M��j�4IU3@-!b���f�GK��1�ak*���K�hZ�� -������s�_�G�XW�os�x?�O��{��G���Z���>�]�A�Ը�V�6���)�c�}���㖮H������E�"�*a��.�!.�$�_%���R�E	'��0��R8:?�ظ�K�H=���u�)�	$�u�1����H������a�hǫ��&�-r'u@,�6%�j�g-��}c�(3�����2��!��	��Ea[��0�e�H`�s��8-XQg'(���ϱ�D���/��z��,1ru�S�5�A�Y1+��߉��5^��	]�^���8�_�$�Cj ��](�k�!�@�1�B!#_2pz��r�����a������a?0���b��g��-���>0�U���et����e>&�+<Vq
&o�Z��2�|[�?��Ch�]1� ��/~GB31Z�@�0�sSD)�~^'�}G�9jN�"�l���iB��j�9�_�P��v� %�!��~>�_ �!p���8(�>:v�W���_P�	�X�A�ĭޙp�L&�c��x��)R`��[,�T��uL|�o�GҦ��p>H�!����0���(z�xFH��s電,�~~lp�!�z�M��@��~�XU2��;b"wѧ�R$�Wn�Ӗ����s �9���C�����.#�0?���$HG�.�-霚�/���v�ؿ����ۍ�}o0XR�M�h��l����/��\r��)@-�@pv���^�:�2Wi��; ׉�QOX��U���'����5�l
��L��4��fi,@?��?���V@R`�}8�,�R��Ag�!u�Xbj �V��|�E�D��1�r��T����l��u���d⟓�9*�p_�M��-Jw�~`��t���<��v�y1+[�hj�]��o|O���=�")rӕ�k4#� �+�hY�ςp��%�4���
^�	|2�s 3q�~����e`H 	1��c? ��B!�)�h�Z�����xN~�)#�A�	�-�0�7/m�=�A��*�)�c�����������Y��u�������$e@�1�S�Չ(w�D��Z�hLz���H�%X��ј.J[�Z�D�
AעItJ���/�>�@�T�7fZ�ƥ`�Ł\6yJ�4���1��]���B�:��jݿ�q�S�3R�#P] 3�s}J0|N�h��%T1w�E'��s�Z)wO�P�VP����,k _�3Y#� �u8R��I��BTFu�ʃ1���ט��	�� �ݰeS���r�[��� ��&(-'q
!� @�;^1�īAɅ&e%��A
Au� ��[��K�l�R�=�_�x:5�~�%_$��%�0�V��+�N_�~�		�l���j4	����;v
��A}Z�]�i�48�7����Q�E��JF��ף� Q�l%�'"X��ç�ÄD8sU`�#yv.AƻaG��0Q�&���X����\(�lT"�	b鋊�:?w�<)���;	}Fo ��q�i�H�_��jLp.�B�/.)t �uH�3��A�o`�Lw`��nQ��.J��
Z1)~�; .6��Q2�}@;���3I����f��޼6H���x�Tr��">�3�h/�^To������i�-)A���Us�����w������_e��SW+[_��C<hWK�D�w��U<ӯm�nk��
^P�24�৹e�,��:�[ATp���.�<�NTp��\Y��8���93i*��p:g��]ǩ|0����9\9���N|��i��-�HB]�Kݻ#~,��� U5�BO��R&<�X�W@���`�*�1�-)�L�����
Z[h�#3���R�S;�=Y���� �Q<ru'k��hA�[����_���97�-Q%k>���"�M5�]��Wpb�uDu�@yZ�|N��o��3I��Ej+�C�?0�� q�Հ�S������TY��e�!}�4`�D����FA��
A��Äݾ �I.�� _QuC�zP-�^��h:?�fy�ZQ����8fgX���Kp�뗺4��9�C�%&1L���ҨZ����F+h�����7U�Ž�3%ZF� ����@���I���7�����qht<�Ӵ'�t�-R� �a�6�\top��1n_��]_����˸[ �2�A@%}8��JM�MH�E�'i=mQ�:�cn]�b���(ޚI، �<�DJ��,"�� �@Q�Q��Aw��;�*_ ��D�!ѕ�U��Rh�oa�����#z靨�U�&w!����1�{��}،�2�x�x')К�P|��	�kQF~ցIr�)D$�
/:�/�l�|L> �z�x��ӽ9�.�g1�^��O!��9+�e�0�p���D�:��j��RTS?<_���Dq+�p5-(8��r��J�����[&�P��I$8�,�ŀH8i��BK�HL��"��uL��S�`�3-X[�}�����R�y0[���o_�v-h��61��0���=�ط�a��4Z^얨hq �3�U#��(���l����J����sZ]py阝���h8}^����Y�;�ow�e0�h%VF���t
ZWVv�pTR�P�k^12��@.�b��R�^�.�N�pM�E��AzNm�1�Q����S/!\I�z�OK�w������w��Z�J
鏊�� TsV��~C�z��7_j�*����1����T�ـ������ku���Z�e�G��5���y8��]_?B���66W�@P_C6&�u�b.	 �cZ�dX{_��ǊNIW��B��B*�}ƿcW�����Cɻ�S�F���ڐ7'�EB'�1�"���(n� ��th�H'�Ĉ����:� MDO"����n���]��>
�V��1�����}v����a0�^
9]��i�ok{&e,���U�;�]���C6{�6D _��>}o^V̳�	�&�t~�?^�͚P�-��N��d8�h�X!��k*a��R6�M�)�ذn�z���b@R���V��j���Fh��	�^Z_^3T(=�� [Yh�D7]�4�ag)�`���V߫��M�!>�>GQ1�DkO\J�/ f�8���`.���r)��G ���w��[Z7�L�0$#�\dz� �7�>��)���`�R�	�V�`�tZ�XdY�1�7��1kQ;Ы� 
KF�B���_���0x-+�Y�0���2>%��X  �4�b��UN���U_-�������`4ZO�������^j�pYv)�M�u�zy��)-[ܵh'��K~�^C]�wv\�uJd��VP���_�f<B��@��]��	F_�6õV�71���!J��a�B		�ʯ���jЭi�h�Y{i�����Z�{���D�Di��~���u�-L�΅ ����{{���&-T�טK�_��R'^�2��z�K�W!?CY�bh�	������F��*'0^�����(�#	�\��_V�4Z^���U�bb@F����S���7�~��^�WkP? A���ݙ�-x˗�C_{ B��� n
���z����:�C�Ґ�����\������'H83J[����k�c!Q׵n��8�4X�0�hp���TZW��� �S��F/w���uâ]d�NpGP}W:v�pyu�u���^ќ2U��X}���S�kp��Z�#�L"Y��B����m��Q�_F��� �81p�)@��|WEɉw�p�hn)�x�����~�ohM{�kK�Ac(w(�hzÂ_8g�0MXo�WV�,;%����rdw06����;�"��)��Iq�c��T-��}kF@-�;	?�3��|���.�	zm/���(i��ͷ�r��q(N �̈́'���!�c1�_��m��R��O�0���Y�_�̈�8IN���1���h�z��ė�����t/�[h(&���a�D�_ 0HB1�^J��Ԃ�:�����Z�]��4�7�#XM��*�	�o��I���p��9�#��\hu�'ZB Os��|��M$L�����A(��L3v-�t@�O)�m5�9:�+�g:�%��ϠU�*-�}._B���4�4���]�:��5{Dh#�m���]���}�;)�/�ĠS��/��~�:~yl�ւ
j��)� ҘC���u"�dR��l��Fd�WQ�!E�����܉I_��/3Z�K��v��_ʱࣶ��,8�tc������[�
(���ϳ���R~�3��/��
�:_���y�^ �w��- ۅ��sF/���[��ӯ��n�#�ogH1��S�`�5�&�y�� ���?�)O髀,�5^vD��Ƅ����N_%I�rt;u��
bs�~�
���\��LK�d!��p�ʣg�Oskr �U'�t��Ѷ޺� �)����$I5��Rx@�M�1�)� ��b!pR�ŏK�uD�O��|qV;	閚�1��#�����HJ+�<@^/h�G$Ȉ�AZ蟏7�`$��
�3'E��N��YdT���G�T_���4n%��eP�ݖ 3�_u�)�_t�� �N��5*���Qw�ƔZ��	��ܖ�'+|I/y����4]����u�[��j�c�{��*m�1\�,8u������F�8�&JH�� i�J͉�1�-{u�9A���@RhdU0�ZVT�z=���W�<�(BE��0���Y1������_���[2����#��_��%�1ط����	�6_���2"��x���/��Q*S� E�)�Y�P��:������M�s�U�YN��ѨἻ.�FJ?��w}V�n	�{>�1O#Q���x>��nSP�)��%OZT������C#�*��l�}���L�y"�s�-A�΄��:����͠4 d[%z^L�j�S���3�$x�5 جnu�	��oV�� =g߈��-aδ���)�[� ;���<N^�c�m�c\�A鬱��B\R�b�����E(�z��z���ϒ7a�H�"n��h? ��gaK���9z�ė+�0f� :�8��Q,FE�-�23������틉PP��m�5��%�E��P�d���]/A�V�c��Mc��&щ�N��0�<����a����/W��C"�������(�µT^���1�eKb����j+S�&�`��mk����b&n�lv��\��NA;5]6:����G����|^<h�;�J�VY;�*���uөЄ�	��O���-~��ښ�!��������U�Iv���fY��P��QԽ&�$�{�Y~�}��AT��P-�K� ��p���W��}Z1;@H�q2l�/%���Rr�.$Ѐ ;A���'�YU��9R$vCo@SU[]��^A�;_7 ������x:$O���P<�D������7@dUoX0	�7V���_�\PK0R�273K+��^���e<j�׻
�
`�f�^� h�7g�!�Y�{#��r;NX�9�@;�-��r0�?�L>�����J����D	���D��t�n�IS�3��JIue��0F90a%�;�h�ͽ�����ž@��`̙z�й&�ԋ-}��L�\ɼ,�#b��Ì�8�J��0:u^��{	I@��~{'�DR���������U�{�<U�O[��!J��!��N.��h$e��1u��T�V��c�Q^��m�,���\��:p�	�]�| �����w=��]d��j|\4���_o�`+ �	G�1�_��������%�cҮ���-S��9*�i
�؎'懵��lW��u� %Lָ7XscBr�������~�օ�ܥ���m_�$��V9h�8�&a:���;1�߇(�Pژ�����}j5�J(�[����P��TH7	��\냼��8�(��a����s�_2p<~	��r��R�YB	Q}�L���'��F�֟A Z4a'oe�c�&�ڟ���K�N�I���`�d���Eb�U��I� �3�1���Ҫ�H.��h "] Z�G���W�U�TJH�a�'G\{`��B%��@�!]lYP��0}�VT��j%j����s	X�:@�~�L��)�����S/h4�(I�%�j*@0��<���~61\���.z��9�:��[��RX�Ż��Z��"��P��-(X%e���.@E�t��;�*-3^�/��[_'�8�e��2S+[#a5*{�!m������=}ŪBU���s
�x����L��"H��} 6?r��,x�JU�� QV��DI�B��O����?i��Z�q����Pe�� ��x4�r	0�@��\-�$���_�!�q�W0=(��%�uc&]��.� �Q���r�Z��%#�<�J9��4��A�P#n�7 N�6K[,�0�!�&��;��J����Ц��h�H�.Z���B�,	�[�bV�D��1�+�&-���Q�P�U錗B�_O ���PS���4����rH��{��aq�]��|�}�hM"��̸�x�ɹ_.uј\�:0�on�
u�E� /;i5K^lsA��)z���N�s�����WP:D�U ��I;a��rc�{�=�d���:���o�����0;�jxO@�w�/�4�J��p�yZ�y�.�)���n��א�A�_�j��s���.pk��S��H����ރ�x��
0� ����Q�>N�����0�צ�6	F '!Ż�<G ЫH��)���`D�t�h ��CwK)'�]׈Q;{�8.|�4��Q��v5cff���/�'z�2�N���1t۝ �?b�;���𡛉rKBS��m�;_���@�����?pv#���)���O�+���g^gХ��K�˾\m%A��>���YV�-|�T0�=��;�[&��Z�{*��F[�A�02��)�:�< RKWu�7O�2aɢr�+���Mu|}�-t[�
3�L���j�0���	,>dE8'.s�O���������%	ZQ�vfi<6���e���<g�&��VA��PqK��A��U�*�^�1��R��ŭ_����3�B�U@��F�]|aiqV�\@9��	="AeyF�u�<�8LZ1_��epp�:C� ��H��m�Ɇ��u�S(�vZt̸_d�&�����
��Q����j�0"��41� _�?F����s)���5�|>��/L���B'>��v��+�N����>� �(@���F�և�ϐ��?f���	��i V~�_��)U�� ��*�Et�[`�Y�eC�t�������.5�N���@_L�(B����Ձ4�(�>���h;'��#h���5��RqT^����vP��̟EZ=�ĹF#*�t��9,��$��J���� �ѨP\�X�ɗ�4*cf��	U����.Q��	m6����Kd��,2d�j��h���B�Wv0@�e/P�3���G*X*$k=b����B!�qńhxu�|���y�Ah4��!�M?��*g��e*�}�q����h%Ja��N�Ѕ�<�4>[����qO�o��[�ټ�:Z[���4+ /�*'�S>~��g�Ep(r��1��"�hNr���(����p�x �,}�&1��%�(_Ǵ?�%�b�o���%W \iY��.�Ih�/��DK�v�/��cΎJ��
���Q#0(�1���W��a�QP��dsJ���^e"�h��H�&��'���Ƭr>�m0-&vG ��tb�	`{Gxu/�ɆUXi��RW@�h�X���&a���#�r�����l/W	 �1C��7a�\������c�Hd=魂;I��h�U!<:�l����ӿtN�r�3��7��K:�"(���������yr?_��-�[%Z���{jD�x� ��WhVB
��$/�(˴����fgc�����(�%YQWfD���&��rڥƵ���Gjp���]� �-�͙-<��6�G�8��� h}n������bLz%3[�A0c��j�,mw�bv -F9׼� ����	)B�q�#
�]!:�6��WQ�b��@�Ə���1�=�(4� ���Q��(ȯ~� �=�n� x)ý	}Kd��p��ܰ��X��l��P���Td�6\��b���-׺��L:'@�-�KS��A�b�� �	�8j\m �y����$;/\�Y<���&�S���0\RI>	|Y�P�6k�.�K!�+0�`�z��b� �EϤm)���YMZ��n��X��a�;Jɞ��� +Vrzw�I��X�q5	8����H�Ӈ!�	�"QA��@�n��{�1���Z%B^T��pJ-a�D !��a$�u,3"%�n�P���g|�%�dH2 ����\3w �Pc�!ڗB���$�Ɇ�;�Ƥ���&�JL�? ˡMk�O�.����*	�^�g�]�6�R�&�N1m�]W��R�w8W�|?M=ʄǑ�� �ǵ����)�0��cu '�#dT�&��_��_*�;�O�����0RDL�8)铘��\�z��S�� v�g��Bt��5�"�\)%�[�@��n����m<�TM(��ܴ3���P4H?�*Ze���E*��� [�B4��r�B�( RX��-/�`� �q#_H�&K���-�#�̺�;mK�$V�N�ͩ{�a�h�YH]����=G�����`�roA`o �:ş�ǈ�!�Y I�����	��3�-�Zw��x�^K� �4�PD�G82X_D R��Y@��4�{`("�L�UyG�_�vև�VH��=�K�8Q;1� �/e�[\��Y30�l�F�HeF�:�mD��Z��w��4����R�^���н����Jʺ	o����[;��*�jܢ���U�_�(u� (|����ӗ�?0�P����������|��M�����(�Z<������}��/ܿԂ�Z�/Bh���\�^~��X�	6Q��!?���_�s��K�B-h]g̴	xp�q ��9�j��Ec\�pi�R$6k�� �Q�W0t]��Ϣ�NTxJ�@m�������(y�.���gK�8�vQ+��\W��z~dQ�_�e�)?dz)q���#�|*���P�U~Y�\c�{�y1���H��b8^F}�I|;���rx��Ն�@��	������p��w�E�N�T��kM�?��-�&?�$;��P1��2�	�N�� ���p`_&����+.�5 �ixh�V+�r	K(�/�v�o8I�P���-H��)���[���	�g�3��d{r�( 4���s��ۘ��x��0������~���E'����CH��-^P��1Q|:�5Ұ��Dv�V�O���*������|G�������R�y�>�A�]P�5=e�|0��J0�y��1,[(G �cj�×�H'!´J�L�-�X�u��9�_B ���|)�v&�w��׋?p���5�&q�u�cdy���@��_Qi�G�A9:n��T�1 t,�(�r˰A�kY1�]]�J:�W���vh%!̸�R"�/�a�X�G�A�h�+?��(�q�	S�j} N�Z��Ƽ]Af w� "���1@LC�0����n� S��E�o- 
�?$,c�9)�	�1���2�R"�����N�d���A^}{ h��1��l.�cqb��E�
��ehYU���D�`����A�o��B�ͼ@|%#�_�uR0�Ly4���k݌�&-�_��h�4� � S��k%p�@h�a�+�,��H� ,)��2�V`�B rI���\���P��'c��42~5���ɀݐ�	�o)��5�fz��;ji u��[4� ��R���-'��0�w��!�_��	��.ݲ4~Jj}�K�����1�K尝�IR�P$s T1�Z!�X��c�b��~�P��)b Y�頔_�;�i�{�G���~�R�Hd�?@����		��7 $�^R���JB0	�0A����0)��lI���(�����!FyHU�-�Q7%��m��;n�	�Uc��l飀裸h^/�{*�*��a~��!�����[����� _W�0��
����w}}�²�fH�LRh�)�6[z@�QW��;�^�?1~ ��Ix��� ���;�R��[�h����.�֜��8�w����~Z>˃vH�Ƀ����0^:i���-eo'k�H:5Ofy?�@�-ni�@���1Y�e)�Z`̋)'m|�&r�.wf�ܢ�q����	��;�@���5����E39,r$�CS��8�t�C������]!���E[�*є��`&�
�M+�0f�^B�A	�ҁ�`WTv��7�Y`�@)/���1�.�2@�w!L[��c ���s�n1N����FpW�_���V�9%6~:z��E��fKp�<�A�FQK������U/�,�NO`�� )���Zih$ri��O��}��O�t�%dWfȲu��N����M	��'2:QJ �Da�uK*�
�򄰈�O^U>��a9J/���cogE�A��%x[�ş�F�)ꮷg�������+��<eQ��'B�P��`z���.�W���R�mw��b)F�YCP��(�ĺ��+g��*oV��
�f�]�4O;pI�:��C���H�Ru���YQ[��)}ye���^ѳ]*��D���Q�|�/��U�:z �-vF��\�]m�o�D��]��!��'qaL�-L�D��PƿZu���iAz����0-�p��	��_�_�*UXx�[j��l9d�3\P��еX��!��g�D���X�E��C�1=�Fn�i����R�W���<��h�%���6��2�{L.�3f��4h=1�K�M��G�"5�~�aj�_	�bW��'�J9gC!ق�c�:A�q�i��0[]��'�n$��c@*��r�Z	���5Q!�����-����1�5;:4��Ұ_�����
��K���#���X���	�~��)]Y	������4��Z,q��"T�1����QgT^窀��Nc�z���;&0��<��|`V�;2']0V��+�e�	$w���>׀�5�$�X3��]���u[-�XL�
c)DY8���0�9H�|�/�Ec����Y������ һ�T�9��s"����N6��)������hbQ��Ї�l$�'!X��]��s���2�RB��v��K?|7/��vElb1�~����ծ^�Q��虩W�P��.f�"3 �� FhKO;[r��B`c��p�hɍ0��8��T��B��	]�<����(<{p]�M��J���n���?r}(���Xh�e]�q�5�n�� ����WTk����	3*�b�we�.W�5��r��	k@��[���r���ދ��1 ��h�6�[,]���!������\5����O�q�7���g�b=��E/6Q[*8V	av%��u-'1���"�X���ȷ,����!�'��ԏ��^  ;��^�o���ߝf��/>�
���w�Z��uq� ������E��M%�D}~V~+��E��!��\�8iJ�{�L��uڬ%T�n ���p$W8w�_5`h2[(2i�X�1�IP��s��)�}T��v�vl/�Q��m� 1��/��\WØ碥��=�S#.�}^�	ef�������XA5����<��ame�c���h�_] ���l�4��c~��^�e��e%St��%�}�Q���]��UT�R����ZLL��]�a���&~+B��v��LS}&��(�S'�ˈ��LaQ�kn��h�\MvZqB�f�4�� W)��Q`K�`6c^���I�9��P�o6F54Ms$��`�9� ;+d�%2Gr�UTPO�rc�,�R��������1����j)D�S\@nXW*p�^J�(�^�: �����&ы��il�围b�LoW���!*J��HE�&�-���	��H�PŅ��t��$��]�:��2$�J���V*�R:�����h�:FL54�C�_md�}/Q�n��u`V�5�F�*^�Č1е��O��1`dc(J�E@�N�Q��[�^�*��R�,XDsJ�q�`�n)�hQj���A�Y�٫4_�/4>#§�|r�hu���`���S	/����`GI�Nw�Z��!�fu"A�W�)_�X��d;J��Y�-�	�:(�&I W$s�1VJ���ɷ!^����[��_�.~�U���WӀ�ֿ�o�L�0'�wApN��i[]��@�"�J
������
�ި/�]�[����T].�0N�G�Jѵf����
H V�vM_c�� (	�t�i{*�s�2 V�9u� �y�I�l��� ��ofX�
 ���(w �1��;V�Ĩ\ro�j� aQ��mEa	O�Y�o�&Æ �hSm��Ug�w��o�]�۲�{�����4
U釽��>�.b���x�F�y��!d_��P�w�H����@����@-Μ�)8Xh%{��X�_<��MR�P&&]E0��2 &\�K(�����kP֕NK��.�Qc~.���O�D˸����b� ]R��1�}:�.�ل�ew�.y�	�R�i����2>.Pvi���0c�c�\�C�������R0��|f?�d��y�����5@��[��A� ?]+�ٷ����$~X1Y����jTr�,2�` ��|�i��ZQFؗ�M�#U2?���E!���uDT'��!������8�}�\�l} 0�(g Q��?�ݓ���PS�������oz������:�\����1��;�[h�Yf�/T��.U
)�!�㇉�� oE?�(��?=�臱NK��phf.Aʫ=�J�V`YN���9�K�&@@�/�Cq�@4`���Q�-�YD�(����zg�JR4�Fu�`����Ҿ�Ȣ����t�$K��0F(w�0�=hXR��]��X��T��f+�)�+�Q�C�u��N	�����[��P�q�R�mkr|�'�EU1w�T~�1<S���Է�N��V�i��F�,0OA�v�=�`)���xW没�\/��ր�+�/�t_?�P��/���Z?R#,]QX`��ᙠ�h�J$�UO�r��X��ֲT���?�m�oSBQ~��^�(�!z4�����T�Z����[!D����A�g��-)�>��S�t''O��1���w��_��p�ubzʺR���Q��&%ZM ���0C���O����ř_ۣ�OW�k@�Y:7_1o{P�@��J� j���C�1�RP è%	���>S�H�'T.�y�MBq�%�l��!
���/~݀ٺJ-��h�M#ws��%���/{� ayYNȫ�P�gNE�hq۳�@��IG	�]�,f�r��j������iH �~�.��t%�N]H=cy����X�Y�P�W�x��mUX�m���_cF�b4�fu��D�l���~�1�{��|��,�Ql��e���ҔDx�X���*��g%�Iu��� H�v�;�Os�-�	aYa�d�.��"��Y�R�T^?��N���i��n<�1�~)�j����2�����GcM�#��� ��O.a����tEр��A�Hw�*�g�M9�S��JV+���@�_f�1@�Gi&�0�[-�������`Y�7�Jl�d 1��s��F}4��cNB�<�Q��1n5
?�c�����=Π�I��H4�R-k��L� I��~d�@/R"V�&aS�-kA]��p<-���~�`��2	H�oL�����Ϩ� `��h����Ʊ>��w(]��߿�=��XF	K,�A��&��`�׳/�T��W�3E%dI���2B���@�ˀʽO�j��Xv�Y���CU��	�E� �x((|`h/)l�K@]hY�,%��g��� f_�P%��XUv8Yڕ�!J{���P�f�����\b�-3c��q1A���>�b[�p�/��зa��C]=�F�[�l\u~��;��+[Z��. �g�|^�j%~D'�7��V����#�|;2� Q�4>%Y�]-��?`eH_��^�����%���|GѺmQ	��t�s�[�˲"��	WOr��@R�b��ߢ��ҏ���hlaj�y@���?6Y���A��/���ʕc���09J,N���1Ӹ�@H�-a�h&6�4����]^�A�N]!���#�`����Ǵ�� �Q����IN�3��^�h|��W��R�'��Kq�V�k�@���mEpb2���H�"�x�e��s/�V��l�ؕ\q@FA8�9`�	�:�D�^X-^��� Y;�4@�.�K����b��h�P�����-] -,A<N�1^YW��(�&��"v�I)�U�R
O�c�V%@Y���<%LBr��2�����0(`3{�,��veK*���l��N�hU���q@��zb{���5�_���
V�0^�{�Y �ʀ2]Z�4�C��{PE�}A@j���ֲ�![ �Q���3Ň���p����>Vi3���&�/�? �� _$N)���\.�!V^8j���5 
m*:1�h�&,�V(7/tz/y�d��3�2� �n>'�]uؼJ�_��	g��(�������z1[|��8��[�~�k��a@>nF'gH0����	�x�-�]�l�b�We1�hkT��Y����f[�. -�=[�� �5(	�3!���6��}��Z�gz$�2��@a'�f�>�/�h��AD�_�Ʉz��@X/�6Q�_2��ybs*V>$Z��	4{ ���b��)�I	Yd�b�C�������`(z¦�-�,��w���������.NcuY�B�M�`�uZ�-0W�����Yߏ��3�+�U���	M�� �f~
�ll�A�u�$�k��U����U1�������W�[q.���\�ʈ�
ƾ�� 0SJBP��Z��y��R�ק\X���a�"-`������ ��L�z�-�V��9|��_t2P��`����A�$,-�	j�)�1H�骄�@�j���䃦�s��ʦBڎUl�'��}娥u e�h���_��P����� ���k��a���r��@��nG+?E���O�����+�`�h�e�Q�r��I��H'�dx��`�	)w�{��N�%�W���Y9A�1z<R�!���@���D����#)\ ¥�'�BC��.pjշ��	Vl�����*I�^i�fn����}��_�K�̲�@#;]Vh�^����%��n#\: �-�jS4���G�&���1ݗq�B�bW�z��M�`��V�K1��)��to R�Yi�K�.���t��7[��Z>s�`_��	&�^�}C~������	�0���Z����)E������`�ZS��r^�#-o����3�01d��,Y���	.�1t5 �T6�9- G�/�!ݟ~A�V����֐K�a,Fm��J����[��ߔ��'� �[�`qx�� g��܅AJ~��uO�& �^8�A�]@z�������х���qA�'Y�n��P\.!я�W���uZ2�hl���y_��w���ꎺ���lcj`�
0��9�WV$�aN�"���1��A@KhxL�X/��_��ĺkj�,�ru]x�v�4�Rheg�X_L(���-1�vZ/}4�'!�+�§ &�NQa�o�=�q@��>�aH?8��e�u� �_�`U��5�V	�]��� �*�i�@���/��aH�l��ۋ7�Gn��
"	5u�:�'e�]l��=^�&�9I�KR���
3�	���%�<8/���>_Q���p/�G���-����E���k��(�	c��M>P(	���2fX��H�1ؕ] �~<?[�<B�a��q%��k{`�\�*�st}T�ߪ�������,��S��GRKP���\��n~4N!먨���?/�Fw�����+~��%	�P�LA���/�dS����h/bet�h�<�#��
{}=	�޹�̀!!Kڼj��������g�1��`�?i�	��}o��q�' �R7�Q����"���>o���J_��^�1�á(@�QPT�F�mN	��` �	���0�.�p�R�N��R1Xu�=pw�n5x���$�!�̼LU� �x�t����,������0�-0@�W��Ϻ�)�:�Sh/y4e��A����(I�t�p&钉��}��Xl2{�^�*��@U��6S�ބ� ��\�e�t�A�h:�0��
���	G�ғD_��W ��HQ+`U~zxS���P�v1� �E`u��AO�_��Aj�=?���[QXm5���;����z���E�`}���fָ[����щ�>��! ��jl�)�f�����R��&�l����^��U��U1鑟�c��x����b7��@� �R<���)�_�]��p7��Y�7���\�(��\��h8�W��_�6~, xr��gPB�v=�� !�P��$JS�7J�Q�K��0 �di-TV%]a�B[�	/]F�[@ r�
� J���)!T�
����� l��%������p�� �9�0�S���sh�$,��'^$c�Z}HT=�	l�p�Uz�)'X��	����z+�".���֕1���*���/(����n �������  '3�����>�rb�uy�*�u [F� ��9(J6��`?���*!�)$/��Ϳ`��B{5���"���B�+1����+Ĳ̀\�t`��|:�	��hq��'RJ~ޠ'�)�0�|���>�D`����!'�=����	A(�[�hr�%^]�~��U�V)p-�SH.45�� �rq]d��u�){f��(ou|�ʩn}B KD�Q�AT@%-�LwHu)�G� ��\�btJ:��s�x��-eBU@�VnE�׬��vi���I&rk��5�-�ʧ�	�Ib|�Io�u��o�e�}�g�`\e�]^��x�%e�"�U��WMe�@�Y�\�G�S�Y���-�ă<�E�Hv�9%>��[�Xˮv� �)vE�!��&�p��o�&`o806^f0Hh�/�^�B�̿[C�˩�.t�pV�	�Txqp�����A
�R$�!�]/ @OUt�iQ�;���}"H'E��t�l&v)<Ne	����V30x=^k5�_C���d}@�h6��[j13)�p�Z�����q�h�l�67G�	S/T�k�Y"N^���I1I��y1�&����ڕQ�r���ӯ"�h@��H��p`�\�c�W�y��k�z_)�.�2$X��5��UM=�Ə������>'���X&��c!�6�H����,����Is8T`A7��oP�A����g����;�Yʝ���	��Tv���l����*��w/ZS��	�]���z7l�GwqS��B=%�hu4@Cx�m	��'jB��X.c���������=�-�ҫ�ǵ,������p��Ƴ	Kv�q2O�@��χ�,®:X��m,�K��Z�险.��:
J��&@�)�����(:	sF��$"]����؎�� �1븭4/j�Ҏ(����io9<)Ǹ�"�� �h�0Ii]�91QYmd��e�I/߹5:�en������0>sB[!ȷ���fZ�VW��w	�[%e������&������X?q���e>B�KyX�kCW����|4�"���L�	�T֏����b��L�Xe���A�(�� V+���=x��E�c]��6k�ԐK��f�b`^�1Q0?�����*	�1Ui��k�|P"�-�e�C���yZ�;��[p��ѽ$tQ��E�[=_�&�-	)�V#SG�l�PAI���11}/�������;�<�X'!W��,	�M�h�Mv�]�)�,�h-�R�������wXX(#5W0B�=��_h�߸��T-�W�(ܨ�;,���N  �[�hrk�(�F[��'���8�����[�
�B�[$[ʠ)��I%�/��Nt���z<�4�[^��'�7�1�����5��8Am=�.�(p�~1�� fS���Ϯ�QE����,I�AU./��&G�`��=�^��R��(��i�p]����s��i�Iv��a��I���*�eq�H�>Ëogx0�@1��'_Q0�BqcS�MyN��@�cI6�q,z��v�Y	L�܀�5։�/1ڌ���zg,�NX� �u�P�2�3.Vcqg?�w �?�M�	�`-�F�b��x'2�y'�`%ln (��yH�����0�Z顷B����@�{G%��u�_K.������9P�v��?Q�˯a� ��6�-�d��c
J��M��Q~��Z{�E����4@�5�Qp�go_-��9M$��nf��������S��'0�62�`d�]����b����d��`/u�]�GL	��m�)� �;��Gns�������-��3��@�_(�(�o8�_�X�2^W	��NHBX�����)�PX	qs�EF�h����� �ؠZ�P�q�WAi(-���ܽE#�� np�Ɇ�f�K������@�]���	�)����OC�7�&]MpL��Z���@/�'q����֗eY�|�L����Ac�#�����/����cz�`|�|V	�U�"\�8����M�G~Z�Sv��<�oQ��'X����M�53��5�XZPU���?=�	T+�mH���),g	ht�G �X鷪�ID?]4I�0uy�Ϫ���|�@5�*�>��-�T[P�(�i�"q�H�"1ȃ�L��J35�%[u��
�>� ��)���3�V	]Z�f Î�*-���1�h8=�����3@ 1��s��H�����*����)��0l��[��uL��N)~��J�m`��PCS�	X��&��Ij�a���s!k(LB@�1[��{P��r/X�^;�ׅqG������G4mT%Wy�>�[�v��8���/ۄt&�
*�E�%�b	
�;qp��� hx�g[�4��o����<�`N�	)Ue^�3�-�JƍjCC��>Y�:*	PގYQs
��P½�8Fp�����
��)4b(���N��4�.� �ag*��(XRYӾ�7�3,� �5�a�~0�"���W ��QJ?���('�Z�NȌ ��@KJ��� �1R�t-5"%�[T�%LW�Ek/L)F	��m��"% �&4۵@1�kQw�k�*;�"	\ubj�_I��5���45��Xϡ�w�W P�x2)���f���f[*	�9&��:�O��A���>QO7�q�`���v�IOۀ�ÿMe�\�� ��ҵ���{�=�����8
�0H�c�լ���x�Bv|�6����p8�C}J��Q�-$��Y�	��#��Y��R�Sb�ž<#�ظ4�_�J�I�qN�Ɗ����I�HG%�h�R9/����|ÐN[��l�^�T��]'��	�/ R_��p&c:K2v���C�MmAօ	N1� Cn"\��)	hO,���{�<�hYfТG�]1:ч�5�
�X�^����dE��A�0�V��'�mg�����g�8�ԫ)�Y�`��	h{l\�fQ�����X�����n�ѽ����l�PRL�V�C�o46~V؝/�hm8�B�ⷩ�yA@f�ٗ��mh�9���B�с�_���hw,LUS�z��i���u����|�ѧ�"�g�8tO���K�&����q�ؼ%����g�ZaZ*�UU�"?a@^xE}d �:zL1�[�H�y���|���G�(h�E�	!�[ݪ�	��՘�Pd�P�0j��)�-�I_Gh�QJn�[�ո� 3'^��%�h>5�1F^b�UX�ߤ`'�6��f��ri�8��fR�??X�����#w��JX� �(U��'Q��5�y�|��8ϺF9�G*JW�)���:�%��-�5x�e4����0��}Z�r�!h<j�_|�T\��x���"�3�1vBbU���Ez-��k%�3vdZq&@Q��&_]���٢���'�`�S� � v�����ԉ�^`]1p(�x�|=�J�AC!��)���� �z��� R�u�0<_��0�}(2)� 1�%��`o�Xt0LYh �zR�۴ �BruxjE5�'sۗ�� ⸝	�I�8�1����Ƶ���_�| �5���<�� 방��,���4�;�0ЬV<Q�V1;C ض�*���%n�/�{�f�O~��3�eP*}�Ky��I��d�%hTg�yY���0Q�%> 	1�s�~�U���8�#��G�=-�}�\8�3�h�#"bX �@���4���Zp���N/��P6���.�7�0,eb1Y$t��;��B%К�Oc<H	v�.'Xֲ��/xw �a�L��e�!� F����� �^�]1˽�ud�w{R�����`$/�OP�"��
w�v����f+6K�?6�A%+�[����J�/W�OqJ*Y��M]�qÕ21(U�|�])���Ch�e��m8\n��3$��|b �LX:�ՎFxv��W���yL/�0� H����xO��X��y�{]\�@8��10���HX�@$P!X5�O8�T�k�t��9�,�X�k8h.�e]���l�%�~��>K�.���Y,�S�:���L����QIdB�NFx�D��k�����@�l).P�'� @ 8;m�N�*1ȹ9w~��P��w��G/xʼa���H[q��!�C���C
�S� oVh�AI^���O���醏���`r��)S��و���_`�ډ�s�M^����8�,7n(I����2XZ�h�9���qa�>b}��j������װC�p��j��49 CX%I@ �e-Q�~ω\�K���sz �kW�f��'�``:�Qj;l��w���	<�5�as� �U�剢��
��s{�&�	��@�4[�>�!94���u���0u�:� .�ɤI�F�:�dva��E�U�����'1-v�@󿭢Yshm��'B�hf�/;�;$�.S�����BDA.�>�����y&�Sim����~#��N��/~�P��1��"oL9v�!ڣK+ǐ-�M�P�5�qK�����r��v���%���NϽ�>��Ő0	no%Uxm:��vP|��(p<��h�տ�����u�A2t������{�ñ1�;�Oj��Y����4�����fJ]���U�SЄ����/J�p�ϖ�!�hbw$�Y�X$��'���F����YiK��z��:\BL\��wi�U��A�D'7�����K�O�?<����i�6���Lڋ���I|Ę���?3� �i�e����q��_֏Zx�	��s^Xh� ��a�b�W�E�']0M�LH�_�e����i%}�#��L)͕��@�V:bh�[h�/04Ac;����@O�>�sLC	3�r�@'^!=1�vDz�30o ��>@f	�b� �[�^Q�������P��B��F�x&��	��@Qe�(ڟ�ߘ�ڔ�Bwƾ���|P��Z~�)��7]fR��	z��j= ��m�?��G��1�R� ��!u%>u#Z�w���ؓ����|��#z����<!�f�ԙ�[�]t�A����\hJi(��,�U[����{: ����m��饕���K1�_q=?����80p�t�ry��Z�,�v۲z�W���S��L�	�CE�1����nh^��{�*�'`�ߦ�s��BS�	/����H=RO�t^��ȫ���Qa 4� �p-tI�a�}/̉��i_)ɀc���m�@���^R����ʿ���S���3��1��n�����P�����$_%m{��u0z �P]1J����AK�x���$ �3Lnƹ�9�׬v �1pJv��(�ۊˏ�Gh�\L쳱�o���e��)`H�'%u���4�\I�R��6�N�x�ꊤ:˭�����|��X��Dk��X��4�6������`���N-9KH���TG��Ȱ�Y�S �xk!	�@&� �p�@��N��[a��iV��;��i��tA���K�8-B���@�#�Vv��|�	^���� ${;��E�	��`Y�N}o]X�`�] �0�-��>a�j�+c�IM�T@���H	�/�d��
�V���(Y��<�]���/H�����)u�(�������"_v�:�h�n��� ���	�����[��Z�N�Ս!^�~jHk�X� G���^V���#S�_T(T41�������kU7�0�B@�0P^_��0p��f&���1B�")�5�XЫ��'�i�S�G_t��&Xb��!��Wh#0J��e�J>���L�%|�ȓޫ�e�����5���so*��7r nL�ډ`�lv�c	.N��~��Q|�?ǚcIR�Q[80`�~2J^�<��Eh%�q��QE�AF�i�ԃ!g����(s���@]Ĳ�opX��C@'�hE�<긐��Q���ǵ�҈9��h]f�EX|R��V���T�����XiX@�w5�\[<�!^i�P�^@�[�K����[!t�Jb>,!�qz�h�`�1*�� ��LG-��V'����i��Ws�~r��j�h�v|�dp!'�U��-�rh_!�q���^�3��F^����s�!�LH[Z��(d,��Ki7�X�<z���lQN���.��W��!�h�hG �4@l:�%����1w�$��4��m;ľ+'Kʦ �B9h'�Zx|O���_jA���S0y��	�[HD ��w�; �#x�F%�{�B a-ws0�D�t j��`�𐞗����˕�ϷZ�)�X���8E��O��c�[�B���0�'�� F�(�a�� �P-����8
`Chci�Z�
Bo�a<�;��9�@W+ ��'���V�r"�L��	>&!誜�ޕB����W�2���PW�	��DdO^��P�Y�?S�չv�ĕ�9-��~ ��\�S���7�j�ˉ�R��9�4�(�������6N3��G�ͫ�L@��(]����M*��*Ǉ^��Ǹ�)����}f��yLb3-Z���/��R��`2+��O9P��^��o��]��z�f�"�TKT�Y�i;Ř�U� .lV)�]!�VBy�9U(�%q����/�uA��˜k���J�� ��TƑ��O����I	�Z���ն��tB�c!y���G\��>ŝ1��=�
4/�o�hI0�����N�Y��Q<u����[�)���&u�8�
�k�Yh
������h�t���P��s���V���:P!�17G/;j�W��{�w�*�E� �+�d^��d�3��+v�w� �P��8m'qAH��p(?�{9el�8Bć��1����C=)	x(2�ķ�x�:{���R�X��0����D�� b���7Fu&1���z�z�C!���*��溞�Xgీ��Z�EОC�&vM�0���{>���y��=�6Fg-@!yi���y�A3B�nsT���B�f����o��j��<-�*���u���N��$��őR�
��� �EP�*U�X�_�d�y=0��Q�Tq�.�����@dOO�YaTn�ǖL�,���u�@ؖ{q����tງN����I&a����@���y���.���Yݤ�cI���o
�h��z�wl� �[�����~5Wt��h/X�[
Q��o�U]��|��"��
,E(��K�H����Iؐ�0�	��X�LX#z����j��0?�Y0 <͜
��K��/S��h�^�-�{��4��Q7�*���+�k� �K�_{�+�X���x|Du�L8�d�|��[B�����6�1�	�9	��擱y��B�m
ʀ���a1JѮ��[Å��X*��H��p	�5 ��CG�`+.A}�V�D�,�ˮ8$>���=�W)����K��b'Ls�ʉ�Z�H�g:�j���.�A�}i/��:'Q����O�c9����똁i�p��HG�?���x�҃�1��[�w?���F�U� w�Nw�E�-{�޽�T���';8���K q�J$0x� ��w"	H�}�(8 ���YX+���?�������Y��;\,��|)N�H�&E���h���� �ө�1�)t���-v��w�\�Wɴ*��S��P:�N��J6*dS� �c=M������V�O�b�]�D�q`�s\%���X`��o�(�nfY���(,9~*��t�oP'���88�0������
�`��'(�h>t'\�rwni��h��n��ǫ/g���堋��Z!sЖ�f�R��[�����b�_)B�@�K�X�w�AjλT0z�K� ;Z}D阒�e��&�+iE<-�U`�Jn�rT�qL��	F#�(�^��qn`�.ZY�:�1�t�������h�/H�G���� �~�4��1%���l����.�SY���fץ��ɪ�x��2Y
S���bi+���1B�h��ŲX��#��a-�"��P�����^�������|V/��ߚ6wQ�Ph�z�M`���`�f[ �	Z�h���u�'��5���C�4g����r�����]h�X�_v	��I�����׀,��}�X�rFo+	̀��V�(��h�A�Iz��%a�P�5��
��HDB\{��@�	3邓#���1���0e
�!j}�Z���[cw�-� ��靷J�����Tx�!���0��uQ���?�у)�Pd[�SU�G;��������_�0\zZrhT�27WwZ���O_���%�����B�pI.X�p�ٴ�	@E^�� )���X�Q`�2��hW�Q�b���x<	{)_q֧о�6��`4#r-�d��A���n�(P���߉�
����|�x�����Z%5Wl���v^��ziA��$��CHS[�y4�|fh}������K$��B_~WO�<D�G9�0j���@���S01�}� ����'*˷h4)����X3*�z��cj�I	�}_���mC�_��0Sۚ��Rn�5$��6�	�v���	�~�`C�r'/܂:��VB�g"��K����/d���HN.%�	2L@��#��N.�ĝ��K0A��c�!�w� �Z_��,Xz"k�؁ ��Z��3Mi���#���S{VWCK�^��U`��m���)ڀ�1t���ux͇�������+�L��B[U�LiW�Lk�W��W�i���ˀ�@2��`������w��+�8 ���r��Ĵ9���yo�u�\���t'�.�Z`@���xE��[P�����H��@-�b��mͽH.�e:�j���3�1��+��hf �c[�M�W�馢��UY�LU���ݐ���e������J������[!��	F���k�V����]�����^�?gh6��c3�}�1?��u�[Z��;s���:���y �4w�sjl
)�-']��n�,�e���h��p3(���Y��kH���!JkΟP��U(�h�� ���M�?ʓ�Un5G�O����6����']YVT�h��;�	~gU ���D�y\�z��k$|�`�k�cP)����R)�p��Dqp�D��%�B����8�q.#B�c��w��c;�=�|@Th�Q�Y~^�ǡ�[~����K��l����T����	Q��_�Y�x�ڽ�$$e� n�;��ftY�(G��	�#�� ��x@�@��v>����r���#�&�"J)�ݷ,��	U]q�� ������F�BX��f��8@��������~zQ��Bq]}z�jSY	�]Z��a�-���ٗ��}mI`�#���֤�����f[��hR/�T�4]09Jà��%fZ_�v�=������ Z��[����O��q���$���Yh9��;�R�`�1*Z����'�T�@��c;��àN�# �vd;*1�	]�	lhX3��qzb�2U�8��x�"��B$qf��	ɸdP���X�P&�4	h\��L_�Q���ZB}~��G5B�4W��0:m�p()ɢ,\�l7��R�ba0����ω�p���JI���cP�8�#�h���*�Xj�Z�f�ꘉ� ���:�L� !]�K�z0�+�v�H)�/]��e��ΈQS�C��.����K����R��h�J1���@8�.L`U(8���#�]r��n�)J�l%�!Y�>���i#]L%|��G�H+�%4������`W��tD�0{���)���$����t$������~��d*�7��+�z�	P^��)��-c�uB� �_���o�IM��Å�U^,�*;H]cK��nHL
N��
G_.��-YI�o�鄃�0������I�M~�]� mR��W� i�y�a���А�^B���V�j��j�v��0'��i�X��% 1�-�.;�h���' Т��9�f[�7>��1 ��4�G�l�xu8��P�%�\,��y�OO#X%E-�MW�e[���m��\2P:d	��:$�T	�d �h�A�+)�+ď���P�߀�@-Cj��q�hQp��![�0�rE Sh/�eiY�&�@���WZh�{���`PV�g�j��1����$�������ˉ�qd�6�샀�OXoz�rx!@(`s�,�/8�K��X8C|���ʾ�M2�V����(�,9�+E04����:z�8w�	�VZR�(��� �pR��(�Z-����&E�:�԰@��a�[��W�B��^��ɬQ*�4w����_����;����t��d%�_MU�7�!~�����?�BT}U���,�_���hf_j�c8O���P�S}����1�/R�qx,���� �}��b���;gW�s�`ΨT�%o��t��{N"XhK�������He�zkw$���I�sqk�Ⱦ�K�?��)蚽=K{��<;M%sa=�6j�hi	E��g�b��"J<�� ��@�H� �U�t�+�)�!��+�BB?�xS`��T�cP��L��ʘV|�@�خ �'_c	�[�
M�)9-���'1������C`D�]W��_`�J��瀠>�3����� ?H@���8��!�ho�)��)�ا-��!`"KY`�rJ�h=�+,&��k��_$��
�Gn���@4��Z�� ʟl���-���4^yJ�A��Y��0�p�Sn�Q�*bC�61b���~QK^X� ��=hT��n/��_p��
�l�N�����0Ro�C�:�M�<[�`�;z_Z3(U�=����sź8N[�У%�b|a S.�����A��[U��?���iK�\"y0��,$�7�U�	I)U4q����j�'���Kl��01��w*���z� ?H��hZ^Ic�Ą�������G�'����hq��@�y��e;>�d��0��B8U&��4 �����)�[�x(	A}�6��5"^�Sw{hm��Za8��&�P ��p�%�R�=�lm}��,Y9X�	TVUSa���**"���t�j��K�t4^��������_vB-zT�-�$�Bn*I2���yHK��ei!��E�̪���ς�@-�a��,�D��	��ߠ�[�K��`�H�%.U��ROZ�i1
����	]\YW��
t/�����p~\~�/��7����ꌿo�֘�R���k$?����ax�0�Y�bZh���i��[A�K��7�B�W��&�J?��Ph�kGS[���=�Y�D2Bh�(�*a�~h͉����%LX"x	o.�O� }��dM辬�~5�`�2P,wd~�/���E��!x��:;Q����/)�TU`�� HrQ �w�k錇_���(��L���`F@���Q�so/�g�[�bYfZ�	EIdf���鰘Z��}���\E�.� 3m1+�IJ ��IWs�k~饛@:���d�~D��w5��%h�՚i��`J�<a9�Tz?�_��U ֐�%4�"_�vb�r!�so���h~��Z��
�0׈�((��P�y��N��X�|���,ޚB��@��c2L5�iy[H��&:�g��/RZ��nH��r	���	5������[5��KӰ�)R��T{6���@��U�b�'�юSZ4J}lԀ��W�z5�%�B�_�6T������h�A{���^k������[g�tKd~��FM�����Z�U�9�@���Q���I(!,0��`'�=L���&!���>x��{h'OCN ^�u�"3@�U��c�fͧ�G��j �.�B��s�52�G$��$<��'f�f,ZKP�� �9_q1U[�s4�o��D#c��2���n����5�X���/k�����>��s�^W�n�n�}v��]1�-h�r�.�M~�% &NF3�PT	�ϝ_�����]ne�Not
'[�+>f)=�y^�*��x�;�I��|�%Tົ;�h�]1_��pn(XQ�}�+�/v/�3�k��T]���A��3p��;W��dX �|�1��0�JD�<���Pȹ-
_�S�%T��>m_���/��k���Bj=���6l)sڨ:��v	g�F�
���"�~�{�!|�U{���!C/�Ѯc+�����?R���޾��8Sh9�%vY���B+�]YM�.�g�����u�NXx���$y�O�@>Z��T���(:?�|�{�'�����g�]A�5�|(�f[���R�8�n�pp��[-Y����"'h�a����Qt�p�(�s)�d4�K���Z�`��b�B!�W���H-2A'�u{> ��~@W颼���U���g�h"~y�$O�8�~�	�h����XRI_���]p�:Ś��w�%"���ż.��]��.��]�
�#$�/c���>/�^Gp���^I��Q����J��%��z$���5�z�/�s��rQ�~�YG�:��^��42xd6��@=�D�`|���-*�z��ʖ+�Ѣ[�� S��P�h龯����	
;�Y�� ��3�\x1GD@#��`F���OBLE�%�U��a'zVрX���P|�a�IA�9=f+)Ȅ��u�D��[�Nf�p_'�u\���p5�Y�;W��@q)������g�@ ����^ObR��&�\���#Ć�j�hwJu��0�EֹZ^{֕_���-�N�g�Q��~����/h��$�]�A%�Db@��z,� w��K��[T[������/��b��kY/���+.ABM�)����'�^��j���X��0�[�F���P��h\5j.��b,��)��42�"~¥��-ݠ��@
ZP����@�`�[t������ xg�j��+B<��%����z��{@�[fP�j��0�� �w�iy�Ƀb����!��Z��1��@���p���+������U.�4����܋ԇ� _ ��?�1��ڈ���A�ս��Iֆ-�,z�szq���B�u���(K��\6���`_{���N�-�|X��Q��<q=����5	s��<���(e���U�K�&�|à������`H-]fuI�\/����/�s�c�����%{�(�԰�����݃�ZK V5�s%fh'o8U!# �"5^�4��[�A	���.Q���B�=��/�502/�_[�!$A@��W-�M����\�\(�'�`N�yK��D���S6 ��J\���m;��z����{c�C��!�
�>�r;���!���>��jmC��`D���m:&��cf	_<W"�zGHXUw%	�� bP]�=kߌz�1O���A9�N�*{1h�����&-_lV�v6�郫��0�3�
X�o$P����y���X�h���	5��4�> ��(-	w{�x~y �|�pR�^�4�VG�t�o8�T^��-�*�����3�lR�`��$��b�^`��?h;S�y�s.�,�E�*�x|%u'↟O����	/�P\�@[Q��y_O��V���h�h~K[)�R�������Bd,�������$��M��)��$�����<�-��U'��[�����f�6�su���C(����W����^�e��_
[) Ny7�n`K�����w�6()ڠ���[���ܥ�Z��b�`�'��`���ZIW�]��eF���<���_�ů���K.&b%^�H	�WeA�j!$�
NZ���Uh�u c|���^��4PT��Qj�=����(i��۪�5�� �(�&�!�Zѷ�E�꜆�i�Z�%fKZ
�]|�3?�:�ax����ޠ�`��F�)@!d����-^q�dLSyr�RT�bK� ��"d-Qr�^�ChT���%�_�y ���w0ǵꢽM���HZ(��f;�%��p\�t)T�#$B����N�O :T8�x~�{)��z�ƶ� �Q�gqM�0F1��S���v���T6a��=�rz��E���B�t ��)���HhF-E4!
���0t�X)!�z��/���@�}-�V$����� G�K;�O���Po]%�X�����?����0�zF�^C�|K��D��-�1�E@�>m	|�H	�w�+RYB��o7`�9J��r�Oӫ��Tk�@�ix"�����-(j*�Y`1C��o�XtW�T|_/��93-&i�����Z<�0�_�@�ᮕt5/�{-�|jA��/�*�Ё�wZ��y�<�<G�}��sF8l\�� ��a���0� �9��PD�1w,���o�d�*�`��>>�?��h�*ɀ#�xL�E/u�G��4��3zy�T/�?��|�Cz�/Y��!�x��k5��_N^��1#:�W�gc��H%`jV�I'1�|�i|x����4�/����*~@��BjW$g��k�]��L\�@�2[�4�l|���Jj�8��^�	ܷ�PI ��+�)��� �F!���Boi��%�X�]��w 4�����R��!C�����`bR�\٢�[^��=�,H�����	����h�K�wﰎe�s���������� �50F�l)����l�����W���܎,T{V�07��4=��,h��:��XI��]�h���S�-lڽ�g
ھa��^���k�Gc��D{�e8Z�|�����`� �(2E�t��BS�X>��`$�
3[P�%��a�#�	�}�)tPz&��kgY	��6�A��-X� ��?k�OM���z�H�� {!��i:����X��F���N�9�j��:�^�	��wA����l����^L��]�n�kTxS�p��mJ�e���p9C �L�m��[�[���O���Oh�]E`��/��� �xFy�`	a�|R_f'�&	lThɌXJ�k�^0�B������8|�
�b�cZ�11ڴK�������}�: �f�x&�� 	O0�4�����3iT\�O��Zh�>/�����e�%�P�H	A���V]W�N�sJ��I�p�(3���mY�ΠNi ��f�XqX�w�iZ[��P�`k,�`0Xh	�1f:���ňeA)h+x7 @*���\^��O�< �k�rM��O��, ���i�2_����C�(��� ǧC�/h&�IT�K�	հ�T[�v��Uj��E
��P�氉S �0TB�ԫP��Ә��=}�������Ƣ�j��Z�$W�%]`��Z��g�*?-�w]}���B��F��6Q��#d�n):�*\Z� Z���R鍗U��(�`��d��N���	g.�}{��?��t�U���t�I�߼{if\w�TI�8@�v|NPB�*,8�Rʚ���>��TZ���B�����4U�'������b�	%�ł׆ݱ��4BQO�
����Q���ҫ�1O�5V��T��e'/^�,�(�4oUC��?s�R(ʢHA9�>$���"& �_D�'�H�6N�S�Q�}�H�MD��7����8��p
�����o��
f�v�x_%��(�~^�h�J3���Z��9��h5�9dQ@%f	V�>���R�8.1#Nɞ�z�^u��B��q ��@���l&�C�� \�)QO���>pO)�C��%[�h@�%Z��Y6����$�^R@��U/o1޵Xh��l����_��2���ũ������,RGv� L!�N0�/��S��92:w�vpp�sX8? ��qh1߸kH�'/�R5U%Y�w�@ϐ���Ĥ��ݸ�-&�i%|���IqS�pN�����|�Tf��>P-���:��°���C��b���(V����0l]['SQ_A��Iu��Y����=5�^��`�P[j�E\>����!@`۰�0�F�7�ܲ�sL�[J��׬�����Jl�/���<ch�u��Q��r�I]鱒<!�ʲ\�^���	;�����i�+�^h}	�p�z��MLB$�҄�q m�s-�	@�rd����{��z���1� E��6�c�
�.e���t�x��U��]���3zX�n�.��P9(�ʶ�YB}X��@ �b�	m���� ��Հ�r�l_1 tYh�E��*�-�8l��2�%�w�(ч1{j��Tg���	����C]X��3��y3nST�=�/��P�w}d� 	����!^�V 	�u���OI�!��M�����(��f�i�SM��/�/�)��:$�Zo�B��lZup�O[�H�a�f���'^b=_�2��,\~��0	�2P-$G��a�!2j���q{��	�T\�� �6d�k/�k�!�k�-�v�-�0�!���[i������
T|�x�[O�_�W�[��$�-V�B�_D a�A��-0o��A�#�W��u.@�56<:�v��gl	�87���=V PQ�b"���cVՠ�n�E&)L�h���ǐ!�a��� u�$2&��雺:�v�2����ڰ�@/V|l4�Ȫtòb	h�Z����&�/���{�-	*v%@07b�+�}~-S)� ���=9�������	�¸��VI�?@�Ho�P���D��Ty��+�[j�,w�؈y��Y�~�������c6X!������ �}^��V�'I|M@]��a8��U���(��:�)-�]Tb��!�5:�kv�����1�]�=Pޫ0w�'�v�w@ O��E^�� 4;��fdb��,&�		6�upU��;��K,|:P��AN3���N˱�pb�*�PKJ���jRM�AW�_U\^H
�X��]Q�~q�k!�˞�b�-���-�Z�����w�O&{$G
+��I�����@���{���wQ�I��1�U1���1���,e(�RS.��*Bz�v�<Kt�$?
�˱&��M	=w�`�h�< ��L/u��-%Y��~�p��i/X���`h2׻TN*9/m68-[�0x�E�J`���x�����G�Q�/%^��!�&)�RY�P���������)�P��[��?��X%k8��f/�?���MW���y!=>K�����(��H&IZAhZ �1 � �Y��R�	���܂�Z^L4N�Lp��h�f�\�L�J
�������/��dPy@X �v4���L@�0����M��B>�(��xSK���sؕX�`��nG8��D*j#`�h�./��1�IA�U�dP��)N��¬Za�M�$2 N�/��,�Ӈ�����	����J�!�~�Ph�N*̉yP��"M�1?�z��-X���7��DAU��7�ݩ�w��a�*�d>�-@�1_��R[�eWT�.?W�I�i�
 ?Oe;5b;�	������z���i}T_�+��U�� ��L�+Tz�����]��0��2�<oN1�YP��M��Q-�|)�;�aOݲ�_�+M ��	tSc����H)�I���� �r�OWZj�����$Sn$�M� [`N�)]��
�\ع�B�.��8�,����U��y�������>�����Aq����(�0��� [¢�=�O?�T���@��	���XO O ��C\q��Ut���kO���-()w�WB�1�J�_쨞{?�5�9B�[��r�� �0�F�-�q%/
~�@�i0�S��c;�:����C�s�� �_����"�(�ۊѧ^�@��vkZ�r�eH;'�_�C�e����l����p �y�ck��(a�^��Wx/��!N¦v^�!V͹v^�C�A��� '��!�Pq�_��� ��ۭ�ѕ���Y��W���/�.hO- 4�5�|\� Sw��P��D��o���~$	����=�|#�3Z،�z�f���,G'�Y��@Y��(}|z���ShN�^"3)�T<Y4�n��� &���C��}[=n��Z-K#�L� �	1��NǨ�c�OR����i)S���.Vi��Z*ΔtOF��:�|-D�	��W�YJ��!�ʏ�ɲ~��.T���mkO?��[���1�z���F���?�s�':���,U�-�x��j)�ˊ[�!��F6A��*�`뻵voKb�%{+���
C�����V\`�$m �ёc�O
h{�`Y�M�ώ\��r�v��/C�_i>(����kh��1m�4/龋R}F��9�<�=��L9�tf�_W�xd�zi���U��,=RQgi�@�*:8P� SE��K��e�$�! ��7�%��!�X����~�����%���ҘĞ��u�F�m�8!́>�w0rf@���)�x`^0��s����<��q�`S~��^n��/a@�%(c �t-b]�`H	�zT�9+�J�Vȗb\���HH��tǻvr�V�F�$�-TmJ45S��~�K<��U�A�1|y:�<�g,�|��I�ws�I���@�&a.)eT=��@�3���=��o���T�^3Bm�e�<C0ՠ�"�-m@�*�����X�>��,���)�ۡ(~�h�d�Z�u��3(��^������r`2��Z����/	�3Q�/ڑC
%��������R��)�K?c`-�f��|�������~<�B7�����o}��U�Jp�Z�>;���U�R�*�]P��:�0f�*�M-�`แKvb��mp�������(�`Si&�\IV�����JT��k�}��=P�9} S�l��(1�[[���hK<�38�nD��N�����'m+���;����1@+5�B�MC����-��
~��+�)�+�����]�~R1"fhD)1-�`;DYa��	�����(��I}E~4����,�����z��>�eF!?+��/m <eH�	Z��5�����_���O5k�^Q+�Z~�o ��?�P�F�z�X(ӶR^˾0�@V� ��'����1����>�'w�;��1�Z��]�C����\��Z�(O�럃�6f.�b�
;�1��K��s�5=>�} �*W��FNG��b���N�E!�l��'��8`&��/DK��[������Y��T���OKKZn?0
e-�꺇f1n��I���N�kr+���g�O� �#5�b�B��L�1��)c ���:���^6��-n`���y�[�#$���^�Œ�����Z��2�+�h͈
P�%(�Ud�a+�8	��	|A��Z⒯�>_hO1=X�y˅'��w�v��G �ϰ-�2�zQ{�n0�s"��BP]ŵ���D��/�"0�^�G 	�J&���a3)#W�\G�KX�bt�[0Lt3<=X
y�	^D�Ph(To�X�h�N�fk���������-ŏ�?M�V>���#j8�<�����'�]�q�$"h�;jZ[�JAy���F$E�lb��o�����#X�h 
y0_��O�,ǈ?N�}5�)n��Ȼ�?\�;�,�o����+�:�l/� QE`�n[?�ȃ^�y-�պk)�ܔl�V��Z/�Ϙ<��F�'���@�G7�l��_��4=�>�r]5�@��(J�1V�$� �x;#�ϟyQIp�"A�W{[D��ث����=N�� )����K�м�,�-�<ZW�g�4�2*?W�ρ�{r2�u�q�7�i�}	@��Q
I^@Q���	�]� �;�0��FCNx��H�z�x�u�3	B�\����B� �Qh�6Hk�%������L̲*21�9=��W��K�˚�v~��N>��ژ�\(J�O����V�N�`
4xA��A�z�y	�鏢S[�$G����y�$g�_�F�
 )O���?H-	1��Wȣ��*{J'��E�\T�|� 3��)��q�B�΀�
=-i��V�%�P(	�.�0w ��{�#)L ���z��y�����S(Ӏ°R��!�%��/h>	҅���Ǵ|R,h�n ���ay)-�Zݑ�X�z�W�g�.��V	`&Po'KTt_�� �<9�t���a��c%�&'��B#|ǂ!��j��x[l�|�~-	�Iwyɪ��'�ц����|aA!�^A:��P��[�OM�~N	6��j��r�'U�����kހ&���������8��0��(7Q�
�Y��� �间_��ǩ�	UEtC�|�(��>��_�2�UU�]!J��@��'��;�.%')\�Br.Q���`(���'V|�^����;�WR�JM_ž���E���/�%8�`�!�f�
a ���]�wZ JE��XM�WFh�u2Ԯ�z/l9[X�l�!X�hF����(���slƋ]��QT?k�d�.�_Z1�k1W`/�Yqg}=wG������/QӥTC��ń����[�V J!��e��B�7R���\��*�/��o��) �l� X�}p��	D�Kc�[*�%�^O�)�1��Uv6~O �΀�lh�1}���wK���5�|:�g�M���`�T��&����?�U�,h*��K���)��	�U�ze�ۄ�ꀜ-@%т]���
0�B�Zh�Oi�2*��:�0b]"�郒�Ҽ���v�l�[x�cS�JsLf��-u��,��j����xj�Z��aƨ��êc-�����?�:@8�J�A/�ދ<�U����5I] �t|V�]&���H�� ��o1-�+�sQ\x�(r�L1u ^5F�_�Y���5�ׄNRǠ�d};n鲦;�(�2� 5��C#Z=�$9���i	��b
:F)�����(SP�����

A�-8�tNK�A��V�l{�s�X��������݉G�{}�8G�X	n��G�il~w��s��t0(�O(���n앹�ٲ�aձ(x:���$����Swqoû������9�i��� Zn�)\!�hy]��O|N�Tj��v���rJ��X*��zm�����8S�..�%��G4�x��}��5�X�]}��<�9R��`rq'@�?�VWn���r�_��|�6�a��G�=����UD�[Y��+nM����h�_����s�e���	w��^
H�3(��~:H{Z�K�^ C:@V ��P��2C����/#�����1úPZ�A�p+�&�d&$?����B0��P˷f�iW�[��Pk��c
�)���%V���bC�� �r�2�s�Š��	�TB��w=k1�tY��6�Pht0 �f <R��2�x�&��Mc��)�:�T;_�buZ~%��;*��@*h�[t��/�xͽY=`S�;I�?. ��
�$� �ٚUVa ���k���xN�o�o�z��m�#aXˬ[�#��J��꺏Xo-�ܹp�����0�θ�'����ހ���Yw`G�+�Zu�1��h-=~.�Q��>e-�m(%��� CRW��|q@��x�X5-�vP��q��(U���!N��V��5P,/���Ʉ>�@��v��{R6���0��sP1�_Þ�Dm~��J���:�f���pXW�k����o��z�忋>�r��q�FWY�fJ+�K1�x<O�JN�g@h0�{��6�y�]8�~f�� !ӸrQ �Jخ ����,1[�詵	;��0t-!��`�H�9�[��;����Z�Q�/�:ZuF:$*��/���/���!��^5�+ �>vY��~ z^S�)sOă�$�5Dlv`�6d]P��T,k7��X��S	��_ �57V=	�P�-	KfkG@Z��*�!�֏�1ǳ�-����t#�o���\5��UU�,�D�S�Q� y:Ho$^K,bE��?-���)Z�6g���<��?�v��<a�?C�JT����8 !�����V��>M<�@ԣB�+�(v+Hi���P���|�$>��z��akX�X�;�k�����6N����g�������Z����'^w��A3� [YJ�GMP�+l�,p�	Xſ��������B��!���<ˎx���%49T)F@Z�\@��o��k��|�7M:���@h�s_/D�� ,(���(32\>�}�|
�%FY���Q�	q<s|��^�cjU ����������W���vDu�-�  ���?�<0�/6|sVJP�;�S�EW��|OP��P�@1- 2*�o���(1�0��%�EuU�2��c�N�P�"d	G12E;��%��[0���\�8��S�\����(H������`lR}�j)���9�s����b�ԧ`��������>6~�91҉h��S����/Y��w�:N=�G���/	�u�6��j@_����ԭ%q`���q�[B�ua�E��e�<X�4�}�l��A%�DU�9CY��Q�n�	ɑˎo¹^w�]�́B��On&zA��$r����F�\i}I�%UO��}o$)��>�����Di�d�>pz0]�M_,x��逯jY�Oir��퀂��5��!��mZD���eLP�`|��1�I0��7�L@��M����@d�D�`>81w �©</^.�v@c�)L�}W��v[Tk���^���&	��y�SC�˰K0@�60}i��NU ^��e���ke|R�=��Ǳi�f�@��n�yػg�.�A��u�)�<��K-k�]�s��Z��B��,�]��0�vH��[�E���; 8gD]��:� q�F��)ˠ��c;%f�<����?%�@���8ñ# -7��[�IW��D�x)vA4��!���@��HO ��pAQ�wC9�8L>�b�����	F<!X]�H:�'�t}V�_�K�8�v�E��
�"!� �{�Q�G��x^P���3�eW ��1\p����Ҁ��ŋ��)��on��h &��_�q/�
~a�h�:���݀�] o��;��C�?��u��k0c��
IKڕ��T8��[9�);:�C�C]��ܠݵsڽ��^��Z8�g��qc-T_�Ӂ6B��^���;���{�+� ���c����T4� ��j�ǆ��d9f[�Gh1!������D�)^�n��0�M(��W{������K��Z�g�~ѣ���Y���*����Z>N�+��6uLA���4��hm�@_1�M�_����e-�[ܟض"h%�7�$�C'�J��Tj�TI����SQ��n��:<N�-�h��`���R�U�)���kl�	� X!"+p�zb��iPm�(&O � %�'4T�h�a?�-��Q�%L���%��'�_�:�|s\�hf�S���&vb��X)���^�`S��3HJ����-�m6!�W|S�H�,�w�.����E����;�VZhL)������Yղ�W^��T��SU?��<x�����X[Q��;I�U�?����*�9���WP�h�|>/wx>�>��z-@���m�?,)��"�YhM&_�i����u�v�'�W�ZB-U�:���	-���B;GR�YT������f��|.6z7�8�tUҲ ��^�}��OˑȀf�YEA1���'�SX�?��>���	��m���P�'�����F�yh�C�H�����up^�hl������h���\������p4u���V���� ��Z<_����!K	.}}�N�?�1N�ώH2�~6�]yPo�,�n�` '�^�)������fO1�?��m�a9z�^��%T	�p�DJ,
��&~��P*�8��[h,K���/��]�#oE�<���q��F��󛇑QZ�rҪ��x��k~�n��3��f�x!����Jh��FvMyV�$��ЕW:���S��y�P��Y�	ti��ux:�˲Y�� Rh;d�0]E4�`l���"� a������$�)� 6L��q隰_��8=|S���03���)�PFRNr-1!O�|��^d=���v:�P��@I�%x�R�̱�*&8�2P�ro~�vzS�lW�V��,{L^
�b�Z���2�J(�Bi!�XWQw[��� �I"k������u3��6�E@;�U��Q�%���x��X��7ܽ�$�v�HI��������p��z!����]a���V�B<�C}
��x[?+�_6z2��"�u0|���J���5��a�a�S���M���V>���~�s>��`��81n���W]_G�����A;��Q������5�y��V�"�'A��������_��	T�	�$(�]KE��������j���s	�WO���x�d��c\-h�ET|zʾ KR��[�?�<�#%�;\hf(��`0�(I1�����h��%�]�`F�)�x9�s��h���K�%U��F�Xt���8�ƴ�!׻I�P2�PFuN���{Z��c����KV�\�0�����2YѸ�oM���  h~t|[CS�$�4/fȮV��ZJ�69j�S�+�R��i�B��1r�[�  �|
b���%���y������)x[(�aK%`�f,iD	�]��p�Ӗ�1�����_�`���C�E��6��b�Q�YhR��h�A�O�R����鿕4�M�Ѫ�tK����k���^��u0�VX�P���a ��j�T�>Z�)�N۳+��hH�S%���0-5�=�HPiA�������p	k)�A60��K�����K���-!�Z� ;]�w����jzhR&�dJ�V�!���
�%�>�?5�)w��������f�Xc+[��[	�#
 �
Q�N�?F[H�tKN/�ZǮ0_�ԩ�Q�Ph����BLd�\������#��2� ����~�	���B`�� ��?�_��rxjU�6��C`VW��_.�O�x��@����	)~W��������#T�0(�^��h�o1�>RS����P�6 W//.=�>pt�@�_xI�Ё.w�	�������n�I��Z��wK�­��5�}���鉺��PQR�'�E�PjyC��c�2'CmP��粂,y�N}t(����<��P,��@�������Y ���DK����6�)*�h���qW`L|i/� �2�{�7ld�1Z��ǔ�i�]�1�	0�X��/�{�$Ɗp $��P����N-У�e�J$�n���Yj�d�K���N8IVZ�V1�!	3� �(w�����2���+~��^�7s�W�d!ؾ�Y�hos�:����zK��a������P��Z��d�"�{�����g�L;�4\Ѐ>K@�'_^q�P��j��FC�؆���Yjd�T���K1��s���'�J'	�����/0��TKt�+{P�����W�V����cM`�<Jg�Π]`�'���F�*�]$��h{G_GӧE6����X����VQ�T�CL� YX[���9����р ��2N������5���f�W�G$�~?�n˼v��ޤ >0��R�L<�v���(�ׂ��H��h)������<' �*�(�߽�3�˃��$һ�KuF�9$Z)���[�qQh�K:kYWHR��
a@ڸ�*yj*���5�J��(c�l[2B `B1��_1�n�pOh&2�r@�Y@%x[�9�9�lF=hIKD���:Vp����g`��ːJ]L�365yb�B	|.�+�ZW��S�,Ӏ�3������U��1� h�d�g����S��z8@�'�eD�-�|	p��(�{�KP�l��Ы�A�v>>�xne @ɶ8���͛>�cn�K7��t�I�Ll\�H;�i{a�F~��;�t4����h�[m��uCDHvj�H�� �X�
����d;�ٝOU�n		��w�pK�0)��k�&��h��V R��b�)��0L,�h4��%����7����O�<��UT��&S�(.�r�K4���Uk�zp���`�6�$L�j5>���V*����5��v�6���^�/��hPK�v�kq�&b!�YIK~�����VU�rX]+m�>�[Y� ���g��U��GHGO�/�w��N���1�!�X�îiuĻ���,�e�������1/{���Q/5Z`7M�_�R�V�R��`H蘟_��}�v��'�0^c���# �߰̩�\��fh:d[JD#�����~���[���K��z����%m�PqzG~� ��ŵW���1�.)T��ڋw�1�����`s��T�2��b4D|[x��K�'� ��-�hO6`�7A@#��B+Aߕ���@L�)�A60�r� ��
YF�>`Zh�{���X
P����ѱ�;�������?�<LT&��k$�����(۽�����
h/����6(��_yNT�&B����7	�X�W��>F`��[r����!�鋪@�Ç�0��+%I\&|Z���QQ������A��X������c�ݲ��EH0���	��F��ӕY?m\i�(U�4�����{H���<�%.��@|oq`rXc�n@{~1�] lJ-�.Q%C_bD�0�~���a�^!»�t��@�(����3�v�)�د��hQW�5�����'�Q�4���@ϑyN|����5N���р}�� Sh�5���j]`Z"!�>��b<�?����n/�`�!����-U<�f�	��Eu;r���(�7�9�� �x�k��)��,�%�w1��D�v^� ��z�>[X ��ꑈ�/ ����t�'��:�%�^�櫀��|�A�sw�y8��������ᆲ��&4;)��}^� -�i��&b5 �R�!�KF�H�ϰ�o�eg�.�'�j*}����^�<���aJ��*�/\fٜ��ЮYS��8>�X�;W�5wy��x��A����@'�#���!���^yP	e{�� ��b��
 ?x_�4+�zGZQ��i�`_���uVC�	)V'wE���^��$P W��\�Q���- �#��Z��õ48�����fY�� �b0؀ÔH���.�(�����!�"9��u ��>B/����Xl�`^^�>�~�|A '�&g�o�%���?!��l��@���o�Y_˩]��>2l���/<8�l�c�S;����N��k��M����ba��UGy�o��Ý���P���<X�,�����*�B-���X"��؝hwQ�>�.�L�]�%�69�{���b	�L��Q���?41���'l�4�X�J�B��Q�_�"�J
2锜 ' c,�GH�?&�� -qU}� �fuv���	�"p��\�`z>)����e9.������Q&Q1����e��]��^%F_����R�Wx���A�Z,B�5�k�0
�V��,o×�����	�\�:�����Lw�$�n���Oʓ^⮃鸻Ud���<��։�)�-�&�f^��Iҧ�WQ  ��y�G-DEۓ@�^��n4!���NH�h��ĳ��]Q��7Lx��,;���|8�� �^瓸ٹ��@n~%PB�`*���8�l���@a}�q��ݖK�
;��8�6I�WA�5`�7��E����˄���:
w	N�� &�<_?��)�f@V�A:l/�����1��!�<�H�P|?PY���,�@	� ���^x��)ms�^ ��:>Lh$�\=�c�7�@��f�t����Pm���4���+!�N�1��B_�f���L�X(Ӹ�'4q�w�z��j��P�C'nS���?&�/�a$R��&��AJz��[�P"#C,��H`�)�-Ȧ�5֫����A���ܛ+���JX�`��Va�Phf^l?�F��Z�1�D� <R�7�9�"ʊZY�� ������G�,i�=��zL���"�|D�<1�4QxܠX'?�����l���� �+[�,O�� ��çW��� �&�uKTN� S�1�P_^�>Ch�tO�󒍘zbm�͌j��syz�iku.D�c
K�T�}:�<�	�w�T���T�ߟ#�� !���W�0h�)�?]M:7�(O�ESAeg K�Q�n)��� ɻ�]N����ք-���՝��']ip��@(�V��K���3�p�{�'8�[h/�5�?�	?���� f�a�>J ������z� (r_��v˥��e�)��0Gh�|�
��i����>�jK�^о��Ru�?A�rہR�;�,�R��v����~����z�����݀�|@1�bZ�@g�28)}�'�B"��|0s[�l��Θ���P�&� (�*�Ti�z�F��o�e¨��9���(�[��Z�����%VO�[�d��8Ʋ]&_��/�l�J�x�z�1�_�����󄲼�P�'�BUŸa��}��M�u)k �=:��x�ˀ�XM�m�>�B����ט �N��h����'�_A[�׵�e}a�'I{�1�τ/���v�iD��t*�u|	�ev0����CTO�����	���l���V��1���v� 0�(�_�	������P��P^�C��W�\ ��1�)���W����
���.'nk@Q��J��3O���qRY_�¡Z�"����ffSSG�C9�Yg�P��Q�.�X�h]��P�O\�'�C���0v�5^&�"S v�A=��1��ڂ�.`X����[�@��\'�`BW��$]pN�)�w��������W�z��jw���p�-��m��b���� ?͘IF)�/�w�-��.����, P2(L'�/��Y�����p������a^+��*�� {�2)�-�h[H����2^/��VA@��]�/��u�E���*A�j�/�8N�7���(R�d��feb��wV�[��D�����-�R83>r�,i:4�|/�V��t�A��6/0.���bk�P����K,�G� �hJ=�wJ[ꕡ��\+��@��''�aP�	uP`]�B��#yk��~�b�UTl�\��z��"J+��	��֪�J�:|N�|�
)�HKu�|���D�
�Wh},0���>̘�-<�HMx0XƎe!N}PXh3��%J�%�tU��l��#IW~���J�����ף^Ɗ<w� ���ɀ��{�?,� ��S%��:'���U�A����i�_�(����j}�ٝ/�z�3����(���_��V�K�Q��b�U�����1�H�z�1��SB��	�m�	A��Q>%�?��h�q�����nr�>�:(�Amb#�@��VJP3�����!��"�M_�GA�5-��=>KNS�l�Oah�;f5 il�C��&��p��c[����� f�>7�}�>V���[��N�
�H#��Y�m-#�w��$|�OIr_:���5��z�=n�J���-o:�_�z�"l�x(D�hj�֢xn��x����"%6�;�=��z!�|�z�}�P&/z �A5M8G7�x�K���.��.J���� ���!y
�`�)��*Z���xZ�'D
!��%��/����g�`�m|�~WRU�9:)J	,axk�R�Z�@O�;�Z�q��`}�.M�Bp^���JE �t�Ѹ��W �-�D*})�Q@L��JZ�sA��u0P�
�e�(��P�bq0 �Ŋ�t��{��p"=O<�!_!/�b�C}��+P!ʣ��6�̔'�SW����?�˼�{d�lK��h�Ӊڀh�'E` Pb����2�Ռ�Zڰ������(	[Yw[N����[�?9h/�p���?*O�o�D
��T��W녌��*��Q�<h�s�KYtD��;��1~IR=tB��	�"�*)��`ĚD$Bn| ~2�I��;˚}C�P	e;SC����1~��|�Nx
j�}���U'%�X�,Xht��4��(�}���J��n�]�5zJd�[w��,��[є���'PB��MA��i�0� �[���܀�s�v�����0o�˭: Z<��V!F�O���N�4��_�� rQ(�)�h�>-T�i��O�|�R��ŕ�8����'!���%���0���;T��Ñ{��=�2��0Ot'.]�H%R��H$���@�*��K�DZ�}�[�P1YXW͓o,�!y�>hC���[��"/
�s��2�U2����� �(�K�+�n�˃#�f(%2�-4	�V2׍ZR���-� ��cP�
� ~�^��40���-����mpU�"�q	����Ť�I�]{}&=F��iAx}%/aL[>�w�n�L���l~���<�1��yA���b�8�Y�	'��D����p	�Qo�/�tK%��l5��%�WE4�P�r��^	CE�e��8�L���~h�R����[�#���`/�5b1U ���Ne�P�%��ax�0��J�|���0�G�Bڡ�	�\j��t��%)�1W���I��Au�0����0�Jf��0ӊkU{�D���HS
(��� �P�)\���D�Ke��+���<N�>`�Q �S?!�1�h%J4�`
���y�N��5i�����K,^��:H(O̽��1�2{�;;(���:�S�t�6K���%2(ʞ�Sh���Z(�a��h�>oi#H����}��wt��w�$�5�B[�		����\L(����1I [Y�s�#ៅ`����#�u�@U�Ds@�Zh*�#� �6O�Vͯ��@�iXP]�	�p̬�8�w�P`�?-`�>.�^� K���:J.�|��.��@����(�ӑ	1�h�_�)��рo�@��H��J�L< +AJ�WT���T.p��B�U���]D����p��O`��nó�`��+}�]��Ԑ���磆�lQ�޺�dX+����=��uNl!�uƎ�{��v�G^��n�d�9�{��
Ư���c�YY��
+
p	�W�b3	��v�	��/� L+be��� �2��RgQ�p@�_�H/o^K+C��@��A�`<J*=����VÀ���mA�NWT_jh�B&L���#��g	+���0�b�nL��EU0#ZPF��<�U�����՝%:��n��S��&|��c�p �������НXf^�P[�/�~��vQ,]#%�>=p^��K'|2~�ɬK�����p����ѷ�u �;rq+$��Ƀz�U�V59Zm�yA<:��4<��D�<)�Z}�]^������Ou����J��5���%���N߫��_���E���@�n2_[]��/�E	]M��_���T	dn+�ܪC��u��4@��x�u^Y�i�������S�3�0��I�ɠ[v!��G��"�T�O/d�?��J2�^��!��^'�8Uged�BUa�k�x}����x��l'�5(�V�!���|��1�!G�y(�h!��RşD
	���wb���L�	[P�B�+/H3U�!���D= �+J\��hq	���'F|S�V�X��PʐX$�6��^��/[�c ����@��~{B�󹿭�	�3�Viw���Q��?�- C�%(�5�F�������sO��͢j��4N�0���*�(9��!� :���G�	5h&Q�3J5�|��O1�|u&]W^:z�o�}`�-e�q��TN1�*�S�D�H�-�Vh�}��;^>�N�Y��0}�QԐ"�/J����urT@��@q)�`H�0|=��O[L-t60D)�b�V�
��TDp�Ƣ-Z��C�zqT�� r�$1�鴣��X�������h���TRb������yRe!!��CH�&5BjY^��h�1?\qPV����f\�Y�I�h�UTW�*�[F���eȴ���[g ���,*�[`��h�&=V]�fܭ�"7�Lq|oe�����1*](X�V���o����� 9ZYO�N�b� �]R�'�Ț$p*=��ڗ;)~�-���P�a\=@�����a9E��w��F�-t�%���Q e�u�~4u1��o	�h�Td�{X[¬�C��v�(����-(uN7ѬQ[҄œ�����1�W�(
v6��|Q�E�2/Ij�Wd�]�!J�ጶP9�'�>o1}�G�n��H줰��.{��Ζ�d;��,>2��w��������μ	<�-V�6��c�@R����:L�G}�ơ�J���(�m 1�6Y{[��/�� ~�Q -Zu�'Q(Yn!����B��ڼ'�\� �����[@-�GR�rX|]H1 �_�ZW�ߗ@&1��
@|w�n~awo�P&���.���9��#G��]�8��W�3��W���//f�h0�[:�ɖ ı:�d^�i��K2��׽0c�hk(�O���$���LXL<0}aU�[�����h%R�5��H��t^����m��	1*���&�("	OB�M��`�h�l/s�,�����y�8�<�d���X婱�f�o��BJ��-Q�Bf@�	���i��%��B����\�A��٤b�yUҽQ{�-	dK���*]��	�e؉��p��_��%��(���~�A�ˆ�fK4�-\.邒����؉����X�N�gb�ȉ�}d��<(���h��S���!�?�:�*+�
��&�X�EG�3�ێ��L�m�+����P��-596���~?G��(�H�:K����o
@R�V	^qX�w���}��J[B�#{���I�-�����u	{�_���YU'C�S}y4�83o�Y�;����-T�Q����L�Kt��4`���,�^�H�XcM�&�_Z�[�,��=h�`���%Qb�3oD�>��@K����Y�f_�w�� ,c��0�'fXV�¶u�'���^T��9I��ɭZyB�"aa#z{4[h10��ڥ&�>�a�ρ��|DF�>�_#��[�~�Xo	׈B)(����<�h�~��y ae�|n��[7� ^����*�ں#��y��'Bpd	/����5J��Zη'�0�~.Q`�!-wX�2ˀ`��uj��J���i�����B���;���Ѽ;w-u�����J� �5��Qo�X
�8�n�cP��hK_q �4,p�:�1Y0:�.��I��l��*�����Y�R��]������A��t�F�Ka�?��H�K�u�R�6�-7E�C-�w�~��ZV��a%��H���Y�''��ߐJh�&�ڷya��\j�IQ-zʭPF���z�%5���>�F[���̊�D��P��	4�$�.>�G��r��5��f��Cq���w�dPt��pW'��� 8���a���c�Q����������Ѥ�����0�}YcaV�SX��0��Dn6�I�oHi7!z&o��4�Q����S�X��/��yg����l_,>��i��PZ�, �2�(*f��-N� �������NPVX^��bI�}~rɆms��5L�7T#�X���xPH* A/������cI����%�tn/'��d�P�P`\
�����f�&�'tBQ�{)�9����%�IY0-����-��5�'�W�wJw`P	!XI5~ΟV��d�{��\��t�m��}�����fS�;���IC�PWv ��}�¶/�W(5��둌i:�A���(��V���(���[�KZ�!Ӫ���u��7s�He_���%p dtJ5cV9-1�ا^4�����	��%�X�'�҇�iw�\h�c�5V��h�A� {P`�4S���\�����F4��z� &�t%����	@����U���A��������]����h�|��d�LP�O��T	^�Q��<u��ԑ\'m�H�� �4��1�uH�� �cG~-B�.�)�@��F Q@~_"W5Ji@-vc��(?{���V�Xa����pE^Ds�U��%�I�f��Ӧ�N]��v����~���_���N�-aX���_����UZ��'�G?M���,�Z�/��AhEH���;&��D�]�E �X􉫗��h��N����pFS���T�H�WbHSF�(O�����{�\t��$�-~�&� W��(�g��P_ѳ��]^2I�v�_�@F�VK��k�V Y�!oy�!�^0hӯ��5���Co�+�h��z�WxVRP>�%}r�#�A��X)�R:`���-EU�K�ɾ�Π�0�J g�R^�1Y|�������H�.��	^�|�U����嶯�@d�,X݌�[�Y����Q���� �fΌ�Y YC��	g��z	|�����'�sH����z\����f��������]w>�H���sσ�]�)!ÂJ��B7[X�rs?Ua��gVYR�/�	(�[H�m� ���x�P��`�v5��1�yY�*	c�"�������X�@�lj#�;�-���~��ȝٞ�B�����. ¡q17�W�^jg����u�{T����?��:�6s�>{���B4_aMA˴��#��ǈ@�{O�Q̧/54
oH�&��e4��	p��<a��ׂ
t�&5E7-�\�� ��S� �[��R�僆���g?��W ���D�w�'�gX� �z3ot5NJ �d-��h�QS�n&���	���E���:����hl�.|K���%]e��W�4Ϡ�Р�"x =zU���0|1]!���Q0bݧ�0itR����Ԩ�XZ�Ȏ�X5&"e�vyrq��z�M�;&%����S��-�mb�w�F�@�o)��SGNM�H���,�\�I_�=�u���J�G���{�@��z�B��,/0w׽�Y����`��A��1Tk�W%���/S(�Q� ,��
�'Z1�):n�G7�V�0��b%9� � ��GDV�Y"�S���QE����
�8�'���i��^y�B��wD� U�#wKh�� ���R]�1�6�"��М���ȵ�i<� B4�h��ɱ&Z��#���^�ðQ�l��|��������(�N��]�: �vR`h1�w����7�P�Qkmi	�%l�/ 1��?{��Y�0�BI�.�}�
"<�_��'0��	�)�wg��p��U \]���A�(:�� -wl6ƹ+d���ɕnѵ�f	�_��j�`�ׄ�ꮟ���u<�0�9p�����;,�ʼ¸�[N�1���D��ʍ��(]\�P�Òh/`�A�H��~�y�X�rx�L�)�6t0������v�l/eS���N��Պ ?�QFz�������Ov4�Z&�f	������C&e'B�L�شG��W�v�YӖV��.��Ͻdv*�@d�m�}�)��U^�����T�����_S֥}E˓5�ʜ����1��-mk.�b|C�C�����8.�~���f��B ��v�@���(~����6�@���S�g��b'��&�N���%V�UG�	zhYC_������8;�	[�s�� X��p�w� �H�;-�W�%���UH��@���vW@��
��p��C�3�n���2e�`-锚Ӌ�1�R��3p_�)��i~����}A��	`] �'�A��	*[�(r2RbB4�.�sW�� ������L� _v\	�=��~�A��IZ/��*�=�:�<��(���Yh�(b6��R1���S�)9��;Z�(��'|��+���H���s}Z��)��~1hr�A+����:X��(�[��Ե����8�^m�M��G�T��S�`s��[��$��p�J���%]�'��Dz}7�����޴�X[��Ӣʃ����fQ���������E��6�>Z;���d�w�� �eY�(���âx��md��a[��U�Bx�̄��:lb��,�Z�!̉�+�8���=,�5�_��ie�h9��	�,��L��r|����[>�1�9PG$Ad��h�Fwn��t���o�&-i����*��y]q�s;k�n�`P��Q����ONy�d��×�T�A��>	X����p��P���B�E�|O[Z����z���k/:��h7��U!ѭ�X�Sg���|u!K:����RU60�_����>;
>�!x��@��j=d˼�R��+��ϲ�w�	-]B��3n�Taс�`z�3��/�^�w�|��	�@� �����~�y���LN�v9����<��	��B�x�w~��x3*�Q��Xǲ�4w ��*0&1���B�jV<�椾�a_�X�lqC_M���3-v���	��/_(B0�?��?���L�%e,�׽+/$�n6�V�_Qˬd�(��ʲ�x�h�Z4��W��R�R2,B� �ReTE���j�=���jʧ
�H�������#.�(�0�6�� 
�f����uX|-&�����?��I�S�h�-��Pعf$��	�g�JR��k[]x昚��^aR���2˝� �[�ц��c�}�ɤ�O��X���I]s�3�Mn�f��Q��.������R�����qj�tA�./{�8�S�i��[�L����5g���s�];ZtK��̐�e�#^�?A������B�`ܰr+�J���������͉4�R�Y�0_3VG Y*8`}KHMe	mo�dXW��P�H�5�P������ ��BV�7)��Cb�~���βH�?3��:����OH�?Vh�e0~;�X'B�Mm�A����l�w=0%��H�m�_:�c�������?>`Qe0������!�X��=��sAl��အ:����P_�V�;S"P	:sg�{��9��-�t$�9n_ ��*��I"бO����x3�`�iP� ��S$��6M�sY3��)j��z,%9�%w��V�I(�.�'�8M���BJ��;]U�'p4{�U�@X*��� 	_����t��Q�M��[ �3�[$u&ç�Z��
gp���u�y	��qYb��/sZ`�bx�#���d(H�gU��<d	�]5�R�C)r�	����$��.�3/�d�t�U��v����	J1�=��$W�=��K��w#�1�������zǯ5��j:����Z
��A|U��
�#R!�ZC%Gw�u��8�Z�(���@�Y7u%�
� �5z�r�㈅o�I��,:!�J�}���既Lޤ�yhj"�-�n������,��uM~eq�(d�E��^�L��M�0f-��dQ�`P	6��1���y��; �ܧx$GL�JyP"�A$��?��g1��M@��w�~�z�?9)� �1�5�<!=r����@�J�Y��覓� ʻ�l�+�
��VH%�`������X�Iݴ�Qd�reƇ�P-�G�)���	zT��G��h�X��]�/��<ԪZ���n� ��(�v �<@	%J���')��]ݭ$_�,�@n���e!��"�lj�5}	�']�RR=\M0Du#[Hs'��B�}����ǁh�p[уjg0YLX	H-$߀��8J����1�!���Sh�Qnu�p�C�Vez�s�8w�	�c��H��A�;�qB�Y����"�Ƴ���1k�T��~������v
�bK}?wx+Q�ly�x݀�3����\�@K�	|��`��(`[G�/UԀ��'�T(m1�A��O���Ӏv��9-"AW	Ƃ�O���a�+�Q���N�<���(_�6�B�k��Z���{@975x�{��%Q����	W��0�Vs �
�<%�I*�>�&A �^���ՙ��� ������5~3��<�Qbe�L�h��/�@�E�ʊ�Qc5�i�_@S��h�+y�"Pݕ�b(&��@5�n�*~m��T�_	�x{ Z-q )ڃ@�8���̭j���k[D-��YD���V�~0O��JK���K���o|�����0�!��(��Jh�-y_�&yo��p.O@��c Y'Rh�94H�gǯ�I9H����:��/|���A0�B��$�����aF)�A	�q�j����;i[�p�X-E �0{�#Y�r,1�r����5JU��zN�i�*+��������(����H�)��#����e�0;6��UT]e�@�'4�HH������}��F0��2�@xhZY���&�N�阀�WkoA����.�?�%�}��r��~?���D�.��٧w��'�*�nU�XZX��i]���d�g��Vb=����8��{b���J����B�ȃ�w��i���<��D:ʶ�~��Q�G�k�1 B�K�l�7�z�QZ�+ om��A{��Y�����sd%z_�Ŗ� 5&X(Zh	8_�|���us�Y���*�f 5eq�]��t�TK�A��?غL0%)�Kr�K]0w�`�6��ťӅ�\H��_�lp�|\��"Z�)�Z�%�ݜ����oRюB�ԭ&��ˁ�����i�V�;�+�}�"���Th ]��C p���-j;���_���8Y!y��[� �H6�`j�Tr)S�={�cp(�Y����j�J{W8(^�-��t{BU@��C݂��o/��\-���]���Da��v�g1��:��J<!��������Y�x$�2�.q^yă,��f뀚��V.U@��v�	����u�ć�N{������*'>R	���� �:�v�c�C!£ [�h|���aA��D=��G1�-�S^|���F�������������T	r}I��!������b����i�@��z!u�p��Æ)�1�@�c,.M|��+ ���w�l���8}%��H������Y��g�$��:��<����b9�b݀�P��^A3�;p+��
@�_�x���i_�-�����$htL3$�ċe���bU�c&��7%r];�M��k~n�sjp	��:d�,�U8��3)Y����HL~��p9�.����%�W������U5��
Z�Oe�?Ы��'M��V�{�6��X�/$���] �\v?ZP��>��"� �rM-�0���5�~	(hy���=�C�F��z��ز<�C�%3uł�܁�c�d�bl_��h�'.u
L
K����@I~����_o�	\1Wٞ�p��?;Ï/�J�h���c��� F~� 5'-L�<?���1��eWlג� q�)�!��*�Ⱦ�n�;	ho��l��@a���z� 0g ���(�����z�5����-BZvh�j�a�G��ݯ �6|h��F�SS� �<ceXPZV�*�|\Ss~=J6a�7���P�����t8��Y4��=���݀�mvw�� ]�>!�1��q$����!�*�	��`)\�
��࿾�Uq؊h�Y��g+6�(nA^/����}#hl%�e��{�}�@�.1^8ƌQ��h�t	�7�F�-��!3I}șSu��Ԟ@�i0e^��J�9�����B=����Y5�) ��CF��;�����5[	�XUT�q�yMe�k�H�|l�|- ޑf)�1�Qh`n~2�i�'Z�����s4᫕�0K(�A:A���\UǍ�';uR�E{��A ���l@�Q���Pv?1ٚt�J��^^SQ" ��2�;<�x
�vE�F��q7+�KQ]�	� �#?�;[�ڭ����dJs���t_ n2K鿐x�k��[�@AGmT����J�5�U+YX-h
��V��<�@!X��&�u-|N���J\`��./�dqSgv�hNd�4/�`L��P"�x�����^���p-�:���k���N�<E[�<2� +�G%U��KWČB�H�?�b�(��� �<sV�1��D�:R%�t�~8�Yp��2����
`�ŏIĝ 
�zx?��@!��T+��c����2���� �w�rX5 �(H,I �KQ�a"�fN1��}G�zxH��X9-���;�Dfx���/�5�≢��F��h�]�����Uf�+��%9p�O���0���v�&��+ٻT�.��n���AC.��&#�!a�ܻXh��RFZ�CN)��,�
E,�s;v��!�P�����������kP�����h��Mc���XJ���,�H�>�@6P}M~��	�h�iF-]Z�0�O�_'S�K� ʤw=aE[�@���L�*���=s1��Ӆ*��т�i�KŰ#:`OJ�S3]�&�0�)��\L�m��HgV�C��^h!�z��P�����ji��j�h�h��tZ/���-yX3�%WH �w.J&�G��g��F�oF�W� ]I̜- 4hX��B[�����!=���\Y�%�K]tw�0_�"Q�R��e��\���� ��5H�#N�U��w)�aUDmP���������hWFe����_�������/R�{cʣ���~�3���� ��Z(���؀�j�k@C`�lE) Z�aNs�v���xйLw^����$P	��-z��~R"`���3+�5@X���:���G �:]��8�<����Bʝ�����	���"��Ɋ[�|��Z ���� �Sh�\=~ЉZ���n�]�I��0{�5��g�eo���tW[bAkR�`��UZ��:�8B��o�.���릤�A�1�@e��D6yS%���n�zh��O���C~Q�^�Xϕ߰�:?�HU���0g&�l���N�/3�8Ȱ�,x$O��������JX�V��UR&I��"��o��9�%`|5��ӏ�B}/L�`ʽ�
/3
��	�@\喒�j�)�vNu�U>1��8m�d`�SQ]d�_���76V���@ώ�r#�*B}�"�$/���,Ƌ-�sY�ż��)�]�z��
�
0�L5��$_d<.	Y�_��W�x�*B���@C�S�{JML��8zf����,���/`�*���v
�T��7N�RG��#�Y��Z���X~S��Q�G�MN\�N� G�bzK�Z3fJ�4B�"j��'zY�ke�a�D�# o�3C�pY��X5�	P��q2�|L]c(��OE�za"�K�NRO��HF��C�2Af�F�K�M�,���U�6�ۉ�9�"�H��-RZ0��@���g8~��w�r�;7�`��B��s(�0XKw���i�1��S�r��[Z�YP�h�F�K(�J�`��V%'�9(Șa��C{���H�����b�X�l����"2%�W�`�%i��̊�OK3�6����-�����l��lL.[���2&���RZ�閶���-Sa.��
�`.���ڽ�{y <�(e�d���%��P�!;��z*��&�	H���WTa��D� ��:�}qI�H��ω;߂`!�w4D@��hPP��1g� ����SmT�|��mGR�a��2E-|�.�J�0��L%~�V;�w�`�I��	��U@P�N��{D >��	�������{���Bw�M� h�p�,YA ��D���"oL�� ;IAU�zae������n0����v���R��ş��&1��SB�$z���Fx��-9P��5��wz��� 9-�r%='~� Z��ÄN�f���r>��� VJ���@�6饊�	s�MB_
zX�^��<,{�ŀv�Wh� �'*_���
(���is���Ģ-��X�-�sbŽ�߇�A�0��G7�9d��u'u�~jO��>[Q������u�Y���\	�%r� �X��(� k�rG�1�ޚ�@#6��\�-�\� ��ϵ�}�R����vO�8�T_��S`�n��D����	�'�W�B��2�ۜ?�y�"��IEл��v9F)����	a�@?Q(8N�*����������w���=��;1�^��X�6p���e��o}=,=����0N����2':|]F=�D�aX|��
1�)�̍�� 4�[=�n���9�h�'�m�46�@mH���ZUP�᝶�H��As=���bd��`��B!�_�mYE��q�![���t��qK�f)�=�.��介�Ԣ&� �%zX+��5D�	k���Ѹ�@�?�HF<:�i���{ �W��Fc3�$�4��!*P���l�+�ͷA'?Ӡ���\�y��K��Nl���-�%��Q����t��"U׸����^��T�i�ҹ�����T���|u�B�PQ���'���'��x�0OH�e[����[�� �UH�b$K� ��v����X�"X� .]K�`W��)���sc�����ʻ�<�_U�}%�ҡm?�!r�x�L�2ouW@Y��h5�3M�b�C�Q����-40�|�CO\I��W�)��\\9%�/�?s�N���t+{�qе� 8�D[�P#�Tm���cSYQ�"35��Az�'�[1lU@�{c�J�a.�f.,�h7]f��� ��v?n�骗]l&LV��A[n7E����nc�=���m� ���?�8^�쁵O�c��6ŀ��J����}c�~��#��`0�
�hsWi)��XZ1vw�f�G.,F�@qR0XP1]�KKx�w�
?h��һSw�5lF�%=�b���=����4
��π��_�` H��j���>��,�0v ������||'�[�u�Ɖ)�Eg�րr�(��%���Y���J6��!���~�pX�(�����<n����C'yC�M���H�vm�q�_��W2���XSt:`Uh�靊�v&��F�IH .�@�5��A��7xP:�"�&B�]���`�Դ�b��	��)�D�j��h �Z�8,* 
^�Zhv&�y��L� �	�g����SP�)�[����2�=��x�d,W�@�ٽ	�h�`���d��I�eN��I�����`&��*	�9��U	ga�u؊�.�ᄅSe��H\ tM�:�����|E�Ɯ_E^�Hõ؋��5�~{hH	�1��=E%y<�H��� �x-�l ��8���JS�*C���r	h�6yE�R��	@w �
%1�0��(Y~��l^���7�D��L?]!�[�|%hg_�A�MjoD�+��;�vY^G��#z�JH����Et���'_�C�D���J	@?KE� 7�0��	�!�U׈O�%Q���ʙ������@�O��Q�S�=���������0��#��A���i�Um�f]�*�ߝ�<���(��oǝ�(�?�Vt-~�QK�$��T�%�,z���Ru1r:��źs��,Yo%�QD	8!���s����A5Vz�����'�T���˝��­��bLϘ��t�H����'�����7&D�.wږ�W��s�C���9��_@�4��^�m* (������ oF �
dw��A@{h
7�v�9��B�+���`�^��y��W���D_T���u�	��T�� �q��i_���{�Oz��AJ�O��{��綄�����8fK1�'����� �s�}����%�WE����6!y��F����}#y4��Qo�݇
*0ʻ��^�l|0׈� �/XQ�2���x_�ܸ'	U6�\q���#5B��|x�fo]�Y���c�N)��y�	]��`�D(+g�ڲ���!����OӀ�)��� 0@�=X+:3O��� ��m���]�`������1�cq��hD0�y[����2L� �)�:F=k�aQ!�.��|B��]^)� ��L�t��7C+�JMWtB��WRxh����Y1*�Bu��)��'>��_Q�1��6�	��ڂ
��u���ʥ`��Q��/��^y � �4��w���i� *��%�}�{��mZ��X#����D,F�غv�>���/R
)�KY0"�K'�&|j��?E=_ �oZq����E!�O��^:�g��P��l�}Ѱ,Pi�_��1V¾)�g8h�e@��Z��{��(�蕝�� �f��]�?����Ad��F	\_%��,��3Zm,X�;<q|`n!�bOS��Fޒ�c��hHx)uY1�c6�.^��d�[�	�z=:�Iu_�.衤��9��!rI�3yd��	2f�	ul9%��_��m8�pD�ѳ�����e���縬�kq�Y�O�0��K	�d��#qC�(%ЏN<y��XA-�l�pkYB�� Sh�;XZH�% E����Ad�M�0Y�DlEb��(���e�Y�����81�.	�3���)�� �#S"&�t�0���=� ?ٸ�h�z E�-�/&@��������e5��^�^˦(�Dx�D��}�o%�!.A'W�'	� ҽzn�\�Q��3,N2�~����g��������7)b�(�l_��8oG�V�6]��\�! ��.?�%}�+����ab�$Z1!ٺ<-�%�C{�Nƭ6;�1-�%*���|�';��&�w u8���Fj�P���-~�Jp�S4א�4�e��Į��+�h)�f�j�
 �G�*{��.^��|��e��)�i�K���냡��9n�#H-�p����?�'r�P/�� ��o�H��e]�\�����P�d h�����N1 �p`z�_G�N�5|'��͑V�k�]n��1�	�~�)�Yi@h�Qd�8�4���^�_�����y�<8�>F&�� �| �����l� U�Q5(S���׬ ���;P��q��'h�]> [;��n�G����L� ?1��aD��n�H�
ze݁�Xy<W+1�a?���/���1�������L��Էj������hh;�Q�4]2W����	V�P��_�zy�j����K��^�5G)���|��]2f�f�"�0��Q�9CkA�I�d�p.��¼�Ĭ))Ӝ�:�I�� �X�� �zΨ�{�J���Q?Z��ⵎ���Nw���5}2��`��v�O��h���!�A��<�l�;v�/�~��� �Ht-v(X����w[ Z�FE-�Sz�rN�	���2�X�:����=ϳf��7������QBm<_Fx �N���G �P�A��.�6R|�}������@S�h;�0��w��zՖh��*_�ҋ������� 
�h�j$�	W�{�0����Ƈ_b�Ѐ� ��g
L��*d?�AðY%d�S�	�1lo77GN �-cK �)5�1�\R��@�	��C��|���(�/0L�4�
.�n�d8)�K�TP�w��MN�邆W+^�Љ5LU4!%a�x�oPh�WU��-<MQ�$���q������P=gSs-�K5t`yX�]p� ��T)|(�F������?������������o��x(w ���0�W0�{XZ�v|P?�R����A���D�!����`6�|����/�%��)�>�<��2Z��oV�~Q~9�W���)Z ��]N~��C�zc	}�5=}����ħ����㓽����F��1|`x����Xw��A�&��e�0�i��ZR��<��4���] ~&E�<���]���qX���s�����3k�qIw��"{�_��./�*<K�wz�Ȁ�X�u%(�}�������X0��Q���H�_��L(�����"�*������3IW��%t�^LP}%�@Kg�����,X�vQ-�vnV�ܘYġ�7?�M���X	镆�����G���b��a�lx?�R]���)���Q�m�ȃ��Ҡ�� �}H�X�\���'q^ ,�(�ý�&)��\���e}	���`���P���\&
F�!v'�jx'1����!�Q��k�sg:��3mL
�c8��]~�@��/ 8��5E:v��q(������L&�]�>���@��xQ���ZA-]���f�X���? ���)��2o�}�y#&� H`*)L�t���T/��}e	�Q�3,	�x�U1�{�4�Yn�.+a�\h�%���	V6iWrY$PxQ-]2�wQep鈝p^K�����yu"P�ɢ�]VW\��8��b^��eJ)4.�,a?B�L.��S��.��|(V�	�E���v��/;�:��z��	|H� �:\�J)�Q�!91�������-�J���Gi�(-��>!�n �Q��Z\:ȱ�pw_`@h�]���� �Q��j�P�W�sA�>�[��g��e����_�7~�fk θ4#����O�Ёx^I0��q �f 8R�`M`j �5<�Lzl>��G�@L�[=쮐��h�<��%�1��h�U!p�@�������X 0]�-	tU*�|:g�x���|[	1�ڮ��4����)�t�c�N=[��	}`G�-�ĺ�W�c�Օp��H_�Ԅ���������Z�/l3�;Г�A�gh����!)ua����x�WT�ɥ�=/��!��g� �S���>���~a"�� �}`>�/^�^	z�`j'Ph_#��J62Xw���w�0y	�>H8`�<x�`>Z������|����3�om ��O|�Z@�����$�|�SS����S���uh-y�-�`��	-j&p^��͋�^��/�k@P�n+B��o�3�T�ٴ�j��-|�ah.�ǃ��Zԥ��+1v���Y4e�� ��x[��"���U�|��?<��w�� Or��ZZ9�5U����X1y�՗�����C P&��SK�����)���{D�?���G r�l�O��QD�;��zd�\��(���.�'�<�/����V�14�t�܀XS�F\7�&�� \R��JB4��)�z�`�v��L#^�Y@�I�E�:�@d�5�q��p�[�L� �=�~P��dR!�Xa�i�D���50gOv59 |3��Y�0��[4P��-P{\I��t\�V���A�N�}PW2�Z�-�3�*J��sT�'yp��_�{꿦���yzQ��A��P���!8=I �Z*���\h�Zd��~�_i3n��p�h:V�?I� {�G����e?�{�X-�1^�'��e?��K�bz@BWP*��y�h��[XD���s_T�c��o�(,K���/(<��r�O���!��N�iZ!��3ݲl�Zс%cE��ʤO85�D;��R�b�2K�����6��.�O
�CA;q��10�t�9�����B��隯�F}H��hW='u�͙0?-OR�� �G��'��X�I���M�Ԁ��g�#o�ӳ��*���;�"����B[VsB'v��V�*���-�~�E5i�I�D@�5�N�K��v�E���D����*���e1f�|�-�)Yye���--Ri; ��դ&� 2�W��2�1�`.i����s�gĻ,$h��]@y�����;�|��n�Bg��_��R���X	�	uH��>4��mz� ��10<f��k''�o���501��Hߵx��Dsr�/�5�һ	@]�
�fz<)�A�E���d�H�H��LAS�G5JD?ǿ�##�X;k�A�_��+7R�V��3~ŹP��yE1��Δ2Q��U�/�����(�-�c`9Rhs��jY���"LF�0x�v\�S(rF?�
�M0S��NY\>4�J�;�vA�o�c���j+�9���ycA����9���Ec��W��Xb�+�5���{Z؅���&�W�w�R��1Z������aO0���?�g؎���a�
� ��)ս	�{�  �s�!�[��(@`�)KB�B��x"\���M�-�ty�I� w)�&M [P�)#"u�̓���'Vg�#�U�uzE n�h�^=�-�V�AP�K�6�>���/1�����|��p�_٬Px��ƽ�T�Y]��@���Ӹ�5���I�.��;*����c�Dj��b�&[7
�9�%�p��^�-��.��e(��v��О06�KM�S܄[V�w{��ev'ג]�
 A�-4�������L�A��e
�Q馫�LY!ź|~1]�	/���	C��ɧB��wĪ����J0т\5_�#�T�L���A(�O��>'|� �-������luI;,p#`�w�l�5�y��h[}2="!��Z\�,�B+���:`�N-�����o'0Oe��ڹ�f�nr+�bt�,���}$�\�;W�7Cz�j/J��#^o�`��tN�B�,�o��$vO�!�)#kwTRp��%f(I��-�@g��K�en���݉e�,i��9��t�Y{	�Py� �uk�T�8���hC��t���Q�q������K���(����E� [Y�5d�tj�� �&�J�1Ȃs�U���ЛŚ�]�-�eB���A�,mD���Ɣ[ >�c�ނ�Z+���	TKm<]�s�W� ���u�F�e��к �B��.��z��5% X��kH�E+`�j?g�-!P	�2by�o�unQ�f>��ph��=n�O�E��-��q/�wX��{��Lۙ,�l��V���F��_z3TŘ����[��q%a��{�vS��N�	��e�֘� l����3J��d��y(,��R�<��?
@�ëxx��-�!p<�)�1�ښU� WY_�P�T?c}��ٮ���<-�8�!�� ځW�`q�(������?�	c65 �49�+/��qr�ߢU!�:���qJd��]�X:�R0�<%S����e� �o봠�Jt1����% h�*/Uz�y��</u8�Y:Z��2��Oǉ��f)�	X���@_��y�M%����|�}h�]��Q9���v�2���� �r�2 S������*w�/�M�� lv�Q-��u3	�����X�_O��!�r�>%�Q_b+��jY]`�r�/����hUV�9�,��`���@^��/�� �,0-\�1;_�{c"��w�	�Z����'�18��V��Q��E>=u�JbF�S�4L�����U�f�r2L�tdV� e߿C!o�"H�T�� �]�����4�J�����;�@'�a�I��N�	hu��*��sz�5{Z6�~� 	�h�YB]�2�wo:>�4�T	&+��}���(�v�,I(�XY���$��^G)��&���e��l�8�@�\�, vyZ����<���J����*V�4��wT�'��.�[àB�MP\e��wi��08��e-Z_�zfK�� k�@uO⴨�C��t7�0�W����?8['��U��Qhm�
��I8�ً�YJ`[hgw�G<l`�7�m����Oب�R�	�� ���MeM)r�!�Z��W�f�:S��_���_j���`1I�XYX>�-�o4���XPj��%RZf�,/"�ELP�[G����yL��/���A��̰-	NH�%����^1$J	�&s�>e��i.Id ��K�C��鍊"@nr5�V[w`O�W�O�P�Y�?�̀��)T{�X��v&�|�9q��W�.�@�R�@����Zt����P��k̂�A5��E6f";�X�U���(�+�1:�X��S���^+	��V�� ֻ(��	��s�W[��+�B��7	�06���_�P�	H~P*u̗�#�]d(��ū3�t���1o+�+�pK����П�<��'�*p�O��(E9)�h�s�A���d����L6�Rs%�FEr0� y�U�Rг����W��4���W�D ���	�&ZU_�!��)�`R�\�;[{`�^�XD'Jqä�Lc����|�����Щ��a҄h�W�U~/RUŨ��έ��^uuh�R8 >p X�N�1�K���{�-��M�i��.�ݟ�.�D���U&�Ey���X�'{�ꢰ�rT\-��fS�-�l�i�:`5	)^���i�ѱ �Lh)�y���s�����J�oJ��ƛ�AsX�.ui.]0���kr��dn0�$E�,O�h&d�݇>�8�W�,��0����i_��xhtOH��o'/<Jn:�;0Z�j��e)�d
������GBw�5�I��a��0b�ȁ�k.^U��ZP�MS]x��M_~���hR�Z0U��NH���(�܉�����K&UN�F���g>��V[��f
jgF����2Ha�5:� N����%�L|%��wf0'�;_+��C����ð�[9q�R�	o�+�iӫ�� ٽkz0�� T���	/I9� �d e@z5 �1�jm )�-W8�(ͻ�REt�PI%���0b!���Wٍ����;\)�%ݺ����f�O8�@[�>cx��X4�{�������B��^)��Ѽ�,�h�h1�L�=_ 0r�~�'9ٝ�`(U���O��'�8�^���V�Y�G]O3=���*�<^�l���v9=�F|f[p`p�Ȏ�D$O�2�0�T���3.���yt|,��OUt��lD��Ų��l����0w��A�S����4) ��j��\�����&r�.1�lQ���y{�
�h3e�i ��mKC(X5�h�pE�H1�����Go7��Xߚ@h�
/U6�,���g��c|�kl:�?	�;iU���PY�IL��Lڄ�h�Xơ� ��`O.�Gr�N�lIk �|�2Z��&i\�� .V�h�r]XX�%BF��{ �QW��Jx83��j���L$H-D ��81��Qt����a��Y݃fR�T�-T�2���X(P�� ^�нq"�!E�29,���~�v�%Ha˭�)�O��N���F^�2k���:�H��!�Y��Z�q� )ȹ�8M?�Oma�;�|�*a��2����@�������W��:��՟ �L?(Yh����A�I�cz����4䘗H*l��O�pc�	��I�j��X������_P�Nr�_$s1[YV	:s	-:��N����n�����>R	^8��.��|Ǡ��J-���G�N�(��X�ly��X
4������-roFb2*���	���Pִ��IwqKp�^ R�i)�_�k�\E��`����	�fb��M�h�:�r�T�EUh1���^3l�J��S1�Z[R%�Ȁ�0d����#�N�:aj��������1Ӑ���z��ӿ������R�h:�H�V�@�)�Lp$:˝��1��'��p�|J�h� �(Cw�To\��[O�>�nB铼���Qd$�VA���p��N���haC마�L& ���o��Y[G���P���C��6��s�
/Pԩ@-�2`u>u4?�/ ���! ��1'@���{&7G�$�/ωx�̓����U%l!\F�@hˇ��:���h<~l�$�[f<�����e��#q (8�\_�'4�qt��Ѫ4D�%�^��L��1�"�@\�Ю7~��8��>�X(�cBW�y�)C� ����[���'x�� ��k"l�iA������ x��[}�H.��ـɻE1T��H���h#^j/�>���d��l��FCs.4���;�8�ȮԘ�۷2,�A�=<�韔�����J�8s|�u���������%k�8�#���޸���#;n�	�:�����{��)�e �h�x�������ق>_�P_�5��{�Lم/�����8A}�@�����hSz�+kN��j8��h���#�D�6kzUe���E:^(�֥p������' �9���_�(�_���xe%�����aq@��^S ��(q��N �-�j�k�O'���9�_��,�twlk���"h��\��뇮S�0�	~=A/���m@������
W#b5�a�ǆ��3��=03��1�|�1VT��^��/k��.���	#c�eVy��(;W�u���~�$�*�?/��	�Gg ]l%�0|&|U��e�����"#��8+��է�0�ƃ{?��`�������R�9��9*��Ze	�(�ZxR��9�7�2���=����0.:ch�Nv�'�
i.?--^Z�09]lS�� swDB���|%JR�����i�?�	�)�>�����/���P�c�x��0�ױ&/�����1�Q,0�� _a�kj$M���A��io91B���1�^�0�-i �')ؽCo Zz�N�M����D&���{�sVQ} �F�J��N �`}U1�X8�Ѷ��Ո߷��[��@��Y�,�����Ϥ�Q�Av��8�gd�/�P� 鼘����k��_�_)S��Vu+vK�.�x��[�,O�)k'�E)Y	tŹc	�k�}Ι�RE�'0�w� Qh�$e/XPb���@A��;�A.��0?]DP3�B���Ѝ|6�u���#��/	��H��0�%:�bV�}���+���	�7%�	4������0s�3>�j-�7�׃���|��u�7!�O���W������K$]M ��z!�H[P� r�@{�q�- X(:�S|�{D�u�{�[��X/Y�D�#c��^h�MX��_!򗖿^R�}Hd��`����J�b��A-��ݒ�AU6>��. X�'WD4̢��f���J���^)���hA����م�]��W�wy40����,Y�UM0�<IW��<��X^,>�'�{q��T��l!1��P[���q�^�"��]z�c��[��4`(E�r����Q�'P )j�7���(3�-�������'�<Ъi�^E�(3���.X��"��ծ�1��Y��נ���ױ�<��7G��<o����Cw�j�p$@��g�����H cq�X-�k#�f���1��%����:d�C'��*p(X�l{1�"�=�b��3K��@|�0^=��I�8$�hi;�˄&w)i��E(��(�ᚽr!%b��9�6/Z�=Y-N�Auq��-2=�K���on�HW� �6�c���'�X�Yo�#=��]u��}){z�^`4 ���S�����)Ё�Fd�H-	q%�p��z�'�w����*�'�~�|�1�����4rr�-ud(�ۀ-���~��קܳNv�:)��!�ZIY��ri>�A_]���M�O�;6����Hv�Mo����� ��t�H�Z��*be"�+]@x����$|3���v[:��[!)(�p�x�;)ͭ6s��9?P�@P)/�[d��t	,�-X���}�%Q�T�@��@KC:� q�-�����`2�j�o���(����	�>�x[k9 �P��Z�s��YQhbyw,��%�|��w��̐=�ڈ�l	��f���b@��X}[d�)��	a�x��e��뼛����:E�+�Sip�PhoZ�=_�6u��b�t��s���Xx�a� ���R�����{9?�g�Z �<(���0�髏v�it�%��X��	"��Q�J�oQ��9�߭4�$`��,�~�zIQw5�
X���G>��I�����b�E(b3BmUA�5�C�[)�V����h�:��N_1�.�^��3eK+Y �-@{V��l�T�,>�,�?�й8!gK��p�S���6F)�kA��~�|�꣋�_s��t�XSh
	EP� @Jn���	�{�P����yN
��c�|qU�98+p͌@�ܳ��I�d,Ĕ=�����bi�rC�vH�Ll\2{�|M�t�J��f~¯��}���-k������U��� ��!i�TU���4�r�DG�K�@���P����z�?	�����p3����h:������:��Qb[Phuz/d �O�YM�9@�z���'�{04��
3����`�i|2'�e4ʵ ��/���4���k�=����P��A�ǐ���.CKU��+�p�a@�z�!}%ù�vQ(�B���;�ȭa:���r�F�JX  A(|��2�#���z�� ;���$!OS{v�������P�6;������n�9v\��L(���� ���i���oB���_v=)���b� HIF+-����|�M�vY�`1XY�L#w(����9 �P��	�q�u�:f}^�L[��7^���:�T-2yFm!�:L�@Qh	vX�B��k%�7~T?�f/�!'S�y��>@K9#�Og��*=(u��8h�D�p��*�Y��`P�e���1�XSW�O� ��3���H��B�D�����\3T��Ţ��p.)�^����8�ǖ>��]KSR��H�H���M\;m��NKv��f�>�@��˫5)�-�%L�ոYWr�-�~�=����E�bNOE}��Y>o=�/eb�S�K�"�B���$#[%�>V(��/�<dqZY��Ɇ�>U���VV��A�[�>�*�����ޯih;��$�Q4>��A @-X]�+�TqM�G)�+�giP*��u�l~�3��`W �1�!�P�%H� �y)`@�N'�>�/���N����y0��
1^�e����,-��WV46Wf�sP�h-BX|r��Y����������9�~�w�	.�(5�#_����!�^5 S�A���T ��dB|�3�a�~����?�;{
�\K�~ƗA_������Ɓ�F��*�j��_�jA-��I��]��'�'jS��F���$�@��!�1�~��_�H�(�he)��@�P��i �F�s4�/^� TH�i[�{g6R��$_	 �,�u!�h2[�v �Wto��QҪ |{>h*�[-��`��ِn$}K`����%	J�X�����V�2(C?�KYh5��T
S� bk8��wOA��	��PG�o��00��Vt��UKuEu'W�4�Tu�����C�S �LZ���ЧS7*@It	A��m�d��p/rq�3��	��z�H䮩/��@�m2S��A+���.��IO��V�("�7?�U��
A1����������\?���68$�a��0��j��s���<J
����Ɂ�A}g����T�ad���Bh�n8�NF����k�z�@��N-l5�$%g�w�r�Q�,������Q����%`؏��(<�'p�&�'Y`�X1�.���L�V�5�	p�RyV��8��}��A���(^? C9U,�5�1�G�Q���\^P���"��g'ZX��^b\J�E�w�� G�B�)��O2�j*�r?U����9
�C�$��):!��Txo�W�9E]�Z�·d_���^M\�!R�+���bV�0���Nݠ���Z�=�� =w��%r:��e=�?t�����4 �-�x�>�_l�ŵxs'Y[nUXV�pPh^Kv=ؓ�7���ZIK�ȷ��^�u��')�j*qS,	�`.��bễ�����q�h�S�-`S���^�6/��D�����3j�Cx,��rUE�i���{�I��%^x}PhUY�X�l��C�@��, �o��' #�U��!r 5�YoJ��O%�?
��T.<Xno_R�1�V} 5lP4-�����.�0Z����sW��!�E1�_�]5ryz���� �+"$�MR�6lY��E��B���@��z�I%�n���q����dM� ۽�L�&�Hr�O��4yf�;6a��C�j���r(�L~p��q;dO��E�Nh�8͍x�\�9`�?�/~��a�')�Z�~7iWwBp�Gq���|zP�)d4l����K�}��U�&^_�����p��eJ�g�Q�`1�y�|��I���MA��(�3��?%S�F)÷�J>�2����R����U�A'm���C��HK֪�0 @�jr)����i}Y���Z�!NB��U���"HOX��N?6B�+p�X�0|I7�]��#�fhCj�u8�[�H�-�h8{)Z�,��0A�4���L,��.80ڶ��	F��x$ӊ��J��D��z �W�t� A��|e@�'wF�Tx>��s�wb �	 B��)��r��J�Ö�ɐ,(�������^hb@�:M��\�r�,�Q�%�1 ���|Z	u<g?t�°���?b�aF���g�m]�ζS���á��r[�f����&5u��E��(�z�V�Tg�� ^�J"����E[Q��`գn)H����T>����]`'�BFU�LPh�H*E���)e�{�����D�����F��E*h�p�3�`�J�a����j����,#U��<�$xޟ�霔���EZV$��J�(l�2 Z#1�D(�0V�'0�q[��G
P�D{U�� �D��1�Y?���!�]�+�x=d�Z�-G/�A_�B��@
�<�'�X�!�H˽/X�[q{�#�\�(4�v��Q�s��]��Tb�h`�~J�$�¡5`���c��G�y�9uzR/�w)�}��	(Kx��3��	z_~%���O~��EU��L�p���nF�5��y�>)��U-D_Xt!�hQ��	�G4�F S�~��w�ߝ��9̽/�"��7_�/��~�Q�:ǳ���oo����i�߻J�y��� �oS��y�ʲR�mBBŐA�6*@���%ɉQ��n_�`���y��S%�q�C�EpG�R��o�[XfϠ�L��o@�(� ��� J�'5~�5����/�� l��G�|!��kd:~F�o�i�P�@ ��_���d(Jh)dm`�<z%PTY��5/�lJ��׎�/9� ����^t��_a\|n-�AֵE�2��鯻 �fS�������[� ����,�m$�m`*a��Z��!�XBA�Ɏ�� ZY�\ #�/�,��E�;�'�Y�vZ6�u���Rw�vR���������A��S/���
n�F������;p��a�����H�u�a�xd6��L���������:>�E��!�z��	��wl�NZ�C��2Vh�HB�H�^U��,�J�����О��YH��&�.%����R���4<%�G�G܈�`�%u�:Eb�W�p�im�V	޳Wy:�C&� �T]kN��KU\W��LGf[�v�!�[U�l�5q�tV򼘴�d�!|:<=�;1��1�`ch�]ΐ�9 ��%� �}'4L��c�8 xIA���-�v%�Dw�f��'��Y��-)`��EP@����o�g�(����\��an7 c+)W��t~��3�q�}���ʙ�`8��<��\o�KZ�hg�`�]�Ru[x??2�� 5�@JF�h�2��>�Vs������i�z�P�k�����a8�k���^$�O�PRPh�$,|�6���g�A�[o�f�����p!bk��K]t,��dF|X6�?����������R�E�����������{���S-Fb�U`���h ��}X�	S�T�k� �96A��.5�c]v@|7aC-
�o��>Q��0X�4G<��;ُ_�'v�Ɋ��?ΘOU�Ok�"GLbP	{E�ޅ�	[�b�W֯`��_��KX0�~dE��rR}qi� �gW�!��L�%����s][�V��uV�`hC'/HXT� �F\�&�-�i=2^
�7t�[��E,r���beA�0���(K��a19bd)�h�REH|�D�v��8a��Z��QK��tÕ��.�'<�U"/�.e�_����;�1X�$��\�5�(z�I�WȾ�9����y	 �{���;,�A-3�cz���Q 
U�B�/��sE �0�hw{Ĺ��Ĭ�ą����y0�|ht[��u������c�K�����EO���s*�Š��U�&��o�|�ʎЈ�6�h��(�4��0��R�n����¡��b���F����߁����^ !�Y-Tjy~e2��1�^M���	8�_^�L�����!��� ���`2�yHi9�����������c��,`�Е/)�|Xb �`�LM%�>v�H*��V�r@F�=J��1��D��9���YR���Z��Z��P���D`���a��y�Y�VQ�����!�����F�k�̖��'3���B�(�,����ÈH8�K�9���S.X1K �"e�j-�k�(�%x|��錻���5��Q�>�	�	����%����_)~�,��r��~��/56 d
�`��-:)�Y�G��DX/����~C����)�`�@�1ݽ�Q��/���y^�_N��+	j��p�_�c��Z��=�ى?�1�R]��'���C��������,*�C�Ŋ���36�+��,��E�����Q�0��9dz.n� V��`- NF���G�.�b����~�e{JȪ���&��a��8�bjв�Fk�Q���!Z���h� ���=1��CS�4��U쿸� ���o��N/���K���� a3�?����)X�-y8d�YV3?�ǯ�zH�rĬ
[����^�8by�%���B/ZXw�6��L2Zf�-��U<���_1����XC=�[�a�F�>����o?8r\[�	�����4.���E�:�b��"|�<��Q>��DI�[��9�05����d���A1l��ʀiC�k�a�61�Z�=^K�g��'�Ag��3v:���Wl��n�eG��bVx�PF/�	�%Y�[,���R��,�(��Z0ð�֍5�� �fZ����\��g���j���S��p��2��('wy�kΧD+���u�Pz٢�'�)_B���ev5!��H�N��Uj��w�s��*.4P����[~���DBfO��#�
[KQ/;��:@�,��k�} �0�=S�u���lT������,�Cj�4�마O�]_�f^��QJ���'Ft��f[(��ڮ�,.�/�m�1�V�7'(�ղ!��[z�f��N-�Da4/�M<{��p;pP*˘e>)ޮ�MA|,�h^
�'"���)��\������Q������0I�[���K�U�HX'O7�V��\9�� �B%�ｅ�k���j�>�X���&(p	fP�A����)ָ���|P��:?���Y���C)IGz�
�?{3ˬ��#'f ��.�Z\K�ݜ�8���>B��!8��N�H�B	���޽��ႅ�u1���� �d��ϟ��-�A�s����ݝ��B�{�-b�x̀�\x�@!��+gT��_-�FRW��v�/�Th	���o���@�E V�oga1+��;�����%����J��<�S�hi�$������<X�
,���d49�~�XK��ߡڶ����t�?B�v6���C��T�8���˄q����x{�W���a]Rff5_��-�?�u��i 1<�� P�5�
�_�N��Oi���$V�3��TUܯ�]K�j�����ou�<Z����U��i%'rcj�	_����'R�*�0�� }l��7�q�0.�N��S��������&P�胙9!�2���O�Lafֶ�堽fNh�s���@��q�`��^�/V�������D}��R��fh��� ʖ��"�y��b*1�Ǎ��~� �D�X@��l�0�-�]b(أ2)��!�1�Q��BA��jA ŃRH��� L=�0sH�@��[�/1�����A��ͳ}
�fB�RP~��X�ZU$
-%�.���e�~���$�t鋜�6��R/w��H�h�}L%]J3@")������u�~�H)ؿ�0v��-�e�
Й���������N�B�����U�V�����pO&��$�)P]@J�2� P��v[2�&j\W���Y/t���S�o-�U؋ ��H�)1�_�^�J6��S��	����[n�Zk�)bZ��<�u'��U� ���p�^�"�#�H��W�� 0��HG >J��$5A3KC9�Q+a�M��%>�2�.���{�G�9���^� h�nY� Ẁ�z���h^��1��զ����4�h��I���?s<IX ��dW��9]!������X�kI�f��<C9��A-�OHAj)�B#��v˟xv�����o����	-��Z�l/ �y���6[�o.�,�\���X�L��S���^�'�j�*:'�1�@��>���X���\���~3��0?>R+B*�64������kd��9(|��x��H(���z#P�%t~ �	�c�8�h'�3zs/m��S�&J���������	����E����]O
�s�0��Q]����[v�����]y�B}�fH���Z*6�W|4���ׅ���^V��y.w ���Z1�)��]�{��n	��~�������Hg81�^�Ps�(K� Q�2b%��j���Nڂ��?��u�}:�Y6��fc�q��^�J `"����'��W�D��I�{�z�_�֌���@�S$���1����p����Q����d��Wh�o�G��'��~��[��D/1ͼm� ?L"d�3�Ռ��u}N1��Z�E;�������b��R�Z��-�P`�ʥe�-�� /��B2T=}@��N�ʁ��^	��Ɨ6iYt������w� ���A��qL>� ��Z��-�_��xfK,#jM��������	)�[U���{|� �-�@��U�\�xR��:�~�F�W �ʟս�3�"�t*�/�O�k��.3d)���-��&(�ti�9o�
`�!�`"�v/1{�c���U���	: �Z�vi]��N�4�X���~��Â�~��6nk>EKyV�T[�^�iOD�j]'+��߆�h������D �v� �9-���/,msJ�'*+�P�#UP[��f�g��k�)���H��1@��>3Fo���_��Z	�`�}�! �(��+à,h�UzO;��RY����tҰ��TcϦoD��q	��pK�W��[_� G�-5������/�; �(�0�hQ�/�v�	�2�`���Ws�(h�,J�t=0I�J��!�'��%סk��$��p��<��+�@K��^�yqB��|���+�P��V8xd���YS�A�k�	N�*�%:�]����^�a ����m�wQ}��������YX[6LR�3����A�t)��[颮C2�QhU`�g�<n~"Baw��R��>�����YW�#}������Wa�&*�!�������p�^'Civ��B+�����P^�\�Z (d5�A�h��&�`wM��aʔկ���JUM�*�� :�f殢 -$�r�HwɕpY�Z �|�vV9���e��C�Ԟ}1J�� ����$K�s9� Xh�au���d�#D�l�Z$��
��m+� ��<�D��2�lC��]��^)U��s�~t��b��A�x�?�M�Rn�,XH��'�^#�h�`&Z���<j@�R�'*}�/����l�7',=���?�%[xq)C���'��@��ϵ	�5~��p��.,TN���2?'/<���>�^ISLu �).Y���e��������;�����uBw�Dn����\�|�
�>t����+~�I�AV C�F[�P��*4������vw;�Qx��!Z�V��B�����@�lH)�����h�S�T��*6\1�["b]`�?{��e>�I��c*�9z��e��yK_������qN��!�U{�%�'�_x$���պz`�n��v�%�u�$��K���b�W�m��5�	I�D%6wN�;���x�Rhs�`Z�y~/�xU��	%d��K]���d�����(��1�50]#o!��TI(OJ�`~8��@���@�e��C'B7@	y  r�t��'�{��0�qǐ���Ϙ��?���8���g������<��7&��CoNqs��B�C��p=�˓��r�^�=s����U��T���'T�`�M}xV�Ub�m�غc�R Y|�YJ�f��'$F̽~ YS0}�4; kJ2os�0'K�AE �z\H�<ub	KiZq�u8�<Ȏ�1�NӋ�}O'�:�Z[�xR H��m��!�1��K'�� A)ݹ�0��/��4�D��p�P]��I�#���/fN(�hD��O,���y�Uj�v��FĜХV�	TE|fh����X���bP�K�P1
Zo,�� �N%o83{�?u5��	(�C���Be~б���﶐��}���U?��M�
L�; )��Au��!�e�� V�q�IZ(���W�⇮d��v���1����p��"\@G!��1���'�pȱ�=>�-��_&�>���-[XMP�K���F��hTp[u�e&i�g_}?�w�����<�ù�Э�W�{V,��r�[خ2P�U��]O ��"�Y���� +� 1o��-G��K���9�3/�4��~hD����^�h��;t����iu?0J��+)ˇ��P4 ����]L��N
�Z�B����W�I�R�4$���%�LMu��H��W�{c%��`�V����X
g03K$�~	#YǙ?�ML �B� �%�3+do�G�i��pc]r�a�$'���i1��	^�_���f݄]| �]3Y�� ��!�J���U��_�X��h���X��N���r%, �<ߕ�0�)��zg�H��:�����ҋ��ȱ������b�|�@��= |��{�,�&�S��YB�w ���@�UԜ�}`>�*dY��_�瀻�6���%�Fl�����Z���Z��P5a&.�QQ�H��v����ﱍ���{�>�\p�� �� �7�JK�OR����<��)��5ST��vZv+�U��1б鶧�p�)��q}&�	]澑�Z� ��J(�0|�*����#�g�ã��$�+��:nz�+�������Yy< �� ��!�1�	�{��@�S�`f`�`�m��$�,�	Aoc~��p���B�Y�-g��� f,>�۸dL����wԖ X-Az�G!��%i:�	�@�"u��y�q,�[P�~%���F�M5�2�� ��������C���bx�Y��Wŕ��W��J�� )�/(Q �_j(�Ww���#1}�7O�K�Ɍ��,�4��kK_� <|�O^  V�ytu[�Xٕ�` �	.�Eh�Mw� z�,D���1��:�)D�-�R\�vH6{%���E�3�ê«(��qz��F��GST�U��E���&��<��{�;4(�lT� �[�b��|@v�נY���  �Sh�4y7X�Q-�ldEvJ O�+5�Xz [����%P��9��Wv�%�e�<��,�J&� 7�4ERdmx���ZAs�����0�!�]0�7 D��B�9|��9'��.�ܭ���,U	��B�s	�=W�: �r_��7nWB�\��w�ח3�d�ia!�XF�VX�mCP�ӥ���PŚ�z^.�X@�\*�W�_� � ����� 5Z�zX�%%�T�W-W�&<!IW �U��ߨ]A;~��w�U�v�Q�0��hl?y��cT��v���;p%��@5e[Aa�it��ѽ�}.��hv[�99π�25�aN&��	u~��T�0��S�A�3���#�L��b�t�/T��H�cYe�.w��X�����+	�#v�S��1X�O@@�|zWYaX�U]n� ��>�HF}-��kըB&K�jr�&�x!�gxE��o�~#���z��r���.��<=T=B�Q`$ט�A?�^��w6G0kt@1�_'����f�A/T��J~>���-D���U��Z���pfQ������Y��r�� ��E&E� �CQ��Kz1�B���WQ�Ä�.Dr?��vt�H���1�)�=�+�j�u��	O�^r�l
��>lI(!�<���9x���	.Z�\t�x6-�Cx!��)� �{H�B��(�P�^	��e��\�^��H���e�����L_3�}I�J�R�����; ���%ޔ���K�)J��}!;D�����!i�_/�*���o������v�Z��`0�(���P����f���X��S�v���ŵt�xB�N?��ר���h �0���`����
��.v ����:"ZJT���f��3a����/@�Rnc�{F% _q�G���4�dP V�d�����U ���ΑN��f���A� -�6)H@s!m>5��!��G�Yr���wo���1xzq�{ �P��l����J9�q)*������~A�~[�B*��}44�&�ϩ��(Լ�S�A�,�z�p�½�
�Z��Z}zL0�[�<0�lJ.GO`}E�f�1���C˷'�O6���IS��-[����9h�|DpyQ�DY�*�&z�*��C�[�Y��XLy����!�.� ��
)��C�J����%Z�k�u�ͮjfN����1�@��~{�`���im�b]V;�����J�F_��cczE�ZJ�.�( #؉���������.~)	;�O?�_�5]*�:Q� � e-�������?z�'A�1Aߧv��_��U����B��V�x,+Oa�Rޗ���J@;��*�tR��������ى��W0���#i$�h�3�;\�=*�*���{��@�8�|�V ��e��	%�f��15�Q��6|�fVX�	L�SGj�J�IE�EQ��,��� <�?U�Y)�>I��W�%��7I��%{u�^��=�Pnbil���h>\*�?F]M���7�E m�N5�?�-}��Ӏ�%�1���IՁ����~ĥE��ҷ��P!���[Q�K Y��j^�e	
����)W�U_QI2��́��nGY*�9�2H^iwC ���4��-�lPo��A{83�?�h�T`3Y�*��k���L+��~1/����hs@^`��B�3�ր�,�O�c'��G\2�Oa�9� ���{��7M�eVUK�.��̠?]�%+|���[B�����HM45�O2�i�^P��@�X��|�M��<�(�xZ�~��x{	h�8慺~�ݗw��]�P_�=�H��׎1�Am�ȓZ[�Ag#2b01���د@�unI-�o:�j1�y0G�/]2����U��zd$��� _U�*V	a)�]����|��O$hy�1�E*�0 �h}� o$�2j"P4� ^v�	-%O��*DF����je��Y�x`1Pa��v���ꀪ�E�Am@<�t�]� 
ZV�R�!���Fp2����h�|�z��I2�r��d}.��}���l�A�:��ew�.q�BaLb�AN*��E(�Y-f��.��k�$�̬�^�R�#T�@��T'x��`e#�M� ����`t�Ũ��!��i1f����4�;R���'*�M��C��!�>�0��/������L+%���i���4�e�=@N�D��K�6h�>��^RV-/��Ot!����j�K,��I���Z��ы�E�������j/���TM��
��8-�^�h��� WhfN� �`���%������L-�c�d����%��Y_)gA?�X�� �	Ü�����+��f�H�W7�+ �S�ŕХ�[R� 0�Z ��8���"��SҸ�<�Ҏ�OTiw���W�{���U�����O�%��]�N�%����S�ep�*.�Ycư��� Iz�N-��Kg5���1¬����؉�_�l�� ��5�X��,
�8Xl�X�-� �߉���y�r/�_�d�����ţ�X>�PE�a6�j�!�]0�[��_o)����H�>fv�-Gס݄�I�>hy>C�[��,��BsJI��
1���K�j��[�>+V4\]�+�����Ē������*�l��[��c���p�T�X%�p����V�Z�Xȝ]���H�~t4��B��~$z@�\S���HY�K7%���KW�t��a��O�u�^s� ��u�qk�x�0����A
<2��ʕ����d`�ʞ Q���|b?�qk�����;^[&k�2�B}eRbDeh/���V \[�7X�NLHy0��X_1ڷ�Q����~��L�$_V�<8DQz� p�6���+��o�T��������{�Ű1��F��m��s��E�� ڻTvs<�؀�!����VXtG��]ٺ��g��^(V��%U�'�]���rf�WV�:s_��댚�Ģ�Ӵ-�C?`j�J��f�)�B�����ʵ�r�
:�N]�)F�RDTHW9��Z� )SL���_����_�;/�8"��Џw����.��n��~BV$��d�j�����aTK��a�hCb�Wv�rN� QhcA2:�&ee�8P;gTd)�s	'Hy7�n���ɍh�^�L��~�������cɗ �Ո�Y��������vo�C�d)œ� �1�h�UMA��2Sv�&���j�A �1��W��\�V-&j����
�/45��ѽ�[׼��4wJU/jEz��06kR��\�-/���=0u;�rN��T�Ρ�?����ߧ�/ԟ�c�^��w��*�B:�a>w�WaED�X�@�/0�=�G)|��@_���;&S9T;���5{ꗈ-'��ND�X�{W�"��-	?D���+�q QW��`�H�e<�^�qDH_�q���,Cc��?�;ˢ.�K���|�4��H8�%Qa���V��3����.�&���û���l�g~v�*F%3-���W�9-}��X�)������,�y>G��)`��ҶA�!~.� ��
����R�-'7��
�#=�q�9�%^�tW���������R �|Q�n�`�P�/�G醇`.t3�~���|	,��?�f`�B����ܡ�>�2�eb��8C0"��' �Q�ah5oL��(�'(��)?zT[:�
�� �Z���3*g���f�>�Z�)��τ��𡶐ۻA�T�D���aIE�.	@;�#_�y4���Vߝx-r�fI_Z.���'���\M�y9=!p�P	{W��)�	��A��ڽ�Jn�` �@�"�Oj�ǻ �Gx3DM �5&� 阩���4β,��������K�b\� �k�|��0"3M�l�Չ	���]�H��Ps�$W�4�|=�/���WW�
�=�R)ý0|z�wEM�H/�4$r.0z�Iٸ�%�?y� R�+tP��v7zؾ�eK��&���;��F�r���P��(�X�6��2���p�J}�p�fL{[�����Q�M	1�)�� ��,#\~��B'�s����uF\p�r��
�Rr��Tw�L< ��\sP�/Y�����h�f��@�fM+��&{��ib���8	�q�A�3E���w��k��u�a�z
����̦�̄
{/|���r	̐	��a��bD�g�������.��ý�b�"�Cv~%8Bp����_�L�I}�>߸U%}3i�в���?���.9��8���!Y���ⵒрp�/�ɘ�!��d��Q8��1�H�>�R/t��-�J�x�ΗbP�9K��6N���-�F�J �VW�aU��:�+��)	��h��;�~/\!Ӿ�{��<J5o�A��SD��P�4^#Uh�$L�%!�����Y��-�?���i�p��ˀ
D4	!�[Wit:u�?ũ��ł'�0�3����_f8�,+�G f��%oߠ=\�.��P���C.`!�J�J�;��&�}!-�f�I��d(���~i��\�ŋ�'����B��qn��J�؀�[��, ��R�hn��!Kjꐛ�����í;A���r~[��F��'R�'�]`�����0��b��F,�0!.rJB1e*�@�g��[%f����O=-y�P j�T'�`71JX��$!iz�3ruJY���]�	m�,v5 �v /�7-���S��?���[�r� �sRdʘ=�%y|iN-0슘��E -?�]k��	f:9��'�\%��hOP�	��VI��I��݈�f[�f�PVв�W R��#�p�=]ڨ)˿��CQ�1'
�J��h~G'u8/�Qd$�&�X�������n��L=7{l>N۹�ԥ.��A/i+�j�=-�7܂b�}T�hL8��� Ke"`-�g,/(�>Q���,A�	�.�(�[��ߕ���U:�6ym����ɂ;5�	�~J�Q@J:8��x<�}߀׹_Y�AI�����E��N�2��D1�=h8+����I]t�P��n�U��1Ƞ�q^?'3� �iF����̴p;�/z�0M��K�t쀐��p����YTl��)�KX� ���>cN����Ɍ�޽-^Z�h7UF!��$�@ ,�����^�r(����0��Z$�� �+?~f�������Av�')�R����p�1)Y�b�.ηQhSG�_:�W/����E@�sw��%$�#��,���B���;�ʖ�����#�t}� �(��k�@�^�)�i&[��,�WL��V+����y���ZY�pO�N��#i2>xM�9YC �aʆ��%�~,'ԕa�z�x���ԙ�g���z�J��d[w0>�#XM]�7��P�[��L`�qN!Gw"+@R�y1Kݻ@����!	��'��OP�Ptv�^*A�0� <1ZѼ���%�_��$;T��R��3נL7�{��w��>x8���5*2��Kl�O���䮕0����H�RZ%)��^�p\f/@e��Y�����i���j�Z}�-���Q�J����V�c��*x)�
i�R�0g�[,�'`�ş�k���g�h�b�:����g�Ra"x��y���R�%��T��^vt��^��!-e��������
�;^���j0��4����
]XWz_:*����TZr����w�Ղ�p�b���`���`,<[F�:����=^�����$ �!ָ�Y]��XW�	^]ы��ѫ �v3=,Q�f�h�L]x����3A��Z�f����d�l�X����-��n�N�-sk�qB[#�)�M������I >�Q��0�قf���0[���\�(����$Ѫ�}�,��<�[����۾[�Fj~l<����Uz��2pD� "Pp�4iӌ�cw��;}v�|\S��X�-�շнR����^�,<�_Mm�`Y�NM ��jq���H�]Y�c�����t�k�i�@��~�n�%��Y��*������֨A� �<i�	D  �9���z�H!�.�q��Q�]/Ĥ�WȀ�L�q	l��.`e*��6�7[��DP룰�mvA[+�� 2
Z��aS�� ���<fh�\�?�[�*�׼�Z���ꬴ��h�,�Lu	��#�|�a�*����5jyK|�Rz�
_�{8��'��,��P�Y?���H %:gAz5	�E>�����n��:�S�h��%�(����lJN��P� xB�:��ZH-�A�*�R���1��`
\�g~V>F'�� �����*%�fI�:�k~��GY?����W��!�<%�UA� o2MA��Ä�a����E4?�͂5��FTK ���K5���ʍ呌h�z�l���� �2�-(п���@n��I8Q� kG-g� �)�Xh$��`q���0�r-�FE� Wh�w���? 9�}��
/�����l!}��*�/���=5Zl��_U�'{�2~oZ����A3~�iӸ%!TT�1$�?Z5��V~� Chu8-;[K`� �`$t@��
����FJ	m�c�3�_$[)O��Z^�*�	h�=�L�Bv��ï�����'����h���5�p���1	8uY-v�w�H�Kubg](|ɉ^ �P�n�c�
&�����#~{_uI�u�(�pӊS@��%�}�llI,�tZi�`�9{�J�
�K��5XD%��h�[-+_ZJ	J�%۵��KQƽ.���p�OS��p�j�@Rh*��'��aP�)J���CJ��9N	o�Tj'N������c�5CX�
��h')	{Z�I'z�;�G )�Ph�Y%�l�� �r	N����q.��`�"�
8.�r �\�cNOp�����AɜH�E������r�9B�T�vU.t�@�z��6��r$�p
@�7��t��|3�q����������[\�k�*��Oؠ[h�v����Fz^w�ڲ	�����
�_���w��S�)�#��g؎��тJ]�DQ��Q_oҴw@��'C\`��x0!<>�����bX�X`-�l���T�q0�2-(�:�P������avJp�`q����t�����(�Z �[RV ��{4a�	|�
)�^}�a�ad6`*Ֆ����o,�jt�\/�=a�" Ռ�HO�)�O�� ~�2L`�iz�OL4�YV� �����\yX.5r��P��`�%��u���q���7����>{^�\�0�dJi��s��i@,gi�^r����$�	�>'u����hR���ǉ�U��0�m��	�ZV߂��T�V�f.�)	�!�[]8J����+�Q�C��P���Q����
1��K���y42��_0ߠ:O�G�٤N�������h!u�_�<�/�\p蜂`�
'y8}�� [�K1�%����{���i������6�-���٭[):@X/��Wd�ծ�dS�ZL ��v�ʷ��'�RM����A��$	h�y����%�u�����,�R'�g�V݉_m�s�!�K_�S�ĉw!�,�D���OH`酆d�ˮ�j �MR�%tO(��-��f@H�B���ޘ���i=�}s��2�ff�zTk����):���0��3�"�������TE	t�9o�0Ms��!Fd��a1 ��+F�5�����W/��g 8SAm�z�S��K�S
�	���
�i��zE�:�(���+DO�1�h�!z��1��ĸ;�'M����+�M�b,�BߩZw��{0!��[�1��8g>�3�i��vh�'�O�<U��b�)~���^A��o�͈��KX��h~�%�Q����f�p�'�%��Kשd��	���70mX5�,(�zl��N7�U�B�4W��������ؤ�l�\�p�H��a�W`X(d\��a!�ts]��fz�q�iq����8
?��фD��4�2�7��Oc�!�-�K� x�Sv�q�']�%5�H�ZY]<�%�� ��\2.z.]t��f��ڄ.Wۗ�	�_h[��2�`�E�fR������s�����b=,�RS^��0Gp%�*h'�%v� ��3�Kj��KR���5^]�BQzFk�'�G�З�H�t�T�i/�oE����[��� �;���x���0B�0$mY�r.X��Y���c0������]h&�ZHR`�!n%N	��J�pK��A�30k9�Eă���j�]�.e%D)|���YIS�P��}v�%�qh�>�(����d��He# S�� �Z��z����;���
��3�Q%���thL�k��>z�q	�&�`f �!�h�w��'G�b=} ǯN�I�<|G����@`κ�>c?|�^���ѹ�Q�!�.�� mkEn��$�\	ChWG�R�X닡��Q�Wބ��y�} ODڕ XW$�Y���(%	8V�,�]�随���2%o��9��^�i�������e�\!��D%kX�]H �a�J���0d�&�[�sO]0�uF}�� �5	�M�1�����_������j�.���dQ��3[*p�-�4
�/�7��ݺ����EHKl�vx�ZU��9C,�:
��OH�)��(⍗�2}���C��(`%���,}$b3X���.~�s��½�éї`�3\��<Ao��c=]���<qD��(9�2��,�h�f�Y�5����hs*U)�1&�~W	�U�����2�O��ӧ�ݺ"�����Ya���9�B\q��KX�)�N^�0$�h-�TzY�!>k�&�_z���������紓�՗y�l�\k����-�0��A\2��G���^k-1j�"/^�yP{���`��P�s����_3z.�����l>V����xc�r��o�5
)�At `�lMw(L&�Ǟ�p0ʀӂh����"~�w^���)uT�p�i�� ��pb��T�:z�}���i�1��kI�T$�����)�d`�*�'鲊Ѓl�r�c��=�C�J�Ob� �n�p�(w�&��t,�-�t�f]�0|��X�-�(��PF&���?�l}{�2�_l#��Մh��8o}��y�BY�̢�h|F5��[���Y`���L�;��-~@�^x���V1�F0	S�U� Mb���X��8$Pi ��J�C��BA�Y�b�\�6�r��.nV^V �)Ƚ�*0�^V�����{�+mE�W 
���ص ��]i�����	���
�S�B���@� �Q	}fC( U�8�N���(� �d!�;��J����J�E�{&kl�˼[�Y�&��ZK��R��H�$.E����6�,��zG��(�@�zM���V�P��X��}��&�W���P^Z�V{�����F�: ��@/UQ�0�]2��ht�aJ�H7�����V���a5 ��$V���1�^0˽M���(�4!�h0�����H�lN��҈� �]M�WuJ���������J1�)&d
���^Qh<X37�U�J�\V��!�r��* �և��`,�
�:�H͐�|)�)��P�'�ɴm���-�; �X3����5�d����&�������N�������wnx�~��pu]C���
�B�����'8�"����o�t�h�X x`K�!1U�	 PC.=X�P�]���o�})#���S_�Hs%�6�%7V��x��cQw�Q��5/�����J-X2W T�o��I���z�1�J��GE!�)n6�L�XϨK	.��PV� &�Pwx_Q�*�@`/�!y]��	�4��u'���&�����ؽ-�c@���A%�3�G��!��q��{����/����Hq���Yh�5�H*�@�/���_H��O����k+6��wP�V����=,oU� �v�(�����P����,�]�nlV g�4�a��h�6�d�-�:�o����0]�Xu�gv-J�߷�.޹+B���5	�\g�}�Y
Q���-��Vos*�[������{UL� a	�9�<��M/�.)��J����f�b�t�%1�[�T�" �g�-��k��c8[1�z��=;YN��A�Qi����@��%���P	ٟ{��__�$QP����XR�����,6]��AZ�
+ E%^<S�]�5@�w�W�����J%a%1��i6B��&��.��*�r�a�ܟ�hh�R j:3-�iVC;Ç�4���,Z.!�ܿ@x��Y)�]�wHn|���W��[̒�Z�(?9���c��+$�B:� L�%���'	
q0�G$@�	l��L�	�V�����L����!���Sp"��/C�������\4v)L�7vSU�	�س\��o�	ȃ��j�4�'3�À�A�����A5� pf��iX!��=-���Ư�!B�� ��[�.?�(1���E7��#�=o�/G���a��m[� + �[���`Q���~��-H��?f�\X�E���P�Е�a$�ɿ�vh�fQ!�q�)L�a'Y�,��M>w`�-�(�5%n�H�%>0_ �)��� P��2|�4΃��b�G�]?6��x~Z��ݒu�Ȅ�*���i���FLtG,Y��#:�o� �_Q7Xm+�*ίJ�HX�d��9�Ƣ��^ )�1�!��q�1Q� ��h�GCJ��S.[�� j�7��N=Y��O:m"�����L!�0�Ⱦ��N��!��F�u#{�I�4B�M�(ӟ�ti���[��0h,1x�gR��p�JJZ���]A�~	.W�Lx�;�֒���v�JP�j�iT� `�W�\��*��d���q�L,,I-/W5@�[�'p�3<*ƻOPPH��a���,�EAZ��� X�t'��PN�28H8�aZe������u1�*�5uQė>�d��G�j����/�5!�i�pd���Z��uFdWx�.��`IS��O`�r�pL;
��'f&_V��l�N1:�tS�Q�5%�d�f�e�M��R4g�v}����Q��M�P�hW:��r:�Z���0����Ȕ/Q!<����3G@�`9�^1�XoB�2�j�qʀ�Xz2�Y�e�w�WR��e�[�lEM�/P�%v�qr���h)K���a`[��-�s�'����%��`�A��)E�K�-�����	:�~���>V�� �!�r���3m^����]'G%�d�_��0��`V������R�ח�'V��
2�4BS"\A_�[��`��p�b�9��B�YA���љu>��1+�.ZA3��54��	f�)�O ��R�L�t.7z��Q���4N�����(�Ŭ��m�Z R�5���	�ME�� $4L6�'�s ��e�K	���X_�N'��~�~J^�Q�߸J��\��oi�x �7�_X����H7m����@�1��r�X|��WU-�%�T>��.q)t���^P�J��5�B-�Q�`��X�Rh�3_���V��^\��:���61nA�AU�[e��LNV����v`j)�!H �]- :l� �H�_O}��XѳI��,]���z��X�L�U�cH�C�6�� �bA=�f�͋�d�>��H�<�* PQ5)�1K��0go�Kf��:�Qi�T��)���|@<�1��27Xm��4�h8ϴ��k���^]�-�o��.Q�h�/�BG�n↓����#�JN�����_}~�h\�)���F[ ~�N���_�G��]��&�hW_�Z~�V�������ͧV� Q,�i�x��}��!b��;�,(����yA��F]�qXW����6`��yIc`�B0��pKa	k�-C��(�\}	�&xN��b��d�A��*�?���Y� tP��7��x�q��_���r�{/NɈ�+[���雗Y�ǨQfR���bb7"^B����s�)T�UT��Z^^eR�E��_�W�2����=<%�a�P�fx{�V�o��$h�"�n&�I=�E�%x(-4N�%�a�l]�@���Z�0�L����q�KL��܉o���������<�(�XR�Z^N���Ճ��[��U`u}1&/e�x.�ӻo]`���:�X���	�Ⱥ<A�'����(��Z��cA��$1�#1���&�z=��( ����n�։Z���c��� �[zeJ�ʻK�^�-+0)��|�,��ż�cWa&Z 1�]R7�;��![��O�s�������l��� �0�����}|�w%��r���$�c�N�}x}ؗ��A�6�7���[-/u`���~d ^����ۉ�M���Y�s/��PԽe�t���E���n�]x����|���43la	(��`_��e^��5�X!���=��o��s]�~t���I<|��!�K�����~�1��_�_ w�{�������f��ڕ�� 8o�����x(j��{A`o��1�Y�N(7���+U���0@���`D���<� >%O�$ b��H�Q4.�겤�� }	bG�����8u��B� �!�P��WrO�����[+/Y����(�"p�_'��_�u{��UN/���#��&��!� Խ�Vc��-�{�n-W��	����Na���~M�V.G�,��Qў?��1���?�����(KV�i��ʼ2�i�F����f&V�Z�{�A�*��Pf�U)�82��ڕ���OWXht��')�2[�h�N�Q[� 1�)���Ů�'f�U301�|�(0ꎁ����0d*��yo-����\H�?�D'��Y �ҷU��_k͛��?������� >���1�ډ�|��뤿�����ő�p~��KN-)D��;^�zy�O&�W��������3�u	�~�����:MK]Dp�FN�!	C��R����;�*�)B����]�Y��qR�y�s��9LM���t`1��������DQUL#��O�(Ͳ-���0�ʸ��^~MX}am��";��?c�7j�)gh+�V=0K���iq�k����Ab!{�ˡ�6{�H��?t[��q��
|3���� �����,:(�x��� ��\ 8^]��?%rKS��[�%臅��ހ[�I��-s����w�^�D�S_�΢�֢PXP�G���>����V�2����)��[ 3*Z�We&K���J߀��%=���G��g��r�WTT�x��T>�Ylu��w�� ��	|O�{�_�����}E d����9~�w�'�y�PCia	�X[Eݠ���Rc`<`�X1к���ڌ����W�uc� ���1shV8%����9r���}�&='|���p\/�+���)��׀8�%!��dLĨ��-1_�����	2�U���>�t�AtVC�,��{��3���^�V<��x^�p�/�v!��`��h�y���P������u���j� )�^�1�z�_��!8��Ac�J̤"�(0���6�!.Q't�@X�< 2b�e�U�ɷxC�g��[��G%"0�Cz-8*��b���80_QnIOU����'T$�bЄk�~]�zy!�/ī�kw}` T#�齦���R�p�������X�ZV\���^��+�:�	�F��߫F}��9��`���m�a�k%�	AS�l�ҁ�T䨳���/�H��-�~yAP׋���"��R�l�G{:<��=�`�(��Z}T����gr�q���L�k!�kw�������� ��G�
h,J@Rd[�-ٻ�,1�u[=�+{���()�	�� bp0s5;U����E@}��qGU�&pR�n�ҥ���%^��l W_�7[����X��%�AѹcJ-��#�e]$//�$/@YW��K��^p	�܃�1Ő�)���-��k��L�D�o�{�H{ ��Bp�N�0bj+5UBv����Br��C��l� � p�^��]���~RQ�n ��!�_�0E�vL
:�����0���\�}��q�OBF\�M�k�����挪��v�� ]Jb�}��_5w� To.���{�g�� �D���6�t�݀�{��9� -��T'w&w�p�d�-�Q����K��P�&Y�%X)���`��[����;��9Q"�*p�&�K ��J�N�q�-�0L.����,��S붠@�S�����������b�*���b�U�*}t"%}N~�&2g?-����]/����J%SK�B�c� R2��������7J p+AG �X���I��'��yLhg�Py�@+�'�"��C�u��8{l����l饣j!��!-`'_���{bwRi��^l��h���p�~�1���.��^�t
�җ%�^����XË���zJT^�.�8��L.:��X=fZ������0p���[�)��B��4�v!�D_?�rK���-���$pqSK�t���{3f�daq�ν~U��`����UA��%i�q>�&<|L^(��$1��q���U��p��t1��V>�C�hdiG^f�L}�	!��a���^/I �5q��`�1�H��N���ZD���u~����������)�OpWA.h(���5
%} S�-�rR�Y z�jΉ+���.0��X����}*�j<����a�v1��V<��/,X���~+��h+�(�J.��
�FK��<΁|�i��pu>g���Ȯ(7�(o�}�bQ�}�N��.�Ok�+~����m�q<��+�l�Tp�����������ו�O���3�Z��PT�	lm	�]�v%_�j�!,�/v�%}��\��:�v @�OVo��)�Ph�4��XTP-�@zr�C� P�f�bh��w��d���L�/~�,\�$�nwd��Q��=�8~��)��hNx��I�U��N,]l��ux�yd"��^ I������o��9;G�	  �
ON)��"IJR�l\�<�Ti���i�.�o���8B�;���1@b@�[��:��{8�XU��drZY�RJ(~�,o���|�)]h�Q�C��7����0z�_x��']�,�uq.تB����P`� B�>I�ɟqK��=��J)���[�< D�%eTr�4�u��� �Q'������˸3�~���R����,zu�x�hT~n#����3T[1?o�-D �p����qzR�)S�I���WQzT0���﯉� ja�U1L�;mr3
�d�p���Pcb �WG�Xa�F>���ݖ�ER*�l�<0��0�@鰊��W{�6]��b9fU�~%�l��]逪�i:G�L�!&�.�����Z1T�2�|`�s������)�1��yQ-#�J�4��t��1�2>v��.Wٻ�w@?Uv[���>� CN��u⍪��j��-�;���� ߠ��_�����eI�Wɭ�vb8J��̣�- �B/5LX!����xnB��+�`3�!p�)�1����Z@��3v���C����6 �8�%KɫQ�qZr��I�!�ˍ��!��}Opn��0��(�ڈ�Y�^K�@�>
�xmq�X�; H�'5�J�=���VF(P��g�[|`$�v	-y�值ňf:J��<�IUk,�R��>b���`k�%_4��޸b� �BS�cd)QV鑅8�/��s���+�IZdz���'���c^rN[��"3#Wb���3��7G(ẵe412��>Uh�mi��z�:.Ŧ�W������.,R�st�/��	�B�}N�uB��U\����`�~>��N��$Lh�0=0��-��A^<�'�������3w^{qaʁ�#��w~���;��X�(D�P��BL8ca�&~!��u_��Ε^�BUV��i�W��담��E���G_�?��������K싦���.{�i�<�/��)��\^�8V��%U}D�[��GT� P��<�&��J%���Ģ�zo	*ZPY�A�[�:~��8;�UG�J� %�^�\1X�:�i�5�� �;����&8�I��P$l�N&3v���-�R��A���Չ�j�t���k� ������߱l��;F�m}�o�
��y�}������?���7�"�I,2�	/�u���{�n��Uk>����u�F��rC�=o!��1��� 0T_���TIgHƂ@Ar$)�g�s-3�f�S�p���#%;@0�(���Ȁ�׀�����,%(�t�ߕt�A�{����6n��[����;t����N>��!@�{�Dj���Vo�C��վ\���_:�VE(�Ҁ�G=1���H���hN��YT�!���J��>^exP��"b�Y�:Hg?��h�Հx�.O4����;��^���.OQ?����Y��v�,�V�p�pE��zF&xq��~u��a^�)���XK��Iٷ8��Q������>���:��h��9�%uL�p���d�_�w�	J ��z1�������E����h]L�|q����g�,e.Y��$���*^k���� I�"b	�_ՙ���A7R�V?�-|�o�����
��p��1Ѕr��42��0*=y�_���0���Z�
�R�u����¢� �`�~K��\�&7�0�=._V�bW�7��Ӯ��J�+�\c�S���0��v��&%;(.'P�K��%�iWT��a�,��v�
��\s�Z:�t�i����OA%3��Nv7r_`���&�U �BX�8��_�{#�}��`�2m�N��a�YA��/E��O�5�GQ��\P~�^#�<�:�X�=���,|�����Q�)`�/9��iZ����l�_�� �a]hom��l%�CR��N��k�U���?�����Qhz�`��Z|��#p�v�S������>
�g�'F��<�CdA\� ��:�	���&P @%a$�:45	eJ+�b��FK�kBW�-� �;���`�51D־�Kt<�,u�w���⪺	�1�V�a}F�1[��Q9���hIpN�V�Z��r�;WpL?�J�|�vd )��R�pK�dX@��LcsH�Q�)L��*���-��^�^��hb�tJ��¸�$S#.�TZ0��O �Y��~0h-?n:6�&{�A��/0�t���SS�[����g_�#DGx�eK���С ^ ��W�#hO{����; �A_54,� �-�d�l�� �KM_������d1�N)�����|�9�3���g~{�%h�'X�d�����u	�=>C��\��2�0�%y�&�Ȳ��Kw^�:G����9/ (�̑A=I)e�_W���؃���0��V�'��'N�+�S��[*ᛧ ��(�ʾ)�u[`�,V3F�)bh�܃'[#�X�&@�M�m�A�|�2A{s�2��LZ���A�~໓����/�l4�A]c1��._@^�*T�J�u�v <z
(WZ��./'90�޵<�Pn�^�T,�<']�s� hTuZ��=�H��X�b����J��Ě�@��2��=�'�u2��O$9ǀ M0�Yh�	��@���K��Tp�n�,���1�-#B$qU�&≙#m�˃�2�Cl�zA�Z��v��q�s��fB�Tm� �F6r�[��J;�#l9�3���e��1�?��|(��2q)�8YS��j����GZ��}���|C����^�%4G��3H�'������j�m���.ӻ	�6_�$_�%q�m	@Q��(N�/9�}��(ƕB�wZ9,��o�~�} �fudv�s�B�����x�^sJ��':x4�����%�u���SAE�,`Woń/�*�@ٸ�-�5|�DF�mJ�yK�3���mp���G�W/���Qm:��B7>�����[GHN��$�^�J�h�}�ܔ>,�MF������h?	�@��(ʀ�%Q��1;o���Lx~Y��s�D�k�+F'�����3��ϰ�h7[��������� �q�h�r91�'���	铭6�V{�5LH��y��ڊ�D+Kr���@S�t���c	�E���gG�Ԁ/Y���n��U��@.@�H��30<_Z'T:)���-�,�X�	T�̠¹��)N�A3�Az�z ,w�T�%������6���RӮډ����U#5��]���Z���[ͧ}�B%�P��Y�����׀P���:"��ۜh�_C5%��[����1+�aP6�OM�dq�%�0~,8	���J$`^L[x��YS���� �o6��YT2�4�z�4��D���U֪)[;�稽/�r��P.ͯ0%A6�'�T�%�4�l���fw1��H�,���5]_oa�� ��K�!�Ѩ�1[RE>��̀�W�`&E�˶��9j.�����QI|1ZU�4g!|R��� t
}�齾��[���(#p����Z&�O�� �)�!؛sA�
*�Q�\h2') N�#��;�[��ya��]���E��$�~�A[��b�ܸ�w-)�ф  ]�$H�Y�2�� �jgL��� ��*'�v��_:`�p0hM���&F��;�-}tl����(	F���0q�jg��=?����Ҽ ��������0���.!� �u�X�3H �5A�^�i��;�ه�!';����_�U�E��D�+�1�݀�XY{��k~����鹲��	�b,��3��Z�k� �/����O���骩���e@�[�#��1�Z�lK@�������9u|_&N��K���ɰR��=�Lijuh�\ �.F\��W�,_h�w�C����[�9��'ZX嘋�G�|^�%y�����`[C��h���X+(��t.O���K�-���C9���!�_�O��I��1��4�梷*�3A�0Z+uF$��#\S��U['WN$�Jt�w`||�	`j�8(o�'1�ܠA�h� %뒍� 1�=�f�h�3���|�`���r`^:'��A������K0������R�,�*Pyٽ�7dz/�.rA��ID5{�_9�a6?0���P�������e*W1�� �_b���� �>���fq�����A����Þ0J�{"'n�}�'x�	_[C�g�]^�Z@O���)i���BS�gd��#>/�|RE��J�U��D;�>|JJ���đZ��3\U�v��QO�4�)�,%�T�	날Ӥ�f��.A �so��Y��H��� �1�i/g�S)�Ƶ��O�?W�@B�-)H��?��2 ,�(�4e���0���p��fh�K���.}9�(��?��Tw(�°Y]�-`HH������V~鑌Zi�w� r�
z.^P�F��~��)���7W���	!��ZI�c4�����酚�� �3d��nF$?r�*`aݠOɺ3[s� p�v��)�1��i�m�c���2��'0|�%W�2��<'��~)r3��;� p;˞m�sJ����/	z�M�d�%Շ;����+� rk���f� �-qs�00��A��d�Ø�Z��a��� ~h%GF���	�)u �uV4O����5�i���	21�^ա�>��,�H[�a�Z����^�W�	�&_��9[��r�'�FʭS�XT4�(d��KD�@��-���h{��n�h������g��C[	�8�^���
W�Ҙ�V�����^����bT\Oxa���W��}o���,�]Qh�zBO?��=���a�;|�$�)�Ⱦ2�E�P�3y,8��.I��	3��`A!����:#/�o�,�h	j)�{�L�U�n�C��:ģ`��4�,�qdP�%Sw��K����v)p����I��֟�T�����x�����c(q��	Y��+��y�['���	�H|v0�% jJ5�C�	%P�8�-�����8EL��)UEuSU�b� 7�?�+	p1��y��Xӱ1;N�J1����"�8��_� S�[{z�Q;C�X�iJ�;�V,>�x������7|�Q�(;�Q	�pmf�`k�F)� D	�YS������QA� �k`�h�3�Y�k}��uiZ�q��^�Y���x����3�68D�O�.�]��bx��&5�r�.�4��`�H��	�r���Xfu:����o�3! knW��lU3�1�����A}0����·|���8;��>_렅e:Y��G|H"5pdU�sZ�S0nƚ��Ƭ���:��'����� �.�c��)����]�50sZ	⾀�� �a_-M!` ��IaI���x�[�D�+�T4j���>]Lm�qh�W�7}�QH��6�)k$\�+t�:��9	A�r)��>��;��~�9p'�cv& �\�/����E�����^��,u�Z�ş���]'1�](@%��iw�aZ���N�@P�Q�X,���	�'�,� ��	h�L 	v?@S�ˑ�g7q^�}�>ͨ�<H�j��Z6���%@g]��c���/��@��_;�P��F�N�pSh
#���&o���0�����T�Me�dB�~fvԵ��n�A6}H"�-��[(Ȥ_R0�ZXH�P�
2��؈�)�[w��o	~,��	la�@��=L���ߐF���1��h��S'�}��dAˮ(!0��!ŵY0z]�v�m���
�b�(��4����h:��������\�%u�'�����IA%�����VW
�Ű�j,�|�P�_>A. �t��H�>Kv		/�+b(��౉�)�'bF2�,S��^���N_�w�Ӌ��%�/����l$c�19�:*���rY(ަ��XV�	��?�(���<�����N
�-�b�W��u[U��!�Vw@��QLh�4���)���>���'T�#�(��.�+��䁚�k�����6�?��T���y�F�) !ڽ�C��.�p\Mp�Y��/0�l���"�Ɗ.!ͩhF%	w�1�<�$XhP�1P�2i��y �~�ϲ�{?�3�!����/�����e���P~]\��;#�% i�&W�i��Y�(��3�h�)'��_%S�l�W �sF�k��w�����,����i�A�Uqg�Qr6o�I�@���Z��g{�=NS^n	u҄X��5v�ׄ�)�XSp	zPFDpH�0�r%�H~��xM;�����KGV]CQ�ٸ��}�-0�etC�?�
��f9���iMn�O�P�l��	͖;Ӂ]� Ύ���ng/�)�ask�,� �r8�0��k��SIo@fP�(v�'%I"Pp�a��r�WT_�JN�H��VBHh�U���|���X�*�,�5A")+�ne�������r<$�h0��������:�Y��,�i�4���c2#mNAk�hJ��b�� ����x�L��"��	�G���6TA-��^V��v��Wq�=8���#���Q�x0�Y{��_���h�!�mX������Z��d�R	����H��	�7��.��"K�]f ��J�z)%-l�Zv� ��i:
z|H���o��;��ǃ�< �[��W0r����fQ�*N��]�����(��vû������h������	~jP]q?�o��-@��
:vg�~�!�h&�F˷���-Sd�N�	@1�nU\j���^	�Ta5�6�$�K��F=.^�Ut�O���I����`F<#} ӻ
C���� ���q)��'�Ҁ~�=c�����QA	���:���h\2�%O��Z�VdzT�B>qB�T��,�
1#��t(��
�f��� ���V0`S(�*'_wPGhX�yˇ\��@�i郼����%.
��|�^�!�Y�}\�'�705��O�
�ˬs�[�`��3@<����������r$#��hW2gҬ����uV���I�u�J�Wi�@0��9�%�%޲�_�Zf0��9]y�Bh4��RL�h6�A+�X]�MbC@o���r�c��*��O�,�+��.BEK�� �TK��qx�R��,ϯ����=Y�;b���47�w�f�	(X�Cʉ1�h�8�ld)a�lO-{��E��AK���f	{�$�J��?0W<�f[G� I�&�j;-���h���2]y4�#Bu�mIQ�b�%l_��\�W�_G���$O��+2�(>�	��˛�������'�B��Ϩo��ԛ��i�)o����V" �~aZ�A�q��T�h/�o�ڽ�D�fM�;�Fw��t'x� ��i���e �_5�a� �-���N髞�咎}��-�����l^��hb5�G�� -�fU�P���(���zU�,i~��^���� ��K�d��	�r3d���@I��(��jhI~Tb�Bb����*zZJ^��@z9�K��!h!��%�9�AB	rUQ�k��L 1Z���n�X�s,#E�͝G�A��:(�J��_Uq��\ Q�D>w3�P1��#jpŚ� ^�OwU%W�=+v ��_�;"/?^a6�����	�jYR�$��!��zg���	�h�U`��=3}��1;Z�g�-����I�@��>� M��f�_�%��(�i(�Q���D����6}>��xy��4 t7I0�`�����[1�J@!�G�1�U�je���49��x�:1� �U��\�F%�=��Y�-xu3!�Œ�B�w1��,�`��nTD	I/�PU!6 �(ڊ8MϘL�}'�@���י��Er����������yvf�V�`�fhH�$�� ������|�o}����[b�@���Ruo�������P2����d�av|�trLH��!�Q+���� �<��eE�eoHqGX�@%�2a(-R�`�ߜ��@�H����ptqN]��} ��2��x��A����oae �`�����Fy�� �DHT߃%�T:�~�m^*�|��(���^^���8��E�2�@c�_�xYL2�Nd{�!	hFV�
�����Q@wB��'��ݠ`5~8:E=�/sv�B�a_r��-G|9�zj���J�~B��P�f[�"ۥ�� �Pe՛ݫ�E	�|Bd�'��Č��c�&��n��)���$`@!�h#^%~���%*�/@1��uP��9��������
��XZ��>82�6 W�y)�1�-	D�/��XI��~��zhH��{�@������Kf�1�O�rkǨ0�W��L��{�U��-�w����/^`, �-PU�yHJtw�{HK����C��tJ�*أ��Y~D���G8-Uo}����Q}B��`}(�Z�ܫ�z�������(�0���	.�/υN�z�^�T���dB�s	W�{�>��2@bw�o�*�l��p��-dc���O;�*�Lյ�}L��w5��of��`������O�qc:���TL>��`"`�H�� �W�|9{q�*�ݰQ�p=�7�WAL(1Ƚ�:��4���lQ ��9j��:�
Hs��a��@ѿ�?�M�J��6�x�D�����TB�u!u�6S����	id_���$�b��+���o[����0�*�l4���c
�R��%�-�'�x����e}c��O�xWj%	�(��,O"���{�VVhU)4����3!#Z^;YE8�~�t�#��KY�u�P �!��a������_�x�%?�Uđ4ٛf���F���9���;Q���P$3Xh�X;�ĸfJP��b�UPM�1jƤ�\��?������x�	�0��C�Z�h�==�n�5D؝� �&��?NJd���)χ�_^���u������6r�_��o���V/P���gO���2�����#����N����,,} t�����gM0�d3���^�@������0 ��6QP����H��@e�M�'q�b3u����Ld9��sn`Q�ŸHf��w�R���+�lH4I��A�lXD�5��&��}�+~��ܘ � 5�Љw^XS�(:u)W|p�HA0�ĭ���.�����W{.����,#�Ց������@D�>,r]h���_a�5��̀������ *0�Y�V�^�����e�Y[������!'�\7%T�zWh�R�f�T	\����� **2d/��.֠�5�90��Q-j��i ��H�X�Z��
O�`1���Y��N�Ă��@E���y�Z�2���ey�	�1d��9>\m#��������Y�P][¶���f1�'�(O@�8����4����|�X/�����Is�[�	K�*'3EZQh�fY��P��$���|CX�1�wa7`��_!��{�B�[��V��ߕk{�iW0�c'a(��e�}K:�).9�tzJCͺ%��!�k���<�$��= ���Z�,S�`����5�4��65���r=�1�X$�PƱ� �ͷ3��`�����]N��|)̀�!�Xheb#�ى�Ud!E��	Fx�h=�Z�r��%��#�v�O��\��6,L�UP��
I��2�2^-��F-{���Y��E�U��IK�NN�)�~���0���(�Q�A�����K��;�A�jA�Aҁ�g_�m������A�)�8�O3dݔ�
�0>��n;�Ak�\���y����5U����K�g�!g[ϐ�B�f:�����5���d�D!�`����t���xa����.�c��O3�F��� �˰�,��\��N�| ��61.�q��@�(�Z�Vi9[���V�ϣ���[\��;���)�!/���|���oX���Y h,H�S]�՘�-g���E\�`��40�Rd|J��w$d\0V��(1���#�W�󀬚F�;��[S[���>)@�U0k��-���R�P���x�5��A�V�U|�����FfZ*(_����A7@��5��t�v��X�T���\���as=(�	�F�6��}��4�Ֆ��=DvN6���]�yx�	�銠��Gh	��hiW�qKV��3X @{Z�*����	+��YYZڟ���џ�h�ps�:���b[L�����Qr�� (W hRw�M���H5�^SP�� FV/�N�'�d��MX��/3p� ��-)?��n��z�	$�P �|rD]���<�@��+H�[uj�c��k������j�\h1P���P��̭5��ҀAT)��ݎ:��Cs�A��݉��S�n��`t����*� q_�wO�� �Z!gH��	Sa�3B<W_�����<�H���X@BʻQ%M��LP6��ԯ,۳|/ז��n��H��V��]pz_]��h�I
��P^spY�׋��������}.�����	H��U�t�@��=�3��9�'����K�������-N;�� ����%}eM�� ������n���0�Z�fY~&%�>����(�P��g�蠽�hZ����y����X0s�SNEK*�����(֞�^X �Wh��z5�� -}�����~�"���5�`PɤN_�������a�X��F�;�i�2؋��-�R�	�HZf�C�I����3\ �0��8L7-��{����UU_"�F����G��	�Ӂ[�O��a�.�w��ktT�X�l�%Z-��?0�o��F�����J��0�%��U�����5j�k��F�ɶ��C��s�Zv� ��J��	e�qY�R)�W�> �th�JI���'|�D^�x�%)�in�8|O��9�6E?�%���^��M,�P�/�0.��P�-�1�`�(ky)�[�(]m�<���DV^H��&%�e�a�O�\*� ,	���]�M�������6���h0$3��>����!։o�����1�p�SW�k �5Oz�4U��+�A�K�a������)Oă�� �
9T����+T3�1�ꑳ ���]h���'hF~{~�X��ŉۭq�,�n�Rd2o8��p�]�O�n���r���@u;�K�e-�g���Pa@Wm�R�v�uJ =��w�1t�`�Tjfo@�&�Wq�^�{��=�d��f_^��?�E�� �Yo�f�\�(�D�����4�s�	�A��.�^�����4V `#��t��>R�	�.���]�O;�7�q1pn�P@"�Xl�U+�!VfV{��|�ׇ.�� �w�!���K� ���k6F��X:!d� �R�z~���7}ch���ʋ��U��j�wJB,	g�mt���6�h8 	1�����F&�*���Ϳ�[������o�&����I����o�뷾P"@�#�P%	�Z����J,�&���2���9+�&[+�����ahHE8�D���b��4�[f�<�A�z��Sh� �{p~��/�붱[��>�%��-N�@�V��s0����d,�L<�^����e��HXK��됵hD��q0P��0R�zQ�SѧZ}V�����i�H<�^�PD.���u p�B���LL�N�'&?\�pZ�:Txo�� �����p�m��uLi��m ��W@�T t�viS%	�E�shO5�'~��/X Jj��g>!��T��u����36�e�Q|�����Ǩ��=V����_�n����#E2���n����.1¿����&?ιi��߉���e�#PG߽hVm1�擯h��.r<�Ï1ع�yGA�(U��b���TS�Ռ�nDY����S�="�~ÀO��?�o�Q�2����x���������L>>�1W\)�c��_;�@��������X����]�&Q�B?Lb"h(_T����������N�������)
;�:}"/a��g��T]�'�\��B ��&�K�����XI7/v��!�p�d{x$]1�=bh0�x,�N���m��<?�I���J�������I��l����ocF��J�>Vp�AaD;�w��>��*�e����.�	rAn���f���Ì����4�u�^������nFa�uo?B�_HZ���D
�	:�d���r�=�ˬ�	���Y�A	�\��xL	�K�u���1*�6s/�FR��~E�!���K,X=�kN]/�_�.`6[�(��ɱ/�P�
>������_Κ7ҕ�,�h8lJ�-�:�xT1�[/���XlKW�"/�wz�Q�r�F(kT�k(ե�VAbZ��]秄�= ÷,k�(�-���_��������=�Ä<"��s�[6�~���!,�<[7�s-	�4�tI��n���4��i��P{�m�h~�FjI*v)U����]��	Şat�/�_���K�jT6�i��%1w��bN�t��*��l9hJ��c��[��5�ua��yHx���l�~������P��0=&�y����X]-^dL=V��n�f�v���HS�RGI�f5b� HDT3�@�)�H�L�?ƀ�^-�g���G\n�Q1�W�a�;�C�P�/���!�ZW������?&�=�Z��׶���h����c�������أw;E��h���j˔X5�h�h��#s ��E�K'u�糞į9�2���$���hg|��?l�0�p��AE;�e4 a��;�4N��Z�72 z�Y�&����Z����O�0[Fj�4P�����,}a�z�w^z=���ͫ�X�����S�oh�����J6��	P���,U$� 2�35HWK���t��D����)��xI�eJ*J/+݆����O�����G94����ǋ4�� �"=e��)��oN �a���]�QDrR�(_������hz��.��N�j!�@�����Q�[0UY�w�"��6������� ��1�!�h-0�ȗ�sh/��*�hp�-�2~��/�r0�������]�AE����S0A"����i�[�P�0	/��s��:�l�� ��,NCH���43�(	�vV>-}2��
���(`%TX��>���;a���}a [ �F�p(�Y	��|�l�1�.�3��C\鮺��U�?:��Ў�	J��7[*����&��a�9kAܩZI,�v�W���[M#��3���%p�PVhEg�*0ڑ�;���hV;8�������u��`G 1�R��N1�+�a+)*ʿ�V@���>����(��S��y	����-2�Q���{b������D-_�����d�90:$��
��Q�����rX[J!�q*�|��!6F�t"�/U�V�-N�I�(�?��_�c-*�[�A�%z�X+�.�%_�ae� $W�8N\F�����Եh>����f��9���ʟ�ЍQW�T��[h�$o�OȴMZ!�rN?�3�UPkuE)�A�wp�'��wP��3�2]���N�=��g(�����(�X<�ʃ�H��b� ��Y@o%1��v�N�k�.�lg�%uh��½�S�j*�f��/H4R�� �0�Gx7.LZ�@	J��`�]|$�zl;�ۏ�y_fS[c��d�.�Wc<��Q��iDK}��O,��N8�Y~8/�aG�%�	'@o~	�_�:h|g��D@�%A?�^�*�x��kJ����wa	�$A���:�ʉtIDQL�O82Y_�I�p�`���z|2X�D'�g��*��� !�N ��yI�r���1ys ")ciC�N`^�&��:��`����ڹ 7:h��z%�,H�S:k��֖ 0�fY�_�c���ݶ5/N��xXi�J�8��!��g�ϐ�8�\�f���)���c2�&[n��0~@iņH�_L��[�vP}6k� �2�H���M�@{s#��-�
*� C�͌�ܿ	�`}�=�5%) �u7���I��q�J-=�h��$�A�N��X� E"�IV���'���&-��l�vd��ȶII��L�t~sw}ׄ�� ۓ^�[?T9�BM❉ �5�X�%�[1�� ��Ks,�����������(_+�lL>�UA�� ��3�j�)�^�����!��u�5��Y+\�P�	O}R;�A�`��YP��=��q1�X@��S�d0�o�1�4"s	�[o�=�yB�$^��D,$��D���Z��}sB�*q!��n��N����5X-=؞��)?�x��$`�O�A?�?����D<-5�a�@޲M��).��	*
�jJ�$�j����[�$��]�" ��]��[����B�d-� �� �m,`݉�`����]�A}X��;���R0h$,�f�~�@��jRZ-�)�DP��]��9��z%Z�?ay��/-�y�Lx UXh�i��~��"B�^�T��+�b,�D�(�Z��z�� �/h�N7�A�U���&���� �a��;>0��(�(���R0��yK�M�$ �l >�$K�����/���	�^����E��i���	��\ �q�����#)�l�JXu� GN�QhOS'35X�w+�2�,%�j��/N�'IY��C��`1��s\�,(��h�9�K]��	U����RF�"�ڮ���p7�;�	Zh0?�J�ۼ�շ(��E@��nK���X*�����N��Q�9��:�;���(g��*��<@�@����	�i�_S��]�R�8�J��%�T��M����2��f&6����7�(X��[�Il"�� |�(�fQ����_��P�>zZz��PA�H�-Eh�a�b@�3w��l�U��<�)�:�܄��.P�{z[�x1�!ȿ,&iq��筙ϊ���S�Z�-�'@P�W��Wt<:���F�]�P�5$��> 7�ޓ���f�̤����_�� �c%%����g�v��	��x&�2 h�|e[��i��hS�|ZR�,o=�X)�-6~�-0�3�^<r_s6�>r;B-E�Rq(�L(&�i	�HX*� ۹^�)�:�r�\����Z��B#�-�} ���gW�L~��X\���ʂ���T���R�p��p�yc`���u�$����˾���l��|I/X�4��`�$j�8��|L���Lp_��S5��E�Q�gs^�@�~o%E/�B�ԱeP�U1�>�-��}��)h�pC�~l��&�
/��e����BZ
��|򵢷ة��{���L����5� �s�!:��rw��t4B�Q9��)��y�e��h�D"1�+�+?6���}��T�:P<h�Q +�=Gk�^�w�N5��a�"+�p���	9)�(���Sn^��<��n�V�J hn-&�����8zh)�yۭI�Jdɳn ڃ�>������ ѽ�e��?d�ʅ�B�hRq�W�� ��5k�I�\օ��O��Pݍ�?lSy�����Ƈ�_���PRh	J%����� �:����)o��9N[�WZ����a����Y��(�����'j� �n���(�������	�W-/Ww�;��I���KCX\1X/lx�$tԽ S�h�	%���I�]0�}&�mW�8J�}/o!9TR8����)����x�{��!
��2vS�|�a
wX5P]S��фػN9�{YF%�����#�hA1���1�u/�,�2��;w@-�@��O4�
�&u�����B{Ah)���؁^�Nd�z�0݋��>I��uX��x��\u���g:r���fh���nN)��>�]�=(~�<�Z��=%)w�{ �V�1�En2XP��l/����z��x,tp�	�7pU n H�J�&\�5�d��� |"�5F�Hn
�� �;�1g�q���!w��h�]�1X��(�#��ճ���L��s�3� ���0쳅 ����Q�c��P����p��0�pY�e�%�E�v�w��*��� [Jt`���n��'�0ˇ.�B���Ö�_`���9B_�6��<wA{Y 7�
�&�8�LOO/��*�g�i $���%)�ٞ�R��6� ���Z��SLL��\���}��W>�]2]]N�鞝עc^�C�v1�ZǴ%G��39�`��h�+�1o/�A�Q�چ����m40����7�5��;"ܘO���C~H�s+C4#��Y�@ع��O^ �{r��<]�ϵ���gn`Zk@��R���/�U9Se��pY���S�AG�o��Ub��!xqK?���	�}�ɦ=+�	���>��T��,@_/�źЕF{?P�A.����z�\�	��[��(��S�DŬ�d��k��<\n�4p�u�/�v�+�%Dh�R�(x ��vY���v�f;9�N�'h���ȓ�N���]D���iU���5�໨v���^�� �#��~�0JB���|�_y� �w%�Tn��B�&)L��Y/8�},c�|�4�Ɏ��d�9�L܀�h_�^p�O�gq���{rH�H�&�A��j�$����ӰH�u>���}\H����h�bL�P��fr��-����N�Y?�$���� 3E��p��ҿ�ͥ 3�ŀ�s�8��s��� �/�\N[�VhW�`�E}#�j��l�4����R�/�e"��է�Sy��T����$R�(E��(E����|�G"E��7����!Kٽ����h�m-���H�fHS���*�!���_��dM 1����G%�e���C�.�S�8fzS� *=zR�?��-�X]�$��/�R;Sg[��6�wK�1�b��#(�%)鉊�E�m�P �w����ʄ1v�8O���JZ��R83PF�|X������HF�<��N���~NaqXF����"p��Rh�l�YZ,1ӡ�E`�R���n"���f�!��Y�}(	8�[R	��H��G��^.*3I�/Kˎ�Nj�B��,���)�S"'�@���rw�	�oWz��������$��WEH�x_�}��͈�� �PRXZ�\`�����a�CS�a,{���MR2�Y�6 W��Bs}��|0�q1�%�o^�#h��k��$�07�����P����_���	h�FX����[��>'��yE��r��ԡ��Z[h�zt�i�SQ��/��{_?��8a�0�ɨ�a���^��2.���n���1
�0���>��݃�E�&����{}� x0'�AQ������@ʀs�")�1�%�a� ~@-yZUv�R����p�蝭(�K��3
�u��	�^(r�H]�f��k�L��W����L�28Y
_U�4�L����=~/�Y/u4/�1^R�����f��dtyd>1\HnQ��@�yĢ�N4F��x�5�t�-�h	W�-���-���ej&�ū�	�sÜ��ܺ -�*&L1|�(�� �C�%�zL�`�6�f�+K$!�����~�5e� U�x��c��C'�<�k:��f�_w-a[L"W���l_Ƽ/��^x�9�:�WU)��7PeW�sP�BG���1Q�W�j�z}3s�7�$�>�{��q���D�	'1���U�2�iB��`S��sS�� �"�s�r(�9�I�x,� �h���t4y57'c�� �YJF��:0 ���[�0�p滴].eq�?�9g�`
ihC�0o�&P��7;lY�$Q��2�����0^�����z�.͔� ���C�j�B�^8=�� ��!��Gq��s3LY�7}���zz�F�20���g(')�4�9h<r
z�%L5~ga�����A(�8|0i�$WXB�q)	X-�P�a��j���<�ɿ�y�F��QKS�k��v��}���ƳL|�1��iS������uhurn?W1����Ů��H@�^�2R�݊A�:�/�`/_X��`Z�q�2�Ka2hD'���1��)k���~r~{��j���(v� ��*2�~��A��>������z����/�ġ1�4��X���������iV_�^�h&}�Q)hrA/��=���4��V��7��2y[>�W\��:O
�4 #�S��]-�xv_Ew�\�c["%p���υ/̎�ǀR���%�Z���2Zx�;��
��?K��~�!��i�G��k8�,�|w"�|}���(!>���'�>��a/@��=l��ݻ��A�����#��@��v�8�n!�qW�*v	x�MQ:��!L�V�>�8����k}��Z E0i3��>-V�	����nA�?�t���9�1��� ��t)O��N� �;~*l�L��4}Mxŉ��~��x"���B�/��/����Ƥ��FBJ$�'t�,W��IKk@��\�J> 1[��g���j�
!�]��_ �!ջ�wi`xZ#�K���vb����lw �1��h_:�3IX��6B�����5g0E;�q �!��*_<�* �'�:)��(z�-�s��RB�;^H��n'f�i�?D�g-��*���a�S��5�`��,;��ut��Lü��X]�%�	� 1.�h���9X6�^�;�2�w,�U��`%lu�%4	��E�Ph��N�\$���A�꣞�a�"��yNH(�J��r	����h7s+��-�v�n��t��YfZ�Ԁ�!��xZ]S��2<�H��^��nk0��f�7��u�"g
h�|MDWC�q./^V�ߩ��@ s�[F��B�g��;�R��$ �pv�;����$��� �mnNː#��@�OLX\^Q-Pzw���!��?U	�x��V%�B�3��Z�m*Q4T��'�v`]�Pk�ѻŉ�p\�i� �1��,5#��N��L����G%؟v�UK����a[:�=\*څMwsW%�ބ���(����*�h��`��y(�f<����ΐ.NZ�x��[(�:��z/��������`8IF�lH�,�0Yu U�c
%�j�I�S-z/	�T����]���4��b�P^b[v�[��A�eJ����W9�M�tL�� R��lm� d��(��d�X��Lj��N�p��;J�4��/���8Y��ٯZ� Z��W��w/�r\t�����辢/�5�ӌ'W�n�C�N�U���Dk�Q�=<@�{��� 
��'�Mɀ0��ߚ�W�O��gd�X��-c��H���dF(wn�Z@��'V��	y�	�=������.�����z�3�c�H?��{w8����uh��z��j��Hy�<B�晅�[™S��KX�<���[6I`��h�� �uy���NN�L����.YPX0�g��q3@Y�T>}��h�x����;�R+���Mԝ1��ab:�o:���%t��,Ю�UJM!��)�v��| Z^�N%L�x�,P�o�j���ZO�eP�����p#cX�%�Z- ;�g�׌�}Z�қ��JΠW/����TZ��1~��i�C��W����V� n��+4 Q��)�8'�e}%-��k���I�#~�,[�*��t�����2j.J|�e�!�wS�@U����u	|���[��	�S^f��#J͢n��RN�bY��gMQw�MB!�uey�ۦ(S��7��] $bMx8-�t+����_}�}!�14���pS���ht_���1%y�@��'�XI�7dg	�?a:����	T������!�1Kʨϲ -�lF�\� *Q��Jf�P�wd|h>m%�G�I_D�0eMrsw_�8{Zͬ�V<�`	�����H�;.��4��AI�!�]+tw��3�h�	�!��e	��Dw|� �O­�t�Q� bڳ�ϸ<Z�|�(-��5�/B[V! �C�)@IO�ip[_:SWh�7��%P՗s��>u;I)�h��EZH����i�;�)$�f����/F*�h�'c[��ek��^%�I}��wV�O��� r/%�3AO@������ ߶�ze�a�	���ᡜ�x� ��j<J�՝@��s�S?飯�(,Ph�l�N:��Z�O����(�}D�[��9h�S�鹄�����b�V��˪��J��[�����g�`���v�$�mc>�\�qR ~��h�T��_ٮge��{_�4	�
_'q�W?C��vQ�B��ꙛ��+ᴥ��P��������/QK���Wtd�ˋ�k�~!�b�/����R���惷Vݭ��	2
Uf��k��@�����D_�C��ZY�y����:C\^�|ZJ�� ��Z�x)r� ɸ�{�Ikn�H�~��P?����h�}�9!.�\���V> ������$"r�(Z;f<�7�(���Go�>�v^�O���� 5�N�I-7e"K�f���͈/Hdx��ok
���Š�Yw���2c=���Vv�<jO��Au,N&��	c"���>���+nS_p%�(�<�J�-lYRhpB^)}	ތ��@�K�`�%i�c��n�"������h���oq���l���8�Q��@_���r�e��"@�X+�e!#,�ۺ	qG1� �ɕ���:�{��c?���������yvH�U�&���R��uן^mA�����	FDy0 3�nN`�%�AJX.�m�t��Z�y�^�5J73釚t��i���O�(�BY��	;3�Mܧ
�)��h���Z7!Я�<dN��J�Ը���ӭa���4w�2���\�;$�K ���rK22U��Ƃ�
� ]���,�����PQ�8/OA|)@�7�u�_'�?o&��� �łN$�Z%X+x�	3S��_���-��tY��l�E�Ya�kG�����.�����f@��� 9sO/šazK�OB�'� �!�Yg�q=��E	�5H�@��wC��d��*)��%V<]��L*�͟�S>��b��Q-{'HFu�U���k�L�K�1!��~@Ҹ(�Q��͏��S��6R�UI0�Y�'����V��g���)J�!,�	�sD" �^
2_ ��3���辢���{��3� \B!M-p,v+�A���,�>�?��3eh
u\]���-��k`��Kc����aw1����$���(-"9t��MG.&5�.^Y!��t�u*�� �#	X�oI��+[���[�&�E���D���*���,VAd�>�;%��uR� ��-�"/f��Q��:��
Z9�骮������BG��(�Y��a�U+�p��Q��b�*�1�C`�����B�wZ��,X���'na���;0�ӽWN>�D��H(�Z3��)�qp�x˄ ��������@�X�F�$�o2A�^�����h/UFz,��9:�){W���߬���_�����-�!����nW��ELA�_���=�t�=��n'\�Ө�}��Z[@PhLr�L|���JFL��w��(u�=��=r-rv��R����>]W���cO�ʕK��l����S��懣��d�,F)/����z��b�P��Dql�,6�@�[M�����ϰ�~��K��J�����r�}������RW7�N F#�,�ם�kX5|8�x��M�LTn[~�D�p�����X�	0_���h(LF~�B[��R%#!%���5�ӂ1������e����0:�����y%�o`�4�"Zu�\� 1�vJ���t�*�� �_�-\aIz��C��E��_D?X�'l1�@��[�4�\d���}��.?�5Khi�1k*�z�7aQ�~�ղGW����'�u ��2qB
	�)�������λ�췡+�{�'��� � f6E�c��T	�^��0�K]��3�}TX���Qv�е��%�O?�� |^�џ�D��@^�d��n�x�&4i�L�%T��;-j&R�BG 1߰�	�}�'�Pg�]8��7u�H�9/��U���@���&	�>�� #�Nz�gg]�
:O���?j�3�5���/;�
�����;��Rj7T�6�J:�^ (�u_�{e6���H L�h%qD�'dw$�U�L��!1���`p�8.�,P�2�Cʓw��n���%����@\5K�Ďl%ր���i��<Z��W�m370���>J����[\a.w�G�ʪyI+�Ee��ynn�VZ!l��`9���wE�h920����D��'�#��鞠�CXh��]!�ܫRt�	u� .��tÒ!�
�j�y�`.	��ܿ%�g���_�p���q'[	]�I~_�x36�X�@)��4�$��nf�vSPh,���_�RKȇ�<��W�(����b0{=�+�Ո���i�^-�}�eE�S���]C�� B�[�r���9�D��*�p1��S�J\�q���@W�
%X�ר��#�������'��(�`_�ViJrv]QW��Y@)S���>�/��|��8ej�Z�  [�~b�U��+�X�k�K$�2��fh���:4������V�Y�S�;`]AV`��N� Zw��v�8�_T	��x�U����YWL���HH�O���
Dv%X� ���	��7If��p| ;�N�/V�$���9Ѹ@�H5�"�~�-<��')J���Q;3F@>O#+cH��*2twz���;�{�^�����P���\+��^��V�w�L�O|K� Il��JU��d-=������;��;���T�dL����@8-�5(]{ⴈ�����{h1^2,Z��~f����K�����6,$�{_�@B�!�@f�%1����0֛"�������Z!��0���P=��y>�(L�u��P�Ŝ��QI����1�݇�����iAO�P��+�-Q��w�e�O�J�]-&�vd���,JQ��bM�0�@J�f�b�&k��_~�=g��@��O�\��8��%�p�0H=L���]1->����5~�YJ�N��rz�Ǡpx�>I�9Ze���GRJ���F��:�P�:���@��m�J1�	�RF ��^h�T[�'�/�K�^��uL��/O)|��2�)�kwu�]+����@l�o�21X�RT1����ȫF����f%��aZ��+�Y�\�0빡>�G�Wh&	5+6_��)�U��|��V	���sȭ-J�r�/�_�Z� (�_�m�|&�����鿮�YF
EK��pKв$�W	,w�x�iPng%X�tX9�-K�������G
I����L����Y(�@o �eL�S%]fn ��%�gH�}1��ڈ,��[�Ú�X�N����%�Ȱr�����y�c؊>_T���_��"ҹ�->�OW �9D����⟎2�#.	��sԤmO�����0!؞�����vX��S��K��tXh�<���k)W���I���&�*��Zlo���M1Z��:������H0˕����������_X�A\�4x"+Y&QN�6���5.D��_�"��Ugؒ���S���ݴ6�(�Q.�kJ��W|D����Y���M�j���KE`^
��.a�=,l7��5�,�����x�Yh�n�I�5g"(��چ��v_�_���r_��w���%��-�� �}�Ղ����W�1gsE���=����0H"�&JE ���S6!:��^����I��T�'l1D1R �oN-4�w�����y�&��G�\�������7\�O����r��|�/OP�q)Sd��A���!q�ajj����P�Jb��s-N�]L�h_>	��<����G���*���[�5'�%��|�M	w� ꒅ>ꪅ�1��h����U;��-L_��*C�:@�O�81�@��(
)�Y�U��`nc_��������Y�f�J�$��z�$Hn.,�Ah�dk�yJ�O�20;1�����{�d��STC%��d�	E��d���0�1&��8�O�;*J��r �QU��h�JE��ٗ5@R��^K�����B�!$�[?8�dk=v���8�
z�����{������v��� ��VKJ�X��MWD	��w�{x�O`هO�;U�P³!��c~�cp�t 1���f�g�Z���aB��� �_�������^�k�E1>�Ӓ���&�L���6a�P*�S��Kv-?�T�xkW`f-��pY	9{�t���(\K?1����kQBb�[���,;�A��r4lH�<w:G`٠;�y鉌�$e�(z��q2��e	���!
d����5��2�7�(�нS��75�_�?�r�bd!|[��n���>��P��s �ധ��^��m׾�����Z��3�ؐ�E�F�x�A~�#����A hM;dL]�fK�@ARb�H[�c9�s-�2���=�ߝD?E.�Rg3�2�:�6�d�y�n��U�P�h1����U��'Ъ-�PY���jh�|���zVl	�-�@���O����-b�tx^�:,��so��#'����OX��
R��EzKy���60���u�A�`�bSEP�]EH�q6b0�@��	w�=iXl�[hD�U��('J�e�k�Z��t-Yl�7Mv0�7��q���·�-�6�f���^�~3���9�퀷-
�8�Y�/zn \�\]�{-&8˶@�Wk��#%�u�M��/�R�����QBU��Iݞ�'����-�@�^�r)����jL}��H|����_q�?��%���*o,���	3#���7�u�%�MB��;�AI��u�׉uXB�/-�Н���n�5�`�(�b!X��&�0&�	9���Vs)�1�:!�%� ��a�x�}̷�/H%Մ�,F�7t�ۍ��(� H�<O���O����A@�4rfs!�ӥS^��%ې%N�ߠ�(J�����޻�Q�MF3�v����Y��}e�i��BtX0 N���\�-EO<�TЭޏ[g��$�	�e� N���Z������}rc;Ijڳ��.��f"7�O��I�K��i��̼v��o��	?vu ��B1A��H��b�noU�4[��	�h�6u��94�F���P]7 ����K� �%n�5�&!s��^Ft-�a�cD�S0t�%���g�YiRW���]t�����OT�6U|�X�3L��-%� r�Q��P+�'A�1�|?���H~� �w�%�ȝ}��b)RF�d6kc����Չ�~�X���K�vUy9��3 f �@}__I�Ma
:�G�Д���W/Z_�>�c��R��%Ei  �n�a�2�f/q��>H�o��	|5Ci?�^���h��_ڒ�x�zt�/�9ߞd%Խ�Ć/�);��؉ø��p���csu� 	J=S3��� YX�4=�%ܬ�.���ux\���-I:�UP�1��ɿ�	�q̖�]Z���V����k�
������?�7��1�+?�/W�`rk	�K�'Ŭ�յ� ���@h��_� -{Z	��R�t�X:|B��.o�C�G+��HW����	JG⦧�U���I^1��[����=�e�^�㟂��אh�?9$y�6��kNu�J1�ͺ	$ �g.(ćWH��)�@���(�Vx�	�f�%�_�k��(h�'@�c#0R�zK ���q�rQ4�w+7���E����՘�b��{t��7�O�@�^6NF�`-|�B��~aI����k�j*�����Ș�n-�2���`�"�������>ފ�)y�}�H�T�4���y��@�� V���!0�4RǠ��.t>#͉)��K��H�WkGqXN�щ�:�P��{t�1Y��wvJ� =h]��)NX��~�-`��* �}��nke -�~%��o6�"� ��ĥv0x�'�جHY�	H5� Z�!��8(\p�vz�s-���^K�vBg�
�{�6�0 R��T��>[���|��F�*��� ��_�jf�[�B|Se_U��ƣ��hr>�|��q��^�ɃٻW�h��{W`�鏚��`��(;�)��V��f&�3s._1`�����R��@	�z O_�K�@��#�}1�-h�~m�P	8!�n���lyx�^%�W��}g�*U����A�2! �_�h�[rȁ� �&����'�4|�x���;'�=^�&�1�I�}��V�P���P�Z�\F&�T*K���A�W���viyON��pU�fJ �����X��K�r ��-�&� �5�mKOD�6P�s+WjnZ�g?`X�]�'��7��`����(��3u$*��:3dL��i��֔���f@��Ag�JT/�%�;CκrjK����ߋ[�O~��	Fx�_����U��c�N��x�:�0
X��\���d`��tCq�h�V��\��Y�� ���(r�'g ��Q���-�)Z	���i�j'~P!��?JC�`���9�,= 	4fu��W	��`��.�yI�'\���E5��� QS4L?���ܕ�P�!����Ď�w�vhK0V�dR�8aF�~�.�@�/Y�V�n�XӺ���Q����7x'	�<�ud�_)�� w0���=���#d�dJ� �^-8�WB&5"��նz��͹��z_XY �Scr�����)� W��Z��`1�-�+^&�l�*� '��U��vi�f{�����`<�����r�,��0��^4q�I��2Bp�c�`��V�,�~=��4�6Rb�V�R�m��4 :|-�r�)% �Z5�ORf�Ee�񶥐Y�Wً���iD�	!��/�[Y:��Xx^ ��mYHo'X�cp�Ѹ�)�|i�dDW�%n�09�Y��k�������8T��.��M�'}E^U��[�r�zDa�N�6}g�d��)]�������/��vV-�hW�]���k6�^n�!�U|:p��e�X��� \�c��k-x]��h2ql:E�!�Vp�# �5V��D�@.G�@{�\Z1�)�%�q%T@��o���Ygq\j��鵀il�?d��?0��x�iG|!�_ka�FP;��'���J��K&	�E�BF#�O�gL��p�}=[-�U�<����&`rD1�5� ��!�ja�~���1��LD�#>�C�| e+L@�Sd&��+�k��
>�[�0˙����@h=7(R_��s�T�&�;��j��~H�V�W��[�&�!�����b�+��`f����<���Ё�;�_��T	hO�4��QC�An+Ä��62"�^��_�]0��N��Ab+4�Y�>�d���y^j��C�� #�t�]^E�lGh�ǚ}j�̒�m�7�H��9�U�
�	��$*�$(��} t�}'�՘��;/t�i�W�^P�S��,�Z�R����>�����߀�h
��[(�@�v�1�Q�(W nL��u���ZH��J���-{�I!1X��!�����1���ߴ�����u��>_ �x��6�]�VP6L�	)�Yj�I�s�n�%���W�mJ)��h��d����؇�XU񬰂��SV�p�('\�-��� �������>1�|!�/I��V�����������nP��^h��U�v�j& ;GXC��.)�X	Ƽ�T�; @��E����ɲY1�R�r5�g�Г�JH�A�͡|x�.R? �	*�f0�b&����z��G�R\%hp\E�v�v���6	SK��L�2(Xw�+_v,��K%}�	�������f�O;h�Bw~'�]U�:��R�Z3�����/���Ǳ��0a�:�����̷��j(g�
���>��S�8޺�pn T� �&�� �r��)П\���^f���$���ހƽ�c$�D�ł���	��UqYE	��P��;�(�@�4��z��S-,�ac�a[T��X�ó�[ĤֺOS(U��J,Qv�	䝟L&'{qy-������C1�)������%���,!og ϐ�ob�nIL�*yD���6WR
| �h)�7��x�n0*���F�Xk�t�`V��0�	X �fW��#���H������KU`�Aӽ��'N�[P���0T���ٟ���Ȩ߸�6�s �VF?oW� ��},���We�Ib�]�O�8o@�OR�lQPh�1Z��0� � �0�Ȼ��1�/k�yi ��zb��kQ'_`�!�_X�Z�	0�݄񃋭n�ea�� �e/�.�7�u|s��W�~	X�w�J[ �uk4m�2���'#X�����gۙ�߫?W�0�.h@Ip粅Q %�n�Z�)T�}银�>��-FgN4��>��!��?�xM�&P�,8m
�� �^����z��9�f�DQ �`�1�_���d&N��3OL@�����D�ui���������@��[X��?��Un�/T��*~��\yK.��G�х�"~�-/�t��FA(�B!`D"�"$`A��_@K��^�%�hŁ��-�kKq��d��t6Ȁ�@;��(y� 4�2QI�1x�&��Lu0�_�������D�0F!m�|�����-W?�+C�G@��!j�aj��4Ӷ��p�3J�ß~�]�Nۺ�C��|�Lf����gd�S���3��z�`���A"Z4<=u-6~�l'?�\�~?�pÂ1�1Dj� )oю �Nd"���+/[!�[˳,��Η'��I�b}����v����d��[��@�@�1��1*�@����P� S�`�G��p�� �7U+�%���*��S���I�|6!�{���W�{���АD�J�}���G�L�u1˒��[#4^���Y�Q�>u`���t׺�'��\�B�~�"G���_�H 5�{�)^��c Y�CL�)MR�#+��ҩ��[u0��{�9�������1\_`�S�<�L%f ���nwNH� �,�gN��D��D픴��
�I�Q�n�* ��{��X�1S���>5��l'\� qQ�,/[��J�qRu�D�װ&ȷ$J��<)��F��߁8%�@`"D�����O�a����b��ȁu"'B
葻6 �'[(���@v�8�t��#�D�n�� ���鶴k����)�1�@簶� ځ�:)]{B�y%�wm��̫�����c8C-'
Ѵ5r����P�	�h5O�c!8$�6TE�j������L�$@���N�����_���g�E��Anġ0p�h�c���~�(lW������U��Kmg)V]M�DK.��8V�Ŭ�p�(	u-�*�\@%�E1�]k�T�J?bNX)���4��r�d�4�q��,h��W��)�R拴 2-FRf�O�P�����)[��O�l'0�!�5�s�Nr�0z�n�ۙ��e��'��pg$[ћ ވ��ϐ�������ET_.���,N�D	��/3v�KwMv����2����> �	dex�&YO��ŘȝVe f@"�M1I �4D)�]V��I>H/�E|�����SB�\h�Y8N����SN�w3�,_J�/<5	[��J�UX`�9+Ov��P��2����Ui	DK:>zc�>t�����ս���1�J`x�c���t�������^�_�%}��G�'>1ʖumŞ����4�cx܅� bs�uV���HUB�A�]k��	�G�h�-�� ҽ�D�{[ �nu0p���F	#t������� ��g��q`R��\�߿!PՐ�Apk�[���p�q'J]E���@�l&��?P��V� �H�3�5��t�����	[�R�:�����s?�ր�0�Z �u(���B�����x��XN��w�g����5�d����Ư�%�����
�W���&�^6XdF���������>OnK4� �uU<(�m��A��Vx-Ոx� ��B���n�;�4�;M(�Uz;{X%�=ߺ
��`��;&*.����ͨ�Z����� ��@Q6YQ*)=�	�T%g@��OX�t�����Ϫ�g����H��4 �2�<x�J~ ��m~4�ꄡ���+q2�!�1�6h�S�u�p�bG�X5�U��[(��Z͘ޕ�� h�{����S�:�V`�����������S����NY�-�h/�[���z2�X}VV ؗUB�"r���\+[X6R�O㌱RV8^�������P�aG��?�/�u��#� (qG��y�~�@7b3-1P^�'x 2�X� %��H�`g��s���Z���	(�fX����u����N���2s}���)WO��,J	U���u�l��\+�Ų1���A2�eM$&hs����t;(�V���7T�Z����Ƒ(w �����.a��/�	[�wщ� �_�xX�>���.�8(���Y������!��`��b|1`�X^�&)�+?H�N�6臋��]�8�
��ڴ2tw��W�TU(O��
�>*���)�lv��XIj] qi���/�P��o%������ط�����*¼��)�-�m'L2�ˍ������@��S�r�3�[?����0��5L����N#�,H;r[���o�=1������d��a�^���0i 1�5WbDI!H��~���ꟁ[��Q�b���R@H_'�Հ4W�墟�TAh�s�]����"��}u�E�g-^� �,���(In��e�}6A5Rg�������Ċ
Xt��g���g�.����@�%6tp- ��&��P��LR�����ί������ez�`2�Cw6K�+d�̃��P�|�-q�/���;��� >O��AhP?�eZ�@��^�,��0�.���$���Fk�lA��>��󪨐;݋b2����%}^���=�?}��E�w0����^��v�+���C6dzST[}4F'h_և�<�١*��lkG)L���	/m,#�.c�;���<S+�>'K��&�Un�Y"<�߀��kP̟ڸ��uP�Q��<Q���a����1olV_�14�@��}=��t��zzp,�.����2#4(�³e�h�&؟W�ڽ��86|��d4Og`5D 3'	��o�z��_��P!��xǅ����)?�j�o�_�B�Qef[�n�V�?/S�q՜)��1#��|�Q݈Be�=O\�H-J(� �/��T���d����h��ؕ��C�]N�o���X�F�tKַg�Ρ�bT�%�g�G�Ngi;6ݿG�!�3Z��6R���	�;�_�R�HJ,�EA�����7PM��_����od��1
��,	�h�#ddW�<DFLWh�Rq�m�T*���V/X-�����LID��w@�X5��-��1щH��(c���$MZ�Yr&����a ��%���I�� ΐP�0Ghi'��!}@u(G �Ao�
��:�h�NM�k��	8bu��H&�0�T��>B{�٬<m�50�h�d�ސD�3��f�.'�߯r��be��q��>�>]��)�V���v�I����p$y�ӻ���I8|v�L�z����R~O���&0�{�Nb�A�H�0��-1�6���	��>��1^�W�a�R���h�*|HY�~������6*�o�P�]�b����[�	i�w�w�/V��\�S�k����[���a�K��y�@WhSI	Ar[C �D@	!��^BqU�m�g������-�<��y�����+,�Z�����1�y����	���l���W@S,�b�7��%���p�|��.��O��^����G?O͖��$��Y[�6̹���j���1�Wv����%�X\�a�4V��2&�Z3�Y��hҢ;���_���sB�6wt7^�בF!+%m��VxZE�^[�a�;��i^�x�!/m���C��m5���l;0�)R��,�S���^���\*��3[�24�����!��_��A���I��b�� ���0/���t0c����~*҇mAx/����~�B �)ý�N%1j|��A��o��O!{_o��]�\wW��X�������|5x�*�/��������)͖_}#J6��%L���K*�Q���k)^�<��&r ;:s��^��j��}��KрN�j=�/!�����J�Übb]�o4��ԓ��a.��ܽ�~�q�rG^��M�HL��6P��!���r���}~.`�7�>�P�kGh%xX�.Ԃ[�o5�w�!?��`�;��L!���[RE������Ut;��h�}�D���3g���[|�m�%kW���o0?�Ka��\B :t���H�h�!G�)��~�U�⅗[�K2X�S	�B���q?˻���v�R��V��9;�7����1��s�Ma��*���	�bD���׻c���~2�I��&wO��imU06��\`s.���4��ە���7��U���{������z#n�e����`.����	��1`��P/nX��!�\4�EL��-�+1;�d %��� ���u/BAd<8�	�1� ��|@m?)���@��B{��!�R ��>�ܑ8��D�E/��3�]j�bj�y��/)�!�s�d�&kݓ�6�˦�@�".���(yH��K���K��cT/�U�	�oa?����ʁ� ���YÄ3f	Y�Y��&,R_Z-����Uh�O�wu ��)\v����iUՉG6����Ch1�~\8��S������V^�t�˒5��)N�l���]����C��f�!��~����oR�͉{���^�L���Jͪ �7N�+��D΀Y��p�,�������Ұ:$�P�}t&;�5H�r��Zh�%酥$I#9�z�c����d�ڠ�3�0p�<�U3��������\�P���������(��O\JO@��* 9|+S�{E���1/�[p@��c�1����o�L�h\&'պ? �!O�Q�4ЌP!���$[��c��q�ր�t1�7�+�! .�J9�g`�fh
{A8DJ�ur�*�#�'GN�<���;�)�; ���R�2(�5�\��K^h�=t]̗3K���Q;��%P!;\Y����?@�-Bq�%��'eT�>P�2z�^�IM:��j�_��l�?����hZ����_K�bg��닯Vr��-�Cp�D��4-r���s.P%��I�����n�uV��� ���j����P"���T	���d�:>�{�L�x�g�3�
����<�&�7E����aIZ#��;�Q�]|+k��)ѷ�&��ɅI�� L�kQ�������?2"q������m�;�섆j��Y�l���K�{�z�^K�.���P	wp����'��۔�_"*X�Z1�����4T�~���m���*.�W�'[Y@��{&xM隴p;����H@���M�G h�ukZJB��_c���(�L��	�U��R���"@���a.�9�8�H�V@S�:Es��;P�-�Ԙ7(�p2W�z�&�
�W��?�<�)L�/J�F�޳��G�Č����P��0�Xߎ(��?`:h�Ddb^�Rw ��UKi�3��A1�� �/)� ��[0��`���Y%Cus[���~1hL��k$�ↄ�D���=7���Y�X�{LpM��gy��W��f��`}n�8�7f0��KI����<E��-�5z�v��1zT[ԋ�k�	]��x��E;zo�B�2��Q��YfQZ��@oh;�R�V�@47/�:���	��:�p������)���	]�|
���\�e,��n8X*����n|հzN��
�-�K�]�xE+��S�6<�P���2ؕ'}�q���RK-��a!�� �ZP������fR�?������-�ؓ����S���~WO���h�w���}�y����(L4�`�D�;����nTX�������D.\h�5������,N�X dP�q)��J+Ž�&(�v'�]���ƾX%�C�]�	 ��i�Ǳ?�������h�}4�AO�l	���=�j�I0�!�|�\ ht>J �v�ś�_ހOq�;1�^��l� �`�h��H�+Vw|1�!�g�*L�Ҵ'��yF�$���/�������*�`I��Mw��.�"�� s�\��AU�|��t�������!�^(��1�t�(�*��[	<�e�B�����S�������_��HO�E`}�Q'�]o�I�UǇ��)�xۀ�C�����H�s6�zW̽v��]�n���/�y!�8�����b"�dA�jp���P��`���7YX,�k�UM���C�x��Œ�Ղ�y����S�[V�a��)���-���]�H�f����@߬aNi6�	��d����iE	2�_�!�/�'���d�����n>e.����1M�~M!O]���:A�?�/ ���PЉ���~`�@\+Ks���R�5;����V��{�����f�$LC��1G�%I�����%X߰��(�6��'���C�Z���Y�e���һ�ʨ�N?�Kb]��B�}�@IA�EQiK��w`��w���Q ܤ"a�vcv��hnEq�z0H0f��r�; 	�'h
�bZ@;W��O/D�Gr�^��X�$�,C;�+�"8���c�@D�:���,Fg�	9^-H %� c�)_�4{�d�,,ϧ�(R����_�I�	ɸy����{Bj mJ�%U�MN�5�$���B�(��
U�ױd�9['v>����(��}���"�)٠t�`Y��;5i.���w��6�=���l\���z���O�_|�96yj���= Gǅ�!���LFg[�<z�����^O"-�A������	p+�'��	�[1�T�#� "FA ��P���s ?���.�pTXv�ѕ"�^*�΀�i��Q�$)�Yu�59��!�F�Q<	�}T�U�Iv�v�����"�59��Bf'�|"y��,�|&�V{�i�I�#i�Y�gj�}��h��*���\��Q�/X|i���E�(�u��況����
�_��C���S�q����V��\]'/�`�J��Ӫ����W�I$h�`쭸VNT�*ƄW�엠�0hK��K��ե[H�hJMw�8,�n]e�W��?������YǇ��Q��]��^�%��H��i�y��H�����:XQ�ʮ���Ѻ�^��������%}mU0^?�T%�3�v�	�B{]p)%�f�F������~���Ԁ�N���p|�����	鶥��Sh�$��9PV��z$4~�7�\��N{ Ȑ��h޶uR��hY�D�-αx'<!���Q�d�������P0:�^�ʷ	S� ��bi)�/l�g��[|x_%~VV�l�:�:�gHV���Z`$I��7N����A����7N��{�|����ı�{�c#��W��w�{X��a�])�-r��@
�x���9�X	 $Tv��a�:�n�n;f�$k���YG���%��pý�7���
�&���A�� 3(XZ��_Z:\�D?d5�xӀθV,sF%�)�}�ع �lZ\��&F�L�;�B%�_�5�|�\���-�/�y����p�d��|И���ܐ������:�F���h=u�X-�z�!�m'�����4Y��P��"=�e���G��	�P]��� ��+���5Z����mj���Ac���0]08څ	��iV�;�,N�N���)�>�����O�0r��}�M)ڒ�b<`�.2$ty�����+�1ג': �G��9�f�+OX�Y����y>)oڊ�v�Q
�/3�Z>U[SԉН0]����Yc���)�B������F���?O6wC)�cz�u"d�����w�YU���'�r|�X�3��ńj:A��*�h��t��[ � �0��D_�ra�M�R�Y����w�Ȃ'7	M�j��!EA,�Ni&N|�~U�+���h���_��`�u
Q0�C�_ ��GJ!�01Ɏ�R�p��>�9��e{m}b��G	s� %MX$@)�N����~`M�*Z��-b@�1���ZH/�2�`�"�;�PNזZ�b�RN�'"K�1��k6�k}&��7�b����1��92X}N�5'yq�^�<����ӆ ��I� $)�	 �̊+�!�,"h!>.$ �f'5~^���%:�k�(��{?GUh�#��]�	� a�1�dL)Q|0�#dhZD��`�c^S��+\/�V�#�Ȏ�}�*�Y��"Ė��%�D.�E7�8p�J�`G��S�@hּ��{��,�g��\A��*����C�B��Q�7E'�����W�8;�6^��c_�9;W��ȵقc�uT$�y�	��v�V����ᩬ,� �
dvh/$g�$H����D�G������hn3�i~Y�^ܟ�	e&޽���0}���(ά��%W�w4ǔ�%��b.��pP�E �+"S��p�#� *��7�O�,�;@~�!LBbZLw��e-�L^W7�`
�bY ���SX�%m\��1f-%��g� �&�L�(��ԜTP����[�D�Q�����@dQh�*3b]���u�P-��>��4ah���[�uRݐ��u� �~/ ��"1IɈ]h��h�L��NX,��pu Q�bV.6H ����)�5�O�Y����=l]\�s	<�����כ=��>��C�U/0<��	�5�+���h�W9��� @�EzٕD�N!���%~a�{�p�/�ox
�����[� ��r_��PJ����XSe` �Z)ڻe;v+��'�D��&R!�Q�ɭ/����!k�³N8�GN�-m�y�W�Q&�HN1���o�7��z'��v��Q����'��1�'
�mۜ� e8|+�0r4����Mn$����2�`yj�
A��!�&A��{c|H. �^]g!�)���<>|w$yB> ��*��Y����	_~��^�t��2Q��Ȣ�$�_�z`���+@�_	`��%���m���u $�bUy�W+,�Sa��*����(��p/�%�[>�7�ѥ��[&X��.ǐ���֫kL.�|}�U�ވ�_����i	!cSR�l�'g�)�;��!�K\t�%V@� (A�I z���4b�a^"~�!�>zԦ�g���Ft^	MB1t����T'� �w/%5��0�3���E��']�P���"�Y]F�gpgN�!R����l�(;/}��g��qp&FE�z��EZ��
��T������v�3̇ ���Qz�	�o����Z����=bNqE~�$y����_L�c��, �>�JM)�� ����}H�]U�hgO`#�3��ؠ[��Kٱ�+�=� ��� ����31U���� þc�6�&K���Y�ޕ�Y��X�_��~>�b��I���$/[I����I��IrNx����?u8�I@�>r|O!������������±r@�V���Qzo,섥�D��|%L�EK�%{#q�G`��T��U:q�32Z�b�YYUb1�+}�Q��K�L� �o
�S����գw��Ci;B�-V]	�TUQ�Y,��+1�����/s���+IN��D<t-�GG(�	�<��� bci1��!��@���	� �-+.(8U�� ��]H����o�2��u���K���pu~����&@�l�POJ�6 ��{�K�%Z�(d�����?����ώ���J�!���=���^ƨ<J靆���Y��Z\�/h����3�|Y��g`>��h� ܟ���[� Z�?`����t)/������2A�w@~/��Eh���<����!�X���&�� +"mYl]�y �!�_��K3�%��, "X\1�%\�w3(�I�)ؿ�{4����K�V�ʩ�\��L *��P������@)'�Ynh�.��`:�)�*�����XL�s�+.X�~��^�UɚnB����֒�kWZ�R�������p�A���6�J{��A�^$2R߂�-�*	Z�'c�����O����Y��;��תA��?p� R�Z���� ��c?���@�ï3��� ��1�"��D:�J�Ւ����9M�����k�Θiw6ѣT\���T,��0�RV|�~�	ӗ��{�a��Uv%\�k/�*�`���yM��L�
��wjQgHw�e[`Y^1�)��	��?��c�t1�� #]��ià���o��C.�}&��<t)a~A
�n�ֻr�+��s-S>�@L��\)�O-/H���Hm4$"���i@�?	W�kwJ��h�k Ph;<�0�%q�|K#��Z���g�}t��=�#@�%���5��`��mҞ 𑏀!�-�
�&�7��Ts��x��'�+Y�� �����Y�iK��@@-#HXVh.@���U1`%�e� ��R7���c����0�-����nBP�L#�������P�1%�P��v���4��pWR'K9�@К��B�٠��x��O�>�x�|3IXB� ��f���Uz�������W$-ZQV�EY���]�����_�h�;x�� �{�f�[��@1ع�$X5��-E�v��^l��������n�� h��c�(��MhF��P���'�����K��As�\Zq]�G��F�%�]Q�dSW�YJ��(�.$��k:'*��ZX�R�EoU��S�lE���@	�o����� ��jqZ|��M��P^ڂ!C�3�bo~@��V�߉s��	@$�3M�*�U�c��؈���@��Y��%�v�0��[D�c����0P������XIyV ��� 2m&�0��3X�v�d���[�	hHY���q�(Y-H=rȂl���!6a��B I�ˀÍ@Wh�p�:bC�����m�`pw�Ӯ'�T���I�	�U��W|�R]�c�a��Z�2ŭ�DA0�_��,/�a��K��P�h����A�H2# #R��>��Z^�+��h�0��e�
ŭf��1
Z��s�h`�yqJ,���*߯Fυ�$��sQ>�W�yT�])�[��m0N�A��[�V�Bv���ȅ��pn�I��v���%�	�м8On���W�'k�x_�38y�Q�9D����fYR��0�Z(�A�ܴ;��Gl����;V�ή,xJ� �a��x�/����K �V#u�RJ���������/?��+��P(��	�Pe>�n�@H��J�VÓ�y�"�'E�}mQ-�� hm2Z���1Հ�gC����`����:;#��	�)6����2~����3=�o@`�J	@}�{�2@�g��Yz����`�P�i$?	/xLZ�9X��u"�fP��p��ɐ�V��6�E�[ U��>�O��`?
)�1�W��.�R*���IqP}D�!R�%~S'��Z.��[�'B̻1sq�/�/�_�-�?�'BB���-<�{=KtX�!Fb{���OY�\����-T�+��W��0Yp	�� �U`�?���y�E�յ�|`�N\�O ��$�j	tY�>�ҹ��4���4�;.@1��vO
�u���O�����g�y�����(��{d<�}�,1��{����)�p��>7O0ҁ�a|<w���8gB���o1|�@5�/�l���]����#���'X` 5b	���[�Z�N�;�+]rcҐ)����,4�]�����%� 2Q���/A�U�{l�>�y���4{����׈E�o�r��!w�9�H�~H�K8����0����d�M�@�Ҁ��f�d������j*Y�հͧ�e[�W oSh�Z>k"�՜���h�[�-�-����JP�N6c|>�vY�u3n�*�9��@h^\7��*�Sx@�z��2C׃�Zf跨�π�e���$m�W��������ŤS���&�����j�(���0�X�y�i,+���
5��-�.�%�J�J�`r1)T��(�Zp���q�m��53@�4�ϴ�,���q� �l�=-)`O6�4S'	��G����a]gn���!��]��T"iJ^���pJ��|��	�uo&�2��=YF��4=����5l�9���'�;�B���KB��q��e�)��:[��r�B�����B�GUO��|1��t�b1��^W����LAR�4���?a�JPR.�����|�4�/v�3��1��a@�_!N
 �4A�f��e	ҌZ1P�1�L�(�W��j*�O/V��J[��&L��H��S̤8�	�fXw@.e�(��NUё5��ZA�/��K���^�	-�)w'�V5�`� g-@}�XIz|@�̚v��O�JVcK��!����e�a�Pb:�.���N)؜���dz�w�T4��]U��x�m�r�,
]J����g�v =��蓪�\��É��ra�.�4�z���#uY&a�2^ N�$�(�'A�;E���������E�b�,�_ȑ�O%�8��X�M�i?IBS�@�U�	�A ���v)�#����� $�����W�w��uNZ�!�V���}��'U`Z���M �q�.�YHkIJ��{�a6�Q|�>M!] g���	�y���Y	�4i`�� �1��[�v �}3=�#'�Y��U&HR�]0� ~)�/��兦�-~�"������r�.���¸i	��1	�運_d�S.�-�H']�)j4�����BFV�ʧ�H��;�>J��៓A^��cމ�"�fv21�.��A5"�[�νo4zO�x gDE阷x~ Q� (�Y�1 f����|N����t�,{B�����ذ@�0�^/�8�Y�D��$Wc,��h�xU�����a\�-AK��1bEr_ǹ�������.�FK_	���ZL1ȐP	�P�}B�k?U����SI<�#�Csw��[�p�-  ��qM�)�ɟ�lB/����<P kOR�I
�`<�~7�GI �yR�HV�ĂR�܋���}G��B��'A� 70���. >d	�!CLV�퇗�W���cI8��R�g����7f�D��Y��˱�(����n%�y&�	�)tM^	2�\�/��l\Tq�uz�	�p���!��:E � K|�8-muO�R�\XH��}�Q&+5��mW2��- {�?�!�1��vW�@ �Y�����G^��|c����0'C��8FJ1��ě��[C���U�jė�!v��z�-�L1L�������/�NH�a'�D@Z�O����V$~n�	�K����W�0(<D7� �s�	V��!0� ��YJK���`���jHՉW�A��	6hZE����F	��v,w'�<]h�V=-��T�:/W -�%�X\���>�5n!����-�^D�6Q�V^A�E�՘�6�a����_|�8'��i&9�������L�G �-e<�y1N�A�鼭�;�����!\����$�8
v���A&k�ܜepS� |.���`.a��D+#p��?WM��/׾��"{�h#2+��(S�@�yt���0�9=���O�\"�`���'&l�a��>1��e������nÒ0˗���P���_O&����Y'�t?�����'�xQƌh�	�B�mR�n��Ԗ�pov�$*�����^�GD� F^W�H Vf������`�Dr#)ݏ��*:�.���w��Q"��W���qx�ִ��sWD���_} �P�Ah(�A$�x�-'�[�Y.	MoE�Ѝ� =)���j���ZC	��E��1�1]�	A�V�I�(���}���H=[�,}�k%W�G���GD((���_&����t-� ����L��-!��os@ 3+[��IBl�`	�F�u�OC����\:�!OU D����霞�y����u!�5�T}�E^1%f��x0D#l8L7�ײ�O�Ҕ�hz��&Ѥ*�z���~��f[��	�<�	�3�Ha5 �b�x�؍��W�i\�_�1Q�^
��8I�)x K�A���8�������Í��S�ȵJ�h���NptE��WU��(��{Q��k���zR(��?5E�������yJ;���@ZCH��\i)�a�Z!`�7|R91��"%Za-������:I )hR���[�4�ڐ\	�P�^�O�;4V"���D[��=��Y��^�̘j2�(��8�l[�(�k�z� ަ��<�����J���&	� ��^�<~]^��YXSƅUT.*�7%D�8fp�?k��˃ J@_��$G_���A���	���tx�iN�(p+g/_bv�@�0�h�uOo��XOVȍ����}���X�dR
��:~`�rOFL�[�p�kT%����^xV�H�iu%)�q ��Â]x���Y��
a@�:�zp U��ϻ~ s���	B*w�1��\�r &Bc!�醕�A aEMf�\K�b	��\� (VEP�C1L�@�9@�.��>��%�h-d����� iyv1�Y5�)m�c?�P�-u�!�+6�9��k�h�����H%��<�q��AO1g@�bw�Py�6F����	�0xo�-�� ݹ�Q�b���p,C��&�u��%y1T��(w092$�X5/	��<	F)��R��YP��^�yIe	|[��B��4Y����WPqh@]l����0Ӝ��2��J+)��
��%����Y��Wq�:�^�]j9g��"[�  Xh�&�y�UkT+?��������%�M�Ų���:N���7�V��k\œ��Zy���s���̗h��G�����3�������f��2=�b�݁�_��0p��o�\�?�"�А��`D�|��|XK�t�%�����(�)�	��^"�
�f�^$�C| �~�+�	�6]	'��?C�U��x�h&
S:h�=�8!1����i(�C�h�x�M.YAN 6�	�͒	+�wE} ��gXv�+/,8���C[ă�]��A��[�
 ��3<�C�b~{��1Lk��PfK~���(��l[��Y���u"����ŗ�����Z���%�PE�$I�: P�akJ	�,�^��\�b'-T0U�\!n���b����I(��'U_�B�zU��B	�?gP�
2�rM��Y��p�N/�x���i�$dފ�f��"�2�%�z+^�FH�^�FSu�ZK^�}ĩ�@��K�j6v 5*HD%�&Z-h�	��r@�G�y��Z����&r<��+� �D`���)��z�,h�0t[��INA� k ��o�9U��҆.Ľ����[+����Z���,�R?��Y�v�qB��R��4���wGh#XX͗V�7��?�%)�u�hJ~��&��ўP���[;�Ζ=�h�ez���]�����H�f0�sn* SÚM����)	�d7UR���_LYWhۥ��h��
���'�>y���!amO���h@[
e�>P�ջ&+N�����ҫP텕W����X\h$�P��ӲY�+2V�j�IUg��/U�~���W��	2
Vu����R���1r��)�dX�6���1�Ϻ�Q��v�
.�Cn�����t�A% hvH -�����z���"�
��� c/{X��d��#srPA:C���q�C�i�J���璀�t���`GuKq����:�S��t� ���R M	� ���!�"�B�p�X�^_x�~�*\or�v߾����O������)-��w�e/buQA��A)�^�Ih�w[�rw[
�y}B��w�	����C;15�N��4�Ɋ���.\���4"�3g�Ӿȼu1-�^^U��vC%��旮�a,e`L�Qf�+��`��Wo��	&�k)���`��k�V�8����"Z�'���RaCT)��_��� ����Ö������4����$��r[�Z3�V���uZU�]��,[�hY��Th�*4H�ȧ�<�Ka�K�J1�@�?�'GR�`�&bzv4�"���R.٩~�O��I0s%�_�DH��Z��)�k��k��Qe;"]�M�&�wƦ��'E=��B�ʂ��ePW ��(�[0����s��D.��>/���
�"��y(�	a!J
4����!I��d*_X�J��1>/ ��\�w����f8 ����ZZ���'��/�p���@3UY�h'�H_�	^ް�y9�v�s���	�/ ����)�\�j��v�Y�̄�XY���_̆P���X��P�+̪1h������ ׇ-h�X}�}9��:�M~�`.{`)J�c@�5�[a�oz~oVD� X^��U���0�j)ր��Bqy�3c�;~�A��N��]�yO4ۻ��^�N	�-W��0�k��B�b���w�'N_����0Rf��]F|U@
�I�l�9@��BN������d�x�_2�U�0nm�钹4����''�C�B���)��1J6o	���6�( ĉO ���i����ʞ�x��g����m+�b����>�3�Xqz��6&t�"/W��W�h�L%W��C�M_M�p(�^c%�:�a�:��A��_�&Z�*Q3�a0�1J�1��v��k���v@YoN�H 4�Ѿr�_�^bP���=6�:��������Z�����Z�r�i�����S�A�&�g�f�1����``�-���2ݧ�^u����R 8E��h09D����)�A�T2Y�+�.�D��ys�͚d���z2� {
�$�$�/�����hOr��2&0~�7C�5郿%��JW���_�+�?7�6��/�|�o.�z����2�A���ـ��
R>��%yй}h���%}�<I�Yr���]B雙�!��h	Z/cN����83?�՘;�k�:c[���{�Bv�Bzu�zz��^�I��G����u�0~?�3�{{M}�VO�w�ł�A���X��0b�;�/�#1ý]pJHI��=����a���T�;_�L�U�iE)���i����_���bQ�Ar��� w�f'���$5=G>f:M�ԛ/�#h�x[�)�:��˽���
Z��I�\��(n��!�)󉭠��avz(XP[S��Ouh�4Q*%� E�Q-ւ2@GB����Yf�H-�G�:b��1�`�v�bnK���BZ�Y�{�Ү���� �n)0y1��j }M~�iP	��uӄ>w��J���6M]����W ���̡���lJ�����J'���H�f��}`��FC{� ���p��_�V��ֿ-{0S�^�#�ZA;)���^'H
�N���#�$ ��2P�.S9����w�3�c���h'If�?�O��-}^�����o�Uu5z(��Կ���ZvM}t'Y��Q�#�F�'���ӽ�GL�@��s�����/8�z|��_!<r�hp�%��ܛ��z�;���wN�4�G�c)[r\k;�8X"%}޵�:ً{���k�XM7�%2{��Y �50l���/���(� +w��a$�h�Tl%���G=���"i([��!Z݀	t�g��Hmh�0��_m1+[��.���Fp$�L��X3�N���_y��V��[6%�B6_�+d��u(�Q�rcL4BRNm�*�c5��<�acԿ�JkT�^n��p,K�迣��8�;0#[�y ΂�N�`�0��/-� ԃ/&H3Еu��sE0�c��@L�"V��A��D ���Z� �fR�E����b���;������
��O��E�j�#N�d��-���P� �����6��C��>�������^��-�@�l�Ed�|ya��CX-g:4}QX�j-���y��R�c ����}H0!�bU��sۘ?�]/�~�!9�g���n�Ns���� �5
+j�������m�^ٱ�/�՘�p��{R��Nih�A��J�R�X��`� �YN��fTA��6*�L�G�x\\'h�F���ga � hfkX�
L��N�<�P�A�:�د�c��,9%��>�A*���L�����I�] �qeO��C^�PA��, �B���X��ɗ�.���@	�1��Z����O!�)0ϠM�{{|V�i�_ 3	X&PhD�qg��_����=��ĥgV�V������?�B鷈�/���߃luN��=�`Az�R����1��CO'P��u&����K.*Qd�&���]M��h�� O���T!m�2Z9��xK�6��p���J����^YI+�L�_W�P�%ȉ{�ؼ�}z�@уi]\ �m�ǖC��^�:0f'$Z!��HQ2z"BցO�;�]qqY)w\�H��(����IRV.� � Q���vcG��P�#�Ÿ�	�Z�_�yEC{uKf�9p��k����	 x���'Ar?���	��pp9�%BP3I^�8	Y钌���N7��I.4��O�����J��~����	�$��\�{$,	�Qs ���$s���Vh�1�m]_Hv�&��f�A�]~�H_ӡ> �SB�H�Ms�)x� lO���;�@w\9��y��ľ�:�� uU!�r41[�D�a���q�!�>�)�|�1��\}-�X"ip���/�N|�� `d_�r|�}���q.��,u<uBz�ΫS��d1Ƚ`-(c �mp8F)��=$R<��z(������,̦tA,G$��G(Sc�֥��QO�#b������i�K�Vd+rw�B�Vw�+wiGYw4�S�*Z��W��A[�a'��T_������T���VÏ�_�m�d)��/�h�h�XC������'j�X)�͓"������$sT���������^#(�I���1�?O$0��h�E��Є�K��l���5�0�o���l�����-��D]�i���$Z΀@nv,�k3�V.���Rh�0kJ����O=%�-�\�&�2��YX/d;8� 	Ng�؇b�U �4�P�� Q,)�_�[*k��V\�d@��J� i�~��^#V`��H\y����� ���z�/tK�<�4	���H5: �{.7���·l6o�ڸ	�)�ڟ%��~p�EY�U �V�.%#D)�������u����d
M���A��Z���$���CE%�w���`���ɦ@2 ��h�d��ďt�jq-�W�b'�-�@A��nL�Sr}fuH�� �0�.5�8� L�A�f��]	M�{��vL|�rH�T~j$�B�q
Z���"1�R�qSm?��QxH/�)T�4�����
���R��5����Tih��ut��-�#�|J�-�גh0�����,N,b�]�;�?�L
,d1��� �G�&�Q������ӈ�Y�Za*�V��ϫ��PRo����u���[]���ω(��$>SEAs��B0R�,�Zp�Iʀ[h��������tPzys�J�����<a)6�y)�� 2ZQ���U��_Đ�U6zF%x��S��hW�fe���I����Q	p�oMc�{ �Ud�ah|��}��u�E���`���4�ޔ��l�𑫗�'��\4^0����MĨ�������[k�	t�uP���ö2��L���Oy	��X�4|q �V}�`�1��̈́wD����'&�cd4	G��&�Bb%���AU�:���;�O����tZ�7���P�2+WQZ����#pُ{�1�v�������B�=!,+h�~<`lY����lT��t�."	�7!�0�	�W �z����Q1���.�8|ϻ��-�6�Qx�>��XR	� ��Iŗ�1�膾�E��[���j�����E0Q�}�
?�ǵX�	���ߨK�:����-$f割����'_@\�'1V�(lyaC�e���Ey�����#vI�L���k�b��9g���QE�Ag���*�P�N{8B�
�*{"�7�~�K���|��4�D���9�`F|	�,��"'�C�
��2:���;�Gu��F�����c�0�P��u��'c{g�~1)�ߒ	�l���Y��}@O@`�M�r�>hTI��u!�bA�O��$Ā�p]N[��X w:�,�r\iL�h��Tf`��G��<ο��Yd��#� �l�tB�ҽ >���i�n_�0\"�y�&/*�z<��6�aE�0�� �×pf7o�� ���M{��/ILm�����A�Z�Ȫh��� �G �zva�woa��W�]�N��Y�g�h{?�l靯�?
d&�J��l�DM!mvw�y���ca++q����%Ǭ�pw�u��H��˗΢?��-�܇Z�}�p��(����S��K�[[I�t���4��)��3�O�4�ُh���}	�J��K�� �R�'(�Z�� ��{���>Fd/�����aL��PSW �t&�v��
	T��K�F�}��h/P�oECɼ�A`�g�#��`<+(.1���h��h	]P��' 5�U-��,��]%P	��'�Z`z�w���1� �P��$l�3���*��s��,A{��O�/)�Z�	T3�7�d��=lM��HjP��1"(#��<^>���]�1%4�y{�&}��>�(��z�ewӧ�F�Ϣ%U�h�po�Eϖ��Ċ	X��4��V�>e���%���ML�ejٕ�nA�?pM_�珠�h�p���Q��qvi֣ɠ�M�'tX��hY[��rk�Bʀ��@��0���:i+g��/1I�=��z)Β �q�#1ɽ���y�Y�j���X���Gn�p�w�8��k���h��R逛�_�닦��`P���ȇ��`�^�}vG���6@�K	<�ꎤ�B]�P��B�)W���`.Րu�8�8a����2g^P\t0����U��)}�5���*���`��n	ɻLt_d�wG�:�	W[�>C��_�AI��(��~��Y���q��h�DlZ��&��@�͐F����H]��R�x���j�Y��_�b&����x0���y���:FIGW_v� �%q}hRS\�
W.��HTja�� ��(�0� �����Q��>��2�LU�A�	*�gE^7��w��'~6xs(�Uџr�#y�+��4�xE���� ��h�{_F�mV<���=�k*�
�	��Ҝt^�������~���SL� W�[S�yO�u����@`0���l�6��)序��X2qE��Yj�)�[�|QR��*�Uŧe��j�H�k��C Q���q�Xb�T���*N�¼��8w��=a~��'�p�t���S�)�>v�:�	�lTR{��\��0帔��O����bU��J�N_3�69 D�1R�?Q�&��.�1�Nڗ ��Y�$< k%F+W-���:	!��ygh�m�5�
2Mu^eVG)w���~�W�A�K*�:�^��/u(��u�h�j��Of��ނ�Ya��b�rg�/��_�6sBlA�f��R> ��2g��ω�Uc
X�ʏ)�	*5Qّ�!��;(3_�<t���Y,	�6��#D^����O��܀Y1�)�RS;P�/q�|���W�3O�FM�1q�z��o���������#�G�NJ�`�#$W�3Y�Qb)���5H]���D��ˮO����!�,�d6�i;qQk������Y"��`�;�Q�+�l;���%��G�R1X�lځt)`����Kܮ�M�\c���[^ �u���W�=`Z0�ׁ�-R�gM#ZN�{�i8p���H�a�b _�����%�A[ag��.رY�+�]�Ϣ���+�JM�Q3�*3������-�1�	3J��H-Z�{�ҥ/�C����	.h���B�9ڠY+�$@:B�HlcZ�!�&�UR�P�O S�u:�U|�t03)��A�%��� ��̽OE�h����ypf�F.nl����y,�`�_φ����DÀ�XN�:��y�%�ѝ\�@�ڼ��U%�и ��(X��7�B��D�n���թ
���q׎I���}�-5��GW�ԠEm��z��Y���*�����@
}���lОtv�Ppw%��Z�a�8Z�|�����%�֭ P���m����۷*]��Ț��>쭠�'a����B؝�����h�Ee{Y�G�}`��_���Fx��T���y�<b#�@���}N/���٧	.�ş���z��vn7u��h���J��j� ��~�]�T1��~�.�<��dS�����
<_Ӭ�����%Z�f`�h.*�Ph�2d��{���P�ryGX^/	��h��*�zr�-rN����h��h������Y�,=�� ���`GN!�sc`E�?�L/����ن6,�Lh��2����
8��i)��.����0��X����W��gZH��G�K`?I�`	��H!�L����G���o!��E`>�?�|�U�Ďh�� DS)˯�S��1�~H�ow`�@-�v2}�����p�����4'r��� �_��Y���Id�'p���A�����b 5���1ؖ�4��̰�XS �IH����ē��,�	��D?	� �x�>;�w���"#��DY�d�~ٮja{}�:�H}��@3������l'0���M��;�
��O�P�&G�+�����\�� �Q��LT�� �#�X�.-��t�`�S,^��U`(ȫ���:��$nm0�)wW��eу�&��Y����XQ�tV�,;��_��q�h��J��H�9?X��rL1e �53Bp��iIo#�A^>6aQ�A��@��L�j`�L�X��$O%�t`�.�{��XcuzP\�^=� ��fE%�X�$��Cð���
��ݘ{����tK W`h.��%��v���	1o>�o��z1��a�R�fh�}0G�z���Q��uOp�'0��r�}�si����f�Azд`Ƚ �{s��M�ݹ�C�ֺ>��s��ѷ"�@�`dC�uvnd���a������L�90k�%��,�(����h�O!2l*�/���-=�Uw����{ KR���O�H%�|�T(E��L���%��ş�55�b-ц u�������w�*�I/xU�م��.xChb�W��!�(	�`W	����wU����m)j�
�L�KB���tD{��1z���,���r�p�v~л��1W�����%hwY�B�y�%��-.H���W��=L�r]t� <Tl�{z�O\ ���wV���kԱ��s��%����"p*�<��!�Q������d�i�%�,ʴ	��	�^�XLq��vTp��G����t/}����{���h�1Q؂j/�X��[�C��-F�o@���1��X���>P�J���8�y���x/;�b	Q��G�h]0�!�h83vp�
�@�iY.�rAn�����������͹���D�}0���]�B�����>��J�Ǝ�����9t���7�%���M)�@,X>&k?$�;�_7���� M����(u���Y �Ŵ����T�o�+��5jLxP%�v�O)�@�1(��0��n'�2t�O� ���Q�t�3���b?�}��z �[��M'n1���G!ZJ�-���d�J��-�!�Z�6��jO�e����7�n &�$A� ��C/J4x8�;t\�P03 	���{x���Y��!(�$i�{s�cU.|�ӂ{Հ��(�f[Qh�ZX�`P}�@��_?I}&�(����0�����Rx�E�E@��?�:��0��6����Ϥ�c���ȗ�P��P�������k��d��'+=�Kr�9z/fh%�!+'X(���|�D(��^�|�[H�2O���PJ��_^��x�%j]ȱY:�n��OW �k�2j�@��H��he~�L	<�X��F�-	�"�Q��r���w��'Hf#?&��L�Q��۲Y�yP!��o\3Ҳ�pcݞ�K�CU9:X0T�uyGV���� \�*_X�)Y��zpVg[�u��DP�>��J�53���Px F
�fr���H�ˤӺ�{ӻ��QJT�h�Sh}'�:�����Q ��/���b�%!�����(Q�j�Q���n�x	��1z��3<��!�_����+����V�q�����4�+�	�E`+�D�X0}*]T�F�'��\I�HR���[�49�ܭ��p  -�h�y�x'��`�������\^RV̞~�V�x����R��<�7�/1Jھ�"DĄ-�d�)`z�'��U��h߸&�����=�����(����������xN�J���)�h5;M�o���[*�n�ӑ�������b0���_$��")�pŉ�ĊNX�$���h�.j^�����,����� ��d��X!�1���`B������RA'�b��I�Y�(��4��"�?�������w|��Q�<Ҏ��/n"W�8�!��F��	�D����1^YW �q��B@޽�4b_�� �GsHX�W)�-���Z���4����B���ג�Dѝ�@����cS��# ����郍	��'ЉZQ�;a�p�؀5�l��w��^���F���������7Y��i}��@��,F{���KiAZ�1��+!8[Pp+���!c2OX�����p����<K�%]��Jù|,[�s@/Z+�@���Љ� ��)y�%�31�.��y�h�w���rO�_z�s,k vHV�);K�E����'�hj�t�Q�+�����10����t����1��B�ܕ�A�C�{1+_����kW���o��_��x���A%��b�5F�AlW�TpVrk���Cȴ�-gZ��)p.��C�r��3���zL ^p��Y�u�䶤t5��j>aR�0��i���X���=�7��sЪ���ձN[A���B;ܸ���v�nl��(�P�[�k �t����'�i�Løm�e)ˠ0~�ԋ���K!��i��+��(G ���	5��c�����)1��M�+�uX��,h;�ȣ�H���H-�U�S���Х3���X��5���~�[-����?��\�>
RAN�d� W]�4)��`%_�r���W�-`S�V(JL��^T�� ��f��V,N�A&��)ٺ�c0�h�f<u�����q�D�u�ʏJ�ʹ����5�] ��XZ�갟Ke������T&v:K1��u�?�[~����d�}ѽ�]���,�c�;2�4�H�KJ_@
0	�Y�<wEq�v�;(�>g�B�������ᴪ�͖I:M�k����)�jVI9�c�wr�	�`e��ܿ��TG�ey��� q��D) mB'�AE�Ek_���#�)�U�D��*`,�h'Ko8�ӕ��6
Zhbz@�;+d��3�0ԛn�[���[W��Z@A�01O!�Oq���t"�G�t2y� �t mQ�P���㹯\>K�Ͽ�Z�� u/��	i>.. N��GU�LQ��&X~P��y,�_�$s�����H��x�<(�����w-��T�>�0��DI ��R���d���k�p���xe��!�"�.'��9��B	3}`w�hy&&�3+��X�E�	ʜ�GPg�n�%`�-Nd�)���o��>��HgpMr[2����Ui@ ��,�y���<3�Y��b�U�BR�B�ZW �tf��`I���-V-<���K�0 �p��;��XWZ�ꀿ�\��X�z��=�Ǭ6�/�P;���hK��A�����hAr* 彺1|?�F�����-�m)��1/�C�7���Q��$�h�s��p�o�*�v���Zn`���&�9����X� n��~�X��!J�Ӭ��%E;�Cu����������K@�")����z-F��{&��/��`^(31��.�W���-�u����?�!��+��MV���.��J`��yv꬈�Q�S�Y�4���i�]�IH�P�������3M|7�β��ܕ��}�*:�ɝ@������%	oF�y���3[�/Sh���5^����[h�N��KH�?��7�fY �^[����m�t	�
A%D`B��qM	�&|�`����(�o]�x�-�c����Ր�(�!N������K�J�W�fn��5i4�cȂ^���`�@�(���'_1p�|�6��� ����C���odw��0�H����x�_����E:����.�U�1�z0?�T�R~a7M$RZ��]�K��@�#����LP6k0Z%�{���l&�H� eD�Q3a��b��`[@�����ԙ�%�Xγ��h���D�'����S�s��I3�t��ũ[��i�4*_U6���g�ʋ\Xn��t%�T�$�Ԕ	
X]F.p�
��͘�s��fm,�l�@���;�!�Y�?"��{�V����HV��^C_3�	Y��U�������b��5�/.ߡ��Mm6��"�	!����,�NJ=h�q\,b���
)h<H��а+��o�V��?/��!�h8Rn1�%t�L��=Z�@����݊�� Âzf9�5�X��:e=|)_Y ���RT �]):h*�)O`=SI�'B `@+J���� U}�^�B��3A*� ��	Uo�*h�3��'P�of	y�ѻU �W�����#/h��bF���DƼ�N���`�Wh�Nl���%z5� �S�1�[��p����`
o��B��-L�om�F s�Sþ���2$@��6Z�!�	�(��/`g�"{�k���#:2Fpjs7�\X)��B�i�ԢU�ֿh���`v�q���l��,��ԻQ�Q��d(�*�t`�+`}h�8QYA	�֢j�w�ԏ0b��6����P�y1��,�	�Һ,w�P����[qYh	cu;ug����@�j�(�X�g1�l��^X. 9E�}~j��_,]����[1�wg�:kmMYP���m=���W�5$�v���Y��p�[�B0�b5� [�P/&��`[��X��ԣA���_;C�AX�+���`I�vʬ%�|�z�����G,d��a�Z%9Jm��B	1��Z؆�n^ֿ�{!�pg,~��/��'zӛA�jJk�̀��w~�m)��Q-o O
H�O��#Z}�O�~ #Sl�-��G�̀�ML5��?.�!�5��-�L�������a�h'��n, ^�@L_A��:C�TKFb��x�	5m���p.!��_�	�邯�.�#�������o�!�:��q�� �Ru8:=�ɻ�&�D{xx�Cu��x�K�� ���TB�V���;�&����>)�rNV�1|���a�9h�I.�}ׯJ�͂[C�~�u��{?��9���}�)��-/��������s�)��A��@��='�8�y4����	��j	��Z��	/���%��t��-47`e�I��Qx]'L�@f�$��D�b�H�8.-���8Y�	K�@�OUm�|���k��n��rV��eFȧ���_:B��B������)_'[_��>�/QT �	�T���RRS�K�`r��)�K� Vf�N�ȭ�l$3O��w:��V�~u�	;2uڭ�xu�&�.fI|���$ݸ7�F V��0`K�Y�*��<�} ��	�1i˸�Z�n�!1%��'���f��z&|��U��!�[���~�
@�K~/�T�u�c�}0�,�����:@3�fO����a-�A�Si�u��^�~Ա�+�L|q ���]���"RT�;Z���{��0@��(�������-Ɓh2�a��F�_��9h���``O-}]	����A	�oA(`[��.�@���E�?�V���%J��z%�^f%�Q�S�D��V	h�-f�/+	B2]Ѭ�����-U�Op�\�H�Db�� !T�C��ye-tB��Q��)�Y�#z*���5�>j��-8؎Ǫht��p�߄�M������.�+�۸���]���!�^��'T�A<!�{��X�vd����1�5��z D����������a��B��w�k'Wdp��j�7�'?�<�)-w���F[�s�{J�^��d�+�&��B��'���fh��r"��(*S���x!S:�_�'W���B5~A!^hiրh5V�0N��;�/01�Y^�t������`�h�� �f��0E0�)"�L!�X4g�����B��'G�-�/Ɨ��#�Y�c����Q�Ȯ��&��o� Եy��&�ynFn��i�����Ph/�\��b�{!�>�:e��h�q!�,K�H���ۦ���9JiP�ศ��Z�)�:.��i��ѿ�X$�h��^��?� Z��%5�(g �*�Y%�k �_@-�l=5j+x��а&qW�.��[g���� E�)߄(�(>�A`Jc kL��r�e��{a'2�x�P)+�xe��`��@�c��!�Pb�
 ]P�6"�����
�b����&����	V$�Nעf�PuF��џ�%0�Y�%��\R�O�@(uPQ	E�vBC���$o��g> ��u�]��/��.�3��û]0���L��\O��B=>��x[���?�_�3���'\� P�-�'?XW���x��c�����v<J��9�:��������m��z?Q���z���QOT��--�VS��V��X��\�`�#QU�Û���B��I[6��<G�N�4����ؤ� >�c)ù
(���9$�����R`��w?�l�*��fk+2�94.铎�p,֍�(ӗ��NW5��ф>xgmq��`9�n��%����-	�D%� �[X59O��� �x>�����@3!Xc�Jr ������)�1ه���H`&�e����u@gT���`���90�b����5K� �~7��iN��6���?�< Q���).�2)���-F/�[�➡ld��	�~�u)&�5�P����f+���D[�t����[�n-S}��+��[0?[�no�P�h�.��Zx�^dDٮ��ilR{e?2�����s�����\�J����G���+(K�S:�s'%WVN������,ZdT��h1�`)^*	E���	|Z$�VD��x9K3��C���i�B��'T�\gqK�Wa��fZ��Xh�"�,�8�	�8�/p�d�~AցX(<SQ�Վ�Y��[���@�PS�@�x�=�י�����8��[��R�����"� a�,*�Y+AMpeRw{R�0C-VJ/Cr�K��$���D���=�ٛ<>�u�o��w!��gkϐ�S��fK,�����Վ���^�r��!�������P�{�!�AS�]¬z� �Q0����v)��[�!���dB��Uyf�@i�#���rZ�[^�w"�|�����u������K��_K��dZ �v
��AӶ��\� ]��2������	0\����<D/�v�*�¨��wu��@q+�!����|�� �5;��2������^Ʀ���}�[/��(�%��J=O)� �9?Dc̀�
�{�w(�=��\^d�5�\'nx~�Y̸�|�@�7X��`�P):�Y*��K'�E�3,�@��d�K U@�T5�k�~:'�X�DK;��]B�k Xr{�PS�!hд��U�@�P�!;�<Z��@�/����c�>�1ؽ`U:�������I@�� M\N�����ǫ�B��w0�\�Չ��4Jo��R��������6��q�.f(=��$���
��R9��o�i"�[���uAL���xp����*�cͩu�A��}Z�.;1x�C���\Po�h�@L�	��e�_�r��"B�,lh'�b�Ẍ́? �KD1��� ���� RS��,j��)��l\���a fq5k�{!?�h))[ T;8�YM'�'�݀uPqyC��V��v~	5A�y<�R�r)]D}��1Ȥ7 �/jM�Ahs/PI��@fj��%1��gk������@��K�z�����Q]Q���R�/5[��L��)U��P�q��#���̦+�O�W�ai��������xg^u�A8V��*��;!� �P�rY�?`E*�\/d�c����X�	�Y�Y]�T��f����J��:SB�	�[U�}�K��^���)���j�� V��~�|^o��¢�FА�9�1x  �(�PR��?���R;��F1q�[u+5M��v�� �)ӝ�+<_~m�L@���$Ӊ`�k?�&�!8��	��T�lJ@�c����1�l�s���g;��@����fN9��W��v^ 0���EV@�	�R &�(�jK���@ŀ1Ҡ�3g%�(��$�?��8ߩ�����]�B&��*U�Z'��*��w8�U��}K�E�:Ԯ�Jh��I~�HӁAp*yYf� h�jr�@_)�ByXu?ZU���Ä��aL����s.II�� ��5�(���?%6�v:��=�G�t��=�p븹�-LO�K"�	:]��?�}�� A�2���sm�P��c�}Q��5U���'��\\ Sh�"X�E�	Q~�2@3��IH��`V�&m�6�fx�jB�Å�B�݁ZcVP�L�U�)<�A�
�+HX� �CR~���
��k���(���.�-IH X.*�3*of�����������E��'`r��f�7|�q�x(%Yf2�F���o�t8�ʂ�ך�d�tX�Fx_�`O(H�;�	��:I��ٌ��20Z���_̔-h��q��^����=��\��;u�)"��/	:�p���3(4h���Ϝ���F}���7[�{��=��Z��H/mz~k-�>�=�I߈ ]�6��H�b���7�%�q�v-�%��Z���b0�,���D'@� Z���I�L@��O
QaBlJ[��J,��`;�ߤ�U��'�bѸ!�ĕ8�����=Z��x{�Z��ԓx&/P�"�#��w�l�#V�����܀���[fP�i�k =�)�&�CgBT��9��w��ߎ�N�~���:��B��nwX=�47�;(��8Oo��1�� �N�� +�W���^���I�K���%��vm0o2�t�B-��@}�.�=�H1�!X(R��a����^K[X�Pm�H�R�������@����pZ�T�"��s�i���	}y8q*�wI	nXP���p�A�x.�~F TLoc�@:�Q�h~$�0��<CK�)�!�]P�u��w5J�Y	���<:�(��2_��W�&�)
k��Q��,:�4�pI&�Cp[	P	0�Rl�R�"B�
�aZ!�|��P[�#�O�$���k�\��]�F;��w�|^��2z��^n����p�u�u���ɯVTc.b�4<������&�)'7!WMA�Q5���[�%y��\*�_��#.��νD�Rl>H�阪:�qb�b0�H�ː��Z��
�����fS��[z��8��	Q���
P��߰�ҀF�K�Oq��{���;��\�-LbTp�i]_Sb�,*;�P�Z�E��06�Z��&,p��z8��U���ڵX���R_n�0/ ƹ	�gw��(��i�u���5�t-v�r�Œ�ՒW�m?�،�j�)�L��'�]yE�e,F`t#�h��E�'�Xc-�0\��!��AO����>t+@��Vd�&0BO��j@`������0I#/�� �{)UJ��-��eX�HO���RW 0�(� m]�d������]e[C1�����h	~�x��
=�NYz|Z�0d��Z:�՞��Y�C�XKV�*t��&R<���cB8&�����N��M�}�0���O�BBbp�sR��^��!,4����4����?�|)��T��ͮ�9�f��>�	.�r����hBy$�+R5"N-�%�TO/��+�Lƣ,n�NY��!P��]� o>@ݸ��|c-uo f�<�aY�������!k�}���&���+�"��&�V�c!���9@(�|u)��&�֯�c��к��P��1�a���?eg�[�w���	=0z��5+� ��':�g,�SÉB�����M_/"H�����b/�ޞ��ë���^1���%�_*�>��qZ��RE]�H�:�k.�`�`�O$��<MM��C	�U�4(8�����fQ�̓d��	��moJG酻�[w8�w0�l%JJ7��A�>��g�T����@��P%[�eY�
�V+�A��35Y���'-��l���!�Cd���O����~7k�Bťe�Z��<�i+�CocK���h��H��ry�������fe�D�	�+�xA~1�����
�U,<��l`[�h�6����c����#��~f����>_���q�(ɓ �t�K���x!�i�}`�ևm���q�{F�:�	@�
��[]q�W	~��==k=�@K�0�ؽh%2~y�	���m(:�.BYU�S��鵁a�Y+�0IW�, #d��wĊ	)����� P-��X0�T`=kh5q��}�C�Z��I�5W~�
�e�<�^E�/�-J$u#��K��3X�Ὴ�WEP��p���v�g;���Zk����F͕]:0u�+�V�@�f�`yp1�_Y��H�l�A�N�rqA�.ci�m�)�_|8����)L�g�t0%��2���(8z`��Y~�$���9	�0���W��+^��~�-xv�/};��8���	�v[��3	�_�V���<��eNSC.$DVq�r�*D��H-��Wk�n+d����\��.��쒵���>�C�Ĺ\5_9��;�J���/���o-��)[�X8E{K2�� �3�/���-5����s;�,R��0�@�P��(Jܼ�����uy�04��(
��g����\���E�P1F� ;���*��/�*�O�$��~[�B0��(�Xطv~Y�z�z�U�D��<]�%3�J�@=c�Y�jE����tB}@9�� ���|#�R�;F�B��� +��7^J��c+5�%��r�4�I)-ȑy��>��%����A�/���Q��4M�;BH,�/½vR�'w�'�^�P�PS�[�l��b(�5[�x�=�.B=�e��B�U��G�.�і��2� +�ep�*+�a��f�$~�!?�?�,�(��CQ������.*0�X���/K�EՎ�Z��I�տ ��Gd������@~�2,	n=<&�)�3�(aM�\� Z��Yh���(OڼVZ�@����6�����2������ɴ���) ۺV5#�:��K	�1�m�aHp���F��I� ��qh3�[�mX@��� �ݾ����1�鶫�-[]�d��4��h�tG��!��U���xe#�
�ـ1C  Rh>@|H� G����UZ�#L�����:Vs�?��
�K�.����*�o�&�wmN);�3���[�0%Y|F���ɷ�i�x��U�J��-��MB@I9;��U���ϰ���J��1A�,�1����f��h`.:���%�-x�$�3�(�4�<�Z��,��yK��q�h���屉)k�4�h=5 �ą��ˬ�&:kE�P�9%W�3t�����]�;�������[8�Z�U1Ш���	����]�^l�
�[Z�^���i삞��ha�^,�B��z
ҝ�~�p��	��������
y�N���]��i��(j\_\�x�^����RϬ�^�ԕ��!:E`�1����Zg�0XY�����5�J��:� ]- �B�%�C�_
�a�����1 �M{u,��i����φ�0g4-f��h1o�Yl�J�"�Ng�i��@4�0�":o__��h]�v�`1���G����L�W�m�`E��zp�޷�S��y��_�A
X�;rw��@([��MH�b���8s�%�VfΈQ��>��qkԦ	t}b�����pqOf������=S,�Yj�P1�]*�yI`�31����Ⱦ���ea�<�1v�����U��%�u	BՔ-���I��<**�c�!��,j�KYh�ѺϺ�_��[����>7g!�����%@����A	F�pxIs&"vU_V�@�	B	`Rjt �^h)�A[��t+�T�ɱM�U�W�Y� ��3kF����lp��D_��y5���eCv	��Ig��A$E+�$ �����!�1տ�ݠ-�M�B&hS({-b/�dZq�<�^�+P�E�W��~� F��#�7O��w��	�_���c��|�u8K�+L�U�ȭg,N	� &���)������U�p�܁g *g��P����A5*��UQq`�	LJ�Bv�yV���$W� �e��MY�LpW� X�yladu��%��p^���G�u�_,K�y�!�c��s{o �!XS��PHj�/�j/� @2:Wq��E����]4�Q�:��hg/�d+��-0�#���ZY`��x0�3z]�^Y���2*ˮ_�� ����?����~gi~�%�&�B-3_m�5sP��*���/gV�ࣿJ1�Ӛ}ʍ���A� ~���U��#U�/�x�#�T+Pwt!A�ݼ�N�ѹ�O�uhdek0�u$cP=�
�G1�)��-�4�\Rvb�{�5���	� /�d�%)�:�}5ʀ�����o PV��m<t˸ݤ�8�Q��9,�S���/�@����©�c]@<��}__"���N�2��2l�hY)���A� !	$X�)����28J_���	"�r�0�-�oݖ)Q�j����O������ݱxā�C�.PP'���`�,?���[# ��Q֞k�Vz�t���x�w�	p�:�����0m��>�o#T�j�6Z�����U�0''4,�!�Bzg.鸤C����6W`�e�[�x5�$bw��?��s V���kZ��_��?MPcR@[��$\��?+ᇿq���0&�R�9������>�Ol����W	�_�� �k'��;�n�|�&��̴�N�����5p���WA�����T^�{%am1n�� �3g�rJ���M�
>�4W�'��Un3�1������4u��/2��o��1�]��L/en�5\�eY�À�̷���9_����#���V�^��tA	��N¨^j`9*|n)<"������G�`��Z2��۹	�.@� �h�/�P_��\حj׶���Ԟ�"	�Q�B�3&�P8;#?g���[)���ؐ,���i�mx��L�����]���:p#�S��Q�r��Y����PĂ ���(ܽ��~�\�5]�=�ZN��U-]������V]�g<��	�c�]}�-�C(܅�����v1%]Qu�QYP��32�^b��kD�F- 5�?�g�2�s��V�Үh)p�Ű�D�$5��=�p�2�L0�M�h���fq���0��6\I0 �OT�M�QW�o ~:m�
)�-%��(ݽ�S�9 	>��@(Dr�������O�S��0:�(o_F���h'1kF�-,`��^Q�������y
e]w�f�`LQ& fiF�=�k|��'zfр']8p�ðS�ϓ�����B����pE�H1��,�ג��ʛ�kUl�4us6���t�	�y`h�W&XQ����R�h�/�/@���	𽱋 w@;��v��9�tB���]�O�O��+�\5 Ht$f�/PRw�NZ�~��[$��n�������`����(u�8�%���ē�[ /�a{�*�N>�"O�(�gZrF�f�V���o� _�w�1�58	�p�&��X��0�@\�
���'��wE��H�,K�n�� lv�x�TA4)�V�F'NJ�Y�*� |h=0�%[���a�`S�>�q�=�ډy�:�`����� ��%�3W��Wk��	��`��qX%NvK	O�^w�=��	h�I��U��V1�����\�Y-��/�/a7^w Ph�)�H(]E�e����R-�p�'����\֐�9`� 1ۥ��� �,�6��2D)��H�9?	m�6V����&K�-���S� ����,o|D1�7}b	$�����Ӻ}����� �	3��V��)d*�w0LS���N�Uuk+�
�fPd�[P�E h�^����tP�}��T�_��Z�������� ñ���	�7��ue��P�,T�����~�����������htf/ֲPo�F�p�@���*��X����� �p�}���hi/UZ�����HJ�4��R[���K�Վ�	&��^�+��*hK'���y󝀑�@�b-�#�5�/���.�H�2�4t��@���?0�X�7g3��`��N�����ǌt�<Z��z@@�6dY�:�����t�h�b�fq����h�0Ps�_��X�
Z��6Fm0��e�0L\�y�U�e�������0=X�2�yo�[��r �xX�� �WP�?ٻ�wz�"�\HTX�ST;h�W�[�+C@���3ǣU�I��-����X��5�J�B7ku���@� М�J�ꌸm<��±��` ����I��=�-r�,�S��K�+�������\	��F=&�/�t6P�M���xHx�-u�i�î�ܬopL��8,�J��A~ �y|� ��@|)֘�����&o���:3�`��ױsp�e�D��b��IAw��+�@��P�?�Y
\������[��/�N���4Q�x�io�_q��޾��2so_��4Ӱ{�Jf���_�8e3���h�\�C���9��?�)p@h'�=���U�l���͖9k
���h�p(�v��wq���6�yߢ�Ѫ�( }M7f-�`L
��h�TW�	�{^� 1�_��U����ɽ�a�%�Pp�?���@Y:%]Ջ�e��K)?���8U��o�]}�a��A��+����N�ph�	�1���M��EY��DJ��F0�@a~�"$��`��:u�n)�I��hB��H�e����1@HؑPn-r��q� ��	f��)�鯪��8?�_ ��)�[U�}���r=H`�p�� hVm�1��>�}��z@y�>5wS�ڤ�MQ�4F��$8��mh�M��î�R�i	8&�V4�&�%T�����U� ��u���:����RX�0{C��ۇ�[JHd���<�����A����Ԁ=ZV�]Q�vH����8,�=�t��fS~�z(�AЗ8�WT`��nV�(U/�RBf�_Z\ ��I-�Y�[	��A*��� )�_���K���
9�@ 	�Z��x��#�4\fT]�)�s�Y�e��	� ��y�N�-����%d!� `v�C�}�c�J��^��	�	�yԢ Z��|�d��C܌��(����	P���R�}Tlt!��(��*�T�⽆P�t1��D0�o�*��Ÿ|�"���N -�0i_�m�r�
�Z��U,HOr�`�ze���}X�i'��]e@eW�d�����������Vٹ�������wQy��Y[��<�y)	�h�]�����[��Y�s�HO��	��Y��:[A�k�8��B�<��P)��'"[f��#@�G� 3	9^E���M.���J�ד��O�j����O��
�a]�p�x�a)��R3���	��_{������آ�	؋}x����,$~VL��Qc~�+�/���슃�M�1� ���5&#�O!G��
�V�u�g��8Fi�v9��o��_�&����_����#�w����}��Y�0n�hrZ�32/�����>w�htL1�
<zb�9����"�F�ȡ�@b-5+&�Q��b�_����Mo���a�RT]w9��mƓ��1|���8X�x^��!]B�48�)J�������#��cL^�#n����_����q��(�?3�!�)ł#P�XYIP�͝�h.�P���E�j�Y)����0<� :L�;
��Qk�D!�\zbh~�����L�{yv@sa�~�b܇O��e1��7?@/���'��x�v�X�Z@ں(U�Z����E�Ű�^���,xM�����ө��To�Ŗ����6�Pa�!��2XZU����鱒�@��	�:�]� sV�y,���4��}(�?�zITV�J��E@�d�>�s� P���nI���+��OxmC��"�����]�V���i)SW����4 �W�a�P5��/xg���` .{�i���<���]�d��;8��d	q���-���R)֌M�G���1�����D���[p(�u,� ʭ�䰜�.V��Y�N���@����H���A1����b�����d!,�>QTE�_�)<�bZŅJ0+�	�|��_�	��}<(Y�t��u�詚 '.1��B�}ш�&���8"���X9?�q��<X�'��Z!��[zW;
�0eZ�w��<�")�-Eճ_�*G��J:�ܴ�-�{����ժ-��9��u(��)���'?4��NJ��P��#�}�Ũ%�G_b�	����.�2T*�+ ��my�2�B� 1�]Wz�?0:)��̿h�22]���_rc�1g}y�>g*�*/�3�F/��v�o�j> ���R1ΐ�)���P���0%Q���x� q�{�O-a8tEв���J�6pM(�#�Xv)�0���+��-��Z���|��u%�4�0��1O)̟[L�V"$����Fg�hTM�>1������K�,hlL�3�� /��9W7ހ�:�Nu����:�Z���07���)��L����:	���ZE���
H0��q�N U�"׹����qx5�B����'b�D������ѝf��ޝ��ϟ!Tk�I�9�����(�U1�*��=ZC�!V�lÄ��/��Q��o�t��rdA�|h�����a���Y������������}��ݫ� Qx� v?�
����ٺ���$|8E�R�V�� �)�h)�p��j�7>�_[�-�~m��|��]��o}[��x���.`�����ۇE����ב�OC�YȊ� �5 �AV�� ��1�^)ϐ�[;���_�����Vp�bY�a�)��0��)��ep �k]�,DbZo�+�%2|���9]@�S�	�L�d޸Iste��g���۪W�V�vо7���_V�"�Q��A:��h%�jy�����O*���7�6YǊ���X�J����.����Zꧧ��1b������n qKJfZ�P'���&�k|ǭt\rw[D�`�V��PI9uA�B ���5�&���S�	<��)!�+��J~fh(ҡ��<><J��S�䅈�;kes�\7�����q��}�+	�^�T� GH�'��z���̓���r)� {3$ �Ši3�m�V�? ��!I��xu_�6��2�泡� :�+��B��陜�Z� ���|&�n��5�k!ԇ>iU賂���l)$K�ց�G.�u/����-<, �5�Rx�8	�<e�K�vy����?�g�� �P-3��!����%�4������;�Ӧ�2�R����<�-���Ӆ(��$��П�!� �{WY>��?)m���l����!cǐ�2���
�4��./�@q���f�e��9�1�`�9,%)�h9�}/v���WӺ�ċ�x�.8=����7x%-����l�g��Y �9L?&%�bZU b��ه�� S�UP�QD]����J���$�
�LQK� �aPAI�`_��\`$�b������T_sl���L�owBj:ؕ���XhB�`��҉���#J�M{�������|�c�$�.p�C@�@��1�"�3�����ʗU�������X�i_qj�����!w�s��`�_��V+�Q�0t�,R�� U;v��%^k	څ2{���WZ:�g~/髈ň	�J�ls�)�@�5�>�a��j21�@�(&�O/��>h�`���Ԇ.�G���#���^&JOG��ׂCi`C�d/�2Z/�(FE(�r����x^71���.�0B��������?���ŷ`�׀�G)���T���0�����fOY��X q��t��k��J���/��g��U��Pq������<N���N|�S"�RW�:~Z-���r��5.�8���-
1X{'V?��P�`�>���U������QZ�:��P�w[�,}KOW�yW��@�[h)Eͭ��A�da9�̈��ٶ0�����[�^���~A���� Fz�sZ���^I�m�-I+:�N�и醈�'����}�Uz�i��C�W\��0�_T-�󽬏��Hpu^�A@�l~ O��mK8������L{� �?�b='N �[���Y�����b��L|�����˶քQP��ɣխTL�_N���eu��k�aא��Pp�`��dpz	�C��� ��9 f!L�N�>�� h�5�]�	�k�2T.�{'[>
3)�-X�5leH%��P��H�+-ik�^�_��+��������	A�� Ĺpj�
��I} :`��)�ʰ�`N0ǀ�N�^�����6�b�V��/	��)�1[{���	��R�ĭ:��<�C��؂":���m� ��Fk֞�T�������!R�ao������WO����<R3�#���	i�8?�}g���� _��X�ڵB�s�� JYXh�[��)����r[3U��s��׶WJX���s$�j6A��@w�Nx)�� ֹ��d�%�C�\H-q��0G�ZB�w��At�9 ֚�)��
#��9˹����|hЯ��n��x(Gϒ� M�_"�ON=������;�zbXI�K�*�^o�2{���gW �';�}�h)�ZB	�YIM�\9QD.�X&�S�}�'����h?JY�Xփ��)�����L	�p-�怹P-
�>�Ҧ�_1�U��2�zo�MJH����։ӑ�Qf;ah�PQϷ�0� O��2������� V�f�O -:75�=�|<�E��7H���C^�1�-�4g#uЂ[�vE�fT�k:��h���rO�n�������J�S��tF���p ��Hg�y)�[�L ��(YD�-�݃o|t��A,�ǔ��Y�_��\ �a����j���/�G��Ж���[���35�¼�8Z�+! ��k�x��q�!m.��UHf8�|�� Y�qDK��A%0����E�����j�4Ty @���
�!�i����x��ހS8ZS�/V�s7�?g�4�؎2���(��s�;X�e)�׉p;�0>�/��U���L�!	qv^y 1�p�<��`7����<�`���_� ��Z�/�E�AXRj��^�P�x5�ӛ��:ֳ�S}�{�wF�^�`��������ui�6n��<^;	��QL���8+f
�ř�0�CT�om�W!�htQ[/^%��$�B���b�/�7C-�����H��u�</�] 2f�	�����I���u��Iu1�����˄ժ���	Bjt}�U0�a/�`��pD-a�dZ<�[�T��RV&�1]�*KZ�4���J����2�a��`1]��2<�w����t4J*W�Z���U�,Of|3�Y���Z8�d����)�hGp�5e~��'��
gyL/���0�鑂�l=#����(����,���K��1P�&�*IXn�(�"��^�v'�vW�W�]�
	��/�b;�|k�d� 58W�X��X�d���=YʿL�4��t���W�DA ��H-)�����$��U��
�gi��V			>��H��S�~�PMXva��k�d���9{C)ʘ� �r�+�G&�[=������8͐^�y#@�)��sJAp�#�e;�������P4?�j7���(�-��
4!���!�6F	)�!��	�[���! �h,�S��Q5@�[���(����)�I90�:��B
j	j"��O�- W��y��b�1��}0�t`6}<+)��F�]�?�Twty�|^��*h��V���h���0�6�( S�ǆ��i�_xNsC;�?�0 �p��L]�@C-#��B�;���q�[���Wɰ��l%vf+�Q��x����AK �[G%�\rS���t�I�L@���%�y� �ˊ=-Kk
���(L�	-C��3)�(��s���N���:�1�"��m�����;XM�;�t�T1�5�qY����(�}2)B��wN��^[�ö_f��-�x-0�R���\`�}�iQzJaP�
��;�/�6Y@;&���/D�v<�T�"a�$�r��C2|V� �lb|*!o]�Л�@nlHVp7�v� �]�S	NH5`�dF.�kI�HL�H"���Z,6�n8��@陟�-]�����	"�zѳ�1�L�-ZkT����!~�g�P	_��V��	X����9��qt���0n������L��>uA��u������'7]�����m@��rjHWT��jT�U�p,t/�X� Y��d�6�Z�T�-na���_�A�b�~  ���ӻד��N��N�N�E4�ߴ*K-x�j�<��5�C����y �k'cA�4 ]Qh�IVw_�xw����`:�A��W>��~�T#�}GDR0�����l�(h�dB� ��:�Q@�AN�38��dt ��m;��e0[�>'��͡3?�����\�T���A-�Mvҁ/�~�eN;�N�Ϲ	Z
Gt�a鴱(P&��$ESFBR��h��� 2)��EF9oKQ�#1^D ��h�N {l�/�S�%��ʻ�:AirP��X5�(�!���jJ�+CX��[�}��f�!��D��5�l�NR��B�$]��Cf���|p��/���vW��9��Z��K����.�9�k���s�In�?_�L"+o`�rj0Z�=��w���&s3ah�/+Ϲ{h�8�/S��d^��ft?)�� ^��w�Y-�&{k���]<�5w6 `[�J�x- lb�8���|�Zj(]Oɝ��V�><m)? ��y��� �!$��-�;`|0���`�[LPy wrWt�-��L�w�n�}�^�#�;S��R���d���L��U�3���4Y�eAz��e�a�A4��V�}�W���2�[�fJ닋X�<Ip7�G��俈��thWn5l	���S�[��?����P��h!���D5g|��~	Yuz��h8��Z�9)�E%�@����XV<",)�/JZ]���	S�s�I���?|p����S^BA�x�l�7?@"a�E=.���&�	0	�[�~@�;)�^�W �N����(���G� �(��a�����j,L+����Y��G�鳨�g����?�Q�~��\(�:�vPL�����������%Xl&Z���	�,z���l���!�}A����m�Q��i�91J�&�K:�`�_��W��	�1��Z-E�H���.�O�a�R�� :')�V���4�T��c��u[�IP�����"�o;� ���N[؝�<��Z�Ǟɖ�)�"����hFf�j[�n9�"���J¼�H�*�9�����f&%|4��t������X�C����z$Z,O���^��fuvY`�G�R��D��w�~[��_��ka�>���^h`�h���!Hj�!d�p���l7+�B*(?�fV�<j�7����������Waeb�'([���!��o�z]p�VZ�ꐋ AK:r��g�K�Ah ���@^r��QxP��Z����L��{�������?��"W��!�)��]�O_�����Xi]:��%/��Pg\��(�F`�Ys3��$5-1}!�~��cg�t�K�����������Е�Nv��	4pG	hjl^	�R?��&f�t;L�lV,�=K���%[��	�������(h��^�^[����Y�O��ID:����S���w�^D�j�i0�%��KX�1>�ه.UW�`M�2� /���1����w�MҹuV��_?�$+��#�겵��e��
9����~r�0�q(���]Z�g 0��%	��R�K�96b��]�-�wP��OY�g��|�y�{W?�G}}w����T�`��.`aj8�E8��_XӀ��sVt�!�P�Y�:�r��%H2L��
���T$i� �^S�IskO'�#K�~i���	yaʻ�����鑸�PV�}���	;��� Ð]�HWh
D�J�	��a�R��hL�����Y���v�����&g�hO�qP��)�1�	�;�N�lB�Y���e����d��-��������*�)>+�<�0�0���g`����E	���^	��J'���$�!��N7�UŅB��]�`�TP�)��̟W�>./P�@zc�Zp��	�$�[�iԤ�9�2�fYU���	g0.E�P��-%�`�J�?��&����ky��f�Cϥb��8O^�RhYW�[��}\C�ݧ�����5�h��?1�ҏ*�Ô�/J�ʢv!V����"*(���%e����}����֠�3i|d4!��jG_Ts'��� �(�� 5���%��HgL��PZ)��� �� ��xo&��W.�5G'N�S�\Cp��y�� (r31^�=��{W	��
�����h��&*����	�}Y�����a�K\�˿!�n��6|��B�%���^��P�� H�'�1kD�p�eq.���=�t�}V�^Pah+B#^���K���Gܖ@RW�K\EG�sC��B�"P��A k�H-#��}�E��S�(H� Z�w��;���A��Ӵ�q�	�1A�:5�*�.�����3�j��9�8��&���oIZ&d��	p}�tV@4�I�2���]�L��v�=[0�¡s��6�j��1�O��b�Hh9y��܀������{�J- ܔv�o����̐�J�iB��0�2 X^�3CQX��.#���7$R*j|kAviB�+W��נ�^c[���BY�������ȝ���������n�����~	Q����l�D�|7`P@Np�G�����/�[8�QA�g7�1�9)�:�(��?<_�vYh9���[���8�_���렀�fP��N�F{��>0؃R�d(����?D�����;�3���?�����hc��R�FLyx������]��j�D �YsRc�Ot�!��-B,_���/��1��B�]Է��yda���a5�@h�xE�|��'w<�]D/\!e��H�`	�_����!��
%��
�t\�$����}1?����$��� -]<�|/X\��	g�U�%A\�B� ��{Pd��b!�#��َa1*Z&\ ��W�r�@8������.*�K�7�.����ٓWO4��b.F��~v���i�B����t�)��EF��[����:qH;�mK J���@ؾ|E�Z��n�?��C�qH�AXz|�B������{�Y��eS0B�Q�h��fv�X�'� Hl�L^oȚT|_k�1Հ �y͂	VyhN'VvX�7(<H���05jX�+%�q�S��~
@!��n�|;�B��']����<��	9YRxqP�- �TaK	'7Z��P7���a������io��A%5�h`��J�����̔�{�,��z~��s:_�-h}�Z����@��RLK��	�T��G��\h0�McY�KJN ��x	��,~��B�S]Rq�����������r �
�5HH�^�RAȶ���-51L�-�B�y�L�� ���ă80�Գ������<���u-��)A�+�/�x�;���`d���U ~���-�%�l�;
�h��/����}���t8�i.�8ʃ��0uE����*;�<�G@ŀ����X(�Z)��M��10�k*]X �|pM�u������>�\��',�m��C�������*^����lp��S�qA��l�K�0h��UB��� PZ-6qsa`1ԻA7�Hk�(l��@��VN5x��_�P2�흌-�[0���h���	M ����^%�j������ɨ� ߀��QhŊ{��)�g'�=�;���D����Uq�p�A�v�x2��u\����c`@Y���K�6R�y5��F���zp�}V�`g6��(42
����)�u���'v��Eb� �q�/e%0GZ�0�y Q�� +��<�O��\m�0�Tb%�"&���V?cV�W`#�a��\�+Q1پ�!��܆��d�d��� b����RL��%)�[��Y�B�ˮ|%Q�
��.���Hc (�f[����ke&^���)����J��(�J����3ZO�$�=i_ހ\�0g �������^eо��r�+[��#�	�1kH D2Z}U��J��+����!�1�^I_p�Mh�l�s�����9�oG�J5;�T+[h@͖G�8@��p�wX4��h���vF
O�=���:��#���z�/H13C�+/C�L; �,>�S���@�nC���"��'N)��&1����]���:�
��䢏�9��3>Ƭ�BCl��O ��H�m[���)�n4~1��r�(���O3qE.�TY>Ǟ=0GtVk��%�[�N'��A��_^���b����LO ?��1n_���ZWD0�m���_�I�	�@��K"�D+�Ņ�(�s4� ��Z|luJ_���K���:	��SF8���6�L"f����g�_� ��V�Z��1�Ix9d?Pp��f�kR�|�����Z���A�:���!`��0D�Ԁ�]�������i�h
��%�>:��GM�'���6���.1�VBk�tN�W��h ד@b�wJ'N����Y��a�&�.< `qw��r^���X��V��
j�.>���۱��7/�c�BAh�d�]\^^%�V�5���P��Ն�y�/��`��}���xz��(������sf�k%�ev�_>��#�(sn��~��e5�x1���}Bh��.O	��Հ�{����_�{�,���w�������	RTZԔ��B@�1[�D!�N4HP��}Q��8]��|t�2P��� Q��z�=�5�^<���x��5�j�I7*�	������R�A��<���UN����$v�cr���24н���K� ��q�h��A�;�b��m�>��������~+f $a��5�_�	uSU���HV`3�U�7T�x%�-���ӌX��ƌ�*�@�i�ߖ��Y�@�WtRiE�V�KX�:���N�ď��@^����2V�bXY�g5��!!�0�0h�f9�0�A�ޥ�I��c�&ܗ1c�q�_�GėL�"9t���!�?�|���J���db(\a������,��(6ꃧd�8�U��%Q�]� �h���S!�W/+��	��*���Rd2韊F�$5K���	���}raz)���:@+�E�R��/3	��=hA^F���j�JЭ#�e{��{ ]:+�h95�y;�Q�����Z%D�gd��j��& )��D��vGSo���^%����';�_�o�ZD�K�Ԋ���S�'��@�U1؉ū4��2In��;�,GNk�f��x�y��%2A~{��T�(��4�X��"S�
���1��k|k�����e�*�@�M=,	��K�v�X�nP#�h/�Ef��g��'2x9<��~:�bc\.��i!_�%�RwT�N�OӪ��k�x�x�1�c�m���p����*�nuY�é텪c���`[u~�r�I�N������4�` �+��q�oqF�\���:�5-�|H�.���[�¤(���*��@7{I](_��nAlM�%�9Xt���B������>�_�p������ 3`1����`��GA*~*cP�h<B�qe����'�L�o`*�4z���.�_�B"~$�UWh�2UdB�f �X��!l숰�/�I髝UH>'�Z)�1����V�P6!%9:a)V��+�u�M-Ynl(K��B�~���!�yT~�Bs�H��W&�u�-0%�u�q ��9����A�Zw�I�G^	Q&!ȀL�?FCH���R��`]�����_��F)"N5��`Jһ-D�W��{ ϖ<vds�'Fp� �+�^���0�Hsvbz.8��ۿ:=%wp<Lj>��|kE�ьo��H^���.��-@E�z����陕��P������x�?9�Y��(���PH� =?ڹ������\��}1�$N/�oGizZ �BK1o�����
V�_f�M��KC1�)w^�RF�}��v�����ў�ն��6Y�5`�N	�r�1S�	���c�������P+{@�\����??>�)�N�� �Ru�k�w���*����,C#e�Wmpn���?;)+�T][����@�>�{�D4Oiy2m��?��_%SA d��w��H5��e*���`}�)O4��r�@4Q�mL��?;�SqpD�;�(8�9`/\}%Z����/
��W��O�G�F<�tU(���MR��y�X]@�^��_�a3��$a�/]�;i��S5�^w:��������Y��	�K������o��&M�}HD�/�^<<hbx_:�,���$�@�P�B[���O"ol�T-/�E��D��^%Wb����8[��nA���:�- @.�i4�l�?PQ�� ��M=�f�ɴD�lWx���e������+�	j�4N�Ć��+R�S� C�
�n�k,��g�2�kV��M�*��I�@�2�\��CI�LL��bn�K��<c�l��Y�aI
pX����gY} ^%��^�� �Z�5ez�V�ۋ�K�%�n�'P x, �}7@-�
�� 1и��a���*��  ���~e�<���������|D_F\�	Wk�)}j�zY�5���`TZ ,�OU�i�+�]��p�K����5X#GD�ˀ�q9n�K�. �0!��J�� ��N�}�ڮb`�6�ʬ��Y,s��nN� ��R�'x}F��yk�}��IP��΀�{���4K�>㟂�u���d���M�Q��sTJ`ӂ7,W��;{V/�8]��J�X�LIK���h�1驨��.O%֗��q#h� %���j̜�	Dr_�T*Y�G��cE�;&�Z$n-@�|�K ��X�j��OA*�<�� l_��&GP���v�V��2�X�RYZS�L�:-/����a���qÕ)gv�'����d�C�_Z��J�	�!�tm� 2[fS���K��^hV�2;���UZן������9�هFX^�����(�!آ��7�Uꁊv�B����UP���%t2^�Z�h��ku.
�Z�S�8A��'3_��`��� ���?��l0��4�h!pN�w�|�ѯ�Dl7 ���N>��1� ?-j����_�9V/BTh��R%tP�:�����_��� �R��'�@�hd{�������tI�ހ�H�_U�t*���������PQˏ`�Yf��Ԙ�|���=�'/���H�A0�fK��v��x	�J�����1���X�Yo�V,���&��^`�h��;�E	�B���A/lZ1��;����n�\��/��ĸ���0�qY������#�����a��7�[��+7#�b}b�abe�����5&t���j'wJ-�  dVR�4� %b@�}	"�0p%-u韛�ʐP� >n�e	��Ԟ���D�C����Ğ<�ꇘ�ͺ#c
�0���
_� ';�=���+��@����ຳ�ґ}dX�z,/�[_��MUbm��w�4IĴjDk���Os@��C�	���Y�)FPP�=�pX�.ɨ�>}����nZiW�'���"�J���3����/��$юN�޽jq�&��<-��@}��V.8)��HC��Y����_)�t'�W��[�ah�&C�������S%��@�,���r �%)�W��r'&v��`�p�>��3M5 ���a���	#� �w=&^Sd������ծı�Ĳ������Y��6�vT��z�^\���Rh	[ p��5���ڴ��(��R�z2�^x ��7�O��į,}�-�%��x0���YM	Eh0F�	��7} ���c�����m.����ͯ�Q�</k�0�j�sg	_��Ŝ���蜔a�х�����H�vF�s�6����{�q�5$�3t|V[��[
��ә'}b��q)�X5	_:*P����z����(A�Nu���}�`U�)X��"_��<���;�)�D��n}O��0DT; �o%�~��V�ܶ|,N@�r_�eW����Y�;M�9��Q�^MIrA�	lG�?	r�4��V��7Һ��Tl��͚�^��t �!�@�M0��uO��O���a�O�U,� g趷>���%�����5n�V@��u�]���pJ��nW���4"Xק�o:/'}l:B���H��'��1o�|�1-l!7�0�x���տЄY;�82#��J��s�Z=!�/p@�W��#�51��=��s�%����w���>G{'s��hI>������u{ω^�UljB!_V(�݋�Tj��	k� ?amQh]q��s^嶦�X���Ձ,T��e���9�	,6�K��Q���:��7��m�|\	}q����}%L�-�PX�y	/58�۴���z��uZO�B�%�ae_@�'y`�nu���nJ�S;��>]�8L�9��ŶL�,8���t���y|a�h�~�E7��3^^�l��G**�]9�/N��8-�u���9^����`�`V1��� @�&}l � %�O������-	c�<��ق�2��hY�ـ�F����p��l� RS�~��	��=���� Pv���=&��1�^h�	g>mXv^��~�	�-ؗ�`&}"\HR�"���X)����_��x.$�(�E6�H�iW���*^�t�cRh�o�'ZZCj��9�/��p%������ڀEJ�$�0���	�
��� �΀�Z��v���� �[��"9*ӆ[d����P��|d�Kot]/�&|v�Q�p��9P����{��"�@���i
�zǓ���̂` a`�Whk*Z4����[U���"��>,r~�%ؠ/PtvP�ʪ�2G��jXh&�u�`�/��d��P-�G�U�=��țʟᛏz�ns�%�դ����x��)�j��^D@QZ願���X�Lg�n� �����O�+[1�_���:�G듃���s2����
TY�@Xd�B��I��B��H4S?+3��=��b:ۨ�!T@�952<�d� RQ��f���g-���D Q��)=Lh՘�A�'³P����۷`�sZ)Sn���������1��il*��,�?z�aP�����bG�9�~��([�K����X=�ī�L���^zKb0��c��'��ߔ�!fw�Zȥ��Bw��:�\�&�ʷ�Tp������(bY� S��	�6������~�?�rx��aj���\��g)�铱���?lC��)�}��t_aa:�k-j�<����4�Gk����h�_uَ��ZNZ�������3�T +�	�0F����-!�0�uѸ�������i�<��)�I�4�n>�]KS�Ww @"�#�d��/�BSS"���8N���ֲ\]�Q�V��e4Hs��5�G���Jlv��Aw�J��D�:^����<��R{�%7$t�!ү�݇�v$ú?��a?�p��3Ռ�q�ƼLN���R��h.?f2��x���ɂB�1]b`x����N�l.��h%�٠���׸B�� kS|(6�p�靵`���;�ϠL�$_]*�O���h~�o|^T��@�&b���MhzŘA�z��Ԓ�|)���&+�	Oh�]dywT��A�����%����F��;`2Hp����8ׁH�	�>"��!L_*VH�� ^o��ʂ�[�w�߃��K�	�`!ׁg"�S�{���C��?)�X�"�_��/~+|�Rh�rU
Z���\�r� �]L�(VT�h@X�׾�Z[�z�(	�;V��I�����{b/ ���T.���*I� :�����S�d)Sc��`�}\���	>Z����	� ���v�TZ\���������'0��@%b]"h��c�<���������Z����}��,���XbXB�Vz�.�=!X,�4����][�2O�����(J��B��y>b�^�n��4G�����CC�	���W��k��z-Xz�����
_��,0����?���^�q��{q�K'���9���b=��\��	JK�:u�P�ա�%d�!e^���hAp���J��� Zh�_�D[NC���.�����q�c+�U&%���e�߱U:�/J�N��2���tJ _��5�)�"<0�L�����*�	�y�`�#3��&,�F�5'�\sG*�P�Ӵ'��F>4��.����R�r�=�Zc�e%tFN�>:��O�\h`��-�������"x�H��t0�O�q'8(�$�	[Qw�4�rrA>� ?�R��j�l/I9x�A�*"���b�4/� ß2(����Y1Ah�I�ut�Q�m�	>���۟�!��aW-��@S��[.�c��������ɽ���Eр��"�)�I� ��A�����!�U6�{�tD�@#�O{2�P$h� �!k>�Ҋ�M�V�^�vz��_�qc���ɖ�͎�2ځ�G$ނw�BT��5	�6�giswΊ
�%Q΄|cw>_ �2YfRS ��I0����x��_����`�f>K�a��8��P �[���0�x ����-�����=�Y.jOlEis�%��r�~��'�Qu%�R�b��A4�u����'R}�V�WIQ�OEEN��e�=�eV3C�6�������M'�j�R	���<vw�LP�"�� S��W[�ÿ �X��>����e`(��� !ѽ�yBQ��|HN�<\�ޠ�� �7�^�Á��T�O�F�;�	�MUgTṇ"cx����1�!�?�2|0v�"H-��9G��(�CZ���r��_"01B�:w�(0���Qti��Xw�M%u����;rw�>�S�v0�f�cqH�| �5�YG�Ƹ�2��	}���Gc�,��p'���/~�U��'c� 5Dk q-�08�(��X���C�Pb	�ynuq�����v� �x:4)�Wh�>�7�÷�l|���I�-n�	�h�B+��=����	B�N�@���@`�^�)�[��kǝ2��]��CŘ��v�8fh��ڳ�����(oK �(d�0=���_h%tS��a�3�v�P�Yl�X�� K��w	\��{]vuP~c)
[!��Z�f��ɮ�0��J/�Oz� �����T������I5`ד8rJ�N'su�]�`N;��m������)ޒ�]�{�ax��h(�&</N�*)DFЃ�P�n�Ѐ<� �l�3���vDm�r�?�w����L��Z��A�<	�}�@�5�����^���qlz���fu�|��ќ-���J��U ��Q{h�8�-�	h������	�8�]�^y�%���`� K�\��۷�ˠ��@!g �.F��?�1` 
�~�>	�9B�4P�еX���:�d����i��-|6Ĩ��%�פֿ��c�
՘�hLN��^�$��q�û�����ִ>��Qp��d_�
t�Q�6�N�/Ū�]r���&���Iz{'�}@�y��i_��^"����	d�=ϓ����˄���/�88�B������̺�X� s��	+wٵ�����%y.�+)v�C�S�`Ȁ�H��`0�[�9��tC�Q�u�1���z"r@�Y��B��*��s�V�s���^����{n�}ǈ�(�K��2%�������+xHf�^��V[��s�4�������>���HTD_��gi7���:a3�9��U ͬh�~%,�aa��c�:_���*SL�E�1�!�p`Z�BT�k�`�y.^
�iuQ�Z$���}����RQ�{	��P�NQ��5�]�lh^/�8��)����o�'�thN#��m�@*�S�_yz�h&%�wU��J����[���������ŀ)�}ĢNӣ�{��o?Eĵ�a�� P��;�d�
�0� �
`�h�[�(]ґr��=&�bfX5-��<)�PS/hdW�c���ģ��'�%�]i|r�|�+-��	�LpEU,E�wT8D�<��_�j��NJ�̕��8��sk(�u���<�1�3~9	�A��Z��c��}`�>b�X)�@1(X9�{���h�T+I��B[dߍ��Ѐ��}�r�A���-"�������)��A$�b��l�[HT�?e�>��\6��<���U�x>�%)�]�����2��m�2����/�,1�'��	$E�*\ d�)_����1�R7�Uѫ,�{Y��$��	�o����RA��n	X� p(-�	��z�e9�P���8��/ua�5��Y�p_��� ��7g��g͂fQ]��;?Y�8�(���R�}��{�� �Z��J���\�F����Q������`�pX(�Z 0�P���[��0-�,
k�M{��K��:�Eo��V���������C�Gd�1��(���N�ȇ�3��	�	�H�U��%[{�!Ђ���G�\	��|zv< �G,İkOt3I���xI�>��G�~�zGh`�<�����{��Y10��A�u�J���;>N;�A�[h9:P>�]	�<JB�lIVU	��?�UZ�p!�%\�&�)Հ�1��7�R�h?��^<k1���$�]{��*��	����^w�WZ-s6q"]�o���[:�$�A��!�>�0L�Bep���5j��0b
��H�ɂx1-��@^��˝RC!��1�B�Ktpm��������fAw���� ���¡�	5	[���:���5����rU��u wk-MS[y&8�T��5�(���pO?��-$sGl,v�FI_s� �L�����Zy@�.X\R�ͤ{aY�2,��gO����^W�4K����O.���]�x��p6uJ@��9fNE�@���%����k.}�g�S(�-�=�8M�t��t	�����A��] +�$��	�hr�q,�4+ ��FY
�)�_��v���0����:�S��-z<
cN�D�R�ȻCEh�EFs�gkp1�&`�`OZ��4�Ն�
�İ�[��c�.�w�V��T�,} ��x[>ʍXL	�^�Vu���N�Fvi]U+����&[.���?6�hv�`��(�Y4K����q W�F� ��4T;��`��\� �v*��H-Y�*� eQ�����$�0t�(�!��&�C`����=@?S%h y���A�t\	�ɀ8YXi�=<VV��,~� ]it��O)�)3�y2(���������&�����2�0ÿ�"� �Vh)��-#~��rl��_3 b��x�Iʂ��'_���5;j��N,c�,�D�%���hxKV�O�;�G��b<3C�'?�O��������9��'רKY�-�6&�|�h�!�k�$�]	���RA0�Y����,R�����2�{��d�B�p)	�&-T�4�F�5�`�Hj��g5D�����c�)��m�0�2rZ,h1]���+�^e\�na�2�EK�P|^�_��B�;�IY�P~�	v�~1�s�9[��QȒS�f�J�Ī���{6 �n�rÂ�3K3��r�bB0����)�	��`�=��<�o�>B�����b�h�@�	Z��Q?�/%[����$�	�X��:6�6� ��>Q���	�&'^%���8�8���]p�R�_ �v.�ھ��%^߂y��R_'����)a���	\h#S�`G4���ݶ4HQSn�o�X@�}�<�y��q�oNvҫ�w�����|V�S7�ڤ, K����8�}D1u�%�=������o�i|�����C�H�"���[��(�AiPlW���$���0���+O���wB�?()��}��H-�w�B��p��
_�-��Ns<����H-����e�����AЀo��LHv���R�D'����(G!��n�+�a���,!���PR�9DA��p��2�w\�H,H��j@� �3R��/WM�N8Zܵ@[=P��]�;��a*�xxF���c�{̖��O������Q�ëgVe(�wY�]U$�6<ǫ��k�\U^ܶG[�0ݥ��?�	h����2�tgN�w�U���2X�:��,�:� ��&E0�L"�,��:�R��n�1��(�k�H,G��0��PE,.=$OϩB~HUc�c���p�q�nUlʤ�Y@�h�A��]��WP)RI� ���l�7�|�	vkp�D�Rst��Z��P��f�!	ϣo�W�:O �h,�/dg��4n�8e����rNנ�@�!���ざ�TH� �P������i�iWN��{�p�~Gca|��ȆSi1&��1�c��-�|����;�4��;h�Y�Q�ً���l�?����.�N�밗��H ��2;�Չ� �w�`��:*$U ps�
)�����x8=h�ʼ���`��5˓^w��wr����p	ͧ�MW0'�4��Q����2�	����h.+=3�q��Oә���*���e*�m���|f|=rԜ�C��;�U�3��-u�K�Ǻ���<rL��W�����F5o�
3�</�f\�TAQ3z��U%��~e���r��)! RK\��N�/�t���T���-G���`t;.J�����$� @1؁�q3�bol��r��Su	�nl{�5�:��Ԁ��0�t�q�Ҩ������m��`;�T����Wa��M�n-�U�?�3�r�^����H��-xfhiY'�9��|���~����;�����|�����s���Ч~!����Ȏ��>�m���LV2e)���ΧB�~�_{��®�Ael*�D3����O@0��O1НnM�^)\���
[X��86 ?�R�|�7��t�'�x�-<�R:��`Kt%���C/�p�(����`�
J�D�,.��/���l�U�Z�D���*�s,��T:�g�	4BXc�JhJ3fZ!��  l{��Z��w��._�|n�@$�rI�S��]i�OA/�8d�S��m��!`}����}J����~k;&\�n�^Y��D�e�
0M�{�'o)dG@�DЏ#}O�c�R��[`
R��[����J��`�^?�vDү�︨-@��=�
lj��� ��5WG��%D����?�z~~�(�
b��L>0���I����h�H_���=R���X���ʯW�&h�*��.BIx�-	���#�/�1J5-���e�	�Z�xR~��
��Z)N��j��9�t�l}�4�ˠ��熯�6�}��逕���qxSZh�C�����>�[V ěY��K�[�1�S��usM2)���F-|	ڒ�[t{���"�N)�1�h�rD�Y� P��d�{"�j��0��4U�E��xm$]�"��Ӧ����<������ل?b����IW���֙	h
�a��bt\/tSR��X�Y��.�, �-�݀�e8 �D��t�9�c��a��Zk�]i/��e�� :0б������;��Μƀ�v0��s���l�(ȲFT�3PJ��`���*<{���f�)��� ����LnHsx[��*.���f����|t+���$�a/�@���Q%rR�:_Ƚs-��,�!<���v��� �{b����[`'��0�z-��������0u���Ɇ�R֗������>�}"B�>ӫ�OZ�U��2�Ru�z$�� ���<�3R�����ϖy�&����>��'@�@��_�Q�!b9Lu)�b� Կ,1K#�����*�3y�/��0��ah�
�]�f\��uY�Kь<-�b,�KYUn��x��4�蒁�
5`d3 -EdW��'YKQ�t��Z밿Kꃉ� ��H�&^n�2�?,('p��]�5�Hԁ�C�u��ʝ���F�w�`MX}��{�+/��^=>�Vۀ��w,@)L��'� ����\0���9�������8L4�
�9�X�F�Pf����vz�'�0L}�p�$���� 8�z�������ˀ�~>i��!ʋ�"��^����l�*�Z�4�}	{kCPL��i|��yN�K��B�6��m�'|��Qh+/cp)_����Kn�x�IWE�7 `��?Qw�,�2��&o�th%"gO�������ͼ��nإ�_�O)� ��r���j��>e�VJ���7�;�X�d]=*X����k��+E�%U �m�[�"�f��PN6 �мU1J˸�$�ms&Q�����"0����;20�&�{�}F�aJ��D9J)���C��(AA5B�[��}z� D�����`��R�>�CP���b]�O_[b	�,Fr�ɺ ����_��bL �O���gcJ��.�'w~|�`1��K[XU���F���;̘d�N#qK�}@c��
��)�#W?3�}U�d'�PۮiH�6��P��K�CRڇ��ãD��������x�һ�=�s���a.i|'�͝{2I��R��%�W�Z+�����B���'�D	5}�OG������=�h!�f%���eO����< \(Ͳ������݀[����	��R A�f)ӟ^��˗n�SU��D.���Ǳ�'فoG/F*�{@}\w���+�a�ÄJ���X�V��;�$�������<���� ��7��8�h�n�]��y�'�sZ��o��\�1�9�<<]�-}�J���zZXW��1�1��Cڄ������u�VR$is�|}�Â��L�|'�>1nol<G	�P_��ۘ �B)ڐ�N��m�J6�W��ǛN	]���U�6��b]�	�	Qwx��'��RYA��z�^������J�W^������O��R/V�Y�4�q��-\��a��Q BU�c]�g�:9�:��d�OV������?x#���-�-Js��-V[D�¬�r)]�/[�|[����I�?	]�^���@�sb$�W;�n�ÝC]��^��
+����1�Yh-Ѣ�0P�bߑ�c*l���!< U�Vo&q����a2z
�� �+5��� �0XZ���$K0E~RPhs{)_s&-������#���\���:�&�v>�<��9N5;�9�1���~j^:��c�J�Ss�UXB�&��{�����1����?���W�v�w��o)�����k,a@�@+z�g��qq^H��i{�Lj�`x5�@� �0�|��Ht�.{� ŹFS�����I�A��j�&��@z(q�)'U9\��o���0���r��h'J���Z��.Y�'S J�=xC<���j1O ��;���"]U�?�^��i1/��T�X�����(�{9"�tP�1�5�X�	�!@H ��}Z&�rZ1��� �p��Hx��_�d�������� ��\o'Z�H���X�r����X�[�a�
��U��Ps/��|��Zk�໌'G��׈,�!�J[��HZ *be EM�~�LCX�I�{9�F��;��1��U�G��L1�!A�~SA����AD��j]|%k�APR��S����[yZ��n��4�%�q��}=Ħ��f��>���X ��Y����/s��XU��˴�!_�wh�߶߾�}�_)�{�wX�/�Fj9E��dZ����{�*�) pV�>����:8�W���K?�(�.a�h$Y�O��1�y�3TEL�[�n�s�M�����K�	�[�4:�һ� x��l's5r1�wZT�����hy3̑�]of-:�ԕ�����������XF0�oq�aQI7�
鳎ȗ0�)�-D���"�	H�I�Jx}�?�9:�,�U?�� x�ֵ�})Q�_��`� Tg*�o�/tiN$�}��h��w�p��~��[\��S�w,rvi�8P�a�.P����X��T�)n��	X�/`\w��j0�\9K�S��=���jA�|�E��9�@�5�C'����+.-?lgF$����S(AYn����.�q�yw*N�*�Jp4����eRlu��_|v�Q����X[y'��^'t�b!�]�9�V�����5,&�&��\��Aq�tP�%?	U�d��g1_k�����Ւ���4'��cY�<���?�^}�O��f#�b Q��t+��wB����:��{����D�1,Q��Fl��#�[h��*�&�'��R��50]��}f�Kq`��$73�����b�L����.Ah{bP8��U�O�5Rj I%(}Q-1����e01&/�+�J�3ԫg[��=sI��BB����MK��^���`7\�y�}bJ���8�k�<P��>� ��AN�Ƹ&��p�U	X�qb[��Y�l!m(�p_�f�(瘿�2S�ٻA�5�hj��%YO��_���_= O��W�3<ړz'��H-�"u��	�Y�'K�E���(X�HCߘѺVT�v�����ƾi��L!�1�td8�|�{�7�����#^��s�@��:cR1�h\��O�Z�5`k��P���|��w ���Js����i�
� h�W��,IF�}��w��ؾ2�����U��X��-���8�^��6O�x�b^�6%�׸�\V�-t>�0�
5�.N� ���_�����(��PJ6w�V��mvU�T�F4{)�w����#��V�8�K%qi����	^�P{ X�f�8��Y.toC�Vw��1� c�-���r+���*��^�v�9�Cx���������� ������i�"J+.aF�ͯ��tl}�匒O�B�D�"1�f���a��v��+?\t$c% ��X���b�t)��*'\��QgA�N� ����W �G�U1�JV�]m�o4h'�/[L2N�Z�,Kɒ����� ��P�IjT�`qo�2P�<�-�
�W�
q���%䑗� �O��i���ҳ���o��y�_�Bg��م��Po�R	�T�q$5y�c+�;~�@��O�~�r����1T��z�@Oҧ�p��9���4w��'�o�w	����PG4���0�7���i2JsWJN>�ͽ���D�X�:6�T�q��_��\Y�3�5d�z�&?=�-���f������4�ia��E񓿩ZB�m�"K�&%�=BUK���4�ߚ�F.�%X�Boi�.�J�
���]�RB��D���%Z^���C���(0t�L�+���ĠP��̀��T扞D<� TVZ�D%9��PN���~�@3����R�ܒ�TEN8�(��1��UaeK��lw(RΡ'��t+x�N#�E�$b�� y+s&��P��R�E���)oW �?�sR�l�bJ��eK����c�q�Sup$�%���-n{2��"Z׌��S� ���6�E+`|f�[^�$����?�\u���	��X/I!ȯ����l�:!4��n�yS/��X�N�K�M1��4ʠ@	�B!�uyM���zg�C�R�8/�9���1��	]6�KN�_"E	�9]����>�^�~�����S��o�8�ۏ�C}��$Ĳ����.3��Z��� ��B���t S���Z���:�S�o�V���)3jK�^�����	h�{d�N� Qe���	&b�v�AZkQ�I�EL���:9�A�w���	�pD�		0b �I;�:|�͗��Q	qcsPlZ��j�6�*�u{���Ĝ�^��0 k´'���(W��x_/�^�c�1������fh�-�P/� �݀�wD`��5�/'Wgҥ������[ң��T�b���E���Ipn^��e�H5�J%�)&�-`	�c�S��V�`r��dO^��hse��G._a�1�
'�Ԉ0����^WN ��Y1��+'�"�.�;mҲX#ŅT�{�gi�K��� ���Hw/8���f��iV���W^��	�y�'UF�,	v)��F����5#:�׾H:�N�5��AԱtq;��(R� �!x���6/�# l��S�X�L)'5��ƭj.��{����_c(y�N���~ ڽ�l P�~y4��s	e�B>��H�796@!H�a1�Q�hwXX?���m���}������Agk �!�731�[�Ԓ �����5	�O��[:�x���d�'��q����R�,�������ċ��p���1�JY����`$y�K�%�����U�0#��>��z�/�U�1�5A>�#*����xd�_+�9E�>FEm)���C�8Z��ƣ���W41��?�g�iV0T-�9�|�f��(w�]`�Es+�|>Ptt���� �!e����BE\`��1'`lTΘ��W���#yzX�A� �� ��9Ih�F�_Xd��Hc0'`��'�Gv�dv�Χ�j�x}.`#��0���W'D@�u��D�Nn	�r0	bk��i	;jW?B�`>x/#+<Zع� SQ�9�'0N���.�[�u���~H�*V��S���r�0��w�&ւ�����3	�-��u�d����=���ek^�@-�RX�!�����^���4x�t #�C�B��>�����l�����W�BD=��41Ș
�I�P� y��uL0�!�Â�2UZ�)K4k�Pj�����(��m���� ��tZ���.�1 �~U%�{�&lќ��5㡗r���� �ox���w\${ ��U��%y=�g�?���:)��������P�p�Y�k�Y^�`p��b'3��><�Qb8(�AW��૘ŵ�:B��@'M@ ro&`�z������#�0����8��y*�"o��K���']}��e����b�[�sp�_��8)>��=�����'�a�hK 	?�EJ�v����[o5�nG���ӛ���an`+�g������'C�����C��V��7�[h�z��Y.pE��^hi_@_��p3�]0S�����Ls�NE�ZLBA���yc���p�S[���h�H�/�zUV�V��4�3��p@�X�+$��c_&���֌��jS1{�d�Y��8n
�%��"�M-�i}7�����})��[=�K[��à���R_�i���qm�ޠ��3B�_�K8�����ɘ	���~%EqV�V ��	�g~�b�O���P �B��Ni,n(t�j?>؝�kf�꺄q*g�9T�f�w�#_h���?��P����Tf�����tF�V%����M��ِ����a�u�F�KQe"�Z�M���0���'�0� JW�N�����$63r�/�^��������`������_2a�k^Wi@F�{ #I	�[��,-DZHp��C��y��,!
u��Әd�!'�%W$;)�NA/�t����N���9���,0ќ-^x%��%ޫ��!V�r!���ͥ	v��P��(ZM�� ץ��-���6)��������ByN����=]WV�]F��f�AUE�Z���&�JOP� U
��{���]��.�A�sI�H��朊W@�1pS��-o ��_g\��)I��(k��lG%� BۃxS����gM���Wrc���!$�0�. �7�_1������I9*�}�8���E��xV}0�Se��&��������!�f����0�y,\[x� ��F���ك��[�o�T���Sŗq�_�T���h_p��2����o�FZ�a����k�h�X
[g!o�j�c U���=�1�]�O�BI�.�J�h�٭-pyƃ���4�	K�/�}�����p#�����߃pP���|�R#,�H+F~hTz��mt3�`� 1C�FJ�HI�+�~���F�t�KI���󘩰��|�fk7
�-U�������:�j��ƿ�y�%6}F���%����0%,) ��Wh�P�(��{T���6<��pYR���=�U�����|0�t��O[�����q\�kPq�>�H��-�A�	K�w|����H�S6X���S����;�G�@A���>I��T%1\���*�S��^(���z��]
3���V?ir[��^˺8���.���x)Uu��:�x�^ȯ3M��"��!��s�u�C�XX4�]��ZV�I��߆P4�9��<��a�������(�[�S����R�g��)�Z(�R�>�z7}���k��v>N�����A�U�<�T�T,	iakȏ͛�z-�@�?-~m�M���� Q��^Ih��Y�>�:�$K>�<���vJ��W'3����{aw���l^G	%����c�;�uJ��z���`�l)�y�:��	�ߘ\�huVF��K�e$J �^@S"4]X9�gc=���/K��ߨ�[�B�ӑ���/�d~���xQy�+�'�Rٻ����	Z+�d @�l����[ (�R������
�ʧ3�$���k�Z���>��)Y����
\/�(��kɂh�$2�Se�.������@tOQ��p�mRx�Д��=�u3
'Z}�	��s����	P�h��Y^x@MwW���D��B-�Alg������ ��r�;%�l w_ ]�?4�OE�d�=Mc(��� 7�V�I�[B_��X�B\�hD>�BJX�-��=0)h'aeI���l�^���!���p�e��n���Rh�3~ +Z�������D*,�0)z�_����>�E��/�����]���QdL�x�2��6R�51-%AW !V�E-Q����M֐;�.�?b�D��|�(A	io[�׀��O1�K7�4i`_P�?0�ZH�/)_s�FP)
R���~���_v��Yzo�B���U:)�`*�(W���-�<L���uX��Z��7'�F�EUUI����/�T%?c$����.K�u���|0!�Th p-X3����RB<�LV
��Ww�������A5q�A.#�P�9 �p��W�`E@k��}��2_ŗ��S��Zd��
 �eE2�b*�|961���U#o���~_	|?[�sh9Q#���f�0�ƚ[HFH	�r��D��R���ib<b|������XNU1�,nP'�A�H>%^ywB�	}�%�E�,-���tyXҟr�UFBP��.��������I��auh�m|���;-�A	j)�ES�	L���l��Q���뀼-��P|�O5�&~*�)�/a�{�Ζ�u���Z�n�(yf��q&�m��@HO�5��>>����	C�Ύqj���~hW�B�����[���V:�\k$�^I]J��H'�o/.0ƺ�G�EѰb��c���^`��=U$ZK*�z6(@~�q'Y>��(��ݿ�~�u��/����!8��H��X��>���O�A�[��3�|j��fF��OӅ�E����+�<���Ҹs��r�^AB@H��[\�Ly1`U��� �Q�l�X�fgqt�(E��Gb�|`��"�e��5�7a��w��L1�_}B��Ѯw#��D����S�X�� Œ�.Ӹ�����x�1��		�Z߲����V1�o40���gO���A�T��V���	�[+ )�xh�"��	\^ ��
��%~�B�k_묰4���Q�+����_6���aA�>������=Q߅�����$����67�`�)ڹ\ �b�|����`K�!QT0��	̍�~GL�Ҕh�xP�" ��(��wh����^4�!��rHK.Z��ˇ�Dl��[7%AQ��c�'X�P�"as���hǺ�־�
YF�
	�fʉ����	h^XF�f|�%/�L��o[*�Y&��-��@��.0�B�Y	"30)�(�A�=p.p�u3�x�h	y*����0��
�Q������:�1�X[f!$'�MX�%��:�/�*�I@��2�X%�ol�_f]����A�Z+�i�E�6/��_���Q��F�{�4��`��Hz,^����t�Pf��ha��vD���סS��LF0w�K�����l}/����w`���x��|h���G�C@l�r �1��p:-�v4���
�e��vdLV��}�����FEe4�^�l�F�����G�������G���Ů_~r��+�%�b�	 80e�d겗������;	{�y�G\�OI �������- ���% N������L�2�p��l��>�q�	��I1ŭ��	�G�E\ �Z*�~�J�� 8��Oِ�:k
|�	/�W0���)�C	�r����/��p�-�7�k	�V8���
<�5�q�0{Fޯ����pT�y���p~L7���:�HE�#�4i�1�B=�bVk�� �g1�X ���	��w�]�\\�\o��I(�w �H6m�o�T,k�j�ny�*P,�;�HZH�^�Uנ���Q�	�� �!�E�a� ?��u�>�.f!��(/@F�N颋�O���ה�>%����P�IB͍>�u�uI�`mS�7b=i�w��]M�Vh�͈?��,	��^U�����%64b���"~ �X��?)��_	�nNt����h
`�^$|Q4���ʍ3+�^b� d��t�V�;q̵)Ϩ�B$_�&��X�5:�C��E��P�xY��/�-��,G6��;�����Kt]5?[>)H��I��$��O�@&�k�`;�-v�Pͫ)	�h�?w��vd�+PaJ�}(	���.�P1tX�	�(���;��m��i�`�4�U�]Ň��!^M��)^�f:@�h/�pY>�'#u��r-Y���@�%[�h�	25K��(��K�����O���	�@�Ẑ��4���s��B�%*!�$�B�/U�?��д����0����5�D�2q�k`x�&	 �W��t��H�������G�]�`�?v�� �ы[������b��Ƃ,% ���Wh�V��y^%�U���z�����v�`��,
rAm,>�hKN �Q�����xy�0އ��,c�q�����H�{���L!^��Չ�1��Bv����N�m�r��!�葭W 1q�-KJU[��T��N�F�f{�0˗ѐ�0�X�,�@���^���J �6/�-D:8m�d#��q�s%5�-bU�Y����:4����c�Y��-�1�j�W�pAWg�'s�.������˂l�=�<���sRI������� P319�I��1�+�;�ً1�e[�ؕ�lK��ٛi�Q�¼y��결�)h0Wv!�������ke�r�,��e�1��v�����)�sN?	��d|:��l;�c�g�v �oX��8Q	������	d1�^�����3r��y��l���� )&�Xeo��J�)J�;5��1�?	�\w��sH����������ʼ_�υ���v�a�By���h�B�+���{�Q��x�Ar�? ��;U�Q��R$�b{V�t4}�[H��7�¤ �bQ��wd�6Wh9�j�b��3[��1��H)�A�Um��X�G �H6��K��������y�0h�"tDB���QKƋ�]�o�]��Fs�������Xr�_�'~����{�D�z�90���x�o�f�E�>�ޅ�R�����-
�±�-u�A��u�TzX]V�f����a\l���|0�E�c%=Q�a��P�-?#�WL>R@^��ǥ�P_�\Z�L:U�-�¿ԐT���f�e:�G�R��k�K���lŕ��A�o���&P�y�|�B%�Vs��f�u(<%NEJ��~䂘'	��l �TLAX�O|�O������)���T=v[����
�J6�#���U{@�`D		K�Č�k��yW2)�x�Wйt�b��u�?A�X�#�H�f�1�Qh|����Ҿ@���K�~��j1���ow�|�>aY�q��O����k\�(,�.y�`��@ �L1�^D4?,��%	���%j�5��A%�|*; ��rM�&��!�B�`-�5����U�A�q5� �@����`^erf*�3�LP1Fw��I��2�S����~�|9H���/��~=��n����4��}��R�*��c3t(�	�-G^ ��;�{��Sx��X�RWH�H!/EHD9�ut�8Jϰh�P��[�����
��XVkJ x���0g�Έ���U�Ed� �X-(H�H��,���b$�? uO�`�[^�7�tK��p��Q��*����Ek'�c'V�����;КY�u ��Xw�� �9]Y-�e/��|���
��[W���Fr����*u �����Dۦ�J���� S�BT�BkV!��������������s PAI��iW������Ƚ/�-|�$:��y�����HrZ7��iaن�-�p�a:� _R�n%�ͺ�1I!��R�R

Տ(O}�[��Q��ϱ(5��1L� �T�_�o��[�xs �8��,=�A��{ȣ�H�Q޸|Lf9s^R�Jx{3�6K�h��+߀�?Z� ΂@����z_UT����]�V��T����%��,P���)��S+.�]����K�B58̀n����2J�Gv63,�Hȩ�g,qN���^��%�X��Y0�
���	��I��@5�n/	%���;oN��s+J�0_���<Y$�o\Ex�>��D2�f ��_�U½y����j\b�x`�!�@��¨�{�& }P��fh�YXB��B�ǐ�-� �ϼ!��OO�]���u��g�a+̃8	f�U��d����<m����X��M��ɬ�;{$,.s�'Y!������%^�I�Q>�+����0��/�L�7| ��z�^�0�O���3,!#`6{]XR�]�w:�aXJ�6	�x?!�j��A�  �i�ڶ� ��q�r��eY}�Gh�ês����'C��Y	����i-7<vW
�h�����O/;?� P�Y�G ��w�)0��
�?{r��R�AD1n��E Hv*��P�������th��=�!�qTn��1��j��@6lB��$p�/q��B��+���uy'H@{^�L�b`m;�jfqO?̴Eꐆpux���U�1�Q��W����ԋ�R��4słh�nY.�#!u�h!>^�{���	H�'�@B��L���.��we��o�W�cp\h/qy���)uq� �`ZJU�C-�b�v����
��g����t'\|��*T�R
Vj �k�M��8&j�OG��������$�w�	1� �;���@�	��=���#�h�)qĉ<Ѧ�U�'�EYI�a&�_�u���� �f[h"6�Wрc�Y�_j��.����1!P�%#sV���!л�	:d�k�OH��/��/Z`�R�:��uVq�$t���N��Z��`԰b,��JD���VD�3�iZ���ԣ[ ���^u4��I�RK�N監XM&&�S�~���_v(�Tv%�E6�D����G�<u����4�P��&(r.	u�Z�����9���Ä��B}��Y�&��_2���@ �e%<P3	�R�u��쑢��L����*��άv�w��B=:H����)u���*�V+�-�^�8�7&��?cB�ڽ�"q?�_&�� ���>{ŝ���<B"DQ�>;�5&��o������XY	�Z��WB9�I��So�BɅs��iK��>[��-1��V~r�	�N�qټ;�[j@z�I��hԿ����	�����(G��3*Z@Y�t7�p��Q�0A��mW[@�6}JA�o��
�H	�z���~����[��;]S��'^4t�:�e��K��^�w��Y�rסT�%���[��uŖ/՚M��8ҟ^��PU~����&�fxu6��3>����`NC�&,���[���->
����UT�9;*�O�z6��@E�u�?��Z,^�'��	��������;�¬}W���0�9%��c��a	]�n�}2�-<��{��0HfhMK0l�����Z��<�P����ƸZ09P�h��w�uf'9�TL�g�	�<�5��(ŵ`��Q:�͗������:�3�~����U!�	�Q���.O��9U�	^�y Q�|t�VՊ䆷-~[Vj����J[0�3:���R!X�@�x*��e�zܪ�O��h��SZ,o'ؠ���5�Z�	�R8z g�6�~��2n|�#�tT�0�30��<�rN�04�Nj1MU��+!т��rh�'|`�]����~�r����f�n�����/�(���l�"Y0� �[IG�j��)�1���/�*�C��T�@�O\%J�AqQ(1�-hu����ޏ� �X�`)�x ���9�\{-Bm�g37�;H��h,�cgU�R������!�)��Ӽ���ٚ`���;����OМ�`��np���@hfZk]��+�{�l1���Y ��%��S_��� �	C1�������E��dc.��SM�Q��b(Đ�;>�a����Z,�Y�=xo�T��N-8�^�'u�g��U!!��%j����7*�q	�X�0�fxUZh[���X�軲�A3U�Q�H���*X	[�d/m���^2�:�H�4'֩[N���<��%����O�ȫ��0�^�&D�.���3�K����w�Qa�~�^��W�W��A�����=~�b���r��͐+��(-�xFkpW!Dh1{�پW�<��3�)#����P�KuHPh�^f����邠��H��9	YFLG�M�>>��*!�@��x.Kv���z1���!'�_FIö�7s��ါ���*a1��_��U@9�3\"���+�c��5�d������K���|aL@{鰜 �cA��y�
�TbT�G��zP�)� ÉȽ�DG�HsX�#�M6P%�t�}hb�1���G���f�),�1*&4�vZ����c$�%�t�¯�C���Z��IJ���J��;H0�@�h	�~(g�AV� މ�\�UQ� �,͇g%T9�-j<���(�^�Ϫ���Yz���!K��hu6�QI
(~}�7�jB�.;�4� �;nWO]�@7پl�=�1���x i��YI���M���)��1�}h,�g��ah������zO�8��%�6p�����d%տM���ۓ"�b�p{PJ�.Ϻ���o�7B��ZS.�"��uV��uX����ܮd81�<,�������蒖�@�LsiL���Ru���=OM.!�1�(�	}TV��wW�@G\��%�H{����V��C^{�&b��1*-��T�s�(�[W�����Eh�����[)�{���s �>�6�����@���!������D�� �U�����FN��x]��� V¸A_�i%�b�J�<��b��X��h6	n9^{��K��exΨ+������y�L3"_VWo�j���P��m��ݦ�	G(�/��nF�zj�� ��逴�쐺 �:R�.��%x>-�$Ձ��V��G�wM� ���çs���K�MZ�|M� #�f]�������a<����vN �mr�K%����?}t@��0��Y�wB���h�@��2$��z[��3�9��6x��-�F�P�w��1/� ����dW<�i���?��o�U��0�:[	�Q�G5Z 	����%c�Q� G�	r&L�Qv�r�J �!�"�#\?����J���5ݣ��.����y�:!�X�6���--{ �m���g�DL5_7*�f�X �F�u��E`j������� d)�Q��[�E����˭II�x�)��� u0oR���K��tk���A~v�\�����$��S������ l1ɹB\ �S�� @H-�*g����3y�A�DCA�J+�������!��gϐ���f���z �r_��$u	Ѽ	�E��|���+Y%�K�p��\W�Ph2%t�u�q�i�y��1���&GY3��5���-��i��l���e0�~��c[�r��F�zH��X̸}O�E��C	��ޡK��u��j����*�DYz�W�1m tgp�_6e��݄�f�x(�,X���(}&C�Uz���/�* ~|-@� ��o`�$VM%�6�����-~��Y�h9G��O��^���)���@�%�q(
V�>��[�b�������b�_�;�bHQ�P �\�g��y��鿚����������h��A��\�\�|G�+sg�����F5澋���A�O��и\HUo3f���XUo3Ne�>�8�V�|VD$�#��)�Z>��kr�{:	�h�>ފbG���@�i(yv�^_��A+�����VsE aD}�H����_+(����I��������5L�@��lא��x��=c���\zs,险�5\s%1��z�^�3�Wa�˚��$2�)��_D_Ej��}S��3�K����;��Hep���?(�-S���uDX��ؠ�M+8�)���G����ӏWr��1Y){AkU��\�B�7�o�W�)���a{9��&��/[��F���1�2�.��_��v����S�1pR��\^\�)���Σ}���~o>]@��Zg�����鉰k0
���h����^r�uc)i��1E�ΠP�X,�3�������WaOn�J�o������~����v�+(� '��J�:�(^hf���Qlӽkp��QvL�	H�Q9�[Z��\Om,�����~,��i2ej��N��CꊴJ��sN�h'y@Y(��h0�G��_1�!�D@�U�Ea��p��r�^?-9N
!D@#��� ���L��%^\�� +<~��u� ��΂�b�y���lx;�Ւ�N��W���'���C}B0C��}�r�� $h�v�0�0��u@�4X�8��/���N����y�(�;�Y���>'�p�`��!+i�!@\�Q���;ͯ�u�M>��c�u�U3$�i1���%^D<FW�QK~���<r�S|<�y*����/��}V��L>
a�^t��&:�u��(�����@�j�\����K0"D��j�7_�E�����%����_� ��)
Þ�$K^�鮺���!?�k�Z��zr��]�t�.!azBK�;�|�a����(�P%���|K��MK����[��N�\�p=��$R銓��i�1}?b��w����)ͺ�}L��|�:P�L6}O����b�B�±_3��P��@��v�0�^P@�-�*=�M@> �
S��/�X7�a����}H����~M-z�Ⱥ '
�I�ڻleX���h [~8`ef@CaYN<o`�˪D�h|Y//*��d�E!û�᥮����]Ɨ_E���ȗ@��4����W�	flkw�Ge����%QT�1���+���Na�O ���h�R������!�l����S��¦��������
ˈ�0�[����|�З`�ϼ��g~�Yˊ	�� f�]IH-Vk�)��S��� 5�dy�t9�D�L���V
��6"�$	2�C"���n�xT@�E �z�l �y�9K 5��2-� ��ú�K�0[*�Jg��4���?)���U��|��5�W/��]��ǣ@ʶ~ �fZ���e"F�w��C���Ae���_Xnv,�>���Z��k�W��� 0�n����
r't�7������DV8���*�WL����� ]�Jg#�	UQ	R|\!��&���z�} X):[�B̿�s�X��Y�Հ�zA�j��r&d�l�������-�(�F�4뼛{�U~���L��T���</Q�{�=��)�K��Q^�!��z��IPh�'�K�����<���p��'���&;��,XM-� ��c�%<�������^Y!#�� 0��y4A�o��S�`;F�l��vOi�U� Rz!.%�[�T57/������6����X��E�u��Ym�X1�+�c���:O{-N�.o��*	k%�1�8<�C����	/>\�&�f9!ف�&�X	1���ʄ��Q`Һi�s����JVh $Y9^)��(���������k�s��hE��*��T�p�H�G�M-`=� 8�f'd`w@���U*��g�6��0�/PD����Q�yJ��8���w;i?�o��I_Q��G/j��A�)�ln��,o$�"��0������{	����@V�����}���B�������r��.!��9>(ڟ�'�GA}F��iq�G�iYG�G�Q�x#��.[B��8��)/R�F�Z ��`	�N�j�YP$�hs�f�	u�_�Q�V@ ����h�T��E�Z��V��)��l���B�!��*���骟x�]J9�[p�)+��K�`U-���l���'����H@ɀ�Ѝ���ǛȭvH�i�I���x�%�g�)gi}B�u^�{�r\WDg�r=j16$�ų��!��,��_�$N����)`ꌞY9������a��YG��>��P� ^��S,5�x!��Hr�t����+��0Z�����\�_�$˃�ĝ�F�/EG�5��l3.��)��d�p��M�������G�&�t= �u�lXTd��n,D���"���Y�� �K_)Ӣ��>*a؍_��m�*�j��1�k��e5-�� ��K�I��������9�(��{~V$��{&"�4n���ז�r���C�� w�4Z�0w[�X6�F�]�2]��h30�Nza�(G�`׺8Z�@l\y�XX ��S4)��p�!l�Oh'�	Vi�I'^o=�)��<(1�����ZK[�F-~�8]?�aDSR��+�����~_�˅�њ�D�5ĠP�	NZ��t�3�0�a}��gmLݥ��-Z}�n-\���U��B*�I[K����|�m�HY���&v���敘y� �1�Z� ��M�u�\� �fR�*���tf��8�[�%�V�ÄB?�Č�x#��78��[�,#��&	��p1(D�������`Z�m�'��C���K�!V�����{M��E�`�g�'� �WЀ1�b'�˫�@'�@�Iu�ݑ�����_P�?���)�������.���kz��i������ �02/�%<��r���� �%c1fl�̺zK҂���fZRY���h� ��%I�����]��W��/tФ�)�����{G.L��ó�����Us~(��^�\2�A ��<����%��J7y�>b'W .N&1�����blc�t�n��!�h���R�y�Ha���?�R����4C�$O���W}u�w�%ٲB��ܠj,	8�Ù�S�ޘ9N��`�jU?��w�
��b��Uvc�>���A��t��/[B�(ͼo-��h�2W�,��; �!�W�X%bpREb�^���b8@�m(-j�Fo�J:����%=�aN�L@�VT^�=���^1x� �y��
�u���rsO��4�cz���#�'P�w�4�� �E?�(S� �`�U�i�wΈ
�h��2n��F���`�t�����D.��ϔ�> ]!�-:�+�����$o�vDX�����A�@j;g`P+�F$Zv���%ެ�.�Y	�w¥X�-��]X�	�w�RZ��1��BP5\��)�)�"�[����L���.M�� :������Ϳ�@ ���g���? o��'�7V,�9���ޖ�oh�n���*4>�a� ���1]�2�� ��W�J[�&��6�V&��B�������Ҳ���/zHy���Z�l�!���: �Y���q'� T���b�]�*�5�~�nS��G@�Z�ýT҅h�3�G��8yD%/�t ��U�kf�6�"'��#S��A�5�a�:�bg��[�����	؂�;�w�̒���Z�?4���^�7i|�ҩ��[6�a
X:�9�P�H��~��о1)Yt��x&��@o�2�v��]n�f��P���[�(2(��0��NY��ӬB�1Z���U@��
�JS��B~z
'x�%���@"�E9����e(��S{��mo� u	e\�dq?x�ŧ�x>� QgaK�0A��Xf;S�����¸(t�Ѐ� �����(�����yh�vtHt��s@^h �$INX��-E����4�Wg��4PV�WH��%&��I��zc���9 �;']��j������\�Q?�����_���[����2����R����>�!���=n�Z��T?��:p�&�M��G���/s�	�Z����(��ߟ~�`�΍�ql�67�јo�+���gy�^��t.���P���|�;��M_�Cpx&4%�h��W��qPn�cX�P5N�UQ�$�vK	�(�?^HBN�̞��' /[S��h�8�
`p
!F�`|�� �M�E��bI8��fU�#-	V�o��&�r��q���Jܐ��P*�R,�7"?���4�uy0�i6U�(J�F����q�Z->�&.	%Mp(��|@m^��&_���Jf�T�������ɥ�@N��9��[�͹���cX���Ж{���4�Ȩ�B�@��j�hcOt����6���ʌuan�$Ge;*+>��#��f ��1�!�	�5E*�Y9�:�'�^{S̆PO]�@��Tŉ�x��V:���ѿ,sh-�1V�p��O"�+	�~<]E�U{3��r�ia���[��j�Ή٘� Z�N7�v%�Ref5G��P� fX��-DV�qQ�b�d}�R����|y�L�p�'[�p�'?	Ҿ7d~!�|\28�11ba��01��RX�0�����h����"���i���v���'_@�);k$ZK�u`d�["4/�z\���ğ��P�
�1F7�qdI,&�R�^1�1����4FNMA��h������o�	a�wa��%X(������:=2��V>����5��Zd�^���Yn��\Y����[X���� 	�kw� �[ @��۽�A'}��z*���f�PR�yw\cD[��(��L��v3�0̶���^N�M)�_�<N0p>�$w)'�;V��~\z��s��TP�<r����?W���K6����1�3)^��췞q,��"`�?��IE���n2B�	aW*k��!Z��*�b�[b��&ʇ:��Y����!ux�|�J��%S���:₰hr��Ef,a�Y^N��?�]�]�%ͦ�����>�,��~���_��ɊG����R�	�*	�j�0�K���?��rHx�z�%����0���W�K��h��,/�@�0��j7h� T���k{@�0[-�e�Z������¬'q�~�H'\����A�0��Q	���]E����!����^m�H���V�h��� _R��眂��<�*�k-p�0B"B�'��Tz���4諕,?)˚ͯ��Y`=�E߀Uh�I�HY�ف�`Eq�PM��u��D��f�`_�ʾۢ�8 V�0)��*�Q�:���C"z0�p8����I �fQ�~��?��[
��K�Q�><X-�	hyV��uy���f[��	[�'����:�x�pQ-֌��1ə���`A�p���r�i'_�`��)9�n�^QU2�^��`��.�[��e�J������E�S1��ZK�3����^�����.�����^�#4�'OP1��\���x�f�Bo&X>�)T���hI��;'5��<.�']����TN��|�{��)-��4i#�����A."�uA�����0?P�d}� JQ�:j���q������95`���dca��2�Z����Q[��R
�H�0P)��$4Y� %�����C�R�zJ �}>nv�����6�L�)� �Bo8��0��bh�~�������@q8��Dm(UƐ �,�����!�(�t�yK�'M�� �����:�&9PW�hdOl0[��e� ef��_ V��dW���jH "��U�zy ��O�'�Zu.	���-�T�S�0��B���#8en�o^!�U����aYt�Pv��l�\_	�N�8ɻA~'��<+-���3�
��
�&�(��x�,x��h�c�N��;�DvMɻpk�C�^1@�U)��6#x {�/�\�%W��Or�20<�:�	[P��,V�=[f&J�haank~��<W�Ǔ@Y������(�"��&�R�-�?�����	A~`���D���죁Z-vJ$,:���A����U:�R�����)�Z%�Y�zGU�Ԑ`�l�%5 <�[��U_H���w��x�����������UV,� �8OK�?)P|��3����&BLJah�F�0~&Pɵ�v3U�<��.!�NI�5�F��&�e�@�Q�?	P�(��:;���� \�_~sM�m�71��4�7�>��sr�|Q�d�zl}�A_}���e�goR߲�=*��WfH�:+�1)J�|���A� O3t��f�0��Zh�}���:^#S�CG,��"�5}�����1Z��4�ũ�:�c�
,]V������������K�����(˧�Uf�E0{^( �(g �(�ֆ	!�4�ķԈ��& �#J�����+ �(%�Q��&�CD0�N��
��E.r'�@���)
*����A�'2e!��2>�`E@�``$#�[��<�o�(�4 �9��V�T 	.�P)_��<Y�Ez-?x*qs)��@�Z���-/�x��H�0�����p%��~��1[k�����:=1 �xvIB��	�tgsݡ�*��/�a�4e?�\�����#��D���+��-D�HN«�
?�XWT�QJ�=��Pi]ʮ	�	�HWnO=K6E^J�_ez�����	��};<�)�κ�aN.��{#-�s���~?��h���2�)|cf������ΐ�10�W�Є\���h���b��5VT���-~phX�L']�R�%�߲a]�|i��WA�o�&��PjEs��H�m�S�|� 긱�5-�*U	@`��� Ÿ�F�GODh���ȧiF-3�~���l�S��6�@����3$�AV�	k�o����F0��_5!�fi8�ˠ��I'$mX�;h7[�k��34'W�u�F�� 0*˰�5��}�
�L���`W�Vd��1k�����B/�X�T��Z��N�LF�h�[s��P���p�_�7e	^j>��'���樊��@R��(�Z���v?�� �0�S���[���p��H��1��0J�qyD�	!jV�iv� R�yv60�(�*�.�\V�'X�;S�	�R`U�/�v��- ý��a�� ��E�L��X��5?{�m�vG�-@�շ�OAhG;3�H�*��>�U���>D��ǿ�����^��=�*�q��`�����X���k�Z��v9�]+��?�)�!�_3��0[�=��:�˯��$���� t^�yB1[��+����q�^;;|��@���>1��0`�5�?}yh��-[���
$��p$^�>@({�^�Yw� ��F���-�+h1-h*�%8#�R�&- It��㸦
*|�Y�a�8�N� -.\`�=o�a2K��A�)�,]kPD����M0zK�{�'�%V�@I�ʔ�l=�C�5s�7�����"п�@�ہ�>��+�"�n|���bϐ�G�e? 8�P$eI�0���/E�V;��d^)���M�6��HW�%&\������1����w/�Q��h-�fwQ:e^���U�)~qY��BA��n�YPݹyj$�3[z����#z�n��0�����u	�5�;]|��X�u'f^=��盥:[q��^��"� X��{}y�HC�fH�8-��Tl�x�BڭThh
�	陰|����#)��yR�٦����+�]G��@!�E0u-�1@f�&ĳ< �^�����x��A�?Y�RC�O5��4p1���6aqCD�rO{�WnK�@���j.He'��Y�p�h�]��צ/�0t	�%� �RZZ	�4���w�_�	w��=��:'6_EYb݇D�.ur81�c!':�6I���j����,�}��`��@%�D�K5��o����.�h(�pc�Y���fXj-�_����+0ŅR8�^�*ZX9�͒;6˗q}���~'�^��%`��b]T@]I���4�BhU���N0�K�=C@�0�1�[�������!�h/5E�r�!�aL�R܉.�X��@�\��Q�k�q�����G�Q@�|���'���1!>�UzK�t�'��kw�q�P��cTSB��I;�~�0S�g(��e4Pd~p�����`B���V�t�����P��fk����J����9?0�#mL4q<��DrD�!Z�,�U�c	^/�D�ٻ�-#N�4�!n����QHCv�d�<���M�:7�X_QC�׫��z��D�ܠP��EeoM��A��|���+-���T|P�Ly,e�&4�Gki�)�j�du�@- �.|���� ��Is�c�� ��DA9�˶�"�V�`?6/�nb{����9�b��|����Z��,�h&<&1�{���_j����8�E�+f�Ld	���|n�V�mf%5��S'�:ݲ�	W�p��$��ƺ1'�]�0�O���z>�#��� j?�(�:�;�ez��-�phWi��ɼ�d�;18&��	?_IV���fC��g.���n�
a�!�)�?}$;��#��)�EN���
mA���{O?�o�_h��Dy�]�( Z�F���vR��F!��c���a+�����#]�W�tJ #�
<�ÞՐ�1ʗנ2_E��1����؄�о�E�X�:�ŋ��O���d)W����_F��7\����Z ���!H�y.����3�4Ɖ��A�U^<ʚ�50;I^�A�o��[蓂���L}�5�*Q[df;�K���Y�v��@�E�p�% Q������9��y7V���2�	�yM�ǋ-L[(®���[��b��T������E�AK@S�'�QR�P�_%$N��iJ���x��H&wX[�	�� �ɮ'�a9X�g��}2,ĒB�Һ���g��PK���b����%[��\4K�2hBh���QN`C5yY�^�br�v%�IDcHV-����!�p�[�<�E� Pe�	*���/�%�S�ڪP���������D*̈�j 1/���������J���֨U��R�i�N�ǬX�z?k�_���1A��S�Z�ׇ�@��� �<K^�-�n r��W�_h���J|�(����a����3�e�a�+�硤n�йL3^\I�J	�me�@4�T��� Y�t	?ZQ�g!��K�`}� 4R���T�\vLr�g��|�@Z��(/���@y�u���?Ck����%���G�4��&���!�LD[/!�P�IlO�.�+���v�݁��6co��j�a���O89 W��B6g)�|VP��$�=�/d�x�ܜ����\��5c%�H�f�N]DN	�a�T����t�YA��,8�C�@?�Biq:���V�R�h�� ���_�=ߋk�d�JD�7�U[
���k�p��"nAH��6�f�~���c9����1(:�`Z/#_�]�@\5�*=.x K�'+�p�0	����~$�*� s0-��\�8��lI@H�%
�jJ�Zŭ�6L-ǋ~8s�!��O0\qQ	N�P�"�B���n���~��p���Wdȗ��v��۸�{���c�_��c�XD)�������M�O��le��즨g��^�����	!��s�*.�luQ=��v-�NxH5z0o3��,�3������� e�o�A���a����~� "�g
]�xğ|��X�/�PZ�[��^��1�6u�11�h�ۘ�U�D�����i�gǬ(	Rw�zyH���g�m~���Y�raz�9�Z��508p:��r�!��(�-(}]��פ�h��V����洂Q��NIWLp1Y�W�����%�tq/��X�uL����]J�����Q�(uY�\_�-��	O4�0�����Ӱ:U�nm�G!�]�V����i��0�CQZ����Pڝ�3m�n�<揶 ��C��;��ֹ��I��,(������i�:�m)y��#sp�� �Nh!�)˽ �B�8�պ*vT5	�<@9��-͘�/5�li���Q@���	��[u�T5>^�x!�	�H�P����~d��2#�)���4�35wsW3Ȉ�)�Y_P`��Lp	z�d�	-��$��,"n��-PmO���$�	�Z5V�./ �*ET)�1�؀�r���CM��	]>�|����Ȁc2�d��!�&���!��K]�T_�=v[X���Xk ���1�H||ZE�t��P�g���`�,$�=� ½jMr: E�ͱ\�%��鮒���`D���l���a�ҦYƝ���`r@�`�n�|U,�ABD���c���A�8<�W@F�w�N��d����G��ǸIx�)U���Sk���E�eQ���UW��!R�?��Z�F���$bMi5`��j�� A��)�����.!��`6N������8����6>t 
��X�*[I�ϥ	� o����0�5?u,�@b�f6���Ⴥ���7/��\-J�v����� �\�(h-N䦇t�:�1r�	�ʄ0-`fV�B`J���`��R};dUh�.��r�4�f\H.�X��J�Wg��ye�8�r ������;`H`�S��?\�����̍X�门B`��[.2*����W��m��1�_!�]:�S��r P��+�R�b�1�]�@�9<�'�3��@�zv�>��3��&0����_�H���#w�E9$�t������j�~%O�`8��'=q��)��>�&�U�Ji��zBG���c���1ʃ�Z�$U�#���2%��<��Y�]�;�1��+������s�_��9gф/�{=�>m����x�R	�4��ٛxs����w�� F�H~}?�(���?I&g����r��Z�ڶ���r�:��y�����{���B��	պL=7l_z�����R����N���N���(:�Q�K�Ĵ念(Z�#��B u���,v��q��@��G.�mQc�Bx%U8n��L>��S�0�˴P�"ClHc@s��j�b��1�K:$�8	P��� ��%�"�B �I�^�e��Z�}�����f�-�+�� ��{Sw���Mj�;��s��sK����O^�q�W|������Q�<FE�����h
��Qh�l�u]M鷂@�5���[�h�]cvLJ��*�<�K1���W�됩h~y �=X%�`�	G�U��ڃ�6|�4&~p��O�\h�ҚW;	�y�R-5�_����^A2s ���P�&�Ѹ  �k驈��_v �p�}J,��^��_���+.���'SH�*O�@�p�j��hi������>�	h:_����	%x�����k�_��B�ݖ��y�i�*�{0� ��%��卭ٯ��)?R*��i�^�m\��	��Z2�P�	�-�+��H/��CK	��e%T�H�~��g�LX�� v�Y-Z���AC�q$)� yb/��J��;-�S�?�rf�^���E�;(�$`�/-�Uh�M+�1m�ZGj��y�ې:6UG)���DsB�.P! KX&�vN���U1Yp���N�F�p� h2�����8�V\&)�%��@Q���*��"�6K��:��@Pz�r�^E�H��q'��t�V���1Յ$�oȐMϙ|�2\O�G��;��P���0��`�R�u1���;�	���_&�n�S#H'V�=�2-kM�@����F� S�h�x��!auSz��j@5/�v3� &�X���d�[���aC���=���t'�X�҉K2��ꄿ/H�8��Z��"z����|R��#�Z��0�[�LI�'��E���1� ��f[B���^�v��0D�uWyq0�$�X{HW �G<*�ܗ[��1�u�fW���P ����$,����p��<:/8qr� {�41�^��b���h9�~1UhX�=u�8>�%G��*IA��>��Q_{TA�J����%02~�!M��|���a��v�B]49X����KԄ��	U��Ew�� �oe�DUX���C��Q`#x��(�{ɧD�_��1����Pc� f�+���#^��F�� �S��Yq餕�u�&\�q���u��y[���A;�W�O%�[������+�mfP��0J����sJ/�tx�q�	龶��3� �}~�7���[KgĮ���	��2AVj}:����]��<aUh!�P��i�H��Z���K�G �>�L��2MT]��ivef邰����F&B^���%�-�r	�LN�Z�2�������14RC?M����O ZZ�q�sr��o��ɥ,j	8J�,ٗ��%���'S���H����!�U��9�Y?��PAT�� K��'AnG��%o�I*U~g��Ծ�[���\P��a6P���S	��V��-�~FNa�V�!�_4�+<]�V6r�O�����)�md�����%ܽe7�C�qB0{Isx��c7�� ;Xh\BL�p�o�QjQ�(��Z^����4��K��_:���5C`~���.N	�u	���y��@�����nB�p����Y��t���(�5���P�Zh�	�ݖm/
R�mvzW\�ˤ������I'�ݚ!v q���/�[P�5�=|���	�j/g��!'�610��� � S�-&T�\}�\U�ƥ�U��@��ʐ��P���g��3C�n1��!��06�
^��!�����Y|	Z�9���+��(�	V��p���n���k�A�����4i�
Qq����D�q,@d)���ũ��t±�A-��"T��M�E hi�7<Y~r����D� ��^��Q���	����wD;TSy»]w�yI}N��uբ#ȉ���n���_���V���%����J+8�)(�R]�RA�;�T� v^|_��=Y��e<2B�hOF�������,.* ��LG�vj�Rt׀ZX[NS�.:P3��̇���>FY����f_B��\�6@�cT�`l�Pa�01��(K,�
�^��� �h+;[�����`��J
2�23�"��pVV	�P̳�vۼ-���'������M���-��tA]��j�;���� ����)�;	�|�"��Rpm\������W�a����@�uI�n�	�kj2��餪�Eh�\�r	ێ�WѨy\~���������9���] �0�,x7�(CfS������:����> j����PVK~������1�X?���4ޑP����>f{J������L�y��3�׀2�]��BX-�Ӗ/}��*	�d�����������-obK!�:�S �*hk6�K�A���?�g0#�WK��5�?u!�®��z�ՂT, �
R�!)�fQ�^��0�CY�ق���� �h�6F��C���	|b\D<2wr|?��d;MyCN`��.WZ0b�$��C:�M'$'>ը�4�*��0��uB~�yh�}l��+����/F_�엎3[�)��0�44�,�og�P���Y�^���$h�)7�n��$���[{��g��/�σ���3�K�����MW�0M�"o2b-W*�L��D�Á�8�);��`�ANE�|N�ެ �;iu�4C�j��7�N��;ٴ8]���~(���q�Y�X>+)��|�H%� �\
6/�� �҃��9	���(^g��0��X� �e���Ь�Z�@)Vh �Fs]�x��x��e��	H	�zJܭ9�����'8��9�)fY�"����z[U��N�q5�Y��S��n�=B�&�Q\�PG��N���R�_��|�`��������v�~0b���^S�0]3H�M���Y�h�2�K�S_�C�����!�:.�90�\���r�]X�-6�.1��?����Z��#�FS�
��L�si&�܂#	�b���6A��}��_��?|�Z|�
a �:�#��-��	�X��#؜�:���O0^I� ;Ɓ�Ah	K��0����;>�m6�����d���
 !1Չo���b��s>>����<�O�O�*��@�0��i\=<L>�_���ay�l1���2fI;�y�)�}P��('�ۭZ�&����n��s�,"@�붉]�!љ�-8��|�� �v�QZ��9<��� s=C�GZ^#�^HG:�J�H��������b �B ��90~�PM�5	���д ��Y_ܓ�z�J�ďRED���Z����?�1�Sp��a`���Ci���-��\���Y ������[R�C�����|A>�0�V}d�	��!�w�eZu� ��ˎ8D�� gL�NP���ײ���V'_E�@��MK<�L�(�� �80�ڲ�R����tB����q��`�n�f[�� \��|ch����3��3�!z�7u��X��9�2�~܍h��5�C�́1��+a��-�=XK� ;h�|Z�l"`��1(�gM;p'Rh�x�^�
�Ohu�����)o��ͫ�@��dBW"�%!�Q+b7����ӆ B8 9�N@��@�%X_E��\L�Y�v�����B�sK����6��3ʴ����<%J>��	&�����]!F{�
��L��/���iqG_k�����KC�&��!���H:��b��p^���`�R�*s�p�EH�3+$�JY�*���>�H���˴:^ґ�T� -�i�S	�Tl���]��rĂ%��l(&?�@'�]~�<�m�;Z�;���Z��ph/�Qf��~�t�^��H��Lc
��Z��Q�٨��h��@�� [�iڐZ;!��\l�&ń�p�9)���)Yk�����D��հA���d:%!p�J����d�;,�����\,������t�`��߃��A�D����|�)��ެ� hH �:Y�Ơ(�hE`��� O�]Z�	�B {�_�E�GJ=` �����B�n"�@������;0#��
��91�Z�8佄'���'/�Ѧ �f4-X�	�+�3CFÙ���x�wI@齰��-�(y\O�֨��a�~�]��ܠY�X&.���>:\���[�ց�W�,1[�&�����h<w�U�/�vx4a�@�w����!�ܖ;�@����D)�1�p<g�� M�_b�@'G$:�1^�D���bPҡ�QS"�X��G�%bB���
oTU�0D��K��	�l��� p�)×x�Z*	s(UF$�v-��d�h�����_�S���!K˺`��	L��fZ�����p;��9�9�/_Xkh�-P���B�2��`��$:��wL�f���p��`0��&�rl)�Sh�?�X(����+/j�(����v`X�� Z�)ڹJ��H�G*} �S�f��ޗh�+P	0SAIuzu�Ք�LrW�m�C�-ԫ<4�%����Z)��o�
Rh�@���Ç��E���ԧ�1��z�I�[�Ұ�#q@�	O����@��_���"wV_hr�b���@5΀��j�)�1�V�^�@(��#&*y|��]!<C�A�@,\}-^���9fSh�Y����H_d(l��v,��Z����:��)��o��^/�Z������&,�� �!�|���3���h(�	��i��`�*���YMw�*3��9gp��7�&�#�:�`ŀ8����8��$�>��]�Eh[� ���i�Q��)a�r�0@ ��Ў�����<K����GH\N���Tm8<871������-�@Hq�*�����K/)�_S�,:�Y�4�h1�Rox���?�@
�l�-��2��._��'zC	I@X� ;1��̕�WGT�F�o���1j�.���_��h-�{|jg��:q��/K��l�(�n�L�Pw�0�B�3)Y��Z �%2X[��nq*�o�n�4�����'�tP_'rD�Q�Z�;/P�,؃�5�u.��9���G�U�5��w�D'1��X�->y:L7t�d�u��<����!A��.Gʵ��� ����T�	�f�A��Pu�oIJ�%�ч�[�W`�}�Fj|�M�k�A���ڝ��1��Pd�!�^ѧbE�{v��'0" ?_����(��hx��/�-�/t���,1��l�댺Cy�b>0؂H7&q>��=�;�����[
��Z�ؿ�� �T6&��E5�!�Z(�Z�x����`��5�#�~b^�`E�$�� ��4�n*A���6�X3�~�۽$\0q��>@}Ō.<_f��1�we�S�������xD�+�x�6�-�����Yq�R�G�䗌����ͥs�w4�n=���YV�ԇ@���<���X��_r��B󪜼[���\�.����鳬^^��9���g+9B��wd�[5�i����T<������0��ƍ��-�R~%os��=i^ ?�J�x-/t��2�0D����/E,����<�V�;�w�>�R���������,1�0�2��8-FP���\�R�,$Q�.���-`ջ�so�*���[����bz!��E!����/}.c�OZc5���/����B�q��- _�U�h�����h@(��KM�� P`y�R'E�g�+��h��H]镁�	���H�ǭ>�b2���T����!���H_��ĉ�뢷����͘� �`
1��,�~'�ǝَ`�Y8I#)���W[�s���_������_%��1;�}�5�v��_��%����S�ӉLZXe�������q����E�\|X.z~������ׅ����!��Q[���h�t:��Խ�1�q�7�3>�^I}H�R������Q��0����������Ӏ��B!g��Ж�`E"h6�<��	��S5׺�O�Y[�e��xК/bS��`� `����ܻ5�}���%��q��(��FH��Y�h[��R�cIx?�
uo���Z�E�%׺T�����;��Z��"����%�@��h�B#pV,�oH-�I'wd��c��AHN.X5)1�A���!�w�1͈�n�xb�H#�v�B5Y`:|�?�Cw��ڝ�+-&r��8�rE}K��5���j����@�DB�1�Dj$�8i�x%���, 	4��]p.A=�S\y���U��.�<)�]�����w�^���Z�}@o`���� J�Wv�iAb�ok�rU�2Ŋ�ôL�ā0��@��/�����fQ��b�8h^zM4����m��n'V����D���1��:s�e�M��C�B��K������pD��B�����M_aK��޺���#�i���D�#C�2�)\Ѿ�\I@�P�-�%���_�}w-z�T@��{
JV�I9��/�����D�k,+��Qf����+�0.9�!��5�[m��A8�adcy-
���䌹	:�7�֠(R9�&��tuIBU�'^+� �b7�DU�YX=��934��^Q��.��q��瀸V��RF+��i`�_�u% ݹWRIA�EN����_~��-�W�����[��ۯIZ�P�,�^v�f�\�ծn2������(�l��ȲAK!R5H	X_��$��V޳L�����ˮ|P%Y��3��	l	H�]� ��@����)Ϳ�O������(W��i@!�Ǎ�.!4h>~6�(q��9K��=���8�h�5���"U�y�Œh8�$`�'�����Q� ��{��v���Y�[��`D=Ce��$��<
0� P��f%&��ehr��9`{SXpG�'1�ߞ�,��A����*t��=�z���G��`GT52�~n	�]�_(�y�/�M��UQ�a1�!٫`(Q^�*(B�Ol�c�(�j���wh��B�|[5��,Y;�� �������f��� ��CUm�$�I���'��Su����%�4����+�X��;��S,�X��}�u!�|� ��u�@1TP��5�U�C�ؓ<����ީ���p����:b@��8Q�允1�K�)�<ϥ��=���ú� ��!�N7��v�c��͂TO`���w�1RB��TZ5@���{�F���X-I� �,j��=ڴ�GS3��M�d��U�j�ȍ��.z�{�gG�X
�ybe���C���j����n]�29�g��G�>�s7�F$G�ȶ�D���1�Ѭ�@��Os@JN`?�"xuY0],E�-�g�
��)Gm���2!��HS�A�k�;����g��	F'��+���U�>��&��:����3x|:��&�ч tp�F��	�� SV1�������-��A��W:G����dg
^H0EY�>�x�L�d2��-E�K� ��H�����f��yQu�<�_�^神]�"<EtP�[Y�Ո�A�(�C�A���"ޣ�d^h�V�Q]@P�	&�܁�NR�C�5�;���P�|e�oq�%7�K�mLV�X
�Gp�	`*x��a�*�$F*�g�j.>=V�,�,s�v�댵W龃�Q��Bj�>����ODj�d�WP8�D�X�����$A��yL?���ޫ,��$��D0�_{�&�-)�/�ڊp8Gcݸ^ ���p�w�{((l*��$��,Aq_��Z��\�16�u��B!�~y�����M0��-`0�g`���j�\{I-� %X��T�r���R��sV�W:f��a��B�f��;a=R��C�.<!PvG	<qλ�"{��n����j���|���{��Q��P>�X���p�x����^�;�S�s/3��Xn(�%(��[h9b=r�DJ��nz� @|��C0=�%���ztX��4���q:�EMH�X�)O�*9��z�jb��U�kx��(�ѵ���
�����Y)���ܪ�՚<]�k!��`+[Vh�\�AO�)���ƀ�-��P�`ȕeđ���LN`�Y�G4�e[���S;�'�W3�E�t�-��\(n^ m�\+ �N�:)�!�!�PZ�h'��wa��u��M�*�D>��{���S�1��HV��T�9�L��h���u�5?z�!p����a��%�R?�L�#�G�	5�/h���?k)jW٤@��L�x�D�aX�Щ��b^H#�+3���lT����0j��>����!þO�ͬ�%ƽޣXcOq��W]ϣ�>I�	�6��F��3]���a+V@��2'Ol@�	4)FLA�U�D����_�Z�h���Q`���un*7,%�h�C^r���&%�L�	Q��0r
�Rm�� �v>)�O-h@��0��e)9�ׂU4	o��K��+��fh�Nn^�}���4�ԶdY��S	�:Ȏ�m�P�Y-J���ku
�!!ʟ|KU΅{��1�L6r.�i���>��vL�raapj�@X�^�-�.��`@+�9\^A�VF5�csa� �1غ{;�Y�L��gs���i�*��ӌ�_�W�� t��(�8h2N���?B|LQމYj�v9�`2�ø�Oಓ,h��)��'P�k��UW۸%5�yE�I �7_aY��G>�q0H@X�#O�C��
tZT��`��P��,�c�`�����?�l�GS��g��C)O���<w��M@4���x�:�lO�-˰�� ��>L!��4d����0�3�%�}�~H1�#��բ�k�Ы	�l(�U�ЉP��Qm��ZwWg���<��@��-C8G.�p�߮#��.Z�í}�{i��!?Yj��L�	d�k�ǒ�w�g?�}�����_��@����sAX	��K'�����\�V-"�����&	 �)�1�h�:0�Do�`BJ�#�N��J��Lc���juh��q,�}@Zh����d�R	f����i��W���pKB�-�$R���2qO�}\C��HtL�h��We�b��@�0�[f#��x����o����}�	�g0����,(Y�h#��=!"-yܠ��|����/^��<�����[)�5�2�-�b:��h�4A�$��d���C��,Ó&�UR�8���Bwh.2S ,Z+�2��o,���A@�$��V	��_o�����&+�Ŭ��J��������M8C-���	)�[�/R k^12��ݑ�
'd_��4�_���~�aX�ގ��4�A�����r��ĴT��c�`�X�IA�U���o�!&)گ���hB(g[����O|��tG[*���i�v��P�C^/���� ��N2���%��v��9/# ��׀�' ���%��Z�8Em�2Zݶҵ� ��� �[UT靰T�N7�ӱ'�,h�4ƪ���[0�����(���d���[���_ho�j=���S'UO��-��Qm���x����c���<e5.X������j	��.�h�G�p �r(�fX��[�h�V�d�N�!S\ _�[[�Ղ�1%��0��-w2�B���(BNf���Zװ7�����A�����.K��S�$Al���S�	p�Ul����n��L�%`����]���@5s�	�)�V� V�p5��OK�@Ɩ���GA6�v�W����Auoq�_eaTl�9�Ҭ�^������y�k�;3}Vݧ�)1�^1�-�9�g������H��n><��n��#�bU��8�F�r^�bQ��{Q�|��;�~���#O?�gY 	��WF�hC��-��_��/�RD�㪎v�|	0�'Z�
"/W}�96!���_�x*��ٻ�|�VC�Y!�	�����P�	�N�k
dzD�3E�d��c��B
jOWje�
�U	N��Ƥ���}6�ZP-
�.�D��¿Uu:���=93�kA`�k�(�H�'|)�h'�	��	)VU%�j^��R�d�h?/�JV*7��'XQ.-�z,PLJ�o`6�`y~�3�����UJρ��[/ŗ��/ �銈�>����/*��b1���(�h-bc^�`��>��U�^� =�6�0E� ���!�x��
�H�^a�づ����*ـ6��	�t)�_��(̩D&�kE+��_�g(�	dwY���[r��y��/�!P� ���|�U�`2�� Z�'�&pX��& ��I 	�����4��j��BN	쇒�zm��L��O�`b����acAo�l�MT�����2=(�p/����""Nt� �?>�muX�Li<i��)�xm4.�������`�/.K��'Ryg���Kaڽ\r�n�@�+,iȠX)���b3P����j����/�<X,Pg�h-- ��u�x��[k��� �h�lw%�B���#/�?Q�`{���	��Zo���}�m(`�|P0:�>-�/=�YT�_��0��n���o�XM%J/�a��h�H�H��I��� �?�ȕ\�!�R��w|~����3<�k��QX��7�@}��a�ռ��hX�J��M��'We����S��)L�W �>+�;/0qFoơ����}��[��-���^B��,���(��ӷ��O������/��ˮ�N�̰�&���\(f9��y����Ȁ�t<��԰ ����pz�w�^��)�������dv���1k�
U���� |E~Zhdg6/����'H$̈́y�1T��}j��@m	���<7^鑯b �۵6���?�ڗ�m��n�P>�kX�Us�����h`zS��N �+�����IJ~Q�D�q1o�|�	o��r�Nφ�ܳ�������߅��X�!��oR-�bj���Ɏ]�,-�raY[S���� 3�c�Z�ȑ�Xz�p��L�K���6W�V>���$�q&J)D�����0��/"�� ^��4�Y� 7!9�������JW�"��ulK��;,��@�5[��a�h} R��%��v�Ƈ�ث]���
8j_��U:g_dc��IW%�Y+k��h�DLXR�w�	�Da����ݨ�k.�^���W�-w���u�A�Og]�	�>�N u�F�9��\�)K,\�`�� 4|��m���q[ Io{)$��񖃩�~���	����ŏ�}e�7H0�\2:�z��]Ƹ$���՞ͧdH��	�2�R" iQR|�I��5�� ��GU��#T]}4˘[��#���k�������.v3��f���g�PXa����_tVySk�	ɴ^�%�4�K�y�X��f�-8���Za_�lh�'uj��!(Tսq1�U�T�k���bk�����%����KP���m�q��^��'��!����ʮ�D 0h!3��FP整�(��x�@`̓Q��v0��
�l����-��B$[4}����^�G�ߺ����8�\Y��Tk�@(V�1�\!�`��7O��k�@GM[��X�ޛ���a��VE���yO��j�KPf�XV[��:�����
0�1и�3c
�����*�O�1\���&�y���\qҪ��2�h�Z��DP�E�
����-�:�m�����t�n\��h@�ݠ�0����(|^褨�p��N?�!�ǶD�y�Ph@�s�u��H7S���I';hǗL��S�a�$&L��e3�xu�/��hd/�tР�Z���a�Q�+���XI�x:=�
	�����+-s��?�g����'u�I�u�@S%��+~5C�i)�	��B_�VQ����-�Qh�Y��U���=�<Z�)�1$�Y\�`^R�i-IwqKb���� ��{(�S ����fR�W���[�`���%����HW�	�Ȧ]�����D	�������_��O�\�~��c:bUH0Q)�����e��Ohq*����
p
��}�x�a��|���Uh�1�F~������/>�i�7�Y^��|�o#� h�]E��!�= JR��&��	 bX����v�*�kN��x�a��yE���f@y�[�L�*~=�������	1��M ��S�VyxTHW�Ѽ�폋P��{�G뾶�M$��'�	�k��!n��h��.�M-^> ZRh�/�� ��A��\�5�9��^c��[��V-l"����\:�	�v��h(Kl� 瀸Ë�?|_�^Q*@/�2�U�Y�RS�@R�j;�G �S�8 �D
+Z�V���&�)��_�����	��K�	�q R�Q���Q�k^%��.��'���E�a�n�r� �S�"5�%&�h�	����-C��.�Ĳ��-�s }I@5q�Ҷ�|�Ʊ4jTH���/|�Xhx�	�Y�@|@7X���br�o��!-��i��wQv=&>R�.7���a��~��H�|I���xJ��!�H5��3CO���W�~���P���@X���4r˔�ͩ�,[�|�4Ԙ	���1�)�!�	�-/�<���DOk-�%`oX�`1���V-C���~���/����I���Z���O�D'���TO��͠�N�֊v)�:�L��[���J��N=?N�����_�Vk��@1�D~���Ra�@_�W�&������K�T�6eC��Y�N&�84�,�Lk#u����`x��h�܏�XO�/�&��O����zz5�޽Ců^X���}�U������J��g��Wej��^�����w�"��u��W~(Z[� �q�w�2}{��r�x(iى�(�,)���[K�A�nlj.�CĒ8�0�6Q�O�;�(��(>O.�zA>�� Yh�8\e�rך`w��(�y����M:5�I�-��n���[��	��*�=�������0ʚ�P�9va�Jxk�@b���T�4�@Ph�,���0oj��	=�jn��_���썒���4�O�r)�_Q��hm|�Z���-R�|��Iz�70�8.�JB����?Z�Vc5Zİ�딐���<B�xv��Ş�C�51�`:�	�f)L<�:�}�L�}I*<ў�K���)�1�pXaL�'��+=?ROA�� ��E�0���i>�f<�Y!�F����� ��`����0�;�K��΄����1_U�
x�{�l},�|�!� F�1VQ��G���nRB?��(���{�G�f����5PF�8[	�
XW�.v��-�>�+�^��.�^ �`&5����!�@� 0��G	f�W��Z[y�%L��-���l"��E`U�M����<��L���n+B����oZ@�S�-E�(��\���Џ��Z"���|@�R��ӛi��N�5�^(�e��~�����o\@�����Ȧ�r��^h�֌I� 7� ��L~.QG��E�"�"�@N»*����V�t����b�"��^�w��������a����.af�	����	Tj@�X-/VZl��5�[� ��()��`��� �驹����cO~��*Pd�[#�W^�0��P�Oˁ(-]Y��D`nQ��|	���;�˘���-�b�@V�:��	�Y`�Exr$!ݪ�'�����o�. ��pG�a�h�No��Y�;���]~�}��q�oŊ̻Bc�s}���8^ h	�mT�%�D�A�)���B�q��񟤥��}ė��)�J�bSo��Q���h1@QX���x	SV# ٽ,r�j�^��'������b?��Ʃ)���"��} J�(E^�Vd$��2�џ��qfh@�h0��>(�[��8�%�Y4�D�j���Y�=�`���c(��B�n��w�RV^���"z(L�	ⅳ�_�5Q0��~C �(�fZ' �JJB�q-A{#�� Uh�	�~�.�^��K��	�r^f��MK�{A����	jY���
��/a�U�	@A�J)J��gʱ*����*O6�F���N0d:�5aE���:���-��QYL�H-�'���u��b�!0;I�	m��x7�Ӵ�x�i�$wz�7�tI'[� �nC�7��g8B��cP�^A�C���R��r.�\���3l�gL_1�`x�Z�ѽ@� �\�l��5�����-`|,0��p6�4X�}��|�x��ULI�U �p������5��������lzS"��(e���d,v���#�	�)ˁ�����j����/a���~r���؅;��h�f�I ���(���Z~�G��)AՃL'��޴yp.G�k~�p��q����%�J��a�]�4����]��i��v�:�e�yl+	�+�������\�Խ^	��R_�6���^2b	�ҩh�¦�8�5ic�U9h�W��J�下h�G{�QU�*����Q l
�9u�$�0����\<X��B%�h�ˋj�{�(wਿ@�hb�B��ѵtR�~B�`l8�]�{q9p�
�5�z�>	s�r��N�"�c�:��E0
�J1�b_�^鰸XQ��	�wfQ����t%%�?� ��(��m����!�} �R0{Ab�� !H�D�af+;M��=�8�� �༹��q� �~_G�������<��+�bLM.M2z'�:	��Ӹ�_��h	���u�͒V.��'��s	�G�u�~���v�'���f).�0�{��9�_�La�Q);�����t�d��9��ߣ���u���\��oZb	�,.�i��&Ӈ��"��0h)�x'T���KV�Ў�SXthO�Zu��,�2�������0�3^�	�H4��A���Ɲ	-{)a5�����3�������0p��p�� ���ԄI �=1}b����zH5�j|���p�%�2�a��b�1�)щ �{hU��;��>O���Q� _��PW4?���a�2wh��g�@S���9Õ����2�]e�X0�C��jR��7�0�,�ae-�l�Ra�!|p=��F���I랶��U ��l�{�����!�!��g���;_w���~x<�������2
�K!��/1�w<B�+�ᄉ�J�l�?"�b�D0�'�h|b���� ��v	��Y�K�y1�A�59+�M	(r��:B=9N��l0�$��\A!��o���3�w�o�@'�q	!�5�[���bx	%�Rbxp�	�˜�U���������؈�^Oz8�����_c�w�M;ć�,5Ბ_��3�(mz��)�w�S�l�w%JK����e�	��P��*�t�+� 7�6+P �}&ph
Z��R๛���,��d�]6j)*�5
�E[���(a%ʰ�u���W��!�=JE�U��P��@��b\>��t��!�B�!TjP�J`� XZfS%��x8���,#wC0���紀�W�����#d����%��b��Z�i	�V���-�=��y��q#����)0�c�t'(��A� ��6�h����)��C��5�'�S�,��	o[�o�o76���W%�(�e����>�w5�[_L���7hD`ؖ�	;�O	 @E,0!��@�'g_�6�vup�X[�����]�Y��Z`�S���7�5����/�b"ȅ���- ;[U�J!Pz
��L��r��'�pN�\�-ݞ*(�u�]E19=͒,���R��y��p�F_B\h�����V��~	9yQn�h�
&�����}��0m޽��a0���lu�:��@�� ���A�h�l�*P�<�[H�T��$�|%�c.�:dc�C:��GHw�I����IT�J�<1)F�H�;�,�P[lQ`�A;&�1�	:�|[����?�'������f�&�H�W^�GX�"x��u���[b�ؐ&��H$N��5�MO���PpY~�h�Y���H��5��#>�F��4�^L<�ӡ��P�Eu�Yd�)va��@+Vr�+���s:^�o$�a�V4) g-2��[<�%��!+�Îh��a���;�0���#gM靶z�yٷc3��(wK ����Jh��@8���y�X�i���iQ��0��u�*��m���Y/�Q\�\@��������O^ȯ6/��L,�h.cTH`�5YyLg�kn9C�]1�Y`OZ��^��Of��2&D ���Q��>�
j�=���O
@�'`�:q�g�|j'�`���"���$�3[>.Ua� -����>o@��F'�t�Z�+�����
��X?�x�K��!r�|�1ɦd��PS�����ZJ�5)��z c@_��O;��~,�vY]�S����w���)���k��/.�ݵS�a.k��z�j���MV��
5A���0I]_1��3OJ��;�JPh�C㷷�b��h�Ifd^6 C~1ѻvs/9�<S'�����1X�_P�Ps�v����5j�����]�'�m?��*�x�Sh��e���a<g�B�:��_tE���	P�,^��K]�+���F�Z��V�\B�S�Ne��Qh\l�4��1-D��+�B�촄YV�m����?/J\Z'񉽥��[�[hUY��<�Z��pÀ�X�����t�]��sh��|N����ϲ~�Nr}������3D��'0r�k�qV�K��]&���teAH��C���[��	UH�^ ��?�g�X�Z���3��=œ�ݳ���VD��i�m [��O� ���d��1���T��E����-�AY0B-[l|5:�8L�wu���pT���i�p���j~L�����!�?�����5�u�1��6������'_��������`��^!¸�%�hH`ZL羽��c�"����Ͱ���`0�D��4�I��C`�K���kA�S�[`��+-G�u��U�)��	�6����T���xJ�B��>�!Q��]P��~���	�MU��Ӌ%[�S�m3�X�'��� Y�x�X��KV�xb�bHs5�m�:�}��;�ʰ�# ��9����`ǉ( �O�����CC�'n�λ	L�x�{�05;"�B>$�5�-0���?����|I��;���'��j9���n N�-���% ��V�l�M} ���ԇ�1����X���?��	���H*|�A��t�3�t�pm5��B͛�	�^���jT[޹�I�{'iY?( �� ����?�l�j�	߉l~>݇�Xb=D�-�,�!`j���Pf�I��~]��H���1���n�_8�\Y�
O��)�����/:�r`Z�ݵXVҭ�����k���s <I)�Z^(����*p�PS� հ(�[�萞~����������70�[�PU�0�h�g )d_��cn�� ϣC�	Q�~U �,{ovq
��M��`C�.��x�}鄤�s%1���,�/��;�PY��4�\4��؂��d9���(M���N$S��:�c�3��{Mo(d��1ۜLvi�,��J�P�Pf�'@�\?AhM;2&<+�6�آ	�i���m�������a�3�qK0�vC%�K��h�[X�ↅ��U�>����&�ȴ)�]��;��N��B�P����≋�s��`S�*���P{VJ��>S�Q��W��~<K�)�:��	R��_xSd9ꯄ ���Z��*�N��v���O!J�7��AY��e	����}�!	�����U[zD�����/�>tf��r�'[��. ��Hٓ[�-RJ0�G\
:��A��c�Ė؟��v�����Z��%�k���P��8K�E�$S��R��{�*�0�����`[J�2@).x�K#�����������y���(z�>9�{�����-�_G{����I�L�S%�[�
���_hdw�s�A�\ޙ'MܒW�g̴<�!6.�o�D�wJ������|�&5�2��}�	w��O�8ذ���j���'��<"�n�#J�^A�e�0��:]������D����� U��	��s�-� �-	���Y�&T�4��Q!�.�1�*�s����H�y�K��hdb�"�_T���k�z�;5"�U�,�'�@1� �z�c�T� �8fhA��<��	����R�h_9�4�x�|*��z���0�0�����{�p�|�,<�c	�@��o��<
 ��¤�԰Q������i�[=���1�~!<�n��k�y�	�`F��'�'m�1�����$S�}0�������˝O����^	�)����G�1�z�-X�%�Sw"ŉ�V���͆�����n2'�}E��S} #/_ځ�V�C)��(k��W}�s��'!�{�%|[�	Thi]p�	2mu;����@3#v	?㫌�]K�?��d�CQ�!=a�����M`�z�lQ	 �1Z7Yhl�N ���owO�����(�h�9���R���斐C���a+o�l��̣��L�EX>ȿ�x���Db�_AD�]Z���q����W�
Wst��yJ�ct�J�{t5lG�A�c@%��w��&�=�i6�	�P}r�K��{j�G���	�� �b��h<�5K]�@E�x��Xo�0�;Wh~zN_����_�����9�
�s[��vC`,�mb�NuZ������u:�u�]+HabxAWṽ�.��:-�	���Y��faD�z�V�AH0�_%��r�w�gX;*�zw�^}����4==v&�c �������Ԝ�-�J�AQ*��&D�> -z1���^�d(4.*�����7�����/Y��d*\	�~?�Աj �WS���q����(�������(�WC�嗐4�#��7��2q_�ia��Y��{�s͏����}ev��'YE����L�	 M'�>����\3�.ls0�v	;>K�?�+�2�N0�ȏ<
U9m��̳hD��^C9e�۪x�A+B<pH��dJ����1��@rEkq�%8���u���+��MA��bf �Q�f���C/@R���chB��R�!�al� �#z/����'�g`U������ٞ������������R@�3}b��%�6���
�� �_ShR?`Z¤v������K��/ל䜶c�p1�hE����`D�7w��B	�w^=I�v��@Fj�u-J�Y��-P��&(�	2
��ۧ���Z�P��,�$���� ��D��c/5HT�d��+�'���'S_��>�}S���� �ZWm���:^�͹E�	4���k�t���!�/I	�?����������}4)�.)�ʧ,8_1!�Nd`�S���KO��h"J,�l[R!�;��@�X��v% ��Io�ɬ�_bM�"1|ǒG��Z�� K����r�Q:�0�]\Q�[D0�i��B�aAH��@:���"�$�������J4_5;H8O�M���� M��!:�M�kw
D1�{;\��K�+9��N� �q]�)����-�mZEsC�X��(k��^��H��y0Xx>=�P?������D�Lr�@L�uk-�fvv YZ}W�%�H�ug(�Ӿ�c�!ɺ� ���0�����p|�u��A�<�k������
�(�X��/1])Dw�	�H��WD
es��R�Kz�k�%Y��V%�D��u�{rN3�YJ���D![��<��&��A/_�E�h�'��@��
�_��1��͗xؽ��c�� B�6!$3��h�7�u��7[��*����8� JG�)���L Rʬ%�H�$m��	!"vx����o��v
ܜL"ĸ	J钩A�WA�;�o����	F�p�i��} ��xq��7���W�3Pu>�\�������	�U�pc�I1�Y�Y!J����҃.an{�k��� �T�h/N=f���� ��5��p<xHX�Q�UK�~�8��O���!�UV���id/$.��g�X�J@����ﻺ��V|@�&$j�����|��v�/��ˁ������;0��_��)�ւB�v�¯w�KA�P��L{N?��8� �۹�^���9a��f@�#%tJ0�6kP,91�~Z��.D:%������8 �z|X){-� �ΕX�2\��@4b@�^�?@ہ�j;G��tY�}�tL�vi�WP06d>h�j&�?Z��4u@��p�HL}����Px�V�+=)��Z1W�� ���eh&b�1dR~�-�M��'!v�XhE_�x�W���=�:w*�`�T�$8�1�Z������d�J	�-��g`�����X�� 20��B����~d	���}�큻S9frhS	L� &M��]�T0�o�qB����	]GO/_����v�~N�T}N��|h�� �'`����0��������A��?��k����Z],�f� #0�X������݀�6;�Ĥи�y���[�`=-v�PX��H���%���{�dЎ/�X�;1��W�/^^�j��4�uJ:��w�{�,���z�('����ӨbǄ_����R�����!�����o��W@R�7b�O��$���>�q�Rhc/IZ`�q�NJ�~O�e���?��+��;���=�(�� ��I*Y�����~l�S��/]��N2�̗�/(��.u��M+�Lz�֎���i+(y�h+�`�i/� 4��	�݋6�Ą�{k"����We�0��מ�6( �T��^��9��Jc�Y�i�:L�m��.z��_e�5M�]Q����� w�LY�J�A��m�u�q�Qb	�.ߏ`}�zK@�x�,���%�|_1� ��}/ #��l�t��j�b��+R���|ynR��ldM`�]50rE_7X{w��Kg^��;�J��Xp��w�%�	�ݠ��%��/ ����DSm`�zXP�6V�֏�b�%!����v���d�����@v��0��r��pb�n�s� 4�g�ݸ'l���a�j�]1T-%?\U {�Wh�O�%���[���J���q�4�����6����� ���-YW��0�"XP�V!Ջ����� Ð/�t�\Sh*
�Yz�[x���.������EN`Uh�%�;��*B�Iĉ�k����&��Bn �QB6!�)ٗZ��^�q[�+��} (}
-^� ����Ҙ�$��| �(ǐ�Q�	�`:e�(�3K��9	:)	ϷOv��(�'ħf�`/[S}4%��PX��sG7��"K~�ɷ:�Z]�V_�D��a�����l��Y ~(x�0Ā���k���(�M��`�{DcW����JjA���>[���~n6���Õ�)ؗۮ����JvLAZy�ϳ��z��J%Y� �^7���f �Xi";�0Q���F3 ����s7a�b)�-B������ht��0�� ��3��Y�D-�~'p�W=d�����@o����_��p�X\֧ vU��K{%5)]�9��n�C�2���;A �W���`�w�.�&��� ]�M� �3+S)Ҟ��bB@
&r%�LWH7��(���K��� R��C��i����L>�����%��Z�ٓk����_��p�a�>�h�e�85�A�pM�P	�� �S0��E�	
9x �`,1�y�)�!��9;�2�&R��@���8cez�N���CT.H'[SPr��S��_���g2L�����x$',X���k��"h$���D	I�0�� D�N�����~�	Y���j�Zv�H���.��S3��w�W0��w���{Ŕ��uGR�	�VPj]����9�qp:X�c >���"v��6H���_�p�e�3�`K�TB�l��E�����1�ʱ>�?�F�1��X�(�W� %�]iG@���9gQ��@�n�Y['��߇y�.�� �bFK�+M[.JW�ߐn�+��Y<@�4�L�f� ����Q�M��p���[���U�W��\;�Ơ�ZP��G�yo����hL=�XCt��.���X��."2��y{Ȍ�hPS7�K�
j�}�8��\�a����`-Zor����Ƣ�nn�L�T#,��d�*�>o��	'�����6��{��C������bm��:�r�p�����}�P�y�l��
���'U��,z�y?B����HQK"
oUzL�Rh�rA�Ţ��O�%b���dg���0/21 hl��0Hdw�7g5��ae>���UR�J_ ��N���[�Se������ *^�˨�!���A��O ��V>�/J- x�k�f��\�]��E���ek�N�B� T�m��iH�yd�	�LW�9��	u�"}���_�xO�.6\�2��P�F�k(�`��/�����[.��&;辷�V~����X�LbV	�����ֆP��eYAA��$�h%�_����윀����sy�5t��)��3�w01;@Ὠ3�@����7��(4�J
��?��C��τ���Y3,�t!-��i����ZT@ĭ]!�չ�'7��hup~�}���
�X�x�ߍ��*�3:�1t����,dg�����^)L��_
�)���iw�3A�u�+�T��N��@�{,r��(���e&��C]�E���f��.�L��,l,S{��C�N��̓KP��0�T0`&�($�'=�j}�N ��W���A�PB�Ef��U6�>ft�� y����!�-�`VI��@1��6��6&�BM8<U=�?o7]%���Ib�x>h0J�2���KZ��B�`���&xU҂��3��Q!�;�D��M�Ա�"���Q`�#Z�U�&�O�� ��{6	�~�K-�>��>����;)����:�t��w����t�������j諨DP��� �@-�T,-1�w�s���$>a���#O��*K����>��FL�-�~G~U�����0-Q��;�8����t�!-�]�^�d��ShvH\4�K��B�X�d�t-hI �smaNAR_�Mi)��O��b~��o�~�A��&�谋��řg;�Y�"���x\@`H��N���"x!��W�|�_���j)��,*]���',�1�
�H�h*/{K+�a���gk~�Aha3({��4B)�#ئ�c,K3�|m��u?N�1�V�i`) ��
@)��/��Q�T[y�G[��H�4�K�&�j��,��:y�鄲�g�H[�x���a�9��X 
�0U-ͩ$�%+�Mk|:x�4��M�Nt_`��aT� �e�"/?0� '^��X{�ݏ)1�! N�N3�M�E�[�0 v���b4n�1n/�lXٗ=0����Z+�x�*!?�R���q3�y��l�ű��r2�ݰ��G"���b�����
���( �P�r���k|h����P�[����n9��P�@X�)A��,^�6���������9<�M�O����z�ʈ�Y0灞(����?�&w2ӯ���ğ+�i��9
?��U�Q0�/�8Z��;�nY �E��������	���EeIT�1q�$RƤ)����s:��������7����,p}�� ��w�Q��gS��B���u�R��1O͸���� .�2�2@Fh��X��Kٮ�8`k�Q!O���_�h�	��/�*�J-_?��N@��Z(�w��
�!��<:�+�=e��M*����_J��4	(�O2��	����f��B�㞲� �-0�$hx AY�V�K}��Q�i [)�Y!�<5*�a������H�K��91
�Ҫ��SK��ӿ�
;wOJ�h7�?@^]�Z� ɳa�P��&ԋ� )�>�2�
;������>���o���g�'w�m}�+�5�Z�������I|� Ӹ�J�N�.~`�&D$T�g��D�J�ӂ��j�}�S�=�@�0��5��$�Y �36i�[��]:+whtڃ3����!���N 
3��>=������- ���1��	8m��x�y�kY�j,�98 �зp(�����B���������bUHC��>S���,c �{��u�_�O��Y0yD<�,�j8[ .��6����fZ��Ő(����K���K�MV亚�V[�%n��)���~=�s�7r�[@�1ەq.���{b#��J?ca��� ��o?�,!��DX�s9��~4d��[4�
5�b)t�1\��&�AU "�,�a%�}��ÉAT�r�4����Rn;`�h!$�*gT��S�(p�����O7L�@o\�aI�ݽ߅�!��� i60!��-�ߙW{pa��O�-�e�=z��	�Y�
��h�8�N?������	qz��Pۄ*�����lz&}�&�<����K�Zm[\���6�S��=hT:�H �9qG���S3�^��y���X��%?U[�ܐ Q
']�o� �Fbh�����'/�uG��2�������	��jH~���B�Z[�K������_O�w��`�g Йa�h�/������<U���_�M��0`m����{h�~���h7o-֦����8�;8X(J��nGV|�Z���]��3[/�y+1L�J�K�D��;����ݩ�	z�0�h�T#Z��z%�R�@�|�`��p�[o�����d�/)\
�=��h�}>Y���	�����@��f"57� �xMLH�nU�"�@�\3!YgD�f��0�}⁵���ac��������S����@r5�d -6n1��Y�`hY-1X�\�ĨN ;J-Y�Q�~*��|s�Z�!�:�:���s(�����]T�U�9H&D�O����R� ���� ��E��тͥ�_ѻP2��Y��hG-.�pRh��.�=�,�����dˮ�
���2�ئ��xL��|uM5�}^4�a�"���0��~�j�(�`M�f*�J��z�p26'�r��\�n
E��I�#[��r�*�"ZW�-b7:K��[Vz��])����J^���|���R�cI�h�Jp���.!aM�$�n�� �/� �1 �5i�H!�'�S�G��n�0��XU�R��A>�6�k���h�>�'���r*X�gk��7���A�H�K'/e�k�[Z�#U��#C�W9����`��E���u��$�����/��;,��-y��j �4C^aغ�UVJO��ȵ����_�k��-hb�z_�J`+��o ��O23?X�kqRf����G���/��	�_�"�W�U��r��~�\#����y7|¾2z]�<a�`�k�	�D滣<ɓU��u�<���	C���]-��в)Ɠ��B�F�\��)�]����L-n�[�^��-�����H�j����?�z^ā�_eYR(�A��Wq?���@�_���'2�H��m=t��hHQ�c�UW腐��=� 2Zv��Y��e.��]�~TJ �F�1|�2�؀YN� Q����_��v���e��?�A�����:tQ ��.-�k4%�$�b�{��P	0��S�]n1/��+�P�w ���4D������{���Í�p�5#�H��P��&�F�Ab�C��o�>�V8	\F��z�(������hZ{�GXC�x:���\_?��v j^��W:�#��ȯOx&�nf/߈$
/��Z�0-�m��>p��T��<�����Q�Ӗ��೺TQ�S���s�v�k�>x���+��t5�1������>5��d~���./�?�g�Jt��i�p��<X�#)9��/��4�BA8/1п��)�@��V�<(����^��e�[��8��)�/�E&���{*�5h*?`� �OU�M�I�w�\�^k�yi_� �h	�}%`���f�}��4!�Mc6�����L�K����;�-�PJ�6N0��XA�Qi�&��gr=�Ґ$>���ּ��L߂p���sSAQ�#��X��� ~�x'G���-ݖ'1�䆊b:ֽ��Fu�-�1h<�D�0�������9��THQ��\�R��A���i=�|R��	��FN��	�.��U0$W��O1�Aa��@ �����1��4��K~	^��^?�)�X��3Q%bKW���%\�/��.ȿhn0$�BE�!�S���@�߄=��<<ԩ�	�q�R_ ���\J!�|ː<�M)��p��E���	hxHwI� ����A`����;�H�Oe�w� W��L�!��{�PQs��K,T�Š}EKod����Ϲ�+�^�veg�$��xv\�Ȣ�W�/�W�ѐ�W�ۀ/��G�˔����k�_�L1~WrAD���.��Rϰ5{� %- �:E�3�Scꢷ��ڝ��WB�܉�~�iT-0J� &�
.��~;C/Ի�2��PL�K)�� �W�\����cy�/6ҭ��`8�hJ�@on����u �t!��>���P�����+��q	�4%u�J�V��]�Y��O�CAC����D���<�S���w�p%�Y�ph����J3�(��%:ń�ӯ)}�鴔���8������wlk����h�.�KH��˹��B�W x@5�n��o,�G��^�ʴ�)����d�n'�yG�I������d�~,<�~t�+�8qZ�(֌��?WD}�� KZ�VKxe�T	hKYKj��v������������ߡN?=¨l!���d�Ek�!�)��.JG2����	��}	�Q���V�R��m�:��=�_�~h;&I8ܬWy�z��H=�>�٘�_��B�i-M�r	a�C���YA���!��[fh01�O�Dۈ^b�[Ǌ��w��6P�&S�Z�knW<@�fR��; �>����0��Sܚ����Gye�@���T�r�H���u�MXPZ�Y�@hG@FL]��U��΀"� �L7!����~�\�nb3wAx���x�����Y�-)���@���/'�}N��|�%���ȫ�=��0"@<}L�hu!�隣��	��:�@�y&�-��}��Z�E���ϒ����?t��JM�2<��5:%l��x�=��'"Q]����/pG-/�[�|W��d�_h��J�,EP�u�з�GC�K �r5�.N/�x�M��ĢH�kx�-HF���|uS�?(�N��cN�a�F
zL5P9�:��_[x,��Smz~H��i�`*8�kK��^�м�/��c-��Rb�vXh�ItL�C�,��K�=@:i+	X��B�U¼���`{W�5��C����+�����?,=���W �_����輵L1�(��rΝ�؀ލOV��pǡX+����)��Q�d?;Y��y�
[U��]h�LL�D�J��� �*��	k�K�!�P	>����]�cd_�t�-(^N�X1��2���R{���˄�!LP� R��	wji]�*�-�!L	_-M���z�!8x��Xx�@��M�-�^JIG�hk� �Êr*ƒ�����y1k�h.�O�⛜�=u�m�ָQ-��f1�#1���^�5&��`
�U��,UvPZ���)����pk�㽬�g?YHOB����?��^�$�2:w_i�/ZpڞUQ����\#� �-���LK�������aҾA��=���񍉹� �`�&_��xB����W�2�(2��8,����(���R���"���;G�_��)���G���N����Ѹ!bSH���p2�[�V����޲'#���OΔF�����O��8�Z"��&2f������6l3��1��O�8�AY�Q��.Ȃ�8JC5��Ъ�T��b�[R���V��W
)ȿ���8�F5�H�7�[;�\��|��%��v���Xi[����~@5#{�I�n}� =;�j�,>Ph	-� ��_cNu����w�Ji�>US@��fK�\�hd��y=�Q��L��f'Ɗ��ĂG�61@)��#e��9�_����!��y��v�i�d����XT���--<Sw��[Y0Ȱ{�{��E�R�6��~���|�k`bao	B�~�VX웭��I�ԭ0��sv�arX5�42B�xbqv$?0wJPWh��}k�� ' ^��Y��M�K����T<�LjHc	�R#�����YXa�О=�_��a>1�{�G��&���#�?9Z���L3�Pf�ko1т_�(�� Z��:�Y�,�9!�m^x@��Ki\_`��o���Հ�����xD�.���	���[��e��o�G��3+�)��\�thor�Q���X& �X��q���P�p4��
?1�$ |d�c)շ^%�\�$�i�Q1�M�C�'��wv���ۑ\QU_��Ӻ�D��j�8WQ|�����>B��j���KLb*Wc ��X-�@!�W+�~��4B�z�p_�x�kAumn���bS�m��-ՖnkRulniF7w�&�+�IՆn#[�?h�n�-g��J��9�~���Z`��=(5���Yh_��U��4���� �;,,�U���k� ��_G�-Z,������7���/��Dr��e���
��p�_bW`ƷT��9'�Z�����+FT�c`�*P��k��Xv�(� [;�R�+հ���zȗ�%��H,�<��O�#���Kn�o�����$ꂺ�U�K���(�1�1�{SA��s;�:4�X��`�����R�v�b)�Pgw���o.4(C��'/)��\�m��	=�"��'c<>�	@?����W��n�����n�q0 e�q�m)��V��� �4��qO���<g[�ʀ����k �Z��C6�S�$!>�^3�X|L�����e�03�{����'՘��Q0�KB-�������o]��)�p	!� PZ��Q���Vb�sw�7Z�M�a.�{�)�x��键A<��`6��4���6�uܵ���y�"h�(�	�. '��?�`��o�J0�/��-��
fR%�|����� Wl���$�dD��[� �Fnj�i8����]�c<1�&�GCg�7Hj�����:�D,�/�@E� b�GJ9)J��N�	�o3���`�!�]�̍V�+��@��T��Q��)�Z:��x�iݩ�u����Q� 7-�2d�� ��.*V��`&�͸q��M��l& G
� �P9`��pw�6 )Ƃb4��vW�~Թ�3�K��m�;^K�Ҝix���%�Aߌ`�]%��f�,�<���$��ō�t�2 9�N�E聖��kv���7�����ጂLFQ�ey˨-�)�iT�h�X����,8p�&?>�kw7W��4�_F�U��-̵�I�_�X@� Nw��"v.3!B	���Ň���*~�-��"�ikڏ��;	|jw�)��QS�{�����G��Zu{0���D��� b1ź�=36���a  h�W()X -�q�H5o$�O*Gf���!�����	��	�������1 "��@�5��er����ω�����b?w�']�?���B</D2Z�=6J�T�x�x��R1�|9��U�}�!$�	��<��J�?7��Er%A%�
�qt�� �3J��·���]���{0u�uc���[d��9 �-�/��en���,���U�>�C�
���\�N��P���S���g��5�8)�]3@�
2�J<��Ap���j�hh�Jo1���A�^	d��[��Μ�!нT�-z�!)�A[�2�S��d����Z4&{v ��;�UP=z�a*T#\��rŽ�$�K���| ZUL�'�_ ٺ�dM^.�ܹ�QE�ј�7�xq^���  UC|1x��9k�.gD%�r�[���='}�}���S�9�~�8��a�[>�#�L��o;4�Z��MN9%ς1�h�~Dp��rm�}�PWLx�S:E��		(�x%MwřFU���w��nZ���^�-a��*���T�K;��A��l�	@$�1V)K���_"Z��,���D��=�-�@��#|D�mxL�}��h%�GOD�9��PU�	fo�a@���(�4���"]vS@5։��emC-�J,m�閰ֽ	Ve��`�.�Z�4n ��|��pVpI�	Uә�u�	4�1��0�/=LK�b8���ٝQx���� �R���Z�uB���)��:�˄��*������J0�r��Xe� �
`��?$�U=�6�(a]�H��XNQ��7G�Sp	���\1y�B�!��G�e�	H�UR��yǥ��i�$�C0>9~��-�d~e�#-$0��Q��>��N��T�d�5�[)йA!��C���a+��zͱz���;S-X"*����f)�v�%\���i���Th��x�B�����T�g��l%scT�9׸B'���/.nPJEW�F,�ԿhBHJ1�	$�[�\�D���T&cX�G"�op��CL7Y_���VG
鷶��E	�C �K¹�Y�cV��l��Q`51��z�P7��;�8_ը�LF�1�H��j� ��;�	F��QY�ߖ��9<g �^�NB� �5�{1\�M4�?�>�m^�2J�X����0���*��4����%�4~Z�^o{����u�̅�����Ke���ݒ��X�Z����bA�d�PZ���h��z�BDd'1�wR�����y%i��)ah{VU�E�.����$HR���PX��(�\5@!���=�d�,fՉx:��	� �S5C�ݫm��h
hŃ�e^����r_m�'��C
�9�)�����}�S��z�,�(����a �����^S<�R���J9�.�x�dyq	Re�\ �~|hQ�G<��9�з��0#�h�X(�u����Q[��n�$x���RU�)�!��a�+�(:)'�]������)-QO:���ˆ�C�p���~��pUh�(L8X�MO�(봇6c���:1P(��K���3_uo�,�}x%�X�"V��s}[��L��$&�[c�4�T���Q�
^$�pRa۫*�!�"��h���^�	h�#^bX��	`u�J42�Ұfh)��Uf�&��-�ƶսr�N�����[��0>P����]������`������n%�����<@�t#��A�=��b���_ܒX��kC]�B�]t�^k(h	G`@)�b!͉�ӡB��g����G	1*	+D��@�'� �K_�����'O�����"<6���D0�fX�ˀ�h��/(��; vWl��0�H� oJ~w�c���H&�k ���4���̠��hOeZ)�p�`��jgJ�]��P!�O^�A⃠��)�h%W:�,�Nf-M�X� � ´�(����Đf��{9��� ?y
�j:�'u�� SQ�1���Tw��	u'�gw��B�Lq�Z�o��;���6��Z��l��A�GX{}�q8���1�!����7)���W�4�:1�^L1%s�`T\��;L(��}?@�0:/<����f�%@�Q�������������3��K��B��U�$��b�l,���0�����������[��V��c��A��� �[hNqGZ9��E�-U�h$�<)�	�!��j%�EJ�Av.����ؔva)
[X-*D�������XTdP�B%p�WM=�굁w� �_��� ��2gN)�]��h�$!4��xc�������ɼ m(8�Y8������y��
;�x	��K�����ç��pOwS�����8�=�\E���ų����R����uq�z�z�ް����;��K��f[���X)-��pp$���@e����q�7鍝o��l6��_��}�����lE#0�5�f�˺'��r�	��N���ܽ�`B}�W� 8��� IA��B�����¦0)`��-'A}Z0�P^h�6�	_�?�q�ۉ�X(�0�u �4�0�6b��wV'@�{/�3�+�9�r�B����h�sTcu�p�`t���:-��($�w�	�,���!�T�	�����u�}�v�v���A"�*�B�k�X�3_��m&0�>	s��?��XPJZ̸-�^��0�8=v�(����0ESU v.	�4�ws��^Z�qs�����R��:$U���a[��,�����7����I�^h8�jR�7`�.5>�'�~,U�0�x1'F��`R5��y� �u Kl����}wZ��Ӓ��~r��$��q�)�+���;E���ǚ �h�d[�Wp����˾��YK'�L�ܪ���̔H���BN�%K;C��Q��jE4�+��^8��۹>�H�-jq�|-hS�P�Ӿ�;8����θ��x�{8mup���y�F��0��PA����X�I 	��E%v�P�ZL�	^�UYx�g��*�D�v���@��L>�Y�3���[W�]�0��qN��o�5	׀ϝ�H	��U��r���N�z���@�)L��A���fv#_@�`]��ph���Wb(�`Ut�u�[�GH�8o|x�*r�$5�X9P1��:�0���b~%v1�P�%Ph"�:�I6Ȇ�C0�Md��/�������y׀1��}G�S���y�i쫤�:�W��fh|�t�R�!�����CB���	Pq- �~��h����MC
#�DR%��T�����,^�MT�/��+_��X���Zv���p~d���w_�`]%�Em��k�`���&�RV �����	�{i8�z��D�Lw~U���7K�	�i1;؝L��_x�eB��\��Ji�Y>��*4+\�/�ל��XVO���a8;,�U��؁g����an�;�o��H�U��f)�b���f��h︞�Ҁ9MJ�����`HBA�%�5@��M���lL톮�/�J�!O����8��H��)�.1��ȴxLl�LD@ʹgTGE��Y1ٟ��=.;�����T�< �
�*��$S�4���0;\����$u8`hTПZ��_�}U��������O�	��j�}����PX���`EU׀��Wg�*�7"�ACY -���g.j��\���Xh�'�	��S8�(�[Ѧ��>���j0n�JZ/�q���j�e;-G�PJ[9�K����Q����M�;_<��Q|���.x�7j5'��/M�:��O ��
�y��	�=���h�:�1F����ɿ��!{�=+�!��K⿊�;�J�̿h�U�X��`�z�*#���ٸ �1Zک��Q��7��7����+�a��;0S��do5� �-��H@Q�r�^d��	op�u"��Wh��k!���i@��"������@}�X4/����˶�p�h������c�xw�\j�   �/:4�l��k6F'�Ny��������%���rYI�َ��Eq�-�N��pB�58')�\� �;�0V��%����p�u~��r��'�+A�]+P�0����F�z-����\�ʼ�^�щwͶ;���,5�/�1h�M�h���@H�2� ��<�R��uӌ �8H8�a�R���u:�UCX� ,iQ�Ѐ�����n���y`�0��zw��?�P�%D1W|�t:2~J(!���0�*f�S�Y���)���<l$�`��T��3Y[�� 6['�0j@�Z�[���f��= �N�z�覰��F~_�G�K����VT�:��4�[�!{XN������UzN�`���~A��d;���	BM�<Y��t:�e!�^�VC��WHB �w@A��I�W|l�B�$X@a��*�h&�)�`��W� x��Xm�s�`��
�Z`EN��S�$!�Y3��|_��E*-�dΰ�T�:�pb�k��	���U2It[�1��O����|�������)��R��_E3B�qЙ%T[���q�Q�t�h%BW�b�`A�@���V0_�D���ߒx��N��ҪⰀ�Fz�5�������p�H� ,ta5T��ݎ2�?�u6-Btx���X]���@k�V`.�H5���@��jJ�p��G�ES0-()�ԥ]��i���1c��0a!�		��=��.GX?]B�W��U���s���R<�2  %��;��h�	B�}�1�8��ma��� �s;-T�taQ�*�zV ��5t&)�^�͘,�b`&�Z%���W������ �;/�~��X3=&���rC	�����?��>h�7�x��#6�-Y\��02�U�[Z1���$h����X ?vB[W����܆@�Q�A�(S���1��I�B�7b�!d���,�� 1Ӻ�HVOQ��xq.e@��D�NR�̲`��O��0���Ҍ��yx/2X"mY�1��4|b�rn�Wѹ\�:��+��<b��xa��g�K(��ĄQS�p���մ��^����P��2�Z��,RVD^l)5��jZ�,(�	T�tur+�H��1�)��u�u/BO���L���+�wHWW�0'4,)��e	��/�Ba-=�D%~��[p@�x��m ��Y���p2jo8����鲨�P��(�Bƫ�T�v� ���E0�5;:U��>�0�C+P9O�(v�	�f�����r0�ZFI3���**"�F�1�"um�a�(�wD�-�U��%W����z@`�P['_Ef��-?. [a_��f:#�2
wvd�(�����cn�S�ܨ�`����=�v�ח�� F'�4�)߯��S6xmH����9lY]�lKZ��T	�<_j^���9^Ѽaq`T���I^
����ؘ��l���b��w�d�����z�R��KDw3�	�5bR.�b�������HZ!�Q� �|���l�0r�i�(�����\-B}�_Y�na!�i^�$v	!��eb �9 ��9.-AY�U1��������������Z���[�ٜ��!u�J���6aT���y��e��G|ol�U	M	�"�	?L��It)A1`�9Y�\n���  ��!���_��A�5x�y;K�*<U�lAdw4R���y�7��n��a0s���>W6�g��+N��@��(\ތVxZ�t�ǽЭw]�}�[�z�o����9���/|K�W:����4>��EDOz�D�w�lo����Q��^_!�9��K��	T�/�~��Hy2��A+D ���|Ja=��u{^�e�qY�bA�3� 7��_m(-�?!�����ah�v9#� �h�o��R¦��d�e�AY�O�6k�C@fLK"� �l ��!�w$1�^Bn�p��=�{~�S\WL���B�P�n��l�T�˧;��ė^���I��)�}�x����"L��٘;l�h�7�uT���q��<R�o�P`�gf��mB�L�R�v��q�����
�/xB͉�I�D�-���/��1�8��ݕЌt�诊����O���e\x����X��f�ق�z����n�% z��x�KZ0g��kۉ�T��f#x���K�u䁁�r�N��9LT;P�]u�lLL@�%~��n���t���`�IE�!��Y�;GL�܉D&P���a��gX/��_ϑ�yþ�?�����YO�p��M�$��&��!��.�^�sPA�=��"��Y� zao�/����݅��MK]D.!�Q�j�W`��:�h��`��-�O�KJ�k [��'KU�N�/�E)�F2�������\��1����lgi��[��Gh��N�u�G���],DcpT�	�ӋL P�}�Z�ۂ�N��$�x�>.8[/�Lz��/��@�wx�7���J�)�)	(��f�R�I����݂���1����zPM�vw�=Dy0�L�Y=�ĝ(�L�,[Q�}8V�����p�CW� ��V�?M�����j�)�뷼���tYb�F�Ol�:�JꎁJ$h���J	�p�w��f;�d Y����HEd�9� �eL;��cPl�w'_� 1�K�\	A�cY_X�-j�����z�5��J*R_X�r9_�qhDꮳL��R�^%*�zh�W��/s:h�Iwsv�ȃRY�^������H����j�W�T�Ut�p�rB�K-`��N��{������'�J��A6>b-2o� �8��iI���6�(���f�� ~�i��j}�zև���?��@�)�P�1�'o"�v���8δ�	Ê4=��t/�%��ͬ��e����F�>�\U^�Da`5�Mqx.«�+�l(4�dz��|��z��(CW����߲�J�AAB1O	�7��QLl�#�����'��#����2�g7''`���ZހT��^�-=��r/\k^W!��D� ���y<��>�TkԒ���./�UTD�W�|�ƕ��C�q9�~�q-(�v�t�����0�Jj���I*�EYHыJ��v
���(�o�ŝ�Qaa�c��H�BE'��A�G�FHh�[6����(U^����������^W�F
�_Q�Mf^.W��C`z(�̔5I��V%�n���<����o 0��WG; ��P�S����� '0C����/1� � ��@��\�G��g��X���N���DQ�(P�#���0������T���V��i�~^`�7uz����AK:r��T�	�֏:py�!�Qg�>��5(-�['Fvp��pO=�"�6G`�gln<��R)� �X��h�k����K}�.��06�Z�����p�Fh��!����`�H�<nW)�q�xh�^.�S��q��YSD�[����	�m��XS�� ?��eT�~�H��'L�>�a^�҆-_j���	e���Z�����"�!ͪ VY�g�.@��K']~���Z
�\�
B���Y1Z:�MYh�5� 2��!�S�3Knu)���_�1���^���:(�� :ک���Rh�#pX�5���� n*.�P�N3*X�&�+'֞kVCbjm���t/��^��蘽Z-Vi�!0�)�c h�<N��w���P?����(�*q� ���b;L�0���v�K\a�j��h%�)�ׄR�����`��~��:�9 �P ��O[@�L�Z�z'4 �J_.1�	 �R��)��ם\<��Y�{�S���~�N��2�%��l6^�a'���\@���S[�^Œ��y�P�Y���t����閹�z����!O(S�eg��x-���h�)�(����;�.���0��^�:� �c�@H-�D,+F: t��1��a���Icf%�\>B:�m(i?���>4��j�O)�W�p������8.]�
��&^'+�4	]~W h�L�"a%"�^]	J�G?YHnX	3t�s'�����m���%.,�U�ZŎ'07Ө ��VS^5�L�O)�.�(�j��*�:wua`�F������6D�X=�L?4�|�{	H�I?��Q��%�<u���c�t����[���wNZ�S�Ni$	��A�-�"��QP�4UE��XH�n�c�ۧ����݋_E���,����5�6�LQ���/�����X�'�P�X?�H	�� �0&��[:�C	��	�> �jEK���F kNR�m!s1 ��ތ���K�>%��t� 9e)�$�S;L5�z��h%/=|ʂ����&#��/J^]٨�[�rU)��V�!�o���G�W�ܞ�BU�cSQt��A��{�	�P���'�0B��=Z�[��]PHhJV/Gؙ_}�/ww�(���{�,�c�������]n���.+�*
 ���(<qv�h �� ְ�Z6�9^*bK����Z��cPߝY�e3)P��o�k��U�>׆���-
��[;bv����EO��8W*��i6Wo����1�;�����&�/�	-~}ǋ	������ۉ��c]2�]X\^A����#.=Sn��e��.�2J����T'J���1Yn��J�4��*�z�I�Mh|F��Q5b���Y�DM�.�\�D�<0�lL��)�6���y���z�����ݐJ<P/��vb%e� �� ��(���\[�1�1
����fz	P�������?yJ3�cik9�XQ-���&�f�1=�_��B8dWh%�Q�coMe�As�@�hwT~��}��I7#��2\4��9S��V�V?	'|�ಖ�Y1W���o�c/��T5�PbZ��݉��4�2��fQ�J,��@���۹J���}�����?��h+����`�9�	�O^>�
����^W�Q^U�_%�Q��M� .�Y�)�Q-<� =31Ph�Py�k(�� 5Zf�{�1�@�9t~�X�VB/gr��@��/�F��\�et���O���_��%,&ݏ��GM��[��L�P�dC~�2��Ns%I���B8�m�_a�J#$���*���$�i�w��p�.��3c��r�����`	�T�B��QT�_��A���<��O `RV����^���Џ�r�-� �;2O���w�l�O�-끶��$(�t��� ���,�(H��6�����3��4���Y[ Q�\)�O���M��L}�J��xP-�X��0E�
�`׊��	f?Lpha�.�l h��Lm@��*X,����N������f�s�U�K�)_ �A��������C���Ź�����x���!ijV�+�$U8�,׸�h��s���,�9�!�X�L�6��	^;
U k#I@� �O)Ὦ&!~�I<8���~d�I(�� $�1)ŕp� S��6�"�ӽv�Y��08�5W�|��u��Rt�l�r��Z���Vh/a�X��9�[A��11W!;��Xhz\��V����C���x�p�"O���!:�=N'�Zض/!�0	ې)N�.�O	-�ah�ܩ�Ђ�[K����V!��R�X>�8p�Z4J����`Tl�ڷQ�8 �Ea6��Z�^����y~u��}�LR20��Y�=�Zhʨ�;~&�t[�����Y���:(���,b0T0C�l�Yk^���Q���c�LQ]�*~�[��[���Ld;�f�����=$�ӟ%qL��4<u(�Xh F�)f�	 ��A�'���3�����Ǟ�.�1�੊8'�K���Ѕ�ec��PQ��]�BhJ�볒����^�	��yp��m�1�0f \#�-�7M:1�	�D^�&!J5 �T	�n� ���&�/���^p�h�pIP��w<'^���p�$`��Q� yg�$B�¾��R�(�9�����M[�*�%N@�����TZ�]�?���T9Z�1,����3���J ���߫���D�.�qȜ��x�6Yh�1%X��A/���<B@ ��e	@�%�	��n�	�pSJW�:.�0��U2��7</z6Ų�U��/�c~�����`��>�V�Ty��Tp,�L?U��IR>�AG��r{z ��<O�w/��b,�C��VT/げ���'� 5
���r���7�|1`��<� �ƽkA�c�Z��P�0t���io�ŝu KH� Q�_J���&���(�x��66i*��R�`2B��`�:dX�U��� )�-�5_����0^�,l�*�O��=�>�6ل�r�ĥ���h:�����9Fs�)�^��P
2�Bh'gZ�2�U}QLM�\ f[(�Ph�lg_���Y�u��ʆՉ�<�+�e�#|�hS�����D��sؔ���Ӂ���e�y`�!}�%���Hfn��W �-c�)�7�v~��;4�
��;/��`!�XR�S�Z ���0��O������]Vq�t�������O��S�W���M���� �i�ʍ=�����]b)��ĉf}�����D�Ab�O�K�_���A�w?B/��7�_�^��X�Z�@�!�h�6���T�E�_��p+(.2�γ�װ��	������~��Z�|���uK��RJ��<h/'�W�oP���z�(�`ʍ�`;8��	g/�n���8n��G���xX��Jt(
ZN�&~�Qh�	t: X@-/;> o=R�)�^*�k��H@#�
1�u�}�U��*��V��Ӟ�,�S(k$'C�)_{�X�h!U	]e\������U�f�B	\�D����Q�J Z1j�_�^ Ou]IU��*�7袉�h�0
(�j�	?`Cr�@��Y��H�� ���=��	�W� !"c�P��r��⡾_��@�}u�n^�ðȲJc����0���4r������Ʌ&��b,$
*Q^��n����<�;�bj8aix^�u������k�0qc��<��V�k|U��٢�\�;tX-�_���kZx|h�3N��[!���P��)����yK+��M�o�Xh0�W��=w�́CcNĺ �1O#`9������g��*�,N~ժ��/�@P��)�E��ϕN���'�T ������,4��P��w$|X%�z�9(s����2 ��Uo�.kL'@]�P��W�DT�@m�ClR3��� ��SsE��`�l�Z.$�� _���������ִ܀�s=�	<�7�6%pp��(w ���{u[�d7��Q��I�#@�2-1��L"r����T��f�\��i ��YV)=�1W��k�R_��,:``)^;;4�<�n`R �7+�l01S�I��>-PW��!��( s�z�	(v���P�]��I��� ��-�8zЧ�>i�B��J��-	qf��Y��E�H�n0��S�q9VȔ���.���G_ J�1�(���jn?��t�w��P �i�J��C��͉U]�I���>��\��w
�D� �9;�)�%1��d~�B
%�p�wP)�z�h���> (fx��ؙ���Q-�@r���x�s���EH��]�CJ�H�.M�6>0��2�I�Nz��*�ثb Z1K��J�"^�F�5��x���ktW��\jX����H)\G=]@�W�. 	`-�w�(�v�Z$�1u�?����� �Yw����@k1c�3?�����q����� ��\�lbm�	u6}�L� ��Y���Xq��)����X!�ťErP�SC��^l��f[�S���_���~���L>]X�ql�_�V	\�;rL�B'M�3K�@,n������Lq9��^����LOKrEB�u@!�Z���ʢ����(���j�!¬�BIH��Z��Ӯ���`o�1. Z!7X��C�Y	
�t)�9@&�|u2�_(�&E�N闓��0��G�-]0�h��wȆ�,n� �q�L��Q~�*�;�	�G�n�_E��HݰV8���������#�g�xO�7�?'�T�a��.���2���=>�n�k��!���*��aw� �[��{�7�u�泈���OYIٳP����Á���0i��� �MN��D�	k����[6�<��j/���N>[�����-k��jq�+_1�R⋩�uah=7>����:;ZU�4J�N�#��O���rΘ�PS����E0[�T�K�bO��7�F0�Ï��T}�b]��S�T���TRA�V{ �?t���Azz�{�횣�k$�%�B�vJ���=�	�t�2W�{�(�&��Yݜp�����b��@]hUv#x���}��Zt�0��?	b[�,�F�Y1�,�/I",�����В����")�W~���z_��f�����x���
~�4�G��͋��0�?�V`�%�8��B��>|�O��i��a�*�� P��q4-�w���}��fx�p4������R�������y����:��B͗|7)5X��U�B1XE�Yc����8����� �)%nkzt�;�fpV�%��6Bh,�#eq����3���ۏzo��"	�:J��pG���%�JZ�Yȶ��P,64��ο�LZ��m�4���QPYX��U: ���6�ɴ��0T���m�h��N[�1��vF ��;����N(]Qoq�?��o�(��(�O��|��/�Y��C�����d��X��� �zf\^WU h�x`:[����f����hg� �+�#�PŌ k'M�_P���0�#F�4��L�.h.k�l%��xY�f���
�<� (�R�Ҁ�l�Χ�#����2�'Z^�����[H�vx?9 -B�NI}�M�iђ���J��/[�1䪳t���~��1_���㔇�X��İ ���F�I��\ Ud�@�:�Z ��J�q��	�.`|9CŲPfɆ����c���hp�E�E��`N�����jI�gC�ݟ���>�	���	�n-,�U"(/)'b��adh�is@ ��a�8��9��v}��o���hIDu4�����eh:;Q�dD1L����F�݂	�`w�R?���7LSo7�m�IZ�{K�,�m���RrH-�@k��a�s	�@��V���CbS~�>���@�;�E�^-��/3��J�1Z`a����^������!�1�!��h�=aN�P'O�)x�트�Cʂ�,�0sy��0C�M"�l%G��x���Z�f4����g�a�TX��}|%��������`0|q�\na����i���N3g�|h�bu����K`���P�%�S^�и>J���U���k�:-� ��C%��~nvmz�-��� �G����N/�}�E�@ֻ�9vX�-X:���|0DT^ �)�h%����Yׁ\h�;k�ÚEO8�9r����������(�)�뒘h�R�J[�V�DI���~	��^����E�)ɠ�� ib,y1 �]58(�	!H�E`��u2��u��H��Q�BPw�r�#�G���K��$��(�2�_W�@`�l[���H�lN�*�Y�����W�aS�9�����~� �XQ��Ft"J�\8�('����aN�~M�~+�P�4y8��O�ؤ�e=䝭R��CU)W�e3E1u�L���(X#/�6@�1��a�����O�@@���A't_l"HQ�ѷ���ؒh$bu�rw[R(ϵ�[��8��$�L8 �EM-�Z����p#���o�G��S)��P7�g�&�_w`������Փ��Ȇ~@���& �ރ�V�v��௉���:�D=+���H x:��i �k��qN'�h�؀�J��oN��y@�D}NU�%@_���?D�ZI8^�b���>��1͔r���m+$UA��x\VĪ�	�hE�����%u��Ѣ�r�9�g����o"�(c�D���R�kn�Vh{��F?'y$L�-E�M� �����A�O"��A���ߛ-S��y��>�OƩI!���\iv$mL%m�&� @(��n1�����-Z�qQ�Lܸ�X^�x6�X,faFpX�U]?�R�S�R�U��V�`��r�i��;�O��Pj�M��	�'QG���5_3�AZM�[�H���	�/q�R�j9?4~ftA�;b)��)��g���<�%�*�! �鷍�ya���c�I�Z�-h/�vq������ ��<'�KP���iq>�+��N�yjow�ܞXr"% v�'��M@�9^��Nvx&�,/��?�C@��*̝ؾ1� �'[>�N!�����I�0�zg�X+���)FTiT��B� !Q�.yq�`nA@Ea� }Q�����c���˖��%�yc�����P=�	��[���܉�b�_S��Z�*p^�h	h�%��q:<��a��KB- �:����C��Y��	 �#��|���BgWd�Y��ecN)�@�(�^� G&gt1�)ڽJT�\]az�&Ԃ��B'�P�/.U⒀WO� ����:J~}h�WMS��TXoR2�bgA������F�O��	��J
W�Z���#f6+(yE�'�_D�(A-ט���+�]�.�.j�����!�c��hZ��$R9���Z���0 Y�[-��y:���2��w�S�2�`Z(�,����Oȟ[��v����Y���*��������\��y~	T�%d���+�I1��
 �%md��: f�c9��u��
�Ž�"��u Z1ع�}!Jx���%4y��n!O��	�C�#��m�I�ʼ�`�x'�C!��d���'BՀ��1�^h�O��GZ�]X b5����n�ICP)�Y��>�Uh����R����`���0��	���:��^�D�S�#�a駋|g�u@�1ـ�@�)�X�.Xt}^�L�^c�wvF�)�1���-M:= |	����h^h�ƥk6�\=i�h�0�+&~��L޳A�|�.�����P��S�A�����SH=��KJ�4�Ka�
��N��i��㙒a���$�� �ETU��$�.���p�lx>1�2KW(w@53)X1�1�$��E�:�>h^;z�]%�gч]��9�P0���۱L& ���Ʌ-�� ډ*�=Ƕ]�
h:;�ݩ\(߁�+�0~ZQ�-�����0�4�-� ��6l���7ܮ�ՐN�#ɌH���-̀�Yc�`0�^�(����R�"��+�^�����7l���d)a���r�@�9� 5�-��Թ��X`	����̱��U��m�_A�
3>p�X}�O�-�@%\x�b73�LZdR<�V�J��G!�XO��4q%��p����}��nS~so�z1�@�Xr�bk�W.ȶ��y�	Ă�z�H�@ZP!��]�Ŭ2O(�h-�,��d��X�Ԫ�	�X�w�@����,����)@k��4�I��<�0���>���<_��'d�q��}�4��U�~�UH��T%"P]-�`h6G�r�W��@�;�ߘ
����Y8C�J
���ctA��7A�u������$ǥ��;žFM���THq� XY�C`%�c��B��J_���	��}��?ė�1����^����4W���u�M��������ׄ2P�`�u Q��m�2	�{�W8�K|��F�r���t�E�)�Y
ڗ��R��/cr�	�hImT`��V���O3G�v��_8�2&�&��|!x-\=�}�W^F��#v7�����<قJSrEU@sK���CjbΣ���-EeSl΃;X��5��0��e ��������R7�R"�Zz:�A��"������@�hL���i�W���'_�W�	�X��xۀ7G����(��;��(-X.4	W����1JV��v+Am]��0���ޖ�'S�Wf��U�Ѡ�G ��1;1�;�R`�"h�v�L��Z�i��p��3Z�r�������?Nf�ł�����-&2�`)�^�y�������~� �H� �6910�.�Wc@~�hڢ��Y
e�%���8ZK+�#�<&B����U�|��-���.u�Mw�PY�l���c�Q;N��K�`U$�o���)�����/� ɹ�S%�J va�c��`��5�w�XK�^�fAl�	���8dR��ntw��;c�2�k�y�~��g�Z��݄��v�`;�l۶���(�0�ӿ`�P�����.Y��y�0q�D�W�PK�o��݄�V�蓉�e�IZp�v�F�O�G7[~���!ՠ�3RWt���.]���
鲃��r��{���@B�W�, �JQ�r���R�x�H�)���L:�Odol�x���Bh�-�߾��%�)�^������f'@��s�{e��V�,- 5),�;�HE�2C�<��F�4���9�F�$!�;̲��q�A�\-)1Y�=�.ܮ�x�?q'V��+�8��Z��3�=�d��龩�4XQ1�/ �P@�%�0L�w1�Z��JHƖMԕ�~tW.>uU[gk����L��\z�_��a4����N�!���&�o�kN#��IUhnf^>l?�/��_���U�s��7�k��A��������[A	�[ŽB&�e��h���+��Z �~xiW�u����;�4a ��f�AH�4���EBQR�����q^]cu��@
Y����NdL��E�����c�`�Z1n� �p�]������/���3(:���S���&�1���ؗ��}�Ftr1�も������[��Z^�~��Q"s���1��^
ZRᰈ��0̸]^��������.@�q)JVٸ$b�+wԦa7@�I@ȍ=�v�����-3��:��e46$�,��(t�
iJfUm�����_�����Y��}��cx_�<Һ��kɕ+�L��8|+�����ߞ&.����c���j=n�I>L|��uWf�2�}Q��B��]ǘ�
�3 2�)�7%[�_�*ӟ�5�k�\hNTt�w����z�������� у���e/I��-�i����'��sdу��C�8��L�����t�g�'��]�o�7K��{/����(����r���� Z���>!*������)� hI�L]��u��3���n��B���Y�p�QB�	�O����N��">�K�8����2pVK��,]��|�A]���	����=�A�ȴ�1� -7N)�������O%u^�/�)a*o�g�P��˘��GP�!_�쫭����-t��'=bu����N �_)nH�����`�h�T0�+N�O-�'j1���
j_�����2]��)ѿ�Fu�CT}���5~��� �������TcV[� Y��'/��tKR����@�$�b�VWY�z}�i��������N��Bbd�ɪ{%��CN�aé�#)�e~��n|+����vQ �#����)\˫	�>�d([���V�zp�?@��%0�P$I�Nz�pZ��%ub?C7��}��	%�� �Y8I}ٻ�u��d�x��I'�[��s�U�)�L�I��m'���h�̣IkT��	I���Y��>#5f@�/*���2�J�ؤ�u��-��z�{�	>�h��1	�abeڸ	�g�{]�� Z��:�u��u�/f��0��Hw��T?'GA�bh���9��H'7�$5넍��|`�	r��I���K�4&�)�h�_������kHuB!�T�q���-�n����i1Jv�/��5MXJ��`�Z)-���g'���R��;����؜����*{oBMIr�c�Q���=�U�V,��Q�!�/�k�f*�3"h��u��U���ޝ:���T��<N�{�����?<����0;�_�N����]�Ăw��y��g���.�����J�d� �@?{�oN�i�@�1�HZ� Pqsh`J��`�������,�1�'ܓ�y��nP��	�a�~֕Şf�9��z8.Q���n]4p�K����ҿ�,Yh*Bv'Q_*�ipy	����%��1-��a��J�l��$��5"L���,!.F��X����abk�%��7NHǻ�����n)R���]��`wZ�:��a�?hS��q)�v�縷��ZRT��3s�Sሮ�,��ޏK['	�k L�go#�kowt��s-3��tK?�^׹{U���n��>���č=jhYJ��JM����R$p7d�n6�;�`uKE�E�XS�H'�d@5�Q\Gbf�6��^�?���	�]�%�-	�h�3s�Q�+}b�w�����	OĄ|���O�`
hJ	�j�V�Jq�@���Gƀ�~ń�!�_�'�_�m�`�aN�,�r�Z� �"�H�� � 1%�&<�(=���ڹ��~0�Y';y�0	���� ]}�4)�b!ӂ��|�7��f��π�R���Z���P��J������J�P�%�.�>��X�h_�$�9�P;��K���`�S@c � �J- ��:��HM/s)���Y�^��r�\�G\2�UH�`�p����4 [?/r�/򆀼�S�|��w�.��<�:`�Ac�#!� ��G����_L�yKj�&�6	)�G�O�w�Z���ɥN %�� )�"�6���;�0��WI�z���Z���<rM Ŷ9z�@�R!�u��������m����0��0��,h7_�;����$/�+ ��G�`B�ڂ ���1�	���<�U���K����i��4N�4B6��'��f�Xf�~K+<	�D(�Q�\���,^X �Z�,)�L]�5- �(	�����2ԡC���~��N�n�o���t�K�u����e��*t	hMƈ�J��^��;�zdY8_����OW�w�$�ՍQ�*�	c�^��g��<�иKޕIà2�0�#��1��F`U���Z:����)w���z.���"8()��%%����h1��M�;�9�<1��+*��W�6�~��g!�`>��8'i��}�-^/Q��UdAW�\2y)������Y�HA�W3�� %���m�������� �R��m�J�B/ |o&pO�Z���������v�(��.[��=xh�]�/����f;���P�p��.)�'`f0ӵt�o�N�p�q/�O�[s�#���( �;�H΃�|�BxU���7����;A�2{�S����:u�0,�	�~Mx��J+\Y�H`�_W����S�)���ѨZ[/��Zع�R))�5_"g��e5�P��cC�(<h&$�\Z�ZSNA�_ �$w��
xr��)��У���0��L	���%�����S�`{oR�L���0��;f"M7�����$�r����렋9@zIƹg��c S�y�*�ΕCi�2��$�6W\(���*����cDC@�Z�N3�|Nq?��]�B�)��:����z��n]��	)$y-�B5�
!hK�:�&P. P�k`�
�u=C ;��D1ƽd�X�r"�h�6z��a,r��^�m����$\� �ۺ��$QB�=�B�<���c�,yPPb Rh~�YI�����-(+�+��!Txc��d�5h��(BTXuq��``�F1J�z�	v�x��4�����)oI���LP����~#�!�^���E��J�X >F�������v������c���\�%��C[��s5,�13����X�ƕ�J,N�:G�;�Y�xM�`��v�{)�-�W��T$�i� J,L �����xD���P�'����� ��)�Li$v~P��	�ktz�si;+`��u�,�1�b3���@���wuXZO�8�_�p��� %�sc -/�Q��(\>P0Xa���-(j~V��@[�$���qz�'{������L���1��6�S,?2�\�kfQ�|��X�v����x+��b[,k��[M�H�Xd+�*�LR-��Hx���"C����<]�N� ��8�*P1��u�/K�*���_��D��1����u�����o(�X���ԵVh�T�o]�G�^�����&`v)��3t'���	��l�x��q����bH&�ثf!.BR�	 4�_ ���Ms̰|Z[�+XY]a�#�n�a%g�V��+�?�*�!i��u�h�T�&����r�N$���0&d� n�;1ݸw6%#VZ#dFf$�:Y-Z{B����G�a8%�]4M����i/'|�����N���P%� �/[�Q.�R��T*X�V��R���2�`8(�6�锬�}������@�)\�;N�:*�|��4~|���rf^Z�)W&���׀��O	�["��@�"�'%@'�DcB9 ٳMA@��ޚ�,�J�0�w�P���M+���w�c���5lK(ċ��� �$���)����d�%muB�E�o&$��w��O\�"�t�h��"	��2�ֵ) ��A�l.ʅ�Ӡ-��O0�Z��Y(�	,*�����>6�9cC��I	m��S��)/�Ϻ���o�5�	_�588D��|�./쟩�}���_Z�*SF�uY�?�� .�5X�����o���s/�	��q������Sd!�{W�/��V%�>�=��pAP2��wY�U��T@��X8=	w^���a�>�t��	�s
?c���a�\\}�{���O���/��������H�w��u���A(���1�Z� ��Mm"/�_	�w���d�ru1A�B1�� �� �Ys�T���)�-�?�ޘ+�>Hqǁ�O��;�QY]�:����{��*�.lyŗ��.o�_�U(��9Z�)�DR �q<���/a�@X,v@�/�w�f�a�@�SX�r�k��DW���9_{�F)Xnȷ�I]ZE��z�Z��<�Ëf�\�&��4������j���)�]�Q)
&+�'�u��� >�k�����h|Q�F�V����W�DW�J�c�SQ����bLY��U[��-HG�zP«vK׺ 9OK5���4�a�@���,�2�!���6�	�U���V�I��0�LB�2E�_]Ŕ� 6	+X������a�!�>@eX5�|�NÌ? c�X[V��������&�����?�� ٘r׼HS��3�u� �q�O���(��8�AJ��A�W�Z�����ih$AdʹA�1k��R�|�L 9C�d��D�:�ɍŇ ��o��6[)�5�R��l�N��@8YhuO&#P�2*~�����{����-��i�0X�5��_�cw"RH%lJ%�2����&H��X�G����j`fn�<b��8 �C�6ã �6rhf@��[�:F5MRp���h1
s�s[��]�d�B���D��Q�kS$��"$�>l�&8@,��3m��ϡ�f1{2[���^H������_�W;�V	�{x�#B�'X�sb��uX<	8�m��]��s[�6i2��.P����=�d3 _�/�	�j?1����{�1F�n~�[��2�W��y�ru"���P�R�m_�)�+	����� K��p7S�O$����؄h��|��X�dI�����3��B�S��f�A���h�8!��1��{;�b.�W�WA����4��K���WA��/Q�X8e&� S����x� ���-���[/�e������$h<���)�^ GdU@�@�,_S�r�t����$���~W�27sH��ݝ�����DQ���d�L�6�R:�,��"m^Y']�~�	Ov Wh?_=��9�2�^Ջ,���X��dfN�	^b�ի�ژhXB�*]׀�/<Y�R��� �q5o�͆�^���C�Z�G�W�nJ���T)(���VU����`!Q�}�P����A��ʂ����_b��vU�]�$�}�N(�snL�h.m3�R�1�[��Z�d��r �Y�?1:�M� +tA:�)�/���!��hRz���x��Ya�c���Ina:功���,h=�o���Ĉ- >��$M��%1��l%��
�և��	}G��E\�7t�g��}��T ���z��"�(��)�᚞ Kn%1�V?@^�;��~� �f�uJ$��� Ph�0�g����,��_�u�	"茽�n
(��E*5+C�A(�_�I��8�� �����������隲_��X>�q�;5�	@�K
�����-<M��CxrZ��lQ0BFY�%��T��,&;��T_�B}�#�ty�'���%���dT:�G�i�����~�c7_�0�48� ���!��Ow���O_����L[)'���"�������f���"�2�a�AT	%qa<��y_;�r��
}�Qy��J�(��޶��kU���L�z���y�uN #�N+�2����q����;��y&�+���{ k�m)���E��b��+ꋴ�[�셞�^L�{��%�;](�1l3ƴ�iLr;�Σ5�S��������	7]�B�Qx=J��V��`�P5Z^�
�R�)�en? cI�z��i�~A��v�N{����;�������I��	�0<��ݻ'N&nF�f@�>��@8�U��(0ti\�~��$���'�~Ӆ����AIuf(w]?JKIG[u�SG2�Y�)>`�����fSW�O�|zd�Y�q��}h�0Lэ��  �Õ���5����A������ȉʠ��1:{A�:e��N]�B�UDӭ���a��/Ce5��i"X�&'�W���2��,4>��CZv�/�`T�}:�-��(�FOk°T���~����R���yцՄhf�2�����&��	�9^�;Q���kv1O��r�F���yr�w�a�30|ROhR[�.gH<[�)h%�ـ�@�[����ӕ�s�*@Ox LP�����\R�D���P��K/��7��aQ>�qBc��1ò7�D{]p<PX�u%��1`��0ӗvEYw;N���h�Y��}JH�;�G�!h�b�>wF��ZQX�;���	�2m��YG/�~�@+o`P��p'1h��X���y�?���'(����h�F:̟��. �$S���)Ĺ���<v�q�f�-�� ��܉�)��0�c�V��D���M�'
ذO�L�Y��Nhct-]:p`%�8/�T�z�d�S��hH@P�Ԡ'�AN\����D
���1�s���1�'����N[6�'����� R�#�ӕO*-��Ds�&�MHӒ(!� f�Y���~��d5� �|�L�^�])ژLo-i��1�h�ckR���),i��.�cm4R����1�ාd����Z��O{-�2H�й�;�\K]t! �56I�u- K�b�H(k�	�C����� }���)ӗҩ�:]h�~e/�9C�;���ć�,�KX#�՗�h!~#W%X]L� Q��S�>�L(��O���a��Ҳ$Q��G/�tb��h�:������NO'=n���V����WH:3� J�8-� �G4�~K�I�y7�3kD9v.��� JKM�Ya�F�èC/���v��w��K��`%Y��w}f�pG�L;h B|�RX%k^�i=oށ�J�A-�ր�G �V�^v�?W�	>��8��h
����P�g�[-�j!b�b�]L�	t�(� 1�~d�*S��[�Q�,�J���!���W�ž	���]ES��ȃ�`����[Y���w6@�fR�r���Y�r�)@��~z*�!��h#5˓���]�a��	: f��d�L�;���"�i���-�/DI@��:����>�ؕӖ��P/[]�R�������@���VZJ�p�w��!��y��Š��/�n�N����!��X��_���f=�yO�7F�zUq5 �<Y���/UN�������E��=����
�:�<!�C��o�	��Go�	�o�A�4�IQ0�o�����m��OuWW��{a��@-(2Z�6���\<��J��b0�'�C�����I	��a�_�p�?�V��g<MY,�:ڋ�+�CS��z�.�]���V��x|�E8`]0��4�@��)�\ir"��'/����;��9^�Ws�����r��(�@ۿ���Ű&�=���ʂ��6/@�1@E�s�D�[�G��`����J�0�f(�����O���L�M�uY�1(t}�$Eq;�&����޴�Vr����z/�i	�B�^W�46V<)�r�]o�\��	�~��X�M�����%��V�G�R����h�ۊ |'[��. ��L:S�LD�I[6�d��3���.��w(R�,�������fP�;0��/�
�q1$2I�K	Us+a�jS�0>- ��(���/���M�q�53���@=kS��}��oJ��=P��H�t�)IVB��	h"`F) �j�1�鄵��]�֖Rw�ډ�ZւD6�`�G�A�qR� þ�u1�!�^����S�bn���U�We�%�x�`L�f�-�_zW�U���'JVb��о����� 3f SP�������������\n=��wz�*"P�˾U�n�~(T!I����������W�J���� D�黕&\�Έ܀�A�֥Ԁ2S��n�8�*��y�iu'p) mX-�5M
�.�Z[ �~S�=�C0z�$����E�U:�`�x ��-���1��F����-!�`�AČt{fk��A
.�<�;N���8t@�Zh/O,0��a�``�r�4�(�	[P�Re��W<�g_����X�:��5����<����`�sCXi�B�U�
w)��hE��7�i�a)o�P�V�	��	�T����yAV>+��)	��r�MWf�Ҭn!YK�P�v�D:�pb���P��wZ94	��q�	�_�W����&,MJ��j#�Lh�;�C���V�Sr�<��^��N�ͬ$��h�1�_v� �#K^-����!ù�h뀦m@bX�>74W���+Pw���/��P{�q�2+�=��K�����0�I��ֆ]���뼺N��ɯPm%Y[�	�Uf�@�ﻃ%�n4^�w[������N�� H~YH#6P?j~�������j��P<�&?e1ҩ�"��aL�w���dA�h�U����uT�Ku6'�W��4�[����΍Z�r�!�0Q�P��W=	g酶 ���: x�ۨ�)�� 	�PwG1N�p�j��L)�A�4.�{9���@��,����	����|ʼmP��i���)��_e�n :�C� �,��e[�f�fn�hrZR���90����%�DB';z�?�k:A���v��;�����X�1���J���*sK)���5�#%}׀�aq�}��l%��}g��W��_S���aф�%���K���|��1��^�� !ȽLZ�m��U9�����~�O�Q��G�`�%� ��c��{�-��:SWD3��F8�����o��������,��nҫ$��&�}I]��nX����4��9(�d�71�(�Z�AX��[(:ľ%���\��0�6�p��([�-hR*_m�/q7�"��C�	��Z<��Y��@�>�X��������*8���!�/O��3�%~r��odnO	Q�:�+W"���qkI��L9E��[�����=m��:(F�	���WY���c�	�^]�G|��zhJ^���P��N`�A�8�Ń�!�s�ҭ��k������E�ϡk`{�_����:���s!��4-�_�i�鈡�א��DZ����V�?QEݿr<
h*J*,�'�2h�*'�:j�o؀����@X�g)�D���K@��_�Ew���(G���e}o��*5[�!`�>'
�`Ζx�\��4���ى�P����
��F��8�F�3��0���f[ ����P��(8�XHH�57,�*->���$��Skڕ��#�➲eU2=U`���;�:�>�!�a��{����r�N�h��:�?D��:wSY���!ќ�2>�t�QY/�)T��d)���fCJn<�=c���t��N(�&-�6Z$�r�@�)�Wu��*�����O��>�B���Ѐ;���-K�i)��9JJ	�SA5�[=�I� ��!�-�:8K��v���>wA���]FZS�JKY�i��	����$��G	_�}��R� �O,37�t�h'e2F� `Q-?�+	��à��5�>3AI�@��$0�rwG�n*e�� E�a&���Q��^c���6�笖�0A"�>�	�̀�,e(�������1�N�@�� /t8U�e�Z��9]p^������e�!�9+�C��A���! >��򾩊j��K` Z~�1�b��9)�%��Ȋ���8��!�_�ل�#�@��P����$e0b��㸁r���	�^�\� ��Xh�	�<:��d��u��1J�3�P-kq�pX�A~}�-
|�X8�� �-�NJ}L��)���Vj���_Y�_A�+�a��5�-���$� �6�i@-9?,��� 5	}hO��u"�-�L�L(���,�-V�X�AO0��ĘH�gm�u�=�%�u�q��W�v�Q�+)��WYpX�KԲ�>0��GԒ��u	��T�����!��Ǉ`�i7^�A�'��h�Y���ɫ3�Kv�JhlE_�-�AFو�P[U'۠��ӻWx�:�p�'�8��jy����ѐ��z���G� ����1�W����p7��	iT ��K�����l�2**�'��x�K,�3�!?	{9���R�i�)F����! %h�@>�ᖲX���*4�=|+]h���m�)�}����:�i[�������'N⾎�du1�~����e�.����o�9��'_L�����N�~c��f��T�`��c %h�u�����*YZ�����we��Cv#g}�/ƍ�Ь�	�XCϚ|�-Ċ���2�1��	�ў�]R$��_���0������@�w +�b�$�� �xC�g!M�l���5`�?ۄ�h���[э��z����xz�V�k�K���������B�U�-X�-�g:$�N/��nqK�@z��%]*�1O0�~���-SG�K(��N^�.��XY|���y���+���s�ؒo�| � �Y�h�V�!����-0��D	�|]���Z���^7�X��v�e�sd-n"�G
"�:�1�?	r)X����}�Z�	b6i 2HI�1-'��R)�X�`�8�N��?�~��>2��](+0�(��)�,bQ���+��-����� ���Μ��(D��.�&BL ;�2{U���t'$~�%U ���~���.�3�Bw����eZ客�ѡ��c���g�hjJ >[�y��ŤQU�3�)�,���d+@)�3"�d������2�T� �X��5=��&�d���V��c ,ڵi�@��D�$�1)���$�Q���Y|�Dј�짜�`�~A 0�!v���AC"�ſ�[4���%J��Ɛ�>F:YC���OՇy�?��2�~��@$W?&eb"CA�\I/�=��vp٢{��]���)�IT^�����*�R��!G~��Zy:�z {�U���*S㓷�RzҊ�~[^����J)ú�c.B��Jf��<.�|"�+��	K����)�"�H&�m<��P��^��F����'7�P7&{��8��s��)��z���D('�?m_�n	�x���| ��TD���.[o�b'	��
���/r� U]$;�����}�ݽT�%��!'M�	\�f 9{�+�p+��ٸ�)���:O-��	�7��X�
��0�u�׉�����-6�] �A%(F$�la�5�DCwi���o����!����'��U���1.'�Ij�	�C�N�)S��u�L4����}4z�[�C{7f)|�47_���lG-C��H8.�H��D�]A���O9�oș`�y��@k��S�6��H�u(��;+��ï�1��0�#�5��`�?������,�'���	�MV
*L�<	ЭP�}XZ� ��b�T��6'�0�9�H)�so����[Hu�:���^)�Tڢ��8�����	�����X!ʘfO.�{[Le��)j�qz0��k-V�J�X���!5�GO�t!�M|����_ʗ�	V��rx�z�<�VL��������{"�k��wZC����!�2�ڧ12XJPQ@�q����gk	�h���WS(?�_XFzP&��A�"HW��_��'�oq�2��Z���
2�R� ����� h�^�J�K���[W��]��1	���¬b�[���Wqr3)ڴ����2����ͻ+�"	��������	���:��1�^�PD�鸙?W����f[NR`�^@�	����cH`<O ��ziO�
wkM@� ���h�d�eƨ�B^護����TQ��M��E���h�vc�_T����H~n�b.�Z���%q��ͬV���)��w��>-�^p};,Y^���K���w�8�x>��f��� ��/R]H�L��pha`���6����4`��Έ�O�"�o�WcnZS�ϋ@��hإ�Jx�o�ad�b�@X+�{AO��ҳw��Xk����n�^�d���Q�/1�H��^�̩�p:qe�]U��1��hK��y�
OÅ��	�zǃ�����5�%Gؖ�~��̹?rL���]���Ta��L�� �RY��	� �	�zZ)ˠ"М?�Z�^Ů�fQ��+� <��"% dv�@5r��bd�O�\��iH�� ��2l��	�}Lp��8f&A�}�$�(�>��7�-IѬ{�:����b�wc|M�2P�\J��'-���Y���M=�I��ӆ%�I>@�?n�Rn�>�O��	��>����]gc~�����e�����n�֪/sP6E C��C��v\�Z��{A�����Y��:�,L8�h`�u���]U�	&+]��(P5�`��'��T.�cd�-[*�n�k�MR��<y5�ׯ��-4���v	xU���*uh���^P�,r���Ȗ��fy���ֆ	�Lw`��p�O���%�#�V�iT�|��I;0�:	0Pb�EL,+K�(�P�;DR�����p���v01r�hV>GU�)z1PB7�����cth�b�Hנ�3p�}���P;+�q<�m�Ef�-A�@_d��k6����DN�&��pDB1�H�vt&�,&X�����J"_��ˣ@��n	�p~�%_�.w��P�K��(����CҚ��?3�	�Z"��DQx���?��R�>����I�5BW_��-�9��I_l����1zFl���Ձq�t�8�^y��M*���4��As� �����&���7�	!��G���[�e����UPi-�� ��o��C��.���pW��o����d���$!�\�W��tk0�Х�S ����rXP5��tMW���2�X`e��\u��Wz�(����>\��C��$h�{�Y�Z,/���fc�P,d�ȿ ����0�lj�pm�@
�y���R��$¡��3"s�P(P�?��&��OS�u��%���(�mP/W:*��Z��N�8k
@ƺP �%�Ձ�h�|(+�`�y�~�@��J(��(m��-�Q�1�0C4�@�h�0~'��}H��J������;�'������|bf{<p>�7��ew�02K�|�"�٪�8[��F�5���!@Rp�K�(��g�U갻DX�cKCg��a�G��4�uj���'������h-�a�1���8�
�J��.jm��� �ShA�}��2dQk4(��?'��q a��{��0E68CS����R&J���g��nk�`Ð��(��>�*��k�cc �t2�,	���[�s#[�b�<���_ܩp�	����k�
�c��ǂb��v_�%��,�b^f�7vb,�Z2$����SOR��2��S�Z,���8�3Q��
�5�O랫�� ٷ6����r�h�x�j؂�10s!P:�w���@�ŵ@M;,)�}DF:H�kZ���� �HW��)Kh�7̵	oה�I�|,]�a駊 �@��{�5:
��Z1(��/�h9UB]@k��/\�w�:�|�-��h0�%�~P���F%Kߺ2a/1k#���O� ���������t�
��=;�#�,K�x#�q��z �͹�G_t�I�T�O 9)o��3"�*��B�-fPS4����`�V#.5��WV��i�A��e3 �ސh*b�2�<�\���M��hPh�b_woZA�]-A!_ܥ_O!�V��Eiz��Q�H�ɑS��9/X��y8��ߘV�V��o���~6�|^p �x`+j�=����a2����lm�<&�� 9/�1�FH�`�BE�# ��h�+-�r-7i�L�E2�)�1����/�}�B��m��>�b��+%�`����S���x���b���������	@RvLkt� �	�O`qPA���-1
�k(�������Qi�L6�1f�!�� y2 �|�L�
���{���h���Z�t �J��dPn��,}�ah�F�;$��P1Ӫ̶<ӵ��g�J��)ɸ$N�2�wa�@�5�����S�N`C��CU�z�)���n�SQ;�D�-�p����>B��!����A�� ʽ?�!���h/<v��,G)9����I�8ʍR��m��!ڎ���/�9@��8�t���p(P�����<w3�u/�C���n�i%np�u��+�~� �;%x�Z.�����b�i @0v~U-��w5�n0=�=��()���u�����p*���	.��I)

)l�][Z��F��|�T��`'�<R hIlZ	���9 .�L�n`
E�S���Q읱��G����Y'	@��+0}p�?e0J����^1ј�B~*)�JQ���1��'��	@�#c%;\	�&孉�`p�xA�WK&��uO�i��)�*���;&��*W�����bx@D5�<�%�_�0�����g��;��Ao��t4����ѯ��� ���^���Z�N��Vh?m'0��x 	�L�uP{�]��Xu%��Q�fG���>D��Rد����������n�e6_f�V?�F�O�lQ��R�H�^�q��O����$J@� �k5C݃��K��w���c�� �_��O���V=�J��PM� �c���)0o܂Q�2S]��6���k� !��0��Աz,�k����z'��d����n⠟Sμ�_�x{a<j�)�u6���剉�CY�%�h�r�����hZ��2a�5�s��NU���-�����]&�r%E>V�'jh�{��d�v����8WC������
14<E��WN���'}|��+X�*�LL-�?��	Ny�ej{	�VX �:>�y6nj ۱tq;�$�5�%����e����V9-wW$���EJ�2�W@���q���n�a�?�҉���É���rYV�"2$%�Qz h0������\��@׵�����T~WY�j	0*�] �!|-n��k\0��4:��fS�1w�,"/���k�#����R�50�$�J������?{p>���)���L���O1�h�.m\�%~0�Q+���^^`��K��LsJ�B��u�
ȝY�`�a駴��`�e���)+!���	k$c��W�F���L] ����;����,����1ݎ���բ��$���{��r^��)�9�-�tpxh�Xs����ʀ6͠�fh:@&L*�>8XXD
gY��� bc�m��e
n�����2@	�%�*Hu�����$�����l��K����0� �U�Yf��]1V�R0���Y�����S'%���ph�q�w�:b�Ћ���BB�WYE�YT�-�i���3�!��z��R* 247W�� ^P%��gH-O;r2��{K�r�#��P� �0׹���Z4��_�35F���A-B�^ X]@f ��&CK�:uU�y��;�}�4%@�S�T�S��� �8��֮��Ot����U�	��ק#��0X0szc�`@d*z7隡}*���@��-tUQa��/�d-!��3+���Y�[�Z���תz#���b����s�h�D)��ތA��R�H�=�!�_h�X�*� `��9x���`� mH��_`Yk����2�*	\���4����<f��l�N�Z�s3�Q'���~'Ws�9zK%�SZ�\�KL��s����B����^@M#�m/3q�`:g<w��	5^����Z�$ |Pu�̥�����[�I8��JLs(�=��S}E鋀}�=�`e��1��E�u$����!�L)��A��9�#� P�;)Iq�gX�_f�7H=O�:C߾�@��6�i��f�ɳ./,��G�.����hDm ���!uO��j��4�gݨ�4� =Rh�5@�Z9��I�-�&ѡ��o�b�U!��g����b��i��A�Zj8G��H�Q,?��/}\&�1�hqC����D�W�X$���7�W�� ��I�O��.�3�� ��G#L�H� :C�9�A3�6���)�n���5�zOcG8A΀,�1�� )Y��O�L�$���$7H��`��HL�Ozq]-)�����h0���~f�$0�-�9AF�pj� dn,�;X��\��u��V\붚7�H�%@����5dp���}��]�9�R�΁)�,���fnQ����-����_V,�PH�`���9u/�F����,�J��ħ-r�P��F���U$2!���e�ݑ�~n�h֜aޫ�o�D���O��6�����X�+L���i!y*¢�
�/���&� �mC�(��a�p`��Jv�P �"@81�D)ʱ�`:L>�n�R-o�/J<�\�cv�HT�Xɝ�R��`����� ���}��5Hc ��>�k�+�[ٷ{�ș!a�f�dvHZ�4%L����VL���A.�x<B�=(�8`���(��U��. )� �0� ���g��p~n��Q�"�BY@�^�"���U�E�f!�b	��a S�:,|��$
�X- ]�S�u��&%A�N�!cj-k���- ��D�z�Аi����Jq)�*�y�R����P0j'�s(�q�C����� 0�%s�������_�Ph'GD2HT.��Wox h���2ƠRW�Q�I¬?�\�ȋ}���K_�b/�C�eX`��`Z�3�{�R��}֭Z�t�pו��C��{U��p����t�h�֡@>�!�yHk��W�B51;uQ�$Vi ��tHa-�hȒ�.ȯ�:K�ց�]�k�����*��!���%UX�R��0\���dU�-]U ߩn~�(	�!c�%�Jw���1�$	�\@�9�VE%{�x�as�-�S�X����>�E��=�V����뭗��`�l��e�uj�\�����h#k�����	�w�瀐����_g��_0��K����뷜ҳ���ʤ�15�(��R<L�;#����k2��.�!�{e$ҵ� ��0�A�<�X������;�������SE'�寧�XY0��veO�;kr�.= l���*�׉����,_p�(ꯃ/!�]�.l�b�~�<-�B�������! �M
�,S�=N�p�`V}_��ʰI6t�DXG��qn��y-�x�D���A�=C!t;� �YKx�Hot~{WQ���U��JP�ki�SC��A��؅�#����$���IJb��*L!1[)�z{PU�3�įZ�� ���4�ZS�
ݢ�Y[�%�;�S��%�nf��8�b����>�����a�
��x.���gC&U
H�:�N�˪_��<�GI��#� �<\L1����Q	A��'p�Z�����	$�;�������r��^��@*4>���-`!v):j�� �?�9��'!���Q2X%��U��h�(N(���{�����N��lr:�S�L�K�0]�_�D���/2H�-P�}� 1�]��%)�JM�	�ru<�>\Q��n�t|;��7K�cRB��^�)�|�m�6�=H�a;�;���6/��� ,��}3���K�;���9'�^��I�8D 1Ⱥ2B�	��%�#-K��~�h5����#��� L�yUW�O'��%�M�Y��s/���{�-������!˕��F@K�1[�Q�wB�W��']�r� �ܴf���w�)�@��/�L��c?8� A��C�� ��#�;�QX�}�܂��l[#�=��R�"?�YD�B���0������,�F�X��W.�k NE114�,���䶰��� ��ȅ���/,���f��O<5�7�7Suz��q۩�����o-0�1KڸY�kV���A���5G��g�{˟���X&�!9��f0G�I��*
yJ0�M>Cl�hܞ#	�*��Lt�~�e�E�-���B��x��R�*ꗼ0KFTh��1ʿ@�����_ 2^0�#�`�ܕx,N0妹�����}2�� _R��(qG1T.�b/π�Zh�u�Q�x���J�Mjn0ּL=�;d)	!�^`8r�mO����y_�<��e�VhSA"�{�n�FlEX5@h+e���h�;\yp!�a���2%Z�Q��4s������z�o�p��p|0�1��p��^|��	�z���}$_����}Lܷq����U��w8��X��~.-��^���!��]H�VӅh?1�����p#�`;bh���spA� ����!��S������q���w������ld�E^W�.���	�05�#.tm�1��?I��%"�-�Rh�M�"�xc�ѵ�G��{N��½	�5W �z�_��B�$�Q`�-�{w�'��p���Y�HF�9v�4�q ��-�V0V_@Iv�8.�(��	g%]zM{�4?�ba@ݶpo)ȰT	P���J[�����F3'�c�r����o�b�aU���#4�P3((�=��{�~�q��h�/������2w0�(��l��A��A:� -�a�������3,D��M������OʰR�MxVو�~��0�5�� z%����3�)��@s�ِ� ��,��0ൔp>���Em�b/1��R(��:��������/��X�;,�M�-J��X�E��A�_� ھ�g�	E�͒���G(�Y�O�
�T�h���D����}�u������iyUO��`��X�����@���N���Z����ubZ� �Wh}Q�|���!Ip� �rD@�e�HpcP��07��)��Z�ܒ|rx�O��B�0³�!�Q@��!?������8�톓)`/��a����a��/�
k՞�v���§���(��J����,��|O&w)�춟֙ �h���v�yW�;'�]�1%^v��a���͠�\i�������QF��Y������ �����H/��^!�^��6"�{8�R����0�M��k/h��ב���7��@QN�.+��\��[/�C��m���
JZ�w���,3)��y_���_�W��X?PU���E������xݘ>�U43�l�K@v(����o\��إX��x�Z��h�s�xJ����xrn"[a4a�΁��P��p~=�>��q����]�#��a0�j�{/�`�QP�P9O尋m`hW���_)yʪ��O�(9]҃���Wo����kq< �_R� 
"xu5��t����<�	�jeR��B|
C�X/_ƫ �Z^?�<�$'�uZ[`]���c���r�O��i�*�;R�ۺ.�(-��
`��CXz�B��Zz'�V���Od���W�M�2�+F����hF7�E.zAȹ�/ �6~���,��*����q�.1�F�f,�J��`�4��%H�!�
t��@�@혺�Voa܅�.�y����`����%jW>����w�Q��q9�k���_Gx-��HoP�e��K�U	�T�v���\�#Jم����)�A�s�^O%�/��G ;�U��PZ��WCB��5`�PIXN�Tb*�N���LSokK锦@�!�X�!k 4�?��� tf`!t�Z�
�����%eY-|��u�K�m�=K����`2��OL��Sxz,���}`�ikv!���Ulj0�#?f_�[�`0��91�0�m�6'���ќ7V��TL�J���Li���Nʸ� �������.����,�(�hp.��������*z^�;��z�X�1��
q�u'����øDn�j ��<%�w1�a��^�K�}���2\j�_�dk�BUq�E�VBf����a��-L�E���nVk�BD��,*C
.Y� Sh�L�m��J�!�p���^�x�N�*Z���HC_��>4N���
��А|��M���}8�ڹ�ӄh�	�{l��~�H�#D��r���(�C�t�	�'4��߱�jL3Y�>�;��� �0;�M���*)4��(�w�Ӏ�������d�]� Y:�LŝuY�*>� ]�ݺ,O�r�-iN�Y�iw�D
Hl�-[h;]\ή���yAfn.l@j<��P��$�u����)!1XʵK�	:��(3	|M���Xh��K�˂1X��*�B�	��4�.��f���k2na�\o�; (+�Z��C->z�'[���vuKH�Go��m%+M��bABH��{M@�Q��j�F�{&�ij��!ڸ�I��J���ţc�#J�e�Z���n���^�� �\Ph}�Xj�T��-o�YK�{���T9��Z��y�9�X2��0� ��0TV��w;`�[�:�%��&�*�}���[4��'�yz�	�*@A^��m	�k��l�P�AΉy�V
m� ��"���Q=��A�ұ�Y� �[K^�v�pڗ�LZ�%�z�D���I���f1+���I�����Wg�[8F�Y��R�v����O�R��.�t-Oix\.(Js��]�H@/�P�&܇�v��� ��YJ�~I~��QmT/!`����� k2���v�x��_����w��g�c���*�� Y3p����)��ݒ��K��ӐpBP��8�q���1�.����C��:�?���+� ��W6O{��횿�+���P�~Y$�
ڀ�;F�B��%�Ԏ��dR�Xz<�^!}��mK00���q�b�	�.�b�xE��ß�M���;N �~-�6��+=��F;hR|ӝ��͹|�'��U�8dS\�^HR<`oڈA� ?�klHCjT1(���&�QZ��~�'�� c��n�Ԧ5,A_C���B�����:�R��#YZS�����1�Q#���L��B�o�}(]�,�[B���U��h�m��ɩ����D����s$k�2���c��D�2�����J`?^�0|KU�� S�4o=1Ӡ��^f�I-�F�D�Q�o+I8��˃�dcj����3�(G���a.��������;b|���X���
k%�Z���f���Zr���D8-P�SmX�(N{����)XK�Jkq�r0/ �_�N�@	�XQ�L� ��'��ݡ�4(/���\��I�_���f�^@���)���<�ЂS��KW�;���,����K͠_7[0�|Z�X1?�@��}�C���
9hJ2q@c����̈́���c�N��Pc��N���7��5 �eH���zS��0�����@X�&|/�=~$�Q]1����[Y�sP��9��:����^�4�%���Y|P']fa��JX��H�<���[�s�׍?E@�ЏS8�0�� 9�-�ӽ��0�� W��G,��~>Kₖ��/Iݖ��!�p�ex,���-��Е̪�:uF����s�)-8Q�_�|t����w�)AԌ�`]����N��(%{v�2�c�Yh�A��.��?�҂h
x_!��?�W�:K���U]=�����򣀍�[� �)��gv�-|+'P%[^(`X��{��"�D�h���<Փ[U���$�*�f��x'��I)ٸb��u�N���}X�Is�W��D*�8-��F�����q)z�������uJ�K���W�<?:�yXLY���\T�l������%S�`���HfQ��TǕ���2j��]^F���=��ϯxo��;����-�F'������h����M�� F}�x)�(�ܘ�	,0Y1�2�Ϧΰ��v[]��0j�L {<����kܟ1RiXZ���xB#5���U�DC�j�J��'���
_|ûS	u��p'�:=/o����ګN���h�K�]!SW�؝�VG@��ZE�#׽/�	����!���M��_�Ζ/���-���\��PMh>���g���q���������7Zs�d��,�07w�3*%UX�gT(���}����#T7��(|�ehY��s�a%���|�s��1a��*��w��kG���;;%u�	��`�1���8_[ -�^&�O}�3������_�R_��{�h/�EtirW���2X[вb�I��Y�\�X��K�����!2��a��TgrCc��HJ�� w�LZ�^�&��E'��81A��89V�	��l� �K�������8�z���C1���(w� �	�D_�#�&/�p�`�FRGl��h{�)`�u�1H^| z��N�-�2���&�`gRUh"j	&��!���P�T�`i����AmQ�/]�4�ʍF'�bHX+��':��C��+1��(�5��x�Vy�{�	]�9,��
S�ȅ5F�ha=�(�+����u�u���Q��_��ǅ	.o�>�}Nx�w�ʕ����  �WHD}�Pt�b)�i/v*p�� � ���4�pP���J��� ���?[)��!�Y��6����(����o
�F�@fYea�Kӵ��Z��P*a�����Q�v�5��h��閄�x	�Zw�ꭀ�s�JR����"��;f9�!��M�	��w�?
)�	��
�-Z�q��?���!���}��@�Jb�m��\P�y'LQ�4���Wj4Tdjt%���=�чy�^_c� �)�Y�e��^�@/X�&��ͧ=�B.�g#a��	k��R�:� _D��.�������qx�ւW|
����c�)�-�	w���X3���M�(O���a[�Xh�0t>O �I�mY ��%?�Q�4J�����O��3!���'�`	T_VS������<�ޤ�-Յ(аom/kE�	,��Y�j	��[�d�s��BF}��N���h���dEd t���y/`U��@%r+U*� �jBK�J�|dfh�%��`��[0�.lB�wȨ�V$3p�<(���B�G>���Z''wDMz���wTg9��1��}�Xj+Gw���ʃ髌�x!��dN�Fw�" �G*>����P"�7ڰ���j6�r�\)]Y��!h�ط| ��Zb�'aW��* .��\;to�t(�'1��{	S�X".8j�=�*���uU�B��a��*�X�	%P�U��eqo��f
1�>�1V���]m�����&!�76��UB�Và�
1�[�:���	v>:fNdg[� ���~3=��9�7�6h��V�N����cj��L�o2�-�\$f�0^N�OR�*��,�;N���cn��X=A8�6�.����!�
�4}N[�0h��%`���W�v�>�ǽ����<eM��Ȓvz�>]鈑��œI���囫	�D�x �vr�'!}�P��vc̈́������+��[�#%�U��U�^�8,�ŀ��๣��t�	9���:(ˇðfY�����g�$�A0� ��,PB���TI�"����0PfP��$W�4�h_j����]����h���C�?��O���Vj%]�@���V]�D��'�w��E!�~ �}�/���3�*-� �w.��t��//���!��(
��߁�� H���8�_fJ_2�o�x fR�*��:(�P�d��x� �|�r�K��Ȑ��!%Ul�d��E�iWl�/TG�E�|�6 �A�"h�6�˂�8avAX�/���򟥾1M�g8TЇG��mT�/��<�H��2��o�G���lY|��n٬U���>��	_�:B@T�%@Q�Xv�,�;�F
��;f �	�(�#'�!~o�.����X��'Е�Qc�D'q�K�$X�R:���(^��d_;�п�}f�%�`�Z�OϮ��E��
��Cfh08YhGK{��=�_�i
�S��,�^�'�-�Rk �#\�Y	��H!zN�/�X���A�0W����Z�ct ^]�`�Ʌ���
�Xω��	�!�	Հ��z����i�~�������P�����p �`[�sT Xu�H�k{���,�:Q�  ���'��uF}�	�;��]�x>Q�ZH3$J��)�B�wq��	�掴�	�Te%�0��A�R�_�Zc%iW���M�(����l��/b`��i&!�O��qA��j} ���W4�>2��E�b&H 1���� UV���g�)��,��]p����� Q���sY���o~(�@HE���{P ��9#��e�2y�';�U�����UHB�VhʅO�+':�dE�	 /�F�^$a�d���,OM�M��v��vp���r1��VG��TE��A�Z(q�)�@z�w�k�AU��<�P��YR�l�x�����p�a��.|����P����q�`X1�f�Q�o�ؘjuK%�;�3��uph��U��� #!�����b�Q$w�}�G�1�Ԥ{qЏ�@�Q��rE0�5 ��O�W)9�Xۂ=M���UxhZ6�>G�*�bF_�Z!,�>-H�;W��
����RS`�6�4AK�2tna�b�j-Е��$A���`-k�m�XUf��W���,)� ��{U0(8h�'�i��햏�u,�6M/x�F;�F5�tE	h=�@�ѷ��Դ ]Ynfh� %0X-~�95�V]@&�튉�,N_�m�8�8��*�@R��J6��M���8\�fʫ/M��Q��dhAgttnx��yZ�3�kQUa�f Y�c.0.Eͫ�Ѯ� �f�@'[�} ��y`9(/_�6ٛ��'w׮�ރhE,-O���H-zb���02��h�>�%Y���� R��\�O��&��Һ1�<�nce���p~&�M�@��Ϲe�t����Y��%M�@6(�,Z}:EHT�D.}k<&���������ꢯ:�K����!�%�Y�m�1C�����^�S���B�+^xٓ`~��\iA����k�߯�$�����z���g; ���hMȻ�\\�5yP��1>��u�/��Ap�n�P�h1-������'����	_h��w&L+m%}�"S�^A�T/�@��n�p[��Y�z)_�Qh%�[W���CZ�W�H��! �e�؊���)����5�G�� ��N�i� ��K����1�!�:���3$��2�w�=���$���Ĥ�Ea�J���j�y[�ZC�7��`2��<Xw��z;ʀ��r���#� �w)���e�`	�_�� �?S��Lx���1%�z�	`�Y��7��|�H ��"#D��P�~14)���d�c ��Qy@{��d�$[�������`(h>U�q9�����3�XR+�A��]1�?�k�(��;��Y}`g"f������v�`JK{��0��t�LD�>~ܿO���@ڰ�R�p��I(�0�^��H
P��4/��X ّ��{��|�4�v�3{�g�0u�FHtHp%�]�:�X�Tt��ogJ�x^��rSq+���z�'��E'Pe�C��xJ�1�h V��cu&��j�[��U�] ��m�H��������0P�`!���,7��:�f�N�E������G;G�E!	��ڀ��〕v��}�W�A�E���0��0fJ��M�n;�l͊y�> �`e�-)�i�d�'���y��`(�X�]<�d������<[2ҶuĔ%#�׫p�o�!��׉�ݖ[~镀���*&�\��c��="( Ì�p�KB��?>d����/����y>�31#d;�@.z
H�
-[e�	�Г@\&BX(W�1���a��r;%�k�?�0���,w�+�h��t ^�Tq��zX��G"��bR}(-���U��(r� h�LG"�y�ܬ�ӈݏR,a*�r�N��3Q�`��;?�
7�a��|���f��V ������N�+��ߥ��(_�J��$�����*�����a@�d5o�;��-jKw!S�.{�	��t.d��� ������v���,[	P�|F(��p���,�MN^����cT)����Q��4�-'z�t�,w�)��e:��z&g�",x	_F|�9\�B6���̄�V��F�fR�ys�q؄���c�X�UjW�C%�Zu���6� `J��L!�H�`m��a�Tp801 ʸX�閿	a]�[�Nj@}TNL�2�}���]����y� ��vS��pFU̊.}	��Af�/�ϛ�og�#�,!��.½Y`%qJ'�5(�%UH��uIލf7.�s "m�۸�0q K5�2�	�&)�*���o��`ٽ�S�BP̨��%1ӋE�㎞�6hyH�B�(�Z��3P�5�� 77~��̂P��Ā��6'KJ�0��[ؿ�(�� 	#B���zCX3����DB��I)"P����:����A�Q�nf؍��b��0,���HJ�.�;w�~��!>�)`j2M�D}��Z��2�wJ%�+�C���%}�פ$xTh�j��9�W��.pdb{�	J,�5v
�9DD�N�Ftj�N1�@��'�2U�v`4 Ƿ��Xr�Z�і�h����~�u�<{)Xf^�H*_`ZB@ے{k@@� Q4 �н�^d�s]@�V�Q(N JYR^�+;K<*�SZ�/+hR!	���.��=�R�!��[yC �eXw1�Y�IS ��x��s�s��뀁i�Ӗ�^�0[YZ�K�J��\�c�(غ1W��,N��]��Y[ht|�o�� �j�����-Y�Х��Z.�?���2�O�P���rk�v ��-e=#�)���-rf4f.� ��*{���;��|�nG+�(ï w�-�݉��5 �.A�
P���qN��윴��������"Hah/;�"a��(PX:?+�~��q^���.	����R��R |\�_���Y+zM��'�3�z[��)ݗSͶt	��@_�=Дt#��AD����~��1��Q �1�_Y�Ah*l?�����}��dP��|��ʐ��v�������Q��(���֭���~@b�b�x7�>^2�-G��+K��1�^^�L�ZR����YSThv�Y����JMc��:��K��1R��Zk(#�����[J<�H-����	�~"��5^�㬉����j�5�>������uR�@�-�I�A�����ו�/���������{y�\b���?����~����W�_b� �-�]2QL��'�t���V|,�H�I ���G����J��[���Go��U�;)_��st ͟U��? "�'2�H����qw.�DsZQ��
)�_p�H�~���3��`��l��[�y�z�p`K1 M	w�F�	�*Jd��MHP%1��"/��g�0u%D�)��Ϫ��P��j��k�x�[� fRP�N9�i�8��fH�! �YT�,�TBuH,�R%Vp`w0'A!�C�W�@�&��>9s����c�Ttyqe���@���i$Gb� �	#���X�p-I�� _!�h�H��rT6��$��ڍ@)yW���^Eĥ�n���	�{� ��"� �� I%��j���`��I4E�b�W(�<��oK�P@l>-t�&�uN�9����v��AO���
)о<��� iat'�P�+��e�P����[����at'��.�H�XhU���1/� �A�r�����˻��H 	�WXU��ZKt�@ z�$���`�_���u�
h�F=!s+�*��n�(�&6�fP:�l�W�h��w�[ĺ�q�v�Ù�΂��(W�4�]�`{�pVo�F�c,��&)�Ђ��Vׄ����_٥ ��J�9H:0;��e�±LvA��LYP�&[0��@U�� ����3(�XY�3�[�o����R�#Ձ���I���v��.�?A��]S�a�2�"����<�	��\�?��+^��Zh[�1�3�f���k���a���
7d� �#�H[x+����40�c�� �W�H/�~_�
Y�w�s�-SQ{��z��ٓ��Z�+���悾U	_� ��$)��.|{���i��)�� �um�7- 5QYh
~B[ZW���ఛN�7�x��]��{u��1��yD��8��j;�o Q�h.G*��'��r%4]��5a/)��j<	�Y�<
Xk�l�&�L��HfO���
�|����5jL�N��:*��:��(5�'N���i���R޷'daM��@ �K��cE�����e�v#��h�2A�7�1��UzZ���[������h�S0���O�{U�b�=��&Ia1���wR�8����U�����lk!кd����}ّ`��+�_d�X�[",�]�<v(���ր�q�i�-O����]>�I
`Q�t�,���ֺ.�i� �(�'u3�]�0�X�`anD�,����*�{B�Y:�]Ie>�Ʊ���/_�`\��X �h�Z���!�a�S�S�d�B��1���
�R�}�L�o�LvQ�{��`?!HX@1
��}L�EV��5��#TQ	�@��㡛[80��n�^�&�ݥ����:�7-:�`��+�.,��9��e����@j�0�q09do �ށ�25?���o�vP�v��ڈ��S����P�O����x�����&��WQh>�;.P	�vRJ��CҚ.Z�����N�*-�"�u
=�-g�f)����Z���� �� &|���(����:I�!�5X�QУ���>�w��e0D�˶R������6���&KY%bq?@Q�:'z5�*�w�|�j-��Հb����-�r]
q	7(RW)wLv����9����Ä)�^�H��!(��� ۹�1Z�u��N��ʬ���0�񱏷P����9+�a��a(����W:�-)�� L;$�J�3w��1)���>��	ܝĂ�-^+���D�1ݺap�K�WShR	(-.]�D��\� [h�"s X5�m�~��o��$����du@`�JD�qLB ջ(��:���̉����X\�/h.c*���ꠋ	���8�迒JKx��`"�������p��j:A���A�/W����p5�X��5�R��H.[�XU�(�t��p^��������sRA \���V�Ѩ���*�50�{�<Pzć�?���~r>2s�&@��bV��-���U�M�p�ځ�^I(���p3!:o��U_l�f�bN�H���Q�zu�ԮC������a�����U��&�����N��(�
��H)�,��Nr�k����Z�AU�A�?.��][��1e���]S�`�������{#t�Nd��,��/�i��a��6�]�(P=��Y��`<�w*L4$�Xd�i�l�y:�.
�[-�y _�!��~����&�bwg;b����>a�(�����C,��2�[�r����^���	����0�X�ɲ�r���9(����D.�����R�������_��=�Ƚ�����N	�/9��.�������U�)T����y�񦒠��`�#��.�]5	�l�}Ԏ 01�4i|�K���R!Dyj�Z�i��'N"���� �jE��Q3�+��.�֜��;���X�g؉���I��\�Hx��^��M�n� �fZA�ǷA~+T������W3|LD1��-B���ѹY��N]����`Ir �
9�c��s��c�JHi��@Q��'lFv<5��(�����y{?A@e�	�rt�vӸ� � ��t<Y%�J&�>�R|���-]�9����n	z�w&���vJg���*�u!��6�2.�^���J|�'��b��\�gyL�	h3?t�h1���w%�R�`$Q�NJ��9��"A)6!:o�B�h~�}P���R'H7�X�_\���P��\h-~4��%���Q՜^Jx .P�XCWPU��mh4�S{]a=�n��=�\lw�?����-�+pd�S�@&��|��å�B��`�� ���o2b�H?��՜�u��Vj�d��������h/!�Fk�ɕ�F�q=.�^���qI�`X��%��	f���qW�\���4�'���Piȕ1��fR8�Z;�t��B��5(�u���U��Wm���(�1л� �L@�p��+�K�#U^eB��	�L��p�ǵܭZ�r�Rh�%�zy���g�8-��|�uu��z�r˚E�j�_H� -�<Bh�H
)���hC'.xd �@�?���X�t��pw�Y�囀Sh	�~�R�+6�M�^�>�̉z�
Kd�0� �r�k�Qڹg`Q���`��s)���B��W��P�R����m`P��0�r�Vm�j��0A�__�A[$y+a�a1 J	�_�����|%��� 0,4��h�&�Z#_�i!�-)ժ�6 ���2�e�V�_��1@%�^��x�25�)���`s�0-F|޳���b)�z�Yf�Z��mJ��?�^"��0yԣ�[��IH�;U����@a�9~u��k�u���h�t���O� ����:�$�ne7u�����wS�yR00K	>�1)ޓ/ވ�W��e)�U��-�x��.
�Uj	`��~��\�ٵ���-K�ʾ����m|Kٮ(�0@�N\J�a	����w���ˌ)	tu.���4ma��Cx�z=�1�N}S_)�������@���r	;�i�ԥ�X� �vs2�	�-�(���I�x/�
|`�5hYJ[�!v/�=�Ҥ�	�W����k!j�_w��!��d:@>�g�^)FtA�nm�K���� s���F`�q�U_R�4�HHa|.�Nx�3�
.*1� ���T4��f����!�Z�7%�X<��j0�'s����|��"UyR��-u|o����w�7��]Gm�5UB
h��|,�q���C���"����]��#��Z5�Q�>�vq��6�+�>�ޡ^X�(\B_U��r���Af]&�?+)�?��%cFP7Zڜ�Tb3�k�$$=�B/@{J�>d��ۊ���o�]{q�,>��G�f	��>����)�֘��3Ώ�r|�]q�J��5J����8��� Ӳ����#'p�w�����̪�/p�zP0��|c�_^�K֨r��N�"�Y�6ym��t�[ŇhNY	}y#��j�/)�+�˼^�2�c�`nܾ`�� ��V��Y�p%(��u "]�zHT�&��2/�n"u����[u�h�	�����*�k{)�͸�'!����^�W� ��D�5	RQ�U�.xinw-#av;p:�`x���R�/�Mrn,�@e�난�߅|q���E�Z� ���\�5)Ī�K}4�J/�H�L�����Y�;	�hQ�b�U�cP�R�q�π��M�E�&Q�!\x�{��3sN�� �]'.�h��)/Hq���|_b�]��Cf0ԯ���G��S~]�s�,�h��n8t�I	;&�ƅ,�ɧ���Uz�A�Ћ���V�!_��ob�7�^b�?�O��g��Zh�_7҃2V�z ����!w!�H�mY�XY?��q,�xC�Ւ�@KaF�����ҭ	�zqA�R1���J�`q��F�n�)"|�����%1�_�����[�À�;QXH	-CH�D�2�_J��_였���>
�hi3�a鷰C����:�(�^��u����cm��g�Z��h�1�_Jࢢ$�,)�I�w�rα��y�oY	B����\�bE����@ ��N��(��{��"H�h�J]�`���P�<E1`���P��� ��0z^Y (^�m=�W��_�aϾ���UgN�f�%8��V�<���ȟg,^�������A�U�lHv/ZM��[?�bj~L��v7/V넻����h�.XYR��J�E�%y��װ���t��pO��Q8T����%-։/ݕ(`���Ra^3���.@_�r�/��T4�����c:����u��5o@}!�)Z���Q��0���bw� �)z��iA�0������%���]�8�{�USt$�v!M�^�g�7�3����\��=��)���P�h�/o �4	��Y��ڗFP}�L"=E��Ƚ�c�P�`���U�Z2gQhhӠ��Z�,��1�D�ɂv�[	Esv��ך� hmq�KO�zj!�f��WP)R�)N�bPa�kj�"�=,�&�Sh�M�A�5q"�,'��@���� �flkw� �S�&`����*���h�4E�'��Uh�d�X]!��V��1�>.}���|A �c3���K!ʀ_(����O� G h�?!Y[=���%̬�y~�`#-�7J:CX$6�%�Hbh˺��1⁀5��b1�*�����3�W~�g�~u�$��U˽��Z��7�i?x[���j�qN�W4���K�8���N��K�[�%�:P �(�X��0N��#��_� ��,�(�(Q�̰�����hZK\���L�jY�&�[�HLC����H�&!��=K®��Z��ݔ��j(C�Vg ܹ�#���mu�qW ��`S
����6�r��y��!$.�=]�Ծ��t��$mfSR�w��?�����P�b%0��'��5T+��=�jt�w 9|]�/б8)K�X� ��?É_ {�O���v�����:�Q�'[�����mJho%[R.	fx� �r+ܬ��Ri;��0�y�kvDz_��H���4�8�����(�q�(�)�%!��i�!����?��b	����_v��a���"��-�fX ����^���l�w��;���� �R�I���n����	BHfh2�
m@v�bX������a(L8�(X�n��7�,0�bj���Srk�s;���T���X�̃�"n"�m��i��_��>��רEu0C�XwQ]�:���H�R'_��^Mh)�Q�LWxZ���I٦�F�~%UOV�zZ.�����˗Hud4-!��a� �h�r/�%ל�����_�_�Nw��n)iq�wĠ	�~=�W����K/�+�@�۰�L(1)L3���ju��vaU�F��[o�O-evë�@"V a1�_��	0=u�w,:@���� �s:��2��J�0�XHR�i�_���ߥ}�~��E�Z�����IR�c ��rZ��8e�@��?�H>� ]*�	������$ʂpQ�6A�-.� ����TM��$���.� �qbm4)�������h�n"y%�9�;6%Yh�5������L��N�+XZU���)�e꿃����E;��0W�%�R
��h�| o�����[�fQ���˴�z�I��8� :Q��$�)�����Y�J7���1x�`���`KN�D�	�e�=��`��6���D���Wa�xW ?�4�( Ѥ��Hng����@6��\�D�����������ץ�-$�U�`D>B�՝��D���	��d���!��㫠��	NW��Q�Uq�T�n]���&���0"�aR&L�)�WYX��J��R����K��[X���[q�s�U_�p����YM&<��LH�ܼX-}�VU���L/'��M@8@� �'���__��t���;�Yо 1�_�?_�{<E�2@�0Z���M1��) �-��n%"? 5����QhkMp	 [�^r�w�t-'��M�"�BUbK�	��H̓*F
�joe��grG~��g��1�e���H2�(��'�[Q� ����}a;��0ug6�S*���؍&d�&~p��t�O��<�f|j~�|��Ui�|��N��7}\ AX�V;P��b^JhA�0pQ���� Q�k�vR�V���' >�ɪ�� 0Zc�3X�/e�~P��-!^]đ��%k3�H���\�F�q���^?�]Bǀ��Y�K��R4�<aA	�s���C�w�����i0����p�%+���r2�n�f����v�>�a��N�<�2���&�����]�x./�g{D��HP:_w^�	���(I@*/>��[��C�(����u��@��>0�p�
�&���J(V��"�p�S�$%('�Z�L��0Ej��?8�f?bQEi05 :Th!+u?A�� �`l�A�y�~I�M�^�ّ�P�Ïz(U��L�^_��}�hp�4	Ά���Dd�0
.��4�- �D�v�*N�v6VhBC.[�����7܉�.	k�V��Co����� �՚��e�W�z�$3�v0{[Oy
��,ƥVeB�2���#����ءr~Fz�[� ]�|��=0�X�/����6O�H=s|y�O�� "P�������>T����8P+hb@h��mD?l8`,3xnO������!��/QuP!
�e)�u�C'Ҧ=�{�Y��D�cD뼲�����#B$qݖYO?�p,�Qw���j��(#	r�v�Z�!>nI�E*��z��Hb_6i@�S��r�����"�(�(ו�1�.h�,�1��@� >�u��_ �a��0��L�XEy -�~�G��r�/�����Mas� ���H2��FGv��@��J8QQ:�x3 w�):�@I�~�&Q'�5t��z, �d�-U�x����n2g5��|vx�[�͆LA�����%<� �؀�L#�R!ȯ!����?P2�[��{@sJ���'�$�_@�l���;�]e����a�o�1+�J����5�ч��0��G�O��"
�����Y`DR� TNl-�1i�)�VǺ	q_Ӌ��'��R$��2��`*� '�sR�kX�5	;��`D\Z]�v�(�V/,!z8��[*�&2���U[D�rJ�P�;�!�%�3�W��xr���Ҩ��� �k#/

顒�/t�G!j)�U$KAv=��w�l>�-�[h�t������K��̖߫�Jdb#t	Usٰv���U��-8Д�O�43���� Л{FO|�0�R%�9�D�>�����5�&'f�����;���X�TNZ�����ֿX��F��D	�
����,�����R�߱���3*X�h�!6���#U���Oq(�~ �%�a�<L���qB�X�$(C�1[�����κ)xN6���p ���!ӹ�%��BA�`�����K����sn���M<����4��ןU��wM�K�	��2Q!'��s�T��f�d�J{eq����/�o>
�ŀIς��)�!�>���j� �^��	\l�q/�<�ޡ�7SP�uP��!Hڒ �pOh_b�n���6	VuTO�b�� `�.�=�@��{q���S�X-P�����+��F/o�	� �z��ev��N��>5��W`<��3�E��g[v!p�?_?��+.}�k�u����%����2�z��Q\��1)�� �����/\�P>S�h�f�,���_���X���v�>��^��/	�9�z2��S���<��a2�1���^��X�vŽs2L�8�VLӀt�d��o�^�m��T�0#��Ca��ȁ�u]`�v�.��uj��E) !hY��0q'���S�	�UZ���1�@ݸ� B�,�7A�����0��)0��$���-�L��4x}��.L��j�q��<�k�qxO}�f1�))�#��S�h�JpL^	�1�� ���:!k�N��Ãg�;4\)T�3Z�W�/O!v�H�kYP�"G�T�1�5 @�%��.J{,A UJf!�Z5+<uG�>�1�-mo�p��e��z�%
�bmG	�5Ҩ6(c	�M1�ł�T(��3H ���t)�]�¹Sv�]��~�g`Z�"0F=�Pd��
�3&���T�	,i	��q"Y�j�<�O+nD���5	'JCQf��zP�\��lR�U(��Q���W��M������?H��%%dM�����u�:DL�>�]���-�e�sje&=��]��b��G� ˀ�Q��Kf�]M�X0ӵ��LŁ���z�;�=��0�됗 ���Q��f��	E���QZ���X�)�f�}OX��v;�Y"�I�����N����iv'&EMb-`��o{���1&3 �h�ٝ�#�j�yf�^R�6^I?0��6@�x��U�����JZ���Ҥ���K���p:*s��k�Do��	�}�0��&h��ߔ��M���T#��:y�v�Zh ���&z�@H3 �P�������]�
��	�^�rw�_���:I�=kS+��H*� �ö�0�[- �)��T^!W������� 0e�!�Q�]c�őo�vi�XV��_6�CNأ 	�hx3�^�����.�1��Ä3H�1輒��$�h<W/x $��R���O��i ��[��x�BU���Y[����p@��zixdk0���m�W`�*5��Ga�7^�>+��T����	�_�y�-�UXJ{�N�1%I�a}�wA�	<	 v%�������vwr�«^W����%��>��ߎAƈ�E���j���k	=�I[�L, �8�P������{�^Y�'��䎔���� ��jU{c �W%w.�@ tF5Unpzy c2m��� ���5�E�8-�u�.�&X(0�EQ��N���Ws�5d~J��s�E���a�{�h��pˉ���z	ad�q>���S�) �1�W�8+���zw���@�3/1�Y���.XlO�$E�J���� n��t¯G�uۘ�A	HNJ��PC1&��X�B {�Q��g�)�P�N��6�{�_��k'Zx�'���:��zK]j� �p
J��h�BQ.<����ߙ�q�.�rHIh�"a���(P4{��	K��L^�EP��{b�w�G<�U6�S_����e�2�xjDA�c��dx���!�����ʅ(���n��� R�nQ�~h��C�x%����z���. �h�r+{��O�#z��M�00�&��f0�)d�E>�dډ�z�U	Lx{�Y�tߋ�d|6�p)D:&]X1]-Pa�߶EN\�����6Q`��9$�m���� *cr=Z�,���?��x����r!�:1� �Uh9Em�`�430�Tr��n������&\)���xX��(�w��N�-h�}˂鼂t��-1���%蚽V<+ ��*
 ��#�O����Js�Z��P)�h0˱��
�Z�	1��+�^���x�>��Shwz>9[؜����#J��{�c����X�9W�~&���K��,~�����`�X���SGn1U��9�z�6>G0� �Q����)0����k�^UO�0�P���M8Bb:�^ -��`c��P�� qM.U/I 6�+s}V�	��$�ԙ9��p�*:B�-)Yܷ[���Z���E�й�/?��@�B}AX��H(���=�t׉Ɂw�;��q���$+���Rh�$k '�t�����(�}���X�:h���K�'�D�6���S�l�?Ñ=V�2`�QX�������h�V^!_��@�jŗ�"�t7h���L�@[�
 �c�������f+��&�:@��hb�B�9Df�Gm���rA��y��[��i��]���\�R+J����(Y���NQ�"L�hTv��3��� ү�&�	�����A���lb�v�.N	"b�h�g-�x�h�l�.}�'13^[S,gN��� R�+3�e^�=-g��}(�trG�6�fU�����E�
�u�-��B�%��$í�:[����kRF�`�G��Q�%\WTP�I^�V���ϡq����W���N���p,$l��	�s���}��A�Z��(���}��v�X����u��[0�=
���6� %>3�@NKc3��Zο8e��j�A�(��Qh7lG/��������C���,,�q g*5Mf)�	n�w:�t� ���+�N޾ɯD' )���^��*�����0QD��@H-��0���9(ޟ�/#�)��U��Հ�*J�[$1�6�e�vw l�w�P<� ʕ���9o��P�wt����]�z�9��5V;˞|AHl����+��֘�53�O�a�1�j���vl4���M'%Й�N�tZ�'[Z�|��	�S��`/[�A�߳��쪘�N��=((���ڲ�c���	st
����F�_���%r�4�� �p�*u�]@	뤿`ȰZV_)�� ��}_��,�͎�GqR�^gL�*m��-@�"k��_b�P1s��4*�@V��e����U��2*��$Zhbj�ŀkY .P��.(0&�� R��E]?=�� !TH%I�H/�@�x	)����{��!�h-�+����~xP��c?#��z�2� �(�Y��kSO�� ��kNZW�2��ė�wY�t�0Bh`c����,�h�6}�bH�:
J�GNot
@�&�[RX�Ä��z����sM����c��<� Dͦ�Ow��.����d��E棩�gv[P_���K"�Ag��N�(�}�}�`�b��o��v��� Mx���QX��O���M��K~�r)�}:e_�� �vS�1:� �%�/] q�t@��������N1o����Cm8��5t�U��^\�k�/�Y�\�@��cAP�Q�f��`%����-)�@zG�~{�Ln�v����'�l����{�P�����!�A�W�m������V+���]ny?3o�U41���h�\5~��9��wi�0s�����m&;7�>����Lʩ���vh@�+��֙ L=�)�Y%1��zJ2� sSP9O�L[`�D'h�;0��!<�R�1w^hu�@0v5��^���1P��`4�[Q�L��	���p�5���� ��R���uhHD���'���^-�+�ܿU���&苿��=	�����
�zU�*>�Z	�3�_Tn��W	ˢ�UO>���@���s҄�Mإ�Vn���1/����e�@�@8B����#�l%�]�S��'�Y �,�������xՏ��$���7!�F��s �3W�I��)�갑2U�sMU.�*��0r?�JZ��X�18�w`D_Q���Y��`�ƥL �B��<Z�0cEh����(G��vJ]�%Jp��!�R��4�i+�6�r���]�_�� FND���m[1ƃ}��xC�`	�ck�* ٯEq%�+9��.G1����PXCJםV�|���2!��^� �%:U� 	-rn�W5�����!A/K�����T1�]B���[�M�z�/K�p#g�_3�W���� `�[c4�dD	҅�S�}-HUD�:hTFL�Y������qrd ��D^.]�%t:'��W ���@O��� ��_��G��νfK)���c����{7.~k�,}yI �)c*\+{�����AZ��|	�@8�=�`����E�k��/���<�Q���:��]��y�L(�z[�5�5��'��/p:��2�z��:�2�
�+�b ��+,�&	�.pv'���me����#m�Opp�3+-[Y���ӡ���h2K{#4R͈
Z�i}�l�<*}��"�g^h�
<,��3[ XWR�5"9�y c.�!T��ZX�r4�J��m	�/�ݪ ���A
{����Eu`
mx��3�0�.�P���ر/��y ,�|hT|r�Z}�]����, �o1e�8п�iCO���f�0���G�J���w~�{�7��p�,8Cx��@qP�����_���	����d}X@���F�i�1�'p#��/>J�=x��I@h�S14d)O��N��7��[�N�� b'�aK¯٬k_���np�7����O���J���鯵X ��
9��3�,�L��<�r��q.�h���|�v:��2Ma)� L��׫:���A�+�!D�O�`�l�w�sג��e�6T$�d�sĄn��[��PV��~w`k�q�jO3)�Wވ����o�,c��aJ�B�;���^�M7L�4=kଈ��.�0����Y�H�{m&�!��~��b��%/91�E�����Yyh�G�%�����@r���ҽ��G������0��h�.���y��
2� 9��,A�j_���֝F-�ײ��M	�)�]<D@�p���AI>����!B�T	�D���#�"���UX�y� K�?�A�h�R>$�D[;���٣��o8��n����u�(d3��f\�iWy,Z�!�sq�*	���7Pz�G���ţ�%��0�0�~�/[I��~ �fZ�̀�����Q��(��Y餻�?/!�}�_��N#�� y�	g�^�������� �X!���Զ�P���pt�	�!\�'tn�*��PR-�YHdT �E9�;�qC�-p|Ւ	
}L#D~fG}��S�D��QQ]�0�\�I~-��l�:�kAO��o�&X?�g�s-E��A�: MT����\�U���y�R�Eќ���M���K��Pr`��.�V��BuX*�	qw����h�>p}(?]�\D7�����3'/1�
c�g�	�t�؍K[���q.�o�G���)���,��?.:�����v����3^������m���H���5Ȁ%;��S�̀�s{�s����l�ޥ#(�B 鼵V:��\]�	�#vo���L�ZUc��	�/) ��p�L:���=ջ�g	s;>��R�넉ڼ���	��Wed V�n{�B��؆�M �� ����1nԀ�p����#�����Q�4tv|Ļ��M4�}d��U�I��U`�!z��_j�7j���&`ݠB !�^[�QP�74��U"�dSQ�<��1�b}e�a�d�`(0��[�ŉ�P��8a$��[��0{��K&�.F)4��<ί↯%�b�]�q�C�	��P�P�h%װ��'�T�U /����������G^��;�	x�1��D�] ���,2�H��k�y@5��+�[k���~ ٜ-�C� Wi<w���	)�^� �(Y��_��۾�cZ����2Q+��
*��<'$	E��%�)F�j	CMl2^�K_1�D�\�b�I���@��x������_�
 R1QtJ�^+��	h�jqo-H�t�ޚ
\E؉D9_� I��n�X�(�6yv�[�}���Pk�B���Y8]_�	5�}r�j�qR�s��ZC�ゟ���Z�P�cX8�1.�zHk�
9�_Kc�b�^����y�%�8+�,e�>�a���/XYZh_>D�%������	�k�!V�GH�f{�8������("؉J�:X;JR��r�QT�s���N��P3O�
^��h+{����>����M�1؏O�0�h����F�j���ET1��)���P��2�_���x8��Z��^�����3Y[��?�l���vi�)]�Rk���ʰ� 1M;��2�P��8Tk�iq雸�u�A�H��O 0��_%�'���(��L��D3�s����DZ������-�>	\����1�T1�wC�q�drj�U-���p���0�	'Rai�uX���4�K������_��C�|+��:���P��f�@��^��-'xP(V�v �ߒ~w�^��E%Xf�&L�f���	y��D��̀�黼�\�e���%��,p���K�5�d
M��Ѓ��	��(�FA%�26@
.
��.�
&�+�.� "\"0��,b�P_�E�m1��B@!R(�TC2]��/���G�%�j�B�&(W>� l�hl�3W\t0�%�T�ąD��n�H.T�)
� ��N���6�^X�WH�g�ޯ�ᾨ�H�2�K]� =0-�1�
���2���T�&46��HV�3�b��h�\�<b�I��A��g�:=��K@��墀_wơ�^X��X-f�_�z�3����]MF���!������S���/,�7��`��Myo�.2�E����@l�lE[�._72��{Z;�V�������sN%?1h[!bH�.	U��H ��識�ˢ6��vя��i0�~�%vW!ݸ�R�
Yg%� *B2�d_����B����L�<d�}0�3�A�M.�6�$-� b"_%T�A>��;͗�� A�5�p� D���� ��U�����M��4@!U �R-��� ��t�駾�v�ZVUy^R}R�	)�1�u�D��@,�b\���X�-��Z�#׮R%t����|�����=n��)�B ;A�h�S`�V��MR��;�����ah�L|��
����[5h�v��3��C)+�Z���2���*�d'�)����'��gA�R�h,�@����QH�?�QX"����-j�bmwe���T�����>6Q���J��������N��J5�]_�!,���-�7������G�ܿL�0�n�Q
��d*�zSm?�|����e��)�@&�l%�s��ÂC�@�U�I�uH���ѹ�><���+Ġ�Gf|8h�*g�tQ8�� 1lR����	��a�\hp(��� /��I��/����P,e����\oIL�B�LF���@xȰ�P��JP�HE=�1)�9�^�:7Q
�a�X����s�K��oSC�僞�	���E��Dalh��t='/1e��� V��Bb�&h<D6p�(�Ț��19�����½�l>
�a�7)��pC'�j\�
���4��]���`� G�f�� ��~7�@]�(�[h`���'o�;�y��YA��H�ѝ��m��S�0�w)KJ����!AC���H�pX����Gw0�Y ��
���}~;yT�?k�u_�wxRP `v�b��%�G��8��:<�騷���1b��_e�t �U	��\(V�:�{*�Y G$��Z�~h_/��P��RX)���к�w2��Κ"���H���>�'=�h�+�>�ς���e ��fX���P�R�(Iе��0� � |�`���J<����V�!��)P<[,�����v�	�!
 �q� ����!�e%?�E RV�: {1�>)��?��K�9���Lz~�ͣn�H�$:l�ޔ�/�����A�`EH5yۄ���c�Q`�!Oز@����U4�]��'��R����l���34�DV���^/���	!� ���Um?Y]����_��ùK�';���5���� �k9�O����R�'�*0W��ڀ�҃��1 �ɹa׾�	z�K���A>�2��G�㼖��'�`�5S�\������xN�7Y^1�	�bR�������d�X��,���J�_��Z'R�N���O����%]�S�%]�S�a���g�����B�
��ⷠ:U�����5>�z$F�"�`[ws��~�f�E4-�N�n� ��q~���XZ�&��F�À���SY)ӽ�I�+@S�Q>�z���;�$��	a��m�
7��\�(b��-�NA�!����X��w$K.l31I��&8�&�nzF`R��k�h'�[�ڒ����H���C�3y*�H�

K�� ���p�����⤪E@f�R�u(�Z���20�Xhw��7�	v>y)��$T�]%QTb�	��� �т �ǲBx.�h�	w���`����@��Ru�kh�}Z[��'m0|Q�(��y�ْ0��^��#����	=�X���<MS��0]+�lK\��j��#/W��RjC�MoW�<�{�/\$s��.���C����t|Q0���X��e��Q����s�!�1E8��+ecb��ʲ��1a~*�4ꢒ�����8��_��6���Cu;eK]������@IY���JX"p�-�}	�o?�H-*
x+	�����U���������J{�yp~�rBZ��Cp-n�d�Γ[�o�-��G�H��WE1�)ݙ+K�(�~^�΂��N<vڒ<�����K�W���DD�L��dA��.�_ �܇H�L5��ݢ�� ?��<�_�������O~XH�
D���I�m�X�9�\%u��]����9& �*N�����#`�x��r)|��_�`f^��W�$l!13�H�-U'�X���>�b���og@�� ڹ�X�
�p�X�l>$k�lv���W�X_#	.�/�K��/Ȭ�,j��n$�c���F@J[^ż�-��N�������i�1�}�ƈ��cr DS��k�k�����������BN-��%�~b9+(�� ����J�Q#�*5����q�X�%��n)�D�_!�Pj�,"a�$�r�=U�ɖPog"c�}��K:�Π�zn�p2�vF�pP;�Y5`%p���[��L�_�o½��W����^p��Ot��εU����lm�^\��t��OS�1�h4�EX��`�I&itxT�%������13!.t��jn*��bQG���d~� �Lx	h�"|Cc���{~㸎��P�e��0������X	��Mj���� A�z]���(�,PA����؋�P�_y��.F�>�)����z������}D�r0�,u�е��,�'�ÃL�.�Ed-�H�[o���!�+��{�
x	�Q�wֲ'���`oS���4?�ђ�Gd��_��A`0�<�8C༯��xoN � 1عu�3_A�3	,�	���6D1oD%O�nZ_�yz�P�R�pAQ7�"�FUj���:��5�b��Z(qg�/��t�^_������``L(}O��01u9:�o�p=b��/\fx�_ΔO������-�M_�+ǸpP}!� ؿ%�mK�N˱؋pJ�'�Z���c��Jm��RXP�%^� �(�	�J^5����]�_F��JD�� �O�B=�C)Qޯ[��f2~<L����-}�U�5��Y��io��GV�Rh轠�-������:��T� ھ'��p5f�~-�9=/r�Z��^L-�j|$%����&������k�C�!�y������#���G�����e�h
B���WP��y=&~ �X��B�L�0��I��H�sDT���g�_��K��X�	��>P�xc,[2�O���U%5{�]:@���c 2Xfh�~�ѵ`=����ш�I���~��_z$[�k&�%�L�s�`]�&pb�p�'w�@����u��1������Ff����r�{$� ��1ݠ��&(d��SB�������Z���Ϩ�׮���6%�HD���Myq���RaR C�	�(�w�����GK[����2�?�������U	��M�)��;(��!ȹ��o�|%P��K@�c
����e�^˫N����]`B��ح���r�L�?1и0c)�,@u�hm&v5��`&��_�F\�[�@k�\��C]C^�0��N4��U �@-�=!��7A�;ݎV3��-=25s����&�����	�[�$� �&�1��PG����}s�X�%��hl;1V������?�J��/5AG髞�|_V���C�����Bʛ8HE?B^���Ц��un^�����F��%V���Q��Ɖ� /S�ӡYN�Vi�_.9�y�z@�v0h�ip�"4�v�OD�>�����9�V��	��~�'Ⱥ��[��$`-���+wNhJf��i ����9�W�G�L����_�������!�R���C��X���(`T�0��:Ŗ^LS	�,��	�|��]��ɏ���^��i�0w�^kΚ^�@dV��hI7��J��5��!^T���,�VÈ�1��:�x�6�Gh�7F�_�t��Pw�"��:�N	��H���/���1�@�-�W�tz�(*�k�|)�$���f�y	�a��]I�P�<Щg���o�ȃA[�w��#C*P�h&�>�j�P�~M%,�22�=�j��dSI%B��X��0v+���̏���ƚ�%6����"�!=H�R%��}MN`��t����h��k0��W#-zp'w*�Yiׇ� �V)�Z]��Shz�oYC�����DHv-n��\Ph0.1я!�-����w��*о�)M&�����.�'-u���㰣H�cN�O:-<ZT��1)z�	�뚦	śd�6_��8������������G�
`���:G'	!��y(�2s�A�FHbF�CwX�
h�N�ݸ��#0���{L��ȑGk��g|r��/�9�J����3Ì/V�ֺ�bR�����k8*��A�{/�_�h����`��l$/XT~l���@P��
�Z�.�+����h�`�h��-w�nX��G�%�` ��+������)]���=J���%�����4�Ѫ|�v��Xa ?/�X�����p�-L'�K�ۜ#)'���( �������?Q��*7��v6}��a����qE9��5�-��;��)���A�U1r �Ä1��0I�
�7�r� .5Us��;uS��<�Wh# 8\�~�D��ۈ��p*5�0�A:�LD��(�(�\G������5y������Nb'|�/��H�w�H�<q(Vd�J��4�����1I��fJ�@1���z�x1�Fc0�6;@Lz���`-�~�%;G�I}�{FKH�v3?�#^&Cu҂�i�; �)�01;��Z�Ǿ��pa��:��L0��,B��`�P���I��	 R�R �m�Bp�����+2�=�o ����껍$53,��*�A�FE�!�)����E{J�]��)�!�r��T�ͧ:�g9�N��T��)W��h=
�3b+	�Sk\��Q�D,40HG5:���aNMơ���  ]��1X���4+ S�Rb(˳��`SPhy5DL+[�j&�J�Z�	�?;h�:��5K�Au/2�)���Нu��*�L
@*�[�,QVY^��1��Τ� ��i�!˟�C�R��^��ǯ�h�Z�Q3�+bkU�LP�V$��*Կr#��!F�'�uW%t� ��bsL+c�d��ʩ!�0��3L��7a��r���b���-n�1(�U �	Jm��/j�)�bEAϠ�.�����i>��m�D?�z���*�E�4P�h aLoj^�� ��gzS��鈶@��j.X{��k�_!�Q�x~H�-,�;� �e$�b��	z��"�)��1�z˃	���D�%�k�� /X�x�ufBP�`����j�y4~�:1���r��_��c7�0 ��i};H��4#?Å�+������o��b;+p��C�S��
h2c�����3Z��߂�w���y=, �h�/E�	��!����dy��_�\���q��w4�����d�*�����Jo��uVl��K &�C�}�X��"`�c���@D���L���#.�嬫`�l68>�Lkԑ��VT�C���_��,ξ\5��ͿxH/T�qkp�;	Å�����DX;�y~z<O��������a�!��ki�Ũ�9�D�����x� ~-�R���h;g�tO%��!{��N@HUh��Oe�[� kE�����-�=Z�
qD��P�>^3)�1
czv� �S��PQ�%<q"� �_9%;�1���Yd��)ˋ�Vu0�o�[h�|Ļ�C����3��o95EV� 	[������w?�m�r�j�:]�lL��NP��g�_�˵!���*g��cN~[�'���8�n�{�{$��,#^��D><�ֲJ�pxR��xFX��$)�4	1� X�[ {"Q5JH-�z[݃��O_�o�T�5H���Z��6��R�����(�|��DS�H%T;ǚ���G�β�{Zݐ/�x�w�V��N�� ��Р��CYNV!�[���9n�Z�YZ1�[@׬!�[݅����b	�R����/Q_�^Yt�/Z��d0�X_(�� }|6(k�3�b$<����f[���t�Rh�XA���@Vl(�?W
�� �Co�!y�5�3��$��i�?�/r1� �]�k鵲&	p�5�}�gP��X���;Q87�%=W��v�h���1�}�~k0�P-��ىآ͐��@��h�}<�m䀾��=�O����� yR��F��n�� ���%�ud[/�ɇ�!�q�-�������!�]̀�5D'3-K(.���Y	���z����1���q�\�:R����˓�%�I�1�$g0� K��|@�X���*�	���!@k�60Yx���oCF1��h�Uo �Q�'��|c�8�.�V�v�y>d�xf(��T7.�X��nqJ�٘�}-�}�I����Y-tp���@酯�n��oBMQ���$$�0� ;sv�NI�4H����wh�C��>�-5�\b`n�1_u�<��&��S�Q���Z����< �{�U���h�\]qA�.��
A��Ĺ��A��|�o TymGO>�;�"Le$ 72�8��r�p�	��@�-]	\x� �9e����΂I�.:���4y�#Z�\��n�<V�t���3nfDO�p;��%*� N����b�u` �EW;g��P���u������3�ib�������5]���ٽ.6�PL�;}g�)�Z1��򮾃�[V���YGh!������� *n(��{M%C���gV��y\���(0^x/�^-rb j~�{!��T���	�3�
pl�P�,!!�z����^��};-# ���5�>I+2E����p�usM�I\UW��g<�\�M�ZK��(��Ns��<b�c	��w��V}K�c�0V�?��ib��O^�ǁ��w+7@ĝrQ�¹C�����s`��6�D�O�q�2ƒ
�5�� O�L�(Y� 5:`�>��L$�1 �� C���a��n/ !�SZXR/���������iR)����	v�KA0�1`�
;�|�R�'Ϝ �~GN[��/�� W���06c��%>=�z/� &�o/�Kt���93�W�#xH[M�UJ���8�����I~1Y�%BC@�c}��\mo���2�^��'Tw�W�c��RA��z���Rg��fZ���A(�0�#��ߚ���V|�+Q@I�1��@Jp�펌�H��~&N{x��	�+��ʌT�a��0�S��yJA�4���b)\cIu��<��y�l)�_���&���XD���	��,1�W;�u�6=h����� Bl#�o�X�0'Xz�ZO��<��Q��sE0!p|�D!�z�#�̞�\�[��a'zР�`��<�`e�JPA����=��n�F��Ƭf�]1�QiÄ����1:�s����XZ��'qo^�i}#��%�WX�
S�t��L�8W`5U�	� �J}�� p�"�UV�a�)�����kհ����(����J���=�!f�f������f�3~TG�x?� ��1Y�$������"!Jw�,�a	��	;O7�蜅���>��m�1n��x�Zd o�龁P���(���rf?�Q�i��@x���UD�'DE�Ih��oLxp)~��,:�^^��|�z8���+A�2BZ]�;iDK� ��B0�4J��0���� ,� �h�H�0Z��8����KV����$���Zt��Q�o���V��ǉrݡ���:�Z��)��ʖ�.�-�	f!+{�^�����'mQ� �
�B<��(�n��9_q1��h8���R�"xQʚ�}�6�=E05Ab�0�C�Hl�!.	�}1>B`#_���Q+�?�BR/@}�ҰyK��+A�(�1Y�Z���AXLMo)*�DƔ唟Ab���[1� 9$��8�0Z%d\hK;>6M�b�����3X�}ͪ08�	sB/� �Kz06��Y)�UT�(3�*�-�r�h�,���c�bv��x��S��q�YTN*�i-��E��@��wHVQ(UZ�_A��R�X6���auI��e�'h���Z���/�XO؃������I�f:��0ϯ�b�N:�����DI�~����C�)JL��� %�tb[u�]�����i�.���< ���*�(��|�E�B�]��`���H$1���d�ۂ!��g1Xk�r�wZ�.��"�0�\Hlu��"�:]�W�ZPmo�O%[�6�����;&Ȳ�j��c$�AB/k@�Q����_@ �B����>�_3ћ�%��ʠX?h�HT�ý0q�JvRG k�#1E��AIs��(<U10�7 �Հ�0o fU[�D��p8Y�mK����s�	Y����5�WQ˄�v@]hzh����
������j���t�� <51&u =>bW]��� �Sʯ�X� �e�����t)���'5� ��QH\=�� #��h�0��.ߕ\�b��t�-�Rq�ɔ)3��s�Z��������c� j��[(�X�6р�pLL�l=VS���k�0�3���*�P�z�[��7�(�-�M��P�����$���'XM�+�R�����V��-K��lҕ�I��M&L	`k�D�%L�j���s�b�,
U�)��@����6�r�Tb��(_N�
�5���\�� 0�!�0A;�-�D�yh`}���N���鱤�����*�	Ff���t�Z����_�#c-^ٍBj����2�L]�i'�5;�_��	��Z	�!�E�v���Εu�=�{�2���h��*���5�'d$	)�w�GB���.؆�D�:S�F�|�Ӕ�Z��p�z�
w�0B�N6����A;�k�G4q	^QTY��@��N[��j���� y���)�1�QX�^��D��	�B�&1�Ԇ{����Aj�e��o���+/K(}�_��Zz�)Wـ8P���L��ͼ�b�D5����߇$=�8����/�H<K'�oX�{�Y���v���(�O�R�q<*�=�)�;���xN럊O�}���C���QƋN� P#�& h,fp?[V�8>�s��^?�A*KI!�Ol�`\
/�GC���(���������D<��5?7Ln��� 1ջ)��M|� 7Z:���_��I_A��1���V��b�<V o��xq)x�P�_���V�|�\Zd�<�Z���%]`&�Z��zC��������<Gw�L���4��^.]ns��1@N�w��v5�A�?��k�rvr�D�@�\n����v��iA]>?BmW��倒[��y.3e:	"U�]w�� �1<0�@�`p�˻�v��S��(�j�n@��`@ <-�Gz%�6/�����[���(�'c��	`� ��ͺЁ6C�^i�%������-׉'�Y@}�1�/�*5�� XP������4��(�S���M�Z>�"�s�Z���';W��Q���*�E?�)��ER�r�mn�I J8P@�1��sf�����i�/H&�B���ɜJ-�R��(��O��#X/Q�.D��+�l��^��!����W~>bqV��]?҂�J��É���ǌ_]�M�|�NA��H	'�M��;��w�-h�Fr��g	�N�Z_��t��3<�z�Ma.X����T��p�Y ��Ә�H�P��7�t[X�PeO�����'�Y8o懒���SW�D�
!��
�2��Ķ��x�e�PC�x�1�^�<b��������#r�d�}eo�@���[ρ��K�l���N�����Dg.!��Q��ߞ��Iy�3�J�!���J�(�4��i�T�6t-q�)��@��&�`W�~�.�@��Q�.`��X6V%s<���9@��v�`I�H2%��~ 5���)-�1߾S�+���@o~B`�hw>���  �����v�903`ԥ�QKA�z;1�-�a��<�� ��lNHM^W��((���!��Q����h��V��s}y	�Y/|��	hu_���أ1��n���q%-pX0�rJ%��M�4�Xqb���r�R-@bx�y]��-d�	Xx� %;����� ��|%1ݠ��A5�p6�X�� �ȉoQ¸��_�	U�Q���!�y/�wp���A ��}�3�:L 5u�O.�2�f�!]�so���	��?����9�f��0�����,/�-Z�%d?�Y�s��v[=.؂�1����oV�A`g]��El��ǞK�$U�v���N��?��˯�[å_�t��kh�o1�T[;��u.ˁ�?�	j�*�����F܀�����%���,������t��x�J��ɉ�9t����ȅ�`�Q�1�J0����@2ZD;�	��b�C�����Z�K�� ^X�F�eŬ(�*e�m���'�1��0�:-�>W� ="�`���.�)gנ��y1	�M_#kwY �*%)���D��$ fh�&e�%���d&��U���L@kt���O�%�7���Z�,J>��C��{ìl��!^��Fv
�#��<�ydqk20Џ��bA_k�@�$������0�F�L�4��ϋZw<	h�U$�4��#��+�E��g���҉�Tqz�S�����Lu�T�s��,y4r�X(�	
��@�S�p|�o�cK��N1�h+�t�*z_8vup�מ"��P����Ahri�#L`��v�bP�R	���&.C �?m���鋮	_L-2�Et�v�<�@��}ٵ^qR`��[w���8��i�)���q�?����	�I�_k��䁈�;���U�bL ��*vDH�Ziw9�9 �Ӑ>$�.�:^�Ɣ)p��㕖��V����@Х/X��_"w`�|M�E13�/�)�2���~�Q��;�8�T����Y0��K��4����J뜕�1.���%��3��K�; a�P�B��~���:H�[9�q���ig�(�@�%X#NT{�U���W�`����A�"�:`v�S�x4
q.���cT�J��`��^[��o�j[8-R���v^��	W�@M�?��>[�:��^J�a`(��AhEz�y�	][%`ЂX%��1Z��@�dNh�j� 1Z��0|{@��- ,NR1�$���3 ���3 1�.n�p����ҍ�@�F��l�W*w�U��g��!�/xu�^Rh�4]���_���w	S]�,�oH�V�\}Kʫ�1������՞���	5�hf3
�d�/̲s���R�-B	�(��A��Y�ZuX�}̟Fm	PW�.�`��Ak�j|�4�	_�� �lĕN���L$ Q���.[�����N���H<T�*B&(J��=J���)1ʇFB܋T~�� cY�l
oXt���^��rP�h:4#R����pc�{�4����/�z� %80�T]������3(	�z��0Í���V&T_>���P�ͺK�\�w_�O� 5P{"��G��#o���Ӆ�*�=���l.��- g��w�A ��On~����?J��\0&5��u�����*��K[��X^�$Xo��������g�)�Z2	}i��V��}�t�T�u��� ^!�1��е��y'���>`$�і4�������k���Gc<�Uk@�X)�*[��d ��Jc�k�JW�'4����(���f0�h�p�tI�-�:ejt1u2����|W��h��N^�wH�������c=��ޣ��P��(�X#9[��<�ݖiTA��F+0U� {�()��nvF �Z �X/�Q�4^�jLH�Z�(�k�;ww��P�d@�%��|�Z�����M�7�?���hrF���hH�S5RF�`��3PR�7/bxOG��(��5"�[��)��P��m8Bر �n��S�����xP%t��	0UQ6W�a�C��+Y�8�fOj��E	�b��5U�P�T��䂂e�Q�����]Xm��8�E�W V\�*T�s1溅A�	p<X�4#)�4	����%	}Z{R>��>[h.Fz�vu�c	�1����D�5P�=Oj�
gx_��A;�������%����y�^� [����`���,8���<x��(���@�oW��U���wex��d:�%�4[�=?�8�_��Ԉ�S7ף/j[v��$f�D;��*Z;htO$[�Gy���ti�Z]Y�IW��]��#w/�T�n���]�pnF�˽��H��_�� ��P$@-vX
�������Һa�Uh]'!�Wei'rY/~��C �E�j�+gL�p���H_o�A���m�k��&7���/CmB
�D_�{5�@})Ƣ������jW#]��0r���fBlx@m�Dc2�}AL>@,�E=�5��W*@k� �1����c�^d�#�Z�07@y~KX���m��%������<Vb�[�5,x-U�*�'|2b�5h��R��L+��f,0$]YA����{�P4����֖���w�Ug�O�����`0��?XR6�&��դ���<Cq��2ܤ`Z�H�S��vI��U���B�d��Q��&1��`t��r���N����J�� Z��6�a��������!���	:3[T�7�7�8���}I�p���sF�1�Eo�@�N1��N ���� t-&npQ��5��b�������|OliV�w�q�N��v��/���^�aS��h��1QA���&)p��Qr�0�"d-�:��)1������s���`"����fZH��3O���i�n��B��� ����6�<@�Kjt`����-~zN���%���vJU�;!a���.� P�,�A��X{N.%���5��jF	�.S��%�%D��wژ�&�#Z]h:�/�=,R���S06`!-/_j:h� ;���Ì�;0ΉM\�D5u���RL� C+t���p�0�p�#�TW��*���R���wR� Q��hi.��GcU��>	���|��Q�h@W�2z=}�����{���
�R�L�FZ�C���	[��c,��%w��LǪ0�����@X�% } ���+��J	� �vN�v����<���0���R�w������ �1��n`�0��X �c᳋/"	�	k�䦄�20�h+;�ցx���;J)�?�ć�a���������@�!ӆ�V�Q����\�O�Gt�3	5���XWt�]� T-	_�]�}u���2��fRh$caD`���=(�[ѻb#P�.�+d!�*N���WR�Ȥ�?a(��3�XD�꿁E���?�V�5\6��Y���&y���<��	�b�/�)�4-
��5"�Z��@��)o�J��Nӗ����B���Y��F�s��G�bj� ��F�n|�����aa��!�hO#ie�:	�@R��a�p�E���P���kB�u�"Zu�������'mE�~�
^����t�O�r4��~_ݞ������� ��
�I
H�	B�x߫*����U��9a��_��P�"��� ���4����Z�	q8��qM���'�-��`븹f>BHe��1�;�]<F$�ai�@��L��!��9�EԸ���z-��hO�	Y�d����w�9z�`*�0rhLI/wn���@V ���,�3Iu�qX8(��N�4���V����=�ڠ���n4���3v��\�[OP���-?R�p��+�1P����T�������/TAS`5��yJ�Pi��w�y�����nf�7T�6��l.�$����c��C���ufS��	D��ܚ���C�dl5�!�	3^Ѓ�y�n�Q.G�U��.�;��"�@*ur/���%]��:�1�ha|b>~^R��ѓ#U� �u+�E1%�_u�ހ������K�t=�Z�a%�i0i�hG8�m&EΟ	��݉�՞�S�P��RJ1¤��	0�]���� ��{u&�?o�n��ªY����/��5m%)ʀ��D�MWJ�@���:f-�)�镺{$�O�/���S(T;���"�e�F�'���绘%�aC��[r�BQ�n*�k�`z�6$���˖8�Q���t���#\X2��гu�D�,p�<�=D�Z������}|{tjAt�R��I>�T��i�S00��.C��1z���^6^M=Qr'!H� D$	�J�Qs�-���'�%XV���Cp���4�-������R[��0�X4��#���/�	����i
 j"�z��[��ބ�܁wY�E���j�����%_�P�m:����M��B�� &�)�^�H��\�rwL��,�m)!���&�LX���K��l�5��@� ��g���R}��)�����P�--��f\h�p�w:o]{R�H�����%��ɋ=J��� �M�y�'�b�w~o�\��h1�>�8]�}�2)� I�u�|	�]WTa������=��W��-���!��!�c� �5�$��o���{Ї�
�XbMNud����"���ir�X(�P�s��<X�(�]&]�!'qY�����m�q�)����A+ $y����$!����g�[���N�d�Y�}~�up��>!���*��X콐 bj{���s�J賀2�d84��t�|��!�����_v��\h�?�X�'aa+�5���?��������Ib
5�\�P-��&�� ��[����_m(<J������)�:�:�a��%�˰��U�)~$y/=>��"�46�*	��=��W��'��	�E3g�%tPZ#��T	u���J�=.���;<Cd�S�+�R'1�p"��:��x�(��_X �Dh�`��b�@�^W���D<(���rbUy�W��-�rv8V�/��d`��$~g{	%8qM�H��"��2�uѠ�W�@Q�������6t�������*���W�����R��s�MJoNA�@*�q?0;Ru	�cq)K��&������p�5�$���a7�����)pB#^�~�iQ�. C�H��,�~�C6	�[��!wEh�r��h'�zQ��'�����5���_��ᝦ��%���wB�k��x�*�i|/0�鋯R�ĉ`�Q�J��P�
2	�[��v�c��YPp�� )vj�։��� ��P��/�0�T�/�J#`��98#��3κ>U�� `�-f�Y߯lH@�'��^��� �+��uˀ�;�D���/����v�H%Vs	a+T�qV�M����!�O�J�x��$�[8��*�1c���OP�X��2������-�Wp���M�p��
>��R������1�W��Gi��}vPRa{���&��. ��b!1Pȃg�-,��յ�� �*C�`���c%�j�h5eu�=$b�R��{P>h3H�8V��!�F�X�E��O܉�,��$l�ˀ�&+{1O�?����o�`��&��U�a0B0ZxJ�鰵�L���n��s��j[�\�_�~RT����OP�-�3X,H��-[�8�>K#	��*�8)Vx��!<tI�YE���\/kX�ڕ
Ei��~Q9���P�,wC	��?p�^Y�3�K���~8T�P�	�YQ�EU����ծ��X�h$�L���Z0b�r�|h(�K��L�&�9����Ǿ`FA�k��*�%AZ_�� m[�
�(�_����\Q��2���uf*����&�ags`����Yi9�<ۋ9: �_�.[S�%���O�Bj�p����	6Tfr�Wj��PPhW�� ��yѼ� �>�� �<JQ`5�cUH@%�i�t)k�]1�l?v	yX{u ���f������m	o.1!�´��A�[:�]����'�b�U��pB�p�S/�����@�v���S"EbR&�%yoI��i�}z��u��0}�,h~H�H����t`�v�BX��`Q�l�%<�U=^�v�;h�!'We{/A�\R3�=�'��P��B���X�� ^tl;C�'z3�y2ZS� �N�����q� �40�/�XD��� n8�9![�eH��d��TaQ���)�-?��NK��$®���,E(k�)� ��_�I�M!��i�*`wbpxq��6�`��`S��b� 1��1�@�".4Ji���.7����2%���s�)p��M?�%-w���"̖0�5u"�D1��_�;��>p&W�B�����_��"t���/0�v��Hi���QѨ-|x���m�$Ph�s����d���OE��`�L׃���rrA��_h]p�V��-Zn;��)Tu�YK�D0��;w�����8�$����W~�y��|��X�ی`~��|�p�i-�.���Z�0+��A�?�\&�%���@8#d�]	�v��L&�g�@6oH���!Ԓ��k���}Q�W���K��i�� �u�}��)����{A��*�J7 ��#mL��N˒��b�_ḝ�Kj�TW��L7 �(�E��)�[��e���%&*l	L{k���;#ud��^����LO��H��U8���B�>,���K���m����RU������	�`��������>E�-��}�.hXǺw�����$�k�?�U�	H��Y^s����[��	+�� {��^i���Ҹ�U[O���J		�Z�N����)� 3�N1Ѻ�l=�F~�m�ն���2��̈P<e��5K7��"�cZ�$V�	�9 ։��PM�	� d
H�Y���d݉ۏ�_>�0�`�PX��	�Ws�Ă!-O�8 �k�������߃�L	)����ހ�0}�r� ���*��8��cH�AO I�ru1����M������C`K�NYJ1��G���0�C"�eb��QׅU���x�`^ku���ʯ�6�������~\�.��eb ��b����g]i ��P&}��F-�(�ݓx �ku��Đ����_'`��e��P�9��L���-Fs>�h�a�vv]�����v�?�	�l1���� Z�����3���<��(m<n��\��g�c��f��h�Z� @��VLj:rS7�6��:�j��z, �i���4	O���?�5`|��0\2�)%l��W	��Z���R���a�p*�����5m~N4Q驅Pj�n �f�[	�h,"L�ى�t��R"���\<)�ϰ��`w���I���>�~d�{1���g�Њ&[�	���!��|��'�4�����$���{Ձ���C�	|h�0F Xm��N����s��C-�UJMh���a���$vZ�J���9��߸7�p�\l�$�ˉ�<ƈ �Y"�j-�0�l�Bᔜ�<�и�
/��5(0>�	�*�"d�41 r�;:k�;R��+@M5l,{!�-�a~�>�c�&�� �Lx9�,Q�.g����>�=� zAc.����������a���o�r��v�3�*�[KG��S{��_����2ķR�,�<����Ʃ���A�n�N�4�P��b(� �Z
�K�5�x��,D�$��"}�6*� )��[K������S�O������x0m_�5':�2�)s�0��	%��~�pL�`�~
��0�ŀ�9s�@y��T 6	�5�4�2?-������� ����p#^)�.[� ;sg�|�:�=Ϭjª��u�UЧj��-M�r!��[��P)I��Wx�7cGh�,�P錴H2�[���c�5a���i�!�dj)�.���7���`�O^<��.+��X9�|��}[Xb)�_� V\h�Ld
�1�s+��.D$�A��&�2v`,�T��P�% DK�EVP -$��W)���	�_�n%��S���B�wݏ�3�<?A�*�# �N`9GEM�Pn�*,�(���I��Pt
��#��)��`�X� S�C��4TA�<���}�����7��B�[��� �2*0�b�p�vJ��� g2o��&�1)1R�[f��+C��Ľ��{`@�0���k�t2��(U�DjF�N���k���S���RhA�_pF�C	^���}��P�"EXUR���N̞���Ut.8;͌p��N��L���DL����L�y��fm6����S���K�⭂�|�Bb]d��/,�a�����Op�q�=�YY��`JB� ���Y������Ap*e��)2���ظ��IL'�	��4)�� �h?p���i��٠�hJF��Q��|S%�u_�F�x��\�,��ٯp��H��J躒�
�a���I�W�0���:R�{+������%�"�`A@(r���^�N<.x5GfF���{�1>���L��]�e�k(�&��X���3BQ��eO��^��>�;��[W�"Si8N^�>y$�����@/��NP֢9d�d�:8|h����� �4g��`07n \��,%=�q���.�y1�^/�4����N�,�X���q�Y�[K}��UK]��_˷�w�na��s�gu�!{��	)t�^�H^C�4"��_���3]p��[_P�Xʄ��� S��aH��1ӰQ ��z���lhd�-���hM+f�\�$����(�d݃����X�Up�I�z��o)*�_�`d��S����sP�{���ȁ4�(�X���N��()K����P(T����ꤶ��rՇr��t��j.���������
�!pb���p��0���(Ʒ�����w��*����#YK��`1���aI8B�w�ދ�Ј~�'������i;"4-e�õ����Kh��K?�z58}(SV��hck���2�n�Q9���w��+��~������U��7i^�UV��X����_���.���h#�"���I@�}~�5�:B��g���7\�U���8�8�C��W�x��,�(���h{�mJʃ	h�uD$��c� q��OKh ����,�;�8�[V�^��C�R���Jע���P=a�`�"@1�h_J�k�Vx�`f*�J�s(���[k�.`ͷ�`B�L�^)�1����PN
8=��ZE���B����(-�7�	�!u�C��/��	<pW8���`m�.c�/�U9GفP���<�9������|}	�k����^�h����6�.����t)v} �P��PmH�,Z# /)��(�J�B�_���7;�n �\is�w���WЬPMh}d}Y��ö%k�vт�/3;����W�y�x�GB��ٶvyZ[�R��dL�Fah�e{�z��+�U6��$��,��0U�������lN���1�[)�����B�]���x�jX-��S�A,�Cc������;k��G�R�պ��w*wJE�{���d�;�=�<�P�P�2$�]�0
2O��ҧ��w5���������� _�g�ٽ-�$����c)j�Ha_���w{��0Օ]�%�@����%X*NX�Qi@�߂NU��n�����]1�,�(��X[J�'�D1��ؔ�~�%��k~-Y���P��������VK��^*0.�r'�$����{�7�w.d`�5�D}Y���}���|A�x_�b����7��'ZUm\(�=*<(���l�X2�@
���fLG��J	�c�Wݤ�6�7�a�8]�X�hQw�i�ؒϿ���)�]���9&���Kq)�Yՠ隐�4�\��ӥ_`>�N�Ͼ���R��Z��4�n4�X��( 1*Z��?'� #��?�v��dO�PxR�
�n&"�w� �
�T�)"0�W� T��@����J���j�#��z��F��!v��*�\@�`cY�����;4�!��K��Xmk�P<S�?��hʺ�[�E����!{�w�0�U�ĸ�y_����V�	T|�0uР����I� .���W���~�I�`c�W��)]���X��m�Eg4bR�l���U}pf�� ��Ed1Z�6�h4IUf	`%����Z��.(J��)�dt��_a�2w��A
�PhIX��� R��s�E�	��@�F=��k�p?�E|�� ��`CM)�1z��z�ur��e�d���pPS�� �_!�)�k@
dv��X^�1|�m�`�	W؏�n-e�ۇ(�?|CH��`~��Iwo������ ��:	6,��J�ĝ$��MS^�.~���	�+h����q�X|29���B�� m2a���=\'; ��,�7Z"��b�c�@���:�1�?��X�T/���A^:��0:0Z��[5c��b�h��{`Qͬ�	�pm�{���-(��静�N�B�.��l��S�}]�`l�&�F[
�<"N����d�i	Z�`��7<o�: �X)��;�r%<Z�����,;i	�]���0)�FRy�"xY����q�ݶ� ���ǘRrLgE\��Y�ו9�(�Η�.'�,���	lA_�s�m�|^�A	�d�i฀�_�Nf��b�\I_yx�ʵ�,�/��>t�-[L�hH�V� �)=�kl'w�;�鴅� �(�
1	�Y!���1'�7[V�W��x�Q��Dmےcx�o�r� �}�j����(w��C�_x�E*5To�B�c?��Z������3?�:`?�]$|������F �K&��o6L7�h�>�?����Y�;O�ح?��?X��(�W��0��`VhN����~�{�����Y�w��1Є���	ҳ�L������_�z7��^�"{�V��W�:�j��	׼��h?C�P]`(�we�X��_�n��Q�������R=�1��~�W$<-��@�i�@PiH1^  Z:[�U��W�b�j�j�?-������l��.$L����΢���xOx����`��Z�ę>� P�ց�Q���F�65�(���p�g�����@��M��ЗU����b�3y%"�֗p�v��� #�/���~�����I BB)�q�ʵv��(�����Yl��C)Xhw7�O��@W��m��ȱ0�%R	^� ��ڝ!��~#��
�c�\��<�O�X�T�����������Mޒ�E����+d8�
��~3����68MW���ŘB��9J-5^ā��u:*ҿ��<$��$sK,ւ
���Py5_�U#�oh;b�I�
K����^���E�� VaS��1X�WJ�Y�������"Giu��O�E �FC�q�.�/�����=���9!�o ���0[�.�B�C�ӆD�~�hZYW����gw��[q�[ZPR��r�y������6�N��la R�����:�ҙ�}R��܄d �X�����	qa�U���}�ڃ�<�)�+���w9pݨ�4���v�HE�_�0��Ki_O��=�
�e��>���?O/���=���0Y�sO�S0k�g�4�c�G�O��h��u|wU���/� r��_N�G�F�%5�}~JO��1鏧[��ΰ��[�A��r�c:ZQP��
Wp�X)O�Y�9�K.k����g��k�&\�^����~�-q��%���0}�T�s�#M��I	 1a�@!�[5�.th�1��2�@�Z��B�~���[c��
E�� ތI/�ؘO&D�g�4���w�f�/�02�Y�e)�S����V���U���Y�O���@v�thy�i1�W@�E�Z�P��'J�R����UVn�p����:(��R�kz�Z� ��PD��v|���5z#���u�^�g��}�����x�k�z�>���^��I�(�V��,)��	�����J\��6�.�9�VP:���X�Ba�n�d����,�w���z}Iu��(jp���r�h"n�>]&���	kO�rW*P�h,v�fQ�M��v:�]K N�!���I��9�⟘o���;�d�r�P1�+��-sP���à�ز�u�n���g��w��`�`�z���HnaRT�)Ð��0b����6o.0QZ�t��H3x���40�$�K�
�u����(���\�7�B�X���x��A�+���tv�=��2��gp"$�	�ֽ�����Ɲ�1��� �pVv� Y(�0�R����d��K-���1���6�@)�tv�7r��Sx� DW�f=�B)}�Z���z�ˑ�c1��r�$]�	����		 (�iP���E�-������Np���0���Pm���6�ɋ��ol�P��%]��҉받� �9U,��\(7M�Ԃ>J�F@5�S��W����/���_����Z�ڒ�S��Ԯ���`�9 J�.OA�Z}e:��)H��Jqs�h��w�	���5�C(�4����4Oq����%Q֓2�:]��?��UN3\�_��[hv�Ys��(-�h\������)]�R�
�N�	��K�ˋ)������%��g%D�(�_F ���@�(0CF���.���/X'c}�����l*�c�^��T�weoK�q߅R�{��PP��b���ƚ��'b�����d1eRaj�Y@��-
Xag�D��n=<n76� �.L;J�� �U�@�>��F�M����zIn�-7���A.���k�\ �^2�Y�e�G(M�����5�Ib���Ul-3�t��v�W�7�q�J)Z� :~e o5Q-k��?�i@�O�P�Hh�-EX����R ���	1շp���N� �˳/�9��_50G0�ڪ	����"Xh�I���0�γ��������x�1��Jg�������7��­�S��[�\ ���c-��u��_�Ĉ����{�ғG�4��n�84�	eZd���T�w��~>gBpe
��=W�L0�R�eM���:ǉ�NHV���nIEW�:�א�,�2XU������(ѕPpPs���R�_0�����5�(!�1�@�)�S�F�S �Y��ڐr0��(G  ��!m�ʙ.z_
	n���!P��U-���U��-�G)p
��`0_��C�����1�XXQV�-b�c�u:ˢS�LJ��90>�ڨ%��V��������*u�YZ�A�]�Z<��8`�:B��5Nv	��W/�!т�zgR��]fD��o�0n���RTZ�L֚x-�l�)�U�����ru�}�����d���i�Qh�e�0� �|�{L�/ %_KS}�):�#��{YH@�_���-�	�E!Q��}����p��Z��A�'��*��J��ܼ�R�#��Q��~	�pUio'²�s��9O�1F+�2�h��@`i��I���u�.�9k�2H/%b�`t�:�}[LhX���2����x��p���^.�{�V���P5#���N��_�S���8y���yh�
��VD	�ZUq���A�����Z�C���8e�'��ע���� ( ����5Y�����b�����0�,�{Ƹ��:��/�|d�*���h/J6�(��%�)v�chf'�f�(3���Vq����o�h(}eL�t �YX-Ǣ�X�Ako�jɤc�&�%�jRx&�F�(�[�,��0rI�_?��C������'_��5��;�|�K )oH7fW-C�^�ĳ�M�����)��,���d5UVE�(}������K���YJ_D�`T��&0I"����>�`_�1�Z��@��c0\Z s�'b�f�_����G��PZ�m�e�Ѵ�Еèj ��J�?>Peh=R}�^�X�QD�|N�� ��/=�釘����_�|��骪��(؁ �{˓����9J�
^)� ���a����.��ę�v���y[��,O�6��������4Io��,���)���A�0ujz��|'b�[�B3X�*'�%�7��`� `�.�>;`,�^�L� ����S����%i"��!�	��`�uf� %���b��
�\����>���u�+0!����/H�%����n`T�@)& ��}��AZYhӕ�N����
��m�U�z ���B�����8�/�!Ӱ�z~�|� �� ϲ"��0�(� �h7Bn㴄�i����ICq�^�\t
x-���J�z�^u�2������	�N�__(V�>�vх��*���*
��%����d���eX!q�=�����^Y����������**�
��/̸	��Q@���[�?˯�X���A��9N)%�C��?8 m��ij����@H��'��=>�W~BAN�4D��ȇi�26��#��rJG�;P�L�U>���1@��73/-\�eLq��P�K�,-��7�[��1�� ah'����g z��ݲ���<2�^#	G�y�d�����u���L�(���;���;��-�r�n�0�!�_+Z+�������p_L�e�E��� ��'�OQ��y#�	X����(a�΀��1XR$v'�)x)��B���j��>a�{��'S�N.���p��'�|p�i!^�?���� �*s������(�ƠR�3� o�^Od��_ӹ%�$hSW`�:����0y3R�	�]no��M/�W���JB�D]����R/)��](=�ƵV; �}�UR�[��鏷@G �o��X�*��c����f����ip%�T�ΐ���� �S���a��P���/�1JHmcd ��;]5�|�@@�B%@�c��?�_���8)��-�Q���F��Ǆ�Npq� U�8W�4v����G��p�"
Q!�	�r&�_���Չʨ�g�ߒK�_^o�y�UT�e������-D��D����������I��Ly_�`���ǅ(�Ű�G�D����h�)'�(@�"-�4A.8�`�mk�p ��G��Q��Ȝ����t��E#�W�
D%I/ܗ�H_� ܸ'� 0Z�{\jh��Ua�/����|���_T�=2�.t-�a�h-��0�{�㞎�,��݋[̔%�QhE('P?׈�-�$e�T<�N���1៨���\�0N��F0�fp0OZ�_�b��C��E-%�G�C�L��4�(8:�a��	���C�b"�.�$��}��7}ɟ�����/$���1�H�?ݠ%GN�]KIu-.A� 1Y�m�'�&6ZTӯ�7�})�K�H�k*W�+!��>�eJ�����V*�1�h�=��v�R@	��~�ݨ/��2n{�`�f���[�PO�	3��M	�Y{���	�����	+^�1_F8#�$�/ ��k7XE�9��x�2�)ʮ�����J(��aP����LX��0(3C�1g\�r��*�a��@��)x�m>�B�f���,�]����.���y�a%�ǌ���P�UG��H�P� ��k�� %�69h�Z@X5�z[x9�Z�e[����*`�?��@PR��}�� 6�f����n�px]b�A��5J ~�M&!�Z��i1�*} *��T8%XWgI E/���C��1q��e���c�m*��[�Ѐ%Z��Y��u�
2;��l3*���g���l E�����I�&��
]���_I�� �E�n�k.u`��p��-!o�>�ּJ�H0�Hgԫ�Nh
z�@��üC/��pu|�v��<'xC��؇�$4�'in���o΅
Z�*L
IWhCX��?���_Ĵc��1�����38B´�0�4J��� �3���T{{�G����~���;�B�����<��� ��%)���,(�<7s0�M��	b)�\nZw�<��(�9��Ǿݐdb�O����G����-NqA�]P�1�C0TX����/K���	���q֊W	��m|l�rZ�F�����꿃���KP��6	��N�q���D#!ӱ����_�0ghU%�e�� ��6�ϕ𛰺L"�3=���AS�6	���Q��4�B��[�Aø����W`-C�Kx��6
J�4 �Y{S�}��J�%�3�(�[�8���y	�eU�e=�3��w�6�HX*Ew �-n�oF^C���"`ӹ�d� ��˘�06|"�+�`vX���0��Kr�78�����zԿf�����o�r}[��".��8{�h ��?( �<`��-3�+҉�HO�:(�B��`��Ԥ�(X�����/��Ӂ�P�O��-z�Po���6[S�_�R7(r�0��f`���S��EMp��9�ao�A�5v�V/�tD�E�'���6�GK���C7�@Z� ����t+Y�K�U.�@ܶ����_�fZF�]V�ra���v�l��k�_����1貰hH��6e�E����!�͇h~+�`�_����C��[-�v�'XU��@s(+O[����$_\��(a�d�G�S�� 
5�Y231���hgC�,"+p>�X3�T�Q�v�����0������&�a��	nc60��uA�� �Y�. ��k��Kڰ�JPB�*-�L�	4R����U�K��V!��G�K�`��NШ��!A^����ؤ)aXV�%��>\���~��:�`=�'��&�A!�Q�/�*��a�>�peqH�<!��$j���N��#PP��X�p� 4O�ŀ��(����fY-h���ָHKl-]On�S>�r'��O��B�����1��]8(`|��eXIZh��.A@ƦP��@[8�	 �:�NH1�P�8�L�S� �I�?P�f�����/% nXV5bɺ����@�q2-�!�E+ �$� �J�,1ڸBuӰ�Z�ݼ�* &�}��Gwh?́C�͘�	4���} }!���]X��N~�X����'`Ym)��[>h1�H�c ���[ ��A�i� �\)mLZ���}�~�!
J�Җ<�l���_��1�h�:�f91�,���m�0`�kG�aNM��h&d0E��b�� :��!�1���x���k�	[��4_uȠCW�[)�E��:V��%	Lw���Y5D� �U��V�_J� f��w�*5!`0~�6|E9M��ܲ^�9���T~��]�R�8(uo�^Z�����<�sf
�(G �x4�`-3s��'k�V��}������S�HN��0=� {Js���/��H���w�P� v�t������c�n^4�3�6)˄��'p�_�<R�����DO���gX	\_��/yϐ�N�1��,��('A7e���-2(B��E����+�"[���}e[��!D�W���h�2���a��XC�+��K-Ru��� ��5n�\N�)���'-��>����˯�Ktm�[�T��k��IQ�h�|�Y0���m��i�����8N�Eh	�W
��~{~�و�h�Q�.�_)��N�*R��0H�'_Үqg�?^��^�5@P��'���'�H���o�j�f��\�@|w�����P>0DT���ր΁�<
i����aP��C�XZ��fo����EHw-�8��@;�r��A0v����V�RGw9�@��B�	�J�r C=���#6�%_����a�T�&���W�[��A�X����N�I�?0�J���N���P�	�����n�몘*�m.�)h��6e� �X!Z�;���4o�Ղ���>��f��tn�r�C�0�����d�t4��A�1\+�'^T~����-X��`͹S��A��D�-UM�1Ȁ��^>*O0���+��b$�.� �?)ѵ~1@���~Q�@��dK��-�>��s���au�!
/�;H��h��!;%�	�)�d�v: q�hZ� ){�^-�C�B��@e�Qm���I�%_wdd�j
�- �_0=P��.]���z��@̅~[��w�V �3 OR���3��ԍi�qא�dz}��n�����
)�~�%ݔ(�r���+SĶ��Z {�Y_2��24�Q-��$཭��b� ����Q�b��-�8��հ�Q7�>�p�[~�.�H/MG�x�O���9�p�@s�_�C�$�s/}�e��@ �T���\j:�v+a0��4n�<R/&L�8[�?i2 �ǜ-`:d
�K��/\5��j�兤DB����S���0Hd��/21 �`��!K�f�c� ��!&�GiVp��:'�Z3�%_�� )�[�h��u�$+�(��aX@��	O�w�T(�Y��� �;����l��� p���wwf=���C�3�\hx	>���5��R��
��f�:�V�zXK7 �����_$[�������ԄZ�a��������B�<�K��%eCc��M���r�0�����F'��3}������j�I�&��!P�hQ�kI
W��{��1�i_V���|�jQ����awC��4�GY�\�����ϡ �U���Xs����
9��=ʉ~��wmQ���������k���������{1Ģ��V�k�y,z_9�(!4a,m@��Y0�v^Pyh�+Z�,X��j��;�������d�s_��b���J"�(�n�LQ� �)�Q[YSKZ�א'�Lxc-:��5e��ެgo#�� 1�xR�2���35@�@�}�.�yj�B�(v�䘙4����z����.��]�r%~��	/�,d�^%�U�����ȉ�#���h�UH*��R�����*-';�����ÑZ�3p`��Y� �O��ŀ�X����4?v�^��r�}������`��?�`J�K�r��M[�\��H�"�iᨽ�h�,�����EȢ�����%��� �	|/)������~�c����Z0��&��2P$�B��~�T��C�wa�1�]j�dE�v�N��VK�|�G`3=� ᘦ1������?�4Kp��<Cgb��'_B`����VU�ڿ=�zE?���d��n��$ �T�1�]h��?�`�Ţp0L�r;��hg#� ���(����h�V/�k�!w�B�B1��$|As�=����S#I�P�$T� �d@B��>}Lls�+~$C��q|s����)��5>J�\w$��ϔ �+[��vh[.�a ��5!O ��w����i�:�DЮ�@'-	�ʅ����tWHh{���1}���d����.��ӯ�K�X<R<o&w�y_��ل܆��W����ZU���;�&�Q�o�oVh�8�㈠ ���&h��}����������r�	TR��1ݻwq�0p�z�t T="C�'KA������Ϡ�\3[���(���o��A��/'C����a�{ G�0�\ ��$5�K��_�<�����&�	��(�]!��ZPW^bcR��X^U	�;��.�����"ƣ΃�w�$�%(oY7G��� '~\ v�rsa��ER���(T@��N{����1��>�;�%�B�}ԯ�#����$��I^�� NX�>��Qn�Ȗ"JZ�N��|D�;���{Ȑ�	�7X����X�@*� ^!�5�U	Tf��/y����q�UJ��~Z�R��X��r[������⶯!Zc���U��	�8�u��9'�wT�X�}z`|T�N=8b����k����O@�����T(�� ?MZ�JQ&��f&�,���&1h/	Xy����Ub����l��1ʷ��`��.X5t��
E�+�j�Z0� �?wJ���ve:�$W��)����"~�4����������y��RQP����X��:Y��] &S�0ds���pc� "�'���;�r��u��(qV.ZW�9�b[�㎰(�o�sG�f��OAU��D�m���%�(�>kPG�7�+u��c��[&1�oջC�3OD���(�HKL�`�ø�^%���q>�)������R='
���	��e(E��4IkU���ZO �>��)r��-���)��$�p(�V[P��&��辄���+��B���&5�6:�t��RJ�@R�� M@��l*C��ɪJhG`�OB;?�X^(������D��1��x*�U�+�]�	���{��I��-�{��{��X&��i��������\ S�xu�<� Vw���B)']bC��	gaPO�R	 �w`��=?{�akX�]� �?�*(��2,�[�hfPU�D��d3?��f`A8���_�����-X�DbY��� �
�)����ބ
������#����\��80�@�#���il8�0�W@ ��`�V�c�f U�(�������N��E躙��ϧ���v0�����Y�x[@����c=ق!�^	�`/���	�$}��Τ���r��SwG*P�n �J�k�<�vH^h.^'wnl�Bn����9����5�%�����m�N�
4�O�0J�xILWrt{�w�0�Gp-��ރ��㋒:��A���~��J�~�>�A3b�N`hM0sq&?oI��[Q�S�A���_�T����/�bI$���Х ��;Kz�\%���������s�ؼ������,�h �y����m�I��!��KcAAG�/A��6XA <��/�lM	�-+KD1���*j�m@1�@(�@�/rx��$M�L����4�,�J���7!�{�UU�8|�/���u��t'E-1��l�	:�) ��	:Rd�i'��B!�`���&�����92@R ��W�
I�6!�_r  ͍���1��b�`]��E��������gF����K_��ey�E�h�GJ��!�)�?�h��Kd��
"��'�dȰ����D�ƙ%��X�{7�v��cXV��8��Z�� �*���sL��	�(��� �$�}�h�m��!�ۀ�	��� ��0�;Q�'�1_'�h]j�Z�z ����(�r@ŏ�\y�/� ��,DN���/�Hx�pt�ED�����9@:E^�9N�Ol���-	�9R\w�$��>�Ug�����x��D���:�*O���-�$H&�=�� K,]�i����Ck�B(_&��'��x;�d5�B���++�9h&�� ��N�z����2��<����%�)����U�k¢b�ĵ�柖���n���Ø��3�c?���P~X%0I8M���	��K	^^�[h"�F	�D��a��*ao>�u������� X5�	)����y�֔��(�� YW�rlM�52�[��H]V���|(M�K(����o��'Z^��Z�ݹ�XqO��A��8-*�� ��|�E�HG
Qn��@�(p"����NWn �<X�a�&"��5�a�a1+�.��A,����v{"�{�o8. DX�D��>�J�ge �Ls�,��[*y�/Y��>r	B
���R�,�����F�28u��`ي{��s'{P���^h�J	�%�X�.��%}�}�}P����ٱ���	�h�y��)������~��y?;��WU�`L(���A-�$Yxf�[���{sW��B ���V)'���2�g/�	DXe Vh�HWt^����?���
�N��*����_m��5?�;u���ʶ�X7W�Xh6�"4ɞ̄ 5�	b���$j�}�-$4A�A���v@��+�[��Y����T w�=�񺨘�����)��Ή�{����ME��i�O��J(�G`aX,'a���ץi;B%�XZ>�v��~)� �-gcJ���%2}�(��
Z@���7?%Jр�t_��g</�#bnAz��h�:�B��a��`��?�p����~Jq����>�wP;�e���Bs}�t��[�K��O�襨 ����=?��qo�j��w�ޣe- ���ʕ��a�\���I�E�lI}І�IN�<܄�雂"��j�Ֆ+KY� T�~\!�ڼ��nj� kJ󊂭!ИYc��ѡr7:%m�c�%���l.��?dXC�2�oAA>!@�I)ِ�#wE�����,{3_���%����b�	̓�F��%��0��r�W%]g\ƿ�C�_�(�\6yJ�"Y��w^)���"	{)s�\�p�j:*�Ya��{����!��+��.�-Үb6�	fN Q�bhg���S)����ƀ�]A�9���C?��r,�����[�)}��*�bInM)Z+�+��hZ� �VN\� nRDs5�c�K��e+Kr|Y,���M{Wo�i\b8� .
i%n9>5��E�² 	�e;,o�G�	zc��6��$s{�+�#�ͱ��:-fҏd����0�\��4�(��7�4kI#�c{�6�v��^h�WT4��x�\z��ap�f����o[��n�+��LE%�]��_��Z��l�-V���+�'nI� �p����1PTzRZ<�z��Xt?���F[�z�� ,T3*��!4�@�YOW"��)��\���b[����8H��d.�dU��sÂahWԩ_)�����kTPbh�9c�țr^-���K_]����30��&J9�W!@+�0z,5�}�1�uF1 ��+F��<�-)������� S��d�-�����+pG<k١�i�x���A���?T������؉R��]�s0�nK/���h�*�^�f=���L]�+���nV,}���twDQ�&!�xA:�_9��e�:�b�-?8/)�@�X R�&iD�F�@�%\~|���w-�mt�B�� ���v��IjtM!87��vZ�_����B>!Ћ;�|$�CEO�������K;��F1�YXh�@�M�[�5B]�`���>k�~�ע"�s�(�K����@Ve�@��]~0��e	M���I�Q �~����~�e���
�>�y��O�4���	[�8�	�k p�&q��Kک��>����t��Wc�n`9fS���ؽL*6ݓ@�����y�W< L�R�q�j��o�wp�~����E zs�1���D�]6��b�u�H�|E\�����KY����!w�a�����j��8N3�_M���0v�n���铐x&Vh~	{p]#�-��l�w)��n^1�~�Y��&� ��/�1�P� '1r���~�	QUY]`���N�윓��x|Y��0�^h�HX���=���'�*#�J�K���){Z^�R�/)�`��j~锫�@�'5�Z7�2a�_��O�0-I���6he���hle�XcZ;(�-��$ �jB�N_�
�5Η���}�B�g��:��#K_�Շ��UN��F�d r�1XU� Z{	-G=)��%I��Zm%���FɕtP�ᨣo8	�<lS;��W�o_�h&Q� �	y�� L�`�����>08�N�L��LB[쳱Ͳ,��^�&_H��ӓ9\h	)�:w���x�������[P	��x�~_&��)��/C׀���]��W6h��e:�ߖ}��'~�V��[R�_{������Z\�*���D�<We�a�����˵D�3��	g8��0�zm^� �-�kS|X�� $��IvN�n,�w�+!>(	�d�W����y���kH!�C�L�.1�R��>���׬����S��k��`O�/v��1v1*��Q+�H��BHqˬ�	PY�l{E5�i�T!��hm\��]�Ճ!LHfwZ���靱����%zdD���9Jn%��F��	[��(�`#�����3�����t���$�bB �UJ �'��k�5c]���f�}oьx�(3	�h��b���ѝ@���z���iO�r�j��!�i��{��_Q�: �q���5@,�&��Kp"�.6ZA�� (P��Nf���߰^�[�fi� �+�,	�W	���G�Sz���,5�tC��Ԧ�!ݰ��l���M��0���4$Q��$
V��r�/�};��ѡ�(��c#�����D��m���wZ��Q��X��V�9��N��� ���A�o���8�� �V(�X#�+�	G�k^��}�g����6i�Pha'�4(m1Q��.�su��UV�ǁ�ͽ^+���.���ܭX�����[�ȡ�k(
�κޔ�%WQ���!��-��|A% Q��\"�-��ׂ�o~�>#F �K��w�oss�[��,�T���)�5��0�Ff���Ĩ-3� V�KH5V�9�h'�%\[X��jU�u=�k�tLc>4L�G�2�@$��\��
h}&K���4@2���Uֈ-��\���9p\O��򨱸0��h�adW����u(��ֺ�ҋ�X��l��1�����7 )�W��rM�^x�pA�C�!1_D���馬����,HMb4�����:	[�Yu!L3�V/R��)�3*.�3a{}pc��� �ܚ؋�%���l,���k/�Ļ�"Vn�c2�? s��)߹�>$@�@�+A� |�Kv�`|�u�	~��`��3Ԫ
�O�� -7*�?1-�)�b���Ϙ�[��5�"��
�����.�V���9.�5dq��V�i������կ9$���R�fa|:�v�JY6�2����}�҆?��¡�Jp��d��+�O��0W�q] -��C�W\9��� �]��U�_�v��:1Һ�۾-n��[����hPn�����6�!����?	��Iaʡ"�`���V�g�vk@���S'�0���wXF�/8�1���a ��"~�pu�'����z%O�����n�p/\F�W���s&2K]�����Ɯw���Ol�wz��i1����R������w�e<����c��;�|�ZN���H�0%��$�;�%U�#6w.0"(ƀVtR%���mB�䂣0���yL, J�!*�_)�1؁M+^>(�뀕�)q��g���*w ��H@Q�:y	�)ȅ��[���6_��]�[A�@V�(P)�$�1@���h_?R���]���N$鿼� "�,&��'���1��:''�f�٢���[���V��J�}�0S��Ѝ�9r[ۅS�\�M>�/�V.�X�r�S'Y�� O�%j��-��^��\�v�,��/�3H�'>��%��ӱ%�n�k�y���5 -���=)� �u�1�Q���UiM��Hޖ üS�i�;�r�d�Z��xkS�"�i�J��:м�O=1�r�TX��'��Į����!�0��������-5��(�-�<�!��T���FXwJ�u7��`\��|�D�H����~�AhUp:�u!�z���7c�fZ��,����B5C��!�])�f�Cyu:1Z��H�`�N�-
2\u�%�v�����y�����ޤ��D��P��n��L�u��t�K 7�3�}�p"�XZ��H� ��Z�4��5�#� %�o�A3M*؀V��M� g-"EZ@� �=e�a3��]	P[���#S���>�H�R�Ֆ5�2Y ��7�5����WM�������Ta�:c@��It?=)�K�����n�=�S�Q����KW��S	D���L]���J�	1����������(2��vUYR�^��{K��鲅�2x�� Y���Z�7-�2gN?�XA�c�[����2��'�@���/u�m'��	�_�H���j �#��X��h�K3�mzؽ�X��e�)u��������{a�*1�R}Fhr�ˎ[fK��G1 ��hyq}-��V�.��pA�d��+5~����J 8>�	\BW���IR�����uB������,�H��&�{/�iUĜ(u�4���xU�s�.9a68�q8�&'��,{�F��&�(���O�Xk�W��%!�]�͟ �<=j1��'N�l��\$k?u�ju(0/`��hZ-zX�3�)�#<�-}1&�Ѿ �5ZV�L��tS�A��\RVh'.y)N^����ѯ��Zr� <m�оy9K �@�3�*���O����l�M��A
��q�VS�pp��$�8�B¿[�0�������������v����`ron�*�+�1��1�0_�E0��M�"}ep���<u�&B����+`��b<' K��#PZF:�-E����%�����w��yǭ���6�����w�͘`����M���u[�ʓv,.
����h�%Z�L'8�����1�0�F�G�S�oE&�؉� 5N�c����Y�&��t����B�0�A*���) ��X��_L�%(�h?4����G���K��<��$x���*n^�P�O��-� "v�I�K��߽$fh�G�c!<�����K]�#K֠�M�����)_��t��н�J!�]?	��JX˟o֟WtF�"�h�2U6�������'w�p6����q:��8�ho_S2-)\>���(�1��ӑ
Y)�z,n��Hj���Xp�q�X�C�m��%�P���ܒ��9m/�|F-�wءJ���0|&�`%�iu��Q.ңYtI����%s��p"��0k,�	�ԇK�yh8�<$x�Y��ѿ���{3b˼P�6C54���k��W���V���_�/�^��n�w�9a@'xj�	�!=�U��AM�E���`���V��� 1����P]��W:`�X�瀁�� �Pǰ|e� y-�}�"�2���WRp�����	�������R&[Pa��!*V1a��S��B'�M��@�^+ /�ox���W�g>�9�|!;�B���QB���|kC�Y���9�l��!z�F��0�mF'�3�cU�f*�	
;�}ē;� F4�����E� l� �;���d'�~�̠Z�Bj;�˺�Ͻ@O�L0�V�qx@\X|FK�kQCB&*9)ֻ�Fh*�1�'B�`�4:�(�%㩍1� �5�I�Q��A�yĔ�_ h�lf"�����J| !IjM�c{Nz�4i,��HW��V�^�-��uX�J[�`��@�����Ԏ�\ �����q�wA�0��hi4`��+�(;,¤�m�Z����+��tNy���G'B$!�� �h�� kz��<�^H�+�a�pD%Nw���M��k	�O`��o�T���p	�W��}���*�:��`��Rd�	+���������[àFhMB�J�)�.�\��աXh�i�|@�b<�D%O���?6)�w�9"�#���P�C�1�龊�8�'�Y*��A
~ұ���Xh�K	̣�,�
�N�M+��62"Dtr�����h!+���"	�1��@��G_}��ϻ"%�I�a�n�/�t��́�Pn��l�udk5�K@���(�Y�X��F�/�� A�-Nr���a��h�^�]t{Y���[a�y�a�(�*�M�U~M�0f���Q�!nF��~.?��6jfs:/)�y�kT?�B�a_I*��A��ّ�K�@���';�e��1a0iɣ�������)�6h��M��� ��Y�)�01��a|	h6��_=�#�X&�zt����%{������v�X=�O��	0O����F�[��)X��$�`V��0��k%��*��pF�U�	�]a��/NcA}�����A�^��KJ�� �`[�{��^�����JlP`�� h8V�5��'�1�Z��
�[�������� ]gm�oB�r7il�~/�v�R^9�0��p �y�z�]��������|%���D 5Ok�+��G��"T�_u��~��,%�h:�M���A �U��W_#��P��0x.`d����K��ݹCZ��1��-KH�l�	�@)����dj� �za`�9�er�VM|�c��0z[��i����k�V8�0�%�Ϻ�u�t�%�\	&JU���D�N��x6�K�h	�# /qC�z�p��:	�Py?�{���	� �r�oXF����l��K��_)�-�#�~޺�8_)�jK��wǰa���C�X@�d�0�5"��1��`z��YH|sN�@�Y��xմ衒��KT�� W��DRh.Ek�?�f��Y��V����2���6M�4�_{ 3�2X�y;\+�쳠~��sѿkt�Q�l���Z�~�fR��$�&���9y?)����'%wUqR)��r:��[:�b�L��@A�^�)�UAv]8�-P�+�6Q���j������rnW1�V9���p��%�l�S� ����I�OB ^�1�o���Ok����;`��
.�_Y�~�yU��<�~��ҋ�tIX��� �d<�L�&�%�i"��>����v�Z���qY�M) X^�%R}`��N�qK��P���}N.Mi�DXp�$��3�߆ShQ�Ԑ�09B��N#���}���\o��4̶>�؂G��W�51:��R7�S�&�Z%U4�i���_#��At!�>h|�F.]�,O�g:��_>UT�7�>=h�W�*���@(#A��\h�4�k��Tf# �H�ҵw��gz
c��̠[���~
�V���`�>0�Z��z�M�W�iWn���6�f ���)(�V�]��v��+�3��?d-H,�P��H�k='L���~O.>��G�R�wa�78M<�+���l�j�E@ ��5蛑X�xN�5�!��:��8V��u7�ߐBm^�đ�THg��q]o=@�v3"@H踡�)��/ݚ���!�ޯx�Qit}G2���rg0�0�� JS+�*mQ@�(	nw�dx�2�b�� �+	J��-�%��߀��90�F�y]�(0�S"O6�;�J��H�.��,�\,7E��6�1 ����^�����S�( P	���-�$�&a��_�^���˂VWhFT5`�C�I��D�zQ�|{�&8	y{��=�TM�.�;Z-�4�,���.���S'	|�6%[:�Xl������hi_���d �D_���.kc{����K_�x��)��� s�h0&&k]�O������tY�`�h6'EJ`4�[]H�"KYe�#����˻�g��~s���}!))�s(��B��95��o.$]D	_�)M �]I��_EP	�*�.��fZh��kBߴw��!�;
K_�kh�����}�&S�]E�8�9�/H[S~�CO��1-���}�w�#d�8V�4!�[���w�C�@��\⬱Y� �1H�aN��-^������ ��E���LD,౻~�߰�]+�ٔ�Hi�SH:�2�����'�Z~�-����[����L@%�m�8C�H`$)�[1�5�\��-�VG@�(�#�Qր��xT��E����{�&g^�I�P��{��q@���*lN�X�F�F�Q8j
����� ����4���{�%F��L��-���J懟eɦX�H�-L)�7Q�:1Z���o �z^�;�W.b�[Y���{�sf'¤�h�h�~+��Q�� *���vx	���,������5�t��Y{{L�� ����)���|*hW�w�HL
c�_�]��/������-ib.�Vi�p!�6&d)&�,
J e�e'�e�dؿ���+�E'7�����'�!�/�i��tO��Ϙ[:,0M���I��+�X&�2�UnO!ٺ-�*��I��\�lb �������{�L�(�V8�xu%|���kv��s����hP�ǌO�z	�KCx�^[xމ��k�_�,��>��X%	+K_�Y���m?�$A�Ap.a�BP���e���Mhz+4>�:��}��@m��Pm`��B&Qa]��tEy�0T���1�/�)��D�ަ�vP��P��Q�g�6�?O_I�P�}L���by���RT�@����9�?��+qaa��D�:vBN��<.�@�X5Cw6KZU�*���Mpɼ�������S�R~�`��D���8h�XS_JV���ׁ���G�S�C=�X�p��3	h�t|�rsBZ@�����WTs�����e�2	��٠<6'�( ���J�oh�D'W,�ԋA�E0HTP_��L����1�ǀP�^-�(P	������]Pƭ�٬C��N�����i�p��Ԡ��-"r�)�*(?�A�Pk��'؋(X-�����׺N�R�^����?=7/)^�y�j2ם]ބ|�3%������.	X���^h`R%�:Z@9�0��_C����vG���*��LE?}˿'�WN�Yv���/�@b�Pn��/��Q��w�c�K��wBWt��V��V��F��f�p����z"ԳL���)���&3C	G鯔 ��w5�Q;�o�I�tYcU��4@|��i�ڽ��}� ��E�tu?$ ��m+@-\p(H��A��b��غ	�D�%Z�e�~��?<2��*x����`tP������b p�5�}�.{��b*7�K�g=���c�)����J!1� h�O��'����fCۛ�xہ�.����f�
�2��f��o����f@���F�S	ft�LB�
��&`_%��Y�> �sA�_ȸ銟'�r�`͹M%Y3<D`����|_|L�<��>��AL��ud%�2��^��!�ҐP^1�����	e
���� P�-jK,�x	*V�O�f���P��Y�ZCW}�/�p:\�o^�g�U��i{0�3����_Y�C�%CA��"��h�k+��a$y!�[����gw�Y��}��x�5��t�L HMKS��2��(����? �L��x^#T�	;�t�[!r@�g3i=9��*j��O
�PF��2?>�R��)�Z"��#�y�H�%vET�<J=�3���6U�U�����'�B�ne�ros�C<�1���[��c���<vNs��*�0�
�p��GeKB9��R����h�	��ݤ�PC�� �jp!�5Q;3�C,��B|� �R�YI:���:�˫��4��K �F��� �}GC�$,p%�m�aTB-_9�'�Z^�zh�Ъ��( ���G~M���HҼ@�Jk�.��OaE|`�qx7�8��
��JX(�)����'x���M^?��C'���e��{�2��6�d�������͐�9!�`e��A��:�^�Ԧ&������G Wh}j�#O�;�A2�BL܋��`o�<�v?��4+�l�2���()��?v9$s�}N�a���1��K`�<�	b�G��v� $$1��fP�N鍼�'@ V����Q/����K��);�42�+M���h`C	���}�V)�2�Y�0ވ����@{��4��`��0�?���4��gp�
i�����9?��-)�u�kT��#d KVh "7)���ew �3�	/�ع܋�S�)p.zD wO�~�尺�>F�qѴ��^�0Q�̀��������:�������]�o������H��'��Bj��\��PlTix��(��*QIA�+�H���$�e�!7��1q��zK%�~�%SK�q��a��@�-��=���t�a������b%�փ�ԫ�����,���׫��(�YGo0�����4�<Z��/B,�n/�`�.-}��6	dm�_ U{�f�\;�Z�
���H߯��y "�;Lk��N	��^6���w�����L�@��r!R1�5ad�eE�S�`z�j�Q��L��,_�p�Z$֊O������B��x��Ɛw�3a��u`�|@��hd;��kH�,9,ht!��d6�j�8�^gPD1�����xN�k�D���phW-��?�n��!�&b�<颡����`�Q��݅���:��t�	��Xq`�Te�k��A�Y��X�Z��������\H��_�D�x+������ԮpX��9��2�j&��i0wu��:�*��PC'}�����MH�am,��ƀċ
�[��8������ �gQbv��U�0}�"�]��
�w���q+e(�M� �h'�Q�:�n��!2���20�k�(*Қ�����"��p�%����Nn.�o�k4������>�qC����~�����1�\���׀�u�-�yI,_반����P%��0XD����!R՟k��(�4^9�XS
v(,�R>W�)KT��tp �>���]@�	<z!�wrU�j��1��b���Ԅ磲@׭2�`.+�TK��^�1�L��UJ) �,�q�1�pQ����?�@�v0Q_)�!U�d�=4�����SB�����@��V�ƣ.ć�(�tQ��h�L�v����4f�nW���C��FOb�8�¼�J��M�V�tZ,�c���/(U�V"(�(���c���_��ߝ�.0��Z�	�� �Ղ���t�ok��a ��*�a��eF ��Ey4י`��GL��>Z�(o��c(Y�,=%�H�<s�?�N
s��*.z���OK���!wh��a$c6O�K��8,&fsA �w�PK�%^2WH^:/�TX9)��'�D1�B�w�y(( nf�l�h�J"�@��=M[�)�:	U	��V�; R�X�$,wq{�@�Z5�Y�_F�zS����-�V����(	z����8�95������cPg��2��f�'bV�وm��>�����(��̉�7-���Y���&4+0��+H['@Yh�}7�O��s��?����)#E�vª�c1j�P�q832s����!��FFܚ�]=�Z��M�y -�xa����$X�R��~���q)��ZM ݾ�Xa�	�6��.�ꢸY_�=.���	�U��9�͆���
d��4 �=�nB�;]}��E��_�X`	�R�,���e���C��p!�-7��%�mt| '������]:����P�0-���v2u��|Bf,^��<���5{1��[R^���rq
�y�*=#LN���|�81ӝxR�� �O�r��5X(�h�JB��nA�5�z�9h[v�w,�{E[1�Q��!}0�i��W�`�u�g���];FQB��L�T�k���ޭ\���x�f���o�Z��-��T�	|..X��������˟`WVėrO	^	�S��h".�_P�)w���-9z�?�\���/_�vXst�}GD<z�Z� "[fPS�J )�$�4v�HO�4��7Tf��N�G���r�sw�3��`����/;�^|%t ���N�`1�v��$)˯�u3����	�<�e��?�!��px!�H�b��.s���R��o_�?`��(�}�+#R� �Z�fF� ��"Q���ĸ��^�y�Ѓ���Y��.�[�g�:�1s�0IB.��X)9�~N�d�Ӹ�3[(�ᛇ~��9����$T^s)���o���jO���fG+!K0K������0?tj?���.�_5�#7�@����W1�l%����凞�*��%�<b#�����GO�K������dt`|�S����B��[�Ɵ��v(�0
�� ؑ�N�� �񷨀%���R�W�W/<iWj��;�a��ZTYϩ%�)/YR	t_���2`�R�t,�x�k�)�X�u%���8!��Z�*`����� �bv}=��A�
%X?����߃��5f��@p}�#[?��J�I{�h����'T�-�8 Z:%{�%���QZ
H5kj^��{��$��	��| a��΀�@5X�^�胎��yZ�ʫ\XW��8d^�lA� ���3&�	y N�"�H&�J�U#�X�F�!���/T�� �2d)���CmE��"x �O5H�/Й�����M�0���U �g�0-�1zϐ�%j��ʧiF�4��­f�k�]�E����(����&�VR[hU^��Z�m�������Ƨ0�fZ �'��,��d���]I�0ߒ������M*�B�8�S���0c���;�/)�`�LS C�3�;��z��i2g�Q]t`�����'SO�:�@�-'	�V�`w'���Z�RB�	��9��+HZ۸�͗�� C�ʪV�;&J���e8q��=u(�ȟQ(��RB�{w�OVc!�������@�W�	)f:T=��7���ԉ������!Oտ)�;��F��N&L�|C2*vI�_)q	c ���ek$;J#�l�,�����X��ѶP~��T(?_�I��V��!� ^U�q�?)����x��*�m�Zʺp��&j/wq`ttÕ]����
j�	g�߫} ��ˉհ�J4K5j�o -���������z�p�>u%-�l����_�j�F�kh.Q[�z��1�xR\��%$]g?��ZG _߽����G�P���ϡ��*�Y���(l�����GП�  �(�h�;�[y���@N/k���S�,V ��F�Q1��7��h�s�8��.3�=��E^M�`��1I<��,�0�*�ϽH�^H�X�$1^9г��?x@`ӽ�af������X��Hr�@ �n7Z!���,x��a�X�;N�@�v���� ����E��EO�9qy��s�!���h��2�j����:~0$���k��OY�ɲ6AU���a��;[ Q��kB������3�_?y�v e+�i)�-SmTa$ZzxN�������_�?1
0�< �,���� �C|I��[����g�i�B9�Q'U���� y%!����]k5Ô���5�r�d����~��łKts`���L� ��M2�f�
)���'�]m6�f��z/�- �	�X��p�!��>����k�H���z�q���z$�&�6��,��KE��@�G���P�y3���_�WvP���{�@��h����U���}F��wb�u���N`')�T=Zx�^I��]RhN5,	H*)�b����� ��˦��bh��/-D:�u3�	)�G�OB�0^\,B�`���%��W����V;��vK�ƴ���*�� �|V4mM��Pj���b%�Dl���(����1*�]�0�X����j�H���߀�f(��
µ��d���7;K�`�^&"���r�dSH�y�`ph�[u%N��O� �(@Bs��2`�Cn�VR��,�9-���8ep�����^0M�8.Av�AI@�^Tj���'2A��a��1t<���oQ'�<��%M�Dh�p�JӨ�O�F�]Ubqb�E����yW�=!�/�]�|��_��LPQ�7� 0��{.,^S-��	����t�%�v-�дH!� �1�R��r0.Iy,OKM'��'l����^� nW��s�	�K!������J��0)��u�b��� ����/�� /P��}�*�^��3L:��?�N ��[0��]/�v�a��`���T�0?�W�Zwp�[��]�����|b�X�vӝ��i�~n��� ���R��GT�&(���N?�)�����{���\NэhX��3)Y��p( ����k�
�e��o����'���_���-�<&?hnF=���j�y�S����AQ�D�:		M�O3K}�o���t�дT���<T�N�Dz�{yL����rn�a�үzt�Ph�?[�����2����� �Mir)���W�+����_٣k���ֻ�	�H%�S� 5&�]�%��}o�hS �.	��u='�n!A�k�����z���Z�%M�ͰJ0D5t_BN���	 ��S��p��w�N%tP�SK��4��� �5 Nzx��� ��eZ&j�Bd�!gd4�s��
�;�[��۽K�G��WNe#���K����<|���ٯ��𒢌]��D/�µBZ��.	�K0���� �˵�(�����.�ͩ2�Ż���ݿ�F c!��]rq��-B�1��?/X�'s��R����8�hF�n�q�&�p�rp�.�����O�>�J"�������s�8pa����L��F�̘�{�)��7%U��3h'<+��5o2fBǅ8��V3)��W�R}Q�E��5	RZ0ta	"�\Oc�;�b��	lfh�x	UZ ��!\:ss);��%~K��L���a�@�W����LT��H����������W�y,��R)�V&M �Q�b�� �����PQXY��-��;!ń�@#B䗙Zy�Rh6i�~]�ږ$��I�_�C(��h�*�uP�'����y��'�3W|�����R�V�9`p�4g�TH*�	�{��Q�}y��)%l�곶�`J��cϲ�����'��}�aa7T��y9>9���?��!�$�
q��9�+�ڡ*Ȭ"+���a���w'_��Qh	�l�O�ej�{�A��z�wvD"���Uͥ�����/vyj�*�@����R�����D�#��Kl`V�+]u�)Z����>5�cfP�1A_H�Z����%�J��G  ��������9����0���o �Rj���Y%~��T���� �Ct.B�Xh
]�	Oj����/ ���g�O� ��d��7o$D��{(n���>����(C2��1��([R*�h)����i����5n����Nvd@R�s��t#4��D�J�W���P	�b1�2�I�Ot-�o�r_����ꢂ )Z�k�N�?,-#T"O�Gȓ�w:4]�5��h�k܅X�+e�
!���_M�h�P����WR��&����Ԁ������
y�<�S#��>��#��:?t˼%�ީ��l�>3���{��1*�װ���ƍ{m%>�D>=��S�&]��4� >)]�6�ʛg|_�~{i�#Q�hCڡ�'Ir��	}���G��l�����=&cM<hrV��)qkx��-r��⥐6�X�_	 �h�z�L��e`Hd�X��}��%[E���B������
�T���@u�Z,y+9�\�Llr�4�r	O(�1L5�%�0(�Q��&*K�����w2���׫��\W�B@��'H�-Xd�pE�O��ȇY��V�T�?����d�bX��}��<���]��는��*#QPj	S�?)bs%un@�zM�H�� H�"dF!�] �=�,��ZE��pu@G1ʓ�vxX�mzN���0����&�k[qg9��Q��z��aD᡾>�IhO]�g�9�fl�ݫNN	pr� Yt�!�4[��Ϯ��������wG+g�0wQ��0�Y �N�墈�&E�%����3��_�;N6�"%Yު�'I�
~R-�YX�㡱���aVx$�j`���i7xzU�[�0'�,-�(�O/�Fa�ADB�UP,=�׉!L�^��W��?(�_��.���hUE0ŊN�ߤ�@���n���u�l{�1�%Y���ʗ(!��#(q�u�]2ߍ�[W����]����80÷(�i�_v	���.;�t8��6�$<�n��	�^�.rc�)��LNC	�3:8e7_����IO�	N
�lL��9�H\dJ(|���!�����?����~���-�ňO��)V>��0�R�F<���-�{�Ǯ7ĝ�Dyz�R p�T% !�ʍ"P��-X{;��Hu���������(p�t�L���ժPU� @`�MZ�� �T�7G.�ה;%Q6p�>�݀H)ͽ�0:*�x�p1�(�;��(��K�_6�q�o���T��>��	\�����B�Vg�ݼ0F3���M�����Y�����0��v\�Q]���$H���}(����� kZ��zf�|�%}qf?�����W �A9����J��شe	
��)�}���[�0J�:�
`b�L?(���8]zH�~Ǎ�3l]m��q�A��"-R2�'��h�\�f�U	麮�w��v�#0H��`V��Mc�hs(W�i�#��JS��xZ&.���ϱp)i�>�@�|;S�e'"_�@�2= �x�ƻ	&N<�(���+ƿ�V�t�7��!a��P��dB��6hx.��F�Hfe%/#b�.��KU��qP�����y�_�A{�C1�1A�!�idz|��� ���.)�e:d�R��b�W�/�N�����5�B?�P](���{Ea3���~����Ͼ�!V��͛z���!E�G��p��E�f���Z,��&0B
�����f�汎!�R&/�߲�`��l%�v(�/��T�Qh���H,C���Um8-݄2&��,��1@_Y�쏃:P�	�=)��?Ν@�IJ��FU�+�D�l�*��K���Wܭ�E8�i9(�	.s�
R��e�(��^R�ӱ��u��w7(��!V��=	鞈��`��^m�"^S�Ytwh;���,����߄��,�}�i����v�c!�_/�!֬�ojvP���@��N[��g�%��T�Z���E�˕J�
׮���1��,��8f1�]8v{���N%��V\fQ���B:����s�0�����&E?�,^��[�@�y����B�5�φJ�k���^��1#��kg�'�ۘ��9iu ��{�� �M���=3���X&�Ru j�U�ߐ�.�(�R 5����\r`-�U,F� %�0�Ҍ� >1[�[�5���~X02����Goc�wwq70֏���I2�%<�u�F�
߃J0��[�'������#�]��V���[&04�9��+�p+X����LWsX�3�C�4+�)���G�~������<z�4>�X^h�:�I���f�%.J� �
i\�j� �Ed,nA�#��1�/?�f�(���hC-�1w/���і$3O��ݐ���aR<�1��]�sWq�iAO�?+�i̞{�KS�� ^Q��1k,�N��)��ذ��މ�p�A/�f�!�=S~�Ғ��n��0+�9�'K��F���,���at��l��:n%u�[��Ǌ��4�y�����Е�A�$$�dwY�3pډ0��E����R��$��1YW� ~7�]&.����L f5�v<Nu��O�7�X-�e�Om��9M
�fZ��19:�3�;��4Ն��.�|X�{%vѶ�PW��H@�r��(��R}��vma�{�H���[��U�dF'���ÿͼJ}��O^&�b!����+�i��8kZ����^�-8~�i��
Y��%N��d�ο�{�	PL&.�Xy����G�i��J�<�Ϊ!6��H~��IT�¼�w��њY�:�G�0�Mq����%Wy�rx�5�����������	JKN���]�����z�R0'�2�l5	��Sh�K_��gc�	]��4 ��?&=���W�r �jIչ"2�9鸉P�
�k�$)JU�{^��G� "����uQ�= -TDRH�����ȝ��%ה>�&$p���/^X��Y�f�m���K���d߶)�U��������� �Y�����;v@�=�����Z)sE4}���/��iX@��+2�t���B%�i~u�, ��)ΐYkJ(U�N ��[�><���^(��;�*����
�[�h%�L�C
~�P�D�Gs�%XD������ 3u]�8�`��N��x���Y���D۪�C�ҽgG�6M�q�:�Z�FƆ�� ��'�y��	ea�  rk��]7�˙P}`�&t���i�rk�0�)��VJ��:�U��@�.%F_d!-!��[7p	�e`B�_�����8�R���X�	g:~ j	p4�/ֈXY�w�1�S��6_���FefHz	:'	�BU�|�aÊ�3�'�%� ���'qZ�n9@�~8��"��LC������1�Zz��OUx=
m	�Y!�	�tGD�,����\ �9�W�����f`Th"(���?:wP�Y%�|,���T����%����r�Sܧ�8˝sF�}���e��X��{e��|5�*�2���	Q��V�p:�Z�X5"��!�n��aɠЕ�y/��'�^Ԁ�S h/�|b��b��A�v�}��_;������#j����P+�/�il"Mp�F�n����i;��c�ۤq��R��4b�~��j�����}I7/��!(w-�|��X��N��4��#n��~c�&K	�!?B<�� ��a��� G@�:�ZI�yp�`B��M4�c���2�;dBD�h/�I��Xm��U��/��V3!�h��ֿ���'��6��N0��@/I�ebMxǊ��/� I�F���m1N�:��Y��I[&�^Aį���K�(������-LD�~;�����6��b�	Ds wND�̭.�e��������AO�z���D(�i�\U2v8�!�?�w���0�H(����u�@��	A&
.��\T��\)k0�d|�_J��X������
�x��;hI'�N/��[p�.	��z�8�0�f$�N)��m�:X�ML|�'1��h~�Œ�,���ВX]_�E~Q�&���R�8X1�O`A8�c�6��P~�_w]0a��Q<(��	Z�݇�.$([����K-6V�c�,�!	=X�r£������&���Q�\�[�ih)K��&�"���5z�) ��+i�P-1X؛���T�KV�dE�R��`y�Kp�[�� t.o6)�1� �_h�?-s[��I� �)�1���PV�]��z� �)N��:3V�'�Ȧ�J�P]���m6���c�X���E^	4J��u��طK�ּMӪ � ��25QKt����|�3X!�U�K�j@����vۯ�4�����Zp*��	O*�h�Xir����>���=��Y1�6u?ׄ�3Z�)B'1����s.��%���r^���1�X;�ӫ Vn!�E�1��Fh������^?���h���~/�:�I	�Ee� � �h�Bk,Y���E:*wU@!?S@��A��m,���+�� @H-��L^�R n�SZB$�K-�e� ��U�h%EJ��]��*�%�L�b2�lO� ˥�g��H���	�/։O�!*J[�B3W�f��a���ϗ�-��������^�W%<d�'MeGl��u!O���#�OP>Ȑ)��mc�&���,}Hj=���)���H������O�'Y��&P���'-ЄZ�	��^ܼ@�ag�/@z�
um�p��|��5� 83[h�&�������*!}�Q���lx��� �]
�P��2T1�\����le�*�Q�⃀'�%n%ku�i8+��Z�\b iH��
�=��L����9p&_D�41Y�
�kI�0j��m{�j ?����H/]@��^�t��?!b�K�BPT�`N�t������J0���z�B�����,P����[�f�w?�9�J�h�>�d �}'PZ�|O�1��"�',��p������I/?t����[�*m ��MP0�H�1�)� 
wXt��@Zh�2����ig�
�ȉ���ˡ�^����f�� v�^8�����a��-��~���~�/�L	Jv�XK=�;��D�1\mK�#*�'C@U��sd��);���G�\����ڑ�s�����ĽQ�aA��
16��z�����ZZW�pJ�F�ּ���PN���`SZ-�P��1�U��.��%������`=K��$�;B*8��[�uj~�5���Ql��-w��s6�NJ��h*oOͩ�X�l
 Rd0�P&��� O-Cs��`6��2YKZ���O)#=�ݯ.
��*��	�{ʅ��?}� 6r:�'X@5�0�8�,\��.����f1��-l$t2�;Qa��W0��?��hOi��e�G�O��G䋜���yI���e��8!~���P�� ��i�\���R67��@&.�N�H�UN�i�"�Eo���h�( ����h�X$�n*�}@�hw�子)_!=����"��.���y���ܳ]R���.�������Za�@*i�&q!�$'<0�B�4��3@��}�1o*([����Pu)ݠ��_�O;@w ܓ��S��Y�S��P.�聍u�a��WE��������Y��_ɰ�ŕ�
��,MR~���I(�ذ;	 �9>T���nS�XO��	�N�q'|�@��Q�Z%�+�J",�Tͱ	wgM���;'�oXc��,�R)�<�@�
�*�LAdڽ�9��tyn]a���n�CZt �" pQ�������tK����o�́�F�o`��R8��(Yė�39xŌ)п /(�%�d'1�]�j`�-�X�΂W�5e�\��_�K �A�v��q	�,w�,0��6��%��Gv���[
d)���$"_��LY���>���AG��Ń�����.1/�)V�>��p��DPy�HV�h<(�0}�Z�U��ktr�hwN�@AuKxV�R0[3$'�*�|�N�fy�v��Q�Jo	ܐhY6 �m@ R�]�[��\�[�m3<��]�FG�ħG�x����HS&�\	~���;ג�Q.qZ��*9�W�%(N}�����.�PJE�I*+����o�U^D�|�o�O�:�/��E�������W�vg6�W`i��h�J#���tcxOپ,�([X�^����ʬ��h��ӀR�Fg�u�n��	Nի�N� 9�)W�`Z��h�P�aYV^�L�b�L��0��jd-Y(XWA�+;�D�$f������ ��������|�)��6�
�C�NY��X5GP�)o:����S���N��)d*4NƱ<�~
,�&73���}' .Y�/Pd�Ph�>]g���:/or�p��G?T
��3�~a�.�*�j#�ZL�e��>�ZI�`���޵ZuKFR[�=��)���Q%ץV�;�jh��+$�BOC�yު�-�
�^8b1���a;N��z�����3AW}g���Y�^}[�ƿ��E�8KeSB�x����绻�͔�{�tL�]w��2|��u�$Y_�,9�B�yl���>�a 	�vq �
x*/V��1�$'���8�Zv��hM��J�t�:K�:���M�"�&	�m�<nB�\�a�ʓ$i�Su%MfKPOPЫ#x~[}��������~!�N`���8�:�ӓd�	F骊� �."�@���	��B�S��K����%�`�fQR�6�ⵝ���Z.�I � \�4�%�Ǟɼ*�I�L��`��:(O ����Q�AiXw�>,}'=B��!���m�!���h�!���A�[�]���؛i�>���[�41��h����7����޺t��Y����^� װ\�Z7�X_p�s��� 2y!�-�[��Q��!����K�u�-�gӦ�_�Z��U^��\~�b��$�Y~�';1W��A�@��^��`�*����~ Q��k	�_P��뱡�����is�0"����0�됞�� ٗ� ��:S���t#-��h���%��W��!7�_�m݀�|<f9�F)�Y	��>k�l��̒v'�3��r��d@�'�%�Z��t�5�B���E�醠`I�7n(�'K���!�hZ��fk���JD[��Ӽx� 1�|x��JԲ���	j
�>�����/��`|mT,d�oȇ���	:��Q�n�]���M��d�#�*S9^[� `Ȋc{��BX-�[P��[�(�@5�?Ut8<�/A��H?H����<��h��5�4~��%�ט��? q��I�� ����HfBA3��)��`a��#�v��� 1ڻ,?i�MC��Sj����&���x�ٮ*��!B�J��P���f6I~Z$��@�E;�;������{��ev���{Z@��=9'�g|�(y�s�\��H�[/,��$�s�-X��y2b'�_�fW�t�[ n�v?n�m���NP댔�0��IXװ��3�4�s-Ua�"��X�]|�O���h�J�>�F�0UB$`Kf�O��P�	�SW[����Z ��R�HS��f����#)10��� �RD�����?���=v�f�נ����>�l��%J��o�^D����R��Uͱ鏂��h[H��Њ�9�>�J�p8���`P��)O���(��pǄ黊�}瓑�����o��������R���JZ�_���#4(	1<��F��ˠS�P����X�����И��_�^#X�B'�9q��h>@�[�� 	W��Ž��>�o��=�-��d" �XH�Uy�תՉ��/ �˸#w(^>�q`[
ǶiK��#�����<娤N�D�O�U5�Y�s 1�-k�r�_��t�� �;d-2�$0��wx]�o^�S̉� <2O�3^��ׁQ���y�;�Y1��f���9+�!D-p���N邶򆛎���W�D��f
(o �<v�&q�D ��9�\V�g
�4�t��w0z!�^M:��T)�Y�-]���1АC�_x-5IL|!� ,	���\�^�p�x׎�B�B�UT|�HX1���QU�oR��X �栻�/ Nw��!m�v��l���r�wh��+�Ah�xP�N���k�X�����^1*Z�%����5c-�YA�9k;�b�[���aJc��h?����%g�A �qL�Kt��(@'�_�c��(�K�O\�_����{�-M�,#���8Wcv���HY�� ��MS:h QN]����@aZi3�z9����Ã�� ��=��0���̂O��̩N�h�k����D�O�\>,��J�C�����	��Fx�-�Z x���>�h,��@��-h��|�Z@���J�@r�"/|��cC(Zh�j��&�����p�V�ܐ큍|�)+��-���A���L h�D]���Mn��H�E���l!�P.�x�տNn�F�d)��P�ʷ�����
��}���JWͮ.�N�j�{QO2�"�����^�!K)��lS:�� ��C�3�������/ ��K��$o"�QUQ�-]]h1S��*V�O��([ր �vk)I�^���Zc'Qz��EB�I������ȋX?�t�$��/U�p�x���/�+��[��)mx�^P'��غ���1)Y��[G��hpJ0[�+�O�耬t']�|��S�������
�����JYI���?P�T���ҡ���;����&O��>
wPri�b���ςm��q����s5J�Ml@6D�^�/x�K��f/�O6�y�s�ZJ�1w�� hp x+]�iTD.JB������U��	�&FO0ƉW��$v���njO�;��r��A�Q�C� �n]\��P��?!x[� �{G]D��h�X<8���$����ώ��'��$��3�,"H���5�v��31�����R�l� 4y�_��b�A@� ;�M�K?F�ZE���&9�ݫ�����SP�><.�ri��;wv!;Jp-���2[�.�	�|�U=L�,6Gpu%^���c��H|R�CE���_��q�������	7-�0j� ��,8]��񉀹
q_>�)xY���hج"S]'���6�-	h%[}�$��	���!�ң@���]���'�')U����<M!K�>F�:��#'������o$��WY.���$X��aƬ����Q�Ň�ãY�À�R;����������0y����0xl��jg���B.�`W'�%�X�O«����#l�����hv2�_���:�,��e��[�������� Uh:q�i�0���Q>��k߰dz�`=ho	-�j�	���� ��Ԥ��c�w��a�5�.�4o�^1��6P'�0��]U�3ƃ�
W���䁽z����#1w
Q5X��	}4�( ���q,'A%,G��~6e���|O$�H�-�%b�`;��iG�L��\7�̆�.�pA�K��!Q���CaL̺4��ȭ:�9��ŬDA鴾���g�mX�,����W�j��0U�=��{?,kdR@I��щ���0)���V��/ �����'�%��Et(j������?h�!vLY$�]_���0�y<��1��-�bV[\5��y�+f�$	�'[����f������h	�< ��&,P��uN���3%&��%;D�!��h�^�1*��=�k���2�Mvh�z%b_���}G��
l?���$�Z�A"8�Ƌ�ι�5�>1�.�a��OX'2�wD��3�+<�Ɉ}<'��H���%CV�@J ��H�^�+�\��9 ��e�3���hlY%_7�@����ȉX�{E�G�^U؀�`� �z�	�fR�����h�i����A�(��T*�����V����[ ,H��C>� �-Z6GU�/�p�ƀJ���hMP.�-���0i�5�[�\���GvC�� ARK�71�@+�E/D�s�	�@'�� �#�LZ�_��*��%�1���l�m�ou��s�Xż	U��|�����vk
�L>���O����"��+�ђ�p�&IOJkJ"_e�@r+S,�Jg�h��"os�,��Nv� t)6j���Z���k�`�[h��ŇR��$���]���6'}0��< �N��'h׎��_2�3+�/]�{C�苀h2_%ɪ��k��˗pN�)�<�	�H�W���_#��Wŉ� ޕ���*����!8����J$����Np���)����VӸ��1!����q�{א�-%�
N@5� q1^��j"S6�p�r4����YX<n��"�A�;%~;�}�jgLU�������~�P��Z��@��Ղ�}a.G�{/���\�|P04�?"ҝ�/���SD��閱Ҡ��V�F)�h?T���fej�9
[�,sA�%r ��d(�S�6B��#�wT�[����	^苰a�����\b�������������n�'���p�,Ya� �Z���:y���us�p�)�^��^�p�2<G �
���W�$���<0������@��xg�ºPc�{!�� �%��� ce*���y�V�,�6��@�}1	_����Py-G�+� �J*Z��%H����'�]������-?Xp
_��kډH�&���)�,�����-T��
�1��B�E�]�s�}uw*d�Ko��90t�MZ=�L���PW;m]���{���W�/X��<M�r~	�N�Z�f��J�V	���_'�����Í��궫!�]���'х��b�uXj�u���b=]� ��:�����F�4,�v�C(J�,:�|~%�`�;,` �'�B�Y(���$�ls̵���WW�������	�"����[�� �`I[�����_�q@/`s����fi��R��:We
/YRdد�	z��R
*܋!Y��T��0ʹ9�$)�IÀ�k�7�t�/'��"j��W��$_�^^���dcs,�.�^ �+o`P�ad<�I0R�8>K���ѭh�J}��F�؇���ܺ���Z,N�N(���_���|��.3@{h�8J^D׿����^�X�n%���eí&�u*I�[a���D���?ӵ��P�1I�(�[�]5 �#O�g>)��(Gś/�H�|�`�ܺ�;�,���ҞF�6��\`��Z�8��`4�+�p]h�|���f���I����x�h�J8����
��
�U�4:�㗁��&E�����	iqCI#,2����т�Y�xA�a!���:�Of��-]�5Ⱥ�Iz���h�xh�!;�{Q��u-/�6��*�����$1���S��_>*���kW�Q�]Nܽlh;���ݥS�����z���9ZH��hZ|�a��@0�Z	�S��\'^��\>���چ�nxO]�=�z.pN���#pz��!@T]��LG%8@��-�g�H�`O��S�a$�ks"0 ����jI`�E(�ZP��]V߅��ҭ�q�	���y"�v-%�n��Q�p�h-�`Ij0Ċ'
Z_GZ�����Q�+F3( U��7g)�~j�D��ѱ�3<��ITA�C�S���2:�+�)�a��X'�
�4r_�UKWZ��f�]\�Y�>��zMJeX-BP|:-e��\�U��,��e����T4�< )o�>���?�}!�������/��]�;p,���HM��-'������8h���!;�Y����s��at[�Z�i��o��+�UMSH"rU�:���hc�u��4^�iZh�[�T}�u� U��H���_�����3[�b��5c �I�s'�r�p��l;5H��a�w)<�B;0�!x\�z0�+m�$�>J��	@R�1�H�A5e�A���t��ZSð ���[)тN$]�OU�5NY�ہ�o^2{	��Ւ��J�ԡ��^ҫ����������3>/.B�-0��\.4�[�� Q�DP!�� ^_E�R�K��
eS�Ҭ&)!�Չ@��~j�2?e�	��]�#1������gI�AwD�$�l�;:�(�K1��>j� �P�7����trbZ�9U��������sA�+�8W�%��H�P鏞� ��k�w�}�Ʃ�щ@u���S�B'|�`��1 �-��z�!�鎕��x$�v~,YVQJ)�r%ӻʓI�->t45�C�K^ݾ��O�����#�AAp%���J�7<�m�4P��q�Q �;1 �Q��)DC�y��k�'40)�:/����w�-2Q�+��+s �rPR鐀���d�(�]�`�O֋'B 
�r����E���Gǀ���1����:�
M���:ɽ�oR������8R��W����tA�!N �˕�Q�fh,+��$�=v�~PY����c�	� ����^L(�%�W�<h,e��
�]��K��P��!}�y�<�}yZY��[;��� �>;'
ߔn�{>{o停�sj�6����uKǷH��U,>����Y�(h�~��%~�40}��R�_�Z�<k,������������ @Q�ڕQ����@�C-���`�H��)y���'l�D�e�-��Y)z����-�1��Z��~3����$�Ln��BUa�grE��<2���Z�� x)���`z\��=�g�$֝��"_�>&z���[%=��'p�r��P��gS[D��B5�xlrX`��0<vd��#�q)���cf�[9��l.���DfJ��@����t�rȃ�P-3����N漋���w-]}��&�:��}����z���+U*�e��]���i�*�%�G&R_[	ғ�9H2X/@%Tco5?g�AA�t3@�-%p"��XA�8�:УR�\�yLS-E����N�3��X�}�6Τ=�@+H�HhO�\��S����� *�N$�L�U� ���GK{�	��w5&%�J�e��� �^��0(6M�/[@��2�,�0��4B��hy�45�Ux?B��z���b2��8	G +��N��ؔ��o"T��@��x0�8<)�r���b�]@-�u�s3����[�0 �fYN��$��I���Ӗ�� �-K"�A�h O.)�p5P]��b�q6���P������0`p�J��{�(}&`�
]� 1�n��oRWeU(b� 3�	�L{p�)�2�K	'�@�C��hN����^]E1�����zw$����?4|h���(�0�Xp��O��[%7x_ׁ�2`�_����F;#	U��dSd`�f</yKai�	�ʐ�+	�^h�2��Ҁ�|�N��Z��V5�-U&�벽	tS��� ��sh�%B/��������w�)����J_�P����^i`�}�V����	�pB�v~%qR@�R&[Kf`�l��(/�8 �1>M��m}���:On�����xhb�)�I�wP���=<(��b<�:;�7Hs�Fd��X7�bXnU�`4mh�D&�x���1����'L��8�(��xX�A���'a\��.C����ӧ���T[�L<1P��V�q:ccK'�P@�p����ɩ��:��IKc��!
�R�tb�OaE�<)����V���
ZWηoA�6(@�:fnm6�e��ӐXE:C=ڃq��8��5Z_ȨH�>�f�zH� ji�(���$���B�)_��hռ�&z��!�Z��=w-� t?�T�(!�����+�����~�a������$Y�m��ã��@���*91�X� �\v�����sB�Zʛ��^�D�G�Q����@Z`ìE�6�� ]�V�cI%�x�>uJ��e�i�� Iʛ`��n �Ey��6e�9ɠ[���h�k�N�j�h�o^���� N�@cL��鹙��z�|Y�j�		՗>�u8!� ]�IU�y������E��l��m^VhPR	UlU�;�̡;W��&Ъ	`F��P���VKC���w�	� 5�2�#�S�Q6�o�v�$���v�W+m��\��[�4�͵���n;�p+(CPNF����[�'��z�h}���xbP_^h/�~w;�j>=�[6^�Ph�o�W��@�?�Y���[ 
"�}5Ax����@��=�1� �h!dO ��!m�A/�+WL@��+�`�r�z���=P�$�n��\�2`�h*`�櫱�<	��Ch钞-}����9ӇuaKX��f<���ײ3�g�Bv����:����9�����"��.@MJ��(+C�����cfWA�������Vz?�X@X�g��g��s$)��p3_�Z �[�0h�$T6K	��@U�%����Ж[��BJ|{QU	@�� ��4o,�����\����րƍ(����4���~�O��+�������]'��1S��pJR���@���14aQ�a��H�2�T��1 轱["a�t�)���
#;> ��o@q	`�Y2�A�C(�Z� �#m1�)�R9h(P^Ƀt�.J��������|��٘��j�]y�v�{|���)j���D�z���-.P�W�XU���r�\�}`��_νSJ|a��g�֣�^�S�s�J�`���:1�_�*�q0�߽	�T����j0X9Fu�1�S�3�E�o�*'�~�Z`M�/p�peQ��������K��O쨢�F�V��e���@n�:�5��$���Iz�|��L�PW ��O�'%H A�k-����;�v$�dW���.e�|�D �/Ld1�@��
��s��W
�:����� �la'�B7wqʖ��|N��u5��	���x`(m0��7�J�|�4:���~�O����Y I�S�@G]�:~GЋ�X��5�U�Y�Ȅ<��>	]Ru�dC?�� jYQ�]�̀��
�!�`a�e���ԁH�bq�+�d��2�4UB�'	5-�y�����l�����!Ӵ��L��"�0�RF�`��w�%���`	h�8�q��"Ѣ�X5H��`-��2��X��ќZ_|^Qn;��TZn��O���<hݳ�K��-�F�LY�t(����a�Q���@!��b���׿�b��y�>K臼�J��?�t����+�~�o��s��!�>��~�o�%��Q�3E�'yKS�A����#��N��h	�*]�����޽�X�Lx-M.
� ��u�����*&u����"���zL�{J�d��&u�dZUŎ�/��&5��Q{��B�	R�8����h{���}�aL6�R.�	���m��LஏOa��������ڕ>
��/󹾘����0�f�S�'�}�]�"��n�#�={�b�2	�b�)���IGX�͎￘�p=��i��?��/ET'���;��Yp��'���u	�}�Z	�P�QbM1!@�j(��%qu]��N^�J�PV�7._-��顺�ć\G`�!�$�39TB����(i������$뻚�8L˱�@l�h�V�#Z��aYhkT(r;��Hw�*�&�� M����x��7&�I���qc�r��#�[�$�܀���a|�2M %����(O�JY�K�� 	x<c=��;O�;��N��ۅ�<�	�w%
��6h8���W�j���f�W;�}U_��='Ω�A�h��5j�A<�>rB��60'"�v{M%�1���^u #[s�l
b -�3�>5���g=��ʮ+w	���Z���`����/{Z(��ȳox'���C���i�9JC��[X6���$@47��(?��@<h�c;�wϪC���[��'�{h:�3�O���&]z�A<K�`RnH����_4�����B`{�u	�_s���U�;I([Zq�^H'N1L25�������>(Ӗ{�Ñ���hYOF rU��I`�� 
)�-�F�v��]!�^8_��b�Z[}��!�MK���J�H/a@ND�2�6� ��R)�h�^[���8�[�l	��БHi�Y 44|�1�� ���.'�m_1YX@����k�w��i�Ę��0�2�,\~�o�7{T�Z	�W�|]�4!�Z�S
��R)߶��J
�*��e�����w�w�zh�a�Ob ܓ��/�+B~�����(�<�$[!�/r����Q|�T~҄���;�	�<��.����N	�����8�������I�^�s5�&+x�fj�F�=��1�)����������!��0a��ϦA1�&��
����+8lbX	[PiE���vL�,3+�W@ɻ��?�x[��B���Y�R��*'2��t�-��Yj Е�R�@J'�5��Kqe���^�B5�[aT�.�Rz������g�ydb0��v�O��&�`��Q���O�UGj�P�4�F��I�T��`47%��0�t���}���hE�O��y�{��3S�v�5X/������QWyv��aa��ޜ
SA�8(�[��;^ ��|�[^�>y���)"�i�u4C�̌�����J�"Y�������D���z�?��U~�
��6B1�}�%���(gx -Tv�>�������`�~/'���)���q��>�A%�un �2��b�Jl�H�gh[�73��*�M:��ܠ�H��^)��F�����,�r�
�^��C���|��
�-\w�j�O�"�ѣ�r�,���Q���jɸ�ӅSMr0  ��0N��E�E���6em2��p�\Pk��(m���=�cZ�:h/i���n�Y8�'�V��>� 0IE)�hg/�d�a(�<�鲅 J�b3�\���YP&��=�r-L��^X-D�
gi�������x46T�ܠ�������P�~�Q�rPޠioI_��g%�@���|b=[��ݲ��Wh�S�Pw��	A<�^�I~�1�Ҳ�xU�dP?c_��R�!L�{)n�j�Vq`�!��>�VA#)� �{�=����e@��v
�/-��|��mID��Flr,L�
��/�z
�-��ْ��XV A�5�zK�W��&�F�����T[n�	$�=a��u;�I�P+��0�>�tZ�A�M�__8@��H�)��"���B����Kkn"hvِ����3��.�e1��+����01����A�^+���b!�U��%�W�L���΋�.{��l���96�T" �Qo�ט�b������#�.�-���o�J�+B�W[�Y*��\C#aE�jS�����k���O�+��HvVR�BoQ;�2귬�f�.�e��P��w��P藓�8-�>���+��.�"ɎY���0��AÉ�H�� �[�?��䀵�V2W �¶v��q�D�+"�r�F�5�p��&J`��A{�9���P��O �Q,u��5����Q=�J��L\�l�2�l�u�
� �Y���C�X Ja(�G�E'��]:����8:[�'1�UN��Yha!��(�	{�Z����%S��W��3�6	�1_�@�R��K=C�*7	J�T�	W��Z�#�P� Y�y[P�� \F��@�?�-�}a9�k�U�	Y1��pl�Jx�B0]j����hP����Y��W
vm�%��/!7��)ex'����(�d���(�y=����� ������%�^�3K|�i��mzaUU�D	�]�5Q�';J��+��w;RfS����p�J��e�����R����m5����Ҍh�lH �jZ��G�y��]WH�N����=r�X_!�.`�����0�&1�S�q_�P�#�\5�(���QAk}�q �cI(�Y޵䡱H��N�v>d����/�gLdc��
��������/p �j5<%WE_� ���
1���tF�y.!ѠKu�V�6��F0�_��P����6�o8z}3sph��"�K�W��*Z	�}ex�]8��)��g�v�2�1��
j���*\/Q��׋nX��pv<�I�����I�F�7@����D��قM@�U¼��L�
9�1���0�`�:����z�:8 ����f���DR�3>2��^��Հ\�O3���Kq�^-%�O�� Ҵ����IO�+�vK�g�2��m*;��"Ug�e��v�h9{̌"UM�E�q�Z��z�@�2kθ4��C�]�/�� �/>��M��"�>ʍ�����;�a����hD_�y� �Wz�/-�.�/,n,�V}h�[r�z�b������o�^)����[ĢZ�DPl�~4MD+�`�`���O�?���tZ7�� m.�_=�'%Y�,��%=���|xC�
��q��	� Z����y��� �!�8O^���]S����\�P7p tD^h��~��2�+R[u����VH3'��j�M[b���s�d����B�F>,T��`[�8A(ޭdԸ�2��,�Ä1�L;	��O�m�J��-ȧ�N��o�N���[J�,x s=a��iD-��Wd �o9�IKxr ��
D������sGـL�V�I;$Z�!�\�-¦B�	�u �?w('����~)��b���*|�h 0tj�S�;)Y��_��'U|�By�-[*��ְ�X�R���%^�:������ac�`�p��ƕ�+�E!�`�w,��C���:h�.İ��[���Z�+!��K���d�)]e�E4���qjaX�#[Z�ůN�O�2'�����DZ/�IyV��X-Y�����'��?[0�R�nx�-䉎<�7=�,�y�����E��<��<]#)\P3(����J�bI��Ñ�П���ğ�Z$v�G�6YN��<��]���J���D8���9k��>ֲ��B�B��	��۝A�o ��	�9RG�)	�a��8 |^15���)�<�j�4�\ �&a�R�u�6d�}9`����k�:<!=f�{@�<�R	��w̫@�mM�� �6*)��'��~Qt������0����u
���_���"o{�2��1���3��hn7�6�,p�	�i�lס�*U�n��'��_블O��h_wJ"q2Xe�D��4*��Z�� �>���+0wB��vcɈ{��A�o���qClO@Z�&-:��_*����	$ �O��^���E������N�*`�!:�$S'�ZP�"|� ����1�&��^J��,�8^`�	�g�n�S/R�2��B� ��`��JN���X�^�`SY��i!"�"���K�H3"S��_}#b݈A�BkW�ϳ.�ɀ9�ȥ�^�/Wª�5�%��.�H�J�*�5�ZԐ���@ֺ>�B��Cd��\�N�m]��r9�ϰ��3��:���ȉ�/
䍗���d����}l�e�p��8��[��ñC�ㅺq13 ���` H�,��U{�NS�]yUP�蠊)O~�� ]�8�X"��&� b0-�2�}�)?�pL�;�'�A{� n0��y[k��"L�;�V�'P�(`��mfk����B�qA�IH W�/S;��߀���C�L> G��-+�2	39�V�t𹈲�<�wϞ�M��������VS�g�����a [�訦�h|A���2uv�9(�@����W�E��¬H݊���|@w)��L5X ~���*=9@�ʥ?����)�^0��O4��J��Ph�U`�ĝ�F�!��^Ҭ���>���Z��t0a�^��O���R�������Ɠ	�p�� }�K?���"	�	��/�gޯ �_u�;QŸ��	���P��W@��dFKH��R�J�$��" �����o y%=�G�T��3���2u8���^k�np�:�l��[����5�y�oh�Wh�E̝ca��<�]��������[��]/Xe�M(n���� D��a�?�O>���AW�RLZ� ����Q�1�P�4�/���C5�A�Sp��-���/ZGz��ӧ�W�����2
����+�u�l8�3BQ���V�xd-��8�JF�,���M�:܍�?�y�uL��(Xh��f��8�&]p5k� �f2�M��/��h^fCx�����!�!S��W�w(�m��Ws�2Q�w����2�^}VT^v�R�m]+1��[���x9o�Z!��ىo�Rş��+�NG���3t�]^|Z ��o�5�Y1��Q_���6��[P%G���X-��&5)` ��*� �(�%�;gL #)BV�I	�-��������gtA�)�.ź�!M����Î]ǚ|[�&k)(������)=^�@�g�Q� X��J�H�L� ���"($��
��XK�˩Q�{�\��=I�P�N���Q�}����� ~d�P� ^R�AoS3���BGf����Ij�Fn��p�<�x��{��H�>�m-���ҨT���+��Y�� h+M%���>|�L�)	!�]S��}�<w���uPh@x�[[P��@�˿y��U��y��EL]@?C�ǚ������z�����ܳ�� 8`�KX��?Éu��՜T%�{O�S�BA��NAh��D��/C�~�D�� �s Z����7<z6���^�I����4e�M� ��Wz�w�)�?�>��ݥQ!Z.:�  _?vD�f%i���U��$1�������V5YA`�z!��=m���K)����}'�QU�D
��E�3Z&y��"Q!�w�R-:�Ul�3���Y��"c��%�����a:J��(��ʯ-V�\�����<�i���O^	��U�UA\p�W-��n�J1�J�Z���tx���G�f ��;[E��A���]]��	�� ��@�`4T�V�R���>�~ �W�b�[�x(�E�X	U�'�0�$Y��YQ��0S����*��%V^U��� �DB�F!X��7=�C�I�ĭ�}�%�>�4^]��"�����
[ᨂ��[:l�pf��&-�'�X�W� ��}h�&�I��0Zf���@\���H1�Q� �f%y��-lB
����(�-]*W��h7K�:	HXO7WL!n,g�r	_��q�''wd'!�����SR��-��sJ��!7&{ ��-%q,^3ɲ����w��^Pd��<�ܯV�鄩'�c�/W�<�	�G���Rn����wh�qF�A�`�S/�1����� D$X����A|��P�;B�k%�v�D��%Ţ�0!�\�P?�٘�'��ߚsWg��ū���;�w����� �@�&"~`����R[(���41%WS�j���
m��4P��0�f[��( �N��5��478���7�	UA¡��@�TY<�1�L��l��|jP)�w�Ļ�Aeemv�������,�ݫd�y�I�;^�z1��sK�QS��ƕw�`z���v������^J<p�u;(�g�2@[����,��	�r���{\�j��T��h	b�%�*ŀk�[�x9����� �F4{��T'wJA�B'q�0W��_�- i��=)Ⱥ*X&��k% q����RV���^q�D�LckS�*��S���������c�h�v����7��p~���nJ�;��E�n�b�[����x*�J�9i��d�q�K��|�U0�f1��2���g*�����Q�&�Swt� NY��
��ɑcjO ��������b�%i!��蟄� 2S��=2`0N���o���y���W?~+�vE�]�'���\��+��w�'�6��1,�(fP�Wп1xr��v�^���ˉ�{�o�,�W�{$3 1�Z�=�n���2��Pܕ�!���0��)���^5* ��aO3�r�^v\$��y����:� +0�X���ϰ	��[�6 � �Y��*yHW�}������{����X�W���_C�����1ʻ8?����2TM�޼ Ipb%	a��/ �>`-�6�`]h���MKE��`�X�_����N�@I�o�(��	,�h�>������dS�?�_pe�Y*�*�_��	�џ��������il��u �N0��mLR��yL���@��^���zs�LY��`~�c���ؾ.!�a	��UN!_���:�����	E	g5�5��!d 1��0�fZ�W��c:��C}%Z(���Z����>��"Ju^�	�\�������@�P��O-���B��okp(~���frQ�J%�4�}��8]�P�U���	-�>���Tj� ��Ph�H�z/��Sv�n��gW���''���i��N�m�NuTO��H��:���t=�jU��b-�S^�@�5�-��M��H;�A�{K�L�B9�)r�H�0 �e\��5�B�FWf��np�H0D/�vf�V���N%)���T������!������<�y���n�Y-)�q��u����"2,�z.�&�к�mq-�b|��!��l�,�j�u��-�)P��?@��͍NvX �>�C�~�c���o�b��h���{�k�0�������u��Z��m�} �<OA[���� BQ�C��/u�^+P2aB��&>�~�a�f���$zYQ�1XH�FJ�8ù>Đ�E��A�{Q?9bn��`�/,^��x?%x�L0PW����(�K��� LQLL���\)�XQ5 �3^[U��Z20����3#<���h�6��a��ݧ��"w}ќ��h�YX'���4��R5�/��e:�-��3�b�T�� �v+#	A�^X�'�g��)�ME_h5a9Pu��:ƺ��!�UD/O��ڂ\$�/_�?~��¨�!^���_1�sd�K��	x>�%� ��=`F�	�B^�p����;��u�t$���;�7�H��z���P[X@zQ�A
�
-��M�CneW}�����w(Zv�?���!�i��]��9!��k|������x���=W@��Hj��b����P����iW�$�:*fX؁^���hrR�x�,l���ny�.�R���tϷ�1U��@|�B�J�{!.|4x�A�;� ���y�2�I��,���ݽw8G�L��/�d��X*��+���{׹"���P�>���ǵw	[r�J�^^�2H[6�nxP��hL�~�_�0���	��]X�Bx�}`�b�A�ND�p���Cq@�-9)��S�.�8�$L&9�Ĕ����s��!��Ĳ�[}��C��H�����1�{�B��2+W�j3�4ScS�@'�F("k�uP	��{U�ø�����c�S�$�{�	�X잴�zy�7 �X�	��umZMF�0U������4���@���{�o�1���p`H<���Z'w:�`�J��Ћ�P9�}��W��c�R�T4^��UߎD{-�4V^(��)N���BAP��(�fXR�� ��Q�l	�C�yNw9i5]b�	�<K]��x�/a����vЯȁ���^�A/G�p9�4��v���E�5��3[RVA-�d�^��Gr�H����_��1_�g�/�@&�x3��s#D?k��#/E��w��WC�o���G�{Ք�4QO��~����Gi����o����~�1�6@2"/4|D�P^�M�К;�m�e��������t	T_��C'�N���6�~^4�5�>([�XbU�u-��|���� �E�Q9�h�~b4+�އ� �(��9ꪻ�
f[W|�Rҕu2d�zd���&6]r>�Qn�`�U3Pg��Zf�O �G�vI� ��ŗ�hCR�������ʻ�0�"_|0�(Q<���W0;�mf�U@~k"�1���ғ�,Y'RM�$Ϸ>�p6\�m�	�]̽-�G;Fcp�R�W�`Y�*[Y6��g�?]���-���+侲��鶬�vhKP/ט�kyH_�5=۟����s�� ����1����N)��T-V�>�H�3h]�
US�'F��Ao�!���¢�B8wP��Ya�$[1���A��u�3� twV��j�Y�>��I��"����q~���)��	�1[/����S�AW�8�5jOP�+��]S�h��_t���,FB��'&��p�j��%B��O�UK��k�
���'~(�StU��1:	ч��� W����I	����l�1�@���Y�躡9{ E�Ph��n���%��Wh��s�����J���@���������Iy�3	ztt6,n��]�zHj{_)� �!�[��-Ar[`�*�&�!Ȅ�_[�@�΂�Z:���J��@�Qh�f�MX��%�O`�-�$�.��Zk
�(������tiY���br� ��ς!?��p5x8�\(��O�d�ȭ8K#�$&�
��?ºw�Z8��p^��
�,�Q�
��7</�cנR��(7�h�n_zj��~�����K,]�c3*�A�NCn��	��0tG,!�6<;��r�A>���+�H�2�%��
v0<�/(-��"�lE*��1Q�Yj�$���4�>��gP���6;�)<�	������U�Y!�^*��}��&.!��+�tR�X�7��%�a/Y������Z���RT�+�/��y���'?o!�)҆X9SU��+�5֫g'_J@� ��s��)�A��,�Z���.%QYB&�;!J]��P�-fj���>�����5 SgH�J��K��O)����%�F�,�wW/ҌB�U��6�l1Ew�л KX��xc�� f2��P�Ks���@d�I�u�-N�V���p�'�h��.�*��\R�x�(Z�	�`j��XI���+���Ph���W�	}ү���4`6�	b˂ہ�VF0�-�/�b�=S��
~���[�󫷸Ґԙ��]�=��I)��G�!�p��%�}�ш��x��9cot)��u�� ��
�m��>�ɼ �_Z�M�z���h-J8d�NR��P�/ZDX.%��V�~���׍�3ʇJ��p$��A�()K��,��I�+]X�?^�Z�)S�ȝV��F�-��0�2p1[�b?!n p�% �����{��A78��UT��pk�^���8�`f7���^h]^~ɋw~Ha�R�>�Ȱ����jv4(����z���(n����4�]�LQ�R�K�d|z�F�hw@!�&HQ� +>������FU�����U�	�vx�w[���-uP�/��i��^��8S�Z}|P�X���������o���˓�鳌O��R�y7�G،h�l�#7��ߖ?���`@	!zu�@o��L�n<1ڃ��"�V��0du?&$S��"��U*�}K���d4|@�y�U���E/�g�1 �{`6�%m������о[C�^�X�~^�mi]�* ֑�~�P֜*�yS!����m�6�h?$���=����UO�w�>�	��w9�p�R��7�Η�%\�H�.})5e X�h*Z:��5->4Ce�Єh�\��6Z�C���5��G1^b�Q~�B���J����-�S�?pD��胮ʐc�)2��,��:�,�!��G�o	�s��I Y��v)���5����gW�@:��VE���_�a0�NwF���X_��0��:7�߷�19� :�
|=dLç��NȁCj �P�.���$  Z,e(��9.��"�3P�ʊb0I�	� �����)\�CG�s��0�;Xؑ��h��ٸ������t'_N_�	�c���ſb��k X�q?ea0�u��1L�X&"U�i^�0l�@�ʩZY�T(�=i�!B��2�\��,/�tmV�E��X8Po0}��tR%�w�&�8J����|g��C�o��+.�E�V�@���L��]�s8�}/�Ԟ8;���`��aJ� )���Shs{W�E.�4c��LFz-_�:�������+�h�{������}�}AA;�hf������`�r���k��	��yOW��gU�p���D-��J��h,�o�%���㚉		�&�^췂[W�����m
�T� Pq6?�*���K<�j	� 01�T�:[G�����]���M�'/����qh�q¯_�^2����V0���_������Rh+y��1��B��0i� 8^١���;��o���&�ӫ�Za` ��^WT��u$��I{'/���/*�i���.F��[t_�*����5����O/VS](�����Q�>,�څ��,��@�^�����C[�^��vw�F)PX�-�j�u���8<ؠ�[� "i�'h7q�{~�� ��D�ER��V�,L�H�$S%joج���=�!.pRRVn>w��/$qt��j�a��X��MC2@�n�5�W$1��s%p (�0�I�~zA��|z�����+�:�� �M�0!o �itg�+H��p%�!�������fPS��� B���A/����tQc�o��By�6_T�����+����Y���Ij�s�.QE��.@���#4��	^�* 7mT�-�#q�g)<�ї���/hP�C`��3(�, Z���?�JN9����t(J_�����C�V1|��f	?��]0Zu��D�)H�n �	J2�H J�B�4@�?��F'�T����P'��N�T%1^A�k�I���n�+�%T� �7��1rՖ��!p`�Z���;d�-�<.�1��������9������J`b$�[�e���@��ZY�`3Uhn~�Ne�	l=� 8�1%�C�!-����I��Eѯ��}(2�(�fq���N� Ӗ1�v�l�k3Vtx�gP��t�N��YfR��]��Z@���#�[���(������A!�`�%p�qA�A4p�ߍK���h<�0�_+�Yf (��Dr�WQ��V��\�p�J>+x;J �I.5���J���92��8��7(��0� K���Ub]@���0��Ԩ/�Y%��/a�!)ڂ[��*�0�Ces�����u�b��<���7�F�pL/Qw��!��y�X�#%���4DO�]� lC���	���ě����f��"�Ҁfh�nTPO��k�}+�y��{�'��P�C��0���&8�B �G�(�,�"�	�M�ul������[��s��k�W\���~�^� ��o��lPBʇ��4^��M� e�݀�x��O�5�3OԈ%F�Whu���rh�K}'����B��i�-]��}���ܰ1�;�q,w@����)��XBS�,һu!�I�lc ʩu�s�t�JN� w��<&@%�Ue
��Z �'�h!�	�	��W�q/�Ҁ6vhQ�~ 5�K!��Ɠh�&z��A�<�Z]l'��X�l�h�W ��k"w�˸��[��ɠ#5sa`4S�8.�|N�H�����cPR,̋�A�,�l�)eL �{�T��v��ݘ�3�\�P� �	�o�����១�������A�	d�-d����,�)�Y ��TP	�_���9k�N9b��fu�q����܂�[@��ڐ��UL�L�|\�eT��^J�-�X]x�QK�>�bwH���(2��#:wd�?p~���mP[�ѷ\,���%�h9]���H��l��L�'��-�D�؍�	Y[o��Ƕ�1Ҏ$]~AX�?,� ��j-? ��6%�$�^�d��1�]��Ҡ��Q��W>�fշ �b?_�;V�I}FfilRe�O�v1�ڽP�KJAO�(+ �=�Q��U��� Z\�$������J��&	F��U�X	>���Hav+�
P�f�{^��aI~��B7�H��'�����(0���fݔ�5$������T��}L	KQ�8�P��p���i$ARI$=nW������J����$�1���,���ҀzR2��]ߘ�EH>s&S2=���X��Q���c=3�	��9 ���W(_E�;�[�b�	��@Y!����E�[=�>����i�*x	~!�� �q؏.�4�*��)��K��H���zZL ��:S�1H��`��*�c��KhX� �_�W�] <��������{?<ГfS�=�`h �-�npw,(��v��t�۽f<Ic��M (�Y0�[��rQ��Z1�xZj�`6%֮��n���A.L/�(��bk�2
�X0KӖ�(,�
����� �q�G1�-;�` h.�l���x��O��;��s��ſ/�P�VN��$�<b�h�W��\�S�ak��6����8X��%��A.����Ѣ%������^O�TW��#_II��tpo^=f]l-.��0��.�ϰ@�R��tC�??��>>��ҭ0v�jSh�+�es�_*Pb.1*��0�k���U�)�8�#���c�)[��yn.�hM4�?+UӛX�
I0��{���A��L)�0l1t�c�>��z�~���)Y�s�L��U 9��Ή͵�)�����^�'[	���f�$,/hO �W�xڞ����)��1@���N��F-�����d`�M&*\�TK��_'��b3x�����[��R�V��S��:�Z$_�L�~�r+�K��JCrD���+��-����&l?�j'
_z2��Y���L�h���!`��3���/��Db	]�jn����(M H5Dk�W�� ��R�S�^$�8�hА��'�ǖ����� �_��2�e|����]D��lh�H�t�-ѥ�@�WhIy"Z��>���z�C�>�=��ױ�����.���G��p�M����`6%q-'��ė^��B2��$�;C�R(�iz���4�`��(1��	M"dI	]�@��W-���Y�O�#v�[\�K��N>��d{[�%Yu�S�)v��I���̿Ix�OQ�����#	��)��|U;xN�%hc��n�����0�.�������[J(�d���X��I�ʎǧZ���%���M�:�f�;+E�a7�+�Jf>�W!E��hJy����Dg^s�S�.�`-�YHN~�� Rh}Z�NO�Mo�eE�a`�sA{V�k�hLl.}AID����p˝ 5R��H%�-��VK�б+m9�ԁx��>	~�?����mj�W�!��.4���*���VX^*��x�v@xlFZ��m�`���h~�`�@J��f3�+ 1,��HP�ki������R���ד���<������!���dF�aS���N�E�鸜�����m^1�h'76�4��AY![ʩ+��K�XZzB�	]��w������^Ѵ9�?z'l�1P��HhJwB? ��|�Tn#�jxR@~TF_��~(��Q?�*��8��;�/
�L� �����IH�.���)�ĺ+�K��0e�V/%���`��A�kb��%{#�n�!��1�k�֋Hܡ%}2?�¿A�Ws���R� ��>�&��~�0��D��J xA��yX7�2->��?�T 5T!:1��^��Wn� N��A�!��֥ԍ��X��C��^2�Vhz��坋��(5\K�B� ���^�1����b�4�R4�|^�|"��ZY� �-_�Sh=�E�R��]�@�&	f��/N(�*��W�cXH�chJ:n �r0�[�*����V�G����Y�	�w���R�vu`uB�o����
�7����A�]i��()�.�<��:��	�����U�Lh�0L�@�c�T�a~R�q}Q���Zv���	CΨ��.K��G0!g�T�٨�V鳮������N1�@��@�N�l��>%�W�DpUe}߃X�IK��������c:���S��[��<���R�V)�
��%tQ��F�GV����.��)C�&��K�	e_�d�F'��G10V��r%�p���Z>жpCFO�l1EQ�Ӎ͸����	2�lB���T4V�A�,�������RF0�\fh�K��u@5ض�*`P�	K(Gi(�'֨P��(�ۛ$�u�VLY٨�^.�߿ /�o��q�'�x�)���5�m���6Q����J<$��D���� ��65�M�	��ω�����	�_@v�w5��HJ�K��#N;������ ]�b�S��U�\7�:�v�L�F�+��Y1�JB,�?[{��_8
��?4�I��H�S� lqd���K����~W�"�I�_��5؊a^�\�I��U�������} ڄs�&�G%}����u٭CS����-Wa���)�5�8j�	�2�G���	9LX\1�/�n ��,�[E�# �i�J1���Z<����򹴻�H��ڨK��H@���\ �5��AcVUI	K�S��餠�J7az�A�����e�K) �ܶ�g����Rx�E���Ay�W{M ������������z'J�����Y9Sl_�V��#�,'��]�������IT6&zs� �'=bu�t ��3N��-q!��Y�qA;�8-?!��g3ϐ���]fZ�)��*�wU�'L8�Z�s��pA%	�sR	�+����	N�g�dH���/�������v4�.�c/�+�	鱜��lNc��3$#Z'�]�d�fA� Yq2[���X�C8���&�z���_�j�J�PѮedz���Q��A�A`�����X�����(�Z �@Q飽���8E�������Q����I�F���E�l���j�K�Ypc* �iZ3����, ��yd��: �5{	���Py�0l+G%&�*�/�;���W���Q�C�1,��� ����·���} �d��ob�����Jt9@�QJ,�Nk2V +}(/L�QO�A��D=��3�T�]e0�l�u4R%��	2�DY���v��2�s+� ����hz@)˫߯(�Z�޾yKOb������32�)+kA�?�;1�Gy��O�+�%V�yDKQ!	���o��Ѓ�@/���c� � I<���ȾA��r�_/�ZbX|Q}Lx���$u=B�58A]KȻ����Xs'�נ7�Lz`~���Q�ѿ~ѧNL��6
^���|�9�Yj�����2X��^S��A��[;���G�B<�6M���M�PL�H�U�.�4m�r�Ǧ��$Tu�,�cm��"�)O��ɔaS3�<B�!��U�\P�vK'��S��8?����*�+�)r��q=���N�	0b2��|e��<��ق�)�0���$l[.�Ƒ=���'*_]k��"���D+�?��}@�6''�Y ��xM-�_�F�tHJYFV8��뵨G�.1�z-d�[�h\!�"�)y�<�����_!���"�O��hMrk/����9i0z�������δ	1�!��n�m[GXp��BW���R��@U��������q������S-�9L�q�ژV�k��M�	\����J�)O��Q��.�%�����!���@���x���]�?X�W�N�2�%��B.�Jۨ���}�@����M���T��ݖ=	�h�B]4"�����e�[��`h8�Z�}�,|_�z[S���	=^�;�9���J}��ǂ���ò�����fyNܱwk��nPB�	����Ա)(V��4�#.�M�,q�:����Z�ph�5�X�Z\��`��x�mY�4�!�A��#L�,~�;3[����i�J ��5��T�L�8 �5����d�J� ϘZ*�غ�	J¡R��-����gn���/�q�f1��<�j�c}��O�ר��e�~}uOj��@mz9� �U�]5�H���ا 
��i�(��+����
=������V��O��[��EQ��������5Ef(�W���p�1r�R�@��j�s����ho~($�:�a[�	`�^/��U�����Z���>�1��)N ���4�zS'L0���Q�kly-{t6Y[�����ǒ���N����@ڐ*	r)�,˽g'�� ��w�
�%��O�P����f�Q�!+������W�+����R��%�Y����7L~��Bc�`���p�"�7�/��m�HlT�-1w��\WB��B��Q�O��U4$�|o���q�Q�X���Ҭ�iIи����`��(]mY�C�ƀ�[�(;��t�R���EM����3{)���w%��zb=�`���Z�����G7*�6��-�)�5|D�(!��-�H�u���Q
B�X����x��� R�"/V�r�^ʤ-$#�N��pu"�ܛ&���|/@��+1�^*%;�weI�ǧ� �Z��,�0�$�(���������q������ �S����"K���XY������zgĕ�����k�'@��ĭ$���7r����O�>�_����X> ڙr�&��l�[��׹@�o�i9 �+��G`���%R� �a�d5ţ�D��q��rZO�?�9g��p��E��HK�Oi�uX�	=o�����B�%�\hD�ғ�{��#�^������PΈ���P�J���`Ұ��	�
�}�m:ӆ�ɵ>B>���"sM���]���*���B�}lF�s&��o� �;0�_邿��Xh�zJ|Y~y�5U�%�ְ�S�-(�{۝�;O�S���܅oK^��j���)�B��m$@�U�pM��o�0�Ű�8w��	�4���_�c	�,��ϱ�-�*U���� �� I�� S[�r�\_���}�pǱ=�����Wf׀�����[PS�ˮE��X�}��x�,�b�%�h���f'=�L�!�
'ڢ0�Θ���,�ES]2 ��p)$6C�'��&|.�@�#�N��ZK�8��/_�N�Un�W�w�יE:�B����Pp�P'TXԻ�1�'E�����e ���:F0�*���4�T"�NCkWy���l"*󯕘��=�А*�fG�]o���#@2(5#�K��,�a1���!~���SU�WA��+�|���%���mn��}�n?���c�A���CS�)�d*��_ȉ�ï�0:O�*V��(���p�+�p)�[ �c-��x�AWv6���܂mMT��qP��!W��F�WE��Ъ�X�K֨��S�?p���(�w&O�['!�|�q�G=O�Y|� �����/��$�?%�P�����0~��_A�������UNX�4��	G����'ˬ�u"w�>F6>2�Z��J��а�? �'A��J��AFX��zy'�( @�kiZd�~+�̨gUz0��B�Wo�/VP��.��~)�^�Aym�Wi�a���Bj�?�%���d�����T!�����P� Q���0�Y���BP�P Y�$�����FB�;�\���X���*=��<�����H	�Y�@�B J�����*a���&�(��sׇMIӋ�Qr^�W#�1���1��$8��~z��uL����곀{>�!�	���U5���\B�h�V�bΔA�cq�O}-C�c��7����[ �
b:���_�u*����<�ů���ٽ�6��1C)�`��-L��O���:�-	`#�f��	2t�X�J�e\����a�0�*��,[o� P��SR���Z�*(����g���4X��,A�{!�<���D�Yrq�
�m��	��[�@�%t,�> ��ƾ՝w�����Q�!��4��~��˪� s��W	
�0%TM�H:�%Rb��f�)�X��!7�a� �2YP������(�N��Z��������W�_�ZD�t�m(�U���(䮁.�~��	�k3��}O�E��](��%mW�
G^�<�~�H���&�O�`h�{(��P�����_.xY /^+�@�xI��K���Y�
��	HԘJ�}f�<L'��|�!CZr�j]l�������ݠ��93��o�1%۝�/��ikK����JX!��;� ���f��[����B��B!�X��sh�"H_�-�����	E�@�1	Z�)��s{fn� �h	\E�%���6,皕\��0�/���qiv�M,U�	�'Uq�R��}:� �*l )�URu�X��>��{H9�Df+�h!��h0�d�- Z����_)��{S]��Zw�l�-���<A �)N3u��%\�fP�8%���6P!G��#-T��-���P0�-�J$o�hM�4�E�^��O �V���f��'���K�E"z��_�@GZ� À>r��1�V�3+���uY�B�Bb�|M���'������ܽ���0r�J�菪���s�q��ko�>����b�(	Aۿq���sP��D_�\��j�	��m�K�����硙�������h�.�lY;�j, L,5U?�Lz}X� 1�]��<�,����~�|b�T����.�_�+F�l}%(�pp
�hoV�_I�r���uѶ�2zFY�(���C݀}ց�N8,M��!���6N6��R�.-~RY�+�o�@������LAB�T �I�<����P��hX;-�.�2��~�B�Pwh��]Mf�^��K.�NͽCb�w��]�J]`X�u�
ʀ�B�}|d��������B4���8k�)��?��Y��<��W��oa�,���	�f�ZȘ 1�4�U�m���8-�%�!~5 ���e;��%*��)��f}Ū[Z��]��R@'���n�hg����IY�P���d�Hf�K��J��-w@��}����
U�ٸ�X�%���T�g�IBW�n�Ը�zf\)|�(!F��B��=' �ue�K���X��,�6Rl�����r�Xt�#�Pz��SV	��w^���0�"��(y�*�D����d!d/�*�(��D���h��jȷ�%X.x�h�/���y�-@[�":��`+E��Pc�о	\dT�U��&L|T�1҇D���܂���i����|�Ȏ��J����?�k�~�Z4�.��[ s�?Y����^Z��/[����>" pН@lr�����bv�� ��$� �#��6t�C �gc��?@I0/���	[j(�Z��z�@`��	@�W	��z��i��"=$
W'���SxN�0'�o����ށ �ඣ��)�t���.i�D��rX\� F4�hIKD�-@�`��������懛ޡB�j�6�<X��^DQ��F�8�@�Z�u�C�����ʞ_i�Vz��w.�D�aFp+��$�n�=iOW�|a�� �Da��h fc� ������ַSL���c(
��� �/�� ���[�Η���U�!����IW��i�^��-0m�C����@�"jz�1Ϫ����@G?/%zU ��ͽ=	ݠ.� }_(AW���Ǘ������i�����k%�h������	>+~ �����U����h!���t.vNX`��Q��_�N���5�@@�P`��V�{H�%���I/��ᢥn��~$� ��v18H����B �*5��=�)�ܑS%�J��2�}��z��ȫs~��ɝ\)�n�P����,��e�E��A`/[��K`g�T����=�30p� npg��|�0�ͺ�u�C��_h��2�W������]z��й��H.�2K�s���X�?h,�yEeA�HtJ#��_*���9w�
�t'Iv�}M]g�J��yQ!�+�8yP	���ElW���K�U6#f[\�����y4h�J����e��	�)�1A&hNM0���@p�S�V+0�i�̞�9xr�K@�cP�-���Hd ��������p��O��sVo䒡w_P�����<#�&��6S����:�`�m%eq����UY���݀�����%�X-�.?)!�<%ve �dI��Qb�6z��|�#��)�Frp\�^�B1	��U�-ά��\-�G��؞�ԟt^b�d@��,��`x��!���@���V��^;��.��=�T2��6�N�~�Q�EY�����:�9J_Ȅ3��R��d�KI��
)�-h h��=[��
�)`c� ��.��'Q���R`ۣ1����A� .=�j��4�L�Ǝ	-:��Ѩ ���N���p*��)��O´b���!/@�@�x,1�)��B_4t ���iW�:���V+|S5R�6&O@��.j��!�UL���$��N��3��^cP�}&�PNX�3%Yv�1����O���)\UP��C�����UC�)~򋴫�2����H��C��R`d�6���h���U� ��}>a�1/Z�b	&B��`��,���~�U��Z�8!}�/9�i������
'��:�`V�/�sR �>*����� e�5^,W�
]�����ljP
�r�-J�"�)�5�:;��N�A�AA�W���z�-���X�߰��C_��J�>_Ö/�R�������2i.��I�. �1�$m�%�Y^���eP�~ ���O���K����9#5`��{^�3K~�NV��8�!��(� h��qX�J�Ƿ	x� W��'6s1�^_��e��n]��5.�%1	�)O �Dg@
H�D�w���f�o�������/Յ_��H��RK�_�s�pp�<i6 ���C��o^���� ��(_���/pB�˜���tX��yX��A� .�C�L��c+�2H��<���7�g�=E�Xj��)K�_kwght2�l�	^�C��^��L�	X�����&0�Xd�)�>U_��G(7��r[}Eۅ.����5�rV	�>5��!�1���h��Q����uT�-��ܙ�\l�/~ڊv��S`"Dh�*�N����������[~yR ��Cx�P~��9�H����ˇB�����}�����\��~K6�T��0�&�����ʕkʬE鬫����fo��YΉ�3$��1kV@S���.���)z�[Tgu�R�'�_�Z�5ࠁ�gM&����5�ǒ�^����OۻC\���V�9�?!2K��`A���l����Mq?1�RQ�t��Jô��!�G�1��Ɨ��1wK�	�M�����ym�5>���¨a"A�m�A�[�F�|�3��S�QI;��|=_�T�`�fF�v�5,��b���1����H��/�zP�T� R����k
>�)���{���	���Z�±ws@.@d������wj�^�B|_WVcV(>ۺ�o��т��`�Q�>�͜���c�Y������[^�X�O��E�f� �h�g�q�A�D���U��l��;��� J�h[��`EkCtl�����u!x��	�;���f�Q������\-��v�i Ki1l|�6��z��p��~ԠVYQ[q~+ �W�Fmo*�J�(`��`-R1�)ѷ����%'��!Bpr�k�������2���&�h�?W@�w`���.�1IK�i�Z˭^�� �E��z�~��UyT>)pB��tUV'h&���iw�lA鳊D��M�:�:�t��AS��~��M�� ����"�<��G����/'��1-,{j���o�m�経n���/��TTq\�{ʀ�u�B���j�*v)�6�$Q����C�u�:�9�m)�p�w��\Y����@��L)���z��(�JQ�j%��2�*Ԍ!��,@�1�S(�N�g��r�)��]=�:��S��bx�Pr����X�@��y� � .�'��re����[�Ňh�5�a.`��Y])o����M�8`asf�z�頄Ð���L�O�;��{���hd Z���������>��:+&; ��LP)���-eKz�5j�r1��3L�G')��68�H}�H�u5H�A*�]��p���a��{��ۻR��Y���P	@C$�ϓ"R٣� 	�X(�9��ʟ�^c��T����Du����N4 ��2M7�vJS �G}����2s0�H؜���eX}� ؾݷ����#L1�<��e�n�o� ��`Y��F������mO�Hz'�T�D�C*�%�]���v�
�6*�<\�E8�����ͯ��zd��G\&��^LF��[h3��=Sî9N~<�S�VH�+���h�.�-��R:�lP'�= �B�h/3�?ɸ/��-"o��wx�(#��\Rh	m��\�@iW��%����� ��Qp^V���T	���@�c���h�TV�b:��t�Z��~(�/1���O���U h�xcX5s�b ^1~�h �@��-�H �)�銃�ǅ���K��Jd�m� �]@_k�P�~�K�h�����i�6*�tHS�_)�q$��k�0�����s����6���
»����J(<7'�� ���r#1!�4d�;�vm�[�� �b^df
��F�a�j�����h��pl_���'�Xk`��Nj� �d��(� S������R �O����C���� ���7y�����W�������.')��uY�wT���L���4^�� ��p|-�$�J�w`��%r��`ғ/fTY	�YaJL�+����2ـ�-Q Z>���%|��������*N�9�|N�lx�!Ю�y{��/.B�}��UO8�}����b� �I�~�À_��Ut�n����(-Cy�c�Z�Q@�G -	7I@+����fQ����j���IzO]8�'Y}�s^CR���[�xAKZؘ���u��|(���"�����������E��Mܳ���T
|�-1��R�ht��1�	���	��� N
k�Z� p�ǹ���Mt�LO��X�B��_� B�:� SZ��R+�M ���HW�V�R	�_ sDnA�)K��U��b��	W�U�Ex)ɇY�
�%��F�.Q�):E�I�@�MWVQcdt�ݿ�^j ���TK�eKv~Tt�	�;R E��*J�_�4v��z%;�B�@4�媐)KŰL�'V���S+[#/�E�E�@��r0$�|��]�R�0���\"~�,����1���	�}�4����-.�����s�K��.yb��|Z��E3X�5pu�W����X�xe��
�"l� �\*��~�z�WK,�)I#\ 4[Z� Y���x\/m��s]�TK��g/�_^�QA�4)�]h&�}MgP��e��R�G|���S)ʝu�8�F�ـ �4�޵�q������`��*R0�1�vS'�މ-VV\�`�h�KY<-�Ƙ/;���TW����x�0�&�,��a�QԤ�W8��3e,:��9%�p	X]u߀��(^[�t��A�}!�:�ji�+��^uk�+F)�0 h�5�S�Yt�{5�O ����)1Oݱ�`��5�pMs�tϱ���n��"�o��q:4=2�N�8P]��u�����,���������1�L�J&QRh�HV���A���Uy�Dh��	��ј'xV��x	;��R��w���,96�?(X�L0�����wTk�p p�%���,|�#�쀖�}�,�k����k;�b�ŉ�����>/�qºP�1��h5L	}nܗlW���83�a��cq�{)��/����U{5��/C�(�bƘ�-��9�0BѲ�L�-Mp˵���h��%h㱺K�=�ۭJ���&D�ˎf��2�?���O���+��|��*<݀X�^%�!�V�0��&)H�D�9�^-���?g8r%M�p����5$F� ��7bd�ot�,b�I�E#���ܧ�!��f��q�Å�Jz�a�G`�9�]犌�� �Kv@-.�. ��I�z�$�����(�(3��:��р� �(�"�E]V�G�P$/v��ݥ&�xIPDY����~�`��}�Ld�`)"����3�K�[�O��Y��@~0��;�B��WP`�L�)��)^��H����:�4��� ���e[�^U@��nx]E%KCt0��s�;�JI �
��P1X+�@�&��G��Ծz���*��b<�Gk�#��xL?)���@����'�N\S!P �@��G.sL;K�^�<�����PhJ-�u���K�%Y�@ 0\�J �:��Ͷ�u�8=K��%8X������.�8��党��6X��C�(�8�fW�(�������GB�{�Ă{��1v�hs�D@��KqB��>�,���C'yZ
�^�2�� !\��) �uk�)%�d5I���Ղ(;XX���R}�NA|a�{|]\������/��!�B~1�x�h
������~a��c\	��1 j�3(X�x�bYl��P{�c_�įАn2{K=_͇�x93��{|���[�Q���(-NS�"�}[iĻKZ���]8B�h��� UhS�#�:&��ނN�	w	!\
�K��� �����.��X1U@�&3E�� �� MI]�	��8ğ��:>���e@H?�P�M:?yhsn]6�Ӱ�şU��+T	_�җ�3��dn$R9�]L'm%4��V��_�L�!	TJ��Ar�.����
KJS���~MN@�����>�����8��	޾D׮�W6��@��K���+J�dA�]飚C��DGS��*>��w\,@��rB?	;�_��˿�!�QfK�bY_T�k����	YQ��2�>��i��v��������B����u	� W_�(�8_��^����[����Om�� ������C����ߏ�t��(�N��������Lv���qD���H#$���V���'��(�ħ �#�m��V�i~Xe��CJ��}�E:�!�B;�h()��������@,Y%��%��'����?�|s�h��4x�� ��b���ߡ�a��gKiR5D�VOY��/�(8�Z\6R�;{_�z���81h-p�A]�Ւ�О����?����,����Iu━a*M0�ڶ8P�#Qo�*�k�	��^Zz?�:���w�oa�{Q�V�`�����_/S-�|څ\���K�^� ڵv������|������g�F��	w�5�(�<BNYy'	��-�w��.�� "?%6�����|����	]Vs�?O��"�tWg'f���'E�$>��p.�_H���Y�'b�Zh�Q^!�й����P�^��b{�6��{�2~�b!�.)�{�������h�m8��-xV�{�2Nn@��!�Su�D��3�ǥ׊�	�yV��_ ����sF$��q17��`%����
��.��"UEM�Ė�>�k�nn�8����- ��{��5�XW��2\0V_�0h�4�h��5��QS�`��XQ��]>������~����h#	����2�D)��=<�5�S�f$�4;<����P�?iX"꧅|�O
�l����1�ZP��(X��(�la�EvD�^�Q�}q��	 zEVh�7�+^Z�@a����cD�.e�!�Q$@�,c?�� ؽ8IF~K1�R�4�o Ő�Ήa�2������r����w/'�ncD��.xy1 @�	�B��@����!�P�_Ñ� h+k��%���D��Emz��C�l��H>z �q'OjP�%� ��sRC�h1	E���~ ��dt2��nr!ǚ`W5�BL�ì�Ը л8'�C�2��!ě��^�lM�]-�s��g.���E��e�� �!��lg��pl;C���@}@%�9�m�f4����x������L�E4�V�	�(�LM��/^ˀ �dmT{[��r��+�~��-�����	�6u
X��-�L�㕘�˯G[�@�p��7�Z��)N-�t �����-z�Ȇ�3U�<��?�r��a�*Ѕ½(=-�K��Ь�������Q��x-��@i���XEK���9����63O��/*3:U��1��� d�r��Z��id�h%�R�u�� �X#�Z��p	�]�Q��E�~�̲F0���U�-x$N�p��2��l	uI��!3����"�-_p)h�b�x�Â�a���D�(s��#�H��v����x�_u�jWB����)�Jݤ����� 3�	�������V`CE�R���\Hj?�P1	�M���bX'r~J��5�[f��W�:{��ԬAw���J6noY��,A�®�J!L��`�^���rdz��,������C�g�M�"#�!�Ї��.	�V@.2�&��l��-�nFa2�fƀ�1�)ۘ8�װ ��%?�@@�������~��:�#r���:�<��Ύ(-�X��\*�k[���(*xj�����Y&`�?[8�hR�#����Β��8]!��FR/����e��Vw8�weK��؁�*Z���/h���<3P�\=9�Y�%0@�������vU��p�5����έR����l�'�%)��H(<X=�[����:�4H�͏9�u
���&°�i�@�8s-�����	+I�X	�?)lW(I �2�Z�`D.��-��"C��6 ՕQ�h���;(�>�}���P˰�f��� GYg�-��`�ܟy�g�����廲ߨ�F�5��S���
v�&l;~]tJe���P��� ��K?Zh #=�A/�Qi`-�xKtz.SZu��W�H`J.	A3��1�w�<�d�p{N\����_���<Q�~H�(M~@��i}�� ��@k��u��Q��G�'�i8�xmP�cQ	�j�q!��<�%�LF�#��e[��j������=��� ���jg?)���z7*Ha�(��-0>U��U_�>��V�r9�N��|�YX%���=�h�߂�)�@�1�P[%�YOk{�>�; w(�s��Z#��q�n�������-�\�� ~��:�HK<9&N ��E�m�s	I��#w�XH�8�[�l�K{� �����p��4���q�ʉ��Q�8B=X_�{�7{
(�`�J�S��#��� �BiD1����}I���%�+�������'�p`� ���h�^?'M�A���Ơ{Y�=�V�ğ�� �Sl��检�^�#Y +��V������u/���� �"�9Nw�	w�����h)�d��D��cҩA�Z]`��l�}cY��G4m�ca�/�E��/��Q�`�+9�^k��� �� A��f"qH�4���`���AqD�����4QF@b]�	>
�?P$�y(���>��/�##�K�e�� fn�K{2"5��"�Y��'T.-�&�ù�_Cx4��"p��q�<u���j�:*�)�Zl�>�/R��X���S�SaRh��I(]E�������.�%8�p���Iu�I2��l�h��'^	���Ad�dP�q[����pB$(��ݧ0w?�:�@R%�	{�1Ѐ������10�zX�:%H$�1���� H�U�.3�O�\	���WF*�Z�	��]˛��}
^SW��jL�Y�'��}�m4��f��m����(J����U�k�{��!^D�j�WM	vhO届)�nK}�F6�~�|�)��O���_]����*�!�˓-R_��d0�w��K
PTh-�:�}aTh�l-[X�
=M��<"P�W�@\K�Q"�k��#3��UW`�]1��ݗCs��U�=��G�/5.[��3�M��H����d_�@�� n<Im�G[\5�c5!�j� Sڻ��L�(�� �Wr2Ph�	ȹ�s�'Rf�;���j����^�%q�w��s��wF눚�l]�}/sMЂ	�ROIʟS�F (��JK�'�	7=cm��b6W'v�[�
C�.�v��1�k�w(�9ф�a���X_�&� ��4�T�d�3o��)��u��:�(�x>����0�+��h`�kn�-��x�-��i��j�d�MW+�E�9|��!��r���ȭN�!�������P�m���g&Wa�R�+�70��NK�����	h�NDE��|J<����`D�L�(��V�휀�)�h&g6�l� %�XrP��[���	��^V���z3��lr;����U�R��]�k�Q�$?˸/L��6�ٻr�������i���/_��"����u ���D���Ru�t��Y)^}�xp9����W ��6�1��1!�?��	�|'@5|�`>�Qh�6'�,��O������Y8���U��	�i��X֥(��ɬNP��0�e�	�X�h����_y\�*���T]�4��������O���w��Q� d�fh�>'�o��n�T��tu������I}<	:]��|�%�5��RɕZV5��h3s��'X�m[wr�Lo�u����B�q��VT^/2X���0]hy"���'W��o����,��y�:��Z���xm��$�D����h�H��L�SATR���P�x'*�ė��^,����C�ày���OP�NiV��G�c)�d|��4U�ͻ���|) ��~��o%�� \c�F5f�Y�)���'�x�;�T6,�p�i��uE�s����X~��@Fh�0?4��cM�w�k�M[�])���,O�d�P��	��E��[������9���I�ק���Y�1����_�GZ�I�]gtc��d�'�|T����R�,h(��a��/��#�l�:�L��>��r	�q^|D�x�2�U����ꌰ�(��@��H�
�3o`4Z��!,G ���AJX�j�Y�������XN��ZNQdx�����Ք(�֑�Eʿ���@P�{�4g%!���>�+�-���0ϑ�D���� ��'�4�]P�=�����܂%�0�F�^	���9�Le)��$τ4��7Ӿ��Hu��\�*?~/Z �oi�`�X�R��AA$Lu@�0��:����W��;D;�
�*� &�����Z�0��&{'`�K���i>}�W8���*����^�d(b��E���O��)��u�QNJ�؆~�,T�@�g�81ջ]:��>�&.�a]K�����Q��*�D?�Œ����F��L�0 ";��7��(g���[��y�����'��#*�K�n�/���8�tWx���h`���f����Ux,�ku�w�@L�z($��^ÿ �RY}F!�]�W�O���[���b_2���b��R�cE�G�t[��?3�YD��f�����
k�x(z���$��.nɁ��"��u�E���L"ee���8cR �u"
0���&�Ϡ%W����aha
n1��8XY/@X(�牥^`Ùi�� 14�&��-���%/3j���9���@�P���U�X�-&h��u-T�P~,."�Y�0�n'��g�R�[�i	~�6�%	�!��Qx�b��c]u{C���z��ە�)�h�L�o�F�_��� �Z%�UG_EY��h+���Z��Bv���u���H���������hY ���BCu�Xc���У��u�P&�MLx1+�\y)Q�Á3 [�7z��8�.	W��.q�����&���w|?E�ƹ�8>MK�p��Z\!��r7l@�%,6�f{EKR��������}�@O�^P���Y yR����0S����������������þ(�[�*�0�R�()8ם�6# �.�Q��M������K՝�+�`���LJ9s:�_��Z�[�!W �Z_X���C)��o�1���@\�IlCh;?�?��7�pa-d�����'X�	1�)�	���I�RxRNu2�U����U� Z@�`1���~�vz�ڨv���h��I�5Z¹	�_�FXhy�Q��j>�4$���錹B�uF���0��/�PX5M�W過��t�J:������@ ��kl ��E�5��T� �
��ڂ��} _H7{EAq����XU�d���L_�K��^�"�V���M�@J�r��[����h0��%�6�u�+�2��@*�^��$K�%���P}N�h�&����'kՊ�T�nF2����q��.<�ca+��:
������`Ҹ�	B�!T��N��Cr锼J�����{�E�V0&����\�@�.D�����¼u�/,Q��D�;nN�����@m0:�餠$ �6k���%�n	�� Zt�&��L�r%o4iiVB�R���TZ��4�����hK	|�]�YIMC�(�6Hj�y�)pݸ������bH�F(6	hnCQ��	 2?��m�/'�����fx��(I����@�]R�qM%�*I�ܘ�[��ٵ�ӲDD����Y^+WO�a��2�YiԂ}��Th@���P�������0�g�(��I^Sg���!��>�x��тd���/����NJ�CB��猖��S �~+���Ԑ	���,�8�"_���@�[�(���b0�^qkL��D�2��� ���,�a�Ӡc�5-)� ���}�,���o�,V��i���<�	�1�{°��^\	@�?��\�R�C�e
���	����H�_5%�M�(�b��n�ȇ���`���s3��A��X���r�p�<�6�`�)�QJR��0�b�B�Uţ@5�90X~���� F�&�adl8ws�Ͳ�\0���?$�u;������������^�A`k��P�BQ��.�H}-�/
E�0�-��Ћ��_0�+�r�Z7AzA0M+�r�
�FSL�� �1�8(�I� �-W<���z�1� ����v�\K�<��?��"����Ј Q3�?�8�����gUÅG.\^���w	mH�K� ЗTG,)���]#�*���|V ���U�	��>z3�s`�� ��Ȼ\<ր��a�=�@ۼ�z:�����_���V��q�X_O�0L�)
��������j�l!�[|0X��O��	��B���P	�2��U[!�:ؑ���J�v�n@c�/=�ݗ�����uFt�I�@-��TV�	�=��f|z�w�[I�A��i!��)�`G�JT���-�A""(U�������	dG�� �r��;�[b.�dP�l�W�1�$�sxB�H+å�:����Ȼ�Vp�����.4�Ol���B��
��u��BJ ���͉`�w]b�^lW�c��6���PC�-�)Ӫ쫀h�n�e�@/�
�%��۸O0�Gv�����{D�ٵ���s�����h�bO]Q3�U��]V|b�<��i���d�%`]8�!ݺ�0�B�I8	-���A��RP=���v����I�A��W�5�\\R��B����@��6�1|$�g@Kb;�����%�<)yx�`+�,T�[N�|X!hf/vvIV���UShcB&`{�R�O��D��)�ߝ���Z�������Ӿ����Kp�H��b'~����
P{���v��Xb\w` fZ[pM�W�Oz��1�90(���I����Ml<!��J@�%@ �+��܎Q�w`)�_!ȪdX��$�JЖf�Ț�@(�Ӟ�%]��BN�$��� -,�ZLM�5��(&��Z��"��	J}vEn�k��Y[�9d��\(�X�E���YS���wl̀�w���hu�g���N'����@Pܘ�hx��Z�K���{$G�5�',E��;&|��5Z����(&�� A4��������Q^���B#�r��0���	ebR" ��I�v���%���@�=$lN8�z �~	*W��@z,U:tX:f��Q',k[���i�)��J=��⓱�!>FE��ZR��HB��������3H#�<w�,�������b6]֝�ΰ���m�����h	����&+m�����Ը�;
D1о�<�?@)�f%B&_`����Ea���vM�ڿ�����T��yPU�J����`�Y���*4$]��a����Ҡ�:� D�x��Ă�Ez0�`�HS�)��	�ȽR!/�X���pp�e'�a��_�h:���i�Ä<�!��f���<z%8�S� Y-Df7h�Qï�|­;��_V:B��}\�B��^P��Nn��{!�LHDV�_��y2JM>�BA����D�/tZ��- ����kT�_�EpRҀ���>��+Q^@5��c����D�5��d.N;w^H= �D#�IA�8���A)��<*��.��qgo؀��(�9u�k��p��}��9�[,����kQUX��3�L���u	�x��읃�[
�uk�K���1���q"=7E/ھ,1�w�F�`�XP���Is�oN�YU��r�>9)�N���UW�k�N�@�gV�
�АB�7XH&�
Ch�Y�Qp.y��HX��'���z	c3N\���}���E�\�&��
�9�- W�&=:'ݡ�{M>�8�����x&9��!����x��'��
4�,({�E�� ���rA��|$]>,؇�@i���U�t�!)�P뉉�u�b���hfg|����Aaa;���#�' �p*A�X�q�To%0і�:f�1ҙ^��H	����%!�t��t���ΉO�Lh�j쵏P!�f�_>�T�k�-��|~u ���5�!UG�-9[����$��a����p,��0�f���}��|�`���@(��+��P�S���Q�T,.��
p��f3��u$P�Y��^����6%��>�J�h|Tx�� "7O��/ԣ'���{���a����1��@�����n鑢��]h�K��x��l)�O�/A��H�/1>0mI|N�?���D�t��0��+3e�b��Pʀ2�ZA~��[>�����ķ��^��v|?�Q��&�˹B����~{/�K���&:��'��L��pvLH�^�cX"�/��Xj�h���.�Ŋ�1H���ah78�oFo��[2
Z��A1{��O����[;`c��H���<���`�^�u	��O�A�S� ~���$��T[�Y@�ޙ���/M"ȁ�Q��q��~���/!������j��N/�z��b�M1� �=���`*"�@���$�tS$�)Ձa@wn���\�j�_��� f[��W����Q҈A���*�\�8�9��f�t��n�h�Q�1`&�0�Z� ��r3�A�����w��e��a���2A2��SW���ӥRhz=�x"��Sԧ_D������ݜ�?�1N�~ y�梟`̮].�1� �["c-�e7Z�|�U�	f��Q:	d{ ���P� ���8�ݝ��'`�:-��r��(���%fZ~؋�~�
�H�-.q8���7Q�Jh��t�?�D��
�3��-M�Ӷ������U<a��h�G�QX��x@��SCՂ=��3�>�fxWAl�@[��D�Z��{�7gM��yu����X^<��\_hS	7L] ~�r&4K!��*���xz;��N���,��k= XB&
!��"���\Q>�8P�)�T���JLlzg[ד�O[�,U�8B+^�4U��� �[���Kg����|i����'��������Ŕ��ٔ~�́��;1�)��I�K��@�0��nd�ıXmsb#� WO�B����F!![|�Q�-��^����$�&&�D}TPUᱳ�2h�'�����&�r �\^_�
[��P�-04�"5F)A
Ö��,���S��ȃ��A[ ��<(y��i2?z�h5o;��%U��AG'��)��}����1�=%q<O_�����)� �&uh"�0�#�u�wIe[ZWR��Y��O}jZ�>�� ��(���'a��0Y�[ ��h���"�7t�./Kh�)V	�m�6UۆA�>� �V%�1���Zn;3���"���«��K�IN�� ��-�9��\�z t/u(��߻M�G\k�dn�Ȥ�R�zP-�)�,�q��H��N�����@r�1�:��ؠ�-y�tP�0���Z�%͏h�/Q��(�Y6��f����4�������=#����h�Tՙ` ��[�\)���X�����	!B�6PXy3az~��m�	��bfi)Ո&Y �^��|�aim�n��(\M����-�󮭗,3�����t������B_�+,��7�f1�.��Oe���S)���
@ �3;=���V�0�������M�Ժ �����>^�÷���3�4D@�V�K��t�)��@�qu�"���)Ӑl@t<�~iS��_^�o�o�G�B#9�A|1/�һ�4φSI�L
 �
�P�]�$L���&u�:N��t*S"4�А(2���J��%�hxqm S�k5-�j
׎5�Y|`�e/P鄦��<1(�]� bS�C�j�.��>��0�j�,�.�-�w�f�X�ٔ��e������;\��id�NP̒�g_��Y�8��:��P��֫0�-(t&Yޠ|3'�vv'�}`�0L�0�n�-�g'|��>�j�vyzN��R�B���*@WF�b ��va�/���J/�gQ��J�z�cT���H19є�y��4RN)�Y�>XULB��� r	��{J�v�W��� � �ws�4�����5٠ቪ{�`O�D!��.I�O�E��o� 1^���b �ۢ�%q���[R��a�C됦�\H?h[�ƶ,X�r	BZ���9���
���ក��0�/��8R��(�Z�c6���K@�������h�3�G[��jM:�ζ���n~B�3
��*�`;fP�Q��ͅ��f�>��)�C�q��\>�xn��#��m�k�yP�r@�)����"����� ��%#/$I��8jv��"�2<!�y��JN�������K�&�0��u�Z1�N���W�W<8�cC-���=S��*t�(��0�S�/0���̀����`�`�i~��Y�n��0w�F�4r��(�v���E�%^4�CD\�����h/pN�u���̮��Y_�*����0{���k�g��L!�1�h"z�3�b|���u pWX�Ni�/O�|<l��;h*T1(z��zlD|#齧�W�%}f��!$ؖ2MM��1ͻ�)t�_l(%�]_�r�yr}�[���� �K�%�(q��N���b;_���*,��&�H3��Z�)J���飀�P�	�	�U\p'����%Hh�ң�@*?RV	E�����ũ�@N껢4�5��`0aT�^�.��*7v����9��S�!v1��*�ZQ�`[�3�� �=g�j�╀W>2y�ܸk�(�5���@7�~ ��\�hRX���@_.���O��X�˒���m�z������\�W8�&�N��h9�@�Ҁt�C��[ߡFP2�ݿ�5��3-K��c: ��0X�-�Чi����>f[y��D�eZ,�pl������9"_a�G���.%&5����/��k�	_@�N�}?����[g��^��~y�c��GL^�_�˔W�o��&!|��U��^.�n��	1�Y]H���B�!%U�̊h�\A&YD@-�G�
���8�,߮C��^����Ү��JE�3Z�Q;�	a�t��$+9��D�]��>����d��� ��Ƶ�s���ȇi(��zQ�l0�Y`�fh �$ܷ(��%}OR��
>��?>�4�[{�'�Rjl�����z�	1i	���\�U/b^�	XS  BL!)�u�9s�B�0��	��V�	��+��X!A]����h#c'fX��}5����*P��!�_�(.��}��)������[�W(EH��Y-�.}� �貏����Ҡ���㠕R!?T�砕_��X3Q^��
�e�4��T�R����%,�z�s@)�0[���ۉ�ޕ�}iN"wv/%��W���yn�n �P~( �`-��Kk��I��j�	��H�0	������� ����A��Ѡ��_(�B�7d�:@���D�0O�P[4j���E��/��_�O9<��,Z�XA�0~�ݜ��wv���E�R�%t��2�S�:]�n(R��"e���v����[�����nɸ@D�o�^E����^����<�Hۙ�d��h	������Ĕ����b%Ķ'��RQ-!ȡ�H�ώk^����pZgس� X�e`�(�X�2�v�uQQa���~�	*���Y,*Z�є<.!:o9�Ae#j��j��d�hQ��~���Z�]%��d?�|!Zi�@5>�J�������?�����k�������ڄ�N�E��1�;� g���]_$���H��Z���q�L�(����8���C�dfR�
���q�ϻ�B0 ��U��*1�½1�n�6�$q��1��A�YRr�� �0LYTfe<@��$p�/�<H��O�.K�0(^9Q;)�WhD%��sW�h��}N�'�s�}O+��	�x˱�Q�c�%���V�jA	Q[_L�NR�v���p��W�����z�d��|O0�&��['(W����S�n�oAy]H��L%.I�M&��� h�\�1]���`�NV�CA��pb�{�%g��Ln��(�ޯ��^�:�N�Zг���N�%�3 [`2��=+0�P�3�P���q��9�,�oR?ݺ.02 �ca"���?����O2�$o��o�R�0`��O����F�L����`L/��A`%��~�� �#0��zSEN�WD���8,��)���:&�_�@��u��1!�h�Ҿ0R�U�S�rP5f��	J�	.\�S�0p��K
��
J�'���|������[󸴨h8IAp�n�u6{b)�X�A����֙�h-�`��P��/I���a�����0�y|;%�	A�/u�g��ӒO�[g(w�=�$C�vl��������ڍ9��P��p��;��G����q�iW�!�����Rh��HF��*�0|���0�4�-?<S,a4n��/mD)pU�Q�(|e��T�ʐ:]	%�����X�M:�0d
�;|��4���Q<�5O���)+!�nm��[��������iA��jlB�=��'�x��y�zx` �s4�������/�����P%h^�i�(zuv�-��)U��)��%Z4Go9͞�zO�� vu>R	_�`�G��eT$7Qcņh���X�LjMW��22�`��F�){LvC ����)� ��I�o���Mj�>,���?}^wZ��(JD�P�{��f�v}�j,���:)�6-}�np�9�8�;�~t�IC��
�[@�piT��3�+��|�-�4`85�?j�H�H��[ީR��	�\8,Q)$S��&X}���PWy��-��3�!����}0 P�iV�`�ka����b)��2x։��@�
o�g0�����t.Р�Fmu��hBhi>'|2�W�Guɓ>_5�2�@MPS�s)��q��y5J� c�IE
���)n�_R�94��`c����[�R����V���������.��O�JB�"�Oŗ7��t�����!��a.0�=^��	L(+��KS[,�C� W��jq)-�_���U�"��/�8ӷCu�Z����H�)��oiyB]�O�ߵ�n��u%��(�n���TT�,de�І.=q`�$Szr���~@:g!��#`:��%��αI�K�N��K�ф(�0�?�@0Y{�US�) ��X���NI�x�2FU�[݁��Ԁմ��(�_�h+"���,���Rwd'���.p-��^��pZ[��&�@�w��XYIZ��?����5�Z:P�x�z�!^���� Hl]+�=�V�%J�0 �_��&�iXC9'b� g�[��?.�|�W�i�Y0���?0*$��(H.`iN02	����f�����Mn4�����2
�K�$>�RԪ概<��]��&���	��b>�p������D�w�룂���z��5L�VO�Vf^���n�]�@���Fqb����1p����4���N���S���ـ�8�u�B&�4�t�qy,��mU�@�<�Q�
V�*� ��Dri��?mo:"y%v@�� ����r��,u�0)��
7\ �
�	#��Wn꽮�X8�&tTO��[�R4g�.�5�) �@-�x��:��= ��������]@�EYFvS�a=�P���v��;�J����?�����,'����(X�f,NP�_8mX��S;���+�)�h3����,�B�Uhb�[d�:�ʂ��ys7k����}z�ch��B>�G�s/�!��e��u��u���f�w�]P �#�!B ��tT I���;
d���0��k����>w���y�� �%s�<�+'.�F�5C����Dv	t+(/�Ҁ���{�������׉� �)s'v���	����-;r�{(!��:}<%�����v�V��@�l��F���l1�X�.Kc�1�r���(h��JR��T�������Q��0�Y�h=���,���@���w�a��{����
qA��=VW��x�Ҩ���)������&Iu�}�hUq�hX�P8�i�w�����(�1Y�)pz����y[��G����~O�=�+����>��[��0��o{
� ���ߟ�K?����U��r^Z����g`޿Ȩ�1�y�S�!Zȭ��٪J�b�SS���duZ&=�m��q���7�B�y�%/��.�װh�9�/�v��zB� ���	}��"����+�8%�E�U��.�y	����_��'�eQ�[���+���q2���fUS�F�V�[r�9"8�����IF�� �J��G��.in:��h.`�f�>�5�@��D �'�U��p��� A����R�v�v�7���I@wܗ�Z��)�nŮo3B��*�'$�{H�_K`\�9: Г��aiF*݀�fh�4���m-n���j�*��w���{\Ba�b�X���o�{��Ӿ�������eq]l�8�31v[l1�>���
�x�~!�]�u��)�&M�P��Y�οa��}i�U��� �8�qoU?����~�pA�_(�Z8�~�^K���~{-��$R��GK'w�I'�ї��VSm`��_�}����п�\Sg^�jv����F�ԯ�,>���)Vt:߄���g�`6�IW�[��[��V:?H;�θ�ܟ:�
VT'��Y�(�q�T��v3,T�#Z�E�*o W8���[��J�Ǻ�Qh*��>�_Hs�0�O2X�Gx��pܿc��r��?�����:�|
L&�[�:m	V�+!���1����. 7%6At�/�w�ͩK�/[�ӌ*C�6UL�����^�n����Wr5����~H
�?	S�⽐`�^��>>��u ,�|_Th�|�.W\+0���-� :�z*G�SV�	)��H�=�<:9�p���W�����L�^���W$��1�[\tdU�ZP��D�V�������3�2���.�K S��Y�N��r�F!j�����<��2�h��.��Q��`�KN)��ұ^�:I_�|�%���*�����Cd;_�l$]�� ��[��<fR2�2w���>����Y�����P��k�w�nE�9/� *���	(��E\�[��@S��lQ�N/��g��5�2��"�4�?.�,�&a.P��C�/u\3O��+ѡė�Q,/���x�p��vR��<������(�0� Z�?tl_0��;K)(��c�x��.�����^�"���	���u`� %�2ؔ+ZM���T����g��P���$2�/$��! |�,1+�n������+��0g��"GS#P;f��<�5H�	¬d"l�+`� pʽPf��߯+$��N��J�5���8�'%z5�"hs^%�	J��٪*�%J��ျ�#iW�jF�v��>!e��E�ԕ-�l��}S�~�A �L�.^[���y�R�j1i�!1�Y"�	'u��� �M�������T1ۓ����18bc )�����{m`�6Xr�pk0��޽�Gz")��@�()��5?����4�1�g��X�>-�L���z�y� ���'.)O8.����s�]x<Ӿ�y�j1���;�5-X�1J�A�Z�kǶ����?�gL`9�3���;�*q���,M`���?���J��-��ܵxPh�7�-Z��@%�G����~�'�"�;�Z'aը���G�i�{J�.#��v�-\ġ������*��� 	~gU�2-�l ����B��a-,�/Y��¨7���eO'���B�]��\� �U�q�O�Kr�+�Ӿ�V�q�-t@�H���2�(P_�4ɛ䕯���k�_�;h~LH?P�%2��X�0�t�P����(��+���h�G1���!{�}Q �tKY�_���!nN	hR?��Q��Sɜ1�fP5�4g�R��8��	_$����A�&��hb�5d�EMz���X���-�(��ς4B����4P#�n=���N-�Z�V���	{�̨�6�0�Z��\��ID����J�؝h�1���l��Gf�V�D%X�q���qd\��Z�!:�*�+����K=_�� �h0�|�Y�
�3��$G��ݠ�F_��n���Yv6���1^ո�[�x�-	�vo��/����v�}>ʼ��rh�OF/�b�VG
��((�@H���%t�̺����<@��G4��*)rz� �{(Ґ�zP��k	?����}��j)u�F6|�XC��D�_���QO��sr?�����R0�'��B+�2N�h,t4��u��Z]	h�C^GZ�c����D-}�2}-�]	(0Wfh:DUI8.�"�R��}g?�s`�B � ��C��R�AJ1{��oN6?����S�c1�O�F����������c����4�d�.#Y}&��E%c����}�w�S����N��3�jy5$sA�X�D�I�v����Z���{[�b+\|����R�qV/@�l�_C�q'�}E�^�*�W�'Ñ���Z��e� <uZ��f��G#�vhO]���r-��v׬Es��NX&%_��&�}u�Yh-\Gf9.�D{/t�XW��L:��d��__0hkTbRP���)������Ģ]�G��9S����"+��Ghn:���������=���sv�	o�	�_3�,_h%	f�
�
�D�y�ZP�ԣO�T���v	��Խ��-��I$+!��6�1��3^�I�p �\8hsgb�'�+�{�eZ�B��y����â z��NF^5�!sU��?���fx�����~u-ݳ���l>H
�-UBbzQ����%��L�b!�Tk������H%��$&��:zH�Qv|
%�� 򻈥/G�����h-wN� ƫ{�_l�Դ��Մ�����%� 7��@
����y����<1�@�dQ)�Z �����fH n�~,O9�� �r$5�j4,g("�*8E`��si��)�~��n��UI^��?��,?+�\�ezG ��3���bBWk뀁�F�H%�rx��|�V�,�Ip��)�`��_	W�;,`(�sqJ�@w�Y~��	�`�2wl� 	6�
�Fn<��!�1�eES���e킯Fq��w�^�L=�X/Y�'�Q%86B����\�W����B�J�{;�@��@�����KX��~tTI��!|g����U�%�����W��\�8�M�聆���� گ�)Ph"%Z@�|���ؾ̀���_�%�xw; {,luO�HJn9��)������xd\��䬸P�k��H��'ZR�7;O"f~�P<����tQtba��hR��)})!��^/�&У��p� ~3X��q�V5�S�����H��̬���AL1�_�8��]�/����d��C�Ho����W�-s���p,��������r�ؐW��J0�[ �qQ�y�#��s���V�o��g��'�Z8�J���o@źp���H=���c1�^7��W!��fM|h]Nz������H�d,���i��v�J�6��v �x�SE%U3��)��?Y���v���s@H�50~�|�s��+��-�ʓ]��O���G�%_��	�Y��xq���/�}׭B�)Y[�ܧW��]�We%%�o	=x�5f�1�K"�|`\S�L��=:��[�u��3�YA�&�
h� �c��Ԯ�?�%	�E�80�x��ܟB�C�24 ���^H�\ ������w�r��D���"� �������B��}p� &5�T[҉���nfz�a`scZE� בKL�@)b�,��	�+���/�-
��.�,�Z�N:bfm��[����2�F�b?�%��Q|7��4Oz\Px�R��}_ZE�o �5�`���!�S �d�a��Ll4\�u�\��>i��~Q�E>I}�>�����œmB����;� Y�#�	I�[A7�* ����	���X��t�d� R�{�(�<R�~}�41�-w^8��-��~�/c"} �h�C���1HZ��?0��M-^	�g�X9L������	G��rMh�~�n��<P
.	#t��>k8_�ni\)�P-Z�V`<_���q9�Y{���BhnV"d�p_�Db��հ;�mҘ�Dw�D���'�$�'0 M���u�/���ї y�]7�\�4 �z�)!�^ ��/+�=�J Gx-�&ˋ�F�1�!��1a��D�w�f���W�}� �6�S�x"�Z�GH�M�����E�D𞺺�`�O{U��%�	�r�L<�R���_Vf�/Zf)�G����Ί�����~�&��4��0RB)ՙC�E��F�0Z]���JO�!����~��!��� 0�Z��[��)W8Z��	A�;��,�jVP	� ^�RFN���'���tH��2�3}�|@q��fhEDҐ��+���?�0 � -i;�*�rT/5�v^�P�-�}w�(J�����;�{��T�*1l�@�)������A�\���� 	�ǉ� Ec^�)�5��3&�d��R�v���K@L�$�,��s*�����1�JZ�i�UwIt�@��QJ�K%ӗ^���J���p��,4�%%�_��-^�Y��^�ߖ��T鴭��9|U�x�=_����l�1	��&x�fS��9��8�=� [ �0��^�׺ xlJ��E����N�H���/�޹��B}I�e4/�"��g�IzO��,�	j%Z뭀\.U��L� J�h�M�Xc��a-�D�W�)Ohe�'&�q�F�ؾ5����O[2��L���;UB |>�J�0�IVe��gˁ=�: V���1�`�صF���	�tP���@���[]��a���~nBגqt�\�b�N�T��[��d:}	[�I��E��nX5B�:&C �aXRh@�a������p~S�d��ٝU���䆝u�z�����N�R�F ����B r�<q^Z��l,���~�U�=
0K��K�E�=3�1y� [�����v�:"���UCe�Kb�;��h�=����,�!� �6Uh_�.�kw�O�10O�ĉ���\�C�:�G�J��v	鸤�嵋�_��Wp�KJ�M�2Io�(*�P�����Y��9t(�u��1y���= ������F��W��J����p����<�F4,�Yy���M��s�5�C�5-~�#ι�/A�"&�n0��x�TTTd������� "q� �������vs�[�C��Z�6W�y:�u�U �+���py�Ԝ�q�G��c�k [�tT�LE�7���S�k ��}�[�����V�r�2��.`�=�Z�p� Y��!�|(έ�,v#+)�hs� c�XS�9�P����TZ��������R���ĩ�][��F��T)��B�B�U��į.�#h��*�U���p���-^	����K �����ր�X<u��p�so	v�'ݘ�U� �r�W�����s�h!�`�,4JܞŎp���Y:$U)���|����t	Rw�H�s͠���Я�cק�����,P%��z��ʔ��R��~�l3V�?1w"`�6I �S����n&�u 05�)�T���(z�-�`w�G&
-�.�B[�l��r�O&֖��$��o�Eђ ��6��Zr�n�3
u|_T�)�����d�M0��	3T����?���$]@[Ph�Y�t�g�`��y�Ka'!���"�A2G{ e�-,h=��쮸 cG�y%JW�Z/�T YrlH�� 5�U8��L�L�/�x�p)KF��8�_��B��vj��]!���UNѣ�Dk������j��}y�'�Bs����zE&�I��!�n�-�\�����t���] }����\��^�Nos-Y��%;����]�`P�r0½^;�!�$�8~dOq�\��VW��X`��_j���pa,^z���~��C��M������R�6m� ��QP�s-�'xj �Q�r��#��� �*=t[�{��I��)@��#R!�qar?����3�ڂ��	y�1>.��;}N�x��%3���:���1ߧo<�^�IwX1���ڎt+DU��*��B�ռ��[��Y��������Te(]��$����%����HM ��xV1��[g=�_���R4)N��D>��!��r�r�S�\��\ҿ��e+�ʁ̏�`��/)�Y����s���1^@�T�3�0�F���g�	�fN���U�+V�	KL���g�����S���gC�4�o��]��߁v|�$��L'I�h&^�����<j�`�ɷ�w{5d^�,8)v�>��N�\(�V��L �e�w��,�O�}�
�tGjXx{�)Β3�)o仦.l�U�_,�0���?U��I�����{E6b��w�Q���+���!��:�[ʽ���L�Vp;L��UH�Qh-1��5�9z�XA�- ;|��8�>`qXY�J�u�]�j��h7&
"
������D�g����H[�m'Zp�u2dS%F�95�?�E�t�G��mZwk����vC��]uxJ{��f
1�1%,�v/�� �'/�S��^;�Uhl���th�Y���������	��S�G�!�|o��4w�0~�@!hK3�H	B1�ǹ����-�L���fS��������h���Ц"��B]�-��	���ӭ��Q�z��y��Q��z������֖\�v[7����Z�����c�K���:�i��$6d̑������|�v$b�wN�(v���Eӂ�&�#B�`">����� ��(Q9M?�����ɅKz����5�;���b�t��3�� ��VD�	�x~XKL��u�^���ti|L�M��S���U�=\]��/�O	��):�A�҂� �Q�.i�JyC{���:pd	0H�LP�_�T����(X�L�-��s���F�	d}`;�����qyba81@�a>��Bp�eǪr���E聽�6�{0�pb�B�`��E@��	�e�_wq�/���^1ÜUw;���O'i���-�8������ ��t\`>g!��_-��	1+�we[��q{8�	h�=�ԌvfK��\��pwoU��/Pg��1�_@�G�Ҹ������Ic6�1�- *9Hcl@oe@$��ſ��`��I{���7�1Ԧ ��ē��?�]��z�)Y}H��f$�7=������y�)Z�k��9�/��|�q>x|͓k�-	���s��V�	���J=��_��ZzMY��_o���H 4;.#_���r��τ���3X���3[~�v� IN6��`��V��㾢#�-�3�k
�-s#�2`�����eh��s�1R�/�|v�*��0{��A	 �,z�`4�If��Sh LU.X��E�N"� ��w�w�$��O{��� 1[Pxt�*��	`�������C%�ހ�R(� ��7�ѣ� h�Do^X-��5��2QS}�Z�����W�QP�j���~�9�W&��
�ұ-0j����ǂX!{H��$�Sڟ��<Z�&l��J��t�x��in�w�KLW�3���_���g�{h�#�O cgF%U�������={��yTr)H6�j�(�pjQ��Re-�M�7)L�S풲Y��s�f|IRo_M�1�4	��6�ǌhۓ�����4b��Q&�H��wZ������f�I��KM�$�	
R�&W�N^�û���D/��Q��j(��Q�qtV�)�O��L$�Q-|
(/_'q�h��S]�Z܀	��,݊����#GW�w�b�G(	��@��3�����#�����U����Ù/HE1r��Qh�������٨˖��� x���l�B��r�Ek���3��+.kmA�®wVP����� f(�S�[s ��eR���@�~�š��KbG���Ph z�	�/b���KrT�'w0��)ϠR���fK�� !�顉�8��v�p9�%��`U�Z��rl��8T�Nڲb�ZB?:�L��5��J�K���ڗ���(qm��3*����X n	�1�h��cY�<Ts��L�Z���*Mp��~�P�K®hu�̕vrT�w:!�9j�� ����$��9�[(��V�N]�nK�M3����G+A�.y@���8&5V�a����X%`-��d!��<1&*�p�,���/��� �5��Q��o����Rs �^9�� �PUh�"�c��������]ԽBle�ǳS�D����R</��C!����/�O��8>�������wD0Y���\�R�QA�l4q��JWMW z��P�)ر��~j �}�Yh[��J��4`=�ײ�҇;|^J�Z�zR�)�N�bz�;cm Ⱥ)�HX�J��s�uj��0-�'�pD'�x­a>2)���r91Io
��8���_��댕y��S�$д%T��U�������L!j�fBhc8O��4��k��!�lh�A��'+�d^� �#\��-XB�'H��V��n?kUȯg�=��yYIOA�f`k���%X��B��{��5x�c0�×��f��'��c0ߓ�X���Iq[ȡ�J�e(R^���9�Uh���ؿ�׫t.�+4�^�s>��s������y->F�A�$�h8zQ_�,��129i��.�b^徴 U��fi0��� =�e1�)�>[�U#���)�91�	D���Ő��������-ZN�s,,f9˜���ş�7E��aQZ[�r�P��ho��/}A8�(���*Z!O`z5��<������k8�[j�w�b�w��#S���,Yz5 \�Q�4�U��{�RW�KI�D�	1�3���*�������=pB�x��^K��|G��2��,O��P��3KG�"jP[/1{�)�C\'O��l��4������_��3]��*J�y�A(���`�<-�tl�K ��H�
���?ؾ�_��v�s�4)A��q��u����Qަ��sw�7��'��h@�E_��7Zh�/R��
�>^\���S�� �o�/�o(H!|?�9��%�h�\k���.�Ny��1���xdA�r]�	�� z��w#�b���������\��
=Q����_)�z�q�8_GL�0�T����3	_���/h��9B�P�8����)�@�WD�^���4�8 ���/1��*��Rby�$+������R�k#�J�~�SE.���Q���q��K��Ҡtt��s@nOK6��f%t���%��S�?{�m1�`��ڣ�aQ���]븜c�Z�ۀ�	 ��қ�hz��:RtJC�@ܘ_,U�D5���]w�� ���ƀ�s��߽����%����h�~=,^s��_��<�������w\nB}uT9t���龲��%),[ė^vJ��ȶl(w0����A�1��w��`���,@�@ @	Z�ϔ74���(��&?�ܝU�+� ���3��0o�2#1����c"�)���o��}�	��8 1f%�>p�~6X�J�ΰ�n�x:�^�����<���%��E�y� �:suh&�`���*3�v���I�������v�l����	�`��z7.M̰,��!`��c�)�'�q�Z�����-N��ͼ.EX�_�IU�����ɷ1�Ѿ!�C	X�c2��?�NY`�����0e���B�҃�Lh�l��*�����P~��CUt	�d�EB-T�k����$O�wv���:�{�\YfS���p��|���sȱO ��L�}��zsV1�C����\H�{�܂�_
^T��@S��`���?/EXe{O�^OA��6�(v.�2ZSh�ÀX�[u�B'b-z��/�\�z��kn�vAU��M���1*�@YP/�Q���R��{��(�!�0[	n��Q�<,R����E�:���c N���Y�c��]�YZP��l
�\ut[ �}aN���ؕX!�M���� ^[����+�L�P���Ph�]ŝ_��!wu���/eܪ��N{�Y���:@,r7{�:�?�N�h��@��	�x�*@%�28Jq�z������� ^_��j,�E�\wA�V�2����Z[պ�h{���Hg��1�)��-����p���P�_�-����a�~�@HӬ �Q.ng�])�-�Y�����!�±��f�ǀɌ���*�-ŝ�?�_0P*$�AV�ZUJ;V��b^��`X@��"�&�0Wp�+�	�Y`M鶻X�և�#	��s��]�^���w�e -���C���Liz��+V%�P���	�W �#l�)�_�� |3�H������](EP�K_�I�o��N�Ay�|�3���j�P!Շ�g��1���{m�~�&/@����=�Aځ�k�LR��]�6:�S�In���踏U�+�K�9� �_"(���S��
@�1����\���m���F���?6�-�o����f^u4Z��1�3L�������sO���j%<�U4�j�(4g[����΄z`�l�}9/ 6��R��~'�Ŵ$�*��Ar��	�Ϧ��,8�EO���|}O(\	�O�h�#��1Сwt�<��I/W������WE��7�~Ap�y!���[Wh�V�sq�~����R���^k_]g�'��.�:�J�q����_�W]W`+@�b�Z��E��(L���<�D�7���HW��*��݋"_h�NX~�ß;7#�i݉߀�
4<)�HY�u�_�6���k�x[G�r��h�Pu���&�.l��a���rq:��	�{p�)�]R�֛��s�AhA@R8Qx�'/<��T~��#<J�V5�x^U ��0B=�|�'l�R	�;����M��
93��}	^vXHs���m�(��	EW��@âXgAP!I��>�,n�*%���X��s�d	�+�`�bY
�3��vc`R�iS8���^��i_���Q�5���^G���&�(�u��0���Z��`�Wس��:@T�/=�<��� Y��
+���%�5S��r���'%`�J>,$�`�颼��[a�=�+�`
nM/XM�^���W ��B.	fI��W�!�Ղ�g!u��)�]�	\�i	�/�o3���๼G2��i]#����m�6=q��zC&G�	�
Bq@XN��\�[�6M�~�cAF��J)�����rvqzSڍ�/�j���-�^_���.!= u�[h��/EX�`�ml�Y�k*��JhG}�e�1��2$&�&m�����){�ޞ�W*Zh��q�н��� �?r�')�W��U�P�Yr/����3�%��WX+�����oW����̉�jz3��Ւ�Շ��hL��0�1�$i���/�:�d����;CZ�f� ^g�9�h�xS��^�T���1Hj��0��N2�Е����ha#����/��_�Y���?ք�_�2��Q�R��#�Z���n�� ��ـ�~g����ߟ�4 �z�$��� ��r.��:Ec|�8C�W���Mi�@����4��7�^$�q�+|̯��k���`�O)WsTe_���ͫ)��b�vHs�LS�����)O����~�a7�;�u������XR��DK���A��x�x�����`�P�5�:����'������*�p%�y7Od�[u���=���s����1H���]f*��oYC-�+�o�'h6N��o��{8�`@�ky�!���9�+)�B�(�VY{c��y<]b&�G�wꚢ`�&�hð�6+��+�� ��W�<�v�_ �%V�P �+D(8�ջ%��t��: �}�@���yKp�Q+�R�S��0��O���p�j��WT�%��ugU�,/']6���A�Y�.����7�4�k�~0��69ohF\���1�G�e�)ђ>�A��k��Ю`��G�Z��j�D|�1?�(րƿ�^��#�������漙�+0�,�A��A���[c T��+8@C@������^���h�{�"@��!D/q)�(e�2]��v�α��	0 �����r0,�[�7m��̶)|�����S^���;���8����+O���x��zY�p=]�9#c�q����K�앨�Z���h8�l��� �H;����Z��T�>$�1{��]$p`�o���z�H�kK�;�kM��D�Х!�)��=@����(�8���I� B�^ng��>P]?ʬ&-��ccج�qI���`v�\��UY��Ak�/����U�^S�T]	3�r*��͠�0�,W0�X�gD}���/��(�YuF������0 ֒W�ɵpYv[4�'��T��-<+b D�b�_A������l!��N0���h!F�f^�Q�T�H�ࢲ�� ����(�J�㓾G�|�NI�I(��{ܘ@e$V�>kD��π������@����4��fP�0��!�Ѻ�G�.�O��!*-�)��p��p%u��`��i�3��_<��������Jq�Q�T���� O �5��v2g�
���fg��0��[U?`�sV[P�K$Y���Kpk�;*�<Rs�#�,��ɿ0�e. Q�إ�p�J��L6J n�?M�	�Bb�����;�V\��`o�aՖ����΃K�!�A6 �X(G��	
]���Z�fhPF+^� �U�z(�x���O�`�I��S�)����Q�YpU�ycO)��!�1.�}r '� �^qX��8�~j�eC�Ͽ �nLEwhGl�M�׋+�]����:g,\0O^�!��S�<=-��?�@�%c{��\�� W��-���6E_1[�	5��*�Gqa�@6O`÷�� �7��7��}�Dy�߸[�kJu�����x���K/�w+h=_�����a�p:h�F�:��E��u�-�<Z:t���lG ���V�ѹ��,��6�(��!V���'S��"��h��X�3�ܸ�u��U�����_<Hy(o�KX$���`!��~�u0=��S�fO�2����۷��$+[�����ՠ��p-�;�h?E�j���[u%  �����1*8�����zFK)����?R�D	�`
H0�*� �~)���<R�_��o�πk�ԓĶ( ��bq�0�˘�d0O�E���pj�n�s#�_"$��Mh�'��M��N䯊wN������\��� e	�Q���n�ƣk�C��0���^1��Ә\���H�#���O,<���=0G���!��H��ӭ��2�dl �����	l�JI���·.��v��c�w���A��+<�[��Y�� h~`�
'�g��m������z����5�t)�Uj�2W\�5�	NE |nq�Ms^$)B��Uc r��0!�6�W�0��xRtKD�O�鋹��hvo;¨d~���.�H2��?s7��4aLkr�ΟԝK�s��.�(�pD�q��3�T_�m���^%��2�iT�� �K�'\Z�{>.4�|xh�;F���	��	��L��(ko���CԞ}n'�GU�a���n���r��@��K��M7��H��	Mp.^!AW��"X�@7�8M���1ŇG�e<@��dVL���ÁMi��@���%-{erU��n��@����&|(*�۷T)�	��E؂>P�m1���U����]Eɫ��]��&(®~�0A�/����t�V�й�S����;4�*��2�#���Y��z0ENf�g��^����}8����-�K	 d�enfI��H	�2b�]���,��F��I��ר�������I$΁#�q�u����b�����_�kh�c�Eۨ'���0J\KF�4@��*U�!"�S�����P�û�'6���/L�Qs�:����[�?�i���Y�6{��������׍�F�ͫ*����<#z�	q�P�<�1\]J��N�8��g�hU.-�V�Xn1���.t`�TV?�w�%��jB/1�+�1Wf^ w����=�'�b���a����ԅ�H��'��ӳ��jE�0<�_���H�?&g��]��[!r��Sb����vz��Zu�����B6��΋?ް�� *L�J����3$�>Xv���G<�H�!� �·�B��2 @��-��Xc;�$�����������s��y��g�����	�i� �!H�^D#y%1Br0����w����h'�eq�#}�4�,�TY�H�[�5cR+����6	$:lߐ)in �޸��a��*e�1�)�|{5����|K����
_@����61WߛҫO��Y�٘�y�C���6UT�EA~]I���鿪4�߳RPf�_~ P-�X'�(DV���oP�U���]��I�@�<@�f���, Sh2[�p	�/8t]b�����1������B�^�>V��	`�D�@�hVZ�?ƃ����K^�<��(�A�)���z�[�� r�XI��/��y%	�m�WE���^Ro0�c�t�o`Zn��	%��SJ1<�ʀ�0�fZ ÷�_���u`%
��^�f�8 ��e�3[�~�_�쬠kӭ�v�PK;�L����2�B/8@? �k�T�F%]t[pM�J-@�9QD.Z��� RE�r�Z�7��1��X4�w7� ���d�|.�2�w\��'�a�K��9_�&����'sYK�5A�C_6@�J�:�09����ݕ�%�~�wE���+�i��>hn�2�T}�e�sd�Za�WRKK�)_�Z�H��N��V>��`KZS��#�0L�]�9�FC�q؈���{L`��C/&��Q-W��A��3�j4>���������Y
*)���~V�=0�PH�Y)��6���|��J�Ƀ��2*�ϣ{N��a03b^5�E�`�Z�T<%�j&�R���}gN0T��.�)��Wh 7~�H_G���#w��`�P����{f	W0F8Njˊl�Xj���^�u���+�)P] �~85����l�i�Hn�wu���@`t	���o�� �(V5�+	��y0:��*�kv�B�6!A&��b���]J�*�
3�%��(�$[RY/h��7$�
������D���S06��%ģ{��o�J`tC^׹�;��s��r��,���b�A���������w�D�hX	�����C=p���v���6$�l��<c3�1�m-wM|���'Kނʶ�uQ�^�q �R��+�J�WNؔYs������)1]�+����U�������՜
��Y�̽n�B^+�^�Re9��C�[Q����`,m1��0���
�<O3K�����������I��D��'���fŝ��dJ^�mA�z�8~� ��+�LK�'����B�,YX���m�r�ɰ��,�`��Y���~TG�Ni�,��"_/)UX�'��Vxg�M~��SĹW@�s�˺%��t鱽�p8y�j�����$�a/�����ӮB��W��^X5oZ�k	�T�'P����.:����(ˮù���Qh"��?܎*�ѽ@��I�&�P���'�0VL��$��Hm�d���k����uf�?�.^~�����ww>O��eԘ1�")� 9,�S��V�����fAU���\��R��E��13`��pZ�*}����h�z�x���ͦ*���>�Q��VzB`BP�	 �Z�����Ml����FK�P�u�Z��4���<����pu��'FmwEt'd`��ђ��������(��`��`q!�T�I��W��ޜ�<`�v0%]�h� �[���̾��Qՠk��S��ս��\ǟ�od$nOCBM��Y
Pe[���H���l�:��e!�1��)ŧt֪�Pͭ�.���h�N�D�-�R��#�|�p0N��H�;��=��#i������@���9d�jC�GHp^ShQ�A�~�Y|��B��G�<�|f��J4d�)��ێP"t�x�Ȝ=O�4�pP֗Q�����,��Y�?-����}�Z�Ѩ:y �&7 \��r��X�	�(��� j)ȁ��FM1�@�Rq%:~�	ͺ|ـ���xHJG�N`� �Y�*1���F�_�
}��~��W�%\pQ�a� ���M$��;Rh��@(nŘ�=_�_�����3')����{�/��#Z Dp�;2N��A��/���f�h�5Ѱ$)�K�u]��-���4�!�ïP٩ڿ�- �Y�`�h,(�F�-g��� Z�~3_��j@9��C�$a�L�X��6��	qztY�V6��XB�Ȁ���G���1�:������H)4��9Va��8�]Q��/`rZ�F��9^����=,]l�$� b�
})q�E���,h��3�-/�����HL�O�� R�|�'��j Y��a&K�3���Cx �����)���@X��iP�!�Z�s2Z�
�����^��7��2�G�]����	����	�����Z�b�s�:_�1%���`����U ��RuJb$h�\10S)�U
	��.��5m�(����L�n�����0���h��}=xC��RG�2��8�M��je&��m�*ߢQ�W@�Y�-T-���tOS�d \�g3�U���K���i����.���h�<�@n��|[��Z��Z�*�K����l�#Ý�>���(�+0��� Ś���1�����	�@���2�\���>V
���zh��|�E�Q�:%_jzp��-���[fh�aI d�(��s8����� ����E�b� ��D}r�P��똭$�� �LBE)�x�(|i���^�|�y`�P�k
�_v'}�K�9&0���1�꙰+�4+��^�C&��6���&�[ndGɆPf���XP�{�Լ���V�%U?o�ȧ�88#~��K�3�͠������Y=[�j�`8�G0н��rZ�_��e����o�vr\}x���C��[0�^$�w�^��AOna$x�N��ҿ�]!!�d���3QC�`F)Z��u�w0���	jJ��VM������{7jr��`�Vh�q�^���O�<r�Z��.K��N�Sh�+`����!L8�/���UUj������1)PqZ��7^��d�0A�_R{�d��\ˁ ��u�9I��يz<x�ˣg���ƹ�b�_H�(�/#*�,�Q��r�([��]@)�����f�_���Vdp�'4wTt��Z@��I&�e��$�:-��>⛡���@����)�-��p�����5l�D�C��Y���6�h	;�J�	�d;�c�>�,�]�N2~u��Tk�5���+l��������>�T ��/%;dpa%l\K&�%A!z��q��K �[1�k�����H깎���G1\D	�p����ƿ��?�ދN�e�a<���K���c����m0+H��q�L�J�p�f��p����)�0�Qh	�<A�lK�� ��b_��5�ը �-,�t�/�e��5hk��������-��\�������0Y>�*e L���}{9.�Vl�'S���-�R �!�'�b���ʾ��mP�+1z�Y� �,� �fXR��:06�'|�� oi���D��G��zx?�HP�$,4P8 ���S���8��:�����;4܉��	S�H�WAU��*�%P�u��-B*��b>'\�<��3ޠ]��O�0��2�	d�q���YZh�>T}A��R����Z�3RwJS|�h� �������Ǯ�>����t ��`��f_��ʻ�g2���\vu�l�&{�'�<oʚ�HW�5Ԉκ�	uT�K+ή���(O �Ҩ�LAk���+�[ ��,_ۀHK��F�� .���N%�,`7`LF�[��P�J�DH� �6~A=�/%'Z�/�x�?2Z�|�+�K̯R'j=`_Js�D)�%F�.��ju_/0<������u�����8�[����41���P��LD����r���ѿ�t.P�jN��dPJ�D��[�Tx9�&�X])� �I;^�Y�l�_�y�N��/�L��q�������(.���~ ϣ*��aR�,�ppR��>Ez�F�mC'A�1�<�X��lU~4���Ǿy'-s\_BX����M&F�� ZR�����090���x�$�]·�߂�h��Y������^�$Js^��xei��*L[l]WV
�!%wEr��n�so}`$�G[�`i��<6K���/u�h-�ȉuN��p��#@���a�G1�/�jR{v�%�cPi/%w�wS���{�A�7W����ha.�������x�6f���:QJ�B�,O~	�9�.�3]���v�%w�S��YR���:�,*�}	On��U���ٯ�	��ĘpW�Â�«�U�2	}iv����J=���%��g�I]nL�yH�}	3s�>�Qڠ|�JY�z�d1EQk�����PocJ���W0OE`�8,Q��U����+�`�h�Ob2���4f�K��<u ���� �вK��8b�@Fcm�dr�h�H|a��h�Tv_���K�p���� �	�rRC��<�o�/z0��(Y1��ym�M<�P4�95zK��4�G�_Q��@X�T��Z�y��3*_�������$X6I�i>:�H�P�9]�ZQ���ǽOm�x`oB�J���V@0�#�-�t&�kp
��1ySX;�mS+�N�/��:�X Q����������/0�Y��PTfP��(��X0��q赘oI���R��de��h���ހ��%(wܳ]��wX���{0���f��u�d8���<���0E�8�eS�[V�Ѻ�_�0��#!h/�:y��
+�=1�K]�=4�;�:R�({��?�Q�`y�d� qX��%�/�	��W��1��y萻]�O �`1�^�~� �6�D����N���a�+����3
�� X�n@N�޵z������j��
�o!Ђ]�*�p�K������h�0r^�t�8���2�� ʾ�͐�}ٯ�Q�C+���+�>�h\f�	Ws2��������k\)�w6�v���#��Gq����\-���'~�Y� mE�B]W�U�C����ԉ���
(y9	�7g��ý�+/�iTz�����	��U���{�0�$`\g�ֿ{�x�K� �q5�� ��@�L=%k7x[�J�d��r�+�W��H�k�-F�^��*��!|�^��-/�4V&�YS�|���	�r�ܨ���#��Q^k,,�Qݻz�αcvD�ė���8�̂�@�/y�bK����Ҹ�BphFZ��KN�'�_�(GR�cc���@�X��[ �Re�^|� DB-ASM5�?�O�@_��L~�1�a	:�`�����)�O%�8B�H5�@�@P�-���	F���]H�$%�}V_i�R�}���i]�̡u@��j;#H�-h6��[�WZ�´d��.k0��j��
��L�%�e���ws��� �(��V�a*�mwj��ȸ�0��y
��V}�u��{��K�LXWyKA�y�`)�N�v]gٰ�h0C�0��_!��q����-#q�e�鑊U�s�k vVo�^]��S����0�{��#q�+�z�,7�l�=�A5Jqs��T�܍O�	��.�d���1Ŀ�.We���S�Hl�'4)�C��3�/XEPUK��A,�:+$�!�0h�j�%[�^�K��c�����Jw^�~y�����0�m��4(�f��U�]g�dY��jV�P��SU�5Yd�髻0y)�u �IO��sM˜XGO` �5�(�� v\!ú�A$�7�KH|	��p �n�a�'.�����T�신h\N������.���d��y 4��DT�z�\�/�.h%<~�	r
9��>���Q��ݦ	4%���L�cZ�H�x�����YTl^���Z��䅋���m�v.��[0�cN;��1xio�'�C�����p�>������
P�^��=n�gvp4O[�)� �!w]�r�Rf�-��(X{�n\�]��	hTeQK&�A��P�=���;����s �Z�5�I�\��.��R9J0@R`!�',}0o��'z ��B�ߢ	�RY�E�.�s�5f â�ҿ�I�)�l��A�:RP�I��X�×p�������/�_ ���fj���Y�'g&� �bgE� �f'3%�� NV��<%yt�N�&�B�f����ŭ!�}��kΔP��pO�:����8w�#T�:4z��|�|nP����)����F�x �5�.v��\�=�@�CR��|L�e!�h8��S1�ZU[�/Q��X�9ߜL�
	r6)ڡ@nͳ�8�)��:	Y�p`�uO�`�t �[��frPhK��|G�؉[(p斄����w{
^�k]� �P|�T@��B�X���=5�yP&W�@L��\�
W��t�M0�_�Ġ�J�����n`~��)�e��GPu�订�v뤫 �&M9��?�3�큐��k	�c��P(��sS��8��?1��6�3�d	�g�4?�B&�� �w�p)͵�[b/[� e�O3�2��j3d),g��K�d��{�X)�x�X7�P�Z�,@+�9���^)K���? ���QA��@��l>�.#�~1����|�Q��~B�^�i��iȢ��M��߀��N��x�J����Y��7S���o��W��j��h$�.�o	8~n\�t@Vr���)��o�c�s��`w$�' G��)�0�v���T�\@����ɼ��&QW�P�� U���]Ż�����q����+�<�Q��G|���'ZA`=��Ѣ̀�����l�=� ��P+��;@�!�[�؊����"0`h�
$}}�:��oj�{�1�G�H�w��$6]h��@��S�5��A>�`MhH�ٛ����MN����+o` S�l	�[�V�/��Ř����s����"N��*8�� ��mo��tO��*_-0�-ƞ8�Zi�`q�׳�Xh%k{�����\)�P0/�g���}$;�b�z"%A;u�� K���
��_o�OD��,L#�	��	
�Ɂo�G����}|�ϼ	��V�U�j�8#%�
�E�Q�&��=
s7��[�*,Yo�	��e��^���re�r��[��f���H��1�- ֡�M�J!�1(U��z�X��K�"5�]�ʹ	o)��z�	�u�Tѳ/�1��E ��rx�2���[����q֙�@~`N�j6X8 λ9[�d��>��U;�O�W�)H.�%�@n�qR�y�_Ë��@^�S�� 	X9�O�u�x���wz*�ԦK���B��󢂂1�7U��%�$I�� Qh��{JZ���ʇ�~%�8
P9��M����>�/Z�;��Y���i��f�B5%.���	G8D�D�����{��!�����4�}�{H]`>�d#З�=i(R��l�Є��y:���ꊟɻ0~e����Ę���ݤ(�B)��*�sP��%O��7�@pS���ޙvX?�a̲Q13�_V�)�,W�P���t����`���
���]��+")t'��pQ�e�������p�p�b�y�<�{�K0�	�@�ح^�~�^��%���/0k�*_�����L�o��nX�8N������XIB�P��I��;�7p����v�����O�JXQ�z�=�\{A�&�D�����̙{�AŨeI.)�O����ٽUJr�ŭc_)�p����:r�W�~��������PK�� QZYh+������	���������ϳ�;5Ko$��Ӹ�ˎ�qw��do|c�^�T�h��`bh�Js2M8,*�V�F�v�o`���:%MY����kT�P,H�
bs��������
#�%�Ta������X�}���Ь����N�(�� G�*(F��.��7�����l~#��=���H�B�v�G	=Y�Qa�����U�t!��K����Z��Bu�o`cקr�@Ľ�>+�P�	�e�a��[o�<�D�l���8Q�r�=N�U<	�����Sa�7C���ψ�{��>�����������<�M_����h�l�fDj��v�0�ۄ�H��]�c��T$z0[��_-?�S�0g����_8�rpd��%�[`�&�����q��}�Q������ut�����m	�i6���>y,��`�u]���a%
8�OUV���[�� ���!���	�+����[��Dq	W8#��OZ(���5%Y�Eb�S�����1K��(��޺�/o��ph��V|]����	����@�*��_���4G˪����Tm��T���U�2TJ/h]+Z��*�Z)�]�W"����h�.����$P-@ OVغ,+H���ld���h�OĖ�W�O)hP���:�(崽��@1�ZUh��LX@-�IF7�Q�8��2�|5���}���QȰ/�9�-4WǦ0(�/%*1W��P�pr���I��K�<~�~����QQZtZu]�"�u��ƯN��{'��Y�]
�\� �q6�OE��z٥S;Az����R��5��c鋄��`����;'�������F�as=(�H6l��� �X�ѻ���\U�&?c����4�B�I�j58Ǥ��/�=^	��_'B�ƿ�HT%+J����j��h^�UEI+�'.�6��Uj�=�`���gp)a��`��OO��Շ1�&�7��
A�K �^m�?���*j�ƽ�Ct&�	m%b�uj' W�w,�3N	_�U,WS2)c��%��t�M���郸/ �ɒt����	�!�{B\ܱa���>�΂,��1'��y�l�~A��
e�){��i�53�R)���J��	���'ԗH�^LD����1���˚R���*��>��l�[��U�%ۥ��n��T)|�LHDb;G��	�$P���h>G@��S�*�Q�t
'}�Nd�l�)�r��}S��#F{�_Iސ��:;�i�c4dJ������K�8$?%��kTT���<6��4�t�� uKi0���Q��(���ӏH�6�h` ��@�n!���U�УJM39�/�GT9�i�e`�Q������?�@Z�iHP�(B�
k�~�m�)Fޠ�>�K���9R�CGt�!�������T`q_[�)~H��/ga_/m��u��~�<�XL�U%�(��k�8)�����K �"p餱A����0+����!`��Z��`E�uk�LG� �bL��ٟ�a�w�@��fC��./��l�07���N�s�yՖޓl�Z����Dz�^4��t�D�i�$��1�c���ˣ�N�ws!��f-��hc�h&�)��Ѝ��, .kU63�C�����.��k�E��hD���f��f���)BQ�T�E�@���zL 1�[���U���b[���~�%H�`�����ܢ��yپ��v�h'�;� ��C��Z"%B����[�qK|�Z�v��=���S�WNc�^u�(�SY��ڿ�����g�J|�����K0�V�m��m�P��F�1��Z�/�׺�!����~�:$M�)��C�uA�IQ�Z��y��.��W{?q)�1Ӻ��Z��yHQ��,N@ ��\;��K [V�ݙ���hpO��.R��Rg�՜K�!0�F��s^��0C�5����v*4}��F{�� ��X���\��4?�(���������T��\��7��f	�u�,V�nX[�;_���@�Md�:���.^؏$�(��**����e)�g?'���]\l��}s��uϋ��=թU��=��W����c�K*��T���1h/,nhK�1�޾�*��s%w� U�c��1���� �ӂ�����{.@�5��V��Z�wZ<�DҸ�	:�u�/�Fǟ��S�� 3In �h�9U��N��"M)���tv,	�Eu4�LF��!`Y@-��.�o8.K%W s�d��\(aK��r��q�~�F�	O#��8�����W+�E�Y��e��6e�Q@�U�E�t���w|<�W�}?�Ϋ=�j��p���O��J(��K��"�;7|";�n����2%oG�rd�BW>H �
� �&��� hpb3-[����<����LC�>0!P�eM���@��=o �&�78,��R�"bJ K/�{2k��dM�D0Ыatͧ����o������Brs
�@1�)mh	�&�N�F1�ǀ�A7g�+p�\��Qk�)ȉ�,I�&O�B-�{Ra��/H@] ��$'Gr���c�~>��p =�x@5�S��b���ys>�"�g��x'�+T_b".t,�Q�S]���=W	���q��\!f�18h'OL�pO�Ƙ����dǸ`	�c�O�b�'-�	m�Գy�$!VJ�CiIҰ��N��u�պ(Z��C����}5����L�/$�A.��gC�����`n����Q�������t�2SI�w��n�q� ]�
�Dy�ڍ6�2�T�s�bd�v��]�	��� �A��!�t+�R��4���(�}���L����X/.4p�� -&�>L7$�K-;�����jtg3��Y�qO��W��RHY���p�) �1ѽ"
6E�&��R��!�����	�{a��~��iX�X��1:������mG���xX#�P���6\� ��@D5Ru���oe(k��	B"������G< ��}\&o	���������J��#P���	���D*N)��L��%����i`h��dY�N���4�jS���k�O��s�a������0s��.Y��v�c)=����[�j��_�0��
}%!�鸼���J��-=���Jz���yi�6���W�[��"���'b>T/��>ū����.���h�s+Jd�-�����Л>�D�?+V�bF��T��@�'��D�Z��^��ic,��rW�z\!W�� �NG���R��X P�Y����,\�D/����-�=��񠫴.��Ή�I�i�	fa|h`/�����c�p�-D�����.� Ύ0��	LC�s��I���!~���䱂j��E ����M�k��V@��2�x)YX��Sf}7�c�S����[:����iUe�ɰY�x� �S�;�-ˑv/������HfFM,C���RVZ^��zw� �Ph�nX�6 9/�1�/v��[����	I��Wp�ފ�۞�c��uxV ĕ����-\K�O����1�r�'WW�0����Yg����!K����p�=��B3UG�h�wu�Q��u��:_^�4ZL �����)���!�ʦ�f ��1�-y>�nC]�����`/*^=�C��� _K�7�A�`&xPp'���~g������O��cR7_ע�$>W!��|���LiJ��H�0���k
�KLd6 ���K�;��n�VB�	�^�#m�+_~�tn�u�:�o��t�T[�+�(�����EX���R�'�7�����{�z/Zﱣy�ŋ�-B8�@�?A��TK�
���mՈ�� ��p|�9)�?Ú?^��ɵ�0�1w�v�����Z0.�f<�'�ǉ�o��P��Z�VX���N���LTw��jş�����3��
l%�Z�\=7]A��\�1l�n�w��@��W�:,� U�]L�{����C%��<�荵p{��!xtN���U*����`��i."o�b�tp��[DP���ϧPi%���B�k����F�¬��|��
������C�yBeՈ�$] �_3�F�.��L�%QuK���p}�֒��t�N���0���1�Y )�-�u�g ��m��S�[]��19������[�Ͱ�����u�vs��L�OS����h)���Tp�t�V�
]m���v���h�>���\�'߶Y���`�m5�<!��1�/�{Q?�[�i�a�Y��	"d��������Vo&q����T6���Ese�[}B�j��*V�	�n����41��X���r��g-��I��uK��<g�'B�hw#��)�W���Q_?V�1��Z���Za�aR,��MC�� "�~S�j�r�Pl�� 
2X�A���P��!�*�RT�y�U�e�����n�;Q�p(�FD;����{�@�V��A�^���C+Q��x-U	 ��R�Y�)��b(P/Q���W����B�����4<���ϔ�!Qu�]ҹ1��M���[:X�'����u�C�-x	�R���e�|Xl� �Ã8�[#��9�T�,�%^!1e�q
LB�'Tܠ����Z߽��y/�'.���LX���0 �x!	�-8�֏iȮ-�R�SPU-_T;�gP�@�K51�B��)���אYs�(���B^ �� �]g�m֚3DLN�j�-�1(�HEYR�Sҽ������#��Ծp5h�Z�ǝ$�,�b��*PO�s�Ah�xÄ��8�}�J�XA�?�D��i��U�D��u��Bd�Ӻ��ߪ#�^	XL�QG9��ʢO{�M�����1�hўxi�h_OG�hUg4�3%_�����5�1��Ք��+�L��v�6'B���!Ou��+��ӻ�q��=;B4)٨���ެ�H�(�̔�P��1�A�����8��ۓӼNX0	v!�6�zmy��jR>*���� �z�6�w^�O�o�S4h5����z5p�bRZ���#hJCC�^�>�'����IZ-�S����R#j���(��ā��?`�A�(vP�N���oh$n#lJ���Rh�Z2�E� �
s�`2$��P5�W���!�֤� <��P�\�Bu��z����g��[h�^�ZR}���a�}V`m"H�r�ނ3�^_P����'vT/l:$�̄'�J/8�h�3������m;�����42>�������X�lhq6�P��`�c��]��ŏ���i���K���u��o���h���o�NG ��K�0!�[s��N���	�%p!����1���zq�<[܂-J�U-tqodp{��5q~k(-'/�i1�|l[��/s��I
�}�-��^Z�p�U��s�c��R�3�7`��7Up�Nf<S���ì��1�_u+V�E�`+A5��"k�P'��_iW@��	�^H�E��*A/�~�zG�����)�E� P�Q���� YX �fZ�h'K0�H��N�dM��t�)�ۉ"�,K��PͿ�oU�Q�d�~���K2�u�짃�`0_��8΃�UM? �� T�����J��$�(�=|�����ݹT=h� �P�j��n����M`l��M�m�e����V�l����Y����FK��(���+�r�^�Ov �� ���:j����]G�&�R:
���	� �0WX)�3&� �(e1֘���M��눎v����P�Y��h��8<@7- 1
0%�&	��✫-S�|������w�)�R�:��Q i!��C$����/�z=��TY -�XL����U���+�P��?���[�;^�O)��ߥ`�1?�
�o�\U�L=��ɵ��H�a+,9`���K=��yHGvS �b�)O��k���0׾�y[���|��I�F�p�7-D���;�8 #���S,���^��a��!���u�X��*w�`h'�&����*�h�|^H�j%�^� �tlGK�Q�x���Fa���
J��ZK�+���<@�	wG{>�Y���k$"$T�o���"{&߮%��@k��F;A ���)x��ZU�g�Ƨ-�������d��؇�'����W�H|.�L)K��S�%4*�V�q���æu	%����S���"y[\���rѠ�2����!��Ȱ�:1�r�%���`*�8�[x�]؀�2�<��R�'.U���wt<yvK1 �3e�~��$y�<��N�J@ܡ��/$]�[��Kh,�t\i|}��`��V�-B�v��!�5����GN�נ��G�\���*�J �	hf�[��}��T&&�>'���C�@L�	9-
F�f��D"$:�ˀ�0x�L�.��\����[�C��nPxJ~2~�r��7a".� #6�)�����j��\���=Y�w��b�@R �Fi#�9��œ�)� �E v �Mpd!��Nu���k'`wT�56������ b����S0"x���(J���
���JX	m���a�s�}*`&ez��S0���1��}�j� Yh�N�/�Zk���e_��_k��1�!�hJ?X������P�r�q�jg�q��2�a�k����s��Rb� 2�^M���W�9�n�����h�[p oT_�?q|H{ œ������KB��hB��ee���p�`�雯�˽������ P��y��%�r���1�a�t�#@��W|���(�/Xd)��/�v�<j��=1�`�[�y��s,~��O�J��'�^�AZRY.���]��Һ��� �)RN[�@�5�?����O}��ء�Qo�����{�١��?� a��\�'!ڤ@� ��_O�� ?1J��c�*H�$�@C-�R:b�mB #�~���-6��,_L� P��h�r���1�b�Հ�Y	"3-.0�B�}���O����V0~ѫ��W�T�F�#R�o
'��b���!�0�z�̨Q
���/ו�^�{J�*��m#�L2[�#�Vx1��CYM��԰q��,\L{�zDF�������Ǖ�w{������l���J ��)�4�ő�G%�����;J�]E�����)�J!��V�u�w$h;�A��x�>,�{<�J^��>S�C2�b"�%M6%9[�QS~�t��j�$z�G60��s�mA[����"�S�b�������}-L���i���dR�0��su
'0)���
����ػ��)�UE�t1������-�!Z�����=�ݺ�U�m�vu����TXo�B9� PU���AOS1 )ʻh2������s<�ȴQ�MӮ]��������%ÆMHb��^oǉ�k�զ�
S�P�2(������xE�!R����h�����>B��!����R�x�']vܐr�E� _?u�
�N���Z�V��9����@W#5�_$Xp H��	�(��d=Z^��!�a'#�b�HM�U/WM��Q�?8|+��ϊ���%vRrW��B!�]e�'̊�\�A��C4�ͻ�L`&6G��CW�L${j�E�Ve�aB=T�9z��ծ[�z'w��8D�D0�����5�%��e����ozA�/�! B�i��a'�~��1�؀
�R���Z!�X �n��<P�Y��A���4���Bu��W�PxH�|J��[��P��4Z��$�\��1W�J)}���~|�^/G��d��hy������v����3]�I �nę��)�G����C��[�In��@]�^��	˽Z@� F�;\�I��~H�h�[�v�]^�;�{^P�ѡ��FZT\�¢v� S;AKX5��gJh�s��8L
��R/�+�K�(!S�u#��"����w��q-:�Xg�(����J1��A���].�zt	;���CB,�}Tt����U򼾳��8E������r����1J��$\�1?��+�\`
�ۂ-�C��.�(�����Ŋh�w�J��{B->�w�0�j1�S��� <���y �}c�Q1���hV�֝�Y�!�,��P�^�"`ۚ��F�`�E.Oz��1幀�C�gT�Va���ژ�-�s���	�Cx�vAR>ME �A�Z]`���HDP��s��'cV�AP!�^n��s6�]\�RtC��p���hAU��x@��U�Q����ayFk��_�qN�,�3+[����h��n;��t��Ch%�����~&mYx@���v�ȹ�{0�k�J<����B�EZEB� �# ��ΒK��I5L{��N��!�0�H%$8�-th<-����X'P9�ǘ�)K#.
��B��]��B@$/@�/��P����.�NE�]c��`i3!�+_�R�}nG��G��N{O�+�`2dP�" B�ZPw?wh��^��Y %)�~?k����:=�čW���	?m���A�%�;���x��%���!Z�P�C!��h E���v�}�� ��,ec-��k�x`l�o)	�h�
��N�}*ѭ%u���흕�ɬ�u��3RhX��(�! �+5�*K���|�e��w�D-�!V�U��^uKwE�i]>{�b�עU���YR`�X���;�*��O0�
5(� ˴�[�R��wޓUG�8q�������	"��g�-�>�N1�0K'�R�2Fۀʰ]�c/����aV{Q��;��5=�?��Ub�N�Z1���S�2���5�Z~d@���paxF� �1K��[���-$I.0��'�	��[�w�XԶ�a=���z�sK>1Η�fH���L�k�W��h�-�l��A�Ւ����0��\d3p.2z���Q�_ą!�[�'X!Z�$_
|A�'w	�E����i���A�6"�ǣ^���mb��
�	�n�GK\��Y!�λ]��������fZ9�(�,N^:��m��_���q���ܛ�wі���@�Xh/Huy��	\?`�<�&	����	a4��wd)�^K?�������Ph>/-�op�8E��(��:U�|_��@N�n�2�<ю���O�H	���1Y^X���id>�ts��ӟ^C
G-:�W8��x���K3��_1p"9H�:-�H�@.�)�% ���b�CH��[�d���2�D �0�,R@!Q� ���ŀ�poK���L����G�k��|��=�|]��hwf�]r[:V����*�~���>�k)
�g���b��HfO/�t� S��Q���l[X(+(���n	h�'�e	ؽp`���"�N�P�}xOH�H��Ij*��	�qz� <SB)ڹW9�ڴ�_C+����052/�z��� �c�`��~����AȬ��������X��2(�s�7n���E����O�'ߗ 9�7Qn�1���$v�"V�	��F���Z�!�o-Ȱ���� dV�G� �P�ET�������+�ss�PQO!�~	�=�ـ��P6c��(�Z����UQIdD��d�@��!]	�_�PZu��:��m�;�/9� g�~uT�X�Ŷ�ф���ˀ�P0!�р�J�,�rZ� ��	]�}0!��7�u1�Q]H	��?�p������i<]��-���<[�
���gkC�ߏ9g�4i�D<����;�f	��<���0�ל%�" �d�C-w ZE��@OB9@�
�3�$^}�Qg��Bk�M	�\�/�'�IbP2 �����v ���	�@��6	 h�h}��p�.&K�� ��0{?(ݫ���H	; W��� �, �S-��`	=0wDA���_�S��d�	�AZ KS��#�M���]�f�� �Kܘ�-Q[\%��Hy����4��X9�㤀)��8w�J�CAuV�����%'7o�'reH�� �<F
�꠳�30�̊�)���R8!:�V�gH{�j-6��� mF5*bc��G$g���	�\l)�׎1�e�, lQ�v��^��	&��LS�e�C�!Kj�4����l4.�cV9߃�P���I"�Ox�1=_�aB�d��]Y/:���{k��|$��U���0wWh�#�\_�b&��IA��g;@��oSC)H�F4$��(\�b���%}���M.�ߞP0��Ph�-dt����*#}�f���9�$o좹��۰	�e~��W�(²�YQ���k���pF���t�N��Q��Ĥ!GRU06�J����J V��K�4a=:�.E� �5| ��nX��זP!~�Ll�@��Shx)�DZ@��$�Q�T�}x�	j>cU��_d���T��x��I1�\��\��V��h!�����,@%�B;vO�g�@�y&-N���C
9�8B��Z�p� ��TN;�#���	�n5���.:X�.�o/�hT�U?�e&ڒ J)�A��A��o�
�Q�T���'�"�I�_������ƖR�Xh�;����7�,PKo������쨠�'�	鰥Wy�A7�>+|�XC�3
)Ǒ�~���V��߈ ��C����hλ� �AjXR �\h;?��c/�}���E���o��r1��U��b�`�@��Vzs��;��p�ڋ�\�.Y�q����Y ��au�c�I��EV��A~��Xh&{�0������G�F�2B[@�lPH�Ž�u�Pϖ �?��&�<�R�'�N��v���@��/Ur�ї_1�h��P�נ��vڽ �#=6J(����M�q��!��E%J�\���0 E	'�Zo���t��J�
x� �ux;[�����9�%?�<PR�9I�L/�h�Y��i!�_�V���hA${F���H�r���mhn4���[�%���q�)-S0��5M�PH2�np!z9y���E��_ɂkl:�O�%����1�nZgW��ת�F�p~'F����`�o=�� #�Y��p�uS�z�@\�4�($��D5�GQ��������p�X=��-h4����aa*��E@��h/�O�� -�#���.�_k/|q? �K�n�M�~��H3p�sy�X	 �
�)<'���8�^A2s˴6~΂LTYV��	�z��WN!�����U����7l�3"�sH��]2?���!X�+��Z! �����wЕ�PܺC�.��1V.j)���U}������^wxpX�E�.2pK50G	� �e�1��w���iS�� �3f>�o��J�=AOhx�v��>S�³���}�������������������.���M����<+��eHW�D����>�
�X� >m��(vj�$-��%W ��(0F�� �tR�f��\�PH��%�ie:nɻ56�0�E9�����1C.A� ���·���V�5����� ��P�(⺘��=zD%�b][[jL	� ��O����ܾҵ�_B\h!��X�	�ZF����8��"��钕�X?��Zhvw��HV�{^/`�i\��J�)yE�^���H_:�khhWE�=�Q8�YUa�[I�0�����k�����UL-aGf�k	�ޯ	��?�#�O�x_.�^ɒ�n�-'�5*Dk���0�$]��µ�ˏ��H;&@N�<�]Au �5�@z�����b[[�+KM�~?�����g�Јh�:�i�3F'D)�\��[��*��CD��d���� �/[[0��+��-��J'�P�!��K#�Ю�n�J������x�y0<*�OKU����b�����Xl�K��Z%f�u��v�9F����a ";GXC�^�d`J��J��f �Y�<�j�mVF>��N똒�1+V�52 �1<-��;���+�ɲ�p-y�`��Ү�e��Z�_�Rq�Y"z�����p��z� �I_QuQ\.D{ȍ h�:�y	�I3�՝ᄄs�"/��/@��ưC�U�vk뀄��M+�:�Hr���DS��������aO1R�ϱ/��Ñy(b�pO��#��4D���5|0VI���#OY�F��D�Z��1:v (�p�(Q�	[�;��('�B�����	B^��`�融�Kۈ��!t�-���SZP�dh�o���" ��GO���E�e@NU�G��p/�I�d1���Є������!@`��gOP~1��[YE&����uX-発	��@�g(�����V�D�����	Г�[�*���=��	��;u�!C鈓��[��r�ː�Ff�"�[]!K�7�+�3���sW0��)�-?a{���?	p������z ��q.�|� ��8��Kռ{Ӽ)��T���W	]>�{4
���{(Q�>A�8��#�r�_��y8K��=��U�����YHqQ��7�l�0z/C�;�fQ4���S�� }Td$1�[.)ʤ���fB. �&4i�2��Eog��W�9�#�����&�5�*���u�R�	`n�&p�7�T0Q��g'tI� U>�������k��UTA��7��
��V>aD!�?���j�����s9��/p/�����>��Z��hQb�-`j�^���V��e�w�����X5i�u_P51_0�JS@.M8%���)I1�W@fYS��U�kN�G�mc,3�v���
�d�ԁ��(�`��r�Pc�}m�VֺO�͆s<$X�����@]]NM��D{)�0`h$� �53���|���{fl�B��)����Rh^I�s]� �`�&�����W�`=��$A@�~a��h�Q������G8��])��hI���`��B�	t�&�Zh��[X�O�޸\�|A`T�S�ƹ+�zHIK���tPp��7�K��D �|�^0��_��o�����uތ��?D0�_��AW:�����5C���t�� �[5r"#O%��$Yi{o��(5�xkwE�[ͅ�����u�,O6 ��gm�MMPC+(H�� 	� %�45��n-�AW����^�{�S1J�#�ɬZ��Ѥ�� R�a�h�V$L�)���<�ͼ�/�^�-���v/�҅�QE���Ծf/R�r	���q�V��^�D����$��_�0���/��Z ВX��B�>Wr)E�+�#d̈́�B48E6A<Z�����R�0ג�KJ��X�@�%Y���R��?M0��zc��(��h�|.�Z�k(#�Z4����/L�6ھ_ ��`2�9����7`�Kg`Q[�J�J��V�t'�:!���L��X���64�V� �odh1p
^)j���CHAeJ�-���5K}q%y˔v��T;�׈�ɘ|A�(�ܹF�ӿ0�J4��@2����E1p��ֹE�P��{ �c�1�!��VN�I����1�Q-��Ԃa=$�13�@��'�N,�g�G�D�:B��t�K��G(����pN=��{bPi���eJ���� �+`�S�63'�v���\c5��E@1�����s'�Uh�$H�	o�j����F�4"�����D��a� �-�y 5�1��[�ʺ�8{���k� ޳��?;�����!	1�����#~k��cMq`$�%$�&��'mS=���$v({N"`��^,���r��C��;}��"(I6K�ǿ�g ��
�9���d�Nu��&R� kat�o����u	Wf����Km";	d,,�+(�h���!�`9��8$�L{��q��� �7CQ�n����H���[
�uR�4yP�/HհE-^~`�<�c7-[tSˡuL��U�x���(Q�{��H�1�0�甁���a�z>Y^�]��1��,t^�*�:�8�,[�P��M�eMbՠ�e�t���$�A(�h�|t��<���-�nu=�8 X�qh�+��oC��E}I% Z������)�%���bW(��"�e��Ȳ��i��J��Y�p��ӖL�;�u�_��zm#/6M1�Z�&5��;�-�c�
:����`�_���qn�����S�r@
h$A*�i�����1�GtQ�;]6�)�U�����x�v�8�ZfXG�׻Bv�*�N��'�r��R_�	m���2D_������J�����UVs��O��:oo)27s�����,����5���Lj!�H�&��Q�4(���꙾~�I�]�
X-EՍ��j���e�Չ ��s��g(�S�9�L2L����˒�A��m��U邜����%]���E]�W3����/����<,��1� 1���������[P�3�ː���h�(-X��Aq=V��i
H`�� Rc7-�1��	�d�uBJI?���\�S�*Jh�p!	�.RU�G��^���|!�Bj�e 1�X��4{	0����Fo!�v�G`�x�(Y���;��b�qp���Eҷy0rh�d�j�]�ŉ��^��I&y��R����-u����Y^���������(&��
yۭ>~P���q	;W� ���)��->�-�z�	h�S�������J/��FWX	a�`�(���u~|m�����z+�)L����A<�l� 1�>���V$O����|��.��?�Z�(��Mc���P0ZV�T��'�(Le\�x��g��`�b�Չ,N^�+��B��1I��P����+�v:	�0��|�O�����:���\J�	�#E a0[�&��Fr)�1݂�,_��2>��E�U�� @�9��'+ixw	�HR%���y�Y��X�1����"������?�e��J��,>��A$��Z0����z�AYY*AA�#A�ST0?�@���{ �j%�l���b\ ���3����p^~t��|�6�i���Ƥ�����T�m��J��� ??R{�(�F�8)��,e��8��$h�Fy�����Q�܀9�Ȃ�+��π�H��-O<O��
n���!迏jC5��'}� �\�q�B���Vp�y��QJ\Rk}j 9�C"�	��E������ $��hS}	UY��F/�]�P�#:�$����(Z,�"=�V��9%�.�U���R�fZ��dA>������0{����X�����h��'�^��h$���ʄ�;��A%1�?ؿU\�hl�%Vy����t�kF�js �C�s1��(R�}�D3QQ��`�P�)_�� 	�R��>d�g]4?�j��8%�,.�e�2HK����}�d%_���*�����o�O.�ꊾ%��e'ߖl]:�eH$x�$����x)Q��J3c%���������^��R�5�ؒ����RD������ $����2�)h�C4	���D�8������1�>u|�X\1C�4T��9�b��0��/��4�]}T�+@ ��U, �b�1�w�[Yh�J*��Pr����ڦ�$�U`!pn�R?�����T<���z1@p���OQc~|�o'��˓���	陘�j��Y:|�mV��C?�}���Æ�vQh�e�1�0n�Ʉ%��T�7oe��@� W���8�"p����RP��_I��Ͻ��E(�;��#Z	���պ-^�cB��1%0����i����rp��?ivZ3 �Y�>W��3(�}���	�*�=/����r^� ��T���@ǁ��;��0V�BMb��,�ߋ�z��Q�^��G��>�d�⅂鿞��١hJ��&�e��46�yی`|� �uB,��C<�l�)_9��R #g���� h�:CX% a�b5p�-�����`Rqdq(�{`OݴF�$@�_�aH�Y���q��<��/��e1P�4C�����0H�`������Չ��1�@�3Z X��*:B�&j�!I���ãBDh�� /�`��R�)����H� �,�j1Ӻ+/G���_�g�Z��3����U�>I��V�u�x�k�	¡���f�xl�i	>�Z�21���u�Ƥ��h9s�S� }��_uM2��1�H����th�8�׺�����H-�(YP�p���9�b��ox�V��F֍���t���W� ;�#����d}�}�/�*[�a4�zŉ!�@Ώ�j��phhU��$�����n�1X$����Q�c:������vS	�T�lW��k{H���[�D�P����l���B�����o�D����k�\^�[6���Z'E%�kF1K./�}h�G�Z���-��wdNr,�^�e�7�{�R:�}��Kc��*�R^EV��,�F)o@]��� 3�0�fA���i2�r����`��j�F�(>;~�!,���?�-���j�NI) XH%!.�#	��<^���1+�hJq0z��]{HV���>E���]=25�����S�k��U��_�һ���@H�/��PZ�y4i�	Q�^���	L�3MS� �{�s�����0!�P>p`_OTt^ )ѽ�3�2h*�.�*�-y�E+#
�bf�0 �7Q�  ��¦s��dWS@5PV��-#D_�1�!����-�P�����)�X��_��4�    )���t(i;�&��s&�~�   �4$^��W��0�()�_��3Q���ҁ�L�Z����i*P�����:t���}$�1݁�Jyj���$�    �   %�h�D5��\�������,#�8�Is��&rS��vs�:��B��asс�^��)Y�A�u�~I�����������Á�s&�~����!�!��    1��wD�$�0�(�3�����O{01L$Y�,$��   �H�����j@h   h�   j ��u���y���j@h   h�  j ��u���y���j@h   h   j ��u���y������yj@h   �vj ��u���y������y�����k�������yR��zB�й?   ���y���y�	   �>����I���������y�����k����3��>   ���y�����?�F������yF��~
��   S3ۊ^
�   [I��������j@h   h   j ��u��)!������y����ыFk����й=  ��)!���  󤋵)!��)!�  �FX���y�FD���y�F@�Ft�F<���   �F,�nT��^�%�F\�    �F`��	   ����Fd�   ����y��U����`�E�    �u�H   �E�X�H�PU���   +��   ��,�	   +����   ��4�   3ӉP���E��>�������E�a�E��� ���y��8�%�5�&�+���1�ȃ�I�������/�%��Y�%+σ���1   U��`�w8��   �w<u��t�G<��p;��   +�w<�w0a�� ���   ���b$"B�3�x��+ӔZ�    �   �%ĝ�}�xTg��g�wi/��    [�¹[  ���X��Z#X��SL#X�   t��\^B�@k��2��Y���>��q�kd��X\f��؁��Uyq�
�   ��P�����A�wӠ��oX�꡸�V������V`f���   S^aO��������\�� A��k���EV��G��we��)��K��!���E�E�E�E�G�Ԭ���E��%/�E�7��B�B�Fx`�k�_�dx�qD��L�F�~�Q0�%���}ّB�B�����E��RɊa���D�Ȋ$�)E�F�d�!�l������2��.��{�S�u���)$?�0�SӶi��7���F�����XѵL��'���A��X_Q�X��<��Q��S��9���b��8�5öm��G)��E4���S�e�7d����ꕵ� ���w�b�쏳�͆=�����a"LЗA��ĶK_�5�d��~H2���|�g�� ��j�{�$ W�guԭ��1��Ŷ�r�?黨;���!�E����;R�ّP�~��1���?~:� r����؄�P���\�9�Tl�jj�b��b�C�*Aǜ�E$'�@��m�R�E=���%��Y�<Goն;��SF��3���JNi=B�]E� �4N��. ��ME��&�E_�檷ض!Qg�߳��D��a��Q�������`�����E�W��V������OF�۶��Xq���C�F��������C�,%�l�l�6���i�kR�����K��9m�h�RS�������_�ӏD�g2��\�c�k�t����A�C��AE�w$�2:����=F���G��7:�&uBȶ��׶���E}�S���l�$��\�K�6E��ut��g��v��E� �*��%��jE7{�-�`5B�DY��=�!E$��f�D0�B�uv7GEA�|~�B�Q�Ӷ0܁Z��P��Mj��Ʃu�MտH�͚�]�i�F�DO�Zd�d�8�|Nwn�E�'�I�vSj����UI���4E0릊wٶs!r5�a�����ҤYg�HE� ]r���gEDTxI��Y�C:��̶L�%5u��i���	��
�����k�=��rj��&��E��E�+�f��t0�7Ŷ�VQ~��X�kR�����V���v�̇gwm�E�*��5Ӌ�i#�o��<��vF�-zh����Ѷ��7�FF�S~��R�	�0�E�F�預V��G�߶ǆ�"��E2�5Dc�Ԙn�@��� na�7��RE�2��9w��E���x���cenS�a�7%�Ƕ��cEB���rP���`�ۑ�EY�E���9�e��iT���,��!BE�t�D��Ȟ$ݒp���9EUΝU��ݮ���G��.Z��Ex��u�'EHuE	����b)�U�ᕧ��j�;ss�.�8�bߑ�*Dǜ�E��a'�<EA8��%���kR�k�h:�V��ׁ��qz7������5���m���tg���?�m��޶e���G/�R+Uaw���=V��d��s�����ж@�uF��OE
G]��R!,A��)�����u�E�$�����9�Q�E����Ҷ/�ESD84/�	v���b/GDI5�#��R^T��H���@G�H��>��+�ȶb�B�ި��S��5�i�(��q�p���L�V�)��&3˜�}�)��昅���c�݇����DѶ�AW��EYF�vy�]g����*�x�aG��iN�
��m3���-� U�W���@�Ϲ�7E4��L�G����}���E��Q�3�D$w�[�!X)G9�S�sv����A�(�{����3�z�w��&y���g��L1�<� <E4��N���U�z��\E�mp�E$v����4GC�EA8��)����u�����G��Qs����t��	\��0N䅕㾬�|L��;�b�v� E7�1N�H�~��O�V��9�V,�B�O˳��T��
�;'���#J�٦��E��۸%Tr7 =�U1A�s%\Ak [(��H�f���KHE�O����"��E2�?@��.�⪎x��S��^+U�w��&h��#��P�z���4C��Ip�5��G�/����
�䙥�L��n̶	�1�H���������2�#��D��^�e�FW`[9����ꙵ�S���׶^A'�h�
�����(遶�l�g{붲���!�ƝGe��n�����>!Ծ�>���A��2.�jT��sӶS��t.E��+N��K�<L�6��8ʁ`S{����C������!�7�Ge�6�T������K�Ԥ5ꝵp۶��7�m�fG�N�LG��q�5�`��TF+���b�^w�g�������J��$�^�U�r�bZ�
R蚹�7,�&��m�G�r�����c�pLF)�\%>�q�������_�N��r0�Bu�D�T/����V��8�y+�ŶF܁������r��G3���!�E��yt�����FE��G�����ζ�"C�ڔ��X벿�̕���E��,�*�@�����wmE�"��J�D;�E�6�v�:TF�� -0�a�=��ؐ DFxH�l��U�xD�o�����v�8��1{�)�f�f��@G�����ѵ4G\����傹�CEЅ?M�|�sY�����Dж[}����V׎E�P�zvZ�n��F0���������� ��x�%��l�zە�M��4�wf�3�d�u�kL�ζ;�V�ө25^�4�d�� �E���طض+Ҥr�R��,�;ύ��3�W�E��\\u��S��R������.��T&�%���l�V[]���ǒ_��_%鲶ϙS�s�%����i�\�v_K#�O��E�ʶtޔ�qh[�F�B��EF�Vk�H��'u�'���D����H�1Ն��E���م��ӯ߹e�u�Ҷ�k������K��X�8Y�!bE�~�ΙH��BW�@E8@�!��RG|���9���X���OW���v���b$ڒ�{E�FE�  Yr��;�b�v� E7�>Bى�΄�a�~� �6e���M�~��',�Ú�CF��\u��e�7lE�LNn������H��Ŭ��mfEN��Gі�$�O������>�V�҉�ݙ3�we�r��x�F�15Ν�H��7=��$�U���v�����ɸX�kء�&,���ٝD�{���e-��F��E� Xõ￈�v@�z�n���sT�K��l�c��T��v✶T+U����E������n� �����Ji�N�r���V����!,C瘉�n_��lu�T��2� Au�Vp��{ζv՘n[u �B����C���-�-TD|�D�5����LE��wP�\�/�YE�D�t��lΆx��ﳩ���z��@�pFg������&۶��x��E�j�r��͖���~�����sQENzԛ,�;�ة@�gP�5�����5F�e�죗�۶|Pg�����K�g�M�����v���E)�ƫ��r�=E�fM����)rE@�s�����Vm�EkM�����B��-tĩg��EE���$�{#��ζC�"����C�Yqp�F:��q,�u��t��m�[��y@�Xε����#M�Vm�r�*a�Ǝ E�i�cؖ5�-jL�BfE�SQ;�h;�� 2���E̶_ꃶ|.'�!BEͫ�ڟ�=���l�E�(�D�t	�	�D�F�W2'���Ni�|�c�k�_����~W��OE�y[-�%Ŷ��P[!�X����5�p�p�f�G�D/��,�Ҙ�c!�C���9�2|��,�b�v�pE+�>O��� �E��{L�öIb5r.nwF��n�����U:7��iT��d}�	�D��&�����~�^�V%�!�\���GҜε�w�3�H&��|Q��g�,��$�f�}�R)�~{� ���n�D�_O�����G�V}5����0Ks�]xg�۬h����U�����w�d�F�i�G]���b_�"�JGY�E��<t��������E��si�uN���0��èB]�XG�XE�A�SseE+�+ՙ�r�&,�y���+DT4�mG7{�%�G�����)��5E�� z����l��P@���in���lꭵp���0�3hYi�cJ�E�s��@y�#:G�W���)�$��G0bC��zE'�EG�NS�`͚�Ƙ���R�&� ��Ŏ�O�׶�`8OK�ʚ�����Ŷ����?U�ic��x��&!REީ�gY�i dE-̶�_A�?h4F��DfT��s�c7�h�,���]x���HӨ*T?��f�%0E�J�d�V�a��I�߷eS���8rrE��{�]�N�/�z�H������n�,$T�IW���l�F^�[�	�F7�9u�6D�r�m��a��*{CI����yh�feŶE�o ���h��&W���?���
M��^+����`�$��#l�sZ�"^/=�Jj�BA��',�~���,�ͶF+���r�&,�+���n��Ն���1�#SG��b�9�t�X�*��VoF�׶!�T?L飡����p����!Qж�[ق񪖜4�}�E�f��(ģE����;��ֿE3�G�^%,��E�
���-���E�؊-:϶E���(��E���
���z�~�z���:�j�^&��?�(/�/asd�a�E���0�/isll̫�Ӻb�����!As�/��)�E�7��E���.IC���>����SFlH���Ej@AF�;a�%As�)�l�a���j�)�l�a�>�VF�7��U�,�4�-]��E�Ȋ�ɪ��E�/Asv�M؊�(��b�����E����~�F��@�E������(��E���Z���z���6�E�)�n�a�s�aA#BT�breQ��t��g����+����!ysdkA��*�El�a��sA��O�7*���r�aFlH���EdhA��
���z���0kiA����-Qs�O�+�)T�)��%Asj�a�/��-�E�7��E����؊��A��.�-As�/ysdCA��j�s�����$���Z�7��E���b�7As���Bv�M���
Inۺb�����!qs�/��)�E�)�n�a���喖��t�{C�C��A��.�-As��P��
�Ή���z�7��E����2����N-�g���r�7As�E����E=���E* N���qs�7��E�����A����-As�O�(嶭�sM���EjEA`يtc��qs��י��j��@b��b����#=W�WP��:�ͼ���aq���/asj�a�7��E����)s�M���a�ikA�Њ�	(��E�)�E�-Ys�O@)嶋��m����+�E�)�n�a��/��*�E�7��E������-���E�����k�^�/���zm�/asj�a����E�',�ݷ��+',��/\�q�a�sM���EdmA��b���z���0kiA����-Qs�O0.����/��E�uA�l�-As�γ\���Ό���b����s�"qsdkA��*�El�a��A�kCA���%r�a@lJ���EdjA��z������-klA����-is�O�.���C�m� W�峮C�m�=�m��$�K�m��m��~�/�m���m�])�U�m��m�n��E�m��m���?���m��m"�g�m�'�m�aڸ��m��m�2�ϭF��W���4���Su�d��a?	���5�Ow����ۣ~Ж�-�t�������u��R>��M �s��2�8��Ǉ�x1���Z���T��K���]�'�����/嬣�E�it�­Ei�E�O�/e�uh�E��EM�E�6{`�+M�/�Oa��T٥��E����E���J��E��.�E��ȍ��^�/As�/qs������^�i���^��ɚ:�ɒ����ˑB�o�|x�o�Wx�NV嶰d�R�)�%�7k�lVS*�7"���B�qttx­��`�Er�
­v�s|\|­�b�/�u��B��7��D�a�kj�P���Eʃ��x�����kd�yީ��kB2y���?s�D��Tx����ǌ^�)�l$�t­����+]��#�E�6��P'����	C�z�n�E�/��ɑB�<��0x_�)�M�Y�j 4�@)]4G�B\v ֋`�`��Ph-قz/BLo/����Bew���	��G��ij%�Y����m��od�i�.��h���Ph-قz/�h���.��h���Ph-قz/��z�j/BN��cr���v-�bG2ԃj1�XG���{;��	���>���bG�BG�BG�BG�BG�BG��G����^��>$��Ğ��M2�G���l��M-�x��ME�G9,��]FP�>$�C���/FP�>$�C��^FP�>$�C���/
{9��ﻖ�|��M2���]�EGC��^i����^�F�G9V��]FP�>$�C���/FP�>$�C��^FP�>$�C���/
{9��ﻖ�|��M2���]�EGC��^i����^�F�G9���]FP�>$�C���/FP�>$�C��^FP�>$�C���/
{9��ﻖ�|��M2���]�EGC��^i����^�F�G9m��]FP�>$�C���/FP�>$�C��^FP�>$�C���/
{9��ﻖ�|��M2���]�EGC��^i����^�F�G9��]FP�>$�C���/FP�>$�C��^FP�>$�C���/
�,��V?G���x�/�M��JM��x�/G��G�B�܋$N�bȍ��<�$N�3�R�B�wM�!��ϛzG��WM�!�B ˅BG�,���
*�	
�,��V?G���x�/�M�JM�r��>$����^�9y��]o�Bǁ�����K9���]i���99$���|��M��{O���<�0$N�3�S�BFP�>$�C��^FP�>$�C���/`M��x��M9���]�V9$���@�B�Fp�>$����>$���KB����M2C��^FpY"�����/G��G�B�|��M������|��M��[&��r
"���^��>$��Ğ��M2�G���l��MF��x��M2�i���m^������կ�$N�cM��V>G�C��^Fp�>$�C��^Fpy0"���g{9��ﻖ�|��M2���]�EGC��^i����^�F�G9���]FP�>$�C���/�W�""�B ˆBG������p��M�������#$N#�r��>$����^�9y��]o�Bǁ�����K9���]i����8$���|��M��{O���<�0$N�3�S�BFP�>$�C��^FP�>$�C���/`M���x��M�BG9���]�V9$���A�B�Fp�>$�?�V3G����^G�B��BGF��x��M2�i���O^������կ�$N����BG�9���G�BzR�B�>$�EG�C��^Fpy0"���x��MM��x��M9���]�V9$���@�B�Fp�>$����>$���KB�����M2C��^FpY"�����/G��G�B�|��M������|��M��[&��r
"���^��>$��Ğ��M2�G���l��MF��x��M2�i���Y^������կ�$N�cM��V>G�C��^Fp�>$�C��^Fpy0"���m"���Nf�FPI	"�C��/��>$����/�Y-rC��/Fpi0"����^m"���4��FPI	"�C��/�Y"����/��jC��/Fpi0"�����/m"������FPI	"�C��/�3"�]�G�B@a�oo/��1�ot��d-�6 ��j/��m�ot��d-��t&�6ڃ�-�hd��o�ov.پF���qB@k׽F���v	݂z�j/B@n/֋s�m{�6&��z��tB@k��z��tBG�B@j�orԃ{/��h�G�B�W��$�B ��BG�9�D��G�B�ī7$N9ڜ�J��;�!��C�p�/��E"�C�F��
��$ ��BG9�,��9
G�C���3�_�B�V0G�]0G�B���3�G�B��" ĀBG9]G�BX�CGV�G�]�A�BzA�B�-VHG��SG�9G�Bz �B��BG�G�]?A�B�����M�G�G�hU�W��$�B ˅BG�9VM��G�B��_c�$�ZA�B<��M���V?G����/@�B
�j�u�BJW��$���hUG��G�B��G$N�BGM���L�\EG���ﻌ<��M�3�R�Bm"�EG�������M��G�G�hU�W��$�B ��BG�9�D��G�B���0$N�BGM��@U�8EG���ﻌ<��M�3�I�B�."�EG���RU��EG���ﻌ<��M�3�I�B�."�EG���UU�BG���ﻌ<��M�3�I�B�"�EG���#U�BG���ﻌ<��M�3�I�BE/"�EG���!U�XBG���ﻌ<��M�3�I�BC"�EG���7U� BG���ﻌ<��M�3�I�BY�!�EG��˼T�(BG���ﻌ<��M�3�I�B�"�EG��ˏT��BG���ﻌ<��M�3�I�B�"�EG�]G�BX��" ��BGVQG��r8�BG`wY�B��B ĄBG�}�^�( ˄BG�}X� V�G�?�VhG�?�V%G��SG��G�B���3�I�B8�BG��G��G�B��G�B��{���zR�B��$�BG���ҺZG�B��r&�e�Z�M�K���<�'$N*3���i��B >���U�BuN�B�v��r43��+��G$N2��+$N\�C�zZ�B�բ����}�����9l��޼jes�T�=$�y��9J_���G��G�&�=��e���|���<=�
{�f#������%2"��wA�BV�G�3�E�B��8ѻ����Y��k�������u����v�~jǇe��`�z?~��졜u�u���h���h�z?h���j���d��ꡙ��e�s��5��u�z�����b�v䫘�����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������6؍d5��������������h��.����C6�~z����bUv]��zKu���D\����9H ��� lV{YM��Nsz�qVJ�V�E%M����i�A=����DD���]M4��� �A��w�{�w�u���M�zK�'.�捠��*d�z����bUv]��zKb�����L[��{ߒ�];����zK������bE-ڱ�L�M��H L��捅���r�L����i�������DD���]�zKL�b�����hϚ�VN~Ľ`R��������rz�G��������������������������������O������5�")����<u�~���j���l�l�k�����z?��?h����˭�j�z!̇+��������$�s���s���s��t�5��s���s���s���h;u�s���������������������A�����������������Ϛ��o���������������������������#��������������Y��-�����-������њ�����������������������������������������������������������������������������������������������������������������������������יȣ��¥����Λ�����������������������������������������������������������������V������m*�������fr��Û�*����@���H�b���������Yr�v�����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������Ś�����>؛�����������������������������������d�ݯ���s���s���s��������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������߄|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�׬�h��y��	�X�|���|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�:�hDIi;�|"e�:O~�Y1�z^�|�X~��E.y�|�X�:�m��9,��?%��+�|��m��X��=���f��3-��F.�(.%m�C!y.Y�x�90j8F:u8!��0�5�i3-ܒ�Œ4��B6j82;w�M�l�K��F.̒&6f�E�z+F(jF�i3-ܒX�n(!̒&6f�E��E(j�/m'/o8F:u8!{�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|'!�(�8�'�k�X�|�X�|�K:j�J;s�t�k&(�|�X�|�X�mF%mh�zC��'!�(�8��,D$(p�9(�'!�(�8�K:j�J;s�t��C���L*�/y�9.ls�z�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|8��2.��4�';v5!r�f�fB6j(�)Y�kC(�kL75� y3!y�k�;�2;w�M�8DE:fF:lCL:j�J;,ڊ;vY�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X���J.py�j�90jGL:j�J;-2;��&-u�&�7M!�F�:3jG(1y�x0c�4�u6�b�2!��9 rK-l'%w'�kG)!yB0lG5,jGC-y5�vN!�A%wG2/zG::jGD/fD�vy:zy0c(�jL'y�M�z�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X���J.py/k�J�oF%m�6s�x y3!y�x�ݐE�k"'!�A%wGL:j�J;-1 ��A;�L0�)!mG7���J/w�E:�'/h:)-�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�˒71y�%.hK!��&-u�&�ێJ.py*jG64g�4!gG7!܎5;jG5,jF��F�kN!�'/h:)lG6;fD��5�FL1�F!gG5/��L/l�x0c(!�'/h:)lGL:�F;w�&0�&L1yG8/r60j���9F;w�&0�L7@�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X����x�9.l�2�f�X�|�X�|�X�'�x�9.l�2�f�X�|�X�|�X��'/w23!mY�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�i8A1w�K7m7'-uM!h�X�|�X�x�90j23!my��6y�xL:�A-o�x!s'%�B/mG5,jGE:fF:{,F0�3-yK)j5��B%iF�7"��'/yG4,fF�i5:ވ4-py0c�x y3!y�+4j�юJ%h�&�7"��'/yG4,fF�i5:ވ4-py0c�x y3!y�:j�4!̒&6f�E�7"��'/yG4,fF�i5:ވ4-py0c�x y3!y�(pF�i3-ܒ %m�L!�.	͚2':py7cM!��00y�70fK�v�E�fB6jY�j�J�i3-ܒx��6y�xL:�A-o�x!s'%�B/mG5,jGE:fF:{85%y!yB+jG��G&:y'�w�A(jGF�v:+wL.�A!��&-u�&��7"˚�&:po从J.py&fE��L+j(/yy�o5:py�n83l�x�n�9;j�^�iK0ވ4�eC/�'!�(��N�d'�v�A;��&:pY�|�X�{�X��':v�x0c(��)(f�90fK�ێJ.py:zy1m�E:��x�e51�y�݈@-m�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X�|�X��?��X�|�x�;K�('���&�]�|�%�;qa,i{t�/<�<s~��>��X�|�x�;F�0'���&�T�|�"�;%l��X�#c����Dfd(	k&���X1�h�]� d�x	������X�S��z�3�Kd?YA��^���4��8����X�S��z��Kd?YA��X�|v�!~ d�#X��p����7ۖU�|�J�j�%ɞ�0�`1j�!DG_>��q��O��p�g���h�Ɍ d�w��yS�O�|H��p��{�X��f�&�[�?�yS�O�|J��_Y�|���^~������X�|*7W��	7�O���y�NP���y�OP�	k&���X1�h�]� d�x����|�X	��ᇤ���h�]� d�x�۲�X�|z��Kd?YA$ef|���X�|�[��ӂ%��X�||��K~7��s�8�UXÎ&���/w��p����X�(sB�����%]�aň�r��O�	k&���X1�h�]� d�x����|�X	��ᇤ���h�]� d�x�۲�X�|z�a�Kd?YA&��y�P�������Dfdq��j&���X1�h�]� d�x����|�X	��ᇤ������{ d2{>��|�X�ը�Ke�Ke�|�X�ͨv�-(xEI��$d<�X���X�|GK�v5��n%��Y�|-K��k�ΥCJJ<��y��O�|"b��^���4��8�D��d�|vށ� d	��ᇤ���h�]� d�x�۲�d�|vށ� d	B�ᇤ�����1� dW��D1�����S�O�ّX���X�|GK�v-��n%���X�|.
K�,Er�b2����yc�O�s@}���Oa�f������Tfn�w�v޽� d2{B��|�X��pKe�Ke�|�X�٨Ҙ���S�O�Տbچw��O��������qk�O���X�|�%�+W^g:L��q�O�s����T{�����OP�Fs����2{>��|�X�ը�Ke�Ke�|�X�ͨ�����A�y�SdO)��X���X�|GK�v-��n%��Y�|.
KZgi��Nx��5� d2{=��|�X�ܨxKe�Ke�|�X�Ԩ�&��B	�q����Tr�	���X��F��4���+����X��>����M��B�pι{ d�U��v��"d$k����w�O�ۭ�]� dȹ>A����J̼qk�O�r����X��A��<���+����X��9�_����B|�Xg��'|ڐE��+�	�q����qo�O�ۤ�&��g�O�����]� d�p����X��A��<���+����X��9���G�Ԗ�o�g���V,��r����X��J�����+����X��B��35�9�ة���5� d2{9��|�X���Ke�Ke�|�X�ب�_1�
����q�O��d���G������D�Us����BJ�dF�H��,A������~��b2����T�4	�q����Ed��2{<��|�X�ߨ�Ke�Ke�|�X�ר<��9%efZfaϨs6�����|�X�NJ^Fs����#&�ܺ,�b��8(�c�a�|��$��1z�qk�O���q�O���X�|����?L�c�|��~Q��ts����y�HP�Fs����3�d���X���X�|GK�v��n%��Y�|(KxⰑ�O���x	�P��b:���y?�O�s@}��8���&����ݤ�� y�}s�����O�Fs����#�CS����B$m�l��?�Q���X���X�|GK�v%��n%��Y�|'	KDtl��X�9�^���k� {�36d&���o��ʏ|�XyϠ�Ә�����~y�c�O�r�	���X��F��4���+����X��>�U}K)�;���d�p��'�&u�8��Oi.v���I�H�~-d�[��O�8ӆ��|��5������9���9f��5��a*ꂤ�O�w�fӆ��|��5������9���9j��5��hع�O�Խ��5}�Qx|w�(Kĝ����G�,����U��5}f�t���Y��Y�m�5}Ĝtp�'W(��?'%d��}��4}��U�E���bҶ�b�'}����Eñ��Z#rm�֟|����n��5��(	���}==�7I�	CemѼ��,��R�m�}��4}��U�E���bҶ�b�,}����E����3�:�o�,yU;}���.�H6pΡ�V��q�8x�x/�,��W�zr�8��Ud�vYF�P�fd	Cem�}��4}��U�E���bҶ�b�+}����E���ݩ��O9�Z��O�8��R�dm�>��,��	fӆ��|��5������9���9d��5³T��bX`���
k�,��R�mmў���5>�/2@Solm��Uw�5}Ϣ�� !�Oh�o��>�>r��1��F�%}����N�D��[_�^����,����U��5}f�t��yY��Y�q�5}ãt��o�uNd�U��p�8H6t5��5}���<�W�O����5}���<���Ї�f�^
��,���[�uW��a�8�Ӣ&d����r�8��Z8���@��5}���U��5}f�t���Y��Y�o�5}ǟt}I��U��z�8U�5}D�ATk@��Ш���W��5}���L����0w#Cn��^Elಞ&��[�,���}���8�H�r*d�t5��5}���<�W
��O����5}���<�����$����ϯ,��Ui�	t5��5}���<�W"��O����5}���<�PE�P��Z�,�	Cϟm�@���5}
	��^�8ӆ��|��5������9���9o��5���1OnT��,��l�E�Ҳ��8�ʚ?d��
vKo�m�5�o���EFg��ξ��,��jcѐ,���
/�,���(��Fg��ξ��,��j�cѐ,���m��5�*0b_�4���$\��Uvӆ��|��5������9���9p��5��h��7A��5}�O���سy��5x�5}����\�8?'%d���z��5��QM�m\U6~��%��5���n�8ӆ��|��5������9���9i��5��{�e1�:��Ӫbd�U���8�uNd�p�XxC�-�Zrm����"ad�[�|�8ӆ��|��5������9���9r��5³�_S3�m�x}��5}���U��5}f�t���Y��Y�m�5}ŝtZ"��aQ�WK|m��*���Pܮ
���W���I	}��4}��U�E���bҶ�b�1}���E�u��y�|Ą4
��,��R�s`�}��4}��U�E���bҶ�b�'}����E�LySB}��@��5}�b+�mѴł�@L�5}���U��5}f�t���Y��Y�r�5}ƞtڴ�®��8��b˟m�x��W���5}�Z[}mѴ
��,��ٺ���5V~�5}�	64��b}K�t`�5x�5}�C���)d��@m�5}�Og�Q�t�8}��5��O�p�N~1���$�C��OE�@��5}���U��5}f�t���Y��Y�r�5}ŝtAS�m�5}��}��4}��U�E���bҶ�b�,}����E;�Q����N���8}yS8}�μ��,�@Solm��U{�5}��c�s.7���U�ٵ��5��}$Zh�[��j U�    ]�]�l$�D$   EUô��qj Q�    Y�Y�L$�D$   AQ�J�ځ��h�*S���/�I_��k9f��Z���j R�    Z�Z�T$�D$   BR���[bU�ԣYEh  �   #�	(����   4�����N�́���@SW��9&Y��f�mQ����	   ���G6��_P��e��L&f��S���P�   �K���xf�Ӎ��%f�}}PW��_���.	�(����j h�   jj j h   ����%P�����/&ƅ�Gh�^����q��k9��j ��/&��j R�    Z�Z�T$�D$   BR�@ێ�   ��&�   l����e=�fW��<`�   K�n�C���o���o�&���)a_=�7  �m   �   �����/&�ڗ��e'��
   �.N�(�Pv�J�Z��   j S�    [�[�\$�D$   CS�}���   <l>����٦!�1G���/&���e'��j �   7�e�P���j f�� �j �
   ��-�)�:W}j j P�    X�X�D$�D$   @PÏ�ؿh��nj ��Ij `�   ��`a��3&f�ƚP����f����`#����a����[  f����ȍ���%��0�3K��)�,j 1�Uj �   ���Щ{�}F*�j ��j j Q�    Y�Y�L$�D$   AQ��?���1�   �k�Y��-R�����6j �   ���ҏ��YZ�Mj �P��y��3&j W�    _�_�|$�D$   GW��x�s�';)�P���0�����E����{   ����; &��}����%j U�    ]�]�l$�D$   EUÓTO����Ћ��j ���x��Y��Yj V�    ^�^�t$�D$   FV��f�����Mh��/&j S�    [�[�\$�D$   CSÎ�Ln9��j j U�    ]�]�l$�D$   EU�VO�?TW���$Z��'&j W�    _�_�|$�D$   GWÇ�0��ld�   ͵#��y�7v�C:�@!.P)��*j������f��P�����j ��j �   �X�f�d�!���jf������/&f�(���R��ӫfY��  )����`�   h�Vf��l�a��M u	��� tPS����  ����k�%��[X��� tPS��  ����Z�%��[X)�=�����Ĭ0H3��ǅi*   �    NT�#h���������k9�Љ��0h��������k9�Љ�9����%P��q��}�t�؍��
&P�Ӎ��
&f�8	u
ǅ=!   ��i%�   ��s
ǅ(   ��a ��Q0���& �C   j S�    [�[�\$�D$   CSÂf����C��)�]!�  `���&���!a��M)��=! ��   �������^��d&��Pf���   "v�kȲ5`j`�i)�A1aj �   �    *�'X�rI���pj ��1*��e������&��=	j�f������&���/��U(j S�    [�[�\$�D$   CS���   1������%j R�    Z�Z�T$�D$   BR�|K��|��P����ef�LB��)�%�΍���%+��Pf����)�%��!��}�� �|���
   xo�LH������Y`f���a���%�   �x�ӧ_�ֽq`���Pj P�    X�X�D$�D$   @P��-H�b�f����)�%S�   S�	�n�0�[��V�_��}j P�    X�X�D$�D$   @PÂ���=�%f�q����%P�   %�Oh#_�,V��U?��   1����)�%j W�    _�_�|$�D$   GW������}�   �#�]ͥZ�҇P�D�&Y��5�%���-��M����%���0Pj R�    Z�Z�T$�D$   BRÅMS�r��a+��)�%�GAeY��}j V�    ^�^�t$�D$   FVô���   ��e)����9�%��a���%j R�    Z�Z�T$�D$   BR�lS���V�f��P����)�%����}��U����%P3����)�%�����}���-�%	�a.����%���*P���&��)�%1����}�Ӊ�1�%���3�Uh  j P�    X�X�D$�D$   @P�+��pa'\�����%)�� P��	�5����%f��Pf����!%������   �р��& �   ��(�  +����=! �   �Ѓ�D& �>   �ύ�^�%j P�    X�X�D$�D$   @P�y��K  ����   �����I�%��P�   6����l)��d����%f��P�   �@��$��%M�=! �0   3�Y,����%`�   ����>hHV�B 4vP��5$a�	   f�ˍ���%P`���0a���%j U�    ]�]�l$�D$   EU��NX��|)^P��*_��	1P�����.j P�    X�X�D$�D$   @P�dx�@���   �nm�UU���W�_��S��)Z��M u	��� tPS����  ����k�%��[X��� tPS��  ����Z�%��[Xj Q�    Y�Y�L$�D$   AQ�p�$�bWu�   �;�SL�(�   �c��+���   �j*4P��-��{d��O���_Yj R�    Z�Z�T$�D$   BR�-4s�3�����Y��j R�    Z�Z�T$�D$   BRÒk%�_q��f��L���I�%orea��   �   ����%P����%P���%P���.��ƅ�DhO����q��k9�Ћ؍��%P�Ӎ�I�%P����%P��=! t����%�����%P���%P���.��j V�    ^�^�t$�D$   FV�O�6T�@������if�2�%�   ������'   f��b(ǅ(   ���}�%#�)�S   ��'?l��=! �4   ��y	��I����%�)   �   �<��O�dt݃�T��l	���� _����%���$�����%j Q�    Y�Y�L$�D$   AQ��f��x��=! �1   ����D& �)   j S�    [�[�\$�D$   CS��؀w�  ��.�  �������M u	��� tPS����  ����k�%��[X��� tPS��  ����Z�%��[Xj P�    X�X�D$�D$   @Pã�D��W��`f���f��va�����#�Q1f���h?  j Q�    Y�Y�L$�D$   AQÙ���\`�   �   ��2N�Nr�D@]Y��aj ���)j ��%����%���   ����A�%��)��-/j j P�    X�X�D$�D$   @P�j~��\����j j R�    Z�Z�T$�D$   BRòj P)�U$Yj f�9j ���%f�ɗ*P�jf�ȯj1��,j���h� ��E_��=! �G   j P�    X�X�D$�D$   @P�I���pD̋�Qf���Y����%���"�$   �����=��t�%���'�   ��"P�׋�AP�����A�%j P�    X�X�D$�D$   @P�N�����$���-�%�   	�1%���>   ����q   j S�    [�[�\$�D$   CS� �~��S�.`���JN`��aa��E�%�   ���?��"A����='Z��E�%f��ż��U�̅��   f�=j)�Q/��=! �:   ��)����%�   ���?   j W�    _�_�|$�D$   GW�=~�=��t�%�   )���   /�Um�4P��A�%�@�:U��9�%�����   ����E�%f��-j ��}(j ��M��E�%��Q��1�%��u���   �   `��%��a��E�%j W�    _�_�|$�D$   GW��~�if���;`�����$a��U�]���   `f����]-aj ���"h�   j P�    X�X�D$�D$   @P�Ջ�"�   f����jj R�    Z�Z�T$�D$   BR�E�K0j f��j �   g�j�
���n� h��Eh   ���	��\����%j V�    ^�^�t$�D$   FV�hږ��f��������/����  j U�    ]�]�l$�D$   EUØ%��   ��9�   �z��X#	��+&j S�    [�[�\$�D$   CSñIm[��+&��  �ύ���Z ���j V�    ^�^�t$�D$   FV�ҳa��U����Z f����j P�    X�X�D$�D$   @P�/�����   ^v;�2xҙOǬ�R��M u	��� tPS����  ����k�%��[X��� tPS��  ����Z�%��[Xj P�    X�X�D$�D$   @PÎ���G��޲�)�%��f���h?  f��j �   ��q*��r�TƂF��Q�)f��2Yj �����"��+��)��A�%�h� �   �e��=! �Y   �   �   �{��)zrx�2�s��⍅��%�   f����5   j R�    Z�Z�T$�D$   BRÐx��6��)��t�%���P�	   ��=�Im[����A�%j R�    Z�Z�T$�D$   BR�c������,��9�%��e#��E�%��ǅM     �Ń�E�% ��  ���*��#�%f��P��%j)��)��E�%��m��=�%�   � #�l�����}�$A�����E�%�����Uj S�    [�[�\$�D$   CS��`��%f�9lah� ��=! �2   R`���$���aYP���_����%��0   `��%��Q"a��t�%j P�    X�X�D$�D$   @PýP�   1ݾt�|:,����A�%`��ы��a��9�%j W�    _�_�|$�D$   GW��� �����E�%�5(��E�%�����5�%�   	��(��E�%j P�    X�X�D$�D$   @P�/"���ƛ�/��-|5��U������3�!���&�   )����y�����E"��a'�a  ���C�%����%f�;����   ���꽽�Ԃ��
j;��   ��/�o(h�Zj �    ��Y�����`�   	 ��<X����G!k�ya����%����f���   �/j �⑥�_��Yj V�    ^�^�t$�D$   FV�21�ɤ�!�������Y��M u	��� tPS����  ����k�%��[X��� tPS��  ����Z�%��[X��f�Ћ�)�e"P1�+�؋��!S������CP�CP��'&��[�   �Rn�rـt�$�
   ���^Y*�Κ��j ��E%��'&Pf���j`j S�    [�[�\$�D$   CS�z��'|S	�f���������=P)�1'j j f���h   ���-S`��=(��e(a�����A��e'�ʀ�����&	�m��5��y��   1��ډ��N���j V�    ^�^�t$�D$   FVî�2��A�@�qǅa    ��m.`1��a��=! �+   ����   ��i0=�   ��  ��!�   �    =�   ��  ����Z j S�    [�[�\$�D$   CS�N��t�5&�   OͶWi�E�-ڙ��M��j S�    [�[�\$�D$   CS����&�v����9+����Z j W�    _�_�|$�D$   GW�\�ڜ�f�� ��j V�    ^�^�t$�D$   FV�F0�������;���   ��c��M u	��� tPS����  ����k�%��[X��� tPS��  ����Z�%��[XP��-&Y�����f������E   W��_ǅ)&    j P�    X�X�D$�D$   @P�譝�ε��  W��_�b   )�����S   j P�    X�X�D$�D$   @PÍ�% �?�f���  j S�    [�[�\$�D$   CS���   f���_�����u.�������M u	��� tPS����  ����k�%��[X��� tPS��  ����Z�%��[X��j W�    _�_�|$�D$   GW�KXI֧(�ʹ���8��	�Q�O  ���+&j R�    Z�Z�T$�D$   BR�����.I����I��#&�   ������H   ��5��3&f��@P�@��GY��#&j P�    X�X�D$�D$   @Pè�й��p�   ��j4��uP��#&j ��M���b  f������   ƅ�VhR�����q��k9��jh   jdj �Љ��&ƅ�Gh�����q��k9���Ћ�ƅ�Oha&/������k9�Ѝ��&Sj(V�Ѕ�u ƅ�Ah�d�������k9�Љ��&ƅ�Lh�礀�����k9�Ћ��&�[S���&Sj �Ћ��&�   �C   ǅe    j j j ���&Sj ���&���&ƅ�Eh������y!��k9��j j��f����u2���&�C    j j ���&Sj ���&���&���&��e'j ��Yj S�    [�[�\$�D$   CSö�aǞ�CV��%/YW���Z���9&f��Pj S�    [�[�\$�D$   CS�����d�5    j P�    X�X�D$�D$   @P���e�K��#�5	���Nd�%    �
   ��.JĈ�5���� �e   ``�   պmN���H�`aa��%/a��i*�<   ��M)��q,���
& �#   ��n6��  �   uD��$=�{H�k$�p�k�3�j R�    Z�Z�T$�D$   BR��	1�A&3�@?d�    ���   ����Jj P�    X�X�D$�D$   @P���   ��������&G�]{�����   ����*  ���s   ���'�L$ǁ�   �������   3�Ë\$U�    ]��:&���   �� ;&���   ]3��j Q�    Y�Y�L$�D$   AQ�l#�JZA)�/��%��:&�   ��V�}Pj U�    ]�]�l$�D$   EU�5��r��a��   W��Y��q(d�5    j W�    _�_�|$�D$   GW���/>������)f�5�d�%    ���!�
   ��UHd���eԅ��@�4 ���_4 ��hXMVu
ǅ%	   d�    ��j R�    Z�Z�T$�D$   BR���beP��Z�   �����   )�9Z�K���   ϔ�c��_�   �   �*N~�"H0l�[�Y��A$��M u	��� tPS���=  ���&��ҹ%��[X��� tPS�=  ���&��s�%��[X��7M�T�    ���:     1.855                             Exception Information Please, send the following codes to info@oreans.com. Thank you.

        (press CTRL+C on this window to copy to clipboard)    

Version  = %s
CheckIN  = %d
CheckOUT = %d
ProcIN   = %d
ProcOUT  = %d
ExitIN   = %d
ExitOUT  = %d
TPin     = %d
 ��m" �-  ����%P����%Ph  �����%���;&P��<&Pj j ���%P����%��9���;&P��<&Pj j ���%P����%��9���;&P��<&Pj j ��g�%P����%��9���;&P��<&Pj j ����%P����%��9���;&P��<&Pj j ��n�%P����%��9���;&P��<&Pj j ��v�%P����%��9���;&P��<&Pj j ��}�%P����%��9����%��E�   ��9( ��   ��i* �   ������  �   ����R4��@��;���,���, �U   ���,��L���<&���,��P���<&���,��T���<&���,��X���<&���,��\���<&��m" �   ��9( �h   ��<&��<&��<&��<&��<&��<&��<&���;&P��5<&P���1P���.��$j@��<&P���1Pj ��Mj��Y���   3�#��w�4�\���^��#r  f���    �   ���<�   f��V���u�R��� J����<�;����_!�٬�<`�   �,=▢*��@fa�Ӄ��KKKf��f��d��������f���y������������P��|�=i���:f+P�De/����NF���}e/����NF���}e/��������QF	���mr�D�������>������q�D��K�������dN��jm�j�M�v�A����r�q�d6������_9��/���T�1j�T_	|��i6h� D`�(�D�\�C�\���)H1�����r�q�9�I(/���E��,g)�M�����_����C�y��r��ù��C����E���L�]����y]6���(b�/|���t_��h�Ƃ�E�B���5���t`z!�����z���XǾ�������N�M����M���O�x���~������g]�a��|^/�W>XĤ�/�������n��^����Ē�&������4v_4G���6���64�,�QրbG��1�����������e4E��	�K���(boD�����ibkD��щ�&cjjkD���<��YÉ��C���I�#��r]*�YÉ��C���ŉ�&cjb�D��ŉ��?�^���Q`�l1R��������B4�J��L���O���Q`�l1R��������B,�J��L���O���Cx7�Z�l!Q���qu���8����4߅&������4vb7�Fjb�F��ŉ��?jb�F��ŉj�?jbCG��ŉ@������%��d?�P���/ЉF@jb�ē��l_���S`� gZ�G�����@�����dG����?N�	�棍_�ҁD�v�7^�f�D�"E�*�S^�lr�G�㢍_���rI�*�˙�?fR0|�ř�?�d�|����?D?�L��^�?jb�=|��fb38|�щ='cfb�0|�/$�����������������97�}���F&��an��H���vBD2й�@��Y�,�c6�4H��F��T38|�}���JIoC���JM��(����(�E��4�)��	�K��A΅B���%�T�N�����3��̃��z#G���f�h_�f�J~�q+\�8s��mF�z��H*�b����.�k*���v���w}.��������R/�IC��^�M#M���xz�'mFϥ�vR&��b;�O��7�h�
������3�q*:��-��h��1��)aW�+G�Yr�^F�ޟ��@_��d���]Y��F?��s�@���E9�ǾzX��0+����O��i(��/����~6���`g&GK�L�R��,��0��I#�G`�fhӕ7E�WHU�_���dH��uo� ��	��d�!_V��3&�/�R���lxH+������F���`��y�6JN��?��c>���h��1��c\�7m�������'����O���B2+�c��<	Q����z�>~ǀ�AE4h:������N��{�.�i��Vvp�Sy$%��*�ˬ��[c�!�T���G��f����i�ۦ�=#�='�w��+� !1��#����z���Lj7��$s�8���7uN���aU4���o�����ƾ���Ͱz�L�i��y���W�Kޜ����&0�n���Cb�T;Qp����.���zc��6���䉙c�%�a����*�����Փk��F�����p ��!���6��9����uT>0{�����^3��!��5��'��X���F�U�.9$�����+���a��s�\L{��6���n���!���8�n��c}!���XW�����jD����S	�+4�VI���Uq�l��<&cL��A��7�����Z�U}���2
���;qdh~B &4𠵖����[_'����X8��9Y�G �t(a	w������`��	��;�4�����.RA*��4���(	�)>+��y����I�������d�5��A��r���-[Q�������-�,��Xq�{+�7��񾿑�-$0���b�V̄O�6c��l����������=�L�A������+��l�荒s������p��\|^�7�����c����	i��F �	�v��ga�}x��&��aE�J��>�ACD����$	'-^ݹ�$A���(��*H���Y�w�����}�I��:uT��7�Ҷ�����Dΐ�<{T�����bj����a���D�����4�F�:��T%���;�.���_'�P���=N�F���QA���	������(A��V�F.����1A���缩q�%�p2	�Z!Ji�3;�6!��W$��<�.-\R>%��I�Ս�,s�(�V,V���G&�f���Q��z��Ti�ت�^�"�:C��P|���-,3noT���w�fj;P�-.�<�i�}{.B7��;��5�󖿱�7��5g����X�]�G&��s���(P\�v<j����<�1��.��i�Z!�.9f��)�������p��=�uN�9�A�WٌQ�|q����������":Je�ב���=#�1d�b�����dD�k�$�l{���Q���,_	�r�﫛�b�q�i�Ĭ'12���ͽ�����"���eA$|fY���n��̉�"Y�*PsU���t0�Dt�9��&�F��g�+g_-�8��
|4���4*��iBG�Y2I�Ů�n���F1��0&o�Z	���;\B7�q�ݱ�&1�7��AƖsjn7�L�������ƾ-e��	�S6��F,��`�P��]��#���nYVI��d(qN?��J��Q��<)z�e���X"t���E_�Y�/�2	'-��������'�0��v�MT�K�\�(	���%^����:�$����J����nשD�N���J$��.����;�6,�����+3U#���f*�Vd+�'��A�|���/u��~��Z����>����1���ţ;��I&�IG���`	���'f�;�R�#�Q<׼\���E��'���^�����j�%�aF�{�r���a������� +�����1��(��g� M��6�8=�*�Ŭ�d-���~8��B`�a�0���
�C�x�H� n�����a?���cdN'��%��'�c�^��	z 
G[�EH!��̳4�8�0v�(�,�7����	�]&�ch��H�
T��DV����f��M��j��?�Q5�G*�"c����]���B�&_���@��ތ���ӎ�-���>X����}P���7�Y�|�D�i���G�&A2/O��� �J(��������f-Z�	^�D��]��.OM@�������d�8L�

y����-_�d���xw�~4��St�r�%�ׇ]�]��^7����8��*}4���t��!͢^*+�α��,il
_�+�6��d%�����O�;Nݣ"��_ �A��s���n-�<Z��o;�#-���t����G��!w����s�X�R��Ph�p|b&������l�o��]�u�8C��^�!V%r��Ak�/���?�	G^�-eRь[�����^��K2�B�-q�7������pJ
�]�<]d��Ў���-�fŞ:5.YRѕJ�s��
:�}(b5�.���-�C�H/&A#
JG��M���.��42����!ks>[|��$�B4
�h$-�=^�#cV������+��V��m��.��8K{~��*��Rܵ� ;c���T���}B�*a�g�E�������Pw�6��i��k����&��=���&K�)G-��O�D\,!G�:������E�&��l����g@_-��
�|��;\��3�:�P�_�Y�'%44�͞���2ǞQZ�{7�z�C+M<a!�W��:���=�-��VZ5���?N�M*��m;�h�m�����0cY�Q*P:L�v�Ʒ��2��T�C�^X�MZ �[�R}������࿵����
p���"]��Ӈ���:ܪyP!;v�F���1_��H�a�
|x�n����Ͷ�۬�r����|�z���0�/��.%p��?M�!&m��3��9PJ�$s�8	ښ,uN�� .�\��Jb��+�V-���\1����2�U�����\������K(",�.��"K��V�՝�-�DG��������G�h�m������bV�6lFK�v�M�Y����U����>��x	G&�������D��������v��tPa�Q��GɌ`��CT�hH6��T-+��J
J.j����
��W��F�����>W\��� �])�4��g1h�h`A^�	��t�I������,����x�� "Dfr(��M%6f>��=_t�I�����~[>�~�����n�J�����cR(=`R(8^%�(��gh�h`�l.��lt�f�hl�ff�hl"�f�h�����m�se������,����fi��I]t�I�}�E�Y(6h
��h_t�J�S�P��n�J�����cZ(=^Z(8^%�(��g-h�h`f�hl�3f�hW
i{E �.�H���]�S�Me��-4��<�8�g
n�I����eZ(�)" %E�c�"�(��8���n�J�����c:(=�Y(7h
Ɛ-�ey��h	������cB(=^J(Ie:�]b(C^$�3��e,��������lH��l�h�5��eX�G����u�������	w������>l�h�5��Y(:h
��hcn�J��%W���)�����]r(I@]�]:(?^(�/��e0������}�D �^n�-<�=z�}���wcf0Fc��h_t�J��z��h���2��0�
&������;J6�H����6���H��5W��rDp�;K��W���+�2qO��W��W�-�U���X��"oK��V��OY�����DD2`��F��%���n�J~���:f+�BD�a>d����"�=�oG���J���珓��|n���Ce̺u��>�
����:H�i||�p�~�4o?W��G�qd�ac�ri��1��C�/�Ŗ�HP�Fn���Z��-��E���PF�3.P'��MbW_!�M��v�.v��>��Z�����nR	���4�˵ŀ��FPGb���w�����;=�FhJ��M�S��Z��Q���TF��E�Ļ>��:\7�H21�\���,�i�&[+���M�A�[�w��ޠ��H������楜1�Z�*b����6�|n����y������a�n�����y{=���H��x��;Z?�zg�;����S�*���v�dr����K}<ݢA���qWv�y��e-��>r'��~�p_xw�?�"�Fz�@a���]{���7s���v��N(�:��"_�͗�dK$�	�f�Gb����!��7����p4�\���^�T�-�������"փ|4����榓:�'����.D���T�����x��>P�Fn�'����!D&��_��Gag�g�&CRb��B}���dw,b��}�Q��e��t>UJ��-Մ;<��4�z�@�xt�]r�&����F���n��9p#��,�\_�@�|n����J�擇��d��C�Q�����r��uC���*��^$�����e�1�xK�Y�!��E�p��9}'^��~>�߿��D��5�V�AIP'�C�lX���*����q`���N��,Q��\��������>slu]�#�H�L��gO��C��P	�����֠ca�XDuBJB��懪�5,����І��
��T~�Z�.�&�s ��T��;�[�rC����@�u����� ���:0J=�����:�������N7n���v�PF���Ӭ����-
�v�blː�D��J�CW����:���;��!,�H5��ZG����-�.�*����FQ���rO���1�_�L����_��[���L��=�/����d�w���V-d�������DE�g������ ���;0Fa�B�Őq�p��U"��G]!4q��^�u8���������\^Ý��G�	����C'-���4�A�?�yp=�<���s�������p��;�_���I�@���b����RN����m9Ԝ8��V��
3\�[!^0��3���p���+�`Hp
�O��(.�����d�S�"C��V���b��B��;[+��欔a�o��p ԑ�<�f×6�A9Rn�#��5��2�
���~Y��.;&�|z�n���!�h��H� ������(:���Ӧ$-{�H�Mg}d*�Wm�;G[�7�Op��}����F-������{��vaW��q`�{��O���(�3��'Q����e����s�d��xˌ���g� �,|��e��X���Ɲ�jF�:�P'��IU����H��2��|��-'�|�ꠜ�ӌ:
m�������;��5��JGd;����C�����4���c$S%�@ ���υz��8����x+i�6�~�6����B���Cκ9����a��?���Mr�����+q��ܕ��&�j����$7a�:1Q�L�@j�(R��@`P�I��^����~ZN�z�?g,f��c��k�TF�;���8��3!�܉#��;�)�x���S�&z�&����/��QĨ���1u�`�DM���̝��H*��9�s������q�'����P�L�[稁7sO���-���{7���AG7u�� �뼴�;��[z����%g����q�1G���'���M��<�#��(���ˋ��A�+��@FM�m�hl�X�|��`��ϖG��Z���f˿� _lYfY	�=���Fۃ��xAE@k�T��ah���	���_%M,��#_��U�y�V�d�����ي�S	q�/�R�*b0aG���IH��.u*�F"�`I���]u���]��X�p�G���<8Qek�$-�����T��M`n�m�Nx(��ż^{9�1���2E[�v�Pc�Xc��g�tL$h<:��`G�G�_&/��WO�q�W^ٲ�6t��B�i;���bp�7������f�'�z�v]�Y��JHREo�X0%;�-Ze�h��^�Tbݮ��X���Yg�����G���B�lD�%������qE$��E�������-4��Gz�Tp�MbNF­��lU��i_p��F�1>����ZI~�q�.i�A�6�3��>�p���1.6�{��ӿ
}�F3��׶��HPTa>������$7y�;1I\�c�a��pg�p���V	߬����,;�&[������NE�=na����L
�3t+"��O���Ӳ�xڰ��Iq�a�_��;�aj
�ڧ�T..���T5��j�e����+qq��Тo�/��q���|}��Y��`���g����6G��<ԏg��"�H���i�됸���wk��N�Q�tU�li,{��Clg����L���wn�gPz9�_�~�(_���u]s�bi���P�)�k|-���HGU��W�)��&����e{�q�����j�[��!(�\����̝q�P[�����2I�������c�A ����gc��FԖ�Mй�H���S��T��N�u_L�,o��Y�6M�"BL;y�K%��V:���e�z:��ތ�T�V��^��FN��C6Yq��g ���Sց�g�h���q��J��&�F�i�T�����^1/͕�p��%�;�aIr
�|OE �-�7a���P"�J�AN���~���*����i�r���'$Ҕ�����A���qW��C��@��Q������|��1֤�G����,��P�G�i�Az{7��AG�(����kJ4�
�J�\����8��g�@��Pe�و��������H�7�f�~�6E$	�-�:��l��Ӫk�O�A�����;vTJ��AդB�瓋6�s����1N��H��;�H�[�D�C��]~t~��W���O9��m� �h|>��~j�i���6�|n�G�"z��`�P�v:���Q��:��#:����N�R��&�����J�G^�1�$����)��S���� 
�I��k��X6�s/��io��BCg	���LQ��"�PGk�w��L���������L�S9�|�C�;�����.��$�*�w�� �
�:$XP�=��]Q��&�L��k:T�����Ng h�D�*=>�=���횱�RBa��%�q H�rk��M �PIa�|�l��[Fb;�v�^���~F���QG������A���qG���b7�H3������C�5#T�J��&���V�s�����=C�	����u�Ob�@G�A�4�I�v7e񆃇����)�T������F���̌��(�.�z;�.���h>��"�����<��g�A�q�u��X�geVgY��*��柔9Āã��ڈ�c�� �p>M"a���ٶ��<$˖����&�i�q�n�G_"�lU��i_W��F��O��3eT�@ ��C�֜���ioW��u'���z����?��ؼO(���C��!pEZI�$����z(�B�\�e��s��Ѳ[�Bv�LP�$�$'}����잤��,*�3i_�Z����G�ź7���������׃y���W���B^#�2��g+B��(�	��
�?����s��h������8�
� ��]^�=Z:y�}����A^&T (E\l�hWf�����t�J�}���t��h���(��@�
&T����-�[f�����CmJ��e�Odb(=?�I������n�J�����h�h`f�h[0����e@G|s��iL��eh�ΫU���&�]f�|Xl�h�5��>�:����[�l�hYf�����n�J���0�
����n�J�����h�h`�{,��l�f�hTf�B��1��h�h`f�hZf�����t�I������Z���C�,	n��5!�� �3_n��C����;p�D�m�9�@�g
Iq^�]B( $E��w��h���/��c:(=`B(B^#�2��gh�h`��*��-Yf�����DpJ��e�<dr(=?�{���������g&h�h`f�hW��ױ��K�j���<f2����������;�����fE]��h\t�J��5�����}ŦB�+@0�O=8^%�(��e-�������t��h������@�
� ���n�J�����h�h`f�hl^��El�h�5����fi��Icn�I��� �[�l�h[f�����t�J����}w��h���/��c:(=�����Y�����v���������c:(=?� ������n�J�����h�h`f�hV�4x(������h(|�l��/9�A^�����>@)���(�gJ(�	x�����l�h�5��Y(:f
���u�5�%p����m��?+* ��c��66H%�c�Dd��2�ctEd�r'c�Cd��rGcDd^��EeGd�>d_��V�Ad�=d��ߢ*��	���v��|�eic�π����n��梏��K�&h�b4��_~���������F�_���q�f+j N�Ft�fM�a��.������N���I`�O<���b����ܸ�)6<a0�4.��>���K���S`cl�7n�_�:	dn�xL�}��M,��e0�2U�jl���SHfIq��V�k����	�������t�IS�a���rxf�k��]��xoD�N|g����˝vV����
�#����D�� 7���n\xf��xf��xf��xf��xf��xf��xf��xf��xf��xf��xf��xf��xf��xf��xf��xf��xf��xf��xf��xf��xf��xf��xf��xf��xf��xf��xf��xf��xf��xf��xf��xf��xf��xf��xf��xf��xf��xf��xf��xf��n���^��x��/X���xf�M�ޅ�K�P�I׆�K��tIg��ϻʰ�=i�X�ؐ�Y��Kl� ߠBk\��x�>�	���N��I���7S�l��G�M��b��o�2���ˢ.��ʆK���֠@g�0��J�����b��ek��uKR���Xg���e���.�;j��&{�F�ؐ3f&�%f�,øW�x4�	�T���&
��ȵux�4�f�^i��ԫ}�3��ˁLO�K/Vh�M�e��:��	����,�Y�JM�C孺���kxf�Ԧ�B�h�]}
�9�+F|�s��T�fn�3� ��֦{���4��x2�qf��f�iH�˱�'x��6wTnx�V��e1�h�:Ga�e��	���˘O8q�hƓ�p��h�ʤ��
;v��������}xO�2fʘ�Q�.e�Z3��˧��P���xhj��h���K��^ڕ���`�����i+U=ذf��N����g1���ˤ�j�*�\�h���gk�ϫ{����D�g������%�h�>�z�f��$C�ʟ��G�/X�ț�Lg�F��QfFexm�YKks0���T�f�߅9�vD��e�X�Ge.fV�9ؿLg�#m���B7�yh�˫n-�F9�(�f�0�f��� �¤Y?]��VٜP�Er�xb�"�f��6RW���ߓ��B���uX�(�<�f��ۤ(�Ig`�(��zץG���,�hٙKz�/x�d���� 4�$%�˘f�*�����`��I�P˩��ʟwr����f��'���e͌/�˟t�rG't�h0fDt>���3�G�o���\�<ً�����f��8L�f��|���Z����1�Y�����fn�3� �צO��M��X�v�>׽�h����?_��f{���v�/f������if��9��ef�GN(�p3��G�w;Zg~f��:��3@V������@���U1?g}�N��%�g���3���$q^�[�@���h�Z$�������~��i�Sʁ�x?T�fz�����h���1������W����mxfɸH\�˟���W��ˢwvTgj�ȡⅲf��N��Sji�޲7��W�$�0V�ixO�.fn�3�˥׌O�ˬ4��x�8�h��f����#YgF��E��aZ��@���h�oxf��Ygǐ{	*K�$�ˣK�Uu���K��f�����ŝ%��x�M���	��ȵEx�7�f���M�.S������Xs�rG��˘f&1�f��gk�A
({w��ˤV�Z��ֱ��ðLg��eEx�_g�b�x���+��*f���gٝ.f���`;�&p����t��G\�c@g,1�e���
��)0��G	�G�*�2������Zxfˀig;�&������V�
�7خL��3�h�˭׌f5���˩�f���̸��y�f��Ui�����3���p��P�F�LxKd��f{_P'e�e��y�e˧�XO�(�Zˡ�h��\mLɄ&u$��c�tcoFy���f,Qyf��n��`]BWI�t�iH��el�Ga�e��x��RSw�"��Y�
+ȻIg��̰��f��x�>��K�����8�Ս����xf�����<�QF���9�P̡+h�(ޞʡf����?]/0^�˃t�rF�&c f�~�h����xKB�����d-�;:J��G���fD�|�KEc�WG�i��+�X�fd����ôfz0L-1FI:���bo�>�6��Ն�/�h��։�K�v{�x������ex^���hn�3� �׫T��>L럑k����f䏅�8{(���R" �N]��Պ�F�yxf�{W��i�Y��a���fN�z�Ӛ�e�Yg�C*�Z�t��	�˟[o.����f�%�Z�?�h�mx����-�O�fV^�.iɁf�ʋ��W]8�f��\��Ս[���:�f�����n��1K��Dp +���Jx���>g��Qf�!-���m��~^�#�ˀ?�\�f�
����x�AWr���>0��U�x:h�Ig����h�A�g'�C3#�G���f�j�f¬pgJZ;�geNg��Bg+E��@����xf��̷�d�h5�� �^u��IB�+��2�h�x�ZW�e�{TK�<��}��&��f�q4&�*�T�A	u˥z�ZA�zm��p�f^��+�3�l���RI��Iu��������`g��ǝ�fQ��p`�S&��|GؔK%��f����L�&��w(��՞[��6�f��(F�3x�A׳��d(�eh�����e���h
����������K_�G%ο�H�:g��w��d�f�b�H��I���XY�x��h��ϧK�*���h���L��ۛ(��cf�28��$�f�bJ���X�c���3����xf�F��9jv�IxQC�cf�͡�f�X\�ʡf��?��>YD!f�˰�b卣�I���xf��Ψ�y�{��g��b���G�W��cf�%f��i��l��|I���_������+��0f�h��5��+����/D.�jx�4Lg�v�:�˘�W
x�^����щ��$�xf�����g������U	��;�
����h���1�wJ���xo�F3l�G����f�f�KFa�)�x��x��� f���
�[)��:g��(����{��*�t��GAY �t١f�ʴ��eI�� ˦jץ�gc;U-�\�h��`U�Z��!�����t�϶ �)�/p�e�6M	���C�������VҢ�F��xfؙJ��EO�iC��/�v�f������(f�[ �?i�����J��8x��Fw_�xf�f(��Lh�+�^iˮG�ʘ�����	�f��[(���c��ʭt��I�2!f0�f�ܡ����f�Sy?�ʣK!��J�Ź��f�1g����
��H��9׵﨓�h	hM�e�&I�O�F5�mW���,�f��ۖ�جsfxL�1�����
���3V� �ǚe�gƐ�\�+���	�ef�+fO{f�14����S�\��I�y�Üʃ�Q�Dg������x��A��H���(���GLy�hDt>��* �G�m�˱ҁ�0��x]���fn�3� ��֫P��}ւS�6r�xhj��e��Qf�C
������K�~��x�%0�e�������W<�˥
 ��є8w��xf���h�xV1xo�6��XW����BG�f�L5 ��e�������/���Z���h������RS�T˱K�("f�����~f��\�X�f�嗒��	X�j���ۄ���>gҨ֮���qI�F5��G�G��h�1�fs3��~������a�ܫ|��|xf���N��<�[w)����1I7���h:f��(F9��A0u�ʡE���ː�U�Eg��J`�I{K�x�i˦���l�.ʁh'��f�����f��|���`s��I\xq�fO�h�\ء��#��])˅��ň\�GH)3f�DUL��%�*�(�ˀ��LhL�+o��cf�o�b���'���XP8_��˥�/fҬ�e���F�6g-�B3�-��7�,cTIg�[M8b��cx�b�K���!���(���!f��ᘸU�e.�-qS�::$�t��oG��xf�TL��8�+��˳��S��%c�xʤfnT3�{)GئP�ˮh+�Q���Ê��h���Z(	�����[o���&��lf��G��B�yL˨���x����f>=hf�3�� ��yI��Ti;Õ����[�:g��hՙ� �>WI� ː��I���?;�/f��k�|������˭�-ZG�78�e.�h���ɉ�{�
�F�
�]>���/�ʐhq1?g����?�e���/�ˣW���5�����xfw�g�����]e5˧�sS�8̎x^���h��x�`~VY�2�f��>���էk��	�f�/����Xz���1������o�˂:�1?g�fx��*���G�˱eE��ُ\I��f�/��$�h������L�~P�q�xg���f�͛a����O؍b�J��T�P�@�և�h�v�\�Igo�F_�˃2��x�x�f��fz�w�����  ��tK|W�ZH�+Fg���P�d���<~ʧ
�Ͱє�u�+�f���؍���^F��ʬcM�X������e�D�b��/��.��(�Jx،���3�e z@����Ii�9eX|��?&וfn�3�˥�֫Q���e룕5_T_�
f����fVL,^��Y�����Ӊ�x�1xf�ã�l�_��Lx�p��YםI_ ��f����효m�G5���XW��
�P1�f��H\�˘��
x��7b�_X�\ʉ>�`gɹ��߇*]����|�R^x���<�%f��?���>�1�K��(8�f�yەeFexf�� ���Zf!t6����(�2⯪��	�xf�4����A�3n˫J�E��;>��0f�Ŷ���hv)y��	���fQ��ڟ�f�&F�O�Ә��-�ʬȤ�վH�Fp�xf��A��T��3ˈ���L:�q�h�H4f�R�e����bx`��`�Z�X���)�j���f���d�q�hQ�ͯZ��5��7g�f/�&f����jf�UxEQ�p�	��?��G;q܈e�Df�����z�<��_MD8��ʥ?�\f��G�N;Rw�"��V˴(��N�h2V�f�ǘ��>ϧi�E����9�����Sؙ�e��&R����x��˅z���zIA�pf~��ؔ� Y�In��?�8�vѯ�cgN�VgnT3�{)GئT�� �gϬfO38�ӫ�f�i��5M_�����`XU�fF��_�h넹G�f�}���P����;���"(f����׈Թˌ��˄I2�h��4h72�eϓP[���R��ˡ`��'fΏH��Sg��h����{�<��T� ����Ie���f�̛��$�אA5���I���f��*)of�bi_�ë=�r��S9������_�hy��"����� 	A�;���Kg��t��߼h�������DV��>�A�j�'ׇM���>g��i�����;:�˵�0v*�[��؂�e�Ȁb��zfI�(��F�=�ئn��]��{f~Ki��N�-� �˴�X�Y�׊xd-�vf�2Lb9jV�_x���U/��I�nUg�f��H���к|�_#˥e�Q�QRʩ�$7g}��[g?f�eaD+�~ŏĨy��GX�h�☧2�����Whi��tI�F����f��h�j�=�&�IF��?0軰fO���۴f�x�����|�c&�������&E�xf�eh���ۨ:Hl������x�Ixg��f��!��w<g�zM.p�{gf��M	�%�i�Qg�E�enx{D���6��htX(g�|f�G�bv�/�}�����U�78�e[U���.f�0 ���(��֐X�˂%�jtk؛F���~fn[3�{)7ب{���ذ�'YYL��h�o\ڽ�[g�����v��T�|�+p����h�,x�e�S�_����>o�nx\��fO�h��Ȳf��SY�/�U�BE"��8F�xfw͛5e��n�e��Z�{\x"W�ef�%fy���I��x��b5˱M$]�-�����en�3�˥�ֿO��Y��HG�KdƼf�k�g�`��;��˞��\I8X�ef"f����H�{ʾbQ˂��ؗ?�Z_װIg��f��E)C�I�M��}|mfpbx���Gg�C���"�FP5� �6��X���ٿSg��tgM3�v(Mg1���hͣ��qfn�3� �׌N��贘��˻�Rg�_��L�����xJ�x~ם!T�����hzϛ��s�b���w�p5��x��Wg��f�rߗ���eX�x��}��G�L4�?�5�e�G�;�%��xK���A���X&��xf���$�5�O�uJ��7gm�
Q�ũ(�fyn\ڽR�h���",�D�x�hV�?إ�h�r�NiX�;v;�FKWۄܮʒs�}�h�� �[vjxd�h��6��XW�+�w�am f|�ܓo�]D��R���X�G��x���.f�Yx����xI5ˤ`Σ�B+���`g�e���eHu/.��~���@hXG%�f̟���GJ���x�˵�g���S7�Jxf����h����d�}�[xV��F�5�fŀf��1��x���D5�fo��T�Eg��� )�F�x�O����|��nآf��u
��8g�v)yK�J���Ֆ��$�xf���bV�~�lxo˥h֟o���!؇�hؤtiM2,�7�dg��@�����%�J�e�o�[	h��,.��
�����F$�I~f�0WI�>L!iEI��E����7�O�F5�fԜh"�#,�]1�4��I.�;Jg��f���`�X�f%�Kj�}Ke�k�O���axf�Ј/��BVM���K�$�tF���>g��6���fI����B\�߅'��L��f�ʋ]�R�'n�fc���0xl��x�Tg��&�W`s�&շ����	�4f��x��f��M."	��( �j�bY٧0�Y��,+f�ʏO֗�h��]��@w��F�W��e�h}�O?��i���b�PWz�Qa-K�lfn�3�˥�ئQ�˥Z�WJ�ћ��؉�h�M�[��n��ex�˴��\I�w��e�e��N��Rmi��$;�ik���qt����fX)�+p���?���>���fN~�3��Yg��|Ƅ��I� ˭mK�r��F%��f��7�ؗ�-��UI�Dd(�
fh�x��e���bQ򛆸Y�f)˩�����E�f�fx=����F�G�ˣGe���O��n3xf�㿗8�h1j�pX�W��ͱs�n��D˙eڍ��U���ExY����\��k��0�f�.|���XY�~3�˯�8�kը����xf��v�A�4���;N�˟7���h��,r��%f��~���xp�}X�ø�i�3��,�e��Qi���)��m��҃��u��x^�nf�nf�ߍrax��}I���k�˅/Txf��R�yx�<6��F�A�?��;z�Q'o�f���^�њ ��Fn=��N�;�"X�i�Og�#8L������;z�ˡX٣�a��*��h�d��6�:g��=��ʀ�vS���xL��nfX/b���"��ˢ?((�h����h�L1�����X�ʤX�G\��(��0�f��������,4�	e�9�A,73ނ�"f���9ʸ�Wx�o˞ϖ(�f��C�ׅ�h�n��uS0h�����˩�6.GZX�eOf����T�6*@�D� �E���N�aiWȯf��?�	�hĂ-9��;iF�K�����gxf��V{�x��+<r��橤�Փ��Rxf��g��?Z��Y���W8�qKg��+���f���6�0i�K��N����j+��\�htHM�7jƜ@����y�dP6[�x]j�`g�Hg���	hK�$��eى��.CSm^�"f��� I����\I�t����p}-=�'�f�jt�׶ui<�G�8˄ ԇ끣J�/�pf��M�;j&�fx�e������Jw��fn[3�{)7،Q��>c(d\g��RDSg�*���
��ޫ�we���p������pg�6I�:�S
 ����XL/���?�U��xf���L#�g�`�}�y�����/�Xǰxf�7I��Q��x˧^k���˅?T�f��X�/�f֤f�Ec˫���oնȒ�� yf�Jx����-�9g�˧�ʭI���xf}�h�ߊgNj����Fg��	��W:]����&�f���3�������˥��(��s�����e�����hlR��˰I�[����%K)�Zg�Ix0��-�G��B����XV�;�f��I)�@�R�tf4ː���(V���n�h�I8m��I���x���\/��O�d��h����#���~����R3��I#w(Mg��f�\x59�X�~x�c˪�� +lK{���5of�
�F*Hx���Z����c�@�֡x��lf��Gs�W�2�f4�D�����>�xf����<��жK�����(��՞k��n�f�W~Kb��5�Mx����m�qsf� a��%f���A;���GK˅t~qF4He.f��h�1�o���_�1P��66q���׷�h��0�C\)��T�x
�� ՅK��U�xf��.ּ4��?�s��d��<��I$�Ztf�����!�&q����6X��4 "��o?�f���ƌ�f1�-qq˥N�φ�����f ��S�w�f�v�o[�{?X��eוJح.f�[~�`��)8��D�����e5�4g� fsDQi ���H���e˥:�˃���f��_�/�*����˯:n�o�:�iKFgM��2����w����]t��=�Ϳ>��e��(q�޹���CJ�RF���f��zr%d���3D��~���eH"�}���h�_g��͘�o���ǀj�!���}wIgn�3� �0��{���J��&��x��IgX/b����
�����C鶐Ux�˗Jgn�3�˥�֓{���%�2�x%^x��Ign�3� �H��{����Gז�jx͗IgWK�����$�����	D.�JxУ9�fpp[�Kx�֔M�����2�x%^x��IgnT3�{)���{���ZC鶐ex͗GgWK���ݷ$�����	��ȵexc�9�fT%u։
v�֧R����{mfpcx��Fgn�3� �@��{�����G��L�͗xfW�3��)�$�����	��ȵmxУ9�fpp[�Kx�֔M����{mfpcx��FgnT3�{)���{���ZC鶐mx͗GgWK�����$�����	��ȵmxc�9IgT?k���QاR�����2�x%^x��IgnT3�{)���{��ɚIז�bx͗IgW�P����W���tK|C�F���Ggn�3� �ר{��]׀�5��V	gޝesai���+�{�T��	�͡�S2�����h����ʞ��K�#�I���;�� 8)f�s�9jV�1x��ˁ�g���bB�n�xfu0:���h
E�ؗ��O*D�B����hpcxf��H\�˟Ɛ�WP��U��������hM��2���w����;tg�)����\�e�ag7��[h�Y����K^��F�&0fz�O?�8g��3=Nˢ��K�ޭe'1�e��8>4�ҷL���dw�`-#���en�3� �רP��v2����{T��^g�����kͿe-�����Bx0r����mf�E�eΐ��
���؃S��*0xhd��f�Ƹe��V�9W�"� ��ͮ+'��}�ʡf�x��!h�z�K�`W�����B�pf�K�h��x3��~;���KF�K���p�xf�dQg ��x�v�ˀK�ڸk�%�i�Qg���XZgU�)�_�;уSG���xgd��h��Ufΐ����,:��|Ie-��f�����h�n_�SL���H.�* �$�f㖁��J�?��c˅�v��O�|Ƙ�9g��h
Ea��;n���P5�G\�;Jg�.�f�fH��)�F�I�˱d�[�}yʥ�'lZg�����qh�˸�ˁ]���1[FxK��]g�ŸP!�V�#���˟�wf[��׿�h��ϤτfV�(���h���{
��Kxf�[ �~�k�VI�e�LcS�x��˥?1f�1���ȭ	�L.��~*n���x�|fᵤ1+����\˵Ԇ��e`j�%�ޥf|�1/�]X�-��Pː����q�����f�hX�+��G�J�tK|}�M8��Gg|H���Hx�f�g����	�4f�nx�5�f۵���2���@b˥3O�e��-����h��!6�稕��4� I�bX�-�F�E�h��b[�6}:�6�˰V�*�wʳ���f��Ԙi�t�*�T���8D.�Zx�4xf�C���v�:z^5˨f�<�&Y�h��h��0���
;ˆ�ˁ
�Z��F��0hf�ʸk`��w��b�=�Wۼ֮���fx�[�#�;]��突ʥt�sxbH)�e�z�h؄agJ��V�bg=�p#'(�e8�kr��fn�3� �צT�˭�R�Dtn�y�ʙe�"���������:&��(o�nGw��|f����ʇ)�����R���9�6�lxf�����8m�˖��˧]{x��˅?T�e��bG�h��wT�W_�(cg��,eqp�e�ق�z�pqx�i˳/�v�f������(fܯH9�_XA���P��4�Vcxx�Txf��h���!���~���}@�����X8g��xf����ig@R�	�Q*w�(@˜���bg���[�i�>t:��ax�Lg��H����h�����|�:�{K9˟�гu��`af�xxf�00���H4q�\���3���G%��vfWAϓQ���$������4f��xc�9fT%u։
v�֧R����<v�:׫)�r��xfY hZ�{)�D}����&
��ȵexΨ9IgX�+p�������&
��ȵmxc�9IgY�}�����6|����PjP"�z�}wIgn�3�˥�ֵ{������Jx���FgXx�q��k�����/D.�Jxc�9�fY���,���6|����NdP!,�}w�fnX3�{)���{���J��&��x��IgX�+p��������	��ȵexc�9IgYō}��aD�6|����PjP"�B�}wIgn�3�˥�ֵ{������Jx���GgX�+p��������	�4f��xc�9{fY��Y�{)��6|����NdP!,k�}w�fnX3�{)���{���J��&��x��IgX�+p��������	��ȵmxc�9�fYō}��a,�6|����PjP!���ڌIgD|�A̺F<�G�p���&
��ȵux�7Ig�D{hݲ;8Hc�f9�}�������xf��j�$ۏ̇�+ˢ�f��q�N���Wg��K�9�U{�xDQ�aUof��V���%f�	i����,����t��IJ��6g,��h��������<��~�SKI�t�hpQ%f|*�E� �2��S����t�:׫)����xf�Gۘ�Df��ڬA�Lݦp�h���(��!f�1V_���V��ˁ�t�bE���i^xfn[3�{)7ؿN�ˤ����f��x��׈euW��7jƜ��b�auwqI�G�6g���h�^l�O1 d��x���G~l|�e�L_�\g��u�Yf.z-qK˲4�x�:���EF�xfs�ev�c������K��ֹI%��f��h��Eڹ+��˘��HO�˖W?��h��x�+R7Ix1��]���h�"�n���h�����˘��]e5�������B7F�xf�o�
a���pix�D�]��cP�O_�e'��f ����I7q�G�ˁ��P�V�[xgj�f�6�`����#�����e�	���F��f�+��fx�n�ޖ�SE�ʞfN~g4��Yg�́޻-R�v<�1��Y��XW�q�É?�Xg��f��ݏ*���V:(�,�P��h�����1��dm��V��Zx7�f��h�d�2�fٍ��e��زP���}xK���f����>�f�^b4���J�BgX������h�/ޭ�|XY�~{���]~ �/�˥�'l�f�gg�s-�bR��R�d�%��>�^GgĤ}eU�1fmˬ�q��lK���f���S����s���P����m\
��ʙe`��p�!��������5+�и�=t*�Fgn�3� �רP���ۗ(V�R�G0f��Fn��[��b-��������Vǌxf��.6%�O�?gu�ʟa�pgƓ��1�Sg~��e�.�e�)=g��`u�oxa�w_g,}!f|��rB��^���3��8d8��hƓ|0a�hn�3�˥�֫T���6�ofV~&��ǡfԨ�����Ǖ�˟���~f�↳��ft<J���S�Dx1��X:��7�̩&��ef��g��6*��o���F��Ƹ[�F;I̲f���.���6��p�]W%5�l���̾��f����b��<<�zLa�k�%�i� f�7x<�S�����=7`�zs$g���{f^�h0����J���wu�Ϙ�����4f��h���I6����ǀj�!�(�}wIgn�3�˥���{���J��&V���FgXx�q��k��
���Ƀ�G��L'��˗�fn�3�˥�֓{���%�2�x%^x��Ign�3�˥���{���]C鶀bx͗FgW�9��P�$���Ƌ�4f��xУ9{fpp[�{w�֔M����<v�:׫)���xfnT3�{)���{��ɚIז�Jx͗IgW�P���$�����	D.�Jxc�9LgT%u։
nRاR����<v�:׫)���xfn�3� �@��{���ZC鶐ex͗GgW�3��Y�$�����	��ȵmxУ9Fgpp[�Kx�֔M����{mfpcx��Ggn�3�˥���{��ɚIז�bx͗IgW�����$���Ƌ�4f��xc�9�fTE����֧R�����2�x%^x��Ign�3� �H��{���ZC鶐mx͗GgW�P��1�W���tK|��z���Fgn[3�{)7،Q�˵\��fձ�����xf��ϣ�d�e�b�H�˘f��)p��Zs�$=g��h�����-��aX��P �%K1�h��:��l$�Ɨ9�{��Eŭ�)���xf�_	g����'۪|��D����e�vKAI;g��/��g*y��S��"{��Ǳ?LxfM��b��o�V���˵��kD/���.�Ggn�3� �׌{�� h������oV��<g}�M. z�a�x�b��
�/��FLĚe߱94؞�?6�,�p˴E׷�LK�m+خ�e팘b���
��pg-ˢWn��6��?�׷xf��"��Χ��Җ�˥�2x8��ff.!f��he��{ʊ�G���Z���k�{�ş�hs��0�\�f(��1U�7i�d�f��i�Ӗe�����ڈˌP��ń��S�x��e��L. �e�ox�b˄�`.�O��g��h�☧�>�	���i�2��I8x(Mg�:�f��h���gKY��˱n֕Ic���h�}�h��+ �e�uy���CJ�(�f���p_,f��4f�0x��Aȳ��Tӡӈ��wxd�.<g̤�h��e�X�Dg�F���H��h�8��xfߜF�;j&��xDQ�OL����څ*)=g�£��~vDfx���R��%I1xq�=f�HN�����eQ�E!����h�8p�xf��F�7�fhx�
f�ʘ�٫���k;���Bg� c�Q��'A�{d1��&��xK�l��fD|�A��M(�I�m��W&��t�oJ���vf`��r�k�֜�����v������I�h���e-�|f�"�����&
��ȵux��5Ig{\��C/i�$$���cZ��C�����U�fۯ��˘l���bI˫�{ZI#�w?gp�%f������b���ő�x�=K�����j�Ggn�3� �רP�ˮֵeh�m͡�L�Vg^�O���ܯ�Wi��27�F�6��hOIg�����f�bxC�b^�ۘ���GG=*3f���2ː�����)�Ub���K�ˁ;�TQgϧ/���[+��K"˫����J(����h�+��_xf�����-v�:׫Rx#��xf��k C��U����ʟ���u�R�Hɽˁfԏ��(�����ʅG��v�1X*�H>g���[�/X��D��y&�nF�א3f&�%f�%��gF9����@3|����3,�{%f��F�9ʘ��x�D˳zץ�껖��,�h����i˞�pYō�Y&��(o؇v��|f���ev�?
��^��*�O-f��kf���h�/�����V������w��x�̹xf���*ڰ�Ux u�S!g������h{Ȁ�V�,f5����HV�������f{� ��>h»'��Iu�qx��vf�h�� �6�f�J�p�����m�FL�f�Ÿ���6VŐ>�d�]S�8=�xa� �ety�xr�xcg��&�ˮ��X�LKk)�֐�h��h��8�<�;j��R��AI+���T�h��G����
g�f����z�!��*�����hٜ�h���&c f����	��ȵEx�7Fg朥e����cpgQ˩fX݇eF����h�0����S�\����Ӵn��{I9���f��a�U�f�fY���E�֋v�'�f�ˢf�����YX\I��0�R��&w�n|ʡfƱ���mH)��*I˘��X;�ˁةEg깺��%�e�̗#�ˀg<E�/�ʡ;�Tf�<F�E<R��x�Y�S���/�����mf�ã�-�F��Nx�f˱<\��F���&��xf�ťG�h�J�p��B���є�����f�1��+s��xA��9V�*o��3~��3�hn�3�˥׿N��@d���&C����h��(A����ҦG��˅	ן�h4/i�Lfy�h����bI��˩c�������))�f���gv�!������|�8�k�{���bxf���9ʘ�]x��˦����w�x�n˝e�difȐ����_��t����E��)�f�� �T�G^�o���S0����	t�\f����h�f�(Z˦1�� ռ��v�{xf�Ŏ�7�'�m����=<8SgF�捲fn�3�˥רU��	��h��E�م&f��L�9j��jx:Q�F�آ��d%@��f�Di����&���z���o-
��xʙe�~	i��!]��o��[�p}�/V�h�F�e��xNH��q�D�^��[�қ(�֐�h��׶u!8�Fn��Ou�-IBh�o��׉e�K�f���͟���Z���N���p�xfDt>��OM��o�˧��P�p�xdh!�h�=L��@�*(�����Mt�q��ʉea�D��3e��|=��O�=�����!v�Bg�ׅ�)z6[�xK��Eح�#�[���f��	f7�}YY�o��:	u�϶q�3�]{�fȁYf��+-[���˃&��x��f�_��IgЏ�/�t����˪Kb�"�v+-Zg�7�`���ؑKx���v2��I�e�e��yf��ۚ%%�؀A1���A���O���3G��f�����9W��"�Iނ��
��I���h��vvLx���q8�;��T�v[�?6ؔ�h�HH����˟����]F�v��e|f}�ev���J���K#aH>$���_g��ۤ)q��r[�z��@�}����O	^2Vg�GH�ˀ��x^5ːŗ�89�x�W@�f��UL�dT����pϑ���٭xI�$f��i���6�:g1�\s��FIxb�f&U�f^����e�uy.��]c�����)�f�ʰ������!��v���cȪ�#�xf��#-{L�[���J"���ȱ6�lxf�uX;���-������h��) ��T��:g�>���rx#��Z��tK|���q&Fg�F� �f��xEQ��Q��2&!���bxf��x����L5�eA�̸�9�6��f�o9���e���M(��B>sR���x=�xftn\����fBE�e˰�9ByF����h��E1�2��.�ƺ4�y�տoVv�Z��p�h��i_�{I������:Z�ʯ�����U�xfʻ�����F����&
��ȵux��5~f���b[�S��-�� �=�\���W$�7g���e��N�F����M��o���Ҩ�{xf������a_;�O����8a-+��L}fn�3�˥�֦N��p&��V��h�E��xf��O?�8iH��7�ʂ< y�y�:yf�6�\�
+��T�����شx~��f��e�םNgU�� ˬ�z�!��������h��u
Gb�h�j].K�� �����u�xf���`v���f���ؠ��d%�h��$f֛K� )�.tx:Q�M��[6]��o��f��3�j���[5�Ukإdzc;U-�\ag���)hV���Ju��I�F2�J�%f�ߘ�ʞ��}^#�v>�e��=ʧ%G,hf�'I�A��F5�m��_��}f��,e�p�h���-"	��Jgx�i�H�������I�ѿ�f�nb�~�ALIAG�Jw�x�Vt�f|�h����u%�g����˰��Ci�ػ���h��_7tOg�{�
ˤt�nF��f0�%f��[�%X1�|���Ia�d�hf��_�e��=���������z]}��P�ː��Dg�`LP��A�����4�5�>')�xf{�����89˖V��tK|*Ԉ��'Fg��&R��E���L��d���K�ˡ;�T�f^g:�h8*f��}о�{�d�e`zy���hn�3� �׫Q���eM�n%�l.�;g��dh�v�f�)y[�Q���ՙK�8@�fד4�G�V���	A�7��.I2�e�f�,I��d&Fgx��V�Rg��uo׿�e���i���ЙiI��J�M�Xe�j`��f�Kii;�N��xf��9g��X��ˉ���f�����h�xʸ�4�AWمש�w���e�=��(hx��!�q�˅�0n�қ�gؙ�en�3� �׿P�˯Ii�����5��xf���_�O�bG��˪���kՁ�%_xf�Xnf��L�={��˭�ː�j*Fgn�3� ��֦P��OL{���˅/T[g�����8A�ʖ�4�����DFee��f{����!ڦ�F��H:X�eFi4i�kf��Kΐ_�)˪l��vXHuf����Q�f���
�˖/��A�U�e`zm2��f��Vڽ%f�m��P�{����M�51?g�Ϲh.����>g�˧�ٶ�e%�h��$f��2�kH��ܻH˯�~��[��l��=�h�����f��w/�=dx�eV~H&�ʡf���?8/yh��tFoxE(��f��f��cgD���(�f��|h;������:g�����xf�x#��a�]����(��\f�ǹe�2Q�G��f�˥f륕\M3�oyXg��h����n[:��c��]�����^
�9g������������8�dLgcGU��_Xg됎QB��֫3���Ds%rGF�c0f&;�f��Xɭ�x8��F���f�U7g����.Sg���ؔ��SbFfI�K��'j˫���Vf�eUf4�#�:�*�����4f��x�f��`���[i����/�@s��x�8�Xg.�if��K��1@g��F��\I�v��e�e���P��P��|�_�˲�S��:�3~�"�f�7���S2x1�˨��̟w���ʍeө��Jg�xPD�t��x�f8*f�if�� ��Q�h�A�Y�De������[xf�����,f�6I���e�q�hƓy�o �e�G�g�f���	˵O�HfjsW�՛�f��`�àeU�)����>0��U�x=�Ig�o��u��hh��;ˀf!i8��%�X��f�����)}͗hA�9�L̯������Ixf���b_�{������˳tKsG]�n%f(N�f��f*��P.�x-���&
��ȵux�4Ig��	h��{��;z�˴�%�LWY	f��h�/���ܘ���V���lͯDܻ���xf�/���52�	�S����t�:׫8�S��xf��x�NQS7��x�"�:׵�_�ʩh�~f��úǉJG��tZ��8D.�Zx�4xf|K�f���>�.��}��!�&VYL͝e�aYi��[��˄I�����X�x��xf�+I�h&r�MRU����t�:׫)�S��xf�y&�]^�Ffr�M!כ�?��>�2f��#��yI��Y���j�Ϙ��+�J�fn�3� �ר{��ր���V	g�e��Wˀ ,�f�a���6HB��xf��W��0i�B�����f3�|���,fy0�����h�.�~�U�f����Ċm�{������C�+��%ǥ��i6RmD��LЁD�����t_?�3Ǭ�~��X'�0\���f�;�����ǩ&��!L���Y���G���n���U�Ǽ����`�����恘hk��������y ��I���0���&�}g[������ǽ�F-�������D�fA�3����O+������3�k������?ۼ�ǐ�?���Œ��F+���L)������ ��ة��� ն��^E�e��dK+�)�N+��߾��3�k�������u:��AL���>3�k����&�D�fA3�bA���������Dk�fAc�J�w��^3�`p��=��Cսt��@{�1�kL)�����?ٖ�ǐ��F���5O���Β��!�����k�������<3�k����ܾD3�f�lXŌױ�>L+��ܾ��1�k�����F*�������Dc�fA�J����^{�J���^k�:{�HuA.�J���^�3�����lA�O3��I�p��C��r�~쒍��>3�k����޾��=�����3�k������i� ��_��+��8�+��+��¾��3�k�������՞~�^�A�bNb��&�9rœ�0ݚ^ŶnC�1�kN3���0}޸X������ШѺ�@�aA� ����H*�=�����3�k����%��W�$����ăzPս�F-�������됅�?[�ǐ՞?x��ǐ��L�B^�6lLsE��(?�F�_ `�����3���+�
���ݾ��mI��^�5	�:�UH]����@{�lA� ����F-�����������Ƒ�\=��m�����m����F*��������됍�H�+�S/U �+��M)������V���
�e_��39:��L��������ݾ��lŌ�=��F)�����@�mA� ����F�������������X�߃�as(�R<�;��Ѹ1�k��Ꝟä�:������@k�3�k��ǒ��?3�k����߾D�fC{�cA� ����H(�=����Ž��3�+�M+��޾��3�k����՞됅�?^�ǐ՞�V���+����e�r�Cjא����՞H+�cI3�(�5}޵N������ݾ��)�O+������3�k�����!�ƫx���⻦{�xR����n_k�3��������+��=��+�M����+���J n��^�3�����Jf��^{�5�������ݾ�@lŌ4�
�уnJ=�aA� ����F�������F.�������D�fAk�J���^�3�k��ǐ�JG��ː)g>D��ǐ��Fk����dK�+�|�����ݾ��)�K+��ܾ��3�k�������%��q�)�M ��+��¾��3�k�������՞?زǐ���#3�k����+�D{�fA�lL�b �)��������蝞��������蝞���p_��3=1~��
���F(�������D�f���F+���'m{���rJ�J��^k�cA� ����F��������k����)�Dk�fA�l�y���Ř�����Ns���Ꝟæ�bI3��]��F(l�5Huޠ
���F*�������Dc�f���F+���'�y��Z2?"�Ze���k����)�Dk�fAk�J���^�aA� ����F������W �=�m>3��˦ �cݲ^������h��+���k��ǥ�oM$��
��ä|�觪j@$GC�cA� ����H(�=�����3�k����� �ơ�X��F-����������#3�k����+���=��+����+�N�KzI���h���ך�'�����^���d>�ǐ��Fk����g�9+	���ݾ��)��+��¾��1�k��
����k���l�����(5v�YZH�i�F�<3�k����$�ŭ�ä�㣩+"�+�N+��߾��3�k�������OC��_�:4�N�.M����lLb�(�0d��F+���O+��[�������������ݾ@k�lA� ����H-�=��ˍ��~�}��#3�k����+���=��+�����+�N+��߾��3�k������՞�:N�V���s���՞H+�nC�3�k��ǼO3�ҙ�1�3���ᐦ��՞� 3�k��������=�����1�k'Av��F����Y����
��?ﷲǐ��?Z��ǐ�F���㏁i$i�W�]+�� ����^�3�����aI3�y���5�B������ݾ@c�cA� ����F(�����(�|�*�g�=��w���;� ����^�+��޾��1�k�㣩r�+��+��þ��3�k������N#\p_�ƻw��(h�v�3�v��'�Vԫ���l���(&�F.aW�h�|�\���J����^�1�����b_���@c�aA� ����H*�=��)��+�l�������=������ ���{wK��R���
lA� ����H��=�	���F*�������Dc�fA3�3�k��ǐ��Jk�`��<��_3�����TC͒��p�<�J�T��^�3�����bN���h0+����F+���	���F(����������ݾ���U��*��&���~�U!���+�K+��ܾ��1�k�����F,�������D3�fA�2G
b���6
����!x�3��kQ��
���ݾ�������+ء����1�k��������_��2��O3C������������$�D3�f� 3�k����(�D�fAk�J�\��^�askK��r(��+o���F+���L)��ç|ޒ��#3�k����þD{�f���F+���'-z�^}OJ��cA� ����H�c�[�����R����F(�������D�fA�JbʺhC�3�k����%���+���k��ǥ�J���+�
���F*�������Dc�f��eI+���'�z����M�r�����u[޼�r��'���E ��u������{�HuX��B���|���\��қ���C�1]�����R��\`@������4Q�B��+���H�PP�E���������a���v���7�Ɔ���՞��eñH����f�����L��������p:��������� �2^(��������D���������N�o���@����"3}����؂���ڨ����f�����g�������}'yU:�������{@������cʺh�����������OwR��j�ŧR[v���'^��ZH�@«
��$e��a�5�>>Q�\D�tk��e3��l�W���7&��]8(��yg�w�hD����J���k�D}6�l���7�lS���7�l_F��7�l�E~6����������Hn��!������^���F��������ej~������GT䑢d/i��j&����zp���b)�r�_ �!�Be������q�b�j���7���]���]��o���W���Q�_��Hƽ)�����*�+3
�3
����|)�*dǇ{��ܞ9HƼ)�����*�+;
�3
����)	#�6j�I��3�U������N������츽x��&�)��Ʝ��9P:7d)L���q�m�j���7��쐕���]��a��ǮN��Z4B������]N�����HƧ)�����*�+
�3
����r)V������oRU�%�ʪ��r��i������������~�k~�k���@b�jy���v(���I�p�-	,�+�U�������}(ަ�0�����7J�V��w(���L 
,n3c�R��1��2����z���ق'��,7��M����iR��H'��HƸ)�����*�+
�3
����s)R{0���h��HƼ)�����*�+;
�3
����)U���������Gc��[�靅MM��ǲ7J�V����	������춲��������g��V�k~�k���[o��� ���*Rߗ�����H'����v&�g�!�����������%�����Nˑ������앲�����������n�k~�k���B`�iΏ�T��������"ϣ��f�ur�����R�m����2y�������a��T�!�q���)�����I1V�*!�oAz����}��2�H��	��R���ǔ}o����S���ls�7J}���q�a�j���7�������]��b��Ǫ���3��G�l���Xú+-����'�����"���D�������;7�
0EKP5�&L����;����/���!������^���F������	����s ����Zi���w���h���Fh����X-��!N������dA[��F��������}�0z<�fϲ����Hƹ)����)�+
�3
����p)��rP ������uz�񙉆?���ܒ����S�������Q9�6��^����z���6���"F˦?z�����y��hD������l���6�p�B��$f����� ����Þ!O�����^S��F���������
4�=p�<�w���}$��S$���'�����[j��Ǘ.�&�Ǣ�ꉲ��7���'w�+9h'����?�`H֩XтԝRI��ռ��H�/�������HƼ)�����*�+;
�3
����)��R^�%��(������U��]�>WVL�"X�{��l!���Ih����?����ܓ���'����1Y��R�e�Ǔ:�P�'(����O�9>�&Y�����O�(����n��Ǡ�G;eiA����n�\C��)�H�Rr�6���p��F8w	?����!������^���F��������w,ϡ�Ɛ���g��Ǆ��	-�� 0$��)����������n�k~�k���B`��'��.���s��Hƾ)�����*�+
�3
����})�������(�G�/`>����Bݜ���������_������R���Ǟ�꧷!�V�����C=y(,��3l�>&v�����:���2ڏ��Q1_�&��S$��!&������[�77	����N��Ǎ��[)	'������EՒ2I�k��@h?�����k	��,�)Be���֫���������v�k~�k���_c��R������\�T�A|�쳬[���進�)���������s<6�T2K�T)r�_I�B2�T�v�Q5X�^�?_^"X�A; ������V%w�_�7�U<Z�Q26�O6F�@2V�@%w�A�J�W�7LJ)t��u�������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������               �R  `����a	�e���j U�    ]�]�l$�D$   EU�:})�q9D$��   j S�    [�[�\$�D$   CS�� _NYz$��`�ndC4��9-a��=! �\   `��)��+a��k9j P�    X�X�D$�D$   @P�ar��o`f�*��Ma�   `��a���   �   �    ��y!��Q9D$�g   j V�    ^�^�t$�D$   FV�9����$'�   ۱?���g6ziz��ǅ��&   j R�    Z�Z�T$�D$   BRåO���`j Q�    Y�Y�L$�D$   AQ�/O�I�1�Y�   ���%    �   ��M�&�u��������&j j���u,��� tj ��4��th�   j���u,j U�    ]�]�l$�D$   EUâ�Sj Q�    Y�Y�L$�D$   AQ�[_3N���   ;
WM�	�ٞ,��+�j V�    ^�^�t$�D$   FV���`f�ÿ�m�)a�T$(j P�    X�X�D$�D$   @P�X�)�`���1��1a���j Q�    Y�Y�L$�D$   AQÒc�brpQ	����1(�<   ��=`��un�J���at$$j S�    [�[�\$�D$   CS�%i��Cf�j W�    _�_�|$�D$   GWÄ�0E���,D$$�   ���   �   �k�����P`�Z!�R��ײa��   ����@x�i����& �p   )��P�   �   �    �$)���D$,�P�   ��A"(�?c�<�$j U�    ]�]�l$�D$   EU����������i&��Љ�y	D$(j U�    ]�]�l$�D$   EU�����
   ��N������@�@j V�    ^�^�t$�D$   FV�3,�� `f��<��a����&j S�    [�[�\$�D$   CS�ymK�n�C��X��pxj R�    Z�Z�T$�D$   BR�,�)����`��a�����|$$   ��   �
   �   ��e���	   <���9�E-PPR�   �	   �a#�ۤ4z�1`V_�    aZX�j S�    [�[�\$�D$   CS�	4`f���   f��a���D$(j S�    [�[�\$�D$   CSØ�9?�P`a�$)�����i&�   �   ����VPy)1��7����j P�    X�X�D$�D$   @P�fD�t��I$�j P�    X�X�D$�D$   @PÉ�)��1��)��=	t$$j U�    ]�]�l$�D$   EUË6����}�   `�������3a��   �[n�y��|$$   ��   j P�    X�X�D$�D$   @P�	��   ��s�^�L�����QP`�θ6A8a�$��D$(�   `�    a�   �P�   `�   b�i ��g�D����pYf��a�$�   �0x��a�9&����i&��Љ��D$$���   `�    a��   �  ����,j P�    X�X�D$�D$   @P�&�)�����|$$   �  j V�    ^�^�t$�D$   FV�eUv ��   (�Cgg[�w��U�ﱐ�   `��f��aP�   �	   � O�CD��j V�    ^�^�t$�D$   FV���D$(�   ���� c������bO��PR�   �   ����bMzަh@B	�jK!G1PR�    1`aZXZXP``f��SPR1ZXaf��a������i&�   �   �    �Љ����D$$�   �   ؑʋ)C{�ԪM�����   N6��d�P�   �?�#�w�nW��(��1�Y(�j P�    X�X�D$�D$   @P��^,)�u(���!��(j U�    ]�]�l$�D$   EU�5�Q3X�`�   �   ",����   �   ol"�Ѳ$�z��\�O�z�j Q�    Y�Y�L$�D$   AQ��CwAhU;�a�`)�i��a1��#1�� �|$(   ��   j V�    ^�^�t$�D$   FV�]$��G:�� P`�	   A��G�Ǒ?e�   �~XJ l݋jba�$�   `)�!!)�a�D$,���`�   �� [f��aP�   �   `a�j U�    ]�]�l$�D$   EUÂ`�tJB�t��   ��e#)�i���i&��Љ��.D$(���!`�   �   J�IiX���YT�)�m/a�j S�    [�[�\$�D$   CS�61C�^����&����& u
3���T�&��V��|$(   wP�D$,P���i&��D$(��ߊ���&��t:uLW2��u�^+�R�3�I��3�3۬2��͊�ֶf��f��s	f5APf��IT��u�3�3�Ou����ы���f��Z;�t^������]���^j V�    ^�^�t$�D$   FV�X�\(�����j S�    [�[�\$�D$   CS��0QI� )�A*��j P�    X�X�D$�D$   @Pô.T8=!��(j V�    ^�^�t$�D$   FV�#�e�U(�   ��.Jľ    `f���	��-a�j S�    [�[�\$�D$   CS�e�b��   �   	�e,f��   ���`���E a)�e%�}�$�j S�    [�[�\$�D$   CS�<��<�j Q�    Y�Y�L$�D$   AQ����� 	�Q�|$$   �  j S�    [�[�\$�D$   CS����   �   Nɍ玈$�6-y,�k���wD`�����Y�zaP�   *��KC�$``�	   ���I�3�+݉�5a��a�D$(j V�    ^�^�t$�D$   FVÂ5�ei� E���/P�   PR�    1`aZX�$��1/���i&j P�    X�X�D$�D$   @P�!�� $�D������j S�    [�[�\$�D$   CS����5���,D$$`��/f�r%a�D$�   ��h���BS��ƅ� ǅM�&    ǅ��&    j U�    ]�]�l$�D$   EU���4��4	1��j Q�    Y�Y�L$�D$   AQç�����   �   �.��\O`�բ�aj V�    ^�^�t$�D$   FV�}��� j R�    Z�Z�T$�D$   BR�@��`���f�a��}j W�    _�_�|$�D$   GW�jE��J�%'k�j S�    [�[�\$�D$   CS�����)��$�j R�    Z�Z�T$�D$   BR��_y�   ����Mv(��7-�7r�~`�   f��f���<a�j V�    ^�^�t$�D$   FV�؂�   ,cX1�,p�dM��)��|$$   ��   j R�    Z�Z�T$�D$   BR����";�)��`#��aP`a�$j S�    [�[�\$�D$   CS�%���.jw^��)���D$(j V�    ^�^�t$�D$   FV��!��   ���'	��!P�   tGt�~T�U�$j R�    Z�Z�T$�D$   BR��Y{�B�r��i������i&�   )�)�Љ��?���`���a��D�&�   `�
   h�:�x���Ra�PR�   �    1�   �    ZXPPR�   �    1PR`a1`aZXZX�j U�    ]�]�l$�D$   EU�����/�`P���"XP�   �)&���r��%~�_Yad�5    )�E�$�   1��!��Aj V�    ^�^�t$�D$   FV�������   	��d�%    ������&�   �`)�� ��a�`j V�    ^�^�t$�D$   FV���
��l�   ��EN�yg>�+�  j V�    ^�^�t$�D$   FV��������   (���\�<v9_A��`��;���q!a���    ]���&�xV4�� t����  ���,�  ��Y`����&����&P����&P���.��aj Q�    Y�Y�L$�D$   AQ��K����+�   �\�\�C�JG3v�$�   1������&j W�    _�_�|$�D$   GW�0�'IK��@`���_b���a���1��> �   ��I�)���   �������+���`f�Fo�   ��a`�����a�   ���"a�   `��3�83aǅE/   j Q�    Y�Y�L$�D$   AQ�k�7i�`�   ���   ���!a`Pf��Y�Y��a��&N�	   Y�
��V���   ��\$U�    ]��N�&���   ����&����&���   ]3��j P�    X�X�D$�D$   @P�Y\����0�Qj P�    X�X�D$�D$   @P�#�7�J���`j V�    ^�^�t$�D$   FV�0���|!��a!�   `��4f��a��f�&	�)�PR�   Q�!�|]�� W�2@,5:�11�   ��Ǎ�ͤ��]fk�<��ZXP`�   �	   ͭ���@�W�f��a�j Q�    Y�Y�L$�D$   AQò�Xկ��   ��NZ͓��rd�5    j S�    [�[�\$�D$   CS���   ���]��Η�u���� M�C od�%    j V�    ^�^�t$�D$   FV�7`�̋�a����&j U�    ]�]�l$�D$   EU��8����$��`j P�    X�X�D$�D$   @P��I�G��   $�q��ƅ�Oj R�    Z�Z�T$�D$   BR��`�   �cq.Og�	��e��9$a`�10�   ("-�ς���ej�wah�
��   PR`a1�	   ^j��i����ZX�$0T�=�   ��8����$j Q�    Y�Y�L$�D$   AQú�1L��   �   �����&j V�    ^�^�t$�D$   FV�/b���bɉ�
   ���{؈�������   j���F�.S�pgʁn7*�W�   )��\$U�    ]��p�&��q���$��y!��q������,ƅ� ǅM�&    ����&���   ]3��j R�    Z�Z�T$�D$   BRÐ��D���\�   �   ���m)��"�xV4j V�    ^�^�t$�D$   FV��~))�-,��d�    ��(��`��aa�   ��jk6��aY��	   V���VaM[�   ):kM��i  �Ⱥ} �3��y�3�	   �O�3�.	{�3�   &�������ٮV�� ���4�^X)��1��kO=3�A������!���e�   ��������~�~�w���(^�)�U��Ya��]�ùYaV#��+^��   �   �)   ��v�t�b�g�TtM̖�X����-'�S������M��� '�}y�@�:��>�u���$�O�@�f3�j\&R����@�i�j�d���d��\���`�C�M�C�M���{5�\~��I����P�z�l҂vz�dA����fDj�d�6��2FH�ZD�a�{��lL�i��!�E�gI����&*�����i�Ol�@�����(�i�@i6qˤP�ĕi�@��lpQ�r�����i�@�f��_=���g}�V�ۈ��.5]�O'�D���@�i�v@��O�0��Z��&�$v��Oo�@��OF���xf�@�4,l�-�-���=�'���o�!�of8o�{��c�)�Gw�,�g_����/Q���vj4�x a�)d��Gܟ�\�T�
�G���L�qQp!|Q�D>q��>r*Ez��GӁ��k�in����	���.f�K�p8:��)p,�)p@�)�v���Px��/,�M\�j�����X��h�*pU:pЃ�* m�)Z̑δfv��Y) ��*�h�b4��i�4RY��z"��z"��z"��z"��z"��z"��z"��z"��z"��z"��z"��z"��z"��z"��z"��z"��z"��z"��z"��z"��z"��z"��z"��z"��z"��z"��z"��z"��z"��z"��z"��z"��z"��z"��z"��z"��z"��z"��z"��z"��z"��z"��z"��z"��z"��z"��z"��z"��z"��z"��z"��z"��z"��z"��z"��z"��z"��z"��z"��z"��z"��z"��z"��z"��z"��z"��z"��z"��z"��z"��z"��z"��z"��z"��z"��z"��z"��z"��z"��z"��z"��z"��z�3�X?�K󦃿�(]k��8�O��Šw"��&dy�ڜG�v"���{ֽ(��d�t�vR�%�x�����������z"ɠ�#���[��(�|(���R��z͎��$Ca�?�a� �Ǵ�����z"i$�e��ʖ���z"��6S�W��[/��R��z-{隣�0���3/����y�N�z{"��c�3ZM?�%�)�=xџ�z"�_�X�'{$�%#� �JQ�q���z"�%���	Ȝ�Q?� x�3Q?�����'R�q�x��#��yH����8%6�zu�)44��̱��q�3eR?�F����s�����C6�ml��z"��z"��z"��z"% �q$�W<�#" �~����Wt��#;3�s�=�{&$��'+��'�������z"	�5�Ԗ'(Ö'�z"w�5��7�%���SqF���:���4r��Qwñ���8���qv"� �&�q��;"8��E�?���q"%��T�qv"� �&�q���(8��E�K(�H�#¿u"��� �'���g��#������I�K��8�O���!yP�z"����� �Ǵ�Ǵ�z"�����pέ��آ������z"�M8ى2z�#��R��z��{m��'�8�����z"DV�r�
EX%���e�R��z�I���(��7���!Ɩ�Ȩ�z��z"�f�$�F��2Fw��L���Út�v
�����z"	�5�ܖ'(Ö'�z"h�58��4��̱�'��q|��R&��z��BĚ��v�t�vȨ�zd�BmLB�s"��*c��P4���M���#9�u"������g��g��#���S�����l"�:yP�z"����� �Ǵ�Ǵ�z"������~s�'�ۈ��u�8��{�2Z�t`7�8Z_����p̱��'��zk�@����z"��z"Q�z"���'O:�(B�j�&k��K��e���S���zx�o�g�؜���#ƿu"��������g��#���T����\�x"��Bm���S��z���GA��y�����󦞠�z�#����~�z"�LU�Z�>�������N;��󦚠�6G��3�R?��:웂z"�z�#ÿu"����&�w��g��#���	�g��Z�j�#8�u"���
���_��g��#���R��.���jP���z"�%���8�O��v ?$��qz]=�7�'�@��'�^�q'�Q�̱�!'�M�������X�N��������#9�u"������g��g��#���S�������������#ǿu"������W��g��#���U�����a�̱ �^�q��A�̱E���qk�����z"	�5�4�'(Ö'�z"s�5����*^�q��A�̱?��S��zBw�t��nB���d��IE�#9�u"������g��g��#���S���?�-T"�Q�̱��#��z�3ZM?�!yRP�z"����� �Ǵ�Ǵ�z"����_�/��s�í��X�#ƿu"��������g��#���T�78�����3��̱!ykP�z"����� �Ǵ�Ǵ�z"������Q���8�O���%�q�#vƯ������z"	�5	�Ė'(Ö'�z"i�5͎�'��q3�z"��9��M���#ǿu"������W��g��#���U�4�2Q�z"�M_H�ix�I
K�_�&�.��G�X�#ƿu"��������g��#���T�G��xA��?�ܚ�%�̱����z9��̱��#��8)����o%�E��~�a%"ދ'�ׯ������z"	&4�̖'(Ö'�z"r�53�")8�O��r!yUP�z"����� �Ǵ�Ǵ�z"����I:��@x�z"R��F��7��4�}��R&��z��B��$�v�t�vͨ�zX�B���d��O�uC���#9�u"������g��g��#���S�$�����! ��q���z"�."T�����z"��9�Þ3ZM?�!ykP�z"����� �Ǵ�Ǵ�z"����'Y���z"����Ѓ �:yQP�z"����� �Ǵ�Ǵ�z"�����庤X�S;�����?�{�q�2P�̱�by�E@R���\vƙ�4�����z"	�5��'(Ö'�z"v�5�B`z�P����p�f�uC��b�3ZM?�!yQP�z"����� �Ǵ�Ǵ�z"���䁝��Ԡ?��-O��y�6�K���󦯒��_�8�O��r!yUP�z"����� �Ǵ�Ǵ�z"����' ��q��z"n9HU�6ZK��0&�r~yx��1��{9P�K���SƖ����T���y��7�TS�}��R&��z��Bߚ�v�t�vɨ�ze�B$I#m��Sy�N�zx"���c���M��S��z�$� �}��sŵ��:x�����b44�uñ�J
�����3`vñ��Ȩ�z��z" ;�č�@h�f�l\%��k�؟@:yUP�z"����� �Ǵ�Ǵ�z"����ǫ�H^��z�z"� �q���̱(�'�S���t�x�%�������C�ɚ�ivñ?U�/�7����#������������O؜��y�N������z"	�5�4�'(Ö'�z"s�5v)'��bȞ3ZM?�����z��wñ�J�z�z"�����v9/ U���:�gt$�����u���߄��
�q�{�z"��/B~��L�cy�yz"���d�;0�������z"	�5 �<�'(Ö'�z"t�5З��x�z"z��z��Hm�Hɧ�3^�!yTP�z"����� �Ǵ�Ǵ�z"������t��y6A>��M��N�������b�2P�̱��#9�u"������g��g��#���S�p��"3��o���#�7�,�k�����z"�-%C�{��(âd㦴R�S��z6�c�@BF�x4"�Q�̱!yQP�z"����� �Ǵ�Ǵ�z"�����M.�nXx.���ܼ�q�Y��@�y��������ea�����z"	�5�4�'(Ö'�z"s�52u��������z")����%8��>�q��z"��w!����GL�x���u�
��z"��Ǎ�!������C����#ƿu"��������g��#���T��bw���#L>#��&���ϟ�q|��R&��z��Bٚ,�v�t�vȨ�z_�B_�%��v�y|"��&M�s�SƖ��(ښ㉘��z"�F8��x4����#¿u"��� �'���g��#�����[�t�yH+�������z"	�5�4�'(Ö'�z"s�5zWF�����£	3��A��3��̱X�q�2P�̱��#ƿu"��������g��#���T���y�c�{_Ǝ���7�}� !yTP�z"����� �Ǵ�Ǵ�z"����� �Q�̱!yP�z"����� �Ǵ�Ǵ�z"����y���83��2��[������z"	�5�ܖ'(Ö'�z"h�5�����s1�y������z"	�5��'(Ö'�z"v�51ܵ�	(*7]BP�z"����}	\�Ɍ�8_o;�\���'�w"��b�,�c��S��z�F?%�C��y7X��P�z"��u���#��bL����k���Z���'9�Ŗ�"��z��؜��Ǵ���n;z����؜��Ǵ��X'��n���؜��'��q|��R&��z��Bߚ�v�t�v̨�ze�Bӣ�g6��ܼ�q|��R&��z��B��$�v�t�vͨ�zX�B�����g�m6�y������z"	&4�̖'(Ö'�z"r�5[Ż
�|�z"G�M��0b�\�_�3��̱E���qk_�;�Ҡ�E���z"�L�S��Nȫ���3J�9���J%&������uC������z"�W��[������z"	�5�ܖ'(Ö'�z"h�5��?L�q'���#��x޶]�i!�� ���&���'�/�������z"	�5��'(Ö'�z"v�5����I�2P�̱��#8�u"���
���_��g��#���R�(}yg�jqȠ�#��b�m���b*��Q)�'Tb
h�UT� �Q�̱!yQP�z"����� �Ǵ�Ǵ�z"����i'���1�ۢB��	ى���z"z z"��ٞ3ZM?�?�{�q'�:ykP�z"����� �Ǵ�Ǵ�z"����n�M3�y���ۛ���;��#ƿu"��������g��#���T�.��Yչ������(��C��}��R&��z��B��$�v�t�vʨ�zX�B��%�zx���7�z"��'�X�q���z"7	��%#8��Ǵ��X�S��z���������#����B�n��o�|8��R��/Q�eX�����g�¢�pƆ'��q|��R&��z��Bٚ,�v�t�vɨ�z_�B�gwF�n�q�P�M���#9�u"������g��g��#���S�eNw�ӀyR��z�%Z/�Z�u����0d��� �31�y�|?9��Ӕ������z"	�5�4�'(Ö' �z"s�5�[<YBq���q�{�z"�:��t�ʂ�\9x3����>����&��Z��P�#8�u"���
���_��g��#���R�{�5���2�3�R?���qR��z"�͒��)�n��/Þ9�&�=������̱,8��z"�q|���#8�u"���
���_��g��#���R�(Lu>�=u�VȝP�yH+�������z"	�5�ܖ'(Ö' �z"h�5��� ��^�q|��R&��z��B��$�v�t�vɨ�zX�B	m�_���q��z|��R&��z��BĚ��v�t�vϨ�zd�B��='���=�)��9��#8�u"���
���_��g��#���R�RB�������-�,��d�?<}�q���}?�p�#��eE��"!��z�4t��e�����z"�5ʨ�z��㊚t��0�7�Z�t�v'H:yP�z"����� �Ǵ�Ǵ�z"�����hK�;�4�>������z"	�5��'(Ö'�z"v�5 ��(ୠ��N.�"h��64�vñ�I䞂��@�س��)�u�����K�^V�����O:yUP�z"����� �Ǵ�Ǵ�z"����b�µS��zW�[��A�#<�k CG��z"�'����z"z0�!ykP�z"����� �Ǵ�Ǵ�z"����7���|�z"zx"������z"���#�����3���d�LV��:s��R&��z��Bٚ,�v�t�vͨ�z_�B��!��ع���z"��iX�Z��#s����z"z|"���5��zu?���q"%��T�H"쳇z�3|�̱���q'E�¤�Qwñ���8�"쳇z�3|�̱v��q'E����z"!���b��kxi�k�?!yP�z"����� �Ǵ�Ǵ�z"����e�I��#���<#���ë�^��47��M���}�z"�qp�����ۜ�(����z"zz"����P)��}�z"��z"�WO�'�c�I�#Ŀu"��������g��#���V��m%��z"(n3��#ǿu"������W��g��#���U�;�'D��q�3��̱!yP�z"����� �Ǵ�Ǵ�z"����ץ�;����S+��zj� g�O(�ǭw,��w�*Y v������z"	&4�̖'(Ö'�z"r�5}������!y�|�z"�,]s��M��SȖ9�f��� ��#Ŀu"��������g��#���V��^�3�y?�!yUP�z"����� �Ǵ�Ǵ�z"����Es�:��̱:�u���S��W�ǉ2z|"������'!yP�z"����� �Ǵ�Ǵ�z"����A<��l�U�����(�#�����z"	�5�ܖ'(Ö' �z"h�5,�0�:y���P�q���rñ�P�q3�Urñ�ETɆ��y�q�~�z"�#��X�R)��R!��z7�� ����(G��J����T�z"��z"��+�?���l���V��)�'#���:�p̱(@�������z"	�5	�Ė'(Ö' �z"i�5s�8
D�U!��z|��R&��z��BĚ��v�t�vΨ�zd�B`7k��"�"�wñ�]4\z"�'�ǯ�����y�����M����n��z|��R&��z��BĚ��v�t�v��zd�B�����q �F� ���C�ʠ!���ڟ�� �{"���#ƿu"��������g��#���T��\��z"mk���1����ǵ� '\y�q.�&�����z"�!ykP�z"����� �Ǵ�Ǵ�z"��������1��M���z"�%#��,
�q��z"��X��Q�sj�5p<��!�̱!yP�z"����� �Ǵ�Ǵ�z"����X�0]�D��wS��zi�V%@Ʉɬ��_y z"���ĩ�y"�����z"	�5�Ԗ'(Ö'�z"w�5>�Y!g�]s��R&��z��Bߚ�v�t�vͨ�ze�B��d7���߁��z"�.
	D6-��a�R��z:��A"��d��ĳ�q ɵ5%z�#��؜���^�q��M�̱�S��z��06�?{�R�^�vƟ�u"�!yQP�z"����� �Ǵ�Ǵ�z"����ՠ`ڂ���)���xz�Xq��z"�"���P&�����'�����R�3����P�#¿u"��� �'���g��#�����J�A�J�
x"�����Cs����v5�z"� <p�qx�������^oR��z-�,G�{�Μ8���$��zx�Jʔ�����z"	�5�Ԗ'(Ö'�z"w�5љ^�6���uG��S��z��5�]J���Ԅbw0��7��#ǿu"������W��g��#���U��O��!yRP�z"����� �Ǵ�Ǵ�z"������t�)���3Wq�����z"	�5��'(Ö'�z"v�5��xt3�z"���&��z���T9覓�m(����z"�����z"	�5�Ԗ'(Ö' �z"w�5�S�	�y�(������z"	�5�ܖ'(Ö'�z"h�5b�����`�z"�!yUP�z"����� �Ǵ�Ǵ�z"�����5�U���i�IR%�=�%`������z"	&4�̖'(Ö'�z"r�5����^y�#��S��z�Uy��F�*�^/��0�5��������z"	�5 �<�'(Ö'�z"t�5o&K�Sɠw"��wm�z
���\o����z"Xw�#��z9���̱;!�u�$���x!��آ�t�Q����̱�h䳖�q��z����̱��^�q�̠�#���ȃ�-X�e�n��96%]>�:yRP�z"����� �Ǵ�Ǵ�z"����R��JFx����2���̱&�7��z3�z"�%��I�S9��z�3�̱:s��R&��z��Bٚ,�v�t�vʨ�z_�B�b!ڜ�Bs��R&��z��BÚ<�v�t�v̨�za�B��o��w!�?\�q�2��̱�5�!yUP�z"����� �Ǵ�Ǵ�z"�����MC���"��z��:yUP�z"����� �Ǵ�Ǵ�z"����T8' ��J��(G��J�����z"P��y�C���%����󞣛�Ȇ'��q��z"�lJ����;�w̡�_�t"���y$���3�ʆ�d�q|��R&��z��Bߚ�v�t�vͨ�ze�Bm=,,i-|@��9�
�/զ�uo1�@k����c"�:yRP�z"����� �Ǵ�Ǵ�z"�������~���I�#ƿu"��������g��#���T��VU�v"��z|��R&��z��B��$�v�t�v��zX�B��i*v��]�q�3��̱!yTP�z"����� �Ǵ�Ǵ�z"����^��1Q���X��XrM�(�' ?X�q|�!yTP�z"����� �Ǵ�Ǵ�z"����?���:y���̱����q�}����
�(�㲖���z;�՜̱��J�q��`Q��
s����
�q|�!yP�z"����� �Ǵ�Ǵ�z"����X�q^2id��zñ�P�q14l�̱�P�q9�5�̱ �\�q'E:yUP�z"����� �Ǵ�Ǵ�z"���䍐��wTy������S��z���z"�o���qx�O��U�̱Wq"���p��z|��R&��z��BÚ<�v�t�vè�za�B�%j��@S�������U!��zN��ﷇz|��R&��z��Bߚ�v�t�v̨�ze�B�?�k�? �q9��|ñ?L��q"z�#������z"B��+���hz"�!yUP�z"����� �Ǵ�Ǵ�z"����|����k>��������{"����G���9R��z|��R&��z��BĚ��v�t�vʨ�zd�B ��I�"��̱��{�q�2x?��z"�!yP�z"����� �Ǵ�Ǵ�z"���䗡q"��qTxQԞ��q��`"�:yTP�z"����� �Ǵ�Ǵ�z"�����*��(c�R���#��1)��_2&��5�ވ؟M�?P�q(������z"���yH������z"	�5�ܖ'(Ö'�z"h�5U8 ?p�q 8%����}��R&��z��BÚ<�v�t�v��za�BpYyFh�ƃz"�����z"	�5 �<�'(Ö'�z"t�5g�@Q&�Q�yFj��uñwz|��R&��z��Bߚ�v�t�vʨ�ze�BZ߱E��y�z"4cn����Nm��S8r��U9�#¿u"��� �'���g��#�������>����2�A�̱�(������z"	�5�4�'(Ö'�z"s�5[��آR�E�$��z��M�̱5�J;��!yQP�z"����� �Ǵ�Ǵ�z"���������z"�F�Y��(VF
�Ȍ�������z"	�5�ܖ'(Ö' �z"h�5�V\�N�(עF}�y7X^�����z"n�>~��lܖ�j�M�U�#��9��#ÿu"����&�w��g��#���	�=�n�'��q��z"���N���ʆ�d�q��?�\�q�'!yUP�z"����� �Ǵ�Ǵ�z"����Fh-iN�s�?zVt�����z"	�5�ܖ'(Ö'�z"h�5�~����6#{"�����z4�̱�(������z"	�5 �<�'(Ö'�z"t�5��������̱qx"���#8�u"���
���_��g��#���R��#r!Vyx"������z"� �q���'T��qោ����z"�;��%`��u���������z"	�5�ܖ'(Ö'�z"h�5���X�|%���g�}��R&��z��Bٚ,�v�t�vϨ�z_�B!L��+�zy>A�򭷇z|��R&��z��Bߚ�v�t�vɨ�ze�B=,��n��z"�!yP�z"����� �Ǵ�Ǵ�z"����,9����	����� ��qcO��ͷ�z|��R&��z��Bݚ��v�t�vͨ�z{�B��m�P���Y8�>'�C&���̱�;%z*!�������=���!yQP�z"����� �Ǵ�Ǵ�z"������>j]�9�>��˨�z��z"��%�AuE�&�i=�8>�:yQP�z"����� �Ǵ�Ǵ�z"�����"/)�>8L�������Z�z"�����z"	�5 �<�'(Ö'�z"t�5���v�{��f�z"�-��������z"	�5	�Ė'(Ö'�z"i�5d����X+�%���w$5�@'��q�2 �̱X��-?{�q��	?��qҰ�z4�z"��!��G���*���uG���#ǿu"������W��g��#���U��<�=}![�9�\{��z"���
�'�q8Hv��ʆ�d�qR��$�ٓ�����z"	�5�Ԗ'(Ö'�z"w�5zWF�������z"� ?D��q�Bp+��%,��z"���B����y��Ѳ�������'L_�q._�����kt��9!yP�z"����� �Ǵ�Ǵ�z"�����H��~�z"ɖ	!��z�O)b�J'���!yP�z"����� �Ǵ�Ǵ�z"����Ɖ�K����-?;��#¿u"��� �'���g��#����y8? uΕ�诠r"��@`!��J��S��z������'��>��u�"����Oy"�hSӉ���z"�l�I�J���z"���N���>�
��SP�z"�u�~�7���%8 ��
s��R&��z��B��$�v�t�v��zX�Bj�K�#�����z"	�5�ܖ'(Ö' �z"h�5�� R '�\�q)��#ƿu"��������g��#���T���JCñU8d؜����q!���̱�p#��=X�{�����ف}럖z"���W�Y�>�6�pZ
�����R��z�W������z"��wm���|�� 8%8R� v������z"	�5�Ԗ'(Ö'�z"w�5���y�T�y�Jآ�@�}���#����
)#�G\s���&��z�$	��+4�yH;��P[0�@�����z"���zvFXp�9�S�#¿u"��� �'���g��#����Y"3�p̱�x"��!�p6:d�r"��z"��ߢ��8�!yQP�z"����� �Ǵ�Ǵ�z"�����jZ&"עJo`��U�̱Wq"���嶇z|��R&��z��Bߚ�v�t�vȨ�ze�Boᡍ#������aY�c��q|��R&��z��Bٚ,�v�t�vè�z_�B�|���X���z"�ک�0ry w"��9>�%�7�z!���#¿u"��� �'���g��#������b1��w��~j����z"�����z"	�5�Ԗ'(Ö'�z"w�5���!0�1K�������z9�ɛ̱�!��1������z"�����z"	�5��'(Ö'�z"v�5-�=�����#���#ƿu"��������g��#���T�<_���rñ�w"��w��n+�2��8��z"�!yP�z"����� �Ǵ�Ǵ�z"����5�:���̱B��ɉ�J@�������z"	�5�ܖ'(Ö'�z"h�5�F��ĩ�y"�����z"	�5	�Ė'(Ö'�z"i�5�e��J�>��-w�h泖���zx7�z��=��#9�u"������g��g��#���S���������}����}��R&��z��Bٚ,�v�t�vͨ�z_�B����Y�q�؞�v"�'ע��*�wz�{�z"���Vh����p�����'%��-�Vt�����z"	�5	�Ė'(Ö'�z"i�5�|*�X��!�x"����ּ�|t����P� �z"�!yTP�z"����� �Ǵ�Ǵ�z"�������2�q��:yP�z"����� �Ǵ�Ǵ�z"����I�_��*��z"����x/��6\�~;��!yUP�z"����� �Ǵ�Ǵ�z"����'�A�,�؜��p#��GV?�~$�O����O�y���#9�u"������g��g��#���S���>��X���������z"	&4�̖'(Ö'�z"r�5��<��V����8%,�(R��z��o��b�uG���#Ŀu"��������g��#���V�7�ԇ��N���u�1�yH��3�*!P,�$�Xq�'�Vt�����z"	�5�ܖ'(Ö'�z"h�5�h%�k(��n�z"�����z"	�5��'(Ö'�z"v�5M_?���O��#���GT�խ�WB&#��z|��R&��z��Bt�v�t�v��zb8B\�6EF�>#�xj䟄�����N\s��R&��z��BĚ��v�t�vΨ�zd�BJ� ^�Hg�n>A:yUP�z"����� �Ǵ�Ǵ�z"����#+s�����!yRP�z"����� �Ǵ�Ǵ�z"����!�X��<A����z|��R&��z��Bٚ,�v�t�vʨ�z_�B�ε�V���̱%��H#��z���>6Hz����C3�{"���#����s�+�G �.�"�Cs��R&��z��BĚ��v�t�vʨ�zd�B
�"���q�̱�;%z !��R��zv��W@G�y�OV���������م̱��^�q|��R&��z��BÚ<�v�t�vϨ�za�BbQ�s�����!yP�z"����� �Ǵ�Ǵ�z"����a�R�u�l>��q"��!w;}��ٍ�����d�z"�u��Sj��z|��R&��z��Bݚ��v�t�vè�z{�B#�����N�����H�)6�^k�7���P�����W�!������z"�u+=�؜�:s��R&��z��Bݚ��v�t�vè�z{�BI�3r(������z"�u�$���Jp�7G��J����e�z"�����z"	�5��'(Ö' �z"v�5��yf' $\�q4�uñ����q'�U�̱!yRP�z"����� �Ǵ�Ǵ�z"����b���7�����N?����yH���t"��?7�0qo��-_,�?��#ƿu"��������g��#���T�1��3��̱!yUP�z"����� �Ǵ�Ǵ�z"������#��a��}��ri7[t4h�p#���zވQ�O�����Hɠ�#��*
�ԩg�	i��*S+��zp�fpԾP)�}�2�bnT��\�qx�O�#ǿu"������W��g��#���U�����C64��ŗ̱���zx7E���1��#9�u"������g��g��#���S�.y=v���ڜ�e�̱��(�� �[�y�N�3��̱;7�dɠ�#����3�f�&��{Mԋ�؜N)l%��z"�����z"	�5 �<�'(Ö'�z"t�5�^t�$�R��z��6J�u��� �g�q�3��̱!yTP�z"����� �Ǵ�Ǵ�z"�����v�0�-_������p#������U����ǖ�&��zx醴������z"	&4�̖'(Ö'�z"r�5���У_t�$��#�����z"	&4�̖'(Ö'�z"r�5ǈF�����3!y��%tñ�s�q|��R&��z��Bt�v�t�vͨ�zb8B=ʜ4�Ok��b�c%�����_�qR���}��R&��z��Bt�v�t�v̨�zb8B,b�'�����#����7�����pxP�� *;!yx7���#8�u"���
���_��g��#���R��&^�?�����yH;�������z"	�5��'(Ö'�z"v�5�q1�vb���R?�!yQP�z"����� �Ǵ�Ǵ�z"�����Q�yFb"E:yUP�z"����� �Ǵ�Ǵ�z"���䯑������t������9�y����zr"������z"�JS���z���z"�o��q��U�̱Wq"���X��z|��R&��z��Bߚ�v�t�vè�ze�Bxus��"��@˘���z"�8�HW��������z"�����z"	�5�Ԗ'(Ö'�z"w�5�	e!� $�硏#����-���c�N����z|��R&��z��BĚ��v�t�vȨ�zd�BX��?W�q"z�#��������z"�F��(�1�:����z"���C<��#���#Ŀu"��������g��#���V�@c�2݄8��z"����R��� �q|��R&��z��Bt�v�t�vͨ�zb8Bpӧ��c����dt3����(�y'��S��z��=��>���t؟M:ykP�z"����� �Ǵ�Ǵ�z"����?8�q(������z"�u���yH������z"	�5�Ԗ'(Ö'�z"w�5B�'+���{�z"e&K_�u��2��s�&������c���'!yTP�z"����� �Ǵ�Ǵ�z"����ޡ�#������Θ��<Ͻҋ��3��̱��'��*!�u[1�Xq__��Vt�����O��#��z챇z"�����z"	�5�ܖ'(Ö'�z"h�5V�Z����؜�5s��R&��z��Bt�v�t�v̨�zb8B����l�IR%�����z"	�5�Ԗ'(Ö'�z"w�5yf�/�S���N\s��R&��z��BĚ��v�t�vͨ�zd�B��t_f�>�yx"����C��^o��������L����z"�j��� �U�̱��d�qQ�a؈S��z���� ��E��r�����ޢ�'!yRP�z"����� �Ǵ�Ǵ�z"���䍴c�l��T9�#8�u"���
���_��g��#���R��O��)�Da�Nk�����آ���oז����z|��R&��z��Bߚ�v�t�v̨�ze�Bƫ�5�ە�(���%��N#���z"�!yUP�z"����� �Ǵ�Ǵ�z"����6���3$HR%�����z"	�5	�Ė'(Ö'�z"i�5��}xSv��(V:yRP�z"����� �Ǵ�Ǵ�z"�����i'r�5٭؉���z"�� ��q3A��#ƿu"��������g��#���T�W��7ƻ(<m��̱�B1F{"�!yQP�z"����� �Ǵ�Ǵ�z"���������q鰇z"6Hz|��R&��z��B��$�v�t�vʨ�zX�B�E�R�y7V^_mP��Ԉz"��z"�	����՗������F�%���Q؟O:yP�z"����� �Ǵ�Ǵ�z"�������Y-b�����Iv5�z"�!yRP�z"����� �Ǵ�Ǵ�z"����>�n���q'���̱ ���q�����z"	�5 �<�'(Ö' �z"t�5 ����'�\�q3�:yTP�z"����� �Ǵ�Ǵ�z"����{�7��z3)y"�����q�3�z"�����z"	�5�ܖ'(Ö'�z"h�5f�,�-�(\,��z"�尥*S��rq��C$Q�z"�=/��C�
����� 0�q��ݘ̱(؜�:yP�z"����� �Ǵ�Ǵ�z"����&��/3@4�����K��C������z"	�5�ܖ'(Ö'�z"h�5'��؜�_���q�<�}��R&��z��Bݚ��v�t�vȨ�z{�B��~:7�?i7G��J����j�z"zc"3T�̱!ykP�z"����� �Ǵ�Ǵ�z"����8'�����y�z"F�^އ<��z�̉�y�B��P���yH���z"��R�b�%��#ÿu"����&�w��g��#���	�0�8�s��]�̱%)��������z"	�5 �<�'(Ö' �z"t�5P{9�;O���q|��R&��z��BÚ<�v�t�v��za�B��Պ̱!yP�z"����� �Ǵ�Ǵ�z"����1����>��<Z�#¿u"��� �'���g��#����1⚍7S��*��q�3�̱%"����ʨ�z��z")t��Y>m(�-�k���%8�m!yP�z"����� �Ǵ�Ǵ�z"����dЧ��Z�O:��o����z"�c�c{^��R��)c���֠'*���#ǿu"������W��g��#���U��>�@ ���z"����䜄z"���˕������z"	�5�ܖ'(Ö'�z"h�5[��1,�m��Fu���>��#ƿu"��������g��#���T�	N@��S�%*y��Uy	z"���2������}��R&��z��Bݚ��v�t�vè�z{�B�+��,�!:�?����#ÿu"����&�w��g��#���	��Le����zx"���?����#ÿu"����&�w��g��#���	���Q�̱���q9䅉̱:�����z"	�5�ܖ'(Ö'�z"h�5���z"��K��l�@�%�eɗ�X8ʓƠx"��ʍ�<�!y|��R&��z��Bt�v�t�v̨�zb8B0��� h�!y'�ݝ̱!yUP�z"����� �Ǵ�Ǵ�z"����>8�P�q|��R&��z��Bߚ�v�t�vè�ze�B�Э(S�y������z"	�5	�Ė'(Ö'�z"i�5��S�S��z���z"�o��q|��R&��z��B��$�v�t�v̨�zX�B�/�D�_�	hڗǾ��U�̱Wq"�����z|��R&��z��Bٚ,�v�t�vɨ�z_�Brt�����-����0�����z"�VSɚ]4|z"�!yUP�z"����� �Ǵ�Ǵ�z"����'����z"�id��c~�ڽ-�ז!"yx"������?��q"z�#��S~��z|��R&��z��Bߚ�v�t�vͨ�ze�B�%�/�i�ڏj�j��{"���#Ŀu"��������g��#���V�K(��tw��z"��0�1�����z"�-{1�@�������z"	�5�Ԗ'(Ö'�z"w�5k��l�K��p �q��`"�:ykP�z"����� �Ǵ�Ǵ�z"�����{���'���qx�kڜA�p#���C5�����gx��H6ȵ5%z�#���*׆�^�q|��R&��z��Bt�v�t�v��zb8B�+8d����#ǿu"������W��g��#���U�'+����B9D���U�k_��S���z|��R&��z��Bݚ��v�t�vͨ�z{�BS����b�Խ��uG?�*!S8�#¿u"��� �'���g��#����O�i��4��̱�(������z"	�5 �<�'(Ö'�z"t�5���(��uS�$��z|��R&��z��Bt�v�t�vʨ�zb8BRҽ1t��:yTP�z"����� �Ǵ�Ǵ�z"����@S���!�̱?]�qោ�����N\s��R&��z��Bݚ��v�t�vϨ�z{�B}ն�����z"�Pb��Bs��R&��z��BÚ<�v�t�v��za�BQ�F�����*�uG���#ƿu"��������g��#���T����p����d�qx�K*!X;%�Xq�����z"	�5	�Ė'(Ö'�z"i�5*�k�Vty�#�����z"ȣ�ۣ(��yяZ'��v��&�y�%���N���zuB���|ñqx"���#ÿu"����&�w��g��#���	��极z"��d}�pqR_;��!yRP�z"����� �Ǵ�Ǵ�z"����ŝڜ�arñ��#��A���>ǟ^����/x��N\s��R&��z��Bߚ�v�t�vͨ�ze�BJL�C^���Vy �#��S��z�M?�$
�Fh�ffyx"����3��^o �=�:��qñ��#8�u"���
���_��g��#���R��5^o��\�z"�����z"	�5�ܖ'(Ö'�z"h�5��6�B�찇z"(E5����ⷖ�&��z�
9��mP��P�z"ze�Q�#ÿu"����&�w��g��#���	�8�y��)������z"z	w"�� w�%� ���̱!yP�z"����� �Ǵ�Ǵ�z"�����ho �vn�K��X��
͠�#���D���|��=򦏘�^B�#ÿu"����&�w��g��#���	�,��e
�Y�k��z"�� "
#���ѿ7��z3�z"��'|�q�빕̱��#���xt"��S��zw�l�m�C��a��_��q��c�}��R&��z��Bߚ�v�t�vɨ�ze�BY@E9�Y�D:s��R&��z��BĚ��v�t�v��zd�B���U�̱Wq"���Ĩ�zx7m.�G������z"��z"���w�������y�B�������z"	�5�4�'(Ö'�z"s�5Ҟ)_7����7��#¿u"��� �'���g��#����Ɣ��>bA��z"�As'���k��1������[�����z!�	�̱�#ƿu"��������g��#���T���4�u[$������z"�YP,���/�����`)��tO0��}��R&��z��BĚ��v�t�vè�zd�B�����a_آ�'Ak�F~��1��y7V�1�`��z"�G�tJM�������@;T����y7�O�6ni���#ǿu"������W��g��#���U�b�>8����#����g��~=�Ѕ��M��	11��R��������y���#9�u"������g��g��#���S�0�;7_0uz�y�!��ZC+|�3*���#ǿu"������W��g��#���U�����3�������z"	�5�Ԗ'(Ö'�z"w�5+����q��q�̱�v"��z��Ivñ!yTP�z"����� �Ǵ�Ǵ�z"������'H�
�1;�(xΩ'��>������9%8�v������z"	�5�ܖ'(Ö'�z"h�5��'9����.!y�N�#�u���A�������z"	�5�ܖ'(Ö'�z"h�5�h����z��M�̱�	��z�3 �̱:�9j�ڵ�w"��+/~���ڷ}�q"���&�� �)	s��R&��z��B��$�v�t�vʨ�zX�Bgo��}�?$�q|�!ykP�z"����� �Ǵ�Ǵ�z"����͋��u���U��yH;�������z"	�5�ܖ'(Ö'�z"h�5����t�@�����z"�`�����|W� E?D�q'3�p̱����R!��z7�[1�آJ�e��U�̱Wq"�����z�덜̱�?X}�q����̱!yTP�z"����� �Ǵ�Ǵ�z"���䥲�U0�R����q�U!��z����̱�]4wz"���&��z�|��;6�0�z5�z"�!yP�z"����� �Ǵ�Ǵ�z"����Zd/����#��1������z"�����z"	�5�Ԗ'(Ö'�z"w�5L�=�"~ ���u�"�{�#�zx"��u�;����z"�!yP�z"����� �Ǵ�Ǵ�z"����=��F��!�̱^�
Y�q"��z9�m�̱�q|��R&��z��BÚ<�v�t�v��za�B��7�y'���#ÿu"����&�w��g��#���	�������_؟M:yP�z"����� �Ǵ�Ǵ�z"���������j��q(�����z"�����z"	�5�ܖ'(Ö'�z"h�5�^4�%S��z��3 ���yH������z"	&4�̖'(Ö'�z"r�5�8�7�/�|�kQ���}��R&��z��Bݚ��v�t�v̨�z{�B�4Pʎ������z�x�z",C'��,ײ	5n�!�S��z���5����J4���/%���#¿u"��� �'���g��#�����)PS�����z"�8\���� ؈�#ÿu"����&�w��g��#���	�6h�,�0����z"�4�ÕEXq�����z"	�5	�Ė'(Ö'�z"i�54�D*�z�z"!�)��Z6�W�lF��ه&�y�=R��z�Q��c�	Xǖ(������z"	�5	�Ė'(Ö'�z"i�5�.X��$��z|��R&��z��Bt�v�t�vΨ�zb8B��v�w޽���'Tz�qោ؜�>`��{��d�B�k�������z"��>.� AC��Y�u������#ǿu"������W��g��#���U����z�y7����uG��{�;���a"���̱ '���q��!yQP�z"����� �Ǵ�Ǵ�z"������D��z�j��' y�q���̱��}��R&��z��Bߚ�v�t�vʨ�ze�B'e%��Vt�����z"	&4�̖'(Ö'�z"r�5��%?�Р�#���JG⾶iJ�2'�4�{����̱��6|"�!yTP�z"����� �Ǵ�Ǵ�z"����Ze�оL^�O��O:yP�z"����� �Ǵ�Ǵ�z"����(��t�6��z"�C�#ƿu"��������g��#���T�q���:�;��?�X�qx���#¿u"��� �'���g��#�����9��kw]o�}��R&��z��Bݚ��v�t�vɨ�z{�B��xӭ�7�]2
魋x?$��~�#��z|��R&��z��Bٚ,�v�t�vʨ�z_�B���tB�z�z"x��l^��W�7(%�� ������#ÿu"����&�w��g��#���	�D�Z[I�$ܮ�lO��_��z|��R&��z��Bݚ��v�t�vɨ�z{�B[�k��l�Cs��R&��z��Bݚ��v�t�vɨ�z{�B]8�i%��z"��O=�轟K&m�)�����z"�����z"	�5 �<�'(Ö'�z"t�5E�����4�%�̱��^�q|��R&��z��BĚ��v�t�vͨ�zd�B=.��.�*jG �!yTP�z"����� �Ǵ�Ǵ�z"�����PG��ӈ'%?_'{�q3�?� �qmd�z"z�#���#¿u"��� �'���g��#�����m7]g���v����z"�:s��R&��z��B��$�v�t�vȨ�zX�B��O?�q��Bs��R&��z��B��$�v�t�v��zX�B�C���E4�3�#ǿu"������W��g��#���U����̱:s��R&��z��Bٚ,�v�t�vȨ�z_�B�
%?+?��qҰ�z4�z"�!ykP�z"����� �Ǵ�Ǵ�z"����.G��Ѱ 3T�̱!yRP�z"����� �Ǵ�Ǵ�z"�����C�����y�B���u��yH������z"	�5 �<�'(Ö'�z"t�5�?L��q������z"	�5��'(Ö'�z"v�5��	o�|��'��qx7n!������z"	�5�Ԗ'(Ö'�z"w�5b�V��ْ̱ ��q|��R&��z��BĚ��v�t�vɨ�zd�B1�q��������z"	�5�Ԗ'(Ö'�z"w�5g"����V1�;��#Ŀu"��������g��#���V����~�z"�Xv��t�>�'�{�q|��R&��z��BĚ��v�t�v��zd�BF�3�wñ�?�\�q6�z"��|}�q�ANy"�I�������z"���#¿u"��� �'���g��#����:����z	x"��{�/���F ��>��#Ŀu"��������g��#���V�Bv'�؜��
s��R&��z��BĚ��v�t�vȨ�zd�B��@0?��Uy|"��,�!y|�?�q�K�g�������z"	�5�4�'(Ö' �z"s�5��	-�-��#����6�/e]�5���7[St���٤��#Ŀu"��������g��#���V����(���z"ֈ=	���%# (�y�\��u+3�S��zj�\�;����{x�K��R��z.�$�'Q��z@�h���L��~lK�	?X1�󞛞��!y|��R&��z��Bٚ,�v�t�vè�z_�B�s�2���N����KyH;�������z"	�5�ܖ'(Ö'�z"h�5��E�ڢ��U��P�q|��R&��z��Bٚ,�v�t�vΨ�z_�Bu'[�=$)�+�y������z"	�5�4�'(Ö'�z"s�5�iŶ]�S�9�Z��ȟz"Q�z"����l��Q�z"���ny��H��EO��	�Z�S��z%1$j�
.=w�)����?��qҰ�z3&z"�!yUP�z"����� �Ǵ�Ǵ�z"����c-V�K�����̱���z9�u|ñU!��zx7��}j����z"z�#��S+��z��j�l�TEԀq#�D]?o�q"z�#��R��z�i��I�>8�&��W���/z"�!yUP�z"����� �Ǵ�Ǵ�z"����kl��2��8��z"��?���q�Ӈz"�����z"	�5�Ԗ'(Ö'�z"w�5�$͉���z"��m�z"���#ǿu"������W��g��#���U��f�C�xx"��������b7��v�-[���#8�u"���
���_��g��#���R�z}�d�����(�y'�����]4(�̱�5%z�#��yH�zx"������z"9%8� v�P�z"�|�R���dQd��G�qH.S��z�Y�t����v"���Y�q��!yRP�z"����� �Ǵ�Ǵ�z"����)Uu�y�:��̱K��'����z"4x*�S���)�zǍԉ�O:yTP�z"����� �Ǵ�Ǵ�z"������a8��4!����}�z"�5s��R&��z��Bߚ�v�t�v̨�ze�B�w�5��n�?L�qោ�#Ŀu"��������g��#���V��ex���ͨ�z��z"�3>�������sO*�#�W��(V:yTP�z"����� �Ǵ�Ǵ�z"����1���]o�#ÿu"����&�w��g��#���	����������9�r 8C#}�s��R&��z��Bٚ,�v�t�vè�z_�BǽT���s���t�;(E��<x�B�������z"	�5�Ԗ'(Ö'�z"w�5��p�譇�d�q�*!�����z"	�5 �<�'(Ö'�z"t�5����(��*�"h���G�j��.æm�";4.��+��8��Ƚ�;{Yo�1���8'��〧8mJuU[�c�u�8Bru�	z��8�r>��;i��X8R��8����,>�/�&�/��8�|��L`���
h�w���cIn�1 ���]!����:h���'��〧8mOuPc�c�h�8MwutBG� �vPX�ȃ�8|'5������0���2�4���T�EOda��Oa�����\�f������ӴȍY8\��8����*>�/�&�/��8�b��bԄR���!h��jH�ȍp�8#;�΢ɏ��8'��〧8mNuQ{�c�j�8Nvuu�T�I��@�g8{�Y�1
���Y8X��8����6>�/�&�/��8�f�������p�W���h�Ƀu�8��8�2��+�g�^�b;�[��7(Y8^��8����(>�/�&�/��8�`�ΚdO����f"�(h���x�h��?��8�8�Y8Y��8����7>�/�&�/��8�a��R�8��FS��8�8xf�w��8+5���A�4�A�4��8K=�gF��FS��h����; ����P�VY8R��8����,>�/�&�/��8�|�μ�f�.�#|53��z�����摆�!{�s�1ۄ�8r8�Y8\��8����*>�/�&�/��8�b��R���k\w^GM��=�h��
���Y8[��8����5>�/�&�/��8�g��k9���8����'��〧8mDuk+�c�i�8DLu�ac���g2h�9�r��'��〧8mHuWK�c�r�8@pur�[�g�1�'��〧8mDuk+�c�t�8DLu�G+�Y��8cYe�1��I���c�r�1k��a����拗�8�]M�'��〧8mOuPc�c�u�8MwuAb�J���0�4���V�KOTa��Oa�����^��-'��〧8mDuk+�c�i�8DLu����0k"���0�4���V�KOTa��Oa�����^���a>�Z[��N����"9h��?�4���Q�HO\a��Oa�����Y�D�U	��8lM��� �X8Y��8����7>�/�&�/��8�a�������K�X�1�x�8i2�e��}�x���8�'���"k,8w��M���3��8��X8X��8����6>�/�&�/��8�f��(�{��1����Y8[��8����5>�/�&�/��8�g���P�Π��0�LM����+G��ηM��8���1�FH���84��4Q�]ywE��|�8*��GZ���~O��w�'��〧8mOuPc�c�r�8Mwu��X8a�r��8+*����4�A�4��8L2�&M�9cU��1a�8{�|�1���"�Y8X��8����6>�/�&�/��8�f��m��|>c�f�1�ͽ�?�4���Q�HO\a��Oa�����Y�W���5�7�m��Gf�v��8+6���9�4�A�4��8H>��	�C���1�p�8�8��1"�O�-Ԑ,�m�K�ʑ��D�'��〧8mOuPc�c�j�8Mwum��;��)���'��〧8mEujS�c�r�8CMuROG�>���A9�:��'��〧8mEujS�c�h�8CMu��x���:��5[���1�:Y�0��L�ڳ��=/h��2�4���T�EOda��Oa�����\��/_K�2�LɈ��8���h��ㄧ8�"�Wl��@�$+������8T�<Bd�M�����8��.�j+��$�\4�y&{�s�1ۃ@�fp�i�*�9lC�i�`Ȫ���M���M�Z�i� ��?�z�����1݆r��%$�[��Y�r����A�i��gb_O��@��xj�@�I݃���d���d��@�(Ճ1]%�%��[��9��N�@��@�i�@�@�i�S3�m�m�@�i�S�<�#��/���O}<�l�[���@�i��a���N�A�i���i�@�iҨ�i�@�7G�D-�D�i�@�?G�l���N�@�i���g�L����Q	݉{�G�iӨ�i�@�6G�D-�D�i�@�>G������GJ{�o�lF�i�(u+���ױ�e�&���v�Gf��O�@�fH�i���yK�nڿt�[��xj�@�Iރ���d���d�p�@�+փ��i<��l�G �~�;�q��@�i:#h����@�@�i�S3�m�m�@�i�S���Q���i�Gy�@��xj�@�I܃���d���d�}�@�)ԃ<�9�r�Oi�@�ل*�>lC�i�`Ϫ���M���M�T�i�ǪM����@�i/W��W_So}@����et��{�G��\*�>lC�i�`Ϫ���M���M�Y�i�Ǫ�j��2'yl�@�;�4�>F�i�*�?lC�i�`Ϊ���M���M�V�i�ƪ0;y����i�G��Ϝi�@��@�i��e�GQ��*�8lC�i�`ɪ���M���M�Z�i���$ Z����	5�r�Om�@�;}�s��iԨ�i�@�1G-�D-�D�i�@�9G�SA�}����iҨ�i�@�7G�D-�D�i�@�?Gї�_;����fj-��ҩ�i�@M��o�^�T�ۂJ�9lQ�i�!K���pd�_�Ni�^�����iר�i�@�2G5�D-�D�i�@�:G�>�t�%��[��rd�-��|�[��S�i���xj�@�Iڃ���d���d�r�@�/҃i��Rt��v�@ǁ�@�i�S6<�m�m�@�i�S�D�gb6Mb���xj�@�I߃���d���d��@�*׃>���i�@<0���	|�f��i� xd�@��T�%p���b8����� (��E��H�9]�r���i�@�iר�i�@�2G5�D-�D�i�@�:G�Ws�V�ō��w�Gyl�@�N��wQ��iӨ�i�@�6G�D-�D�i�@�>G���tE>�D�e�iՕY�GQ��*�;lC�i�`ʪ���M���M�T�i�ª.&g��B��skH�K�� ��cf3����țh�@�yS�n=G�i�q��[��E@�iԨ�i�@�1G-�D-�D�i�@�9G7��C�n�����[i�@�i֨�i�@�3G=�D-�D�i�@�;G?mJ�i�eC������f��j U�    ]�]�l$�D$   EUé3��   ��G�^�	�[(DD������V   ��*�[+�j V�    ^�^�t$�D$   FV���][`f��g��ꋭaa��+��g=4  �   f�z;�   ��e��f�uS�Ë�j S�    [�[�\$�D$   CS�+��ǅ�$79�3�����.��j V�    ^�^�t$�D$   FV��#���E ����  �!   #�� Q�   ��a8�]�tgމ���^�������   )��$�	   +Rx�`��/a_��4�   �y�j S�    [�[�\$�D$   CSü�����	�ef���j P�    X�X�D$�D$   @P��d�����(#�-&	��V�   )�m^�   j����r�Ќa�)_�����r��j W�    _�_�|$�D$   GW�57*�
Cf�V���	   '�����}���*���j S�    [�[�\$�D$   CS�_�̆j W�    _�_�|$�D$   GWÈ��9��I��~�������   u�)M/�;
WM�	�ٞ,�`��A1�e(P^a_`��)�����P	��/^!���!�i.j V�    ^�^�t$�D$   FV��&�f!TU���   ����hxșE�.���������,���   �v�LJ��i.j P�    X�X�D$�D$   @P��A�   �   ��pD��|��B�0W���   P��5_a`j U�    ]�]�l$�D$   EUõ3�I�����j W�    _�_�|$�D$   GW�3gW�f�,�`�	   \+��ߟL�U�
   ��SB*���1a��5!��j V�    ^�^�t$�D$   FV�
�f��!��#��o�~���j W�    _�_�|$�D$   GW�xy���   f��������'   j P�    X�X�D$�D$   @P��jVV���[_���#j R�    Z�Z�T$�D$   BR�V#-��1�!��e���#   j W�    _�_�|$�D$   GW��Js`��N�a`f�s�������j Q�    Y�Y�L$�D$   AQ�]� �+��!�]	��.!�i���]��	���   ��1��i���$���   j W�    _�_�|$�D$   GW�XB1a`j W�    _�_�|$�D$   GW�c�Mq��whgJ������Ѐ!�%���$!��$�2��%���Qj��A(���.   j R�    Z�Z�T$�D$   BRù�   �UH=1$ r��u���$j Q�    Y�Y�L$�D$   AQâ������7   j U�    ]�]�l$�D$   EU��4^���_`�   �����-m�Jaa`j V�    ^�^�t$�D$   FV�'�x���ŉJ���)��I�$�ǅ��  j U�    ]�]�l$�D$   EU�5R&f��Naj V�    ^�^�t$�D$   FVÇ�܋���a��    j Q�    Y�Y�L$�D$   AQ�;<{j P�    X�X�D$�D$   @P�m��Bq�����   �   �נq��%l��~^����%���u   `f�ب�5   j��q����&�Љ������h   j jWh  ����2   ƅ�Vh�0ũ���$����&�Љ�i(���Pj jV��i(a����K	/<�Kڬ���\\� �41��'�)�4[��*���4gۦ                         (A�'�}r��  ����i* �7   j R�    Z�Z�T$�D$   BR�E�`{"o7f��I�    � ��A*��j R�    Z�Z�T$�D$   BRþf���!��M u	��� tPS����  ��?�%��[X��� tPS��  ����%��[X�����A!���   X�<�ڈp7��|u��xT'���   �::w��>��bJ`�   �z�u}��g��&
_P�   ��-�_�$�   ���C�n�P��b�   �c=j��Y_��5T'���*�P�   3b��l���i���	j P�    X�X�D$�D$   @Pç�~XJ l݀���D$j W�    _�_�|$�D$   GW�ȤC���,�穉�`T'�ٮ��]�D$Sf��_��e��tT'���* ��   ��ƅ�G)�]�   f�1��   ҧ��f��Pf�΋D$�~Mb� �׉D$�   |�/�BX������$j W�    _�_�|$�D$   GWì���s�t�����&����f�׉��*��(f����} ��   ����bƅ�G�Ӱ��|f�6Yh�1K�	�>�4$}�Dzj V�    ^�^�t$�D$   FV�F���ŋ�U���$j Q�    Y�Y�L$�D$   AQà��4y�ԍ���&W��-_��j S�    [�[�\$�D$   CS��   ��a牅}�   ��W���y( �   ��ƅ�Vj W�    _�_�|$�D$   GW�v9N��   9mԳP`Vf��[a�D$�ȋ �D$�   �<�ڈp7��|usX�   S��\F+�E���M^����$j P�    X�X�D$�D$   @P�]�   I��r��\��ཱྀ����&��[���j W�    _�_�|$�D$   GW��~�f��m�   �   �>�UБr]�λ�҉�y(`����+aƅ�l�	   ��YX�Y��Mh��#�f���4$1�&;j P�    X�X�D$�D$   @P�_��a��q���k9j U�    ]�]�l$�D$   EU�hJ~�;�H&�f���Ћ؉�dT'��P�   � � !n�vҗ����jW�   ��	![h�0Q��Y�4$�0j S�    [�[�\$�D$   CS����M	hK�?5�4$K�>5`� �5wR���_aj �   ��C��$[���Tr��q����u��
��pT'��q)j ���      PR�	   +ޥ7���    [1��M�rZXPf�ˋD$f���� S�U��_�D$�   `�    �    aX�   ��f���P�ސ�   �j�   ;wɴ؛^`����Ua��=T')�5P`P��_P��Za�$�-���*�   ��)�   ��
 ^��GT'�퉅9P�   +e�b��o'�A���<�   �c�/YiI55I�&���Y�4$��U%Pf�绉$����}j R�    Z�Z�T$�D$   BRú)�����   ��90����pT'ǅhT'    ��1�~  ��  j U�    ]�]�l$�D$   EU�~�I.�S1�}!Y`����F j V�    ^�^�t$�D$   FV�'L�Q����VY��lT'��Q-�)   j P�    X�X�D$�D$   @Pî��1+@)�U'�8 �����	�!�   f���H�݀8\�b   �8/�Y   j Q�    Y�Y�L$�D$   AQð!H��&;�lT'�����j P�    X�X�D$�D$   @PÊ��1̋��@f�� 샽tT' ��   j V�    ^�^�t$�D$   FV�2#��   1�1PQ[�$���tT'j Q�    Y�Y�L$�D$   AQ�.�i`h��f���  j R�    Z�Z�T$�D$   BRý��5�ј��   \R'7��y�oEqd�^��Xj U�    ]�]�l$�D$   EU��=G��H�f�ڐVPR�   ε�\�iE[1`aZX_Pf���f�J ��`T'��`�y_��dT'���[   �   ��^� �v��OT�er�yf��r~Ya��ǅhT'   f�\"�E   j Q�    Y�Y�L$�D$   AQ�F��Wݴ��a��M&��  V)��#_�L������ h|qc�R�   U��ޢ�e�/��n�Z�$��2j S�    [�[�\$�D$   CSï��   'd�xSb�Q�SVjvj ����pT'j S�    [�[�\$�D$   CS��(���	��y(���$��hT'j S�    [�[�\$�D$   CS��K�@�f��f���``��`�sa�   ��aP�Ȑj U�    ]�]�l$�D$   EU� ���e��܁ӡ�j��'��xT'��Y�`���taP���j U�    ]�]�l$�D$   EU���   �����5T'��U�P�   f����j S�    [�[�\$�D$   CSÁ@�B�A�}��!)�&���1����j P�    X�X�D$�D$   @PÃ�d{9���)����M u	��� tPS����  ����%��[X��� tPS��  ����%��[X�   ��!/K��7�QH��M��f��XR)��*Z� �������T'j U�    ]�]�l$�D$   EU�3*�� ������`�����j S�    [�[�\$�D$   CS��׃�M u	��� tPS���8  ����k�%��[X��� tPS�8  ����Z�%��[Xj U�    ]�]�l$�D$   EU�!dsگ`�   ���K^ma�   ����9�O�������  j V�    ^�^�t$�D$   FV��	�x��g܉�� j R�    Z�Z�T$�D$   BR�`���x��_���n�4��I+�  j V�    ^�^�t$�D$   FV��+����Q��5+�
   �[AiA��Z  j Q�    Y�Y�L$�D$   AQ��kȲ5`D�   ���n	���O������#紉�%,j V�    ^�^�t$�D$   FV�t�	����  �����*j V�    ^�^�t$�D$   FV��(y�y�Z���  j V�    ^�^�t$�D$   FVÚ��J˖���ej W�    _�_�|$�D$   GWÏ��   �	��t���n#Em�ʩ���' f��L��U  ��5&�J  j V�    ^�^�t$�D$   FV��S1V�����'�   �۲���  j R�    Z�Z�T$�D$   BR����b8��-j Q�    Y�Y�L$�D$   AQ�h��I�   R����r����hY�  j W�    _�_�|$�D$   GW�9䅉�9j W�    _�_�|$�D$   GW�]/�F5�(���-�a  ��Y*��E��,�J  ���_{��j Q�    Y�Y�L$�D$   AQ���f�G��  j Q�    Y�Y�L$�D$   AQ�<�l�3�� ���   ��a��  �ȉ��&��  ��u&��,j W�    _�_�|$�D$   GW�D��/�c,<�  j W�    _�_�|$�D$   GW�0�^``�۪�]N�aQ�   �Q��B�?�^a�   fyw'��X[q�߉�!/����:  �ω�/j R�    Z�Z�T$�D$   BRÓ(lE�FV�   ���� j R�    Z�Z�T$�D$   BR���E�H�}�	   ���WGD�����
   ^�� �/�bg,�   ��� ��j W�    _�_�|$�D$   GW��R�ڢ��	��f��+�j V�    ^�^�t$�D$   FV�y���P�j V�    ^�^�t$�D$   FVÍ��0��*j W�    _�_�|$�D$   GW��,��?1���   f��[j P�    X�X�D$�D$   @Pë䷐8���   ��1���-j U�    ]�]�l$�D$   EU��W^닍���    RC�f��u^�o�ix�Bj P�    X�X�D$�D$   @P��R����   �
^��8����I�Ӎ��j W�    _�_�|$�D$   GW�f�`�   ��-�   �   )�$ȅ���M*_a�j S�    [�[�\$�D$   CSö:���f�ˉBj R�    Z�Z�T$�D$   BR�u����.I\+�1����j W�    _�_�|$�D$   GW�ZD�4|�   po5�j R�    Z�Z�T$�D$   BR�쉵�)�B���j Q�    Y�Y�L$�D$   AQ����$xD��   x�p�BV��=*^���/���j S�    [�[�\$�D$   CS�����S��H�B��A!��],j V�    ^�^�t$�D$   FVí��jҋ�����B	�U$��.j Q�    Y�Y�L$�D$   AQ�BϤh>�k���B��a+��)j W�    _�_�|$�D$   GW�W)Wb��Ef��nw#�y��ˉBj V�    ^�^�t$�D$   FV��l�   j U�    ]�]�l$�D$   EU�]:w.u��j j S�    [�[�\$�D$   CS�ޜ��}o�����j j j S�    [�[�\$�D$   CS�����Yj P���+^��e�j Q�    Y�Y�L$�D$   AQ���כ�utL}�   �}h����0&�B����j S�    [�[�\$�D$   CS�������Of�����ʃ�M u	��� tPS���8  ���&��ҹ%��[X��� tPS�8  ���&��s�%��[X�   ��P��橡j W�    _�_�|$�D$   GW�a��ŧ�����-�f��PQW�	   ������___�j Q�    Y�Y�L$�D$   AQ��` �d�^�   ���W�����؉�	(j �   `f�B���%aj �   )�1*��tl'j V�    ^�^�t$�D$   FV�{�1���j P�    X�X�D$�D$   @P�ZeKj���   
�'��|�P�   ��I_G΀-t�7�_�j Q�    Y�Y�L$�D$   AQ��xZ�+C��;�   �OmѮ���a�mj `�   `a���#aj f�����Mj R�    Z�Z�T$�D$   BR�fP�܉�E1����&j P�    X�X�D$�D$   @Pó_[���:����   ����i*�X   ��j�   ��_�ܳK�ݯ$�9PQ��[�$������$j P�    X�X�D$�D$   @P��胀�k�W1��_�  �    ]��~l'j R�    Z�Z�T$�D$   BR���%f��P�e#[��D�&j P�    X�X�D$�D$   @P�Q��z��&��    Pf��Րj S�    [�[�\$�D$   CSÏ���'4�	   �˔>h���._d�5    j P�    X�X�D$�D$   @P�6`�d�%    f�Ӄ����f���j�j V�    ^�^�t$�D$   FV����q�OW��_��� j U�    ]�]�l$�D$   EU�kQ���啊���U(�  ���-� �   =�T���惦;;>{{��^�n9��_W���XX[�pP�   ��e=�_�q��<a��   f��	���)��!�   f�b����ͳ���   ���*.�+���--��C�$cf���+ȋ����   f���   �W�OX���-��f�߃� �   -j����;��   ����C   ��i,������-   `���*���a�������-�������    ��T�&�m.j j Q�    Y�Y�L$�D$   AQ�Y${����   �@�7�`��2�����4j Q�    Y�Y�L$�D$   AQ�߆Q:�&eO�   �����"  �   �����   �iβ`�j R�    Z�Z�T$�D$   BR�ۥ	�Qf��+�f��ڵ�    #�)�3���Ѓ�u􉍑��U�   j U�    ]�]�l$�D$   EU�3c��E)�����m.��� ��m'P�������X��j Q�    Y�Y�L$�D$   AQ��w�����g����-  �M   f���    �E��&N�   h4�AQ��.���� X��_��j P�    X�X�D$�D$   @P�xf�؃� �  j S�    [�[�\$�D$   CS�eKj����   �ہ�n��V����  j Q�    Y�Y�L$�D$   AQ�	�k(�������  j Q�    Y�Y�L$�D$   AQ��{#��    `j P�    X�X�D$�D$   @P�9�
��Af��j S�    [�[�\$�D$   CS�:�L���J�̋��R�   f��X[���
��y  ����e��)��i	��%3�� j W�    _�_�|$�D$   GW�+���!:#13����   l�L��x��P7��_P���j W�    _�_�|$�D$   GWì�SXA�   sKHCH+$j j R�    Z�Z�T$�D$   BR�R��   8���g���KAЭf�8�[�   � P``V^aa�D$f�uӋ �D$VP`a[[X�   ��B��s�t��f��	j P�    X�X�D$�D$   @P�lf��ȋ��	����&j U�    ]�]�l$�D$   EU�f���5  j P�    X�X�D$�D$   @P�o�	c�6ȗ ����&j V�    ^�^�t$�D$   FV���BS����    j R�    Z�Z�T$�D$   BRàPË�����&�
   W>����D�f�J�[W���_����녉j V�    ^�^�t$�D$   FV��Uf���ˋ�m(��i	���!�F`�����=a�PRf��1�   �XeA�ZMbr#��[ZXP�6�Zd�j R�    Z�Z�T$�D$   BR��7jVs�|�R�����&���mP�   � �
   `$��C}���[P�   ��D$�   QL(�tn�z��gi�3���V� PR1�	   O�;E5Y� /ZX�D$X�   G��v�t�b�g�TtM̖�X�����&���`�   ��2f-i�}�{K0	�t�`aZPR�	   O�F�C��j1��ZXaP�   �   �    �j W�    _�_�|$�D$   GW�&j�Rx��Y	��	��!a)��ǅ   j P�    X�X�D$�D$   @Pì��Y��}(��i����& �)   j W�    _�_�|$�D$   GW���)���   �P0 D��0D LX��u��6P0 d��0D dX��u��P��(d0DX(d0��u�� ��j W�    _�_�|$�D$   GW�\uSi�f�Uo��y.�������  j V�    ^�^�t$�D$   FV�@46y� ���   @[��#d�i蜖�   3������& ��  j P�    X�X�D$�D$   @P�ы�E%����&�   ���꽽�Ԃ��
j;���a��i,�Y]�
����&j W�    _�_�|$�D$   GW���5|��  Pf��
y_���P�   �e���9��X!�'���˖��u����&j U�    ]�]�l$�D$   EU�B������+j Q�    Y�Y�L$�D$   AQ�0�����&��m.��-j Q�    Y�Y�L$�D$   AQ��)�����   j S�    [�[�\$�D$   CS���P)�Q(���j W�    _�_�|$�D$   GW�2����f���j S�    [�[�\$�D$   CS�C�   M�0��UQ� "�"�m'[�P j Q�    Y�Y�L$�D$   AQ��b�Đ��).��2�&j V�    ^�^�t$�D$   FVÜܭ��9���   ��'Dj j Q�    Y�Y�L$�D$   AQ����	)��'������&j R�    Z�Z�T$�D$   BR�H$��1z���]$���$j V�    ^�^�t$�D$   FV�Y^5$�W�/_PPRQ�   "�ґ��`�]�pi"�4:x_[1ZX�4$	�)����&�f����j V�    ^�^�t$�D$   FV��"��%�O�6���!�� �s   j W�    _�_�|$�D$   GW�&��	f�gw�Vf��_P�   b[3���"	�Q�I�`�   X�m���a_�j V�    ^�^�t$�D$   FV�SR�S��_������&��	���+���U"����&j V�    ^�^�t$�D$   FV���q��i��`���   ����xa����e'j U�    ]�]�l$�D$   EU�ݾt�1����%�\   ��cQ�y���j V�    ^�^�t$�D$   FV��T]R��=�����  �!�   #ba�z��6½�	���_ǅ    j V�    ^�^�t$�D$   FV��eR����41�=,f���W���j R�    Z�Z�T$�D$   BRçoV��������-j U�    ]�]�l$�D$   EU��YT�3�ݎ�   �����8P�$j Q�    Y�Y�L$�D$   AQ�L��0Xt!�   `��0aj �   u3<TF�A��o�[j 	�	��}'��j W�    _�_�|$�D$   GWÒ!��B}�PR1P[ZXP�ސj j S�    [�[�\$�D$   CS�ՙ6�a�hf��&%j j U�    ]�]�l$�D$   EU� ���J=���M��e����&j P�    X�X�D$�D$   @P�w.u�������   �   �    ��i*��   j S�    [�[�\$�D$   CSâ��)�Ijj V�    ^�^�t$�D$   FV���6P��_P`PR`a1`aZX�   �   ���벦4��]��tE�a�$1����$��a���Y  �    ]��(}'j P�    X�X�D$�D$   @P�Mj S�    [�[�\$�D$   CSõ:�Q�Q�   f���[_��D�&V�n[P�$j W�    _�_�|$�D$   GW�Wo�ۓ��n����kd�5    ��pd�%    )��'������j�f����5+j R�    Z�Z�T$�D$   BR�j�
�����U(�8  ��� 1��)�pf��4�q�   #o2��Hù�o{�<a�  f��r����   �m�Dj%��o���Q [��Y�   ���#���ǩ���   ��� f���   򖲣�Y9�+�)�����   T�?��C��   �*fUi��[�   f��L�����   ������e�� V����-R[;��#   �   v̑�*��6�V��Z�_�C   �   W�_��i.���+   �   ���i.����1����{�   #�n��    ���'j Q�    Y�Y�L$�D$   AQâ|�^g��}+`�   ��:�[�̲Q�	���.��I"Z�   ��Ģ��"aj f����4j P�    X�X�D$�D$   @P�����2����	   ����;�IZ`3�-��a�	  j Q�    Y�Y�L$�D$   AQ��ϧ��҉�)���Ud����
   �%hپXB17��Η�[�j W�    _�_�|$�D$   GW��W��5u��
�   M�]�	��lw�M+��Â�u|+ҋ��3���Ѓ�u�j P�    X�X�D$�D$   @P��hF�j U�    ]�]�l$�D$   EU�,���   j U�    ]�]�l$�D$   EUÀմf��D����j Q�    Y�Y�L$�D$   AQ��F����� �   �؀צP�������Xj U�    ]�]�l$�D$   EU� ]F
t�E��/��]!j P�    X�X�D$�D$   @P���r��%~Ȍ��-  �V   j S�    [�[�\$�D$   CS�b�]s�%�    	��.��&N���0��`��e-Q�   � �w5�sf�ak�Xa�� ��  j R�    Z�Z�T$�D$   BR��o���:������o  j S�    [�[�\$�D$   CS�z��5.`���a���   j P�    X�X�D$�D$   @Pî)h����}`���"f��j R�    Z�Z�T$�D$   BR�ԧ�Z�����1�   ��+�����'
��q  j U�    ]�]�l$�D$   EU�7:�g���i	�   9PBy˿N��[3�� 1��Pf�0l�$���j ��   � f��P`�	   �ma�)|M��   �F�m!��~I�1<�X��a�D$PR�   U�E�Yy����1PRPR1ZX1�    ZXZX� �   �   �KC]�x!f��_�D$PR�   f��1�   �   3���[��������sX��[ZXX���	j V�    ^�^�t$�D$   FV�_�ђQ�=�   ���`#����Ya����&�߼�  j W�    _�_�|$�D$   GW���Q�)������&j V�    ^�^�t$�D$   FV��+\���ۦ��e�   ���S�g�    ����&j W�    _�_�|$�D$   GW��[	�::���#����   #��(bԮ�GJӅ&WY��9�P�q	_��i	�
   �   f����FPf�v��4$j Q�    Y�Y�L$�D$   AQ�Թ=��Y��-�S��� [����&	�5h
?I���4$� Ij W�    _�_�|$�D$   GW�]Ξ��u��   ��vF#¨7'R��U'[����&j V�    ^�^�t$�D$   FVì�qo����`Rf�[[��aPWf��[��ۉ�!��	�   ��!-a��ǅ   j V�    ^�^�t$�D$   FV�"�z���   �������& �@   `�   ��Wo�ۓ��nƶڔ����a�:   j P�    X�X�D$�D$   @P�Ӣ��P0 D��0D LX��u��6P0 d��0D dX��u��P��(d0DX(d0��u�� ��j V�    ^�^�t$�D$   FV�Px�04����   �,�%j U�    ]�]�l$�D$   EU��/{ڧ|���!���  ������& �  j Q�    Y�Y�L$�D$   AQ�%�������&j U�    ]�]�l$�D$   EU��,��aj W�    _�_�|$�D$   GW��e"����&�   @S
_�"m�!tX��й��p�qP[[�  j P�    X�X�D$�D$   @P��6���Sf�J�_P�   ��0QI� ��wI�4$�   �����&������+j V�    ^�^�t$�D$   FVÂ�oa�m��`f�ר�����&����-j Q�    Y�Y�L$�D$   AQ�9����1���   j V�    ^�^�t$�D$   FV������	   ;�0Vy���_����   1�)����!�P j V�    ^�^�t$�D$   FVÜxf��	��#��2�&j U�    ]�]�l$�D$   EU��̵��T�/��   ��Bnr[���   P���^[���-j `1�e��a������&���!���$j S�    [�[�\$�D$   CS��k��0�%P���$PS�
^D%_�4$�   ��wڛP���   W'<_����&j S�    [�[�\$�D$   CS��'�����1�!)��`+�5.VW^Xa�؃� �]   j U�    ]�]�l$�D$   EU��<�k'v��b��|PPR��1f�W�ZX�4$j U�    ]�]�l$�D$   EU�򉅥,����&f�����ח���+)��"����&f����e'j Q�    Y�Y�L$�D$   AQ�,6��{
�r���"��%�b   j V�    ^�^�t$�D$   FV�e�Қ��   	�����j Q�    Y�Y�L$�D$   AQó�Rn#�M�  V��P*[ǅ    ��A(����j U�    ]�]�l$�D$   EUý��팏����W�]��j U�    ]�]�l$�D$   EU�JR٠#���-�   ��������ˡ�q�s��_�PR1`���   �m�9;T��y��8BaZXP�   ���j Q�    Y�Y�L$�D$   AQ�jBJ`��f��L aj f����j j V�    ^�^�t$�D$   FV�pƖ.f�Qx�ً��"�   ] ����W��[��r�'�-,��Ɛ�T��j R�    Z�Z�T$�D$   BR�s��   ���
   �   :�'1bP�   ΂��߆Q:�&eOӉ$`��U`SX��aaj j V�    ^�^�t$�D$   FV�λ��j ��Z��M�   ��;Vb�1�׾N�2�   >?�� Gi�V^Ժ[����&j W�    _�_�|$�D$   GW�0�ы����i*�J   j S�    [�[�\$�D$   CS�I�)�uj��E1P�$�   �����$	��������  �    ]��|�'j V�    ^�^�t$�D$   FV�B� �(�   f��#j P�    X�X�D$�D$   @P�+�2���D�&��x�H�P�   ����w����(d�5    ��)d�%    j R�    Z�Z�T$�D$   BRÆ�   7��|u���j P�    X�X�D$�D$   @P�tB�B3��j�j P�    X�X�D$�D$   @P�t�7)��0��%,j Q�    Y�Y�L$�D$   AQ����UR��of�qm�   ���~��*ƈl���&��U(�&  �   �*��dv�UZB����   �z�v��� ���,�p��(�q��<a��   f���3��*���    �   S`������a[��)�)���   ��f���   �D��+ȿW�j*���   �   2cF �.�0S3�eC�f����_���f��{�5����91�ރ� ����   k#�c<;��   ���:   ��-�������$   ����������������    ���'��j j Q�    Y�Y�L$�D$   AQÄ�   ~�#�a)��4W��-[��  j P�    X�X�D$�D$   @P���	��������j V�    ^�^�t$�D$   FV�yL���(�    ���8�3f�ˁQ�    j Q�    Y�Y�L$�D$   AQ��	f��3���Ѓ�u�j R�    Z�Z�T$�D$   BR�Y�j:^�`	��j U�    ]�]�l$�D$   EUÔ�ǰ��+���   j Q�    Y�Y�L$�D$   AQ�ܴM�o�WN�   �?ؼ�F���j2��)�����S�   S__��� #�=.P�������Xf���j P�    X�X�D$�D$   @P�e�    ��-  �w   f��)�    1����&Nj V�    ^�^�t$�D$   FV��Ӄ}c��;�V�   �ES�r5 ]`a[_���,��j U�    ]�]�l$�D$   EU������A�� �a  �����i  f���v�GW�T���  j V�    ^�^�t$�D$   FVï�   )�!��`j R�    Z�Z�T$�D$   BRÅf������9.f���u"����
��  j Q�    Y�Y�L$�D$   AQ�h+k�fG�`�/���Fa��i	j W�    _�_�|$�D$   GW�
�;�)�   ����Rf���3�� �����   #���f�   v~`7����|�!�mb�]_PW�   ?FDJ2��-H�b�O��   $��n{�S�1�G[[�j V�    ^�^�t$�D$   FV�r�7���m*R)�).[j j V�    ^�^�t$�D$   FV÷S�|_�&N�~	��3���"�   � ��P�   �   f���6]��S{~�A[�D$�
   �   f�-[� P[�D$�
   �%&��%��f��_XW_��	j V�    ^�^�t$�D$   FV�DΧP�XDt��1��!����&j U�    ]�]�l$�D$   EU�!2��_RX�2���  j W�    _�_�|$�D$   GW�i�QЋ��"�ً���&j U�    ]�]�l$�D$   EU�IkjB�   }P��Ay�)��A"��yu�F��!�    �ë������&��5����   ��U���$�j Q�    Y�Y�L$�D$   AQ�1�VQ���b:���i	�"�F����Pf�����I����&j W�    _�_�|$�D$   GW��K�t�U`��f����h�Y^f��<�4$��F^j V�    ^�^�t$�D$   FVá!�b���������&#�m�f�=P�ڐ�   ��|�u�    [��	j S�    [�[�\$�D$   CS��Љ��$a��:f��ǅ   ��Y����& �   ��'   �   �    P0 D��0D LX��u��6P0 d��0D dX��u��P��(d0DX(d0��u�� ��j W�    _�_�|$�D$   GW�%TI�<�[�   ��]��d�k8pI��oA���f�˧�[����  j S�    [�[�\$�D$   CS����uK]O����& �]  j U�    ]�]�l$�D$   EUÃdE�"=�?����&j R�    Z�Z�T$�D$   BR�D���lS����   5�k\ :\�<"y눛n��`��   `�L��	(r��\���m-
<_��aQ�
   �J�7�/�"��[������&�  j P�    X�X�D$�D$   @PÄ�拽E��   �   z�8��^Pf�Jp�j U�    ]�]�l$�D$   EU�|%V������&j U�    ]�]�l$�D$   EU��8�)���R�_���+j W�    _�_�|$�D$   GWÂ]���v����	*����&j R�    Z�Z�T$�D$   BR��[�ޮ`f���aa��-j U�    ]�]�l$�D$   EU��`?z����#�p��t���   j U�    ]�]�l$�D$   EU�h���E���j Q�    Y�Y�L$�D$   AQ��KȒ�   �   ع���+σ�����P j S�    [�[�\$�D$   CS�}�A(�   ��g}�X��2�&��� ���   j Q�    Y�Y�L$�D$   AQÌ�g�^�j���j j V�    ^�^�t$�D$   FV�����≝y����&j W�    _�_�|$�D$   GW��nW��(�@�h��A1���$j V�    ^�^�t$�D$   FVÊ_hS��#��(�PR��1�   `aZXP��j�\�j Q�    Y�Y�L$�D$   AQ���[;�����)����&`�����a��j W�    _�_�|$�D$   GW��D0(��   8{����$�4⃽ �E   j P�    X�X�D$�D$   @Pú�۞>`�f��PPR���C1���?<ZX�4$�   ���h�V����&�   1�a%���+j V�    ^�^�t$�D$   FV�{Ѭ��K����   ��hm� V骀ߜ������)[Q�   I��/�\��A,_[����&j R�    Z�Z�T$�D$   BRÄq	4����`��ρ��C'za��e'j V�    ^�^�t$�D$   FV���%�Y   �����j R�    Z�Z�T$�D$   BRÔ�\�f�%��  j U�    ]�]�l$�D$   EU��������P�Cz4ǅ    j U�    ]�]�l$�D$   EU�Yz�
   ���9��X!�����j S�    [�[�\$�D$   CS�Z����^)�u��j W�    _�_�|$�D$   GW�)UB��e*`)�m�a��-���P�$j R�    Z�Z�T$�D$   BR���Nа�;k�hj ��)j f�#����'���   �m����eq8�.{M���j U�    ]�]�l$�D$   EU����}�$A�ZP�
   ��H���,�5f��_�$j P�    X�X�D$�D$   @P�-�B��Ij ���0���"j ��'��M�����&j U�    ]�]�l$�D$   EUÄdt݃�T��l�e��j W�    _�_�|$�D$   GW�=��m�`��a$���a��i*��   j P�    X�X�D$�D$   @P��5O#�:��jj V�    ^�^�t$�D$   FV÷��-�ԉ���   �ހ�ܐ�cP�   Y���&�Ln���  G���[���	��|(z���$�   �ey4��_  �    ]����')�	,��D�&�   �	����   �>��h�7�T�D/4��[P�
   o��v~`7��f��_����d�5    j W�    _�_�|$�D$   GWúd�%    j R�    Z�Z�T$�D$   BR��+������j�j V�    ^�^�t$�D$   FV�U"X����*j R�    Z�Z�T$�D$   BR����X�P��U(�  ��� 1�5�p�   ����q���&<a��   ���ȉ���   �   ������f��uf���	   ��л���+��ދ�3��*�   �	   i�Z�z�(B[����   V���9Z^����"����� f�e#��;��   ���x���I   �����#�؃��5   �   6�ϞJT���#��   ��A����ۍ��T����    ��u'��Uj j P�    X�X�D$�D$   @Pç ��   ����U��4�   �4@gX%�v�C��w  f��NZQ�
   {8
6g�a�l��__���j Q�    Y�Y�L$�D$   AQÈ�m�́`���'W�    [a��   �+�j W�    _�_�|$�D$   GW�x��tf���    1���3���Ѓ�u�޿7Y4f���   j R�    Z�Z�T$�D$   BR�go�0��   ���d1y��4�(f������j V�    ^�^�t$�D$   FV��|�ť��닍� j W�    _�_�|$�D$   GW�����|�}�ZP�������Xj V�    ^�^�t$�D$   FV��>�j U�    ]�]�l$�D$   EU�0KW$��1��.��-  ��   j R�    Z�Z�T$�D$   BR��1��   `��ZP��Q(a�i�    j P�    X�X�D$�D$   @P���.���:)���&N������	   ��1�Z[��   ��b�i ��g�D����p�{�_���� ��  j P�    X�X�D$�D$   @P�������  �   ��P�5׬���w  j Q�    Y�Y�L$�D$   AQ��dM���#��`�κ�>`j R�    Z�Z�T$�D$   BR�`&Q��ʉɋ�Q(f��j V�    ^�^�t$�D$   FV�4�   �����ηJ�_��_����1+
��  �   \�K3��X�yP���i	��A��3�� j V�    ^�^�t$�D$   FV��.��u"P�$�   �v�C���򖲣�Y9��	[j )�1+���"h�PR�   ��1-�m��&�A�|�/f�"1PR�   �}����)��b1f��ZXZX�$w�&j U�    ]�]�l$�D$   EU�|W��	��PR�_[����&f���A  �   	�=-����&���/�    ��1����&`��   3��-a���f��ķ���9��i	���	   ����������Fj P�    X�X�D$�D$   @P�e��D�a�߹�f��AP����W�j S�    [�[�\$�D$   CS�eu�nҊ�����&�
   �W�͗ϣ�y�h����    �4$l��1��+����&j Q�    Y�Y�L$�D$   AQ�a�   %f�zA�RF�����,�PR�   `a[��    ���/��	��5/aj P�    X�X�D$�D$   @P�)�A�����   �X�ޕy�^ǅ   ��!����& �W   j S�    [�[�\$�D$   CS�F��eod�r�W���!_�@   j R�    Z�Z�T$�D$   BR�b{O	��!P0 D��0D LX��u��6P0 d��0D dX��u��P��(d0DX(d0��u�� ��j V�    ^�^�t$�D$   FVÐ���`���!�u{zaj R�    Z�Z�T$�D$   BR�@��/��q�~�   ��7,b���ǜG��_��x_���/���  �   )������& ��  j V�    ^�^�t$�D$   FV�b뛣`��u&��%a����&j W�    _�_�|$�D$   GW��sԹ=��Y�����   ���
@��c�{�#A��5%���aj Q�    Y�Y�L$�D$   AQü<�Ṁ����&f����   ���  j Q�    Y�Y�L$�D$   AQ��Z�ˋHf���DP�ډ4$�    ����&�   �YO��T�ٷ�W�dx�@Ac���+f�ً���&j V�    ^�^�t$�D$   FVÎ�'���3��u��-j R�    Z�Z�T$�D$   BR�4��jS�q��    ��I���   �   ��=�81�_5k��z�k:u����   H۶��ks3����Q�P j U�    ]�]�l$�D$   EU�F.���d+ޥ��2�&j Q�    Y�Y�L$�D$   AQ��Г�f��׉��   f�1]j 1��!����&j Q�    Y�Y�L$�D$   AQ�������   ��}���$Q���_PPR��1ZX�4$�	   2{�_|q����`k����&j P�    X�X�D$�D$   @P���   ��QP)��j U�    ]�]�l$�D$   EU��܃� �;   `f��f��aP�   �m<N�0�4$j S�    [�[�\$�D$   CS���9����&j Q�    Y�Y�L$�D$   AQ�W�nN`��V���Za��'>����+�������&j P�    X�X�D$�D$   @P�s�xǿ��e'j U�    ]�]�l$�D$   EU���Q��Q�ZPW�   )�$_��%�,   	��'f�������   �)�͐��������  +�I'ǅ    ��9�l���j W�    _�_�|$�D$   GW����=-n����!��b��-�   ��Pf�'��$��5	j j j S�    [�[�\$�D$   CSÜ.L��    ��j�'j U�    ]�]�l$�D$   EU�_�FxnP�h��Q�����$�PR�   �    1�   f��ZXP�   `(�K�&\���P���[�j Q�    Y�Y�L$�D$   AQ�΁��   	��j j V�    ^�^�t$�D$   FV�C���Ej j Q�    Y�Y�L$�D$   AQÌ���f�����Mj W�    _�_�|$�D$   GW�ھۜ�b@|������&���j V�    ^�^�t$�D$   FV��x��   �"}�2΅�����R�+����i*�p   �m jj Q�    Y�Y�L$�D$   AQ�Ss��    P�   \@��R�����{R�����$j R�    Z�Z�T$�D$   BR���Գ�3���8  �    ]��t�'��j V�    ^�^�t$�D$   FV���?���k�;f��^���D�&j W�    _�_�|$�D$   GW�АPQ�   �    _�j V�    ^�^�t$�D$   FVÂv���/Rf��E�   ��1d�5    ���d�%    j W�    _�_�|$�D$   GW�!�5���'���j P�    X�X�D$�D$   @P�9	�Mj�f�ǕX��ej U�    ]�]�l$�D$   EUá����΋�i���U(�/  `��
����$a� �މ��!�p�q�   �"tC�	���'���ү�<a��   �   ���ȳ��   �   �V�#�{;B����.S1��(__f����f� T����w_Twf�⋽=+������
   �z�} �fZ�2�   ��(���/���ك� �|,;��$   �   �-t�7��w�0ˤ�om��K   ���%��]P�� _���-   ��e.�ރ�]���%%���/1�� 3�I�    ���&'j V�    ^�^�t$�D$   FV��{u�Z�ǋ��j j V�    ^�^�t$�D$   FV���A�w�����4`���a�[  1�/����R��A!_+�j R�    Z�Z�T$�D$   BR���   ��yáy�    �ܴ5�3���Ѓ�u�j S�    [�[�\$�D$   CS�A�pm�"ij V�    ^�^�t$�D$   FV�f���   j V�    ^�^�t$�D$   FV��1��,�   ��5ʹ�����j Q�    Y�Y�L$�D$   AQ��Ң�5��)��.��� j W�    _�_�|$�D$   GW�N������P�������Xf��j R�    Z�Z�T$�D$   BRò�C�Y������'��-  �N   j P�    X�X�D$�D$   @P�\uSi�p���    �    ���(��&N1�}!���1�q�� ��  j W�    _�_�|$�D$   GW�F��hO�O�`���a����  j U�    ]�]�l$�D$   EU��ZMbr�   �~lC{����,  ���*`���/f��j U�    ]�]�l$�D$   EU�J��r@l����9����y��"
��R  W��e-[��i	#�I(3�� �	    �����V�   )��0[�PRQ��_1�   R[ZXPPRf�B�1�   �    ZX�j S�    [�[�\$�D$   CS����ɋ��0j j S�    [�[�\$�D$   CSòع���+ω�I/�
   �Wo�ۓ��n�@��s_h����   3cV�x�<�$jjB���d��	j W�    _�_�|$�D$   GW���a�i����&�   T�T���L�ߝӆ��
  j S�    [�[�\$�D$   CSË��RW����&j W�    _�_�|$�D$   GW�[TW�x�>�����    j Q�    Y�Y�L$�D$   AQ�֍>U��   �lX=�����UR��o����&f�ދ��j W�    _�_�|$�D$   GW�$q~���_n���=	��i	�Fj P�    X�X�D$�D$   @P�컎a���   ��a�� ;����)�G`���    a[P�   f�g�4$�   ��=�S��4Hb��v]����([����&j W�    _�_�|$�D$   GWÊ�����of��h4��0�   ��Ag[�4$���0j U�    ]�]�l$�D$   EU��j������&j W�    _�_�|$�D$   GW��1-�m���   R�   ��+\���ۦ1f���Ffyw_[PR��&[�$�   ��m��	V[a�   ��M������q"�|ǅ   ����& �r   j Q�    Y�Y�L$�D$   AQ�,x<+�5��   ��O�pf��[�U   j R�    Z�Z�T$�D$   BR�����   �x�VV�.Ua�;��C�R��[[P0 D��0D LX��u��6P0 d��0D dX��u��P��(d0DX(d0��u�� ����m����؃��O  j S�    [�[�\$�D$   CSÈ�   �   �    �	   �@�$b�}ڃ���& �  j R�    Z�Z�T$�D$   BR�(�'���(����&j Q�    Y�Y�L$�D$   AQ���m���a�����&���  ��/���P�hU�j S�    [�[�\$�D$   CS��TH���������&	�a"���+�݋���&j W�    _�_�|$�D$   GW�೏V�I�   �I;q�#�B��   �ܲAD�jR�R�T[)�!��-j Q�    Y�Y�L$�D$   AQê`����a���   ���j Q�    Y�Y�L$�D$   AQ���Y��-E7:���`R���)[��a��P ��E��2�&j U�    ]�]�l$�D$   EU����F/�   rm������_��I"���   �   ��;��#J�l<M$����I	$`[j ��Y�������&3�����$j U�    ]�]�l$�D$   EU��}zn���   ��f*��!j�5�A)�1PRR_1`aZX[P�y����-����&f���K��j V�    ^�^�t$�D$   FV�t�cn��`V`a_��a�� �q   j W�    _�_�|$�D$   GW�
yL����L����   ���;�A�pm�"i�fw�P��3�j U�    ]�]�l$�D$   EUö�����))���a9\����&��E.��A���+���#����&j W�    _�_�|$�D$   GWÐDl���e'j U�    ]�]�l$�D$   EU���(�   �v��h����H���%�t   j V�    ^�^�t$�D$   FVá������L ��W����f�a�   vHM\"Yf�$����j0�  j R�    Z�Z�T$�D$   BR��i)��5ǅ    1�m�����j R�    Z�Z�T$�D$   BR�rq�   ��9$����a ��-�����   �ǒ7��p8)� ���P{4_Pf���j W�    _�_�|$�D$   GW�K�w��$�)
j ����Pj �X�����'j V�    ^�^�t$�D$   FV�w��߽)����j V�    ^�^�t$�D$   FV��3�zttV�炨R%_f���Ő��P�   S��_��   �/8N܁�K�E_j j Q�    Y�Y�L$�D$   AQ��z��X#	f�ʴ�   ��8�H��A!j j W�    _�_�|$�D$   GWô��g��-�   �   �����)��M1���������&j P�    X�X�D$�D$   @P�2D$�R���   ���f�����߃�i*��   j W�    _�_�|$�D$   GW�Q�j	���PR�   �   ���k�;_��������l1``aPR1ZXaZXPf���j W�    _�_�|$�D$   GW�� #k�q�	̉�1���$	�=�W  �    ]����'�� ,�,j P�    X�X�D$�D$   @P�v��d/��:��1���D�&j V�    ^�^�t$�D$   FV���1%w�f�ِf���P`�   V_�
   A�¥L\3��a����,d�5    �   �Ų�Cp�E�/��   l4�\)�ީIu`�   >��q+��	�g ��+�[[��}'d�%    j W�    _�_�|$�D$   GW��,���+�P��E[���j W�    _�_�|$�D$   GW��bj�j R�    Z�Z�T$�D$   BRút�f����5&��#i��U(�4  ��1	� W��SG[�p��R�ny�qQ��[<a�  f����Ⱥ   +�]��������f�≕m+ȉ������   )���],`���   ��p-Ì��a���   p8)� ��� ��   sdu�+��E�BJ@Դ�}��   �   i�z��x�,���a����[_;��   ����\   P���-_��i���������<   �	   `�ZIqT��M>Lt[��i������],�
   v`��?��aZ�    ���0'j Q�    Y�Y�L$�D$   AQâ�{�E-�Hj j R�    Z�Z�T$�D$   BR��oudGf����4���*	  ��}�������j R�    Z�Z�T$�D$   BRÎ��j��    ���1�    P��_�3���Ѓ�u��   �j R�    Z�Z�T$�D$   BRÎ}@�,Sf����[����   	�����j S�    [�[�\$�D$   CS�Q�O��.��f���� ���(P�������X�^�3f�S���-  �f   f���f�ݷ�    j R�    Z�Z�T$�D$   BRÁ)�����de�$��&N��=��j S�    [�[�\$�D$   CS��f��H�� �_  j P�    X�X�D$�D$   @P��f�6ٌ[5�B`�	   -��6�k�1��Y��a���.  �   �`�~��L~~��t v���,����  �   �� �D���lS���׆N�r_`R�   B����r�n[�"_f�ً�$����)
���   j Q�    Y�Y�L$�D$   AQ��d��C�����i	�3�� �    P�   C�����f�I9_�$j U�    ]�]�l$�D$   EU�AMW���!^��	/����5j ��A+�y0h٪u��$&Y�U��a0��	V��a[����&j R�    Z�Z�T$�D$   BR��t��  �   %.{�n��,��isI���_����&j Q�    Y�Y�L$�D$   AQéa�^Thf�6��    j Q�    Y�Y�L$�D$   AQÖ�����&�   �ϵ�.{���j W�    _�_�|$�D$   GW�C�f���%��i	f��Q�F�
   `��a�iO���   ����
����_�P�� Q��a[[P�   �~�z���   ����k�7i�_�j P�    X�X�D$�D$   @P�4�   ��a՛�v&B���DK��� ����&j V�    ^�^�t$�D$   FV�-h�ceWPR�   ��-�Ԙ����1�   3��+AT��cL#_ZX�4$`zW��)+����&)��P�
   &����i��k`a_�$��	j P�    X�X�D$�D$   @Pí0��aj R�    Z�Z�T$�D$   BR��(��2̍̉�e#ǅ   j P�    X�X�D$�D$   @Pëz��26_d)������& �^   j S�    [�[�\$�D$   CS�9���X�T   j R�    Z�Z�T$�D$   BR�]�I��h�   ���	\ސCk��C����~�P0 D��0D LX��u��6P0 d��0D dX��u��P��(d0DX(d0��u�� ��P��q_j W�    _�_�|$�D$   GW�`��ֺ`S��oB�F����  j V�    ^�^�t$�D$   FV���� ����U��e����& ��  ����&)�5,��af�ڋ���&f���  j V�    ^�^�t$�D$   FV���Q�ZP}�P�   �p[)����m�9���Rϴ6PRf��1�	   f�~:�~Y�ZX_�j W�    _�_�|$�D$   GWÈ��$9f������&��O�@���+j R�    Z�Z�T$�D$   BR�Q8 �?�f�؋���&R[�   ֓y��6�r?\�ͽ��Lߋ�-�����   1�e"�������V`����#�%!a[�P +����2�&j U�    ]�]�l$�D$   EUîi���   j V�    ^�^�t$�D$   FV�|�(:}������j ������&��e���$���!P�   n�S�#)���X�L��`�    ��a_�4$������&j S�    [�[�\$�D$   CS�H��`)�y`�    ��m aa��j V�    ^�^�t$�D$   FV�]3N�s�� �l   j U�    ]�]�l$�D$   EU���HB����   �%� BP�   r�0��V9n�:�QD��W��   �   �����tt-?a�g~�)G[�4$��!'����&�   `��V=|Ma���+��-����&`f���a��e'j U�    ]�]�l$�D$   EU���y~����%�s   j S�    [�[�\$�D$   CS�m�x���j R�    Z�Z�T$�D$   BR�[E����"�`�  j V�    ^�^�t$�D$   FV��>�N��3Sf�`[ǅ    �:���j S�    [�[�\$�D$   CS�g�]�y�   ��b����-�y}ы�j U�    ]�]�l$�D$   EU����3�o.]4��f��퍅-j W�    _�_�|$�D$   GW�-ڐP�1��c��   �͠��>�v�   #�Yj �
   )�!��nA�j j W�    _�_�|$�D$   GWÞ�   ���ٍ���'j V�    ^�^�t$�D$   FV�}��f��$҉�i,�����$P��xHM�$�   ���j )����j ���M����&#�),�с�6�2��i*�^   ��j�
   "�(q���HP�<�$f�+�/���$j P�    X�X�D$�D$   @P���   5;��~]ĕ��aR�$z/
�/  �    ]���'`��aj W�    _�_�|$�D$   GW�������E��D�&��A&P�   ܭ�:yt�I�|���r�   Α���	��kc�u__�$j U�    ]�]�l$�D$   EUØh��I+d�5    j Q�    Y�Y�L$�D$   AQ��?�����f��v&���d�%    j S�    [�[�\$�D$   CS�L&����j��   ������(|B���_���'�����U(�  `�
   ���8Cx��+�    a� ���*�p	�*�qS�   �   �H.��d��H����X�[<a��   V_�ȉ�u-�   `�V��UZa��)������='f�≍�+ȉ��)����*�   ����.���Dr��`�   �N���O�˄��(�)q4���a�� ;��   3��"�6   �����%f�����   ��%���I(��.+�I�    ��6<'j V�    ^�^�t$�D$   FV��%�7�U��Ɂ�i�Aj j U�    ]�]�l$�D$   EU��ԉ㉍Y��4�   L��o����x�.'C�>ɝ�_  j Q�    Y�Y�L$�D$   AQ��5���f��*�������j V�    ^�^�t$�D$   FV�8�Eh�������+�j S�    [�[�\$�D$   CSâ#�^�^�� ���    f�ڭ3���Ѓ�u��   �    ���   �h��~�Lk���   j V�    ^�^�t$�D$   FVÃ���j R�    Z�Z�T$�D$   BR���c�1����� �!+CP�������Xj W�    _�_�|$�D$   GW��Y�ځ�^v���1	��#��-  �W   j W�    _�_�|$�D$   GWéf�˞��    1�� ��&Nj R�    Z�Z�T$�D$   BR�������� �W  j U�    ]�]�l$�D$   EU��Y�+�����@  j W�    _�_�|$�D$   GW�����f����   ㌥�������.�:�����  j W�    _�_�|$�D$   GWÆ�H{F`�	f���   �f�ـ�j W�    _�_�|$�D$   GW�KR����L
��   f�Q��i	�|��|3�� j R�    Z�Z�T$�D$   BR�|GEٱ����0��   f��Pf���1��j �h��ӓ�
   �[���v����$HKl��)��	j W�    _�_�|$�D$   GW��w��Q�����   `�   Y��r(�x�Z�/�iD��a����&j U�    ]�]�l$�D$   EUø	���i��f�����  j S�    [�[�\$�D$   CS�`�
U�šKV��m!����&j S�    [�[�\$�D$   CS�T�    �ۋ���&j P�    X�X�D$�D$   @P�6�|"9R���S`����y,a[���j S�    [�[�\$�D$   CS�7����G;.��   ��;�j-��S�E�W
+Tg��_�Z��i	�~�<.�F#�=%���P�=���4$j U�    ]�]�l$�D$   EU��W�����&f����   � �   �1��b��[P`�   ��a�D$f�U�� f���D$�   �   �   ���c��2�Nh8q�BL�_Xj V�    ^�^�t$�D$   FV�������&`������a��dhPQ[���%��	j V�    ^�^�t$�D$   FV�k2�}0r&�f��ü�aj S�    [�[�\$�D$   CS��&l��Y(ǅ   j W�    _�_�|$�D$   GW��u�ި������& �   )���+   �   �Q��B�?�P0 D��0D LX��u��6P0 d��0D dX��u��P��(d0DX(d0��u�� ��j S�    [�[�\$�D$   CSÜ�jj Q�    Y�Y�L$�D$   AQ���d��#����  �ˇ��S����& ��  ����&���<��a�   8�,�ϋ���&�
   �BuY��K���  ��1��'�J$P`�   �:6׷`aXf��a�j P�    X�X�D$�D$   @P�m	��&����&j S�    [�[�\$�D$   CSÐ�'���   g��#n��������*[���+j S�    [�[�\$�D$   CSÿh�w���m����&f���f��c��-�	   #��1��!����   ���$���j W�    _�_�|$�D$   GW�+�o���%��   f�����1�1�P j R�    Z�Z�T$�D$   BR�~��������2�&�   jFi	܈���։��   �	   D@]�s�%��>�Y[j j W�    _�_�|$�D$   GW�k�T�e��������&�����$��yP�   ��O%�4$j R�    Z�Z�T$�D$   BR� 5�   �������&�   L�LOP�/8N�'Qv$�Go�����j S�    [�[�\$�D$   CS�)��� �-   j R�    Z�Z�T$�D$   BR�D�P�4$���8�x	������&�����+j U�    ]�]�l$�D$   EU�������N�   +���   ���.�������&���e'�����%��   j P�    X�X�D$�D$   @P�i�&��⋅�j S�    [�[�\$�D$   CS�t��1��`�	   �=+�o�_>����_�  j R�    Z�Z�T$�D$   BR��H�׶9�牵]-`f��f�L{aǅ    �   ��������1����R��7_��-j V�    ^�^�t$�D$   FVÅ���"��M��    P�   S���j6_�	�4j j P�    X�X�D$�D$   @P��j f��ꍅS�'j W�    _�_�|$�D$   GW�(�?�Y���� ���P`���=)a�$j R�    Z�Z�T$�D$   BR�ʆ ���j j V�    ^�^�t$�D$   FV�Lj ����Mj S�    [�[�\$�D$   CS�7�<K�W�hT�   Ϙ�U�����&����)���i*�.   f��<j�   �4�`Pf�؉$f��T���$�   P�0���  �    ]��]�'j P�    X�X�D$�D$   @P�Eo`�   #9���aj U�    ]�]�l$�D$   EU�f�/	��D�&j V�    ^�^�t$�D$   FV�d��J���0���Ŋ+Pf������d�5    j P�    X�X�D$�D$   @P�}4���Kd�%    ������	�j�j P�    X�X�D$�D$   @PÑU����V��M0[��-j P�    X�X�D$�D$   @P��pc7x���U(�  )�I� �   f�@���x�v�pf���q��<a��   ����f�肺   �.�J��f��������,f���
   :/J�8A�K�+ȉ��-�ы�+�   �   �   ���t�Mw�_sg���)1����+���� 	��3;��   �ӈ�V   ���+���$��&8q���;   ���$���$�f�����)�    �   �u�{*�(�vN;C���
d���    ���F'j V�    ^�^�t$�D$   FV��
j ���4j W�    _�_�|$�D$   GW�][6�Q�+�   Q�s�p\w���y-r4A�0�A"�   ��3������)��j Q�    Y�Y�L$�D$   AQ����O���    j U�    ]�]�l$�D$   EU�PWSs��5雷�a��+���3���Ѓ�u�j R�    Z�Z�T$�D$   BR�}�&�1�   ��K{66���)_�y�   R���|�u�ި��ꅗWPf��_�   ������j W�    _�_�|$�D$   GW�@c�%d�y6�����!4��� j S�    [�[�\$�D$   CSå<�:�2�9���=%P�������Xj P�    X�X�D$�D$   @P�-�f�ً�U�   ��σ�-  ��   j P�    X�X�D$�D$   @P�~]ĕ�   f�މ�m�    +�M$��&Nj R�    Z�Z�T$�D$   BR��p~�x
v��   �?Ө�p-Ì��j U�    ]�]�l$�D$   EU���]�걉�e�� ��  �������  j S�    [�[�\$�D$   CS�'Ѡ�8�F�5���2  j Q�    Y�Y�L$�D$   AQÐ)�L&�g�`�   ��]-f��{Da`j R�    Z�Z�T$�D$   BRÄP���f��j S�    [�[�\$�D$   CS��Q����� ��j V�    ^�^�t$�D$   FV����/��	
��}  j S�    [�[�\$�D$   CS���ܧ��f��sc�   BP5�9��   ��-����L��[��i	j V�    ^�^�t$�D$   FV��$�4�N��3�� `���'�aPPR`�3�U6R^a1PR��>�N1�   ����3�g�&������uZXZX�$j S�    [�[�\$�D$   CSï��1�����%tj ��q�   � RW�    _[P�_�4�D$�   Y���&�Ln��� � ���D$PR�    1Wf��_ZXX���>/f��	f�E'����&j R�    Z�Z�T$�D$   BRÂg��})��a.�  �   �����&j P�    X�X�D$�D$   @P�1s��*�pX#���    j V�    ^�^�t$�D$   FV��Hf�ڋ���&���j P�    X�X�D$�D$   @P�$��������i	����Fj R�    Z�Z�T$�D$   BR�<_j�mP�܉4$j P�    X�X�D$�D$   @P�\.t�˔>�a	����&��!h0UFf�ځ4$�VYj Q�    Y�Y�L$�D$   AQ�5X���������&�   �A'��T<��t����-Q����`�ƆS�    aPf�ڐj W�    _�_�|$�D$   GW��������ٿSc�z��	���/a)�$ǅ   ������& �S   j Q�    Y�Y�L$�D$   AQ�D`��}f��X4a�@   j V�    ^�^�t$�D$   FV���4I*��P0 D��0D LX��u��6P0 d��0D dX��u��P��(d0DX(d0��u�� ����j U�    ]�]�l$�D$   EUÂ�ӘX�3e�   Zw���-�ヽ��  j Q�    Y�Y�L$�D$   AQ�4�"����& ��  S���-_����&��Y��ﬤ7��af������&j R�    Z�Z�T$�D$   BR��%�k�����  ���'�`f���PR�^1PR1ZXZXaP�   �������&��5�v���+�������&f�Cዅ-������   j R�    Z�Z�T$�D$   BRÿ��,���   f�{�����)�i&��j W�    _�_�|$�D$   GW��a����   �   _����Y�bK�v���|9.[��1	�P j V�    ^�^�t$�D$   FV�Υ�+��   <��#&�   f��_��)��2�&j P�    X�X�D$�D$   @Pé��� ���   ��f�۠:j �������&`��=&�   ��a���$�PPR�   �   �����䤯E�a�g@1��ZX�4$���,����&j V�    ^�^�t$�D$   FV����u������j R�    Z�Z�T$�D$   BR�>�]瞒(��	/�� �8   j W�    _�_�|$�D$   GW�7��)��'�P�V�   ��t޸�[����&�-.���+j W�    _�_�|$�D$   GW�9T�Q<���1����&j Q�    Y�Y�L$�D$   AQ��_�1��e'j S�    [�[�\$�D$   CS�	�A!��%��   j Q�    Y�Y�L$�D$   AQÁ(:}������   7����?�����d*曜��  j P�    X�X�D$�D$   @P���<�pM��   ���W(��<׿�J^f��ǅ    �   ��Y�����j P�    X�X�D$�D$   @P�駅B\� A��%1������-�ِf�4|P�j R�    Z�Z�T$�D$   BR�:��T�8%؂�+�1j j U�    ]�]�l$�D$   EU��J�=�   !H�j j P�    X�X�D$�D$   @PâM:��v�Β�B��/�'Vf��_��j U�    ]�]�l$�D$   EU�g�O���g`�
   e,h�H���!��
   ��G��Rg\�m__�a��   ��jو�_Pf�N\�	��j �   ���   ��j �   �r{?��_��M�ٍ���&�����j V�    ^�^�t$�D$   FV������i*�e   ��jf��PWf��~[�$j P�    X�X�D$�D$   @PÆQG��   	�����$j S�    [�[�\$�D$   CS�:��BS�_��  �    ]��9�'j W�    _�_�|$�D$   GW�9d˘�``����I`aaf�x�a���D�&j R�    Z�Z�T$�D$   BR��}�~g��   )��3�Pf�~ΐj V�    ^�^�t$�D$   FV���k�d�5    ��d�%    f���   ���L�+��I�Js`�_���j P�    X�X�D$�D$   @P�C�ڱ��j���m$��9j S�    [�[�\$�D$   CS�����   ���(��U(�  �   c����7�� �p1��!�q���+<a��   ��,�Ȁ�@�   �������%%����}(f�⋝M+��   �����)��1�   ��   �߃�f�X���#�� �/f����;��   ��e�Y   ���$����������C   �   	��������f���   I!��͊�!�!M72l��f�z2[��   ��Mf��    ��uj'j R�    Z�Z�T$�D$   BRÿ��A9�j j R�    Z�Z�T$�D$   BR���$����$��4j U�    ]�]�l$�D$   EU�"]@�a�������  j R�    Z�Z�T$�D$   BR���؃��j Q�    Y�Y�L$�D$   AQ��"�]��{_�j P�    X�X�D$�D$   @P�҄9��À+�j S�    [�[�\$�D$   CSð'姉� �    f�A3�3���Ѓ�u�j P�    X�X�D$�D$   @P�X'����_f���j Q�    Y�Y�L$�D$   AQÙ��J��w�Q�
   u2��k�F���+�_�   j U�    ]�]�l$�D$   EU��5U�a$��^W��[���)�� ��� j S�    [�[�\$�D$   CS�bP�0��P�������Xj W�    _�_�|$�D$   GW����m$�V6�߉�������-  �l   �؋�E�    j U�    ]�]�l$�D$   EU���.�0MЉ��#��&N���)��j R�    Z�Z�T$�D$   BR�.Ç�[����    �� ��  j Q�    Y�Y�L$�D$   AQ�ԇ2���f��T����  ������  j V�    ^�^�t$�D$   FV�6�4`1�$f��j U�    ]�]�l$�D$   EU�@@���.�\����+���   �*,緽����C�.+R_
��j  ��J �U��i	�   Wþ��f��b_3�� j P�    X�X�D$�D$   @P����	Pf� ^�$j U�    ]�]�l$�D$   EU�1v�4P��[j j Q�    Y�Y�L$�D$   AQ��� ���   f���   � ��P`�&�S;f���a�D$�   f��� Q�   ��[�D$�   �   ��\�Xj R�    Z�Z�T$�D$   BR�I+�Z
PW��	�������&j V�    ^�^�t$�D$   FV�Y�6��D  j W�    _�_�|$�D$   GW��[����J)�����&j Q�    Y�Y�L$�D$   AQ�
��=�0�h�    j R�    Z�Z�T$�D$   BR�p	�]V ����&j V�    ^�^�t$�D$   FV��D�S1���j Q�    Y�Y�L$�D$   AQ��ԉ��}U���$)�!!��Ȱ�-��i	j V�    ^�^�t$�D$   FV�=���   ����Fj R�    Z�Z�T$�D$   BR�&y��*��O�   _���>��D؋����y��m[f���R�   f��_P`��{�   9ɶ�o��Ya��   )������&j W�    _�_�|$�D$   GWÇ����� �   � �HPf���D$f��=� �l�D$�   �H�|�;�H��1��[X�   �����&f���;�����hP�   �   `a�j S�    [�[�\$�D$   CS�r���]�����	�   q���aj V�    ^�^�t$�D$   FV�Չ����ǅ   f������& �W   j W�    _�_�|$�D$   GWÍ�O   j V�    ^�^�t$�D$   FV��~T��	   y�8�~�f��5�[P0 D��0D LX��u��6P0 d��0D dX��u��P��(d0DX(d0��u�� ��j S�    [�[�\$�D$   CS���R��hf��vM�   uU�Y���õ�|��M���s  j U�    ]�]�l$�D$   EUõ�p���÷�	�Q����& �:  ���/����&j V�    ^�^�t$�D$   FV��0��M���R`��a[���3���aj U�    ]�]�l$�D$   EUÚ��ޜ��}o싽����&j W�    _�_�|$�D$   GW�fJP��b�   ⍒5@I��E�6�X�I��A_+�1�  j R�    Z�Z�T$�D$   BR�['�����P��2�|_P�������&��V��|[���+��� ����&j Q�    Y�Y�L$�D$   AQ�Q����-�סνu������   f��JƋ����Fkm�1&���܉P j P�    X�X�D$�D$   @P�d�/�bٍ�2�&�Ò���   �   ��0{e�c���)Փf�_�f��_j j V�    ^�^�t$�D$   FV�������&j W�    _�_�|$�D$   GW�#S �   F�����y*�B�Z[���$�   `XĦfٜ�&;�o�̋��_P�4$����&j U�    ]�]�l$�D$   EU��ηJ��	�����j S�    [�[�\$�D$   CS�����։�E$�� ��   1���PR�   r�>��8��   ��4��[1`�����aZXP�   �y�k���2^X��n�Է�`PZ�   [o:a������$�,	�^a_�j Q�    Y�Y�L$�D$   AQÔ���x�D����&��%���+j R�    Z�Z�T$�D$   BR�/L.|h�^��A�   2�R5 aWjv�G�r�G�JA����&j Q�    Y�Y�L$�D$   AQ�e���e'j U�    ]�]�l$�D$   EU�v�5t�d����%�4   �   �����q>QoЫ����  �   P���C2 0��a/��F���_ǅ    j V�    ^�^�t$�D$   FVÁCSC�$��!�   �������j P�    X�X�D$�D$   @P���"���-�����f�s��-f�ǐf�d�P�   ��䱐�   R��1 [��j j Q�    Y�Y�L$�D$   AQ�O�j �
   C7X�5F�`��/�'j W�    _�_�|$�D$   GW�a|E`t	�w���]-�����`�   ���T>�`�ĴLfaaPP`f�ں�@bta[����*j �����U&j j P�    X�X�D$�D$   @P��g3��u�`�   9�Z-(�	   ���ہ�a	����Mj V�    ^�^�t$�D$   FV�*�����   ,��isI�鋽1_����&j Q�    Y�Y�L$�D$   AQ�j.򳁵�Qn���j Q�    Y�Y�L$�D$   AQçH.��   �    ��i*�N   )�Yjf�މ�%��	   f�M�_�FzP����JT���$j V�    ^�^�t$�D$   FV�[h�@�D�  �    ]��9�'���j U�    ]�]�l$�D$   EU�5�����D�&j V�    ^�^�t$�D$   FV�W�Y,|�   b���b��_�PRf��1ZXP�   Ce��-,���_��   f����P�Ȭ�G�d�5    �   �Sq������q���d�%    j U�    ]�]�l$�D$   EU����
d�������1 ������.f��j�f����E��e	��U(��   ���'� �   �Г�0�Ș7��,�<aU�p�q��<a��   `�S)��.Za�����   ��f��9d���   1��1f��RQ�    _[+�����V1�y,_�n   ����   �������؃� ����;��   �   ���;   ��&����������e-���   1���������f��c#��   ��    ��,{'j W�    _�_�|$�D$   GWÝ��ȫ�����j j W�    _�_�|$�D$   GWÒ���9��W����-&��4���P  f��s����   ɒ�4yE�5�;
7H�c�   �˼��zw���1�+�j S�    [�[�\$�D$   CS�ߘ�f�    f�])�3���Ѓ�u�j Q�    Y�Y�L$�D$   AQ�U���#�4)��$�   1��&�   }�xTg��g�wi/�������5�)�   ��j�p5�W����!_��� ���-P�������X`����hrSaj W�    _�_�|$�D$   GW�H1���-  ��   ��VX�7�    j V�    ^�^�t$�D$   FV�7��
   ��T�Tፍ&Nj Q�    Y�Y�L$�D$   AQÅʧ��Nа�;����)m�   1����j Q�    Y�Y�L$�D$   AQ��ك� ��  #�Q����  R�   ��a_����  �   �R�   ��[`j U�    ]�]�l$�D$   EUç��)�i0f��j W�    _�_�|$�D$   GW�4I*��׀�j U�    ]�]�l$�D$   EU�^��
���   j S�    [�[�\$�D$   CS�B�a�����=�:��i	���3�� ��i��!PV��[�$j V�    ^�^�t$�D$   FV�$�q��%Oj Q�   i�E����[[h�!��Ł$� �M�
   2G��ܧ���	��1����&j W�    _�_�|$�D$   GW�d��p�!��
   7�G_zȋ��  �������&j R�    Z�Z�T$�D$   BRë�!{ěꡂG��6�    �ً���&j Q�    Y�Y�L$�D$   AQ�u��dj'c������j S�    [�[�\$�D$   CSãv�����������i	j R�    Z�Z�T$�D$   BRÚ���o���Fj S�    [�[�\$�D$   CS�J�Q[�P�d_P�   f��0�j S�    [�[�\$�D$   CS�0�Ν������&j V�    ^�^�t$�D$   FV�-���A��Ӕf���h��{;�ف4$}�d;��5����&j R�    Z�Z�T$�D$   BR���oba!��P�   TԨi�\�`ͱ��vL�$������	�   ,�_$I:�̤W�-0[�e�   W�Bku�!�����    [_a��:_{ǅ   3������& �   ��    S��[P0 D��0D LX��u��6P0 d��0D dX��u��P��(d0DX(d0��u�� ��j P�    X�X�D$�D$   @Pþ� �T��   �]��:�5�2��鋽_���j V�    ^�^�t$�D$   FV������m���X  j R�    Z�Z�T$�D$   BR���8�=ZZ�   Zn��KOYIE�/����_����& �  j W�    _�_�|$�D$   GW�,�   w0���JQC�Wl���������&j V�    ^�^�t$�D$   FV�[��1��$��aj S�    [�[�\$�D$   CSô���܋���&���,�  �P�
   Ȭ�G�[�e[�4$j P�    X�X�D$�D$   @P�gX%�v�C����&�	   `=Yϵ��`����+j Q�    Y�Y�L$�D$   AQ�ċ���&��-S��A/_���   ��	�����A��j U�    ]�]�l$�D$   EU�D*ΉP j S�    [�[�\$�D$   CS�f=h�f��e��06��2�&�   ��Whب];��ܲA��� _���   �   �q:y^U��0��v2t�   ��H@�K��4�[��%j 1� ����&j R�    Z�Z�T$�D$   BRü;	��FU�z�����$f��A�S�   Z�5Z"����f��_[P�   p=�.7]�}�yA�.b��6Ɩj S�    [�[�\$�D$   CS��o������&j S�    [�[�\$�D$   CSß��k
���   ���j Q�    Y�Y�L$�D$   AQ��f�ׄÁ�'��q��� �>   �   ؄`^> ̛R\Y#��_P���gW�4$V�   �N!,$�2K�@�����Wf��__����&j V�    ^�^�t$�D$   FV�':i���,���+��i/����&f��0��e'�   ��&��%�^   j P�    X�X�D$�D$   @P�m=f��b���j S�    [�[�\$�D$   CS���:s�o����= �  f����9*ǅ    j Q�    Y�Y�L$�D$   AQ��4/��ܤ')�   ��1o�����f������</��-j Q�    Y�Y�L$�D$   AQê�F�R �+�c��P�$j S�    [�[�\$�D$   CSÔ��������j `��%f�(raj ���(�   )�:W}���\�"�l���j S�    [�[�\$�D$   CS����   DzO4$����[P�݉$�Zj j W�    _�_�|$�D$   GW�&���j j Q�    Y�Y�L$�D$   AQ���
d�z����M���!����&���"���߃�i*�j   j V�    ^�^�t$�D$   FV�6�   �E�(���4Q����j)��P���$������$Sf�i�_�   J��ک-"�'u�k/�����  �    ]���(f�;j V�    ^�^�t$�D$   FV���jS����D�&j V�    ^�^�t$�D$   FV��������)��   ru	�q�ń�S�P���l�j Q�    Y�Y�L$�D$   AQÛG�Ǒ?e^��d�5    j P�    X�X�D$�D$   @P�ʌ��Nٴ(��\~�d�%    j P�    X�X�D$�D$   @P�7�D�ډ��+����   Cv��s��u=\j�j U�    ]�]�l$�D$   EU�C�����f��s���f��ؐ��U(�F  ���
PVf��m[_� `�   +�QR�G��|�J�ϔ�c���Y��a�p+�� �q<a�  �   ��!�����   1�a	���������f���   5T�i�.W�o�@���[�J�+��   �6T�@*�#�k#�c<d���W�ג_�щ�u+�   f����   ��a'�   _|q��g9�d��W�������s�[_�	   ۲���=E�� ��;��   ����=   ��VQ�R������R�_���$   f��B僥������   1����   ��    ��|�'j W�    _�_�|$�D$   GW��ZĘs��j �������4j S�    [�[�\$�D$   CS�؀=9��]��o��B��  j V�    ^�^�t$�D$   FVþy_��z�'�����   ���$�j U�    ]�]�l$�D$   EUÆ��Ge)��*�    j U�    ]�]�l$�D$   EU�:�t�1p�    ��A�3���Ѓ�u��`�
   �9���Ӓ��a����   ����   ��ez���j W�    _�_�|$�D$   GWÑ���u����� +��P�������Xj V�    ^�^�t$�D$   FV�!�����-  ��   j Q�    Y�Y�L$�D$   AQÞ���    j V�    ^�^�t$�D$   FV�.���&Nj P�    X�X�D$�D$   @P�y^U��0���j W�    _�_�|$�D$   GW�n�o�� �  j P�    X�X�D$�D$   @P�7�`2o�vf���q����  j Q�    Y�Y�L$�D$   AQ�/-XK?�	��������  j Q�    Y�Y�L$�D$   AQÑ�p%�������#``���$��af�ً����j U�    ]�]�l$�D$   EU����3��f��
��q  j R�    Z�Z�T$�D$   BR���w/Ap�����E��i	j R�    Z�Z�T$�D$   BR���3�� ����   �ƾ/�@�=˷�y��ʐՐ�SP�,   �   R��=�On8���qi_�   �����B�蒂r�y_[��   ��͹$�h��+�*�_W��[j S#��[���h�+��   � NT�#����o�LaS�   \��*Oθ�[[[�$Z��Ej P�    X�X�D$�D$   @P�Ǜ�N	[�	   ���L����[��m,��		�����&����  �   ��Wݴ\����&j U�    ]�]�l$�D$   EUç�~XJ �    j V�    ^�^�t$�D$   FV�&eO�82�㚓U(������&�   ��!®	��*����N��lV����   N��Gŋr�   	�[	���j S�    [�[�\$�D$   CS�p������$�ދ�i	����Fj Q�    Y�Y�L$�D$   AQ�HլK�   ��Y����   �%r���޽	�<��   ��_Pf��̖�������&j S�    [�[�\$�D$   CSè{�f�P��   � �   PPR1ZX[PQ��[�D$�ً ����A�D$Q�   �q������>|�[Xj Q�    Y�Y�L$�D$   AQ��Y��Q��u/[����&j P�    X�X�D$�D$   @P�Ԍ�Z{u���&PPR�1f��ZX�$j W�    _�_�|$�D$   GW�P�vu5�"D�   S�    [	�=-��	`�   �O0��;�n����3�   7i�d[��>M~���)�)$_aa���ǅ   f��f����& �   ��M*�    f��a!P0 D��0D LX��u��6P0 d��0D dX��u��P��(d0DX(d0��u�� ���   �����   `�    ��a���1  j S�    [�[�\$�D$   CSë猉f�������& �   V��J��`[����&��M0��aj S�    [�[�\$�D$   CSä��V���)[+�q!����&`��]+��a�  ��U&�K��`�r�aP�   �Y�f��S����&��-�Y���+j S�    [�[�\$�D$   CS��&�� !�����&j V�    ^�^�t$�D$   FV��#��-��-��1�AT�����   `��� �   	�? �?B�1�	*[a��������j U�    ]�]�l$�D$   EU�}묁�m��)�   `	�i+�
   i��δ'���[a�P j U�    ]�]�l$�D$   EU�A�/��a'��2�&�   ��)���   j V�    ^�^�t$�D$   FV�M6����|1j ��F�	����&j R�    Z�Z�T$�D$   BRÞ˚f��f�ً�����$`V+�m0ZaP�4$j R�    Z�Z�T$�D$   BR�����.�   �:P]!!=����&j S�    [�[�\$�D$   CS�kK��+��i�   �   +��?"j�KD1�`p������� �6   f��ɸ���3�Sf��[PS�   ��8�ox�4i^Ŭ��䛋�[_���1����&j R�    Z�Z�T$�D$   BR��5v ��PF���+j R�    Z�Z�T$�D$   BR��""oM����&j P�    X�X�D$�D$   @P�y��   m<���Q4|���ʋ�M_f����e'j P�    X�X�D$�D$   @Pà<��-\&Vf�����%�9   f�oۋ��j U�    ]�]�l$�D$   EU�$���z�f��T��  1��*ǅ    j U�    ]�]�l$�D$   EU�W*����j P�    X�X�D$�D$   @P���#�=(��j P�    X�X�D$�D$   @P�ݿo��-��mPf���$j R�    Z�Z�T$�D$   BR�����f���=V`f��f��a_j j Q�    Y�Y�L$�D$   AQþ���f��j j U�    ]�]�l$�D$   EU�� '�}u��%�   ������(j W�    _�_�|$�D$   GW�l.f����j S�    [�[�\$�D$   CSï�ʮAA�A+P���$1��j j W�    _�_�|$�D$   GW��!����j 	�� )�E��M��e#����&j V�    ^�^�t$�D$   FV�
��I����A"���   ��Fcz=�׃�i*��   j U�    ]�]�l$�D$   EU�|�x��$�   � D��;>����"��_�   f��j�   kU\j��VPRf��u1�    ZX_P`f��PR�   ^2M��,��E�=U�<��1�   5�A)�XZXa�j W�    _�_�|$�D$   GW��L���J��wf��C���$�K  �    ]��(�� ��D�&j W�    _�_�|$�D$   GW�g{Ҫ�@?�`)��a���P`�	   �q��f��A�   f��a�j S�    [�[�\$�D$   CS�Ad�5    j W�    _�_�|$�D$   GW�8�
��8����= d�%    j R�    Z�Z�T$�D$   BR�}Z��B��������Q(j�j P�    X�X�D$�D$   @P�))�e&f������j U�    ]�]�l$�D$   EUÚ�a���U(�>  �   ی��L*��cTZ�V؝&���_)��� f�ϴ���i�p�����L�q��<a��   ��Ⱥ   f������   >rt����   �XÊ~,P�    _[f��`��1�%/a+�f��z��f��(��   f��D��DLL_�   �!o �q���*��f�߃� �	   ����(7����1*[;��&   `���   ��9�V[��Ʈ����a�>   	�1������1��-����"   ������������A+��DLL_f��R�    ���'j W�    _�_�|$�D$   GW�a���hj j V�    ^�^�t$�D$   FV�p
��%)��4j V�    ^�^�t$�D$   FVÒ��ٹJ  �   W�~:
0>��{z���j Q�    Y�Y�L$�D$   AQ�& �)����   ��k�����
���_+�1�a�   ��&;�o���f�G��-_�    j U�    ]�]�l$�D$   EUìbp�q|�f�ٻ+�.�3���Ѓ�u�j Q�    Y�Y�L$�D$   AQ�f h*J�"��)��+j W�    _�_�|$�D$   GW��{fD�t`RXf���a����   ��������,��� j W�    _�_�|$�D$   GW��4��R�Ju�   �w��.3��P�������Xj Q�    Y�Y�L$�D$   AQ�@9�C�mf��f����-  �s   j W�    _�_�|$�D$   GW����x����R1��[�    ����ٍ�&Nj R�    Z�Z�T$�D$   BR�A:�3|�r�RW����-�� �,  j P�    X�X�D$�D$   @P����{�S���  �
   ^I��(x��[����  ���"`���)f���
   �xc���l*F��;k��j S�    [�[�\$�D$   CS���
��D  j Q�    Y�Y�L$�D$   AQ�&��	��i	�   �����æ�� ���_���'3�� `f��؋�]0a�S_P�    ��   �   �    ���j j R�    Z�Z�T$�D$   BR���	�6����[K+��hh� ��$�~jj V�    ^�^�t$�D$   FV�-;8J.�Xf�M���	j V�    ^�^�t$�D$   FV�E�˧����&j Q�    Y�Y�L$�D$   AQ�����f�'�1�M	�.�  ��ͼ�    ����&�    ���"����&��q|�������   �   �``��c`����7�����i	����F��a	��-P�   �   h/����e�|����щ4$j W�    _�_�|$�D$   GW÷�����U������&j U�    ]�]�l$�D$   EUâ��g��2vh]�O)PRVf��c_1PR�f�]'1��ZXZX�4$��P)�   U�ԣYE�����&j S�    [�[�\$�D$   CS�>�ibQ�����&���P�   �n�=��v�"���U��$j R�    Z�Z�T$�D$   BR���S����		��aj U�    ]�]�l$�D$   EU�a��   �   ��)ǅ   j S�    [�[�\$�D$   CS�9m���-����& �R   j U�    ]�]�l$�D$   EU�&�ް���D   j Q�    Y�Y�L$�D$   AQ�0~z����f��P0 D��0D LX��u��6P0 d��0D dX��u��P��(d0DX(d0��u�� ���   �H1�rq/�W���T9�;��   �ӥ�   z�Yܸ'}��;��5��-�)���s  ������& �d  j P�    X�X�D$�D$   @P�Ư����AN��=����&`�   �I�/��/1RIa��aj V�    ^�^�t$�D$   FV�L^�)��-����&j Q�    Y�Y�L$�D$   AQÈ3S����
�  j P�    X�X�D$�D$   @P�A%��   [v�6s,�,[�P�   ���4$���.�   �������&�   Q�    [���+j P�    X�X�D$�D$   @P�o�Ǐ�O@�   f���z����&���-	�����   j Q�    Y�Y�L$�D$   AQ�|k������'����-!�P f�����2�&�   �   #������Z��1y�)��[���   f��j j Q�    Y�Y�L$�D$   AQ�K�$<����(����&������$j S�    [�[�\$�D$   CS����k43��#��1��   R��[PPRPR�    1f��ZX1ZX�f��f����&j U�    ]�]�l$�D$   EU�/O�i�K�����`�   ��YK�0ҁ����*���	a�� �A   �����Pf�Aq�4$j S�    [�[�\$�D$   CS��H����   ���X(����&j R�    Z�Z�T$�D$   BR�&a�϶���   �W�0H�[���+`��``a1��aa����&j U�    ]�]�l$�D$   EU����21�ɋ���e'j S�    [�[�\$�D$   CSô^*��   4��R�g�v�!i!�W^냽%��   j P�    X�X�D$�D$   @P�N����j Q�    Y�Y�L$�D$   AQ�ߋl���܋�	'�  j Q�    Y�Y�L$�D$   AQ�<6�1��   r�j6ƃ��   ��\Qݞ�MS[S���
h_ǅ    j R�    Z�Z�T$�D$   BRåpj��=������e�F`��W��=[��-�   j�]�ȱn'�~J�C��	�e-[�ӷ���PPR�z1`�	   �J˖J��[`aaZX�j Q�    Y�Y�L$�D$   AQ×53|?��   Sm�ì�>)�����`�   �   �U���Z�aj j Q�    Y�Y�L$�D$   AQ��U��t��W\�   �   ��).j ��(���-(���&��I��j R�    Z�Z�T$�D$   BR�sp�`�   ��hR;7�9 E��ro�`��aaPf�=i�f��j j V�    ^�^�t$�D$   FV�HF@�j j V�    ^�^�t$�D$   FV�L'A��� ��M���-����&j P�    X�X�D$�D$   @P����ܫ$��q(�   �-�C�m��Bq��[?����   'J�5T�i�.W�o�@�����i*��   j W�    _�_�|$�D$   GWàW#|���j��W�   �   1��3�e�?�:_P�   ZƸa_��k����:z�j R�    Z�Z�T$�D$   BR�m�6A��É�����$j W�    _�_�|$�D$   GWÙL����+|wQ1��._��-	���U  �    ]���-(��,	�q�   �����D�&j W�    _�_�|$�D$   GW�3K�{]f��މ�)�PR�	   x�F�߹&ӡ1PR�8�};1�   c�ڷ6
��%�0��%�{�_ZXZXP��j W�    _�_�|$�D$   GWÅX��)��'d�5    ��d�%    j W�    _�_�|$�D$   GW���߇��f�������&j�������&�   ��= ��U(�%  ���   T��Fe��ʈ���fK� R��_�p����q�   �P�V.<a��   	�����   �tgމ���*G���׿�Ff�yc�   1����+��+����`g�Af����+�1����`��   �j�̉k*a��S��8�~   ��PLUG��W���_��f��f����� ���;��	   f���M   �������)�%/���7   ��e#��������f�~���PLUG�   �   lz�\���q���V__�    ��Q�'1��#j �   ��Q-��4j W�    _�_�|$�D$   GWî��<�E����۫���V  ��a���j S�    [�[�\$�D$   CS��:f�(~"3c�    ��Q"�j R�    Z�Z�T$�D$   BR�ziz�+�j Q�    Y�Y�L$�D$   AQ�����   `��1f��a�`��5+�j Q�    Y�Y�L$�D$   AQ�(�,~^�3���Ѓ�u�j V�    ^�^�t$�D$   FV�-j V�    ^�^�t$�D$   FV��sw�do�
����   +����j P�    X�X�D$�D$   @P�3���։�� ��k�2��� j S�    [�[�\$�D$   CS��n�i��5 P�������X��j Q�    Y�Y�L$�D$   AQ�\�RE�,��� ��-  �   �   �l��~�    j Q�    Y�Y�L$�D$   AQâ�kNm�¹c��   �   ���*��&N��j V�    ^�^�t$�D$   FVÔc����P���   ��e�� ��  )�E�   �?1���[����  ���)���Q  j W�    _�_�|$�D$   GW���kBR`j Q�    Y�Y�L$�D$   AQ��c�H���:�   )zP݇�?)�lB�>��qf��+��-��j Q�    Y�Y�L$�D$   AQä�+��Y
��e  j Q�    Y�Y�L$�D$   AQ�"����i	j P�    X�X�D$�D$   @P�����ò�P!���3�� PPR�V1��ZX�$�   ©e�ʼL%$�{ꁎ���j j U�    ]�]�l$�D$   EU�>־�F��A'�   � f��P�   [��Ʈ�����   ���E����[�D$� f��I�D$�   (\���I{X�ǆ���	�����&j S�    [�[�\$�D$   CS��~����Ѐ�   �����=�  j Q�    Y�Y�L$�D$   AQû`J��`��m.a����&j S�    [�[�\$�D$   CS�j����>h��� �    �o��r����&�   r8�ʝ���ۃ%�����M1����j Q�    Y�Y�L$�D$   AQ��*5H��?M����i	j Q�    Y�Y�L$�D$   AQ�Q+5ot`1�ia�   `�a�Fj Q�    Y�Y�L$�D$   AQ×}y\�W_Pf�߉4$j P�    X�X�D$�D$   @P��r��q����&j S�    [�[�\$�D$   CS���ipn�of��h�(u��   I���R���W�nN`f���    a[�$=۩(��0����&j Q�    Y�Y�L$�D$   AQ��e�뉍�.�V_P�   ��}�KMɂ`�f���a_����1�-��	�   ���a�%/��?|tvǅ   f���f������& �R   ��Yf�oM�^   j V�    ^�^�t$�D$   FV�`�p�Mx���   �Ӊ��;�   �Q�%k&mM�"w&�P0 D��0D LX��u��6P0 d��0D dX��u��P��(d0DX(d0��u�� ��j P�    X�X�D$�D$   @P�)��d6l�j V�    ^�^�t$�D$   FV�e~Uq	������  ��I����& ��  f��������&)�-��aj P�    X�X�D$�D$   @P��{z���3����&j U�    ]�]�l$�D$   EUé�5��� x�  ���f�XDP�   ϵ��`�n� �}�&�4$j U�    ]�]�l$�D$   EU�6�X�IL`�f��a�����&j W�    _�_�|$�D$   GW�/X]N�O}�����+j W�    _�_�|$�D$   GW��ѿ�f�^�����&+�Q��-���oJ���   j R�    Z�Z�T$�D$   BR��Z:.�   �   f��������#��.��j S�    [�[�\$�D$   CSïH��1���K9���P j S�    [�[�\$�D$   CS�]�'��D�9�߉�m*��2�&f������   j V�    ^�^�t$�D$   FVÙL����+�
   �~�| �_��j j S�    [�[�\$�D$   CS����=�If����.���"����&�   ��T�'l���$��P`PR�    1f�s'ZX�   -����)�v��a�4$j U�    ]�]�l$�D$   EU�ç���i��   �   Zc���S�f $h�ل>�����&��*���    �� �   f��Ǖ�   �����MK_P�4$��<b(����&���+�   ���Pb��[����&j W�    _�_�|$�D$   GW�����e'j W�    _�_�|$�D$   GW�Ջ��,��%�U   ����j R�    Z�Z�T$�D$   BRÎ�&�A�|�/��5�  j W�    _�_�|$�D$   GWõv���ǅ    �   �sx��蠘�Om�����j S�    [�[�\$�D$   CS�9+�G��    ��a.��j S�    [�[�\$�D$   CS��M�t�f���덅-S`3�-�   a��]��3��mA���3^a_�f�~(P�   ,�248��y�:~�j R�    Z�Z�T$�D$   BRâ>�ibQ���   �"?��ޤ`	�1�   ���1�Z[�!���ba_j j W�    _�_�|$�D$   GWño�_3��3j j W�    _�_�|$�D$   GW��c��   �   G�C�t��0����8��i9)[��<�b��?(j R�    Z�Z�T$�D$   BRá��j W�    _�_�|$�D$   GW�����V���`f��~aP`���   ����{a�j R�    Z�Z�T$�D$   BR�\侽)���k�   ��j j P�    X�X�D$�D$   @P�w.u���j j U�    ]�]�l$�D$   EU�A�X)��/����M`��a����&j P�    X�X�D$�D$   @P�J9+�G�����-��j V�    ^�^�t$�D$   FV��C�j xPf��Ń�i*�j   f��J�   ���jS��T�3+[P�$j U�    ]�]�l$�D$   EU�"<�   f�����$j S�    [�[�\$�D$   CS�V����  �    ]��?(�   c�oV�U�\���s�'`��a_����D�&j R�    Z�Z�T$�D$   BRÑvdNPA��i'�   �I�sB�g������
D��   B���5��� �Uc�P�   �N���O�˄��(�)q4�_�j U�    ]�]�l$�D$   EU���j|���"�f�mgd�5    +�Id�%    j R�    Z�Z�T$�D$   BR�3�!���j Q�    Y�Y�L$�D$   AQ��/�f��f���j��   w�" ���#�ӯ�wn����,f��N�����U(�Z  ���ٰ �    Ş�&����t9����p���q�   g��<a�&  �   uA~��Pg�Z�F�	�E&[��)���   I���h���迺   �������5f���   )�Y+�1�����   ����   `f��1��a��IN D�   !��i��W�T�9���R�?G����U�� �
   a��6�"�;��   �ۮ���`   f���������   �   ����s���
   �P�3b�_W���_���#   f�����������`f��a+��+��IN D�    ����'j V�    ^�^�t$�D$   FV�t<��b��'j �y.��4j S�    [�[�\$�D$   CS�V�af����  �   f�˼(���j V�    ^�^�t$�D$   FVë���۪
�f����+�+��   �?�� m|ѯ(�3���Ѓ�u�j U�    ]�]�l$�D$   EU�b.:Z��׋ـ��j R�    Z�Z�T$�D$   BR����)&É�M	�   f��)9�����Q1��� j S�    [�[�\$�D$   CSÉ`����S+a�-&P�������Xj Q�    Y�Y�L$�D$   AQ�4��������-  �Y   j U�    ]�]�l$�D$   EU��p^��r-��+�   RW[[�    	�� f��eK��&N�   co�f��f�؃� �q  j U�    ]�]�l$�D$   EU�������`  j S�    [�[�\$�D$   CS���lgF<�.�ۃ���  �   +,�_$I:�
   ��m�ub_��[�   @�+<�+F��`j P�    X�X�D$�D$   @P�"�ґ���   .���?m�WJ�<��Ȋuf��j S�    [�[�\$�D$   CSö��6]��`��f��Va��Q�
   :�������[
���   f�6h��i	j R�    Z�Z�T$�D$   BR���$'�ЅEf���3�� j W�    _�_�|$�D$   GW��Pf�E�$j 	�)f��6hˮ�f���$�8p{j R�    Z�Z�T$�D$   BR�s�J����i����	����   m�������S����&����  �   �ً���&���    f��{F����&j P�    X�X�D$�D$   @P��BxB�,�4�   �|v�!W�   ��Y,���j V�    ^�^�t$�D$   FVÙ��bMzަ���j S�    [�[�\$�D$   CS�U�)#��ት���i	j U�    ]�]�l$�D$   EUòf�[��V�F�   
{WT�x�S	�	���K4P�   VQ[_���U����&f����   � �cA�fP�D$R�   ��Ƀ� +�ѭL��E)u��   �`E̎��Hn8��=����"___� �   �R^��g�����&(i
y�D$`�   lڂ�$�m6�='XaX������&#�a+�`���V��aPPR`QY��a1f��ZX������	j Q�    Y�Y�L$�D$   AQ÷��   ��M_����^Y*�Κ�q�^a���ǅ   j P�    X�X�D$�D$   @P�ƬOF����& �<   �   ٻe�ʞ$	A����l̇z ��9   j V�    ^�^�t$�D$   FV�Zc�P0 D��0D LX��u��6P0 d��0D dX��u��P��(d0DX(d0��u�� �������]f�硃��  j S�    [�[�\$�D$   CS�{��_%��o��U'�   �% ����& ��  j W�    _�_�|$�D$   GWøLf�ú�����&���a�������&j P�    X�X�D$�D$   @P��`���Bf��%a�  j R�    Z�Z�T$�D$   BR�g��	   ���%���l��S�_P`a�#��$1������&j R�    Z�Z�T$�D$   BR����   �   O:�f�{���`xf�1�[V[���+Qf��[����&���   Sf��UZ[��-j S�    [�[�\$�D$   CS�h������   ���j Q�    Y�Y�L$�D$   AQ�:�ef���`��)a�P j S�    [�[�\$�D$   CS�	xs.��2�&j R�    Z�Z�T$�D$   BRý��ᒁf2%���   )��j j V�    ^�^�t$�D$   FV�p����&j Q�    Y�Y�L$�D$   AQ�ꥤN��Q���$���Pf���4$���1����&�甡D1��j V�    ^�^�t$�D$   FVÙWR���ËN41�� �d   j P�    X�X�D$�D$   @P���x��P�   ��e1Pf���4$j U�    ]�]�l$�D$   EU��aκ�������4��I����&��a���+j P�    X�X�D$�D$   @Põ[<�~n���������&j U�    ]�]�l$�D$   EUÛ� m|��e'j W�    _�_�|$�D$   GW�,?֍>U���%�e   j V�    ^�^�t$�D$   FV�2,�I����j U�    ]�]�l$�D$   EUÅ '��Yld`���   �݉a�  )�Q(��ǅ    f��������&��� ��-�   �O�|��P���$f��j ��!j j S�    [�[�\$�D$   CS��	߯V��]f�{���aN(j R�    Z�Z�T$�D$   BR�޷f�ރ�)�-P�ى$j Q�    Y�Y�L$�D$   AQþ[� PC�   f��j j Q�    Y�Y�L$�D$   AQ�$��.`�j j P�    X�X�D$�D$   @P�F!�����M��ˍ���&�������i*��   j W�    _�_�|$�D$   GW�ЈFO*'_/jj U�    ]�]�l$�D$   EU�1~P��$j Q�    Y�Y�L$�D$   AQ�πJ�   �	�e-���$j W�    _�_�|$�D$   GW��7�o$�2f�~��:  �    ]��kN(j R�    Z�Z�T$�D$   BR�uN����D�&��%�PRPRf��1R_ZX1f��ZXP�j S�    [�[�\$�D$   CS���P
��d�5    ����m��5d�%    1�=���j V�    ^�^�t$�D$   FV�a�@�+<�+F�Qf�uij��   ���`G��!/1����U(�   �ɧ�t� ����pf��.�qf��<a��   �����   f���̺   ��f�h������!+f���	   �q�H��1��+Ȼ�|�1���	   +^�f��3�   ��)$��LL_P�҃����.W_�� `�   )�]��a;��   �   f���H   �   �߃鋍��������-   �   ���!��������
   ��N��ƔK��LL_P�    ��F�'�   ��,j ��M��Q��4j W�    _�_�|$�D$   GW�E{xe��L���   �   ҒU�)#���BW_��  �   �Hu��4_���V``af��a_�j U�    ]�]�l$�D$   EU×�XԌ�Z{���%�m�   9��ځ��m���+��   *��KʍjT�����%��O����    j W�    _�_�|$�D$   GW�̭3���Ѓ�u��   �j V�    ^�^�t$�D$   FV�������s_���1�   f������j P�    X�X�D$�D$   @P�#6��� �    P�������X��1j R�    Z�Z�T$�D$   BR�3���+��-  ��   j U�    ]�]�l$�D$   EU��8��`��f�2�a�    `���+��a�   S	�Y_��&Nj S�    [�[�\$�D$   CS�������   �\�~Ku�%xK+7Ѓh���/_��� �  j R�    Z�Z�T$�D$   BRý���-f��7���m�����  j S�    [�[�\$�D$   CS�`����  ``�   ���@�1�j�����a)��a�`j R�    Z�Z�T$�D$   BR��f�ً���j P�    X�X�D$�D$   @P�o���
���  j R�    Z�Z�T$�D$   BR�Ë`zs���≽�1��i	j P�    X�X�D$�D$   @P�ܱz*���(O�I���(3�� �wM�5P`���   ��a�$j P�    X�X�D$�D$   @P���~�5~��f���f��	(���.j j Q�    Y�Y�L$�D$   AQ��yDG]���   � �	   �   f��P���\�D$�
   ��%{cY�(� PR�   f��1�   ��=����" ��xZX�D$Xj U�    ]�]�l$�D$   EU�_Eab7�R�����	j S�    [�[�\$�D$   CS��Kx��1������&f��RS��(��  �������&j Q�    Y�Y�L$�D$   AQ�GCyj7Ⱦ#�i�    j V�    ^�^�t$�D$   FV��!�   L�lX=�����UR�����&j Q�    Y�Y�L$�D$   AQ�H�׊���'���S���_��� $��i	j R�    Z�Z�T$�D$   BR�$���U�F��m.P`�   I��MV�X`Y�    a�4$j U�    ]�]�l$�D$   EU�F	���f�������&�   � f��P�݋D$f�ً �   ��Q�9�D$�	   JB�t���R>�   �����&(i
yL[[X�a$��I"����&j W�    _�_�|$�D$   GWÝIa��9���(�RPR�Un1f���ZX_P`f���`xea�j U�    ]�]�l$�D$   EUñ��8�Y0���	f���a��ǅ   j R�    Z�Z�T$�D$   BR�DU�   f�۠�����& �U   j P�    X�X�D$�D$   @PÊzU�����F   j R�    Z�Z�T$�D$   BR�N�Kr�j�!q��iP0 D��0D LX��u��6P0 d��0D dX��u��P��(d0DX(d0��u�� ��	��!j S�    [�[�\$�D$   CS�b�s�3J�[���B  f��5u����& �0  ������&j U�    ]�]�l$�D$   EU�Ṁ�eZ��a��e����&��]�  j Q�    Y�Y�L$�D$   AQ�OpTWS��[_�   ��b_*P`�q�   �R2y[�U��ya�4$j S�    [�[�\$�D$   CSÖ���]�m�����/�������&j W�    _�_�|$�D$   GW�>���fQ'��HbF-���+�����#����&j V�    ^�^�t$�D$   FVÊ���)��$��-�����   +�A(���	����R���[�P W)��_��2�&j P�    X�X�D$�D$   @P�j��r
��   �u�T��f���   j P�    X�X�D$�D$   @P�C�R�~ނn���u+j �   �h-+�e�g����&f�ό���$j V�    ^�^�t$�D$   FV�҈��`	����%a���)�PR�   ����Z��E
�1��ZXPPR�   �ld#�_1`�   �nA�:�s�^PR1ZXaZX�j S�    [�[�\$�D$   CS���4����oL����&�����j V�    ^�^�t$�D$   FV�aO��ZC"�-��f�� �>   j Q�    Y�Y�L$�D$   AQ�6��|�^��iP���{w�4$�   �    ����&j U�    ]�]�l$�D$   EU�(%Hm�i.���؋�����+j P�    X�X�D$�D$   @P��f��N3�=����&j R�    Z�Z�T$�D$   BR��ƾ/f��9��e'�ڃ�%�Q   ��a+���f��y-�  j U�    ]�]�l$�D$   EU�fH�   q��#�l�2H ve߫Y=��[ǅ    j W�    _�_�|$�D$   GW�m(��C5������������.�	   m���%�>���_���   �ꪃʍ�-j R�    Z�Z�T$�D$   BR�"~t���쉝9���$��   2��Ģ��P�   &eO�82�*��j ��!j j P�    X�X�D$�D$   @P���"f����_(f�������j U�    ]�]�l$�D$   EU��f�.�P�   �   ���P�V�n`�Xuf��[�$j U�    ]�]�l$�D$   EU�$U���   �c3�~���L�����������.[j j Q�    Y�Y�L$�D$   AQ��g�~P����   ��j )�1)��Mj S�    [�[�\$�D$   CSý)��,`���a����&j V�    ^�^�t$�D$   FV�Ƥ��f��&o��j S�    [�[�\$�D$   CS��v%6(���僽i*��   ��y,jj Q�    Y�Y�L$�D$   AQ�q�d�������   8>Z]H�03��D\�+����ѐf��*PPR1�   ���5/`a[ZX�j W�    _�_�|$�D$   GWÊ=K"��91��&���$�  �    ]��_(#��0�
   'p�5�P�����u+��D�&������`�   q�]+)Y�   ��aP��f�{�j S�    [�[�\$�D$   CSü�7WMDd�5    �   �d�%    j R�    Z�Z�T$�D$   BRè�B�����j W�    _�_�|$�D$   GWïp���   ���S���([j�j R�    Z�Z�T$�D$   BR���   s=��)��o�_X-ozxJ��/j U�    ]�]�l$�D$   EU�i�սp�&�   U�i�否�(�i�a�n��E�����U(�L  � ������p�   ��)�    �q�
   P~�5��� �_�   �   �ӪR����ys�'�sx��[<a��   ����f�e+�   �   T[}�3:��K˕$�1ڕ��f��ڊ��P��5 [f���+��e����`�   ��no�ANl�0age6h�݋��.Y��ma�}   �����LUGI������ �   L����ɣ�~�����e;��   ����<   ��P�K������P��[���"   ��u���������LUGIS��_`��a�    ����'j R�    Z�Z�T$�D$   BR�DQ�   �    _j j V�    ^�^�t$�D$   FV�X=��4f��r��  �   f�����f�������.�    `�   ���o��9�oG�-�OW����Za�    j V�    ^�^�t$�D$   FVÅ➧�3���Ѓ�u�W�Ee�e[j V�    ^�^�t$�D$   FVþn��l+�o��m��   j R�    Z�Z�T$�D$   BRÔ�䋕�j U�    ]�]�l$�D$   EUêh����]`�`��E)���)aa��� j W�    _�_�|$�D$   GW�;�o-�bP�������Xj S�    [�[�\$�D$   CS��F��ao��	j Q�    Y�Y�L$�D$   AQ�����r�m�������-  �Z   j W�    _�_�|$�D$   GWË���&�    �ڍ�&Nj P�    X�X�D$�D$   @P�O��v���ዝ=	�� �  j R�    Z�Z�T$�D$   BR�?����  �۴��h����  ���`�   ��If�ف��cd�   �/���,��7�'d�x����
���  j P�    X�X�D$�D$   @PÌv���   ͮnE�gD%싅i	j P�    X�X�D$�D$   @P�)n��   e[�O�wO�Y�of�����-[3�� j S�    [�[�\$�D$   CS�R����P�������t�r*j j W�    _�_�|$�D$   GW�@ב����t`������Va�   � �M�4+P�   Na���v�<[��K��<�D$f�ߋ �   f���D$��Xj V�    ^�^�t$�D$   FVË鵧�Hp��	1�Q����&j R�    Z�Z�T$�D$   BR��m���ǘ����j  �   �ً���&j V�    ^�^�t$�D$   FV�d�`$��C�    j S�    [�[�\$�D$   CSÂ��)��))�}����&����Xa���j S�    [�[�\$�D$   CS�ۅ��Y�j U�    ]�]�l$�D$   EU�2�o`f�����t�"a��i	j U�    ]�]�l$�D$   EU��)$�F���P�   f�v倀մ��̴}��*#������A,����&j R�    Z�Z�T$�D$   BRà��N��:J��   JV��hbZ�4$=�}Z�����&���P�$��	aj V�    ^�^�t$�D$   FV�B� ?:f��6�ǅ   ���W�W����& �F   j P�    X�X�D$�D$   @P��Ҽ��=   j Q�    Y�Y�L$�D$   AQ�ቕ�P0 D��0D LX��u��6P0 d��0D dX��u��P��(d0DX(d0��u�� ��j V�    ^�^�t$�D$   FVð��#��.����  f�ZnQf�8�[����& ��  ����&j R�    Z�Z�T$�D$   BR�Y �U�`L	f����aj R�    Z�Z�T$�D$   BR�f;�t��-��������&f��ݎ�  j U�    ]�]�l$�D$   EUÓ�nGW���g�af��aPf�!+�4$f������&��!���+j P�    X�X�D$�D$   @Pù�Tz�u����&f��f���-j R�    Z�Z�T$�D$   BR�Y�   ��u�b���   j W�    _�_�|$�D$   GW���ƽዕ�����j Q�    Y�Y�L$�D$   AQ�o �NQ��[�   �-c�?�P j P�    X�X�D$�D$   @Pü
��_=�&��2�&f�ډ��   #�/�   ��j j Q�    Y�Y�L$�D$   AQ���{)������&j Q�    Y�Y�L$�D$   AQ���@w���Q+���$������
P�떁�O)����&j R�    Z�Z�T$�D$   BR�V!��   cV�x�<�f��[f�ד�����Q���[�� �L   j R�    Z�Z�T$�D$   BR��Y��   x�m�#>�]瞋�A!_�����=P���_�)��������&��e���++�	����&j Q�    Y�Y�L$�D$   AQ�e)��!f��>���e'j R�    Z�Z�T$�D$   BRò�Ӏ��z��%�Z   j U�    ]�]�l$�D$   EU�=j����{8
���j P�    X�X�D$�D$   @P��]���P�  �   �O�j*4ǅ    ��9+������]
�@��j Q�    Y�Y�L$�D$   AQ�X�)��"� ����   �����M(����Dm(Pd�5    d�%    �    X+�% ���f�8MZ�   �P<Ё:PE  �
   -   ������ȉ�9@<�P����PP���)�   �Pщ�aP��d�    ���   Q�L$���      Y3�Ã�� �$   ƅ�Ghҧ�����$����&��j �Љ�A���   �%�ig��   `���!`*��aY�   ���a��:+��d����f  R`����a[�z  f�2
�1`�Ѷ3a���I�Y���9�K+��@9��}9K�1Q�   f��[��iN9�ׁ�eN9`�
   t|�:zE�`��aO������   ����M@�p�o���V�E����~��l����`���w�#VL��V���4�@D�~�\*~��V��<��BS��iw�̚�#VL��V���4�@D�~�\*~��V��<�A[��l��(����s���V�}�=���V��0�5!
�b
���V������.��D����ofXew�ޜ��oa.�}w�����o���V�:����#�"���@U�|�W��s��B���j�8
V3:�L���x�%ic�H�bP��Z8*'9T'9T�bP��Z��w�>D�B)�lf��P�zP�b=8P˄�f��f1P�b� P9��⃏þ!�z����F}�"�P������f
}�bP���6�QE�#}��E��m��P�zP�b=:P̈́'�f��f2P�b�"P�r��Zl�̟�N�ʑc�f��Q|i�n,�������Ji���1�@�������J��C�������@������G���A�󶷶�t��ҍE��O�۵��Ƕ��l���l���l���l���l���l���l���l���l���l���l���l���l���l���l���l���l���l���l���l���l���l���l���l���l���l���l���l���l���l���l���l���l���l���l���l���l���l���l���l���l���l���l���l���l���l���l���l���l���l���l���l���l���l���l���l���l���l���l���l���l���l���l���l���l���l���l���l���l���l���l���l���l���l���l���l���l���l���l���l���l���l���l���l���l���l���l���l���l���l���l���l���l���l���l���l���l���l���l���l���l���l���l���l���l���l���l���l���l���l���l������G6��l��}���l��RxCb������
{�l��ћދA�|�8���̊�\�a��e��H��ɴ���l�ͥ��� ���o����������aQRjK��;	�ʚ��-�'������ׅ2�8(��mD�&���ۖ�EL�?�l�����\ݯ�R���YXn&�i5�' ���!�L��S��2m{w��^�i��Nm��l�Y�'9�}-�^J/�����.�]�/ꍔ�pF*� Δ�l��� 3��� l��o��klTԵ�/�lG'�Ɠ8g��� :��ŔZ�sD����x���]��s��'��O����=�.](��@+�4�[s�h����a���˓\I�����6t�`��^����[^xGv1�����3v����\��ը���@��}ie�a����N���O�����h�dU�1H���fU������>�lA&���'���"�.S��Wd0�����hw�3bm��g���9�}=���\K����@��Om�0����aC
��lc|��r�M��l��o����pQz��&�r��T{�l��ѕ�u��I�^���JAmL�̄>�lu�(�5�x�U:j+�����ʛ��7����g_��lJ�Ng���ҙ�0-9�j�ݔ�O\;��� I������R�/M�Ѧ���Aܔ�_�JˌJ����r�q'�G��S����]l&��X���R��\�%�m��7?�l��\�$,���Hs����5��o�&�
;�.�ޘa� ���\�~R��L��Ѧ ���{҅4�֤��l���U
�7q�\��p� 8d�D��wY �<�Z@�Gma����
5V�ۀ�O��ABа�����&�kDR��ck �M�Z�6-�p?���ȄId~�����N�1�ӎ���n�8�A���CZ���b�T�l�� ��;m��jN�l�Ӥ����lMݼ�x���Δ�l���į��l���ތ��\`�RG��xU2���Nk �`�R����l�l� �l�Ӡ�ݽ��Nӭ ��l/lS�d���3���ՙx���5Sa����U�Tp�JP�\���{R?�0��.�����l����2R����l���`���X���3Sa�����T	p�jp��yO���R���Ob*�Ƚ�R>�2�� /߂$���l��jpU� �������X�l,l��Ra��љX���3Sa����S��l�h� ��vр�١�L�a�ӌ��ҡ�L�y�L�@�uM.�L��L�\jљ����aQ�1��?��-�Ѽ�}��֣��M<���楳��P%�0���I��Lø<������|��3�R��'
t����������o� ���˜b�b<]���I`�%����6��2�l�����읞��lKgR{�h����e����|������	���\l�ԥ7�	���l��V��ԥ��	���l���l�Ӏh1290n�11�>��I���\�u��e�ӦD���lt���L�`��`}��lѦ}��cH�J������cR��?���g�{��l���l����S�j�p�R!p��l�Ӓ�S�u}w������J�m���lF  ىQϮf���
�{�F�����ۖ�ֆ���'��'��X!?�v����{�tA�AC��}��7}d��uS�.��H��ݗX��l$5���0���G�XEƗ��O0��X��=�R�W|b��t� *�O�X������ض1μ<�)���?���C�������bצ��}��6�E�~b���g��������Y�_�[������D9��|�W"����CUq�3�	�=�F�>pE/��|6��;�0�/.���|�
�v6D����I�D+��|w�J�
�X�\�*�D!��|�L(���\�?O%"�\|�������A��8r�e�Tg�?�� �(d��+�'������HY3��6�I��x�ᩜ��R d���
�0��44gU��t&1l~Vc��t��k�`�|��E2��|ig�2��Ph�%�X=�]t�E刭{��ⓟ��;�h��X���s��u> �f�hŞ,�?9z-����k��i���/z�	��]nN��ˌ$�hս1yW~|1��ե������hաL�+�k<��?��0����,.��	�v���Үo��0�y���i���r��7	��&P�R�Ѓ���V����8('�h�M"����h��N�$�Uɥc���h�+�\YM��o�:�P�Ӊ�����{�n�B��8%���������8���(%�E��� ��]�o�@�]��6���8E5jBeY:dBR*aB,�8E�WB	�]��B�A�|�]��E��6���8E5jBeY:dBR*aB/�8E�WB�dw^{G�<(gv���8E�z�gN��x]��8EI�V�9��^`9E��ݐD�0m ܃�{�8Eե0��,9���9Ѧ9E�"(.�gr]k�_�E�.tr�g�y��.��]�cXDY��!Z���A���I����I�K�I��x���a����L8bM�a읆Z2-3ʸ^2gc-�Nɜ�I��I��PUp:z�Zo�K���gt�)恼�ʻ���nE���1�̒��K��x-����FS�I�nE���RK�I�{�]21�1ʫPU�=z�Z�(iҝ�Ts�PU�=z�Zo�K���gt�)恼�ʻ�����@�Z��U�~λ�I�A��E`��m��u�I�T�_9�9����h���I~��I����3���O�K`Z�(N[ފ�a�_v[!�%����nN�K��Z:��1�Ӷ�p�w �&�+�T��\�I�K`l6D���Z:��1��T~�Zx��I��>j�Z��K��%jN�ԝ����z��l6����ʻ�I7��K���ʻ�ڱ�]��J��N����(]Z�����M ��x|����M�r2��|S�H��M�j��F�Zɻ�I�l�<����	 ��Tt�Z�-���M��a��R���I���q���I15Z�G �I���0y�d���f�K�lR���ʻ���`������u_K`�k�����l��ċq����γs����8n�c�ΰů���8v�c�ΰѯ���8�0n�ΰM����8�6c�ΰ�����Tc��1���m��m�B�i��O&��m:�|����6�������m�Bg~��'�Epf��~92����m�2����m�2����m"<N7�{&j���s�����Y{c�7Im���	B<Zц����d����'�Qc���m���h���m<�/a��� ���ۏ$����"�R?m�m�����aҦ����ew��rj��$0S��%m�
�{-i��T���Rj��0m���$��ۃ�g6���j�����Ҏv�g��{Mf���m�����|;j)�lc�D��R2jIu�c���e�jI� c�B�� �)A:J#A'��y�$P���w��X��.4�p]%�xc8EfK��!�<ٜD��b��G����'z2�*�1}=X��`�-��׳*�I��b�b�*$So�QN��!Lɚu[��c�2�f���l�A.��I��u�ژ�|/�v&U�/N ;O ��z� 8���"VIa:l'�H6�AH&F {>�Qd�Qd_H&�8{e��j��J}/s�� ��e��u&U&�0Vo�E�ui�W&&\ߙ�K�\�u�!.Y�-8�A*/�g�l^"[�U��S([��}D�]c����E�`4�_�e~����R3+ʀ`���[:�J�
0yam<��m<
�J=��kᅩQ]ܪ��a7t���Z@�J� j���)Ǌi2�Mbz��_6�X5�F�w�J%>�)<4�Js~(���3�<�3k>�J�M(��ߵ9��6�8A�F4�J%>�/<4�Jsp(ĺ)�3�<�3i>�J�w(�y�uB��FP�E;x.�n4��I|So��I4~Py*�0c~�w4��l>�J�~�p�������M�x�X��=4�J0Q����F���J<�r��1{�y��3��z��B^�����$h,�w��������������������������������������������������������������������������������������������������3��
	��g��G�����wev5R<�>���ՠ�G�<41�bШ��L+������*a���+D���_Euz9����Duf�<2 ���gd5 A������͸T�~Ea��
��A����1)��$H�(���L�
����籷��{�^��d���k ����6�G�t��ӈce"�Ӳ1 ֱu���nj�"	eБ�h=6B����؜�w{Eп��wЏ1��W��Z�����é�Wr�>��J��Ԛ)z�����\@�^��d�v���O|�ߗ���[���=Y�԰��g�x���ԉ�w-��J���p�g����*��ͱWX��z�8���nsտ���J`}����ϯ����q�.�WHP�ҳA-C�x���&�r��[U��������qv�������d���e�Z�6 �L.f�R��k��/���"�YS��ժl:�����ʪ垪n6�G-�/��ͮW ��z$6Р뇽�a"��^�}�չ�'ж������sb�\"D�C�g=p��Vl���	��=�/>ՁW��,����`BB����C��5��s����%��o�G�����s)ӊgt�����ԓ�%�z�����<��}�m`�a���|��E�������9��dL����2���3�ڏ��Z�b;v7�S�uS҉�}�aa�1��J��d6��-���i�j�e9��k��%���<�R����F翋�~h�Gߐ�ee3���0١�~ƺe����	���4	��U׶�����øa��GD�Y���Lm`�k0�ya�JJ����f��pO���̨���4�o[�[Ў��B��8��N��*�ͩW��Ӛt�ؗ����B�嚊f�﯇�l��dn��7�&�͓@Z�y�������(A��:����	������y������0k�dFp��(P5Џ��a����0��4��bȡe�ֲ������Q��h個]��hN��"��������۵����D�����Q�g��������@����L�m9oB����}��叏�M3Ӏ���4��g�A�{�5��}$І ��g�Tny��a�<D`����NCYX��dYIҞ����
���Q�<v�i��V7N��]��e����}!�����}����9`�ܨ0��I?�U�iո�vqA.��\Nv�YS�nC��}a�R�~Ea�²��D���Ju�OӰa���R�~�o&YלA�����2`w qa�OP`�Ul�=\W���zv��0��Zx0J�gRvq�����������ʰ���J8u�OӰa���R�~�o&YלA����ş|�*�g�OP��Ul�=�T�C�zv��0��ϣ�a�wqb�|x+�($����H��J8u�OӰa���R�~Ea��zלA����ş|�*�gENP��R�~�o&��^�1�I����U������;�������G���[!��i�t ����4�^ׯQ�S�ʎ���:��kk"�׊��R�~�o&���^��姷��I�!���ׂl�?����Ǒ���ψ��D��}�.�����H��Q��5�~��S��0��:a���gHMq��(�&Z��rx��*��0��Zx0J�g�Iq�S�s3��G�p����M�v��
�f~���R�~�o&Y��+���r�@X���a��?b�(!)Z��rx��*��0��ϣ�a�Iq��S�s3�/Z�p����MьVi��f~���R�~�o&Yל+�>�Ne���:kVa���(!)Z��rx��*��0��Zx0J�g�Iq��S�Gi59t�����0��Zx0Ja�wj���X,�[��(����K*�����/b����V�|��y+�!���	�A�t~3�*�f�&�R�~%�����D���Ju�OӰa���R�d%��IלA����B����g�OPa�Uv�%�-1}v��0��ϣ�aRvq�����������ʰ���J8K�I�a�g�R�~Ea��zלA����B����a�OPa�Uv��%�k1}v��0��Zx0J�g�wq��|f9V(4;ި�H��J8u�OӰa���R�~�o&YלA�1��ş|�*�g�OP��U���%�?}v��0��Zx0Ja�Hq���WO䍶R�u���D`������?�A���B��Ĵ��0�qO����n�n��[��Z�$IP�����B�R��0��:a���gHMq��(�&Z��rx��*��0��:a�����Iq��S�Gi5	רp����M�v��
�&�g~���R�~�o&Y��+���r�@X���a��?b�(!+��իG��*��0��:a�����Iq��S�s3�/Z�p����M�v��
�@�f~���R�~�o&Yל+�>�NE�����g����(!)Z��rx��*��0��:a�����Iqa�S�Gi59t�����#cc�ۆ�af����Mo��n������_^()P`�a�6z����h���o��)E��\�c��cH�삝������^�/}o��G��A\�=@�A�4�������գ����h ��b�8��>��"	�Wץ�<����G��Ǒ��˧��S��Je����k�*�����*���qb.�����n�ӿ�����2��p��Ϳ�2��5j��]�@<�c34.b�b��A�b��͆v�0��9��L������3�	PI���m�a����?����j6��<f��3��ge�{a�R�~Ea�²��(����D�塋���|׊�Ӂ�h,���9ń���a��iк;��	�g��
2���G���g���b��:��p���`|�
�a�2�׫!�H���>@	a�M>��Ŗ�;w�)����\!ǂ4Z�ө=�K�ֺԌ�o�%G��>$PGb���u��:�Jò=q��6��0��Zx0Ja�Hj��Q���(�n2�g���C93��������L�^�җ�[�����&�!���N�l¨6b�KBȫ��|_am��0��Zx0Ja�Hj�h�z�.ޒ��[���y�8r����������G�k��-UG��U������?����iu9�����MQO)�:W7�g~�g�R�~�o&���D���J=��I�a�g�R�~Ea�²לA����B����g�OPa�Uv�%��}v��0��Zx0J�aRvq������ea|�ʰ���J8u�OӰa���R�~%��QלA����ş|�*�a�OP��UhK�=7��}v��0��Zx0J�a�wq��|x+�($����H��J8u�OӰa���R�~Ea��RלA����ş|�*�aENP��R�~�o&A��D���Ju�OӰa���R�~�o&YלA�>���2`w qa�OP`�Ul�=\W���}v��0��Zx0J�gRvq�������ea|�ʰ���J�H��.B`���R�~%��IלAɨ���2`w �I��OP`�Ul�=�T���}v��0��Zx0J�g�wq��|x+�($�K��H��J�H��.B`���R�~Ea��zלA����ş|�*�gENP��R�~%�廁��A�������� ]�ɱ��%��X��5^��z��撷իG���9�+�E���S�����0��:a��X`�vha�雰���^.�6h�>wb�w3�Ӛ;J��%�q�1+#7����^��؃k���v�����8r�r�:�ӗ����Q��˻�"�y�t�h�-n����w��g�Ag������dЮp�é�g�HA�N��Jx�H��.B`d���jqE�
�H�������� ������[��Y�F��BEָ��?�]9vB�m������ɽ�^Zk@`���ݷ�NPz��#2a�t������:�a����M^�v�☨�*���/�r�oz���G-�⃩�4��z�?�������G�]�3����v�^S�K��-���ؖtu��C8�徽¢��=)��v������h?^�E�B��՜)�ә���Ã��w7���f▱��A�n$��kpR��6�&�g���ҳ��<�	1da
�X��5���J���8T�Ě���uPs [����pN`�`KKJ�aama�ۍG~����1�0X��I堨��b��H���~Q�  ������0Z�:臵�%�Ϩ�/��TaB�ְaew �w^al�O���oay��D̨���I�dҨ�+�s ��8�X��ި��
�b���_:��g��Y�p�ؙUڐ��2'����屿=]��
%����_;�����<?��)q�	.���y0{�g��g߰��ﱗ���B��ך��@�e��G�0��|��^��@��g�v{X�t�o��D.�Ũ�������d��I�6+�t� "��g<杉��W`���	�M���Z��G+	��3�1��NJ�YS�������,�t<k����s�	�w�^S���J�g�K֟�b2*�טW�{ǔ����ݭG��'�,�K6~<b�a��<A�}�!��
���D&�"��؎�@	������*ݨ��l*�.����`�����V����g�v�����0��agL�7���<,t�=���a�O�K�q}��;�¬����0��ϣ�g�vj��?����Ɛ�-zU��T�m�[����/(/���y,=���	�v�.����:���!<R�"�L�����������IӚ�����e�T׵��喿_P���囦����Q�`i<D!�e?.��0*��X�~�x�8������Hꝇ�!Я��� ?�x��T��wЄ��*�7�l�siA��U���C���F���R�ԒZ��V���f����ean	�=���:����Tr��-���g��vkIb8̨Jc�:t늦O`����s�因w��j�m~�������ءUĎ�e����]p,��"8[D��������c�-��ڢF��?�Pq�A�l������al���}���\?��h}	!��Una�v60�ac�G���>��$��.?%�������_�Z�3eV�g���I�os�к9L�����H����Pטd&��H�QA|�|.�����Mf���fu�5q����X�4h�2�a�	��W����&�ם��b⽼C��6�g�H�����(�q�S5�u������dq��J����y�e�����b�{��5��ȇ����ཚ����%�U�������QD_�׶O�	ĳd|� =�a����J�[�IR��"���'�z�����FԳ������h���b��J����k4�����������J�Q�J��k����k�t�����^V)M���6���7��8k1�m�0ͷ����͇�O����㙘�?���SU��_-����g�ix��բa��O���#�O���B��'������z��u�Gy���ʲH��@��IP���Œ��O���EZv�2����Ϙ�E�$e{�F��?"���8M�����CsF*Z�|*UD&�*��05�ʆ�GD�Y�0��g�G�5ȅ����u�?ϝøazh������u%���s�'��*).���R��H�v�P}���0��a��!�{���m�䵇Q���!v��	�Z���~!;��%�ם�G�*��IP��4#2����&�L�`y������<v��g�#��,	��3��ч�X�^����������R��d��g�oj�z�W`A�����zЇ�툩�3��z�����M��4��
SP)i��ga�6�4�?�)�7��0�
�;�BX��,5����v�������D���a����p�Ta�xy��w"���L�Q�=��v\� P�w"�w�g���g�6l2Ө�����!N�_���i�Xh�,�R�d%�����^�0��S$I�կ����>3Mi���٘ʿ��CSvmare���a�N� �Ԕ����R��_p}��.�����VЏ�Г��H���屻�+zd^��`��9U�{4f���$(��&�H��1��������h?b��gW\�K���A,��'�����O"������,ը�<,��Ш%b��	��~����g$�A�壘�=?%e���}ٹ�,"��\�h�4|�A��֨��9���׊�����s��%�9��0��Zx0J�a�wk�r[��ZJ��W���?�)FG@��X��gٝ[������ΰQys��0�͆g�A�� �Ӡ�����Ty;v���K�����Yd���������RO�������AXq;WY�d��r������aa}?��s����Y�O#��2�3_ͮ ��>�d�oq\�b�R�釄Б�iW�����B����qy���3�������^0��&������'���U4��#�^D�3��g�2�x���KwF@�����w�1�*����G>����ƨ�}����&g�x��_� �Z��g����*맱�u������@�����ʶ�H_^�-尗i�����-!A�7������X3V�d�z����8�A��.�"b�[�2���К��<V�����Z�H����uJ��J����HR���E�9��}$��.�G����E�N����������-�&m�����x�����z������Ƙ�O����gʋ�D��]�r�+�P�����_����ۄUH����l���?)��O�Ը�דJ����G��x��x�eo��5������f�`�����^a�8��ea�6ǅ�������[�ddѨ�Hb�����X�6����:�װQ�������߅[����������~���5�bW�DL��z�\`�x��٘�9�"��o����'�:��ފ����ɦ�䈏������r[�͌����1V����]���w.��{���Χ�������;����!%�UT4���2����\X���  ������+�
�?��j������ү���u�:Q�gB5��{J�YSn1�\�g��떓�%b¨��������-s�v?�O��n-걕j�oaʑ�Cv�YS! `��,��@`��D
��g����K����5-��RO������H�iVlП�2J���7T�׶ �)�Z���)��ۨ���w��]�@�U|���mz�6�g1�K�G�?�]�+�ޙ���_���D#�Ωa����sQ�g@Gʸ�h���7���=����������W���芺����0ݪz��z���E�䣻����]���
��術���]��Ds�-,��'�6�gYA��*	�A�D[T>����ACYX��dY�����qQ���:���g���E^pWȭ��g¶�2��I���F����x&���Ww�o���aŀ�SЏ�~P�Or��5� ��A�)�������g��h���huI2!����ڰ}a=��JIӏ�ɿ�F~�W�-����E���%aШ���P�����P����&��S�����b���)�~|�}�����'j��+���S�]�2J���>g�����k"��2k�v4�(@p��81Q^�W'8�����������n��L��&ve�������~Q���HY����X�w�|�&��O74|J?��O�4|T֨�O�>�"�|.�hd*?�Y�ۘb�ܻt�K��!�7W_}`����?�p|�Yv}����om�@��4A&�J;81g�Сh}�m�������S�����I�4H��4�O�����������I�4H� ��aL�'�^�uS������&"�����gl4�(l{������S�����I74HH�4gu����D G�֒tT�݈��ZE"hMcu�{���v^��D�I��r�s�1�wT������4�O�R�����M��n'L�l���������_����'{������U��z� Dl{������S�����I/4HH�4|]e��O/4�!��h|�O�Mw������{���w$"o(0�>@��M1��L�,4�O�R�����M��n'L��8������U��z�D���~Q}OL>��y7�1���]��f7�1���1jKr���1ԁ�1�������1���1�Է(���1y��1�aQ��p��͸{��Ψ��Nh =�c���U���qѕ����H��7��W�1>����������Q��ק-�㱳1���n�)z�@�pKe��K��a�G���E�	�G0���H�d�6mB}���U0�!IR��E�H�1����?�|�hE���-����>��+${Q���U j�V�KT�y�cI�	�L���� G7䩆!�<ܱ����gȻ��a�_dQ��<3J��(Eg��l�^0Xܾ���(E3���C9�q�:����(EK�Cjҽ��Վ.ik��(����:�P�j:FvEo�>9g"N�rrC��:p	�x�j�%�!헢a�7��(E:yA�W��Կ8M� 6��4Hܳ�Eo�(x�J׃U�%p����q���3-u#oB����N�s׌*�R��"KCo��p���(E�(y���(Eo��V�W�^�Ա%�M�^�WEo���4�?�_;�����`w��W��_ϻvǷ�wG}5`5�!pq��΢��7@�S����a�S�:4��	�۹����:�&�j�h��SMŋnI[�9��co�T�P�I6��g$����S�>��`�Z�1}���Zn�o� �{���&*�w@�Ӛpߕ�S�������/����Fw�U�O��SE��❥��k/�?��� ,�́�^���eSX3$�A���
2�	��>��T��T9O{�O�@�)�"���U#�$�K`PTV�T�um�l}^�7�$vb��l��kǃ�Sr6��4���c��;U�����c�@�_��=��6n� K���<s嵨*�h_ҸAST��^��Ӷ�u�T%�I��1F3�5� �S��d�����s�~��>�k���|�S��p��^	�U7'���`���3!TP���S�9�k�n˲��&�7�������T�?�f�
3+���4����^�j�T�G.��́��fH�l��Z�G%��dRxQG�<~��c:���T��Z�5�hl_yC ����ӆ0����S,moT�5?�h�,���:I�iJ���J{$6�SxQG�<~ڎ:@����Ae�^��"TE���L�r��?U�2�R�ھ�AS��T��)�TMƆwS�w��S 2�b�!P���zo�O���TV�w��1F������SB���u�T��i��%^�1�w�k��:GS:�T��T�ӄ��5��B��
���b7�0R@ǀ�T�ф���bEZz��:�^u�?�3���c������dG��,��T��]"�o���~8`�?T�̘^��j,�	Q^*� �M�̿�u��Y�/��C����S>3_�:��F����h����S^1�b����i�*��(Ȏ?^��D��`4�S�Mq]	�U�Q�x��Vc`�����)M�_>�gh����,[/�&V��ߔ���ۭ}St�sh�j �kj
�^�S[`2���^��@M��Q�:�M?�/c�St�>WR�Ɨ��5����A�1}�T.��0�Sr�5���9��k�3/b�ʥQ�#�7�XaPo+�_[�չm�0��o�����t[SxQG�<~:�:����:l_r{�q�)_^��Q�$UU��UT�S�D������jbP���C��M�|S8�Xɴ�2�	+C��^W>��Y�����cI6��V��\��ST�ס�U$TzC���r����~kT�P/_o5��Q�}��4��ݷzT�~�� �S����ɪ�'F���.�ߏ�/��S�S���I��c:���|��S��]cځ�SW[{�ؖ'1���쩴#w���=�^fÄ�A�y篠��fu��~�c��)k�SgiZe�X�e�s��qx,p�^l�Ga
��^�XYM_�*?�
 ӈˬ�6�Ke��R���J�s�&�8̳b��M���l�|S<WRk���S���"�h�
q�<3T}�\e��qnt�C�f��{Sr�ơU�AS[�鏀j���o����(���ĉ!�f.%#T9B��´r��c�p�$���~.�^,q/_o�˪�՝^F���X�~�:U����s�SX	��oC��)]���~_��n��S󺵤��er5��_�|��A��9PNi���c���LȏO�Td6|_�S�g��x�S��%�vJ�	�,�Dn�l�S�SG�<~���s��*Fw�w���v�Ty�S������I�cχ�^��ɰ̖�^� )C
pԃ܁��|��Sʸ�3^7�S_��ؖ��+׎�d)i��-Z���!TES'�
c��sҎe��nyi��"KBNS�x]�u3h�{L��^J�S�Q�0���^T;��&#?͝^i���:U-A��ϝS9`���k7_m��#��c|n����ю�^�ƭSl�_+E���}�S��
?�^@[���8(��/��A!�ҭ��^o����L���M�1Yzѓ�T�?	R��BHO��ܮ���Ȍ5�͡K`PT��T���k����ʐ)�?^��L��nJ�Sd�;{�"�۱j�.�_P^�����SX��F���;EzШ���A?�]P"�TRP�T �O'�f�Uxf3[' �v=����e㓸^�W�^c�S΍�7t!2�}�e��S�n�SE"��� 8�Q}������M`�'�T���%P�^�9����N��S�dJ�UjTEx]�$��c9�^c���@S�YBT��^����������� Z/z�r��S��S$R5��S�����(K�)��/��u�9��v{��0��++�)n|�s����/���x�l���/]OI���Έ�Z=��Q+{���S����scgJk�:�_$I5º�S�4l{I?�2���4�S��ԸPPp�0f͢Yx���S��Q<��[D� PS�#�����v���Årg^r���B'��<�9S����N>��f��8�[���j�{��8��tW<S�2#����p@y�l?��?�UZ筞٨T�9�o|ͺ���|�T�fl�܎�3eM��ź�?x�S�P4T1}K&�X�P�M&�\d^ē�ۀ�sW����S�Pa�4}ׂ�S��5�Si���~ �m���j��IO�Q� k�I��w6"7B�l��Vq{B��o�>Ė�S��S��S��aln:�{w>���dz�>7j����D�`��(�{K����*�x�qP��	�����u��<7j���0�����?V�SI�������S��S�9���gz�>7���������"7J;��T��p�Iu��Y�SO&���dPI=����S��3�󐤖n�{�{K&7\dD*7@�����A�"7J;��T��g��{�?�����w���"q��$��dA��������MHә38��{�{�
%��_?��!���<ű�[��4h|J�)�^0�S���P'�S��u4PS���FSS�㹐^նL�4�U��>7������9j�ř_@���S�S��S��R*���S��S�vGV���d�2�{��LW����.�k��S�_@���S�S��S��R��R��S�vG�ڛS
T��1ɽ�^�SS0�T�6�2�{��^0�S���O���3�7����7�����H��w6"7����H%&I6"7����H��H6"/�������h4'/�Xi��I�H6o�_��9L���\ք�S��k��d5}��S��8]��S�l6�ȏ�g����SAri���{�3��#_����SþTaTB��l����H���s�p����BǯH��u�>�X��̍a�<�6}��RaF�1}MC��dR>��:�t�ovG�_5X�v\��㟔z�ao[ؚ��.rF�{�)�BnZ~v��_��儼���ox���z������r�	m8�)�a���m�"2����a��m��7������7��K!���@m\@mn�7�O�!������7�tң�*��tH�aF�RDڊF5Gs�7���L�#BPȌ�͌�2��2�����7FڊF5x~�7���ͩ$B�Ȍ�͌5��Y��� ���Lo9jI ���7�.86ӎ��+N�{��W��9��m��48m���
\u���!F���6$��IcAN�G,Ƕ�*�����&�i0T�GX/��Aj���ܻ�b��u�����u��ԛOlӮ���o��1�<�)�d���h߉-b
b���fd�Њ�e� �*�
���J������g���X��U���%hp�U�?��+�67�l寠��\0}Q�.�;���[�Ųޓ���IkE��R�	�(��U��m��5C>1���.n��G��� ���Js�sj#�J���������
J����ڸ��p��Ae!#����ǧ�ד��6Jx5+�5�?h�=�1��߶z��B)���#�1�~ܟN��}�M|С^0�;�1���v�7�ؗ��L���T�� o����1� �lHpg4jf�6j�1� �CJn�<_��NJG�P�O���T�1� o����1� ��H�G)jf�6j^1� �/JǷƩd�FLaT0�B�1�To����1� ��H�W+jf�6j�1� X%J���T$��?��>��z2Sý��� �1�6 �ç���H��(w�0��f������&�H���Q7t���6\͌7�đ�!9*��u�C����P�����Bї�����){�[nEY����8w��D��biß�����g����f�b�bim��T��+"v��
��&�!����t�,D��$�oU�j뮾}��MGW�,4�Kݗ�	?�$A�,ŷ��bB��$Ը�x?|�B������N���B@ Ͼ`Q�N-S(;��z�w�Ĥp{(�zW<���g�$A�m�g��+i�{lй��1���zF��J������^��S�&VP*=A���[4|ɋ#A�@���}z�[��j?S�n#V  ;���gy�\�G�ǀrUc}w�[��dyaj�i��LuU��m��l�����uU�q��!��dm|%�S����r.t����Z�W=P;u���-��r�U��ލ�
�WeĀr��������m5� �|�[rUƀ����O|�=���[4U�SƀR�8|3���h��Tƀ��8���Z͐�[4U]sSƀR�;8�1�p�h�hTƀS�;��s�Xm.�[4U�]�X�[��`�X'l�JT��K�[�
��� +}T H=��>��,/����A�~i�c���c�����2�_�2}��a'-�1����ѽ'���`��ť�&��?W㖼`��G�BC�1�׷m��|��Bc.>�c�j�{� �`�
�b��X·�s�o�=����Gb*�41�_���7T�k�_2)�Ɗ��"��d��_4�~0��)���r�C����>,k��Ya@�m���HIw<�S��>)tfS�Y1
��l���;_2,�N��A�
�Q}��e�f��%'���z�[��ڑ�C�7�Zᦢ&�FT1f ^�F2�*�W�H���S�<5�|4�'F2Q�!/�b��5ą��U$��1�OGD&��A�_'^�F�A��dV)�Gt�E��)��{�����7�5��"^2�6�6�~��W��U.�$̍�����y����h�G��2��bZ)F2�&K|�_�d�Fp���AI#5fqʄ�U�9<�?";��(��)�b�!�E���W<��2���O��'�p�T��:�jB2��]�%���~��2�6w�h�ex�vF.ة�24 ���VE�hF����Ͱ~+$~��vE2v� r�F!�8Wƭ�k����!%��2>=�4�%<�}��Q��qQgn�|U�2�K�'9&��`�P�j���H��2/3m<P�c��F������:�,W�ǫ�g�7+б8CH±��2p���7v�3իF���3��-��� 0�0�r��ùhF#�J"<��gY�mJT�rq��U�~�+7lEB�H2�}%��@��aCU�o�ކ��S��Q��5�7�M:�PM�}=�݌�O5�m���K2R�n-$��P�`/Q���4���K'��t<ޑ��u��T1��Ꭺd^����_D2�@�� X�#�d��\UkB�0�EU )7�KP҉�[UFW<��j��G�<W��΄�<
2�T��Q�Tzr����F����!+i<�[���'����^�r̓5��?�_2+r���4�TcY�d\�F�ª2��w���K2��7r��;+Q�R�Qh$�ߣpzhqZ��2i��j�����(h��'�4�$����� �6sv�w���H�C�l-ﱿ5�+��, E2�7�M:�PM��J�V6d4G��.6d�!���P2_2�q��J����MD3H|(Y��2?��;�<s<c��*��6�Kr�뮦ҹ2߳5.	'�l���U��MSG
�Q�[櫓�2~J�B<�"�2O�e�]|	�	cQ�KJ��F2J��� ���>��2m��$�ak�;��-E#�2��E!�}�^����#uwrꩱ���|�!�����Pv�w�,=��m>$S<��%7���mo^�r
E�g�p��B��?e4m</�R?�VT���~�d�QHB"�>F��_�2�� j�U�|7F��"^F;�c�`�<�28q��MA��"��.i<_s�0
�lQ8�2��k��*-�1��?���/2�l��HD2Q5�� ]_b뀽��T3���.�;���2*�+5u8��(α�a�i��(̄��h(M��j�A��^VQ?=��9�I�(�DΣ���2��a�������P���I3·7��\2Oa���F��>;B<���?߄骾��t�3-m2~�K�L�)���˺f�ƭ�'�3	�}��R.�hVtV�S��HNW2T��<��������^!�}�6~.�pOl<O2,��&�E�:cA2��O�,?�0�O~J��2i����;����٫�5�I۠g�2�3Z����2�F]��o�O5�m;fE2�Oq��w!�����<7�n��IP
J|�U~Y'܋�n_���Pi���F��2p�'	'a����P�4��g.�qu��_D2�����lQ��};��aI#}~�;@��h(�4=��;�=�j��$"/�kQ�X�p�9'&�-�Ӏ�^�4�^�Uz��/2��"�Tg�2����j��^n�r=�d#Q��&qY�(�>�=2�1+>�}f��%��5�>���K2ܛ�<Ҭ�2�������i�3իF����2��G�,�ӆ_��ԁ�.f�;�K�3�
�?=��j6��ҬF
��Λ� |Z�#rJUE24m�r��̰������+������F2�9��!]_�8F\���	`����5���(Î퍝�6� 0�0�Rr���%��#Mw�$�0��@���1�W���𷵍�?ecV<J�i�1�i<���O��eo���5r����K2WM-!nT�E��m#�dCP(�2R$F!qY�2&�K��_ǟ�F	�����$�'�nT�!��B�Ʈ����B�O5ls!�fE2K
J�N7$xc������k��α�� j<��	&[���H�d�A�$��^��X�3�!�t5<6'9�4�4�^�h�F���9Fa���<<�{_���`F?���a��zx;\&&(��(��4��sLJ�4^��?I�2�KO!ϽG2e�����8{��J7l��?_�PUB1F2��ҟ���3^�F2�)��*�$^�F��bVq-���F�)��l>�$^�F����2Q<��i�;�C飿ng)�)gၥ�@U��*�2Q�Ew���5�6���͆�c����2Q��&J�F2��ړX52P���H�RA�����Q�J�C鉔�����5P$^��(Ka���yI�j�V��g�|R 7$y��'�R�T�-�#h�j\�o4��T�u;�v<����@�ɻ��W,WK?�҇[�+-�p��V�1�%V�=����s*����΃:�Û��G����f�F2�I��I��I��I��I��I��I��I�_�F2Q�F2Q�F2Q�F2QE2�.F2�Zu�.\u�f'���I��_�F2Q�F2F2>�F2�Zu�A�r����=�v(�I�(�I���Zu�A�F2Q�Fj^�Fj�ID2Q��$�I��'�F2�I�I��_�F2Q�F2�I���I���I���I���I���IDj�9�9_�Fj
�r6�r�I���I��_-y(Q-y �I��_���Ic�_�F2�I���I���I���I���I���I�9��Ur����q<_�F2P$�5k�M�_�F2Q�F2Q�F2Q�F2Q�F2Q�F2Q�F2Q�F2Q�F2Q�F2Q�F2Q�F2Q�F2Q�F2Q�F2Q�F2Q�F2Q�F2Q�F2Q�F2Q�F2Q�F2Q�F2Q�F2Q�F2Q�F2Q�F2Q�F2Q�F2Q�F2Q�F2Q�F2Q�F2Q�F2Q�F2Q�F2Q�F2Q�F2Q�F2Q�F2Q�F2Q�F2Q�F2F~F2QF�;^�FK�5���f���>`9�F2Q_�j늪��F2x;���H2Q��GU�F�ˋ`9"j�S�G7Y��2Q0:x*$F2Q�+_�HG<���sjP�S���ҹ�a6���K���K�c��5��O2�I�(Q��M.��M#&�M$��?_�F���K���K�
���l��I�XB���)_K��ͧ�f�2��%F2Q����!`9 �վ�Hař�ؔ�U�F(�*�3�+P$�)$�z�P�Fv�bbZ�F���K��5P-�5Q��)~�b^�F�
���
��ߜ��5�Z�2�z�.�]�����5Ѣ]2��7P$Ɲ"��MH��R_$�Ĺ��8Ŵ����t�F2���)_K��tH�8��$^��$^�F���%�%F2Q����?`9 �Ց(Ka��2�M����B�$d%.&��I4!^�sRt��9t�լ'�#�}��sv+!�F�K6�4�>ـ0�;�I�(Q���pE2QB����F2Ѣ�2�ֿ2Q�Ƶ�����F2�z5�z/�%F2Q���u:`9�,��H'^�FK]CD2Q-�*Q�beZ�F���K�
E2Q��9"m<_�Ƶ'�����F2Ѣ\2�I�?_���	�s�sI����H�v���<�F2�R�(
ɐ	T�F�K���Z�F2�j�s�F2�'H���2Q��9:��8�I�<_���	�pB=�XSw���ju6
��{=����l�5PHz&����K2Q0��<�?_�.֒bT�F���K���2Q��c.$�2Q�,$62�j*��Ӊ��H�]Ϫ��F2�B��$�F2��H2�$��U�Fl
�� ��F2QK�+M6�cQK�5#A񮕃|T�F�S�g��������QｵH�'�5PD�j_t�#��sZ�FH߾'Ca\�qs�F2��1��D�ү��scZ�FlBv�ـ�F2t>�7Й~C`�F20T��$^�F�T1�F�F2Q�;}�~�@"�~'^c�K�;��K2Q%3Q���{�G�΅A�C�M�F2�V�1�ZA4וTX��皐��Ϡ���F2���2Q�h�C���b;��E���W�܂�3�2Q��q��e�����sΟE2Q������5���U�2|��2|��2|��2|��2|��2|��2|��2|��2|�퍗��-�ޜ�<[zV�?�e�ϸ�,�.X�!�UB˸`�cp��2|�Y�_�ޜ���{V�5��V7|Ç^���)�X4�{E�� N5�ɳ�*�2|+`0|��Gb�򗼛�3|�X����tB� �ޜ�<[cV��K�I�6�b=�+�[�?v�r���i���2|�cp�f�2|+`0|�s�NY߸c�_�|��q���2|�Y���qB��ܻڸ�~�2|��k����� ��ۧ�}�ૺ��2���2|�ר�,����� �<|��2��q�����'�/���˵�G��,�2|�L#|��a�Iz�G2 �t�T�u�x�2|%��T���>:�L�J�n�2��:1���>�ړ,~�1����l�����m*򂚸�2|�"$|��aB���`�2]��e}���r/�2l,p���������S�PZ=d����1�1��O ��g�dxWE���'����!���f
��긔�]�f����1�O��OZ�0��ϼ�✡
@��!��ad�D�tJ��ٶ�]�����f����1I��Oc���n�OH�����FDT�.Z !W���c�*��?��9�~�Q4��Q������8���pŮ��&��.W�c�*��?��9�~�Q4��Q(�������g�*��]�f����1�O��O �0�]f�a�'#o����o���b��]�цz��F��EC���ِ �� &O)��rbd����} (�'�x%�	��l+� �3��3��mg�'�[�f��T���´��~���[��
͞HE��-}��?�ѭ��ٰ���o� ���W�;+.4J�5����dMq�l�/0I�T2yQ�����Tp����f�8/�:��M&� ��m�g���ÿ����ĳ�{��֊�Q�.ڼ}ܬ��R^���uYo�:Ԣ}�?��F��yEfMx_�$��I�}ܔ�R�eY^ʟ�ˌ��ޘx��~��_�K$�\'� ��.�j�vG�%k�:�S�%�I�oG��.������e�ĭx�_Ѧ����G`����I���h���k�����X�4����%�O��/����I��ᐋ�f���k����;U��U�uM��,�t��r/��r�W�-���t�GI*I��G��I��r�������k��I�,�e�z��Dy�+c����qv��IH���ʽpVʽSI1���<����Ϛ��<�絳�q?��IH���ʽpVʽ�I��"Yy3k��72�/S_O��wr\?3�U����s�%�4�|_�J%�0�ϔ���Y$fl���5ɷ#П���QL]�qu	9��BV�U�ײÂ�О4]Wwܟ��L��3}���8���~�Zs�!/��Ͳ:v�����|/�ݞ��Opi��4[�lU<$����}-E�h��mU���/�}
�U$�}�m��W�" !�"��}r�l
l�P�I�j���0]��n"����L�}* ��&s�Dpس�}V ߤ"ԓ����n�!�����^G��N�//� "--/�#p9S�}! �p��IP>g���T��5/�� �cc[�#z��P�ũ���]v�,@��L>^��6�h��c��ǜ2�W�6�N�o�1J�%<8U�1~;&������J`f�:��8V_�q�{'4Si2=�e
X/�G��{4Y�����PYl3��-1�p3�e�ޮ-���=9��8��y*����5l�ST���7+�S�>�����7+zwsPm�U�m7%ֲ��@�*ҵc����2՞�O.g�����"���6���Pą�!�Ȼ,3+�3ڮ>lR�Dd����Sˡ������<�]
�V0�'f>�>�.n�t��Q���Z�k���X=����C)���,�sT~l�{6Y��* ��f����|�~7��y��sn��sn��sn��sn��sn��sn��sn��sn��sn��sn��sn��sn��sn��sn��sn��sn��sn��sn��sn��sn��sn��sn��sn��sn��sn��sn��sn��sn��sn��sn��sn��sn��sn��sn��sn��sn��sn��sn��sn��sn��sn��sn��sn��sn��sn��sn��sn��sn��sn��sn��sn��sn��sn��sn��sn��sn��sn��sn��sn��sn��sn��sn��sn��sn��sn��sn��sn��sn��sn��sn��sn��sn��sn��sn��sn��sn��sn��sn��sn��sn��sn��sn��sn��sn��sn��sn��sn��sn��sn��sn��sn��sn��sn��sn��sn��sn��sn��sn��sn��sn��sn��sn��sn��sn��sn��sn��sn��sn��sn��sn��sn��sn��sn��sn��sn��sn��sn��sn��sn��sn��sn��sn��sn��sn��sn��sn��sn��sn��sn��sn��sn��sn��sn��sn��sn��sn��sn��sn��sn��sn��sn��sn��sn��sn��sn��sn��sn��sn��sn��sn��sn��sn��sn��sn��sn��sn��sn��sn��sn��sn��sn��sn��sn��sn��sn��sn��sn��sn��sn��sn��sn��sn��sn��sn��sn��sn��sn��sn��sn��sn��sn��sn��sn��sn��sn��sn��sn��sn��sn��sn��sn��sn��sn��sn��sn��sn��sn��sn��sn��sn��sn��sn��sn��sn��sn��sn��sn��sn��sn��sn��sn��sn��sn��sn��sn��sn��sn��sn��sn��sn��sn��sn��sn��sn��sn��sn��sn��sn��sn��sn��sn��sn��sn��sn��sn��sn��sn��sn��sn��sn��sn��sn��sn��sn��sn��sn��sn��sn��sn��sn��sn��sn��sn��sn��sn��sn��sn��sn��sn��sn��sn��sn��sn��sn��sn��sn��sn��sn��sn��sn��sn��sn��sn��sn��sn��sn��sn��sn��sn��sn��sn��sn��sn��sn��sn��sn��sn��sn��sn��sn��sn��sn��sn��sn��sn��sn��sn��sn��sn��sn��sn��sn��sn��sn��sn��sn��sn��sn��sn��sn��sn��sn��sn��sn��sn��sn��sn��sn��sn��sn��sn��sn��sn��sn��sn��sn��sn��sn��sn��sn��sn��sn��sn��sn��sn��sn��sn��sn��sn��sn��sn��sn��s�k�o�k�o�k�o�k�o�k�o�k�o�k�o�k�o�k�o�k�o�k�o�k�o�k�o�k�o�k�o�k�o�k�o�k�o�k�o�k�o�k�o�k�o�k�o�k�o&`�&`�&`�&`�&`�&`�&`�&`�&`�&`�&`�&`�&`�&`�&`�&`�&`�&`�&`�&`�&`�&`�&`�&`�&`�&`�&`�&`�&`�&`�&`�&`�&`�&`�&`�&`�&`�&`�&`�&`�&`�&`�&`�&`�&`�&`�&`�&`�&`�&`�&`�&�iQ,�iQ,�iQ,�iQ,�iQ,�iQ,�iQ,�iQ,�iQ,�iQ,�iQ,�iQ,�iQ,�iQ,�iQ,�iQ,�iQ,�iQ,�iQ,�iQ,�iQ,�iQ,�iQ,�iQ,�iQ,�iQ,�iQ,�iQ,�iQ,�iQ,�iQ,�iQ,�iQ,�iQ,�iQ,�iQ,�iQ,�iQ,�iQ,�iQ,�iQ,�iQ,�iQ,�iQ,�iQ,�iQ,�iQ,�iQ,�iQ,�iQ,�iQ,�iQ,�iQ,�iQ,�iQ,�iQ,�iQ,�iQ,�iQ,�iQ,�iQ,�iQ,�iQ,�iQ,�iQ,�iQ,�iQ,�iQ,�iQ,�iQ,�iQ,�iQ,�iQ,�iQ,�iQ,�iQ,�iQ,�iQ,�iQ,�iQ,�iQ,�iQ,�iQ,�iQ,�iQ,�iQ,�iQ,�iQ,�iQ,�iQ,�iQ,�iQ,�iQ,�iQ,�iQ,�iQ,�iQ,�iQ,�iQ,�iQ,�iQ,�iQ,�iQ,�iQ,�iQ,�iQ,�iQ,�iQ,�iQ,�iQ,�iQ,�iQ,�iQ,�iQ,�iQ,�iQ,�iQ,�iQ,�iQ,�iQ,�iQ,�iQ,�iQ,�iQ,�iQ,�iQ,�iQ,�iQ,�iQ,�iQ,�iQ,�iQ,�iQ,�iQ,�iQ,�iQ,�iQ,�iQ,�iQ,�iQ,�iQ,�iQ,�iQ,�iQ,�iQ,�iQ,�iQ,�iQ,�iQ,�iQ,�iQ,�iQ,�iQ,�iQ,�iQ,�iQ,�iQ,�iQ,�iQ,�iQ,�iQ,�iQ,�iQ,�iQ,�iQ,�iQ,�iQ,�iQ,�iQ,�iQ,�iQ,�iQ,�iQ,�iQ,�iQ,�iQ,�iQ,�iQ,�iQ,�iQ,�iQ,�iQ,�iQ,�iQ,�iQ,�iQ,�iQ,�iQ,�iQ,�iQ,�iQ,�iQ,�iQ,�iQ,�iQ,�iQ,�iQ,�iQ,�iQ,�iQ,�iQ,�iQ,�iQ,�iQ,�iQ,�iQ,�iQ,�iQ,�iQ,�iQ,�iQ,�iQ,�iQ,�iQ,�iQ,�iQ,�iQ,b���h���h���h���h���_�I��H6b�X�m~���_2���'-�X�'���R<!Z{W k�?�Ū�|1�q��BRa��h�������������1�W7�����R_1��:~F�g���b�u��J���*łz��o��g�̪㢖����,�%�'�
�"|�����8#~��q�J h(x7�J>��h�%�4�r'x7�J>���}?�N�Jv�^�����A# �������z��#��Xy�{i�Çc���/�r:�/Ÿ{��1��-���1�5��h�-e!��R�������h�c���cb�����|�rXl�?�Ū�5"��+�O��1��]��
�8��h�Y�cরh$������yTΩt� �h���&�1*"�������% ��vȰcC�F EGT���C:L![�QPۼ2�_��s��JFX������p���v��t�ӸF<�I����JԴ�C�S��@�&N2-���Ng��H;A}n��������+�~��>�������8���`CPT��Y�h.�n�֘������TJ!I�J�+2�Z�:A2��+aCP�0S����#�B{"���R��PaCPg�*5A2-�}�Ogʨ�O@�P��p�Z�nTԠ4�	�=n�����O�H��-�\
�4eǃ��؊���	��n�t�`��S]T	��]
�A5������Ny�*�A�����)��ÛJ������N�:��I^�ۗ���A]�*��?�;j�8�&���t9On�qT��2������'PCoe���A]
c�H\W�Gx73�s�t�?�Dx73!��t����j1�#�}A]��*��(�܏A��Y���Q��t��N���Z����K�A]��D�$d�������\
�'�bȑ۪s�@������B�=-�~Ska<�⵬�'�C-��O��M��6\8P�I��!;�)u���0�������=-�iRhaGB�⵬���C-z�F1�ޘ�<v�E$�L��Wv�����^2"OO����R�:-�~r�:-�� ?x��ypٍyp�
-��I<�2Z ���1P��Z���p�3����D 1�u�n��1���A"�g���f��Br�"M~������05�ĸ�a�o����ƣS�y;�8�V���Zl�SM�h����lX�B��Zx�Zx�Zx�Zx�Zx�Zx�Zx�Zx�Zx�Za|a|a|a|a|a|a|a|a|a|a|a|a|a|a|a|a|a|a|a|a|a|a|a|a|a|a|a|a|a|a|a|a|a|a|a|a|a|a|a|a|a|a|a|a|a|a|a|a|a|a|a|a|a|a|a|a|t�l0~�h�N�]�W���yl��k��Mm!���`?`İhl8SmD��j��i%){~-�b!kgŐv��Zk�~���d������#a���U�a|^�	���od3{i�}�g�1x��|^g_�GӤ�zy{���dD)�o5y�c�Gl�Da�GP���.vW��ш�.��ⱤP�a������y\�>y�����1|Ί����w���H�}zL�Ͷ��bo$�{�`A~$Q5������,�\�]T�`5�����U�,�|`ͧ��%c�\��b����c�D�baF������ =���Z�;����`6t2���ϋ�Ws�0�N���� �_2UѦ<���}ɠ�F��3K�Ӧ�<��;��փ�eg�ԑ��ﲃK�rH�Ҟ��C�E����Ro�P�`?�k����� �_2���=Ce�yp��c҉'^+o��-$�Ҷ�2��?�%���ӭB,]A�N0�r�V�B��Nи$i.p\颅J#vR��~�\��L��ӍO�6X�==��U��c�����#�J���(��Ρ�01Fʡĸb��#�/��-��f-�gXCg?��ǋ٩��NI�Z���,ʬ�����w�7���+�.�E�/�!��J/=LN�ۈ+�&kp�5X��^��1	-h�HL2����!����\y��k;a�D�5O��N+-s�����8��"c��,r�/Ӄ2�׊������6t0�=(gV�@ص+�/���!�S�6+��Ƶ��즍�7	/w�^�h��z����1��6]�7�̦+��>J�|[,���~����c�;tl���+��흝�)� �ҋ�Bݴ\I �m�+����P��������Y�ڬD��R�.��5��X���5K�Eڲ0���}8N�.��א�|p-I�����/�˴a�\m /�q�,���R������<���3��"/B�0���ʪ�t?�;K���`�L��1���R�?��>.U�_�+3`�'�T�5j��Ѡ1I�O��Ʃ���>�`�D�G5��t���۽u6���^P�22�F&�������4u��436#浡�IK6Ý�	x5��6�^�wư&.�c��1�W�E9Kj++��k��౗;R�K6�}� ���ș����,`�QE�`v<2��M�|�gV�.=
I5Ę�T����g�*6KH+<�����>����h.d6�R��`5��4�b)��>I��_�+>TMTmc2=jg9G�~ahK=�|�lz���{M`h�4:���l�����1�����3�U;y43�=0k�ϫVC�M7���Z�:ځL�;��t`��`��l>�)#�޻�ș`5v�f̐~����ٓ�EG0��G�X�9�a31�e�9���[iV�Ӛw58͜�1�2���2��h2!�M��,o�Gm�s27�Od>����f^��pn�Q�M̶E5���c�L_c��'^�.�%ߒ;��1�IRK{�4���J�]�Gk�C:lM6]s�t�4+��Y(���4��Հ�EYM6?�`a�oΰ�:��|�#�2�:�?i#3
�a�bϔ::��� k��,tw��	�2F��wc)r��fH�M�z�~mO�/m!2��(d��4c�'�k�RZ��A�~�2 ���r3N��nMa��*����zk�1Cxn6sv�jR=�����;D3>ۙ�RF�1��`��t����9 �ݶ<��U��ɀ�4��m>�ؓ`�<dW�4��gή�9��1'}=�gaU���y���+K_����E5��M�|�o;�@aj���Ӄ_�X���4j�4�b��Ǉk?����=��� �5�����L�;�I��3�d��LK�>�6He	�Ţb�E
*,�.y,E����M6n�M���a+IK`+x$���`�RI�5Vv����F6�wMV�*�s�1#��b�>b5]����5C��9: 'd�[�M���9��w�`���V�M���n��b3�A����`5�9�?�A(��G6�(ݢ�A#>{M^N�`5�i;��jH��6z��/�'��O�}M6I>33H�[�U$; /�2���sF�E9K6���:el�Bk-8��/���a%��U�;����.C�:cY�K6eF{m]���2>�I�����lM�ɯ���k[
�UO�2,'b�?}4Ӫ[Nm�M\�������1R���6�5��jV���d�2�Ko�UA�2$��i)�x5�l|�Q94d����Ϯ9�5a�}��R���B��2Eՠ1i��O�9M����ܱ��M���2�t��N M�|5p���jo6<������UN��55ݵ1�.���nj�J*��E�o��lS�2)�ޤ��sY)�_�U���n�}�]'.�1G���q�\���a���C�(Rz,��х37`������Q; pcńs2-�(�4��1�[�T��4zN=-��M�XŹ��"����a���ZгLȋ'��ן���<�w���cb@�_!�g�>���ý���U�݁��@D��V�%��w��ϵ^��	v
�e����y/���G=&��{9���_��w�? `�>[	�U�iG�SZ�|�	Y���̏К6d���n�� un�d�2@%�,x2��j�� 8@C�C�s���$����O���F���i����_��$���@�T�}$T�O�DOǩ��.(�}�������x��
5���5�<��Nz_�lަ�z�2���z�K��qS�8���&�X�RK��2�ʅ� ��(X����<�����5V�L�j6��4
2����[�?���M&�@�ԋ���^�~��U&ۄU���ܿ㩚��w� h�����}n+}%��U.|g)�[4�����t���W�0���
������^V���#��bU�	����u��O�Ϊ^
���{昶�I�5Ǣ����,i;��:#(�wP�az�>u�/�����{AY�
]�c2�S�����k���l���uE�R|���drC����!����4��e��U���k[:q�j��#d#F�����F�VP_�Bm���[�§r }���5�D��)V���\"F!䛦q����,�0S���[��&�R�;cpF�`�ҩ0���_Ռ�O�S�� ��B�[GX��}���^rG�u�}�_��,Ssj�?���ľȪE���^ƅw�7y��{�*	I�nIɪ^��owC�yϱ쵢J��k���M������_f�%ϒ%�G0[;dI(��?m��n�xɵ{p���<�p����I`�L�LI����gԆ�w��4�_��N�s���r���n������f�R�7���*	��n~�	|�����`��}
���7Yç�-�N��7�9��ı��{��[]�a��}�#fO������e�����9�*Ϫt,��F��r�����C���@nh�O�"zF֩v�/`-��#����du��[�}�{��K�Fڽj������\�Իv�W�[���NJ
����m���=��~��ާ�R�pluT�^Np�0�~��}�� @�i�ϪCEߙ�^�[�'����wu�d���Βͱڰg��^rG�B��2._���v-��	9���̪[��M���@=��q4I�
�آ�4��Y�pN�P��t� h�r���C﷿%C����²���'��V��y �J�$��[{��\�Ge�}^&�Yϵ8k�S����W��\�E[�w����������Y�W���@{����$�_�-y��ZJ+��CJ⠍�}�l��Ɠ���S
����3`�� ���ԍ�%��I�,�4��@ʂ]��t\���u��_�=�-Ϫ�k�&F�	s�↡��3��L��n�짋�ˡl2L!�[��?TDU��,;]�B�������b�	Y����R7��R�'������T �w0�����TD?U�?����}	�u�����A�e��Å }�d2I������ϗ�]��	X�da�|$7�~nn�ɪS�ɰ���g�O�T��Z�D�����m���~���%+Io��o�Wa�տHT���� ��p��R�_����E��:�§�%�`�_�ƩJ�ٲ�����J�}�\���o'}I`UϪ��F��p���좡��ߏ+�։GϪXU7��_U�L��w�[��q�n�I�}�a}�����}�_Q�*�8Qr�_
�n�������*�v[���ZoQ}/����dr7�p�i��ό����c��VS�(��/�[�]O�օ2t��~A��w�Zjn���DW��!�]
FtB��D`�t�U�l�il4y��U������\��P� ߉�C�֢D���T~`�l�C��a���g���f��w���佶�3����G��#�E{!����_\���x`�BD��%Q�[�����1�\�۵-��s���,�\(t*U����:�6�IF�Ϫ��ƹCϋv��Jn�-������ז��� Ԭ+������M$�N�O`����Y�j�,gY�M��T�f������Uj�����g�߭��4�_���4�\G�F��w���V'�I?��q��̏К6d���n���`�uG���:j�w��@�/�+��Ϫc�
-���[@���dl�$�̋�QDGM�w�����ԵQ���H�����r�����T �w�۠��r����R�[�Z�J��ʬ�m��W�3�˺��}`�\�<�J��C����so��,Ssj#>�(�ľȪ��q\J9���I����p"��.�j�xӧ? [��������F�vy�o�xt\�����]�z
�χ��V
j��rû�^�s��\���>���W�w�sO��A��Y�>L�M�>�����t��z���17|�<)�y�f���|ߔ��;��*�@~��8�Ϫ}���o��z�⻴�xw���t����/��]k�\��\���C8s�Dt�o��Zhpy�~�x�����P�� ���;ڵ���?�������vL�M�ĵ�}n���
]���^`���ҷ�NڧL�g!�b!Ǩ�}������]7DB:�EݭU����§*F�����b��%�����r����{�*	��&n~�̸!S��-�e}���=�+}A��x�F`��x��v�$���X��K
��g���.���G+smȊ��9εou\���h��>��}��v�h\L���<�V�f��lw|}�~�ߧr�E�/mFO�>�@q\ U]Ac
ӄ�ާm�t�F8�6�\�8C�Cs�@�9��+}�[��[�%�آʎ�������wݧ�U��T�tӑ��=�Z���HD���܅��uH��B�\2s\�p����G ��N�E1�H����@̙��{�*	��}o�Ϫ��a�@���2�w�u�<����S�����L%��b�YI�����_}o��,_0��%�Uj�b�E���0�E���XY�l��d�#G:�k�nR�rD	��{�*	9�&n�ɪ}��J0Em������YT��y��X����OpB�?�&�H�ʵ.�����ݎ�f��-������S��eV�ܕ�o�h���s�X��O��Ϲ4�c�C'�9E|���̪�䆂3�:[�U���t�SG�l�݁k������{�$}%�� #
1��A��t�Q����;[�/Z9���D�m�W��!����^`�eGu�[��[��}��	,���yS��Ϣ:�r�E2w����R�
�sA�|����u��(?�B\���v��cp�+ϪG�`tS}݂.diϏ�FY9����M#��(�-���:�\o��p����pΩ ���CϪ�x�0t�L��f���֞���\�����l���vK�%�'���aBA[Q��-�~�-���:�\5��͢���}VL����,����T�0mC|�É�U��G�m��"���3���+֢{�@u��ѵ����a:I޷�A������Lw�u�i�L���v�s��$�ȪҖ��:�v2�����%���#e�o�F�1��h�T����_���p"��N�؀xϪޓz�~4�T�I��L�COǩ����$�~�Җ���Lw2��i��|%���ө�o�F�1������������8�К6d��S�x�2�����wյ-[�O�COǩ����$�~�����,lw2��j��\���W-��՚F}���k߿=��x����X'@4��[q4��j�Rs%�w�N2���y��׻��o�_�\��N/>ע�a���g��Ϫ�ʮ4#���Q\�����4����(����%��$��g�5����o�|���˧�Q�0�]��"��D�j� �ݝ_�}�S?��.QՓ�7��R�`�rk$[M�bK����IU.<��Ϫ��<�;Dɽ[62\��x��z��X=⩈���9�圔[_��D����G��!�X"���\�^��c�ə�F�f?���k�p��;���u]�w��_4��ԓ��`�Ϧ�ǩ�r�Y�eNn_�
���줗�u�4��z��̪PO���%� ����W�[ȸ�'���[}��xHUB�a>�&�H��}￦F�b�-���c���@�B�jκ_��򔕡�_��<dt�S��a\C��٥v���do�H���=�� ���]%_n�ʚj?��%��ձֹ`f\vA�U��]h�V������bw�G	�����k0���|���ӱ[���ʘm�"Ⱞ�v	FJ�̪Җ��:�v�u���L�COǩ����$�~�s���,�w2��j��S���Wݮ�o�F@�1Iq��I������h�*	9�؀x}�ޓzy��2�w�I`�L�COǩ����$�~�����,�w2�����\���W-��o�F@�1�����=������h�*	9�S�x�2Q�c��wյ-��L���v�s��$�Ȫ����,�w2��j��4�.6d����FϪR���j��u����K�g�TE �ǅ�)���k���w�������Y"���Ϯ4㷧l�mW���^��[A`�JR��Ԭ�x��w�<Q���,��Sw����>"�A�J�שl�&����6�LbՀLVH)�դ� �	���	�P�b|	�`#�8���|�g�G�	�O�p��	�j���+�w!^���5��	���x�	��W^��Pc���juU/��q7���C9�g��F�{&�3�J#��#3���̤�$�Ӹ�֊�����~V!�#	�ՙ7��S�_�������t��Tq������p�̪���G���9�W<W{�톞s6:����-z��l붮*��9�n	��XS��N��XPKh4������#8��S��?����T��*(�e�hv��Tc�Hd.��W���0<�yx���	3�
	ǳGSY�W�?S���C�0�~W2v����	�`t
��[j��p^�̝64� �]+	ww� �#R�%������S� 4��2���>���CΜ����&cn�R�D�F���&�-?�*��~��)��>�>{`�m�x��y�RT$�͊��F���*�p>��q}*�	r���"�ra�#�y����쩚4n^�&	�R�,�o�X��l��4�tD�$����N�	6�-�;��ѧWL2�9��h�*'V�	�pw��Ģ�f�$��k�$�w��K�ٺ��#Nt���Z���2 �sx	�xr�N,�|�7��B���B)����վ�5\�S��pȫ�����P΀�>3��,<Ճ8&�k���0�L���5=TTzW�c�$f~�W{��B��KD1����,x��T�`���d{��춡*	YG��s��tnXF��c���	�6����?���$�/���;[Z�՛/Tv<�D}T�ο%{�8�JەtF�	)1kW0Ď`�@�q�pD��A԰E��mrt$�H�����ھ�x���������	��W��8�;��P�r���v*K:��|����,�	W%�ç� (�����Y^x�t��G�	T����g�F7�W���;R3�aA�$~�8�����,8Ŧx��J�Ɋ�Q��j��.���UH���?%��*�H{������#eT#,4��i%3�5���X=c��������TӞ�UZv���]��+^b�O ����yc�$�����)X¦w��iYy����	c�I�yD���V��#�R��P���H{_	�3�"�f%��c���?v�:����*�)�	I<?Eí$������pF��l���c�t`6T8��|(K����Y���܆�eO�:;'�"_�� �o�����>By�5'T�A\>$�C�2y�v�+p���Ri쩩��{��춡*	��P�{���c�^{{5��X�It �r�o������_���� ���o��֝���\§fV�h՗Bg��	AD�Q�I#sIX�7@Ԩ�	����t$�<Hn���)�T�?�pT[�x��P��l�tt�����H�R�>��V�# z��{�n	���~r�d�y8��P��~T%Yϕ	�^	�~����m$S��hé=4���TS5�!�!��	�6z���x �E���S���Y�-k��8�4��X��Ӛ�4i���o�Z	�-pjx���U�����0�`�+Cy���	�?:fo����S6�֜��m�L��+yv��j��	� l���N�i
���K-^Ck$Cu���r���J���{��[U6}�����%�����־���	�Tl�$���F���y�7���
����G��%��a;���TE�$������W/Ŧ$�"��n� ��k��.�+�oۋ�o)�$��WV��J�	��%Y�y �[%�xi�l���y�I�{l� t������29����Eޙ����#�,���.��:���"$��5Z�����I���w`6T�os>$���w�����?y�W�ӨΊD��$��q�?r���i��s��vrTe*���y�j�Y��S&��ڐ�����"��]���������z�8�����	b�yx�W$-Z�AH���T�����+6e�W�2�-$�q]n���a�׺n�4SM2;���8q$�<c%�"����۪�<;"3z�~M������i��i�C�m�hLtN�+�0�	x��e3�`�[x �C׀�斅�nb�	q�$�D�Lcl	��>��8y'�y,�v�	��\�$��1��κ��7�
��3�M���&	@5�]R�	U{��~��`�O���;�$����5��T�*�I^�?�#���Q{n�q�sN*z��z-�"��\U�s35�oƩ?T�*���̳R���k�'l	+���N��s�|	�=�%����B9[k����ٝ5�ީ(��ic���Te̃]g�=',��V��$�y��U�Ro�YU&y��Wu��l��AT�M���H$���N\'��������P�+ճ����	��q� �0�G��sY;���X^�yM5�n��Q��B%YYH�$���b3TV��{�
	#���x��26��$��S���V��q��9y$�msڱT�	��@�k�t;;�F7��4@#�(����S��� �Q�׋�$�	�����FFT��P�������W3�Oܱ�� *Ȼ�,���I��(!a2#Z�CX�0y��¨i��X{O���T�����`E?}��ԑ/ ��G�F���	�T��հ	�xH�p$1VW1P�ͷ�6��[+�x���$�5��(�!Ty��|�{N
�춡B$��z��-�%)TvP���wB��"�t8�>�#��S��i��ZW�'	�D�R��6��A��P�;i(�(M[�T���	`�<,/dճ��,���t�E`���H"g�	�4�I�T�\:�s.�4�G�h#�3{��춡�$��P��Ƀ*)	��7��3�	�+6���4�:���֊�^g'�!<yA���	�o;�"��N���EC`S>U��W\Y�������l��Z�I���D8ӂ	8��b/�m��#��I"��_%	?�\�{W��Wt|`���E�<`��k�#R�,�M�b��_�֌�v�*~��Z֛�T���=�I��Jk����̧*�y�iayV����p����/�����\o�9��4{��춡*	Yz��6�*ե�o�t���Tl�?�$��؎���?�(*�	�٩�g_���ۓ�3 Á�l�Q��Wl��*�W��g�7�>$�@����v�HiT��y�i�$�G���,���B������Egì���c¶�La������δ�k8��a}��&UtC�|�oS�@�£M<�a���h��Wv8Zڭq����U���v��;iB���BwIB5�7{O�`�}ER�R�Uw�����S�K���o��-�����ɽ��������e^�G;lU��K-ȑ�W���x��P���l#�	�w���b�c �d��+>䪥3��p$�Ƚ؃������ܤA7	���#�n	Tf�JD'������1�	YdS�uk�/�u�*��<����d$y��Td�$�5ΌEl'�����Š߽|*�S)��	T
�nVTj�� *���o�p��@�e��xł;��v�h ���N���T@�ww�$b�	�GI�¾�����G¡�$��E��x�g��	;��:e�Ү$��o����< �5��"$p}�����P���fc���T��(�5ا��"���z�	�-��*��By�Q@\!$�^t�,��q�G�JT�tR�	)�k4�tAe����x��BBT����:�	A���5؝xL)�h� ����x$��#%A�(�lB�ϩ���"���NƢ�Sv��T�pT��Zo��*� PX"�_#�W��!
$obb��|	����96�x� Ux8�e��,yʾ$,��?�^�i�'TrjT��o-h�>y�M���t�	U% ��	ҧw�c���d/�]}�,��Uk#������W�#/��	���lo���FI�"�\^+]��9�����s9²c3�n���	3	D���0	��#�Y��7�ߓ	��: . $��;��Tr�k#�K����	�P Z�
	&�4u�q���#�p��U�7o��&y��$f����	,�Y���qRXra2 s��K9 �=����@���		Q�N3��	"�	7�TͿ5%3¡\I)�d{|W�m�$����uHw�E����W`T$�G�#*?��݈�P-W8Tڏӧ���	[�$�54:3�Z��4.�E���SB��~�W�(�H~P�u����|s�����)�	I쳢�^�	5�Q_�6HϞx?¨H���$�	se(	3.�H�?7̉-���6�f_с�����E�� ,	xh!�4�E6X³�fc	O�T��W������l$�Bء�cV&,�	l�l��s|����畳����` =	&�ZR!{����W8?���T�q	h��	���>���.=c���"��F�͆�xpT�#��e�g�/��m�)������7�\����Q�	C� ���ȖnS)Us�f�IHm���و�y�>�27�XX8 rT}y�%�����%����?������56��i�,�ӹBè,����k6���T2qp$x�x�P����&� ��v`��$������A�#�������?y4��j���c{N
�춡�#Q*Pé�b�p�NfƔ�U����7T$�C����������,h~�TI.pj$ 5�T�*�xWC��(�
��W4O+(! W\��k��F,�1�����	е��+�7\��3���7�)N=�J�9#5ȷ"l8�(�bl�8pi��;�'70��`;9�i�3��^�ǔ>��@[$$ @72j�iQ�²38��s�/���2���T��)��`IYy�[׷q[{���2���
�T�7tīXꟅš nnD2^���~-��-ڌM�Ӝ�S7�����uZ�}��@�(�w������P�^M�V�Y<���!����������p��󈕝?Xm��r-��r��}������0�cE�#�z��T��#�x3�t�MR"�!���������r��K��Ѱ`�Y����i�ҭD
�R��)퇢��Г�[j�S��@뙮.�f6���ޑ��S��5�����Uv%�_8��y҇����C���Q�܈���[��B*�������R{�5ჽQ�����
�p߇O4*�{9�'dv�*T�������f}��������D&�+B4i�ڀ�m����<m�ݱ(�b�$Fnܝw��ݜ��X,p%1��,,�A��}�8W���	7홏��s#��c�*���r�*Q�<4�D9&4ݜw��tk�{Z��}�|���cP\���US�r������z6�r����+h��ݜQ�)^�Ԝ���� �2�L*Jt���zݜ7w�w� ��� @�V��o�C�0����^O=��g΀)���#%}�������Ve�w� �r������������ڲJ)A���є�P%��`>���d�M�ful�^��R��^�(/�_}��%;�>����wZ�~�Z�Έ����j)�lU��K�O��5b� �g��^��[���ㇽqϦ�O�6LzS��1s`\h*�^�!�y���}�M,��
�����b����7|}\���SK���D�����3+��i�_�qD'���B�2d��Of���B��^�m��kZ���c�j`�e[aZ��
�R�'��Y�`-^�[��*X	���������tQ���
Y֭5SHĜ-
�綧K�^w�Z���a#�S956rZ@�&f�Ç����5EZ�u� s��d�B���B�x� �m�Ƞ
�ޯ����c:�ć�-�է�XS����6�qD���-wbݜ]~/V�2ć��ć��8�Kpjx���B=���&�<�G�\�;�S��Y��]�w�[a
�ݜ)����xc�^���S������\��O���x�[Z���H�.9���fx�8c�DT��ӀK��"�Soi/��諦+�M��5T��. �M��iz\>�^� �+�	4P��Tݜ-�ׇ��V�^azd����j]B��Y���]I|�rPSoi/����fx�8��5T��.��q5+}S>� ��+�(�%P��T��-�ׇ��V�^az�����W��u�@�����]I|�rPSoi/����fx�8��5Tߜ.��q5+}S�>���fx�8�AQ�ۜ����T����jm���az������݈V�À�5����e����6>�t�H,��@�!�X����4�v�K��4θ-C^��rAڜ-jׇ��V�^�a�[��&5�0�������1�xPt�^�-�r�f�rU�~I���s�M����:M����Ӆ�bƇ���:-y�u8����KI|S$�Q{��~�������^���T�����6L�E�~�O����ޝp���v@"R��f��O�w������K�̀8����A�p��/T�H������W�Od�hM���{�����)�Ӵ�!�����Ѯ �~����Y�/���J�<��M]����K9�e�R�>
f��C>����y�9�М�*<��2��r���yK�A�p�QK^��d��^,Zړ��+$�%����绞1�#�����r0[|���l���+mm�3��R�W�n8�đ�.��[�¯3Q��f.�k���~}ε��K�U��z��9����)�=؝�a摼��a�`�K���C�x�h?�����rG��Q�tK�Ό2���Â�b���`{��ˋ�ɳ�w�K#�%.��C�����j��[���Go�>K.o��_�oq�w������rG��Q�LK���J������-�Ү��~���ZY�/�����1�h�[�ѳ�_]6a�	K��7H�o��!��������Go�>.x�_����L�i�9Ϯ��~���ZY�/�����1�h�P��&n�=1�.k ?H�o��w������_G1�d��K���0��$+�yh'������ѮJ���"��ìH�ƍv���Kg�� �`v�SŴؠKU9��y��Z�"��s���Q���&������K�;M�H��e�Y���U��&{�a������kT�(�|��-��,��2�T��VČH���J�<��]��<�(�L|��Kщ��������j�X>D�����&�8� �RmK���"�L�/d�y���̈́�6���J���m����E��),���_G1�d�UK��H����@��t�
a��,O͓:rR}K������I��b3��O�E.��#���@��K��j,/���d[׊���*�b��"�_�Ǽ�u�ad�6�YxJ};�!jA4�����-�ml�a�1��Ba�IǊ2�_�C���dKԓk���v��5�J/����kw'n@�IC�MҤC����X4��l-�0���n���몍b�x�늊�/�L�p�,ȇ�,n�=�T�"z��uV��QK�tk��=Tjm �~Af�ʭ}�H֟Z�����;�Ѳ�iS4v�l��᚛��8�ܞF��8��#O�������:�.R����V�&�k֓qut�u�z�_Un��	��p��e�M����)�ĥ1V�X�Z!����Mh�B&D�����ϤôI��m�)���8�[��i��n�e�o�#^?"����B��g�-6����j��eY�犡K{�4�)���/�zp+��δ7���DH����H����-��|zĥV�)�BG@�u4�`��N<e���3�L!q��#�/�,k�D������5KT�6���VR�C>4�ybХ���K�-b� �Z�J>��{�d�wM��]�%ʿ�.n�С���L�v�8�![�+޺�y�:�!B�$u	�!���J�����C��V-%��.f�V%��f@����m�HG$���ۅX�K�E��
�p��&�|G`��kV�]}g�
Ϭ!���\����m��/�Ms�/A��І�(��7��ٺ_�!7_�v:҅a0ކЄ�1fg��GAj:'X�����@ZύI��[�_���2M�ͻ����𗮴&�A�$Cl�� H;���*b ����RdD.�xt�!�iMM�PJ�ܣR�
�6�lՋ ��؅�f��9�wK�M��b<�	F�J���=��9��9}.Y�i�!U�A^����)8��"���5���ۍ���J�|�y�[�`CU?�jV_���'��A�����_g�El�d��"%{O]����\ϒ���Hɥ���dѳ�b���(�t=j��L���p���%��U�0j�����=��o�Zg�Elg�R��Rw �T1�O����(X-�p���L.%��I������}e~{R߇&0�I|>*�s��?��	�zz��&xTS�U�����V��v+F���BD���0>v�t^�o���hw��Q�.��lÅ_*&��E��G$م��d�8%�B�A�%%�/� 4�R��}����U�R���1�1i��R4��;E��� �.����"����p�uգL.���Zv��?�l��>��9�9-[2��*ۿQu����sRr�c.~K���\b@�B��.2�>�M�r���E.қ��a��[= �-�u��O�f�������+;��c@��'��5gn����n-�W��y����������.o�p|NV(ҽ;.3��5�X������[	��xb����0օ���c��Y�r�%�t~ԩ3��(�O�.T��.:���e��n�i܇�ATU~�х�׶���&�.G��^�d���^���vh�`Q�)�rb�Zރ]����`;C���J��y�3�<����}A������.1U�@?v���c�Y�Tm�֣eNz~?g.{.> �PK4.��?�v�/����{3<���$+Ab �e�Jv���-�QN������ڼc8Y��B�UP��Ѡh�|��#v�K;��T����|����ȇ��.�E�$X����*2&�.�~ӅD�[�ЏÅ��߱��!ӹ.����ęM�U"A� �?+PbFf�-�N`���D���?�J�j'�Z��B�Uf�LOL;<�)��I�'��*=��E���>�r��.�F����j{4j4D�
}<4�v��5����v�l����X�a�
z��Q^��ZJ��s��������xM�U�����R���V��\�@��r�.��-����RŨ'�`������.FKh*(��z4�����E�����ơc���-�?����*�.�Ӈ��.K^��9
0�Ps8�[��4��$c�v��H$#%��Q�l�U���?V����-�I4�癦�za�b����i-�u������������#%��%�t�ef�/�Ś��".O�'��׃� .�	�'���.���JII���H���D��J�����vdg�.�<� �.������/�,����c��.��/����?qU�3=*_��Un?T��,eǸ��m��m������'���"�^�'y����w؁���ԩ�u�=����U�3�i@ڸ��/����3zUCʶ/��Sc�I2֧�Н@v��ΌN��Q���U��
/������.���� �Ȯş�.ˠ/���n?qU�3UU2��.�6y��������/T��˳��$���D9�D3 _l���("y��.]<�Sv?�����U�3��p��l֒�Ssn��?hU��\/���9��.�������ˮ@��.��/����?q5�Rg;������Xs���J٤3��.�y�����	��.���	�*�����\�S����ʩ�u��.m"��3��^�d�����L�����⼮9��.�\/���L���^�.���@v�V!���'ov��.#�3q�ي�.]d��]�(v��.#���?qUv?U��f&	�J�.7���qDI<r���m��6��.���i����ˮ@��.��/����?qg�3rS6�����!���ve��k��X�l>1jVr��n]��S|".e<��nkCe�%�nk���Tc?-�>ͫm)�5��5�ݾ�;�xgz������>C�n�2j��cgz�B��n�!�1/��2�1�D�B�n��Ґ\Y�o(9�SQ_�mjer��n]]�S�".D�"j�!j���|"Ac���T�[j<a$[R�B��3B�Q�k�KW�rE��G��5.����W!D�v´���Bs��g��^~tqP_β1�]fC��nkKj�r��n]��S�".D!j���|"j}�|"� �Dy>��1\C�.�z��ax�W"���>1-�D�C�n��ҐTYȳ\���"��;!*��4Sn>1�#Qn�5���n�2�M�9b�����qo�K%�HD�6J"���qҷ�i��2��6�@ݱ��캼����<��b�)��2�D�C�n��Ґ�Y$�|jbr!�nC��nsʷ���r��{'�<U�^�h����BP�n����2/3�1�D�B�n��Ր�Yj�el�okK�>C�n3��T��[\��#�ҷC7|��
T�"B�p��n�.��2/�5:���ʇz;��,�D�C�n3{���?s�C�q³��yCsz��*�׾��z��Lkì��D�5�)�V�"��gz�����f�\�nkC��n�f�&+�3�1�D�B�n����S|".n�"-��B�n98�����B�n��ՐD�g���V�-¼G�;�-�ۜ V�c��� Z|9�p��,��-*�]��wu�A��j��cn9�#D��b�-��zq;vF�f���w�rF���Y��wF�;�q�b�E�R�Q�TF��b�\�I�LWvF�A����W�觏^�����U%������G���*��;v�5�vF���u;vFy�j�\�I�LWvF�)�����f���wF�;M�;w�o��V�-���8WvF�M�]��Qr\F��2�\�I�LWvF��A��;v;�raz���!'L]�)l��~��_�9JWvF����;�J��a�#y�u��a�uwF�;i��;v;��rS"�{�MWMe�;��a(��)�a���5}�2^�'|>H�Cn�dxU��V��-ΐc;va��._;var��?��0��!�-�*��;v��W��MW΂�;va��q(Z�A*������[j��;v�IW��Mm�<v:Ae[ �ћ�v�Ð��;�-�8��;�-��d��wF�;�Lr�:�E���\��_�qy�V�E�WF?Z�}L9w��pr�����MWΕ/:vaJ���-��d���n�qES"�q�MW�-��Y��wF�;�yq;vF]�����S�r�Y��FF(!�c�vF����VvF�V�����7�<var��a�H��;v9�VvF��Z�E�:�\�,s�y9���ؐ~�����E��J*����t�s?n!�rxLr��S��f���wF�;���X�DwF�;�xq�Z�E�+�W[�����љ���4�;WvF��L��;v;�ra��a�H��;v��V��-�-��[��wF�;�Cr�R�E�Z��t��Wd��������g6_k�Q�2E�����V���;v�Q~F��2��"SF�VC�r��-��Y��wF�;�yq�b�E(Z�F�*��;v�EF���p�	�)]��vr;vFWvF��j�E�Z�����8WvF��M��;v;r�raJ���;va��xG.����zq;vFB�:��wF�;��F���A(Z���*��;v��ya�)��;v9MWvF����E�-�W��]��9��k�Ȯ�]�5wF�;�Er���E�:�Q�F��:�_���OWvF��@��;v;:�raz��;�dy�V�k�|98�_ra¡�;�-�j��;vF������n��_���r�yq;vF��wF�;��-�-��zq;vF�6�S�:&[f-�/���r�yq;vF�wF�;��-�-��d��wF�;�Lr;vF���g��avF�W���:��}���x[�a�xU�@T�a�F�;�-�j��;vFF�7��;�-��W���I�q;vF��w;�rS"�p�MWMU�<��b<���Dǂwػ;vz
\�ǂw�.]woSƤI؂w&)]wJ����w�^w�C!�Ղw	^w��hf���w�^w�
Û��w|^w��ECՂw�^wF�<�[ւw{^w���9&�w�-]wjk�˓�wc]w��b��w�,]wpi�]x^wz,]w��&(��^w�/]wY~���^w�]w*��g]u^w..]w��t�^w.]w��,��u^w�]wxG.��P^w]w����J^w� ^w�Q�U^w�#^wS�W����{⣘ d_��Ν^�/F��>����o&�wS��%$f_�kκy;vSC�qJ�w�Q���;���w%�]_�(l��N��}��wFw�kF�;�5�^;��9SF��SF�;�Fy;v%�d�N�ͣS�*a_����ĂwG>vF�;�9$o:;vF{��<F�DuF���up�S�h�N��eL�`ܤ%�'�Ø��ڟ������~^��۬"�I�i��o��.����D`Eߞa�J��������[��jj��	J��K�5(��Ơ�왶a�Lܳ!��ԃ�F<M�i���a����>[������+vF�.��v2��(�I^��&��5-m;v����ԒvF�\��0ղD��C�����.�{Ə]��,vF���3���PU�B�9�ۍ{B�aqCbF�;皘8L6/,5��j*��R�o E�3E8��[�l���p9@#�z[����R�mE.�Ð�	~�d�\7� l�U1R�������ǘ�q�R��Y�G��Ǹ�͋#�x�bC��܀c�<cˋ#�7�����M���#� =�����ϴ f�SR�=Sf��WR�da��mx�s����vM
�:�/���OԞR��ܯy7��!����ܽ�%q�n�X/��ع9�f��16s���>`'.��^5�����v�{E�!���xg�|&	�O�2�{�����^E��ݨ4����5)+�`,�Z��m�e������e8�$~��>NE��e��df��e������d��u�Nc�#�܃g��e�=� /�������(�f�uX�e�H�,�fM�H�΢fM#L�f����o[��� ݹf�K3���+�a>$8��e�?(�f}�D#H� ��f��
d��u�I�e����+�a�e�����:�����������f����NJ��pg���B��e�н~����axN*8���zUAM��d��7e���@�o[������� Yݹf���e�=�j0D�K#��*��d��u܉e��+1�#���e��#���b�d*F�a���d�8B��^ma�0 YVu���e��l������>�:uH�*����nB���l�������&���i��jŦ��`w�'D�ɇ����C�2�ឰ2Le������f��������-�=)�ݡ��/���9�n"{�Ԁz����K�=�a�mO���m��WM-�`�we��~�1�#*�3�ي(����^j<_�P��1�F�,�n4�z����
k��g�������*��J��+���V0e���:�T��2<�=��n���)�a�C���H�1i���˩1�`�6�[�����<|^\Ͼ��g���ܹ�I����e���b�Eұ��a���/��hz����=�b�4w(vE~��R�赸���l�[��a�iq��8����e�r#r��XM��u����-�����ڃ�5멇����x�~u��XϿ�C��K*��:���&�we��Y�,� 5��Y[�����E�����>�O���#��.������P���{��|�<���x&~U��l���w��������^�����e����ʡ����e���ې<��؂�ۚ�����e#��bT�
���h�Eҫ����O����X�(�2Ձ��Ex���qf��P�=T�Ce��0i���</�����,+��PX�Ev�7���U����f�Б��7.��
M�z������:�@�}��1��4���ȴE���T������j:��B����D��0����j���%�X�Tqe�j�쬐6eݟcF�0���s�J�p���σ���ٕ���G�\F���Y�F&�Fe1�V�m5�b�m�0TT��	�÷�L0?͡����T�W|������F1����f`#Re��ߊ�5ژ����
b���Q�����Zq��$~­+$��e�ve�Ck��H9�{�|���\\/���y���f���ʥQ��S�����N�Y�z;�V�^���>��.�p�ڿ���,����u�=e����������;�k6�А.e�k�e�x�~u��X���i���K���C?n��X���'��ؐJ8-��:���q(�ue=ApB���Ŋ���-7�+u�K�?B��|t?����x�~u��Xo��t���V����SF�J���7q����D���VN���؎&��k'�#��h�ML9���8e�3�h����w��ӏBe�ݹ��TI�p�e�O�A����Z���(������J�UI��2De�v��UơQ$2����C ��߾�VYv���r	�&��!Ro��{o@?(��RuN�/uz��r��r�y@ͭ�qgp5��%{!('��k�g1�6����Fm���Cp1c�B��l��@l-/�B�	�$�jI�L<>nN$�gt	m$Ǥl��~��Y5�R��'��g0<��UhGe���C���$P8���R$�
l�3��s�.ᦕ`[G3�G�A�Z��g���Qhg̑�U�FK{ �L���h[g��O���Ze�������߿RK���$D�g1�l�����ͽg����dWc�ְGJ�h�d|Yk��f��f����M`ý'��_�,�AWD(�~�b� 4a�=��Kix�	0�� -��a&9��-,�"p�ǭ��!B`�a%�L,6��&��`�b�0U�'�9"��D�� A���>�_���?�DIb�I�}ݚܔ\n�[��
�k���?�S]:���\V��@\��K�>�5��&���?�2:�Y�ո��x�� ߼4ݜ�r�?{q@�I�ȴ�2@<hl6�o^uƅu�����?��"֯/�L�Pv��ݒ2�1}�?#u@�������@����Ɣ�n��@.E�����?�e�{�sA��{ה�]�?�y��͘M@� Lr$Q��Y�ޡ0�!G�0/Z�"2V&��r������[����#����P0�����ݬ�0ե-����^'v���;�줉���{�-C����d3m��U�6��Z]�_g�����.���A����7��m���}���ᮐIգ�9����N�W�}��;��}u��Y��m���{����3��)%�Jۧ��@֣���	�-_�����3�@�V<5F����ֳ������j�S�'Z�p��)����f�[����xQI6�⣃X],���w��5�C3"lDr������B�����/������,�~-�0��"��yx�������0�v�����>�/�nE����	̿h
̱<]�*�&(�Ԏ�6^b�g��$��/��$�jIm�T%E�S����P����FmV��p�L8Wu6���(4�o�xWJ�HmGt	ko�Qm�G�w	kok�oWB�G*�o~��69��Wg*����z������i�:��h:~\�^�<���c�9z0��?���f�C�ڭIڜd��ާ�Yw�{zi���(k)ؐ�t|�U uS�v)IS�k�Z���c��,��n��d8�&M��	����$�F�V�#.ouG��^w�HmVImV0�zVIXl��lVI:�+KU�J��p�k)�y�h	pImV�<�F�
�3� �b�XlW�asJc�C�{.� �lVI{.�	>P�ejsoHVP����G*�o~��P��7�lÛOlV����RlJ��RG\�Vl�T����Vv�<?���T5\���(;�Vl�lB�i�V�F!XH��"n��hDE��� �tgVj�R�UP0bCxlvC\�}jV��֢�lV�%5U�!���Hc��n�j@EHIaV�\��%)J;1f~AF�����-�~Vb�����L/��Z;�ڌ1}l��EVy�B �a���E{�<� iW7�0R��V���Fvl$HR��#��\FQ�qwiV��l'S��$mg�Nr��l���fV�s�V��jF�8��h1V�txY��V�3�r��	WVdd6H���wŃPT��~���lh��'W���}I%�����Px���#���I�tVZ���1�c2��H	���V��2I�V��ܚJ�YkB ƈ�VG��p��)Wg�J�����H 5:��,`�s�Z�^��V���}�Lߙ��S�H���a�I	�V����$�� ��Il{jVi~rN�	WPx�k���!B0jIpHr�ԈE�v�I�"Wbjyk�ɿ�"�G��}�\�}I��Vz�N�{jVF(i'��V�OlU�M�F�V�)`��k��~��I���V����c�MV�-\�3*�'���3;�Vl�l6�jlVeo:$\_���l��K�?R��Hyk�oe[V�� ��N�l�[7��x` PWhM;�X�lVtU(��Bh��l��Kx��j��zNV))Wb ��ǌ��>+�{�g���� ӷ�Vnzj|w[�f�{l�P�"��JO��H��VU{9Vm����%] U|��3d 6���V�z�{��l��pl�5���VI��V�B<V�՘I�ll~T���r��m��fV�r�V��l6��a�q���PP5��	"z�IA�V�c�gl�+�UITC���_���V��=V��o���I0NO���B�	J{W�yy�X�HVG ��2`��Cb�"-V&,V�x9lj���rAIJk6L���	2cJ�nVVIL��+��Y_mFl��M�>kH��V�;�}�����Y!�+ ��ߤ��VU?���Jl J:z��PM���IB��HMVOԧ4�����l�Z��n�X��VU�]V[R�I\3ko�l{�n���V�7�˺��V���+K�7��hq��SmjTj�V��W&j�VG"Qa9��P�~v�B�I�V�ɗ#B"2�H�6�F��G��H�l�U��VD�Hd"�1J�8K�nV����5��o� Vn�2?�N�l����qxX�W��:�F�VU��)]�V����|G�����i���7V��ak҇�eɋuVDC���l#m�V�Vu �!�����)��qh����YA~V|�6nO��lUh62��l.��2�V���T9veXX�0J�)HV总HDxVI����BlIT �g0� @W �eFlVouUUUAnh����5W�}�&��lV���z�9VP���v&�����p�G��VR=�lJZwu-o��V��k�}�V���j�ɪ~��G��W�W(=P�nVm��$Z�VP 	(�.�;W�����lVuZ̚,[a)$nb�.�Ox��z�z�H��V�{x�X�l���trH��:y�)�lI�jmVv:l<y^7fn!l�l/Hr���H���H��VlPD܊����ox��j{91+V�	W�2��N��n�m�w�ʞ���l��nV��T�EP�{e�l��YJDb��	�QI	W�H�v�MldGtOwwO�\kW��:2�
�V��
O�X=kc ^ɿy���m��ǉV	��VH�ok(�q�&0VhEFa�
6w}lV��'�f��FHXl
�c�m��
m�cVG��d5J 5`eB�9kV'�׎~��V�wk;g�^�2�MIO��
m"z�#WY�VV�p����X}7VTABr��I�`�I��VC*3$�:�UqT\�]U�y�.�3#��V��yk_��bM�In�)��V�7�����V��O��xkpד(^}�H��V��ѻy��Vz�ml�SX1� :VpR���m}ɘ�V�V�*B��#��l_a��M4��y��0J>�V���v�k�=~��~Kh�Q��v�U��V�2>�I�����l�d;O�V���H��V_��I�l1#��xGG��J��|gVk��VQ���hRZi	;VW��,�V�+<���V�����:y�)�l6�j�V��j	��V~���6Nr��vM�c�I�$WQ³���T�Ĕ}yx\pW�M:Ƅ�lVv�mlh����vIM(@���Hl�eeV|��!l;Vh���Wk<���o ��hp�V���I�b��p�+���j�h�vN�Vw�k֬kw��ms�z�C���BXJ%�VX�ks���:zlI��~U�m�	��V'*W�n(����z�V�tzF���y���H�%W��h�S���}�V�"��l�\�V%�V�B�r��vk�2c�j=V��W	�V�*����hUbi'����1�VO��V�V���T���J�He	J�VcoII�V��6
L�V��kCCr��o�V�zlgI��"�Is J��V3�{H�)Wk �d`���C�-#�2�K���y�`J�nVX�xƃ�l���|�G��Wk|�ϟdW��V�+�=��m�N"��RPR��I�QV���t3l�f��lW�d�rq��,�yW���*+��~RAUIA�� -W@�f�lVǉ��>���I�9�Kk��y��D�LV�J94H�,�'���GV��x�01G�RVM�fI�MV�/�`k�o��m�p�EV�ܗ#B"2J�7�BrT��K��lb���VO��6wQlIt�wOo}� �W^M4�wlVP��`�.����kvC.HBʆR2�dI��V�U�V=�GX�b�I.�G�Gh�by J��V\�O��skx�m�5��#jj>PV^V��9U��b��IwC���_l���VQ��!�V#��jdh7ML�IYV�%�T����HyUڶ��S��NV�njLHD7,Dl�5+<���4B+nZ~`VO���N_���  H��V����HxWLՔv��l�Ht���S��jMV��~.M�V�J11I�,����Gz��Vg~�U��[VG#3:�LV8�?L� PW���Ɠ�lV���h��6=lJt�/l��)WUs�V���#\_I�l�B�l��MH�V���a�G�	�V��ruڇ|��W���97PI�HJ^֣�m�"ek�Vj�9Vm�o=��:M2PC���Ib��H�W�ܗ#B"2J�7�I=x��l#��V%%W`�3���jU�Y���Uj���g�%�0+ VI<8�Q�eA_i�b�?rӣI�mbW%�V��<|m\%�7g�E�j�!4�Y�Vh$q�Hz|H�XuV����U��ӥV}+�1-=*�l"&�v�oll��y��eV�����EI�6Ę@'��xV��U�VS�sI����q:q�L�PW֍����lV��nl�K^1*O!VfUi��V�[����V�����J�85�6KŃFИlj�T�V��J�I��;r�m��ٓu�ɨ����JlV��~��A�HmV~<�݃�jIm�%��reyP��w�VI{`��� VI{x����]�y`���p�,�lVI{P���PjIm��Z�VI6U {]��Q����+FmV��p�\8�tA�#��jIm���eF�:�L���O,lV��P����/FmV��pVI�eF$�eL%IɼpVI�@EmV�.P���P��'���-{ʍ�-cM���_��$��y�ID^`m�d�je�lVIK�BE{���C��L<�(�pVI�F}p��y���{��	�lVI��jIm�|8Mh�W+�҇�� KlV�Q�݃�jIm�%��reF?��m�TD�m�|;v
��9�c�%�o���_�Â_H��.Pط������K3��4lV�P�Dp����VI�+�1sH��C�1s�4�|>�"��jIm��lVI}`��y���{���lVI��jIm�L8M���W�&�����j�{���lVI��jIm�l8�\D��m�|<�(�pVI�NF}p��{p���7}^e`��/I�	yp���p�,�%�e�p�EmV���j�&P����eJ�*FmV�&P����FmV��p�T8M,��WO�DVnm�DD�jm�LD��m�T;�[Gt�q����1�֡L�>� I@�T�*FO%"���VIn%�5�B.P���p�L?�)��jIm�	��eF��*�p��Dэm�DD:�m�l;�݃�jIm�%�lVI}x��{x���,VI{p�Iwg/P�$�%*�N#se��jIm���%�Qy����p�\=�'��jIm���beF��eG�*F�{HB}��('����)FmV��pVI��eF$keQ%L��pVI�CE}x��{����VI{X��ğ�mm<�8{���ZUiI&�e�p�EmV�P%M����sG���=�Չ�^�h2Wu7��lVIy���{�iEmV��p�D8M�חW�u��U�Jr�VI��]��U�Je�J�Vz�3X�J�d�J�uV�J,e�J�'�w#,�J�e�J��iW*�J_b�J���o�0�J�b�J����.�J@c�J�WB�y�p�k);�e4�[?���GF��\-����QzCuW�0��Hp�Xs��X�a�&�t'�dIm��
�Fﳴ@���D��˟�ڣVIo�ʎ2C��|���DGtd6�ɻ]��EVIڦVI���zr6�R���T���reZ<K��Wu $T�y��%��g����Z�%aτ(jIm�����n��e�cIm�����I�Q�h@;�D��LE�'����A��_mVRzlVI�wIm�ׯ�w��ǥ"���s^OM��W�O�E흮�:�7,#=��:g�n���:UH&[� D�v0c	������a5��I���Hk������ݚ������Co����M9�
��:�M=J��fv��A��桳��]Fk�G��d
`���q��E[K��+>��K��z��Q�]t�!\���{ ?S��F�w-�¾	�������:2' �&D�N,��ºhWh��BFL�H1�S��9�Ntg-��/�������.��Q�嫳ܒ�y������K<ؤj���$Wﳲz��s0AXI�C,8o�ɟ)ޓe����N���3� ���.\8<�E; k��?�#<#��ŲXm�5��`)/q����c�����9�Ղ�l��S����~Q1W���[���n����G�u�e����B�5�\J����R1o����d�2�L�!�V(��G�Q7zj�ɬ����Ī-��vC��M"�sD�}L�Q���W�6N�?<!��q��P�S�:kTP��[���¦��a���mΛk�#�L�n^����8�+,b�u_��;O�N%ԉA��7�� ]��ϵN6��8O��E�y;OE��2��
�<ւ՞y��LP��N���-�T����h�&�#�	�M�	O�`�Ǩ[�I��/
���Μ��;�SP{�������� ��0c�F�[^#Mv�sP#F�L1�;Ȫ�Y%�ԫqz<�Pڝ����P��\�J��J�Pki�)-f�9�'��WAO�ƌ�'��5Yaku�ձ?��O$��O���O��߈�*'զ�v���V���%6Ĉ�8O���C%�	XE���Ժ��i����t<O7K�Y8=o#���ծ�i�,I��?���P2�Ƒ_�Q]8��Դk�Z�S)�^PsWgPC�c�X	&����Z�t���~DO�R�?��(��ն4��O]f֖;��N�8?�����k1߱$�)-����������?2%Jw�ݱ�7p](�j.	L��f�PȱeA��kd�Wɓ�=�%Xh��냇�����[IF��!Q�i���E�|�=`$�w��������a�5�mk#|�k�F�+���,���P�U��@$�H���������:�^���|�n��"0�#�Nv�E���v~�T^�����1�Ot1��#�Reo��
�Qv���pz���3$i}�߱g��>E����+t.����s�}EJGܿ�u�S��U��`4r��3�Pg@`�����D�[㗍����$�����2̋��N$�(��s�L{��1�냞�״) ���#�mk#|�k�j�&�¡V�0�����1�<��u�Y����냮�`�H{����A�p���������0o�ى��]��T�7ϱZ�MQI�[�A��]��O,�U#�Hٱ�'1��"R��v��� O\���xO��-v���ִ^z%7���H���T���.$��/f�^�z냢He�C�r"���#���{���
��� J4!����ı �2[����m���X��1S\���-G:&��H-�K�5��;y����/H����f��c$��Ă��"p����%����C���7$��fG�?.���@X�4\�냶�UjD�J�U���^�-��EY���9~�W��A�K�P�m8SѱF��;����	�N����wJ4!"Ż����9q~2�8����"�������K�L�Ёa$�N�ʁ�b|k0�ga��YV/-�m�o�t�Q�ܛ� B!�"$C����[�6�/w7��``�Gt�N%�a��y��q�[f��2Y�)h�\#:�e�����#���
!�[����w�2���V�D��8����� N߅#���бs����0m$�����.%"�҈�ٱmK#������c�-���#} ��f�߉��#�G���X|ʄ�tfo���$j�s"�%��>�z��u^Lۄ�!w�\S�$J��(W�A�ؓ��"���Bb�J�O���K��B��H=��(����2E�\��f�aIּ���se$����a�u!H$�	gz�4���"�A���"�J��ZH����Q��"����;���f�냜h�ǋ�x$�K�d�J��`|k����B������CIf��O@�m #<�4=R�h�,��{�o���2��L�,!r�#����/��/]������x�H�b�����3㝷��ڻ���
�1랯�U���ńã	6Q�ʄȱҖ���O�Һ�ԅ��N��Y�ؘ���Ml�ᕇ!�2<8�"S� ���$��������^�C�U&����ބ�����Ą�+RJ��p��ر��e�酔�N�l�]A�%a�#�J�۱T���k�˱�����Ĭo��I�΅1�H��"Ͳ�騱��O������Y�B�@�N\vB8�*��K����d�8)wD�9�$�p���j������
��1��#l�GV�� ��7p]��z=K	�G�1AQ$���#���F��������냎:���#3�Z��[��[� �#��߱�Z��[���\�ֺ�w��lGG-4Ɯ2�`Y�֣�����w�ӸU�U��c-�����z�ڰ��4��"��u�#��6)��t�*R�ۺ!%�#z��4��O�"�����#�������1�:fO�zU�H�<�^u�7����:���H��>>2��#����#7�����2��#��l���pDR�*8��%cD�����;��#�nm�8劉:7��:ˉ߱����#7劉:���nA���;=���a:�������H�U���#l���-��@-��l����lxu�G���!�ޣu�#�����j]v�#�lJ��Z��;Y߃#���[�lF��^��
��W��c{�����Q92��#��1����������C&���2���E'8I5bܨ�{	2�3ӑ�2c1�����l����#=?ܱ�$�;=$��$��������h]t�#�nH�8�����4��<�߃#`g��{u�#����X/��|�#��$��i�9 $�~$�YD���$��	$����|$�y	$�"��l�R�ڴ��rX��dZt�O��7�!�M�AԅTM�a�V�{ng�����4f�\a@�U醨�������Y��{�׮n��6(�ɜ��.�X�+�}���>xI���"�#�룈tH������#��ȏt���b��X�����:��#�TH�:G��2/����#�<HˮL��T�D�2�\E�KY����`�#ဪ��KY���ڱ�#��9Y����=m߱����[����ϱ냝��+ڀz��6°�����"�#�룆tV������#��ƍt�Md �i�gZ4UF��Ƹ�ٱ냤{�mye�"F�Ÿ�E7��ۉ(���}�)-ܪk��W�D�26B��rI��Ms}�#(+?��k�s�_� �ϯj�'JlR����k�m�I��[�k�$P�%�f�	r�ߥ^% �ϯ�	@�]�=�k�$��(E�������^A������d�$�k�-��yyw��P����ϯ�.'�x�$��ܲ�5�;R�u�N3QƏ�P��7R%�zJ��jD�%��ϯ���-���T85���cw���F�o���o끿y�o1*B�E��E�<�o�1B��!��}4��إ,	�k��o�7g�o2��Κ�e���e�+�o����h�@��F�9�4?@k��8g�o2��͚�e���e�&�o���&!��o��k�C_d�-	��k��1g�o2��Ț�e���e�)�o���G��`~ISU�A���&�n��R�s���=��U��V��"�T%M_B`4�*X���t5�Yi5�Yi5�Yi5�Yi5�Yi5�Yi5�Yi5�Yi5�Yi5�Yi5�Yi5�Yi5�Yi5�Yi5�Yi5�Yi5�Yi5�Yi5�Yi5�Yi5�Yi5�Yi5�Yi5�Yi5�Yi5�Yi5�Yi5�Yi5�Yi5�Yi5�Yi5�Yi5�Yi5�Yi5�Yi5�Yi5�Yi5�Yi5�Yi5�Yi5�Yi5�Yi5�Yi5�Yi5�Yi5�Yi5�Yi5�Yi5�Yi5�Yi5�Yi5�Yi5�Yi5�Yi5�Yi5�Yi5�Yi5�Yi5�Yi5�Yi5�Yi5�Yi5�Yi5�Yi5�Yi5�Yi5�Yi5�Yi5�Yi5�Yi5�Yi5�Yi5�Yi5�Yi5�Yi5�Yi5�Yi5�Yi5�Yi5�Yi5�Yi5�Yi5�Yi5�Yi5�Yi5�Yi5�Yi5�Yi5�Yi5�Yi5�Yi5�Yi5�Yi5�Yi5�Yi5�Yi5�Yi5�Yi5�Yi5�Yi5�Yi5�Yi5�Yi5�Yi5�Yi5�Yi5�Yi5�Yi5�Yi5�Yi5�Yi5�Yi5�Yi5�Yi5�Yi5�Yi5�Yi5�Yi5�Yi5�Yi5�Yi5�Yi5�Yi5�Yi5�Yi5�Yi5�Yi5�Yi5�Yi5�Yi5�Yi5�Yi5�Yi5�Yi5�Yi5�Yi5�Yi5�Yi5�Yi5�Yi5�Yi5�Yi5�Yi5�Yi5�Yi5�Yi5�Yi5�Yi5�Yi5�Yi5�Yi5�Yi5�Yi5�Yi5�Yi5�Yi5�Yi5�Yi5�Yi5�Yi5�Yi5�Yi5�Yi5�Yi5�Yi5�Yi5�Yi5�Yi5�Yi5�Yi5�Yi5�Yi5�Yi5��O5�Yi�Ho@Ϡ\���7=�Р\��[`B<=�Р\Q��YiBYi5��Р\i5�Y;v<�{�+����o����B�;pp����pp�h�Y���Xi�Ŕ�Ѳ��*=�Р\�(56v<��`,���_]�;�Yi��]i5`Yh�Ld�8p��daBp�2ޅР\����}1�\i5�Y���J�8�ii5e�Ȃ��ܾ�'<J8��g�Gx1Jc�v��Sx~ij5�YTk�y<�Yid����2��c�Yi5p�R�eBp���ܾ�-=[��56���z�Y�c�Yi5p�R�eBp���ܾP�aaBp��&��d��ȋ05Fl<�k$�,�<br�����pp4�q4�m��\T~���=��<�\T�h��c�Yi5p�R}eBp���ܾ�h6�Y|����56=�]ɠ\�ze�i5�YC�ߗ�ܾ��L�pp�]R�ꔞM�pp�<��վ���uh��Y�;�ׅР\hEm�;FYi�Ŕ�eaBpp����2��c�Yi5p�R�hBp�LaQ��Yi����Р\�2Ie���j5���z�Y>��جpk,<d�Yi5p�R�hBp�La��,?d�Yi5����2�>o7��ܾ6$�z�2s����ډQ��Yid���o�6gp�0��2e~ei�2��w�,?�j�-t�Yi5��Eɠ\j5�Y����?��Р\�ν`��PG���?=4u��lUc[��x��Yi5F�R@:�h5��cd�ݤ<�Y�r�d�_�Yi��xx�/Yi5\�c��d��Yi�މϴ�d�>:�h5��KeE��>:�h5���Fxa�����ESn��&�IQ�-^oG��ܾ��F|a�H��cI9ς��Oe[�c�{�l��XaBp�@e�:d6I��]�8v��HaBp.�IA�u�)�pp�2�Eɠ\"0�1�(�i���gi5ƀpx|�j5�Y��$56?ttTIt$NLd�ȱ��s�k<a��ιد߇|��h5���?t��FxY��	��W�7ݜ/5�Yi5?��{�� <�Y�v�dq���K@F��fZ���Yi5�௻[T�[�&�5w����=\��n5��9�]�v�4���56v+h�56���?����56�i?��.h�56a@�f�3���Z�"��d�d����SG`;Ihϳ��΢[�w�[�w�{Z�cǈ���/B�f���.�e�i5�YC�߷�ܾ�-=�Р\�|]i�2��w��O5�Yi�Ho\��\���Yi5Ɯ-p�Yi5��΂���HaBp6�Yi�H���LY�r�d��Yi�E�R@:�i5��r�d�g�Yi�E|Y�H�x���M5�Yl��l7��c�ݶ;�Y�r�d��Yi�H���ݢ<�Y���c�ݝ<�Yς��KmE���~�&1J'�-�%���3���HaBp�2s����rH���[��މϴ�ڨ��<o7��ܾ6�������Zx��Zi5?�}1�\9�G��ܾR%,nd��Yi�V�)���56�UԶ�b5�Y��(56G�Р\}���/v��HaBp��IA�faRB�Yix|�k5�YT8�a6�Yi���ܾ��TaBp=L����`<Ie���56�Yi5�^�s�ǺD�i�d�����;�Y�5��P2�an�Yi��^Tw�IaBp��HD]�Yi�Lmmw:�m<H��ܾ!����/@�+`M��_M:�m<H��ܾ!����/@�S|?j]E	;�ר:Yi5�`����@2i��Zl|@q�~eT˱o�Yi$����g����/@���{l�T����c�Yi5p�R1\Bp���ܾH���Yx�Yi5?\hⱔ�v��4�Y�0G�|d��-p�tpLah(�5j5�d��Yi�|�"7���;�Yh����7�p�Fei�ǀw�Ɣhp^i5ƈ�c����w�Fio������?������?�R�����?�4q�7�ƹ@>�.}�feQ:�n��w�����?�4m��^l��/�8Gx<IZ*#���4��gpƔ�1�Yil�?oƔ�|ii�2��w��O5�Yi�HoX��\��$56���.�d��Yi����?�p���h5�m��lU@epLeh⽔ dXYi5X����Rp�Z�.p:l5Ja��Y�9�c�oƔh��Yi5��SD:x2Jd��[���/8?4ud��/8?4ud��/8?4u$e]�b����i������Z�oƔh��Yi5��S�h���.�e�-�u�P.KXad��T5e��@�.�:�d��Yi5��a��6��S@6e���ܾ�'<J��.�m��lUf:l5Ja��Y�9�ah��د߰��^�>Gx7Ij*�~]�α��~]�α�|�~]�α@�7G�n�Fil��T@5j6�hp��m5�Y\���Ȃ|��zu*<d�Yi5p�R�]Bp�/��ܾ��;�YQK�Yi��P�c�X48���� y4jdǀ}d��ĳ2ip�q�/y�Ŕ��p1��2�Q5�Yi�Ho��\ɸ��ܾ�-=\���/8?y�~e���/e�������h�8{���g��=�81޳B�\hEw��aBp�ƩB�Gz�ܾd�����ɶJC;���pp��);d�Yi5p�R]Bp�2��6�\��s�)g�n.�Yi�Ɣh�@��6�\C��);d�Yi5p�R�`Bp����oƔJΊ�yo2��ਹ<*�ܾ���2����6=�5#�\���6=��ޢ\�<�Yid���Yiw<�{�+�N���o����B�;pp�)��lf�8u�k��ii5��!
�\hE2�!
�\l��گt�Yix~=	<���g�8?Xtu��m5�Y�;=m��%<�ei5�,�w�F�i�y5�Y�0ӎ�Ӂ��k4����@�U�;�� r!�<�Yi�:��h2ς��QO{1i@���U� 2����=ud�N6]y�2�x��Yi5ud�;�Yi�Hoy�w��Yi5ȿ��ڪ@o�ʕI?����n�d��Yi��xi�g�<�Y��%����!F�,��V��*�GaQ:L�hp��^�ɸC�����
iT��@b��$D돾���3�}�3����E���$zH����#q5� ל�k�3����⢃��i��rGs>���B<��3�{o���?��Ч��09�[O��U&�CN�J��3��b'���Τ���J�Hh��(cK�es$N5����3p��ù��3��py�׻��s��n��B+�bD3�U$��3���3��<�]�3�e���ӽK��49@��o.S��)�3�̹A��}/_|Q��?���gv�x��I���t�7T�i���I�����Sw���0I��lI����>��qñ�`ID�nF������s�I���#�B�qēʊ�i�p,ɵ^�,��K���I��`�i>�=a��q%�r��p��j.���q���IQV�@=���+j���:I��i5.qؿH,�¹���,��'���u����.�JB�hy��H��򷧆Y���f7�?�5պ@�rd�	�?36��5�?��UO{�=1m�n$�#�q?+���5����䰄y��*̟16֥��91<7����G�5�?�hr��@,-��
1�@�z/0����`q�
��@u62����7�:#75�ӥH���`�}�����z�'��ࠥ�=~�?�͝Z�z%���g&n6�	���L�ύY,��?��48���,#u#
�}׿>����}Լ��������5�'������t`�K��	х���
��|�J�@��(���ץ�Mf�D:���G��j���_�����W�:�l�#�>6)�����M�`��1��ԑ%5�?�q�W���@���&J��%�NB6���W3�	kq;Ԩ�ʯ�l�ﺐMo�F؛]w'��
�"�~����j;�?vױ���3�A��]��I ��U����F�a�:�5�"�,�$�uq����z-G�<�(�<������L����
���6c�a�&�
���6�:�f:�6�����Z�u��|���g@�r�ף���H���Ԫ�D��5��#�_�qK	6��빺��[�+��pؖK&�@�ͩ	6:���4�7�=P������/��%�����0ִ,�f���SM�6��,�uҴ�&:b6v��J$=�)���ɔd�o�����4�X�@�91Tx�8�c��0�#{�v<�6��4ڨoG9((k6"�!����Г�,��
�wS���`� y ��81���D�̬��8wt|q���2���}x��6Ն2�CF49�5:w�������fTk�S����M�ƾ쨑͂��f�}�@�
h�H�Ծ����τ��\����?�j��(IN�����
��6j�?1��ǂ2t2�BY�h�����v[lc��8~���d���w��o��	����t	��(���?��96����"�^6ƾ� �?���n�a�����ל�^׹��5��������6�5@�w���G��嘛!Z����b�F6��m$�����Q!�Q��5�]0�91Tx�<��`�?0ՑFRk�%~�����l�j8ŗ� 0�nR���G��X��֨�U�3�p��G; 6ո��u}���O�6�~�o}:Q.8�f6"�!��� � �Ž��?��� �@���x?1���F�̴43�04��|��4��5�P�����o�h�(wp�O�I��vV��f0#t
���FSR��6%d���N�M�%�}��DؕOA>kIkk6�y��8�]���!�������(��N|~��ƅ����Q�a��+�ХY�����@��^�9�\���D����䝉���6�	�o}:Q.8�f6�#���ׄ����:)���әz/W�\6�m��
��MӨ7�C����hʒ��0��>������>�T�ox:����5��&�稛�ߺ.�Bk!�2����N�ԒJ�gS ؓP�	���Y���� �ل���$�6�-�F���|����8��W�A+���"7�F��6G=Eӳ����_���!�wS��SؾN�c@�s{�5`^��A@�ԑB��
K(�ܴ&I6"
=z�[��*ߨ����d��6�Ӟ�RQ".nf���
��\��^���p���4�,�`�]<����e���̨��P)�?�5��������	i]Ї��IaJ���"�
�dؾ���u�_0���
��b�̍@����66uX�ն�6����K����]���?�6� �,�nW⶙R�'��/a����
WOW�2�{���y�-������M���;�xל�55*�5d\�T��?�,nR�ȶ
^��0�ա�_MM<B�7���5�5��߷e����QGx��4�u���
�ߙ��w���9U6���%�?[��5�� G��ׯ�%^Ě T�h6�Sir,�f�i ���o9����5��#6՛��ӡ{�:p�0�"��K����Ϳ���6���zR���$1������D0�/��{�]�̝�כ�JƂ�"�~������ɤY?O��֟�[��l��7c�!������\�:�5���ԗ���t �x{���I��g;�����\���Y�	&l�ھ�Oh d6�ݹ[���� �Z��\����X�Ԥ2�ּ���
`{���L��5E���Q�L��~6���y�FSR��6%d����N�M�,���S���U��ԥ%�:��������ʼ�	ӈ�7���/X|�G�U�&������:N�("�|�(G�{澌�E?���剮Rޞ3�9���X3�@���@���m��x���c��9S+��������
36�T�ݔM!6����	��Sa��*SP�)���oG9((k6"�"	� �N��L���A h������i��&�Ԕ���P��ͻ��A@�	���_��#���
7��g*�k,���luh���|�
�w�ޑ%�S��V�\%iZ�����6pIxJ�l�Sir,Ԥ�F��
�Yy's��6ۯ�����?�ױ�?|��_k�G�?�5�r�o~=
@��}v�[�?��}=�5հ���������6Ղ���g��h0m���>cGuw7=x/�yVK�TC�I���@�`�?��.@�5�
�x����ax���,�}}�^�?���5հ���8����`�?�*�6N늝�%�5`(����5`(��_;�?�5XI�5�?�@�
@���?�x;,bT�%�}y�3�U�xC,@Ğ�)�5`(���,ɪ'��܊����t�����ax���+�}��Z�?��!@����?�iD̨[�h~Orڿ��Ҏ�Z�?���6@�3\�?�x�+�}��Y�?���6�@��@�/��@�`����Wx�5�?=��@�x�+��8����`����_x��6��Yԛ�O��6�6Ղ�ᇃ���5Պ��?�~�+�}�,=�8@�x�+�h��|�i��WF�QZK��A���WIfB�	З�+B���ܼ�ᇃ���5Պ[�?�~�+�3�+Fo#���?��
��1l$���?�+�1l$��l$�S�%��e#� n$�| �h#�yl$��q$�p$�m$�6�?�m�����v�U��W���c�Z�X��׈i�K�!�=1�Zi��^�9136��5�?��zC�@�5�?��!��^]q!�,���?���/��?��E�}�,���,���?���E1H��x�`��4���?�5�?��?�55�Y�_�� W�� �?�5�0Z���<-q{+���8o��,�H�5Ձ�6S����b�5�?�W�ELӴ�O<w�;4�~�0:136֥��91v�z��%�B���om�UXO��� ^!8�m�z�r?��)��٧�h4ZN�4�A�g�BxhΕ��x�?��*&IYfT\���ɖHz���КOVш[:���ʷT�\�{3)�э1�ҍ�T�\��3�6�53̎)�vE�'�����\�T�w|Y�HrO�Hơ�T�w��-QH��_)�-�Z��r*�;�x��-�Y��r��;�\�T狅
�Y���[�;�J����T���%�-�#�-�Z�T�b�C��;\v%�Zє;��%b�Y�n�JT�\�4���ҳ���8�\����ۚ\�����by;�)s�̂<�:y���P��X��Q��QJ,�B��A���T>/t�LM�0�,���7����ìvZɱL�AY)�f�G�RyX�����%���I�BĦ򫔢�N����(�â�)u2��w�����^h�|�T1�{�)Ёͯ[\�AGuM���tq��)К�d�}gJ �J ��)�;Ve?/���"�`zl����b(�����ͪ=M)���)��O����)0ͦ[�?*S�?*1�)�̦�[�X6#=�!M��_�o��*�����%���IB��򫔢�F����Ļ	���:<~<���M��e�����T�)�}`�Ɇ�N}JM���xq��)К�d�GJ �J ��)�GZe�`ă�5��t�7x%)_�*��M9�d+�k�ކH&��$u:Ẻ�!,�QW�ĒH��"���BM�s��$���r>I�i�U5i+!kf� ��Ԏo�����ޯ{��@��7����M_B�X)t�:6*� ���T-���8UL��F{��Gd1o�e�O�#�TL1|�]-���9g���F{��Gd1o�e�O��TL1\��/�Ȕ9ƨ�)��]^k�~�8�lAY���g�~��T/�w�/���g�@�A$ r$��m��´�9-B��4�4�#�?�;�r�G1�����,} �;��=��q�R������-���&f%<��.w.��	C����╂֮i�Txw�N���¡��='���E�<F�;��6gU�vE�eI�<L�ͱ�%¡� ��hYշ�;6M��$;J�UN�CE�k�U&+F���B�Rl9%��͡�k4���R���Ϳ����5�����O������%|CE���V�M�`�E�B:G,��F��ML,�#2�w�lwhW@4¨�����<A�L��O�� Z���!摁��*�,FJƃJ]�mf��mc�K�϶�P������?3Զ6��!٫��>��-�
}]%"�R���A���T�, �C�!��.�E�o����	�E���D�	|�Z��A,�0z؃����$t�Zn�Ts���(݃A���c��,�!�	�.�T���!�ߤ���sq��ӮW&TKo&���U�����8���z�3p�·
��.�]s��%�i�,"�_���ҋ:ă���D���f��'l�K���l�A{a�H�6���`9	�ҋ�׻��D���R�%��s:	�F�?H�D�Չ��_����D�ֱ�E�mU��o�^9	^�ѐMofyx�8	���(�Fo��y:	z�No�\��F��!�o?x�8�����F�9!x�q[����K݃*��{$�z��`oj˾L����
c�񙁎�ETԜBY��9��4�h��������;�����q�`v�~�'K�܎�ew�s��#TA�9ο�-%�hc���E��8QOSA��,����W�KD�{A���B�&�L/���\������V��w����\=�wx��h�T�b���E��8R`S���,����V���|*��>������^\�)��d�����ۉӿE��d�����?>���Փ�-���$Ƿhڕ	%�Fy������:�X����猟�>BCF\'A[����Q\��|��0�~�H���Dh�=_7�_0¾\4�b,>?��9�ۍG����i~ƶ�ѸK.$oF#$<?Ș!�pbJ��dJ#<?c!��N��@h�=ʇ��B���6h�=tޖpH�8����Y��Ȯc�ăA,>�
$<?lO�-�D'�$C�hY�yvE|�=?�9vpâ�	�����!a�Kh�=?.$aF#$<?Ȟ7��gJ��dJ$<?�'���=#�V���7q�IwnH5��=?hx����_ W�h x=?h>w?�j����˄2�{�đ<�Dh�=_�_e`4¾\4���+>�/���ެ��nHD�#�X������������H��.��J :O��Z"Lh~,,�3[�0J�j���AC~��Yv��~m���b�W�)�]Vc��"�|�8I�˨Lo�<�"Ad9�g�}q��>�S�y���ֈ�_Iy�AI��'c��Z��ڑ���
�=S�]ӽ\^��A�`X�߆�Z)sqǺ�@I��ЄYɩU�m~��P���~�����8�xS׉���rgb�uA��WY��3I�wٲ~{��J9mG�I��1�Xn5���ew���v���I��/I����3@���&E�:��qEV�W"��l�U���x���ݤ��W4�!��/C���bp�l�l�E�������^��p�E"����/	n� `��Tb����Rɳ�o�E�<��ԇaW�a_�E͖�<>� H���@��Xb����u�b�l�Ey�9���E�l$:�j�b*+�QaE���E�l)��8�A�J,A�_E�l���v��h�i���l�=�=Kp���ر������lvHv��s�.#3&i��<�o�^���#������Tb^�*�o�E��<<��aW�a��E�5=�Y�K���E�lc|)bwE*���Q8ʾa�U����ܴ4�0�\�d������ޮ|صψ��0}�>�ج���g�3��z�Ad�ɭn4�=A����n ���M�=ցUA��L}���{�M�ǘ2�E熖�a������|X;�_a���*����0<��|cy��Vr��傐��,f�/ށ�ӵ�`ab�ꮼ�����>i2�=z��0ޟL~�����������ݤ��ѕ�F�,��w���X���`�?�t��j����|���`a�����m�����Lm\�0<�|Y��
IR�I+�.`�}3�&��G�τǿ���W&V��k�����.�?�dL������,S�;aQ/�΂#���:��������_C��
<���Z����',hQ����a��8�&)S�I��/�L;�}���a�&V�h/b%i��s���&VU
2�&֡t�P�&Q
3Dr�I���qa��sV��/zF�0pMRL(֜�z�I���	���}Y_���x ��ɂ����0HR���6-�V?��?<QM��T��M�>�M�t�a������1�k͇^������"熥Q�O�J�ʭHR���OQ�6��\��ͅ5H��<����5�-5z ظ%K&���]��/9ؗR9e�����H\���9e�8l�b0"e�֎��/�-�I!��������c����0�90"8x��0Ȼ����,"��R�o;��y=EQ����H�-Z�ө �7g��9e��e�/S���9e�
�x��f�֓�/9,�>K���e�/�9:��)�G�5"�ҩ'V�xC�iU謯��w�%z$@e9��)�G�5��ǩ\����N!^S9e7D9e��R��i�)�+��f�g���o�,��oe���b��N9��lQe��eex���L�e��@��/98H랗5���@&���~�K264&��\�tz��R9e�eE��*p���sm[���s��]."�����
�.q�vfvyF_)�� \��H 09B���[�/s�I7}��2'=�&^1�a"�&;�e��W��6�P��4�BF�^Y��f�v(F{>~s�H�ӫ��9��߱	SA�����Q�CWuF�g���Gρѐ.�1g�p��~�8HtRgU]A�ݭ<N*��;ρ�J*�^%Aov%,�B���Ƚ$Y*�:9lH��6��%<�H�G���> P��7��2UsP����uq�l	���IZ�h�ٰ�A�9���I`��Sa'7�($��-��s�8Jz>7���.$[Ջ���\��@\�Q`Q�>��S+�K ��y�Οh>�n�c�[Q?+"R�R:����}M��?���
ݾj>G��>c��>9�hq�W�)��^{��l84WS�9r��z%�Q�S����t�0�V���GU�\�Q��i�.I�tN�'͛]��3��F�7J���^F��'�n[/ v��2=Vӓ��r�ǩ��	C�W�u��m%d�X݄�(�G����'�|�o�/!<�N�'͛]��3��.:��1�z�K�()7H�wYn�� H%���?�9U�E���J�P%@��:�sI�Y�$F�s>���mMn1����	ֻv9f����D�9�~�X�nfF~ �03��=�Dc�s42MH�9�&�Dҷx���g뀎��<ʟtk�{�G�[ʙ2�3H�I�]:tYL^��]�М6G#Gf��V��ip�p�t�mF�4bG�%	��>)�ۗk;U��`뀓ݝ��K��]H�=��5��3R�/r!����@/��4;t�;�ےxXHn��R��s�\��en��)E�:�Ȣ��L(�M��4�sL�z:�>g:4),��G���mMn1�H��4�s����c��3����Gj�y��V'0�H�NHm�2$gੳ,Hg��3�M�A�P�L{��O��3),��9����L(�M��4�s��G5noՃ�����G��^�fH��+�'�NHm�2$g�ԯ$�k{�Ȭx�HU;��L�z:�>g:4),��G����L(�M��4~s�@�yij947�-:�3�6��s��S��^�)��js><�8	���@b^��3u�_���l����b�,H`%�>OpJ�.�;r�69ly�µ�6f�����MEk\�s��)���x�g}���m G�m,T@�|�R��l��J�bS�K�[ 2�fA�rIB׏�&�N�'͛]�h%����y���chwplv>�K\P�]@�<vPל#��9_`�C��S�wPd[Q��>D*�j��rQn_�V��9�v�a���~��x�'jj?z�c�U� �",�wpN�'m�2$�4���֜�6��\XU�ުl�փmC��7yN�4H��; �U׼���%��z]灠���H�ߜ���MN��'��4}sL�z:�>g:4),�(:����L(�'��4~s�IFyi������(:ԙ|�����,���N�Q͛]��3��G�Z��4H�A�&�L�z:�>g:4),��G���mMn1����4�s�@�yij94���(:��^�fHO�/�'�N�S���4ѯ9�-�@�\�6HU;ρL�z:�>g:4),��G����L(�M��4���@�yij947�-:Зp��Rzs��M����΋jp��w�▂�'�_�ԓ�
(^pU�M�[� ��G��;�MN���H��)偤>�����i�J��2d|�M�SV�t�S*�A���=
��AH�>�9�g'3J.t@̋sD�5�>~^!U\����\?�vd���x��r��ڍ��v�JCk>�;�MN���H��4�s%��4�(ܶ�@�9�w��2q6��(w�W�C$�i�x�@�bv�Vøa��]H"�g�(��Eh�A _�4��Q>���mMn1���4�sL�z:�>g:4),�(:����L(�'��4�s����c��3����GjmS)B�y�
�Q�N�S���4����Z��3�M�A�P�L{��O��3),��9���mMn1����4�s�@�yij94���-:��^�fHs�
�'�N�S���4ѯ9����,��'U;M�L��2�(,),��G���mMn1����4�s�@�yij947�(:Зp��Rzs��M�Ҏ��>�i�(*u�?Y�������>nu����1�ղ=�U<�>�nʒy��Q���1H�K�9���Ʈ�t���޹UZ+ɏ*,S"�N�Q͛]��3��[�bz-�j@O�H>�Q�N�'͛d�$�\��8�1�����p�C�Ϯ=l�Z<��>�|"N5���'���;������$(ޕQ��@���_h�^�����M����9����\W���1����p�C�Ϯ=\�d�A��>�|�@5�t��0�J9�>T��#z�Jg8,3{״)A���_h�^�����M����9����\W���1����koC���^�M��L��;-A)�7�9$2ʍS-����C� � ���ўD/�n�J��^��D���"W��5˺-hF*!Q�
i���X��	�L6�͘�	���95�t��0�J��;��K�*R1��[+0�9�N5��T�,��4�;�ϤP��p"(��]	(An&�e+�GP�X���M���d3�\������2���@��K�∫Eψ30�9(A5J�t��0�J9�;TϤGO�p҇3�]	-An&�e&�G6�X���M���d3�^.AsY��9{����B��K�ck�VCN30�9�@5J��'�4�;���GO�p҇3�X	-A5J��'ŏ��;��s��=�9����3O��ʼ�/�G/ĺ���+/I���--��o�E2�cc(�Cu-y.W��:�;�D��Su�]�:Tv��m�������v�&��X|����m�E��e*�������%�ݣ� �9���'�B��~���Y�xP5��ˀ�ٚ�+R�w�iĠ���㚣Qd-cR�.A��=�g+?�-3��7�?r`�L��c��N��G��S��)�1�W�򆔄�=޵���N�Fӽ���@��	5�TSS��J��9�ɯJ���۷��JЮm�h�@*�)BM�B�@7�f�q�	$h8Ț�@h�8Hq:�(��s���Jp�ITcS�V������{��^��;U#v��E^Tc�WoNn�J�˹B�@7� �Z'�+B��t�@7A�J��W�e���3�@���Z��E�J��%n�Z���Z���@�$�醧)��j5l���g������Avj���CF9m]�^9C��_���Q&�,.H��@7Q�(�MHw��>Nn9߾��-�!c|��@7N5*�]W?eY��Z�8�o�?y?�|�����l4x����j�XR3A�ٍ�;N�^�jbz(	�&���j�as�l��j��vƆ�IF%��q�G���2���4,ۊ�d�OU�I��
08;�I�,Oz��cq��E)RJ��b��ޮJ�'�&Ǳ��8U̓��i&5G�s��⩢>�L;�I��Z8�(b���bI�%b�m���b�NƮ.|.fe�G�9�'Ʊ�l�§����$�2[���#��w�纙��Hv���|�'��'�&�ರ�i����Ʋ�H�W0m��0���74QW������W�H�	
�I���T1g\Gf�[���B�ͱ��к'� �)1xš-�=V�C]y�`Ү}�3w0�2�E�'zE{;�]o��@��8��(���GD��E����x0��a^�kw�4�?�;�/b�1iat���珦y��̷]�}��>��<4}/Jm0j����\Y̝R�*�e�z0��r\Z���l0�������j�p��'��NC��,f���ͪ��E�È�rm��S�^�̝+9��v��⺛�I����;4
�~?I�������i���2�"�6E������7̌,����[���j"h��A�'s�`d����V������I�����W�fe�2���sС:`������.0�L q(�CDqR�E O�=(����0�T��=�0�	��s�v�/{����j�2}!1���I��5G�lp���o���7���Ѧ0%��>h�hP$�}+�
X0�j0:+��Gnds�'�si��}�y���jĬT�?�&֌�4���S�E?�k�Q��ۧ�b>�~A��1�;�:����1�����Ƥ2���70��~�
����ծS���|��ǭ�L:���ɹ��E2t�X�Ρyn��+����',����`��'��i�7���ꈴmr�d0:�-S�f�};���_)
�Bb0�3��I���Ч��ǝO=��L��呑���/�M1ڌ5���gc-`�����C}�I���g=��۠�ǔ�K��Y��1*1UD*�	H�3O�G��� П�]�C���3_M�)]g�~��3:Ə��mI�ۙ>Y���C@���ԣ��F{�ƲGzq��Ujq���b0�1Kp �	�w4��}�ɡK� �
E+4i�lp�I���
R��Gm{���Gn[�'��Z{�͉���_=��/�JzH��0t��B��� ��I�n�\�Tƙ��o	�zN3�����L1QW�ؐs�ƽ�9O[E�ַ����1��~JP�Y-�1g����Gm{�B�0,�'���!c��尉d�?v,V~��e�'o���뤛#\���E�������z�CJ���DIh���0mF���gnPz߂Gt�E`�#g��E�*�@��H�t0��$�R0�3ur���Q�bp2ͬ&�a�C!��ᆲ�_�
>T7�AXoC ̒�H段����!�74k�՛V��`"�3nƲM�	����Jϋͽ�{	�%#�r���C4�?H�J��n�	�J�s�f�����Ǚ�&�}R�Z�T�z0Њ(6��_ϫ�'��΁�T�T�@젬�iU4a��gs~���X���r{���O�0�K�>�	˧��[Ym-����hIr�� �Y�E�C���FWIͩ�QƄ�h#1>G���H�K���VI�'����0b�n	%����;4�`3��X>��J�H�+n`�2��ˣA#�� ܑEa��d�6��YI��L\�Jei�'SL5[�o0���g���lj^�~�É��l5 �k�fg�>;�Ԝ��(4���`4X��遬L\�C��Ӥ�����a����&H��@��GH�!��̀�##ķ	�&}>� ie��=à�IE�Ӣ��B :ArJ���3Fq�q��Wx�/	>kԒ���(o���� =o��7�}-7k�0\���OeS�'~[G3p��E��dO�YI��L\�J.W�'�]$c��>F�u�͘_�i#�"�=�B�'_c����0���zGɃt�ǒ�Pi	���>>��`33����kI�E��b�O�����j����s+��F<�0DOӸ	F�I�众*���1�L�iV|<�fiI�s�0��`3ӹ��'(`�e}˸��X;��>7�F2 �Ս{!�L�Dܘ̪q!���� ����:���������B㵉�d0���'*��������'���C�I�'iS%^)�����.gYd�g�'g���D���P�q�̰KH>���V�ND�����%OI�E�I�*����G�H>�,
�'��$D�eF�I��I�v��y2��r�5YR�g(��I�E�T�g(r�E)v�I���K���=1�:��J��Z�˃���&����O�ߕ�����R���F1����91�}��a���s֖�����.ܥ~c|�k�Ov�H��f�}�����.�s3�
��?�g���bq��#'('�I���˅b'�I��X���v��>ݮ~���d�:��s��,X('�I�%�X�˅b9;�I�Ҡ�1��ͨ*�4����4R�I�Q4��B�ș���I������3�e�X$���6r4�bt�'�R/�I����ZIW��b����}�'�iPC�%���%®''ƴ�Ã���I�'�87�:D��=�Ik�Ȥ�t���i&5G�s�I��᩻�c���r��qCK�Ïe��T#�e}��\/����z��9�f́� ̐���o����M��W��Z���\�t�(�T���z���� ́� �)���>���æ�@�x:����¶i�b����^8��h-��?"AHs5X!�\��(�O���z��5�X́� �_���r�8���r<�I!HA�Q���?C�&����P��a���(��������osm���r��_"k�y�"�����7vMP3�Țx�X�	�Me%�$^��G� �eY,[��`;��d�L���?e���(6f�?Q���Hg|�p�>�5��i��~jρ�"���!���M��5��"x=u�3G��~�_�g=u0k�6R>�� ջ�%�x&Ƒk�(I�8<������^���mI����S��~�"�N{�Ar]��n.[��ջU)��h��*ջ�7���l L��|���d��r$��2�Cu{.�(�.윬l��l��E�?wA~j����(��6�6?��l����e�}�o1m��m��u����>�)���R�{$�nXS�FOIR�pK~ii�׵%�}��}Sxa���Q�M�/U,�(RK�!T:�����ëeC�Q��)!��R�Ț�XS�FO}R�D��~-���4�P�����jF�O�	���;U:k$,�Q�c���e�v�e��Q��5�	�TǛt����/UK�\S��z'�L�5U�� (dh�1��_�K�+$tY*��T���<F����V���m&�	�ۊX]	�N`#��COt��KE�Hhv���t}{[�$<7�0].��L]�^�G+�K��-O���=���Sc�&6��հ��&��&����_��yK	�zK	8����T^@��J?�{��$@؉�X�N&���&��&����_��yK	�zK	5����T^,_'�/��8,J����6��O
gY����5�6X���6��,7�(J�Q'��
���)�1���O&S*�.���x4��x,=M&s���Z  ϛ��{,�%ix2P�;y�s�jaã=���r"�x06�P�-���;�0��bi����6 ��SތFא�dp�E
"�� y�bc#j�݌�ˈ*Pᄸe�cH�a��B@3�����	�����?�Ŏ���{�f辣A6ZV`��XANFV`��_��J�$�Pj: )�$���]��������?;�f���'�Q�l�m~���*�Q�<�fc���kGN�b���s�$�>���-��_���#��Fz)�4m�������c�������ɠ�`U��aV{?�SF>�c��� ,K֨�"�dZ���țd �Z�8�!=���ؘ��s�K(EԂ7�L���'�V0|9~+]�("&m��7�����K^�(�,my���sǪO(O��{�V^� (�@61S��^�(�4$_�\%(�~������I�f�(��4�����J�|(���SSdvT~�V0|�~+]�("/m�п]����K^�(�&mZ� "���b�SO(���(�^�m��g�EQ�nY(�^J�e'%,R��(�^j��%h}�i�d��M?�N	�se
�`H��뾫nK�k*d���,���Y ���f�7�����JK��Xy�-y�X���xF��V����A��(����^��[��E�h�r=ly��I='
�ؽ?�s
��g��T��a����$�D��������=��=���q�++��$=�
��o�;��$=�Ct9m�E�U��d�4�xB&�������?:��clk��l�A1�)�����������e)2�6����Fa��5NG:�F���j�~��0-�숐2-�R�1�P��1�1DF��TFfJ1�"�|S��SmNU@7�P�,Gӽ��H-i�g��q�A٥Ol��>�u��o.ṯ�L����v�-\�Q08K1~N*��;�O^�	�AUl���08y��1D�1�P'.8c�1OnJ�l�]PU�z7<%�	�AUl�ap58y��1D�1��U�.,O�1On&�l��Q�z7��<�	�AUl��S'8yq1D�1:��&.�Q�1On�{m�U�T�z7�<�	}8DUl�5}08y=1D�1^��&.Q�1On.�m�qQ�z7�# �	�3DU@Y%��1D'�Vy���IO�m���58�P�'z '��mJ�Q�1�O~�Ϳ��O��W����T�w�t��UvO5�$N�R@�C�t�\�F��dAn��m�\�QfNE����68!Ory7���Λ1v��&`>�1V��&`7�����DU�Mv5Y�~4��Z-/��A���I凸��8�@�fQ8�χ�!(�m(������$2c���z��ipY��3um�?9���@������<�O�ʎ1DU�v�Pc
�7 �mn���T����pNU�1}���:�$�Mf���/�.U���1DU�;Q�@�@qc�(���I� 'v.^QDˉ:�NU�@�E����A�l�����]9w���ɼ6������x�~�TW��x�����8~S���T��7Ec�Iqjޠ���ymQA8�b�׫�r�]�Q��,\�Df����2�3_AV��x�feԇQ3�Qw&��dm�QF=We<^�w�#Qw�=UC�}���[��=	������Jc�y� �HW�4':��w��zQ8�,���S��fǣQ{`�\W��1❣3�k#*Ė�ߝW����S�`�f��Q�2��?=�=�arp6qQ>��	g�#�D��=�Ao ��*� QaM�;\�b���q�<v���<8����Q�[÷�yb�!>����K�w���Q��U�7�$q?�1�RD�:tM��"�=�Q.O����2$�v1oQ�f�QY�R��uQGf�
m�d�BU�1|��w���j����AU�w��T]u"�1�D1���>]B����Q�[Q��2����;핆�}�=U�D�b�T��o�����1��W�����+jvQYA���WVZF���1�)�j��6q~���Q6m�]���T�J�]��,���8w�M�T����&O�3~�"�$�/*Z�B�<��T;�(�16R�=s��8���K]9C;*�T���;nP����1��r���r��)OU6�"���z:_��2�[0yg�G="7�^7f�m��4��r�1"��=�ı�PD�[���)OS�f�K89���e©O�hԅ��G|1QKa�x�3k�����1�Bw=��h�Ł� qQ0	��g���4���=�*�ֽ�@�V.OU]^��ݮ��+����2�I|��kB=DU��"m\����(���*�4��7gv�C
�Q�׳��jMR����1���6��s8hR�É%�|B)fB(78�eO��4bEw�ѫyQ�a�]�+�Q}�����)�j��6q~��<U���Wt��Q�T��k1@��"����Tg�gR���Q�o��\x��1��̛]�y�Q��Q�?nk��VN4q(#��VB!�@(}�vQ�X��׽�4�>�-Z=�R��cm6��T��R�y���x)�1���/����VR;�bR�{��u�5ȳ���3�,D�8+�NWrfu�sEPU�\��P=��&w����ܫ�Q�dQ����������X�#O����T¼���XM8�Qk<�����1�)O��&OĔ��-�8VEgf�lq��^���wIc$����=������<!��H�"ۧ%���QO0�m��~���1������>=��8(OE��%,ImE8�&8�&�ad�ky���T�#�Q�ol�h��o1e�A���2�1���Q�}'e:O��Ui�1�(0i�#B��=U{����T�a=.Z=����kߗbR�2��?>p\hq�)��x� }������AI���Qф-���-�t8�5�2��9��}`N�mL�T���84�06Ҩu8=Hw��b�?���vQ���z�Vd38^��2�O?������[m��Qg24*�8�w��G���yQ~����Yc���s���QQF�pJ1��8��h
���wQ�=�w�0@NG=�j�3�QD�V�A>�2oQ��:��}�T�|���=블H�N����mQ��i���D��<-3�Td��)���,`Q�dQ����~�9�2�_�[�v���WVF���36��l8p�˸H��o�H�PW62g���;�s��8��-�y�a���P埍����~�Q�1���{��=j����|~*��\8�q�68`�������BU�����*ꈇ)��@�S����v1qQTD��d1DU��ћ+#�/-���Y�Q&�Q����T&=ȉ4!ۃ@�Q9�1�x�Aj5�c@��N��RV�L����N*e�M�R��<DU��L_+QI�QO3<ϝ1DUH��t���
Z�N������%K��s�:�fe�1&-�:<�fG3MfN��y���ͷ�n��O�����l(_�E��sP�x����~��}w�0���J=h�h���S�i)O�μa
�6DUƭ1�Ξ����w.��s/tQ�1Ȍ���f��M�q쮲1K�LzJ��	��AU#L������AU�Nz�r pV)K-�LU�1D
�2DU����4�/%�/t�a9��e���W��^��1D��:��'[L�j� ŗ�� 8̎=DU�
�2�OdqރyA��͕gJ#(Җ|x�y��DRJ��\K���k�Y.��	�B�� XV�O��ж�wt����i�Wx]��j�g[��$KŚ��L�Wp�(�a��K�,��4֓19n�`�����O}5f{F!)Dy�������յ����P�I�E!)�������L�oq�����f��a��0�1Ն�T=	!R=��Ev1���|Aa��FʯL�ll=��h1|b6�q~�Qs���12ϐ+����[��y����*o���cp�`�5�+
���������Gu�X�)���zKEN��L�7g=��m1�b�Qs~�Qs�.� ;n�,C9�7����BQ0���"+o���~g���5�W�c��G:瓛�؃zc�|j&o�z�����>w�� ��ޒO�L��������� �K�����	:`�Ƭ5�u"��'�Z|l}�DY�/ �?#��N��}>
�OaW�hpa�<ؐ\��������-�w���*�����"��4���?e_қ�����ASփ��8�e�7.6�g�Lw�֔�� �>n��:v?��"�iQ"փ��D�K�%�6�U��g�I�< ���g�I�Ӄ�MJC�V�.�/'�=K	�&�Q�[v��B2z� ��]��� �`چ��Q�7+��}�֛�
��ܛ�Cjt�̰�V�ʏY���L�ƎE([�݂����cs�gdv
��[���ٍzOʽ��"��`���`֣	k��B�L.���岐r������,N��h����,b��F�* mv��\g��i۞68~���z�6��~�Q^�]�
�6�s�����_�.Q8�)u�����\��ޏ���я��A� z�U��|0��`��st,�@V�������]��x�[`�*��	��<������&<O2k����h�@���*�&~�g��?�DS�1��5��!J_������nѭ�c0geb�J�w��T@iP��_�m�fDֻ�P	�Is�#r?�G����ri��Y+�[_Z÷+&��[w�멦���̛U��'?V|�
5��U�wU���VZU���+���+��2��i2��:m���y���{������|��7����� ���5K�Fl@��v*q�ϐ'��üQ�������&"�!��W�;5�(2�!��Y�A�c%2��N� z�&�5r����������z��S�yf�����LT��{rĚ
���oG��Sβ�	��K�����rT0�ޫ�.���u,q���ꡄs��)�
���E�gB-7��Ms�mC3@h^����
5z� ��,�Qr�ª�E'��⤿�����}!�D��9@�A�vA��~z�;�}L������F���j��M���P��x��2ܠ!��!�U�'a�:���Q�l��Υn�e���nZ��U��zP~�M4��a$DR�~��/r�V����6�"��ڰ�+ٺ�����G����1��g���6n�(X�5ɦ
}K��{�4x҅�@w
g{�-K��گ��c N{3V[�4<dm��_������������\-.�+�ѯg1(���*�g7�I������s2�%�1�	v����M0�הɓ����9��4�J����L�Tcςs���)����En4��!���q'��Yo�����#�7T���2�u����
���?U��!�(�c4�n)�*�)�x!�|�O�yA����`��V�����%�m�z/��i'�������K"�.���Jc�{�aE��Wj�[����Q���ߝ�U��mn
��fę.r@����+�ü�B+���V�OL;��s'-���ړ�ǹ��{�hA�b������7��]Bݤ"ʈ!�5��������b�a7,P'���' �����J��(�� غ����Y��|��z��'��ؙ�EC
@苐x!�Ç��`B�&��}�D�︗�H0O�V��9'd"x�77 ��Ջ���vE8���<-i���C&���8�* #DX��������{V�+�67�yF��ʭ��k���^)�!Ω;���)��������m����H���������Z�����Z�i(e^7#W��3�y���kp�?���f@��𕮠3H*1���^��&��<���o�/���;���!R����	����\�d��կA���$%�����
ټ���'�l��4�!�+�L�0,�ݓ��wzv��|���{!�ti�	�%�	ԦX��\��r6���D��0f�-�5��Lį�������@e/����z7�I����R�h�b
�Z:�[y>�#������ǐ��T�I��b�p���HȦu���{b���N��FZ���;7���^!��_�0ec��*��K="$�oE��Y5�4Lm�O8~����~;e�݀>�`�a����-_��	�Kٓ�:!l7�9���M��v^�07㠟�Z��;�8�������%�u��,����d"�W3*e=��z������)Pb0����V2�肋�
0��1��uEv�Yx2�
�d�n�)H�!.7!�YK�w�V����:�_x����j8��y�Tm!ۛw��3�:�����R��
�+7��JP֠l@��Y�X� �W���yA��}�T���(YS+�#�J�xgL�f��]cx!��nw���t�vk`B7��/G�'���|���\�t��a%x�Q�
��B#p�R��J��!ۦ�\��6��v���iB�v�{�:�k>х/�|��4o�~w�E"���F����ޗ�u�wy:��n�}�b�+�[���y!:�l���k⾝��
&ITɦ��4**�������}���m�4����QJ���*�����qHڐ�:�9�����Q�)�#ܭIό�cE�
�?�)9�{
<�&���6����� �j��1���[E
E\2*�o$���^��.=�����/7����OϦ�Uxi��0{1��̡Z�'�S:��g+�
��P=��R&�¸����C.��dQ 
��5K 9���+u�]�4*���:�y=ɰ�����&)��'{V��/��U�K�<-: i���
:�l���N�6��	�P�b���x!��
���<X;��������AȮ"9�sD�a����!}���Nֻ����Z6�Mk��O�ʰ�r�}>�;��#w�Ƴ=#��Qƫ#��i�bxm�'�S����i(	
��%}���e�n�S�K�H�ap����%�c�f�	��%��Ĉeo/|�
�� ��?�
��'�b�0�Auj��T:y7~�9�imy7~�����r뚟4�;�*�y6(�f*�_�����!�(,�%9�k{�ӻ�'S�'����%�HZ6O�ƫ����ڈe��@�hƳ���c�!-���&�y;���w�)�
0�~Y��LV��C�lZ~��9P��� {VM\_5��=L{V�1��� ��s�l�(�ꒂV�<e���vU�{V�RvV`���.�Ru��|�{VKwV`��.r�x���ք��.����f��A�{V��{��z��%�U��S��#�{V����T��p�Ew[�f�l�2mL�|�#�v�[�V%l(�4�v�!tb����Ct�*tQZx�zJtK't/���	t��	t��KXM�:�}�f\e�@�z���*~������4is>U�U&|���X�z^#����$ޭYK;��K\6�U�E��c=Q�.<�S� }�ˋ]�b1{q�VoN��V��\o�G���gھwə���Q"��ZI]�*Pm~uЪ�}ʱ��={)�@���',��C�����s�V�,�!���noR{�[�b�g.k�z�dGwy)��_]�Vo�y����{ڿt�-bg% �z�OSuy�'�{V���S��,�h_%$縊�v���V罸y�V+P�NW0/�<�t��Z<���K�W��\�)�t�T��e#�ya���Q�] ���q���1��9�Դ�۳��0�29��2��_|5t�S�x�/�a_��b�=�����v-r�����_������?�~f�L@�4Ԏ��	�Qu?@or^��x�:q`�n��F�C׷��<Es�۫�_�M��:H��Ō;�q��޲�a���Lx��{'���gc�]�6������(O}7^\,�A�������>h�>f�g�G3�\W���H�F{׏����9Chz���uC����άuW��S�1^�I���tά���0X�/�z��e�S�+�ޥ�G&��K��Im�0��$Q/�gZ����^�h����Xd�g��t �\����kJ\���h��Àb���s�8M��Ӽ��o���&�����ՙ?}qp�K�z������c�q>h�(�n2;X h�u��G�d��Ɔ�^^��b}�g��v�\q�3���a�=h��Xh�F��;WȞ��z֙{d��J\�\u�B��Fh�����\Vm{�
��4��{�g+*y`���BG��[M�����?M5��,���h���h���K�_��d��'uȇ��4 �g����:ᗍ�p{�0�b�.�*zp_EZ�g[WC������z�J�{rs�\n��Ӎ+�R���fj��TL��M}^i/J����.����Z���<\O�q$H�\�+�$"����D�d�ܘ'�_�J�{�dfUvaz���Ϛ��}�(�_�H}^i�Oh<���.���/�Շ���t]\܇
b�J�\�To@�g����R.�po����׊�=¡`�f)F`\U�O�њv�8g�+u�D�����21�N������K��e���L��h����bh�Ù��z�SJ\�+_���st!�1��8�
Xz���Zh]��}/h��������BKd��.۴��~hM�������h�:�GM��O��7�!��g�zd���A�>�~<�H�kh�zk:��:hE�#�8�X���"�J̭|�0���C���e���gQS�f��C�h+*�4Ŷ�h$,��Ao�jUz�B��ܚ�L����u�����v��:��!�&^|�V۠�ʫv�Z/�� 	W9����\��!�o�cPqg���*��jbۖ�~�q^i�Iyz���F���l8"ٟg;�:#BM��p�4f���/�bٽJ
�]]Hڏ�\T���=�?�
�h��Ԡ����_4�h1qZxp!͓�Ji���gueF{A�]]X�#�M}^i/J�r��.b��0�����r15qM�5H��s������2����@]\m#f����K�N�u�h�hA��MɊ
e�;!�M��<X|�M����g$�#��J"�.^\!Cy/�*��V���Fh8T���z��a�F/���2h�u��&!^h�[ h0�+Qc��q�]�I���?�ih��J�!��S �_��S8�Tz����k��,�^El��z}��o\H݇Z<��jP�$ް��q�zש�彁>�Z�����/� h��&ZCE׋�ik9�'N[&�ֺ�Dv�4s�x�s��4�m�h���D�9��g����{��u�����r֡�K�V��H�ث��_��t��pp0
b)��KD}�Y��1��K\�_�g�C,��
��Ҩy�L�0D��Ng��}ޕ��/�0r����oA>��¥)�7N7�jqx{G��?�:ۡ�K�B�&��<��j��k`�u��,��7�NQ�*v���7�����Z7�ا�J�o��]�����2qU���u>�T�ug�u�~g�}Gaq�3n�S�/�^N��2�b�b�cn�FV�;���/���!j"��y��ѿN�h��(b2Ջ���q����@��T�q�d���{��q�Y�u���$j!|�&�v�#����؏s�{��MMf�g���|�s�z��C	{�ݐN��"�e�]@9���[���!�����C�SJ����>��U�^�m4+@k[�k�8)��c�ƌ�ěR�d��2 LYo��c�S���^��놦�����XR��z��,���iR�*=�����f��ыt��d��w�=)į!ӎ-�$6�}�_y����y��ڤ�؜R�ܕO�stY��%j�� �f�O����͕�q���]�߻��p������_rքW���#0�o���}vyִu*[���������	K��q_��p_�,�_����%�_����Iq_�Hc���x_u6:Ox�Z�\�}n�.�
�zq֟o�9%à�V��3-j�׶��`��`��������m�����P!�_��6�q�_��_,����NջѪ��`���y1 +�vp�_SnI�E+Ǿ����=�"�>q��&�^�K��t���O�J_�ou�`1��+�_��R£Q�[YB8�a�_��}:GN_�[e�_���[
����=���/u_�ר�P����,�,j��J\��EX�_6��j��7�#�H����\�jX���u`C%q!�VU^/P{aGT���̲�ք����+��?<Ô�q݄_�c��gmz奾������xFE�\[�Z=|i�N<���໾���Y�h�Q	2|���z���swTt�ź
�~=��4�,x�龻�ź�X#�����c]��F��?�@Y,��ר�LK�r�Z�ף���ź*�J��$����+�ź��6<��1��%�\L�޾�V3�h>�%[�-�B	rT��p]吷�	�0[L<3�Ŝ,�!���G���ź�����źwP�1ֵ�B��F��X#���.�E�9��h��bj�3��RMV�����ř
E#���J�EL#�{J��"��U6�������'�dz����'�/'˾�e��R�ԷfwS�p��$ٝ�ZN��ǼY�j��2ؤ&m���jC0˝j��$���wZ `���x����K(�{�f�g1�ִ�(`N�n|S!su-��y��D����Uꃍ|8㢙�R�����B�*�O���?��W Ԙ�R����R!A�e�����R�R�҅�ݗ��S�����Ș�R���U
@�e�㟖�R�~�G��^��?�R�o=�0�*���|E�?5���L�
/�
��|�W���ݪK�K_��'���{
��D��ȉ����`6�;��ġ Zi2�#�l:~����77`6�;��d�mYi2�#�l:~���$'� �g
Zi2�#�l:~��gD_�a6�;��$>m�2�#�l:~���$ 2�5�;��Dm�2�#�l:~��gDD`6�;���)g
�2�#�l:~���$o5�;��I|
Zi2�#�l:~��gD�%6�;�逤�m��2�#�l:~���$���5�;���m�2�#�l:~��gD�>6�;��d�l��2�#�l:~���$Ƞ�5�;�逄�m�2�#�l:~��gDb`6�;��$��l�2�#�l:~���$ �o5�;��D��l��2�#�l:~��gD�H?6�;���ۅ
�2�#�l:~���$�w�5�;oX� GwUo[��vv���6�m���_�w�����v�[��vv���6nM�Ln^�w��� ��v�[��vv���6�m��_�w�����Vo[��vv���6nM�2{^�w����g��[��vv���6�m=h�_�w���`���[��vv���6nM�y^�w�������[��vv���6�m�5�_�w��� ڥVo[��vv���6nM�3{^�wb�@6FwUo[��vv���6�m�y�_�wb��]Ew��[��vv���6���� ��[��vv���6^ڵK�_�wb�����[��vv���6�A��_�wb���Fw�[��vv���6�g�b�`ƥ�[��vv���6�����_�wb����[��vv���6�i1� ��Vo[��vv���6[O#�_�w'��@�I��[��vv���6�Q*�_�w'���W��[��vv���6���Nf� ��[��vv���6�#-Z)����Fw��[��vv���6[t�t�_�w'����I�[��vv���6�#L�_�w'��`�FwUo[��vv���6[t-�_�w'�������[��vv���6�#���_�w'�� ��v�[��vv���6[tU��_�w4�@��Vo[��vv���6�#��_�w4����Vo[��vv���6[t-H�_�w4� GI��[��vv���6�#��_�w4��'��[��vv���6ƴTm4�����[��vv���6��N6y^�w4�`����[��vv���6ƴl��_�w4���;wUo[��vv���6��t�_�w4� F�v�[��vv���6ƴL��_�w9�@����[��vv���6��>��_�w9��^��[��vv���6ƴ��_�w9� 5��[��vv���6��6�y^�w9���:w�[��vv���6ƴt0�_�w9��L�vUo[��vv���6��^�_�w9�`����[��vv���6ƴ���_�w9�����[��vv���6���_�w9� s���[��vv���6ƴ���_�w6�@�D�[��vv���6��&ex^�w6������[��vv���6ƴ���_�w6� ��v�[��vv���6����y^�w6��Y���[��vv���6ƴ���_�w6������[��vv���6����y^�w6�`#��[��vv���6ƴlf�_�w6��Q��[��vv���6���nx^�w6� ���[��vv���6ƴ�S4_�w��@K�v�[��vv���6����^�w���͐�[��vv���6ƴ�^4_�w�� ��Vo[��vv���6��>��^�w���CI��[��vv���6ƴ�S4_�w�����Vo[��vv���6����y^�w��`P;w�[��vv���6������6N���mP��%��m8�r ��B�5�w�ܼ>���z3�5t��	��V�ȞP�Ԧe��m�"�~z���Y>�� �ҹ�#�&jq���Hwժ���2t$������?fP� ,{�Ӳj(B�@���Ӳ�m/�5��z�?���`U�v��F����~z��>�-V/�iM}e���4�p�����V���i�H�V��	���Qy`1�Z��r��mP�=�vչ�0�gPzY��8�iIl�5'�F	\�Y$v��ܘk��
G��]FM�U��z/��@@b�4���SkVf�s=��{��mD��(��S�a�����.;��@�x������na`>S����3��`opmfW>U��z%?Pʄ]��Kto������	�]2m�;��X���j��~��`˫`�V,C�n�(�Ϋ�;���?�]y�9�G�YlNG	J�`�;E�7W�G;��:�S�o=����l�0�j�(a��\�q"����6��Ξ�9�S��=pdU����a>_ݵF���,�wr�
z,@B]!mstϭ�y�oc1F��-ϚȦ��o^ڥ]W�{�\�c��(����r�G�gF��抦��'S��Z&�F�Q��#l�mE��V�����G�gF�/����'S���;�F����O��A����:�D��y	濾��u�`���86R�~�-���b�ƚ��@����pg�>������M����I�ÅD��Ф�d���,iu0c���((s�H��ċ_������e������{Ӳ��������7�L�c��,��.Q�k�V\-@�$_(����4��C�ȗP�k~Hu�g=�ɳ���g���υv�0��8�zj�h����� ^o��W�F�8x�?k���V����*^V��r0����xӸW�7%�4R�Z��N&vJ"���~d#�xyU�B~^p6�>�xq��ɚW�@�������I�̞B��0��;�f��p���^�y��������J^�/�O[И[�-w�_Y�d�~J�ñ����8��-����a־
��o?NyP�EW��,eQm����I�6���9�x���A;��$�&F�j{{\�H�u?^�/�W3�Ԙ[��-w�_Y�d�~J����Y~	8��-cRaVo�G�xǫJ�Q�8KK�e���:���A��^�sO\?�v��x�7˜ɼB�1�G�����+X?1��.���r���$�N}?e��!��<��ı����8˜�-H^Vo��J�ǫJ����k|9 ����℞i�[qJV�C�<�ñ����8��-#r_Y�ǫq?�Q�8KK�e�� �:eD�>�y���=�<�Q��k|)��C�:eD�>�y�t�=�<)����o��ј�$G�N}?e�q��O1�����<�A|{�ɲ T�����J�Z�9��W�z�lP��"�:eD�>�y���=�<�Q��k|)�J/��-w�_��J�ǫI��W�z�lP����℞MG�#�c�C=����Y~	8��-#r_Y˕��$N���>P(Mz����$G�.�j{��!��<�
̙�Y~D;��$�N}?e��&a�O^n��LElИ[�-�H^Vo�G��d�J����Y~	8��-����a־S]��J�!�FY"����%Ŗòn��nS��dZ?��X�z�l8 ����:eD�>�y���=�<��UNKK���} ˆb_l8��L��٣<1w�8k~{��:���>�y��:J�<1��z\�M*�f��ɖònJ�4V=�Z?L�ޑW��f�d@ Ŗ{��k��=Ѱ<H�q>u��^YL�ɖ�d�Z���y�d�<�Q��k|����h9���A��^�sO�<�v��C~�^Šzf@����[6�º<1��.���r���$�&F�j{{\%���$��ı���A;��$G�.�j{P��A$1�����<�Ar���$�&F�j{{\'a�\?���e�����:�F�!��v\�:J=1��U�8kc5Ŝ��ݔ�(�W��3\?NyP�Eh.-em���
��O���Y��JN����<��^����$\�ntz�G�!��<��ı���A;˜�$G�.�j{��&��-<1w���r���$\�ntz�G��H�=��Њ+������:����A��^�:J�<1��U�8kr��k#G�.�j{�!��0<�
̙�Y~D;��$�&F�j{{\�H�u?^�/�O[И[�-�H^Vo�G��d�J�ñ����8��-cRaVo�G����2<N��ɝ �Qm��$G�.�j{ƶ!��\?ʨS�*����Gh��:G������f�> ��୐�r����x~�:�N�����as(�tS\*�1k��X��fR��v��`�[��p%^Rk��z��f�i�M� =B�52��Z��o�;����֊�HtSR�S��2"��F?��?`��北N���g�ܚ;"G�L�����`@
P��X7��K\{�;"��?}�
���F���suM��)�;Ot������;��P>X7��،j�;O������'�2��ͤ�2k��IA������7�X��U���6Ƥ�2k��*1��2O��`+����'���S��	��-�Z���AT[C����m�ךL��PpE�i,�،jf<O8%y+�Mb�$�����p��B8{{ m#e<"G�L�3���`��P >X7��K\{�;"��&}�#��`G
P���~3�.��`��yc�0;�q���+����Dk׀�IA�52���7�X��U���v�'k�pc+1�i<Ot���Q�'���S��	��-�Z��V;T[C�=�ưךL��P�e�~3�.Ю�j��O�In�]���?���R���͒����;��e����C`�����~7�y%uJք���2@��7�XΡ;����ͤ�2k��X���2�˩IJ �������f�E����;к�7�X��M����&N����ۦ�;��e��֊���t��6Ƥ�2k��CA��2���7�X��U�����Dk׀�X0��AO��`+����$������Ķ����p#�2"��F?����`��P��X7��K\{�2"��L�����F������9�);Ot������;��P�e�~3�.Ю�j��O�In�]�$������Ķ�CYn#�2���?�К���0��v�'k�pcDA�52M鯼 y�uU����ͤ�2k��X �A����`��pp�8� �6q}�����J��g���T���8��dL �"q�JCٌ!=G#�C�D����$�u��.A��U�3�?�Mo;��E%�$��.�+�-A�y����� Mc������#0�3��Po� �:Y"qU�����е9�K��5��N��Moa��E%�$��.�+�FJ�iG������lzS2 Z��+�h�+A�O�|%��5:YpqU���^b�|�9�K��U�3���Mo;��E%�$��.Z��FJ� 2��'|��XU�!�����7G��$�J�ꋖ���l$Q�5�*�&�$��.�&�FJ�N����q=�Dς����:ۀ�.AKYV�]��lY6�g�El�Ԫ#��;�:P��\���-~����a&�$�N-��-A�x��j��)5�a$8��dL %�
q�GJCٌ!�aH�5�@ 	�-@-V�lXCFACٌ!�·�%D�a�El�+A�lX�An�h��{�O�I��y窅R}5��,�;�l�_����eR��r[v�ʐXE��o7G̪����b���	���<�X|��0��2z�2������j7
ݞ����d��26�{hR��� �j�������K/�D��;շ�r��2�%P�����d��2���� L���-���{��6J�<C�y�;)��_���>���_s���݊�U�*e�Sz��
Vݹ����%�ƣa/�5��h�[�C�$�f������e���0�D�{;us}��D�8P�����d��2���{ L��[O�v��{��6Z�k=y���~:�P����K�,��QҀ���t�x�
�n�Z4�Nǧ���|ƀ�d�qF{�2��>���S�u��i�{0�|�I�\}NOt��x��ѣ�At(��F̽��h�vFߧ���*��q��4F̋��r'�5��S������q����r�/�|�{����Ot���Bt(���r˽�|�I�\}NOtq��x�-E��p9! �q�Ǒ�Q����tD��
�n�Z4�Nǧ��-j}ƀQҀݍ�������B>�P��5�K�,��QҀ���t�x�
�"�Z��vF� �,j}0�Q��=������ �B>�P��5�R+0��s���ڷ%VNn�� �7x����	@��Q��=���Y�q�h��[M�jċ��ϑ��r'�5��S���1��T��4���~���c�A�nv�Ts��B>�P����G�,����qFߧ2�t���\�?ě߽K�,΀Q��=����
� �Z��vF� �,j}0�Q��=����q���>��� w��i�{ƀ|�{����wG���Z��vF� �ǀ|�|5�3Fne�1����.E��p�n�2r�Ǒ�QG�ݍ���
��Z4�Nǧ��-j}ƀQҀݍ��ѵ��3�B>�P��5�K�,0�Q����tD��q���'XI��{b�������qFߧ2�t����g�r���R+���s���H� �Nn���Bt(��F̑��h�vFߧ���1��T��4����g�QQRrxv�Ts��B>�P����G�,0���qFߧ2�t��~:�P����Kf���F�{۝6�.���B��W�J���\������Ϭ�4�[�Z�Q"�^*`�f3,\q춝�LB'����:@�Q�
�%��%�3w����%IT�34���Sy�B��F��<ґ��g0�	�#5[x�S��䧲&F+��3�go���3��[x�oPȎ˴�%�g����gZA;�3�p�!ʐPyvTv��ʈ3ґ+�go���3��!��SyvTv��ʈ3ґ��gZA;�3�p�Sx�oP��䧲&F+��3�go���3�p�!ʼQy�B��F��<f3������Ϭk�;o5�Z�Q"���@>�3,\q����LB'��� �3�Q"�T�@>k3�w��ɵ�#g�U�<�G�SyvTv���!3s������%E'��뽏7@�SyJP)���!3f3����&\�o�����ZB"�^*`��3,\qH���LB'��� �3�Q"�_*`�V��w`S˵�#g��L�?�G�Sy����b+s��<���%E'��뽏7@�Qy����F�-3f3�E����Ϭ�+���Z�S�
�%��*�P����go��Q}T�!�IPy�������h3�<����ϬO����Z�Q5Z�QSo�ȕ3X��&\�o���'�ZB"���@>�3,\q���ϕ�KSUg��3B"���@>�<,\q���LB'����7@�Qf��<�F�3\���go���3�h�	!ʄPy�B��F��<f3������Ϭ�X9�Z�Q"�T�@>k3,\qr`�LB'��� �3�Q"�uE��3�v���|��r��{�y\��J!��uE�-3Zwq`'p��]c�.�Bȕ�䧲&F+ ��3��h��r�L�~\�bP"���@>3,\q+���s(g߂n� �3B"�^*`�3,\q���LB'��뽣�3�Qqҡ(س>3�6ߞ�go��Q}��!��Sy�������	ӑ<�gZA;�3�p�Sx׼Q��䧲&F+��3�g���Q}��ץQ���`nC�33]��4��<鹷!5ʵ��Sȅ�y�$3 ��4��h��r�L����IP���S��6�{��g���Q}�[x�B��䧲&F+��3�go���3�h�	!ʐPyvTv��ʈ3ґ+�g0�	�#5	���S�n�1�3��r������KSUg��7@By����F�-3}�W`S�^D4�����S��v�Ѡ�UG�`���<����bMvB�u�%��%Q� ���gZA;�3�p��׼Q��;"+;�_��3��<鹷!5ʵ��Sȅ˴�%�g���h��r�L�~\�IP"���@>�3,\qr`�LB'��� �3�Q"��uE�-3�vq`���r��{�����J�Y3^[aE���F��q[m5����B�q���MM�z��go���3��[x׼QȎ˴�%�g4���ۦ)g{3�G߅3�$Z������=UȔ7 ��8%����e 2�/��%l{�"	��7�e��F'6�^<n��d'�S���׭�˧��n�ÕXj+�)�)��_�T��)�p���5 �����Vn6�~U�@X\��2Z�IUB5y��s���uy�T�\�A�}�Ļ�w�B5"=�V���W��+n��Nc�9��?Q��7J9l����P)����d'�S����p|ͣ77c��U,�W�f�0�l��4�ݶ�l1�J�L�?�8�Ɠ��p�Ed�����z1xL��u���J��-��+%S�	����b�J�Ġ�x����@0������%ye:��z1�J��u?x��F��-��+%S�	����b�J�$u���5�-0�78kA�kx�T`�J��:^�b��u<f��*k�G�H	��b�J��3^�b���=f�X��2P'���J84)��V����A䔷��������xL�v��?�G��F�+�K�?y9�ګV	�K^��1*�&AE�p�<��(�=���`%�ͬù�]�E,�?�x�o�o�����JlV�͖� ����n�0I�d�L<I ��8�Ʒͣs�z�������,�����'V|R���ʖl ����+�F�op.j���dHlV��a�����[��R�<�sx����|`%�ʬù�]�E,�?���o�o�����JlV�͖x ������F�R� X�O���	ʣ�~��Uk����؄��vF�FR�ľ͖B^�3%u+�F"�o�G<M���>�U�l�I�E��u�����;��i�K.����o��� _�2�"���y�@;f��?sQ�U���/0l��3��G��|)G?A�]h�`~��BfEY�%4 ���5|��@���=6��|�Bv5���Eǔ�G�*K7Y�2s^4�`~�U60�GY)�Fq��g0�|�)*2s��0#C �Ղ�3���G��?itQ��-�Z��l�����'����|)G?tt^h�`~��B�GY�C��ͧ|[�ttg83|��BK�_�Jǔ�G�*K�L�2sgS^�|��0T���tT�B�|����t^�ĐƉϢ�X��Eٻ�70�|8Y�}t^4�`~�U60f�X)z\Uu]�D�E2s��E~�.<����ó��˴﵂`�2sg83|��BK���8ż�70�|�'�}tQӋ�gȟ50�x���t���v2�|i��s^h�`~��B�1<���GE�Jd��r5sg83|��BK����8Јv�/t�'�|tQ)Z�gȟ�0�x����rig�f6���2s^h�`~�忭������TGj��.�x}�5`��S�	]�Rj�a;�ǝ�A�H��.�� w[�ȅ�ҩhm��@�H��gWs�
�EϽ�L7:��8dr�A�6�V�~u!�
q�Ee'�L7`x�Ύ/3� k�a����@	����E�� L7�ȅ�ҩhm��@�H���>�Q��{+v��E7��ɫ�P�@���H�~u!�
q�E�uG7.�Ua�.F:��甞�M�Li%X�#ÍTK7��+;h-�L�@v�ǝ�A�H�H�� �5��I���Ms����:�A�H�ZE�,"K7p�g��)�@��F�~�i��=zx�.7�݅�ҩhm��A�H�~QX�
�nE~��L7���944=�ͯݞ�Ml�;���@��T�5�{���h-�L�@;������E�� �5�xc���"f;Ns�;���@	���n.� x[ȉ�4�n���Gw������Ea" 6�ɫ�P�IX��H��2v�
�Ď�5��#���z���Ml�;��"�e��T�5�^���m�@&�����2v�
����5�YH~�m栬5��H�~u!�
q�E~��L7�����j�@8�֓�i��7?@jE�RL 6���H���A���~��k��=e'��5`��S�d�%Ӄ�a;��B;Duz-.�M1B=7�����h�W��8�MT')�	��ETT�5�YH~�m栬,��D���0���qE���F7�4']�k�5��}�~�i����c'�.7`p���hͿj�aH�BN�$1;mEdK0�5.�r`�* ��攞�M�Li%yI*7kTTK7��ă]���,��������Q9=���E7��T�ҩhQ��s�H���l.|J��F``��5�I�#鏮��z��w�MT')��&���T�5�����j�@&��w��2v�
����5�YH~�m栬,�����2v�
����5�4']�k�5�ў�~�i�������.7��ă]���5�Ѷ�~u!�
q�Ee'�L7`x�Ύ;�I"k�a�������E�� �5�xc���"f;Ns�;���@	���E� 6�iچ��>�:HR���@	���fE�� �Z��I���Ms�Q������E� �5�I�#鏮��G���@	����E�� x[�xc���"f;Ns�;��:�A�H�ZE�,"�5p㩪ҙ�O���Fw�~5���E�ZEzx��5�͔���"f;�A�;�~QX�
�nEe'�6`��S��he�a;���@	���6H�� L7�ȅ�ҩhm�Ms�H������E�,"�5pU�V��Da���FQ�~u!�
�nEzx�=7���H���A�Q�~QX�
�nEzx� 6��c��C(�Ms�;��:�A�H�ZE�,"K7p㩪ҙrXQ��Fv�~�i9�̕�4�9��Gީ�x� 1,�u0x���-��ԯM:u��{��Ջ��Dx-�Ի��ԯip�u���Ym,���u�x-YԻ��Ħ�����3߃	D>��d��w-��{;wr��R���X�uG�i&��tO0xC�(���믵�������t+7x��y�&͵�[iš�΋�������"�u0x-�+�;wr�������3߃	D>��d��w-�+�;wr�ip�s���Ym,���u�x-�+�;wr��ip������x� 1+u0x�l��+��D��r�Ӫ8��ѯ-�x�/p�F��0�M:���{����2��D�x-D�"�z�ip���B�]�#
(��u#x-�+�;wr�����r��3߃	D>��d��w-�Ի��ԯR���X�u����"�tO#xC�:�,�X�^��y�����t+�d��w-��{;wr��R��Y}�!�=��tOxC�:�,�X�^r�y����wF=Ju0x7��M���������|>��x��w�&͵�UH�� ϋ��|���%Ѡ됡x:�7�#���y���Ym,���u�ZZ�`���j�?"��^�Ƚ(���uJ��UE'���E�i'��S�}�|�&�E�� �6�
�B���Pk<��hd�ꮓ?��'��#�&Hm;U��%Ws#���)��עBW��9�6�
�B��Pk<򹗾���!:��v9�NV�[N�n�����VJ��rB�"P�����V�
:��"��})A��;uBE��J�H����0�O�����8)��|�.CVZ��0@��r��9�����S�}�|�&�E�� �U��j8���Pk&��n[����v��w��� &���]�L���<�ډ��Z�� �x�5�j�?P������!:m�u9Z�� �x�5�.APn|gи�T�}u����V�y�5{�"���^�Ƚ(���vJ�̤�V�y� &�J�]�3�� -o��KZEQHu�j�?7��[��l�u�Z�B(�x��ৰ?<��hd�ꮓ?��'��#�'�Z��t(��?�/&F82�ܮqTTZZ�`����j�?>�[��l�u�Z�� �x�5�.A��m|gи�
��}v�0@���5{�����^�Ƚ(���vJ�̤�V�y� &�J�]�L��8�/��T�)R�i����'F��]�L��b����T�̤i���*��]�L���"��������^Z��*'�]�L��S�ׅ��TZEQHu�j�?#�[��l�uSZ�BHu�
�#4��}��ƥ��1d�I��*��u#.�3� �<��"�@c��I�gݦ��
/�3S�<��"�@c��I�2�����7���F|@c��9A��O����"�r
�,i��J۰;d�]9���������XC�X�=�G��p�g��u�>�#4��J&�{î�1d�p�J����
/E4��e������]�I�]9�����m
ŀ����Ī�ƥ�ÌN��]�?�-��"��XC�X���V<��p��CLW��:�|
X�tؕ�ੇ��c�kc����{
P%!�l#{PE�9A��?)�h>�E
�jq%!�G��/���d�c�p�h�d1�%�8c
�Υs�Ŏ��2������&v��Fiĵ A�í����1R_��sa l��#!X�tؕ@Ĳ�E��c�g��u�>�#4)!�}��ƥ�Å��`V�epY?�r����Sc
�z���]��=�-�����XK�2���OG���gݦ�J
�#4S�}��ƥ��1d���J����
/E4S��e������]�I�]��=�-��"Ā�䰇��Y�c�Nd�]�0��ΘP
	Z�"!ʷi��J
9Ad�q)�����r���F|@c�ٰ;��]y�3��hY
	Z���A	{PE�6A-�d� ��|
�*0��Ī�ƥ�ÌN��]�0��ΘP
	Z҆��F|@c��9A��?)�h>�E
�r%!�,I|@c�ٰ;��]y�3��hY
	Z�"!ʷi��J6Ad��d��!>
�*0�䰇��Y�c�Nd�]u�����m
�Ԡ X�tؕYs���c�k���0Q���
P�,i��bI9A��O����"�r
��F|@c��ٰ;J�]y�3��hY
	��"!�SE��"ދ��B��2��pKo�7�l#{PE�9Aq�?)�h>�E
�jq%!�G&���Gq�d�p���� ��P
"+0�<��"�@c��I�2Ve<j+V��'v��F���=�%��7EJ�kc���&���`%!X�tؕ�{*>��cఄ�T4����#4��J&�{î�1d�pఄ�T4��m
/E4�����i�I]�~�]��=�-��"Ā���Ī�ƥ�ÌN��]�0��ΘP
��XK�2��Sz�>���J����
�#4�K���Y�c�d�`V���ma�r����Sc
�z�J�]9���������X�tؕ�t�Z��cఄ�T4��m
�#4��K���Y�c1d�c�gݦ�J
/�3��\x8zQ����~ఄ�T4��m
�B4 ��O�&���+�d�l;�h>�E
>�p%!�X��"�mc��I�2Ve<j9Ĵ��7��,i���I9Ad�q)�����jq��G��ѻ���d�c�>����
�8c%!�<��"�@c��Iఄ�T4��m
�#4 �}��ƥ��1d�I�'�T4���/�3��<��"�@c��Iఄ�T4��m
�B4�荳�+:r+�q�l)����>�p��ѥs}�Î���2����Y��\7��,I|@cW�9Av�O����"�r
�A	{PE��6A-��;i�d1i��8c
�<��"�mcg����(K�F�qLy?yH��'�5A�o)���J5�$���c�NrH�c��F�Ko��Jx��LE�p=�G��|��z���kmٲ��~9�� p�ŢyH��.�F�KoZ����z�fV��=p�b��G����`�M���_�
�&�p���G��iO�O]M�g����(K�F�q�2AyHFP_� �n���}��hK&;s�r�cH��io���ٟg����(K�F�q��AfH��>�@��ay���ڭ�K��p���G�J�P��f,��JuM�LE�͟NdH�c��F�Ko�����'K�F�c8t@yH��͎h_-��|��>?eV֑�c�rH��iO�O�M�gs���(K�F�q%t@yH���S�O�n�g��X��9MjTvr��spH�J�P�6x����(K�F�qLy?yH�>� ��M*�,�_L%�
��{��X�GT�_4��$z�?��v�o)fBp�ɾ�G�A���/M����Jx��LE�p�NdH�c��F�Ko��JuM�LEWp=�yH�j>� {�)���J��$���=p��rHGrv�66�n�s���(K�F�qLy?fH�>� ��M�g���.�̹����}�G*���I�r�n9�O��J��$���=p�NvH�c��F�Ko���JuM�LE��<��G�J�P��f,��J��$���=p��vHGr�tp��s������KnSpLy?�G��'�5A�o\g���d!Mv'�%��vH��P���o۹��JE+��͟NsH�c��F�Ko��J5�$�����<��,�*$�5A��\g��d!M�L�v�	vH��io���xM�g���(K�F�q��AfH�e�4��-�n��<yB��/Nop0 �G�J�P��f,��>�����f�"W+9����6[��z���L�o�u�	�}s�5�dN�AuNݸ�����̀���$�!Q&l�w@,D��z��\�u;�e�Ps�6�.��z��O�@֗�;1^�y�9�6=D�I�zY�XX6�A1^��y�9�6���I���������f�`�Vq�OR��6�t�ݸ�>��������"^�y�I�I���z��;ҫ���fɝ�Vᤥ�e���t�ָ�>��������c�r}�@�b�4ӟI�YE����֑�j�WFW��e��\
�ָY�����ִ*i��D������n�ָz������;�e��ss��/0�Ye0�;�ؑ�j�WV���e���t�ָ�>��������>s���OB�I3ӟz�Ye0���>��j�W������6"
��Y�����>��j�eM�5��=?�.��zF�����;�e��5��=��.z�z<�\��>;�s�eO�b�6�I��P�������$^�y�I�I���z��>������f��W+9����6�tң��;������c�]2hu���I���{��P����֐��$�خ�;��I��䣹zY����A�^��y�9�6$ͷ���*у�S�ި��(��`k�3��p"ָq9���:��rR�����1_�H��q��4�)�IrR1�����c�I����;ҫ���f��Wᤥ�e���t�ָ����������$^�y�I�I$ͷz��*уZ�)�ڨ��e�Ps�6�.g�z,�XX6��;1e��ss��/0�YE���1���j>e�Ps�6�.���7�X �����"W������6"
ң�Y�����ִ*ic���%�#]�I�ݸ�>�����֐��"�ˮ�;��I��䣹zF�����;�e3���6�.y�z,�XX6�M:1O'bFW+s���ݸ�>�����֐����ˮ�;��I�䣹YE���1ִ*i>�������I����>������f��W+9����6�tң��;�������^�y�I�I���z��>�����֐��"��<����6���ָzY����A�^��y�9�6$ͷ%��*у]3ڨ��e�Ps�6�.0�zF�����;�eM�5��=?�.ָ�z��O�@֗�;1^��hi��?D��zi�\��>A�^��y�9�6$ͷm�+�vX(�О���e�����.ݸzF�����;�e��s+I��/�Ye0�;��7q��ɿ�lG�!���ݸ������U�f��W+9����6�tң��P�������`�r���OBu��5ӟ{�Y-���֑�j�W��OR��6"
�ݸY�����>��j1e��s�6�.��zF�����;�e��ss��/��Y-��Y�ɴ*i�����Aَ�I�丰;����f�"Wq�OR��6[�ݸz�VX6/�M:1O'bFW+sO��ݸYE���1�7q��ɑ��p��o�ָ�*у�G�O����e���C�^TX����_�x��QtLz:�>�r�X�,���_�x��QtLz��C�^T�х䌔^G��P�+�Lz:�C����х����~�f��wLZ+�I|�G�gY���X�/����Lt�lB���pT3�/�������/���M
Lsj�5JTh)<����X_YB7x��ALt�lB���pT3�/�������/�L�M
LsJ0��L������^@%�kovF�>{Lz:�>��X�����_�x��QtNLz��C�^T[�Y����?nukrtLs*ӧ�ulrTm�����_�x���osNLs�1�ռ=���2�V�
"'� t[��L�/��tDN�z���������/�t��wLt�lB���pT�J(�����C2��tQtL�lr��Z�4��!\g�f��LR<Ւ���rG�g���%X_YB7����Nt�_'m��^T3�/����X_YB7x��AL(���m:���iCW����~kSi#�wLt��B���pT�S(Y䌘A�!\7x��L�"T����W���Y���G�Շ%&�NL֏1d��t.W������X�/����/Ot�lB���pT3�/Y�����O'�c�MhLs*ӧ�u�h)<�W����O'�rj�L�lr h9���܇��TO�ostLs�1�ռ=�*<�N�����O'�� OtY�{��c�4�/�����O'�r��hL(�;n��ZWgC㌔^G��@wi#�Lt��B���pT�S(Y䌘A�!\7xf��OZ+�I��_�H�g����X�/��j�wL��lr h9Z���ۇ��TOQttLz��C�^T[�^����?nukrtLsj�5JTT��o�����_�x���osLs�1�ռ=�����^@%�TN��\�>NLz��C�^TX����_�x��QtLz:�C�����&�4��!\g�+�Lz��>���[���	�*_]�u�6Lt��z��c�S(��X�=�~kSf��LR<Ւ:~�I�g�����O'�r��hLtY�{��c�4�/����X�/��j�L��d�z�������~�+�wLz��C�^T[���	��ED�Hu�6{Lt�_'m��^T�S(��X�=�~kS+�
Lz��>���X����=�C2��wQtLz:�>�����㌔^G��P�f��LZ+�I�F�%R�gY�bw�SQ�Ag�{LZ+�I� .�O�gY��@�C�����f_�%��qq�օ�T�Y�Kl�j�7�(�`U!X�%%�T(�ػ�GS��;�L,���<m���(��gC��(_Z"��ּSZ�	�Ks�T _�(~5��ˎ�E'�v�-g^�l���[\|�Y��N��<[K��`ޥA��<�Y��)�cA������9�� [<l��cf�fn,�%�A=�K�����^��h�J�*���A�7<�ޥtfQ��onD�@��hާgYꞿ]�u���/[.���h��T{�V���6���5�@ΛU��j
�c�i���"+g�(���7�m���q%��t�h�9�:��nk�Ҟ�ԷF�/��hk3�d�J�'�kpaӼ
������h�I�
$�I��n�:����h����t���Z�u��b�5� �5�v�эI'���q�fV�~'繿x��O��5�tTLh��
�i���_���:ჱ?r�+��h������f��W�g7O�����i8�x�w�i0��XU�)kܷA�������kR��紨V�Kc��XU��VWNV����NVhNV�'s��B��ǋ¬��hx%ܦ���M��>ߗņW�e7�h(4D	��gWY�xX�M��|���\X���6E�*q4#�LJ��U��M�9���E�9FU��^�WFaY �H��b�RFV���4��c���+�a,>b}���),poR��4��? ��S�_<�3M^�[ew
��CPF(��1�\x��q����|���ke�������9�Α�%�;�v�O�~��(���k�j�Åq�Åq�Åq�Åq�Åq�Åq�Åq�Åq�Åq�Åq�Åq�Åq�Åq�Åq�Åq�Åq�Åq�Åq�Åq�Åq�Åq�Åq�Åq�Åq�Åq�Åq�Åq�Åq�Åq�Åq�Åq�Åq�Åq�Åq�Åq�Åq�Åq�Åq�Åq�Åq�Åq�Åq�Åq�Åq�Åq�Åq�Åq�Åq�Åq�Åq�Åq�Åq�Åq�Åq�Åq�Åq�Åq�ÅqB����e����#A)hڞ���{V����)�7����qښ�j�з����B��/���зk�=p���qښ�j�з��G��B�ؗO���&�ä�Åq��G\۲4����W۲4����_�����I@_�̔S��`�jqdS�W)h��-)�u�g�&�s/��(h���q��q��#�SGh��﬋?�Ih�����5���Ӕ$�SGh}�}�/?�Ih�����5���X�#�SGh&�n��\�?�Ih�����5����[�#�SGh�K��?�Ih�����5����[� %Bh��
(�Å�Vl4��ά4�O�hO*��6�xuI��R��%���Vl4��׬�M�ehO*��6�xuI��R�ܹ��p��q���_������@_���S�%�hqdS���nk���_���J��G@_���S�%�hqdS���nk���_����dq_�$�S�%�hqdS�߲(h���_����'�p_�ƔS�%�hqdS�[)h���_���ID�Rs_�$�S�%�hqdS�{�(h���_��s�Ԡn_�̔S��`�jqdS�:*h���_��Դ"��q_�$�S�%�hqdS�o�(h���_���\]�Ss_�$�S�%�hqdS�F=Zk��>\���U��k�M7��з+[��Z�v�=��g�����Eii�&�M7��з+N��a�v�=��g�����Ei��&�M7��з+���v�=��g�����Eiq�&�M7��з+L�&��v�=��g�����Eiq�&�M7��з1"@^���v�=��g�����Ei٧&�M7��з~#2�ç�v�=��g�����Ei�&�M7��з~#�R���v�=��g�����Ei��&�M7��з~#�FD���v�=��g�����Ei	�&�M7��з~#�����v�=��g�����Ei%�&٘�:�=�kT�SGh�<����?�Ih�����5����#�#�SGh�>�50?�Ih�����5���)�#�SGh}�|���?�Ih�����5����%�#�SGh>�vv��?�eh�����5���e��#�SGh�P��?�Ih�����5����%�#�SGh}�e��?�Ih�����5����#�#�SGh���+�M�?�Ih�����5���=0� 5�)h���Å�Vl4��ͬ�O�bhO*��6�xuI��R�ܭ���Vl4��ͬdt-ehO*��6�xuI��R��]���Vl4��ͬ��� jO*��6�xuI��R�����Vl4��ͬxC��qO*��6�xuI��R��e���Vl4��ͬU*WNjO*��6�xuI��R�ܡ���Vl4��ͬ)�:!jO*��6�xuI��R������Vl4��ͬs���hO*��6�xuI��R��	���������̧��_����n_�$�S�%�hqdS�?Zk���_���y�q_�$�S�%�hqdS�?Zk��FĔ�~�N7��з~#|����v�=��g�����Ei1�&�M7��з*"V�V��v�=��g�����Ei��&�M7��з*"T'�m��v�=��g�����Ei��&٘�:�=�kt"�SGh}���=�.?�Ih�����5�����#�SGh}�����?�Ih�����5���U��#�SGh}�f�c��?�Ih�����5����$��.⮑ԑ���䮑���n|����5����.⮑�����F��䮑���n|����1����.⮑�����0�䮑���n|���������.⮑��zv�q��䮑���n|����e����.⮑���i�,�䮑���n|���������.⮑��؟l���䮑���n|����a����.⮑ԑ��5�䮑���n|����͗���.⮑����@2�䮑���n|����z�l|�.⮑�*]�5�䮑���n|����)����.⮑�o����䮑���n|����՗���.⮑�	�",�䮑���n|����ї���.⮑h�%��C��䮑���n|���������.⮑���y����䮑���n|�����P���.⮑�	��0�䮑���n|��������.⮑�֧�p��䮑���n|����i����.⮑h�lP�1�䮑���n|����Y����.⮑h��8d��䮑���n|��������.⮑h��Gd���䮑���n|��������홠����w�;�H'�l|��L����Դ�����y��;2 ��+������/����b�l|������Y��;2 �>+������/����jGl|�!�����`2�l|�!/K���`�@l|�{����2}���}�];28�yL���b�l|gO�;2u�5KgJ�<����t�*9��#�'Z�����x6�0��sJ|�;��>2?������<:D���w�;D���a�7D)B����Vu-������5����e,-�>2���B��9�L�����e�B�Z�0۞�D�x6�4�H���h��o	?=�b�l|�32���(ʣl|P	_;2���|�)�H=�U����8����;2���{�B��;2�Yl3S�;Q	U;2��`�o����J��Gl||9Ę���.�d�>2�2�噰�0����!j��ހ�������9�L�����e�B�Z�0۞�D�x6�4�H���Zg8D�1�+���a�T8D�X@��;�z>���>2���p���{��=��nl|�`��0�������m�0�cr�0 �I=2�p|1��;}௲Y�e8D��12��!Hz>��Z��MW{�Dܾ+>��Ι0���|Q�;2����P-w��;2��;2������nl|�{����2žï��6Cߙ��ݑ���l|�ɘپJ��\�ɗ0���K��(j�l|T�XU��;}��ZP ����X��H=�!��ހ�l|eM-~��;2�~5�H����;�)��H��)B2����s�d��@*B�����݌6�:�� ��P��/w}�7D�:��`�6��Q��+]�?�nb����+]���nb�y��+]�Z�c�m��+��A"fb�����M�.?� ,��se�	��/��+�1�+�������.�1�+����ih�.�.�+������=3�k���ڲ������+��e��H���=3�d���ڲ��A��k��+]�\!f���+���쨱����2���+�1fX󝘹2�2/�c��
�.Y�k�k	��k�y�n/�.?"f8����nb:�=�A �=� �ę�b�2/�c��m�.Y�kak	��k�g�n/�*\!f8����c:�=�0B �=g��ę�u2/�c����.Y�k1l	��k��n/�F\!f8����nb:�=�0B�ڲ��:��!�c:۲f��7]־>"f8���@�c:۲�$�7��QF�c�a�k�I��k��n/��>"f8��5&�c:�=F3B �=k��ę�ރ2/�c��}T�.Y�k�m	��k&�n/��>"f8���8�c:�=^�A �=���qo�.��d#��=��A �=C��ę���2/�c��E��.Y�k�k	��k���n/�J\!f8���A�c:�=�#B �=���ę�r�2/��p(%�.�~ �=���ę�v�2/�c��i��.Y�k�h	�
1ߥ���/^R����PC;M���}��4�ഃj]R�-��Y�3/
gt���
�/���e
����4/
gt���
�/���e
��}�4/
gt��
�wt
��LiMI_�Æ/^R;��PC;����}��4֨ⴃj]j����}�4/
gt���
�wt���LiM9_�Æ/^R|&��PC;U���}��4�ⴃj]Z����Y3/
gt���
�wtJ��LiM���Æ/^R�]��PC;����}��즦����11�o:��/	�wt���LiM�Æ�0���/
�/�:��e��Y�4/
gt���
�wt���LiM���Æ/^R�F��PC;饑�}��4ഃj]~����A�4/
gtq��
�wt��LiM���Æ/^R�E��P3-蓍��/~��.e�Mp<������/e"Rk���z�[.A;n��v��/����������/e"R�-�y��[.A;�@���4��/@;�@���v���/~ �.e�.e�/�M4d��T]��-�Me�����
y��*e�gtY��D;�/e�ut��~�.e�M]������/e"RN�y .X.�u�,e��ӫM�e��zD)X.��q�2���D���@GѫM�f���V��,��)�y��/@s���0��/@)�u���/~��.e'�x��Ю�4/��/ev����L^���[�5e�uL|��o�v�[.�D���q����L��[�4��qt���&�(&���"��I����/e���A�4/��g�[��G_-"<����/e0�~��/e"�=�����/�e���A�4/�@�e�w�����D����݀��bt[!׻[���-"<�o�Mty�ÚmY3/^Rty�À)#zF��� R����_$Rty��_�\c�[ �ewٔ#ڤ�/�~��e�D�g����3/�ME��T��R�g���q8�.�ME�Ú-�4/�oe�����ջ�o�4��⴩u����4����/e��Q\��/e��)s�[$����4��qt֫�λ=.�����4/�XĮ��4�T��[�z"���w�֫�Dˤⴟ0�DG@�U���/e���.���=�uB��\��q��-f��/�DG@�/*e�M�g�����E�u�M�g���/��/e0/�DG@��~�[й��uB����Gഩ��L�.e6#DT���/e0/��e���ȸe���Ƚ����4/�듖��/m��.e0��_��/D<�/e�uLA?��o@nT�De���o�Pd������2��/�%T	��.e��$�6X��:e�/靥�e�De����ؑ-"<s�wt֫�u-z�yK���/e�Ի[x��4/���Yy,�X�����4/t�e��̰�/e�/�_z|��zi�[.�Z�/et�e���q�H���m�7(���`��>�p2(
=��\
�>5�(���S�(�Ğ��>5�P�xU��\M\����\M�����!]M�����\7<�����\S�����,]7�����FSf�����EM~����Z7�����GS.���Ћ��>,	�Mb��>�w����>��3��>K���z�P�0�!��GV ������Ou���;��>��#�(��]�z�McQ�>�T�S)�
o	4fY
�x(԰���
5WV{]{r;��P��� !c�ʨz��>XuO�z��CUSO��`�z�~���IQ�>x�Mc��>��"��B��D_I��{��IQ�]{�?���J����(^[��}̼D_I���)&6P�4��>OŴ$e�֗����BB�0? !���8��h���\7L���EhT��\((���[��[_��>�����Y�?���֞��>Kݴz������TZM������EM�����\M�����pEM������EM����[���)fᾛv�����>J*(g���N�J�>���)m��Ob8�>��LM��(g��"������(�&]M�������>fu�<V{�<���^W
�Y��a���}�lᾛf��P��>�\��y��>����h�>�������>������>���#��>��B�V;~?�%�����uU�l�1Kc�>�}��^ !5�D0e�P�c��N����Wt�?���%Wx�=����c��E�~���{'O0���[������l�A�y'��?�V;~?�)���uEIf�:Km_�>��RT@�>�u�=��:����>��P��^ !5�D0e�(y_� !�\M*���E?Z7��|iF���A��|Y��z�BY��X��4��w4���|Y�v�|Y��AQ�p�8�|���^k�)��z:��q�.�8vzwZ���q7Z����u97�vJ���Hq��Y?Kd������	���\����[*
Y����i*��������[�vJ��� g���Ϲ���i*՜�ހ��DY�t�z��[��X���B��^k�)��z:�ɜ�x�.��RXE�|oF���|iF^��|b��7���fZ)9�8UX���|YF[�)�8�||�mЇ��)o��x
���RX��|�^7��ٶ.�B�"�ź��������%|B{�F�>GY[Z)9�E�|��F�H���j�X|Y���]|Yw8�����|Yz��_��کk*
���A!I��C��|YޡH�F�\�G���|Dh:n�|ٺ�)��AZ�U��:�*
�O>Y�����[*
H�FY3�H�X|Y�HO|FY���g�ΦK"�y��A��2H�^|Y���|�}�vF����z�"�#�	
G�m���u�/���|Yu1Ƌ�|Yu�/Ƌ�|Yu1ƃ�|Y�A_vzOY�����4�v�|Y�}��3i�[|YlG��|Y��*�|Y�|Y�1Z����`�(y�(b�"�G \��"'��(b����A޻c漺�e'�p�(b�Ϩ��&,1�l��l��x`��l�a��l"�h`��l��p`��n֘�'��(b�'�0�(b��'�C�(bq臒�&b������XЏW����(��Y)b���
Nux���Щ4�c����Λ�NZ#�pX-���;$��GX����;$��xU�h���A�� KOz�Gx���Щ4�f�(b#h|��A)�#_)b��ΐM�O���)⭦�l��l�Ah���'��l��)�`���Щ;�N
�&)b%�H�W���0���A�WYF�l��r�6���-�>��%�� �Ob�l������4�a���W�����n�6��G��������u�u��֛8�Ou�\n��n�)�7��m}"�� �B��"ub���k�Ou`�a��ۦ�O��%Z��"�W�X�l��:�5��W+����g�n�A��#$)�a���W�������6��G��������u�u������Ou�JR��n�_���m}"�� �B��"ub���X�'Ц��,hQ��A)>���uml9n���?h�����3{0A^KO�W�C���Ґ�So9n���?h������J0A^KO�,jJ�>ۦ��O�����?\���ND�G����O����N���l�A�᭦�l]#b���[cB��B��B�a��b�c}�b��Q��N��A)b��'u�(b�X)b�Ԋ�@[m�9��yyKaa������N��-<��)ܦ�(b��-Kܵ�'ẹ�(b��-�-:���Y)b��g��ώ�u��<�%�h ����g[���+�~�G�5w�S�����!���rkrO���iheD�a�<���2�j�XG�4���C"�=+�YW�������/�i4��W@��z4�@��C5�!��1H���4���1�b�U�3�x��0B$?�3����X��B43��!���(�wN4i4�~X5���M��\j��C��\�!�=�^��L:!���ύ�A�1HӢ�D5�8����/i4����d�d���5K��7h/�i4NZm�(��,m$W���BQ���N�1-���}*��*DpE���=lJpE$�:��vE�o�ds
�Mʉ6+�6�#y��3�![S��v�;{ �����E���u��h�L+DT�Z����vE�Z��8/�5�R&���W}�~�P��H��p඗�n���vG:����?&��J��ެvw*a�a�v�>��(��� T�� �яF�Eɟo/�-S�1WpP�{��+��qw����eB�va�%9��!HP�M	޿��`\(���w#pqE�I��qX���E��f ���u��*�o R7�/R�,�uxݧ6E��p���pTnp�Z_�|��E�"M�-�E�7�oCxt|~�fű7����ӂI��mߍEop����u��o�:�V���C��L�,R@pKjdL�q���$�X�a3�K���SI�oRz=r0�c��951&�qw�\/੖�vVS �ݎ�5^2�&����}���w�Z(qP�{���C��e��H�C��Ǖ�p��{p
BD�oE�ԋ(�R4�}LR�qET�o�8��V[�L{���d�yK�>��
�:RW�y�Pv{b.|��?�x��L�wv��Q)���ny@���{�Vى���.�C�c���t�E�2�͆�JP/�)E�w�26.��-�5!t{��x�6�"
�Z17!�b5w?�e�MΨ��d�뀿x�>� �]s}����Qb	^����HC�#��~m>�=y{^�;?y�8��-  P.|�蠊[ƈ�[���}��	��+�Ϸ��$5�𵅆J�>)��:;?U*@�-W�ՓφT�F���y"55�.0U$,A�y{�\���6��`��(�w �{{�<��o���z�0���k<y�����������/�߇�X�z�M�\���=z\�ΆV\���f�СP/�ӧ%�{yM�u����y���('0K�,<c_�
�vA5�p@7��i\m�wQZ2�,������V_qn}�o��(M)�uo�N��yR{ǆY
2�WE'�yN+P$��B�������J4mNf�> �odzE}��~$y{dZk�*��f��>Vy�S+�z��熇�>���3@f��AuӔu�-h6y���.���I��y�x�6gZ�����x�6�u�]�9�!���x���l��JYKyɵx������~�k;jy{������fĪRg"�tM#�D2|��x�6u�^`N�x�,�=�#d{d)ѲZ県x߄]��dz�{��x{l6SP��xp�il��L(�A�^����w{W$	����p��w���}���e5x{sy70��E.�xsY%���tdUG�p���L{%AY�~�x~�`��vt���z*z{�B�^8�X��$�  m�N��r.A{{��ɉ��=D�w;�kdz���e�y{�y��^y׬|�m���v�P�"ᭅF��<�_{N��\=���$l�������T�]�:�@wt�s���|4�9yF��P{NI �y(c3��7��.��Y�̤585�8��q�µE�f7@M�[]������� �`����8�R�4#l������UV�:�@Wt���i/�xB��M{�C{�����I{>�k�z���y{M	�ᐢ���Q��!�P!�	sƆ������)�"��4� 8(ʽ\�H�+jy{��h�
f��P�W$yh�RKD�$B�U~���Z%��v��6��}��D�+{y{IE��J-QK��x=�v#����=���І�o�y#� ܃{a�g54���:Qx{l�ZyM�O�����}�����gy{�	%�Δ��[c��~��
y{��,��`{�5őKCO���n�A�c{t�����W�tP�òsmF4�~4a�y8��F+�x�4�W�z��),~ty{P�5k��)`����D)���~y?��w{[^�y��ӔF��zUt�b�y#�u��F ���w�&{7T@$���Ny5�{��v���7%y��T�a{�xF\�V�O����,,%yT�"�.�aI�6:Y95��L����K)y.ow��x�Q�?�V{�S��Ty{yӪ��!y{B�t�`y�d1�v��!y~Bss�"t��`�X2+W�$������A�@�3�K(v N��̊t��!�guW��u{i�m�N�guW�m�9B{{��!݈T���T��!��y{��u{�trIy�����!�vj�3.]�P{�X
`�3.]>+/]y{~~��Kv�v���ȸ��T��� �6A����e��䮢��
�{ɜ5i9F.ک�ڲ��hv_0�Ӈ/�@���AL҉3���
��J-9�
����MK��	�C��/)�S���o!;+5w�Q{O{��y{�{�8/]�~\�Kv�g�.oX��y{�1L�\Q>p)�N{z��$]�o@�mC��y{nC�UWs�_"IWW�	���.#y��.x�wey���w{��V��T{6�k��8K$H'�K�݆�\��6����IJhQ��
5�vV�������v�)���3�
ۚ�rsy{�m�w�o�՝�Y'Q��LŘ�n������0�C�{�P��_���f�y{�\F�mlx�B2-K�L�rW%%�݆N9�Z'[�cN�8x-F\�[�H��$��m��on�h� �a�Sf���tM{������EC�;c�H_xߠ�R{d1Q{b�x;�_�T!y�V-�X�s��$_N��R�΋;&՟lA��t�%��JC�}�K��$`N@K˜���7I�sԬH�dm� x�b�w��=v"L2��p�t�ch��c�x�k�����u59H^u������ <
��X���Ɍ�st�
~.�d]����%YԮ"�\QEu�#� �L�k����̔9��r['2Hbu����' ��@�� �� ���í�s弄dzguj� x�E5�
!+�*u���g-��Ȳ��V֯�Wnw�t*��t��\f��Z�r�ꑭ0-���m^h�s<��sZ2*�ʠM�����B �JOm�s��N5X�����n��vČG��=�t��Ѯ;*�ӷv�Fw�>�?�Ö�IK��_u!�5�9�JX�F(�Y/W�wg�%�iu�,tVXPh�t_�i뤮v8� �A�tF]I;�d@ �� �U�9 ��Ԯ�s��NTJ$Q�ZVS������~���wu �9ou�/�[� �xd[<d���s��|e�w'��XW~�Y�Ӥ����t�!��
�dO��VW��@�X­�C+�uډ�+6��e��Gv���c��s�D6u���$��Bl�<uJ��,�����4u�2���]�n��~�Y�Ӥ_��*�t���>1nd�	�SEuEh�ɒ}�s͛���]q��d+����00]��s�-=��
�N��9�R��s�3���)Su�1�E��Ć&�|�CN%�s������u� ٺ0���Q�n֮o��	v�τ���t�5\�&��F��q�Խ����I�"�s���>i3u�z~�<�3�������m0u�4���s)T�nE�w�����Zu���C�!�q�rmo��3���t�F�xj�`ug��᤭� ������u,��s��V���~c�.�o)��Q�4�o�s#����������K����� �s�����!�	
����u�|�����t�w>M��)�� �RL�vb�bs��t�a �R!t�m�s�����<q��(1�s�#1�̰O��������%�H^u���C�!� �̥y�ݢ�k�yu �0u�����Inu��|��g��<X �g<79���hB��+'6��S!\��nh�h27��}c[h�v*[�z����:O�5�gA��8J�q�o�1�nh��hh��?�Ve~cC.�z.hYI\���|g�g���EU;���k�h��h^���1�����ۻ1�DL��T�:ht6�����C��W�<P<��VN/�h��h`Q1	��_� ��S ��3_���x�hB���IhX��1)�u��de��n��gҰ�g��V�@GV�]���tq���g*d��D�c�(z]�d���h�ahgl�`��dH���f�18ɮg��Mnhk�hC��_CXVh�0�g\hw)�hH ����Y�R\@8�n�\h��
�g��+;b'��h
,�C�hw�ؠ6B[u�h�/kl���hU~�l�Y!��^k�{�iP�)�g|Nh>��
L_g��O�<_e�g� �w�gQ1���h��+<�s:�2vSDҖƮgr��_-��J�J9���X����gX����3�g��\�� �l*�T���\���3l*�$*���q�g(�	�[|b����K������C���&�2��)�-\*�g�>��g1Y��p�]�2�5��V�!�=���\���3�g���b[|_��\��g�n}��`_�0�g�u�,��`_i�`_��g��F��g�'��dp���}!��� ��b"Y�h�+)�/�̪�z��	�n�F���s|����C�q�ЫYNe�`�2N\�"�dY�;IRb{��D��btkl��
v9�&Z���k�O��.���T�g�܎Iv��+�gtH��g�-���`_�+U���bf�#2�i��G��%7�-V�Gt���^mT���&�	�g��"�I����hr�H�\�=V�j�b��������� �܅������,~Sa-�\-#5�]ֵh�X�Q �h��%�=f��RE  ��J���R4��9K�M���d$���>oh��_������;����7%����k#��祅R.���h[�}g��h�_o��j=h	��V䝄����i�f�^�:>�N'�\	�WKg��Ǯ1W��r}Ţ%�'l�̓�N��h���8hEū�8����֔�������6߁���_�?��R  ipz���W�}[]��h6"�a�㮊a������д����ԭb�	��7X�ц�5������uj�- h�X�b��j,��w�0�$�^�'�"�ծ�-ƺX�Z�{�������a�
�?5Ű��.�������#G���[��~|�����{[Hr�(!������),�k����`���v8=���)Q� op�$����L�b��@�/�����Ϯ������g�gĎ���|��R��ic��"`:�k�/klmy���N}�?������?���Tz����8-���^��o������^���gj��g�'���G��F�®y�BPO�N�nъ��QUӮ* �j���#���� i�XG�.�hcS�}�\�1�Y4� �+��~x8�"��i俈����~���5�̙�V�7����P:8�k��A�L�$�1�>) ����S4u�h������﹫�Q��I�_U��^���Ų	?p��8|Eک�1`��h��:�Yu��MEX�e鮃t+�N+zZ�c��Hd�4H(��7Z�>�O��A�m�����-�Th�=F_��^H"h���
W�ǭ7:,�k�2�ɕs�l��6��2�^x���W���実Uޛ�b��-+���h�`h�L���ɮ�}^�h~�Ch�D���x��g�%�ɜ�G��(&�j�_��d��N�FQ��HUѮ�20���ݷWh
[�f�oW8?	�cl/��7MG��kd��������� �_�)IR� ͂�e���ٕ}����
H�)"��h�?XW���C���*�iog��j`��j��m��N�4U�^�ic������-��h�0^�������I_Y-�[���3�ݕ�h�/. �g0�a5�V���v̮jO��X ME)��J�����`|7M8���g��g�'���E�0�(����M�}Ѱh� a�G��h�Ů�z���&d�d�g+���u�UO�T�1x�y�Ou���,�y7һ��5��}������hF�����Ͼt����E����ƭ���]�h�>��x�����j�y�/�b@�x�������h/�S��D���e��D��h�R��� �T��Do?7��� }��X��O�fm�h���꺭��U�ʽ��\��UJ(7�I�g���>���\����U������hh��^�����|~�h����U�Q%o�>�h�z�_��gN �gp�L*�LK���	��2x�i�-[\�����Ķ��qj��?�(!�#+rE��i���+j�k��ȅ�x�(O�p�I�g}�R���S啿��m�]h�g8��hb)�^����Zl�\�h)
o��u�B<��{��ugot�kP Lze���_,+�e���`d�h�\ٌD���YY��T�0k�Ia���.���K������	)�� ��!����V�!5_~jh  �?䭔�[����8�,n0�9$h�6.�GB�X��8w4��٦wm��\^[
h7��D����g�J���bm�k8�jyz�-������'��������q�����#�_$��ɖ�7����Dū*'w��A �Y�����֮gD�$�-�E��xh~��w��d�h���i��H��̗�Z�Z���,5P�=�����
W��Gh���p�z����d�d�g���X���lO�=�{n���>h�YM���X�������;.����J�`�Y�ѻ���ah�'�T`��s��*}��=�Y}��8��.nh�D ��P}��g�%�ɜ�G�2�%��*䑍��h6����ЅU�i.3�m�����)�D�jc!5�]�Ah���U��w �cB��/��Tr���H�h��x�	��r���Ü�O��UN�vh5�G����A�j������#G���$�=������=K�h�D����)���u� )VF��%����#�i���(��ye���;h<��d��8GO{[]9�j��N�������j޾hX���C5h�yxl*��ul*��HT*��Q$J��0���L�M��-�:�[����a`���]#��K�g|*���
�ge��\���L8 T*���r�g.�	�g����E�s��]"�g|��-�mϧp�Г���3l*����3�g��\��v�vh�s|v�g���XYV��-�e�6��  l*��\��3���3�g��\��A�(���Y����3�g��\����F�s�g�����p���2\w�ׁF[����3�g��\�������Q.�	�g�I�gl*�T*�-�*�&�m�8�l��Z {�c��4��Q���:�!�-�	�gv�kh�{��7�g ��ǫl*�-�	�g�+��?�k�\
�g�3����g1�-�Z�-�	�g�J��1�R@[5�g�ۊ�Q.�	�g�I�gl*�t*���$����-A7���&>��xq�G�졀����-�i�@�hV����3(�	�s|���1�9���\���3�g�c|b[|_��\���g`*��Y�`u^^T���;�]n^T��Z�����5R�?Z��Ji��P��Y����[]�/Y�f����`_t��6�Ag�W���lo�1F<P7i-}��|L"TF��^s��\���\��cU�1�&�g�ZoM���)��[q걇7��S܋op0��yv`��6f��J�g�$�嗫V�8�g�����|�+�gȲ�[#2j@u���bP#2��te_�o�d �^�O/&�(*y�Ԉ������zR�����R����g�� �X6�^���'2���b2�#2(f**����FxR�&���g�ΖR�*���fݶ*�+����m��qh ���^��L�52���ZM#2.��.�g�p�⸚�R����g�� ���^���'2��l\���`_��6O#2�Q�`_t>�
�g.����k��k�gM��y��m���N�Rr*���|�=�$��.�^�g���_#2��h-�^t9�
�g.���Êk��k�gL��2k��̈́4�^t?�
�g.����k��k�gN���s���^�_����C���&0$��G2�����c,L��|>x(]8壵f$����x9����]J����ء�7�{ZiAĝ�x���S��BpU;�E)����v����z�`�nT��:=���E��ҏ�G�7D���s�Y�:�w��~r�9_8��Sa�w���[�)L�s��B���s���z�����z�R��Z֩���9�!��G��Z^%p��=�:0�:`:�hԔ�
����+Iҟ�;�c9<L����T�ͫ�y��5��yu$K�F;�����.����
;�S� Ԝr�5J�:D� 
&2;��C�F"<N��:Z�m�1p:#�ph�r:ER�n�9l=H�Mu�� +�:��Ĵ���k!��!B(��::-�2�:�%d��{
��G�"�Κ�:c�;e���u����j9����m:�L8>�:x��bQ�F���>���:��m
�-����I�_ ��7e<�E��:���C�Xl�ugu�� F�u(���r�:8��چ�?w�r���:��?��:'Q)�e�8
l�?K��7.u
�� �:>j�s+]GZ��]�*�$.�\��:��:�{G��td:.�8�=l���@Ŏ@�y<9�!��"V����v]@A�Ýr:��F9G;'�b?؝]�-�X�>P����:nA�	�:����5�JTF�RHv:��V��:�㾱�l'=H�O�ZJ���:C �{��:b����'.g�:x��:[��:\�1ڝr����w1d�@/� h�:���:�h����h:�67mZr�'�k��9�:r����T��I�YpJ������U(�(<'gP뫤�9K��FKx>��D >�i};����ˢ��n�W1,֯����t�:u>�l��u���)m)����:4�"�:&��*�Ud��W�d4�R�z�B�����:��:ٚn����!- MLbF�F��:|�H!�j�;�jȒ���2XF[>�N�:t���`:4��ڥWv�7��f2� ��<�ϋ��j�c+��dsM��z=�:no�:���ߝ �j��,IIjsؚߺ���:�d;��zP��&Q ��H�"�:s����Cr��	�W&4��m+7<r���R��"V��s=M�p�ǚE��:��u
u\��N��Ț���Ɲ�:���'���9�
=�f<��N<�i:�
\�>$;��Ω�U��;�i�gn:�L�:X��� :A�q�8^Ko����<<.Ֆ:��=`���۹�FS���B� �(�JK;]�:��?�:x����k�ʀ�m�H�V:�AE �|�>u%<�<=�����Z�:� 0�z��zW:wr���:���>��:d�V8G?�/"��J��i�6�����:�� ��6oC��G^mE���w�r����:R��:�h�?��}�r1�I�@���<��:��t:���9��c��A��y�J1Au:� d�
_PsB�U�?:�v�f<��<E������qif'=H�O�Sk�:K�c��p���5�r*��r���V{:c�;�ȼ������B΢Ƥ�P��)m�:l�B9hlEl�� �>{�@����$m�:�t3:w
�����@0C귴� -R�'j:n_��mF���L>0�!�V�R�X��V:�E�懤�UyAQ=����^/�:�L�:_r�Ӕ�ʸs���C�$(DH�Py��:�=��q�ȝ ��nWs= H�ju�
��:�����l�ԃ����[,*�Ʋ����y:�����*���Y+.��T�O�#�:OW��w��?���]�D�u��1�a�C�q3<��;�½������AL����*'U�:o������9�(\ϟ��60G�n�:�����@ A���D�L�t,�C�o:���IɝG��04�����䳞��:h��%%2*�(�?�?.��-Y<��<��3X���Q�¾^u��`�y*Ew�:��?6kM<���U�<�>�X���m:� PHs���i@;�2<�d��Wѹ!<Y;�n�sn�a:�8+ �{]��\d�:��<x��w��,�2p�K���D��"�:�%�����w�Lz;>�:X.����:��97d�ҷޝ��pH��R�{(�:B�Ht��;��!�Z�@�8=<%�̰�8\�9�r���:���>��:��J<G?�/2��c��l�6*��Y��:������6o�8,p�fE)��w�r�5��:K1*��9�p�JC+�-�dĚLH�y/<�O�6|Ý�=l�'; 53[��s\:p6�Z��� ��GG;��$�����<�9��ٶ�����2�8�<p ��~�:1��&<���f�5������<�n�:~#���l��^"�YM<�>�o^lN;g ��(%��"_u9�z�J#�>�{❱<�mqh�WTe��6�in�9ذ�J�#�:������	s%�r꞉�ʸs��>��:��S;��� �l���i�66�J���:YG9G�%�b�S�aE��wd�j���:?�	�b�s'~�td:c|:6,��t��:]vi������AQmr��픗�k��:D	`v��;�V�b�a|=��%�W�6$<wnbs�nT��ڋ�C�$	��-v8��:I "�w�U�]��U�]͝)��<l)m�y[�tu:��C'g#��K5�<��@��$�T�@P '���:�o}:]��ڝp��ܾ�H��6N?B��-�:Dl���9���1����ǝ��:s�w�p4K����m�~>�:�7��0�:�kQ+"d<ΪT5�Fs�J�dg/���<J ������1�$�i�p䊗��~�چ:�{c_�?�I�$�`:QU� �V���:����2|;�i&���㊗�Z۝ŧ:�Y$�4��#;����V���T���:"z��i��9	7�W�3�g���k:���8�����A8��Q�ݟ�R�� ��:A��V�d�r����;�:�
�l:o�ߏ��#�0	���r1�I�@���;�;c�:�;� {�C΢�����)mr:%�KCZ;P��X�fH��N�w��:U��O���-?��\BU������y<M�>��n�W��	!F޷�:�ބ�:�(|8l���mhJ;( ͸Jsy�o<�Y:9@
��[�;g�a (`"���?�E<��:%�zJ{�!�+Cb:j����<@�B:nl%�r�P�"zR��c&m�:U�J1p�?���� MMΚ��mB!�:[�|��l��/l���|��d�T��:_��;2:�?���������
�YF;Y�BnW'<�X7/"m�҉�����!m�:�S>�����!{y��@e�:Z��:=�:����ǟ�[���Eec��:C��g���.�'����'����:t�����YE;lZ�*e��Ɲ�a:9�� �ܶ���� F��J�����:��)��ED�� `�$@�\�<��<9�F��t4u��8-
LԎ������:���IѝU��l(��(![	���:P�����2���!�vC󦮵<�y#<_"������)�u./�)ؘ��b���:i?;!o]n0:<�H�A8��}=�:��"<�qu&�
�z���r�I�@X��>�;��gh�:������X�>_�ʝ��:�{K_��l� '��;���x�����_::�:�tEN�-%`�@/����:��:a��6:�TzsA��QT�3�a�m#7<���Iɝ#U��6����ip�y<�8��K�=��8��{<x�Ev� �:��75�������-���_��\��:��3X������i�����:������:��<��փ}������Q�ݟ�R�� ��:r���R��U��)�Y5I���t/<b?���8e�
���m�:�M�:DI�����(ٺ�d������������:}����۸(���&�C*� �b/�|�:w8R�:M�:������ǽx�:xގ\� �:^	뱾i�:����]7�?�HL����:z�K:G�Eo2m��3��픗����:t���2���n��%g�2�h�U[:���:�
��<$�U6Z\)��V�˺5
�:Er����EZ$����EA )�wT����:SQ���:�g�>'d��l.5�����:�F���������r���:��?��:I�J�{TJ��!1[��y'?�?C���:�Kp�zS�:g���	\�(���]t�qy:B�ؙ"O�:I;`R3�d�:`��9(��:t�B}�?jng�:���:�&6<��:��� �#U���%XY�c%����)<R"���' �	V��Z9N�:��?�:�7rEf�8����p#�@M�UQ+��:�^�N�:�� 8��2�\�u�b�lp:l룾��:	K]���\VV[9+ �:nI7�d�;@�t��(����º�r�:�h�����:���Dn�:~#�,=�:|n�����f"<��Кp
lp�m�f�:h������+�љ0g#��b(��n�:�<�:'��x��Ν�$E��ÿ*��aO;@�W0�'�kI�v�J)����<7��:�kQ)Ȳ�9{M)$Y��HΕ??h���:�����Q��w Zz}pT�Ne�S�:W�� �p�m�h�@��2��N�:�L<�^���(&��`NB�$<* ���|�:^[�:=� K���̗r�I�@X��>��:m�;@@�zP��� �//��><��"�	��X�9�W� �h�/�:�O�:y^C9�%�r�P�7�h<۫~;�R+<MI-<z��N/W:�:M< @�9>!t:4�!��"V�� B��O;n ��><"�$�)�n#Z��r�!���z���::r��3��ʻ���Mti M�nUC�ˌ�:��3�s�.���h��J�?" ɝ-�:��A�N�{8R�|�*A<����W1��:X�85�?�¥�$�*���֗򎷞T�:[�����?SrC�>���.T/R�:�J6CM�8���q-?E��Òv,��a!<�����t-�<��Gsn�@K� �&	4�:nS����pw�8�
�1����/�:�l<G����T�ډ��h\X"��>�:֧�:y|����`>hF;�QE:������:���H�o^���UGQ�S�R���<M�%���N�<,�s0��=g�:��:Z�j���u��t	��z����ZB��:9�Q���u�qQE*k@���uE��:w���2����{�-����gN�:ֿ;��@��,<�X��dJ�E�Ha?�%m�:�iO7�$V:��v�rv�����k���:w��-3�`>��:��M�VJ�mD�:���:m\�渒/X�8�1�E۫r;��<�A*V�;ï�&H]$���:��v:&~<���oRm�X��(3�{�g��:r���R��AU��1�7	�_�C�~:��-'o���A$�h B�uú˜�:]�@�I�E��N�?>�^?�:�� $�(�:'$�0�������NS��:���6��:h�85�/2�o�H��B��@���:���IѝU}���q�T��R��z:��/�v�9�P4� C�~.�:�x#<�`��m#k:��6�lG*���/�\d�:��G;G���R��"C�Ei�'3E�u�:r���R��"G}�~����,��<rI9*��!<�`��&[�/����/<�L�:�}���V����Θ@�V(dh���x8<��	�t� 9E33����{p���:�Y��~.�X�v���v�m�<��Ϟ���:�K��A��ʝ{�����ߖ��k��k:Pe<l���"|b�_.��YV��<���:R�m���3�I�M^Y =�7%�:��:]���Ą�?�}�r���:��?��:<�F;]u��N(�m��j*7(�:���:S0*삯wG���OF=)�wTsڼ�:�J6C�a8�>���b��l����:9���I��G��^� ���R�D'�:����7���:r�o8��]�<��<���8����Y�]X3�-�T��R�~�:�)_9���~/*<�6<��3���W���:~B�
�py��h���9�T�a�Н{�:_nlp���0x�[f�0�?҉��-J;w^G<@�E^"|��5���a?"�z��:?�u�8�Ъ�5NO ;td����z:<8��E{8�����@]܂�I�fH*Ԣ:`1�_Β�z�n��1'��XZF�Zc:D�5<��i�M�<vl>d�:��m�/�:l���ۅQ����_��­��:�O#<���ڍ����p��< �%����_:��=������#ke��.�����:h>
���
���f��;���$<�N�:8�D�Z�`Q�ȓ�]M��n<nG;�u�hރ�J� ��E�>�[(����:K�䯘�s S��ތ^�̝�E�E��:%mC9h���^��@{��>,6��:"�kK�Wgy�+�y$AnAI;2U1�Jh:���IɝG~�9_���h�Ț���: >��0<~��ug'�JT;>�R���:��pԔ,u���mGԁ;#��aM;��uj���r�	�%0�w>>X:��:q�FΒ�z&���V��0�p>>X:�o�:�d�
�sb�f���3������:�+�)f��Z����Q��I;3�:E+o�:w1PH������:�`R�l�rYK�J;WG:@�un�NX�r�I�@X��>�;y��9m\���弝��F~ȧ�`:��m���ӆ:�IPuiM�m������:y ,��6o��#At^�c/BŎ?��<9�!��"V��P~<�8�"�0�:G_�8�%�R0��h\����ne�z���:�)�8�g�d�:�o����S��:>X=.2�i���)3o��:�� �]<M������ܮ�a;r�,y��
<�:_uC;G0'h�!˝Q�6������:� w^?�:�V���=W�:0��(v:[�]��W:�oMl@����*�خ�!:<_"����' �	V�ڀ ���*K�:F�!�B�$tJ�9U�p�$�B^�Q|:����\[|;�i�74�Z������{:SB���i ��"C�g:h"��|<����`����iI�
��k��q:�O<xj�@�<p��=Ya⎂��R9K�]�:�<ί��h����J�h
<#Ә�:v��3�V�:~����],�:�0��Hv:i�9�d�:�b��6!���O��Bl.��:r^9��G8}}�M�:~������:�Y��~��v���r�I�@P��;��:�. ���E�ۓ��c]i D�su�ꞝ�:>�t��p�o�؟}�:��]Y���:������:���$y>�:_ �
<A��6��T;{��@Ls= M�G�?�6��:k%Z��&��U��r���n�nB�<!}E���|� ��NOe$0�4�N�:�1���9; �&��)`w���}�:(�:@�����V��l�R;�uщ����:m�S���fa���r1���:�.��<��:8[�.b}����\=r��M��:��v:V
zt~;�:�Sϱ� �n��:�_���<I:����9�O���-<����}�:Ӈ�:j��63�UzT��&+�����k�چ:Kl�^��� ��*M�D�G�E	<�K9�����ڝ$#0$uy��4}:���Z� Y�z�y�xa;Y ��$��Wޕ:# :�������C��8��]�:��:B
�F��'<�K\_�* 麏 ���E;E��v�t-�4���e��(��^����:D�w.>>�:��~�`�x�����:�os::[���Ǳ�F�=:����?w�~��:9��^���:�Bķ��F�����|vz�(V<�� (n��G��:���:�u�&B�(V��v���4>�K�r\x+�i�(6���?/F�t
D�H�֬������6����U����:�+#�������m��[���GfT����:���F7��h�һ���:���F7��1�1!s���:)�Ł�Gĩ�BԚӮli[�ֻ�z,A�ų��y�pFz�I�EOױ���z�F�W
sx�I)| (@��F��6�:�ۦ���ު�W�{Fzdz�5�:�s��:7��1��1#s���:+�:�}nz�zvz�[�B?�(�E��ص��RM�Ɖ '6�:�@©�r��:kY�:��)1�x^z��F�����@ĺ��F�����|^z��Vz�r��:�����Y�e1��b��:1�d���:1�ds��:1���{3=�����p�fx>z��F����
�:��Õ��&6����T����:��(E�ϻ���:���F��ő�G��/��읧����1"�F�����|Fz�z&z��&��=S�{>zdz�5�:�q�u((B� (EO?�>�=fxVz��FV.�:��((/�����U����Vz�r��:�������~6�eXP1�m��G��:*�ř�x&z��a�{vz�z�C�:�q�u�&B��&G�{���T���c@3�˻`6���1U�3�����:���F��éՄz���&i�ӻ���:���F7����6�:����������gL&�ۥ�̣{q�� (1s��:�ŉ�G�1s��:�ő�Gđ�>�ԃ�F�����|Nz�zVz���Z�:���`\���j� (6�1)A�s
I�Aķ��F�����|vz�xNz�zڴ��:���:�}Fz��^���fm@���zVz�޻���:���F7�E�ϻ���:���F��ő�Gı�CĽ��:�q�u�&B��&V��:�� '�F㓊ðj��&6����:���&/�����Aķ��F������:�u 'B (A��F���*9��1��uA���~���buA��w!��@�]�A��� ��CN�Tv>��r ���6;G�9����� ���eV��\#��U���YN���"��a�	��K��s"��l*�#���"�����҄�G�7�������0!ix|)l��x�5yWH���U!�����y��B�R���ۥ�E�gjk��
¼��[��`�nT��:=�����Ғ�G�7D���s�Y�:�w��~r�9_8��Sa�w���[�)L�s��;���s���z�����z�R��Z�����9���I��"V��k8�M�:v���3�:p�B9GE&o��Q�(�����2?ȝ�X:@
/.d�:�v���J�U��e��Hql9<A@հF��B�s�c4�����b���#�:P"L6C��9�5����!0���0�:���ߗ����ԯ-"�X.�n��:ꧺ:p:�I���;ҙ��lqC���2t���:`t�gz����+�7;�1��y�S=<u�/��sL�$�@�$��\���<l?���60�_"���;�Q�:�Z�÷�(/>d�͊�:v�a��:tn�_Epn�Q^ԝ1�$�j�w�:��#�2�'�R�5���Y6�:"�:A����kXpI	�|��T���:�&�J��\���	�r1�I�@���;��:��F<GFF�"|��W�x�n��:�њ:�?��gb�N�l��
��'�.E�y/<9�!��"V��5+H ҟ�;$�<<�{<]�V����:^� ��ne�Z�|�:\�=4�p��WG�$V:�8���0v:J=��\�~�X:�j���DLC .\Z�:Β�z q�e1��6{??B^���S;hk�87z�C� k�K��X:�U?9ӌ�:9��6����Q+�c&Q.�"<:E��!h:%�E���oRm�a;��se��y;�8��y���1��*�_�&pI"��C;�&	��,��h:<���u�ácw2V:b�L�$�uw��(~\��wO�F�h�:�� +&2<Ra�> D.d�:��l�-�:�W����-�����| �ܵ����:uu�9'�B?��Kk6�Ժ�@a:V�#:&�o��/�6����@�N旱<9���I��"V��L]= M�n���6��:X轊!�(�H��A��:�d����:U�t�b2�(�؟#�<M�U��:g�֪x/��gLT��r1�I�@`��<��:EC�V.r��júmް�:�;� <�{T_��C - !���?�H�6 c�8<Y��̙�E[�d�㇌��"��Ɵ�:{�$��v��� �k�{�:�L<Xi�-/7<�к�@>#�[w��.<��|:|�Kk~tM;xR����E�B;����(�:�A�9ĳ>N�<��]t��A=���:E��;&�h����G})��T�
��:��k�->H;��y(*,��us�����:���IѝU��'Xt�b���u:p���0�#��D�C^Y =�;�<l�N�:I0�nc�%���
C6 ���F`8�:��i�={+<���*[�݂��DnX,.�u:P��8��8GG�Y�r�I�@���>��:Dn)���T�:�Q�L;�!���*�:�D�Iq�X�9�t2x�h^��:(Lw:QD��b���d����B��	m�q3<���IѝAU����B�� ><���:O��zAN���K6UZAq�;���@�:�� �p��FJ6N��#<�w�	͊:�!�!`j�����l�+�3�p ���'*<;�.@��F����@��r.��:���:n����:�R��]_��.�)��<�M#<|
+��ʧ����cp}#yVO9��:|�n�>&N�:�e�Hd����4��:4�!�	�U�������/dh<�w�h+ Ix�#B�-�g��\�g�:���:mjt��F�*�]� D�ig��#�o@�:t. ����9���q�R;��!�ʞ���b�:��uRA<�g�C�0<��)�r{@���:��挞��������j�ӎ����:1��b!��:�\�|��y�>���:��H=�z�@�:�q��u 'B�(i�ӻ���:���F��ű�Gĉ�A�݈H�"X�{��<���V��:��(�H<ezG}>D?� (G�ݻ���:���F7����6�:�۾��Y���p_�G8��:0��_�G�wG����co ����q�d���B��VNT�_)�gO%�
�:P�Z��:��rNtG��� ���3�%���;���s��ąɗ�)�ZP���	G9)ٲ1�[Ҙ�:1�WZ�(&��;R�e�A��5��9��7�������_¦�q����Z����F���pv���|4�;�Q�����ϝ����{3�A"V�K�ȡ4>�%<��ѻ��"�{���A�9�6􏷯�%�]��=T;���;Nt���rǃ���1�|]�K�{�:����׹��?��h�B�Ý��*��- ��n^�b:���i�2l��:�R�/��;�i�$�^d���T�A�kʭ��|��y_����F?TX���b�]�	�!7q��s0��������S������n�a:��������P��W�Ҷ���WS���T��9����)`�l|f�;������ϝ��`(Jy��z7���`Z�e+<��"��s�<{�@���Q���8�j�f����N��3�P�~�)�������%<��U� ��Y���B�M�-:�hhU� A����2���Ԝ#��c�
 j���:�������KZ���~�f���%��L�N�0<���}D �"�:k����~��:կn8��K���zT��(���R��Kd
�
f|���g�R0���ξ�I�d�4�9^�T���K�� ��w���H_�&��}#��]�<�e��rڦ��(4�g�A����F>p�+�����/���l!���i*��ĳ���$�D��G� �ZV��d���L�G�$�ZZ��Ý��������:�����*4\>i�b�6�&���5qrB�.�~�D�K8rヹ]�����K������s�����i�@��g���;�Y���^�6��\�\��Vۯ�|L�9������K	!��Xl�-5��a` ���tEN��26z�;)��X삵��@��^���l8ѭ��W�2��ǑL��q6ʁl'@
��U��\�����^����`�t��l�dƐ�ۨ��'�ʺMW�!���7m�2�]�\Nw�[S¾@�����z��.��KB�o!��ҫ:�����ݧ&�3���ț5�d���tE�A���6z�:2�l��H�i���N!�"���59�A9�p�r�ؤ��=�M�bQ�� s�!%���8���c?]�)��_`����4EMLO#36�?7��.�����C�惸-"^�������~����ĸw�7Z��R��>��*S�a���)eC�ܮ"�V��Ŵ��V���no��ѣ�=���#������[Z�q�s�,���J����(�H�����Fy�o�O6���ƞ���j^����R�)�6��q'�)6T��i�r� ����F9�,w��&T�H�Oc������㞂��j��]8�����4�$�����+��)��O �����EN���6��?0�����49ó]�T��\F���C61���b���!T9�$R��Ǟ�Z�>�+M+Pa��p�������o8m�o�(��<���U� �AdZ��$�����-��hV�߸�7�����=�J���	���6�cPޞp�����:q��:���7�����#�C�/�i��4�͈/��x���5����iE�A���6��@2����FN����7�)�:�n8���b��F���ʸ
��(��e�눩���i����P������U	�<Rk��u�gV�"�3>�*W���ʇ�r���}�J��P]�a�N���Q���3�v�PA��6�؞a����]N�����-�
��%w���Ƽ�؜�	N�
�����������׳�%��Z�|)�1��!�C�ǖ�6����V�0�X���F���>e���׸�"��������EN���6\�:0�����B(�����}����gu�ɻkyNʞc�.������6�8t���h��j�c��g��X�]g�����i	u]R���[�V��স2I]�Cքh��{��Nxz6��7��U�F�^�������3�x������|,;;6b@ <���t�+�_�6�u�5��������la�����%#3w���6+��n�1���
��KV���6��*(���%��ݦ��6&��ݽ��6&������%TW�#���[��6��*&����M��KKO�6��3k���6(���#���%!3u���6A�6��Q"����E��("��Ŏ�)��p4w���ŎP�Ŏ�A�E �1h�5ZE��_p����deiYz4m^�w7?;%�l�f�x�k*A������H�eN
�K�(�j2����]��]�+�?��j63��6����W<�Ŏ �6h�5Z�M��l�(T��6�7���;t߲]��j6�?�9��S]��K��6��K�Mt
�o@-��l
��uW
F���4EMLO#6z�=+��	V�T6c�f\@��f�_���(쬂���V�n���5k�~ǐ�2s�ֱ��� �����'���d���&�������l�z�F�ָ���*�h3_bN�$�Ҧ���)�
����-E���;�<؉�;�糉��U��6�±eTE�<�X��4���)�?�F�-?T�6���,+�����Ց���ːMjY��:��7���7%\>	��36[W��q�؛��71������2ê�>�4�d�ѝ�es\i�g���6���=�N��ꂸ&}���U$�6��CО�K����(������1NQ�ً�u��+������2�v�6���o����3��fܞ�̓�c�W��#K4�+�����ޱq/�$6���� 8��{��Êj��p6��(E����w��׿�b��p�F����d�3� �AdZ��$�����Η�b$��6��U��V�r���ҸJ�L���ೕ���w�U(6��H�ٌ����6�ϸ�4EMLO#K6z�?3�����&����Ɯ��c��i�7�h�I��Z�t�7�������&�
�������6���O����E��{�xM�ߍ�ӡ��wU��w-��'^�����2��Y򂭟�Ѷ����.�Rn�����D�զx�g��Ӟb�$ҕA��z�\���"�Ȟi�˞q������ʐ����.S���)��7�"P��H%���)/�N9�R�6� ���%�5����H��	��8L��S����l�Q-`��u�aٞ����X����Sզ���	��a��`�6�ғ�͹���X�ك��|8��E�)��zS�����RZ̞�K<m�����^J�v�6��(���|��4�c��mb)T/`"6��-4�c�-%1ē��6����Ⱥ���H�7�x��Ĵ����e���Ɗ�����%8�56�
|�'N��gd������)��+�s붟 A$X(W&�����?\��n�U6��4]��ֲ�&����Ĝ�	�6(�P_�@����9�l����|�������*�R������� �|��n����-��G�TP|���)eCt�7Yч�޸?:�tڞ��/k��F�ۈ�l�����\�p�-��Kܞn�,OKP!���7""n�������2m8����5�������ƻO�
����f�� |�46���~�����Q����C��>t�]J��Xi�����0�lG��w��(%��'��)��au�F�6��x��M�Œ�T ��
v"�AЃuv���=�����6�踴iE�A���6��@2��]VbD����m9�s���6��������tB_�x6Ԍf< ��^ƽ��Y���6��j��b�3��c99���f(����z�3� �AdZ��$�����6�����Q�_�f6�������5*ó]��&"c�	�;a��t6���h�����$�����N�B�ʶ#�6������	���4����/EMLO#C6��;3��M4��R���?��:��:𸔿�ݥ��L#�������h���X���O�������0?�%*��]�*v��Vcq�I`*w���4(�t����.����n�i�ǎ��E������37L�9�p6{'�3���Vb��f���L�q�u0�M5̞�|���ۆ����͜w5�ŕ}�T2�1cwƆT���,�<��V�r���Ti�j�l��}�/��QIȞ �AdZ��T�����!m�<��I���6���vub�7d�5I��@��52�_+�����N�oW v��͞O�ɒ��χ�6�$��̀�jP^����5�۫ӳ�=9�U6۸����ǃ�ݟ�C���?�c�u��a6n�����#�������h���3�ց��G�3���
'BP���D4i�]�y��d�5��Ө����5����B��k�9�����1I_=6���1)�I���W,���	ZX��26����j��#�����蜸x��2��7�}:���$�Y����t�+�_�6�u�4����Ń�Q/Ì��% 3t���6��6���k��	��KV���6��*(���%���%!3u���6)���o\��o^��1�������Vޒ��6&n���n�6��W���6&����?>	�	��+���6B���n\��o��}�*����]�Qں��ٗE��g�j�ʝ��n5�(���6�1��n5�(c=�(�E�AWv!��A��D��ZP��+��OCy�G���<�=�6�w��=��u�~ ����)0"����"����+�gE�%Ar�����:A1�L�M�0Gs6h��P�"&7�س�j6�*�6����[�K꺏3꺏�5��x�[�̴[k1"��6�+�6���r��+�d�CMOK��ђ���i��,���6�������6�bWu�l
�t
���6��_uå���`u&�O���AJ{�,�������6�bWu�l
�t
���6��_u��z#.��籹ѷ_k���n���A*��-�������6�bVud
�t
���6��^uq�Y�J�,���A*��,�	�]�MIOo�/ ��r�b�W��2�y��=���EI�d�*���<�X�ϑ=�B����T���S4������˂�^�0�co�y!g��@��^&m6���(�]6QU�b�hm,5)�8l�?L
�y��SM���܊}�x*��܊'AW�����ϟ9p0��y���k,�q�'��q4�/��/%�*}��28���B�$�%�܊�(�b�~�݋{�+�kTƿ3݉⺿��AL�׭o8��v��y���	�&�9X����4 �WeA�xd���k�'w�F?72X1�,h�܇d.�֡�8��y5^'J��*����v׊�U�f��̴��~��u'�v�'Ǖ��w\O�ܹ�^�2�٠��'N����ꞇFڊˮܝg
��%s��5�f'��j&��`Z�IZ'��W��1׊�g܏'r�+�z	�܎���*������Qԭk�&_7&��@W��V��D%��k'�Cy���&%2�ꬻ:��ܾ`m܍$Ǩ���/�='wQj���h:7!m%��dd.�=�����5^'v
$D�(�[L^3��Gp�L^���n'N�X�<�̭�6���l�$Y��t��Hԉ'ߙV���&lk�lA�a�3�z�`}�'"�'�8��ܪcI��$��G7��@, �&R�&l
p���'��,����a���7�A1�'حqz
���"���>SA��]C��%�'2A��c8��==�-���B�,m�I�'*����l���{7��܅M�ה�����'�z�,�'B����T�<w�'��u��!'r/+�	���ܞ?5�*��`
Kx܊S��k'N������Oܨ[-�j��iKδ�bW;ي'����
F%�n��I܁�}��&����Gߋ'��S��x��[4��xy���B��S'���&�*'L����o����{��~}�OL�ѭ�'@5��꽊a"1�W��@��fv��'f�
����(U֩7`���G4kw������'x Tl'���ܜ)�����L0���&	>���bf��m��vo(΋�l��&jSg'	=�%�����hE��|��v�ǭ�'���&6���G�P$��0sg�-D̒�B�@���'��j�ˌhխ�n��܁
�V9'��#�.'uЁ������ȥ'��'h@���F ��o'*ѕ��@��|4���W4#���c�ܟ'��w%7�j���-p��=D�!�f'���k�&�������M
�Ih��2�܍��E�e�^�'�򭯬����ܪ�Q�-�&�`������X'*����l���|4��ܞ+
�����&Z�&v����L�l��؝��K/םM{��Њ'�θ��z'8�9��D���<&��I'�h�E��ʭÉ��u(�O��ך \[�&I*j���`:��:0��e&�v���
�Rj.' w&7�T���h�܁���p�l���`�&
�Wg���7<�$0�VZ\�V��>'��#G�-p���(���^��y��ʞ��&.��W
��ŃR����@0Aי���U�'���T��'$k��Xܒ!UqGߵ�)@w'ӷw%Ǖ��<- ��a/S�����&Z�'�f'23'�\�5'	�K0Lט&�����&9��3�% ��L+�ڢ\�a��2�}�?�'*����l���}5���''C!gF��;'��&
��7��Fc�����6��M�������'umA�.J�$�H��܆��_'��t���&p�����n:�	"��-�ݬZ'$��s<��&<Q�O�'8̔�<9����}�5'��'�9n���J'��ʅ�܃�������tY��&�ݻ'Ǖp�\^����\o1��?1�rb'?�GA��k���������GB^��H+�'ٝ���W(,��&�&G+��܇��h'A&W�N�����ܐ�͏�&	v�~'ŽJo�)��I[�C&��a���E��'?�A=�[ӷ�������GBn�O�'�BA�ö'
k�k��i9�x��]K�&(R�&B�-�L�&��
N�wC8x#��K&�Y�'�Z��&1�`a��J�C>�BZ��hE'|.ؙ��4|�i�؆�0�\3>�o'u��:�5'�>�l?�g�A�]э�V�0�'�ʹ���2!���a/C�����&Z�'����(���2�v�$Ǥ��"z���5'�ڻ�~�i������GBn��O�'��7&��>@i�F��"�ɏ����]�}'�9-��&��˵�/;8�O���B���'?�L�9'b��s�bU�a�M�Lp�9'Ռ�;��)���w4=����܉Ӿ~'r&+�����܎3=�v�-�:�
�3܉'ҘF�4,"��������h�cv�}�'`�n;�%�o�����?����܈'�A�J$�5[�p�y��W�"�܊���+8F-��'����܊'W~kU�~�Uz�܊'-��'��S8+F�`�mrt��M?3��Wߒ{�a�i�x� _�j=�@��'U�~����l_�U���578�A�h��'�a�C_��m��'�Y�"W~k����x��p0"�'��M��p0<9p0������<����C^={���\����=Kf�'U�h��KP>���hM�mS*5�����m_'���
�0y����5��ڄp��Z1t��Qj��3�4,��������BjM;�h���Bjf=s�*ɫJ�K�=J?�a���ٛ]�K�'Gt�Iu�=ۖ�w׽�5d��]S'��+�F�����O�F���S�K=��i�K%�A�3D���B閩9ɹO�㵴B�]�gb���N!2�m(A#��E	n�p4LT�$���S}������V;8�2<u���Н��'�7;t���&���U����DGՍ\��n�_��J�靂�>���e�Y@o���x-�2n�Pnq�<����n��|��B*��=���"Ӝ����u�!Q+�靣!-�kÅr\��Å?��!�����P� <ɉ���> ���;�=0Q���#�7���"Z�V��������6:�Տ~�������*��w/�R���mk�y'j�ݛT�׫�*)v�(m��D���^��i�z�0�������IK鯔�i���zr�`�����M���ȸI����~�d��#_�a�u�Uq�4��+��I��o9��N鉟q���G���������MNh����x�ov��}��@�'0��������{7��Wo:t�'	�^����r�_F�1*����y*6���{��ԝԬ>a*�ʨW��V��Q�	�d��-���m�ȝ4��=0��rX��� w�0ҝ�4�)��ܝ�n���X鄸�y����zc�ԟ�}���g�h���k\��|2�p�����b��@p��3^_��X��\�]�j�Dn���N��Ɓw)F�[}�����p�iҮ��M�����}͠e����k\��g��a�搔U[���Q��ym$�Z��}�fj�	���ʓ����؋+�F�\���������$���#��)���+��X�8&���q�Вb��G����wh
�+�+� �#�P�ץ�������)���^�7�/X�M�� ����j����#���S���I��K�~O�;�Z��wL�?�����4� ��r�,�k�}������Ok*�	}HRH����N��%��W̚�'�$�ܹ�������ur�`���	Q�����]��_c�,�#��+�T�T�3t̖��ʆ+*v�cm>ɻ&���+�H��!�݇����C{O���/��q��U��i/`�i���k��$�zŕ�3��ă�����@���)β�����ɥ1�0�8������N��Γ:��� c&7o�_�7[��_n���v������e�������1��8���΁�5�v��)����,�78�+8�O۩<�[���J��-q�6��;������k�?�������������<1�8��ͥ����u5�Q�������w�a$58j(E6�����-��	�:�a�F�v*�������\���{����w�:����b�8������-��H�X�D���W�!�����<	I��~W��y��0s���X��Ƌ��8���{8���W��:h��|���i��8_�� ����.}1o���yQ��I������2��/�����A�wAm5Ԑ���+�!�88��x:�Мƚ��W�����8��Oo��m�.����NX���nm�2��o�2ѽ5yחd���.��X��Ap�f�i��&me�TZV��6�O̩�	�_��	O��&���6��;���[���d���c��h7!�����.��X�������S:аM����� d���o���F�8��r��/�2�@�ʾ���Qk���a8��y7��Z��Ϝ������"���M���Cޕk���x����ͮ;�"�oT��]�PH{��������`��E��6�E(��=�����F�޲����/s�U�ϑ2[�f�O���H8Q94I!z_8,"��w�tq��8ۣ�{���q��^���Z�{�2�`��w�8j��I���"1~`�?��,��,+P���_��78����fE��=���U&��1��_a��8�Of�\�V��	J��[��G�����eǚ��8�ޏ��P�.�'�V|�ѣ$���kJ����q��"�\���6i������}���~�Q�ةp�,� <��S��o�������{5QO���-�l7=��8�c*��kP��8��L����=
d3�f��Z^6�e�P�d����y���Q�N�8U��cz�U8�y�P��i4%�i�F�8��q����8X�^�� д�8^Ւ���il%B�n[�qq%��O��wNE4X�	F��8��iT%P�T���8nP�4����=�g��V�ThXϷ���8�N/4XŒ���F�8��ɡ���X,�1?��8��eX,�1�5�1����@
^��-�����*mC�/��x�dm��o/��,+yw-'�I B*��S�Oo?~�LۙAK��6���J���FG��P��8����8��q��4�1��<^��-\<�W,�;7�����Ʋ)��#������*��1f��^�N����8^�Jq��TI��7}���>罷�5�<i�ǥ&���9����p�_�Ř���-������|�1!��8e����X�07ӈ�V��&���8��~v4�%����7���w����iK��������̈́����8��з�����g��a�����������
����%/�cX�f�F(���iW�5��LR��[��+��AL��� �p��_�����=e�|��7�����5�����aoQ�s�Ǒ%����m�U���ǩ���?�}���=8��H���0ĬUJ�L"��i��.�'k�R������� ]0���J���O�V���77�c��ۚ�7I���g��7���A�6�z�8����6a��q�����d#��6��_���]8��3����:�F���`ɏ���48���f�p�Ǿ�J�bf�������A�b+�W8�w���/��_��0���Y�'����\#�7�O۩�	�_��J��niq�7��LR��[��?���h4��HǴ���<P���8Ǐr}��w5Wo���kJ��1�[6�~Fћ��O۩�	����J������8��ջ�ݎ_��*���^�+A��]�M�{{Ѧ6y|�d�x�ՀV7����S�&���Xb�!(�*�s����O��hl�G�����A��u�Ɩ�"��t�<؁��V����F��-�K*��ѩc��3�	~����8�8�p���A�Wt��T8��+���Y�!�Y� �3+��N�n_�Ѷ8����QdGE+�]����Z���O�Q�����vҨI �p6�Z��4�T�f���<|W`�Ib��v|�ʛ���4��oM�����:���&��Y8L��Y�f!/�5qH�����O۩�	�G��
J��@#������Y8��V|}�����X��xQ���G��[���-�UH���D����Q��b�Ѩ{{�����P�I�9a[�8�W�Uub�Α�H�t�wp�i�İR��F�`H4ŕ����Sg�G(~DG��"������k���i8��}3��T�����>�'5��m���@8�����F�C��&����s�4@6~c��[��;-�@�&e��]�r��>�S�h���?��������86�j��9�4�5��J?8��"���0nAf��*�i79��(ј`5�Q*��W���Ϝ5թ�4K���E/o���5�_*���ȼ����2b{b�Z�F�8"-���q��2+���[8x��1�m�͎��������S��ֆ����S��08Zуe�[�p=x���7�̺8��]����.�1$8���Б�P2c���+���������8��~@���K����U��o��,���р6��d�q� >�{���J�`���
�Kc����8����*��f��'.�b�PGx���5J�X����?̟�O5m5,����+�!�h8��{9����k��	�цG&��y� R���I�[������ �k�qn,���5(��1��_C!z_8������=�d�VK�����2���^��Sg�O̩�	���3	I��h)�7�n��O�����Hxy�`�� {���6��`ӧ�拒ћ@���Q�hTV�FF��}�kw�Eخ�{��4�������濏��ʷ��Q�����@�;��ʤ�q���$%_%�LR�����
�O����5�"��^'�Ϫx����;�Y,՚�K��0N�����^���x4~����3�ҕ���?������n��F���-6�a��������8��x4�y�6�8g�����h��&^��R\Ζ2�t���|f�Ǧ*�x�1 ��A���Qk�8��<��p&	�7�4�4DV:�W�M��Aa����?����`�J�<,��+�Q���8��S5W����-�6T�%�/dv���F4�7�E;ع����n��(�%�k�e�n)j7�e�P�d����8���^�qu���8D��-�Z�%�s4%�N&M�������P34�������8�J�TmX�Ty�^8�X�T�޸}��@F�4������[XJ�q�a\��^�U\������8�yuI��il%R�@\��^�qw���8D�ݭZ�5�W����8��`��<c�,�k@[M����*���\zeU����!������H<�1���m�1�$��T�k�J}<�iM������=91'�K��<*O�L�I�RTF�?�H8j��8�і��i%�q�%͙8�ѭ�n�0���qk�ή�1\Tg,�Q�R �M��n5���9�/��ћ1mv�8<D5[,�/��ޛ1���8Ѧ����8!�3^��4F��4+��8�3K���E����E����W?�\<�������8\L)1,���Z��1ѣ����8!�3^��4F��4,��8�3v�$�C8��Z��M�/������5���Xi^�����B�������8�р����kه�G�w���܂M�V6���� r��/���ö<�Q�%j�����O�����(�w�A1�J+��Z[7���q�f�I���Q��I��a��-��`��P-%�f�����g*� :P���I�������� z�B�uT]C��-����_= 3����i�f�-�P���R-;�Q�]e��C�xt��QXu��˖�@�Q����p��"r@/K��y���QoB�^Isi��!��7��Ah
�	�*16�U9BG�_w�|dw���L�«U��U�fw����L���Wc��d��ew�ĭ���˵'�˵kew��U��4*r�t�sSj{�y�
�e숀[w��>
�lx�!ԊH#v䔥ew��_w�|dw���L��3U��U�mw����LB�Y:H�>�vlx��&���q��e �[��UNM揤qp����t��e��f����qj��qe7�i�;����2�:��d:s�!%eE�Iߦ���6�C���],�P�``�(��й��VuB;�ۻ��U�}�5�]��ݾ7bJ�� ��^�yL6HN�ַ�}�3Q����x �!�+�##��+99�~�[���~�5D5KQ	WV��p/����M�3����������6���#+ހ��=��W�$���OF���~��K����t"����;�\�"{mMh�v�',���
�Ǭ��:���yJ�������V�5j'��<�����NF~ޒ�!�o��?�7CC��}��X'�2�LE��2+���X��~E�ǰj�R��l�E��|W�B~�wu�'�Ǥ]*m��Ǻ�/^���8�z��|�ǟk�1����$m.!��q��ަ��D�Ǿ��*�p'��L��7��z�ǐ
��5����/���97~ޫs~ x���~'�M�y��(��+����oX�<߮J~�� B��&�@|�{ޞȮ�d��u>n2&��h����c��%E~ޕ�x�?wC���n#ǧ/1����lN~ޙ��d ���{����s���~>@y~ޑx����Z�A�p65��Ђ�~��~�ہI<gz���#ǲ^���cQm���ބ���u��܄�ǰ7���li����ޢ�L��^��~�a��������R��Z�ޑe%���,�Q�k[�Ǯc������{�ݨj޺�2����8�)��Ǔ3��Q��f���~��[�3�3����)�k!
Y+��N*�#�ޠaX�L߾�a~g<ǭ6KY{�:�ބ2��ڑ�4���3GkK��Q2�J�L��M)���
!�2�X?��	6Ҩ�J-���޳��~��%�/ v���*��~��jބ���u}��ܝ�	05��7�e��~�1�����h��x8���^�/~�^ǐ��޽ʀ.�`~��K��Ǥ *aުAp^%����O�}w���~�Ǒ8U:���~޺�ހ�%ۏ��.W~�����R�XxZ��$�A�2ٸ�O|��b�0�Ǿ/�� �~�?���~޻�T�(MG��~s�ǚ%$'�T������{�Q�rw,׵��(mC���/
�Wޮ��	k����rǃwh��-�Bkǌ�
�~zǞ�L�y�u�p����8K9��6������Ψ~��'V^�&��G�X���@`LF�~�~ȸ�{�s��3�J�������س��N�~5pU���v�E�@�^�Eǜ�2��T~ي���Y��NSf�
��Ǚ�tG4'�wd�u�~�XD��*gQI�ii�����sS�<f��M�|�n���u�����6���Qs�Ml1�ޜ�)����8�����\Z&��\����Y�ֆT�ct�eZ�r���{���=;���#�ހcX���ޅ��Ǳp��ۛ��{��/����n"���WS9�'ǌs�X���G}��%���N��������K���$��~0
�b�"X�ޡ�=rz���3Y\�ǭ��~���ۄ�Xޫ��G��/�)F�ǫ�rtW��W��v}ބ�c'�P��ߖ�Ƿú���]�XHM7���sK_�ڮ��B�z�:BF���#�)�������${���3�-ǮZ��wZ�޾c~ޟƄA�]��֔=��ǐ�i�'�b��,~��R~CS���]6�#���έ@~�����}ޒg�8�]~���0=����*\�fGGO��^��)�z`d�Ԡ��Ƿ_����Y� �{ބ�c'���ߝ�ǿn�UNe�ǚ�ځ��[��A^��0��wk��8��N����e�^���
�aǩ��A-l�TP+,���*{��g�P�fǦ�-HW -)�iyބ�c'�P��ߝ��lۿ�%}�+��#���E�*n�e��J���OAs��dƖ�u�ފ��G��.BW�l��A>^���>�s�����_ޅ���ǁ/�Þ7��yI=	���g&u�Ĝ�rQ�ǿ�����e�Z~������e�c{�u�}>���Q몑�0�����z�Gߦԁ�l����ŧ�QI�_��%ۏ����'C��Ǽ�
YCޮAp^	�ބ���u5��ߐǰ�3��Zƴ��Q���V�S���[�-Ǻ�uƧe�>S~�@� �ܳ��w~p���Q
r���#��+Z��E3{�0���97��j|R��#Āe�)ޛċw�Z�.�~=b���"��L��M)���7x(���x4X���"kx�%~˶~��~���#�]�ي9jm�Ǩ�$D2��~[,#��z��#��ɪ����Ң�J���JҩO�+}�)�9Y9�-��t��J�y�z��ǎV�~����փ#�Y>#~���j�<D:2��~��Y>#~��̽�g�>ٕ h��%)�p/0"~����p/�p/�R�A��=b(�֨��3 ]Y�^KCِ��X}ţ�qE��ñ�B���k��S	�r<�g�kV@�7�.��%�/%V�.൤��ƨ����ֻG���v00�i�ެ�N���~���~���~���~�:���r�W[UhL3ǭ!{�i-s"~�rw��:�u2��٭�ң/�X�Q�"k3�D� �/�s�u2��٭�ң/�X�\�"k3��M�J3�E�,�/���ޫ�{��Ǟ�<���#��#���ǻ�<�1��2|-��c4�턨�s"��8�{��Ǟ�<���#��#���ǔ�;�z^a����Xr3�����W[�O���~ރPu�s"ڣ�~��*?�O���~ިD`U4�E���W�Ǯ�i��W�:�h��ǃ,
Ӫ#��E�n	������ޭ�{��Ǟ�<ٺ�#��#M��ǽ�;u�^�m�w����p��W�Ǎ��~��;�K�2yc�2q�~޽;����O��[�Dky3�"\p��}\�3��q��W�M\W3�HU}������W�~� >K�{���o��U��/@��w6���~�2�桾zY�z?��~�7�G�-�ٽ/�/��!�s"����p��W�XM�s"�\�wJ���HNd�Y����s��8�{��Ǟ�<���#��#M��ǔ�;#��_�|]��/�����~��;�s�2yc�2s�~��;(t@+sK�TU}���J����MI8����Q�5�}�-{�O[��~�w���X�'s"nw�O���9 ��~3oR�s��~7�����W�6���~�5�塦zY�z*��~���g��6ߡ}pr3��������/�l����<��W���~o}O3�~�������W�w6���~�2�桾zY�z3��~�7�8(��ZӼ�D���D="�/�*���~YDX �?�����Wt�~�2��J3�ED�vF
a�D�{��~ޚ�Y�����?�6��ֹxFT���kY��փ��"s"<z]�s�,%-�W[U�K3�O�T#~ެǎ��~��;��c�2yc�2x�~޺w;O��٥�	�/H�i+s"�����U���_�vq�B2��x�Y�2���ޫ�{��Ǟ�<���#��#���ǻ�<ɯ�m=s"6!��~� S{g:�3ɠ�)s"�M��3���t�WU}��,�E�W*I~�/�~��'�2����D����~�����S"�U�b�@@�%��1�z҃�Q's"�U�(�/!"~���
%�BQ��š��?�{��Ǟ�<ي�#��#���Ǘ�;<e�DdCTIz�����/-~���e��G�@��E`������WM<h3I~�/�~��'�<����D����~�����OT�~ރPi�s"n�Ǎ��~��;�K�2yc�2s�~޽;��.C��B��"�~��g)��մ[ލr��ׅ-~���%]�W����(s"OX�~ރP�6s"{��*�&��~�P��s"�YO�~������Wo����gO��~ރ���s"�D�p/�*�J��~�q6���~�<�࡮zY�z*��~����?���m�J[O2Ņ�P"l��C6)��~z�;"��Z����%�9�Kw�X�����1�2�s�ރP��s"ӭ�p/���w�T���ӽ��/��|�"ӽaǣ/�bV�M̠3F�ɰ}6s"/�f���Ǎ��~��;�K�2yc�2|�~޽;R�V�k�OY��~ި����.o�#���ǰީ�{��Ǟ�<ٚ�#��#������<u�ך����~����D	W�6���~�@�ܡ�zY�z=��~쭆."7~�����8��|��\=b��Y���L��;N2����MDr3���~��;i&����?�@��i��+٭�ǣ/��H�"6,��~B/��]��=��W�bV�q6���~�<�࡮zY�z0��~���\ R�}:�J�����l�DWz����	s��Yڌ���~�L<��ŻN�����ډ��W��C	���~8�3��L		m�Ft+=�N~X�,��
�e`	m�����P�U��j�4xrL�2�K��t�
����������m��
m��Q-����ɰ�m���Q� ��ϛ:̾��
���	5�� �D�\��U�������e�	m�8K��g�0ꉶ	m� J�g�ޚq��.���,tm�9�3>l�	���A���r�	���V ZD�X �-m\	m�~\r���T
���	P��tm|d���P�Ltm]�L	m�#�,�|����ͩ��	m�2O,)��-�~.�[Htm�������	ٿ3�T���
���x���\�+�����?�ݡ���
���x���\�+��N�A75w���e�	m�,K��G�0�c	m�4Kx\R��T]�L	m�#A,�|ͩ��ͩ��	m�CF,�φ�k	mO�	m��������~8T��׫f��	m��L	m�8�b����\�<�mL������bn�	�����n����c�����2��1��	m�1�H���n���;�aZWlS��P)���,�	�kS&��o#��0��dF3�[��E�	Ǥ:8kd�b����B����pz,��4ە^2Ӗm�?qg����2O	�����enh������%3|����a	s�,ȕA=��m�W�'	#>�=�FY�4�r�����m��S8�$�J��	�l�*��y�S���D;�&Ӱޔ��>�G�z`IЂ)w���}	Ü�cfk�	הAl����}�"�1	8�t�_cp?��	t8[kK�������؛��Yȸ�P%	zy�Y����D��(S��+F#�
�O�	��%/n��{���ڢ�f��"j�)�	vtiSk����sB&���P)���,���	��c�n5C�������18�mn7��  �	�W�g��m�M�L�E������	Cn�	��vO���l���P��	�C)��	����l�c�Ҕ��F�P�m�L���ڨ��	�"
�j��/`�)R�>�ej�s&	��)zzi,	�t�*�n�н �		�۶����=$��m�d��>���iG$�n	�e��D��!ie�8c�K�"Sb�+�nX	��gr�+q	&�"��7�B�	��	��;+�:����j����
]�p	�	��.~��sf��ڴ�N,�ٿ�H���mU|	��#VDt|km�7: ��=�����;bO	�b���*��oƨ���=nNrNz���	ͤ��k�����V��(�������A�	vh�Ë �������� ����>n��	>#fK�%cm� rk�P���6n�b��	��-ϴ������}��<y���.m�	l�J�� ,m �Rn���P��	�C,��	��cm?S�9��������]�	in|	�|c?�J�
��̤i�Hm�����	���_l�I�>GB���P)��)��	���)m�n��#�8�6^���B(�	���
x�%~��Om�4�,÷'�!�k��	��+_��
Yl���@Cb"���N�	Կx(�JO��Bm�2@�gk��m�x	�.�O��w�6���̶��v	K�	�9�j�Y/�<��&Q���mi���	o��-�	F��2��}.ȫ�)]24�	�n3	+��zi�"�M��	#��Ƃ�	��B�m���0ڬ�[סc�9��J�	߷,��;�$Bm��nb&��i��	ަM)7:�_�Bݔ6���:�����	�J�RU�-`mQ:�����n�=u���	������ө��l���×�^�	��C0]�+n��ϔ�8h�O�e^.'�q	�B��K�mn��M63xq��m�m��	�.PT���؈����Y�DOn=�)F��%��R>m�9����k>���d�m�w	yN����N̄B�m�!��]�p	� 	�G�9:.�����m��7P)���J��
	��3� �o	ٔ!�g�	_ �m(�	��x
��3߃tQ�m� s�U3���m�	��6H��	rćt��]r�I��	��(	�C���
����m��7P)��V5�	�!EJ-B)	k �Ք�a]�	��%��l�	s�5m��?/�_�>���HNbg��l�	r��ݕ�	���2����~�	���j�	��9m�S�j��o"����>����b'q%	����%Ik�QM�I :��ĵ�m#l	���vfM�=��	� 's�5R$�\	�		k�Dȕ"�]��bm�P.��ER$�\\�	��R��+�	�p�w��7P)��V5��	�h�_��DR��n�2~�~�#\�9�	���l��9�W
?�:����Я	��	�9aY�r����:�d2|����1�s	����Sn�+w�GB����.A�+�$	�<ԋn�Cʉ��v��Eֺcĕ8�T�	y�;�m�}k	k�y�-. :��l��Su��e��X��߆B� i��)�(l9	�y�t�DQ|m�	n��5���U�	m����:��h	`�w�H��	�O�7���[吣0@�H����	m�5��1��G���ޅc�&��GJ�W��	�*�7�y� �j�m��J�	m�'�O&.P�`囷��%�qU�m�m�ֺ�qU�m�=�m�P���9��
J���V�4���g����U<5%M�NN��%bS�X3�{��O�m�]���	m�D�Kf=�m�7/��
J�~\����	m�1�}��4�2��]P���tmd3d�|��\	m�|��-/ꩰK���g��xJ�����\�LuEݔ�	<��
m�����U�"0u5D�s!��䔹vm�9�1n{�P=<���b�������
m�%-rR;�iqp���ߴ4��mNUIm����E�����8��P��lCK���{m�l����NF���_�mT
IW�m~-&BB�>&k'�K6��rf�m�����P.$:-k� 7~PV�m�	m�7�K��)�_;�/����Wm���a
tm�D���55�i����S��
-ӑ	�<��m�9Y5��Y��I���u�ʲ�
/.�m��l�ڪ�l����n}���.	��m���� �nOD�G��)�sU��	�{��m���s݂~^�n���ꂵ��:���m�9$�]v�lo�;~P"���	m��#�T����K9EK�NP<�#=�	m��9��:�R���Qfj��	l��*mcyU�r��j�k��+����Y�	l��2m�wus�%�a�7��d�	S�V�6�m�D�#K��D�j�,�E�{hl�o2m�Z���qkx��_�����
��B�mFmc+O�qI�_3k+��l��#U�J�6	m�D�#K��O�fn�Җ{(�	m��Dn���!�%�
����y	�z]m�vz	TK	m���G�&�
��ǵm&Iqm�Ǫ[({n[����f�7�]�l�|{m�oz$k�Bn`÷'��d�,m�͡tK��mj��}�\�m+0��͜��I�����m�@k�ڟx,3���`ѳ���an�m�0(}�
	��3���D�|;m�(��
pm������)�2�Nq�m
�4��m�hm\�����<��4f�F1�Ҫ�7�^fmd�%��s��mb�3����B|� m���Ju%�Rw��4��!���	j�@m�9G5�yٺ�9���`^��Δ{	��:�m�ɍ۰�-rJ UЯ0�
��l�m$�tmi� ��Pk�:?��4bC.�-�I���m�����	�0Y+�x��?-�S]?�	m�wvsn8�#���Gu�m	T�m�tmd�9n��K֕��u@�vCE�{��rZm�D�#K��D�i�o�k��mt�m�?��	����n���NP��_�	m�)���-��)u�d������<m�
���ƺm؜,ܺ���~+=w|	j�@mb7�+�y)[��+�E=�Ul�
m�wO�r�_�k�E�xSJ/����$�
m�n��(��O�k�`�l�ma��nI�m��![�/�m�%���Go�P�"9ݔ3m�9t1����@=9/�Hq�*ckF�qm�㪐	�K��N�	믚�M��	��w�m�/	C� ��{hܐ�\o0�-S���\~m��Dn���xc#����l}���C֢����m�V�Q
m���g�T��m��8+KwmirDl��x�S����󾢺��]6arml�.m�8�.d/�m#�_|4n��#���PKmm���x�Pu�͍�@�)��&�m��	0DS��Ϭ	�/��SeV�v�m��D�#K�ƶڑ@l���\�
r+�$�m��4��m$<������5 ��nJm��Dl��N���Ē��ۮ �ɰ��m�
����\Ĝ��G�%m��	h�Nm�i���+�s�����{4���_m��ymP���l#���P8�TMY.m���Q��u���8�<�m�Xv<	m��D�#K���b�\���IAhLm:�1�xy�MM�7�tmx�sW��mٛ�_)d����p��R�d�H9�#�mŭ��a/�l�Tnc��{;���r�	�8��ml�k�ڸ��#�ǔ��NP��^��	m�^�?[|'�v:��L�n�~�Y��<m��aVyA:�>I��a�;X�eS� ��ym��y/�S��4Hu����y_�0�R�m����b�ƶڔ�n-�:�{�'��m�yBm�G&�����S	Z-3`	����m��#�	nc<�	A��J������}m�y2�h5lco���K��B�I�@(%dm��&6*�]�{��+6���$:N�m��9't(�mV�|���vCʉ�G�rm8��&?ü���Pm��5�Ҫm�	��Ym�h�N�m��f�r��"�h�m��`�	m��������,�	m�m��q�7���5`�����F �ս|9`�I�	m���m�|����3���Ծ.��ޅ���WG�l-��:�I�	m����f�P\sz��E�r�<�mam�dI�f�<�mHģm�P���/��
J��>�&)m�N�	*�7LPOw���ɤy��K).�Y��WgTd�^������J�
|Ik����KWS�=�?�
�?�U%2�\���hA�V1م�>�ƺ"���d�onU3����Oqm�]���	m�D�K~6�m�e��
J�~\����	m�1�}��4�2��]P���tmd3d�|��\	m�|��-/ꩰK���g��xJ���������~+=w�	j�Mm���A�3.	[�������+mtTm����C�^��A7�k�&Mm��΢x6mԔY�(v��چ�̯��*�Ym nPm��y��%^�=����P����	mgu)$`k"�9�������`��mi|Rl�n�s?���\4�Rm�H"���Hm	`ek>Nv�k��}�����m���-�m<��dnp���)��8m��?�S��B�mm�x�KP����	m�Dn�xJ#U!��_<��kc8۔m���fIَApN��o�*On�m������}�?4�\m�n���m�$Dm�ښ�"�U���@�m	|�lQI�m���0lmX$|t�K��Ҫgf�2�Smƿ�}�#���=A���	�t{qm&��m��xk��*�����qv�Bn��r�
m�D�#K��O�j�v�NP�6]B	m����~�U���]q����P�rv�hm�S�nr���	�����~+=w|	j�Mm����mZmm��4���	�t{qm&�m��i�xk�y�no�n!�]�#����	m�FAk��@��{c���#����&:pmy2<ڌjkF�l�䃳����H&s6[m��R��:����	��`ٌ��m�32��P;+�{Ț�3�	�8�m�&�C�B�mn��;�?P�u]�a	m���@?��5t#���~+=w�	j�@	m�9E5�wY#�)�+����Rm��I?�6m�$@m�����3����,����ؽpmk���tRVmV�<����{h"е|�Hm���h�k~�ޥ��E�up��	��m��B%�ynN����M��#�NX�F�m�D�#K��Dԑ�i;~P�"���	m�ފl����$%Cm�����	���m`�m��Ĳ��P`�}Pk�S�j-6�	k��ml���&m��O8��4h�!Ս̲��m��Dm��x�S���FdmRm�(�ė8m��lmڐ�4ݔ�X�%��v���	mʣxѐ!��T�
����~+=w�	j�Mm�x|+mؤ�������	wt{qm&�m(�](�	����֯��xQ\mt�Tmn�h��l����l��2m�יP+��m���m����
^�4��!���	M�Nm����#�R��]A����P��	�	md�Dn��҈��%���l�	M�~�.�mZ���?c��H?�n���B��j��m�� ��
�mk�0���D*�i2���m����]7k���U����xd�m ��m���)���O8��W)Jz���liY�m�/���mHX�'5늬���O2�m����T�m�@����͆	x�MrZ�.�m����b�ƶՔ����Bd�m`�mе�9��k�W�s�����\m�(턇�hm�E{9聩˗���J�Imu��}#m���jq�=~V�[�r�
s$ �m�x�mc|k=�V�2��������ee�#F�mas�1V��"	�X�Ñ����	͔.3m�c���8Rm�u��Q%������vmms�mj�<���	�o�g��!��}	a�Kmb@k���5�{O��PJ/+��}�Fm��Dn�ھ(�� V��C��)�:��n#m�m�H��msR�!��ٗ����Ӽ*�F�m��3mP���8�w��g��!���	,�Mm�/[���?�	���l-}�3�
"���m��@m��xc3���ތm�M���J\�\~m�?dl�m�����/�l�����JGm��	��Q{�0F���PkbT��Vm���n�82.� �m#�! � W��u�= m�Λ�����{�m5�lԈm��<k6m�	�v{Q�_T�Fͯ���/�mFTmk�k�J2t<�G�%m��	h�Km�9[1���=���\m���<K�vm��{l�x�N�Q�mcKY�70Qa�kI�?m���Q�rQ�A���;T�p�<��:�meS����P��=-7�i��P6�%=�	m���Q��=�)���\�u_y�g"ym�v�i�����m�����4PM+��m�����Q�	�2u��(g>�F�6�m8��";���	m��q�J��	�I�q�7���[�����[Rt�����j���B;@���	m�����4Q^������P���	��l�ݩ�M�����m�0��V �����0u)l	�=��0u�LP�������M8�ᬰ tg������N�ab�r@Q�++����{HH�~�Rn-�͗fu�iת�H�}wK�m,��������ա�S�iL�I�N�N15l	�w�e�	m��4�O��������tm�m��ǌӗuf��kI���|z���I�A�[nn�	�g_ɰ�չ����Q��e��
J|Qk��bd��Q��s���H������m��@?�Xh�X�����c�����mɜDk��=(��{S�ٱ�	*t�$mFmPm��f�ܑM�U��x�q�3��g�(�	mզ,�Ƣml��s��Vm�J�tm܃Ĳ��P���~h�n7~P�m�%	m��n��(t?ϔ���2mVH ̗Pm���ԹfmV (�z\���O���pm���ʲ�{�H(p�&�$�$�f?wm�k9rn�I��3k�� �]G��Ҥ�wVm��3]{	g0�������D�kmL�Tm�Y�{��kʁo�h$��ma��ni	m������	�h�j�'��̗��m�Dn���ˣ�)��S�ڍ6v	�8��m��IP�:g2^\��nu���󷷔�m��	�JQ���	�ױ"�	��{�m&x�mc���a l���]���Emn�f�w6m����	���;F���Pi�@}C
	m���`��b���]�MP�
�	M�j�n�m�D�#K��Dԑ���Pib�mAm��_<��
��=I����
�ĸ�m,tm����ҍm�
���ڜ8���n9�z4�
m����Z��D�h�*�|Hm��/��+m�S�M�M�	�p����Ҫ��So�M�m�Y�u�^

��o�s	��/:mL�m�	�wRm/�<����w�	p�ymLym�'&1m�pP��C����	
��|Om� nڙ�'Cʉ��n�F曹�>�n�m�� l=���%�U��F��m`�����6m�s?���P�`�~4�Me�'�-�<���m���m����@��Qi=D{	��J�m�9�5��ٺ�9��h� �m!\ym)��m��)8ۺ�\�mS�DD춲��A�hm�ɍ]��-r*	'Xa���P�(G\I�m&�'�in�����]���sI�]qmcߊ��a�m�� ��Y~�ճ�'!���	m_�� Ns�;��$����G40���'mg�x�|%k�`8c���8�7��I�x<�
mV�sd����=Dn�4��!���	j�Nm��lY��r���X��A��	m޳mzBq��������ͨ��	M�Z�n�mZ���'c�>�6?�FS��MD�	n8/Nm��`.�m0t�Nk��eFӒ�q�m�cAK��	A(;�+ѧ�.��:Ӵzmmv�k�?�D��m��6nh&#(T)P�(m��C8�F�n~4�~y܅����
ڸ��m��<m����
��G�%m��	h�@m`�rx$����#�]�҂�	S�<m��%�(G��	p����PA��MY.m�vI�Aݲ�		F���i�c�#.�m����S	��O&�N&g�Px�=(7m�$�m�ڏ�!��@D��m�����-m�#�[��n�����	=�J�"۝�Tmm�9pOoMr
	̝Js�#W�j��pm�s��(�ƶڗ�k�:�i�-�m�y�q�>F������� ,m��ח�m��DnY��x�S���
nG�]�_q�m	m�É�m�'�c�t�g��!���	,�Mm�yBu��Y�	���l�� ��Rx;�m��	�5pkJW�m��'�3Rє��#:�m���Qþ��A9��nh��T���8m��<�zc���E;�BU�M�~&	k���m����<ܒ�z����NP9�9](�	m��c�	���Bm��E4	+�N�}��"m��i#fXs�l	k���Y�e�#.�m%k=�Nȧ�?��G�%m��	h�Km�}x9��n��Vy͚Tl�m����Sm���m�P���Yf��f)a�l!?mdwXK��)P�;oѦ)>�&>�%m�Zs��t�$�m��]�_k�f�唨~mX�i%�-#m���S8�{��w�4�
m8��&?ü���Pmn�5�Ҫm�	���2m�|*�Q�	m��2������a�	m���	m����\���h4�.��@���m�|����"��UQΗG���Ʌ\�޼���q�J��	�Q�q�7���4�N�m��.�	m��OE/P���BOMm	0��BO"GP�������M���x�p#Dmva~\ɤ���8����'���폦����N�|���<�4�һW��h�z��G=�Z�'��k{n���L��4۰���|�t}�Ǜ���ݢ�m�鍃��E��vm��[2�
���W�`�L�	m��U�K��)9�4�G�Pme�9��
���	ܾ-A��d50��ʄ;��2��ع���m��t�>yT6���9�fh	m�I�	�Vl$��2/Ֆ��>��=Y��鱩9����
�m�	fo	m��>�1�b�d��E� �P�
���-Eij����P�{hhE������±H��/>�8c�8j���d��/+�c���8j��8�x�8j�ھ&
���}t���8j���&F�y�i��y�8j��!�5������/�U�h������/Ā�f��8��Ι�$�4���4���8���y���8�=񄎗�^��b�F��Oo_�GD-*��O���T;�u�y¶��Q���ɖp*6�����b�ͻOaR��������r*OLYӾ���я�"���b�F�ۢ0��Sn�����nq�C��I�S4'#���z��>4P�c�{�c������a�ת�����d�z�c����H,O��5��޼c���H'�#��\�"���6c���4�Ԟ��P�.&�����MU������],�2=���$�6��O�拲�c����-1�����1�"�4����O�4Sުc����z�c����١�����ݪc�����'�3�'�˪c���ט�Z�MV���i��/�)���zr�.���%�c����ղ�c�&�c����2VH�%@�waH�ɪ4w�c�����ݪc�����'�3�'�̪c���d^�`�����c� �5�s��SeJ��I�c��ŕ�_�c���6$�6�
��X����ݪc�����'�3�'�Ϫc���պ�
��Q����@4���խ���M��MH���C�ʮ ������^���l䝜��.�z�%�c����V�M��{�c����g�M%<�$���Q^��j�o���1>�գ�ز�c�\�`��i���Z#�y�孰#?�`�����ݪc�����'�3�'�Ϫc���W�L,�������l�,��{�c���.p��wt�.�
��,1��ˈ��c�!v�^6�G�G���c�v1�T�!�J�ͱ.0����53L�@�#-,������ݪc�����'�3�'�˪c����h1�&Ҡ1��ˈ��c�v�^�G�G���cv��$��`�c����ղ�c�1�c��.�6п,�'�c��L.���e�:��uti0���M��MH���C�ʮ ������w���l�}4Z��c��:I���4��c�`��j�c���d�z�c����H!,��5��޿c���H{�8�����˼����Ӳ�c��4��P���4i�r��M��c1��ˈ��c�v�^�G�G���c�$v��2n D���ݲ�c��9۹'��fc>��z˽ԭ�`�����ݪc�����'�3�'�Ϫc����1U�c��)c����5j�����r��aZ���첵c1��ˈ��c�v�^�G�G���c�#v��{��mbMx���5*Z6k��j�Ш 슋+�.
1��ˈ��c�v�^.�G�G���cv~yօ��@�1��ˈ��c�v�^�G�G���c�v�m�/f���#�VU�[�ݲ�c�O�U�!���L�P�˾��󆷲�c�!�d�z�c����H,���5��޾c���H�YQ��W��dz�c����H
,���5��޳c����HS�r�jM�MH���C��8������]����坜�1�J�� 5jo5�.1��ˈ��c�v�^.�G�G۲�cv�Z'��ʮ�{�c����a��E�:����M�$MH���C���������_��������U,\4R��c��0e�����k�c����ز�c�{�c��;H6KޯPv��Q������c��˾rԯ{c�Ա#`���4PϪc�{�c���*ȹ�Ra���ݸ�8(����,�p�t!NC��/b���4��c�{�c���������H:�o�pE&��dz�c����H
,���5��޽c����HdC��D;��\�dz�c����H,���5��޳c���H���G�([����F�M4���U����	�J�y�����<��>��ˈ��c�v�^�G�G۲�c�vG�]�c��վ���{�
�N�MH���C�����������_�����nոؚwx=�P�ن*��N�"MH���C����������^������c������Բ�c�jh0���+��c����Ҳ�c4|`�)
�d�z�c����H,���5��޾c���H�Sk��/�08���c��m���fVmM�MH���C���0������z��������c�����J5k��[uQH5%�Pr,�L��z03C|VZ� P���I2@�M�
Y�{�c��3-�P��h�nΌA���޲�c�'�c�����˭I%�i@w'�M㞊��1W��c��.c����5%z�QZЭ�{�c��i�|�M����GP�{�c����8����j!�^�c����*���(o��Yw�Ѳ�c����_�^�4�Pl@Y�n��e1ծv��Բ�cY��8�w��۲�c����!�W��W�d8��`���Yw�P�'7�z�c��C�ϝ_�����ǃ�ͪc�B�S_}v�A2��u�[���@.��M/���gO!6�I{A"�Ѳ�c�}-�����C.8�!�ea�Ӳ�c����+�z�:�4Ň�tP�Mw�������Df[�V�K扌�_�j��'ZjP�'��`�c���F$�ز�c���zm�!+�۵I�X���4U��c�{�c��o���ޒ�*&.�z��3G���@4 :��ܲ�c�z�c����c������@48}*:H�'f����Y|�Ҳ�cl��9��5%ziPy4��v����c��RN���X$��i@.�Yw�ղ�c$�(��=4��&D�2��܁|�qk���٭�o���?��c�'%JU�c�B/���g�,%li�Y�ޅ�,L+����S[$ڶi|n @4Οn�&@���F4S�c��5c�����3�c��˼����{�c��%����<\��_%pZ���1Ly�jG,,Φ��c���zh�����4��:�˽�8��b3K�vػ�����l�gh5%@�ز�c�4*l^��U�* `u�n(6�4T��c�pX����c�J����Bұ�A���c�m7Йeڹ!?DC��*�ա���c����ht�L��Z�4Le��@��@4��Ԣ{��4P��c�%z�P\5$X�H�@.&�z�c���6�,Y�p�}
��|9D<��1c���iP�Ԣ�{�c��!��ЖEhu��j�ϓ�.��ͪc�9�OpN�-~kX6
H����/c���4Wݪc���#5l��c�x���V�ie,��1�c���Ĺ2l�5l�l���53T��Ճ���в�c�ɪc��D!]�y�5�5�����c�4i�$m��j�5x�2�2kx�����@4��(��5%��߲�c�m�Q���yNA�*�a�����WDL1���63��7�)��<](�z�c���Ru��
Rj��3l�/O�iG���ɋ��c5k�)�1�c���ę�0J����	����3�c��LJ����tv.���c���8Xtk>��"�MJ���;.ϭ�L����m��jP�4Ԡ�G�[�d.�3z?����53c���41����޲�c���@U��Q�5c���4	ݪc��j���۲�c�p�p��9x����� ,��P�Lw����}���G�5pT�X��yg���޲�c��N[�59�j�+e����^2j��ߪc��ۅv-��ѵ��V߹4D���ݲ�c���c�v���?@��Ұn{�c��C��BM�{�c�����K��O@.�53b�H3o�3W��۲�c��x�UQ{�U~��2M����4�c�����(����s���b.���-H�����LJ���hc<��k!���4ɪc��4f������c���Y�Y��6�H �^�C{�c��4F�>Z����4�����@4��*�v@��Z�˭�����Mw���l�3�;~S<��R4Jo�(�1D����4�c��'��c��LI�����`<��@.����c��(	[��%�iG8l����c�yV~�M�(��=�3�c��Ճ�{�c��U4S}���"A���.��#�]�c�����҆���c�E����%*[��v�u�Ϊc���D�vo�
z=���96�x�1c�����x���/���c��W�\%oriPy��5%��Ҳ�c����M-������'��w,�Y;���c���l((U����^��y�:4D��˦��cH�=���	WZ��,�I�#���@.5%l���i�*0���c����W��gX� d3u[�?Y�P�.�Ϊc��y�Α#���rC	��	(piZ!�&�c��˾�o��a@��P�)1�����_�c��4��f|��@.9�����c��ן)4 ���ێ4L�4��D��'�c��.	5%o�?1J���c�5���D׆5��{�c��n%W65�(�c��խj���T3o�k���Ϊc���U��p���BJ�WT>���ʏ��c�]�c��ԝz*�BC5�Q�3R��ʵ<z�c��!�b�-�|�PS]���dԭ�@4':�_�c����Բ�c�2�c��Ճ�
4,�b�Y��53h�9z�c���(��j����m
�E���h�7��I�c����Vڎ4Q��c��)I���4U��c�3t��i��ݲ�c��@�"@�%�,ht4%x�|�j��'�c�������c5j􆾥�c�je��ũS<���{�c���m)�g�ײ�cސ�d(������c�����:��Ⱄ!���3� M+����π\�	�ײ�c�J&�w�3L�/?�1W��c�K�ղ�c-���M,���X(ȭ��ЭI�j����c�QΆ�y9�ڲ�c_��l�F�ZF<��%k��{�c��7P� ;(;����%������`�iN�iz��@j������c@,0���A-�;��ĝ�5e����`���@.���c��K�����ϑKm̑���޲�c��s�\��p{�c��*����q��^�^H{��᱒5lKZ5%�i�5�@ZƊ3Cԡe�5%si�`̾��c��.�A3��)�GVˇ�z�c������|�����!�G���c��z)i&�5B�iL���Y{��c��L1���j��"���	�yw{�c��e�آz� �����c�늖�o��XBۈo�P�LJ������Q���aai���܁jiA�<�N�7����Ӳ�cW9J�����sy�݁�����Ge
@4��v��g�j�ͪc�c���L�����[x��v����2�c����aMJ����sU$Q�Ü53bt�{�c��ټ)�jC5�l�*+�Yr�7@4ъ8jFD�!��]�c������d�O4��c�˭�2j܁z�i* ���{�c���O"ZdFi
���[EzL��z�c����^��'D��Yv�G܁��53T�{�c���]�*\&peE����`̏i\�U�z�c��ׯƽ!�B�0H���4L��4WӪc�z�c���\��߲�c���=�d�^��gW�����I��Q��1S��c��40���4Zߪc�@4�w9��o���5%b�Z�5	ԃ@|�K�(I����`�#�@4�xŠ5u�B53ۤ�j��������c܁�izNK5%r4RЪc�L0���(��P)�?kv�j���#Ԅ�@.�@�L����ڲ�c:���U��e�H��3~f���i�iA�Pi����濮U�뱒Ph5�Vv�T��c�X(f�Ұ+��K�0x��`%s�����<�3�ho0��ܲ�c-�!>"?ݦ|�Ǜ�%�Vk����Ҳ�cAo�����ղ�czSvO���cM5��T_�@4�o�ā�"G����Ph��G��Z�u	j���jL?�1Qުc�@���%��޲�c��W���5�{�c��Su{%O���&_��ܲ�cp�JvȈy��-�y��<L0���WsJ�yо*|�խ�3|�@�;�odiNN}���L/���&���\::�*�P��ȏ��c53b��%p��|�c��W%��3߬12�iN�Ȅ�%@iN~ӆL�_�:�����cP�L/������З��e��M���(�m�3�B/����o˧t����.�ײ�c!��rXj��6V���4T��c�{�c���A�rpi5%��m4Q��c�{�Pú�OLw������)D������5GG��6H��ղ�c4��ў�LJ���e9��k�@49��4�t��5%k�53{ �M,�����ǳaSPĖ�
�4D�M,���`�8��N�*�iLw���>R�+�K���Q��K��iL��i[�45x�53}�T3k8q�� ���Ѳ�c��ʵ�x�wa9P��㘋����C��@�|{
˭��/J����/\q`��c��4e}035%xiP\�����������VB�z�c��y�C���V�8Z���ز�c�OB��{^n���~="`��6��.�(�c��5�R{�c������r(\ �7�>t/k%��_�c�����%܆53lHLJ�����s[53;�L1����s\�5zwy��VO�@4�֡�53b�dL0���F 6��A��MU���4ū�V��V��v���j��&�c��LJ���,��z��I?�ӝ!�h�iP�L0��������*\ �4L���5k�����c���D�%�D/b�53PцL-����j:o�|0��˭g�j��Y�4Z��c�p��ڲ�c����m�L��:P�LV����=�b�(�S�|L`po���Y�i���3x5-5%z4Q�c�3PpY����#4��?xI�"H���4L��乃�ɖ��c�@4�^�D���e5�6�{��)H���iPqʰ�3G
p��@.	���c� ��Ў7�=��iL�4L���(��ղ�c\l���B4����S H6KޯPv���2�㜓Ҡ�'�c����O@4%i�4��( �P���m�Φ��c2�gm�'a��bw�6T�z�c���Do����ßǮ1~yu" @�b~���e�L.���h��I�.��2l� ���c��ە�R+�4|�4]��c�z�c����:@kn�n��X9_є�j����@4��*럲(e����l%c�?�N�.��z�c���R7����7�u����o/���N��M!��n@�⩉�>��Vql7�F�������.�ྲྀ�&IBwD���G<x�.���.��^[v#��~�P�U"�k��.xY'-m��F*�^P��d��.��w�%�F�j��.iY^ְ�����z�
�0���3*��f���]�1����*�a_����;�q�ˑ�y�.�W�m<1���	/�8��.�y��:{!���.���.�����h��<`�]n�ԅS�P������g��j�<&Y�b�vKޟum#�G�����������O#�	�Ƶ5`�t��{�9M�5ɖ'~y��RijOP��.��T��^���6m+�K�&{�&)\��G!��.��1���Wa��b�/n��p쫜��.ݳ�.���G��V/���W�	1����~�1B���J?"��3��4l��AZ`�m+�N�&�9���oՙ/��N�������i��.md1�డބَ��.S�t������c[��2e\�L�l1���F8Z�����.��Z�zp�%Q�kꐎ`&�`���Z`���.�A�)I&�����y����1��J�)�l"�I1�?�;p{�G�e��.P���S< ���/��G��.��3���skZ��s�촃��.�y����.��E��8���0oޯ֚�����.�����61 ��.���.��~�s������݁{�/�1��X�F�EƑ�,� ���D
�b-���P�'hl�yŪ�?�P��f��.m11��{$}^֌��.qt��}>�m(ڰ��-��Ge��.��!�;�L�m�w�`���.��y���x`6h���>��f�vy����hh�y�i/>�K���N�y�ذ�{�&>d�._���.��Z��켜��.ڳ�1������b4�졁��.�?�O�/h��y�<�p��Z�W�m+�F��.�	�@bi��7�Wܢ?�O�4���P��Q!��.��춲��.��.��/�?�!�� y���4��f��.��.�6�sZv�+������Fm#�h��1���'�W���I~4+�Һ�m8�.��PO��.�*6��(H�êU�~��-���P��nyۆ��.���V����H���.�����T�r�n�q=�y~칁��.U�K{ً�f��u[�� �U��$ҕ�� ��՜�Oʔm�0�#K�+i�M,��Օ�Y|U�ձ�}�l�#U�9
�ް�e����	�FvD�������:����CX|�t+��!$���V��>�g�u�W-�������S�����)c��Ղk����M!���Ά�P��Q2���Ӌ�?8]�m��A:�)��/ ��{>el����򖑉�Gb����JQ�vEH5���F2��%�%]M#���fعe�Ӱ����蘴y)HM��R�ѿ�M/���HX��՞�������[�|v2,/t(��d�"�F�L�$ڛt����>���2�9�b�SB�Q
]t����,��IQC����C�~������e�_T��#d�	IT��v>C�A�J*!���Kl��/�H�����N*���"
�p#۪���YL�q#k�ȼ�y����u��,n�q)�z�������-ߢ<̋���n`�b�$�
����戔�6����~`$.K%��_���1@�t/��(��<R��Hx�#SԷw�M'����VK�γS�Q�e�zIz#kCZ�$ҭ�U�0�$����mpUV��>J��J�{(z{�����_)�����s­G�M(���V�ĀHlf���I����#Pc��N&������吡V2�r����w;nY;j��N��s����+ɘ>��-m�q�9Mg�V
��jqdEd�}�k�^�܅�qW�xt)���Ñ�B��]@Ы�M$���\��[$>FW�񻭵�V�^��|*ie��R����ښ�M,����^�e�7�m��Qhʂ�����|>E����EV7v����@��sF|��V鴅m$>CSH#x-�)�$�bs�������0a��ۘd9�߁v]����ܝ|��'V���*a����U
���Φ�t.���˚ًWY�ަ���)������?�ͱ�/�T�;�ދ��E��%�$ڝ�P%���*&�����L�}'.*Y���������O�*qYM%���<�`Љ�N��t����;M�i�%���n�.5���v�����G�dS�)�j t����J����S/��Ax|��r���#bMG�J|���ӣ�t���CMɻ�M ��եWZN7 D!`��M/���5�*���5v;�#�������s�U�1a�P#STJO�N/������K4�E&�F���}��B���*'�1}奆eT�GT{���1}���$�ݙi�[Ш�,�8�5}����vjȃ�1}�\zq�����h k:|Y�&�%���X3�X�@�U���^@��1}���O��G|q0�_@�a�#�x1}�V��/���r�����S�'͖1|�1�BXIed|"���W�T�x aX�z�p�������r�U�1}9z���ځ9��$j?�n'��6�X���;}� ~	~;��/��1}���]oIQ	�%��1W	ǆs��R3�ÌrV�1}�pDE�5-� F�Y�G�y1}�4������!곎�N��ÉU��%���c\���Q���_�j�\�HK�����)}�b.�@��1}��1}�vVJ��[^�ؔ ��g8�Y�_ԗ�l�� �1|Q���6�C|1}�Y�*^�|!1}��7}����_4��)�����ރ�1}��;�;m���M���8}�#Lx���k�u��;�S�O�(��r��̩ �-Y�@�E�CZ��� �| 1}��6}�>4ͯ�%�z�1uɧY����Y7�/{�1Ep_)کIP�j�>���_@��1}��@}�|���1	��0_z�M\@��1} 
��ꎼ�1V�1}��đ�~�������1�V�1}��{Diņ�Ғ�M����1}��\�1�|���#`{�1+3|?����g����%�@��1}X?��-��vZ��r��ǩ,@��1}�5-�5\� �%�z�1��BH
����ԧ)N(�|Q�@��1}�����Ś���1D��'X0�uэ��4���I)�� �m ��c0@�Zz����`_@��Ȓ�S�G� �� ��'�a�Hj�?}��3���ޤ��1}���N܏^���~�1f����1��ޖY�G����z�Pԩ2}�����=}�(�dye_����s1�V�1}��~4a+���Z��1}��$�Ǟ�Yc���2R�#|&�1}�,@��1}�j��(E���w���o�ծ�Y�<��6}�ܕ�����7@��1}X�l��:}�?6`a����R�OΓ1���q��҈@�p��(�v|)z1}�Y�L��1}�M��^��7��3}��>�G}��1�B������m��3":$�Y엳���1�R]U�1}\+-&>��=�x�ݖŃ�1}����ҨM�o6��Y�m�X���f���\�V�1}��������7v��ɳ���D}�q����8�l�l�%L?,�TV�1}�&�B�s�mR�f-��Y�e�2}��b%��P��T2��1}�wҝ���ei��2�kT�Sq�f��1}�S��c�'�쯴V�1}t���|2��uf'-$�t�Y�̭E	+V�1}���HR3p���=}��e����*�&w	v�1��{O@Q$0���w�U�V�1}υ2��ΆY~Gt%�\k+�B}���-����k����e��V�1}��h��ʫ�Qp>Ð'�#�%Ղ�D�_<����1�a���A��`Ƒ���<}��4���buP|_>��P��1�����8Y�_یV�1}Q���Bn?����$����vf�o1}�("2�1��ީ�!f��Y�S��1}����#Nh��SJ�&�g���"�R��݃�1}�w��-�qФ>�1�N�©	7�v�H�!Y�' ����z�^��20|��1}�+]Vj8�6�X�C��@}�`��_�p� W�-�M�4����� ��2��D�V�1})-�$���Eds����`=[�|Y�&U�1}���U�u�Im��%�; ����w�1ݩ
���	���V��XN@��1} �ă�1}��|h~����_�Ȗ\�|}1}�����ނy1}����`Ր�X�Bȩ�͂m1}��ܠ���"5����?�/�����7���cT��E}��S�,	դ���3m�Ʒ���J�1$���ڛ���#Z��۳Y�m�T��9b�{�k1}�rB��g�{�7��1^�D���OY�曎��1�%��i�l1}�Ứ�) ,RP(����q@��1} N{�1��֪�̾��vvև_�1�(k')�����ͩ�3}��������Uf��A}��vX����^��'�x�1�3!�� 4mz�Ȓ�cӗ���N ������Y�ACӒV�1}!C7���еx~PP���8%fX:K��A}��<D��Ά�ۜ�R�e��Y��_���.�K��G�C
/��1}��_i�8�ku�S��Aw%��PY�G= �"[�Y�F#�SU��Ь_�|(1}�4�1����ɮ�wQ<��R��i�\@��1}�D}�|�1޳=Y��<�Ee��g��oC������1}����ۯC`��k��1M�1֍<zJ l｣!��
0�FwAϩ.�Y��V�1}c��#����Sm���4}�@���:}� ��AU��S��^�Uh����=}�f��G����1@��1}��1}�|�&6̴�%�����@��1}%ձs��8}�/��ScpXY�T2����st��V�1}��/.5<U�����|Qāf�,x�1fJT�s���?�(��x����̽cI�[��=}�K�����z`�t��&�o%���}`�X�\���Y�q.y�M5���Y�M��$�*����G}��1�=���E��f�ʅm���d��<_D�+6c� +�9���Q���6��˲�2A���=ܩ�-'�-%� �����=�Z��Hs=}��g����~� p�����l������=�;����x��2-ґt�z�=���I�]������1;*C�B���U�q�a�率���m�����H�w1@����_*
<-��=��2��V�����=���=��20�s��
�=���?x�-a��ʤ�����=���:�����\�����HU�e�w5@����+/k:W$�e̙�|�/:'%+4�7������q����=��k�lZ�Q��' +�+U2LӮ����}�=��Ї$�=`0<_-���=�P��H�=�|)w1?����wh���=���6���nA�X-c��<+��=���}���s'����ߞ@2�:�o�@*�B���N�~�*N<+O�rcGϲ�vZ�<_3;1�nh��ծX�K=j5�n�<"~�=�������=��q<'��=��<���=�s�^��0�8.��F���c�����=���=��#(��g��4��PL�c^!OsA�i<-��=�w=@����+L�â��=�立e�=��S�����ʄ�X��ywh ��y�`!��+4<�w2C����i�n	�wh!&���O�����R�"k`Q� �:it��=��?J�c�ww%X=�����8�����HY[8��:����r� ></��=��pOt��m���2���=h���j�6^��|6���=����u֚D���:�`�l�/�:���t�I��"꩝~k_���=��<�����s&��Q��� /=�X�ѣX�O���=��?��eZ��xx�������=+V�����= &��!n{ֹh�2k__/���������=�G{4�������>���1�^�o����m</ %�)��p�! e���P����Y��߰D���=�B�a�n�6���z<A�� �X���P���="jZR޷�6f�)g�<_Np�����n��K�Й9���{�Z�һz}=�k< ��=�����=ѸL��-�|~ �'���=��!���c;J��N��Q����w3=�����}�=�yĵ�E��%z�y�f� ������=+,�!L� ��+!�<W'< ��=��< +O<%���=�c������kY�Z������� �p�w� ��)[�h����!��*<�;����!([&�g�`|sϚO�����6��y�c�g4*��7��i���<_=<�|�=�$��וk*w<W6<�*O��x�=��K�!~���mv"���͌��A�����=��m��_�<_;b��ԙM���&c.�c���
u1���Z����wpZo`>��=�����+wl�'lŨy6������b�����=D�'QI��<&����=�xܴ��<��w����=����_.������=����������=!O�k�o`���=��p(=o�<+��=���7�����)�&��M��1��2��T �=���T������+{	���=�%GT��<'x�=�����=���=��맳�M��r���=��=�"{�P���@�����h�Yٔ��^�����i�����=����b�F����=4��G6<8X8�|��/oRV����=�o��߀˧e��t���1�wh���=��k��q�[E�]��}�/��6�C����F��b*f�rb%�lKж#��/fU*1?���G[���=�ȝ1��
0�u�צ#�E���=�J1N0tp��y�=�O����[�1Ǒ���i�n�2X|�����2�j)D F�+D�:����X���E<6�!������u��~�=���V�lz��2 �:�����!�� /�/���������X�&+E�Ϫ<_F���<���=������A7>J�oҍ�<WV��L����=�������g������=���=�3��I���\�9�|�=��3q�e����+����y�=��-5C?Sp^�H8<_K;��lm������v��� 4��u1����=��1cDՆx����}��ܐc�w=@����aU��~q�\,���=d^�㬥W>'ϡ5<%��=���C���xM_xh 2�Ofƒ�lBiϚ9���X�X��-K}������2����ow:9������=d�
L`�j<${�=�w4B����DI���{�=�����1@3����=��ci!E��œ�����=��=���Lg��}��E�#���p!�ԓz�P������=T��EN2�J���w8=����+,i;�G�<_@��b���f��<.��=�w7E������=$�	�ǭw|b)�<��
<*��=��=��B��ӗO1�=���Ɏ$�G�~n����|���w?A����U<�!M�ژ| E��<W?�M������%���>4H���j�j|6��2���=���P]�9�nb�i:�ӛ���y�=�+U��m�K��=��;�|�=��@u�� �NFK<_(�!O~>�u���=�� JR��(ȥ[4�U�X��}1-Κ<����zF3�~>�̃��aO�Y��2+5�B������+.�9�����p}�u{�������X��ģY稓�}�=�7�O�Rx�.�k����2�g�B���C�,���窣[u�<!��=��k/$wp�炓�w�=�R���FĚ�[��왈ч�=��U��{�6��<"��=��,c������=/��\�:T�_�ڀ�1 7��w�=��Dd��n�5¹kr��pqN���"j�8���b6G���O�i���x�=��`P��Lޡ�օ�˚8���<�@ތr�9���¡��=*2/"�
G�����=�N��$�hx��=U��{��w:C�������=���)�e�i��b�iwδ5���=}�Wu�X>����a������=�V茟��<_?	&�Ϛ5������7�_,3�� �=����vwp,!$����8���lŨy6�����c�C���-(�LIH�20�f)��=����~wp+�/�w7@����`�����hw�k���<W-�����= ���!e��*�`��R�´��=���=��p�a6�S�?�*|��-�P���M���V+@����E�BjՑ�r���?�wh� �2�c<4�&�.-�/�t.�C����  CT�����+-���=�������2�e�xT$���8!�jc��=����`�'�^�����=i6�Te3��=��BzǮ"��������=�����6$��l�M��$�mb���<� ��y�6�$���<_5�C����C�v�w�<!V�ξ2g.� �=��ϱ��� �H�Q�έ��e�0�������66��;��<"��=����+5�����=��<WM�7����A�(N��c7_w>?�����������=��=���+Sk���<_P�7���}�� �~A@��%+f��sA/�����=��2�sZ[�����ѽ��=��	ɅQ�lt(�?6g���=Yt߷�����=��o^"#��^l����=����^�K�ޙ�W��,�q�~���Y��o@�r�2�/<��y�=�֌k��Y�W/[B<^4DX���ihs������Q������=�1���<���2�A�-��������x�Zˌ<.��=������=kLH?�,9a�|���<�R¾��n��=��f_��y,̚N����G��V4����r�Ȯ��=��c�������=���^�Ȣ���iQT��C.�bw6H������=��_�i㗣�d	��<&��=�͚7�����6��$'���������=�����W)����6�����w2=������=�iv������Z(=��V� <'�w>F�������=��<�����ӨK��iѥǋ���=�\K�w���ɗQ�]�ІW5�2{���͚M����Z,��wal*T��WA7�+M	�^!øow=F�������=�ܬt�H��U잘�9�"���z�� ߥ�h4>h�����=�.����!5v!?pb�o�����¤��=�X���fꌸm����z�!  6.�
���4 �=��]T�t݌)���jh���=���K�ϛ��>C�ʃR4�
���k�=��ބ�Tv_kSJ���Q�+3pY��~ڲ��=������*�{�<*��=���bD㾆��B��23�+D�Z���)!o#��X	!�!TYή �=���6���\����2���s��20�6z���=��2�y�6��=����w�eqꄅ�H <%��=��k>��23�����=#���	������%���AW��i�������xmt�w<=���� �=��ę&Dc��<_H�i4��b�o�C�=���Y��^i��w�(h'�v���=��b�Ln�"�h(N$&� ��=��~w��hG/��3����W������=��q���=�@W� �=��֝�<�q]���7�<%��=��Bߪ6�� �=��yq^�F��,��>�%���R�*3���=h�_&���f&o��g%;��<,{�=�w7B����!$󼇖�=����� aY-�ml½�2<,@ @Ǟ��=���D���$��QRh�A"e2�=���y?w��z�=�'B� �9P�W�G�<����Yᆷtw:@����+@�oȚ6����֝�#���{�=�7��.������+S���A�o�;�+,�P����e�q	Vʰ����i��@q��Y�r�+C�v�N�`��������w:@����+.pD�g��S�n�}�=�����k��1����V���=��}�H�p�BE$7g^dMC����=���K�L4�L@l�w9@���<W@<%��=���M���_+>,*���}�χ*E���=ǂs�ٝ@P|V��������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                        sharK 3 xpupdate.hopto.org:60123 ��P��P6�[%���C�(UH sharK Server SharK The sharK Project www.shark-project.info boredcoders H sharK Server SharK The sharK Project www.shark-project.info boredcoders �� 6  K sharK 3 The sharK Project BoredCoders SharK Server Server Remote-Controller .exe .pif .cmd .bat .com                �� sharK6AT8XP1TC8��       	   	            @�@��         Z x4a>iuPsilNO>p_mrD;PzU3>bp0JAA0JS3Au@^FX=`fx1w\DbVWpxfsuLtG5=9?>e6r_1Vj[]bgb]2qv2IQsKu7xQ=n x<`Vau:rC@HQRA^g8jaiq>[r@L_9[G1dq\vk:MyYW[^HU85AC]NsTMnUEUGwK6LZT:<_AFk]p1yC]xhA5d^nsPp1qG;_thFxe6OZINA7=kZj@_ 0b50zthdzf96rtwjxwd��������������  ��      �� %defaultbrowser%����                 �, 