MZ�       ��  �       @                                   �   � �	�!�L�!This program cannot be run in DOS mode.
$       ��2`��\3��\3��\3��]39�\3��O3��\3��P3��\3?�R3��\3��W3��\3��V3��\3��m3��\3Rich��\3        c��e�xʥ�I�Uo�1<�"ɲ
�I~��CQ�PE  L �E        �   J  �     �q  P  `   @                      �    D�                                P                                                           Q                                                    .text    P                          �teicgs00     `                    `  �.data    �  �                    @  �7z8mc0m3     	                    @  �ha8shnwo @  	                       �nc4p7fr1 0  P �!                `  �                                                                                                                                                                                                                                                                                                �P     ����<P �P Q     �����P Q                     kernel32.dll      GetModuleHandleA    LoadLibraryA    GetProcAddress      ExitProcess     VirtualAlloc    VirtualFree   LP `P pP �P �P �P LP `P pP �P �P �P     user32.dll    MessageBoxA   �P �P             (QL ,QL             �qQ     VQ�Ɖу������tu��ȉ����I�Y^Ë� @ JC J     ~q� D=	�n�����̩�Dukb�X�ÿG��eA��'}e�5�����jNN�K�ƿ�wn�a&�c�j{�ʾh!�C�~)�B@"8n�Ԉ��"��"���!�E�JJ��'\���N���93�3�(`�h��DDᏬ� �MS�nک@䥁�S%�N�EO����X�}K��W��J��(L�
���C�;���ۙO����sƌv"��/ � ��%����L8�pM,�J�����15g��^��0Rj֬~�C�(/�?C���e��c ��rBv��t�x1Tw�F�]� O�q!����"��9)R�F��Dl��ġ� �]�(�V5a�*�}��J���p���]Y4���V�_-�5<\RħF���c)�V!,�~,Sdy'��b	�#���ŷOb�Ȉ�<YF:Z�r1eR�9�'�%��mvb��������c_�l`��	�}󂉭�n?=��2�6/*6d��[�����XoHTkԞ'S��)P ��B�g��o�	�1��S� �񕬶 \�x|�H�>�iR�y�F?3˪A48�����C�9�(~�X��=�oy0���O��j��o�����,b�V�~���05�T�S-�2�� a<���2�q��U;
�0����@�)�/|�ar婢�����<��oѧg�gqVY�D�1)f��CZsΩ^ L���hL�Κ������x~�^�X.7Ek�.� =E�a?��=������Ƣf�0<���V/d�$D�)&�.4��7O��FkTr3���V/�qWEA�Ф$x>iX�P|�Ԃ)
Y�^��(,�8kvN1?�0��Q0�M(sT�7]�O�́9y�?7�~���<l2�㖣�3�����d�(�H�珛�P���3%4o�F��3��"qBh�7�6�Z��8#�͛����D��y��n�iu�h�'�F�Q�?y"G_�����#]��Ug�H*e*rKZi�U_���}��Z��J��lo�	�c����#�L mg���t{$��BGC�-u��ВQ�(��B�!]kS�>@Y@*	L�Qң:��6��*M1����&�Ҷ���ϱ�����fd鬞/��=����� ���4݂v
8�V3n��S$ͦ��@G\L�Yn�eϦ��/�a���(��F7B>n���� �v���^�(���8.b.fg�%�����aV�0ABp��v?n �Ɖn6oVnd%�-�Ek�č3�s�U&7��7�C�2�T�:̪��^_W:�^�~���[-������8��$|C�( ��gd&��Rm��S�L���g��P6!�,��-�j�U��j১��L�Ҹ~������c���,k�O�,dI��l|1�Y!��~N�m�]�TV0�I@"��JȄ$�&��}�%�Β.$�eeT�{���@����(-D\�IF�b��ʵEi�U� ׷-O��j� ��%zЍ�q/<Z� _����0�]�b�`�,��6��@b�0�!��k�� m,�F����"n���m,b+L�s��we�t�1�^c���}uHaNڇ�=��1"�Q���(���v��q��z8-��^�q	�SAe��,����Q��l�1N�"e/�3U��S���`�R2�x	l�cM������Rԭ����Z��A�o����u�Ł�7���/(=��X��X��"���;{��W@à��f�:5*ޤ��M�y�SU�)�U����y��?C�_�\~� �P@��gH�8	|�:D��@��H��|5�-V
Rf�[�
�3f��3�����A��~[Xbk�n0����O���nwR���w2����e�Yq	�@l����ԧ���Ԧ�"�"ܘ�+��|��v-��u����bX=T%:�n}S���=��P�n0&�0��[��D{�r�E/f�(F1�������
E�߬����9oY�&��f���vb]P�Ʌ&ʨ�{�k��^j���d\"G�s��?��{.�xT���S����}��&[Q+{�G��y�L�t*broE��8����N�ۯ5�t���$K.���61�Tޔ`��F���ž
��2n�K�*bRL�y��F�c�ZDk�T�(c%�$iE���Y�Q�gZ� ��P����>�o�NОܳ� �Fp��i#z�׈X�
^�w�Z�q��/}��������}o��{Lm����T/�(��jXP-�����{��ś��S����^፞�O��2O'���AC7�@�|[}O��7 eFN�I�����y߄e+&=v�1;�!��o��$H���J�`��O�ԡJT8+XV�D�n�Ol�E@� ��Ge��q������J�W�K����]��"��YEl��N��s�zq	��ͣ.�������|�><P{�h�"���*��Ӷ4K�����Y,�+Φ*�/�P�S�U�UVG�K�\6lVM��cV���n�rR�.n��p�� �}#�޲�v�y7ʧ*�B�����î2ҏ��Y)��C��r����d#�.\T�G�Ren�&�8����3m��_aC>����_���C��|�b�"���0S*o�O��-��LH����� -FC�V��@�˪���=	�]�
�h~����R�8��5�X��Rj���}�F�	F�.U�a�'��&�r���7���ocJ=e�h�rC����!��b9�ȭ��qȸE�4��_0)  Lн�̞*�.���(��[��$�S�RpK�����V�����$n5�GӲ��S�c JB'£D7U�A}0�e(����qP&J��䩆�MC"^f@�>��5gvX�K�� Lac}wjjh����A��C��Sd+�3"Oyt���0�r�¦J��d�����);�<�1p��.�h������$5r܈�:�*Ao��(R� "����,)�4*Aç�Q�₌j����ܛ�spn��ۋ?���}��
���,���f�� �3�V%�BTZ"[��-�R�����P�Z�֯�u������Y�귔-�\U�{����B��^Z%潣�(�*^���Cu�k�*�D�ֵ� z�2	-���La��]@��b�T�A7�S����*�FY��ť����)��*��b<�XS&<��?�1	@;���E���X��èe�̐S 3�>|M�+- �,��xe�5��6BloQHЀ��Һ���O�?�/b�� "J�?/,��X,Y����k�aa�T��'�RQ _��I�\~��u��m�O9�6�j<S��A��kT� Qփ��o���qWv��䞪�P��)	��{j��c�>e�{d�%GQ��ۤ��wJ(շy2�U㩶�C��t�ZT�$ܖ�i�u�݇�O���gy��|�|�^peQA
xao�Q�:4������S�M�3K!A?W�h�ZN,K�]�ߎ�'�`}����/�@*����Z�:��@��I��0R['��p��X��|�P#�k3�Ep���Fh~vi��Rgv)�2�l�Ы�]��a�u ��7s1��f<[���#5�J@!w�g�:<��5��(X�.��TL�M��;i#�h3Vi�`��A��C�x��y,��sE�\�̕қ[�[���^�	!g���
�>D��_@>�z*���F��Q��'������8-�����Xr�>k��4�r"��3�f�D�*�h_��C�� �<Y��G��\�SPx�1�{��5�@M��Db\ty�,q'�t#���_���⫣��䋹|�����p@\9S7�C���s ��7Z9Bn�^�S=�aX�$���������B�@15Q������.�<k!ܩ���������9�+�>"���-��΄�]��ADTept	�jfv0|kĤ�MP���\T�}�ƾ�#���;?`@�x�eT��[���G
��"�ś���x���A0 1B��Ep��@�����:4Acz�ʼ�Ȃ�$Q����	E~�).)��jui'\�4�<���A=�P֫��� �1қ����%!�6A(�z�����?�rl<>L�3�C/J!���N��1��^�[S�(�� a;n�4ϲ��Fa�����fƐ4�`9� ��2�!xX'���P*~CT��y}��L��s5�c��w"ڊ�?�%X́A�:'�N�9�� *���v��@M�P�;P-���1Dc2*�0�MP�@��jU�:,;�ᇘ��Ƃ`*6 �@0!�[	�!����Z��ƌ֟�oըFT-*fG�bF��iq���f�]�`@9����p�h(�5 �_4D��k�PuA�B	��;N�}��d��S�lJ�H
+Ј�4Y` p��0y�ۈ�ɨ��e��ɡ���	 �(��&��}��7"����S� �}��[����n�A�(��P��Ǽ1F+���h�8�r�Nȝ��3,�`vh�������b�@�b�	��w�y�3+�;�����rGxG��W��#AXt�֯\@�; �.�H-WAd0�y%�DQ�]C��.�e�G�z���h����`�����_
Q��!ҥWv2hbc�~O$|��y'��*�(��P����T��x?}Q�a���"Xzl������� ��4#��b
|��t�T�cХ	�YFVԗ;��o��
�h'Y��i�o��t�1�f������W�jc���3~h�D+�����"��*4�+���#�=~#�t���я�1�W�)����U):]�#2�KLp6D\1���>@7c��x����W�TN��$���@�zyQ@�/`�8��ú���@�),>��;~μȝ���Ģm8ʔL�014�ڝ5�.��Y�N�U$�Q�@��L��&Fݕұ���#1�T���9�;^%�>�ARFIh����J��L���xBf �۱���&1�r� ֊ڂ-0q���*���|�"n4�]�2�.I��ܿ��4�h�N9�(��8�d���n�1?X�i���M����X`~�������#�!D��0��Ԉ\B����� IKp`=� �wƃ�}�Ǣ?�,�&��؛�0+vZ�,�x�-��i�n&r��E�������U<b{�����5)q.&�Z
X~����:e��V��M!�(.99�*r�2�اUj�.�<�P����y��T[)Y��¢���01Y��
 	"GP~sZ�"�׻l��T�p���g�==t�b/�6)��b=kk�N=%_+�wFv�����5'�D5��jH�9�WWBHvt��d��I[W����Z�<�#3R�FQ�኿��k�K�gV��%�� <�z��h����~�-h�Z�i�rA�T���+�o�����U/���3�I�
�xS|�����&����.�aX�J���~9w��<�:������˦��V�~��'�<82o�W��~�K�ی��1кP^X�b�)�/���`Eԝ!R��8��k�x��S���Sד��>��5�n,���Wa\�=��x�a�o�!!*~�x������_�R�˿~�۲��҅i�a��H5#�l�ز��@�h���[[���ʫ�݉�#
ޥB�L?��Ȇu�HyW�7�9=�
/T�E���L�q!��A�̨�1��8̈́6p=�@H��A��ٜW��#i�阡9��7��

t��#DS���+3p.D��(@�~2�sh�aT�݁�ڍ����Οv��R�F\�� � ��R��%���Ԇ�������p/�Ꟃ
9��[F5�k��q���j���Pt����A�c&���7��!ɗ��	�A(�S�L*��u~�)�1Ή��J��gZ�0M*���y�.�IR�F8�ί��A��s B$q��`����q�\�\�~s%���Q��=!4�N��~U��#��6r��GBL�9�	��:U+L2�h���~���E�3t4Sh�1Um�!"`bݥ]�<Qv��H�+�;���F����^��^dځ�������,�I�W66*)S�����q��bhuRp�X5��s��&6]�u)��`��hcj.�&��ئqV�T�d*ǳ�*���|�6�Ɲ5�#@}| ��W��]�B`1�P�C
����bʄ�Щ,`
#���p�A*;���
L���Z���[閟�H�p�oT���L�]�-=�;��k/h8� �P��Q�@Cm�� �bY�S5�i�T��9��JJ�Ǟ�T��<a��,A��wM�>D�aĝ.d[bQ��#hօ�Y.`O2�/G!z���|�
1e��d?�:���^O�I���K�v̢���/���&��HS��Z�
@�*o*�=���2g���"�n5♳��7�����Y�wH]v�E�Ʃ�#��%����㶩�u�Z�bs�}Z�*|�:�ۂ[�f]m+����),����j�0�-ž�WoX�U6ɘ��F�"����t"�TF;ED�V_�Un�ڵ�1�p�R<Gi~��)Q��X�B�韌����Hxto&Gq���$�K�i���s����,`̩�/��&�6��+"����2�2+q��*����ʹ�u�����e�x�s|S�3E5�}/���}���Z��6b<ڂjMZ����-��`�'�ت�S�lP����e����ZVhW*W%
��]E�0������\�ڏ9]�7��`�>Y�,<ړ-�Yjybo�~9a�"�v���	-+j�z83(1S����
6����8H�<�e2�
���Fi���VKxS��!e�b�Iɞ�����7�|<\��c-��e�~� P�@����A��2�Rq&F�B��B	�/����[���tZ�Y�&Z�*Z������(X�%}'�T��,	.@ �Wh��Ϻ�R��r�)<�H�v:#��9���F���^��HqA6�+�a�@G+��]P�P$�t�Y���3[���1+���*7Ơ	P���*�}��� �vC�ҧC�)BZ�]%!��_�p/� <7h�P��1ݥ�XY2�w�RĚ���Ť��ǿbc�C9��x3-�($Z����s"F��; c���QBi�֖Gx��%�ʪԹ���WZ�M��s0q����YA����G�$m��r�K�a&05�����;}�te�m��.%ZF���ڍ���!Y꺾�TǱ�u��U��3�"1=�!�詅�ztր�s �����V��KB�����RѻDU�hbN��aE��Eۅ��(������n����Y�>T�����y�Y��w(G �Z��8�T*4�����לNhNH�~�[�T[�~��N	]�?=[$�j�Q�@�-i��^���(��^j6L�Uf�y}�Q� d�6Ue#���SQ�?A��Ia
+-�Q��0�"I�^�!J�$�С�a ��(��NA�B�1�w��1��~���F��8zw��/�Ř��ҫ���+�2�
�\�
Tŗ�~E;��R散L�
HR3%���㗫|S�W3�Q(�iL�W^�A��a�V�Oe�>�Ԩ�l����4_Ǉ��nV�Q���2@���$�K�bd0���U��B2���)��ʇ-孲���a��A����)����/����ȭP!AĨbx�w�J4�Y#���jW�(S�~�J�y�(���h2D�Y��t5�6��:�g����z�Ě.��z�(����L��4���洄�@��_*����u�V�Whd~�!���|�BW�WD��!�	�X�e�j��=�h�,�CE>�-�+�U�{;"�#�uk�S��ʢ�@�F�
ݲ�|�?֐[H�C��G�=�.|����"�[�x@$�³���l�?uy����Q7��u�Z������N�ZW������K%ʌ�����x�R�\��M�^`��5B��H�l�Y��&�3,F�����eCg�7X%��27�Z��O���¿�ۙcc[>���5��ZS+j.�	��J� r�e����)s�.ڼ��k�A���M톍�S�¡.��=����h����Ƀ4��Ea����^E�tE�sG�<�c�;���K��*�r��RLSm�G��X�T7�x�<���EZ&�+�w�/o@�M�'�J��WL�#E�����a�:�)���8g5Vڌk���Z3=�ҥ�^�?���=���EhTP�ʊ	f�[�K:Ѭ�n�S)�����7�@�(�j���(J*J�g5*a�P$�|����t�SQrO��x��_TfI�EE�@E�TT�4V^�Z��Z�2ʋR�7����Y+!^mTED��gN��uVUo �� �D�嗒��Woo%�陃Y�cj߁�Rrj�u�r�ח�/�u�����7��'�0�<7�N���R4�9�ϪU���ZY�B�R�⋀a��=D�x�N�B�Z�M�d��D�sh��F�
s�c\f� UKœ�2.J�{�ٝw�JB]5�+�pR�r�����e��X��J|�G9���mE�ޓu�*p��N������K�8��E5�$��`��D��-w����������u��\���U��;��޴������@���_�
�����a���GkA�P ~���"7�Oe#�U[T啣��h?U�o�� ���H��	�� ���C���B���\�"����wڟ	}�Y�(R�#fH4w�&�_ٰ��G���[��"��O�~z�5��K10��VX`��]��h�"mq!���TE̪\����k������t�-sd��3��FY
WTR�מg$ft*�)Jb�����H ��+ ���ƈ"`��;�Q-�S �%����J�o��5
+��z$���_G�
�¸TRpc�Q��ȸ�M�qEƅ�ʅ�/������ٹ ��M��I�q�84j���)�NRb��Aŕ/7Hs�V7���#1:�(R�K�?��T��+�ȡ��,8�EE��s�D�R����kJ=�����j��*��E�۵���[n����i:U�;��\C�o�����F�iWC�Cʸ�Z�5<�h�*0.G�Hp^�	��nV���0\���#�7�������8|ݧ�������Y�E��4F���2��8TQ�����X7_�S���2��Tx����v��_\zƋP���S>�v�@T�P1
N�$�~EbA��b�!�B�'�%Dϻ��DR�]0�j��������G�캥�Y2�|'�`P�j3�@��Rl�c�H\O��b�ن�b�#�?8�	n������ĻP��Z�+��VJϧr(�WIdUYŅ�(u�T�|�BI텕yx�:�(W�6�t;����Ȓ�jU���YbU�����������,�̥smT9Es�>�2y���#�@�\�qњǔ�-�N$}��tA$��ǕBP�*��pZ+���A�D�mĊ����A�V30ڠSZD��:��@�����X��X(d���0���͇~�<[�hH9rw>klT@��괰�q����WIb9#��%<l?4)��]+���z���r)�To�ltH�f�p̥��a�U����)�gU)]P <K>B�M��pc��b�2(�9@�a�|�+��)�p�該1"�����G�B��T�|3��!vc-��]i��a�5�hZ�x��A��i*��K�t���B��e���*E��!%Z��,�����T�\�=(�U�j���p�KTo��c����*u�u�β�BHا �~�`�����:�U���J���.�;Je�����PPC�z�,@5>PZWH>�V��+L��K�#נ�4��.M�&�Rz#� �F>���G�j�O�F,���-�ta�k�F��!�kv�I�4�
WԈ+�
� ����1$�E��S�����֛3��XcT+��C������RF���R�\�	�gbJ~"������ ~؝	�V�WX�>��	�^~Sک�ީ@��A����x`�7�\��{�x+|a���N� 8(T�<�:���#�!���s;>&��U@2�}v��vf`���S�:j��ζ��>-�AH	ؘ��a�	}ٵ���"JƒĚ"T���S�*N*R)�ݳ�L�Nҵj�c�$���5��6�V5��bڍr�U{V��"�P(���>)壺�~���!��]�X$������˚"Nl��.����(?�(G������e_�,�~���E�8M��+��H9P�r���*R��ƼYD�UySA�j?U�Zۛ@��Vѕ�E3��D�A�4ZyH�o�B��|�%tQ������GO;&�z��0�!v�a�佪��U	kF�U�q�@�5�BAAz���K�Ek�mT�����ۂ�T�ue.ԩ4N�I�!���ue��\Z24F�+Ѱ�T��j�t�,rN�r���>�	�X%�Jѵ����4��`[�*�@�L�������dP�.�(���7U�;d��x����#Lޣ�(�R�� j�ǁ:��t����-��v{*�t�s�LƨG(e��:򴐊��irTIE��tj�]���u*cVɁ�UMH䜧لN�5R�@I����diԾ�*�߆�ZX��Cw�ƈ��Fm�T ]�k2űxGK��ؓ � �abQU��BF�*��W�X�Oh��6B�vn1�@y��@ٖ��"�bY���I˄���h#�/��c��"�1~��w5C���P��ZV'!�"A����P0���y�*D�}��~���!�r�}W]�������U~sk�+Ou�)�Y%�v0��.����4C�����5n��
	"��4�h �01C�hkN���4
�9J�*"���n�u��+�n�4��:&�"� ^W��ءu):l`���O��KhΫ:��l՚��V�_�H�瘳�}XA����1�^�j�ݧ^=kH (ș")
;������p��f��[n�wp~]0�����yB�\��G�$g�L���"��J\�O��(RN�`0 	#��y�*����dy��Z��"�h���tE��2	]\�a����!(����Urd���m�U��;�D�/����t]֌s�ڜa�f���-�V�Ǆ���8����A�xn��!`(P�Y��{p)uP#��J oDi� �NٕW4�0��/u��!g�� ^�x1�ʹ!5Z��(�Txe���$.�6I��@�Fal��Q>Ub�D<̉��5��1]D.M�Z��B�gz���u����h��3Q���2�9֯�1��R��m��J4�S��kN�����r
q@�ï)���ׯY��|�:�F����c��p�҂1��`G�(hk�^���ΙE[	BZ�E�yxi�>�dN[��J�RUلh��\��Y,3'�k�Q�,�<j]~H�Iԫ�H��
<,T��׳��^en�:���a���@'��/>[JWTjՂ����,�"��;,YU�7Q��M��҂�d�Me,�+�ue>�<�)!�l)]�ҍ����<=dK� �v��|���**Ŗ�[��vx��:�j�;��E�����C�8�m�;�.x��#C��B�][�qwv"R����r�5��QmZf��&Y��b4�@��:�J9t�ztsv���|�(��xf۟���"�W�%	�TGǍoJ�v���צ*�e%C���}�#v���J��?>|"T%�ȫ�D(�� [�T�a�A[.WeU��ԚҠ�gf�T����Ҧ�$Ӝ��
���I�Z0V�Gu7N8csY'�fD��V��N�%>4P_��4�0o G����0ȓ�g�ϔh}���7Xï�qS�SZ�u�_R=OD��&Z���(/�G�p+�ހ)��]�����]��Y^P��(��;��I���x� QUl��ĄY'���<9�
�-�<*��5���l=�R�َ�
��7/-Y_���1���P��Ye�p@Svo<^�x�T���'�	T��a��K�H��"R��Q�ő.wV튆�Y�_M��p�S�˵�U���蟂бH��A�)�5�#ZӒz�+V���{�A 9�>�h	qA ��߉���(���g:��(�dP������!�?�����6�0�W�y>�e|�McT*~2��i�a���9�,H1t,�0z�_Ց�v�GB����ӑu���Af Ƃ��ܕ'�\��y��oPQ$���.`і O#�# ��wV��u+� ��*�������Z�6UڋC�8��� � }��o�C���V%<eS� M�T�|�6�E�
��tk����
�ήҫz���n �Mjۀu�����\`[�f �F�1 9S�)_��7��*��Z���Ņ�;kQC�Yu�jl�c�09Ls3��ƀD���u'27�Ş.~�<q��bOѽW���`�l}���d0E){���U?�«VL��X,���ɒ�~#�RPJ}����)�-�t�-Cx��"��l���1�wT ��(+Y�%�f1�h�kN��]��,~D��@�z�Q+j�&ğ����t��/����h�pC� �fd5�OV�S>�Á�b]��r���Ђ"��&F)��)�D�0 E�$���@�A��PJ�k+!ꐨ�Ѽ8�O�(����`�D��eD+y)�f��w+Z�i��~dK�j�i�|�/~�Fg�4g�1�u%L�O�Ĩ�cY.�bf~�߱qբ���E�-�w��"a$�"~(����X���⨥jg��,(Z��z�;"�*�<�u���٨ 1��R[��\,�TTF�O�(�A�=����ndv�Ųi!gH���4/�u��vMT��jL���U���� )�� MC�mT�b�J��N`�"�D��J�A����@��-�pI\��<QF���ŐE��k�Fx��*�s_�!Z���h %�l�� ?�v�j��`휟�.=��]�&k}"x�_F˒n�j�!h�����U�v�A�+߷0��
�
���N�<���+C27��#��ㅒ��#G��7�7,T�+rA��H��!�N
����b��>	>�[���9�J,�­��ɭ��>�A徜�+�㴦/0?b:;ۨ���؇��p��Kd(%t��G�^�G�=d�#Q����������b�\��_��,�ؾiLeYV����ls�t٦/����ɭ���%!�e��bu�")/ᢁV�u�b�EX�O�t]����na��aj��8�"�f�e7�bJ�t{�0�N��⸒RE�KAr�L��}W�;�B��F_?6��[��fG�٩���
���7;+Ϣb�����%/��]2\��zfl��GV�k�e�*��Y���,h8�#R'�ބ��%1��(�:�f�F�uV��?l$l��z"���^�*���Z�f�_4�E��S����i"���L��$)*t³}�;���
�ҩ:DP�p��hZ��wb ���>�'�Y�ґ5	��C�ş(��Xf�?�	+�k�)�_��p�z	��ϟ�BPZn9���v�"xw��Ei�P��*26�2P�:*ԭE���*.`��I
T�q�Zg�:�M���lQ� �-�ꇄY��H�k�l��8r;�|<�ʼ�8��X��>�����|�p�*�kL(��-
k�d�LCWQ(���|Y��b�K����G�Ǒ瞚�lTNf�I����'�����r|�,�������ڀ^,���[�U��x�<�������uZm�0�!��V�0���vu�_5�g�2�.��)��0[X�����}�TTe-��eH�l�x#���"��;P�]�+D�έN�bm�	Eт�Dq��e|ؼ�u�jc8�(}�"eMVj�U�Qٷeg��H����f�H����gT��l�F��+�������:)�Z#А�<te5���=�o��jtf�L�ʿ���p�� �B��ة��rr���u������w�y��MH|!�L��Z=�O���I�UI�T�Z�u}1��Y����F�+H�:�犹h�0B�w�#({0�ٞB�E@��fe�dB.�<���#Os����̴��g	Rk��4&�ۣ�=��MwY>�����_V���S!X��cs�TSXF)\��ؒj�;���� d��>ӠO�/��0��?}�� :���d��8˻ʞ�Z�c�X��J�HT��f$,�p�e�b��	#k!c�A����M	��vF��m�UZj4���D '���	����|WT+-=�^��U���$�d��7e�[Q��ob����y��ZQ��+��ڭ�9�
�Z;_��a~1���C7�%�
A�:H�� �ǀwT�H\�Y���~ű�ܘ���*^�l@�H�k��B�E"yyu����>L$z��������>�8�CJRJ?�m:����8�F�"X�G�8#h;U�nW@�jP�S�J���`����Mb���SOo��2�U��-|N�JQ�{���C�p��,A7� ���οف��[���x��Ǯ[�(9 �.�79��ϐA�P��bƴ��+[d02�_�$�1�H�*��QKv�;�cW���v�Mؙ3�KEcV��,�2t�FF��Y���і� Ri����o]�ty��h@����C��𧜜��<�-�C�(yU�|cU�^����A���
o��w�]_�)_����E �0� Hx��=~�Pw,@�R���^,�`*O&��z�N �9�ě*���E	2��g�"e�WbWE��ܩ3�ɰ�Q�G7_�?�4nբ)���K�$��b�Y�%��e�r���;���\>�}72�[$�N�����nI��g$`h��ץ��[n_�af�}��f%������R,�#��/x��!�ޕsuTTm����@�s��⠌�-�*w^BH}ZS���"��'�0S����i����ī�¾��p�Z2;���?yɰ.��(���aB�+hȻ�`4r�1%��P�~��a�� �t$")])�Bւ����*{Mډ���\�Ki;�1�ĆZ�鰤7�*%���Ր/�	�+[c͈�E7+r�C�9�y���%y�h<��=\ح�$���@A` ���<e��N1��w�n}]f7�NR$�D���*r�GA���;����;ږ�[A+
gU�BW��d�p���g�m+�Tpsْ
Ϛ?>��~�v��+�?��wz'��6�
�0%`E(���Q��od����u ���P�AOb]���0uZj��eG��e1\����8Mbe������x͡1�Ge$�����C�+��0���3h@8|�A�)�kHص���(M��i~t�������e�uv[u��#�`�����a���Q���.�X�B�2��cU�Z��p����� �o��A�_C�+���M;?7�N�@��>>����L��E+B���H.C#(n��8�67��e#�F4��I�FD�CN�h)������[j��͟�_~A��K~�4�G �Oޒ4z��Gܲ��K�iZ��Ll�'�:��/~Y������g�yupJt�c�ʴkc$|���X�6?p�d]�m�j7��wj�?�"�{�����7�\c�^�ҫCk�:�0��'�!�K�UM��	�'fM~�i�Z����� ���*7��	陌Q������U�:a��������:��/0,�Ha����T�B�J@�@4@ \*���]�h�W��$SI�Y���c�Pᾈm\O�_0���9�BD|D�m��*���~:��{f�\�t-�M���/�K`�~��dWW���qy���J"v�;q�L�;����2�$�H~,T��6�g�Kw9��:h�W���%XyEfY�?t����4�It��|!햪�n���Ieݡ�U��z�|�mx�>�"�� �U���/�v�;q�W��������|�*�j���P�/IC`Z�Y
W��4��SC$ޮ؀�ռ"�dI4���Ѻ��}T7{���ݧ�>:#�N�TaƑ}Ť[�Aހ�\{`}�bݬ�e�2Ub@<O�$̂�����ډ#]��M�-Sl"kԃ:�,$��&ډ�/�`d��\^F�b���W�jN�M�B�1e��R�`�0R���3��e>�=�+B���&]�ݤEUҕ��x�������{��ՙ��$ �t�B�6	$c�S�6$WM�HĎ,��pP�0��+�(#v�zư.�$��c�h�X7�2��w5�J���$d�z *������ ��xk��k�b�Je(yl�Ьb&4N���W9[��.m��?Y&�;x�]A�����t	۝@���� D��kPy�,�F�����h}��Ш�&qZ� ]m���U�Psu��8��#![&�7$�`4�jE��$/�
3B�0�~I��@�M��U@�։x���5@���xU;PR�'`}��YNsR7X(	z;�9��xZ5Ңp�����"2���h�N�f����j+m�OZ����/���S�]o��pJ��e�v|E�P����b%0�����D.���$I�l�
�P��T2��	e�N�JC����Ч0��")���w�\�P$@��C�����t���	#IjT (�`&X�Wh}�b��[�q��}q
����ʅ����f@�[*fT+
�sq���^��@x���	�,un,��::�ѿ��f]�8�p

��c8� g�L�v#��5ζv��o�e�E��؍��� ˺� 0���W#n�qz��f���t�A� T#8!��� `'t���*���]o�y���,�Ҧ:z�:|�gMI��u��M�Ҝ�p*��׫�����@f4�x�R���ٲ�;@E�~� �/�{5�,���	�@aqT�!��w&�W�!�s��kOu��7"��Nv�O�큀Ջ� EG��)�a���M�dW��Z#�����t��g�j��QF]�8��]�0q0G�x�>���z�r���;�Msƫ�k���;�:��V���X�����71�ͨ�ZwɅ9���@76��J�8	��D@9Zǲg��a�<���j?�wm5������O��^�XW2�4)>d�j�ͦa������a�wh����$��S�$uS���F�_u1^���F�ܨ��H��[w����RQ�^��Q�1/�`Z���U��GȬ3�P2�g�U�t�gT3nVer띮k��+���˩QvR�oDh�e{_�v�$�5��6c��3�&�7�4CH+�P݀�h(��P+��^��
�U��l����ȺH�P��kY�d�!���i�NW��� &�r��@����-c;!�y���r<<
�Sk��0�ޚ4��W���4
�}�(�n�V/~kƑn�[��� ��[5��I���0�!���&W���������.��K�pD�OWE,��+j��%�� �_�����WCt����F\�	���j���(w�=Gʁ��qiB��ϡ��Q�3j�FŞ���)�#��h��Ѳ�_B+L��az�^k��Y�S�it������J�aq���>��*CJXҽ���TrE#�Q_Շ�.y{����!�<�i_?�M�u�8]�$�U5�U�u-Wy�_�~�E��J�NV�ś��E*��U��^��\����_q������7`�p�e ���o]�Tᢰ���-]D]�q*]n��@l-�vtb� +y*j�0dv	� ��t����	 ה}/"����W�~�pA:�u"W�%܌P��;_��u�I�@�|�U�2;w����:�9U�X�a�Nh��b�?u�L�/2)wLR}�G���G^�:#�?�� ������z2���1w؋*�=��Bo҄\X�P�*-�_�rF)}&���d��mվj�
S�X;.�^���Ycp�qo�S�ѯ���T�|�e�qxE�2�n6����?�8_�Ȫ�O��WQ�#w��*T��0~�ߝRXb[�~��5��Q>���X�i�$L���;�Ϝӡ]�5&���@�\�`�u!�T���7NU(,*��ڵV����WE����L ��4F�l��F��H�./��|�¼s�(G�v,(���b ��Ežc>��#f �݅D�M�s��S������	�F�-�d��n�CX���L��@�@�n*��4T3$����b��,�o"�K����#FE�C/��!r�yz�hő}�	������y��r�1V4$7�� (Z^�8K�K����6=[֧�J*���/!��)�!G�)�	��B�76F���A�޸�{fW�W�&����P���Q���@O�)���*w�wA�w@��%��Ƹ�Pؓ�%�z�ZT�\�;W�+��`�8]�^U��Go�,�χ9@�����!$7_T�>�>L�Z��m8@@H�hS�IBd-$���C��	�eO�-=S���wg "IT��v�<u�\�/��B�X��� i��8)���V�
��5n��lCD�\��}3���d��^��t�DP�Q" ��u�$(�;o���Ցu�%t�r�~�,QED�VT����X��JF2�MK�����ү���n���	��c��1�~���4�:B���̒�����#4�����Y*k�ʓ��֐ґΨh�C߆Da�*��:���7���mw,Y�k�#R�� ����?�U�%��
2�_�iWD�W�ϖ��.+x�_`��Ϻ��J�K?ǽ�˭ �\�]�Е�T$�>}MN�iV�F]E�J���M��"�[��3�w�Ы'�j�:z�a�&~���MyG�c���W�����v��U�X�.����p'�W�B!Vvi]PpI�Վ�p�u��#����],�"gB%o����U_�`߿
��e��P�!SMs/�0fB�(�M��j�Ą��ʧ�f�����%M]ϔ���텓�E�XHˍ��3֭���j���N��&�\+U:�4ʫ�#_�E����E�e�@�E��]`�Ž�]Du1�k@hFP:T��w�h�_@ÄϷ�r�fV���څ<�O�OI����7��ԙ�ˋ�Rk�$�X���T��A��ţٖz����R�ux_Lw�i��f�I8���_*�*�*>h}q�z��5�zʃ(�_���N#�P~���i�
h�PԶ�����N3C�਑���`
���:5h8?q����Y�\��֯>굄�ע[���}�a ?aZV��_e�w[Ye~��{�5�՟
HWm��*��H}DF�s2�*Q�:l�12�$�>DA���]Z��5���x��\�g���~�w�x�pZ��N�E!a�YSV��4ŵ�7�e*���U��F�sE�̴
j_BY��o_ݻ���j�21��ރ�6U��ra뎆#�h��,�,ܭ��m�p�AC�>�
Pr��ԪG���BJ�jx�v��N��Y���7����T���^��]�|�Ņ�eS�<2��
S��u�"��өS9n�ܟ���Q��U�#$F�ú̠B���ٻ|�OuA5���ӥ��/Z1ܬ��巤�� Y��R`J�%�F!n�#a1X������@X���K�"��E�b(TNV�;��Yn����b���¬��]�����V������WD���ȥ�.������wd�p�5)aU50����*?���0[|��E"�rY�uau8�����T9�:�:5�r\E�S8��dk�;�|����MSD9UϬ/�_����'�3�x���U��(�#�Ǯ���8���J*���|v�����ȸ$����3.,�gfhn,T
�4�6��(�.�*$��֓���U�O�`On�b��>����UA��e�|�'�����z����Zۍ*��-'I�n�Iu��ySv�I�"�v ��	]������.�,PH��;�,�/�+b�,݆&>NN�7!��2t�h{��|��F�"���v��,�8	h)�y%��G�OC���Ϧq=��g�(Ve�y}�bc��0�v�\�s��<:��K@��E�-)��U(��d{��x���#:�$��O�*�:#p��74:k�H��@Z�48���.c/VoK�ᄦ"�c��v�P��'[w��x��4�F�H�]�� �� **��M!���u�_kOԫ�{3%&��ީ����O��Uƨtٴ>(�4
�Q�AۨP�Mv��a�E1�ޣD���Zt�9�8JW}��(���jU��#u��"řKU)���_�֣�X�ZN��x���=��0�@QE�<�r��28�����P�,��$��[����$B
�kk����6X��ܨ��`�(+�Z�G�����}p��,ZSb�����=�����!
���)��<���`����l��.���IahB���i[Α�jq c>�G�w�qZr=�`&,���.��OG��z�h)���{V��F�qœQz^�wś��K���J\Nڗ4WG�_E�{\�ņ�q���-]��;�7�r}��P�,p�N����ڬg����*��;��J�n�4����1����>B���5�[�<.W�<21N����SO��^7��hr����X�������ٕ|"�V�x�����q��.��%��UA*��*����~| ���\xSc�8z|+ѫY��?�]�������0�]�wЗ="[r�jF�J�+(�uQ��@��BK�qD�ӻ���W����e8g.�jw�Q�����B�G�|�>��*��`�8�
i&�O�n��hs�rژ�*�k�%:]A�]
��˳N�J~;����>�V�7���h3���j��?�cy	��U���Y��m�q����}��T�AD[+��mq�.�c��6K�Lr��`�	�ўXB
vD�+)�������l��$�~(��nøh���}��Aׂ��."�>ШVD��&�!uUА�5�F��V��V Yż,����0���8,�oW���߯]�I�>{�x7(�J���>���&����[n�!W�)�D�Y��k��8�O҅�>�/ϟ=���י�S�%��ްŚU�Y��e\�tgg��g��WK_�_�z_>!��W��̌
�����UI����+9��)�����S�.>��wTp�
� ����](��ƕ�!a��8Sܱ�9�A��+��4��S E�WV��t�u�}q���F�y[2�?���0���Ӯ}W�:����/�$��Ys��rߥ�7%i!w�����?E���_�K����/�L$��N��w�R!�xWz��j#��ԧ��C�hS�������R@G�m�kj +�QL��ޕ,��D�c�`'#F��t+����a,��~��������.:�����V_�.���A��1��v��`q�ү|�h��!���]�����	,�<a�(��d���//^}hŢ�)��8ľ[��M���߈��WBLy�Xb.��H��@��<�F�35��H0̠�y�,�1h;���CXY�4`��&��=ޣJ�Z+(�^%�+C~�z\�a�����j�zȈ�P�����$�X.פ �B}R@A�.�u	I4ʽ �ȥܫA�$�G��`?�Jߌ��*+���6��4u��^�PT���o����j�t �v��T0�L���o��Uu�2� ǌ7T@G�Ҁ�����H �6b�F؍�p&��	�#h�oDcjĘ7 4���>:(tk ���a�hA���H��(����.� 'V�/�P���(,`ѿ��h�ԀjUq=�u����b�@پ$������'Z-5��3|�ڈ$ӈ"1"�D�7��ad����3��DJ5���]��i���Q��M!�Ș�����fz���fW���`��h0�P"� �8z�R)d�(D����bZ\]�Z�vfF���$-�b3W�j����"5b�F8�F(i0��]�KZĈ��ȃe�:��p3l��M�b���Rx�"���f�]�1jX�"��n�r�	�W�k��`�o����e"2M[M6KȂ�a�F�;e!B3e��L0e�͛�״D�	�[�t:�Dփ�Ai(f�,�q4������L�`�%L���g#�K�8�6�F����91��9�F�{�CI��A���!��3��H�.i���Eh���\��N䏶�Թ5�.���ш8��pI� V#�Fva'c#4Ԉ��&���`_�08��`0�T<���L�hHQQ�(� g�F䙺w& u�̙��91�F0�F��F�i J(#�a�� 5POx�י�� &�F��c5l����,��ʄڈ�a4�15B
��x2��X�2����E�3���)��"�a�/����+�����>	��<P4F0g O�� �b7*=�2Qj<�A6]b���B./~(�t�Ҋ �����������Pm��ݦN�F�j˔	/]+��,'�[˖E�����1�]�Ddo��W#�L���.�f�haf���X	2�F0�Fp�F\i��u)�����א���@tr83�)PfdI�,�����,eX;q'� ��L� ��f/��Q�K/e�Օ�ňjm1ȯs�i�ӓ�d�C�@QHo�6������a��ӧ=Qy���o�s��L��3��L��p.E#�iD���%rb̍Qx���܀���e�!e��V���WѲQdʀ4�H:�WE�)��)�)ß#�\��Ib�:k��<$1�AV�oJ�"��(�>E3Y�{!e�#Lx�'�Єو3YɐSN�=RO#К7�g�\&Ep �(���C�#�\�'Kh3��FD�@�2���h)BmĊ/G8E�)^��`�����!VXu&�7���$t<y`=CV�\�)l#ں�'NL��_�G��敌��p�
W_�������i9��9���J:�Y��/	�%H�z�U�*W��+8��q�	�"�#�N`-U�p��	�*ځ��u�K�4�;�SE�G��d�"爲ٟ�9��@SE�8G��j���戵v�M"���N���D�#��jb�nN�bu���H�]V�B�!�������d��ŵ@��B(�+��+��n��^8�竘����A�Uw�"P��J�
W�$	���ߑ�� ��}#�j|��Rôݺ���e����E�RUVtubk*�~_�a��Qc���<JY��}�w�x8T\_S���������)� ]�������"�����"�1�+�5-L0D��]�?���͡7��N�G���Pu��a�*6��"(�����$`��� rS^=���6�6����C���(��f%#I��昼��;���� ���fU��5,ϟ�,���
.\[x�L�7�r���X���T��#w��{@����J�>�ة0�������l�c:(!L���<aW��G�0�~��n&��<#�/w�as�"���)Q���WԏKЉw�Cʮ� XN�v��)֠U�*�V��2�f�T��������u���Pg���/~@��0B�
���R������Ic�\�0.퀡��z�^�<�
�U�ԇ���o��
�Bʢ�����EVO�T�3���ì��W���	�"`��1����ru�����LA��}�Raы襃�dD��L A���"k0������� ��(���S�T�RR_U�7� )s�?��_D ��a�T	ЭU9�~_�M�F��B��@�ƾ�/�]7����5Y�)�	��E^�*�Ԋ)]�(~���ff˃�:.�H���B� U'pSW60l�"F�Q[h� m��
hA�h��o� N#T,��ell`.�8��1�C�"�k$\����*����5� Xe�D�J%�������+)�{������8�*�P�,8�Bd[��c�݅�P�"1���������L�
u��-W�u�Q7]z�*�MW�.]&���1{uv�}%
��V���$L�f��:�����5#
 z�1�/Fn0X�uUA�M E���Ja8��*�D�f=|�h�&N�:��-ȶ�
�]wyb|8��o�1��w1s����s�*��#�t��E�c � �0��T�����?r�j*G���S����BVHw!/�º��� `eJ������. 6�e�k�I7 ~�@
Xp��E�_���KKz�X�덶`��{�"/��Ds�ߠ�>�Z� $svUv���+)���>�����*����pY%�������izr�K
'� �������_X�wC��+���1�8E
�Q���"���%�D��W�CJ�H ���m"������ b�!s_�0�k[��n��#n�?}��Dz�Ķ�	Hژ�>� �����Mb^z 1(�X�DD����(=�D1=�%���I�1���e�.�l��B��͢`�m ������0� �݀}x#@�@�`�LJ*0X�2�A�������yǾ�}:A\���9}6)� �e}U�G$h�R"���`N!�2����zf��°�f�ю9�Y"4��*t�H&ē!�J�,(�X�d�/m�p�y .6�p�6�@��5�C�5(�ֵ���l��;+Y�-�N-����GQzy9��+��!��=�j�-�0�-�w���z��LU���U����>���)_�)�r�t^U[j���r@�;�jq֍Z�U�$���SX=�Ll`�c� N�E�!�RR�c���4e��U�a�)�HĘ��=� ��b��k!��$I�A��!�:��\�S����v�W��i�/l�PqA�׀4����X>�+
\�m=�Ch�jv��iί>Z!kk�������h��wAP@��x�rFE3��s�U��
�e	K�)|�U��ʕD�@�;�P]�.����tt�����Rd�ę{�nК���ԫ�U�Cj�o�hc��.�S�b�D\uP{��uY�Utʨ |S�?]�{��r\�WH1��$�E��UXR}
᫴���M�!h�?��EuR�5Z�;����B���I��t��Kj�~U3�Jʴ6��Ɋ!_�>�O��nf�]�/��Q�q��FW���h�&A�������d#%�=H1�V[̻J���Ayk���+ ?dUffK�
�]����aR��)wb�;���񕞑�e��kgq`pz���Ɋ�8�|{g@�"/���.��	�f��Z5����@(����{*����:JSCN�5�J�?�PH������'��4�޷(rC�bo\�%�{Q���'^Ŵ1�����	D����;z�
.? <��ঊ����Pg(���rF�Um�� �ʰP|Eo-K���U�%�d�	.3�]�;��s������+�9\G0��t�rcC4�!�FaY(�'�N�AP.�S � N�c�����H;���1���� �$Ę1��ĝ(z�bfd'�N�:����?ť?�tWDщ��	&N$��ZE?OܝP!w��v��	�?�)W���؉^'�Y'�\$(p���J��X��
#���c0�tX"�E�ܻL�
5-��y���C��H������{�c<����;~�vp�(�����$��o���=yҥ�rp��H�%Y�.���n��Z��eF�}���v�C�T`��5A{H�m�G�3*�����s(���R�-���s�q��iʱ"ؤ**�&�Wy9��F��_�e�'��"a|�\G�E^�z�¼e�н�?uO�n P��bZR�XɄ���^��+ㅂ�$�0����)p��S)BmdK�"�j�5��))H2Z�uck&���Xb��s�W��͕�$]�wh��R���*"̺��$ �= 0�Dd1E"�����Ma������8��R�F=d��Ü\R���C�(-@�����p�bU���^AEO{W��տ�@�ߔ����-�;PT.Qժf�M4��_	�J�P������o�X�$�ybN"�)a�
Q9��+I
̍�ĉ�s�"rI�����,�͇.��.��F�NŻ!7yaz��He_l���3Ŵwu��U������%�]mJ�D�J�����Z�d?��jq�W�T?Z����%���&�(��/�!0���*��wz_�J�A潦m�yy��3�^�Rj.|�QI}��8���r���vQ�����H�`��IU4�Ơ�A-��<���Z�HUb�������+�@����?�?��`�~l�U�(��h���F!�u����h�~G��?���ѐ�}"��˟��b��@گ�T����!,� KV�>������31r	�o��I����(�G����)w��LU]��?#�}�u*��_,"Ǩ��f�t��` ��\p�橶��w��������M�����'�}w;�=��-(�j�d�Q��ѯ}n��pU�U�hN3���}�V ��Æ)L"�uxО�_E�n�٨+i�k\��ه��;3r��+BI�,���16񄾘�꘱DTk��	��An��.H	�y��$u�qJ�9��X�ę�Uo��A��$�'���z}lb#�:�h3�F����q�	wРغx�&�
%Н}$���j�(�$D�����,��ہ�Cn�B�~�{d]�;�1us��I��M!d�y]���2�<a�O�J��?!�O1��5;z\�TBF�q���OY�՜����|Nkԣ�"
����`bYJ��څ� ������m.���Lk~���h�~`�܌��駧u��I�����[�+B˟s�zl��STv���N#tջ����̹W��be[L�o��DرK6�t3��0M���.�B(�کVq+�i�o[�JÇ��*�
��O�yՊ��f�z���-Ny��8��9;[��6�������:��л�O`Zz�������3��+������+�F�����tnݩ��p��u���2XQ�(� ��T���B�q�;��0�)Α�ZVtΖRU�U�w9���z�FW�KJ���|F���OH\$I�C0!���{�H�I^�l�Y_�)Zw�ئCcvP
<�ud�
��W��[�s���hY52���M̡u� ��r�,���(~j�����a~`y�/`0�d���cb�`���k�`]|���zi����¥�J���=����I��1TI��*�Νj-
�4��u&'!G�ҹj��R (��1�*3�D�5�A�o(|��8��
�H>;�Su�4�w��>���
z���o}T���쳮���=`���gi�Z1��)N����&��\p.���� ���g�����}Nݽ������<!��ȳ+�	��O��x!���J2���*�o�M;:J��wO��.Q�������巏�Q�<렪xq��Z�(���f��-��rX�8�P���СE�5��AwG%�R���o5~�t� 3IXV� �<}������[�,�K�?F�k����3�2�4n�z�4��xd\���Z�� �cZ��V�6Տ�Z�� ��Ԏç���� �ii�դP21F	��;����P��O�G]hpT���kD+U���*rQ|�j�;����S=;�ZU/�h��w0��y+h�@��gJ�i�����Wpnw���ْz�+�7�Z���#� �ԋl��ܿ����`��r�|/Ws�� ��A�6�&GZͥ���;�t��׬�;�ȁ����ΪuK�~C�Q��>'�˺��)� ����(�/�"U��c��CUv�*+����$��P,N���:�̋�������2��+'��P-,��.vlw'�2���z��C>|2�w\�v�Ι�B�Q>~�}�YQ�\�3vG���Ϣʙ}S�+a�*�V?���F9��C��0��Ijˢy�M�T������Sj�0�=�Rx�=ԯ@�
	]�"��҉��QM�0vXs�/#]�f��I+�WԷT���t�+�0��`����9�4ZՌ��!��0�3-�$S4Th!�=����XGELߺ"5ދq����3�gJ�.�UBYnN�ʮ�����&�Ga�F�W��2z$x�<��5�r^c����om��+
ژ*�
58��G5ۘ#Zd.p��?�J��k�)��Fr�*��Y��h�g]j� n���|�D���� \@�?_���U1J��@��1Y�V�"�7tR���w�+�u�~���X����H������%�|�n��7�?��[�/�:�נRi��8e@��ѳ�Ʃ�˕��H�`e�p�S� ��	k�31JJ��()G*X:�����Pv¯�l<8��Q��k���U�*��`6|�gm���"��]%]�L�N����0����XrD3&R�R�yQ�՚U�Tm�z�n@u'��(���`���ǺK�8�T_6-��2ZeC���;D;�	�{M\%�VE�����e ���YZ�ũ`pzP3Lp7hm73�UQwu1W�]X��
�2����B6 �z}�2�n�g9�o����"�l -J���.�ș���]�]�D�^*M���+��i`��kQ��ӕXwm�e���1.he����.�g�3��n\Sς�~̥�vK�ͩ��_�R�/�������#I()���e��mܤp�asAR���~%`^�ݶ�Ǭ�B)�E>{*�qK�4�?�g�������VNE魍 �"�p���g.qp�9N7<������6=c�F�O��.lTk?�q�E[�]sj��2����������RM忬 Q��٢Fs`T U懼�!/ߠ`�`��y��4�G]�n��	�~�Л��c��?�o$�^��+R��4�A�p;�$�0(N_��g�֏j��̸�.�bg�M"�,[K��@����G��&a��m��N0"T pp)ϫ�3N
;�mp��� �l��C'r���jk�2���Q�Hޥ6ެ����Qu�A���d�w	��;��J�-h�҃T�`�Lg嬬P�������.��R�CQ���B���h�_5щ'@p�Ve]�m�����oQ�b]m*���J��7�vȹ�}iL�[fMh4%
#�6b�v*�����s�ӱL�E�
tu\f��OeG_#N*�\�K��8Z-��Ge\���5�	F�-A�� (�G9K0�k#�,0|�r�q�@G��m5%�J�Ɠ6��_ufc_Y}���m���K�sȯc"k
n,�&�6�ke��WvA]��<ژ#�	C΃0a)�]x|D�`ߤ;'s�ߍZ�~>Yf����Ic 6g�Uj�9�2l�F��2����|}w�m>F%����La�w+~��b2����� )�*0x�n��C�>���}j@�0vF�z�-�:��+f�5P��8)��_"]{����*]Q�ed��d��h�(�T`%�t����q�����q�h�/%�<��ϣ�� 3Z'G�P4�S>�Nt�0�d��:@����P�J#�?v������Y٭+�LZ7?�(X�^�k�C�&,`y�*,X���zd���,�eRW�"h8�d�"���11��Ҫ��첃 ��$���M�y1D�6YI���ZO�l�}�V���(���U�����Z��I�`XT��>d��u�_�v��|�O����5�D�z|
8�T���V	����wD4�Qq^���������*a��ZB%tcmoh���T��ơ�;lDb�u6j�EHڍ�y��*��ؚ���Yi�HTu6�Z\L<{����e���	�|!��&8����%�7�<�zҶ�Y����)Z��`�h,32'^�
���.O*Q�2$\L�Jx�-�w�0����7�_��}�D��ъ��+�a�����U�)���GA�h:ZO������@�)68�&�*�8
��D�"�)�1��ɜ��2�:C�F��R�� M�&Ov{*��40^���N����그ӂ�	cE)�1D`�(���
�h�2f�����Oo�F��u���*\�Ś�EU����.��n� ̮c��P]��#_���ǳK	^(�ڐ}��EM�W`e��N���|�|�Y�ȥ��*��-���Al���q�$ym��J>�<ì֋e��f=D��)b��uM������-�����KS݂w��9q������څ��/���T��e��?��:ћ��^�l�عB�I�c���6�`��_PSʰi���RF�+	��Z(�#?��:�8A��$�y�q�Y�(�2=�. �y���P�t�%��/~w��EE0�hܙd��޳�,"Or��w�`��\��o���̬i���f�W�yરФIE�_�60G�&�T�	,!_��7'��������I�� qV*�j=�V���)�}U� \#�3�V{�E	%�����j~��2��>���l��y�G�+�d5��j>���w9�M'(VWe��b$�Z]n^�P���И0 y���fsv-߉0d��$|K�-�K�U�?��wC
&������'�DPbmt��Fy詆'F!��m�
8��H
���"����f��غ<a��_��5���J�,�����>�h#e�j)����1%��� ��hr9b�4��G$A$⠑�"��G-���Ў8�1G�o���h��j"�C>bLD�G�9��u,Gl�k�	)�0e�k���-��&W��D?O,I�s�"WC�/��#_�h3E�R��)�����^4�m�l#�\6"���<��	3Q��'��h�kT��F0y ��'�	n��!'�_kt��0ui@L��Dq�HXz�F#V���G]q"�]��'�#RPCErg0�DG4j�U��<1�	!���oTQQ�6��	>]���	��������D����7O�P��
O���j#<�6"ע�u~��	�H(�r�4M��؈0F9f>W��	/���'�k"k䗮FiyjԐ'��y��/S"� ]f)��`Zd�����҈]��b��U I'/:P_ ��YQ[灈���|�	e4��vʧ��+�l a��%o�{;�
��'�F�"n���FTym��'��y��k"<q6�2QO�U��r���hOt�lK�3-FTyb��&�����(ڋvّ;����E�� �I�S �V�x�Ҕs&�\�IL#��t��(G�P��^J.{u���0{�L���<���G�<Qt"C��t���<D�7O6���{��1����F�rP���%SB΅s���L2���'NyyBSS�:��	�}�X;�)f�����I4O���"O|���'�L0Iⴛ�:�櫓L�:m�es�����OD�l���7N�y�d�'�_yb�'�N4aj�����R7O��)�My�;��	��B��JO;�)Y��Ə�uZ�5+4��/�����x�����V^ZJ��:
L�[3!d�N�&�Eg��c]�Ǹ"�,�r��ZΥ�VY�\�.I��Y̧��K�����GIC��&�w~i���Q^�)r$���N�V���G��m���^�z@2�B�6���+4����.��i������I�F��v�m��"��#"W9��Y�Zl �B�2��4;����2�{	]g>@����퉯�ejG�H#Y��##����Ҋ��,(Rz<�c73Ԍ#�ͮ�d�0k�{e1H�����6�˯�9�͇�e1G!�j���Ұ�a����K���[��W�J��_pj�\�/*��7�<Y0W��QN��\	�"�� v�Z��aZl�O�3�a]^Rha`v3$�/��N���$Qt��&���8uR5���z\O
�YR-��U9�c��S�0���c�]��"�;	r��l�fPy�
ˉ�t�v4�1E'1a��iOv`\�z�C$�81��kG#ڃ4P�*�ժD�&Qw�trG	a.e�&��Tq�<Z#9��g����,u.�StF��&�����֑ty��l&Ŭ��H@�`���K�H[�
Y�Ɠ]�y��'�Nqb줕&��y��b2<v%O|��D�I�L��T�'���IN,y"8�'�<ae�T'�2u��x���扨c��:�	��h:U����B��I!O(��ң��ቌ�yb�
���d�&��yz�|�<�w	<�E�;U�SK�;Y�bA���S���UtB'�7����nST~�Q0�vr�./��/0<�d�O(�,���-)�.0�L0;	�	�{���8O|�	/��:����i� �Ė4O`���Ԑ�N�ybH�'�<!e|�̤8!�NP&�2!|Λ��xy��K���tZ�'�<���G�(2�&N��z�����E��6U$�������r��]�;��oE؋�N]�D�L�!�A�O%�b���w��]�aY9����zĪ��< �Sp�y?�R�*�00;���w��甇����L��Zu�р,L~Yh���HfML2L��s��V��*���-t���W��E�%�����U���F�"��c�"SU�0t1:o�)Z��&����b��<OKγ����>gS6�%�.�@�zo��3��U/Ysֶ����B6m)�v���C��s�~M1:E�l����,�TϽ�h�A���!66��Bgq�G��M������@@$�}8Ē;D�Kh�;ƠT�44k�ԣ�4{�Y��pc���Ko?T�u�i�Ǧ�ɲz�(�E5�����SP�����;!�`Cp���i+M��-���'q�E��}������1�'2�.������Z�pY�-�-btN�qY���e����O\�L���/��S�N8]�V�Tǁ��\Q1Ƅ�Bҥha�s��U@R�rZ:;��86B���:,�S&��B������L���8���x�#�UF�hi=t�:�D.$�@��$�Kw	�ⱚ�h���Ż��U`����"�ҚwPT:X�8�;�����E���i�%�#W\OT����N���-��Z�u�.�JM{cNZ�b���?0`�%O��U���B�aR��һ���(j8~���d���b�:U!((���ʏ�e��i�~�$��ǂ��E����!�9�"�X-����Re~UiryQ&>��~�\�s�L.�.IC�/�Ku��w�JQvl>��}�a��Y�^���1#uf;2o��Ů�o��ɀ��₋`R�:��z�˚̮�:��΂�@�1zJ����$�Y�.1��VJ ��܃��>�����B�)_N��WLuC�6S�������(evׁ��s�'=�ɇ��/@R�H�����1E�u�d.�E�*,��=3����j�'3(��^גh4� 8y�L����ፌ^��5�L�\h�3�Y-�&��3��Zi`�g/a����/�Ǎ���49-EWwƹ<rt�K"� �1�D@�*�s���+B��&���W�1��I��\�`����ZU0m+$������y�on�*��0QTQ0�
�(,(|Y=^GvEL�>�~_�qx��������g/������|�kƎ{[��=�.�Um�~��X���H�e
g�����al6�K���ݛg`�y+�W�Chku`]�|_s��q�Έ�&���*.N�0,�8�Ֆ(����&V L�����"w��Я�1G�GP�t�#UU��T�~�5Urԫq���U�3�˷Ԭ�)<]q*��QZ)�-�J�zC$�aP�6F�T�0��i�	���ZXpG��@6��e� ���9t������	(Ak��Rf�И��#i����Hw��Iλp@|sj0������.Z���+���v�����m����d���1�i�p��gd�i�}9�������v(>\i�Z�u��&Y� ��;�]�{����{���p{��'��⍻�� �5��Ē"�d!��<�Qв��'�]oo����j�\��*w7K�֥ړ1�͢A}��+��1TK�����id��ok�P�5HL�,u蓐=�cd:�oF�����>"����=D��hP�D�������[��E��[��X���$0�ơb�;1)'���Z M���Q�;,)�������.�D�z��Z�gN����~���I3��H>i0$�����	R���(;\	%_oh=��C()�E�!�ړ��#������"�z;��æ��,e�*�����<��2<!$2R�y�2c6�F@�J���w�9�W�Q=��0d�e��y��j[���B�cE�Y�{�����z�?���Q�4�]n��떷�*A�d@ݏ���c��$�3�O�9��4�3O�9�3��b������3�9���g�=i<e#�R��H<f�2U�H�oI�x�j��[�h�W��5��l��"�D܍�jz�ny�n�TK����cC������F�N"�R�5�s��e���\g]@5X���L��-EK�E��z����N���K��D�5?�#�,��(ap�����E�(@~V]9~����e�V\�r&�S~�GMt��g4�������E��~�'3<f$6��HJ�^�m�{~T�X��Jk��ڟڅ�9��H�,5"x�j�Ds�<jK�
ב��A5EyYe0��Y��^��:��K�<ˑK�YQs잨/�F�ȵ��V���Zh�;���,�B�!zcem破6��3�+����䇦��=v�N�����+����+��|��ks�cV��!5�"����et����b'#p�bRY.'����i�̪Ħ����ǥ\l�0�R"Up%pt�9�5�<*���7S��HqG��ڀԌ�.�ּ�uֱee>Y��@�g�m��O���)#�M]�����w\SlI2�,����Ơ$l����J���-a:�sWܦ��Շg��.Jl7��.ѳ>�v�;��iW	�R��W![����bP�_�-{%x�b��ͭv+Ч�mb��N�r��-�!ߢ4��2�
�{K׭Y�zj��h�!ᓊ����!��}\�^l���5^��eke��-�䃙�cc"�^?P�R�9�U��!U~�R��f`��O�>�g�]^�5y�oEM�z�2[qe�6�l:?�<�"]�)��y�EG�d��R����J�]	b���h���ȑ֐P��v��0��MX�aW�ӑ�M��j-M���<7����Prq`6��n���p�>�\/��ۖ+q��1���G��:���1 ��Mٹ�#�q~+���p곈7@��6��?��8���*A7+LH�Ԓ��XE'B?N����\[��rU�ܽ���H^]p���G��ռ�@�@��	bT�4="MidE/E;<^f����^�>�H��a[���O�JXj��	t\+	kY)�Z�ƍqλU6+�XF��֥��L8&Z1�=T@��11A��̖8Z�����.��Q���(��>�2����̜�:�%�OB� K�S�0oKK�c+*ES��(�Uh���ጲd��K�cR��_�-#�x,3�Y�&�[ �W2���[�y'��)-S���r������tR��<M�]-�W��u���9�]،MI��UVV�2Պ��6|/�3�m��0��Vi/�ދ���2Լ\lTe�M�&�&hF�Q���������ҵT���މ�|�o�z��&t�:F��UM@�̸�[��37ƚ��P�����Ub֕�3���A�ǽ�����JK�fSũ�EO_F���j+�\2� q|+}�q��*�/�K��]14�wx��*����<g���ӕ�q>�:^�=9�cS4��jj���Y9(-����B(-�M��,xt��69���Gg�ڥ�jF������υ"�z��(�r��2u��E�1!�}�W����se�=g�^]�Z�Yԋ����Uz2K����C�>�Y�T�ʑXM��#c���<���9˙
���52��ҋ������"��xu\`8H�/Ƹ�xl3KR�����U���˝����) C��(��mӁ"������_�"�ྞ��e٣uU�mp8���v�$໡e%>�r)��y\y���+��c�%��b�!2s�,�x���䴳��(�1WIUƖ��&���K�pt�^�7�&��V�Q��5�,�SGm���tGw�ǁ���#N��j���`��W^�a�3�уy��,cf�|�&�S�]2��p t�|�p�7����oT���M75j-��>���B�,{x�'Q���e�{,X� �梎���$kkf�W����[��`[Wr-��E��\�8�2�Q����FA"TA���u�ESr��laQ�q.>����+���jb8+��~�F���L#����F/W'/WԊakY�(�MZ��8���RW���(\4��k'��p��6����\V�V1�?��yT.�u��ԑҶ濎��
.����U�H=�\�E6v\|���TԊg.r�r�~��e*"�����؛/��J��������\)�G��e���_}@�S�F~l�ͪ�$�`�Sm!-�p��gI��E�Ѻ^�-*��q�܇�n����^�0C��õ)���<�au�~%We�ԏxb?&ܛz����}����'��w�m����h,i�lV�%�T%tgiќy�ˏ$�����U-X��{Lc�,���3��v6���h�T�
�î��ʭ��Gp�{�Пj*�0���?��6�
��X�Tc/���5�8����ZC!KQ3���}ץ0U
�Y<�P��B��k)TjMQE��YYT+�_=)�����NMx�`;y�Aހmfu�J��b nVT\�GH]�N?O�Ѩ���Ģ"�zw��M�qY%_�����	���̌��2�����>��87k,Nn����̷������g�Ix5 s�n�b���1�!�JE�"Y�Ȏā|�*.�.����X�x�F�Vpa�:���@ױ�'�o2�>���#��S(QP�����"�(�����Ui6n���:$1t*{3WF{Vz����FmR�4J�qv��)r$Q�|Z�B1�BU�=$5���X1!=�c�b���@�h*Z��>
��~g��_z�.P^������o����+�7
KB���$��,���W0f8��/� yF���{�Z��W��u`v��Hw�=�͝,���C�?��c5<7}�iQ|g��U%�{Li�N�D_?j�V��~Q��,��F�#�'uf��y����X7 ������`��X�����C W(aEv���BgZ�@C�%Z��Xz��{#��S�1���hŨV�Ƴ��
�f���ߪ?A��6���`�*ܢ�(�)����"���|s���	��M@��j����h��(X�f�q܏��z0�0�LpF�hwF�o4uqYMiP5ҧ��M_Hcg�M
=�~��>wQ`�yV�x�q��N�=���r�PE�i���	�Mk���H��]d(Gd���h#�d4�i��¬Ѫ���,���M�D��&Z��gd\@��H�0"�0\��oi�����֣���)r�a��Q�M��z�+w�9��'8E|[TW���T����8��E���ҌH"�u�俴�}��Z�E���HJ&$���^Ԃ�5�<d=�����L��h��+�:�@s?M6A[?3�z4~饯$�\_�T�M�"�;mwAjS����$x���y Z��ܨc�w��pw� 2����|���1v:��8\nit�׵��q8�4�����:,�@"����E��l$;�t�S]�fjoBK*��+<�;��˚�p���(�X�O����ZI���;��b�3n1�t&����rs�u���2˝�F?5��Y�şBE:4u"<w|p{^ْ���J�ըT����
�U0|p�#�l|#]�8�(��T�[."�G+Q�px��Qđm��h5k�p�=��,j���b�#�b0]��+E��sl̙h�0�NS����AO-a�u�[-&I��L��g1d��

,u��:O��lF��/��+��0:/W��w�W��(7�uH��@Vn\�-�������+t���ի'���s�?�]���s2�"Ū�H0~�[!6,�\rET�"��Xu��1���*8�Q���u꛵�#wg�_��r�"5>�y����A�hZJ-F���H
wQ�f�U7 �z&ν�C����R*&ھ�z�t(�'��WS9��q�𙀳�U�j�'!�!��	ŁJW%nGQe�Q]���U��SG]foG_tk�
�zU�i�o*Gn"`���UR(E�;.[Gu�~��bދ�wb�� ��w�h��j���R�sn���!�,�����eۊ�#SqvE��U��yVwB���::��	�Uq�.���Y5���>g�ۇ�{b�/o�HԠ�Z=��R�R�w�XY��31(*ftHPT�Y{_q�n�����y��1ڗ�9���&��\����a݊���
���zMG��Ƣ��8t�"�U�⯘�Uܥ���L�z�@�.Н\x�a&��(�oN9��y���T1s�1�6��|�Lp��m��J�ؠ���~����7f���#��B�N�ð_�(�j��1K9�n�3��lE>����m��&.��4����h��������3��8�a�u��d|��$���b���S�v�y)��=��<��m�}���ڍ��|ԺN�l��1�c����=����(�@��g�@�����#��ʫG(��f�>3�	JS�v�E��̚���Uuܓ+ݨ�~�U�I���rv��ĺ�P7�ss�q`b�F������S�Ug�#F�����G�g�������,bqc,!QX���L����)0�}+�%7�k�*�}�'�1]��������?:�=�v�
��(U1|��>�R7y<��(c�V�%?���a�`0�b�>1�-���:���;�k0r3��T���e\�O�hm"��R0�/Z��2��ת�Y-3ELPU�:�|?�G��7�8���bx��Ϥ�
?C,8n���8z02��NU�aWiWfAq�?'J�][({1�T]7>��cF�b��1J���\Y��%��8j�W�s@.��� �1̘�(�j7��b+�hb�fQ�j��Ch������S�����6;�������`#Z�nN�u��ð�V���\π?�h �+�D{������=���[�Q(*�
���"�ٔ�H��F�}[�/Ҍn0��ؽ.�&Xԭҿ�Z?K��7?����q��(
��F�+��(֗�b3baG�b�c�~��!�:���E�dEE��p�g!r "�J���mH��yUB`p�?f��}�'��$	C}���o�#L]V��RN��2��u�/z�J����*
�r��uCb���J	j�UF_6-�����oF�?$R�L�c�@�&�6���]D�2��0�z"������8�	�<��K�T�p���G�ݍ?�k|V9z(_&��^�$����P��ߨA
�Blm�»�;���"�JN���zF�O��9J-M}�0
�9
�N�@�����^��\՟r��;��s%?���t��F���J�\~tFK���k/�R�%X����Qj�`�j��k�W��C�����I�k�hfO�oZ<�.�E�ֲ)�R ��--1�H
.��h���ܻ�x��R�G�E-[��Sq���I�*�zc�9C�G%fA䄲WYP��ćƊ~p_bh7]̢T������h���+(W#�����nvT���"�cU��j���8V���*���Nz�l�P{��������R�<���dA�D	������V����=fy*�2�Aܯde�a��wG���G���Ƚ�q�k\e�/4��t8^�%�	6���h[�v�Fc<���R���Ѻ�/l��D@�$�����#C_���%�ˢ�#E����y2$9�,i��5� ��U ͥƿ���t��t#p�o�]l�qM�1�8��@��(��E�њ%0�;a��%��(A��<8NHp��SbY��LnV�κ(p�x�D$@�/	XSW,7�3�#�u���U�	Ҿ�21�o�uƓ\�-H&�Fq�2M$&(� ���hI/̯2kő��5B���4]�� e����t XGu�MQ�HQo����ZV|�`߱��}��W�2z��.��Pn��+��Jj�7UV���3À�æ;;o��^H��eu\.^�C�7��o����04���0&�/U�B�%�pd֥_IEڅ�HIҝ�;�ш��"����-DU�.��@���J���t�.���Pԛbk4g']�۫4������p�hoW��F�q�<	\���0�ֵ�����t�ɻ�|s|��͹*X�|���W�Qϊ������.��V}v��Q>�}��Wmgu�����9��8*��9�����e��o9�����U�
�싕�vWtDA%Ȣ{UZJQW	R�`t�
�l��f^�Rq��}F�g^Z�����{6�E.���va!J*�>hE��&R\��	L~���P�� w��r����*d
�j]#��	mv3�5�(���m��ZU"�b���A�&�2ʈw@��9�&�=0�hK��+�i������+.��BG[U6+�0ݼ��';�ĊP�L��8n+���T��$���3�y}����Y`O����*S0�ʆ�\�P�U���F�+�t�5�.�A�tL ��8�����c�Bu�*�܊A���{��]V�1�(����}&i&�e� +�n>�`�����7�u�50^_���lZ�"�ۃ�Q6x&?E�$f�v�7�v�r�+W���7�ˀ4I�9"�jYi[�<'Uu��
��A:yf�RU8�j�e�UDr.�JS��8f�E����ޏ0x��V�����4�ES)���Z �����hG�Z�gM�]dw�"kӀ�+Q�?m���kg�k�x+_cd�9�Amì޹����Xd�%-�lʣ���/����#�	π��h0������棵:�߭8H���
ę��(o��x��N�?���{�����
�Ԧ�`6�e�J=��F^7���_��L���bҾJ]i��
æP&�p�Ly���:&����Dj}�d�%bZeѶy�)|e)�u��z���Ve�\�1���Mh���U��:���F���,�8����GVF1�](2WVL=m�`֥~�!�يv)S��g>���	 ��e�Z'*� 3��]!6�@�p��M�2}Hk��>�O�8s��K�9W��3���CF�"fP�v�B{i@`��4���M�W��J	E���(��Ȼ�ʳ�jǩ�֎��Jcy�����~)x�UU_[��I��æ�1��BNڟ���^(�TD1��(�P���z�~�^���"0*��b��;ؒ�g&���0�tԵ���G����u} ԁP�_��<�3��߬�RX��(�D�JQ����u�PQ�Y�z����<C�tG��j=�Z�
�d  [<�*�����.�pg ��K{y��
������:��է�E% i�{S�3�ʊ~�
~]Jĉ�e�fq=�����Y�G��8��ۊ����za6;����.���&c�*�䆳���[X�xB�KA-H�@7�͜ c���\�����S������]i�&�	k6��;D5-���xH�%gq.�%�_E�s��F�y�vF��Y-b�7�~�������i�]�) �ɹJ�>�Z���XWE��]�R���Q�� %���K��
�Cis�A�'������3�Q���i�x�+ɠ� gF;��"���	��0�@�1ʻ65U[�"��X�U6�zRUfY��Ѥ�ד��K�^?|�%
 q
ЧJ�oaP������W�9�.�&��������!�Q�Ze�5֢;��*+�+�v�c��-�QeF1��dK�q{�GK�I5f솙�G.���b�
f�t�L�
�������E�[!�q��붠ڎAy���	�#�bk�4 Z�j��<RQ�W!%؛vv~��)��VD`��Y7�\���o�3���]("�qfT[�]���z�����㬁բ� 6�([�P��5�� �qLѾ2�ќ�/�Ձ�[^D[�z=�)�rMN���A��� Lp_`EEbw�f틢�0��W
V�J�����1��/�h�����Z� ��s+G��fI�	c��Ę�B��P<��F�wT�?�a��c�hWz�9	*Q��p�J
�������A����ڊjET�.�A�����u��L�^��\�`Xѥbb���>+��ER,�3U���fl/��8*��r��ʟ�9�jm�ʿ���B=_��6e�~���bW�Tk��ҍ�we����R|��T�>M�s(�<"_5��"
�J �:��bJU��Mx�������^�e�O<5�W0#��%���Bi�R�ؐ�(���\��=�r7�)/�X념��>^w-���7����ht�v�;��
K�	B"����&��`�ꄌʋ
�P��XZT��$�I���.E��GMj�c�6y�i2�x�3��G�㡘�Ɇ�Łސf����j೬�+̵��gL}6+v1�#(� �'Fi��4�Sw���,$bx�~��z3.Z�w�+�i�uh�C��1����BT+�dV(F�n*u�詔���y�Y���Yx�Ee��I��2�M����Ǟ�GW�X����j&FQtڽ�%�Wf_>F�`G����1a^,���~�g�Y�t���Wa`^]n���D_�E�uN�k��4�k���P�rN_A�N�=8xb�u!^E�r�� E��Z*a1o�����cǸر�"�c4�U������2i/-P�>�Y���Z�ؾ�ʸ �� w��������Yc��+�iy�S�NQ$"�V��s0}$�sg�<Z�T-���(k{��h��OAWя	W�䏔�^E���Q�pUț�h����ѯ%����R��
N��l�1D?��G�"�=z20h�B4��0�$е��\P�� ;!���C;�/����Uy�,�oUL���X�ʌ�+��&�_���Uqo�H�G�A����ea�;���b�U]�
��Q���܏�w~>��wpUl#L���ɯ�pU�O����"���9�F\��-��O�����V}�i�rUQHRb=�G�p�\"�$�*�܊j���+C��y�'��I]�M\2>A��
��أ�-¾m��	;K�E�a��E)O�m�Z���Y�����m�1C�щӇ��	]�A#�n[V4y�rX��t��4����^[�����p �i����4��P��m�I��W�b�tKL�5���o��,�kW�_��#�P����|�I�\�E�T�U��Z�?Ʊ&/�ܭwh6�,Uk�%�Q!��N&��L�&ђh%��)�dQ�H�$ZȔ���*��`�_Y�8|-��U וD�i��p\���IY��ϊTF<;�D!�Dj��FDԐ�l~H��O.9� ���D�AQ�2Q�@'����fJI�Y�d�t�*� �]e]� Eɇ�|w�.���_���R�f�.��0����BN�ZJʨ�4�i5�J��EBt����cU5$�$b��	e}�x�8�aq��Qs��*���y�tF�>����]��@u�"�'�$�ʊ�S�s]�ݘ�X�!,�qa��cD�x��&���o���V� E�1s��XE����E{ǅ��Z�̬1jt�ch@kKxʍWK�ss�.	%�S��O$�APm=y0iW��d��'�ℬ1B?{
*�+c+��Q��3��UON'���܉Ki�NY;2�H�����VuT͊k<��E--0�h�5��=�����4��UE׃�����B�Ott����CƘ��q�ZDp��Z���bԡ��N�$����������YW,�����[d��Sϱ��'�9�kgv`ayh�f�A�X�?�8��޻4�oژ�+b1 ��0��a,�>��W�:5�o��aeY�&�r2���Cb�)?�@`b]7%�Y��T���o�jgF�"i��З�Áv��ޥ��=VK����l�BG+�K����1X�{�k?��K�NAד�t�^�Y��t����
�����&�y'�H�G����gA0���h.c���≰�S����|��f�1�^�c x�Ւ�8��d�� ��4�Ҝ@46m�}$)��U�O>@�'��u?�?�AϢ[�B\ԣ֋�/¼�I>��L�FԷ�u'ױ�$�lD}�~HZ}�w��yDA{����״�E�"�D}4���(]�&np�*Q�uKbT�D�EQ]�a�Ѡgkqvˑ�9Mߔ�}����li���
�O�9�����һ�L!ӽ�ÀѻX&�.|��cֶ���K�9A`H�lbv@��1�c���c��t�LA��T��I�M�@U�7�Ž�jH�ﺹ#ŧw��+}�_�J�	����{֕u���K����c�9@��}9F't~,��8��G�V�3`;�>�� �Z��۠$u��LƠ;��Be,P��U�a�@��_^�	�k�1�mwC�|����f��*�}���!��B)�$��7:Ȳ��H�1��S���6WV82
����N� �c	w�'���e���L�+��cT���|#�.{�&�H!4h%M�B�_L�]`�'�8}c�G�X��G�4�����ԛ66�52cT:7��`mj���������](��峠� s �S���M�[�5��PZnFP��"�H�b(�����Jvˋc���3�3Ar���o�w�L�p�$9 �@�*|eB
�%�j	�eՇ1�>��G�Q�,2*���f�Ns�Mb2�,���91�)�6�5��8��0��[|�����,��7�yΙP�
>Py3����ղ�4^=#�����Cj�;j����UOt�{��/���3P�Vx�F��7��,���`%DTx��0a�Ӏa�%N��W���S:K2nsÚhg��4���+�C�<yB�q��<!���o^}_Ֆ$������%]$�"��82��:�U9��Rd˳=	R����
��L�V��S��j��9m�4 ݏT`I\=g$�"� �;�J���b����C�%�S�{�he�_�
|�W�_u�ZbT�[ǡcU���C����b䲖�aŐ�1�@�3c�k�f����Ϝu�����M���mh(K�s�;LfV��g���3`H�_<!x�	��i�L���;cҒ��,\J��I�W�<a	N�dќ��:���L�.g�1p_G����E�f�W�q=��!��)Y�s�cw~�[TG��af�uA�=
��Y����� �b�`$1�L��2F��_Ɲu(�q@��ހWϷ����32c�baX�0���/�y�.Ry2K�%���� @VyWĝ��3�}�����u>�:��-��.��O�!ع�y-�q�e?HQq�Ԭ/��᤿,h2Z�a��k;*��.�����򹨖>Mr�C�"��:���HjPT�j&��-��N	GV,
fuC�3��?�O�*�n�n��2�Q�&�v�m�A�i����?�N�HST��qy�����E�B�qr��9u.E�O�x�bj-�+�������.z�� x�F�3���D*1����Ү"�5��a�116�]�I��J� z]��i�`j_� <{|�Y\�N���l��-�����|YD@�� �(�Y�|�q�WI#�
WX��9���O����W}q[]�F�0(;�Nc���+	:O# Al2��Pz���{ӯ��q�����9�f�x��g�Ɇ�U�y����C���Y������Ot`��\�D���׿3���E_���UGW�Uǽ_<�ɕ^�U(eV�ϑ��:�UdP��I|9!�I��4��ߐ����[�*�=!�J��:LP�ɲ,w�=.��5V��^�q�"�z|���c���oI�3�c:��$	TR����wJ��9���ʐo���ԣ+��d+x`��;�������;\���;�?� �8B�]r�8>Z�1A���1T�M�0q�Ձ��Qk����?�������P���]�n`�/�Pe�΢�R]!��J�PS�`����b�q���[����ݛ�x�US�*]���lV3�ʮt����XZT����h+�����IۊQY��W䚟ڧWs���#^�U�4SLn�iŅ`�C���I����d�[I�ô���0�����8�;�hB W?}C*�0P���꒐���T������u?�͂�ظ�
#�%d���<I�:Rʓc_�0��sM$l�F
�]�Db�P�����ؕ��01�^'pr������	[e@g�
x(�Egs��옕��YZco�r����D��I�0J
PHt�����e1<F��Ip�xO�$:G�Q1��N�:;����Ǡ�1[WWƉI����F�]�~��J1�!DN0��u	�\E�.1��D���M��I��Iy��uLi���9���s���DL��<�HwZ�������_L�^{�>0_�k�ZĆR������#�*���l78�\"�y�a�6֮��XH�л�k1�\^24��*S�(��b"��U�v�/r��e�?�퇥l_� �4�3/I,�J�ui����Hæ�zΙt��RI����ܿ�b�r�n���b��IÒ��]� �
b6��0�ѐ �Ŵ���	���L(�D�0���ZI4s�\����i�cWPJ�$Q���_y��*c!�n����) cp�[(�>��{u
��./�͘d��$	���{�
D���E���(�)X���ʶ��A�ी�b�t�!T'�ߚ<P �����h 'R.I�.%�x�@�< c	J�(]酢�����kKP���﷔݁�1��!�G"�J� ���V.A��m��l��sIi$n}�X����\�᠗(Ћ_�Aɯ���>������Ԫc�����O=LX�:Ih1������D|/\f�6n�|�V`-�o�bN��*��4t�F�u;�N.v�ό�W6?^�#v��`�(Z���g�0��̥�ke���
�l�k/��%�\-��:�� mcf�
 ,u�G 늣��F+6d����(\!����[e��]���6�D�f�@�7E��(����`��w��� ��b)ь��DR$�E�I���Jb���/�FLK� `R%�/U$��RE�W$@��&���e(�� �M�,�����}�b�Sc �!�F���tUr�"��C��r�g�����>���Y�<�K0?��0y�O��-� ���!Av�I'sj�!����_ai&F�:�;={��16��0Ȯ�L_�Q�6w�
4Z1�$\�S�Hs%����K�^�.1�h�t��RE(U$$�REEB(UU$�R �� :�a� �fVa)b�b�!f��fC�f*e��*��B5+0E-�Z,l�~�_LaI�
 PL����K5�(u�=�7`d�-y�x܀Y\�q��>�l �,(A:������������Hc��`�"�C�Lt�P^H��҃���T�����1@7��|�w8C���X��y_T"��Be�k,�
I��7�$AO��vȇ�ȼp�	b&�0F"�Ưk����@���* �($F-�@���%<k��|�Auu�}&�����a"��W��!*�
Б�'�W��Fy��>ɨ���YQ78�i�y��}�A�Z���>��A�X���!��gN^�������|�/T̀�\�+!��5�5 S�,�&4��U]X�7����=ӽ�a��X��]X�CI�Щ?Aŗ��c��*��N����_'"䎆�y@,����	�*�L�_��cn] C3. ^�*C4ïJ�4TӺSMzP�C9��:��RP��.����l#�L��y]P��B�;�7�>Eĝ�7a>}����n�4�<��-I�^Dz`#/����ܯ�*30����MZ�[n(��)@m� :?�.6P�1z3����I�f�L�}�H4Qظ����������	�	f�d��C��.��Ig��ȑSW�dz�֌S����#�L����̿�d�) 7E���PD�2�(c{�0?������Q��3�:�>Fv�5x�Z8Ը�RxX�YA�}�70�O� zX�bҳ���� ?�$D?�H��M50�.	΋N=-e�",����I�Q/�~�ݡ�P�.IU��y���6�D��H��#����jul��F����G���;@��,�z�h�M���zr���/w
��ú���o@��/R��uAD���(+����i{��ʌ!��v�$n��	:?��<{�|c�G�����/����c q��%�(��nx	�O���}�o2�s���k��0�~U�oQ���-�!�ĐC��� ��������}n���u5��a�I��X�?!�f<�kH�����^Ӂ,g��ե��t�r��������`����.�9(	*��P����DH$%��5?˙(5O��,L�+�d�ml��H�!��H�(�ꆿ���6��1\p8m#Q���������m#�󬗐pخ��W��rCVW��<�L�p�T+�F�za /T�GB&叺�����}'����^ 跥0A�����"
��r��ChQ�]���},1�=�r
s�@�(�V�2�7�gv�9�X��s�_�~�w{����E�m�h���<
��� �Fd/$�]��u#�ԡ�ڌ�� �R8'0^:���$�D �1�.y3N_�̸�|��|�S�R��*6��Nf����g��,��M�cQ�jx�)")�@��F"�a.ã;�B�� 	��� �X�EK*\]AU�DW��"*OBZ�1'�3H	�����+�!�ˈ��(�%�6\j��&Z�;�+!C0`�TD"AM+�l��l����++�_0@Z$�I�J"~tpA�����$@!���Xtq��&j�f���\�HE�!�,bƉ(��9S�;�]3A,��Z
��ښ�Z�10��b�� ۋ�5�{��9�zK�>&ֈ9vb<ܘ�V� G&�=
`�y"�����vAEƳ�0r�@E�3{0r@El;�U"S���<%��a�*㛨[�eL!� �\�D���$Mﭡ[�FiM�- �1��� �B*��FN8R��
��
.0o��].���. F���K�%b��\����� 
W	i�+�k�Өc��DH�Pq�e���.�t �Z�W�+e'�H�9�������G�H�\V�-`�����%F̰�ga���7w��@�{�R
�4Z�k8�;�/�a�}���ֈ�΁���B�>WI1n����E��hQ�� s��4�GS�UI���ĭŔ]�(��2H\鲐��sut�cv�p\/~�/%a����)�D���ϛ�d�����Vq�,ź%�2��ĭ�@��,xc���RIx�k��؏X�Yu6��7���KAJb>����Υ���K���P���n� |��$3/6�F�K
��M�f)oq=���[9�J�İ1�6C9`E_~����hAzC� 3��	�c�~X?�_�m&2u���	0b�d��P44�9�\��2�ž"#"�.*�y�#�lP�ۗe��c�������Z�(`�/Y$�9ڧ[U��3��*CqV"@�߷_nVp�EŔ�~�#��|c����r�!C��2(�VE�A�Sx��Z�[�{���N
��_���t�h�����^lDа�$x?+%f�	X���^��"1�i��#�R~�ܔ��P?�`����������gXT��(
�B�:��榒6�lx�O������+�;�$�ً}'10ɻ�j�*<�,�ܚ9%�?�p������"�+1�@`�P�6%|�D(���{Xͱ��r�����JOo�n4`b���I~t��������{��:�@4Ƒl��S`3i8�R� J�0�X�z�����+�@�PC���Q�b��9�k�U�� �ӟ��������:�� �X��K��eh/�e�:w�.���BjPqH]i�2R�$�G:��tuE����<8��_w5-)��$�*����{�}�k�/�AW�yN?����%���#�N�ø�0�4���M�t@!V@0v(v�_WV�B,_y)�T�Q�-�����u��XU�ןgy4�T-�F�!����M�ZhEË��gr�?��6�;2���Űބ��pfF��+5t���'ғ�P�������b_���a�H�*�e�f���Vj��������ce|�Y���r�KQt��JK�x��0�a��j+��.F�.v�y/uf;Y���a���
�&�r%������-,������E*��Z��w?�Y���FY��)�p�(�K��:�%qЖupQ���䩌f+�(��n�Z�ߝR�_a|v�*]��ETlu*�)��nұ��hPL�8���b� Rm!'j�Z�[��7ű������~�͘��� �<N00���������{�	W\ƅ����G$Q��K��@w9�:	��V�����B��]����"�ax��_d���w^��2T�bO��+�V�M���u����r���a��H�³	඿��4��y�8�76TC.����2�����.��E���H�]qGX*a��.SX��ܱ���Qب��)��dF]��u&�x�d�$RwM�\ڵ�����#�ϟ�]�v���Ơ62Zȸ�gSX�z>����"�vC����*�/2&�xdl� x��|V^����ML�dT��zh�B�T[%�ud�:���<$3�]�)zIF\|���P���e#�,���ԐJ�w��ZN�Wr]^��0����`�]�t���:]���&+%��"��~�ɲI�d�,z�a������HIY����\y����S�W�z�I6mZ�Q�7��L,>���*��Y|?�,%���K���Xъ�[J��_��i+G��~�hוu��ax+��:��T�9/�|!�R�����SaǄ��
�Ll �:=8�6�H�<�bD�
�/D��U�������/�i�ΐyRԧ��)O�n��ϿD���7�Pn��P���`���B��	���à�a�0b�qߪu��`(A��-%�A��ȑʆ�݋���h�`|1�0��v�HeS�^�����;
q��G*�QX%
���#G��N2��dQ�q�h�2�k>Y�S?ɋ/mF�$D�"�>u��5�}�v��+��汘YQ�n;d]�]A�P/�/�y���V ��[
r���B_W#��ήWL6��-�*[�*�������⤻'����-���`��j�eU�Q��F�R�U�A�S��WG�@� ��.z+%��\�RˤK��8�>��PQ�R�#�8/NX����UJ@��Lʧx���=��8_q8�]%6x�Nm�N?'	���_��.`X��H�kAs�#�?vT1<?��X\L��q>0B���c�c��/TeAة�Vsj���8�'��#�hPM��.��x��G�%�s�p,.�"��
�qS�蠯7N�>Ŧ���G �+q��a������I�<���>�7k�0y�S�xB��p
I4�X�����	�V&�H�rj�肎A��X�A0�+
�-�~C�C��{1��5Sz���rߎ>���Bg�f�쏄�Ť��M�|Ͳ��Li�<s���Pkcv"�.r�c"�V�U��z�T�x�0�8�@-��Q1���!T�L:���g~���lT�z�����u .8��Ӂ1�s����k��X��?i|p�D|�i���� �Eo�n+�� Y*��P���[-�����8�B�X#S<���C�Y�|��]e	�_�QWapgE=�^���M;�\%�z�@���D�k�.e$�C$]�U�\2�
p�6�1+ѳ�9�{�;0�&UA\�K�Z7��D ��F��ZK�˫k׮]��1Kon�Ѽ�!(>�3�����|�<?oYm�|��\��8ty[N�%\��4�aPM��S���hU�B?5=	��
��$�:��}g�9K��4)��H/+��B#���ʋY�������F# ~�r�BaY��)%�J��P�"�e�N��s�E*��J�w��q������L�υ��Ѵ�g���6��H������<�n�GQ��"��F��|�S���M����^�r({��+��[�>��tƔ9p$�LL�#�F��� �Ģ4=զ�D��ml�\�;1��k��`1���I��\T��D��"���g�0G4 �ݺ!��=9Hu�v���s]�hܰ�R�'�h�Z����=�����s[�.8��9L���`*��>�G���Z��Yb��	��ߨgGu&	]���}I�m�8ўP���@���
��R�V8]��xO�k�A�n����T���̊����@C��H�(�g�
Dq��
ǎ �;�Fb}N��n�˹�.�$�
��H�,��A|pg#���_� 
�8��c�s~1�T�����a�`��墇�b���>0����8v�� ���g��[���ye�KMYV�gqT�_���$�1]C�t4�=�-���r]�<+Q�:,(�F��@B�s��|�b�x3<�Q'�V���3[�~���Ѐ���M8!f{an�.�L/K@��S��Ѵs�r�
(��\�
��1<(g���e�*��i�YY�V���(f^0��C3@3u���[��fi;@���b�'�*u�ٙ�
Jj�,����� �Ka]	>�je׿��V꼥,ݫ	����>,���J��~	^О�;���nK��&|IȪr��ŗ�?��|��G
1��Ơ�u� �����@�X��`�TqZ/m��Q���S�WL)}sr�A�_�?�ᇬ$p �!��Ɣ���3ń�3�> ��(��i����>2� ���}՜(pg���p&�9���ŔM�c�:��?q�@��z����I����?��bU���T% #v�C�!�Eq���W��'�� D�:��YR�G�"݊��Y�@
��^@�,�Q`����(r?�@H����Jdr�Q�ͱ1��"�&
����.X<��l�J�%��C����7V���#?��:��C�,�A��T:-�[��Q ��	�4���7@R�]�?��bux��P�v�e͂E,;2��a��/#TRƲB��\��~a�:��2��/9����q||++m�KYf�z+��gR>��J��pq�z"`̗p�7B���0F�.T�Q�Ri��X/�"X���"
�'%����2HN�r�;�>	N���N���u~�0̕"9ܽ�N�7piL���w�§���<�v�ҥCTJ�v����،"w�}
�dBK�����4K�Pi��T�n1�j BV�1���q@C��Zظ�3��� �E��/b���}N��e�s�X���y@����l,Rݫos�
�a���w'/&Z�3�� H�//�ܜ��"�Kc�_QE��=gf�#�)�`���w!X�a�j��'Q/�v�Ү2#�5��!���c���b�N�����!��]�N2�����?D�D�a�]%o&9|�ٕ���z*������}Ƅ��}�|!��%pBC��)�� ��J�ҳ8(�S=Ŵ�E%1�d=I�Pt�af5�3�q`�lB4��o���&3�����Ca= ]��W��!��B�Շ�4���3px3+�>��ܖ-���L }&�F�j{�/�s��������HϐZ���+ ����"����ϟ���/��@��mB�����y����� WxǡJ�L�.�W.�Uq �\�0�և�!XҢ�s�W�@�⹋z���(j�� 5��z% Ɯ�.1'`2XS�3+�!�4@��`�
{_�{a؆��O-&���SǸ���0 �PB�J���k~f 	�.	`CYcH�.�"OR�U��K��3g�襞���8�;)�����`����a@P����6�:xg��T�Ё���f�֢��5m,ac`�z|1iC�{faטr_Hkfxe��%K�/����_M,ܶ؛5~��7����Ji��X�;%��b����g،C�}Kqĕ�D���@UPg	����oW�L�ex�arW��˪/��iQ�ּO��F����dp�sX��0�Lr��c=��G2zմ�(�m��wL7ب���)�Җ��Q!�`�;0n<wz�.�b&jr��C����MU���:`�ϩ3n�*$���K�=�Z����R��T�(�O����AWsP�Y~=���^=�(����)-�G�7�����L��DT��tI߃b�Q��>l��&L=P����~J�1I�ӓF5A�$����>�%�G���CI9����b�wKV̿�� @=��Է��%���KPBH�Z�(Ƴ�����d䏍1Ѻ2x�l�� ���Y%�=�x��Qu5��ր�eEȢϲz`5�\a�`�fp=Wc2�>X���zj�옃C����U�2if��2E(ɱ��!0s��2����3W�?����;�B˕`.
R_�0%����-=g-7)q
ABe$^��ڲ�2��XVS�m�ȼ� ��$ƨ�m/SӺ�g9�"��a�����4�WAgv*��EӺ_��@_�zۄiU'@�Bv�|���W����+ �L����1��ץ��ڭ_�P�t�F�u������j��K���zu>0�{5��l]�y$��@|+���Ҙe����C�n�D���(HY1P�����t�H&���ǉ�h@F�f���mG<��/��(�Eprb		d,|\
�(7��^=�)�$��	�C��}�=����T��e�����)�f�.���ܲ�}
�w����zu�*�HC��Ki@���)����6G'�=�16�C]���썀�;��$�Y�
�Y���/�TӘ�7Rm݌�[�y_��q)`��?0�`g�o�&T���byG�>P�1MU�h�(�N �Ѣ,Q
����`aTʩ�>`�¦�**yB�3�Ԑ���(�D&)#(6y$B:��=��9�%x�0A�T.br��fd��)O��l�z5��P�C�Шe#7	�%q������p9�y��:��B��D��`������Z=��2΢�K��4�膕U���:���L.�ayd�
B�cI��B�u3�Z��I��pY�t��A +��ud8P؅i \�n�e�+�0���Z�t((��f@a~�T���Idg$C�+��\)TZ�+�HB2�:- ��qUT���������I�WJ�!��,v���P~�kW��Fbe�I�FWmX��[�ڠo��^�����nan��y3����3�A���Y�-pUc�^6�%Q� �p43��.,x\��V�� �6�<3s��D$��Vw���"��;(���SE]�� �3��S+W9A�����ɻ�s���i�ƍ����h@C��D8�*�~ȟ��Ǥ���)�U�p���WP$[�aW����`�Q;��.�ZRvv�uS炾�0��OW��@��s����Ae�
�G ^ic�}`�  ��L���&��©"0��V
51}�ê\�H����Ģ�����:�^b�����L��<���wz]e�@�:�D�""�$��X��/��Ԉ�/�0Pn�#��O_�nH��T]b&��>&i��6��w��q1AD�hb/Dy�� WcX���t��p��F�*��U��ћ��B��H!@A\��vb�)[�	���M�ƀ%N_�%��8�0;,Q�-�1!������2��`VM�F��r1�����щA���&G'C�O-�܅�Ȱ!�b5/9�p�5��0|8�`�[����?�Tg �jB��`?����l1�?(�6�����$����� X[x5K65-���x�UYL��	�����N9�"S �c��>�qEq��O��P�@B���Y��:E�m��F/�3q"Ot�����S��\�0��~�E�gd���� +��s��Ɋ�z.�L�����~b��_�d�h��%��粟r(�l?F�}�����]=��-/�[7�c�
�T�̯�+!����s�@�~}*D"���sА6Kr?>�6W�^�ۣHE�����!�R���{�N��y0S�c�*�����x��Q[�#��0�M*"\&���Hɍ�h=rq�"�u�߭�U�93��������?��3����0���ϰ�u+�Zo��_��^������­T����pP�2ة�|����yT*lEH������J
�]{nNb�3=���d���>��^8C�o�q��V����%6�Bѳn@�3[02�d7��HbZ��d&oH !��UQ�K����
#`E�J!'�� ��ɺ���A��ppL�8��#	ݹ�bv&|?!1[�^1���zN7�T8��E����nl���̈́�*�E"Ӊ�K�?��d���_���"hA�ƈ5r|۵�;�	������Iq�'Ί�А6C�*�Ӭ�q��[�mPU	#?���1�{|)۔"��d�8Z`ax1`�*0M�^sA4��� /a�#vE��a�vW�����o��/r�1BA�B<F�pǭ��ʹ��U
&(b/�}���цKC�<i���Z�A&�@���d ?2�p8��~|x>�S�S�B«��+�B�F.7տ��nx�Ǐ<�#��|���x�����C��"!u=����I W������q���t�\��d'|��2CPJB�Y 1�A�3Jj�e�Q�9كN����7��kJ�&�~_=4����﨓�1�L���u����:է�n�5���R]�Η�+,��Ͼ:~��)�	<-�5�}`6E#x(�����<e�U�����$�QH�"�q.c��?�iJ"�$#�$�g[�~
2n��S2�	$,��:_	�
>T;F(����?8C�E<%�e� &�+�Oϱ1}�ڐ�@�E �4U̵.@i2bSĸԑijE($���,##���٠ BB��f`�a��R]ê�&���ol�Б�Í;��T@B-�T�E����[쪧\--R2ܰҥ�L�
�,�"0Gdv����+��\�۩Hv���%�,���+9w!��S�-�.3ȑ˸���]��@�9��a���;�e�����r��q��,�E�C�:�CI�	PƑsN,��!�U�ȩ%��=���S6�sT�.�>�\�'_�K��} �v\���$���/Ɛ�Czki�Ԃ�2�� �!ҭ4%#H�����T�k����u�)@"0�p4b��z��6���Q�	M�&�aJ�|�À��r�4�a��@�Kn?!������t�;?�%�H�d��(XJ(�3��MϗE�����q.��y=�����$0;�	Z��	\�;	�:Y1��*��ڳ+�?�F����+`�%�c�U�5s:^}�M0�)�0�H qH8�Z����Hd�!�3jj��+����e���b�̾��	�.�bi_�ol 5A5���W\�}�!݅'ڐ�^�G��#h8~�&?ʰ�����s���w��X�%h��r��d�V�A�e�9��$�	�{#1T��Q)�5s}P��z�/#{L�w*��]�A�)���@.��I�݇�ݛ+-f끧���ʕ��U�@�P\g9�J��D�x �)��T	B����+RF���CD�������!���!C"�	A��)�Kc�_ f�~�@j�����iva��`��篤B�#j_)���;;�cx��.�9����S#�������6��*`��a�=\@�R
r�ㅌ�A��!:�G?;��v�_3���.��h�����	�a�<ߝL�.��Ĩ�t�֋��1�$�Eu��[��\MGj$.���!�	�\u�1�0���V��p�_,��W2�p��=�2��8f�D F-"��B�p:�4�� �s=�
ը�H���h���Ep~�_4��R�R�bFwyF:�5��0��l���BPMUM�=�d֙|�y�d��3��nlɜ�t�s0ù���䯯���b�@��SJ
��d`�e F%�?���<۱
1F�d���J�r;hѠҚPS^.pc���Z�駬ڜ�I�(h4*s����R,88/l1�&�b��s��2vp��p��=PQx�r��xtL"�ƇΝ�;a��g�Ywy�`�A�R_ot(t.R܇���AD���p+�R��ǩ̂��H�tCG݅��fz߹��,����� DePyM
�&�R�<CK8X��[�YUd�HÙ�qLD[�p�
�Fє�g4�#�����Y����31�nf�=L�Ye%n��$A����U�
������x��!x�oc�$���Wj0�@ķ��`��EA�S2�q��H4VU�\�.0�K�gA�P��y:�څ_Ynd�N���II`��_م'l�'?#��Uc�@H�4��=��)��~wd�K��X�N���\����l�&=�ۤ��]q/���!�����+���V̇�(��1K	D������A�>�i�-��;��%�dc�fuK,�j,�u�	���&�_?'Wr��_�D>�C�`�#Q	�Ո�CSɸ�3�-ƣK[K �(f���C��(gt�X�
D��L�A���ZNX 	L�)9��R&�0�	2E%��O�fj���
��GF����!�[@��a��it؀�X��_<ܷ�����c;�sQ�x��%���V�	3�`�"äh#�w�U"��B� �'oc�3�b��Y"���G�W�'M���8�B���W�X�(�/P�l�ɵ�G�c�$�&�9��������@��� �(�O]�QlZ����JQ|�)���<17p� =��x^cdx�� b��b���o��n�(V�UU�xe���H���!�(@���IJ���	�����s�}_���u�� -%���E����������3�3$f�����E��!�$3���N��e�z*�H#)A��咀�ڝ��"h�uuu*���)�Y@��Hw+XźS&���Y����E�3� 8; }Q0h�x��̕�%��"eH���p#�v8��B>�<��`%�'J	a�݅|���ߑ{�����࿃�]�]B��ǻ�R�sJ@h7��j�`�`��Ȩ�&�N���H�"�GXwQ�ژ��~�;�֙iQ��,�E�8�cFP�M���E=E�n1Y�XPѫ��ӏ'�����U�RC�~Q����N��5���Ǿș |�� ]`�0��������hP��T��y�u�Ŭ�H��C*ffYt��[mQ�p�Rchq��g���_7$�������HK6�'�V��
��U�̟�W���k�B�f@J�:�ER��)��w�EWiu?���tF��~%<[QB�@<�˜QTH6��m$Ҍ�U;����*XRø���,,�T����rH��A9jϗ�NP�LPoA���j+����L@ Ӛ�;���@�85�R���(ю�B́t��I�����_0|`G�@ �0��̩�_Ԭ�Q
�k}��_�V͙�5,Z��ƄJ�`��q��]���;3Hq�O�������q)��� J�UfѬ�XJ��L�4�j�JYP��hT� 
5%z�m�d!i q�G�}H�7 !	0,�@x�4�!���_��;Č�46��Krǝ5��p��9���$��ܩ�`��#��}#�&�`&}=��%����L���o�)9�4��ȡ�����n(m!;	S����.�]!]8�Aom�t��6LH``c:bH�m���B�&����~T�6���qjfe����]^��/��dA(Z�Q��d��_�;[hJ��@��/���#��5(
���W.�YX&����u|P ͆C��}�Lz�`gS�%ݬ��g�j_d`��u�|��t�`n����K+b1����'���q��&P�c��W{�:�n2����v nx*e������wDqr�r*�907��(Ј� �N8w�>D�"��qɥ��c�.�R~��߹�,�Z,�)�H��
:$2����>�7��L���1�	��g'4Į�g� p;�x����9�Pִ��Y��J��V�i�ß�@���8TH=#�AR>� ��P>�>��ss#ȝq�u�����(����Wm!�
X�c�Zp`��'�J�a�	r�u��.��T�$C.sE�,(�z����K	P��~~$���ȗ�������2(�o@��.F
��	��o
 2* 
�$[c�]�xPC9���'9d5�;|�|����yĘc�,`��>�2�1dj�o^�9�B��8���}CEuƪ��Z�V�)V`4��V��@��V��@�wqc��ʾ�������NvB�<��C6�΃���Ea`�(*F&c�):Ҝa�e��l>�ڦjL��b^��b����5h?!�*qp�큪^�@+�ّ,$_Y�ؗ+D�8����\yMy��	�"jnwY7~�e�4���~�pV�~�9VzB+��+���ey\1��e!R�f�L� D�":w�(��(9:cI�*���	,���=� ��F��N��
�������/�ʝ+�U~�.���93Nyg]%h���|陷�fG��6m�`�Y�Нs#������s��D��E��.��eڲ�9j�aG������T׀/�C�
���A�d 0��g��~?�l:z�X�(���_����H�2���:Vb�?����^?:�򫊗�Uc��/�H/�5I�� ��>!hԞ�oF�#��uJ�F`�"�S$��B�r��&��v��������j��T?ݻ���G�
�##�7Š����]\!���~~��OF��m��+ջ�d~�MN2���N��c�o��)U���a�šp�4s�Er�d h�0XFi"w��Y����G3�p3	ҵ;�T��+��Ŭ���S	�;�8þ�թ�u	�؞��_�ש� �Q���n"�8a���}Z>si��|~���At*{��dd4�hi�A�TǕ�.VY����:��0q:�LK�������UGi1���6������F��2�I��L� I4h_$-�
[E	L��w��00�$ү�@�j���<�`�������\��¹���|]^1H���*]��~iϛ���G	/����;�T�܋��sh��]icO�~{���ψx�04�!)�o���ZL����ը��t�T7��Hl4*�X�t)b+���sd�!o'���%Ǯ�J��@`�oSe6���*�Z�(�1v�E�b0	���z6U��ϦRǒy�\�������ԋ�s���R�qXS�!�B�I�t���+�)�
�,;���3(���C#��L�P�)�FOY ��S'~K��3�eH=b�y��$+f�_���e��sؖ��&Ǝ�yδ�g�c4�~d���3D4��������xc9��-J��N�k��m}c]�3l�;8L���q���;�e�D���!U�"�(`]3E�5��%� k�t,ӛV�]���(�v�K ��(�$��3�~%yDb�xse�m	S:iD B�y�@��)�&�n��1��(B��+���\�b�(u E�4�*����bcK��U�ƌhpy.Ya;��/]�L�¥N�?��Ak:��e�Y�v}�l��B�bJT�����M���:��KҘx[̗�ԈI��"�G^&�f�~�,�p,b�ͤ���5�(��QI�N#��2,�9�.�V�� d�PQ'+��@��^S2ij!C
�>Q>�0�y�_<���U,/J�����>T���(���٭��k�U��r֮�P8�X{9Ɛ��Ȇ�|Y4��z��(����f�i<E���芫4VO1t{�5�$S���~����} Օ�v�4Lge���`�?��Z�N��u�Q�]�v�_T*¹�L�bo�
w4 =w���";���O�Q�gG��#�7&Q���H����-ݫ���U<��?��_R�-������4�`���ꖿ�k�=zCx5-d�[��,��Ы�&���kLd�/|�!{L�M�*�*��8^G���ψfIo�}���Y�a�f�t�)�#=V0Z+��d�K�BW��@�[E�v�f�#�������)x}�S���
9б�����M�dC\V�I�������wZL��Ó���r��GVb���� Ϫ�W�����|��'��g�_3M�b�j<��`�508����n
Lȱ�9?%����2룮��nD4iM5���4zY���M�K�0�®�|���fS�l!B�4i�J�vi��*�gZ���Pe	ʠO�R-c]���;غ"������,�u|��"�Kp��<-ӡ��S�D����p���bL��+\��H�'��x��SdS�L+4�:ʌ~�r!���´r�٪R�*��G`��.,nYcX3Y�W#m^�8�b�!���<��Y�1Dc�Hg`�2� ��̽b�,Ħ�-A�SW��5n�;�a�@k�JT
��&���a�jm\ :U�b�W��g�aS}ڱӵE&պúc`PrdnG�^����@�p�*����$�u���	C!�ORyx^�| ċ�U��U1����E�y맷�n���(�p�b�XΤ��q.'`�[_Ih�+�"�6<fl��#�X`�1��
�h�:�L*�<�!�(���#.
�]����Dۙr}��)d�� o��0�[\�#T�j���A:�	 �4��W�����c@Q�b�}q�@��ɷ���\	�x�\�B��	�H7,�X�[�L�[y+��,��Ur��b6Ϊ�~81�rT�Vmyݤ�@�i���c���K?�X~&�R�b���Ԃ�iB���#(
���f���� 2�_ܾh���3�7�B�A<��9@���*�n����N��0k]اҬ9)p�K��:g$��@�[����N���@j.�~c�Sl��]�/01/���H�L5� ��H�<R�C-�Ν�d���!�J�t����ئb�/�0R|V�;݂ȥTE�g#�+�_qW�W�q·���H�����P��+�?׳���Z��<��b�	���!:�C��y0\�x�����m��
|P���#��#P�m�2FSqۋp'<�R���S(ω/��N��%I
_�0���
��#��9TD9HRJZ�ڕ�*j �q��/+?����*� ���á1�As	� h�Rf{G������7~LU�����ݫ{"�*�e���L�v:�I�%0�O��)��	C�GJ��� ?3#��ǀ�ُ���u�ٙo>�J���2�BM�g.��P��>�N��!��t������S�^�Zhϔ�Z-|��ͺL)�!�f@��1�%�hc��HM���J��N����"�]�� l)�"h��\B0@<8j1����i*�/�V�{>�1x�����4�ĎQW����	b��
ML� ��������(a�C���D[�0ht����/P���e\���
��;�F��	Ϫ�FU��Y ��yˤ|Uy}�z���H KD?D@��N�gt�R fn�����lP^�b#�@v6�m��U�c���%���*&�V�{I��x�n�6�A���a]$� �&�/��L�z��n��>�Aň_V��֓�J+*s}�N��?�̣�	+Mw�.� TDL,�zuĹ����P�Z
f"*�����U�$cV�(�2Vy̢�4`J����Y���Y7X�n:�3�!V`�$BB�aa��)�-��n`bL���$�ݴ)�b̝H���IsPf�N��*�J���Rx�;�Ϩ �����8�+Rj�e�1��(Ŀ=��RG���M��C^i`�H@˴!Q?�  sd�$�9�6�>��Կ��Y[�.DWP�Tb�bqg^�/��̽�� ?�qI2�rh��Hc�����M�*�0������]/��i�
y�Vqd\��-bB��}d���-6�-�
Sxm�Q�&F���xE�xl��i�s5�����V�r�1�uvBKWY�hE�z��-��xt?4OK�ѯ(��n�PqO&�F�y��;�����������g �b��WX�D�g?��u8C�u�
����=���|1t������$Sé�y:e�@�G�����1^�94jd�__G�"�� *䋚V� ��+,�r���rnȔ���gs�nR��\�R�h�"�#���^AV{�va�s�熒	�@a����ĨA{"��:�b6����kRMC���I)�.�D�����8��z
����U��MHl�P �ה�|I/�V#IJ�=��I��pbS���v����J��uS�QC
t2/(I}7��W��%V�j����T��OI�����]�b߱.�Q��0V�¦���L�tݘ���aϿJ1P�f�>��+h�֪͖����t�ӎ�;�;M}�,��!q��cɇ̤��2��K?��i����l���~��y6�}0�7��������c^N��k7�#�V�����V�^�^��1G��ZZ�Yi�K�.�;�Bܥ��KLL�����p�����i���F	F�~��_VU�Ql*(�����C���	+����Ĭ:�������i���=���1s�@�Jf�G�d�(��(�*��9MDN�����C�S�v�ի �� ��z%��yE�`2���{d�y5����&!^_HYN�uR�(����_熭��<f�>��HfP��Rt��S����߯i��!���;��o�t��
��]@�"�g;cq���Zmۢe��^�W�@�Ϯ��q��ʁ�����.�^�yUL|��Y�OF� fGZ �\%��&w1m�)U�rc":�+>�|픀����eO�*�FX=Z�PqX�����)�2�b�\��ji<uut"���گ7S4��cZ�67گ�U�=�Z7m||��W�.Ø0Jc�B�Ǐgn�N�YHw��2��sFNU�9_q�m�L,(fq�o��p<���?��k��	�/Ī�>F����p@�*��q$tLl*$r����nF�����ڏL� �R����]��5zڃ��T?���$(��[��ݫ�z�|1��y0����:^�3c�\�+ )��}�I^e�]L�F���|Lf�ʷR�oZq����H+Nܗ�g	Z�h�C5�,ݠT�aa�v���6�����qwbJ�L��lX�#? �J�Ƀ��v��1�u���}=&�F�_*lB�q�JW�h�4gnw�f�������+�*mk�a�	�q��B�\K
܈��D���� � ��%!.3�3?�Lza߲+mlU�Z��1P��J��|�+^�!��7�a�M�z�^C�LC�9�����!m`�P��	����K �t��R�/"/
�+$�\�~�7�^Y�v�~Y/��ԩ�Ӧ�t~�zB���1��Yƌs�I�c�"|��MS����S�z��A
n��'���x8`O�Y�=������?��j�>���9V�6P��sǙ|-r���m��)���4���qc|�]xM;i�Q�D����E�gr�^� �R�Hx��Qt����*�2���C�.❯_i0��<��<Y֥­a���5�qP�_<ܕ���7�����F�h�>K\b V�F�0�\LP/
x�>���%�@�N�_�"J���%SJ_�D��J�T)1;fی���8�+�ޅ�>�X�]� �!%�S	2��T��K�e�'�IHR@R4�V1��CYG����V<�a���Zu��_P9�\�:�H��|���OuYT��%��G�'��G�e�g�꿁��U��h�;�*��x+_�Y��;"�:���ϛ�%�*�~���v� �DK	��>�����e���;�Q�LP;�PF�\謫P��E��P$r<�
�e�Ѿ;`g����^G�5���QՐd�r����Iee\�8zq��0F�#���ӌ����he�Z8�1ȆG%��n���T��wҲ��lhHIh�Q°�3�*!z;[�$Du
�8���ڥ�����V�����!/^E�oܮB��o�Eǈ��D�b4.��}C7kz����ih`X�5���*�i�4s�����0סq5̩��bMHX?_O���9)Il�p%
�G�{v�����M��M��{���$F$2�D�{��b&���g��A+�}̳�YD�rl�;	}�"4J�w�/ң4�*�{bC�9�۪��1�QGv���8bN��4�_�&ݝi��n�����w��CZ��^���x�d&���m��A"Pk�koԼc>�_h���B�������:<}����-T���j�:��U3S"��X�ɦ�W���o���+ry8�c��5���H,ڗP�'�ݏ8�Z5'���u�L�H�fЉ���*��i�V�&�������+�t������b
bSm�%�/�۱�ٷs$S}1R�B�FF�����M�ޙN���殨j11=��`LET��ؕa�_�@{-���tbR��o��X_��J���![�A����W���������/�83�>U1Q�� �R�WY��h�;2M��b���oT}�8_��M�]O������р�f�z�r@u)$PV ���HT�;��gҿ�#�̫��Pj�]�����b�H��Ew �C�+#l�%X&����ϒ�JZ(F����6�_LBl�Ф[���c�G8�����j���r5h�K�ŌO����R��֫ b?]��(�I��%��cK$3��C��zA�� &���z*2�N({�|̋��"��.6+l_<[\\^A�7����(�'������)����`��E���%�����%�lsU a�4K�ǌ{<$@a寋�+�s���.�L�] �C ^?M�D�_|���teX3I"�_U:.$<X¼�Y�s��N��Y� Ka��-�)Ɣዹ�ɓ.%�|��Y�����JW&�fZ5�$�ϽZ��']Y�9<p�]ƍ��J|"�w':/�ئ��"���l�q�>�@�	\�*ik�f��ɸ 4j�[	�6��%�^��52K�Y��ůűq�&Ta�@n7A��%��
��91�m��s\��R���i@������87�!���
��z;��ߕ���j7�?[��E_�v4UlSK�担�͝LM��<ZY���/��,z��AZ�.n��w�Q��c�ɺ����p�&H@���a�*��+��eQ���R3�z�������u Eg>t
د��(�= 
aJ�f���\��uNn����e�:(�0!}dI�]	*�Tq3��,g���Sa(���Bs�AU�M��1���E1���NU���kW�\b2�'�$T�Yc�����P1Q��A��X��# ����A1B��Ј�Q�Ն��.*]�NT����rA')�B T�V�U0h01�U�fl�̞�@.:��!���th�ŗ��b�r��"$iҍ�|�N�Đ.ĝ6���|k I�Ֆw4�I�ڰV�����7�"m�!��/\U��zwz�|^����]�kY��u�u	L����z�>�Y�R�����Ќ��)���$��}kQ��9�.�
c��W���#�WG�mʫ�Kj�	(��΂�;YDe������1P��l:���H�g��tT���
q�W@t�΃&NUxfi�c�\O�y/ZD�E�NT�UtOpsGaS=;��m�1� T1}�D@�C+�p��VU���Ep��u;���^_�.5��mH�OV!���+1�{20���W!��Pb	����$pH1V��������gO���L��|���'j�$1h��,W��0�&n��=�i?����`W�� aйNl���ƿ*�ڜw�T���5m�9����1:�ݮ��ޅP��:��Z�1eЃ¿���a�����2TE]��g����)=�^()�"(�xar��5%=��e	M��Q1��*P.z�Q��"i}S���7����'7 D�<���5�׆����SF$BF��+���KՊgc�������Թ��r�wyi�	�ʓ�%h���
�_�)�sUA5O�"�9E��TQy^y�d�UN~���a������f���w�QU"�\t�XP6*��$�����h꒬�L�{��
�$�u!��H>(�S#8�m�G_lu�H�|.�V��V��u������;+�da]�9���X)^��C���k��e�� ������~�b+Ē�"|�a��"f�%�cb�B#��3�$�QDL��|+7Sv�wJ��+	+�Gú��H���>Z H���N`X֫�
MĄ¬�[��A��Z��Y�K�>,�V��������?�X6��`�}���|�`Wy1���l�� ½���	�`6@H���t�ev�̻�����SX*Uq,  |_��<��:΍���K�+]��Wס+�;#�Xf�k�Bnx�B�AEFhH�X����s�C��HsC�S�]�]uHįR�s,.,B�dA E�|'P�����Đ��hc�+������`�b�|A�f��U�Q�~^�����xԥІd��)?Qw��i�)E��"�,��!����Ich�V;�<.��Ѿ��ɳh��AO\?Jd��<q)�'k1J�{]�@��a��e�����Ԙ���|е8*
"A���¥h$������juatn�$}��,��?����]�>0�Q�^5���|p�z��� ���S)[GٟI�l��������ue5��%�C
�:�����A��lE0�w���roh@1��'§+�x�}\O?��w�7|��=�����B��1�� S�Z�`�ɢ9�`b ��[a(�~�M#������@N�, �8	� ��/�?Px�I�#X�_8'@����`2���$�B�L��hπ�W�R
����B�2�uA"�bv�
'Z��Z�͹T,�U\���$v�c��%OU� �WƝ{Ղ��+��a2;���QJ��6^�A�9����&�9�:��C�t�/��b�0!�"��E��%3���sn$�-5v�3B���_��>�����;Un���"Ʋj�ubW����N�p�m��`�E�T*��k����$>:vy���A1��S@v|� �]���� �p��#�v��*k�G
ŘV�����I���t���blõ�)��+���UI��<c|H��2Z���HnP�m�
�1]�D�ӫ�����z�9a��LLIr�������xh�y�/���0���W�}�ǉ%2l,_L�\h��/��N|�Ҳ����
���A�C#����B�x�OuT/�������WZ@-�[
�Ry�D�;��`�5hX��L���4,��}t6ǁ�S^��#�-�j-����/��	$M`��lud���J2�Ճ��f�pZ����q.�|���)���H���j�R*G��^�@z_�	9c[]&�%g���i�
�Ů�$���z�������lW��j�Z������`��&�X_�X�����(D���FW;u"d��h��>#�}��b	��䘏���i$;?؀\V��*wZē�#�v�d"��IVb�GOD��WQ�#)d!�
��B�80�-kǷ��8(�盕��	Q��(F��O��Txbɠ�죖�E�!���>�qI���F��ew"����z��*#���q�^����������"����� n'���x����b���	��6W�]K�ê���&���2�:�#�ZJ2Դ(	D����~��K��$�LZnİ >%�;-��+fݰӭ�}n�~+i/rZָ�[�,�!f=� OI ������[͑�ω��E�.!��B�K2��C�Tw����[�˼����t�>���ξc����JU�dP�B.0��"���O��B�Q�R��rf�x�vtU��-I��F[>�j}*�.zpۊ��g���d�!%���yV�um��rū�Uy&y�
gf�f��4�N�xH��'�9�[@��Elw���o����9� �ޒ�ٗ��Z�����[��s!EbE�s}S������_5^%d��2�qb_�{���^w	W��"-,�2�R�q=�g<����s��V A55]Yp���"�5A+��\�N^&�������t%T��:�"Xm��h`ev�
�����E	&�J�\ƅX4��3_�"䊆����UV�@5F�B纷���&�W�c�j������.<�0���G�K��K�CrM.���%��*���#�4hI��K?����6�Z�71��	��F�?��*���X�L�3�K�ğ#zip1W~�aC��x����?u9_<̂�j�$0"6$A��������`,<������u���NDD�TTB�R�L��P�.�7�aR���E�Q+���Ud�?��~;�u�H��k��(�,O�
�l�F��_�XG�)袯�GL@����������`��V|g(_�@�)E�kt1��bѢҵ��j�B���;�����G
��~9����������	$B�.�Ghl�TX�X��+}��څN��������,�q�VԈ�_���K�����\'s`40��2��k�zV�T����}�R8NgK.�.�jU���W������b�'�KE�s%ݕ m�!sf�с=��~`�u~e��� %F/���
�`N#��QH����~��$�r1����`?&�-�rT �[�T�^9�ΐё��}�Q�+����u�K%a-�Ȉ=�yG��P�F�&���
�2PO�C��]"�N�S�c�	�JR���B%�(0��`v���_�D��T��%���P:��u�x*�L�N'��Ȧ[Q��<A��	]A����b@��A�t�
�{%0�c6��\X��O��
������/3~�@�]�n?�(�\�ƾ(��\"�}��B����
Д��!�$�5�.t���U�˒Ϥ�Da��W�H��i�3 ��U�*D)�R?���oRʹ�u��0�����u�"Q}"m<T/�i���1��T��`;�%u�gFP��k�r��,b�P�ʃ���3���9`
1RyκF�/�$m/V0h����e�o�{���!'�Z V�����k%yYC\�<F7�B���X΀�����aUw�8�8�BA� ��`�����w���tD�#� UA����}�(%�*�3���i�l?$0y���0ъc]C�� �y��\y#�|r�
W�'M���ҥ�Z����Ŗ'45നtUa�%ZE c��ԣ ������Hn����MS�ߧ�'5��#SJ������CU��!wY �EOI]��6^�#ua��)�)|^U�WAuǴ.�@ ��S���D:�DK����C`T�i��]��	��d9md����u�o�Xec�ު��7(��@�i�W��U@��mW�3̪bG"_���'��kl98��*�!���͕�{}c��l|��J��㠚�B,��x�p�t���I�w:Q�T�������N�yB��16U$
@Ǉp��l��)�&���I���s�!���������D��GTs��� �������|D׉9w� �<�`�&@U�K#}\��>)F{V�%��N&�E� UW����+��4�Wo�`|* ��= 0���J���<4
���G�1�)��dخX��+�w(30ЂC�i�nXP�<��!%�i��J��_?�?|�|O�a�̰N>�t�X�O�[�r�=�C@�qui�H�1�V�@��/L�I��a�E� y:D��~�@a�)]�+a��2
5��jϯ?Q�W��O����.LR4�B
.��8b��o��ߜY�5U:��fU�&*�:݊��I�!�|�Q|h��R;J�v�N�ǨޓJ�'<k�Q�oR|��%��
�IwKKK!����C�b 0XH�ߍ���~�5eT�:a��~2�F`�	RB ղ�@V�vaMN�Ձ���
U1g~��V���m�;MT9\OnU^ԝG��s3b!��*�P>�#b �$�Ψ������-H>@_Dj���3V��a�GA#�|��GSDr{��Z��-���
H��2�����?N�"����UM�1�Q&�^��� ����Q��z�T��ɢ� 5c3اA���aa��5���p-{�_'j���X�D���GW�J��m�M!U?j��AA��?�����8���
A.����-�>��Ĩ�J����q��!lk:U�P(B��0���J|���88𥄊���|�~_�Rw8ʇQ��]�������|�W�hH黣~�aQ�NHS���q�u�m@�7z�:�/nV���?y��<o; �Q�cf%Ē0֓�_0�B�E� �����R�Q��3�PYv'�C��l�=��A�_����a�Vdn�'	=2	����|ƑC�a	�$H[�HD����v��f!¦M���RƠ�ؓ��TDD��\J(4G�s�?{�.�PϑRKL��,햢�U9�;�A��X�F^iaE<6k|$,W���d^*=z�P�5%� �!^b/��߽�Y��=����8�m׷��d�G��+�H۔�������@0�&A(���6�[��W�O/.8��>�??�۸z������C��^bFL.pE��uyI�P�<���KP�v/�C04�5jU�h)��;0k¯�ϡ�n1="R�<{]4�e�T�	2�VU��4M�i{��w{�����A/����}wf>ذURE���7������Ҹ.�z�����L���C��l?��"@ioE��ZQ;����������koS��r�����rl�g��u��_n����5�KS�ԁz況jc��ĈdZ��%u=�Hd�b	��0
jʟB���P��f\Q��!GE�"�@W.�ut�*F�,����k�	�/V�T2���_�o��F����UC�2���u1���Mb��R�M�e80��*Ei�M��q�Y�N�6 �\����QkQ	�`DjQ��Ƌ�R�S��-��Ѧ��$�d!�]��H���(��� ��lD����h�_�T�'�[9^��#ZHjב}4�$�DD\������SL4T���B�FjH��_�3���c�p��]e��!���PR���)��Q���p��a�^���U�2��H-�����Ί,rD@�Y�َ>H��Η�#��	b?S��:�DI Ϸ�Uj�����`=|B;	T��S���ѳ��o��.B�zw#u?�w\Uѽ3������I4�}*TRP6s� Z���1T�+�u���1D}����.�߅%1�U67'�
�F��	N!�����U�����.HAc��_lB�ϫYKS^����oG=+K�*rn�I� z�^z�PًS�x`����	J���T���U;M��n��O�Dp��'t�=��b�۫
��	qm~&>w\��V�R�

��ӣL@�w~�B��;J�#��|`�z�����	�����p���_����Z�a����I�"�w�bF��+��� �e�f4'1hY=%�Uu@0�<"��"4�D:���@K
9aW([�AL�n�=;�_��$����/ �ml<���.\��!9��W"�1d �傿�$2D��,*�7��� �I�跭�7�T	��lVE��`����_�$"RbE�_�/�>�Ŗ�Q�
��w��� J�h<���  ��,�)�/�a�m7�RNP_�<V��~x��$,�.��K4�;!��$�@�Ru��̷B�dq�p�8�p=)pd` �����]z-O�2X�n�\�z��/:e'D�x� �����|�u��t�4�!��������~ �븾c釿[�y���h�B�@Il��:�x�@�7�� G5>I�����!�0�k ����YF�UD��RƚO?@�k�����������U�A S�Ƨ9�"�80�Ӻ7�b����t���"�&�s��}�DJ�U�p����v�pU�u�����cU�.����/���A��Ђ�e���m1�J��"��a*/N�j�T��M�<�  t}�_L�K������6������m�����

�G��۰�(�W}'����ΎL0B^Yy��ԥ���"f�t��X���Uc���0���C;�kE�g�d�.9a���I�*�����5'E�v����h�cj�YCU4��b�c��o���V�W���a�cUEB����6F���e^�T�Z���@��8��AV/0�(Q�8c�(r�*��t)]q�?�����+���EH�v�W[���j�$_��'�1��2Sg��F�*����~ 2}�
Ĭ&�W�sװ(����L��֦�N�Ԓy&gP��C!4VI�D�\��c]�D�)�y�֡�(<�eY֕�ɦ�ŷ����Uؙ�̍����j�%ݬ�	���pRY�|��@_>����j?tߎ����?$�E� 'P���X����JB�Ղ��g$�y��S��J�.�]�A��%#N�^�U>5���,ɋ�f�ޝ�9P��L�`�B�_�o���Lz��J��:����!~e�4��m����³-�S�(�п^e�?��N���>r%�<u�
�W�23�	魋 �Pm[���N�p,g�`]�iwl�d�Bv0�X,B�t���1�*�A� �_Y�~q��*���+������+��o��\G���Y��c���8X��d�
*G���X����T�$���H��P����J΋���6@���9Nn��<d������ .VH�Kx�:�j2��1Oѡʽş�\'J�}��|P�]�����+�������]K�C��a����˞�*� �3"�O?�`T�+�+ *Q֪Zќ³>">7Б@t�Ue��e�JE���0`i���W���Gc����Y]h�c�9���*+\��Ģ�������E����C��u��2P�u������[�1�M�
������$p��[�n����0�)Υ���.�����Pf�4 {���~m*棃���/t���$N�lI<F)Y}M�q���wA����,*G+�DK���,7����#���|Da���,�541�4���0��0:���`����dF����Y�D��/�����l��&�a �\�c��p����fD�4f�G=���\q@q`��3L�0h�m��۳��b�G�y�9#��"+���G[���}on������9��h+t7����m�
��j��Tm(lxKb�KPj��ŋ< �]��]��W�(�w♇'lc�%]�
5��8���K����3(�N.`p� �0�x���#�.�����D}�dr��� ��Gi�6�$]����
v��q��2�I�_}xz�\8��ꘒ��j�?�	�[�� �h�IR$�E�H���N�3vZn�\�QG�Y}����L� v0�<G��Ma w���+w��~_9�3�ڶ�83����$�`f�"���.U~�!P�nv"zܧ�M*�2�L����f�e-���J�D*$\����9�>�*aa8�Y޺��B�Y#�M��٠�;4�uP��$���}ɣ�* ��S�U]�@�Ҽ즨��%CG����1��O��/���SF5�_�Yďm5�j�fL#,��Ź��O��Aw7��?~�*l�n��*�;~��+(+� H�A���%�~Κ��g�1!�~�t&�W���%�H� ŠKgn����:��I9B>��q/1腛?�)��ޖE+ ���"\��$��a����_���Zד���e꣑]����0;��i�e�`�S�z����Y��U�tt��;q��ʁ��F-tA�u���,t�q�����MMUE�Fi�}���^Tb��]W�E��s.�u���'�V=���
�J��@\H�.XE���]�]�!�sD�&]����
��u1n�����_Fm��ӿ�XG�Ǵ�����<d1l�Z�R��|<�-���<�
T��UӠ3d�EWF`Q�F�BU_��0�Eޠ႒.&�*��4d��c����}�d�bu����YHRj����J>�G�a�6DsUY�@�����r�*�ޟ*U��#:N4Z�cèB��Y�#MJ#���;��v2�fT]��9#]�/P>A �N"�<�c�i���K��2�M6|�����BS��6����M�d'	����,0�{���"�Λ�`�,�Z��b�F ��B
����9��P���{f/�ap���E�*�� ,� @$ J  `B JC       �9� =
4��ۏ(�,#I � ��0m�@�z@8�we�t����x(�8A�ؽ �6À�	�/&�e�@`B����B��.��x&	P�u+�P�u�P`�i� �Dh,h%c�0�>!���.���l��P��h�C���C�E �1B�Ț3ٵ>�J�`@ĿPC@��CL�k�l�o�և�`��� �������0�S��V�+���_?D@U�@�UC�^�0�iC�Qz#C�T��9: ���
�w<�*�l �T! ��!,���%!������)b Ȑv ��|,0�)�l�n0���t@mVVkb�!C����:$���T
X�P����[
�@���R�A�$0�AiJ�J(!�i��P��CEJE�r��%H�T���e��(l�t羀�$H5u���r=h
&��e��0g�:`h d����9
2n�+~ U,S_�r��Y�=�{�a�9!x�ip��~l�����;b�B�&�p�y����S]yY��	m3�76��q�<�w��nC$� �_�ZA��Ͻ/a��k�Nj���N_S;��>�-f�֢>�%��������l�SO�X����a�6��-HL�B�lP��ƕ[���H�(υ�/%{����VX�5-��PB)nߝ�k����g<�s�+z��E����L֫��i2; GŒ�ȯO�zX!iӯu6�uW�lw��8񌻈�]�ׂIg��a����-�X�2�<l��Ͷ�{Pȶ�5h�H��T�Y:��C�'v��]����K�M}��񢕟fѢv�$f����!��6��mϑɲ�~,׀�F�o=a�J,L�qZ�Vn/��z?�ƀ�
FHx��Ė������7h�s#�{����+�{�W�Ӳ����:���b'-���;BW�a��tP�+_W�'����IG�v�u��Q�no}��`qCJ��\;�'��י�&W�.����Z0O
a�%L���hk���웥�pX�s���y䘽z"2e�ӆ����Q�:��]nvo�;�f���� ��m�=�5�閁��nl��W?�Κ�&��d��-?v��dwV�Oʴ�n���Zߙ��'''�l���{�s�?�0������A��=��5����p��3����Z��S�h����j׫5w��!���l�K���PǾR��m������}�؅�]�T�����R<�`w�m.�Y�v��2��p��
7�3P��������I�&���7�ٌ��qy�y�o��[����9ûw/<:�@��4�R�^�����e�Kp%m���VS���kCevϋzwݑd?��V���Gsf?�ºj��v?9	x�C��<[����[���R�{�k�7���f��7�,����}�����ۿ�<]:�_�5�����m��?j�5�o���6�-��x�(񳴚�C�pܩ���\�ֳ&b]�}\�t�b^4�Zx-�}�B�7��)��T�-�Y�as�x���M���=i�J}���ut��[�����fb�	�?So�s�ԟ���c����s�+���庅z���I�mt��u�z���������rd��g�(�xX����S�ەi/�}8Cǡ��q����5����A/��#A�o3�����@A��		�(̚D�/ Ě��oF4W%0Id��0A�+�K%�$�@�H ������z�L ���|m	O���JP�TKQ��T�C'4�H�X�Gh��6/�Ҥ��e��D\d߶��E;6�n�;#�6f� \(H�e+ɕlҖP���o;+ �v]�q�
�J�&%��!�И�.��.3�Y��
0A��&�Eo�v�&��h��(�`���;� .�Bs7�R��3�0W��XJ,$��%7Q�<�" �@������AQ��ߕñ�Yd�ߓ�e�dðJ`�ӄc2�JhD�"  �HR]��۴�Zf�l\&<�k�*(L2�!N+��:MO�F�1AЦ6��� �L�	�-I�Ŕ�.H�)����0(�8��\6%�)
>�N�g�R ܹ�B�;*<�K{1Z��cM�o"Kw
.QM֮�M!���L�H�X$4pf4E�V�j�,y Y�F�F��i`p'<���,06��u��B�p:��R��E�&�E�[�nJ�N���`����c1n�`�M��1@/[����Td(g	a	B��ee9%<QD`j�

�^ ܌5�Bݳ���d�0��7��A;�w�`@�J�jʀ6(���b�Yt��l���CiwZR+W��)��\!X.(B�(]�HҤN�6 .��3B&T�R6��B�C��h$j�F k�֔��*��vV�Q̅���^�
�b�vIE�J�b ��	�bn�S�e��)� J����L���27,S����ʱ)��enW��a�Ȣ��xM�P��f$(^8�:2C 2�"F/I�FD�'P�Ї��_��c����
A��=D�e�$�YԄ<���Z���Hᱰ��!c�L8��y$Y0)�Fl���1�Pk�]��3���=� ��ܱ	����q�qrAU��L�P��ՠs�`�UzBXi�,3��*b0���Z��؋��H�p���Rh5��Q�Ƥ03�_�4ð�z�4�R^�B�Cr����S"x@>@s�[�R�V��
��d?'�"�a�����<H�"�7b�BQ�[�	�,p	z�Ԝ�Go�`TA��-P	����e�J�T�@֕R�RB�8R fB��� f�S�Pi� �@)# tp|�g����Û�:2.v�,+Z�ބ�Q�$�5��.Tg5���3��H{nM�ŝ���{�P�=GQ9\3a&=Pqʹ���i���qqXV�}u�  D"    �B JC �     {J� ��?QDhT��H�MF�t��%�����|2� ��0 OP���22C:2J���_�c�/Rc�[rkdftv�[�x����-�u;��&+.����E���� �
�"aˊ-�
۳,"�H��p��?�`��ۇ�R��6�|��~�A_p���Fp�3M[9�2͓���OJ����IPoQ��|�"֒��n|�r���ƀ�����n�S-5�D/��^�  w����j���X+x��?T��D����;[!��jt��I-�|\�2Hp�}����e�	:�' ��O0w
�6�g�T5IJ�{��U���;m�@����`��^Wc���J!G�ދ���E١����w�2�<�4(��x�������i���cM�G�=�$,�	|�	��Ί���{�x�����Ǯߢ~s�ОY�=~{(��瞽c�}�S��_d ~r|�z�CQm&N!��ߏ�R:c2�����@
�I,uZUP�>��� ��ӤW �)@��e�{�����$lɺ�s����°c���]J۷�4�-i�>*V�z�~:N�����AvɆ���p)`A�g�Qtʕh��m�BOk��Iu��ݷ��n{�(�za�]i܏�k��7ŭܲ��&����^��,?[� ' ߢTn1p�2 a�|RܺS`Ĵ Ú�g9�M[�{�HR�a�[7.�+��Mi��1��h�Հ�
Z�9��J�F;Up�o��K�
�F.g�a0a��bM&��xtY!�,(p�������	If�N: FB4<�	a�~,�|���T�`@��B �$�.�ditK# � �*NbP�:�p�+A"9�W���ɸ2��"�@�AQ.�"����A��Ec%)3٢���;)�t]w
V�e�5�"�|[,MUJ��tD�}2���広6��1�R�~C>j�6��m*��W�����@�>
`rA��29�1"��v1���9<��o�F��$�*)�t�[OW{� �4'�>�T��ڀ��d	k %����Jc�L�S	�����HR3��i5�	q��&� �5�å8,�ɘ�:������6,���N�Hv(S���N���Ln�<�b�J�;���������y�Ѝ�[�(�ڱ�%H#�h��u0����4@�Bk�DR*�P�pq@�$0 \�CG ��$#�Ԇ�ԌЌX،,|Pl�m����lF-�4��J�QJ�n:���< B#N��6�f�?x�,G�� �n�;����(�Q�[	�T���m��K�R�s݆�+.���i�����Z�K�I��m+�'�BX- }xL����_��ě5raR�������0��
�7�� ��LS��� ���*������.|�Rd74m�iO��N]b (���4��stB>"	��z����b[$e��s��?x���Utt+A�P*I�u�z�q�7���I�*gr�'�@S��ؽ�"�ͳͽ�W�cF��f�.W�� ��j� {@ؘ���l�,�\ى�W�S�r��?��?��?D���x~�Ҳ@�ű��W)�,%Jq���G@�
(&���Ҽ �����B��ϡ�ZrI�s"2 �� ��K����)Y�Ts��^��PU�+�&viY(�OG'>k����,�h�fa��H_��L�+��*~\&)��j~Q��^��ʳ�rJ�y'v]��Բ��L�ui����Wd���/DU),�گ��O�.S{���b�k��B����a�(�MzN���)��گ�C#i���></��Rݱ}���.��G�����_��_��F�a��m:�#��	�
����#b?�P��R-��R�O�^*�3M�R��W18�0}زn�^9��[ȵ��Щ���g� �Bؘ.�����*@C3V��)d ���0�F��4�Ka��@�V
#���("iA%S��LkVP�
��_Z���n�.�<�a� �*'�Mj���U�5�^�@"��Gځ}��%�;*�zTE ��� 
��yA�"������cRtK�|m�Y��վ�k�K��D_H�S撩ΈMb� mJ�E�'�!� "��\,b�%~�����(�y���[�����zV/�p6�(���p�<~P�y| ���}Q#d�ڠ�HtE
�AP�ă[,Z�fD���sA�9"�?���.	��G5�A�jP�E�&6�s0�xb�4�$����P��	�kX����2��.
�"L,�����������e�A�%���r�W?�E*�9t���K_�E�ؚ	(,�aj�?��b�F����E	L!RP)<�D�aK�fSƔ�Q�5QW@�U�Ϋ۴;	e;�\:��x؆�Swk[�nG+̕� J�6�C7�F�ʄ�$�Ξ���h�yz�`݊�xLc3�ј�"wx�b+M�cإ��Hŝ��V_ ��\7-cU����B��A��+������B�!~@E���?� ������74k"+�?CF���p��!+�B���ҡ V��ń�������r0�2�P��H�V�m�Ҥ��SL�J�
�ժTj͊�ٱb�=k�,�jӢ�-ۥ��}ݺt�͋��d�`�5iΙ�M��\����S�ڣ7�hm�3ֺ��1p�t�тv�@	}-Z��(_g�������������c� �xb���]lu�>~�Jz�P����J ���G�Xz�
`����H�C�D拵1�<��J��X��%��s0I��@�H|:e8>"�CV���C'n�����~�@�ѯ�>&��XӋ����Lx���9*Y�nƜ�'\L7�7�
r4Z�X�r�D�؇�(憀�T��J��Gn����A+(I���E�cDA)�^��Z���}fB3J���a͟��<`��w�_��|�@B���bGX�;,ݖ�PxX)�'ɧ�����ky��^��+�g��-*�YI8��K�$U"��"m�&�@�0�0�5�C����Eq����0=B�M�~�"�� �+O��������r���?f��_uo�{��F���dJ
��}�Q�B3~0�.Te8��}Y�Q�K�m;~EY�u����_/ؖ%�`d�R��־8��J�LJ���F�}��`-�¶��r}E���#�8�H��+>��ċ���*T�J%{V>Viԩ{��n�dv�%"HҪbR�h�W�K�\iے����DЕ�v��ĈX)�#�-a����d�+���Łr��S*%Y�p5H�
�%I46c��rny'�3�*�H�0�c	��$P�V��4��`]e�u��Q��C��!Ȼ�:/t�!%-�CɑK�2�;�1-��czs�*^mn�m�n��ůk0����i`0��j��0ᐺD�@�ݭL����͘bR�L	L�=�������j@*�d	�+���4��pb�C�>�FS���)�)����8��1��\�T^�@c
���G��y���{⃯k�W�����=�	�e���Y	%�_0Ղ��y�2sCN�.6i�Y	�x�Ue��ї�Bc5�>h�5*�W��@

�:���J�t:����5t���[	��4	�*��H�`R�B�"�P|"e6#c��n�>L��(�N�9�=Xlu�
�a$�����o�Li�����x�9�طCj�u	
YY"fK�9�_����#�r$����G�%�l�\-a�%���G���>�(qm%�D�����h��.G�%��k	�)����\�G`%��f�"/��J=|٭O�í���M�����#�A�ȺD %�[����z4$��� ���JL#�M�����CX R�A���Dܣ%���� z�Sb���-QeI8=�2�Iu�8��"v�g�b��pk7r�mI�=2�J����%�"jQn9
�Q��J,H�E�;�ё�H%�=�*m�K�#�D�Ī� sY�T����z4^B͗XG�%�������Kx{�[�`��̆hP"�Qh9��S�K�#��H���)Qn��#�r����	77f�pp�		7Z��pC��	7Ny򀍞'���y�����۔yy������\$y�������y���''۴yy����'�|��A a%+�3M)�E�3e]	� ZD�Ą[���������  o!�(���(4`3b ���R���:o��h3��^	հaXLL$Ӧ�/�Xza�L�L�h�d�H �Ctp�n�$����ْX����h�C��hY *c*I�Mśb���rz�7��7ݭ7�zo�xI�M.7Q��zaX�ѭQ�ٍ��~��#KCE�Mo>i�I��&�7�4ޤ�x���Mo7i�I��&�ƛ4�?���H�G�i�~��#�Ə4���{X�#?0�j�����ěfXo�x
��&¥8���[o�Zo�Yo��o����M�a�ܷ~��~d�GD�G��G�~�&~$�`�?���vu�qE��K�b���0�Q�x����0���^�����4���/��E�x�LqL/R����"��Ȧ��E5z�L/�ċdفHGł�$aG�"�e�Ja���PM� �Ӈ�Y�������������]�ì]�f��`زw]���E��*U�1�d# g_���L���i(
8���I��=�U�E�-u�����R؛*��x�#�����0U�Ѝ�#�`�E�F�g(�YT<��V���1��Z��`D��OMk�y�(�Ǩi�\IZ�/��$�Ħ��f���7<��,�%���t�ӱ��`f��^!����P`�)�/�rS�
Q��h.�6�d��5H��0���*�T`x�,�}%��`�E�R�Q�
G-N�)��+X.�c~�^�ֆ:�ꐛ����Ⱥ�Q��-�q
�*D��4hd���l*v)d�۴
0�	��0�T6d�c<^t؟�mX�UU�[ �������S�$����"�gݘ)�R�(SP��M֝k�`7�
0���N�k��t�8W#�QU�ԥ.�u�?�qXf3p^K�)<�(By�A�}>���MU?��P�(��؊��.��WeT��8�Z�������(���n�e�f)���c��
F����F�ș�q�Z+�8��0��[� �d�M+�U����bi�nџӠCԌ�m�����X���1v����%�c.�Dn���붑n�$�r$Tk��ئ��	UB���L�Vh<�`D.}lWc��l��?��*��D1�Z�����E�B��23��1�Ũ#NA	P�2j�r���H5��P�U���׳9�mf0Ƴ�������*+��R��U�	e���R��T���!�%�f4�hY�-têi,	�c���]6h[sQ�@�E��REA���%=**�kY�|g֨IcTfdf5v���^0� w,�͇-U�`10��@OJ\���TK�	A%����<]�2]�hR`:M &��V`�V��M=��n�l�"� 
��#2��t��z���h�0U
%��pKS�S��5(v"̍�h`=6�J���0�s��=��0�}����Jp%�>Q�(J0!�;t�(Û �,	�F �L��'���N��)�X�8;��0*$:a�I;n��)���0:!�);wA�)�0}�8p�"N�	;:��)E���ۧ��Pf��N@y��'y�Pf�JT{�2c��$<e�>q�G'�3QG��<e��g'>quBC'�3M���<ex�(�t���4��0�IGt�<1��4[�;� ���QJ%(:r�(G o�+�JL�@(����DQ��L��	6O]%��v)5z��[�"}��ʯx�t$�]eО�Bʥ*S�a@�Ӕn�V��@@�Xʵ��&����y�j(��_Ŝ��'w��Z�c�\Ұ"���-S(�
;$1UW��8�����T��ʬʹ�L�ʅ��	ܙ7lE���0&@\(6$zCd�%�+�bZs[�wE��j��%��X�Z(Ha*x��Y�MU�J:�g��DN��8��զ�ɷ����$H ��c�\<e�hƗ4���ZQ�Z�X��Wh�A�mJ����u �0�����h`���br��rQ^�b�0��@� ��0 �.V�,�K�+`�Ǡ3z�1�ȸ���x����ӧꅠ2f7��B�`i�Pg��{�����a��B�`c;�tc��K��� O����3[���FC�<�^D��42��/�b#�P���.q�y��Lp�7�ed�&���Q��s]�bT!b@��E���I����
�����Q(�(���y皢�=��.��p��)\��x�Sc�3}i�.2�L32�9ƙ���8V�Fu�@���(g�c�h`F���/\�2���x��Rf�Q4{J�z���.�+2o#�ߦ>\�@�����Y�f��d���3���ʷ���A�U��kQP��Oh��KuL�p� N�E��e�l��Y�,Teh,�tq{)��b^�����]o%�=��t5̗Ő�Cfd��=�mT�7�z]p�zQ�K�gP�|�;_�_�ӧ�ɘ?���I�G	�AE�2{��d؛e��Qmn���,A���+�����%I�pR�W�ٿK[5��� >g��t�Q��D�b�d|C	3�ۣr�L�,���z�
�#b�N�ɬ%:9eO�,Lk��4�z�����/�ܫ}IBih�L�e���v�0F��GG!|�y�Ȏ;����xjB�H�ɐ1Y�i֠�f�r�'�]�?�}�^��x�F��hh*�8m�Κ��_���3O8
�3��v(5��p�(��bu�|l1�������S��(��0�"�L�I�j�t��l,ʍB�;yy,58skU�%���L��R�|���{:��ᙆ1��&�eWCK���1 ��s�9��J:{*���� ��X�"�e~Y6��7�c�p�c�A��F�f��9IVZT+�Uo�t�e�F�DEϭ�Eզ�yZ�J�$h�`/flMl��c�]/?����
�2L�d�أ�=�;q���B
K#;*Ad�(���1œ��b1�6~��2W�:�if1Ͷ��C�����8/^!i�m��TB5�ᙓD���|@�0��q.���)R8zd;��9��cƚ����J�(��I�ߌu ��F#泾<��+y�b���؍�.@��͜1���<�����T �c1�,!�И�:�F��ٗ�WP�p�T�C�;v��^���5$�6�Huᣭ-3Ok� 롐B�y�=����{�]pՠY	X�<�v&vӭ�R��P���"������߆b6�����u��Fᘓ��=�WN��BS�Al��)$��i�f1^��Q<^a��e�[���ј^fn"=l�C�ѺPx�z!�[i�˝�֎E��.{'��c�Nd1���8.�5�-+�1���yZ����(�㍪��{���!�;���{e v����U#��Ҹ��~�����y[c�.9>y�(��#Ŧ��\X-������su���;:\E�ʸ�(�6+_��� �c�bf�����;~���,�ʧ��,����8��1r���m<�O2�V�]I�_(�4#�NS�=�12�3�`���R�>dd�抁�5_�0��gT����ӊC33�ҡQ�F�}��hѫ_hn@}Ӹ�W5��s���6w�82s`���0�C6���� "���z'���ݪp�^���"�8����P*�s��فq\��k�s�'�)R=�Ƙ�r]�r@�\%��"�+�ԳOdV>��|=e���������t�X�0 �up���M�ARb� ���)8���W1$����_ůQ�1y)�uѫ&N���U����E�嗥zV��TGT��Z�$Q�ov�w���U>�QZ�hq�D&,�V�-�W�$��K&BZ��jԈMI��YS&
��2������R
����CT�W�	̖��c�f��x��T�)n�-&��B��� ӈ��S��Zlt�mm���b����hR9�[y�ؤ+K\�k���%AjjR��,e�|����-�P�BK>Lظf�/�y�R�AYt5��>�U�*U�E�fAެ9V��"�j��\E�I��J����Ū�X(N�w�Q���W��yݘY�)�e�Dk��a$�[�cP����/�d��ʏ�8��ѩU�g�T	
�ѣ10��qu�*������/v�8R�dH��nJ��XU�АC[�Z1_��\�:�K�����B���Qhǆ@W˲�rA
,�`l��[2,m�^0{�	ȅp�� ��C>Z=� O-�� f�0��:����(	൲4�N���缈����y���Z�#�1I�k0�\����ao(�ְE(Pt�y�ވ��ۨ���Jn�Ej^@po
��
��COW{�/Q��lA� ��_)�8b�PС+��
Ǽ�B�kK����22ӫ g�4���+ݪ\��W������y1 |��A�����fE{� ��N��
b7�p0 �@1��&~Λ��i�e�,4E��h�	����d������0���ڕi&Af��_*���ƥ!�b��Ɖ� 0q�U�؎;1W���ur���ͣ�SY�0�y�YW]�s����U|f��ٲ9m�mm���{��g���ή,�m�}�Qk#����ldX�`E���7 ��S�,L����	i|��}��)�F H�ђ�p��ph*Q��$PޯGS�Qoُe�Q���+K͋�'F8E�X5muQ�S�K����������"?W@M	
4H�0�� �r���gn��	�~�����-V����̉���`�W�#w�Q��u8(Z��p�6U�tXXl@W8��������'�	�Ε\��D+�2�*ی����lڛںL3� ��,�@צY[%�	���w��"��/S���W*L��u����Ba*�H���UFP��� �А��1�}��4Ջn��XסS���iT
��ȼ�����Ӏ�3ys	�桼�����@]��ylo�.��<77p� |`��]��I����Ln�% ;�G����Ȅ���`��]�7@`�S$d�.	L���#@`4�"�dH	��S�0�= �M��Z@�8�"&sI`�r ��L�IY ���,Xd�n�YY �K�uEÓ*؁s|*�:���wݲ� Q��sK*T�.�3X��z �r��c�Q��/XZ�� ��6�R,\� x�Fܶ�(l/k�Y���+k*Q�cj�WDw.�!̬�R>���w���� ^0�m(=�L[K������@��`;#މ�t"�NJN+E�c3qXz .�Ծ��p�Ɯ���
�˘[��� /�6 ���p���7Q��譔~�?]2�\%�NN�L�[���T*՞��mtU+;�]���LЛ�`I��J*T)�Ӂ�_�	�R���8:0�B���فu�H=اh�aAJգ$nt`�D=�;�ӝǂ<�0�8���ǩ�cA-��сy��<���c��aL���Z<t`�1�w㶦��80���(�uBR������[K��<+���F�"�"�E)�p$"Gc�pD�Ge)pd�"Gg)�"i)�p�"G0��t�V�q��Z�߿���0[H MW#���������!�Q])-_R5��X��a�*���VpG�7��i:�8
�U��I`,-�Atp�:9,	\�aR >l �� �"���9z�J����
B@da��;*�E6Ƨ���b��{1e�K[�	��ؔ$g4�l�ӳj��_䛝R8�k�x-&�S�ݵ �w���C�J�`+��$�I��00���૜x#|��k[Q-Z�Q�E�WEɠ3
C�݉)����w8�BWtn���`�eb�d` ���f|��<�LC�D��]a`RG^��F�^�a��T5F�Lm�F�DQ2��6-�
X��w彮)���b0�ppW��?ÇO�(&Xa��wKX��!���x,@�����K�*v�&��fT:�U�D�d���R�NF�O>��0��G�SX�IX�Y!O�'����R|Ga�`1�EL���P�z�a���_���6��#j?�~��6 )@bU����q�A�@��큀B�gU������� �8�Z�q@�|���8��!�NT� �;�i�"����9�E�M��I훘�f�]Ǔ��r���w���#f9�#���	o�$�|ˇ3b����d�$�����&A��0�)R!_�!��?3aL�B�� (�ta@Y|=TLb��p�s���M���CE4Q�RP��P��ؔ7-<08�s!�;�bK��e�a&��X>{\U��-U2r�E��u��W��NHe�Xa�m&D�|�Pae:��&�D�0�#��urJ��g>.X�7
�b�wf�	�A��\�ǟ�Rqve�F�ŀ�A���PX0~�a�S�%,AA؃yFU��X�@,�S�����,
8��:j�I&̑3*+G��g�K�&<R`	�2�l �M0�Ώ�C�Կ��\��[0`j�6T�y� �����}��n�NJɫ��oQ`��[)�0ƼՊ��h3l����s�cy�W$'�"�4�4��}��Q��Pl��k	4�WP�vY$EƋ������\�*��rQN��a�R0[	;�K��sx��s�U\�#RzT��
^A� tq����,/-TN�(c�׸`=Zi�\�й�\D���Q�8.�UR��4�1�,
��wՊӷa��Y�(���rU���i�f��Z�͎�1�=���u�DTR�v�+K����)[�n]�(*��R��5�\JI��_�� J�xfI��N�%, 0���/
"�,P�	Q�ٴ/@���Xg�r'F- �Q+�X�3�TF�B�I O���h�t")�t�(qP"(1T��#�>]B�j��uɤ�3ٲa�ʃ`s3i�o#H����@0�Fs�i!@0�*���-%�
�ɐjQ⨅��K��M�jW��uDf��6@$��_���)Y>�T�q#�۠���C� 5�!e�EpTx;%�$^�TEe�����)��.@̕�8�=�ⰪM�]qTq����T`8tZ�nU�Z@������m�7�p�W�������s5�4.BX�v���F]�b�ͮ_�V�*���N�����������J��;���@așQ�w������y�9F�P�o�S$�D8&m�<��Ӏ�?��*{!�C2.��8B�d�*������,�v��_ɗ��'(�*=�b���"��ª-K�F.��<����A
����x.�6�.�4"O-���ꀂ*��.��Z踃�D��C��HuXEU�e'Y�Fn��9��nꚥB��v�4���gEpU�����xD�8��ʄ�+��B�+�_͜�m�v�Yp׼ED�C����R��]UĔi;�����͂c?;)��P_|�Tp�W/�l�a�`P��`R� �a�B&,��J�a�ˊ�(�u���u�:��F]t�K��T*�!�p�T�� ��T�cp9�y�V����i��v<l*�6І9Uy�~ӕc0�d*n���A�
�l\�ދ
0U0��+�|~��82�5��N�و���({��<�蔯l��ϻ�ج�����h*b]R�fZ��?W�0z�$������I�.�&����X~Е�Q�SV4���L�vE*R�Abn���v�C�*�۳��������4�ʍ��0�ւ����vES�ҌzG�ԯ���ic7�/:Ō<(��4�Ҏ;f�E���w�bHV��V�g	�V�",3�z��:g�
6��C����[����q)��c�b�<�����S���߫E�j�qT��e!Ce�饠��_�w�]��G�28���N�1
���Ɓ�1�zϣ=Ⳳơ*�/��Ky�\+M��=��T� �:(�q԰h)z��-Օ>|��1.
���6!3��zمfŏ�y�;�� �{�c��=�."�Ū��y��[A��!i�Vz%���	K�X�ԅ&Gn�a��v�n�j{Q,o���e�ܥ7QUyQa9W�P$j!6vccdԵ���B�T�-�i .u-p�j�����C?�,p+��/���B���83��p�ֲ�,}���9�_�v�!�/����2>�K�3���!OW,��	�+�Ҙ���f1��P����`�7��@���$'ova�����Ҟ� +�N�����\I�n���Q�.]q0�S�@�@�+Q̵J��D�n��Z2
�,�^2�,��#C}¢d	�DT%�J_�H�	q��K�%�,A�8�DW"��Չ�Q	�D҉/t�b�ĉ�^%�r�@K�WB,QV	��D%���pJQ�('~�����i�s	HK�% K��+��"*Qu��S%�F�!��A��KD[".f	�J|%�*���U�O	(J%)"1�x('|q���%�1�8KDW,W	�J@%�(��P�RD�%�N��K�&�P�@	��9%�^��J`L�"%��J.��n��\��l	 K�%�+���DV%�Q�0J$d�v�<K�%�,��X��X��\�xJP%")����Q|�&�%����K�Y"-`��Jh%�*A����S�G�!��%��K�[".Ah����%����JDU+J��:a�Pf�/����]%�n� K�V�+U	��<%���`J�P�(�쥈�K�!�-����Y%�X�PJ8_b(a��u	�K�%�,Q�@��WB�D�	�R�@J,%)"A�y&}r	��%�Q�PK�W",X��JH%��D�x�E����%��K�[B.Qi	�Ĉ%����JU�*M��J%�\�/�����]%�j��J�T�*�L���%��J<���t	XK�%",q�	��W%�W�pJD_B(�wH�K�%�,q�P�Xb�X	xJH%��D���E{h%~�%�і�K�YB-_	�W'�J8%�(��X�DP�	=��%�v�HK�W",QU��D<%���`J�P�(�𥈠Kࡢ-����Z%�b��JhS*1F���%�K�!�-񖐲Zb�b��Jl%B*Q�%��S�(J ��/!D^�r��K�%�,Q�@�DW"�V�XJ8%�(q��DPy	>d�%�і�K�YB-b��Jp%�)1����R��D	%�PI��K�[B.Qi	�Đ%��K�UB+Q	�J,%�(Q�8"�_B	��%�t�PK�V�,qT���8%�q�PJDP�(=4��x��K�%�-�	�DZ%�c��JtSb*aH	��%�C"�K.q���D\���Z��d��Jx%�*q�	�DT$�K��/ED]o	�K�%�+� ��V S	HJ4%"(Q�I_t��Ĵ%�a�HKDW",V��J<%�(��`��P�	=�%�w�`K�X�,�X	�D%���pJ�Q")#���|�xK�%�,�����X%�\��JXQ")����C�K.a�ȶ\b�i��J�%�r%1��-ͯ������Lf�!��/�\�+�����h0R���!�)L�bu�_b��� ��>r���@���XMW%�$$���¯.E��،�mi��O���K�H�b:4��*P]�W$laM�d��4c��T�0zq�I���@�0mʩ~��O'UT���e*<&<�P� 6�S��6 �L`e�&sGX�4���K��,4b�мd��5��1������z�%h[��L`Ԙ��z_��	�axDfXy�!��m�7��aԱQb5�F�6�0��q(h
�ʂ1א�4�a��P8f�0uĄX�9�W6�wf1@��S�ݬ-ŪI4���n��6�:��Y�њs(5��3LMɚ�Ab����6�̚�(���a���09l�
�?�W�
q�8�Y�-p���X�}�Ȉ� �a0m�RC<�)�1�bg`5R�@�Q1��61(d�1� �'��f���`�C8F|-B֥5X��UfF���7�ܑŲӔpm��alP�5�lў��Lp`�C�,3��t�q�,�~dZkc��:@��6V���*6�|&%�00&��!)!�c�`n<`"�1���h�j�
J�g��>����\�1�fo"̪Xk,R��j��%�a�j�e!��6K_�Ȕ�����9�r��h���$Y$l��a0!�r7��1a�3X�r��1����;U�3�ŹCn.�xl�4(�y�轚p��50`a�j�����s��doX�󉚫�I3�,`G|130�XV@C(U�Ѭ�M�]g'��̦,�	j o�*���;Y*�B��@�h@1�,6��$�Z)��2&��j*����BcI���X��FfT�%�6;Ks����;T��d�@�{6�b��zx�Ȃ0���i��"����;�fɍ���.SҚ�b�B9��_�>je1l��$��9��Ġ��<�8���)��LB
fφ�r�} �p�SS����L�Q�\��&�8��a@Zǋ<E��;��Q���O�20"�� ���f�<aߵ�\m��X�&ys<A�!�� �U�,��?�b��r��6Vb ���0s�A�8�&�Y�R����D$0�Jp#P��h�"�0jblV��3l(y��͞��ɞ�yL�k`f�`+\�Ŝ|}�C � �1�hִn�b�[nSuX�b�@Qɰ�:~o�eK(�n0`��P�9K���atU7e�������4 `�`]c%���c1s�������j���d�0�P��ͩ͡X)�f`�#=q��V0��X�h�o�������M��U@7Kd��yQ�w���6��j��6�d���ZO�Y�l���F@�s�X"������ �ف��$��V2\r��.Y������%G��3:�'Y��,�Ӗb{�@n�6X)�Ur�)[;���]���� ���[�a&�]e�f�('���z�S��*�0�+�z�	>L���0p(]>~�:XG�0IS�A&:iN�8��v�C�'A�E�gְ��&\�60��a��"�ܤ�sc�a��PC�ts�kj±c�fb�Yi3nCE���S�+̊� �9�,)�k��@�1�-Sa��Ps�Ɛtxz,mX�5�7i�,@� d�@�Q�@�R��!��QB?��Z��"K1I9��XfTqWBY1�5SQA�����}.�d2@������*Q$&�U~[�VxCGP# �*�FQ����0���������!1p�5��$����36�k��`Lc�Jᢦ��8���Y��a����=aO<B��W�Պ���Y�C�yi1�M3�[ݱ�J;��B�P�i���mXBa  �8K�>F� �.c0��n�(��T7��L��d�B�'\��8��$
N�xa���"�$�"6��'\��b�������n���zV�t��$�: �8Ѡ(8�u�����TG$D��4j�j�6���Ʈ(�	�ʛ����
Pʍ�����С�10C6��I�aE��'1�I3��@U24VE �54>�C�1�\� �PƄ V1@3��P"�ԋ�/�b�,gX��`{_a1WaD�cE�:^����K�L��fz8)H��,(��<7H�.Z���D'A��fl��&���j����[�[����@(�Q�f�yq��L(�Р6l�0����hw�gmF� �b,�4C�)�S�(������f��w�0Q�&��y�S�~0@I0Xtǁ���5H{Q��M�o8�%3�Tc�	1P�R��1`>Rf�!S̄�Ի�2�x12�~����X��ŋ�S�(��0, ��p��B@����b�V�82`<�(
�P(�`}��L�z1Z�ǂ�0@��Cax�`��IG�����3l�/ �lv�E�5-�V0@�uҙӥnTY���E1`�Q��~6��E	[���\����r�e�<mLU@�Q՜G�11P90c��XtVk�Y��la��(rdTt0�c.icIĕ�������vC1�`�49hxM:�����" ��!�j(`#7d��l�H�z:���T�vH���_�fQ;�h@��w��|��1��ڂ�Q��q�n%���#jc��W�G"�PjBUO[8Mg]C�1*!��O�dyE�Y�`d�扳Ø#�?��ѽ���q�]�F�6��\���Nf��NFY�%4��N#Z	UƜ�T�4+�9�b�z/��B�+h0��������b6Q,�����/���'(6�
�c��d�$|"��>��P�v�Q���5W�
���>I�h�Jae�r�lc�6mX�=þ�IPE��t�^��0�To;X�"W������b2 �]��Bm��c4�_����������(���9�����i��8�:�������φ0�c�-.;�a̬�0����NwK��cN���M�1FT�rG�i�DX�	���aPk\[E+U1f���r:�a��ׄ4'l���M�)a�3jfK��(C2آ�c�:�K���F6a�VA�Ɓy��7VѰ=1a&�4�L�B�?+ �:�0����@0�N�b)�����X����o�Ƞ�[�Q2��R��~P�TEL<���6y��
 ����r٩���L�&����	������ ;v(X��qP�\¡���ʘ�2d���/!�  #�=@���������ͪH��b;l#�E�����T��&	X�*h����IY�^2��H[ѕV�a�@T�޹}�A� �Y�C�YV��0{x�v���&��.+�d@8(O~�a��m��b�s�<��TS������"ވ��������	���+� P�Vpx�e��)��쮺��}�k��^�~�GT�G��G�~G�~d�~���GG�~��~��~t�G��G��G�~����BnQ������������Ѫ��������ѯ������������0�؏BԏH�����T�����Տ�ՏV׏���~��������ߏ�Տ@�(��Y�������ռ�cU�^��Rx��`@�R?">�w�"��P�R?�q�\�T�G��w�|�]L*el���r�B�"��a�G���a0i�C�Q�h��}��`�?3pY�'H�03xV~8<�1@��Ac0f	�MW�u�0�S`��r-;�÷C[�Lڵ�0���E�|E 	�n�FӀ��Ӧ��}I�r�+J�Ch_�q��έ���i���j��}bU����Ki�s�8F10q&�2���}�_�4E#0��H�_C��Q]�����F٫�E��F����{+1��1-� f�͡��4�K�1�b9ņZڳl��n҄�y�HԕQ)�%���¬`���M�C[̛Y�k��Hgu�����όvM��4�[�� �*�RQ6�ޕR�� ��Ye	k>]m�0̐V�JP%���]�(���J*	��q�hJ\%�/a�\Yd	�D`%����JH����^����J�%�.єTQ4��N	3ȐT�XJT%�'A���/�N�����q_h����7B]4��݅��pׂCe�l��������[�8���K�,rq�iy��r3� �ZTb.Q�	]]� ��%�ZBc��x%����J�VA+	ҪbD֋�L# �ᔈJ�R�)I	�J%�(1�(��_"��%�v��K�Z�-�͘�� � !� GVV�+m�e��Y� �!@b*Q����T%�N�0J D"(1�S�RK�%�.Q���D\b�n�XK�%"-��	�Z%�d��J�Vb+���U	�JH%�)ᔀ*�R�	�R%�D�!��]"s����%�іxKZb-q[��!��+э ��U"�
Q	C�'38ei� ��
�C�"_"Dj�z	�K�%�.1����["��Z*��0(�')�v`KP`fU��NX�YW��V�]��Ъ�ipAf�Z�r@k>*w�����\p�y�Ac�u4�I_�h+V�Յ\�`p��Ka
X��]b�"�� �*I`\c]C@q0`l�<��`�V%�9#f����$��<gx�5�V��bҊ��[h+C��́��� ��Ew:��
��7����\�f�օ$���ˈ� �
 ����Jt�ilq ]�ل2�D@^�ԋҔP �pЎ~$�3\�CW���qeč;�͙�F��P*\ ��8#���#2��ץ��᷍��[�eY>��7�bT�	��Y"Wŀ%�.#�vLXs�P���.7�H�W�F��&��];#&�����(w���4�zB�\��ܪcdو�(�A`(��'J\�w0 �.wc�`���f*�b!� ��$N����1�3��$�1�L�0�������!@(L*�2b`?�%:���*20 ;vFQ�v�3g�tun�%T3����M�WW�d@"(��B���车<�0���t%n#��Y�E*���o�Vb���L��9�̆�����优l��<���X&��3N�8j3��\��ߥ�4C������Ċ�B0]���&$hRs�l~��BS�6�;Q��0����>Z�T�����p�PU���j�r�h5�ӫ�@�U�x��ͭ+اc�+j<���-�����l�b�<�x;���	`�x����B�&��1����� �t��S��A��3ǎ?<졯�|�V|��OV!P4 Q��}:h@���]ZiQ�.`{�|z���X�2��h��i)A9	�#a���
�:ȁ(�x��#����eə�:��n�7���7�h�~���C�KQ68؟
�^I��?|��*����q^G�ul+�-
�#�FkQXS���+�*�rW%OT�l��v��ņ��my���c��f![��Ĵ�{�'�v,�;��K��!����� �
N2d>L>_(P�� VZW9���X��~���������
�P�b6Y�(�Ō*��V����(�[��W�Q�%A�]��J��'�
*�$H�Ӫ��c]��L��>�}.;b�r6.HV?�˛�"):I��)����n��ރ�u�3�.sd�>�g�+ȱl�@&�'$5*;�t@d����_^���A��	0�N��)�=s���]�dg�L���F.:�O��$���h;��Q��d�����0w+f a�XX��R�-�7�aX�K��~�9�X��ː�nR�-��ÊC���iͺZ�SGP~�Ec��M(29�����ya�W�boYz�XD�ի��L����CK�ڳ��	6���L�
L��Cf���^�M�IE����$�h��ˌN}4�2�4�Y��$�-[�eН���D���vU2	P�N����fl��*&�'���NE[�ye��ܒZ^KҶm�<	�(�p�Q4�V� ��c1i4ܼ���P���4d�e�f��E</��e�r	*�P|�v�"���M������~����04�CZ���2�Pb�z�Z��dWJ%cbۖ�lZ�m	�l.��MK��_�x�xY\�,������ɔ�j%�
L�+{��_|�Ȥ���S��Յ#���� a
�aJv��B��rw�PuٝY�X�y�&��2�R�^��̜�GJb_V���J�3<b���QP��3Ct���TF�c)LƧ3vP0�1+���J{l�$�F�%m(:v����V�Jiy�r��hvY�zp�׿�R,�^tt�,�,  }��{}���h��lFA�RE�ܬr_/������Y���	�+p΋Qr�������}�1c��������46~���~�ȩ�0�a\eL˰��ھ|N��w�D���3捂�����y 6|���3bb0Y �每����`&���1�J�8ŕ���*���T���Z���=z9��*q��J-���Y�;0�HU1Jd��aEC���zF�*�7�ξ¦��{b�����1��=��0^��,�t�tg�u#���lHE��]�a����ֻD�{j�zA�Dͅ�Sׇ�k㾸(�6Mp�:a0���P�'�E8�>_�}U�2Q���H7�E�G��J�rV8-Bp8w��a��X50��`��f�(T%�#Èaʂ�;u�ì���J!��*�j
We}�q��6�X�2�rNy8G;��0?��Q3�a��	2c_��ru�BcL�g��ƾ��AI�e��c�,����ƾ��cK��̊D${If���0X�����9;�_�1L��V�tv��r�6�c�����.�e��_��ҭ*�J�a��(�0W&��c�\K��4p��9��+xr�,��N�(�ow�����r�Kkg��
7��B7�P
�e8f̍��)a�W�������W�߾)����W�\��������3WeGET�E���r����\]�_����'`��ś�K�$�Q8��zW��Q���E��,�H�N�g#]u^�,
�?Uya�@�N�<G8>F2\�H_�ϗ�0n�ϖ�TL�X.B�9#n֞s^�4O�n
||��U12�����b旽�ܪ)7NW.Fy�$x�5��T��ɛ1�eL�\�:iw��J�ϲ�p�+k�讕�e��ꏚ/F���:��1~�00�>�]%1�$���CAQ>�?��n��L��Ŗ��(NV8��&��3�dkwcԓY���<���,]M+����f�_6���(پ�hu�38��	ۣy�g!�s@9z*�����09i�j��Yr��/�=|�l`����1��m}2�a��=�`�#Wq;�h��s� �4ϼeQ��Q�"W`C�хet(�-ɬ��`ܯdV��Î�p�fK���0*���W�Q,�s��fq���9�Nê����9i��Ħ���wt��QO���˂�
��Ĭ2Nh]E*E�\���jD壢dw���Ɛ�v�Xɷ��w�83���q�
0��.��;�V��x��P���\������`a���r��� ���.��3�w�ҔS2��8�:�`R{FgJ,�ح���p�Z8�*׳��ga�JB���u����ɕd�q���B3��<]���G�\����>V�0��0U���L'u���C����B�UA0�_�W\����RW�T�&�_E5��͛��\���QP������SU6d��Ϯ�sʯmu֦�0X;èx��R�&	D�]��[ﬗ�Y�	�Q��ȥ��8�ql�Y����i�T䌌�b�T4C��֕sf0340#g7�,sΆ�����3�hJ�[W����W�?x�����cG=�����}�8 �3N�_Ի*�1��Q�����^(�$P��W���y�%?�����T�SU ō�,E=�����dUaQʣi�e���p�F^1s�z;�ow�k��n�v*�i�[]��M:�񓴊�d��FS�;��J�.d�5f[��Ne�|lY\��ǋ2����^����4^��t���]XT��r�>?p"�1,w�)�G2i�,i\G�99���+ζiHf.ZԢ�0��0�x��r�l��\޳<Pf����J��nr�9�"��Y�BW��v��C�'K~q0�V��j�N]�SX��n���>U�Y��ܥ��կ�"`�>�����/»�y������Aw���8�Ĵ���.�#0�7�2�>^��&�Y�����>��'إ�)Ŧ,žQ�`� ?"W�t����	�B_qhV&�����蹔]�$ Y�UƘ_�OL�5P��N��"� 	�|W��?���À١�H/�B}�!p�V�{Xb�4f�`�Lo����c�/Br9,B���:��Ʌ���-èwe�O�l<ϳ�i��"$�fd���� ��	�љ0���$��:��v�K�X@@WC�w	h�y���� `֪ ?�-�M$>M�M#��U�SQpN����a�@���~�"�b4v�ޟ�Z�]�v ���QQ���̣I���a>/��s0����D	Q��q��o��g1�3%�,�ƨ8�{�<%�(�p�?��X|�ٜC�
U9@� p��Q��uO>N��q�S%�9�������]m�Pc��U�������W�`�b:qZ�m� )HzW�����9dp(�VeGa����0&a����s�i�Nc�$99F���2�Ռ�Y�)�E oj���)ࡎ\ �0��L�Z�5�����  �T��c1103ab'�.�#~���1���;����K��� �1xXQ��ce���~,G#,�,�Ed� ��O��Ľ*�\#@Fi����+D��VY
L�=c�^�������3������O�*q�9��Z�>M`�������!u���3B�Q�㖠�#�x��6~"@ANL�
/�%3A�^~[0[�����]1/�*_H�B�A����3.v��O�L�� �~Y�ċ�S������43 ��EG'xUU�u��0R�.�Ū xS-��>+0�g7�FAZ\I�%kc����٧���2 �Y�@���>�pGᅘƌ�`	�,�}�`q���5��z�QL:
�ʬ]Ց�L��/`S7��	�˨X�Q"`x
C,V���e�eL"�cf1%�"`����)e��`���S��?�yr�ͅ�G���@6�F�H`I̥`1'�1�E��
��(�"�
���Zy/a�V�z^�Y��,��s�O��3��� ��luQx\d1���,��q10�م�|��1wP�>U�`�������Q��1��>��v1@m���Ez�F@��F�;{ I_ϒ+λ�e�ƞ	�.��RRW�T򎔇%��hexe��������4 2��V�����^�d5;��At<��)�V��R�9�q�]�1f�m�rk����cgG���S1$��Q�{`��o����s8�1��3�̅h/kb_�@�J<@�-�����7�,�?"������E�=u1u)t�D z5�1��I�S��C������p���#l�>��#Ific��"_%��REjuY��d��~�݀�hW�W/�*뚏�,�	�r��ۚ�>`�.���ü��_�-�����|u���s����/�֌���O�K�ď���(��
��Y0[�&��6� ���h4�]���]�EwS1��1�yܬ��9G�K8�W4M㾩ީ+���DI���42��`�a
��)]Q
�a��ٌ9���qm\��g*
�dy�5d1�N-%K�c��Q�u��ů⽱��<,���f�Qg��x����k6~��0h��5���T��Uo[��b��c�
%��(��JU�f:���@sA�xEw�
t[T'!Y+^1;^����(�r�svUw
����.
���(���U�	k�%�T�hJ<Q")�C����%�K�!�.a�ȷD\��m�8K�%B,A����W%�[��J\S�)!I��D%��J/����^B�s	hK�%"-��	��Y%�a��JtT�*�N	�� %�1�0J�_"(���v��-Q$���Z%�g�K�V�+�U	��<%���`JDQ�(7���{�K�%�-ᖉ��Z%�e� K�Vb+�S	�<%���hJDQ)A����o��K�%�.a�	�D\%�l� K�W,!Z	��X%���JS�)H	�J%�z�b/ч��D^'�u%�p�PK�Y�,�`	�p%����J�T�*O��J,%�(q�H�DP��>ě%�z��K�h	�D�%��K�V�+V	�JH%�)��x��QB�C����%��K�\�.qm	���%�!�(KW�+X��JL%�)ᔈ��R��F	�H%ҍ_x	��%��%�N��`K�Y-a��Jp%�*��ЩUQ�XJ4%�(��	�Q��K���CD]/q��K�%�,a�H�DXb�\��JT%�)����R%�G_�Hw	�K�%�-��x�ZB�d	�J�%B+��	�V%�S�hJ<Q)�B	���"/��n��]B�q	PK�%�,��	�Y%�`��JlT�*qN	�� %�A�0JRDB(��m��K�%b.Q���\%�j� K�W�+!X	�L%��J�R�)F	�K%��C��.q�	��\%�m�0K�W",A[���T%���J�R�)G��H%���_�	�%�x��K�k�"�%�� KW�+X	�JL%�)є���QB"C��f�^�/�u	���%���pK�Y-a��Jt%�*��Ш�T��M	0J %B(A���_x	��%�ᖈKDZ�-d	�J�%�+����U"�R	`J8%�(����DQl�A�%�Pq��K�\�.o��K�%�,a�H�DXb�[	�JX%�)�	�S%�G_�H��x	�K�%�"��j�(K�%,1����W%�X��JPR�)�F���%�C��K.���D]��p�HK�%�,��	�Y%�`��JpU�*�P	�0%���PJ�P�(>䚿�z	�K�%�-񖉴�Z%�g� K�Vb+�T	�D@%���pJRB)D	�/E$����	��^%�v�xK�ZB-�d	��%����J�U"+R	�J8%�(��`��Q�"B	�X�]B/�r	�Ĵ%�DZ�Hd��J|%�+��誄U�R	`J8%)����DQj�B�%��1��K�[.j	�K�%�+���V��W�xJH%B)є��R�"B��T�D]/q��K�%�,q�H�Y¸_��Jh%B*A����S%�J�J��/�^�u	�K�%�-��p��Y"�b��Jt%�*����DU%�P�@J(Pb(a���Dz	>K�%�-����Z��f	�J�%b+ѕ��DV%�U�pJ@Q")�C����%�K���.��غ�]��r�HK�%�,q����X%�`��JpT�*�N	��(%�a�@JDP�(>d��z	�K�%�-�	��Z%�e��J|U�*�N��$%�Q�8JRDB(�Pi��K�%B.A�	�\%�l�(K�W,1Y��DT%���JDS�)I	�J%���	>D%�z��K�[.!h��D�%�� K�V�+V	�JD%�)єx�DRb"C��Fӗ]"/�s��ĸ%���`K�Y-a	�Jt%�+��ت�U�S�XJ4%�(����DQh�A�%��Q��KD\b.m��K�%�,1�(��W�Y	�JP%�)�	�R%�D������K]�.p	�K�%�,��X�Yº`	�Jl%�*q�	��T%�M�(J_"(1D�y��K�%�-ᖈ��Z� K�%,!�	��W%�Y��JTR�)G���%��_�H����w�xK�%B-�����Y%�c��JtU�*�N��%�!� Jy�/�D^��u�xK�%B-і���Y%�d��J|U+�R	��4%���XJQ�(K	��C���.�����\%�n�@K�X�,a\���`%�A��JTB*L	�J%�"1�(�3~)%�|��K�[.!j	���%�� KW�+X	�JH%�)ᔀ��R��E��/E$^bmq	��%�q�PKDX�,[	�JX%�*!���DS�I�J%�/�^�iu����%�іxKDZb-c	�Jx%�+��੄U�R�PJ8%�(��	�Q��K���C�]/r	�K�%�-��h��Y"�b	�Jx%�*���ͫUڹwߎ�{���0�\uA�,�6�Wo�l-�`mX�#a�f�0@0���j�*`�t ��q>+Pݬ�k-oq��$0@l@b6.�pe$sG�CF � ,��bAREa.3�Q���6�
4Kl��Fx�c�k��\�*�pA/d!�J>�-���Olb!D<Đjl��$�V�{6-,1B�B����Kk�䅊ŀU��i#�ֆd��`>@��9�@=�"�g�A������Oٕ� ��%��)W,l���k���I<a-w�aVv�awcKPe �Qb�:�a�*΢a�x�`$n�:�@.�!@.�� �ĸ�-��pQ�j
0̸ڊ3�A:��2��H��E[��h�.	��8i �8�q��1���t��	��A� e1q�מ`��1=�����J�1��`X�F��{�AL�$$�@�^��>�1��X6F��!�į0�L|�k]�䥵C��4����t��iL�Xx}�( ^y]�������P|@�|����+ct�|���;#�*�6����`/Y(�R@�(T�Ԑ����}�!@hk,"0���7t1�{�@�xh֡���£_�x]�ǈ��2'�@X?^_[�9H�X�v��è�r�@����+��tEF$9��u��]x�7�ҝ���0,<#����L��[�i��%a���	5^�0*� `)�t����+�d���Y�!V ����A'\��>�=NT&��>!����Q�'�G(�*F�|M* `t��>�;0�u�-���D�;�J��^�{�bb��(X���F�����[�e �S��>u�h1����PĆU*3,I����03������,ϭ$���V��k���C��-+��1���(��ȫ��6�CV�����
� 3E�CX�ٳPW3yM�"�)(� �wc�00o��܌&��h�"B�5&��\F���|p�� ��Nx��1������W������ �8��[{���;�n�{)0N�:��D'(X��L{� p�ـ��i
a��
���RW*��h|�=�"J<�\��"�	k��&�����@`��
zAO��֮�_�!K��鎚�Wf����KL��ۋ0ʖ�e���&����!@� �w��9P`Lf s@�*A�9(����U��#��n�" #���AAB�S�� &.�F^?P�@b)����A�N�db@���$��6��b�(#U�=cg"���1�fҌ$�305J�� �
EOt���/���9�`bEUe���3]`eRt
(B�t��@��_�&b`"��!j�� �n���c���<S�qd:0~�S=� @YaSe�A�0B��u�E�	X @`Rq�i�0!`1@�G �P�p� @4��ab@����c�d���L6LTâp<*�|#�{71lH\�q>�$e�/�^!�[;�A�����Ժ�h7P�Hv�e !Ņ����ŠQ��0&(��(	��AQ�C� �h1?���RW�C� ����:�4�8�a꣄ Vm�|yLʬH�]�X� `&�Ej�=�RzG_T�(
�{M�N �#A>��C��� \�"�g��2U��@��\@�J灱 ��h�dA����5��"@Ā=h�A4ۮC�P����A�p�z��
�h�D@�gYF����g,�H�ue@�%>/�p��_�F�ꄒ\DS�ӈY�`h,�r�W�BG�;�30��|B����0�<�ÍALleP��ј~��30V8��({����@y��B��4���7�����3�;�.+o�)r���a@�̂�ؑ��}�薣b�-���.���`\���E_l(����PY:P�a! Y5�?����F	H��}I8O��0��8ށ�)��g��2��6�����C�b `�-L����|A����<�C��-LƢ)Y����+C9k�q�}��H�u陽���"!���CgaS�&�G<:TzE�y��S�1�p�A��~���t�2�X�c#T9�!�,U�!����[6��0!�-} cq�\m5�j�nb��Fd�!�.%A:�S��	��F@� ʒ��Q���"@�,L0��G�Y�'��L�*���,@+pE&��4x�MA@p������g�8�0�� ��P����As�>w���I��8��5}��>,�8 Luo1�������3̌ddǾ8L2���2����b�02 g�3�:@�����عۺ%`b0�� �X9'MA=�b��,���D ��M� K����D1	mXaS��Y2R� `@�;��2��f<}Q��9(	 ����:��OJ|
��`g$��qO�^N��+1 �(t!`�0�qF8Qd��cq>��zl���3�q��[���8pFV�?u��r��0����q���E��u�<���T�As�����tp���-#��1n�4��B+�X�+rk�L�L� �%���8Pr參�Lˀ�f��@�gjCř.X����Y��f� �F�Y��3̀^o��! ���4V���l�`^e�1BVP�\~0���]H>�A���^��A�@�at�7�����t�(�o|�}!�c$k&�w�N�a��S� ��~˒��Ӛ���N�P/R�q"``�"@�Pl@�U�@}̀IyX{�B98��2bfXDa������{ �bq�!k��������3'&ɧ2Th')����B���@�J�y�~�`^޽ؙ�G��̶�8����A��D���Q�Dy�&�@"(0OF��+�)?�w0@���B�B�$�a�� X��`�Ӂ��- �0��l�K`�a9̷a����� Fus'�R @P� `�=Cye�]�`�XK��k"���r1`F -� ��ԗ��P"(Z�1�8+�4��C����Il�C$� �A�`(����'	�Ȉq���=�_9f1q�/�0."��͉�zF��b �$�]@�ޕaf�!�
����)(bȿB�%	O�h������b @VI��MH���`�X�3r`2�BM΢�ǀo;h����<�	L�L�Ib���+��k� `�&#��w&�.0p,�O8�yw�807L�d��ӱ���E�ׁ!��,�2U�@U`�
	�RGq0`	�*��1��a��2���s�3��%B�Ĥ�B�(�!�pF���Y�n�w0�d���STv�2�A@[(K��>�*��lH@�l�X�]f<���Z��+*C^�C�(X�3��� 1@�RU��4dJȅ�YǙV�`��!��CeM����B g�A����+����d�x�Z�>0�Ѐ�81�
�ư�<tZ���O��A��끀�͸������c��W�"�-b@Q,������٘����r
JL�G w{���vȘ%*t�KB@��ϴ������A��A�;����H0U�|d�=�@L`�� <[@a��!@�XF�y�L*d��Q�D��A�� 6ra�@�����[8H�ɐM^���f�X�
0u ������2�, #��j=�-�.��̀oq�zL�H} `����0-.�
iI�.$j��,Hc� �B�qJ��f��y^�yH�̀!ȱ��gځ�pg��M.#<��ɀE�́� sd�h��9Qŀ��w���T�UB0��zL�Vl�"&,Mlj0�� ��=��-}@OhZ }�DK��cER���o.*�^.H�=|
hL�q��ޙAkV��Ѐ�ߖ8|���$�+};��h@n���J�V�T�T�M VhlBu�������K�N
,#.�F�j6.����:����)��'2���ؘ0.C5�u{�]X`�b�j���Ӽ�ڭ���b� ����9H6�@�c�9
-�(0�@��2��_T�0�&E�9��F����?k�L>u�^ 8
P�t�i��+��DS*[ɋhy!@8+C�j�B@�T���{ݪ;�I���DLj+�AiO+x��u�t�'�K.��wb�� ]�F��2�>h�`�+ϯdp��s=4��`�*��v�����"eO�f����x�y�c�"��c�D`���詉� �2��vx_}͖�P�8�$�8�J��A���|�Av^ǔO�2�*>��%a^+�2ǨF@���L��C@l���X�!dF-��8v ���3�3��d�Z�~�)H�A�+-c�R�,.��|`غ#*�},�,ٗ���>�_�e�*�q*m*����%��7�D�!,z�Lb\0�x8)�q���%��1��`	��{��cX�
cOҹ�Ju����SZ�����/�!��Ո��vK��?x  �e�j�2G� �x��f� -
I*+`�a8�CDY��4L'}}���0 ��FM���
k�E�B����ϜZ��HN4=z`��
7�y铇�D���;B�@}P�t�7;����|�%F�`�&��V!�7O�JJ<\���L�x�@�@`�+`B��e�>VX�2$@���%{�U�G��b?�����@%x�i�!� 9��T&�V`�+%�1a`ƀ���%P�����&��.�%?L#�W�5�/.�D�Pm�>��0�E`�BjX'�SSa�u"`��m�m]H��f�Q^ Sf��⍇))�2�`�� bB���I��Al,��ÊJ�c��`�_�B�|{TX��1����Q����R��w�r��q�ª2�/�b����!)���Ȋw�:��T&���'��[���j*�`�@+\���g�QY0r�������C�ؘ`���aj bЪ�̸p3��H��������d"��jX.� 9r1���D� �`e�˅�1���r=�˿w�� e�� �� MG����#���e�V���̼�4�l�F@�B]B����H�#F�#�W)XD0,�B挘��'���:o�&v�V>���%9'r��𒄀qb���F��)���1�"����a�,`dp'�=P�q6�L�L��F��,[���V+�t���f�Q"xL��l膬���A����=�UN��ˁ�1j���pOV����.l��*�V`��n1E��S͵�E����2bAz� I>-�V��6)�q�E����s J+�-��H980z� 
��d�7/ 
�B��p��i `��g�c�����yVBCՃ e?�h6MEC�s�#+��SL�m��� e���˱������ .�� ��q Ce��Z��1P3�s�� g���T��7�����<i�Lv�vϘ7�,���B�
���g������1
�0�4_P��#0�y�UU�~��3�A����ϩ���C~�@�N��S��X���,�'�󌖑���pN=Ke(b�-EZ�&�VO��8t�*Cf�@�6���Ø4��˅(�{9X��x4U�p����3�@�h�uF�]c���� ��2���}-)NF%+�����:��U~�DV9������>z�8�!t(#]@�6.=�L�DL�3��=���;�Z��2_j!#�k|e`h�H�_F�ǻ��Ke�T�hS)�?��Nʘ��豪�����#�ʇ��\QV���Wg$ u�TE�E�hXJ0���2�U'Q��+*  B� ��t�'�:�9ԍ�|
�����i�c�\�/����Yt_TfE�}y��L-/�	C�Z�ͥ	�h.=����?p�%��������+l��A��>Ġ���[�]�eE�M�q��F�����	��j++kZ�Q1������<�H0.0QϘ/�o]Q�|'[g͠K��W�c�$��;R�3;9�d�����F���TF�f�.,B�g�>*�l`�·26ʲM���,��b5�Ө1练w/Ws	�G���W>��ݑ�^�Q��1F��1���a�`�#�^Hцyx�̓Y�W�UQQ����]�搾��B��_T)JK�����ʸ��D�z�Ϗ�s+r�M8������ma`��,��g�@�]1�=B�Q��p _Jc�SxbQ^��Ej�S@��f����6��a���NL���Fw �-�&B��_�2�W�ӵ�W�U���%��we|(i[�2�E�����(����	?��b��u+�T����|b��1UϿn�j��+�*���T?�*�[�xa�W��7��\�9�t��e�`�at+`�A�yV�^Թ�jt�~@Wi�n̓�D��bu(��˛�)� ���98�?R��;0�a�a�H���p~%
���'ܪ��96�����։�Ue������&��@�T`ewy=c��sX^'�_Yf��'^�0�x����ӐA�2�!���u��e�ᝥ`�O�x��Gm�1`ڮE�1n�B �}�)~Ǖ.]i�d�D�vGi6!T�Sa�����β�P�#2��#%�V��W��;&�"�:Ư޷>�#(���}�>T�޻޷>��i0)�*B0�NۇϾ�$s\e7�G�9z]\���q���^�AA"��<��>0�}��\��A~����[�:���6��#�3c#���:�������'�w̥UE��r?+�(
����3��L�Vи�0�;J��P�����T�0[_����e�k��v�[�?yw�mȞ$���2�n��Y�t�Em��js�	 "��%��(�ɂ�`g ��.wZu���kb"1��e0@���(���w�}��l�}�Vb�_�(3��}��*:����&�b��@M��B �AKߗ&�##b�OX����R0Eծ��г!�,�8=HZW0X��j�����ҡA�s`�%��F��GjW '��a'� `W0Xmd�)�!/��)�8�:A_h 1k��@x��W���̉��اsL(?x�o�.�"��Pگ�zE0��E��G�m�D�(�=� �E�" ����t�a��O�P�`�����? ������^����H:´��>�zI>Jग़(a�)�]%�r�J�[z(�j	����q�<J�Y�(e	�J�%�(���W��]�"Jl��(��ɢ�U��U�DJLT)!P��DI������ ���%���l�
�0擯"���������"ޣ�����,���U�h����a4�Ēȶ�*�2g�#��)tJ(�ʁ�<�E����R``�p�*�W�м*�U5$jK�5�E4 �!U�U���5�UeƘ�"^�BīyH��h�XB��(����]
=��8N��d�0�S�^U���<��Cb�tZ8����`�� F-�d*R׆p
�Ql!ى�Ԕ{d�;!���c�G�=M�H�Q�������(c��$Z �fB����(d�l [������e��m��Z����nn�S�A [(��hy%�Bh�K/���RS� ������E�3�]�U(� Z�W�sk��uW�f�2H�fjJ��P��j�4�l�dx(�����Th�(5*TH�?#Fu��j��rޑ�ῌ*
�1Wy�J+aF��,����Gd��1ɡ�F L����Q:�#����%����K�2nl��
� r���g����jCI�S$�>E̖�I��L}�1�oC�t�s���t�p{���pk�\�5�B�c���g|�Xq;�״�u�t8���)
�w��'n���u��N���tx?&7��C�����hr���������7�y(_�p�{G�;��U���͇>��v~�RJ�&W}"�[\�~��O�����ܟ��z�g^���#��k��]�=�b8p�"Mn4y�X��9�{ٸk��gj)޳k���C1��Jdh����
��7Ѻ����>����㯬���'縻��3u1�˛��*P�u%� ̛K�O ��=�� w�u���}'Yn/7~��`�e9}x��3���E>�މƣ�G�8���q�im�ٻ�kv��P�=g�^^���SI�H8�s��ߍӗ�o~+ʔ}r'���sjF���ך?Y�Y�[�I����H���-��1w�JG��<k�|��z��n6~��aɾ ��b��H�$%gT���Ь�nK�7�ݡ�w�ϪG27���T��u꧴�X�Y�9z�<�3�#�/����7"Ċ�x���h�B�67��]n�Ycܙ:�)������tN���}����/���e�����!��J|Ғ,Ҵْs�S��1g���&�_��{4�~V��=���������)Fg��-e����/��g�D.�*즕�V��O��-k5�w�(��WY~_�r����0=@W���@���Y�*(f+_����8��+G{�W�g$B �   @      I JC       �� ��HЎ�aPB��F�]K�l)nB֥̣H��۔n���y��Q���)Wl�
4��"�$�3�-��EBE�1�]AZ�i�R�غt=`�m�d0 ���Kp#"-Q� �0LV�[�4�T�r6li�}+��Ӥ#�H%�� � �D�         I JCX2     ^(� ��-zK����T���n�a�@$b��C��xk�ۢ�0�x/&��
��9o��W�/�����mJL�0�\ #/�ֶ4��L}"���B����:���zE~���]�Ƴ�Q������ۨ�H���̣2}�Z���@h�C������!M)"����"aG6T6��|l)Ƒ'~τJ��	�.��{ v~�]o
�I�"��D.�ST���ݘka+��fa��h���R�g�Rp��j�o�k_�k�轋\*���$n��p:j�e�J��@7�w�+5��y5t�iGF����)�4�V���:]:�_2P>\��,�>G+o�PE�(<�V����ts�jG3���{y�������(~tM��M��r����,�OJ�a��/��)�J�����N�� )�����vʽ1<7_L�tk���h�,��&`�����M�mS$��DY��ݺ�P�����"�P#@I
��%{�� y����ך(*��[����
�g��]���D�4�O��%cje�>>�n\���$j�|������ucK�g,5�l�z`ڠ�5u�%���T���70Uw�' �2H�~�����P'|vZI���QEkU��(w�N�גt�D���I�ٵ�@���P�Яc���B�Ek�	�+�����R��^L4~��܇���򋩇���8+I�Ƭ؄����>W�R�+#ą,V��zS�s�F�h
�-�,#�L5;a��>�c��PuB�W��c��-��`PF,�����0!��OA|-���%:#Z#������7�H����ܳ<�yG����@�Уߌ�����\�E��hr�1��w�������CH���䷅��ݨ�g�g��3���b�=�XC�b�G/O�HQ-)�����&q���T̒uX8�E�5���$8��_�(�I_2�R�Ҫ�f"���d ��P%aE�P���*uȉ��2���]2�F��1J ��(o��\�Zڬ��bq-�!ǉ���{+8�_\��>q|�F�����B�ԟsiR6>#� X"�ux�.�^G���L��x�J8�F�&F
�������'�C����	��?4�[_�Io�D!�nz�Z"�5��み���,�r|)|��+nIԩ<8�s7(Z��аdx�K�)�V���dNm�V?˞T�D:���o�M6m�=p{����[�5��5v@�S�rZ�g��闛(2���S�������+4��<�mi�l�e��X+�� R��2��_���2Z��=b����u��J�h�j��~\[���lP�.&�P�p0j�@/X n�(E|c�RA$h��5 �6'`gr!��AR���MY�.�?l�R��,eRA���i;v��� <!�R�7<0X[��,(��Kc-(Jw� bǭ��V^���п��
 }�h��w���gp���q��.ab2K�ZÀ�R%�M���>4Z�	�Դ��������{T�$-��*-ح��t��V�es���*��ع�"�}𡔁�i�%,�ȵi�ںĚ�o�8���J�*�⋟B6�����뗤/���f������y� ��\�F6���ݾK���R����"�����4�4��B��(�\ّ���2G��u=7�D8��Ugw{�H�̪HX?�X�5����*���J��i�/u�<��QR��2f�E �� Q�bL�e��!�n��i��A�aᝏF��f[���TX�VC�?����,N:���~8�~Xg_D<�^�<��K3�½����{��+UVAz|���X�r0��0h�Q�z`�d.�L���G8���<8E�ڸ=䜓�=��)֒�j�a�(x)Z~1�[G��{��&f���O�Y�|P��@V��-'̽3�H�8>�a �8����1�"��񺍏
ټ�I�5l�j���n����  R��G�fB��0Sm����0wx�k#_�[����� $ ��g#��n���lsΉ��%>S�љ��K�їJ�5�����ߧ���OD���m7-8bIʰ����cL�[��0��o���z+�/j\�y��'�t�RםJ�Ώ٣xk�u��_�J�s ��/&L���d�WC���EQ��s��E|'��I���4Gr[���%�`�[d�}�_���U���a���AH(>Щ�ph�ؼ�1�rNU�יF�Q�T+�t1����_{Z�E)㇡�L�z���a�@�YlPۨ�ǌ�l���9�W"�T���!\28��%���m�r���`��@A�TL5�Tb�F����\�Y��
=���8)��5xȂ\N��%�mé����0��n�=�h%�_�Slk�R�ǒ܂���[�_N��i�4��zq9'�˄�5��xi�&���6�HݯėV����p �5��B)ck� �l.���i���y)�B�PF�z����]��Y�,��za�M)Zր��l��I�hBTW�~{�(Okcd[!��u���d��@e�O�]�g�]�h��>,Fx{������Q�ms�x����u܋n��R��0�_x����ܞ�̲���h��I��G�6�D=J,�7}�� �����Z�����ōI]S�������V�O�������vq��*����a�<z��-���Y��cvU��'�b0�v,��Ow��Rf��s0}��Z�+H�7�}���x�����?�We
��
02@��Fj�۵����w�"��߹�I	q��- ��Z�|�N��m��tqT��A$a��Q��?QY�/f��[%��Bmxr)1�:�e�T�:�L��p:v�GWϧ�ͻ�N4Ԑ��pq�������Q|WR����f �}��p*N.gY��?Q@�
O�5��7сǳ��;u��r�#Gπ^��� ��������C���=�^e�w�Bޝ�J<�3�O��h�ʍh�ߏ�X��<�����<�f�ґ�;3��D`���f��+b��E(�Uw&Bx���	7n����R25���d���*|o���/YJ�~����g[K���db g%"���h�����k���_���`�(f��%��X|�󴥳���y�60}��^@��/��1Qv��t��H�E�Y߮�Qvm�3�������@(sq�k�Թ�}:�����=k���r�M�Z���|��F˱���ޞ� �7�Jg���HS�F���~�#f�.Z��8���n��t+iE�:n�>2Jc��x�֬m��ʨs�N(��+@,_T���p�p��Ǎ:y�U�� k�&��Eu�B�;�[����z���}�S�b�.���Ā��.���hd8��R\7�U��±�˕h�5B�T�m�����؍
?X
��Y��dx�#g��Y�o�*R�1�2m���4(�����N+Z�"��4�� 퇙߆#�0p�B^R3�3H�n�XB��Y!$>�&���v3�9eT��2�J̇/������?�g�x;�:�\��󗅉��fϣ�L����jvN*�ĉ�ʡ�|fR�̉��@�c��S}}�e�t���i
�{7HT��ZN :q��l��ĐX<Sq��Z�8>yx��m��D��}����6�F;|T�e��(u1R���~�)�볿��l��B��d3l������dV ��6����%nbo{L��pɿuqTI����>	|��:X9*�;Շ�ɲ`�C��y�~'��Q��<6����l�.����ړ&��9��-��2|J�m��(<�ʶ5<��p��/�X)�a4���
i�I�*�����wj�w��iƅ�}��.X$>�Lo'x�1���%
K��)�@*���3���W�/�F�1qV�Ɨ(합G���I��8Qk�JW�n�z�>͐R-E	��Z�nY� a
ŭ�G_11ֹ��ņ�R��-�c��t���m:J�P*����ֽB��EV�F��y����+'����/�J����/�[܏~��M+��>n׬'�ԃ]ҙ���l*��ݬ?k���7H�D��lz[�u~<Bp��x�z��6?���h��g�~G�eQl5M�qa4]�g����+ߔ�Ci��G�8�2��{_�j��虊ѐZh��=� .��=����%n	�
����Ma���Ϲ�g�26��9,���<?v��$��X��8d���(͂3p`��2�!��/�Ĥ%������~׽f�䒗ݣ�U���J(MC�j��ړ��h��"t;w`*i�T4�d��J��+��{u�
 雸)�\8���I5��Vo��xY���4-�T�Q�q����!��@�ֈ�e�1�l@OӪ�6����t/m�!q�(�>���3L���Q$�9|o��:�LJ7�'�|Y�]u(6�>����^>"�h/��Q�ӟM�Q d��#r�ʶLQ��b��C�p�h��Aφi���Y<5�K;hu_8���>�
8w��'�>!֑�n�� ���S|WKޅ��� � �'X��>��;^��ڿ/vm�%��v�Ƒژ>�ԕ!d�����`(�~��R�R��	���c���T[%��X��3����I�q��� ��o��٢I�F+��\�E�Q})���/�ɼeo���Z�d��.�>yZn�� or���e?��(6�ODv���*)`*�
{)6��%>�츷`�>�-+�r�lV�Q;�EB�*D�q*_���TX�"�%�����b-��+B�p�f5�u�"��Ys:-�@x�q�qJ�雓�`b݂ߒ̧}�����c�PQ+�ad�	�������K|�_�v�
� �9�+�Hs�B����-s�~Nu�hw���a����������/��=���H0���U��9��-�}ڒ�UE���cH�.�h��)�5���!���?�yFZ����X2Nw(���iEj��#��*�Dw�'6m��f�h����*R��[{Z�O��ƉV��pvF?\2��zrm�	�+d�/��R7/�aN�������f_����������/CA9�u�����+ǌ��`���.���2xc��_���2�bu�Sϒh�J�b�m��4�j}����G�jtH7�d�k�m�s=J�K��A������2_;`l�|����6����]Ux�(��8J�B��Y���q4�,tJ��w��(��>�|^��	��^}�D��i$6���y�d���/eP�;��ʛt��1w���k��yq�ύ�~�~�V{���Jz{��/�&�0��j�:���tZ���Q~�<��:`#n����_�}M�8 �������ņuďs�K��2���j��:KJ���1k��h��R��N���6F���P+	%��q��+��#�fx��@�͒^�6��"d	<�3N���-��Wz�[%�/Hҷ���l̮�"��� o94�	g��$����{�f�V�{�o��T��]���>/3���*�sO�R�+���r"&�������´;��_\`EL�����D�?~<a~��Js�)�n��ܭf`zl�����'��/�&Ze�wj��M}�H�>�3�:{���8���oL|nҧО���h����H�qn�v��F ����'(��rL�W#+6�
*\]�/��b]	yR��(�R�-�cp���ŋ�)-{��;6\�y\͋|T�A�41���-��E
��+<V:UQgz�fJ��s�V����W�'G>���h�:������ ����> WϏ�Z��������<��򊿰5,�9E�~�]����f������_�M�GTwA�s��j��1���5�)m��B�/LI����Ǥ`"/?L�� g3�pM����������ܷb�/���K�TRjP��)`ܟm_��7���N��	��!eo�!����PS�'Q��Mٕ
�����V���|��4��w�F����ܰ$n��/�k[2�[d��-:K3W?h�_-��ڐ�aZm��������1����N�'�P�_@v�R��Qa�+������	_8������┈���㊐�Vqc�8E"+�JZb���:�?+�|"
�,���h@��Q!���ܴW�I v�#ޑKcK ���%r�R��1Ģ'��F�!�Z$[n-&��E�� �j`��I!�KTS�%�C��*�Q;�M[Jt�4�'���I�A+�Ͼ<�	)F$,�[�f.D߭��2��_������"���\]x�;(��=Z>(�/�&J #���#>z�Ɛ��2X),�=q?�s�ND�0��u��D�*:ͧ�N
���@���.:t�N�b�e'���nv�v׌S��xJ�Q8�����w��C����.��w�&9Z����ξ�����k2��$Rq�i�a�ƾ�Z'{A^�� ͦ�S�����bnt}��q�2�'u����hO	\�۴XpE�� Y�N���Z|��o_.:u��re	��0��漯��R�5��Ǒ�/J�t�X�	��TK��=�q��$�~�r����y���!z#����5]��I��;[ղ�Cf4ф�v9��o̴>ڂ?q�?Ĉ���:��-��>x��� ����R���?�ҵ*� �f�D�$�<�y*���*��(�zi�vR����59��s����Z�[{k �q+�ϋ?+�%���J_� k����ñ���w���	�տ�u��Sl�\ !;�r�K^n�G���m�p��0s�	>BֵS���ó��p ��A}�wTN����oȃ"���LD\1j���#ؙ
.��l�T#��"�	�.�O	_��Ğ��V:{�0DH�>L�<Mŏ|�$���MhͨnEU�����N�X�Hc�?,�J,���UBq�j���lk�9D���PV�r[�ե�"��-g��F�\�3*����]�m��j�?*�Tվ�s�Juۢ���|��q'*�{��Ϯ�N��8]�q�* K^�d#
�uD���V��a����'��ޫ}��R�]��S&�� ��i���UQ��Uރ��;����땾>�A�L��J�8�UIW�ƺǇ���4������/>*�O�-��E?+z�w�پjp�/3x`���n��\LfTuyY��vJ�TR���sڜK\�-}*�x�k���&���ף]��t�!��na�J���*����n�k�3訶��6��Ι;�V�<a�O�jQ�<��7�L�A����T=�,���G@a�pW�v��
e�bM���p�=�\�X�WH���^Ou��pz�n�=���e�C"jy$ڵ�<C�2 #M���/��kV�e�{�mL�U� �����~�a���]qc��(oe�� �)����͎��oTG����dՍ��c�cᏼ��4R�q��WW��vH��@#���H�O���Q��TdF>�oϝ)��*��Ђ_lS��Z/�!AT7'e��S���<Mzk}��Y�'�̓��j<�vcH����/�'_TX|�\�?�m���;����9R����jo��)���,~��B���]�!Kl�h7W{z1� T1$�[�C�]S4J* (Z��H|�zh�`*��6~�P"z�%����jm) $���c>Yo��Z{5�y�=�B��.��ꉉ�θ�V�*��k�B��s[��V)�m3h�w�ˠu��Y�l��q?Fָ����D�/rx�0u����ظx����h�5Hi��+���Βs��[N���~Ե�k���΅��hU�b(���z�Y�L��8"[�D�������(�'�bAӜ�`e�]��ޚ���G~,�j�1W~����O�fI����-��/f�^ZΕKRy�>F����0�ӉOH����C�^[0#B�~������z`��JKH>�~+������S�
ا�e�,E�M�>u��瀞v�L��ᡔ��[#z�6)�#�FbqL��M�l�U�jU4>�}���R�v�Z1B�V�5��Ƀ;�	�:ގХ�CR)ʀ�s�t{`�`��Q����t���\��>^/�O��T��)u�.�
Jja��Ԕqm��9-�e���F�����b��U�>Qf���<0�����Ւ�/�Gja��n>�A.t�k�U�P�lh����!{o���s��TP��:yl7���r�U��;��G�p'L�f5�Ԯ"�SE�u묝��k�˒Z� 
�#/���\�9y��SoL�Z/S�la�`�EB��F�]_���;+g����\��|���i���1����J[�T���!��t�HR��SFE�� x�-�.|���sM�`.��� O�&*��+��H�ʞ+(Vp��0�s,O�҅?z�]Y�L��v�/L��O����="iZ����
o
��Ǌ>��%��*�C��yD�(���}^�soy���:F?̃.��d�nke^QS���E��\G
~8>���h0'(c�� ��# 쌄�|+hӞo�j�E�,�/��������2�+ܷ?�}]�_��DK��jKc%7\R��r��ٷuh�H�͙,��Y�̑����������x����@_���;<^���-�"~�[��#3g��b����p��3xZt�$��fX�(�Ȝ��C�y~�k�h�2Ci_}��^	��O��v{-��CY���P'`�{�ۇ�B��?���ہ5�(D��\o�O�6Eޗ����Z�ں��\�\�37n鷾h��oJ�Pu��%�tx`&�_V��IP������`�e�a�m_x�;�'���r� ������)��U͝��5�2`��ɤ�o���Bй�Fj*CO���d�Df�'%�Metۦ-ws�醮S��l2�B�1K�7�����atSjޝV�)�Љ������, Z�qn��:�{�0��JOWG��v/��@�M�P��й(���?_f�+�K���Ӌ9"�a�����u+�m�����S�o�����  (�wѭ��A�M�"�ZƬ�ܞX:�����
5��W� ���A<�h��Jl#-��V����x���3��-i����@����V�	���ο��[=4�U�5��eޟ[#��3��D�_x�q� ����ћ��L���0}�)� ��eny�~x�S�#\y�U���	�B(_��Z��#��7
�I�r��|aej�l����5��#���,kI7��.L.Q���fx��߉=���oqqʬTP������v�b���%+3�_P���ڃc78���{��.�W��kz�]��p
 ڝc������fJ�|�-.�K0��q���($Z�-54T��J�B���fy$M�(z	ӵo�2��85����J��_�Uy����Hs)��]Ȕ���|�m�� } H�����n���ޕ��	�*�7�	lD���>�2��ݧ���bdUF�w�b�g$D����\VAş@N�=p��E�ts+�]=�d�HK}
g�*�9��V[D�qOP.�"���W)�BeH�����+��$a���hV4kH����nm��({�_���LQm��/Z!����z��>�YbM=o��}x��fT���c��r��[=m}�7�k��b�E��J�����{�a�ήB�4|�	VIO������^���7kÔڼ�T���-�~t�'�#�V����������KK�4c����|��L�r��26��U񓧰�Ov�<�)�`pP��)��ݾQ���!�1�dƦ^�%�S#+�*��r��g[�?��nc���A���E��<|��Y(p(����ג���;S����Y���X9p}�B-��H9S�/�]:��f�.��~�f�k�܋�sB�]~g������1���[�E����ݼ���_� ���|�n�\������LL[�n�����z��<���(v#K��(��X��z&�o�Ο�A���Y�﫹Q��]Q1fi�U��j���l��o��<8T��ϼ���US���ђ�&+����+�fS��K�5�Ū����J~�}�Ʀ���dz�a�C�� T���jAY �Y�G��P6v[a�"n�r�QɊ{��G������9~�n��mX�z�E3�f����o6�UO���-����J���Jh�=u��*�Ս�y��-SdS(c�����bB��f����h5�����Ѱ�N����D��~��%�
<�Q�E�F\*��E�Z	*�=�g��t���&���=�$�v��[��Ӑ��?�U���>xnI/���_W0V��QB4�l�by�L��Β�k���W�.�2-��V�v h�����*~N��b��:�2g� !��/�z��r��h���&�Κ�y��;<Q�'~\�����,<�K�^�������d8i�aO1e<��[�����JV$J6枻��Rj�F���э���*�������q�F�me�q��\B��� ��<������XP?���}w����Ѻ/?]\>B��$�~_����*x�q�x��+p;�O�|��M���W�AP>e����UQ]Ye��R�=�����
��-�M:ՙ�8)sc�;�csW� h~ؼ����|�h�
K��zo,�%�-�)%��tz�E	߯ϙx�Q�[@<WL���<2����A���Vu�ٛj�
� ��Z�vŐ+P�P'�\��ReH	]�[锒a;d|`S��k�]�W8
��}���l�*��`�����M�(jU?x"��wo��N{���Bo��>F[��g� ͔�\>�^M��)�TC;53c�%'G����N��p�Ŭ4�/�x�CG VX���7�Gɠ��G
4���N�B��C���Y���I�nnƜ�q�a[�;�WH	_Lm��m����s�\:��yy7x�N2���+u��婞`_��.�_��S�Z�'�5*�C���%<.Ӗm��F�&i��[M����n�p��ar�%~�l���x��s���*?Q{��
��:z)�Z��"0q��=���I�b_he�zz\UN�J�ux�������V� Iq�;���
�N.&���W�ٜ��X��|�N�v��(0�_��yX����D���Ã�	2T�[��P�(Hq��$d��$���'nxZ4�B�I�������6�sݥ`�ϢPBnq�^(��|%�}X� ����e�aB'����^�u�F�Eb���@A���&JP��n����
�H�JY7�Gc=���V5ȏ�@�^�p�W��,Xoi=~:,%ſ�h�J\+A,���s�����R�������l�5RɁ~?��t�����|	�/V��Z��]�U�1��?Q�/vM�fN�����-�&ڮ��k�K�-��	è��]���E�f/	�4@�mzʸ%�|�]͋�v�?7�V4'�^�p�m�n�
�kٰ��눯�W4%�G�R܊�{��T�f�~�ՂT�G�>n_hOE^�W��K@�&b_Q|��uO��ˤ�e��s�5Z�d����lj�̃����F9c�Ȫ�/�a4bd>���\Q\�����F����n�!�&!�\�$RZ�Į�LU��G�]$�ŵa��yM96=N;R���Y����4�t�8��$��n�����K%�����/�)g�����	\&��fͬ�.�_�Ý�ħ'���*���X�;�X��*St�BKo�/��ǃ�-�~8�nU��
��/���w,���v(߳Fc�
���T���"��r�^KΨ�ǂ��9��4]y���;(W�-���`(�RH7�w��9�r>����'�M���+%Д��Ύ9ҁ���1�o�I�uX(�y�}�z�-��]5��I�}�~T<�Y~X7{k7�T����<���)��M��@��gc�4\�D�t..2z �0�j�]�U�<,|!����K��}���g3E=���J�F��b��0%�+��i=��l�$�o75J���S�D��%᲼�m��c�֔�@��+9�-���%emG_|�|&�k��ʉ�w�"�W7ė=��tcQ��8[�$W%YY�"���p����r��>p��rGj�^�J���V$��`ST+�F�Չ�!d�+�6bq�oI�2����r�|�5Ka3^�Q��>��D���m�CH�(ݚ�-��`��UU��q���5L�� Ҫ�
2�4�w/��6;ն��!F��/A?�&��D@k-�{[nWO��ފuiپ���h�C���]��_�5S�[^.�#�r_�Vr�,K9E����_٧n�ʜ��)�l	\���	L@o�՛m���4�)�o�ﳱ��ǝS*h�rj�Es�t}�ŕ<$�EnRN�p�M\	��j�*��\���`́�ORjs�{���0L'T��Íz�J>��b�?]��=��A��Vn� i���U�ɏݜ�K�I�v�����j��?ᣅi�Z������'��(7��W�Bk��Z0������)���W��N5�>�U����AҦ�`���������7Xι��>+r��z�%!�-l�&w*�PB��K�H;�[�x���r�����@lHj����GV���������V��R_.!)�-Z�{1o�~`�䫰�č6�K9�-�~��Œ5n������U�6*+'L5)���ӍY�r'GeS��,�|d���!i�Vx�ˡ�� ��T�a���h�;ȹ��=Z�_�v,�#Tqe\�������C��r��y<���o�K���Ċ�����=:'|���B��@�$�"S[����&͛�ȡd6k[�uG���q����z�]7�5��6�D�ُ{���cÖ�ǭ�ډ�µ����1���Q}ݿT�r�����C6��rʣ�0Z�S�W)ߓ��k����_9��>����&��o3w��/���v��*�nXd�D'�s��M�//�<B_�����ᮘ���"���:���ɢ*��V"j�4����T������{���%W�aۙ+`�W�%�7�,�l߫Ć{s�_�}0�է@å0�=p窓�_jG�}$��C��h��!]�e��73�h����+(��^?�D/� �,��ˍ�����~�4�|k�h%�A4Ϝ&�^)�]*t@�/�;w��y�9�w�=H�����bd���j�����]���o���WQY�������$��Gga�Ƴ��mj��'��	�a�4(���J����l���Q��x��3M^
Ĥ�<zJL�� Vn�/g��j~<IU]�g�0��$`ȓ�9sM~�Ȩ��*�E+I�f�{Xp��^e:"n�F��u�!�̫�#������p����>�_�D*���ܷ�|��nL?�6���M�V��xG�>p�/��So8�o�X0J=\SP�ߵԿ�e�s*R������ٴ>-�!�r��NiP	CX�Q�xnZ��#��� �5wb�*U��_	��(�+U�遝2\i�i*Fu3A��t ����w�\sK�v�Y��3�I[4�ʶ�9�{���E�nYc߇�[�MD����t�Cs�7��!1������3y�W��$G��F>_/������5A��|���y�zo�7�c�I��sUN��R�Z �]���`ET/�,
�R̫�~�¯��ػ��]O�)��JM|��,�cH�P,N/Pb:>}� ϳ�oI$.�C���<U.y�U������/k���@W�"s�*�Kl8o
Q�"j�<
y�'d�w^24�B���^1A�qG^3*_ȍ�Q��u���4Y�8�w�&K{]�J\�'"T`�SF�*ٝ��ך�/T`�v\�̮�o�pi�����j�������
��qE[%�#�q�}������1F�P2����BzM ��fz�����R��v����ϗO#�';%0rdW!ak��X,�N=|�Y��̴�����e��� �u��4 �V��O$����(e�&�
O3�W_i}:��	Rj�U�3$�n���/�Ɔ��֧��W	��f��J<���xԏ �v��zKZK���w�?x(��)/R�V�-�	h����sѯ�sb5�W��5ۤ�
�_�6mg�-J��V�Gm��O�/��|� ��C��M�Q�������6�W��8-�D9ʘ8�:��꽾1����M_��V�!�Җ#�@~���p9-�Ż̤]G�m���~>J�816Bu���
����<Z��!��3�&"m��yI 6�wC�����-;y�W177��h�C���TXʮ�.�9AdfL��<���I���=|7OÌ��Ҽ?�rG�Ҿ�c�B�o]S�����0�m���f�~8���`J1�> l�]6��ږ|d�Ќ_	w܈��r���ܴ�jS'm��(̹KC	V�����6�?i�/�D���P]6�'"W�A��[�퐌A��?QkJ������P��T൷T�"��-��h�W�⇈�:�qch�g�H,m�UQ�21��_y�d���h?(�w��M�g��v�G��Bn������
�ܱdQ	@�}��,�9�ۦs."T�c�o�%�3;����>�3c�Dತ)a�ʙ0 �*1T��f�J�Gŗm`�LK�9D�5�׳�o-j-����*uU�E�����>��ò���-b�FC|�M�Q��Ą�D�>8Keq��~u#�`�[�����ăjȃ��YN��Re&W^����Թ����"]�H�_�ί���f�g�8{:x���uz���Ex�yf�P����H��Hx ���&��^���i��z^�g��&ܼ�Ap�}�U�/�+%R�^I��T�H��H�'Y�T�Qx~࣒���;��eؚ>��#���P���4o��Ԛ�s���?�?܈2���\�ߛ�KV�1����� �9W�骗@�	r�����z����j�[�Ԁ���H'_�������ks� +�]gw��Q�Rl�g���4�RzCh	�PӈV��J�Cn%�?�UR�)����4B��6[B7+qêx̄l5��Ce�x+�a�����6�t��tN��x�C^M�;\P��B6Z�ίV��Qq_�h?<>�|�� ��=��%�}{� ��ġ����d���� K͈_�Ӯ��y�u�t�+�5ȿ�]r��N�i�[^���<8
X��\B��5�mNGjV���yR�W8��+t5N�̛,:"��Ei�*Ku}���bʌ�>^i��O/��9U�/J�`i�%B9׵���MjV��^��ǎE���ypWL^�3=�F�_���[v�O�@�NQ�՚��h|N�k�;��c�U�agG�v �L���ĝÅ�������k���-�2\D����-j.[�|Pޟ���u�XAI>��ß��k�@�</����/����+�{�E�����#22Za�O(�Z�p�^J�CɈ�J݀��N�1Ϫ'h��A�Y��H����/ˤ�}4�yC(�- u,7��A��xE�V��X��s�sm-�?�ZW�oU�-W#t�	E=TXb*u�Mj�!o[���moO��'��J���ş@�����.&S�	��(��'�ZyՉ�t��Ο��j]e_�1��[���G�����a���� o�3�����qe�d-^��[B��qLT˛y@�0>dG_����r�*��wz��!\��u����V2q�әXi֎�r��ιQ��;�2B�y��N�\p����)[:f:�=~	��k�9�@�ώ�>�s���}����[(�����.~����ǜ������p~�� �l����Ͽ�\Q���1����WӖD����?��SH�&���/T^ٶ���a�+"cq*��?��;���tf�90�HaSd	���m�p9#t��ǹhc�����ş���WF���YA>���U� }���K��)��eIL��	�\��gn�����l�gh,G�l�u3D��aU�3R�!G�;n�������7��T�'@�?r��5�a��ֆ'.�5?�ٛ��TC�ݞ��2{�+O�R����v�,��)�Ѐ.���W�7Ol_ɣH��"���F�$͑�'_A�U":?܈���l�Q���,#<�?������13�*g�k>�J�)zu�K�A��S�Ö�r���w'�V{�S%6���>�~�U;P!JҨ�R5oOYV��h�6�66���b,�,��B�髿XЈ�.>>D�\�^p:2O�x�)���h���/͛,i&�	��zo�T�B��q��雒<Z�h�~;���s^��&D�NK�CP��ݴr��̡�u�OY���CT!��d�����:?a~�t`�xX�R�1k}x��_Qm�L�͊ud������ŧQ�va���W�����q���K��HA�
�˃�r��پ[�������k��Ǽs���G���d���C�}\���7w&�&X@�!�p�I��U�
^���~d�>���N2$�q���U���9�ܝN��$�m���~���}�6�A\�W�2��9��t��58ҍ�M�;xR�x�n��zY9!��-�|Ǹo��E��B��딎��d�A	��x�<���=�FŨ*����%���}0"p��]k�v:��Pn�L>��K���)�
2�'9m
|pÅ�n���x��%(���1W~��{I&x����r�"ԥΉ���K��~������jر"d>���,����>���'�j(��7��pc��Ӎ��
�wo\�/>j���%�\��8�"��λ]Ϻ����T�.V����m1�!���/��=����H������E���j^W��0T��52�4/;��q�g>�H��y,�vؖ���~CS�Uk�BX>�ݼ�Mt���k7H
�"��N����3�*��{da���]TJ)I��߯bI�i��پ����m���>p/�g�#-�/R���e���s���j�`�MI=��i)�=�|���MG�hX����m�3Jma�m:���ԆڐR�"����r�=Y���#�Wc��Յ��M���u�������nw�����&Ek�����?�ʎ�գ���%��5ɾ<�|N8q _&�~8˓_0�e���;��o~���c7��O>�����=���x�R�h���m�,Yq�9�h1O
��c�����Ų���G�r��ݑ !&T|��IF�e7=Y8n�n�
�˱$`#����z-[
��h��[�&9�j&f�O�v왔>UV�����,�-*���,�;�X�C���a�����M)�8r�N�*��U}�&��_��Tj��l�vT>�L�_(��/��m�]$x�	o�aw�����i�a��/��j�)殍9Q3�~��T��%N��<�6�уg�.����� :J�\�?��S�ե��d��X;�����ѝ¼d_L�8-u\�?�KuL`#1���oE`#���6�e�PJׅ�����*xaUA{�|�V�z�<Q}��p��Ō�\"��G�Z?[��QK�A��K�箏���wS=��3t]�m�SJ�Ý���F�0w�8�>9>�V)#,��/&��B��
ۚ"�A^��@mҴz�G�ۿ��ֶ��j0%�{ֺ�x�T�	��N�YL{YW�&�ۖ��h)O҆u�4�E�w�H���C�X����=�-(�İHe�m>�u�b���B�*�5�<,"�1u��I-�;\���鐫"�}��f'�&��-�j��~���g��NY�����_V����T�A�L����������ᇳn��~f���A��H�d��֫/�!y*�́�����ve�h������08W�mp�}L���k^x�B���&�����M?�X�FË���$�@:4L��=��M�w��8����Z� ����yV�~#g��>qZ��ĳ4QD%����8�Dӭj?��a�W�ZJ;bc�e�~��̇�=���_����O�D��hi����a���ϯ�p#��ĵ����s[��s]�E�bړ6XA�<��7��Q;��f���
.)���d�l��r\�5�u�f�ʎ�T�^�qE�CڛoCä��C�7K�9�^S���T��g:����,|$�1.�x�i����,�+��s���}��z(w�U��W�--VQ��cŗ��Vca�IiĦf_{� ������1qyUe���R�B��R�N��E�^���~��ʁV�k�ѣ�c���I]9���<�^^o#����Q����QhT�>��8d՟y;3c�W�X�A�d��%�}����-�ֵ�|w��O�+��f�)$�~"�M�J���D��sݴRX�K�k��W����w���S������ڨg�;})�J�Ңt�0�����vYve_��-!��Go��.�2��x]�|�_�voȄr�n�u��6��1p
�ڵ�9DS�m4K�ޟp7<�Kn�&���
�d-[��7�O}چ�o��\!����/W���ޮ���{�����V��߹o|��jN\ݲ�_,�M�`
�3O�x-.<RP�j���a��fxu%0�BM��A��}CE-�T�38�+2�
?uļ+��x����-�+��:d��f����|-���\��~ߥ�˃���?<���i���N��[�~X@=�H��߹�͚SS�,�7����U���[]P�)��� ye���e�5N��fd x�1'�%���p��$7�>�t�����������>�����K�舳!�E�">��o˾�>�!!ݝ�Ժ�ӿ{���v�yQ���OFHa�aڿ�#�6�����]v.ꅼ�¿pba)��+�L��I]k�����*P]zl�!��։o��>����FO.N��s���������d�����=�2s��U~�XƊ&O$�?V1`���W���IR��s�$-�/9ܧP���E�!�}��ۤҥ�22�EE�~K�14A�n82<�"B�[u���05p�V꽦���L�g��Z=0�t9���h�US3�`�L�� �a`x�a��^�^���,���ڄWL��]���C��D翕6Ӏ�U֏�QC�o�x����i@)}�H�yf��l";6��Kj��Bֽjc�5!��ԇ���)p�͇z��%Ծ�V�h���;|>!pw�,(�q;G�@Y���(��+��5&Z�����;�뿴�.�4�������s~_���3l���� d`��{þ|�;�w���y8���=�e�+�/�`ɗ~V��d��|N��h��lN8�N���7 ���_�}ؽ�I�Rb��i�_Q�aP��핽u�9�j�=k���b�a*#�[�ł������XyJ��JM+���$�$S���]Q����O�\�.8P���.&3�=B�;�^�$�����]�J�	�|C�,�5�(V��kZ;5��;cm�(��h�{r8)�ҝm)�XV�_��T����b'�^.�(��Nǜ󗰾=e���������`j�֑hDH,�T�*�:�}��Nuo�U�и*�aF燋���j_n[�8X5^镻�
�@^Q��Y���)gU��،���ρ�X�#Ex��J%�
��c��޼r$12�6�����00���8��M~��=]��I�"��ڲr8-U����1�S	�+]�f�m+�Cs���Ř��B凥��2��Y�PR(�V;'��v��f?\�T>��E��7�K5@u!��_&�_�U���Г%�*0��j����թ���h��Ր�-�ê>��=&p�_�x��~���̡��)ɥ$��J����-�J��g)N}�"�Y���)'s��Z�0T6��!�E+�Aj/���ؖ@��S����D����co�}��}�+��Wk���?.(�)7Zd��G3�>j��,��;����a���(���*XU{��O���W�{�X}����F���*~M(�)�U�`���BD k���/�+9,E����Y�YŠ��*���wI�7e�F$����d�i���G���ZQtp��n����w`US���r�9[I���&�Z�=���e� ��B;���جe�:m��*��B�m�z���7��}���L�G�hہ"����n��޺*H�`�MPb�WR�%é�s��"�k�x�m�r� ɠ07� TJ����<��(���5U� ����k�W�����?ӱu&��)L��g�od���Gq ����|=�|զg�LZ�Ъ ��bw������5��.�/M&WN��:��!��&\���O�tR�p¥(�W�֮�R��h>���=>Y�d�J�\g �m�l�͛�q���E���g׳���۵�	
K���n�l��u���:�[�r���JI8�c���� m�Խ��,�D
1�2*q��{��s�������,Z�%�]7XdJ](�є١T��K��׫���<&'��՘����Zrb]4i��yMN/�� �F�m���D��3w͛:�Tm��Ź!����056�y�{˵.��Z�'����v�u�:�?_:����p��ڜ�@�ºv
i������n�_5�w�SUN"G]�켉�Ԍ�3d��hO�U`A[!��w�esq�Nys���Pi4�����D����
l�"X�SL��"�\��0Z�yj�F�4x�uݛ��v2���a�w�&QkKei|�Gߴ��Ӵc�@���F�+�ͷ'zxA�z������I�m��n1��R����ϥ���XQ���_��L�\y�g�O���+��:��M�VUg#�彰�a�X՗n�Si|��DK��������*��S�@�Vb���-��(r8 O�P�F��k�K�/_b�k�o��i*�D%+�����b���m���p�H�aLEz���պ���>�p�'���/4!@?��Fܥ���m2���&����c]�*��ܟW�R�- ��X���F܊VL1jJ��)��=�ԹOL9���k`��D=���3� �!9��D�*�r����R-"����G�
LR'�7�W�'[y⥾FU����͟�����^�D�1?la�4�>Ū[O����C�y��#�2��[(�������	��C\�h����UCe���
��h����2b�w�G�S�Rjo�uŧَߙu��so�d�>�Y�g`&�W+ijj���A����J�
$C����/���!�c��B�a�����{1�g�=���B�O�%[����'�N����h5��~��7����*7���T� >�R��0�@��(F���G���=��g�[�8f]3m�c��2���4qca��{U˥;Uޑ�� ��{�^՝>t|xJ��g_�?�^���1��,��V�~Y�O�0���ʁߏ���� ��E��ࢅ�=yA]�e�># ��1�3G���.�g�����V��w�
�����h���F�/���|���%� �6���ѠW��̈ ���̟�4b-վ?#���(���~��L����Z�.�;����0	�#��B�+̱U�x���JT�����s�a��5�����h����x!�o�&�XʺU��B	�e�y8�>.謨�Q����� ��R7]W����z�t �h�'�79w����QbS�Ӈ9ȟ&v��vF����v�}e�@4��4��� �g[@�Y�B9W��PU�خϴ$�W;�?l���K�h��8#�(��hMZ�:�v�x����ی��k��l�~�3{3��/�U5��ۿ��`|�;�ꄌR��#�?�߄,���&�[�����ל,̀��;Á���#��cǢNx��9A)a�B����d�c��n	�[���k1Z���^4���0�26ZR����[����)>�/"љ�w'[��ݤ�AL�,�n&�IM]t��8%��&�JV�k��EmD|��UPJd��M<���\�H�paU�&~��ߺ�U$n�e��r�D�8��������\���7vKՌP���g�W̯ P1: ;,�D�,x:bLu��Մ	+V���b�ݶwh�?��#D����Q�L�fI��Ԇ�K|'������(��\T�saK��m����X��.3����?���@�O�uٷ��8���-��dc���Z�ʫnU�Ⰺ���]M��z�?Ľ=��푏��+�&�[/l�uI*��/5-6�Tl��AS�5�r���.�Wu��E�m�O�ވ��{!V�-<߯�˭Wu�pC��ʅ���͵vC�7mU�o����5��y�Ov� UG��c��p1|-D�c,����1���dy}�Zy_dJ�G]��2z�aP�|9_f�M_Ťo7��kS��:���'_	�_/�3fg���U�eU��P`씳u��ӗ�[�WZ�����{�����q��~� ���� ��Я����y���e",�F�:����5���?O@��_PwJ���쐥'�1a̖�OD;�mv���se��f������_�DN��s������ \L/~H�X�i�}b��l<�)Aɮ���x�E��]ᔎ�3]EnJ�|��/�!�6-TSv��{�b�J)�.R����)�o���޺���.�mY��o���t�ǋ^Cж��E����qGZ��	�.Q�E���T�DX3'���%K]m�o�iIr���������_b��G�����´|�?��y�?00�-?�w�	�5��\\ε�X�����Z���4�%�<���aT��ٓ.�^Y����`M����{4G�l��l9����$��5���J��������.��D\>s�,3��pR���,d�k՘|~���2ؕ��/\�����D��+�w���Q�'����de�6!���������.� B[�>MV)����uP�r��2u/��/yuH2�}uR����$s{����kq�E�Oy��zU��7��r���Ta��ळx1f�n���ͲWp85<l�`�3\th�11ܦK��@��G�M��J�0�Bs���d)y���/O�_%7�ߵhY���BW����?��e����AXz�uepM�G����%�P�T���z�uc�>���=���c$p�_���#��ڤv���4���F���V��%}�������?���'�.ڨa���g� qy 3w��œ]��h��e^#T�Y��7JP�0��'�UZ�+���E��ҏ�>j��tF���Y��<8��X˛(��Rk�����Y��۫�S��>WR�������o���[��黚ux﯌�/`��ٗ�5!]����R,!�K��Z���k���s�B���u�aS��d�V�ɀG�(��0Q�h�J��f���O�ԑ�}�'��S�m�8����>�k�ePq{��,~�Zsvnb���)�*�wm��>.J�}��!�����Y������B]*�Ѹ:y3͉^�B�I�]�g����9/���9�x|F�7� �̮+�^�����< �`nѠYLŋ��~J�5n4Y�����K�|,"|M���/�|3U�ϊ%/e�_����x��_�.`���Q�3T���sw�޺˨�_��4^c�rv
�T�M��h����������A�m;M�8k�EЪڭv
�},�yw*�\#\����	?+�Jzُ�&�4J�BWa�<k��e�=v��ҟ#��G"�9�?�l�*�P��0��	�~Iedf�4`��������U|��\k��q?� 7�&c��7�=V���~H��"}�Ɋ���|)���)^ ����9��Hg$M��0y�_�sM-�?��<T��9�)��*%US����ݚ�/��@-�Z�B��ozD\��"��j��Oy���!+!s����u 7ֺ�qq8_`Q��,BZ��Z���v��m�!�S��˹4��K��<�zP��DԸ[-�!���A`d�_滕e�s�+�=�X,�d\���Ny?oZ8�N5������%{
:��Ut
��!�t�L�4��B۴�Wl���-����'F�8x(���%�W��A�g�`H�]���SW��w���7�cO*�tt�l%����� �J�_�kM���r0 �q�7z���x=����э�+���C�����HD�����������Q�3B���2w��:y�}h�x�����5��{���wei�,{��0��\5�-���������A��}�)tK�P'�C�~jG�H�|��e���Kv���/M��'���
HZ��`�;���꟠"�ֽ=�9x�<�����و�q�5~�@�>����I)�T=��hTFF�=0.���*��wj �9v��U_]��e�k9��2K�ƍ���S�X#:Z���0�*�`J^����BW�Z)�����R)c�p�#A5�1|�%�_X�>�����hwB��j���_,���S���t�`o�Ad{���z���_�p����R��g�~�̙��TM�X�*��s��)�?��pw�}u~��L�::�%{L�v��oW�t�LL�B�AI�a��W*Rcފ��(r�߻J�mCN��f�5�V���L�5�)�?��C��h�Yyq����ۤ�O��[�$,ʩ[�.i[���0q�Z�L>_:ܸ.�/k�|t���.GK�(
�]d^Y��h	���� �T��nN�t���r%�x$Hu��TPC�Ԅ�{Q�U��%)vV�dڋ���r�R.���6����u�������L��g��ğ��a�m��hW���C6�Y,q7K���f.�/��4�!�fn3'�l��޷g/��Y�$G��-҈<x���՚/̀��;+d�B/��/�|'����d�v%\�dc���>�!e�|�F6&A��h쫩�#�2xNI�0��~�,�h	��z2ħ��S�x�L�8�:(��WaJ�U%���J����j�u�Q�V/*�v�h��Eu5���3�m�Y7j�9�M:̯�x��oT:��˿\#�^���ʇ���ڇ,�Ub�GK���>+�U��������Ni���U
�W�֪]o���i��w��_�
ʏι9����b�N�L�� �?���G�.Y����/[��E��8����Kj|@)ފ����߭�O���q-���A,(b�����~�7E���)?P���]��}8���A4��:�Y�XxaՖ񨅷��*Wog�G�F��̕�����^�����[@<P�4[5�)��P�W����n]@U���Y*7��ѝ�����,���]QWU/��>�}����"{	��n Y�a��+�%{�/�P����)�J���az?�3����W�3C�h����(^�� G����ԡ��
��:m]�f򔔫�����2�>u�݌H$]O�e)��\vJ'D�4��~����Z!�J���M0ڨ��j�{ ��6(Լ���q�K˃�2��U��N7����I.����a�&$Z�
�����T�h	��o_��η\p���~~�oh!�������jwY-KZ�~��p�����.�-��k[	��Ah���w�W��+��R-x����Lq��ν�-����$ޒ�:c����.�fQ��݌I���5�Ѫu
�~��U!+S�LJ��.��%+���.�
�yg�bw��M�͘CToj�2'��ې��u�0��`�,
���`�ZZ�-�������I`���S6
c�<�7F��쓫�3}B�_����n�=�m�M���H�1O��t�-Z�)�0-�$a�T�����UI���ElR�����0b׾�C9�}$J�������4E���)�>��;O!��
K��T���������H�*�dX}Y3D�����Uy�2%C�:��fEѷ�+
�M��r�}ܙE�����.9�@���i����b#��?���{v����;����<V{
�3z:�d��T~��9��O�����@F�E�L�m���+Aǎ_L.}�ґyZM`�2��զ�v��=�_���
_/�ե�A�J�7
�"Z�w
z%Z$0��|u�rbtg��o�aM91^�7�?�E
��Z�<�p��������7��Ci�R��kMo蚛ٿ�/9�g�~ק�A��0��I��حKS�Nؙ8����WЁ�_�V7!48�S`ν̍t����z��ꀿ�Ы�Y_q�O�-��B��g�Y��p��<���_����>����p�O�Q�B�w)p��N���c�S�������n�gU�E試��qU*�W�|�x�ڍ���y�J�.9�+��6��	�`�s�������W�e�*����iw*�}�65�a����THԬ��Fg'�}:�3�Y©���-��+�G�Hdu|�F�Ul�4�7��3A�I*�`�Xȿ��N���-�n��u��&��Eܼu���|��Ǌ�-�6P샊�.ݟ���P86���g�Oj���k�����tP���͍��o�q���{w�.2LQ���(���K��l�������_}W!�W6q3dJ����~�1EphI��p(B-PG��^I/VG�zli��������8����EM���GJ��U���ڶ���<	Ж=C%^@��iK4V���q%J��0t電F.呵D�����m���vng�9Zn�<̔K]V�w����z&L����m���8�����&`A�c�	���q���"�X>�?�qHIz%-ڕ/�N���9O���JҞ�Fh�܉�AP�M����(�ڥc�>�wt��/��3����n���9�5�Dx��%&�X<��`��h�K~�qY��!Ź�������,�X�s}>@��Ɖv��mI�>�6�m�ǾW�0O��n	��~Ng��V�i��k����ݥ���ZKp��[}XQ������
o0$s�m}�I���U�6&L��wێ��)����x�(Q4���?��7=�㇄��ڥd����](����Q��fs�����c����b�����?���ŭ}4Bq�\ӯU��>
�
@&A��854j<&.��_��-Z�|����)PN�A�����t'Z��O�f١P
w|���0�ղ����s�Ü�{���镵UƜ��ؠ`��)>�U{��*�dM��K�}�_�%��'��(C�Ҭi'%r\��\�V�P����SJ�䑢�]�/1)���h�σ�I����b�w�ߑ��S�{6RJ�9V��R9�!�N;ۆ�4n����)�Ե#H�P��W��n�����~O[~���K|���x�=����N��ͨ5C��ro����5}���_����<¥T뮙Z�H��<-��r�8�i������lH�ͷ�7a"�w�.q	s�}�~��طE@_tn���*^z�M�Xo��35��\��÷��z%�Tj�+@
��
i:�57��oO��Y��&ځ���$��PFs��4W�����%�F��&ξ)�%ꎩJ:/�H�[ĩ����	�J���Q_e�?�5���p_�1\|h�v|��HY���7��J�ϣV%5��u����sAy	�@5�K��p��v&����U�oN�/�#_�Sw���~��qU��d�-ž��������e���a������R�*���'�x�֔.������[@>�Ş�X��ţi�֕�����ōV K��݌vܔ��E��O�n�CD^~�E�>+;PF���հ�;K������_�	�R��$F�����W4&u]�>�)�Pzi?'p}����.P�yK�Z9p�����bI*� �D�.z"���Ӫ�ƿa5�V��AŹY�%hTr�wm��~��)~�w�W2�5Ԓ�d���r50 �g��2{����������/Z���c4�ix�Vqd+�7��_�&�ɦ��A�a����,e�w����ܫs[c�V[�s��o=1�V�2��I�8W���,��zr=hdTY&���Ջ Tb0Y��N雎4웃�AFI�D�C";�r%��Ƀ��'�S�qI��I�K��U�!�^��h
P��`�%�C�mC|(	ۿ:���;P��hV��V��������C��2x��4��=��+���0����^��F{>�m�UH��:��;�����@��:��*۩�3�25;�+cF�*�ڰ�X����G����AG��Ŧ��������Gn1Ǟ?�(�|
�B�wWWJ�������?Axw`*��f����ݗ'�*,å���[^�_Ǌ����m��VC*ZdN+��#Z��3(�$T
�l>g
U!��aˑ�9�~h�u}p�'�|�	j*�z�?N["�_�]��{�6/����ͻ@Y]���F�Q.e/�~N��{�e��Â�Ru�x;h��UY��;h��%�>�޿$�j���˪��C�¿7�����T�ۻw��x﶐u�����mO�)?ZL�ˑ�ܛ��wXu�ҩS6F���_]4/[�S!x�:/4n'�攞���~��w�(Z��ƃb�ٽ[ͭ�C/6���v�e��W��
n8x��M���Sf��:�_��M���C�]�o��O�O�?�(�njW�~�+����B�"�ݡ3���a7௨Kޓ��Of~9��p���4{�i<z�}��l�y�fߛk�����w.Z�U�Fe��(���acӝ���*�e=H�,��_�CÇm��R�<R�%�d��Qb|�`d� .5�'�fp!��m�5�Uӑ��}�gEg>�=/(���5��_����:S_�+ʛv��
�/\�����?��.`�=E��)ьן.���gk�0�� 	*����F�%D�,k#/⽥É6
x��PO���b�~�%�����ϭ�ͻPڈSq)_am�&\�dD���!|:V����n���ߩL���=2�����ȵk�8�q��w�r�K�-�ހ������WЬ�<��v�n���Y��=�=�4@&�-��Q��K�Ö�c���~G�҄ظ;�>'�2q��e���0X�N+ ���.�t�|����H�c��k�"���P)�"rD��������a+�����ֹ����⇘���{��ݮ���\S��"������nD�F�@?�P9��<����]6D\��������Ų6�k������~[E��B���ӞzXcc�>���e�Hh�*Z>W��J�{FTW���Am΍B}��b���>�!	����Z��xw�dU�h�G_�D��v��b��>~�������7+3-��i��͎��G"Tc�y�[�ˁ��@IS~M�
�T�Htɺ�2�ϽF��֝~f��0��X�U��w5����v���@�_L����T��C�e�����Őά�~�`���_ӗ��/;��/.S3�+9�������+�R������#7A�;�<��M[�ǐ6�ȍ���S_ShӲu	K�P���e�~�rͫD�o�d�m���9�����
%�J|�8 t�2�;Z�%��U�C�8�F��e�/�*��t���2�����Sʈ���\���g�uxV��L$4"U�s\����S�*��R���~�V�
�8{�"��X$§t��8�m�4mj	�{n�O�uR�v7�q+�,�)�u�vr�1V��@)�gC������M�����W'D�j��\UNX�.�a���e�"���J�Z�.��ֱ5�y���h�l����An��vսHĖHD{�^q�&�*���T��݈�cy��Ѻ�����V�-JqL��#��o�����LC�꽘��C�aN�,Ev�/ԏvju�)[z� �_)���y����x��'o���Arct:�I3���*���W�X��3fs"��/� ���CM�����FY�eP a^�(z��Q5/J��lD�j��}�I1&��:d�����*��L���]���M� ��~�����R�N࡮�^��m:��w�:�P��%1��]fCK�V'��8���va}x6y�����;ԅ�:�m�àtR8�v>��	�7�T"��+��Ɲ�����L�����N_4��P��ح]��Z��s���A,Ů��8��~��l���>tl���X�3g��DG'�������"e��l�vtW��>/�{�O���É'��n�Sv0����i��!���2j��daq��e`q�IJaĵ#g��:B�X��_5�8�2'TX�`��B[]C�v��Я����8��B�fqR �������u7L^�hLJ/¶��6�6��8l/�q���u�x�J��B�}�'Rf\B�Ů�����h����]/��CZ딎U/����|5Ψ�eto���'=���K�@jg�yo�z$��Ie�f�oŝ*�T]��{/9��~glU5mu���r��UQ�W�0�����*_�n�ɾ9ɛK��|��՚me��E�E�Tr�D8�(wyQ����~PQ�IY@]�ǃLpJ����p��w��ܻ*�T�hJ��Jb��x�Hu�Z��Њ��\���.u�I���-������֏2�\�+'���Wr]�S���u�LS(>��E��|Q�T�]<�h��w!����'���镚Y]�OQ�\���o[�0)B���(�ˮ�[k��êʅѮ�"l�]���rUBō���p��Nz��Q7"��yS�Q�3� ͒iu�	�!#�r��k�5b5sN��ح߬��C��j����~TB���@�`#*?w��ү��+�[��XW��)��|�(!=�1}P��hw�Å��|���U���;6�q�.��e�[�R�d8���^������VL,Q��x�z���]]��R�Z�П�\:�ΐ;���������\:��'u��Gߝ~qw�k��R�$�f#��z�a��O�R4�]�ѭ�k1W������F����_���_�h��<XQ�v��5!��ψ)r�A
ՙ�!������Q:	-FK-��xB�2��e�s���|c�9Y>�����&�W�]�%"ZU�ί��|��sDO]�b^Դæ���e��v�E�/����^
M%�	��PL:��
�Lp��f�~K��L�FRж�q��H_��(�n�z��!#��#�٘g���E�`��pG�V�˰F�@�;ɴ*�q_��\�9�&�ּ{Gk�-�;_�tL�9����;�xWq\Jy��d��ə���5�Ȓcd�����`���l���X�?��O�hSܰW�A�#���H�݆*"�'�IW]�h߽a�Wљ!M�䧶�����Hy�6ܰ8S��:�0�Su�7���U��u����  ~�h֭��u��r8�j�?��0��?ug�s��k���*F]�U��-��mם_o�b\7J��}"Y�̲hW}eA�jr�T���tPc�s�+���U�T�3;+?��1t�W0$.���j5�ʬ�.<DH���^�Xx�z�Z���{O(Cqβ��:=Q�|&��p�H|c����?���mJfA����1�ݠ\�W��$r�T�e�Q���u�V���<\�Y��^	�����o=�zx����I���#�Y�WѨ3���h|׭:g���ݚ�$����-qKD+ 4�bU�3�*N�/�m�<�}I�j"�f��h��r�PE��&���ש9�����)1�����<~�>�G_�ZO���^�(����B96��Kl��r��ޡa�����*A����Z��۴y���h������?�/b��'|%ŭu��*x�΂����բ�p}���U&!"F���޿^�����Y�Ioד�f��Ê�������$tVF �u�z=6��Jrŋ�(���J�Fݾ�
�!�C^K��D)N+����ג�+�,�T���c��Fϋ��,��?\�������(>E͕�/I{���Á6��?���G�)�;�Z�E��e�-l��W>~��BQ/�VW�
�Q�"�]{��n�NDiM�w����U�`b��4�U��b�H�x��O�"l�k��@���d�A��ki�^<r]]�<�o��/�e�~���EpD�uV�>���_�[w:���[ q]%ڙ':�z����ƥ�n"N�=@��N�2�J�B�����H3C�z�u_ް�s� �
����+����W,5���g�z������.���Xf�h~}����u�g���@����׷ӣׄ�	m���}~�r8��Z%N�U������v)�P��S�m��<Y��j"M��M�$���}_ˬ��;��h�ր�`�OMu�9���^����/J�X��bP=�!e�4}aS�oc���W��v�,�B1���pS��P~�JEV>�R�������/��Q��Z8��q�B2�.:qt��m11eT�bI��CC��f��_rsX_&�;6�[�H尹�b���"Ng�1��_��H�y�\�t)Y 7��տ~~������\5eo>ѹ���4�)��L��рHw%�RL�HX	�ݨ��8z��qC�M4ҿ����,�����{`���i�<�̎{BRl�p��9>�l`:�9*7��J��-�ֺz��s�o�橄	����c-�̿Q�;~��v2��V���{.�ϔ����]����d��G����M���b���������a{be��Z�!�*��H��o8o�_ɂ��犠��Ϗ��u�j}�0����?�NcW�vY��ߜ[��W6�#��'A@S��ӽ$z�ỽ{v��ng�~�5`3y԰���.��\�8��O�B.U�C����Ř��9���x�RRĥ��K�;|I`�w}�Д!�ܵ�|Elt˽4�f6N0)z�I�C4EV�Ս�!CԿ\��%@�+�%B^VU�յO����ڏ������s�i�a9��}�}�f}D�J��*�O�\o%���&�Ah��H��5�tߺ��Ls/����]�A�|	�4��#�|͟\��dUF�lWq;��%��Z�0D�RwD2>7�c+`GO/qD���tlG5�IN�N��@�����>�\̀�_m�����q��O4��C�H��[�f��,��ݥ��(��i��"w�/ۚY��cu��h���A�����i���&fߟ��duU�������Bu_�����rcW�n�/�M�C����ս�jfB����]Yv�aų]�7��k�W��I�/�U�1��f/���[
Z��gf��M�Q�tC�J�5���m���� �[����i�j��]ź�4�����!x��MȒ��r�d��E'�^��r���n	�f/� Y���:4T��˪}��H��z>�Ƀ_Uu�C5z�]��qG:,�mp:Y�Ӂ�'��fMI� �/�;r�*|�a�(�*�]��F��D�o�/<�`��(x$A��_���Ҥg�x��y6��E_}��PQ�Q��R\�RU}Ƽ��$k-Qp!+-����&��Wl�:1���}���bmS�w�	��ʭT΄�����ĂR(>3�@��d6����b`����x�_QY�������+�������.�C��7�O|��_pa����>C��>����<^�S���BEk����M�?�N���xX�y�Ͽ��WMQ��(~�r�#4Ք������}{(!��%qs���/�Cm�7���Swh/jf	�����������:8�,�r��Sg�yFA����Cރm:\ehzr����Ý���������rJ������=cߖEZ��C��b��F���t��;I7s�S��*&�=��^L�������VO)������r-FJ�-�gQr}��v?\�N���Ϗa3����:�9���2݅�>�0*a޹u����S�s⬀l���������9�Ѷ��ES_��HI��rR�L���
0���� K_8;���nt���t�Mk�gҐ���wu�zz$L�E�r��7ط��է�~��LW���'�-Q�h���k��s�ؚH]�|�B0�����w����>�6L�7��P/i|ϢI ��LD�9t�a@["�w�������@�LP]11�c\.~�(����~u�4}}�̪�����ָ`9u���z<q�������]��q'u���K-

�>��w������q�!�{�:�U�N�%n��Ē��w����q���-<A9k�D��d�:��b���>�v���#�2��z���(Y��5�!��ViH�v&(�'�^vo���0����П&m�Ɖ��h���H69�~4X)�����9�w��J�����@!�yTh��9�3i�H��T��6$ܮDWeRne�,�v
�����r�_�룅)ͤ��^�Ĥ���<�Ƶ�ʾՓ?��u���e�O�'����«���.�l�(ݖ���v`bw}t���S�x��1D$��;�Q5A0�`{d��`�Wg\gk)�%khԛ�������>�������ʰz���距���=c	�$�,<�M��KԴ��.6ڨ�[޾�!������	�ai�� ���}c*�}�3�%F��m�7T�rp�|T��e��5|����.S�"�O�������tU���R+(�WqI��R﹫1�d=p���S]ޟ�m?��A9�FJ���s�_!>�-5T���=[����K�]��R����mvh5�+W�%K�I�J������2���|�"��Y���pS]};�K?�\�vx]UQ����+1��Uخ*��3J`�8x����~a�AWH���?(W]�A,Y��6RW�H�E)�TӨJ�{����3 ��PT�k	�cu�@���]�e}��&�_T���}��<�4�1�t턚��:�t��3M���O�-��L=o�LG�/�������JH�ԴEȩ������������:+b����y��	ƔHsWZ/�{W4~��L��p@}�/�'2_&b��a������Nh����~����G�?��y��ɚ�>'�H�D�f�SFV����� x�+����V��h�\�P��WN�ш��r��r�ҭ-�>j��������H+��&�#vA_���Y�y�h.MT��n�L�by��
z.��l袽
qt[X�J.�����y4���g�vh��U��xN��7`�l�$��~�Ͷ����b}�f��̫��m��*�����&�_��t5�:�zQ��O+|�̋���]��=
oo��)C���8��:�R/E_��i�F��|�=��6AW(�o�?���U�A���l�H`	�}����j�\��P>�T��yWk�)|�*sڝ(	���#����J@���юuS�)y4�>ȑ�ˀ�+g��0��S���o �YxW�_�pK1���+8I�_������k�ڈ7���2� sY��cp�zYy���K��P�G�u��Ѿ�.w�����^.,P��R�6Q�	�2#���5: Uh�����ʰGZa�(t]xPqꯓ���� ���*N��b��.f�����Z����8+mƾ:y���$a����}��@��7�K6���;�x�c
�LD��Rs���@ʿ��O,� ��>=����;����_a-��En47�.g�)5�v.��K�j���Ϊ�$��"j3�@T�o�����_4�߭��?�pMg�<:#G��p��}�Ӣ�|��{��|	��������4x�k�*c�S�����՛��)�YܗUlq[%��:�D����s5��{~٦ڮB�K��Rj�u���0~�*"U_,�bo�#_.��F;B�����K�t�J�ᄮ�[Z�JU�:h�'�P�[�$�/ <4�)�OM麨�˸Bx�b!���D#�ݶn�6�X��X�T>,]���k��w���t�W�^L��߶�#�1a9J�5�8� �H��S���Q�ݝ�-`v���Xx|"PiV�LZ<��l��/'�彝���*{�/�7YJuUL���jlҶ�2�������ݖ�R�����6)Pम�1�MS�w��{���pE��{=��E�\�'I�x� #���H��˘��F�?0L������>�6��71�R�[W����h3̣(�ܬ"�
 Z1�}>�o���Ew���sS��w7�ч��z#��1�.�aU�����;.��	��&�>-��sfo�vG��F��xQ���
}����~�9���Eд���zP�A�*���L�sn�y�lJ>1�V�8@֥�ӊ_%~��ya1H��r�?篭XO�{������^�97J-	�S�+�BDuW��_Pe�F�%�U��_�/����(�>����c�w^[9Z���s-61T��4YUN�w>�#
�I����)q)�>	�����UQ�2m�e4o8G�M���Z�a�׾?���:�ޙO�	��u}�a!��`h!]���NHVk"�����[�M&�W�[�a	�W0�$)$(-�ϟ�,2A��A,f�x�D-߆e�HJ�l=��)�,������=�L�E�*���"���Ϙ����^�=0�T��w�|=clo��Z�h��JfR��	��9�0�Q�����[��S�(��?4�>�\�1<�p���
��K�P1×�8hp��2�ê�V+���H�O�����VWV��H��tg�vNջ� �_A�K_J�a��,�'S:��%�%����zT�\��N0�
m���=5�����Py��T��a�.|�6ˡ���g�"�ģ����S몴�t�_qݩ��N�V��B�2+�P�4��-�#t�*��C�a!�<6�pZ���7j��
���E�$6�șؤ����kv�������U��(��K� ��̪ ��j�������~���&.*�U�2�|"�4 !�`�����%��<մ�P�X	�6I�=���%���]OK�7S�
��C� _T�������������w�����=��34�XT}e�'�F�=�둟�|(�6+{=�h�:�^��_�y���~_7�>˩�Q���(G��m+ �w�*�w[ޝ��l	�5|1T�O�t��y�UhH�Am�W�����,mY����~�]�{KJ��_�H���K4��ҦV��������{����廢�i��ݲv�`�W�~g-|��s{t�>�)�/`�������Ҷ�P��u%���
U���q�}��WR��n��<����>%��N�~��˖ ��P"�?�b���W����(�����E?_�!Z�dku|׭˨W�g�-~x�Ә�ݺ�:�bK>��H%W{�{���$m͖�C�����T�]�>NR-S+��������R&k�x��Y�>Ԇ���Fy��<��-o*и��n���'gU�ͣέ�w�b�[�53�MO�r�ɩ���P�5�����<E��rp������j�#�oq���a�שqz?~vm�R>����e�6�����ȋ�'=g��U�SM���F��JƫC&,q�+����k�S�u�5Z����\-!��і��1Y�_^q���V�c�AW-������������G��>�ax�V)ū��H��I�
����j�]��`|�����yϐ[%ZjE�w�F
j�z�/+����/�K�j�Z9/�<�$��8�'Jv��+R�)���V��F�J��WT"3�L����.���^�]C��!r���,���O)��7� �+�#�a��C���jri�uMt)��ɮ�/ͬ�Pk?JZVz�QB��g�}������BL�{��y�-�2M5*⪴�K��|'�ٲFc��
M�����-���7��⟮3`z����)!l��Rh]��4]B��2�"b��T�y��un'��)����l0ݜ�����b?X�����;(���h���u@�9�V�Ws"�*eQ�m������C���8f�X�X_޳��ګ��[�[�%)���д`6e��ړ��i��"�P�h�l�X����U�(�`A��*��FS�����O���j/��h��1����Y�M�}
�[��	��ʽծG��27�Z���O���H��J�0�+�>���܃B�)��M���{�% l��. �[C`�B�A\~|2y�5��|�*�-�a�P�g�l����}l�]��z	G6?�ܯ�l�1Jh�jR~_�.��P!��%بz��[`�ߴ��#�N[kc"t�z!w�@l���T-'�N��4բoj���Kƕ3�lY)[x�A�ޖ��AѦ��$�
���]�PS��B���E����ӻS����y��K�Du�=�8ȗ���v?*�/Mo�ѓ���Ko(V���vh���h�V���Gf�����^_?�%�ҫ��=�3�4�®+�h+
�C���a��$�&��V�u�w�����L1����S�N]�FUJ���!%�7&}pPu2DIb��7^eM	x�5��"k-�;�-x�h�k�[���k�<b��TM�>u��@_�劫�|2�Gq�,�7خf�v�l�<�	RyWz����B/Y��>�_�l�+#n��^�)Ud�	���;{�{�s���&q�������w�`u�<ڨ��C�`c�x�����/K��{iy�E��ѫM~X�ޙ'����~_h&z~:�*TGLם%�O��C������_���>���h�R+"�
���j�!_/�Ͻ���;��}�G`5U�0t�?�*]K�Dw��L���kE�VUp�d��A�����ݢ�9�N��,��9f_�*�s�B���.�%C�\�i1��tK�W�*@�-��0BTl��S�,�V� �럈�q��I���-�����wv��R/jé��WV�7��i�?7R����œ+�)S��"`}T����̧�G�_i�$L�9k4�.j�&���\Q��D���K)u%;H���}��؜"&e�v��Qֲ987ed��5��u��X}���o��s�ۻR'����z���F����}��}ä$KD��e�1u��� lX%;jP��oI�#�@��<�X�g�H�L�o��f%o+a C*�@����ၑ�+L4Fձ�Ak"�%���(���2�"`���A;�bơ�_4=����|��v
ԸQ�Z��R�-q�x0E��S�F~��m�&Uj�k�2�B�����t����u�I��%?��hj����nÜ�u�dʯ��/�.Ϲ��V�𒷫"�T-�/�O�I�骣׼ �r?� O������>C��/;Yg�P�5��������db}�I���l�Yn�]W��B�\w=����m9�
�ۜ��{���|�/n�)G%~���G��^�Я.]}��~�x'������_�gn��a��+��y�dI:�؇��h_%�^�v���.xѷ�P7;n���<�f���q��ײ��>
-�B	+'�]�wO�U�?*�o9�]e��ž�y������ȉ7�5`ڈ�V	��j���߿���:�ӟ-V�\??"��#�9���K���\DUK��K��� ~��ɤ�;�z9�_P�����2`�%�Rr�w�X���,�>�:e�g��dm��7�4*�0�Sml�~�ǁa�Wb@m�����:}��W53�Z���I ��Y�z�
.^Ǣ'��������
�n=�y��|���q�"-de��B�{��D�X3-�Z��a�(�ػ�ly������3�]5�2c�E��9:[�b��F�C�5#`�X�����}a@�ڕ b���R-��ߴ����⋮�O�2p��!������V�a�\����p��hI����MU(��>�t�ޟ��q��dТ�(����b���n߹��p|���Ȇ�\ĕ��R?a��cX�Q�z�>���HP�*�?)=�VB��,)�epyp��	H��:�%i;�Q����-�_2~��C�5��Kn��c�Ak���z�h�2�4K�.k�S�g�Jx���!stS��������;����女��a���}�ɁؑVB-�w b�ư�׊�@�-�����h�k�HI_�HȜ�������{�a�~m��A�Fj���pA�n��P�Z$�#�uo��i\)�VF�����ҋ�\n����j��+��Q�(�����z����.l�ڀ'Di^3�8;�e|���3A��d��2%���~ђ_]f�}�����U �a"�V�N�[��@���>��.����:щ���U�" �����i�!PW�eT�3^�h����}��bE�E{�]~q��q�e����W�6_5^�U�WNg7���/��H��ٻ��v��^�s#�]�צ�sܿ�KD����ȲN�@�mw]J��ޤ*�b��g����ԅOy>��ҭZ
>�T�?d�����*nE�h�v^�-\y�;tq���ѷ�U��6�S���!F���� vt�@ϼ�J8�Y��	pi�"��0�IZ��!�����(�g���Sn_��]W��h��H}~��f��4�X�jo���6	�஌y�s���.�}����JfO�]�`�KwP�3 {`G��Ō�2>���W<x�)J�y���_�����򿌠�?��?��0�n_5��ll�k�h4�z]m��fM�֋_՟cw
�mh��S�⑎:kt!��լ%$�a���I���ĝu���R[{�.ٽ~�w�gՙ.�L=��K������|$<�~XY��KUAEm�Ȋ��[���w*8cg�T꠩�+�z�X �Ͱ��wd�X���{}�[_��g��>G�������X�Pe�e8OP]j՞9a�$i)�|�#%�����9�3�~g������} �;k�F��U��zjsc ��[�11EZős>)Zfqo�A���r��O�b�gn������ͪ���۽��e0C}ШL�� �킆˟U���z��y�#�;��+�p ~h�aU�׶R�H����V�)������*�ui<0�4o*���Ɖ�?�T|������"m�S���KlbE�U/�ފ��1�v����Ɏ��ȃUj��/Y[f�����6j���/9�"}=�@д&m~豣R�{75g���%��_R΃;�P�|�A��{RZ�k�J�\��lέ<���7E�
�bkA���5=��5��
i��Aܷ~Ĺ;�~j��۟�/�zm<�����^t��fV���o����(MKHT�@�����P��	�=b��I-N|iUz�2(OGo�r�^hkU�3�9am����5p~��:�(�Od�����]�UY�.`�'ݔ��u���;4�=�Λ�p�^�Q�~���v�Ѣ��'�S"��LQ����V��]�P�5��|�sMOK�;�$6�������E+Y-��w�h��o����~��Rк�ydM]��!��N���u�`���!FLj#=\��<��ӹ%k^�&ھ�*�폖�~E�f̕�6nY��ېJ�xY��wm����:v�H��}x �+U��NGV"��!̖=KK��>�=��}ASd^���8��F+���oJS	�-��[Y�X��[��#�Q��V�~+��<�کR{�]<��n!�bS�b=d�+�.�=��r*o
u��np�_��8a���P�<��B���E���*�oA�P��{0sv�S-�ڋ�P]{�B��IL��B6�E�ޗ}H9B]}�����3�eKq��xJ �3�8����F��H�D;}f�&�*�����#w�l�+�p�hG����N�	~H뵠D�{W��+�m�����Q���-���{n$-���:jn��3���L먃�c���Pm����^��7�|}�l��kOHFR5�:g��i��%]i�SR���vLF����e�q�[u�.�O�AEŤ�'}��o�X�6�����7���W��e==M#%��`���Z)T��D��Y���@�&��j�9��ROκS��~��3�����~n�D�����\p�q
'QfM�h>[��+u<U��{�o�������s��?��$t�=��q٤��٢�*�H�&8�#�u�m���O����"�M��R�j	���mC�I�?Ʌ��͓t���t��� 3Dcg�m�y.K`w[/��2\u�g\�X�}��?9��~A���c���>s��f��ʁ#�~F|�]7|���8�(<�@�/Q�k�,eӎ�ƃw<Z�V�b�_��@��!��3%aC�C�Q�\ހ1tP|��;_�S(�ӈ1�j6�M@��39����+����sj�h�k��EͰ���l�3Z� .�k���kjc[���~�T�A�K�u*���}�U����Z�H>�Y�Ź�@F�h�;a]�R�2�����\�sX9��J����<��uu�V���ը�δ9��"�ݠ������ ǽ���A��o	�n�s�|5?D_X�:`s���_x�����Q֬~��X��Ze�;b�Թ���Y�|�zT�����)5���Ҡi�p�O���J:ck1�-jF$�Y0�"��/S�f*���0��tN�Ľ2��7�\	��:�3���l"E��F��	%v��'[��쭯��/�?�`.Kt�.�%�5C\��ﮩx_J�ov��';��aTM��/��X���KU�k�@�K�j�B��8�����21x!��5?��&��t�2
�a�0}�z��ߤp�%���V�~�z%!x
�HV$Eů�˘�f�F\�*���5_�I�����*�q+�t\�Ӌ(U�e�#���HfN�x�}� ���Ϛ4Z)6ɻ�n]=��}��Hhyz�~�*�e�;i�<�-L)D���Ek��Q]Ϲ+]��K�Z\1���m��_��vl���T��ѵ�m�Ys�zy���j�8�M�N�3�u+�01ć���`�0����&TtK�Ƕ�p^6f@VzV�	2�
����m	���1Gb0���:�uj�J1��1eǗ%�d�Hw-�̹i���sƠ���,�@)$�K)B�'�\��/�^o���T��mh�Dq�R��EJ�f�^�fHc����8����i����0�|i�;�����c�;���`Kh���+J����$�0%T�6Z+��Ø�}[�;���=���_,[Y��5&Z���>����aT\crR�/BCu)V�o�DG/h׬RB@�Ĕ2��!����~e6���k��-�55�h	%��.�=��xm�U|�>�̹��s��4_�%y`���3� �̖�O;�\�u-�_g��/����E�,'4����_�����/���M%��0�NS��3��V\{=�}�Ӧ�7}���ء�
�Z����}��>�����*W^�#q�T1�N��Bk�d��D�qqK��i[�RC��x�q�}	)�ˢ=Xkܱ��Wx4��:��]�x׶�|w�hS׏~~آ9� ���%r���M�[?�ѝ\˕uO@�wA��u!���1r��H���+�h�@�j*��s�(�y3K��H�*�T*7�<�.�z|~v�b-���wfぬj2}w� ��I��w���Oe��6׈�YS�(����zs�g��Wk�!ܛ����ZDP��pF�( ��N�-4:z(7Mg�n�o>�c���b��6��ٳ�T��jD�L�m[�U*��;d9_,ǁ�m�3)t+���\��X*�u��ɓv/� ��$z�M	\���v)J��5s��p�!i�y@����^)v/��zۯ�=->:��`$Q�/R�&	[c�qw�:M��#�s�'	���_6L��h���
6~f|1��,��	��C�Mri��Eh4Ͻ������ہ�f���W�&�tU�����`���w��#�u��\^�E�XO��fv��?s�ld��~�z��������`�?��]}x����=�DMR��J�IM;������r���T���%��J%�Dŀ�"XN��u���n��e�@�Qo=R�x[G�D��O�`;aGG.f���r�pI���)d�f�3o�~b������@�h��[�3ř�c3q�ӛ�k7؝����LL<���^�Mi�pd�	!��6�/��2�h\e�ۅ
� ���k�������G3vK�:�*����N�?�hj"��\�K.\n��q�%��D�3����>��ף�����!����y^h��:Y:؉hi�"��WE}��I��@-�S�2qe���]���������YXMWn<�˗��t�0� ������!m��"	0���<�=M��{�P
��n�f��aʾ},�&��$����Y8\��dK�����}܅y�y'�a�EV�֐\������J$rw�מrB�.���5a�l;��]�E��u/�-w@Ti�g�?7�����jBW����%X:�%iA�/��r���V[�~�V�/%
��#L>{9h\ś������}��e��}yK�˩I�pa�La�����!�k}����ܛ���s�3��Ǽh��%�V�/��+�'#����;|w�,���y�]cd{F{�M�ϐJ,�_ڨ��ۛ*���h8܀rX*M�<��ڐfGUE���4<yI����OUqj��w�Ӓ�w���(���M��Ǒ�F������>B�7��za0Ra�?����v����ܵ�~�v_�����1ub��v�/�`�]�⫶���{�+	�����f�$9�٧_Bk~OK��w��Ю��Ws���3�q�Hy�DwYi7���S��P��㪣��y,^��2��@VX���wi_eK۳8d�l�5���w)t00,Ƶ��?�ɢ�?Ͻ\�&�F��>=]-��8P�O���5��Z��W���죿Q�\��D��|���#�}_�F��)P2����N�eTi���}�d�&�V9Y��@�VQ۸���-:��U��KY٣��L�L}E�1F����83y��k)��k�|�#����P�;\$0&t܎N�R9+���T���~����F[Y+��5�}Wfh�E��'�����0�*~t��E�_;��Y3�࿺���V&�-�ގ��b|*؅cӀ�����;�q��K�-{I�ot�����?DkH��W޺673�V�o�J?�b�F������l��<\�������þ�XA�u'�b�����jRp+���y�)��Ԟ�lW�;W3+״������J��4�-����z�3�B��tp��.<���][���=��.�����
�c4u5\������*�4�qq!ɽ�K�G���9�ѕ�y,S+ĐD���yUoq_dy[�.�r��Kf�뒎�U�r���Mv����m���[|~���fn�d�/X?�����<lU֊C�=�9�9.�d>�񔬮[�lb�O���Ew'�����̪i�_��Y���$[��� ����'6�W�b��HA\��qU{� �[���˂a��L3g��Z�S�sÙ�l;��jD�������Ts���*ѱ�-Èo���E7k*z)�H�F�P?rmzv>��]�e�A��UvI�o�.+�YB%"ȸ.�}��kf(�n�����4�T��$f�T��,��u�_b��D�u�m>F�o`�3|l��jyt��&��N�=e8}��q{��_��7���Ŷa`)ŨIԹ�X�~��o�]eΆɢ��\m���꓿���|�k�2�m��7M�̴S'Ov����S9]�Å��a��/��8�V��i=��
׵(�U]���K������YA��-��Hc-W���Ǖ�HlH�%C&]�c}/�2�d5�k.xG�,���m��x�����d����� ]X�hSO?fܦ^VZ;?Z{S��O�z�Y\x�g�`]�)Q[>2�r�:�8�e�3�Y�ѧ��x�H���a`T��]��}P�\cŕ��ǌ���]��b����^ʱY�ϡ�(�9Sm޽;�IIϪ@�s,����Y��f���&s��'��||�P������
�P��/���O��0)��a��W��9}ӌ�߱l������8�,T;�4���DdbݏIQ����_���FsG��<l��c$���{q�U#]���&k�?C�z�*:����y4��=fnѳ�h�mȩ�KQn���B����j(�?w���;�|���O͚U#<���OI��V�[��w��מ�v�����ܨ:�=%�2��)��e�UMW~�q!pV�s���:MW��i�hyaEX�k!w2ݚ�d��]C�?D];�ú�^�|B�[W!��Ś���L�i��e�]I��`@!�u
��O��δNꙁr5m����d[��mw!��P�J6�*o(����)��v��*y���u�Q|�����Ss���{���Q?��E�˗l�bbS��K�L���(e���������ct�j��U��LhQs��9��m%�l�b�ಀ��=���୞n�qW��
�W���.|�Ƨ��E�3(5OJ�K�f8��x�f�gF(����}Ǽg�oo
XӸbӖL��F�Au�KV@Gs�U����`�Q�ʨP����o���d�w��BkJa?���P�̌�=0ӝ��}��/�)��ij�N@��5J�q���omI��aBȮ����V�*����1ٌ*��肋�c�1����_�E��n������F�N�Q�l;`�*���/�v*���6|9�}�V�_-�+�m<P��Lx�),򞼁a�8	�^���3��`�h��?�����7Th��{���Oݏ��8eh�������:{�]�̇_�U�R�~�N��):��U~��{�J�S���Imv����Y��a���}z���\�Z<����g���Hr`�����~��ɍ_V��ߪ�U^5�U���V��s�S>h�2V�aq�ʕ2�g����_bEN��!�Z����*$�Q-����r����BW{���v|?p}��K	�7��a��3���z���8�^��sC��x��c
m�j��r�{UW�� 3ri4�%�	�kB�I-�y��EQ&��-Ǝ��
�����=4*>.�6�5U��&Șʯ�K�f��$x��9���:WO@�k1$�>M�f�8�6���	����>G#�W����ؔvޢ'���"�#���U�NH�S��
�3#?�b14+�U��2v�6>�иr����[T�=�lN�oAѴ�\��Z������sD>o���1���qa5�[�cd��x7\�P�,Zh̩
���Х��Ka�k�'��X���ug�ݾ��v88e4TjoL��>��Í ���#�Q��/�E�.N�Z��݊5Ҟ^�E�
�O��:�(��ms�u�E����;6߄�t;Uk�����t�Y)�^���FìZ�1"���g�/�)�:���œgJ�dg���կ{]�Pu�J���b=Z>b�6Q�su�z;~�~��&;�m�m5g_�/�B�QJ��j;��ͩ��+B��_���hv�6
k����fP��@>!��g���qHP�7�Y:M_�h:����8u���-���=J��;G�r;�
��ުN�.C�u�Yw�����-՝�dս^����S�;L�YPcs��J{J\C_���\����*�q�Լh��
��>����_����(�vg�%)�r��l����-��ݠ�z2FK�O�B��M+3��Z����.��y��~�q���ҋ�SfW��pѯ�����tg���[T�%��������<6�h&Nq��u��:w8J�](h{w�af�Jc.�?L�]gp��*�"\�����u���?����k̏��^����'ڸ^��)���� A�u� �o�䨵�ِ������֟����8M,L��J$W��?f��,98V�[�w����؃s\�ѱ��V��&rC��;M�(9eN�آ�f�9�B�1�������g�D�K�� �|6PU��GV/y��b�N�3�@�fqݬ��a��M������ßy�7#W����*f�ă�=Q��g���R��|au��%��X؞�E�4����z9��߉iS l�Z��&YHap�b�u�n���[�ة~~�&�&*>����q�4�v����)Bz_�c`h;9]F���aB�����$X��s�s�W&�C�S�$�pw���F��[�I�;�iDI��T~kV��9����J�XT�5��S��樥S�_&�Gʍ*�9Z��pխ�Y=Q�ΛU��ⲽ^�>��p�}	�m��JU0_F���u��zF0�1�$PY��+�+�`�1Ljiߟ�Xv�F���β�?ρeɧ�C�93J��I�Xb�����\&f��<�0 ���S�Sc�|w{!�G��!�1��Ӈ�C����4 e�x�B�8^xĥFU
?<�fdا��W�s��=�~�7'�i��yk:%��0x�6}��%ڕb���Hߥ/���'ԥ��+�Z�
�,��-�I��M5�M����U��f���:���%ɔxI=�~`��t�:��tZO%H{��Q���>Dx�qW����|O<���Z,&������R���@�U��fY5�����?9g6��
�M>vq7sl�%A��-��/���=%��)u�y�C�Z�ɀe����{�0�5���Ԏj`7�&QLS�O����!)���ˬ3;׉�V����e�h�X�U>������~)�?����b���"M>���m�RJ\ahtö7�������'�9�έ�.�2�p���WZ[/9*?��@���v-wJE(�����������̏}RS-҇�V��ɎJy+�����Z��فIOe�$ru�fOy���@N#�����I�mױ׊oE��~<0�q>���/�]�"k�̅�"��L��/A1����<9υ�v�]�!����"WԘ3��j�Gs��DxK�Q't�U��k���Ye&N=_�"]��_/"W���w'?�����g�� +?}݆�m�����EK��޿R�`kKq�k=���bt$�k"�0e���W�%���L��t��G��ر�@�"��p����\fW��ϝFD}�S��V��Ʈ�����|IU��6�H|0w�����&�#�~���T���YT��.�ힳ��O��fy��?�͌��"��E	��b������U��-QM��j��6�Go���u�t�ۭ���h9O*q8JW�ߖ���a��'A��E���;�4g�Xg��hmǻ"2���J�����q�.3;�6r�gӹ%�hN#�N�@��./J?\�O+�����]���Hh[_;��'ET�ǿp�+�}��=]� � ���J����V4�ɫ2> 0_�X��Ro��o�k�%N�R�.��3	�?�"{&��Lt�u�y=}g^�ɩG��]R�2���hp��"J[���N:A�5�ԢBd����V��a��	b�2�WSH]����y�s��<D�Ž�u�i5u�"�u�����sU���'a����2W(�5T�����Ɋu���;WO+�����q70|˖R��}��'�zU��[s# �CWy�,'��G:L����2�qNH��\�u�xȎ/L4+q����a!�����&�<�� ��5�uB��d+ �*j��9b�-���L��]���m�U�բ��7gEXQw0��z�l6�T�s������h���'�kyy����Ȱ���TS�Hvd�!©xjU��HY�J]Eﶗ�xWF��BD��n�k+�͘}��@�v-̹�Uv螅ߝ�O��{`�l��2��<8�"�P֣ߟ�\�$YV�>U:�*�'�Am_�M/� ��>M-n��UG��*M��cb���VP�$g��a*�cL�����v���a�Z�nY��K:�!Ö�,��Z�w�GG�a����;��
�&B}7��9���Ǒ3�����-�w��I��T1�'$į�O^x���~���_$��-7���P��1ٻ�E_L!�2MUz�ӧ
�=�/�6��t=[�L��������3D;�L�c!Y��F�u�*>���3V��0�-TΜ�.��J�%��ř��D7�JE�*�u�?u��3c��b�6�,Z�w$�6uS)�<�$J�`W�a׆U0=D��8��&�<��ϓ�
z�}Z�+�w��1�!v���W�-�ԑ׀~sg���6�O��+c�A�Ù|�B�]-�C��{�>����G��,�������"�<�_�{2��6�U���l��z]Hx��W;��F"�YJ�`tOԒS>�W(]�����J���}-�r���ߔ�h�R5Da����/�x�s��|�r�kv��b`U|�W���r�{������H��}(�:k�r0��ҮL�]�2(��:�,�wŝ�ک4*��c�R�kyǷ)5�������8�Z��N'_�"͓ґU�����:_�	!�
�2>H�ϰ?��~7+�mJmnںL|cBk����{�*��ܡ��@W���D�>�^GK�?�=�����(ΕC>u��*�_ϵ�i~�OF�W����y��uMC%h|�X�����"
l���(9���Ǐe����K�oap�{��4oj��D��+�Mx Ok8M+����tEbLm
C���1H�r.[(3,�g���U�"��3�-�/��u,q�ƺ��/�+۶���r7?�M���/o�L�����3!�������a��(L	�"B�U�n1�g��#�f[�%���}A.h�4�O��1U��y25S�:��}k��*�]H��K�h����+<PZ���:��������������h7�������)���.O�>��w�r^�\}��ݪ��t����p5�
ц�_y���~=к��� ���G��GQ1YJ�X�
G�5�'��qfb۬?��}�ɄNW�sކK��=Zt��±�_k���E�/wi���f�1�D����ZhUt
���}T���j�.�V���{�Niv�&���Yn���T�C�=�����2N�V��Z�~�Y����/�+�r�#Ü��Z�����L��)ҝ��������#A�;ة�ߦ���"��G�=�
f�r @�_�T��U6�z-��e�yu썆�����6�k�a�������������ҵ.Z�]�~8�J7�b�g�YLE�
J$c�����6�U:C[G8��Y��Z��7l��u�Y��� ��i��E���d�B���L^�.�����T��i`%�T�����C���Y�C|,,/sԄOP�I��b��=(�vp���ߑ�u�~�Oa��N���il�D$f������龯�\`���:_��K��	MU|l�a��s�Cv��_��P%x��"է`����dRyێ�M��5n<�7<O5�bD��@�-�L�����n6��Zq��������vԶ�,3�������Z)����I>��Ťٹ�CƗWH���ᬾ&o�=����	���=w< e�_E��Z�(M���+�*O ���his�=dz':��%�6[U�����N���C��q,�V�U	=����Z���:�Nt�Gޯjvy��v���(����e�o��c�k9�%���GXm��������M�sDK�V���.��%���Ҏy�?���ڒ[����+�����ґ��p/��)����ҙt���ma�����ȿT��\s.^��&�}u&X����kK�ܹ=�������d�+��Dp�&����%���
���:���q&��-���?��H+��<�j���Yh�ā�(,������K�A͈�~��h�mF���C��@P�N�4�!��n�Ȁ8.�H0_ݷy���Cĩ�'&���a3���O�2+���01�n��<�/uEQg~�o���Z�b��+�w`�cU�U��B��+�ތg�����w�$��a�d�.�Z��#�ts'��,��X%���y%�W�}g}�B[�Y��~[��g�v����11�;��/K��qR������=�{}E9K&�
ݟn~qڕ��'�^3n<�'Y���WĨ�"տ���`�3��T�\��73^�K��9n��|ɰ���Y	M�Lzr�w���A���p�,�p���Wmv��C���+�]���Ww��e3�`}9Z�J�����8�;���?�S�����?�{(�T���P����ʦh�f�s�5�zl����-�W}eI��v_�l~֛:]]i��d�M�ew'�ЇPPٵ�q.�E�	}�F���[�{���@	���a�������ަ�MW���;i�>3�_�J��C
Z��U���)��y�W�%�3G�K�;�Y�V�D�vw[�R|$�� ���:/�z$7/u��tF��G%.����=s�����e'�(��u=/KlzH̭>EMfe����^�~�}1%���I(|�0Zj坤1x��Y���,�#��r
דE����q������/��U~h��C
�&�.�҇�S��}<0ǺZ���O$�"�_ü��B����u����;�:E�x�e������$���}[�����<�CY;KV���]�l���K"��E�����݁@�xYhcH67F���d�L��Fd�A4�GWuZ1P�����Q���>2�q�>0B����I�P�$?ֻY�r��Q��mR��	���	Jv�&R�D��F�MFx�t1� �H��j�b ��2k&X�3�8�E�y��3sA�f�jE{5��[�d�d�ݖ{�C��3G�5��x���5��CWYﶉ>�H"}����T��2R������7�w-B� ��tP�fC���̹�����v�4o,����3d���U��Y�H�_W��,[� �bH�s՚_�f��D��^�1*W�a�e�[�;��zV�]�n0�����W���x���H�Z�d�%0���8���{
��*�Zc4�Ɔ!��|��1�����;��G�5�	th�"�����;K�`�a�#�c� ﭵE^/�5�2��1.٢�8��5y�蜣j�JD��C����:��	Yb������S�W��|�`�����Xd<��e|�SIq6��K����~��vWrJ�l,J���=նl6�s��N��s�;`�l=��~�!zlƗ"�^��(��g����X�����Z���qrfZ��*�洺�����FO���(�`s��X�^�m��}���;�OY}`��W	:ϫ!UK��.v�x8���XZ�:�J.����	w�_��h�p��z5T2�B���h��@�A���W��&|v�7��]�>PS�Dzm��������-�j�t
E[���&SG����kQG2HJ�F�ƥҋ����wF��Y�7����"�XR#u�Y�@��%�{#��5��!��cW[w��#P�[��p���^����Z_����3�M��/m��p�����W�W'�<C@{��W�ldkF�L���?h޽CS�Gz|���Sq�b�*!��7/A�p~o��|~�3����چ�c�����FLCkl����Ԥ㰆)�W����}�;��_�O���;�����+�̶6>R$�:7�h�_)��W~�����H�;V�K��|��<3,�c{s��	ON�!���|:_��_�C�SГ�r�����b֣��v��+�ዽif!c��ʭl���r�N�zl���B���B���lo�|�ǍG��5���gD��q��]RҞH"� Z����ʑo��@��˫���Ƶ��d��v����)n����5Yԕ��m.g�}�����A�Ye�*g�%�~�W�h���蠻��-I��c~g؝')�Z"��f����m�-��-f���a�_�]��B󷴲R��&�
�� �
l�P�B�Y}�Zg�bR �?�Cֲ�E���X1q�գ�Dk_��ů��D��<�"��J�$�7�%̼��&X���s�z������X�8��L�l�'�<#!B!��R��NN&f�M3b4eG�è\��5�V��B��p	�?fA�î�vf����e����Àc.q��~k�3͙IF��K�v�m?�NO�y<+�t��s����&�F��)�\��S&��Flo�\�a&��O�,̂ga��y>e�G�l����M���dh��+��v8eV��>�q���ر���l�was���Uj�����jZ�t���D��?��r�y?#��@�I \Hih��T��*�|���R��%El���*ZtI��r�Oqka����O|�ģ6z����޿�bɻU��G0�]6��U�<�=w쿮G���'2i�+vz�������Wd����S��|���(Y��,VY�6C��ၜz��� mF��}!l�l-~e�L�Nj�`<������T0CP�u���JQfx�ym�OZ��kո�>o�P��b�_|nG��\`+!��k�]������(���X�z�_�<+�'�B�����m�Z��R����u���"�����Y��E~)�*	��f6G�SЃ��mş���l<dJ4���U����s�ݜM��sD�C���b��us|F������muxN�\�$Xc;ԭ=0T٤Lψ��s��1�*|��bȡ#��T�쎜����G�U��<~�,�]�4�6��{�8�b�(�mS'[�ʞy9'nGC���r�k�o��h�o�\����Fk�٨��#�lc݊G}W��u��'���%yD)o7�A�3�O�Vv����c����ƕ������ݒ.�5�+��a�Tm�N./ۦ�'�Z���������E����U�O����͚\�
E���§���-}UE��;�j����Z ��D%��@�������E�z�mE���bTǻ�����=_��Y�W�)*�����$��_`M?Q�rt���#ٝSl>�
$}|4��OW�4���(�O������Ѣ��uK<i�}�̾��8�'�sa'_��C)��]�p��	�ve<2�~���V�@�O��2����t�V�7?���/�|xU��ϙ���|�<�5��J�Ԙ���̏�� y�+Z�.����j��4H�֙5Yb����e�<�X�iYt�7���5X���U_�2�c�^j�jk�p�]�<�yT��PAH2ӁHq�Yb�h���l�З��f8�U=��;�m�[G~�����3�Ѿ;{�r�u3��ec�eA�ǧĵ�O}J��V1��
��2�W�(I��򛛐�����r�b��6�Q��D���J�k��)���f�����/��Xq�%��Z��0«��~Կ�bc�mm����\y`���f+�X�_������Guۧ ��Uy�l�ZҦu8��]��C��ؘ���,jQd�f@��1K��x�𮒬p�ب�L�'���}��d�r,q1[X���s����2�Bҗ�o ��='	�l��Q��x���{��|�_R�cԫM��ǰ���&�X$� d"�'&�ְ�w�f�����\y�W�,(1S�>����{_�vG�x�6f&,1R��������%vx嚭���� V)#@r����^|z�ʩ����t��
~��`\�<�.�2���9���0�z�_%����/����O�@���3���'��0�qTTOS��*.P�?�xY��Ń��N�F�ڤ�[S��:-�IӻM����H�i��J��j�����A�a
j����I�j��0�\�l�-����7U����?���6Ue�}C{mU�O:��-�CS Q+�3Ȝ�q9;~Ȇ�"�FQK����k��K��;���^��r&���fb4��R��Z��G�&�2��c�o,�f"^����	��^�ɘ��T��	<9Y� �gj��*kk����Z��heV�T*�h�P���?���[�Ԝ4v����>j*##$of
��?F+q�z��=��y�]V����7�0�i�fR��STi�]�ߡ�6x�F���N�̄K���%0�����luy!�}�.���u���j��h�RW���P5��;xi�rx�U�	����@t�&9R��l�H�*��S�_�ОyI�T@ŵ�	�3�۪����l�/�;�(�}+A�GC�K��b���8��������S"�66LЭ:Wh�KAɡB�������OQ��ձ]lh�J����[X�>���"4����IF�s����tk�Y!�X�@��L���'��]�!4W���<o��ū~-��`k[�b���2�e?F�w7s+�V�"	lW�zTAm�]T,*�n)�S��Y�v��5�wtp�#ɿ��'1�3�a���~6��G���D�e��ǜ���H��B���D���^�@ڧM�X��WBJ�M���~Ym��G��R��������I7+/�t���?������߂b�Uф�U=iLOK~�C�X���{'o��ڨL����*��K�ä�!���W�V�1s�W}݋\���sBv-�Ə_��<��F�/�����z�?H�o�i.ٟ�c�X"E��&������Y/��~����8S�1�2���I�������pX2��X�b�@�
�H��W�Z�9_��W�R���2̊�/����Kʢ<�k�+?����Z�$G�ܫ������U�-�J���m�;�c4�*�q�VAU)�>/���-���y^�H	� `��a։�	����w��iAɖ���o��%6׼	R��N��K�Dp�G>`2)ۅ�$��/�B�^WU�WNEF�h-{Y��z�oEt� V�K>Y�b�)�Ե>����Atx�;�L'��ࣈ��r�=CN�����4�������#����6�����uy��R0뻟"~Y�Bя�fJ�Ĺ�b.&�:٪� �di�#�4Q�'s��/�9�*����I(r���'H}��GyD6�
Gx�1�1��!S��/�xH�=�޹ȃ���.��oh^�|��ZBa��5��i����3�Ǝ�Gq�3�L�K�`D�̸cx?\��c�;�J�-�M-���xI+����/l�|w'IGG���o�Yڲ�2+��4��G۽�,Sĸ^�}w:iB߰��,��e�w�r��N-�J��'��F����2�^
}����F1�+�ŋ�?��ɕ�Z�a�!]\�p��3�q��J����D�d�}#6/�3<-�(t�X׵jݿ��%�_
J�G����'�*��3K��<#�a���.��Tgs���X֏�)w1g&Zk��j[7��GM���K��rZ�u���a I��v��e0�+���J�䝓MXS})���D���l|�u'�x[����c��9r�c�UJ���6q�@M��b�g�*V���{o���Ɨ�y�~y]ޜ�p�-(+�o�<V�1��C�V�����?r_�e-&�/'Z�^�<=2��z��lI~�٠�S��1��i=�Mţ�_<�L���|��DM,�ޟ&��/�;2�/3�δ9�ޭ���E��7�\f����<����DH�m nZ[�^qUwu���#�.�t��tT�e�9�J+K��_i�~�lզYf�;Bک��ڶ��j�Bd]d]h��Wa���+�;��C�,p��Q&G\�d���L�� ���9�F:��f��(<x_'G;������{���'���v����0��HX�<�:4�;�4C�e �o������P���`nӿ���y��D�@=����W��-�$_ߩJ�;�?�����vK'Z�E�{�"��k&�$^��_ө�o���������k��U��삎L�%,{�	�1F[�e��$����:3]�f��ijx�	�R�-Q�#Ǹ+(�V�OX�]R��v�3⭡S��_�q��ieլ�H�%����0i�������"P���@�󐺟��z58)��j�E���Ko� U���TUO��d8S�Q"`���aW�
�?����!W8�U��=�s�X[/�p֍�J�Iu8�}���WY����8�U�tK�L�m�Y�E{��p��{vx;f8��m L�-��%C���Y���ǵ�>�yI���EY�&n���,*C�O{�ALh����� ^-���8c��W�T��(�_.��X���n���E
�����]V��6-�a	.n��+����K��[a�+1���(G��䌷�v��\h�+jڬ�UV� �g����Ts�1v�pw�u�Hr��vO�1�%u(�q��B|�k�4=�+J=��8}��jF�<f^�6��Ѹ���"+��a�5����B㎴���m�{m�a��5;��)��$�T=�je���p���r���Ws����;�/E�sd���sY&��������]�RS��+t�
ZU9�Z2�x�v�'<��s��P~��ᯬ�yph��/��J��������Z�Zҕ"�U�*'�[���6T
/��,�E:�7Z���%_T1wZ�O������@U�]��Ծ>_����R���^ML�y��L��W������=��%��B"�M���P3w���|��
V'�4�.�S���wuI)�����1���Q���;�6����ٟ�c��U�����Е���[9ᄌu=�pX��i9�Ͽw,�|�'��&/^�G��ì4��~i�du�-�����j|��s�%m]�?�}��D���T���}9��}Y�"�@z���\9�U����X���\y��F�.�]Y�C�ۺ����9���}`��7�ְ�ɹ�gl�L�Nd}La���Q9�y9i$a���PѦ�W���b~��c���dѪH�U�wa�%�Xw�W�3U�/s[�~x�b-�v���*�u�M�o�t��f��󗘼�`�s�RqQ�sjlM}U�1�
G���}a���ZWBEt"��)5;���⊭u��o-��0Ag1���F][��v�걾$���E�5x�/��|����}�S׍�M''f���ѓ�f���Sa� ���
�b�~�q�:��'�Z�	�L�f��������CG?Z�p=�,Q8m�����}�Q|+5��v�3VMu�Ԃ���};rRpUF���Q�h�ҭ���؅�d%���N?��>�]��́Ń{|	��>�Ķ�,w�9ן���P�z:����3h��zˮe�,L=f�폑	����}p�Z�Gѳ�d����M����L�oEuLS��n���M�W~�!��I�W~�׭[��D�J�h���U'�C�h��SR�-M5�"�1hs`�cc\�����u���M��K_���ƿ�0�����cS��ͩz�c�'��o�(P�1i�Y\^}4詃Fk�J�x�?Z�yi�h�i��cDo�)���*�&�֡�"�r�0����뾻�=M�睇7� ���fc��0�%@|ǥږ�oa�V�]w�k�ǴR�Q�2f�wY�if�8��`�t�B�D��͢��y�~6�8�b�=���Z�wI����n�T��.�5]Mͅ
~K{�[r�=�Fi3zHU�=ݤ�y���n+�����P��m�(�rc������[��=�ٹ4Za�sQ�:p+{���nvh�qJCj�0�=�t)�W,�ϸg�U��z�H���fJK����"�|dTs:w�7�;��T*��,���s��;�O�µ8*`�(��F���ݭ��t�%�>�T����Pf0�ڣ�a�V
��T�3SI�Bsq���
~��D�q�}���'�*�/��B�]���w��y⯘���yx
�q<@ۙ���"��g��L~�RHTUN����,�x�r�M�)�M?�V���K�'�<Ӱ��H��(B	~؁�*j����������E؀F@��P�E�[��mU73�04�Q!�p�aP�;��{K�Dr���s�a�cFv7;�#�s�n��������/�f;uX�!�ڈ~�%d���)b�v����{cU�^��\�)~?�\��;)cNQ�]ax��*��uO�*
T>���t�B��rކ�ԭ*���C���U�_Q�V��>��p	�3���B�H#�o�����#�k�&�zA��6Z㉔��T�I��������W6�xp���'�mJ���J5�V~����"��pŪ,)����KX<c�c��`�IQWv�ݵ�K4��:챯���j�6�KҜ����@�W���˔VM��0gM��Rq!թkj->�Y�fܦnq���z���u6�HѬ�j刃
��k-�X���c�]!��t#�y5M��%h�@�O�!�_烗U��OGo��Σ�vW���фI*�O�fd ��/���ng�Ȃ�45��H�e� ,\G���ѐ�(��u&��ۄ�gG�ʮ\#%S>Qus�\�-|b��5��\� <��m�5��*�÷#J�A�h^(�hZ��p�T�.˲T"���Z���h��B�;���YPE+R�@�ŴG}����ҎNr�Ua���me����ڀ���Jg��2��7
n]WU�Wc�D�q��K�HpԾ�u���x`X�w_A�/����ھ�Ąl�7.>=[��I��K)�6��I�y�#1���5��v��h��2<uF*�"�v�3I�eN�������7~��fkf:���;9�]��;�ӯ���7ڛ�o�ĥ6K�/�]�ŵ]�0�骮�j�\�M���y�{q�Rjk��X�C�+��
S�:,Z����w�p)�'����ω�>}#��7����+�Jû��{�U#�֪����N28z
��]�LJ�����<y�>�}ԫ�$ڎ��gѦ6,�c �Aϴx<8��!p>�y�����so�}��n�Un��	N��~��w��I	������hV|�E���7��=�#O[K�!��э}Og	,nйFԪ���h����i���R�V>?3��&��
"��a}��ї
�,�̺6uL�V|$���!%Q�Â�_�!�j�l@�}�ߙm��<�7�ٍPߵ7�S�:���
�Ki����`��Y�̅7T4��<h/]�d������hZTJ�I!�c�L�\�)B^�j�p����_uf�QW�nb�m�p��ry�3}FEn܅���9����V:�c�{gW��|���c��Zj�(�T���V�[ذ;q,���u)��:�Z���~boK�U��^��ڜ�O��9.!����%߲��4�����+K�Z)�ի^��#f�UHƥu�ܷə�+�/ߋ�}[�/w������!z�_,ņս�����^����,�|uQ�G�CD�ʈ� ������^�Dl	I���QC�����3��U������>���^~�ep��VJn-�~1��2�Q|�s�O�mި�!�%�Tݟ�M�y��>�Dn��d��\ůU;�J��+���{���|�����b��}˒ U�M����糆u%�Y�5=\)2�wxD����p��5��'������W�Pc=��c���</��̰���Y� ���ZO#u�ګ��wLX6��݅��_Ԇ�2g�p9ٿ\҆&�~����3;�/���&,ܱ��o�@�Z��ڞ�u���p+D��޺�[����8j��Y���D�
�?�pzg�9�Q~��u�X֕�O����K��]�3�|��nYTւK�VFњ��=d����X<��g�r���.�=U4����i�J�ZݖX]�sd�gE�T��Fo����氛dj�F�0����x��5������w__=�#��}u����?7M���s�$������N�Q�<'Ѻ"�N=o%dR��̺h"��B�-2���,/�֍�hU�B�?��I,���l_��3���]�gHT?n���"�����/Y�M��]�1_CfMHã}J^#Ä/��I���g(7_zL�0���y�\BQ�Bz���zs�[�.�\�+��]?f�R��/�+��f���:�`��ċN���j���5m��*��)���za��~.�'��Eq��E_����u-����?��+��y��؝�~q7�B��@Ĺ�^�u>�w�Oq�5���Ń�XP	؟��q[�gF�ʠ���\?NAuj����m�}�j� mGT^A��T���\��o[���O"�>_EW�m7�?�LRz��}������|�Y�zC�t'D`���o��{/O4R�%��}���E�"�c�a���\��j^��!���qT��͔�^jZ���';Qt���F�bD	 �;e��K^+Z�WɽU��nO#R��5@A���2�,f^�,�f�_G?v�V`%����ɞ�E�3�$	6�R^q�l9����W>��ʸjĶTe��S��(�
��q�P���'�=�Ys6���T%0��atU���VN�SA�������S��v�oõY�n�D�}���OVm�ADDK��$9�қ}ك��<8u�w�X)F���T��������?�������`��K<�%�uQSYk{C�V�63��Qř�K�z�)�t]�r�SMlIAk"��q�:��>��	?�Z���|�Z�_tu]�,
g�h^U��vI���A��7Q��U{rhr(b}�*��1���ah��ϊ^}.��O���h��J��A��%�\M��c�ISi� 5|\��&��H*F����Z�4c���RAvC-�t[����,��]�K��C�ٖ�K���K�fQ֚�O��q��;�x��q�3��7TG��DpO��WjGP�}��v�* rߕg�W<�p�4���ћ�͞��)�QE��,{���0(�Z��?�D�e�m��Wɖ���VM#*%�4A��	Yl�]��z&�������E��/0�T.k쪽P�U��������tM&�v���c�V��b�ԕk^����K�%81tD_���Ze4؂�+�mdn�wqŊ�'���A� ��&+&X�������oG��D\@w�r�@�ԥ_[zGH�']�[�S�3NH;���by����̪��<�>����)W�bFa��k�m�¾���r��Q�Q���{UB聵�{f�v��[����V�c�E��|�<�>�=�۵ʩ�B %.�4%@[w�I�}����ՙ��8W<��?'�Fii�*�ƽ�C�V�_���2��8Z�>��T�2f�#�g�lY`��O�/;��뻙��u��o�V���K"DJ�C�aε{`�����K��Io�E�ێ�L��'vJ�Bض��t�7N�j���JSy<u��[��>����ޅ�i��+؇�O�wo��Mu�ew?����̱�<��Dڸr�n<�?l~pE����U]����<�;���\��8�/�I��Ԭ��P)^B�hū(�;�M�Zu�y��^1�$�F�p�`���RT����")�39T?���F����o��D�`cv��}�ϥIatC-�+���mv���_.<�`�yv����5Qɖ���i,�[��M���U���rǕީ-P�}r���q9��0���.�g�u��NLE߇���Zw��q�0z���i�����h��>��E:�ng�մ�_���n�4��x�����"N��m�yp�hI,����նG��=��Ɗ�i���� ��*�v3����1����)ZW�}����� �1���1�l��,�6N�#[�-���_E֐��>��[�IױJژ[dA3��?���(�\����9+�vUc	gs�.ϓ:����;�/���^����㞘P�j�R'�-�����iTG���ӎN������54Ek���<
;�(�Zo�zNa�|};��(9���5V&����K�3�Y��u_��Ԑ�y��>�Ј!��,���X�t��].�*�}���G9S_6�SjlApU���ᗢ�w��'��ڻ�/�d��k^�;�t-1C�l[�4���Cq��F£�g"�H_k% =7}�Q�/l����u�y:�- ��a-T�E�"Uک;~x2<��VA/�-c|������E�A���"-c�!�ȹ����mwy`���.�����!�#�;�rVXm5��l��B3��9���-�S+���0P̓W���]����گ2�.u�/����iMx1����x��Ubթ��E�2]�����9�z&ܔ��hj�
R�#9�2-�y�u��\�zi��2Q�ӽIV��&�
�J�f%'����~�y�{_�i��z3:�C��R{� y�����m��2٩Ӥ}�vRU���aW������T;ײ+�M8U� ��.yPT�8��;nQ��n=1�뿀�d�S-������F���*�ك���
1��Iae-`�gڑ��6���r�U����R��32b
�lT�a_`�'qR����#�ay�W2���,\z��KU�"�|�	�n)�fvfx�R�<�w��X挀ݎ7O��֘��
Zn�}��=������q^�D�:��?\�ET�R�.�t%^�_��s��2�Hɢ-�9kҿp8����g��.-⬿qG��,Dٓ��I�:b�nnϪ�dm������p0��~�lη՗��pW��uX>���n]qS�ޕ�����%��	�?�"�ѽ���H�QA�q�qe^�W��N>�E�3���Q���/v�+�OGN�����:E�񖲠h1�X���)W���� k��yT7����D�	4P35���eڱi��@=V�BU|2�JCv�&��̿j�p��
���o�t��|t��M|��͏6<xƄ_OX�Ri�~���nJ9&�&����_�P���8Ҙz}=���P<�3��k�W���tUQO�i��ًNf�km�L����_:vڑ��[/	w'0��V�v�xk��v�"M���efn���7貳�7�r.���k��X�ȏf;~?�T����K�;-�\�uf�+���@;�,u��J��㿋�՝�bL�c/o9�}�*V΃�k�Gv�rl����
�8[\S2�������m�F��S������ը���^�]���̥5�][n�G���b�<x݆���5�|�.��L�ec��=t��nܵ?��L���+��~f���7+���~��fV}#����'��-���&�@]Cu{���K�	בc���_�d^�Hc������¨\i"���yX���
5�Ҍ8`ѡ�ڷkl6m_�3��4��?�+M�!J%sI?��0�{6��\}���e�0��]B��6���4��5��B=&|)a.�K�6�}�XKV��T�_˘����R06.�~vW3R��ht.;r�������K���U�U����U����3�[��k�'���b:�R-Ɔ�¹ѡ�C1�3*��W7��gv��%�g�~G��՛H ���E�RO���`*�B��4S)�:6֋ѮE�P��ew�*�i���\>5u'�\p���+'��le�e��La�Ft�>���p�n%������?.��׶xN�1�EJ(-�xM+�T�r�C��;�U�1�ۛc�V�C<Z:�Sݏ�/����n��g
~qG\�w��׷��*�������F�2�$���}ː暚n��\2��9��s��#k����\��s�@�xV���l�N�k����M?7���َ2�r��	VQ�T�$bVǡRFkX���֏���,Z�;�F��9ѭ�����p���yR+��x%j�0�`yx�!�L �aW�/�Ҋ�2tV=o�Fo�;��a�N���>�]��!Ҋ%O����َ1�BH݇6�j�@��B6�v^��؍�v.�%՜�yܳ��.n���)v��.YK/S1�4u¾���sZdm��B����
���iK��5���Y9�]%���Ӹ�}��u��� ~�v�E�y�K�bGS�f�En���ǵ�4�؝���y��&��Vd�9�i�8\R�Ȏoćvg�?�aY��-����=F��?[��i8�*U{�־&5[l�V^������؏�j���	s�Ὓj��?��S��;_$%X���E�u���S��8 �-e,ǨI�=�?~��A�?)�Q%ąը]L��½*8�'�wS��D�^��qD�U?��u���R��K_�dL��&�䬺�l�{�#���v�PY玎�Nŵ��f�H���̽�K����	�`Ds�>���%8<{^��aɇ��\�
G�w�͋y�u��+\r�KL���]����%hնH�Z6�h���Ǚ�XhW~�mq0�b��>Sy�ɱԱ���)[��a1��'vE�����1SS���q�~���o�k���qr�ԕJ���b>oDɢx?4������g�v{��UPЬ���AA3�����5c}ҎE|]s��3�|��/����c��A��;+�$�	����V�E�/	�#�U�I���O/	7��U#�7��&�#L�� �QM?��P��_G��r�%	ε{�ɠ�S�꛷g EZ_�RX�:3�ʭ)���odXLIV\��jzu{A0/�x�7�O�~5e�m�(�W.�o�O�*�$r��J*�[��$����l�1���1Z��_T1�R��4�;�-~�2-J`�G�����е*�0�Y��`f�b���&eGQ�&��@�rS��[B�	��:yOm�<�ZP����N��V7�,��6�a4��i#�zB����6r�V�{=A��R�#N6{�ęCS��O�Z98�Ea�U�\k���Fr���'���돿p�<��W�%ک��ɚ|㨟��)��*W���h=�9�)��+Ω�0m9[�P��B.ˍ�b��+�]
�b��[�0����XԱ�.�?r]01��{�]��Oi\����+_�����BB[8���A�4�[p(����<F���TX17u[+:��U�I�Oj�E�y����{�~�39l�>~I�h��kD������,��.����IH�/w�S�P^zI�ɔ�������V�H
bı�M֦��n�t�������FAW�td�����<k|t�re$��%�I[E4O�~7�e
E�~M_�"���Zc��w�Do�4�*+�\$1
��������;llՈ���|�-	�m:���=�B�\��$����z���B����ρ+��F;���ݦ�1_��V��_���Xi��=�`�UA�N'l幺V����%G�%)X�E��*Oq�Z���F6~�܊�$ �b������/#���Ҹ�q2��?��\��b�t)_k��������*�'�J;XR�}��UJGyY�ٴ~�#��1���xF����֝�F/͵�}i�l}#�:bU_��ݰ���<K��}���p�݈��B=���'�'�o򀀿12be� �{��Gƞ����c���m�����QzԲMN�Z]e/j�ϸ�L]��}��GF��
�n�Iڗu�g5饰[�o��L�Fٟb�Zgr��k�:��g-Á����������9�'p&
K���NV�<��6�)���'M ��A8�<-q�7��֯5"'�[���M��H�;�>�\��;/}�N�������
�Z
�sy>��Zݳ�aͯ2y���4*�y�����p� Û��]��ue�'���m�j�*����-}V������WE�P�ٳ1[��c~��kQ:*ͪ�����{��W�31�:�@�3��̆g��KR��|v\v3�p��c��c+������N5�kX����$�dp�Bh��R{((�W�B�OJ�ȋk�e��PC�*y;����8W!�࠭�0���!}p$�%t�Գ^d�t=]%t�y=�������L_�dZ��U:r+T&��]�J�N���zӁ��J?�6�Tԩ��n����!����ǭl�90m��,�S�Z^��;䲼Z2�pm.�%$y�}�sn�ʋ �d�w��#)w�%�CÔh2��BJ����N���.JK��ܽ���V�b�.I���j���x��"�t��~�1UF�Nzq�0V��Bp��_X���X��F�����-\4��2bx��&ek�s'q|1�uť�����F�.��hb����T������D�� ü)'��j��;V��p���S���W���bJ�����l���m
H�hC��_��_u����FLUŶ�*��*��`�s`b�ʰ����Wv�΅�WC_Q�����8rƈrIDf|'���[ȵ�4'�WmT�]ӒR�u�ԯ��e�s�RW�����6^��d����!u��3��~�}54��KV<Od�}D���w�eZNiXJ���.�wՌ] ��ςO6C�U��\!M�q�r8���:c�����,�8!D�YI���/w��%N�'�˜�3�;S��i=��n��?�-��yӣ���73z-�P�h�k���-)U���I'x?c�eX��E�Vt"�_�/c�C=�U��|�
����`2����C�}X/�[UU�u*�~d� �zj��V����_%�+�3��W��?�8C�I�����.��k{U�����GoPL뷧�V`O	q9/Y�o����	�?��D^���`�K�����֟��B���X����>�n1�K�IYj��s���"!�jZZy_���	xs�h1�<|�+l�����*��bk��28�ő{�*�t��p��ͪ�ҫ�ک�v�\B�L`r�.�E�|�_���vÁЭ���m%\2����
�/��n��~���h����-:��T@@���)�1�P��W�ɾz�wY�b!o�ǿ�K�XfZ�p`�l~3��Z=��ృ�;W�b��e�52����1���~��)����L�X���ǵvF��hM�T�v�A���>=�f��
8���W�P�w�ƌ+�N��i��~y-���>������YE�艓��C�3*���~�gd���S�����J}I�y-����x���~�J�w\��K�Е�%�����H�D^�G;�l���T�x��Wr�}�(�B4�t\��W�п�c�G��5���u;jb-aMZ��N����+9y1��R��W�0Z��b��?f\Y��_�7qh��N-V1�!��']3�^w�*�b�5..GS:����u��o=pf�q
F;�`d�E�`p��T�~�y���"�A���}IxA�o��G2�M�?.no+�ɱ��0z�w��]`�B�'�V&Gg��+|�6�B�y�c���1��e����� xݤ��J����Kh�ju�mڂ���@�lܰ~�:��i>��Wax�DW�(�-�>������c| 4DʶO�:P|�_|P��e��N�OҨ�E�������՗<���?h��+귺�KCFԁلd���c6FW:<t��(�g��I���_���}닐+NbR�Jx��6~�ȇ�uy�ǌf��4m�
W.��i�/>�e�y�X�Wu�=��3����hx���^)h��:�l�A�Rɑ���l��Տ�bl�3��"�Z�q�)0c~�4��b�"��k�����=^dE\ ��3i�s�U�1�{�)";��m�l
��2�.B��^��;|r��X����	��-�{�1<E���2�^�MԳ�,Â�N�Lme�z��5�[G�X����ӝ��}Zl]��/��ѵ����͙���{=��f�8��7��Uѷ��6Wђ��v˫yμ���Q�O�c�C�:�+��"9}}`�^�n�}χ_����B��ߔ�?ZeQ���/��k��0s�/���o{P�d����~��㇗Up��M�8`�Ԏh{�D2F|��h�\�'#C��bes|�[t�o5�ȯ��{(.!s�y������1�&���Ct����D�Dk;Sn�^e�4Z��ɞ���v�5a��k�Gy\T����M�D�\W�g!̎�=�3�������W�������F��*�G��f���Y��F'"��W�����ڷ~`��i,�6V��CG���/ٽ
j��gJ�_�l�B�)��@�J��2e޿���R���ԗ˼�ѐ_�_�?��u�V���
�^;b�qGy=
\��<�A߮�c�G�1�Y�fw[7���ӹ�|��M��(�^?�k�[?���p�QI��|!|!d��?�
��W��Z5�7���&Ƈ��3h�Tgo��P:Gt�O�L��{����\�|@�r��۬��BI��X�W��FK]c��[G��BC�{�{�*o`�s����{�7�Ǵ�r�$E3dz�g珖�����q�����'����e��t1�u�"~�?v����.9��eК�gϔ�/p=P��7e��E
��_|�:�Kхw�So�>���*H�j�DD��9����k��?3�'�r�o��Z�G�G��U�>���hQ�i�?	2�����U�+�D��-A�;��Á��>-~�k��e�>3"(��o�W��9j����%��R�[�)�4�4��gLb�Z�|��qp���ze����@3����%�M��R�L:�����:����i�&z$]��<�Z�������۴�?��c�ж;*nه]m���d�-�Xw�b�%�"��]��zY"��j�kݒ+��-��m�;Z+����}u5;}*�������j-w��9�ۙY���S�D�M�;,�m��'��]�n�"WQ��Q�����.Cy���,�XR�.�?�076\����X�g���tG��ɷD=\�X�U�%<h��s�+�8�u����	�%��]T �聠h_�v�K�{����U��_�}@�77W�v(��^��f�����̸���6��Y}lW�E��?	����Ot~��_�-|j3�=�jtOaCQ�zCЏ9�KLV��'J�r�N�
e��	���B�S?j>v����l���m϶j�������TX���!�*��d��Қ/��m�>|6� M�vE�a�������MF�v�ߣk1�`�q{$��tj\��d��۹��38��fI��y{���u#}�m��sG��S]D��J4�`��U��gsM!l�ìNg�)�WD'Xv�D��<�ɚ.דa�V󉔴��	_���u�����#)p8 Z���t��%͜(i�mVQ~�"7]	�]|���)��m	������X�Ռ3��S��ޛ��
m������ͩ+������3C�4 2���x���d�*��&vUdi5�!+Ô3x$��
�=�	�U�e��Շ,���Ce�����0R�*u&�0â|����w���LO�
u�v	�%�k��4r�Kw;�T4p87���j��&�i�>A��Y9yg�Lx��ê���O;�����4�����e�gk�*����LƸ�� ��2#��t�7]��t3Ԟ���]��qg�`ճ�*��P�w:�� ��!��ݯZ�!���>��h��[�įU��ܛ��-hBvթ�(�qQ�Y01����^{-,��L�h�W�7����i�9��9 &�L1�J"�J��t,��ar�hA}_�9J�sD���&���5}I�{&GՖ��&A�]>ٰb�E�X��4)�g#PzQϯ���%���X�nr+��2`��J��QY�^H4��[���d�yi`�G��.��e���v����z���"
7)g�LǤ�$QWoy�>��賰�G��锳8����/�$���������T&V�+Z '��a�8�֘��P��%����+"[aۿ������^�V��K�<�*���܊��LXr��(��lHN4^}.;��ш�5��Pd	�ǃc>��B�>yݏ��}�����il=�����)�,�侙�0�(���W�=æ�O��W�^��Х�u��r_���c�J������%��k�Ja��S����b�ӀW��
j�cs���e�nxZ��E��Z338��M���H���v)�l�3Mx�!�2���Qx���^�Ơ�gb	��z}AUVמW����?���b�߄��lV�FZ#~8v�_5��� �V.��b{T,�N��"Tu-p�6�ë��?�g3}��)���ȸ��3�)�==U���ԕa�Z���ߙ$��h��^C5_�+���ZA���ey��dX��}q�yC����j�b#��EF���z�+vİi5|hn���H8�l%�Nx>v��ﰛz4]�wpb�^�:�c�B#���]�w�|��N��Z�̬��CIE�r�a��GF���~Y��Y'M3D��@�xq���X�ے� 3ZE�?��㼒������Ӛ����E��au���5,!����*�Y�<k'��Qk2��$L��nN��:�͎�(�s�^���'x"ܤ�Z}ǲ�$Xg@r��ENq��-i��6L��5�D(�9�����A�x������9@���l���`���c�����>��XB�.LD���`����e���&$��H�[��G0��źeP%
;F�So�*�x���	�|�p5��td>��u.���]�׭�˨Jd�bZ�E�.9���˿0�Y�N����Kh��<I�囍�RpSy���?�S���<���ŏcw�V7.�y��u=��GMQv�umJ̽���>��B���1�W�j�^�6	o��RY��Q�����}�6h�� ��<J���Ɯ?��	���q01_���_����TB�2��&�`͟l����>�SD+��a&�Fe��_:=e�QÍ�8ǔ��c��}��t��Ǡ�!���VU�Q:��Q�L��$~L-\��I�תDh��� #��;�|!0�\M��`��z�S�B�9�֕����ˏ��۞��?<���yN���)�ܽ�'-�	-�n�FW�B�_q�z����N�a���vE19]���p�:o�j(L��F>��Ϯ�5�_��ooa��c)�����
����A�����w/�ȷշ�*ݫ���oa7J�7�;�3p�Ama�.I�Hֺ�+�@���~h���=�'�g�1'kȄL�0�=F���b|�tY�V/jX鏍�gj���b�6W�f����r5�?�?���"��)�|�)V���{��kU�>p�o�l�����&��C���j����M���*~(��R��b=����Ś�������y,A�Q'}�zT���x��~QV�F��ͽ��k�����:x��_�n�P�W��e��%��WF��r��s|W��P�J�JbK�J�+����m�������+h=��g��:Vr� �/B�P�`����*��e�����`�����ó����_u��'=a�8Wd;(x/rp���Da���gy��V���
T.�;$��Q"6Sv����V��e�]�l�tj���4<��>kO����0�@d�;���+�O��[��Z�橔ꈟ�R�������_si�/�y��K�C�?���ziA�ӷu1Ǖ���lsFb�ӊiJ�t��V�V����&wձ+�����]Y��ֿ����-xx��r?2��TZ�����;����Xb��J��++��S�j*���%�'�O�8	��
�T�o�1����!���d����:��n�ف��9#���*U���ݍpɕ{Wj�AY:�:�N�9�� �se���x�ЬTG���]N	S������ �L�D��+�6��]'G �O��x�op&�q�Һ&ϟ>�����X)�!�;n�#J��e,1��O9�V0{I�w���RU���1�n��ٿ���jp�ʎ��Gu�t�!�t�n�T[�G�3~8ލ�=k�E��w:�7�e��t���*qNxrZ���
�El��]����C�t񽓣�*�g��m_ޒ]m���s�U�`��^�Q�%�r�{�9��FB,��U����Kk�bf��RG�w��_]HU��!Q?�)ɋT�օXj(������ �[ɻ/j�u�%ܠ� PE��'���c�)#��y��-�up�D�{j|�*��S�Y�>�9��2�5:��r�DI]��.����ř2�)�ه��PXI*��
Bb��x������Vu*kI�=|9�!��N�q��wjp�v��L�#	�4�58EsM1!;��v�<W����Ta^�5w0z�n��[���I������b{6uD�bC�o�GJ�JD�u�����[�S�F[9 �/ɾ1;��A�W��]��CXR<ӷ8K��0گ�D�ZԯM�8d�T�G�o݌�k����R@+ʤP��b6.���~N:��Y3c�K/Up]z��vB	~���ԎV�sU�k�Z��f�ff�i�m,�]]X��Ѷt�����f����}�� i�B��(��B�Q�0��tϫ>�Kc	5��7/ڝzxr+��-V׷�Ej�X���ծNARC�3�'Ys��
5/������y���_�x�2�n�ʭ#�hT���z��3O&�r�,'��0gT��rDC}	��������F/#ں��M���W7�"c6�_׶1>��x��*<Y��i��	8&� �,,.kUiJ�Z���2��v3z�����dﲤ웸~|��?�f���w�?E�{����Y>�2���v���
��[��Fu��&�Q_]:?-��R���H��%�=?a�&���Ě������y`�]�����:�/�p��b	=A��)���n��/ٴ���`l2�3qbwT`4U���R'��vy!�w�����Ń���y)�h�F�E/o�*�h`+���\��|��z�����e���-=��s�b�*���b�J�b�2�	�⮀�4y`�6�Te��qv��\���:P����ؖQD��������h<�4#,������g6��$�Nʺ2okP4"}n�t�+�cq��>���Y�
�Z���I�L�XM�#$6�	���'��[���GOD�٨�b(�:����\������m�U�;�c_�!�a-�J�����*���@\O�@���<��*�I���t�f֠M\�=�a�J��uGiX�����pC��a�pU�����G���:�����g�ھ��D3S��^��O	R�*�N�2*�J�����&�!�#Y��{�����_xkVB��g����v�t~�LE�`�@)M�
������h�~�<�}�N�A	��'�bW��0w��y�u�%z�k����n�j0y��m�r���ۆ\(wXڒ2��:���{<Y�����eU�|Nt���0v����xX��;��W�'�h��o�h�S��Í-�Do>��3�ܺYf#�ʲ����k-��p�d���J����v���4�<0�L�6u �x���c^2��ٿ�<4Z�b���t���V �o�CG<�;���@���fq��+�7���|�1��4�w?��2_�6���'H�Y�Us����ʹ���>p�p{���T�׺�K�ڗd
�Zh3�G!�����͡�o��b��h�S��~<"�7I0�K�wn�6�ɌJ�3/[4칿��B�����>���7B�qa-�~��bū.b[o��#���H���E[�$b�׽�2��>�^�e���]`Լu�O�j+md��tg�Jc积�C�p��,�����	5�N������œ��]�8���]�>��+r�h/��2���/r�Q��~~Y�轧��?�j���r��:���t��g���߈���zb��i��a�į<��0x�~��,}��R&� �ݩ��S�B��o��yM5�g\�sv����d3$P�ݹ�d��7�~�ȩw�"{��#�� }f������;��ԕ�/����^�Щ�����
���f�2�������Z�����Ua�>N ����K$|]5'[�����ꫲ���!�U��|#O�����rv#iU����;m-����e���k���q�%2�Q�-�NӔ�����$�[����"�T�[s�뾰�fň�s�X����7͞�+��j�B7/kI�ԉ�\��@��WW@�Qtgj~j�[�����*ۨ�Y7���y�귎,��(��w6�f$�������g�Ә�V��;vHm1�X�\z��,^1U�x�eݾ��Nǁ�G;`�sx�f����g!NK���W��������
�����0x�y��;�o?��h�|%Yh�K	��9X=[���#ƥ�/�����+�����E��&9�sAМ���GG�ƖU8�������;[GS�n\붕��J�{�V��6?Z��P��[�U/�+�}v�@��a�œ+�tu�\}F�>��Y�P����V�f�=j�J=X��d��~GK
���":�FC.�	�/���>����WT�y�p�e���˄��̻B]�o��6�ԭ����<�X���o�:�uF�z�#�(%�7�$��*�S�k%u|���ǥ#��f�ͣ�ߖ��Ucމ�@vpl�s?���A���q�����c>�"��]�k:���R �����*	?|�n(�**�)�VJ�E���4;�dJ���|��D���ƾ�_���~x4�W�i�}��}��F�-f���D�vZ�ޢ�������;��S�CW�zNu�grl�C�k&���ј�+�!J����랳�w|NZW��ڨ�Vt���V4K�F�P+w�gI�����s�]&���LC��γ�7��Ki�C�kq������UD��Pk��gd��/���-`�-%K%>�����^��gCP4|FbS�h��F�m�}���YSb��0JYj,�CN�h�#��f��ȕ��鯎�,?�Ѳ���w�]d�H����~�{�OI,�:�#nc̛�FX�:��ɩ�a�g�����6�M.T�Q�7�t[o�߼���Fh���.��,��B�h�ɫ�'d���f�ᔯ�E4K��L������L�Z�_���W�#��م@�h^���aŢ:���<FTM*py�9�n���E	��!KdƎK<���9��{�v3z_��'�P�����}?�-��lxR�*�fw��`��fCK�C"�;am���cA�.7P�Wt�<i�^�w%u����Ɠ�ܳf��r�do�7&���J���F��n{��?��^i���Nxt+�d��k�|	u^ɱ�$h�Z
L�Z��h��l �hj_1X8���hA��ejW�MͤqL�ov7pQȧ�K�m������O���`�S&Z{�t��s�������BIW56�[19��OV2Z�����z�&��Ѝ&Ǣh��<��"2����^Y3�}�Vz�'�q��]�!{U,1�B�FhG���� 붼�J��=:Gq�(�@�^-�W��&���{~���2	5���#�A9���@�,S'j�H~������!�A��@з���.���};x��V�Y�Lz\���������$��ew	=꫚��fG(�U��g�r��76�\��#��T��r���|�t��@5�q!����}�W%�\y��|���ȹZb�{Ѫ��x��b\�h��������l�G�|� ߈����������ψ�g⡍���t�w����~��9�[~�^_|�.�_�,�����5V�������'�ȑ���e�a�a��Ps���*598\��oX�0g�3�+�"-�'+�$��Ə�}�~����E���c�b���cC_���c�s!��L���9״Ҧ���τ"v6'Tٲ�M�����	�7��e��J4K����bi���.׸2n�Ε�6�Z��)�2�-�ug�Rlޕ7f��hʉh9��
(~���K���uG�\߱���/�,������:7��2�q��fVy'5BE��D�m�/&L��F�8s^uD�	��ϻ�3���I��>��V����Iٛ�!�c����Z�lq>�\���=N��\*�_�9�����X�2�2�q/;�����a˔� uUI���j�E���Re׭W���J_=n�Lj=�������ծ�?gxu����^r����d��F���4e�S	s����d;/��gS��Y�����!��hx+��kf�0�q�Jq�<^�Ԟ,�~��gq�2b����� j��=]gh�������ZeJ�{��3����~X�ZO��>1��79[*�l㌵D敏C��MV'w�X(�>RUl��M��0s���FOu��e�Yfk�1���+�������{��r��e�0�^ή��`�06���v�{�q��X���*-֜]��sʶ��	��,�w<K�q2Q����>��
�J���ۄ�w0��H�I��/կcխ��f����{e\�g�x�v��%b��ʨ��dq��Xl�h�F,��=9tC\���+��f�BR����1��_B�$�Eg�ŋr��oM���R)����O��j�y�z�꽃�c']�ࡨ��6��U��5�����}V�o]�E���'4c_ ��~Hst�C	s�t0��y]�u��#X��A�z��1ڤ綺��}e㟫lx�>�p�g�����/�$1��X�qyVT��A����Ŵ	2�M�B����ً�v� h�#���Ԋ_�y��;�s�U��JE�W��T�GS�F��E���"��I/I��
�ۺ��-�j�H_&���c/����`b�9���-U�E�1{#��3����
�+H�{�4��oM�"ņ���u,��J�M��z	HO.�*���Z�����2�+�0C�����<��y<U��;��]O�G|A�����hP�17$�ר�Kt�~�h��&S-�^%�7��x1����̨�8�GՖ>�&�w')�ݗ���'Bβ\v�Ma���U�ܿ+z����0@_B�ϖKC�گ���n��[iO�D	\�==�CjE���D2W�����]h�1��,И2�+�	�"����i6:�_oJ�ٓ΢��"!�n�[�s����C���q����#4>��2��<�����"ϧ��z��ǲO�T���T$ߩ/������Múd!�*��E��U	P�@��[�TK� ���h+<�����7(x�ýJO�<�����r�R�j8�ˠf�r�����(%���`�u3��$Z�mx�����Y����,�h�����bۊWb}Z����p��{f�{��?�&�$=E�z���ٳ��J��T�Üot���']��o��"K�z�efF���¢��։Y����0wU���ۿ��mЫ (��è�A�����w�d���m�)K)1�L�\g<Z��œ�S�{�˼��z���s���~�E�"1V��Yp�t3]{~J�I�j�Q2}�����b��[�ɲZ��)o��i�*��4�Cm�NIXM�]?+*�t�y;ܢ�!i�

�ޚm��XvD��R1��j����Ü⯝L����*�`w��#�F}gz����7���u�bư�y]�/��`����h'�650M���P����N��nǪ�?��/��ػ�]�:�>F��Je���,�W�����_��)��;�tn�Lͮ5�;�C�y`�Ӛډ�>�u�9��_P1���\�7m{�^f���C�af���j����l��l*�q��g�����-i��`~}�+N�O�!W:����.��nީ���6���`J�[L���.���wߩ�ύ~Zʃ�����TD�չDn�ϛ�����Y*�"D���]o1v��~崬��#�S����Jt���@��Nw��J�ǯI04�����	����+��HO7��,O,���D�@�<���/f�Ca�>p#�QUE��&��c��o�*O������Q��[��O/�.�������ư���!e�Y�7O���F��}�S�����'�/*kj����}��1���F�F����ҵm9�u�C��|+�\�����FH�,ވy�O���u������xC�%A�]�ŀ���0]�e��6�X��qg��
�s��������p�,V�f�a(rpq�T+Mn=e��>�xKr����TPba�`a{U�^�I�/�X���ŧ%3L���-g"�|ىThY��dYz�|p�Ű���>��k�����K�PU[�G�p����.[��ЇY��y������8�Q���B�8UF�>��)p���Źw^mn��������2��m��J�v��'Z��V�4QJ�#_q��D{U��)K����S8���E�l�Զ�y� �EK�M([�e������۠�=b��&F�)c�牺�/
�n�f��h�O�O���%��Au�CZm�Ӛ>����R��_��dT�r��o1��h_��9^�@��(�V���fK�YƊGE��1�,Qͺ�;�X��8dL1��YW3	:Aˆ�y��ٷ�����]4�-y<�)����|����<����'�/5N�;�]�y��:�
׬U{�,q\�B]�s����m�=�p�G�FH�4��A6~��<f�h��-Ӌ��h��.���vJ������N�a�]�!��Ua��^�HW�)�����k��i���3!��/�l ?��N�PW�q�����~ڏ�-&�ZDly��˳C�z�r�A
��|����I�]����u����Rh�U�Ln"C9�?M+S��Ţ�ׄ�ugCv���;��e9��>1	��iDaDτ����6N�xg�B���H���^�X�����%�^,gN�޷=��A��&H��-o��MʇZ�P�7����_x�䶷��*�*�[S'����{*��.fIa��������i�ԗW�����߻.��8~"����c>�A}3�rK��e�r7%�#5`�oOO媝6�aa��de��[�&t\�,�7�;����o���Y�Q�bT,�U^qSJu|�]�:��?T��8�}(�����Ea�1�)}e[��>W��e��(�o0o��b�oHs>|Q���el��^ٽ�ųV2��v\�"D;\������&#������V���%Dԝ���~�|�Y"��b���Y���^�O��o�K�h�m�!���4(	^v�GH3�ri��:N	���^��h�.�T.˂�d}Qg�&�"Z�OI����Ky��E�X,a�-�j��ʍ�%+}�ؒ�u���6Z`A��~�Nesi�_�uk?0��¬&���p���L��|�pbT�3�?z� �M�Չ�.K��zZ�5� U80���D�/�G9=.�?����>�z����p
�����u� 2���W��v�]U>�R�+~��e,��Sް]�$�Jy�<E��L�4�q�uI+��4_Z곾Ő�uW�ę�ͭ\A�]��&�h�Y$cC0�ҕ���<�_cT�v�亡��3����X��E��'�f��,�T�Hg1�Z�.�y�����[���LL���cW*e��"9�?Ʒ�������s��3S��.������Jv���F8P�udh/V��R��]�D1���H���dTN�=_	���pu�ç��
αk��Q��ASE�we�U�{�Ē����K�#�/j62��[pU��W�����B4�N���/H�1��ƶ�~b��hM�'�qMډ��W���U��Q�/6��*�J�|�9��$;�Y(����u��fM�9:����R�Z�
T���5[�ŋEh	9r���x��p�=pg�z�J�UV�nt�\��Vm@���Jq�m��k���K��7킕��Ϛ�D=�E�5(���� :hΚwX�o���l���0�[�#dI��[��i!�*$D����R���僕�L~��������ie��Y�X�����A�y.N�E�u�q>D���7~o�}"�m�I�4Q����}ͽ�4��(��Q|�h_������јe(>���rl�o�r��e �=p����EݳARJg���d��_<��ӂS4�{ճߙ�!�uR04�*.R�g�!��a$h���/UXt����/S�q�}l1U��x�,�$�Ng0�G1�-6��.��Li�<�����_����R�����.����(�~앱6W��B�����w�&�N[x_�a�_���R����ۿ�5W��M��z��-X~��s��NW�"�����{�4<W�	*�VZ��g1\�V9�S0ҋ��j�S+i��*�%��H�\0q��k��=|���^-Z�n#�8:N��
�H�>Q����������!�B��R ]�;��O��W/ϧa�1�ͬ0u���k �M�Q�U��z?���5�_]�pcNZ_�^����T�$WQ]��v�1c]ӫ�*ᇪ��R�0��]-W��X���{?����g��3?�U�9GS2��}��f�У�z����1����tu@��l"���5�QK3��y��i�
��@�~_�(y�Ą�
@�����m��љ����fG)Q��U(�[��w�Jqvͬ2C���-�?����=�O���b�q��J�fc�5��!�չaL��=NR��7(k�#�d� j��Y?n���z�2rT%-?�f����_Z�m[�]�뀶k���c���<�(���S$��mmW�;B�P�CE;V�f{��$x��fg%�,OPP���/���+�4W��bj&2�eE+��2{�z�Z��f�}a�g��������dKq�2~�9�N�~��b��+��r.Ȓ�w�"����Mm�&�u�<f�V���ؖl`Y��y5\Euɲ-	aM�<8��}�{T)���r��̈��6����P��V"J^��y%�|=s���ђS�O�]��(�̠�HH�&�E�I�A�o�rˣ%�L2S֩Oŷ��M�d>�5Rt��%�vQ���zz ps$R���b��k�~��/ODQ:��55~p����:���E�XQ��4�n�	��u�K�o
�T�{I1���ݠ?�����.[Z�~ف�6L��f�Ư��J�$�ha��[�ʄ����,���<��>�\p7|j�bT���>�����qU�퇯���Y`�N�Ќ��>�ö�!��)h��֢R��>��~�[t��"��oC�C�#V��U�6�dV+rA7��뽷ǣ��Da����L�r�Yc�E�5�:������֣㿒V_T.���GE?8Z�`�d)[?�M�[6ݦ-�i\ JR���������yXӤ�?O��G=���?~6 ��R��M�iS�~���L�=�����T��6'9ːD�sZ�\X,�[��� f~�P~�Z�]��.���u0��I�Q]`߭���tUɭ[ݔ��\xzW���/;AF�bYk�*0l/ldQ)@]��I���J��}b����G�dj�;%˞�5)]�*-e�AM+��d���mt�ΤҗHb��'K��W$,Z\T�JT������{�W~W]B��,6��߸W�}�l���`������O���5�fd�j@:�|�z�?<�:1�z�㺅~�aK����'7�>����W����Y������w,j��i�Q�^'��a]v����ylӅe)��ކN2����J7X�
C%W�Y�t�-�tM�Ւ��Wc��X� ��R�>��#�`�V��ҭ�:�~��'��/�7�KS6jUr�h��I��d�'3o�}3g�X�(��`�A;:8힧�恳�z.���s$	��N��U0�{P�<s�Tĸ���je�pZf��|�;�
'VXf��F��o_��3��������/>$Ru�G�s��p���r��͍�i�;Un�v�N�������{�󹻟/��f���InFwQ�ӎE�[(�6*���/a�*�=D�c����%���g�]g�p%�������z�̈́}k�<�1���[etY�8�����=�U�Hz�U�#W�4��#��ƟM����g6�/C�tO�^��?i�j}b�cH�CwT�<hOk�����7��I�Ս
��ֈU9Ec�r��:��~9c'"H9�Ç&[*�����������kyq(�&�"��|�C���Ԅ������Fk�3��T�&Obe��Q����uaN�c ՞`� ��vWR��E�-�X�͌Nv�5�c����⇷T ���<E�[K����j���b*��=\TB�{�Z8>gNGvu����9����ЈsB��Q���h��!�r�����X�hC�ǘ���>��E�ά��rAe4$~RY��������^soV� ���&���%f@�AT�p��u�ᚙ0~E��'%F7ۭ.��#�(���:/����e��z�0}��5<����^���W����/z㳧;��'����B�ocB���y�G6sn	±.�N�^h5Ι2*}��M�z��9��仧���N�f�dn0a��{ʤ�G��gY�ަT�䭲�@�Ԏb��-.Hb"n<,�gΡ O��Z�p	!r|/?bi7���et5�Y��ʄ�,Up�܏Qd%�_LN�]�����`.�����O�VH�S"`�$�V���eRr\�G�U�	��/M�Tj%ݍȿ�E�9P����_�⫥��k��S��i�h�3�,�]�A(w��3ka��_텵�qE��|%�eD*R�.M&����M�o T��������7*��U�b�
��u����`�N���*�9.�2z�#V������ժZ`�֬�}Y��I�|�q��K�{ZJL[��3Q��������`JU�ì!�TL�e�`�\�fJ���'�V@���5��^����-iJ�T�t¿-5/�Y���0tN�V�~��ή�����h٫��Q�A�riy�M���FO�2L���4BzT�{z�Z�����ŷ��
�[*K,4�p�Mת��2J��R���gGϷ�8�����VdZ����d7����]�g��g����j����D����'~7I�Z���+j�#`-W���;6F�E�tZ;��f�����|�E����-�	�.�B�5�S�ϟ�mx�%��K��+���3n�s0V~8��pZho�q����8b��qM��	>�s^
o8�Zɕ6���S�/���xxGIu�v/;�C.[[pm`;_{��z�_+? �C���!��C�|`��ZW�����Pզ�Q�x���X㙚#3M�
P�/d�^�Bh�E��a�@Ӵۀ|C6�Wݟh����Vz�u_�6���������&&OE��=��Qm�2�+�G]��
��Ls��7���]đ�zT'`�F�$1���e����C�D�31 Rv�M ���FD��?����W؛�U�s�n�vDZ�[�k�������r�G��8�uҒ��w�OV��D�IA�[(��Y��ܾ��3�"/���)�M�rOv���{\(w�{y���Ժ 'ؙ�~�R�[�Th�1�R��-B7��vv�9�C� ����dJ�O�g"EsJ���#�.E�b����JZ��;�����
����3�l�<b�s�ýb�PuK����cP7�ؼ�G��'~�BpO]� �l�ύ�vFeo2{��a�n�3�s�ŎT�:�s��kW�OR,��l%���%��7��w��ކ�5^�L^4|�lgݠU�X�	�Oz'�˿�C���u�t��R�jIe=��+v�?t��VH����\5O�S��;UENdG��$+k:1+w�D���j3O��D�J�9�.o�p,آj:_lZ�0�;�C��SKٿ
�Ec������g�)c����^��RU::���}�s+/_������3q�0u�g��<\vL�k����_�K��b4���ް�[�3݊1�rP��:��D����X�,�&�-?�}���^-�B�-
r�b\�}��#,����%��qߒ���	F�]�33�����\<�w�=�U)���mo��x��H�Կ�8?d_Rv�h9�ד+A��>aG�p�uF���Q��gBM��9e}�˗[���ZLje"�M?�t�Gz����PG'��aS��]�5B�aU$d�p9��L�j�Q
Y&�"���eGr"@톦e�_Z9"xz�ڳ�A��.^	�Ir�H�9����W�+eճ{fD����0G�Zަ������}ے��e�=��"K� �T��O����%��&;�؁�Һ��?~��^��%a��*�38�H�)�Z���O�����,��}w�㜱0��6#����r�l��@�N���GG�!ռ-�h��d���u��=`���B���gG�Bz���{nz�'F���� "m�]�Y��a��q�	[�`!#ł�Ŋ'��3�[&�Lkuxo/��,>4��b��d��*I�:���ӆ�]�
��E�_:�E��ee�c���;��~+�( u��_�����ȟ�BG�nT#���k{�o}˙�o��`��eʯN���\i�66��U��3%4�����z����޲td�J�ޮ��Ӄj�Y��[s��.��?�R�*o7X��w��`�d�igS*�p3�q���a���6[R�N0�C��X���[��<8e�[���q=r��ћo_�2�-�+�8X���bq7��x�q�f�����(gt���.��-T�Z�X����!�0�@߮����ϊ$��`���
|X��*C�b��T�������������*{��VKY�|�/f�\�Z��p�����!-�3x��7Q캔��n$_����5f2,�?�9x�����JWn��\����j��ѓ��_d��}O�Q��=R�p8,�Q�����=to�p��ﵐ�%$�T2����
���Ϫ��Wrlڍ�-|o�$k��/b<�TI�G�R������%0a��0��m�dΐ�\��-�=�U�9�mz2�dZ�Fgy��X<;�@#�ߑ��{U�|�#��s��uf�W?�ڏ�S8�N0��%����3W�y���
��hMЭd��^�h��!G���M*YM�iN�q�r���^�J-=�����Y�+���dY3���6m������8Uj�SD��	��oG�!�sْǗU"L���6�>�b&���/�/:�R~`���T}J��i�2�>���C�V�Z�9���`Q����u@(�]�d��?|���%�#_j��;��f���Fǌ�#J���S�C�5)�αh�s����Ԉ��	؛���q�ݼ�����B�B�o�7���<.��/-���n�XC;(�����c��t��#!D�L���joA��A�$*.e_"�,����kXS����z��M��r���?M����u�-��9�š�]�b����Z�XBg7l�%^�Y�>�U��
�~o�;�۹t�J��%Zߤ���a���<��!��a���F��Ta�`������yO�m�a�$ٞ��,P]V���\C�!P��c���m'%����wr�ޕ@�hgr����'R���4:w��?��\�5r�������	�V���X]�b}���.9�3ǣc���ڙK��ܪ��-����W�9\75�V:�.]��;�g��N�%�/w����ƕ�:B�Qp�ԝ��+��g�Wt�hh��Eu]3C
�s�\d�q���e��V(�s�ԏ.dU�"5�zj��y_Z�َ�<=?�I���z7Ar8z%��6��\3F��{���'�|�J]9���:�%�[���{0O.{�s�"��4@8���ܢB�Q�֘��~G���&��g4��S���@�ʊT:�5�:�2�a����rTJj@�����Q�M��u��|�?�^�u��p"W��-*���%�{���m�\��Ŷ��$���S�D9��a/���		;un�&�Pz����Y���4�q��(ue��#u��䁭�j*}�x�k�T���f�~�iÉw|�+�"��ҙn���X��C˭~���4eUu���Μ��1V<d֪6=�'��%��ր��
�3�9K�����xi�Ъv�"5M�C��j}v���]�8�Ԑ1�����[�P���v�KM�x����fF}�-�O]ޱ�;���GN�i7�:%�����t�v����������^~1��"ݤ��5,?<y����M�e�8m&�f�P��/k�/���i�тx!|:�&n)�6J�m�� I)����м��(�0rw�v#���kP�ݗw?Jw��;�M>zV��rNa3Ǚ�FQ;��|q��Γ�����������7rF&X�榥cwdf�s�Q�Je�vt�W��v�3B�$���|���{(�|������G'B#�uE�ʑ��:m�62"���r�K2�	�uk��dRm�0�����[�U#����ˀ��ò�2ſ/���a��|��A:��Ɗ�(��eu�%�m�|��Ӫ|1q�ΰ-��u�jv���f��+EOP�j��r�(�^��]�����8���ŕb3��l���S]ߟ,��Ґ�N��o�|�ع6ms���S�����Wh���h9O�?#l<���_~0�l����_m�H���q�x���yc�����ě��?A��Z��Ʋ�j��(������jkA���w���oƓI4m�!=��^�,W��z��8N��X����h��GU�U���Y#u��H; ?�UT6�)�8��L��6��VW���Ӓ!x$	�̽�3]�9�4UbJ��?l[�D�@A��Ә�NCXȈ��
t�F;�{�<i�8+�U���Ġ%R��rܙ�p�J�ݎRfP@ΠB���L��Z�(.Fxq�K����jI���w����U�o�Uk ȵ6�Ȭ&?gDs��4�/\+1[��>����I6޺��s�Y@������ ��|�)�]���~O3�d��}���s�W��"��#�e�@���4[ c��7��l{�A,������B�7�֛�.S�w���;�,��̓C���K��+���V���EZx-����]I�0�w%J���ry�:B��2л�ݚK��>�#
�x�(�{?t�ؾ�I\I�j/X�~m70sW���o�:5�RV��@�a�ǖ=�V�IB9?[�2H2�_���Sɫ��7\t]�k+�K�<w�y�#��Kt�|�hq��q�s�}͛K:}�>�Nk�
5�et1-q	�O~��Q�v�6���澝�k�E_�t8�N��ȶ������~�s����JU���~��i�I[���>RaF������Ѿ�:N������b>��i�W�Ѫ��{�����~��*-g�D3&�5Ih������g�B:Ũ��R�_"z��+�E���(�X��zG&5��,�E�2A�ܱ��R�6Bn��h����>6]y��_���=��r���F+T�����pz�2V��֮TB-"�� ������枻����)O���B��Rf�+k1�}�?e\Lڒ�U�"K_p�W�poŦ����T"+eTn�W4����ƾ��Ùw�S�7��ݧ����0��=�{��@W8�/��b=Y;�]��*��G��u8�E���8C8�mҝ�E���Tng����L��<@iB^o����w�?���s�o��qE��!�O:WV����&T�A媪I���Q�T�^�MS�~��*f���m�:M����hC��f�S�=t$k�ܝҗ������;�ݥ�O���>ګ:0~�0��N47���vEZ�j���]Z��JN�[H|����<yi�'���V��,dê����^��L�$��M��3;t�F��/v��F�o���8%�F�T8��`�(��ȷ�%��A	
��@z(��?'����&��?���>�|�w�aP;ˬ�p�+�2G����[}1K��եܝ��BoO
rW���@`���u�W��0H(�N�Wq����uΖ�s�葑2����e]�3f���:���$�������ޒ�/hY0l�-��n\2��快�y�F����{O����U��C�v���_��g.s�_��Z}���0�X�U2�H�1S��z&�^��ct���Q��v�V��Ml~�0�:Τ#,�lj�D�P�H�ltFGk�+����坣��o�k��T�V��Bg��J�_��2��q��9?��EU�;�4��۪��Hƛ3�-1s[����,*#|�yP�UJ�¶�M�,���?wpe١�_9<�/���v����ܕ����j��v9'�m���Uf]�&�U肟�=�d��i�Ѳڅ��Պ�&/]�>���'~�7qk����!�K=�\|��l��}��m�W�r�U�$��T���[K�����]���` �1#!֚����8�cr��j�ĩ1TY2�6P��j�˛�'jvQeRX5����=��{8��Nyh�n`�BFT~$%�;u�}/T$s���4�ѫno�Țp�2O`ȟ�m�O�=�r
���?|j�*$*��!���tO4<��\�󿶾ۮm�}w9|B��}ا>�6�wҔ�V(W}�R ���f��]�#Z�I�Q�I��o��yU�Tֹwx�H�SxN�U)1�� ����NdTuLS�.g�xCfV�y����)��MU��������Y8�Q%�>�?����c�q+)���g�\��Xl��:�q+޶�WU����������.y�GV�C/$��z�(e0�N+7#�[[Um�U<�מּpIgZ�2�p1���N��M���č �,6Vĭ��o�������X�WYo���F�M]�aL�=��I.;>�N	�o6(�R<,c_��.����/�N���,��qk�Z���p��q�����?�hL�KGI+�+3���*ӓ�KHߣ)F��e �Ug�r�`�M�7�r�K5�5��99B�Z��������w�����[:qb`�<���t�0r~Y+�~��^p󯓷<[��c��J:�40x�Vٚ~#�~;�7���)����WU�3&P��=<5���v�/�"C�K肂Tf{)(.+���t��K��.!�~�:�����@
J��k8O�ff`��)�6)$p���Q��7�r�e
[!��n���Y��OMU����6"���H�����.�Y[��s�H>��لlmm�N�~�;{b�w�C��+���ȉ�5F,��Z��v��bO��7�0:��)rSZl��q�{b�BߚG��I��N�g����!����b�j.}�_�~Ɂ��K9���9�l^��`�����(c�������,�g	h�"x1��ٸE�p����xt�&��W�LQ���t
]���\%/I�Eߵ]SgF��e��>��[�(bw��I�*��|<��p5�{Vx99g�^�L�(Ń���JM�6rD�����奔��E����~!�w�
yY�?yI̱��<�;S�����
K�d.躧��D�ƽ�Z�<���LPʹgh��ݖՔ�{�^�V�FDa��Yn�vu�m�3�p��/.ۘN4��(��T�ם����(�rvAk����o�.C��ug��e���>z����3��H�ȷ�\�Yu��F�D94IEU��9�Z+�]��No����l�u�W������:���<i���K�K���z&��yU���8���ھGP��/ۙ���8�Uy&���w�=�T9�ρ���}2�ں~h��	��'?�zſ�L���uY��7��mC�G���K��O���OGgA�~�q�T1�*�D�'��s�v7O[�$�=����*��h6��1��`*_�r�������z�j,j�Ҡ|u!�+�>pG���&#�]�X<`	Q4��W��1kwÒ*���F��{��*��!~Z�6��Hc-	�0�?�aF��N��Mw����.r���Z��I�%�2�~
+ ��k�8{��+df���s�����T���6W�gd�u�k*J\c�Sn���Cj%V$�+��JrC�U��%��R96I ]孌�#��4jI\��rx�'�:%V����]��Z��,=��Ͻ]�,AT�'n\��8�^
�.�F��\�A�+�c���ë�z\ҡK�rw�h�0�J�<wW>�8r��/`YS����-v�6������[}���[%�T�4!>�b̤���v�}�B�
�$m��=��,�_�=��n�d�^���X�[����1����A���߫�gx~w����G>ٝB�ݣ�b��a��|�L���5�w;����n���{.�.\�2oJ(��ڨ	M���&Û�	�uśW�����q����������k�]�LK$~�xU�٣�m>3��A���a��m�����z�[����8>x��OL�����c���Y+.���=pkz�;�X��Gy����m-���ylr�pYLG��!Ɋ�?*��G$3']����6��ߺ
��.Y�z������8�+&V��B(Q���u��1H%<8G����x4��A�Yz�"���b��|���u���s1m�Y��F�ܲ��9[k�C���%�����a��;t�InV@���b��kJ�v�3���d��@&���J�����[���U�&.��;���b��R/�.�1�Z�3�v?Eg{��%*�ǃw�㇭@�k^.�Z�s��ޛ����S�R��Ք�i���[b�P�����WՎ	e�}j/�X+ؿ��Il`�p� �ysɛE�e�,����~�aY����al��ߨѨ�k��"�P;��m��&?�y����k�Yh�r�(s]D��O�����oYLw6���&��t�K����JTrU�k�T/�w�%fu	�i���<��;�S�M��W���J�
wY��M�(��|!C��!-��"O���;6�����
�u�^�d
�p`f����u��}g�B�$�vJ�|壉���~9l��ЫN�gr��q!'��W2���=�$倕�c߳鼪��G�əك����9|W�W͡�R$�l�����3�X�(�0����;�����V-}K�O�s�~�FEKV���Ȋ(��)YG�;������R	���� ���O����1�yĭ������V�Oeڰ��E�������!Sy�4�?F?� �;�bk%��)7M��W�(���3&l�:$�L��.��۰;=I0�-:�d��ќ]6 V��G�6+�޾t�e��ж?�hϨ��gX^��'q)���F����P G���������� `vՂSuq�C��O�7�n������ng�UEe�9�k�l���D�����Z�V��
�"��|�i�����ˎR��pzY�2.�[������T�~�s)�	�f���=h{�|�]t�tю"a�(� �:��Z.��[�3β���E�����6;��e���I���S��1�Ԍ�f�-^��א��z�Xn4��6���F�Q~2}%b�Kҁz��������e�j���h�$)�/��u7���7��v�Zy�y�;V�&�N�����"`��D��o4��B��b��qi1���%"wgJ�_8l���}�mu���#Ƣ�#1�<����8�yT1拽�(�J��"A��) �o!�h�/0Z�o!��9V�Î�rU4!�m�*g�#�"��]�0E�%)�D��*^��b�0�
Q��������}�?*t���sMuD���,�.�g{���y�9���.Qi�*En�1و�2�y�SL1'{����h$���a�W�K�>!�:�mԘ�{n+��Y�5o�ةˉ�r����G������Ӏ�&A�:�N��7��;ޚ�b��F_�C��1r	���~����֛�$����T�ݶ�P��/`?�׈�u��;(�?�s�@��xC�-�^�7w�W#�h�_6;�x���4�l��a6Yea->�$L�yC'�x��+ʭ����鶌���x�޲�:�Q(H��.$��hln(.AC�"�o8�r������m���g�f�j��mNd�A�x��b�몪M�4��MrA#�)�(w0���̝#�����Y���d���H����:qYU���_�c+��\%V��!�`FG��5��bP}��ɧ@��j�L��'�\`���\%��'��t߃���e���Kݤn���W@���GL�j��ŗ��G+���R�z��!��X��� _[�]f�P��:}q�D��ܒ�o됝�a ��/h;gm�?�ruϣ{�c�_�v�VͯH�-&�-4�ӿ�j	����e��?�e�7B�忸E�������ټ�^A>�m��n�(��4+>�(1/F=U:���d&���S�?̢����U��q���y����@��<~�!"�>L�R7��%+\s5�,��Nj�]���EԿ���}�w|�}X�W�1�;����뵍·w�K=��?h.k�K,��W����gy6|]s�&z�l��
"�YN淣w.K��jq��E.�+�tE�5wU�|L'��Ր�jUK�2���<<c�O������4���zh�<Zӫ�L_}�a�`xO
\��\+�{�ϖ�/qS�S��X��g�N���5�ny`���F�	ĺJ!��R�P�����;�;�;Z0�2C��'�;m��:��J��N�:��	Y{g���nR�WC��t��*?i^~󯠏s|qL��?x��B7*�:�w��t��?�'��7�6I���W�[�U6?��gpF�8vBc�
��(Z�I�����O>9U�9KY��K��ŕQJ5��Z�]�v����¡VX��6�B�b$3�\����"6�1^N����BZ��)��c~J��=��^qP��Ff��w�5�R�����&VR����T_U�C�PK72����z�Ucsx^�;L���}����>p��y��q��<����E �$�[+������*"S�u�^Zb�,�����*�gr��F1�N�͌����U�RLԮ����D��7h�>Eq��Ի�ti?j��iL;������G�&^=���N��M4~IY��v�SϬHFhW��@!��,C�3�<O��`}s�0���V�����QG����G��`�����>�Z��B
���MRU0q����*\�h\F�]F�4��]�Ɉ"�g�rRາ֝��sL4-��-�R��������3
64^=��w�3|8]�U�/�g���YBT�_h�q�KP��::~��AgK�+�B1�(�*J�����6�lu���E+52hg7�$J��9��`�M���4a*;7R�6"7��ku�_~#�!��-����a��̯D�j�S ��Nv��Y+��eGƂI��|ݍm�&�:/i�����I��%�~؅8b"u}���+�z-���:�	����t1�}M���=��6?�Ȧ��[��	���L���������ș��s?�,�s�;~��ݣ�B�P�4~��m�"�l���:g���:�W�C)�x��N+V�}'��i�l�����Z��+��J �#�o�mb�B����c�<����YB2�g��mwgqM"�vN��G�Ҍ����5 �6��k^��|��c�Oa<�D��|��u���S���K�څm�&��Mr~C���ߦ�C� ���6�}����2� u�Z��H��œ�ָS��&�#��kX�����H��R����!��#n8ж̦�b��Ӿ�1lp�h��r��(�;\�{.�Nn����,�sIk��}�`h�%3 S���P�]��M�?�����^)s	b�������O=���9ys68����bb�VcK�)��K���	���W���k�����fIX��l��_H��/zw�4�a�D�t&�N+������a�)��7�`
�M$�q��]>��Il�r��ߌO�&�<C���K�/~׆����Oӧ�Z1&����	9ϱ��m��<�6⻾Djݵ��׷�bƪ8�?��#��9YR���/ɒE��7}�Z5}T�4uE-˫8g�ߢX�1��gm��.L��5)�3D�1s�1�\4]a`���^w�5���=�ŏ���y���D�����*ӛ����D{;a�R���Ӽ�7Ua����.��hC�>p#~��R�C�H`��ٻ��X��£q����e$��:b����R�������[ A{;͹gQQqu��֧�$��>"�w�/�N������:<��.�L�e��2EO�( ���i��o�s$���߿Kf�Ǥ�Qqk]ZWP�:ʉ�+�0��Ubju:?���gu��M�Q,	�����x��d31����Y�^r�é�3�O�C����'5�0��IT3��m��q޸�S�&m�'6�������܆\�٤h@�|-4bؓ�Mr�7�V�����:��/��wW~��R��zA����N���^}��2�v���K��[{����(:;��F��*��1mq��_(G����S�E�ә�)�"UNd%����T�~BY�͍ &m��le�z窣��7Z�k�^��� ��cO�t-܍}o
�_ECV�P䣇����x�N� ����_�Oɜ�/�A˧��!��F��5�s���&�����Q��s$���0��E��Q���1Z�V^[(ꭢ�����k1-Yf�a��m[Լ���Eh;�ʖ�y���,�d �"퇔3�c�ɫG+�⽎���#E�^�$k�΢� �t׼�>l�>|��ʁ��y��?tXϿ��ZBuW�Ҫ�^��Td�l[�Ф�����~�!��k����ߐ�:�+�,i"��m�(A|.
��Û`4�jd?�q&2���B��y�VU��0�X�R,p��v��Ĩ4A�2x��)���(�.%��v^�f�������L���<q��Y�<�_�/\���w#i(���[�5�t���#{��I5|xv��1��(*�ٿ�h�_J`DQ�-`�UҞ�3P����r�������kn[I9_ET���9���%,�d�4��f�ގv����k���j�Px��e�_À��0�0rl�]f��-N�dZ�\7G�`�o&�U�X�I_"�j��V�Ȉ����}���4�Tx��_\5eU�3uv�����@��U��XH/�]ɗ�
�)��"�U6��а��T���=��mMi;�*8�..����R	�f|�U�	���*���Q���3�������_8���~`�wb���F���_���JC��Y���t�aV�Oc�;Vu��|�`�b㹔�H��F N��)�~O�`wNP��R�7MB$�8�����~Sb�_�bY���[=]N�ʗVy�7X���Vҁ
uRB��ym|���\}[]���P��3��q7J�1��h�����1�L[��f��!"eĂU�<*Ň�R;o�����O�b|�DK�-��e��ߦ���[W��~�������ɂ�a\�,�Z��'6q2�\���k��:e&�������q����t�+d�ដn���i��	�����\~;��4}��$�ߓ6�_�2	���"�j��:�1u��i�T���^j09І�	m�!oA��~9,Kd��M��ɿ���$�e�f�ulo����O���sd�R �W���Iw8�%�	r�E_�3��[��Je���w�J��ʜ(���-�A���n��_�75��X�(����\
k���E�����(|o��o������|�ɲ;��J5W��{@d���0��CfY�M�m��CA����юN�)n�M������9�f�9��/�Q�X�
���c ɟ�����v�_i�u��!~�����U�U�SĒo*;�����(�V�SL���'{ ���?�ҧΑ����*Z��!9��f��������>�.Z�7�u8Y��td#V�7�='H�mU�1�y%s*��-�����"v�]��b�$r|���W6�LsW����&iP%�^���_���x��:dR�L��쾇Zs=���{\�<a����M@�PQ/U[=65�����E�.�u�x��g��٦�c�Zvc����$��A�]�:�d�kd"�o���'Cm���9B���)ʵ�Ī���r줖�|(Z��)$\=lnJc7B�ثQ�vv1�u�E��%��0q��[2�T�r8�pX[`���X5�O��Zk���qx��{M�_���3�� ���Z��_��=Յx��^"3O}��>�Zhn�����+)y�7���3VK-'�{��`J�s��+F�]��� �}�D���B�Kv]��Oir�蟖̳��~��5��T�>��l_`�Wc�<pŶ��2�L}N�Q�EÞ�ȳG�h�?J3[j1��;��iXɨ�}0��-j��N��I�H�5��/O~���G���|��EM����[E��1���L��˩�j�?l�P7����xL\�T�no>'N��Ck	����޸�B7ö��Rټ�5����Z�,�N�s�����~F˚����Jp����z�:�?݆4�諕5a���<r�χ�^�=?8	ZFZw:����O�'�)�Ŕh�:7�rS�u��`)�������*�O+�R��cO0����9���@L���~���<��Q��u���ҿb�%'�;�?��yp��~8qO^�c�,�ZF(��Sq�U�H��.�9���%:,��0��Yjy�F���u`��`������WR�8�D
�{��i1�o�/#��楓�Ȫ�w���e�.f��*I���d��<\}c//C���ް���6�Q������y�"(٩5���]j�1���ʯwG+�:��,~�e ���̞ݜ��۸�<����f\��i��[7Q|p����U��u�ퟻ��B.1��r����
`dd�̒������G�c
1�d �;����U<Uld��4X�X�F9�R�C ����ZH�y!��
��n0I�hk��>�9P_)��L��p��,��G��^��e�KܻR[�KP
#��9Q,�������iH���9q�s��M[��:��RYRh��m�v�/�<�rz0E�\ ]p�����Y��=�$�4�KY��>�b�L��,V��^;P��������ՐA �ǘ��#������n9K����|�Dk���gT}*����c����N�'����I�>����]�����VK�[��Bǵ>��z@�S��K"��x�2��E#k?5 �R��Պ�?G���"�/?"��)�����n�e50�>B�˦�<�E�QKG���2Vd
~������ָa��o��A,��"��9�3 �Kս����MI&&&L*m&F�ߺ�\/}l�\K��ڤ�?<�_�bĈ_'W�a�[ɞ-��Sk���7>q9/�:����Wm��6R��`W'C�ѹi������\��	<3�t�vҧd��ۨ�˖&Z���D���k�����ڽ��_۵awCº�J�P�Z/27�I
�?�9Z��e�[9�/��Mی�er7�n/�Xz14j��U�[nMoT�(�(_`M&�DQ/n^�Y��'�TM�h-ٮÕ��ε���3H۔��P'~<xW2�1(�uѓsͦ�g6�g�l3�}2�����yE��ef�6��[��=��s�hy�k�9RS_K&�r�/:�m����s�Y9o�� ^�K(�N�k������G5��7G;�p���ʤxppꟲo�Y��C��c?f������"_�~4��6��hX6���Z�ԉ�;?&�XFQ5vӒ�NM�/���ʠ�d��0�=�^��a�����:�:	�B=����Xo�I�����f��(��՝�ڧ<{z:*�[�����8K�8/�uN���������y]���#����AF|�f7�N'��y��<��J>E�	V����PV4�'1³`���C+�fH��c�I@�����`����?$�2T����m��nv=�����֡�������߳�� Q�`G�M� 'ZJ��#��y����l�z�D;�+*��(0w���3y�q�*Lw�+>�u�����9���Ŝ�׃ ��`�(�����D�h�#��}�WÂ�3J��dWaiZ�5��it�ޕ�(�j!�����3�5�(xH�e?������/p#�e���ü;0��I�M���U��

��)1�|1|��Oj��%#����T�¾�Ă��K�h���B��z[疧������gDx�+΍6徔��Xխ��٦�` ���h\�ȡ�f�Rqh�;,[8�z��ޛ�?��]��x��$3�4.y3p�je����᫋�:���Zp�}�u �Kwa3�g%��}�?���*��7g��N��;�kz��fz|\�/�+�s�_����Q�n��p��X����R�<x�fd���s��z�"d��"���!S"u�bo��#c�-��f�%�����������Ɖ��q�Û��Cm�.��vf~e����'�!f�V��@��a����ר��5������oԟ�S&�Y+�#�wY��]֠cC�Ř��B�O�ڨ�G3ۓ33W!�:�&���1�X����M�Fk,`{���)*c��d�1dGK���Ĥ��o���"F�����ɘ6>R���S��]��h��b(���clE��Diu�����뫷���	a��Ql�wX�ɔۻcn��n�=[/�+U��k*ҋƾ��l4�t}"�����^� ٔ��=16M��z񡯖kl�J�ϽA��+7�g���F1s�`�E�uf�Uv��������a���}}��@�����{w��c�]eu�e�"PU��+>2�����G�S|)�%g��*������D����R�c�n>>�����8��&�Y��m��T9����:ڟ�u�W/<b\�������_8���Uu5/xhJuѶ������H���m�8��O)S����ǉ�>��6������nJ�F��Q՜w��׼�Ǝ��N$1F�U��Ϋ���f����X����[��|���S��^�.�Z�,A'��.�j�,�?SU�d?���:بN_S�������ʛm�v����Z���ݓd�Rs.�;,���/��+'��2�M ~d���9��6~6\�L���=Xxj��d�*^5Xpc��۠.����S��-��M���#���X}�Z��¿�o}�׸Mv�R����;< ��(�D{6����A߾��>��\�@�[U��EQCq˕� e����M�*(�
cDP�]i���²�����uԎ���x�"7"Z�7=tB�Kn����~��l'��t����U�?��[ ֌7�g֟��+��B�.䃓=�᪼���T~��Kn����]`ӊ�smW��h���.�I~x�9�
{.�_hq���<9�/k�&�ޝ��B���	/�r��:��"�w�n�VJiDr��gl�d�����W��*C	�[t�0����\��]$���*��~�Z�m�~����Kӯ
t��	Y.Ϸ}����x���W���c����F3��=�Y!�,��y���w��)�y��}ޣ��l.p��A_�
%�e�A�{S���;*Rl�]�4T�3~Q�^�#E������uv��/܍�VΞۻt��,~rq�͇3,}�Eg��U�W�wV[>�t}�	S��h�/t*�C���H�����1��!Ǒ��j�9�T�j���B��͞�p	��ټ!�U|�Y�]\���-����κ��\+R�=Y���I�2Ž��e�%�%����*zA&�-P��%�������O�.�T�C��/_�X!�ౘ_�x��,��<���J�� +�o�Z'��}��u���9NF�{���b�)c�I�"6�S�ݥ�8  Fz�~\������[&]=��+��sr��U�*W�����p��;Bm�=���N	W�ce�8W_��W2�gMi��c{|p����_!�f.�Ƒ�+��ȵ��1/�xS��{��*VǳD+|���jsF;���v�������������oJ���d�Ϊ쌃�d���C~�!M��]#�*�5?�fG/~6�@�''랙
����F
ꜻ�q+�_~���iq����ņ�3 <)��>^+�n?u��aa��9��1��5fqT�����j����e5���_�Ϸ��z�������ߴ�Q���~K'zrЉ�6M����_/6i��%-p�'ک���^�F�xD�dv����U�7��S��mh<�W7.�_J������@�N�·LDP�W�㏇��v��(��ܡ���?`�zC.Ց|�����Ƹ�VD"w�
�n13ܽ�$���H���_v����svצ����o_�NgP�k�b�������F%��,��y��1&!�31�G��Uup_و� �6��2Z1,[^BT���A�zW��#�O�/�hڰ� �n��F�D~�8^�}��c�㧎��E���C���z�0p�s�����^�]�/��[�H"1_�n_���S�LC�@�է��X��y��33$S
�g���6+mi������:��,����5ņ�C�5gldf�/j���9S�B�˜mf�|_~b��)�n��6{]=��3c��L����K�0)a�m�w��I�]��\l*���N���;;w�A'�$�>�i��SU{I���Wa�
���y6Z9>\7],���H2X�� ^&|��;N��ڣ�G/�<�<+:z����"^�c��t�z�P�Utܨc�"3 �vQT|�HpZc��=hl���8�
\�=�)Ǩ&�A��;=2�'e�����zֻ
D�����=4����3�v�Pb�ě "k(~�7������J� �Yk�	����'Zܢ�r�/p&�bC�T��)����k�ecA{��|��1a������%C:��?�͒�he�G�������`�V�\�ꞡ�h=����S~ɷ���}�.�A%I��3�X����/~%�-�����'�=��3�Q��VS��(����w}Q�g����3��O�-������gN�t�sׇ�Lx���>�說�e��~8
Ʊ6E�b���On�U�V�&�tY3�N�h.+�Ҋҥ�$Z]�ħU���[�"m�?��İN�:���<��������o���w�.�շ�.�J�}�U)�i��~���(UO��P6R���B�~#��=��HK0ΘX����튑椗U��+���L��̣�^t�[=t>z�����x����R�� ��KN��L�B�E̷O��z&Z��i~ޫ��������R��("o}Ȳ)����A贬]�I�\ �YLF6/9�z�C1�p����]yr���֡�\�a�����+�&��X/��P���vд��G��y�����-Q�wDB�F�6ͫ�:��FC��:.[0�*|�uS�h�0����!�3�\t�A�H��Q4����K��υ�W[�>��wB��>�Ҟ��g]������gґ��Y��#�\����ZJ<�H:�%+�"��N����	?&�����|��1���ē��)�^�%�xϻ����hv���'��C�H���Xz�����E�6��ob��ƨm�ј���h'�l#�����Hr�`c����K[z��C��~�F`]X�]K���q��1K���c�����3{�{�E1����c�~���ff�g�������� �?pl;�t~���l08���}�)i�.|?楶S+}�����2|���������X��G��* �غ4�����y�� ��~�:À8 �p4흰��x��sU�R�;�,�@a����栣��.�NW�:n�����:w 5d��*S��R�l#�姻�E����ٲ|_��3(ĝ���)b�:��0UX�SF$��z���b�cE̽Pg�Ӯ�K��%�+�9�_�{�i���!��ǀ�Z⁭߲�m�g9dM�s.=p��q�͹0Q�����$��f*��<�g�j���z�լ�0��r�nXY���[�>��=��(�yѾ��tw���A�ߗ���)���8�H>�~�Q	�h��m_���&�rR�O���Ż�_]�h��8��3?<�ч��P�m�{��V�����|��\6����x|��_:���E���������7D��K����r'j�&V�]��+,�]1d9��6�@��Y��@�?��f�W=w�L��?Y!�+R���r��*����l�stG�N0�!��Ti�+�؝8�LT�����A��dk�����~�'�F/�TÃ=8��*$7#{���y=�q7k��~Y-bK�s���I��#��$K�v�-R�+��0�z��~��������)|�%������	����?��G[W���U��Go�z�v�7e��4E�K�JRޫS��O�m9"�&��4��-u2n8���UE|����(�!��K��1��i���T&t��/S0pt��Q�H��=i>���e�
��Y���791�U:���B��Z�&�x\UQpk'�8N	�K,qm�;w-�-�����%F���ǜ�M�Ȓ'�*��څ���+b0�S�0]�Z�:p?z�ĽJ����h�/\E������o��
��iF/�ljތ-��f���wp)��6v÷~�5�f��\~��3�`z�hZ�~�T��/��sTfz���.-H�o7��~Z_��{�n����6f�~|��ԋQ2�qx�D7E+U�����*�|�ǿ��fR�ڟY�"F�ŗZ+Lł���C"4����]�Mޑ��<�1ݢ`O�G�H�w�ep1(c���=0�ܼ/��b�t�9v�+>��ًᆭ%�q�1���Фv������x��羵�ttE����hZ�)�亮��k|i�p�D�u�V��dw��5�n�6ױ�_��w���������p��ɼ��;�:���AQ��)Ǳ��*V��\�A��L̫��6�܃9K��}i�hR�E�����kB���p�qA[����J�V\%�e9�R��W���H׻;��j�]R���Z�l�*�/?��B����O}�����-�Y=�y�y�uz�H�9C��@D���f�MqhW^F�+������#k��e�;_�X��c�#x�~�2]n�Vcd��zԋM%�=b��n=X��q��A\��8�!��~�����;o�L�D|MJKK����O��W����/+�N�df�K]���n��r��"�W%M�J�Я������F<�-RMUt�Ht_*�0��V�U��<�(N�T��9W�^g�~�+��2͔ۯ��'���#��x����2qۑ�'������jD��,�� �`�����;,`��r��2݅����	j3
Wq�A�ل��c\�j}=���A��a�Q45�H�+�&�%س�e�g@�=.�8:�#y�t�p�n�;��]��"�&?��iT��nNH����*r%=�ޑο%m����_�|f�2�i*k�Wƞ�kA����2�����|o�R��0�(�*�M} 
L�{�"�?%�!�M��A�ѱ˟��o\C�tQ����W����r��9j�X���|�����"�L��R�-��S��k]�p�å���rP�`�%�sD{�:�(��& �_D[��)�J�<��\/��Id��O�y$,���s�8`4���dJ�E�[K���%NWx��5@����]D�r_|w�\���|I�eLf?��Ƀ_�>���-t�GF|*�+�l�Kڂ��{Pت��;�l���*�N��"]�k��%���/���k�d;��@u��K�݆2��N�~�[��jK����6|vs��*�"?C��������/���LA��{�� ��^1�;>_�f��ur		5ެ�bX�������e��m��C��_�b3�k9>����o�K�DH�9�/��H�\�ڲ��B�|U�6qaJ��OV��(h�Z���85a����ܿ����5�������d�זoÉD�a�l^�>5�@�a��*��|�O�s&�Ҫ�=h��!qj$m�O�Aug��յ�g)��n�\<�#�&�]M���?Ya�L�W�J~@�+�+kS+�%ښ�������u~[�T��o^q@ɷ�v8��:{�R��Ҥګ��L�-��U�{�F�}�{F����AI{V���Y�:�Hܴa�I�Pz�&���y��R��:�6���]l������w?ݶ�����R�����%��Hܿ���v�o#��k���s���M�{(Pzՙ0~�J���N��i|���U+�/x�<g�f���s�ۚ�r1��l+�<o����-����C��9[�x�J�Mߨ���_�����_?��+%�V���3�~��v�;6�/�"��q��.mՑ��R8mO�T\%�0�]�xq����0c�^��v��![�Re�h���VI@E��#q*uh�v��1=�'Fνӎa��}���_�6ԭ��/2sU�J�{k,l��нa5Bu���(�b�> ���R��3������셒����"i?�}���&gJ	'*ui�Z3�ʼ�/h�)���7�����*F�0k�f�VE��$����N9�m�5�4P���4I�X�yF<�N����L�]���gĎ�L�N������@�[��I˃o�RѨfr-����܇������k�ݾWqY'=��S�B����ז�������*w������C���4�#JLŝ<g!����n}�T�u�F�Э��HR�Ũ����N�k�%��5Wɿ�r���	$*a�"��Z��m�����Χ�<A��FJ=�����W �G�3���0gG>�sɝb=��p��.��8�;��	����쟣�	�Y��??������gU�U����j[�E;���c�N5,k�4�oc�+�%��� G�s:nǔ{�����2����]^\�,#��V�U�'}D�Vs�h#���؟�P���>E!>����Z������DwX�O����
�]j�1�hd��Au���jmxfT�mJ���%��a��ZT�h4c^�X
~��3����3�[|��O�[�-�@���O����[~}x}Ľ�+e"Wd�J�N�<@�w�8թ�y���H���t~��0�2��G;ա�Sd��מ��Ψ�ů�O�����Yh~1Tȁ�lA�D�F���8~2}�����b�F(�n6�x�R�
늠�p�����/��	�B��7/S�u��8�k �T>���⮵)����V+��S8Łc�������'d.�,6�W*���L��?��:�����lj��꯿R�X�{�׍&�ĲN5,U��^�:�v��Y٩kL����n�I�"h��voo�Ĺ�U���y�^���>�(R������s��l��m�kJ���ϕ$���P��9Q��3������џ~K���(V����o��N��L��x�U�k'�,ז��ߩmLJ�͡~d�)o�d����@�dOO���k]mS	ǵa���4�9�&�/M�U⃴����وn���������ٍѮ����z�'��7�U/��J�$�g� ���ha�����^g�J��X���d(��ﻺ�lҾ�w�Y~`ɻ���W��N�E[U)zƏ1�������,�=?�ە��ҝ�+�hH�L��C���ġR����a��_܀)�-�U�FoG�D_��K��\<������z`����XD�-C�Q44S�}{�G�RX�i�\ų������$��V��+� ���]�*<z�߂����=�ɼ&�7��}���o��5W���\��P��n4�,�n���MM�i�rU�{��4|�7�Ұ
��ٯ)������i�w]�/��t��-@>��ݷv�-��ZϽmT��.�m(���#��d�$�q�bn�K�_�L�ޡ|�I(
�i�B��9H��o�a�L:kf�q+;Ů�ǭRC������?��+�����6�����+���U�4��+Zk��z��J�Y����.��gRx?�C.B��r̷� +�T�T�(2��Ш�	��|p�S5q�5v=�y\5T��i8�������c]t����?�7P\+��`�CXsk��ݩk��y�d¸1rt}ҥ�U��=�^E��-�㦏�% "/*b�iT��*��f��^�mR�|"IaM�/3P����^��[���5�Xҷr��Qh�R�7��*����%��gE"�����?����}���θ�ꝫ��V&�T$�@�ن�jɳ
j7X�G��v������T��{�W���1��$x���^�2�hꮪ�`w�q+���ܧ�pT�b�	+�����{1��|Ie}�:��f�u�F��j�"�q���V9pNY��,Xf��6q��^�k������L��#Į�CM#\�bU�۪��x1q*��SxS��ЏxC.&sU������獮*�����IAf[^%��e�^�~�c_'����:^��hDK4�Ƞ���������8qh!���*��^��?�9[�2i��׽WCU�� ���EP���+�@'}ъ�\�{pQ��O�í	zc�|������P��mܢG�2Wt�k���7̛?�p������L��0��Mڴ_�C��8�d���F��"��O9lҀ���߆��.�M�x����}���?"�u��TȾ{.�m��Zt�vx;薡�����cأ�ͣ+�;2�U�8��([k����^��s{�I�7��r�W�0�dL<�W��Ֆ��,$�0�*�67*s�親P��gf�>��.�B�Sm�	�V�)2I%yCCT���݅�a)��3fh�:F�:ko/4���	�l[��ng�#Q�ym8ԯmR��_ނ��t<s�'�<��v�i�����[����=�f��}��������P��]�21k1�=�_��g<�~ea�w�;L��jfqR�>a(7-kM~,�V��!4�<�i��7m��6y��h|�"�}k�g��(�����Z�n>�ά�	��S3�9x|�U��fǄ���E��N�2O�g��G~?��&5�>O◾�4�;�k{���EL�֩O��G|B�`�D��c$�����S��H�w��7�:tP�#���d������I��R��@)�d��{�u�eމ�d�5��)T����6HFY'9Pe��«7�3ӖG����6�o�����A�k+T^����p3%DP�y��֗�*�����W�M���^RD�J�Ο;�h�a�H��e��OTm�#p?ܽUWt%>h��L�]��j>p*��2�K��>ɞi�h),N]�oYU�/���[i���2�ʺ<�Ɵ��z�ܚ�]12l�&�Ysq2�2��_�YGy�~�S�~�z`��R�v�r�q^��2 ���_�5}�?n-4�qފ��z1x�c�0 ���f�4��RП4�"IoWϗ~}m�5�E��r���A��byh�$L�|��/N�h�vM�N��R�tP	(�I ��5�y��:��eR��R>pq�͂�d��0�N�?��kv� �	��;YU U��y��14�l���Y�V�#�/dY_E���!Y��K@	6���~�������\f/k�$៭��*�@��/R9/��=�Cj���&�=��зV��n�>���-�T\˵�_f�X6�"����BY�\�'睺��[�j�!-��5���%k$������1��2���aJ�¹F$9�t�W���H�M�t��@��'V���W�	W�!я7��fO3O�.��\9	c]�t�Ӽ]�.�ܘ�=�R\7~�d8��q�Ĉ��.�'qw�5H,R��:r;7�?~8�4m�!F��Χ˯t��H������,��&Q}�6��N�&���-���d�4M���`	5�N��>0�t��J�*����j���%��)C���G;qa@,^�]�)�;;�`R�ĩc�7�a�F�'G��Y����DF1|)�G�:������c��W�߯�/�"r�/��*�l�6aE�+��kx��ˤHƞ�cq�DI�p���#38.��6��7��D�gD�?ݣhk	��dH�Ժ���y*Z�������_��H�f�9�~��*��L^j�ŪN��d���4ow�UB�pM��B��=UU�bF0����qn2�f��`]ElǍ��k�>_�����L���C/���z�2%��4芷]�%������N!��>)65>Z�S�t��d�k��e����U����4��h�c]{��w~a�o�짪�9V�J#�OW�٭���$��Qϰ�<�J,|;�r����E�,ΏK����h�*ڐ<�A���κvCb�����A���i�:T�zEa�[w\@cM��p�;w*��ƭE?�>Źh@����'�����W4�5�k{�J�c}�H�ãY=��t�Q��?��i� >K�o쫜3-���^�G�9�B^�~TQ|oK+~�'//�K&k�|�?��e��T��:Zдڞk�āV��?p\]�y�V=fhK�?�8ݒ탪���(�䳛Z\����Cq[*U�u;[Vps����l��H�,8ߪk,C�P)O̙2_w��c�Ar�hbLu5����=��F\��:�����Ñz�R��ȋʬ���q�]A�$a��m�F�]?�-�(�j	�Z�Ś���)�&�u_��듍�K���J��ˀM�����!�Y��Ӧ������\�P'~����A��Q^�;"��n������|���o�V��)|사(k_�Tݤ��![Ye�"�X����[�e%u8LÜH�9�n篃���=74~��!�Z��Ӫ*��b���՛���)t8"�P�+���f_Iʚ/���s߈�ui��@���p'�y$wGyK=���e?/!:۲7�7�p%�
oa��{��Ч�E`�h`pǨ���8P��*ځ�g�.7R&3�I[��8���<k@��ǂ������7
�&��X�4)��9�u]D)o����9�O�K�.`�~�$`�f����һ�L6i�[k��A:�K�1�J�-]�[�Z�}�1��.�(N�@e���t�_�#�؍?��M'���h�K׻��j�~Ue��}��ZU�I��ʃ�갎rTR�K��/��2B�_!�dg_�Ry����W3�����g���K��Ίet���Ȧ|�ί�>�a{2H����J���ze�r��ӕP�%���eB��:(���ر�����h�s�����G���Н��D�+�W(AC���+����E��h�Q�rK�W���D���or��fdN����xã�#���?y����/�/[��b�/bo�)Z燕1/r�dv���r��~�D�(�<_�p�v���)�ʢ�7��6��2L�QB�8n�w}��l�Lc�F9t Үb��Dns�F39�eK�ln�'Կ*�Ƙ
�]~�a�1f0?��H ~=��ӢM�PҚ
|*k�G�+������$�K�BiۦY�:t��fʧ��CW�۟�E�nН��%�Dm0��]����EKU��޶�#����8�;�Ħ���*����(~��V��\+�EV%,*�S���[��vqi��n�K���'H�$�����&����]TɶK�@�����/��[��O<i� fP�2a��w~��l�̸?�����)[��/�2���*`��|�����ņ���j_���B�t$��
�|`qV�Ͳ�+9�js��괤c��0\tr�[ڞ?�C�LށaP��%=���ї���Ȍ�R���c{�p�Vj�RVۧ9MhV(��YU��x`�4C�zF�-�h1'�pU�=�BI�V��O��B�G��t��� ��+���g�4��*L��ǔ/,���ՒX�\�p�&�*�[���U�fd}��*|��܊\3��jPYE����/�����|���$��j�_��e��u5���w�G���,�R���nyR3�P���Y��NÚ�kK�b

_�lM��p[��{,���ףz.��y`˜��n]E����H�����:��<�mDAm��������MڜԌv�<���ǐ�k<Ԙ�.��ӥ��p��	e�7bE�b;�p����a�8{*�@ �o�3�;�n1�fTUJ��B7��
�w�mv�d5�n�}"e-u��>��2)\��A��1�v?a]8�j>~���+�����ξL~y��
�,A��&~ee��V>��i.�����U��bǁR�z��������z�ID�uÚCƽ������e���m�hq܊�wjN%S�e���=����oW�	�}��
�)�C5n�?辰��Ka����Y{mWly[����;n�+��B	���s�!� ���������|��뜽-����w%�Nު|L�I�F�^�,jqg�3�.HC�n�c���y�g�B]��=iKW"V�Nz��F��ѥ���,?Y��%�Os�,,_�u�I&�H��]H�s�������d+��n�����U���':����|@���O��&��J�\���բ%�<�Ŷ�6,���h"7��]���m��n'z����� C�u�*y��R�V0�uܷ�ҭT�a+ʯ�/�u��x�W�y���+[D������GƊ������|�Z�f���r�PطU�w��m�8�v��R�C�����,Œ��de��Yү�q�0a���:��y����)G-3Kp�]k��,0j�}�"��Պ�Q�6T/+�՚\�KwX~���qE2Ѡ|��r��a"��6�@y�� �m�OƯ��Q���
!���(�[�4鏋"�[����5:"v�bA���^R�⭢5��`�Y"݊.��F���q���ZX���UX4�46)�]�[̓���>U~2�%SRb�F�����Yԏ΃�8��/aGMm���$����:ړ��9�Ǉ����r�2��&z}�ލc�]Z����J�~��G���x���_�6��[sC��/�9��D�6�א.�xc�m��p]�X��4��]�g��t�h��YJ�x[9�_��S�k�߃\��򯋶nt_��N����G��*���w��
�+����[��'�p�ʹ�Xv�uaQ���Z���ֵ��Y�2~X�G�T�4G�<x?I#��r���"8�[GG�lt1�(����z�_�X����������}�|FV/�V#�	�ޟU�@f��˽�o�Ow��N>��]e�S���])��Ť����7C���J��r#�"�ɵP�׫,���R�"p@�_z;Z�<-�['QՖ������0��9Y��V�֓!y���y
����Se���/��.P�k�]4�<n=O�f&�o����hý��\veֆ���VHUx�!��5��G���Ϧ�q�`Yt��$H�\�Np��u����=.d��_6����w���xk���vCB!�A���y#Ty��]D%�ԽNG+��fg����)y2����Aez���<d]UF�xwE���9�n�g�2���z�u�S�R�z:�K룺X��������4�C�Է��G^��^� A��o"��L�Si�U�K�\y�3r㪮�Z��5Dٚ��Y���#U	F��`��\����2�&NR@�"}?�
۫��������v�Z�Yʘ�V3w.�]���`�����򷓠l2P���"-
�����7�U����6���c[|w�N��*h�uϟ�ԙ�=>������l�NC��m��uH
�62=�,H}���N�����3�s4k�ͬDA����}�r-��j�����0$h�b�ٔ�$0:R���J�B]����ds<U3-��iU� b>��]��=��J�k���:�~d�1�7���z�95ZŒ�w�H��'�J��T�����s�[��R�
��!��$��3ή> �Z�nVI��^1��6���k�C��Jb��M����'mW��.�@�Ҫ딬ȵnj�n&����ڠ�����m�y��8Rںn���*��+-o��pw����!�^~q��<��pAj7�h�J��uG���D�`�d��O.�����
y��'��=��z�����
kl&�i	���TIU�M�?������볾����Y����VY����Z�l�N�+�œ~��������w����6V��K���!@��
�Z���/��nR:?~�����6���!��ah��͑�#mkg�Ǎs��)�h���z��Y/U������f��E��eU�^�u��/�y��-g֙�M�<>� T*�����	���.G4ۡ�	O�}�3��%>�P��T�,��L������!��ѥ�^�l�~��D�<�j�����7×
�<������@?������&(mj�-sWx��E�{K�wD�yճjvϩ�~�=����ё�΋��.xZzMC�Y���,�"��N7��D��J��YF���o:U�0}�����ʪ&��H�h���l_��0�=�H�Z�ă/����f�Z5t^�D0l��ȜDd�R�?����a���|�b����%�����p����Y�h.����m�.5:�ﴨM�Ju��^5�G^�D��l�Y��43܌���Q�\_%U�W� �ٿ���H#�����ʁ�m.� P�y`��E�i��a w�2g��fap���i֯���\�\���W�5b�������������V��Ś_�s!���~�X�N�B����4IP���l�lUu�5���8j�J�3i��Z���E�>�6���(��Ki�iK�p9y�@��X�|OsW~���IS�����%��*I���	�ԏ�}Hɓ*�NJ����q�~��F�bD�b��>�ߋgu)kg���-�֚\�����ңk���i~je5�qy<��0��5�Ѱ^{���8��\c\UF'�^�m��"	`�i��&5�V@�� |�A��G�w���b�Mh�+�bַI"������9'c���WV���+Hvʃ��X�1�K���i�}�3���;̶��=3�������n�kp2dn��肶cF���I�����"�^�V���ʻۊ�F+��~B s�,6�X�z��N����������>�R͉n�d����'(�?j��(�۟��"�5����,�7#]�����w�^��X�����7ciN��\S�d��2�S�x�lK�|e�f���2ya��f�E����>���Aږ⭯{���Vu�%Qp)�۪���H�Vb1�����3���G�}�=曳c�1���2�x���Ո���d}�k?/-~.�����������`�o��	����D��	��~W��H���9��*'�v=���[3��8��p��V�+�T�۟+J=�I$��o�ԍ�Ȫ�}���Ee˲q�^��0tV6����f���:M'Z��u�G�}ꌌW"�ГH�=�1-��C�w~�;��oz�q���*��w��0��T�zs#�h8W����`p��DP,�cU�7�9<������Ƣ�>����>�2'�Q���-M�D�r.�~���-��)Z�'�u���jQf�=���K8⇵�U���q�{l�.���Ճ�UR�-G��X~5(�����h��3b��*�g1�\МЯ^����A{�4�^���
۽)��|Q�����K.M��ϡ�W�m����3���'�)��#�ꥥ�DkޔAҶ�m�F2���կ��8\�֝q����u��=�Cjԁ�u����zScֲ�ˉq��3J�ݢ�����Ͱ��E;��7����f�?�\�!����{�1D�'�_���焅�_$�%%=�& ����*��r�[�7�Zb�$F��YWO��p������ʇ*��{ޔ�Om�K����3�������t��[��]�]ԫ�t�А]�FzR���yz[������.!�YU��?�L���TKv���rOh�N������xCrXD��:[U�e&��7Z���WG9?�wمM>� Ƒ�Ɩq8�J�H�E.��޼c��� +5K�gH��=�2W�}V���YWvr��~����dt�6���N[��V�&��o8ʎ�F륧'��C/ W�W!��h��8��lMѣdǠ�!6b=�|%(���Z���M�V)��g0�Zֱ�F���q�G�F��Tǎby`��܋�{�P�ϐG��o�o�jm̶&\lS���x�X��k�;䈃���&�
m��+5�;��aH1�ݨrcH׭ihӘ�:w�������>h��О&R,V `�R�����\��#=M��F���d]�Re��بʔ��~�׊����J,c���K�B��_]c厊�2!t7���W����2q�q�~��[�����\��� �P�cV %��H�i�'�muý��GQ_�
�˽)�{?6���yO��9�����%_�EYk���>+�_ �87�)ߑ�`�f��8��+���J�5�m���>�[$N��]��g�1�/�+�]K�'�;���?�.;׸G���=_Wj�������5r*\z͠�����\ʠcͪ�WT8\��(�\�����@�������>��I�¶�D��{��^F �K�RѼ^�|E�iTfSp����%&Υ;�ְ�������2���=�	�:穎�dU�YYy��zV8�b���W��'����*���tA��tG���dݺpta��K`�\{�95���_k�*���G�.�lf��&X�o�F�rT���bEg53��'���1T~��M]����:i�UM5c�)�Qi���?ѫ�������վ��!R�T��k��5x`X o"	x�ݍ�[�e���s�os�AK�L��5�x+gH*/)]61���`b>��Ϻ����?�7�U6ϔ�6y*�'h�<�uU�&'��q~�3.Y��22�<��G��S¼+Ê�����՗�j,m��؁�z3Y��LW�����lI~��x����S�o������|I�{���q�����s�����6\�k��T����sa��
��s�����I��/�T���)"H�U���0��Xפ�_�v݊�w�V�3�w�Ĭ'_�m����k�\�׸�q���01��HG�r�\b}�"T��LK/���e�k�����u5#⍑S�)���=1���T���l99�6����/K����|��������7.�%�AEJ��w�=���v=O�g]a�l�?7k�vC*��/w�DY�Δ]�+^�U��GI>wrGR��s��D��)�0>�������f��G8,��B�C��@��mq��4��/rv|�L7.�7Tvs�FǖB����J;�K"�ʲjt�6t���{�c;�+c>��x�hG	�%=i`�^�/��8��3��r��)�;ռrB���+zajX2M�Sq�$�p�꺵J�.�_S����6�f~̒�Fۄ]��mW�C�m
�d��b_��͛}U�Ps4�eı?��X3<��ҎR���{	D��by8Wj�&��R��t�E��N����y���D{d����_������vYH=�GS�V�O��d�A?_Z�/G�̶��ރ,��tTJ���w>�^��3
.��Fs���{l�31������g И82�#��۟]�RR3�Z\�yӎ��Vމ�����ᤲ��'��V���-�h\�\eB詢��i��wb��ݝ&��L�]�8�]�a�k*��*���XҔK���f��AA�G�K�g2R<W�,�&q��v�-#��J�a�_�>Ż���ݑ���w~�Ɛ~��
wR�[�N|V�$����&��x`�V��(ՔP|�	��劷�0�������µ�E�v��p{�ͥ�ʞ�����O�r�X.�D�BZ����m�C�S�(�Kt
�'��)������l.￦���c_��L��Δ-Y�O"r��̑�*�t��]����F�o�Y�
�³>��wn�@�ҏ�V}�>�K�q,I)�������R������� �㍚�i-f|nRN|��68�M8
������z���pμG�[���ݩ�/3�\�큣�Y�N�[s�e���:�!m����Q�ށ���n���JN2�Q�]�Ly.
��p_L��?-�|:���%
�ή���4��j�M�/m˱�S�@j�r��fb˚���J�N�K}�M=n��$�Qt��;U86�C���{,�j.L:Z�R�s{36Q�����*�\C)<�4/��b��8Co-Kv��M�
�/��]�}�����>>pɇ�F���/�0�������%�>������N��<~x��\\��	)��.���$����!��a���uD�u���f�b�Ih:5o�q�<�����O?��/q\g�K�V�%9�)�Ō�U�#�U����8��n��,K\Xֶr〪h��V*.QiU~�[��夝��+h���r�˖��Ҹ�9?�5&��%������=xʆ�
��k��>As���+qP袖���?�g���B��TG��U��_�[Q��ܟ���ruA5�~���
s���տ�������K$��aG�`�Av�7�-#ʇV�V��7;+ ����pE�+LqYǪ��~N��7�0���k�x�/����Dc c�?� ����ǒ�zצ�i"Zpq�أ������@O�T^ɓ7��e���]@�[>�����t�%(d�e�t����ɇ0�e�?S.�\��7���Ÿ�l�{�)�gn�ϸ��5h�$P�&ՀE'*0�M�P�}�>���Ѕ��T�$�-Ɂ��M͌����c�cV휺x�ؕJ(����}�=a�n^�Hb'f���Dg�
AGUM��+��"��):�q�N�nW�|h9�/�3[��|���c+��2q[�F�2��}H*.�>r?�t��v�˯�擮n�]�|`�(�D~j��W��j-���Dj���K�d���F(�!����c0��>0�q�)%f�}���Ɲ=?o�,f�K��U|���8C|r��Q�k���u	�<Q�.�4�<�YX��-��5�)��z��0r�j��_*��}$iq[���s��%�P|�s�S_�~������K���w�t���\��u���/Re�za����$��R�_��O��W�0��֔�KTD
�P~E��<�bץ�}}�JT�8���#�VV�Q�s�ز��h��K<PA��5BX���ay�X�H�[H�P;vE�^B�a��(���RJ_0��"5�_)�cx�՗��y�:ʙ��	Qam�:7L�X>W�J�N*�s��6��`j/U�cB�]� Z-eW��}�Ĭ����z͙~h�(�&3��kg�+�%};��h71m�{�Ōݓ�>��N	vW�/J��h���_��$�r�����t��e�W��;Z��sB��� 疖�sNL5�����Ը-���" �M�Q�#�U�o7t����]�qb8kQX� 8_�/���Pm;��q�J ����d�5SR׳�D?5��=C�;�ܣ-�Ɣ�)�C���PY~b+z�Dwy���)s�!���u�O�Ltl�U#���0q�RGm\<�w;	��9[�W�B58��2�]��[�Y��Jh̍T�n=�ǋ�Xd�sS�r܀��1�g� u�.�\���5�q�?싆�r� ���ǩ�����Q�:{:uy8����t��'>GJ�K��%�Kx���V�T�b���m͡\=���J��0ZE��لm��ZR��;�-�
������P��J���3��/���V���{Ȧ�S�-e��%��^B�����>E�+$
� �,�vR�JFVCe��(��I�������Vڝ�K��V��k��W�3?⻁rc�N��<SV��_����M�"���=k����h��\��x���WiM>����?�CE�������P�����y9}����v��>�>��J"�p��D�[�7;��{�&s��U��j�r����9��P�Ǉ�.�&w0��x����4�xJ��;�/n;���T��*�^;$�4������ƃ�u�Pl2'�~:��[�Fs�A���[��Z�������x����O�A���+v.��$�:Z_���/�@Ox[^��� R�X�k0c^yx����H��s%x#�=��m2�@��}�g9�+��܃�g�̫����ӑ�𪪎]Rl�or��.��=�����Zpl�Xrb��#w�dI�\d,�&7�Ψ�"�V��[Ҝ*"MU���R���K~��".SrU��'�rh��)��}��֦���u��c��P/-T�x�v~�X���!d)C����?�����kĚ֦�J?�	;�b�0c��?�O䏖�8�
#�4Z*�� +o��DK��-���6[�q�^bP�J��2!Lc��V�s�Mjs����Ǔ#��g��c�>S2�,U~�c��}��r��OAz�R���#c�y9�:)V���V���/~��Ni�X}F)���
�%}pR���pSքT(`~��U��ED��~�>`�J�l�R��}�'�kA��*[��gJ�xV�Z�,�$�c�i��A�����,3N�e9���UEKz�i��*}� _G.��P�K�9�9M���B--��@t9��3����LK�Q��;�_۸��/x�cT�(�	ڥ����O�U�H�[� �/����"�� �<��9L��}���8��S�V�).�h���j;UZ���1Q��D<x�Ϛ���W�(�!�>�����p�/��̣�)S/f~*���%���١3	�����rVFȎ:k6�Fh3�w*M��̈́�d�������,��]�<ɘ*�*�������7&}��T)�h�_AY6�!+�:�dN�ϱ�8��S�~���Tf5!v�ݩ����{�EkZX�[O0 6%�49�|���0����I)��˓:U��[wo^�<;,��ъ$a�	Ē�4)����Kg�ơV����hX�d#�E�J�s�e�4Ő�/狀���.6D����u�V��Dw�N�O��I�	jw���r-ͯ�=��û�ʉW��|��JG��!-��<f/ˎ�����fy̓�0!k�o?�_Y�W��?���r���_�s��T�����Df#a
?_��-%�xX�@L��9 ��4tD�?dx���n-�T;�t��,��zY[qQD�?4�&3�V���iP�:��,�U�R,�C�˅�_zcf��\��ȵ�
�Q����}%D��eXǦ6�J�sO�8wX#L����_*������s�0euM穻жo\��E�BW���wҐM���M��ڜ��ݽӎ�`�P�ms5P�ǺqN��m+���[�i�-2���
	��kJxiO����$�7+u��3o�����J,���0����s�Tg�2�����Up�+��g���n*YJ��jW��N~l�qn<�?�B��&�q�F��ڥa�'��qf�2����<d��Z���6]3��T�*�[��0R~�BO��%ս�̗��0A��x����[����E8��
��4l��`�;����)���)�\��W��+�Y��*k����:v�Q���8:�{Q�u�śB-�=�_i�e^\	�ϔn��91EH���M�?B���c��v�nbe8��=�^���N(Q=&�L���E�3�2�������S����������t�t��O��y/ً\P��/��i���QrP�R��s����~�KL���n�]/Y���g��R�N����g0��S]^x�q6��Tտ�/�h�'p��� ߚ>lZ�H����ɓ�r)�Tm��6x�r�ꛓ۳쇈qa�:�4j�:��E���$�t��_�5�U��%7ԉ�K�)�>����*ˆ̦I�ǷO�^q�Q�Rˤ�������PqgV]\O�0�V�����7z����ƃ��`���C�Y�"m����zSڴ�.�v�K���*��l�^��JdXJl�Vz�����bY�:+����ּ�_����K~��-=�U��qߵ嚫k�+�6��D���;'c&E��و������w�����.����G��:[��[�fgc��^鉌3�y��><xŞ���xGB��7�p�"�R����#[�KR�m&�8uR՘!�d���~PL=J�~����^|a ���n�T�-��¼�?ϩ���xl�>6?��I&�Pt�����1��/T"O@��O�?l���h���b:��ԙ�Xw��$:�'�}����,i�߻�)�|��i^,~X�BW�Lrqs1#�Zl牐�����F�T��9�ё3���F����c牊��:�Ƚ�e�T}RZ��qh󺓚� ����i]س���ʁ�_]��^7^�p2U���W�t�e3ݵʽ׍�YY�uo��,�.�����˯�l/ջ�Tx�C��5�Y��yͼ�9|۞�3P'��.j�85Gy�⯺��h���O�'a��iҢo�ft��p���ǯ^Uٔ�T�i����ќ��qsqُK�&��߹5Kƞ��֥�U��--T:��>�~�+�R�5{Xæw�}�X;.Z����g��w����)\�jR��,UK(�h��@է���V�p�{e�W��n?K��/��[�}0_�0�E+��D<\"~�57B8嬟���a|���*�ODh���:}��[�F?��Z��0��x���1��S=���#Rp�����|�:ɵ��\;�U���L3��.0-�x%y`G����R����KD�����L���(���ߛ��M�En�ɠ��"��n����@�1��4����_I�kl$/𥊗�@}j���b�S�U\�X� �ݴ�WJ^��\6:d��ɩ{1��mJ��g�{�ݕi��E�;5K��J���Y��=���^�-j����eD�{�n�K�6j��,���^"VE���#5���"fYW��W�	�?�?�7yG}cFK��"�h~���=r�-M�X�+���8p�����$���jHV^�h�/t�'�����Ό���1��8C%7wF���Cvtu(ȷ����;�;U�*��Ofv�X���q��5X~xu5x��M{~>T�"������Z�b���j�%#)G�a�V:�q|��)L�
i�h���}��ې9x1�E�,�_�Y��>�>�t\wI�_�t�F��#����g���Vh�Fm1/��w�E^犯�7�����8�Q+�֯��������$@�fg��*��I�`r����F��؀��;��u�g�3��x��h�܅�t��U�A��v�z��n^��LW|�3�YS�?7:�m�i]�9�#%�<�k��:���ٲ�}��O�j���,Ȃ�x��/��F�mMZ�4Zͮ���.mI�<���w*Ӓ��&L��,�%m�׆���0��Fyj����_���.���l���F�S��T��kN�D$UR�`ꟼ�����ѭ�
,�Q]�ӎ�3Tp�s�BH�yo7&9�e�k�
�z�]�嵰9�dU���f��0s4M��uN���O����t����/|��::��鏍$?�gٜ���M���G]p+��tM�PƅU�V���
f(���>��@��#�S@	(B� F��U?E��B%�>L��b<F|¹'��2�a�``���za`�#����`T ˟�R� ������S0�``X��0j���	��xe
�"�	8f4��?����'��x^�"بĨ1�@�f�{�o�;���
|̛p!]|P�{�	�/��c̹��8u4Q�d�QM���,C���|�7U�k t,���G)ݗ�Va.Y���)⇗6Z����wE:�lꊻ=�+�7WIU�ҿ?T�^�内��n�e��Oq��DN���h�C��w��`E�O�Xߨ��?(�u����Y1�����3��/�`o����-��|UU+��VyF��e�h�P�9f7���5��y�?D}�Ɗŷ&bX�^�+t��p�?.?.��Ҡ�,�P���9SJ���q���O丼�e��U��iY�i?Һ<u��
�5�ºZ�A�T�+~��[�Éi��w"��=�˖U>��$	�L����-�y����k���ꥢ�̭-"�/tUe��̣6���롮�]��P��.
d����u��cW�m�N�PG�����8���K��E�h����+ZF%��U��_ф�я��=܂�>��hޕf�}��:�c3�g��W�%v��h.z���xB�v�\B@I�mN��F��#�?B���ȥ�z���Ώ�����|��ԅ*%�K����c�?8cc��g)��Y� �%�q�XUY�R����efh�c֭�Dޭ��<���3�V�|>i�P�u+�\޵?��*�����A�C�WG��F1G���� v�l����}W%�¥T�\��GM<D�$�����m������[�^��H��34ůN�i6���\�V�,��\���]Z�卮z=+���Ik�ϨZ �٫��e�p�bҫ�>gC�F���&*g�Oy�*�vN��z��f�յ��-�ژ
f^��K��ޞ���Z!Zӟ��;�,�ۿ$����)��So�p��z0���6VO���waɠ�-Qຊ� �I{���F/������îgT�ԙ�6�()���~C3b��7?�Ä=����LM<ʗ{��G�����d��f�p�th7~?}��i[Ƭ���f�gd���N�Xx�ɰ���E��#"$;8��^�u.�<�.�aA��������\�͙9��2V7w�\8�u�}�/D[����A��� (�bjɪ�1P�3gz�Ў��c#�q͕������]�MD���}�W�߈��$���b��=�x`����cE䣉4ʼ��j�~��;��(����-q��HNԺ�� �H2���,H}����������W�&L�"�*0b��*h#'#�D��2!_I�ڑ�YuG")C~`���A ���g�·Y��P�틮|�����a�b�-:ϿQi*�~4�כ'Y�|Fq%���n0_Ύ��:�J�
u�H��e����sM�Jz�1K�Y�ve=dI��Wg�6��j�,�g�C1�@�%ɑ[e<�<�}y��|㑢M��:�}`�/%/�
�ZEXꆺ+�*t� #w��	���^�1ev#���2��ӆ�֤Nب�RE�k���Z��9��_�T%�2��5/<[R��,bH��i?.]Ȏ[#4J5p�mS�V�M�+}�vt��礍�ҳ)��W�Ru֯y-�ט���4�Ե�����8u/đ���>�#-�����4:�	�T/��Btҵ��2�s��_�ơN�ԅ��J����֥�'����C̡��ݱ����@���E�?�%Z � �g�g}�9�z�>��q<lS$����;B����B����W���\i,iZ����]Lh��-\~�m}Uo/_1[�����'���,W3��]�C�Ӛ�ӹgy����u�Y	�xE;u �H�����_ ��C�1��������>}'�� ��Q��<C<�z)<�o�}�}|=�$�v��(d-?W.ǆ���U�^&V��D�?�ί8]7�WM�C�^\+6<{��r�nd6���.�����Ii�`���$�M�"��}D@?���{�a;Â)^"��X@/W�u�bIF��4Ps']�d��y�ע�#�e�+��=�h���b��h�05z�eq������� �c�iy�h�m�D�z�F�1�x�M_����� :�%+-B��_�p2�(n=s��
�����&�M�J!̺�wQ�/+S�*tHc�-Y4Z�bt�E���X��R�����9���*�ge�"mi���a��k�H�E��B���dtA ���qh	Ҙ�0��;�u%t���?����Q���v�O�?�r`�rֳ�D����ϫ�)�WA�۾X+Ĝ�&NTg_n�,��p�����o
M\��E�|��Wj��W��Ԡ��IΜ���P���Mzث8�un�����(L�Wu�Gd��@��)���O���Կ��iU�,5�&��v�c3��=cΝފC�ƄR�-��n�����ܠ����JE+��ۯ'l>�N%/�M:"b5�r5g_�r�p���>��̙��C6#��	�(X�j^_B~B��<��+d��	'h
�`�)�0�� v�fՇ�OзUl�w�M�E�_�V�e�N�/5����c�e�W�8z���u��u�n��M��0z�md���eT�d��pl����G+�D���,�}����X���v���7n7{E:�nn�G�,�k�$�BZ��cD�Vo���;�"~�Q��;U�t�T|�:�����h�/��9��e͊�E���u�P/����s\i8������zl�*�k����=0'�&�3��+�eU�b�}�$��[bT���|��,i�1�H+>����X�b"@VtDu��Վa5^��њ���#+I8��=��(ْ����Iol��v˩�\�ӥ����F��7vn��J����C�[nT��)�Gs�SM^YGW�l��F��9�e7�y�BB�Y*�|��j��0R�h�~蘪t'Kv*?�ou��ß���z�%�L����S.�w��<V�-�	�.کx��\�%M/���Q��g���Kk.=cB����~����z1k�@��3�P?.��x#[EqWD��ګjJ�p�/F�o�J�s��,.����3^Bi�^c��R�A���g}� �q��}�_�1I��q�w�%�i�fjA�ST:>�=|�(ș$����$��i���}���UA�%^���`%�r�1�~_�}<��,S~r����^�¿��ųJ�Y�/�h����n��6�<7�W5�b=�#�<
X����:'�G�.�K��Ц2�=w�s9���1� Z��_�T��R��'c��_�OREr=lyA�FqewW�J�!_q��������-�Lx��ޛ8(t�Q�_��^�U�wѼ�Xm���s_1�xoY4�~t=~Y��zX���,��~�T��2K����k_��~=nե)��'���o��~A�������惬/v)��\��!�C)���$T�����2����� ��"Nۂ��?���z��&�~�F3X�v{�*1<p����<�@��228��B��ra�jd�HR�L�������ng���sz����%��|�룅�O?�5�f^4ذG����\Y�c����w�"l>����h3B��<�ǅ���1���mq��50y��+ɂJ����&D"N�h� ���k�Rٟѭo��ʊk"O���.N����C�m�[��w@��r�GN��P{wBu���/��<��j��f��z��dU�X��i��Y�1g���VQi��
�(���͠.>r�횀�ǐ>EJ�|�D�m,
z7�_�5��.�z{�1{�_Ŷ���'B8�~��"|��ѫX6�l�D�a��Ǻ�c����U~���H���*�g�W�m:|���ɜ�5N�ָ{�:����;��>p/���4���h�;N�rM�]~xv0�]q�:��"�X�^[��r%%�($�8b�rʗ;��IS��@0>�2[{��5��W�W�eRm�?�3g���:���Z^p�_)�O;�@K�K|�Z��)���}T�hSu�ޑ��8<8}K�N��0���`�����%�x�>�x��x��)�����!yd�F��������b������5��b�-�]���Y&�������3:�J՗TIUV����_ҳ%�ۻ�6�=���P��"�Nq��T���g,����~�>�.]�&$T����*]gp��Z�ϑ~*Ij��:�,)���g���. �Y}�I��
��|F���F�z��K��:HhǙ8k�y�e������JюH�����mT��/]^ϋ��`gr�����o��W>-��	��n��-D)�����۬ 7t�AQeX�T�ɩ�.�/����B�Õ��n�DX��3�s�UM1>��9�	�B�Pq��1w��Z��d)���k�y�ʕ�9�����ށͿ�/�m�󁢍�ZXu_w�M�}�M+N��i���7�4"��"�\kT�(H��tM��[�e���f�����TOҊ�i����i��~���y��Vt����3��.V9�ԕ{Z��B�>��j����Ȓi�be>[3���\�]�%��WQ\��~��'6[U�C���w��=7(�͏w,���J\��)6�J�#'�Z�{!��,�٧D1�V.�a(�ԯ�����TD��y9�*H/w�u-?�Y�M�����	u��z9�H�0͝.����*9^�ʌ�p�S���T��;o�h-���/�
�zn��[��'`����A���]���hW����s���n}�s�����d�,R���y�ۻ�4�ce�Ud��	{�'���s�~��L��j��H��d�F��tR[�L��!���U�b�oF�9��
���?j��y50&Y��E�����!��R�Sf�V����)S�E,B����l��XLe���z#3�n"����ˠ��Ί.I>6�⮘ɟ�%�����tf��z�yK3wNU�{jAo!sϧ�����(e9C�ʫ�#�C�?��q�5q*c���˺���8C����H���~�e��E�7V�]7���pmx��+��
�������G�_���ɯ�"_u9T���br��_ �	ⷞ��d��Xm��*ȼ)4�+���~o�{���F��!?�z�L�ðk3�O�,��8����@�uI�ySkM��/�����J���-}�F��m�a3�h��5L�vm2��&T�h�`�9閞�x���X�*�Uh7�������l_�=�U���%ܵr��jɗ��]�.��N�UG����#���&򮨆��Uv8J/��큿:fq:m���VU�x�$�m1��u�hP��m����U�~�v�~77c�/�ץ={k���j,�׋�^�0����)��r�t`DI��'�I��i�2�\�м��2A�Ll�1�iJv�����c.s���ɟ�����kK]�=Su���W8u|�4� ay�E��'SJ�w��n�����4a��F�8)��PE��,hҏ�sr��OR����њ�(	�/�!p	P�e�o�3�>I9uI�}�f3a�[��,��5M�S��%�x>����6�E'x��?a@®���_�%�J�qڽ�7�}zwg�����V�X/�Ŷd%��k��������ل3S��K��ň�"�����0V�<�->���pr��K6��yE��t����� 0 �H8\�� iq��5s�,�+��+�X�;r����}�=����n���ڧ\�"N�GŬ.�+#���`����.���ӒA��VAQ��w�&;f1��<��s͒s*��ݺA��b)R��		T���3����l#z
E:����jZSt�*��,i��E �U��b7V�D6���nT�D�UgYU̬��Rk�����W��S�/g�gO���t� &��������x�y �eQ�Y���
�<����\m4 ��XW�o�M��3Z�Z�1�8�����Sk��*��}~���U�:o�����X�!�V��b�3u�U�(Z���#f���m,+�!~m1V�ץ��LW4��O̔B���˳¹��)@�Z}a��]�+���ź�.L���VV`�	%u\Ǐ���U�����Kxwz�G�"���0�*�����HVЌ����2A�	������	%4S��TZ���ӔJ!ct�0��d6EC��vFJ��d�G��V�{�����3���W2^5�U��M��K�!�����Gy��������߄@� 5���/�:K����IR���+�-n�[�R��q���;�fKV���Ъ�L���Av�$2j�x��"c�Ǣ��ܖ$���_�V����^A����F��X,�����B�V�ũn�K��3�D;
Ⱦ�B:mTC�wC��=�I޼H�I�(K�տ7�L�c�z�[X��B�Y�kYV*YT7���<�lI�W��G�^N���"�MV?)�����m��Z9U�3\./CV����	9��������G��Mg��T�E[9X�]�2�T.I�"�/���`O���&�X����}���F9��*��a�VK������z�@�֘x]�E��u�l�!8��'���)F�_�P��Ui�&o�ֿ�Ü�����ct����v}��� �oǶj�T�.��a������~ӓ�څE[T������Hcv��"�:��jH�R%X|���b���X�h���3sgZ�E�B2�R����}�-Q؉�z�7e=)��	�BEcY���5?7��VvS.�(�L�B�؝��Z�����oD�A/���|�V��$JY�CiwP<������+����[��n�&S+�$�B���^m3E9�m�4O�ZBR�t���_i=� \��q�P���;\L�o�~�ÝR)Tx��bI�F�ڮv��S��1�����(�����!�o�,�������:谢)!V�Y���z
8R3��>�����Z-`�E��go����?̐���MpS�>�D�����,O��Lq�m�x\�E�<��~*���2����]d���}�|e7.5Hmr�G�ȥ�|���+l�4��<�ƨ�A\Y����/�muyy�Ēb�e"����0�	�x���ş*#̈������j��JL<B@���Ѹ�f�z61~8�����ۭ�Q����������>SwVtS�E����Bi�:���PQ;��]ڏÔ]=�穌�彣��;k)<<�'�gcՈ�qrC�#vAV+
�lE�J-E������ɟ"?�I���o�
���U(ޒr����Юx�����"&��D %X����) ڔ�Lɏ�96��O�%��e�o�T��y^my�������RY�p΀��b��Ւb�RY��%1�Ltt�|����t�0X1(_>sz;�{\�6���AU}p�}>�z��F�91�*h��@����?��-R�"~�O���_0�6�'�G`1�|��NW	�k2O�C�N��T�\)wg�kn���С̓~�S����)��ȝ�z:�=[��F��
�9G'�EZc��U��Q�]��iRv0��~YŎѧ[����N�,� �����_	EC!&�,��h��W��7�����}��Qߘ:�Y����{ק
�r�h*��PךӧG�*3۾�$he�|�Bڣ��0h(@�d��L�NY�|�.b�Tr|��=�Bѭ��}����WX�������x���v{C`� Z�>�c���/:���2�Q�D>�q�a�pg�*�^*��%���I�-��#��m��q�i�6wy�ᗱ�6y�dR��ݬ�2�Bbم^�J�U|�^� f�C����de���h�L�3/e�/hGE��5�?u{�{|��Q�l�����j[̰�z�[(��5�t�]I�Ǣ��,7�6.,(ݝ�??q�/Ĺ'8�m�/�/4V�)��~���0�?�li�,_�ef�tl�C&�5EnW"�%�p��:�L(�5���fvݮ��*�|�b�L��7;�e�q�x�>g��?��S�2�*�Wjk�ڇVԊݛ����}��
DK�5�t<uS�/\{�F�,X�s�n��x�<�4LeNrs_[�N��@����d�<���B�~a����D��_�1z��Z퉫Mj0��w�p��r�U!���t��e(��u*?�zZ���Q� �]-9>0=e��z��/�&}��,BY��-�e�`����8M�1���k�Y_�p���Nn�
�J��N�'�O,:�Tr�̏V*P]X��y:�xX����S�Wi��҆u�&B�/:aeɨAʷ(���Rg�Q;�>K+��f���T�g��I�4�����f=6ַ�����d:^�_\��)�_QL9t��
�QRߑT���IN�$0L&l?ʘ
�� g4�D��3M6M�RI
ߔ�麮C�OQ7ָX\�"�?�L����:�p���Uc��mn��@��Ւ�5� ]Sr�@v2k�X��n�F��iAf\ee
W���/���<ɟO���_�4ۮ��@yЫ�3��B1����|g�p9�����L4���T��?�][�΢�eOe�>P*�����x��u�e��-� �n�Rgm�gF1.q�'X�!�a��~�W����y+L����Vۮ��S8�r&��b�hU��/|�A�.D̾�jE�X*�=Zd�S�T��~g3*a�TxɁ
e����S��5N�u�J��b&�AلU/5��]�OIo0a4��I���؋)�P����N	�bʎg!&)��WDr��g�"����ﮂH��#��w�i��$
�)Z�(�lz����8��A����쿮3v��'[�|��z��Ί(W�Iǵ��U��n<ަ�c��0}z�-�p�NZwᣦ6�{Q�%N9' r�jT���֊n걬�9��S4�ƉܵR��Y�2��erSO��J�t"u��M��-渎�=�h#���:��*�Ϻ���ݶ�]a���$z�]�[�?�h��vO���pmA�JG�]T��%�f�܄_��k@���59�"s���L�27�vIq��>�����v�G�*�Y7QXRd��۩�B!]=�U��|��S&2Ow��d_?0�Q�o��-a�)��=Ϲboi����γ�̞�8�қ0ӝ�iU~p�@���0�Y5��C���X�y#�Dn�Q.�]l�/�����T?�բ��I�p����m�e��VR�u�#ٟ��>�ĥu5��y��Ol�o��ZΈ~O��oi&����xm��g�'%�B��ƠZ�L��~&*����<�`�������/��	�������A�)P�Q�u=ԥ�����/�������F
4�t�����K�[�W��I5�ᖪ��x���u`Q?�+��߻Z4��f�����yi�<R�Ѣ#�R�J�i�]�T���D"<}���KpF&6ܡNu�J�D��<pe�0��.�'2˓f�T��,/�v�h	������v�]����ni�������+Z���wE�ݏ�%�j������B�p^#}7��%��B��+*�����%$*��k6vPx�o�έ��$���Ie��Ŝ�hY��Ѿf�G�Ap�r�39�Kl���)�]�)����{KD�.����J�UM��_��>����1���2��,��txF�}��ԧ���~��
��l�{-ʽ�0Q�i?�Q��mj���҆�(f�:T���S��L�)�7�?�{#��R�םeE_{��q����y0���%y�J?9����M��1Y��2t��uP�6����P�C˰�/��fV�	׳�!�/�5Z��q�d�+喩��2}�u.����Ȕj�sL�0&d5��Һ�/�,����?ڟ��r�mf�'��:�2aɍ�S*�V�Q�>,��E^��Ӑ�F\�]����"*��P]E!��F+�V�Ls���iK�3>HbZ��ZUWy��?~�(�i������L(�X*
k
��K�{.j,�xq"ʵ��Њ||�+�h��&Z�^AJ����:d��˶4y��7�-�^�r�D�e�^�j:s��d�^A�0/�ꈿ_���gC�V�w��V�u��_+�߾�bЅw�W�y����/&���^��}K�w�&�#���N�*�bvpT{�f�+\�pv��_�N���KQ��v�Z��U'^~x�br}E�����ˁ���~�t'��,஽��������˒�U0H������j$軞:��:����$ʛ���<��I�
�0\6Bի�Cd�� W1\��Be9����E:�J:��+�.�l{Q��cJ�� ��/	~����j� �א�Ål��H�
HyXiV����O�mݸ��v�硾��K�:���5[W3}��nEɵ�ou�#�4��y���c���j��fR�g�����r`�$�c�u`�v�C�{2���\�iY��f�R�����w�X.蛁;�~"b��)?��OD��?�U�iֱ�UYy<暍�C��>�r��,u�9 �8Y�=ئ/0_��?n?Zu[��o�2�9}9�yR�u=�=J&Y��25����Lq�z}�_n��*�*�zO�dI���]h��e�zu��X�([Η�Ǧ��.������H�#�l�!;��ÌG"J;��z{X;h��
��;%��V�g�h�����)@���t�<zC�h�;wl�Ґ��1���m�q�����趎n�bN�h�=v[�FW�+�S��%%J�Lqj��<e,�JQ���~^){В^���r�_�Eml�/�\���R��+H|���7|c��\v������J�B�0GG4��J�v/���¿� q[�"AQ��єjCgԀ�l[yMM��!s��6��K�;�Jo*��L�WM#,�)�g>�ű~o�/Wb����ro�{5˃�VSØg#�"
�Fr������K��/�P�u~��c�m��YL���5�D}.����i���hm���a���s�}�}�h�vm�慮��
]$%�͔�Q�3Uadfwf�нS�E��gq�̚�h΁� j�H҅aZF����˄V/��o��� ʙkw�tF���R,L\/S��Ҙ�6�ְ\@i�ֽ���&2k���\�ǡێ�a��:�ߐ�~F��-?������/�a��û��$hZ�~�cDn�+��'(�lA��X�U�a�.�-�=�[G|�������"f�{�ߩ�H��@];<���-�۩��s��]�I�1��������%{���:O���� ��*R�J�%O����C͂�Z<�5j��T`�œ�'+�p ^��1qD�H����g�S���㏂6sf����(>��3~�X�b�bIC�b���h�?���Җb�r��:����Av�S�Z���u���EK����{+��/����5�5�S]ֹ�G�KkD>~ӡ�=J��Pb�ݍ��U����ʒ@�Jx�5��'����_͙+:�9b���%�fz8��N]�����pa�Y���4m�v�#a��/��J�J<޷b�h9�����w�_��EPxńD�:1V*몗&R�>��#"�y`iuEo�ߩ����W��j�<�|�E���=�hˏfJ����S�qaM�j*�q}��tTE&�-Sw�Ţ�����=��~!�E�)tD�e��u�6"^��5��r�?[��%IB�_��)3ի̏��Z���Z��"�k~��R��Y�@����ɦ�H5w���#�#�_��R���4n�Ia�"+�f�X݈F��r1ܫ(*Uar�U'�?�yw�ؐ��Q�e��N[����4��r��>-�����.��ЫG�6~��._6� �v8�X]��%5j�!-��o3-C��	nm��4~v��O}��cJ��>��p[�!x)��^ָl���~��ǔ�k��l�lW$��a�E�)#�ϗ�Fi��6_F U��e��msP�s���$����`�P;�����(H2�k�����4��k�{	%rE䬿ό�e���j�[��� �6�n{���wAC�^�)Qh��3��|_��Y)��bΟ�ԑSB��Z"�������K�����p�y��&��H]@���-�a��N�Ԃn�t��C��W	��y	�y���Z�;���_�-қ����v����)�>Zj���:��^��6�|-�z���%��T�T 8�:�@W��_���*i�sBȿr�d\�
 �ә�eӦ.y����ٞ��g~.0��J>F��A7˶�*)Z񐠧ΑC(3T�:+�����}Թ׸�tE��g>u ̃��?���MxBܶ�L&[��Y(�P�C�+A@�і*�#H��NJf/�0I��	Zf�˭�S�J��6۹�Aw딇��>r~�̪�M�hg�i�aѷ+�`�O��`-���_�����C���c���3�V�h�Jrr��pU�J�+��������D�E2�Θ�b8��se�KQ 	��'7Q1��:�+�����#J䎖��^�<pi�Ə����;o�&��z(f��۩	.�����ߟ��7m�	� :�W���fl)�}����� �����q&U�,�Ԯï*F���qڏ�lK�תS��p�6�Qj�*5E���L���Կ���BR��paƺ�O�W�SJ��i�{��)�t=e\Q,�r�1�U�*�\�9������tM,������ъ�#7���]]�	-$b�sW����"��+�y��g�fv���d����M	�Hw�|����,��t�wV6|v���ic[�TG=Ʊ�%]U�ߙ5�g��,�d��%���~��+�iW:��ù\5m�r�5���GE�I >�����M����C�f��D�0'�'�J^�}#�1�-��Nc��>������[�h�2_���2������ O�x��.��
*�z� ��x�!�u#RwJZ$,�(���"�eNў�����U�0\��TY�E��k)@C{&�_��20��t���Z��T�^�K�U��3���&w��4g�fq��A�֮:{v]b?�2p��,�Tֈ^ܬ���7"�О.���CL����lh��MNC�E.1|�����[�g�����01�<��d|�D����X�q�q¯R\���̐�!Сx��ϗ�(�ɘ�P$擕���x��U@�l��s��p��َ�/�edM���I�&m�l�r�E��(?�x�c�#(E���0}�_e�n#�����>sA�k�O�B�ح�����Q.���Ý^;�|%�oKO�fa���=��3Z	�`�M;��>gC��*���c�n\�݆�w�V�h�$�T��ў���@�5�k�eK�]S�v�K��=������n�O긯�u6�-�
h���W?2����)J�����yڱ�{�y��+�~_G��۔�����B��7kZ]K4{1z�9(+� ��m�L�Z9��O���V1|�=� ��c�g�~ҭ+Gq�T_�:~�8�Sƭ�H_��L��X�2�j2�)�W�����I5�$'����74˾-�ـ%ԜC촃����idVF1"iu~�J��_W�Y�|�1^��_�w��~hK_�$�.D����#��2��F���ʎ�F��sz>A ��*E� q��EYh�qb�PU��Wg�^D_X|f�t��<��~���gV��+�_+���U�2�X�(T$�1H�Q:��¢��vMA��0��;��|)}b�W(��ءしk�w`VѺ�Bz�q�	��e~��;�13�i�O�*�B)�_�x��,��t����sd~�s0_�b���}͠�ɕ�\���}M����m�����M���mŝ1��#wģ�����)�j����E�>&�H�����yD�2&J�Iƃ�'}�g�>Q�0��G֭�NEs��ؿ8<o�Q��Ԫ5�˴�C���*�{ܮ5/�ywi�P�A��0�Fۛ@������Z?^m��+-C�~݊��/	��Tf3�	�7�	�-UB�[���b_P��"�UE)yU%�����L�\Mevp�g�5U��aĕAs���{O��/�I?��}?�,�V��_����b���y�x�
*lG��Gh�v4�+�.fW:�_���9�"�_��x{�
�o�pN��Fub����i�ӯ��1�g?� �'g�]��Cz�?���B_���S9��I_ɘ�.�
�o���:������#K~��Kf52�k����^5��f'
E$��;��j�oV�3�/�e����D�����"�	�~(�ک���
�5�OF������G疬W��������!+�D_x��B$}��֚}����68�8�%}U`��1B�8d�A���f����z:<��uE��J�]A�RS���N��CѴ<BJ��d�c�K���{͕t7�YNW��?����Z�Aݛyf��T>8H
�b�ku.�Z)�p��l�T���^�sƳi��iܒXuł������I,ǩ�è��p�P�\��}b�jC������
O��f�eBċ��D��1�Ed�a�.W����NMr]X��U
�P�#���-,��
�)����U�ԅ�|rn�V��>.\�B��j,=cw����J'_(�^T@�v���������0����z�,���z^��̨Y-�U��	������=��2�/��؝��6k2�Jy�+��w�L�Q���w��.���§)/�yzw�$��9��~m�q,3.�����*3U���Žf����T�/�h3*!]�w���<����ۣ��؇�>��0�i�5��R�4.�ȏ6I2��n�����d���t8=�+arT�_f��-����U×��������.�i�VLs�6�8��.�+�_h������0J�~�>�h��?m�b��l?�d$��f5��ow�A1.�����4�k,�3soZu��ӿȂdA���P�&F�'j���K88XS~h?�����Q�n~�bõ�s�f��Ȳy,n���Id������b�ۢ����]�ӻ��5Z�#��JTu�b~(x�y���8��+�.��Q��C��������@�>�PP��8�[��o��=�<�[��b��"��c�hj�v��t������� �����f&������Iy3�۟5o�&�-��:Ω���PA���� :,u�Q�C�3G��6�~(�1���X�kc�0�����g�����W^�yN	��7���/v�MqdJ>��Ow�WN�6����/�R�8p�'��U�B��.��&@����s��2�ʥ�}�8���L�zs�����ir��Ep�ƨmB�7`����Ya��~)Y`�����fA�
��o7y�ӧ���Ȇ�Z��.S��L���Jͺ{R�ݞ1�ܔH�R�6�ՙa}�N��F�ԙ����cf���F��`~5E�y�S��B����V7T��7�˕`�U�j���U?�R�I��~���d����$��`ttß랸�P�Τ�m0ZHJ�R,d�?]�B�E����w���]2��Er�v���.�i��Qςr�{n_�Bul�-���糣�T������R���;�x��5��]�_�W͢@��?������Hb�wit"pU�k�uqӗ�Rnup��]2]�'˧(�e������x�rb��hg��'��w������R�b}�m�m&��U�j#�v7z?�U�Kh �T��ehu̜m���c���ֹ����c� bn��7���*g��6�E.1����$�(X��3�fo���n��i�}��ܡ<��4�bh��xd�u�]P����bi��}�B_	�Sz[�_i��e@���%�ӟ,��7YM�\~�&w�A�����ɐAJg\����+�����%;0&;��*����5�TN^�Q��[9�K��;�[��������e;�;vZ��(5�ʹFc���!>9g�4r�p����Qym�9���.�TJL��!��zs��@�!{�T'�?{��Ƣ$F%�����N�+�썬J27�������^�a�_���ŝ8�|�݇vs��|���x��c��27�u������/���[��_��s�Vu�p�/��!�ԢU�2}�U�&���2�>�h6\ʄK>�o`F��ƾ�.�N�����o�%E��V4/ǎ�.��xf���"������K6�(�hCHB�b,�T-��(_Dŀ��P@��fQ>�;ǯ��1߭�V�y�f,zZzVq��S.L��ki����T�i˰$��}�/��T����mԊ������]pͩb��ON���� �����W�d![H�w��m�$���9Z��˸zS��B����z��Ѡ��gh�����νu��
f�u�b2�6��8�%���.{�"��į�(���6���z��	����TE�h�oÒYGa���Wo���:�=��M�ԍ�Ip��pc~o �c:5�ez#W#Z�nT�_�O�2�>z^���?>vҳ)�גCGćBUZg�h��f�#kR���[��W�M�Թ��sT��.�E�4Z�A��E�mtJ��簹2��v~�u(���nA|�������`L{9�c��"13�Q�R�N��l��d+;��|���V�B��}�UT-�+����>�$���rd����2�]y���O��ϋ,My��\w�k�*,|�����d� >�r��/p;�49ؿ������ye�0ǹ]J�5���޿��w��<d���c�5���!�M+��/��3\?��DP0�Ƣ@]Ltd��w�p�s |�`�r���dL�?'���A�'��d�~�<��@JZu�k9ܿ�Ud5$�r�%W������J0D��%�l��rG>Y(��hAwU�A��I�=W��u'�_3D�^ҝ����,���<n�9W���>ܶ�yV)e�OO9_1s_�7�b���e���"�P���3��v�T�f�t�/�au��}�����g�"ګH-,f��g���)�5�q��5��/|����y<��Q�h�"��*x����������?�([o�W�1�U�1������I.��e�����{`�T��jSK8}{nNGS?:�%)�nsO>���~s�:���:�g5��dtEY��%C��F�|�VK���Uց���	����oq�n�9���Ҩ.is�]�ͼ����Y2B]ﲯ�M��^��zy�Z�Yj�s��(_
a��1.�$Q�$��Ac֫^\��G*U}1���� �B�Y��5+�o�r���CDnZ{�9jTm\�cp�{�Ar-����i8����y}�#}��R�φg/Jy'wI�,/U5\�h
�F3��o8�M�u�E��
�S/���rƔ�_������0�T�^"��{�����y}��g\������K�&����U}��g{E;L2��m�����7$�.��Z�h�Ã�m��oG���?g�ؼOO�G
j.�u��5:��$���r�Uu�i�����yXT����:}��hY/��l���~g�)�Lj&ԉF�����B��3Z*���B����d��k������Z?	�-� VxCR�g�WV�V?B#��(�sI�NK1=_�Sӟ��¶��a�l
�q��yL����i�/�x�-��Q����Z���%[WX�`f���K��&����!��TŘ��`��w��g��`�(�2���ΰR.-#۪H��cx=���ڎ�Z�w�#Q���k���5��`�+����W�5W,�Z�n:��jʘ,b:������3[�WM`_��#|҉ݢ7�����xZ������4쁻'�&���ȅ����J���4^ȁ�?�J����*�pἙ 1��V��1�]������sxn%��ʌ�����{~&�;N��ۭo��x���P��E^�"aNC���� �%F+w�B�5�9���/�T�Q�Φ	3
�"/K��iKK/�k�����O�6�r�<�gD������X���
����MB�>0��û����/��x�x#Y��#+���w%�j�4w��k�3�T��B��τ�'�/��Qc��M�O�	݉v�xp�B���oم)�5IO�e<�T�|ZS�^���EAS�r�m6a;T.��:h��b�OV��#̯�ſ�4n��6$���q�zN��?o��:}HQ�~*�O����a]�Q����#�����-�(|����K�S�\����'D��A��a`_���������x�Ѓ)��(Q��Rb��0+�ig�2�t��&�i��R��}�Ќ��	lW���h��RҘ��u�ϴ���\Og�����9�{�*��1}�nop9>�F�yXU��QO�pǷFΔk?����ϟ�����P'T�Kw��㏹�?��pJ����8ٜ��7�7���~��*�!���̜��t���wY�ȓ��ݜP�
����-l	��r����/=��5�e�ĭ�a ��P=N\��gd-�j�_�O0{ݫ(�c�h��5>�>7b������fe��c �`�k��JY��ǔ�_�^g��>L�����/�;nU�.6�v&�~Y�:��3��FV�8�EHt�S��~t9ǉ�+#�^�	r�*F����f�iHJ������|�+�:G�����;k�7�.o�ix}��d�����QZ�Ġk����}V���E���K���he#f:>�yK?ss
�ggz�1�%c�r����ƨ.�=�*�M�����V�v�յp02+�\��ʇ�aL�w!��e��Av�s�3e*Uv)#*��'tRNY����O�w�V��U�@�;�2�{��r��V��Sl�n �&R;:��}�V�����
��J������D���p`�9�ru-[�B����W�������g.Ƙ��㏄n!�����e�v�-�!�4W LR�5i\2SU�M{WKl�h�,�L���/Oӵ*̪j�\R��������`��ʋ�>�w��e
���MPU͵gx�{�Ԅ��U��:}���C�Ug��f�&����hs$>����֛~�xA��~`�ņL[ߟ_�/�j�+��j�6�@�;�?��$�[g�����e��t��s+� ��[<Z�\i�{z��@�X��_o5��aCe�g�C�P#�-i������ev��9��Э��}ʾ�_Y�2���=�__��o���-�C�p���s��Sjj~��)��o�����?˲o���p!먡�Q���Q5�h�M.v��a�^M�?\�o/�d�ֳ.��H��L��D�u�+u��ɫ�
mA�d?0G��o|��nj�0�	)���0~xpf��C,zt��«�-C�R����H?�{j�W�|�SE}�7T��l�g�c-�TXG���l��� �+��㿌K�#j�r� j���,M�Q���T����d��Vb�=_l9��ko%\}�{��-?��>�r�h�
9a���-����{�ј[WT[j���E�,ʌ����j�/PwnNڽ]C����+I��>ZC���6���������m'2G(B�]��*��;O�O�`��+�G+)�Ǽm��J?�Od������%���op�T�A��,.Dp���uT�7۷�v6�p�Ep}������p�%�����uJ�)����t�t\�U������44.9���O�N�4ߺ+r�/!( �_U�JE�J�m�
���ܻ7����r	��_�?˖"�>~� I�`����3��P&AG���ĺ�~	�����6�V��)��嶬,��>ը<
�:�gl�*ós8&Vu����6�/-��l�����?`xU&���lM�A�E�Pz��F��ڕ�8�ͻde�.aFi�e,�=����9�Vj�Γ�J`@���F�N�{7L}VI`�R��K��T����\��TI,���m%���;�����UN2�*�$��ʐ�շ��Ju6s���'}���&$s�N���8�R8�{��pj����.�sS��	��iy�
�$��}�\W��͘�=p����<����k[����\�"��U��q�f�<Ú)�s�K��QP/�o���U�����;�3�'X佉�`Ioe�A��ji��b�*.�<7��V�^�*��"�|qf�L{�2�ULӯ�0"�Xp-EX�7:��Ք���C�1�vH��	�E�����_K�I�B��/��N{���O�<���x��ņCR��w�ٜq��	�j�b����Z���1Q��wS��W�! ���9<7p�G�h�ΘMC��*�V�|�3]��;�8[���S�Ұk\K�����z���g�md�ֿw�y��K�X?�T��,<�ZcS�*���2%��O�\�	�!;n'�VJ��%4�J�G$P}t�:5�Ѧ0̻��|5U��ӢMb?R�H?��4�<�N�C�m�R�j���D]cos�"�3,,�9d���ō/
�b���e�����kST0�f��=�s�y�:�P����~aVU��ϙv+��Y�-�<�Z�t��5�+v!{҄3�Ě�FQT�!��jM�
^N`�P8���@拁c�bU����-J-�\�6�� �dq�OY�H;��۟ı�ux���2"�|�[,x�x	��OI,AٔM�6�}G��s4�}�
@���Z�|M+E��V9!�FS(lG��h�^�D��|��]��«�@#W�,m�?�aX��y4���+dw�t��G�����o�L�����܉/;�1����f���=X����MI5k�֜m�C����(tb��5��B�:W8_$;��Ӭ���Ph�����,3}���߉�D_<��[������V}�(���(�$}yz)��쪥V�R��i������N���"�7��3u���B�1:�����)!_���n�s��nh���U1���V��YѺ|޶�����	[�Dj�t'��h�CQ�p�ä����焹C��$���h�j��l�s�~#6�hB���h�߸�	���l�y�Eß2�:���}z"6��h���|��!3[�0bu���ڐڥ��HTֈ�Y�Y�� �C�s�N$)�R���DnEZ���s��'���};i�H?-��ҜZ9F�Y(��G���$�����w7¤�#a�R�����<�(�_DjwS���� �*1ʵc?�6�|�N�{@5]�>��}!D_�k�θ����''�������RR�cWu�r|�训D��(=�q��T���j�� ��"��o��锉���&r-��qq�����rV��Z�@�e7{W�LU��$�ԕwQ��V�#Q���݋Z��ec�:����b�wp>�}��}}o�)��l�?:���sԭw�>���v����,O��PɌ���ə2��[~��	����7`����`��́GSc�Z��ZYʉ<f�h�z_M�0;KӰ�a�?�h��_����f*��7�C�8q����=��
޾�"f�{n��`h��Z	��6y#��jS��#w�/<� ˁ=�������Mœ乪�*p��+ d��.�;n��=
G��>�8���*Qk���&����o� 詵�\��-�.�g�P����&�~z�h5<�|�3��jdgfx��h�"��Tw�	YS���n�1�UL����h��F��i��W��P�hjEe:�aZ����xG��y������e�5R~�#��NA�\�ڮ��H�h��]��a�$��ΰ�(�>�z�=8���x`�L��d9�����uK�v����S������r�ˏ��h�-��Z�-���Y�
~U���r�ʝa�'��11�&}����[���S��'@���h��x�+T� ����'���I>���[�?�1�8�\6W�Ǯ��&�����;�1�/Z;�E�h��ժ�����]|�fx[����u@�^����MR�ChfŸtr���p��G��L=�L���i��D��,O&P���),F�$f�o Zc�G��i?d1��Q�=u����g�����8�ߏ�:��^Z׎�&q��UOU<g�ƎA�r��Qr��kP�a
4�O%&�&WA�ju9�R�qc�o�PemD��RT�M�7�b�;�5_�	�������qŉ�wY�@���W���B�1?gk����x{wd��*+Q����t��`,�aH�M9���g0E�媈���>?{O��W*I�W��;��Z��JF�����������_Pӭ�C��%Y�"f>8)ٿ�%���*����������Y8c�P���IW9AldV�_<��n�ć٫����}�_oA�����Y��:1��x9%���}�]L�?��-Lt{
��
�*�W��ߦ�%����K�B���pM�Y�����֎��9�j,����-nf(����?�C�j���5�&�A��RYFx)i�T&�4K��m=�;�8�n�R&�
���Ϯl"�ǽ qP��2��5t�3�>���k�}�G���uL��B��u�,���`�vd�qư�"�ٿ�S-�HUmKA/�o�����0�v���ʲ�V��xD���',��WCȀXq��ϥ	�˥�{:�����x��SV���
�֗��
�)h�B���<�i��*�pF\�='<���v�bE�̇�u�N3�?��m��y΄]$B�7������q�b�XN��Ճ����p�a]3��$��?�(��a�y���G��{�d�Ap��{x�����"m,4�~c���������J�ʃ�Kcܩd&��u����E>_�߂�(f}���4���/6ǣyI���H�='�~|R|�)ک�A�ʻ'/�����o�T;c�Yo�'��@8m[����V��T���J�U��l�k�fV��O�<�kg�xԱ�����@�*��$�}�ɪ�L��e�<�0+��K/xV4�\O���_�$|��twm56ד)�����'$����]4�*h���m@���'�jӍ�K���6�R������gvɿ�׹K��dy�Ϫ������K�c0_֜��>DY����u�.[����eU7cuJ+�z���j+d/n�(9��['�Ҍ��v�X	O��U��=�D����گW��n)=��E*�el�d���w˦�z��m?�i�g8����t�ݖ���h������U�W�y�TG��i�y����*��=���N��"�;�C��ޱ-Ϛ4~�AР��ɖ��^���h�dTw0byi�i�*�_�[�i	���䃫%_!�y����,�Y4��	��4�s���镔�3?\v���3�_w����E��N�3�>�.��ה�S-g�4ٓ�2.���܀!�v+�f�YP�Cz�,���Y^�荘_�<�V,�2�'�	O�l\�0�b�:�y0��/DeUCuX��߸�&t5f_?b����2Q������D�9�~N�s�?g}����|�{�?͡Q�\.I�,e}��_��kU>��>��3�|��e�tMƷ^aC��:�b�A	?��YyuN�}��Ͻ�������T=�����E�z�y��<7P���޴.���3�����N�M1�̉ڑ����������0X��mr{�*�{>�����%6D�5=V��_r(X���Ǒ`y�3z�G�d��n-�y�/r��vJ�Q�L|�U�K��Kk����2t��oO�7	�&U��!���'W�]�GLS�=󂟫���u��;�P[Ҳ�z̩k�R[IG���u4	�[��pY��0�T��zy�K�j�?�w����v#Z>Sa44^)47Oܼ\B�� �j�=	v���e,��D"�4S��͓Om���0�|�C�:hp��ؙ{◻$�v��E���I�y�?y�ꏑ�G7T[)�Y�Y�u��s��n*"�*px�$[���L7�;K�c�e�PR��ILMAUXW0������zW?��{����5�Y/~BoIYK��� �<�?mq�%�IM��.H6��v�����\��|�
"��V�WW�����G�/I�rа�$�A��Q.�s�3Q�s�b^�A���a5|��0�&�p���5p?�q��1c�V� �U��������H�#�m�6w���Y�G/�]�ˀ~������a��zT,�i_�}:ڱ΁M=�R��E���r}���ў�#��%|s'���5Cb嵥��V`A�XVx�KN��:]�_2���G�����?����)�s]\����v�����s\2�\�o���/�^�Z!���{���
w9Z,�@k��P��M��wf�_�L�W͐�uFP[A��NK;���ܒ
��Ψf�l���� P�h�'���=T5�+cVT�OT�������.���0G��;T�s��K&K���n0�m�ұ��(�"V,�qe��A}�n"����Z�Ȣuu�	�{;�G%���>�J������ڣ��'e�N=�M��F��i���.�N*�ѐ�J���yN��a׶�x�򪱭S��0�p������������g�Ev����m���7�Ìl����J��Q���q:���h~���b�3Z�������MbV;��w��ZK�^6���^�t�$���Tag ;�Q�
�^:V���{�/dP'D��Đ�C�Ҹ���r�c�E��/�\N2gs��Rf���"��o������sy�9�X >QM2��?����]݂��T.�A�{�t��d`��ks�� ��<��\��f5W��ɊҔ4��v��:���	�æ�Mx�eu��*��]km��y��#���+�Ta��=�ٔꥳ�1�Ǌ3��r��6lڨ�|ߏܓ�b(j��¥����kz���,M�O���2�'Zυ}l��a�p�:�!��R6��֫&IF�*p?�{�/���Dn��#����ɃI�y-DC�P���K3d��B�-��9��hO~��t���1��y@�]<���Dӹ8��r&��Qz����b����o>1��_C̆퀘��Z�}L���|��X�j���3������'��e��;!�"J,U10�u�3C�<�'��k�=���x�7%�m�`TD�Qh�/��.->�a{���Cz]��;n�bm;�Np��M���ٚ�{�P���}����~y9�XZ'-����_c��yI'vW����sr���G�4��r�%�X̩(Ǵ
�lJ.w`��	�jU~����)$j#��ޛ�eĀ�f�^��*������+{�V ?pn��4\�����*Rޛ��gv9�rsR�+'nsxKE��j�V�������^e^������x�4;��	�ƫ��yV��b�|�W��Kü�=�(���E���#�u��<�S�KB��[|-��vX�1�È!��9�X�<h�̝�����Ir�l�J�����Zm��R�%C�A����rv��Б�_a���eu�F&�w*5��,qJ���J[N�>�:�cF:d�ǭ9������XS���
So��5�9��orf����6ټ��̛m��"9��"i5�{���0>�/�; �Gl�}��.�⪶�G\&&>[n�⼥�ߋ��Y���)0��\�0d��m|\>4d�wRǿT�L6��ۈ�ÉY�qE�5�u9�|B$V��DLϪ�h��_ý��g���k���}���<�tqj�0Bu�:�3�^:Z~�8{os�cu��hr�k��?�J��J��z��3A.�2�����	����L��b�)�D;�N���`	!��y�W�{QS+z_�?n|��w�wk	�+cV���-!b�$�U�ũ�{��ߔ:�b��W�Ps\�%Ϫ�Ld�M}fq��[���~�3/�N�\�5cd�r>I�oЇd/�ɮE�q��T����������|�NUi��$rӭv�qGX���~�p���S-�����u�A6��@^�h���Y��G�F�E`{��?��5��i$��Uy�"x���*���K/��8�W��r�ud����x�H�����J�����kq�6갫}ף�z�������k�:	_m7�c;Z��5�g�T�Qw�:=c�V0�;��Z���e��`k�ujy��G��*�,����x�ߏ����+h����D�;tx,��-g���/���Wp��a���d��:_8Kt5��r7A�)�?6�\�u�ùv�����S�LQ��`��;Ń��yS���V�Ⱥ��B�T�����uk�W�0���0�A�.�m`GHg�Q*��FlS>s�aMwƱ�IX�	��4�yL�V��-
S�/�AXU�����5����B(-'��:\�k�V���T���\��!��,�i�i�7�]��|��-MVV��@)X��4�`x��d��Y.ݩ�3��7�hw���:at5��;/��&Y�CdA󒜞*��f3��5����ْ?u4��H�$ĸ�>V�I�UPj�ײ�9C�c�ͣW��i��Ԫ��r�l-@��x+��A�_嗒�M��Һ'�*�Q>�P�r��n"
X]��=�/�v�2��U�R��7:�Kk�͍�s�r���?��a滒+���2g�!������볈��C��S}��JH"��
~��SN�W���\39�,ays_~��W�	[��$����E^�����9��WL��)盥�9��/�p���>��m�@S�K�%0�fl�����i���p�oŊ@��1��?ڭ}. �E?Ew]<���K�݉J2���9͗K����]��L�γ���}��c�B.3�Xd`��y�>Z~�����w��v�[��76³+TU<;F�NH�S�zcE�C�ל������Ft�,�z��Z����{�U�\i�~"LA>�k ���F�9��Z_��b�ǋ�M�sK2D{m3�xhh<�@��0#��=�s�牢�w����7�/��O����T���|�Z����B�2��L�g���>�z��Lq[c<�,#�TmP?'"S�/oy1�s�m�7�g�'^~H�\����^�*	�}q��с�l�Rmo�pK6Zʃ��9ۄ��r��M�#�-�͂D���!���{8�:},�֎Ԉ�3���%yXO��E�Ƨ"�Lm�|���K�L�]s}��Tb���/�_-dV���ѶS�-����ԛ��nwT�fjU�?86�G*�E��d��O��PAxV���Ķ����[&�D��$����Xk�.�!�?U`jX3I,66�CN��{u�W]>`���O��^e^��F�#�b���6[���(�2��J�:o�a)�^�K����:3������XA��"�o=��OYTq��,!�3�~�1�5�63�ẕ?+����ҨG�������2�Vs�!����֫��������.�Ll~�5x��ȳ�����*Z:��yͪ�a��L�����o
2�j|u��1̀h'��緊Q�!fU@���@�h��Y|��7<',[]؃�gj>`	����[�EM�?�K���2:�U�����=�mTi�2�m��[?O=P�^�:L>��%����q
A �@�\���:r�������f\�dtg�{�e.��p��΀)��1}�3�����E��?��2t]}4�x*�¿�a��C�������_� հG0[�Ӛ�1��I;U�B-�h���>v�A��Y%j��^��d�s������e>�~��u�o�xD���4��qj0�X��	�2�?ʥG�Ђ�3�������ܶ��N�S�=w\�.-*�!ٽ")V>.x���;�1*9���U�*#\̀�L.j!��l.�ûβ_��o���H�dl�k�Z^����]3���ZJF�n,@�,	�K�
;d#��Y��s?l��������bӭS�AY*&Mx{���!�7.?�YUx_�b�<{n����#����C���x*ڨ͙L\�������8|X�j��Z�+h�F�/�W�M�a	}Ј��K�?�؉�B~��{�F+m�rR}#�ҿ���c�Z�T��Ra;�=S�e�Ȝ1q��5~��P\>�3�6���nߪ���3]��fC!¥�c��(i�.�7�����wb�jb��Xtr�Q>��׆>��%�Pv�.��ߍ_�ϝ��z�ŷ�-U�#W&���<e���.���l*X!�k�<_����^{\������?�Ѝ�6͌N�I�O�5Ȧ�
ߢ[�R��~���q���#�V�����-���-�0�hc/��
11�������3�&Y����u��p|p��g��*Q���C�H�lu-C�~A�&s���UE�u���U�Vc�,M��e~Z�m���ܖl��Dԓ�>F���?p�����l�2�\�7+a8�*�H]��Z�)-�<gD�*�L�$��4)�
��ȉ���FP��6u|�~���6}�3Z�-�V�����]Fֻ�l;Q�����7�j-���
�����_(��G�~6m�c����)��wB�_��WTTO�v P�1��й���fۗU;���*��zY}��4����W�Zza��>�3~m�iM�tG���J��Z��d�P���p*d�z�"�wPaG8W�`_0r�A����>Q��P��p��M��jW+�����h�������D�e|�f�?���������P�Fj������p)���CZ��l�XcVo������������K��Q�E�E߶� *+�R���v��ܒ��!g���=�DR�Z_8�Bv�c���I?��3�yK�冻�C*����H�cUY�v�G4��~��x�c�eWb�xq~�n��n��Z[1
���kW����D��Z�gZ*���Yw�'^��5�8��l��.��e,�U�=�%����h+vx��ri��������%]m���]��֯�Mt�U�s�v,Z���+���ť�x�g�vB��lU�_:5�\b�Zs%�\����lp�b^;�C���+��u����r/�>܈7�GՇ��\,jGO�Gh����ט}b�Y${��R�G\��o;���zH��h�X��q��	!K�UM`֖�?B�mIpτq51���1����cqw�&� �|�W�Ѩ��+�*��ކ"`ٺ�H�"*�A������:u"�����{f1xǆF�uA'����4o�e�P�� �(�H��Yw6r�ԗj�h�⮿��eR�Yв����,f|_V�,%|��>�C=���HW��<�<���1�ï
���D�N��un)���u}�e3�$���e;��x�Iz��43Z�R�B5��9��)�-��ǹ6�"!�[�N�n�[��z���4m�?����4:��|�X!*�sT�
*�� ����l�J���ب�ޔ-fխ>���|�s�X2�)~Ë�����S�'�N��}��d�}�o�d4����3�dK�y{���=�r.X�xE���[�>�?I+��ޔ����� �}3ZԢt+��!nLJ$�z�x��3�.�>Z�O��%3�Ү�����*ʨTl~��#wӼJ=��.�e-�o����~mm�zbA�R+FŬ�c�1k����y�杁�X��c|V�5{���'�J�J}���e.K��?�>������U���0ԂդU��ى��4�o�.%��+q�����.h�v�Яk/х�6�%WUc�&U�����:7�h��q�;�e�iS�^�ת�s w�)}bLO�WS±}s���w�=�[��^n�����V>���-
��r��5B�}4����x�δK,
�Phu��#�uY϶;t�Q�D��+�!h~}���*ȳ��+�(+~���F��/Z��wc*7	��	�T�DjH��+�Y�ɪ���
/��9Ju_I^�X�
�ZX�~8c0��2ژ��@��r�%)�7�����A��G��/��eOx��S���eV��m����:(�'�-^n��?��W���<=�7����vc�*4��xl��uo��N�Pq������1>��Ɔ
���l�a8�OZ햃>�6��|s���b_������eK�%b��ο�Q��:��o���ۄLc�l�?��̾n�ݙ�}��4ڡ��W�WE�`�V���I;�Z%���X@�z���u5�W�����f�)9+�����'t�!��CϬj_�ߤ���,@;ST8Z����a偵f���^� l
�+"�j���zqm��k�s)�HMY��*Z���jŒ)�&��G�gޛ�U�#j��;�r��vtQ�$�&�*5Wn�EK�P"����˹]v���Q���K��l���:��A���Z������_���H�s��u�FF<t�y<_��1�6���=��nk�}���u����Q�>�<������Z,�E��_>���p׵Nī��1�Yqܢ�^�|��4�pD�+�#���w�+A��W7J�*{�N��qY:���cV`��B�����'so�������L�U�P���w(��R����9b.1ZdW�O�ǉ���F�@:_�2���8�»��3�^��T�v.�/�=�%A��˫*�[�U!�^��;�Ǩ��)q=��R�|_<��o�3}��B�l<�T�Is_Li4��ۉ`>��Ĳ��ӋL�:�-��ّ��a��
(_��*?��_;�V4��~֝:;�T�`�K�~���<�?��r��F$�Jr��;��.�,��F����zJb
�8�!������U���N�S��vn~4Z��Ծ�q���D��O��JMy����~8*A����h�Z��A�*o��9�Q��ܕ�ӗ����7;��-`�Qa,�?4!�+��?�mڳЕ�~�t.NHj��Oi,!����c����xu�U�MҤ�Z|��P���o[V�������<p��{��œ�/�WjH��F�+���C����ػ�D�K�ZL���"�|��V=;��Ku;FZ���j��`���2ޥ��E��qcc ]!VU�c����F�al���W	��s���zw�fg����<~I��Kg���|����EĻ8���E��,�j)[�~�>�*��z�:
�=�f쓎��.]����.��Z�ܸ<\b�Wy� >]V��@Z�㌍��ڊ����g���,vU�#}�#�|N��j�h�V.0i��"{���{R��N(|
x~h��~tk.*�GƀwO���K[�i.�z�AU%n#�ejK�I�:��I��Jg7 �TU��(nO�Y��Z��	�l���P��x�j��V9-9yr��<ܶC3�Y��/�\:_��ȹ�����D�B�V�F� ��_��u���- �����f��О�<"̮u�Śz�>�e����88R3�ڜ>��ʛ�X0e&���=���YPRy���m����*�>����lKo�Y����}�Su�䧞;�x���9�@����4"{1q!��Mj����+{H��s����ȓ�3˺����!�y�mM���;�M2r��l�z֕#3�8ÈW����i#(�:�wjf��u�$IY3r�u��h2�j�si�i=���}芜��{)��S�N���r5k���ږ2�r~J4G^���g���Ӛ붽M�pc
���Y�� �|���'��=��_�e(_��2���J"M���R�
�J%A����b�>c��J!��C�i�?�`x�*~x:J_HWp�hxi<�dC���f��i�����C��V������&�P����D���>�O-"X7lV����<���Ѯ5�������������pu�
��m���&��>bD���琥���xW�~H�-{3�n=�z�o�@��t��ӣb�%��о{,��1:6U�5ʌF�a��|H桮�_�������W���L��%�Ev��&���C3�o���eY��N�|e��MP�2���z}��#,���O>05BI��Xun�dc�A�����lrTh����B�0#E�T'x��1?Yt�a��Ûa��P�qw�7&�(�������>!X*�ݱN4���t��iU�a���g��xt����LKAՉf)V+`�6=:ݼMdT
�Ӹ�UF�E���*_���W&O�[���1�1Mj�v��.vLq�V�]�!$;�`�Oy�}q�'��&3T?uY���&�:�Y�ک�U���?������t|s,�Mn�2Ƙ�����缚����D��]��\G�rj�S�o��>�]�t�#���2���&�9�R�.ǭ3������8����݅�=�f{�og�dt`nU����W���vy4\9#�A��QW�!�Uĺ
k��D��_ddO!�Y�]�o��d���C��Z�2Ù��Y���3�g�x�p�Yo�:$��@��-����;T�}�xk7'_'��떬��=
%ㇵf˓�����jџn�OJ���i�JL���_��f��7��;��f+<���J
��g�Z+�?�.�E�3)[j�~�¦_KO��
(��Q��C�vJ ��pR)�Af�R�J��=.Zu$K?���=��C���Z��]%3U�7�<�z��i�f��)N(Z��,�	�j�Ŋrq���M�i?�]]�3�ԙ̲���y��n�}ϟ��3�
Ts���ȹc������2�e���۷b~�a)S��-K��P��<ϷC��b��=_%}Q��L�t��C%t��/U.��s��n��t5ݨ�UYc�t�r�z�������]K����V���v�p篮�ۓO��W+y��o�W�]����UE��oc�-�PvX�>����U���cNnѼ�<�<�f4��4�7�����S�[r�~����E�,�/*H����t~��3��x��zʿ�n3���p���z�����Ϗ��@�91�kt��Al�����I�a1��������7��[�v/�M�s�F~X����d+�=~�u#'Y[����>WI�t9�z��"q[��b��!�\���Xu��?i���-p_�U�W���-ͪ���Y����ƹ��b�}ؼ�{�A����"w��W����������Ν�U}e�醒.͉=���W�:	���&��Bn(ZK\wS�0�`�G?Y���������?�(�ÿM��0a�lUs#��~Y`�0U�����Ϳ��^蟯�罰G��TTR�5V�%��P��[�N�{Q�^�!H�����ߞ>|��:�J�A��W���R_���
-�>�ܯ>Eb	�n`'W�e����
�n��pO�Bϩ�Kr��Z�%)�E�l_�q���CG^^s�A��^��2����٨ER���ل&~��ں�����4gRJf��[(��
7�yV�y^��R|���_�9�Qۨ���V���#��MYw���Q��<u,W�o+P����ز��E;7B���6a����#V��	�w��__���7�#����*�bGw�R[bP�ԩ��_�ds�ك�|of_�B�8h;ZtI��E�XYu_���/�_�#���l2�OD���w,[�q=�UD�hHd:�?k<������������)�>P�~�͍��pԴ����L��b?X7��v��r��('; �m/��|	{�g?o�o�zX���u�7��< yYsU���Jb���t^ز��4us�ţ�K��;S���]����q�����UA}���=q�%g��1�N�yM(��"�ӡ�0̾8��
����A���5���\�8�7�~�թ�be���yr\��ޏ�v��7TQ�pE@;��e�
n�b*��+,w;y����wJ��.��:�F�3�꽌��U���3O;�$���ص�h�Tn����_	U ��Z�3��Y*�w��O8ǵK�E�Oja�#��V�4D�9��c���L�WW��^���-*m�F~y�ǃE�z(9kf�[v���˧6����v�7[�U��@^Y��N��u�K�� [�p}hZG�D;�5p=]K,�|6G6b���.�يd�vUQѢ|��P�Q|_H�_�C��ޢ��`K�k�SA�_�D���^��b��髺@RUp��Z)��x}�q��J-��*���\s����XJ��#�^;�h~�K�����s�}�ܤ2��:�|�u�	T���ȔSu�w���!�S��?�x��J��ͮ�gޣ�)�."ۘ^�&j�pK�Z��ge����%�f�z��V�(v�pI��:�����ob����|0>�+���Ԓ���P?%�'|^�k�8Kb�=	�h���(r��3��کi���XK���Lb!m=���2ʪu���F�>�<R7�S�.!�K ��z��g�ecTƗ��n�X��\��������4gp�w?VX�g���O���1'�������,<�#�sg@�I[���Z���'Kc����ї>�}�>��W��lm��Y(Z��y^eN8���v1�uG�.�?e3��7Ų$Q��6h�avN�T��>�����(wY�h�n�o~oi�Bkl�r�w��&���Z�»�x����x����O���H�F��	_3!Z�}ꛡ\x��
��.m͌����z����jx6z�ˎZw֩�'��0xPe�ѩR�x���͎{*-h/�I����V8��:s!w�
e�6.B�Kw'ZItF�2h>X �����@��Whh���j���%��ǁ���'�� 3.�茒;�Z�|U,��%6��M<���w�+�������������tw�]º#�K�vV��μ��ڵLy�2�]qfi�=�6f]�z�?7zt�*�D�J,fE0_O�o�{3�?������:/�ܡie�������lR�1J,~���9���{Ǥ��*]�U�աy��G����u������̫�*�Ohq�1��>��a�6Z��q4w��9/��a��/?{��WF(+�{�˗�~�4AW��(�<:O&�\�OxrdUE>��� ]eS����\�"e��M���S[��&�CQ���8G�/�⡩C�$O��`�����ho��U_��yېi��L�r��1�Y���gUuRc���L`���'h�KC���MjUՐ�/h�ج�3�:רzo�"j�3ܯ��fn;��A���"S��|���)m�5-�,�^�z$��.Kr�ӘŻ��ם����I�@(������}ra��c�i���s�����6$�_��d�-uRHA�R�჎U��bp���E|�-����)<QO?�+�p]�I�ܷ�M�FE�����O_�j?�.�p��m)��s��Gn��3���0[t������D�M�v�.>��X�?{=ӵ�����5P�Ǟ�p�V�
V]���Lh:��~�w�`�݋6a\ܙN?��k,ڭY�Sꙵw�̈������%���#�vJ���;6�?�_��ξ��o���4��E��P��2��I�֒�a���Rw�Rt��5+�#�eI���w�z��<1~n���{���=,�?2��C;��ߛ��2�v��(R�u�-��$6WE�/D	[=.���K��HTz:�ƾ����>mGJ�ݬ�3왅%�������0�ŐT'0#��^�N�r��'���	��m�燷-g�f=7@�U��}RYC!.I�S%�;�,f��a�]�C���{-U��_�-�s�u�_��(1.����F�jΕ�۰Y�v柋���h��V�|��Ϻ�bvu��Vqa ���p��VXV?�-��#}�*JH��{
�����)T?Bt�*�ì��O�<�J������ٚQz�u������������6�e���s�tߨT1���+OU�>�bPD�z�vb��&���ژpkoҤ"+.�Nq����hc�����}��Ub��?b)�6a.O&BS��ߚ��K��EbQE��:�����A�aq�ZnIVU�?�e-�������#��1Y gWS��
��<{�k+ -%�'�9��^��n?�/��Oj��fv;+/�_��u k^��w���?�g����q��8o `��    X2     U�����SWV�E��U��Ɖ�f�>JC�#  ��
�E�   1ۺ   �C1��  s�M��  E�����   ��   ��   s[�   ��   Ht���   ��   sU�   ��   �GMu��   r�]뢹   ��   ���E��E� ��t��   �E��|����   �   P�   �   ��AAX	�t���^��tfA�   �E��G����~   I�	���t   �:I��U�M��1����T   	�]���V   =   s=�7  s=  s��wAAAAV��)��^�������^_[�6�u�����ù   �   �1����������1�A�����������r�Ë�]ÐJC�      <{� �#��C�����(�>�*�7f�|`��J�A��� Hԅ�����dF�g��5����!��$�Hhk?*+�����'`���X���s؁�|	t�@X�iY�g���k�a��3L/;�	B����B���ç�C$i����j��"~�O������3ۏIe'��h���]��S%��+E�_�Bl9U<|XI<�LI�8�5��&fx|�Фg�Lp�9Z�"���q��BO��qB
c������i{ĠybzƊ=j)��L��m@�}Z�<�t1�Uڒ<'I���Wk'�/%e@�	����G��8!H���u���|�}�f���O�]P�)��g�*\\�&RA%tԠD_l���gF���+5��-@/�ď~�-��b����Lc�.�8G�$	�̋���6�gz����]��
��Sa�
T��4ӵ�ˍb����7Q����k�� ���X��I�|.��WF���C��"�&e����2���4�5����n�/i�✁�;�g�������JeE�gӅE7��4Ӑ��o����?]��;!|B���I=B�Ci�(%�s��r��_����*bsCg������Z��/D%�V����bA�\�5�(`a�G�A�=����P�mh%���5�p�BVUM(�i
�(�!k��!�8^+�֋����`)�as2�$"˔-�z��S� M��"_�D��L�̆�b�)A�`�pPԆ@죐�Sۈ�4���S2Ng�)�0�fm�3}X�7��ٯsS���=�w��>�G��TC����7��3QL� w�:\�ة�5�p_��ɫ]m�ga���KQ{
��?�����j*L,�-w63��!C����>Ϫ��2�{g���j�Ӗ�0 �#�q�ɂ��L�ƴ#�^��ԘB^y�g%ƟQ�Awm�[�/��ؿE��&�ψ��i��14/�1] �/��!������!P�'�n(�4%������Us�wi������~(�T��MO��Q}��v��^ݔA��'V���,иP��:F�E���P-A�̎��c�J�)"j��NtZ^{;5x�ت��vڋ6�>��u#bˣ����z�Ϋ�����v�6����Y���jK����Yε� �7��|�x�����#| y�%��8C�)�FҔ�[j��c�qT]�"�*fzfc�V���U4}=���ĊM2���yp6j�g�݂����U�-��~�S�b8���?��h�K�/��K��T��8��ӕ$GK�4����Ph�"�$�:C�𑳂x`P�j�&R�nQ��%l�����ϼ+�r���D/qܻ5��E+�/�,������Z�	d�O�
�&nC�&->2�9�3�Bٜ�(�'�"�����e�<.�!�-����������˝ɄZ%}n��=c`-g������A�0���ޝ!"��*�����/	ޓ���O��o�͇�k
���4�T鰈��n�uT�鶤�j�@*�����Ϥ*�v�	|n�hCT���y��@��xE��k+/�r�Rv�s.P�5�gj���L�ڟ�A�`N���\
��U��~���ѓ�ި�J`�kz�ܲ���K�4��S���ǣ�L ����Q��*s��M4s*���9�GIEη�).A[+4Mt��%l��ѓ�{B��)C�m��~���@O�K.�C�G�\8p;�
x3�������u��Ef��.n{�!����|�}CVt̘���
�x	�&;bw>�X⦬-���Aw�@�����4����A��8��Ik���A�Н
-�s��Br1�كxy?N�:�<��)�	��oΈ�w������I�cZ�6���_/_?­=b���)09�Z+(=]�5�>���y|��/��!��3��ÕRT����_��Y����(���r.�U��j��o��<�W�C�1���3�)��O�f�dUN������}Ԫ6�?�8�n�4M�L��|e�:ت ����ǅ=)Z	͒F��)zz�N9B�P	�����ܱ�Z�],�˽%Ziǁ'3\�E+�t��]�>����o�iSK�"��H�����- �&�l��C���1Q��6��c�Q��������ʈ|��[�^���,�͵�Q}��C�	U2b�~E\�-�z��;UQ��1Z�D�x��ә�q�l8&3h�ga
Z�����){ZK��c� ��K����͚[�_�>���y�BA%�1�m^
��6a���Y ��6[Fւ���]� {�Tݭ4��%[��v�i��@ԥ�+��l�0oG�l
Ե���FP�W=�c�`Ou����V�9��A��{]�(�}��J���Æ�d�Q�郙f8�C��+�����N1������蹆�o�����G���7p�������\4.�@}r��cy��^�A��(��B�w-��E���=w��_�?SD�r���0~ij����_��(Lm�ݲ�����w�׈���oG��Ze߯j�ќP��]K�킈����&k�����W^*5,��l<�
|�;�cK�>����=�X�m�oBH��aj�܋�ʶC�=���W�+��E.NO��͇�+鰛��H���<�t���~�xp�rnS���z J��}�z�߱ꪠAd��|�U�z��c�%AgAn��_�������T�B���2;��o�|>U��5*��I,K��Q�Aؖ���ժ�G��[��^j�҅T���iٙc����1ǏxpoF<Ο^�w��ٟU��y4�{��{���T����3���C�h���0��� ��3^�wj�G�5Ӎ�³ƀT���o���d�
!���ܓ9�bV;��]׷\O_��}b>`�À�V�4�^%I��OO�Y�lE[����ϣ���th��Ѳ���}�/m�J��0�g姈�i1�ny�P�h��C��7'���۶�qk���o��V��!���~)U���K��[�ޟ��S/���õ�E7��0�}ak� P|��ytɬY|�[H��p��\�Am�����>�\�;)�b
@�����Շ�l�Й��l���
���SLL�V���tkd֌v����C��!��ՅK����;*�ecDb��踾>@���TUF�>�|!E�'.%�5�۽��%�'*-l����.�m��oN U���*ŴI��x���o�m1��;�s}XF* �"F	*+tw��Eک�=,�T)���{��s8��ޓ��S��lMB�p{l^:�s��V{1Ή6��_p��З]�J)��N ~��So�B��(��-<8V���%4�\�W&ܷ�΁�ӣ�7a�ц��\B=�+���'=Ean"�0w�g�o�AggDHvz�hm<=�wL�X%Gn)靲�`�1�]dz�S����4�v\��v��\@�-pk�5Z�E����bc	Z4O���~Z���I`��N�]��^G��/N�1��`�4����}$�@���6]Gז��8b?�8��r��'"[�q�g��'ㆺ�8[��ȶ9Zd���̢]*�G�"=^ �MLs��U�~˸�c�����4������5�E](+5ȇ*�g�t���bzڋ��(���=���h��r���rTE~�}l����A�@��*c�����sgUx[=���%2<nJ�zJ9�{���"T�j+"s�0)̥}�H:=�1�X�nd��iֶʜ���&ћ�{���@@�O3���&!�
{=9�@�শo��+0{Gk:݈	=
��F.���bb���,��,�5�5@*m�%ɕ\p;�1�x����Em��� T�KF{)m���r},�t��m�D���աR���x@�����׋�����g�`a1l�J=2	]�ھ��=����z�nN�~`bH|�Ξ����i���b����	*;�����s��f�+�וe����0���|{�_�0Q�M�!��r�j:�s��͹��/�K&lk�~�$N mQi��M���+?z�d�e 16��o��3�0�S7���T�n`C�]Ѻ?��~m��C:�>xE�.s�sH��W�k�G8�Á�פ���A�F���䖎���e^��F�g[�8j��*aYy�߮�
�]�A:�\��"�l:��%g����R2�b�q����Ǒ2ޖ�;K��� m������4�O���k��hr�Bd���Ѽ�}�ԯg)��<(yÜp ���R���c��	#��s��:<����r`��� ���n8�g7,��ۿ��՞?�՚��2Y�Љ��W��3�|h�W�A�i�F�P��O)e��c?�P���\�	1y����Tz g	��2�[��:Q<4х��ˇTr^Ej��|��XY«7�<W��&{Ђ�Sw(Uh�Q��n.�y+�E*�S�7U��Ey#R)�J�|��g�a���5;�Hi�����U���(q:�6���{e��"En=Ժ�E+�0�y�ǌ*���!�<~�e��ׁ]� �<�A�,g�XS��p�NV
�Y�|���/d�eᝎ�O����f]?�Iـސ��k��J�WC:�������lx�b�|���^I�+h8��P�1Y�K�6u�	�{@����ETd!�������@'�5�D;���QE�ᘜ��e�)���Z��dͦ��N��kZ|-��~:E�ќ��m��R�^d��'���^��aW��n�u/�RK�^����b�b�<f\܌U�g8<��ץ���r'�]h>�F=�t�[�hӸ�ԭ*m���N��G�؏�J������E����X�A�>����od���J��5�U����}o$ 	W)��s�U՜���W�-�C+YϸC��䒉勣����FR�)�ͯ����z��[��h<�'LN||�Sm�򍎛�M"���b{잸V'���� _����/���A��+�8>���7ؘ�Sÿ����b��.	��)o�x��)���b<�F6~,�	9�*xX������e�g�Z:����/�Z3������EPf�R��
��ڮ/��� �]��ȟ�����T:3A����?L
ڂh�6W�cw����56Ԥ0��we�y�X�-ض́ψ+5�	�T�����GY8�dG�7zo��r�W��m[�\��X�c�Cr:�s�� ᥌�RZ���i7h(`&�a��g�@ik*6�֔lZ�˪�q0Z�N�9�����_�+!�#i�~�C7����:�]�/�nN�Mv��R�^����o$���͡)��{�k����ON�������
�_S�~ȐGq=GQ���=���Q�[�iO�4���{�xl�k^գ\Vх
.&K�Uc�w��*Y��3V�͉l�k�Y_�9�X�����k�LQ�S�{�PTKU#?��WU��)oq�)B�q���S8�h;�2E_2��8C
t�(j�>���V�5(+)��u�gI�g=����hs�O]?r��x	.�R��q����C��6ʗ7`h,�����'��!�n�cpT��7N��7$�}h �+4C�K��?�ͼF�/�]��钶P�Rɋ���a��D�&����k��j�ޝ�1[�2�yz�(]D��,��*�f��+\e��3�_��J#�C�NmT{�!�7!�س�/���T[�T���u�a�zR�^Im�mcA{8��]��J��vo�\�N����h�e!Ooٕ��TX�J�ԓ�y�%�X�/\����Մ	b���~ �Z�]1��ƇB��/���4z�̎��O�❋����F[��ӣ�V�dn���y�e�6��?h�e��P�ι�FP���N��kE&����fR�J��\�d}���R���h�@�2}B��؇\}`v�睶hh{;��V3�!��k�\jx�����@���1���r�iY�ev,����9�N}q�����W�*���t��RT2�\�m��w��W����W$�3��r�w�Z��`*o�a����ݫz�kYp5�p?g�e3���7��l���p5Xr�T�:q�,�zp��]�^��ȴ1 2�B�$pj�Ζ+ �����/v��i_��ak�L���8�?�|�K��ef��W*(�Z#l��B������g�fӶ�hq�4m�9�� ˿3���?���W�6������g��χ�t�gc�L�b����~���`�!�#��!������&��W�\�,�F������b�nbGq�|�ыG�Ӿ���٩��D�0�Q^���~��C��F�OI ��љ6֩Iz�u���,�j���7�>�'��)A�,V���#�@�t(�w���;�l��B>I�*��nY*-������B�q�7/����OMf�*�~Hdk��5�ŋ�(˕z-�l���5+(�+�F�|K\n�D<[�����9�*xy�\:*S�8W�q�D��go�q:u��p�8�Mmf����V���v*Z;ه���ȇt�pр�!�ll���YF�6��I��R�U�%�o��������Pfj�Wk�v����)\�����:;��w���4zg�x�����M���Q7ݾ��@�Q\&��|qB���<uK�.Q����7k ���K���١�m��Ңo��MZ���Tс��p���Ȍ���f�[lz|������OJ�EE�nI����J���.V�g��q~4�h4��ǋ]��3�%�Ι�ûҭ�mwR[�8��ڙw�:�/f:6T�A��Us�|���T���j��!�����W�N�wY��21]�K�X�,voa_��2L\\�f� a�������4{-�[�W��ڕ�S�=�����Nwb�F�=Ex�+ �&S/�yPnz�O��Ԍ�&?�1D�WҠ�V����]`��\����%�ooD_��>\��H�K$�)O�A�~���#gњ�w0����o�t-:�4���[;����7���=��c�(�<�Kr��&Zo�f^���Sͮ,��I���T���F'+k��`�`˹n���e�(��*�F�&+���kN?�BM~��'�����",_��C�dыO���LT	#�>M1��MN=��/��[ϯbo��M3�.Hz�wy�r�ĳ|�W��Z�P{��I>��$'�
>��ɿIM��%&�s~��4��h�%Igh����,c�V��~�5��|��zE�F+ߪ�u@13�a)��>-��U-�W��7R�#*;L�|[�o����c��ڠw��"j���r��TW�� :��4�6����1L*�g�wب�a�(A�A$��6Z0��ԒS�ƅY~h�^|X�#D���*��(TTmm��Z���p]T��Ro`Y&>MO/���4z|�i�\�߯*L�����Z��Ū�-j (��>ӫ?YڌD-�W�Je�{@�fl ���v�k�e�h�����DW�ݷE���lGjc�%���|��˓eH-��$/*���ԉ�Io%`U��������ȥW��b�e��0A�8���*#����,��ټ��S(���
�/?p%3��۪�/���b}�p�B=<=��Yh���^���P��zpܯ<<�ѽ?�b&8ƥ��}�^�7�ũ��Yw<nt��ơZ^��;�m_���o7�+���Y��C����9O�P�>`U�V9[��]�+���ɕi��g�;�`\t��5)����������Ϗ&~���j(�ő�Ş^��pi6�5����p���Ϻjfs���	~Q��$��:�h(4�ڞ�=���#U�g`��vE�j�5�wn���R����
YQ�w^�+H({��s�6o�9�<�C��
�)!��W����mA5cvjC���ĉt��V�A4��	�^bH��E><��e���xS��ڑ�F�"4h���N��P
%��Y�̘�2����J�(vU�ݥՁ��������%[�i9Tǭj̬?W�b�)�>��	��%��EZ���r)]���j�����l�t�Y9u����V�[�J�O^S~��/1>�m�1���a|���F��{aӯ��Y�!�3f�&0���g���yi�a7x^��N>dy��R±Q�ι�ŏ���};���+�b��l���_)��8�Ip)�wn�Pڸ�M��[��������z�Y-�V�N���_�o���=�������,��#H������Sr�`����0zʭ:���X[�����>"ʦ'4z�7��$t3Z���g����B7T�Y�>��tȑ0���������d����~��I�Q�5���������ҵ�3���K�����!����h���\x5���c^.�8��קѸ��o-�4y}��JP�+A��`�0.�;�_��z_섊F5۔�]^݋���mD߽1��Q��{�b��媞�-�l�cEG���iG�"vS)�3�� ?�'NQe���]����}A��ǐ�K#�>|Qb��V+�~�>���c��ޯ��X����.����T�WA��ށ��zZe���Wm�#�w�/��X�\t�6����N��=.F����P�=�j��*_�y_
7�����!��!Iʿx����%|��$�C0�j�&�4�M�FQf����&�{����3�X����N�l멼����y���?�2���ieX��lM?3Ny�np��#�� ¡����1#hm�*|���=z�j��@�r������8�J�jMC���"|#����Z�b�W�E��2�	�vB��@i�`���ڊV~�R�#�JΌVu(��N�_�B\6����~m|q�K�;�ڡʝpE����|���>8�RVB``��Y�l3i��^/���^Ը��лZ�X�5�H��4��~S�
UL���&?�齂���?�,�L���8�D뺪�։_�f�����4c�6��89���
hQz�g�?~�m���&]�M��z�tzzH��ۯg�-i�`���
��4��z�L��]t�U��9��#�B�>h���[��ٞ8�ޡK���~��Uf{�>ʗ~�_����D�����&�7�i����t�7�o+��ȡ��j����h�]1N� 8?�I9����+�(%�F��B�}�D�G;=e���Tc�Vɕ���R��K�M�����ug��8��y�l!.\
m�t�RO�R}��,���Y�)(���J�r8��n�������(�{��~P;��+g��ͩ�W��N_N���P���o�.����p9'�bՔPn��/0�n��}��6�Y$����gF�/�&�������1;��=E�Eģ�4�ӵ�*�ͭ���K��*���@%��_ �/�Ơ���h&�7S9#b�m<��!� k�Fsi����msc�!<�x����ŀHY�h��4_����M�v�]� �V�~�Ӆ^?.=��UX�)3� ���y�krz\��Ǣ�2eMTr��­�2Q��D��揅���!eC��+��~I�x�д�|_
o�9��5���S�,�j�}5�иZ���UM�t-�ː�pRuetY�I76}l��R������樫��zv5��hM�=�vLI�E��Zj��]&#eer&A�f3u��?ԏ��ۛ���W�kj1'k�����Ј���,֚�:���ڊA8��&a�k�eUM�5��{R�[~=�N���=:ڜbzS��� �1�\`�h9�ʛ9WO�@�G/p�:'�@�sË'��%�5�#�� ���H#��/��?6*��n>h!�h�6�!���SR���:q/����+C/d�?�8���-Q�/�R�P�4z�iL=�~_���P�O��(�l$s�o�,�Z����f%�u��BX��"O�U�{z�qk�? �� �ey�閭��s���քo����oN�Nf?�#W��xp�3���w'؜ �uӢ���G��y�F���ۭ���z�����9��E�Q89��~y���5
��v]�~f9�~}��r,�/f�21���ߥ��H���m$}AW=_�޳y�TJ#���M	r��n���h�y�,h�5AVE��Ĭ�3Zx���T�~*4�l�I��{����7�L�|XލVѿ���Ӝߓ�C*�9ۋqz����gU/G]��~�%Z�T��}NTߊ*��3�6��Bc��}�Ԭ@Ȉ�H5�J�T~`�sD?z��g�Nܜ��3�f���/�/�:H	(�L��-\ʉ��pfB��*�R�3~u_���H��R��c���Iձ��+X4�D*W���.�����G���g�g�h�m�_o���[N��~�-�U�4�o��喻��"��z���ɥ�8��PX�������v>��/�̟/^U��K�M���/����OO�v+�uv}����Зr�6� V�fо�O��K��^��N[M[_���E-���|%�ܯ
+~f~,��]���DA�X�U�pa�!{[�n}�Ѻ��`�"ɡ��gA+`Vv�j����f�L��/�S#5�LݠH�+���c&�&�58�3
vd�Ci���[�v�3��{��D�D���(;e�X����+ttE�JuF�c�L��37�Ƭ���x<`���~A�Ca�]���+��� >~?!�#�ϼ�.��,�;�wK�6򮀠>���LR�<��şܨ]����4[
x��Cş����\~�]������d/4���م!��z����ۥ���M���"�w������h�a�&�Q�wD���0
R�h�q4�E~�~�?����2����s�Ӹ��J[����"��0Jn:Y/�˿|��h�yRE��w>F_�����I��
����Ξ%H�Լ���Ώ}l���� O��ۂ��^^�Ć-.e!Ž+:ן�/g<�u�,����N'OT"?�xpʲ>��d����&��V�������o��V��2�uo��A��/�>4�փ/�[y~_$τ�x����!�b^���l��Ֆ�6�݅�fn;�pI#~��IK�{��_M��.=>��D�G5~ٯ���c�Q���a�tß��T���
�+��3�Xj�l$8����ܛ�~�W
â�c�O�����$:�,تi%������b����5ӡ�ߖT͞�>�gtP2s�F
L�B+[��Xi�cO���ix��V��UO%4�? ��\�� ����u�Y�=���l�wK�{����A�����㗣'}r��Y-�fX�*:#Jиtz.��(��WR�[�
j�u*{��jݪ���Bn�&g�T��C��{�;f�,��Ω���uD�q6vE���3S �Q�*���/�e(]+�j|��$�{_G�kʃGs-z쓢�1]��\�����_z�o�ˎ1a���m�q1j�.֮�����0בaz�s��4��	ճ��	�^)8��Sݍ[��-+0�g�������>�"��	����U.�+L�f��X���r\ƪ`��:=ϰ}��s�2T*Wy��\�/)�P]����4�Z����}g�͎P�[�^�;Ư�Dl/Z�v���;�����x����C�?�nS��
00W���K��&+����WY� S�U2�*f��w��˟�����l���SJ����n��X�*�	>z��u��mƝ���~@O�rf�A�L0z��>�/F�޴h������ҝY:�!/+_���kR	�]�T��s��,T�h�䉖k��w��cW���G�d�[Z���+��h��#�,�'y���Kw�	~4�#����w��&N~ȹ�L�5l�2�U�@�kC�!�֞�e�y�����&;�}��^�Tʤ�q�tԪ�Ik"p�\�
�{�f�t{�`d�Kj�VJ����_�^�Cw��#;�w����X�BW�h��R��~S�J](խ<����Ӝj)K�14�K��l�||c�֣���W�lRo��Jgcg�|��a�¨�57͇/������tF��(���vzvYM��[��rJC��@���'1qpZ�:�h�
�J�arg�թӪ�^Ǯhd�3Q4�}����^%��M��rQk����X��GRj8��W��Z��)=���G�E�elaIC�o�n艩T�5F�)F4?*���
\7p�[Pը�ɚ��U�:Օ�_8L)����_�cb���r��E�"���{�m�{����.�s|ԭR��*�A��[s���[
UY_;���Qu�z�����s���B� ����B��������� /�I�����M������W^>��pnzQ"hѦ�뮆̉P�lB���nŔ�nW�xkU��5�?_�G|�N������_Ƃ���b4�!�w'���<�M���Y����:����pȯs�����ߪT�Aǽ�{��h�26��G^����'e_�J�
��֊�Ѭ����4��i��Y�o�3�W��a0�eS�S%��C�j��V���D��E�Ll�t:����S��<���������+��U�M�b�/2��<���9�e��-A�O\�����TE����\Tw���rBV(-��/�ߋ��[C�jQ��-��⹒�����ND�j�8�g���W��q��U��N>�����z���x5Fι���ѯ���\h}�2����R`����sQ�݉�C�(�㯘!iG~�)�g73y����_0#��/0v7��TǕ��[W�R5�!�P��ܢ�\�⹩2�RҺZcEw��{[�-�^x�;���K��%K��\3��轒��^�7w!�P(+�jco�y�L4�=��`�A��
�&�n'BU�Q�c"��1���#��$L+y��G��-��o�T�pz��>_�mbZ�~[����s�Z���9T`�2���l�g$�>����z-���Uf�V�??�h��uv���n��YN�a��S�l�ʢa�ʻ&C2ԁ���lm��W���ƃ���(�/-�!�+ġtźF��|A�\΍���f��9�N�v�_y5�A�����{�3@��q/���/�E��c����OB;.�@;�	6st�ӽkΫcD�_�qhKF�Ȩ�����Ώ!Ƀ5q���/Ol�����y��P�Q�g���+}��	�|��'��"l:_��4��4�X��SeM��ۀ�u����K.g�~V+�zڍN��$�
�I���`f-�Q�4�K*d��ޞ/)z�ɳ��ylg����G��S�I����*x�TN4��B��3�'*=1���������0lF�b��w�W.a�����9+7<��Ú�Q(��D�]&�`l����o��=-�W��w$���ޖ>��f.~��QPm��䧥��3��W�о*���-v
)��N�ෟ�#WF馼��H����&e��j��/1%��m �H.
ݵ�U>��3
�=����\w�Z��NO/R�i	'Kve�6��7#��Z�����+z�N�h��h��;�ԅ2�U}lF����֪q@����֪qy�W�>�7=Uܝ!�a�k��o�A`��U���ǩE�m,�D,�j�3�v�i��WՅq�3�o+��ǣ~`�۪.?w|�_΀�I�K��a�����i�L��0z�v�/��;��Yo�.�q���O�/����
�uc,��"�C��`�m���.�i�R��5��_��)�W�;Yz7��XN���e
"W"�z�N�Keav�������E�W�PEŚ�:�E�0;��v����v�َ|�� ���N�zXOp�/�@�6\�o_ǘ��1��G�z[�v���O�lVm)9-I�q��p�8"���{T�!Vy������C;����,�z|W�F�~�Mω��$�����[�x~U���b!��[7�ۃ���7,�u�12�ђ�u3M�x�M��+��M���	8���$kp'�1rDy|�ӹ=<����;W+��N2�v��i�dU�Ԋ�������j;�.��6Z��1{��B5���#��_�,{b��R�)����~���	�"�B��&Z}Vd����	����\D�Kʁ$!!Ć�I
�E��ɠZ���W:��|Qw�k����>],���̓�ѯ$_���Y#"vz�����Ɉ��4�{(��xp<�V�F5N��nY�0X���r'��Ȳ~��~k�X��*�G���ޠ����Ȉ�D��Z+ׅd�_\5+w�����7.U�hգ�C�)X�bQ钣:QT��υQ�e�_�4\�=�^]�w�|�L��hn�~&�2�t
w7�D[5�LaT��Y�R7��d�E�T<�:�ܩ��"�9�|�B�5)/��}�����?�v��ۏ�H����ѥ�tT�GW�WM*�f���8��6?2���v����&Z��*0Z1�՚�0��I�Q���/i�E0�ƞoW�5ś��R�3��K�>�Oj�Ĳ�ʥу�g��~�K�rk7�r��۟�[ �9k���ԟ���]vN�v���+��I��`�h�Qg�����.�~j��K�������3R1:Բ)F���P.U
�5.�މ�G�ޑ���3�$d�O<�R�@;=��Y�H�9ϘVs�.{�����5��}��+�$�Q��K��0��ձ,]�\C�thһ���"��/�Z�-]s�RAYyρ������r��_@(��?�Ar�?�JH�~�c�m�N]�Ѫ |���vڬ���z�:mp;Q�����ײ"�k��j��%�T��FX�4~�P�Zx�m���G�s�r0}��Ƥ�0�?��N���GO#��m�\��,%�ȺH����WaMi��w����xEU�Beu�/���������3~�j�^�����W�!F5�4q*�8x��z5�N�h�`~W�2p^�,Qx�S�H��F���SF�4�4��=�>.�8z�+�x���o���Հ�����%u|��9�����MJϏ��j`w�,�8�����I�͠�9W݋�]a��!7�k�</�����2�������j��aq�+G��r��?�f��:��iXy5t.�f�	f4���lIb�7�v�dWr��R��Ӯ H�FB�7~�s��ֺ_��p/ ����|��<�����x�\��G�*�U���u����R�?��U����7Tvz0��ޫٛQ7UVz�U�n��z^�Ue~R�U�S�kN=�=Pɕoظ��qڅ2wTP��S5��$n�X�r˕�"~�w���"?��X\y���)g.4/ȵ�=+V���z:�wi�"��@I��
��B�x��M/;��YxW����{%��u��xZ����W~<��;j��:L�
�������������5䮥�jݷ�i����	����_�.z�{�gMg��:�a�\����j�rK�r���I�.�Y��M��dJ�F�_*[S��F_�c�f�`�Djs�VWY�R8Ӫ"(Ztz�r���`Q.��-E��S���i���	#f
	�:��؋M��st�M��o�Q�"�>3�gu�����|\���dT��	�
�Kl���e��^{M<����|1	s~}�
�r7����ѿ��۠����6�z �<Z�|�e�~"�SM�fY�aN&�����ZTm��ש�<�"V梬�Э�.DV�
�[&��fܿ mnCI�A`@�<����ذ�Pˎ_�!��^8�O��8��1EO�>���E�:�D������z~J�K@��vL��i-E4��\>��'��8��Ro.�׏7�>Ũ�+���ۀ��գ�gM���|�ڥ'��~_�v*D��[��xV4h����}0�W�R�3�G59����cA�����[i��N��po7%Z��� ���ul���&3QCu�8�r����@�{��9t	���޿g����$� ���l��v�Ǫ��@�e��"����;�¿�4A�A�{�tտ���ȎU
%��g��]�i�A#\��`wA�Yҿ�P�W+�P_uxQH�g�F��B>���5X�l�*M����c|�.�P.]���%�zjG#fo��]5S%M����U�JAk���B��=E�	�Z�8�����U�z7P����u��l�J�v�5Қ�p2Z��Zm����y��1W�D�L�]k5'�~�;Et"�����3U:��;\<��p��X����4�Շ��zj��߾k�H�w�o?��ǐJ�,H�E8+�V�7�8�����+/����@���{9.�,��έ+3���Ø�r.�,�0����s3$�>�/�/+<���x	n��v`�'��켳;0�U��Y܇bXu��V�7=>&�c\F0(U�K=�CB��񮵗Ekź�yq;e3lz�a֖ �����ea�(�n�V�d��Yֈ�r�o�f{���V��VȰ�V���u�L]j�C3ƴ@���-���KU���;�UL���P��Ѫ�C�h���C�P�^	���:�*æ���Y&Cg.���,�a��հ_[c>�#*$@�+�b�q�������UN���a��J���ݕW���-��7�^8�嘍�S W�rX�T����~^(��칬�Cwo*9��4M��w�b�EM���i����1�6N�!.��RD=��ӱ�����'�TQAU)?LWOC�O��������"�m���雩�"�\�NV��S��-S{��&`���b�tH�@8l�P��\k��rxý�̩��)JÙ�������D*u�
��D�Q�`x����-�]�(�x��!�׻&t#�vO����.GG�}��.�TY=��������qz�g��Qْ4��	gG�[�ٿO�9�Q����ə�$7�˘~�%pZ��h���^�_r�{�D�J�������z��f�G~m���:�@���~���8��P��0I�X�H�+p{m�L=��~V��h:ӝ\�R�\�W�߻�X��C9��˃���N�����z�v��/9N�����Z�mF�9��:���?�����_\��Z����ĭ��zrGh�"�	��u��O��UU����1>/�S�@b�������h!�j6} ^KR�vq4����x�����0X��+��z�*��n�G�������[4?l3�������'8�=�U������(F���?���'�3���L��/�Un���OlR��d|�Fgö��U~q�U�����x��
֩��f���J/��Rd�2�"�ZhEU��s��t��G�U��B��'��pUoh�����<�^=N����V4�Џ���H�a�E��rL]:^1��!Ѣ���5�V�L7?��ΎŮ�U��wWg�k5_G��Ӣ���]X�������xL0A�� �v<�t?Q�s�D+�fA%�%�Ö́�wE�'�����?���˞^�s�����
4X�}b%�[���^*GH�M�yH��hK9�Uq8�.��}Ԍ�R�x���y��]�Q]�Z�8?�������R�� $��T�#��Jta/W��5в�;����Z�B+s��i�I��0\�r�
�F�;�o�ڽו]	g48�2G-��[b��h�q����3��f�;�݃�:��ݠ3��>+j3�>�������nRih6�V����ˏ�GI0{T�mW�nE�{�_-�̵���B�n��J�'Ji�����*��.a�/�E��#8��&����?����^6z��%'ګԽ7
9>�fe�?Ɖ�B�QR��T-b����I_�j��k2}����q'xx7<���ev��{��?�vN[4嬷�3�vJ��G�Gu�<ce	X%�Få��L�&u.�5�2�Vb{�P���)/}qN��E�F��i��u�k}�@*P�-��9�#�&�%�;�˧ξ�جge2�g7t��cFǮ�y�~d}�p��g���vl��L�d�3�����G�t�Gk}V('�E��:�I���P�n�WVW��E���QZŽf�G�|��Ej勚=���|NU�/hP�����iߍ�9�������d ��z}�׍N��.�=�1u�zX?;ٺy���e?����w&����O�j-w?ΰ��Ӊ��;����@�s�`s
��u�DL�z���91a��Y6U�6ε����<|Z�{�dk�(ZH�m'��a%���"�+����o���� �m_EV�H^&;�tS1D͎���;(�����WatF{_�O�t�Ew5E�m�Dx~��K	/E͋׼E�_�.Z)�~>�����I�d)�v�u=u��!�,b8��Vx���n��cI��f� W���M���k5M�f.;=_�(�og�M��|$�YO~V�p2�Iuk�Ѫ���^>;Rpƒ���i��ǈGM��HZ ]Kk/s$��,���&3@�_A矇��<In`�vy���T��~�<mk5��(��������,�Kp�q�}��K-��wD�O���G��G�����:��N��1�V\��[�ꖄ�I׭n�鏢���x�O�1"�����p���pJB(�*����sm�R�N8C�|S�_6�O6�/��21o�V/��WGp��"��GL��uw�پ���"���>��P�]r2)�<=�\�$Kj ��<��c�s���*�Jw"���8��F��ٓn��ǃů�r���J��)N�J��n��b%J��u��-O\tn�~#w�j��y.j�Tj6���5:.I��ݵ��k`�4���r���r���OYn��my���s�_(�Y��͍r�y$t��� jo�(��~%Q����������o�l��櫬h�;����N��0a��&ZvUH}	IS�
�r������d�:4�kBj*u��A}�g_��(Z��>m�;�`piq|z��*��/_#k�^V�w��ċb��4ˎ�X�� �_	�J���ICI�����Z�2.o
��+��Ӣ	[<+���}T���+6�)�2�$]�B����m�+[� 览�"��I/P�?��\,;���v3xz��B��?g�ܺ��VEU)u[���@��Ts���_���5��%eѫi�TaE�^�U��VHzܼ����=��<�+�W�u�De����{k�����O2Z]J��^�7����E��v�m�-EY� ��U���A
�z���oj���}]�2q�^ͭ�=+Z���]b~��.)���%�4�������()�7�;:F
�Ul{>��WƜ~�_��.[�`i���98!rrf˳���!��G�.��4�6��{����Z^W]?����A�6d���v��U�L����i؀x�n�#��ؙ�C��9иZ
���*;�̇��鷻�%Q/��CqC�qh-2B�x`X�Bm��/Z!��u׌'H����s�I�᫙'rݱE�4螩�e>���((��x@~�p�}o��_1��Gp�[=D"��}���ɛ�1��m�&����ȅW)�ӣ��_�^}A�}фQN���m�ں��R�6C"z�F1V��N�T���-�v���F��0N*�j3���P���׌L����	���O'{	"*�DUCm����?�,������?g�tE�Äx�~Mz�|o���x����!=�.~5͘��1�w�﫼L_��Z;��Ᾰ��Q�M�N0�#T���H�.�ִ4����[��4�ؐ�s�������4M�ˁcJ����XW��H��+�&rµ��_��JLYd��k-wz�་���G�	��w's�Z��i	�,���.ڔ�`����"*#�6N����e����,�?�N�3Tt��	���Ws?����/�(G���\0�(T����:���l���jX��`=&l%���R�ј<����s;\�緐��?�s�.����:�����������^z��;�.ҏ�N��R���ϴ7
���P���,����>|�Ѧ��uz[-�#�s��=�]���Q��r���}��^��Bg���%pA�_�2�4WUYU��s%� Z�a��o�r�K��[��:#��M�c�Z\0�A%S�%;�*A�K鞴˾8#l��N����~Vr�+*�d�x���D@c�
ҋ����9����o*�,?�[�*2�zJ,�i��>h3�UN�*�.yt�-\��h߶L�P
�>���A	��:'��3~Qn�
��3����a��t������_>oVM&�(!��?��K�g����]4��,��CZ���X1u<��V
�w�06ܿD�Y�R�in�Eg�+���qN���Vr��'�oδs��"jֱ��+����H�%e� ���l;|�S���I��7��#B�n�R#��D�M?����&j�ڕ����f������{��o�^֫&�ļ�R�~ �MD1��gݤ��LVY��=�Hvc�/N��� ��{K>��`�E�������;զ�/��[-�r��ƣ�·<L�����=�Z��o)���m�y��JUB�r�U��ϼ��U�oǪo�$P�I� �S����������ps	9�.:���G՞5�&�7NF@�j}�^IC��yzȰ�¾��e/
��O��G�X[��F����
���t��8���"j^E�(T��w�7�ϙD����f���r�O�X��dTH*�#r��t�)�E�rz��U�~(�����ɴ��������q�{��_����z�*�e��ƕ���?��3���z�-<���K�2ʉ��g�������z����m�:�$�&���I��Bz�KW�"���i��t�B4��q���$�6��?m83��;P���exMD���3�DE�珣�zڭM�I���/��������*�*�]�R��k��GL T��1�DOe�å��x$��o:��/��#/f��	##���!c��c�Z����ϗ�O��1�"V;e���l�t�$@l�U��܉q�����b�X_��-��u�K��	<�˕U����(7� }Ǟ�OS�a\�v�b���R�UX�~x;�b��ڊ�f�M.9����jXP9�"4f��'w��j���Ʉ����O��d�FN�����2�q��K@�Ï��X_r_����!����Zͽ���!��;^�J�3ٔR-2��O�"����QܫF�d�\����ۙ�{��8;݌"(Gv���I��^��%;�+����B'����-r^��@��mlO��t�+L������!��s�X�9��R����L�K{{��j�X��'M�1��(����(P{�N���w8�S����~Pu�os5����Rz|��Dr��;�b�����|��_O�ē��=�Gg}��PP�����e7�2�GR�|"�D��[`L���?��F�qg��/Ժ~U���EV;3��g�n��N��@��Ҡ�T`�v����[W���"TJw�~'�Ĉy��`*�o�Wc�{Z���]�6�e_�<*�ȫE���>����T�6���a�Z'��㻧ٻ�Խo�GTl��#H�q;��ۓ�=��}wl1J�<sm��Hh�S�ϰ����i��p>�*���jٿg�l+�}I�C��[�m��"�H�}�c.�wں�d����&fW����g�k�} [F_�h��X~�vJ;�rf
u�����X�Cm�w�s�B5���D֗D�ĔO����I#����`_�:0Z����Ή�Un\�ve��e�č�%����_ĩg�Do7Z5�"Z��;�G*n�[��M'��oz����+7��	,�F4���6K�&9*��C�}�K_��u7-Zl� �܌g��sX���^��L�"R�������Vm+��)��޿����`�;gS3�m�n]H86�:۩�A�X��ڻ�����9��{r�v�/l��ヤdv7T5_Z�h��f��r���D���<e�{ɑ��j�¾P^̓��ۛ��i�X�����m'�U�����}Be��l�[O6��w[��dvrk 1E�~��F.�8x8�eK{77_��׋��+"�a?$�����jg�;���;����5Vx5�*2��J�ii�([��.�V~�\3�v]��\��]�r`j���ھ�	�������(�[<;A��|_���p�/�Ok[^OF+E���$J���w�[צ�j�]��l1�תEl�t�^`��_��>>|���߿�M��[7��S�8��SO^�T�M/*I�|8���Wʓ��g���T;�LO���قԂ��|1�#7�F�{�EW��WZ)t��qz3=bP`�렮�Y5���;���7�D�lf�J��/��s�	�@c���5�)�7������Vȥ��<V�4<�W�	4c>��^�V�Vy��AI��(S�,6#���=��-����.�T��ݹ�o�{`���5=&⇒B)_�l��I;���~��ʪ��_����H�M�8����Zm�1���4)�Y��(� �D?�lc�}e;��ʺE]�ۇ���ƺ?=Wo�N�e�X�-�Pn��Q�'37W0��N�l8ze���/�Zk4��[�Ot��lؿ��b�O�
��Fk�{WX�u�ʹ�Ov����r�J�aJ���z����ER��T���|����g� �����3}�]I(\Ѿ��E��W��'76�H:��w�1|�ǫ{{1���U�Lu�wRc���I���������U����L�S��q�ׇ��ݔ�^���G`$J��^4F�0_}��*/2-×pDժg���{�~���sY�J��J�T�,pi�>�8'1^l�t��H���Z؊�y�:��4�z���|j��X#�\��N-���i���:5� ���ZO�+�W��1���A����Vۮ��R�]�ҪݴsyT�t��2� ��-]�C�|e��O�hi�$w9��hΪ�[�=�?���D���ӂ��2C]����tR���pG�ݟ"���u��w�X��R���L.AO��,��c�/���@���v�_J%[+�o+]�Y�y�J��������g���jx�S��[=t���)�[ ���>�!T����#e� %�PVŹneok�����~�Y�M�>^��Qm��+��;�?f���R�;����iug�<��д�;k�bm� ��iڙ������ڱ�d_]�z�P�����ܡҭW���*�מG�	 ����(=�����]0��7�Fx�:)��k�cBv5�������׃���Y]af�4� �Z���q������ls#�2љ��&i����{\9ul������Ӗbɉ[D��R�Lv�Q)����s��~��U4�B�B/�?�Hn`���
'�Zd*@�?��\�wk����F=���e#++�C�Vg���#z�����7�ɥ���z�.�]��yiñGO��
��
�?*+ܾ�z�����-�l����eQW���>s绺h�`m���T���ɯ��*d�N_�b�Z�xW�U{ò�o�?������;Ya����b3�5�ҝMm�_ʃ��q�CV5r>�źN�~�lP�N��S]�}̝gO�*��_9��}�͎�!�>|�?3������:%�"z;�1�L����JS���8��M�ƙ>s�r��T2^Y��J��MO����B��㰈gU[U4=S���ʌ���@1��+�A�*˺��S/�^��e��7U��S����d�:Y���_^�_��K<�r�^�:)G�����hb�g�4A����iU/�+���˜��|��?����]��|G�˷GU���*���&�b���@�9LT<�,>���ª]s�J�tN���oj�!��z�����z��URV���o�_���?Y@>̤)�RI�]�)b%��ɧ$l�:o�J��O��[�/g�S�3��X�xm���a��(��ܲ�!�x���,Y��-��$��0*=�[�h�ӂ��/�UAM@��w�g�+M

<F�#N7w����
'�����9U{�l
�Yn��Q��5�
��dF�o���V��F�r��_�oލ}�Lh��;�փ^�0Ն�+-�>����^3g5�)�;_���oʪ}uv��Q�>+��T�9�ؕ��DK�v��G�F��n��$8vh;��
/�GJ�OG���hԟS��[7���'���O��qz�(1XWa���Ǚg��a>���V�a��D	�'ؕ���YG	���Ϩm������q&�|��ak��aܭS�*�կ��_Erp�w�BW˟�ͣ����anRzm�5���r��i�3�����WU�V�8a�q��{�hi��Ƒ⁻>p�\1��-^��uYߧs��w�_���)
������K%�5��5��a.\��:nK<��<V�N?%>�l� zV�wͬ
��Aļ��W)�0�z���@�6��6�h�i���T����Fb}���x�ܧ��n=��</�1������V�`��r���UH�n�%���XE��RS�s����V����I���aۈ�F;z3�aT��J��~�x�����'�X9X��9D�<�w��i���!�ę�y��׆U.���>��0���Y��*l�7{&|�S|�<`y[�S�}Z#�,�������`�s�:OT$�[��<��ў^<�������}
�K����*#t�'��v�w_ş\}��@5A6�Yi<�! ����,A24����k�����X���������Ǵ>�*��^;ϗ�~飆E-Ч-.�pI�[����iΪR�1v��"��EL��̬�'r#�+(��ޮ�m'��W<x{��c�8��>��)������Z>�h���.;��]Їk�Ƣs��@S�Kpi���^���,5N���y©������u[�/n��50E��Ǌ����]��-�TbTw���%#7��S���4E{����S�/N�6���,Է�AK^��=�c���G��"W�<�����k�U b���E*ď����0���V$w�t��3։0�c���A���&���ئ���ϊ������d!�G�b�Ӈ.�Z9c�(�~U�rG��H���i)��	.��7����zh�BK��h��7�E]�2�%�+[G��\���T-�1��Yu�#g8
O�m���^�.�<mD��<�,Wro��<�Hm���Ћ����ĭ=W�w=/b�Πz��W�)Jj2\=��/���bm�����F�Zݯ��/9�
{��*K*j�l����!���4M=�gE���	��h��WY���i�~�~�R�[�0l����x�QS��+���I���*==��( =�����/�d�����C�
�<'g������o���ʱ&�J�}����W���e��"���qJ�%��p�-�r)�Xk��;+�eo�Zv�5���2��a�<���QB/ke:�,�uzT�j]��W �\1�ZƢq�]���w������ �5�o����44��z�/��f
�ʣ�y{R,�ro]2c�WvOo]���h��nDj�|<�U�G�F(`������w�X�|AO.<�S�F)���*�����Xz�����<��#g-Ҿժ$O�Z�H��L�ݤ�R*7���u?=J���/� ��̮��0�ز�V,?�~��d�
�G�N���E����M�tU�����.ˆ�:�V!�h>��{���C�Z����O.�Ezq�c�7fƽ`�M�6z����1PGj�a��s_��W�\2(fr�$<�4U��P)yR}}�7�LOMF�:@��,觙G%G�9��_uM"'+л��i�+�c̵ɂL`�%�����qS?�e%�Z���ᗍ��8�p���b�;*�����C�A�!RR�QWpd��G��|�'1e���!��Γ��-���K]{��dч�"��R���IR��~��g�(W�0غ�}��j�����5�]�"�6��u�1k�Z?P%[]f���	UЋ^<[!h���_�Ct��ڃ�h�
"�>��fȊ��0,W�պ$����
VڒF����V�����m�Ȯ�`~n���=�l9�S������E��6��`�	�W.֖7�]՝j��ԃx`�b�>��_ޮ{��2�W�5\=�_�`��o����3�!O��t.���oA��K9.�rҊ��x���t���8�~���jD����o�����`燯N6z�T���n;Q��e�����{���������M�.�"��!�J�*ߩ��Gg��^3Vt�nqQ��']\eZ!��t:8+Ѵ3�J����i����\�Ʒ�����|�`��=Pl����� \�|&�ǟ󎦛��'ˢl�j�pʥ��6Zش����E��HiY�?%�Gk�+f}8�]M��=m/��fh�V�U#y̖M�"=z:p��bI�9�]��cq�)v��.���7�Ņ/�V����"ӷ�o�m:�8=�&�B��Ĳ�d'�5�u~��گ�-u[�j�L]z*3���3����I���ஜs�i�~��Gc�6;���~>&/�ɟ�>V�!����6�3J.�Ta�Zًe�`}���o���,���R�~z��_W�+9Eբ�|s<j;�|�r���ʅ��i�(-�$�i)&h_�.�4��2��)Z���ϴ	�f�)�U�*U.)q�~�dV���k7r]����KS^�W-�7Z�����=R�YOoڲ!�SM'��狠x�j!�+��#�}�O�,�+���8��w�X�u�ӿ��\�F/�n���q��!�1\�އ�\}����N/|#�.ۏ�,�x�ZFK������d]I�ْϗ����k�������C�?,���kO���;����/���@.W�Ά��(���p�wv!k�溺9)s�� �6��U0Au~�M�v���yx�q�;�Q?3�`����Q��7�.�PĊ+������?��K�-��
�˴���hS�������}#�g뽊P�I�]�lʻ
�a��u�[�ɛ�S�ɭ
�}~��ܮ�Th9_�P�݇+��z���˕BT��/�񣵆=q����_���
(�g���/�,̇_T�<����#K�E;U%1����U
�;{}W ,e�&�[�A5N�����%��v�:-� �sz��������_���T��j\}��`5��]+ت?Q�;������J6u��:��<B��{�پ᫸Ri ����l<0�!Q�%7��=����3y]��8��MU~��."M"��Xu�1��ܑ��D�>��-7�Ŗ�R>��d�� '�E���;2��oB^͝�*���wt�����8k)i�m3�?0(R��~���>�1>�����ez��]�5�d�u��.jG�^-^��G8,��Re��~`�(�<T����}��R�n�LН{�*?��[��ߪ:��j^ue��oͧ�'����K
�=�GU��z�|8]��}�onL�	�O�.�*��v��J��+E�J^��O�V��� ��\ffB4� ��&+�i��u����U�#�n�(�&}��Vp��B|�O�����k�}|Y�
%�64X/��|=�[Qq��SBⴓУe�(4��~7hV�߾Z���i���N����XX��-�Rcɚ�vFT^*�R�_�4nq��v�D]�W�
�/�:���oa�O��o���m�.hg����63�ʦ�m����	H�R��S�ˤ�&>��a��;����M���*%�{w���9+��yX�Tr?����b.��)m�XK˂=���<�>�>�(:�W龘/�����AF��$+.�fY�I@��PqB�K������E�[˶;܍��0R.۸���U?��Lۉg��/�N��.^T���7Es���O�mwAL���J���*��Υ��&m�hZ���(��>ZV��4	��<������r/���9e^�(�-�NPo���2�[�7z�!�Y�G~G��Hm\�m]�+��Hkչ��GR�ۺ����߱@�I��m�l{=^�>�n�ʹ�<��|��M���Pj���˼I��0`t7�p~��{�{VΫ8ER&'<|ၵ��:����wۡ'‶D�&�����:�k�}E������U؛�������^r�_쒉�"ySɲ��9Wy��??����}A�����ٗ|�Z}�#i�ωwd�еCQ���:-�w>|�����Ҫ}���?\�?UW껃;BP�^+֕�����ѓ�4.�e�^���(�[a�:�^�ffT������s��hVxK�mX�K��v��^��f-�=C_���P5��s�X�#H���7!�G8���f��6�;��_�D�-$SR���u�ue����W/����Pbz�2=���gigU����k��#-���{`�D.�������O~٦��ZE>�����J[7�``���^�`�|c�ޞF �~�k5�ۈ�����+��i�ĭ��������3yczW�)�2kT��bϨ\g�,ް�y!8Z��m�����	�W9��բ{EZ��I�W}��$
���1�]��t[��&��U*��.,�Le�`��>S�D�g��}��˝�E+z��z�l2����p`��W+��圻��e���]�����s�6�n���l����iP�ih�f5�=���_Q�2=�ȷ���WH�{��dg��d,�t��p��Uب�*�<��D
��s�^�fN��n��;?k7B���R�N�
nA|���KR�f��A�������g���d��H�Q��]ᮽ���5�����Z�.��j[�!G�Ϥұj��Y?��DC��8�'~��Dt���)���,�4%�R�����/�򛞡M��3�Ҧ>�/Yʺ�ԯ�r*����X��a�eȪ2��I���ź��E3�(���+���O8��L(.�;���t���nX��r
e���e�
�V��e�ʡ)�.�v���0Z?���������'=���j���
�W�է����F��lɄ���9�>�gw�|�R�����
�� L����Bٺ�/$�X_�{�������_�+Z��./��G�P5Є���͑jm�͊��)��%��QM �#��sv]�^���N��`�S�U#UD��Ź
�Z�4�?ݝ6<P�	__'�����/hH/�7�ܤ��+~�Ϊ{�X�k��sYi������oU>����T�����.G�Ey�B�����B�h�2�ː�G(U	V/��w�5�\����lnm�+Cr7�|�o��w��M�C�+�MKd���(��e�z幭�/�zV=��-Y���[f�Ģ������DY\z�2w�����}�D�H�L/���zo�g��|�[a��W�?kn�ehU�Ey�6�SA�K�J\�vиN�e]<�+�J��1����_+ٶZ��N$B�6o�Y���^.��}��ʇu���R��,?:2���L�*�v��;��0��Wn�+��n1��n1�:�V+�/��~��b���=�pX����,3�'F�����`��1�M�}�=!{�O�}����@���}��}��0黸������|rڽ���F���5"uo�⍻�^V�*m{�R��Uo�mgu���e��j����݉Qf��?-��+�&A��L*�UR>�g�;�!���睛mO���~��E=�a�yu�f=��B~]SG+�=�(D�>���/�+bu9�9Ӈ>X}��~e�v4L�/j��Ns�r�h=[�i\0V
�E��d뉝"uډ�i>Sc�
�4���U��ɧz�1֑M̬���Rz���2)�/ZiWg\��*"B{%�2z�L�1qp/�_%UƩR[�)S}�~�Ŝkߞt���u̷t���ar~e7������V��
�~WT�Q�7.��1F,ǭ.�QO����`Uu����o�O7�%O>�]��3Q�1e�O9Y�E֤�<!�U�j�hu�I�T�P���r7W�}�8�o1��E(���xIc�8B1�hͫ���^<?4�%��F��Z��A�K���/o�k#{�r{)i5@W.�I��mX�-븮*���5{� $}`���'դ��݂a"rT�Q�:���ER�^�r<��7��}
���I�"%ϟ��$u�.��_��U��������Fl�=N|'3�+�g���p2-Nk�d�wl�u���рP���Kh�OO�6�qv�5������`C�s������j��tw��Z�)d�6<8�	��_/���@0S<@��^ʩ�^��|��.IgAO�Z�+)��;����}�� X�{�P)o�Jnu����ҟs�d�U8�`���ݔ2�{����-ԿQ���G�����`�1���fNUhT�5.���kd�Z�Ĵ ��z]���ҫ7WK9]㓠S�(�յ��P��q��o�T\��_/r�v-��k H�@�%<*�J�X�W�$�,j<�/R�nӗ97}g���
�u�F�{#8+�vu��j��ƙ52@���:�ו'ߖ%ҫ��4c���f��n#U��	jn�4X��P��L��^m�B}��G3=L�	��:F��"���rWl��6K�T�Z	��X{|����
k�)�/��@�Sඖ�g+<d+�����ggJD�r��!�^ï������0Z�v�Ǩ��2��q�F����_��4X�I����X�V%o�.I�ē��E�P�K%)i2=�5W.h����^������9_���]�v�j"���aڻ�0�ry�X�$��m������Ym����o=��2S���@ڰ�R�MRrm̽���%� A7
�m"R�C���hT�:%z�����i����L�B5z*���w��&NП�0��r��(�(�������%&89dQ]%Io�j��H���o�ʃ*���J��HB�nCꗿo|�������`�]J�PW���\:��;��Q�|NJt����T���\�����I5=��d�r���vz���U����C�3S̚�u������}�3>�)I�D�Ϊ9�̩N�ӓ�_�+�l�����PtZ�K���T$�b/Kׄ X�wz�8FV%[�=l@m�K��55<oM�_g�o�_)�+�km�FX������wK{Ve����,��=X�TD˒"Ǖ�dD��<PS��Sut�^W�E�_}��:ã�te�R@�9r�N?��f'T�D�1L8��.��*��tO ��g�u#0:���٢z�E��D|i�M��|2���4ß�p�P�[mV������KVf��H'\�haLU������]IS�hܾ�{�^5�%Te[�#���5L=�w�q����d8E�l����>r���1k=�R�ʰy �.��ɯ��Z:�a~����*�4_&�b$��T�7^�N����vsR�c�*���j6�uV�o��޷e���hU���׸�SGȢ�wb���^����;1���K�~��S�œ���O�Z/��S�a����+;�/���1z#�Xw�́j+�(��,N`EV�*��e�Q�yw��� P������:�&-�V�#t��zO�XiAo.��qz�Z��S~��#�bF���?�ϙ��|�MG�e�n�+k^�7�] ��:=�7�/ú�+˃���C����3�Wq<��`��5�VKZ��=�ۇ���Z��n`���!�eW��k�_%a�]��|օ�e�����wR?�,y~6j�K���XW�T��.���W�g��/�����v��ge��9��}������ �^9�����KJ�%�]?>�TǦݕE���"�!b�I���ci�mŴ��q����-`?�c��G/�hN��a8y�u�?�k�_����cy��Qn�Et���hл;�\�V8�R�#CQW��u��W~7���ⅲ���?�[��Ϲ��]$����gƶ�E&��{�.ī�z(�B�=;��Zr�Ϋ����J Z�}D.��`<é|q��%����z�nn��eJ�t8v6>-���Pq��`�k."�M�}�)o�A�����Tm�����)����Q�UO� G���J�e�`��9��+����9.SGH^7S;��5�}�I�|6;b|L�^����j֙���F�������@m���d��O�Tr�p�9w�hG�|-jrG��h)��:LB7ϴ�M�(��E�D�2�z�A|8��s�5������M��"��F�ֈ���W-��
?݌�朙>�rb��7ݭ�|�r�ue����>��+�k^u�+}!P�"n����N���+�梊�Q������7�W�+պ`Ɩ.z%޿�:L�|�A�x9	H�(�������wr{��Qju�+wi�����`]�Cb�q~���2O>N��a�.��*/��&Zc~���!�E	z�����y��Ul%��}vn1oe��'ryS�Pp H=�|Lݥ+S�R��P�Z�Q���jj\��¶S��U�\���BJma�ѕJ��Uh���` �wz�p�%�^'��Y��=�S��y�p�R�TY�t�GZ�S([��$w�6�R~}�Jk���sw��JYy���t�o��*����
��Ak�*���4�� �����V����I<o�V�Rڝ${)��ܪKy�[���:�X�Y�sg�o������X���u�Fۭ��;���X��zgY[ �x��h�r�:8m���O������g����y��׸����P��8�%��b�ոn�C��]N�V��I5�p���\�^
��]�f.EKz�F�e5�gv��6���;B�2��-�/�D���N�Y;_J������:�Q5��o�ֲJ�35���ǍX���1`��\5���_i�y�dЉB�Ka#q\�<�ʪ̮�}-w��lG�f<eT<��,U��OT����h��S��R���b�9t���w�x����W����7��ʶ��&~��|a��G��f��0ԯ����@b}�����.d�v��{��~֊��ImtV����նB��{q]kB6ÄNz���m�z�H~�_��j�gU�%׏�\�����Yn�i����"�)h�w������������^i�@+���Q�����m�4_(���75� ઞ�/��*X�:+7�l�%��X��3����?�r��0�.�YcHU.�O��FKR�QEc�"�7�1�)�h;2��[ZZW����>+QS���{������?�a"{�-��:9�O�|p�z�O�rNk-<��b�y��~��_��/>%�M���򑒖��O�WE���WD#,PL���<,��������fMr�W"���3Q>�|Zi�C�\�?S�,�f�j�RiF�A��練�r���*��7��t�̳\��ls�P5��>4��t)ݘ����X��n�)�g��Z(��q�u�Q�0��V��Jhf����$����R��1e��NB�����m��]�aEk�3JCV��CW�d<ժ���7=�太:T�p@����nW���Sx�!��ѻٌV�._�"N���6��������FDp)���(��j����>�w���gz��$f��s����<�$��F%�}9�0C=���p:�e�~���o��ud��u� ��پ��h��{��}��en�4��{r�kz������~.��Ö���]mCj��	�>��%��-���o��o���z��+5���7�\OM�����g�|e�<s�ׄa�2��R��e8iORN���.�l�t��Ӌ����.NT��K�;"B�i�l�	#	�}�XZ�kT�A�)����L���ʯ�i�-�륜N�W�0/i�	_�D���ov�n�/U���?�B�_�E8����9��PҌ��aXP�/�#p�Gf���ԇ�e�~�3ܑUAy	6TJjDa�����;A�MiΧ8�f��=�'�w/u4g�ڦ�_��>]��/��$m+f�4SIb^L�����OX�k�dIEg��W�+�[�Jf��9����2n����7�ϵv�n?���g
K����_�a��+�8�t�U�%��hdN�1=U�3T��R��E����- ���=k�M����ꖮǱ��ޯ�U��2��Tz�z�Ҋ1���)w3�ׇG(X8^��R-za��<F��L��ί�nK�~��(3RdǼ�#���5{��Z��sBEr��Uqr�D�by$�����*=p�:��.B���by�FO��>����r��]Q����IY1\���"V�B_	�{�	����	�&�t��.��$���
.�V7]$����P?ɹ�N2Ue��?�E�����+�xp�ЧM{FclW�(���Ȋ9R����%�*�RDu;�:�W�U����1�բW%mؘ�?�E�2C�u�ϧ-��ڙ$+��yd�tͨl77�J���GO&�m=+Âˉ����<
�=��P�ڍ;]y�T_�`~$��Y�񬡧ךt�@��UT�M�ŔɯzP1tj;��W�I��������u�B,�s����w�hL��U#�K%��t�|�XW6h&Uy�C�p�x�3{��0����v>:o�s.(ܭ� �\3�*�k������2D�]JƸVNi��]b��Q�^͛��ǥ	A���Rg�s�A���Go*���V�����u���=�o�t�qsD>8+g��$�����~E�YE�?�L�>{�j/���a���ٵ�q��{�Zf�v�RΏ�ae ��[�t�h����b�e�\���������e���J5���]��S���(&�B����+r�Q ~�f�{3����+1�6�]T���G;%Z]IFO/���hh�7n��bN�&��֙���Z[I�sR�R�WH���zඨ�K�B� ������sȢ]��2M�G���֪�^�@�'!2���D����;7%_�߂�	��w�H	}v�^�sŮ��;���ϸ����*�y{�S ��i���յNL�����XXE��r�#m��B�zvE��iDW�_=8B�e��U�˙l1|�z��3��D�6��`ۘ�{g�J]O�(̅����ґ���.��i|S��Ev�Tp��c��wԉ.$O'=Z���4^Fř2�H��5�ko����ǋT�������j�N_PS^������%*�����H/��;���j�ިŞ*룘�|�_�2��n�gM�/�q|�^�����8<8�u���~`2D��(�ft��Wޕ�qD�}��&���az�#A�Nzҵ`#&��gkPQ�%X�{ݠ����p!�^����ʤ�v�*i��ݜz�~��u������DGN��t�Wq�k�h�\K��'������{��Fd������m���#;�tQ�GO8~�kYq�P2W��S��ղ�R�	�j��*��B�5��g��u���y��N�f۹�d�/Uv��z��r�>;��ۻ"��&7�ս��-��U��Q���	�8�������e��-��ǔ/}'V9���,5�<��7�l�'l^h�*�Q�&6@��T�`�k<��oh�%�*�_&>�˟g�7��ϊ���.0%=�]l{��xs�W��>"��ui�����-RA�_��z=b���>x�����
/�LX���<~T���G+՜t�I�b��No�3�p�����Δ<�L/�wMx�=�a��+��m/����o�����ha�M�M<w�G�9#pMP�#��5Gz����]VR���t�ŧ��P��p�V����!�0�ӻ����V;IU�~h?�i�aI��6���i��h�bՖӾCct&�ZVg"�*ޫ&����6n��,��î��_�'�;�,&r��U��gkUnެL���3�zR�K�
��x�V�|z�{6�o��\(T���9��u316�Y��E����^��|�m�#N��;����Q�/A��C�Lj��\u�7��R�*M����z�s�A'�uν^���gg��6�_��=z����tE��SZR5��� ��n�BB�j=R�lJu<,oiŃy&�D��0��U$ӫ���DN���^]\���+A�Jq��Ҩ&2�h^U$�q���_��/�a%씟f��݀̧�}��||�C��s�Q}�ь��U㲸p���ŋ�rL��@�?��n�b�+m6��rv�꒖�ѫ�ǝ?��9Mu�Hq�,��9ubb���W�t�d��H�oG�`�X��ŭ��}DK{��BU�P���,~�C���{�k�7".pQ��c���,��ْ�b�����`ޢ$8BT���WLLy����3�^�A�"Zw�ō�DX|�1R\�T�94d����>��[��S�_��V��I>�֯�x=7{��p��;}�.w��fg)tJ6��Z�q6���h����ڟ��Zh�B����	��
JoU�ɴZ�gkF5Ġ�����tu1�ɦߊ�cW׼�g����O��u���Sd� ~p��n��1I�%b��I��_	}����L
5QK��l���~�L��/��L���a`�����d������xR�sd��ϣ@v���(�W�k~��r9���d�}9=E&#�bG���;!��'(�u3u���W��n
��Z�4�5��w
��p�K�G;�5��9�&"�|`I���:g�_讣D��6��
�z�+��G���٨�M�y]"��h3�W06(Gv����c�vOy1�Z?~��4��|�]�z*5l6����ج �w��O���k��z��hQ���#�l���R�C�1$l���֭���dP7�C����~߭�ޣ��\���k9��7 8P�P�v�M ������o�\�7҅M�]�E�]N(b�e�<�[�M�	8���� �Y������V*�����+��K�(�^�-U�2�����XO��+���o�O_��H��.��e�z�����e�p��Z�ڍ[�4�Rp�YJ���]�t��
��-@���K�2�W�&�w�Е�Q��Pp%�N�v災�}�lK��<�����az����q�w>��� ��e��0|ܺ��I������������e�߻�8�F�VK���d���mλ�+:C���>s�;�[(�&<��rj=�3����!->H����}1Z�r�6�^M�����T�Y��O�/��XL�G�������w�Ke�	|rHǯr�]�;�V�[�V�;Ln���'�y�Vk�<���yGU�>��%�V���.5*��94λ:�7h�2�c���Rtz���/}TV���u����ֲʶ
�Y�a�6JpbrP�5�[�~�qr�
	��O��R��)fy��;��~�e�!A٠Ǭ��_����o��BR-U&	v�W�
��p���KL�r�՜_�{?�������k'H����ϩGE�O�͛�*߰Y��r{�ԅ^�1f(�N�0�� f�w���ݞ6Z�����aH�ű���,~�_v�K��*TgJ2�|߄��P�P����!GG6���K%A
��h��7
B&��;\w�r]�!����h��h"kG;��^e��EQV�	����e�Z�^�sسatE����D ��f
�U�F���T�M)e[`��Y�D���ϼ�!8_AO��^�ȵ�O����1R��[{��R��*M�+P"����%|�"t��`�ƲuhK[~�
�'R��>է���{�^��S���o,lW��2�����m�~�.(&
��I�V���q��v���ջ�ׁ�M0䲶�P5��|�����x�WLi��2�E�	WY�(��L�>���Ry��E�Y���G�b}`�b���kI��c\�l�._=�� �0�!fH=���[Z;&�e\�e�}�Ĭ��S)J��$��T3O��3�$����\�3�o�+��W�\WF��^~�����-B��8�F���@&����s+�bs����qP�-I�1��m�]T �^2���Y�3�W��Ee�+�_��GP�9(�bx*�T�����������%��}(m�1+y,Ue^��Q	��r$:����09���8<����`�zU!�]�{&D�5GIsH'�\U�*�B�?��d�é�Ԁ�QZ�j��d��r�>���Ͱt-�hU^^9f�`�%�O�(��S����3[34�q�kE�����P./��!lF�$�VZ��S���٪顅$��`���]��������ܺ֏���e;����nlTx��|�;��Gdx�(h- ޝ���n6Q����u�R�/���g�8��z<��	�ުR�tϪ��_3��5l^���V>��q�e���]��iu�z��[:ۇ����j÷��~u���Wy�_����lie�\��_h��jh��'J/(��f���Č�JW�_u���y�d8!�˯��Ph���*�� �@�!)v��p�<0V;��,!�u!�4��_��^��m�=�	��������U���E�޲fd�>담]2[�d��~~�����{`�QB.j����%�\]��"�w���m>�W�O�>il�Ll{���i�P?|H���~%��f7g��,�~�Ȍh��
[�d#V�D�*ʰt2��M�=�n2�czs�G�~�ۯT���D�����[o�o���˧���_�F�H2o��أko$��Cѷ��.u-��;�b��jqu3�\��Gy"�o�o�7�^/&�'�7�C��x���:�5�����FU����w��D����0�����ud��[@ֈ��_���;�O|K��	JO���
h�'S'�<z����eߜrgg�W�iW���*��$��F4��Mt_�)-oO���U�+�Z=:�EE���d_V׀䎀�n�}ǙC�2�L�L8��@��6GRλ��T��[�zƉN�E�81��ml������P� ��٣LsD�FS��j9�������M�no�lQR�2��%��<ݿ�魛^�<����]�h�~�7Ⅱ��m��7E�*%� �����j/�S��Ȩ�UE�b�'a�BK�?Q���̬�c�.٩��v�.�hA���� _"=�����W���F[v�����b�v�V�����V�P^��S+��Bn<���_��e2'�5�V*�B�n^�nz�D����63��O���nT7Rf{�
,O5������2Nᖸ�l�vA��H~`�Q~�I��h	��j2����	<�R_�yi6���@�2���)�Bͪ�Ð�	�nUӗt�[��2�6�:�i��乼����m�˪�؛^8|�?~=�/���Cԥ� �.�=v3.q�7u<�+��|�τ�rYk���!�( �;��)�c~?�)�M4�a;�U��gyO}��N��1����������$�F���1t�-� �3-������|,S�;�Z}&*=�n��(u�R�����=�Z�������*��˒�+��Z�-EH	�~����bS��V5Z^2�5��B�^�s�zF�t�%��-O9�cc�h�ߊT�^�E�S�`(�<��p����9���'j�s4c/q����*λ9ڙZ���)~�@���2�?hL1�ը��ྸtNj�W�<~��++�w���é�k~-Z�A%s���9���˴ßR�C	��� �(Ls�иҽf����
3��d�L/ �$�K�ƾ��~w۸J���3�o����i�����l�j�ż?����ԺJ�A��OIh��R����:V�@V ��R�P0���a3f��퐟ə�C��L���W������YH}Xm�/���%]���j�^���|��^�
	4�nZ.�|E4�JΡ'��Q�l�� �*�xV-�72��g�������a���M�.�s1��њ��nu	?��L,r6nG��Hq{{��r{GXs��W�ngD��JΫ��t]�p���x�]��n\��y��S���%t
�9ߺ�(�
v�c\~|�V�����6�.�`/sG�7غ�ZQ���O/u��|zZ�W�ܿ'Zʵ�u:Ag��#��8��ؿ���-�˿�KM���Ц�%���盲���Ӕ�Ndh�7��9Bu�޸<�{`w6����h��d��<0u?Sb8K�z��a�'g�d�t�g�o�%�~�O�y���ʵ�e��s$��1����I岳_�
6݌���*{�*���m /�?�Ӛ-^}������O����-���&_�v���^���A�ڝV����,��R�ʏ�_io��"ɮVf�}[?�oQW��;k�5x�>|'��w]?��h	TU漶[�X��n��� r��_D��o!VT��6L���_���{nP��R����}��≞F��?���tE%k�Z�h�:}x��_`�����X?��TIm����2�1�b��v��=tq�ek��K���
oի���@%�����p�n}�F{��J�@{zl�'Z�j;��~���q���
���m�d��#v.�;f
����jZLA���+_�
��z�,)V^��?ߓ�_楻��^�\�Kۜ����6����n�3�}, YW.�W�>��~o��o�Qs�0�I�mU3�iޒkԹY����qfp��g���B�5�n>�M�W�п�hϢ7l�w���5*��z}��}3�\�A�j<R�cΐ��rb{/[��/�A����,�����A_�^�19R�f�<��TF��Hy۝^eʎU�Ϳ��I8�+�v�Q)E��S�3��@�Cx�He��RɼC����I���:[�f��EDR�c���k�p}�6K��UK)�m�F�z�H*D��3����7�f��_,8����
Z�t����t��拙йI�y?쮜[��Xҫ�~�U�8�Uw�$���EaZ��Y;N=����1=SE�;Jh�J��}�#�ɨo��U��*T�ݏ���n{u W��r��d_,��Ը#<�[��~��R�'>���W�I�P
�)��b�������b��"1mx �E�iR�	p��T$���Q��oy	.���j!��
4� �w�����(�������� 8�h�%��M�D��?�.T�'�\�� QC�o�0�V�]a�L�n� k��^�\6�y���pbؗ��;�"N���D�e!VBT(�Ȓ-��	x�b�A��̈́��C�+@���(I��@�w�B��Q�@�D�
$�ӿ��C��(�@�A  �}��锯����є�?��y��D8-��D�X���5����/�6@-����-��<BF�����������s��?�W�ǘh�^��$��7Υ�J��fz���$�6́>\��ؓ%?ॾ��R�Nu�Ί��'J����U��x�8)dvO�/F���m?
�̃� �u���1�r'�U�z�[�������5�$�v��!m��&�1�����B[Ib*zYX�AD@��DU��&rm�'f����Nd]���~Q'M��f�:f�I�@|��J @'ʞ�,?���k g�~ !�]]$Qp�MK�_k�/�T�����hnܲ�I�k��P8~p���p-���6�-�#S���[B.�~q�6Sjʲ�FN���K�o$IE��Y�ᡝcҬm��#���� I3�kQ�m(��SR��%�Ui(��yןដ�_�Gn^'�̌jC/`Nnz�' 8�zj��]��,�wU�o�1���#O$��Ŗ�#�,����^���M���cJ�Hqg�쵋�P�&|�Y���P�Tto0r��e;Q
�A,����/#�5�&���C�����N��q�����_tqڶ:��z�D�Y���(}k~�+�D�|�|^�h��n�cs��G�e;F� ��dOoho$L�U�[� Iv~���%�^y�TL�6�\J�:�s���<���ر��D8�v�
�BJ�MU�풚I�E,�tY�s�4��,t���8�^8�S��h�t5T��{[��1��݆���Ɨ��Л��&�vO!�O��s�T���Hx�=�<�4^�Ç2�?]k� ��8���i���/xU�`_{�������7�-#�αR�}�H�C��N�ΫB�9�
[�xf�1�sz�������>qBI� B�j�S����C����a띔N��W�Pu�ց�HƢl��O�Y�Q�.�/jz4�pz�6����zC9F'�k����ⰑCϟp�;?��6d��&���}A�A�g@%��R�w�ԘIi�5�-%KW��x7<s�[j���2�%Gbx�/���M?�:��6c��J8gNw��
�̽.���~�yAI%���p�da������������x�R�+���'� f�.~��hVc��0<���X'	�N/�r?3)fʱ��X х�<�.��1�P*�~	�n�������"X�ץ��U9N��"�� 2$`H!6�ˎ(3����;�~}�<����M�U(�xp.eN<�b�c��y�!��F�q�!s��zC�� �*�3�ё�w�O	K���֥{�5���V�W4�z;�g��R>�GDU�OjKoϺ��a���$�A]�|	��̻G�7A:e�����r�~��2ЃC�'�=�E�!�ҩ�!��T�[��)Z�k�(��D#��~��c�=]ʶ�Y_>�����o8��B]m}o����k�h[>䛶/r������[t.�	�;�Q�����BU�Z��S�aL��𞖣���V�>�hS�G��*�F:Z����0��(�n
5��Rf�s��%��m�� L��#Y���5��r
w�%�����{��F�}!�]���;_U�o�_��	���#O#@>�l��d�[2ˍ����K�p)�2��a���0��*��Tq?R�kإE�!���h��`�S��j����C��F^L�$%�$���R��Y�U�7B�7Rc3���B.��ƽ����b�d�&�5�t͢f�
@���k��'Lw� ����?�ʃ ���ͷ&�6ݺ���.Y}<�rjӰ���b1���w�q�C���*pG��y�Ѻ�ۡ���grB�>��G"��R�[�������烞��~|H`8����T�w��iR����\�<?v�S�|����h�#<p���"��
l�%��������4x�uY9>�v��zJ�S+Gs��&�^.�2�,\9i���t�W���z��B�	 :�>� �2�e?�� q�u�$�,T	B��Bd/�{�5�O��ϷӟF�)��D	��F.�B�I�Y���("|u�@6��RP{�+�^���[�܌Y:�{�&�c�ՠ:������;��'Z� �ʩ�-�k"D��&pY���8W���j z9_��$�C�a-����(z�~�3��u��{_��d�Y��E�c82ȏ$ Z��Og�:�b�̶�W#*#���44.��F�E�K��q�s�[Էx�oߑ'��h�)2[̤Kܬ�?�(@��(Y�F Fx������3������99�:��Z�њ3)}������l�o�m�&�a�	:��߆\���I�/��?�Os�[XǞ�m����/Q�������e��	��#t(��TЇ�r�\w���g�������̠\,�0�����^��ha'��tg�5f�/`��Ai�?��3Pu@m�x���#}�;0p����?	0G�4C��	`�dj	�w��(�'o��:X��t�0�����:h����~&�~w�E`@��xuAQ	�s�3"�&��T/Ţ������g�_���zqx�q�9z~Eb���
�y�#O�w�\�[=����B�9Q�q� ���nB�}�j��Ew�����qh�n�;��M����"��h��"t"��8���Y���]���nL_�QR�xj"�{����\��ү���T<H����Y��XLi��ɓ�sP!�-�P$�s!:)�G-��P�i��+�l���K"�cK���`7�q��L-ԗM��P����H)$���F�w�{0֏�����h-�i�k3�����#k��L���$�������]�gB狱'��Q� �LX�����A�0����m ��E&W&<�J�G>�XO��S��&P�/����9��V�P���1N]r���k!| '�^�x]\Oz���6s8Z����oX�K6S,��-��%��d�M�M^�i�X+,���hQ_6̙����?̅�e����Wp����� �\Y.�?5֟��MEm���hH!�x�t����$th��C�����j���"km�����#�nx �0!7�l��s����;ɂA!4	��R/�W�Ca,9�#[�#�U ��44���ޕ�!L�j�M�xe�8x�Ye�Xr�%�4;bsO�{���@���h�+|C|�J�t4�F���R; c�	��������p������5VFr�/M��K�6�Riu�FB$?�XÐ����R���~�INjr"6\��$q��o����G~��.�f��،�nM~t/E�D+��?�,X�K;gX�˱�Et'-���'��5K���T�o��kb��k�y�*'���a��y�����+f��ZXjd����u��Z���O48[V3��}�/�K�7q�߁#/��뾤�X�]����{g�(�K�=$K)=b޸
0M�z����)Z'�H�j;[]�q�HmrA��5➑��W����S�b/G��w�9�$�n�)N���������B��ս�`��ؑ4�ybxH|�Hdm�=��,������0�\���)An���i�1��.dR J�[�,�5#�8�B�
>�qp���A)�BD$�T��NV&�2�v��=��My�����AXg�-�e�{�q���D�J�at�k#V�
�'}FTg<e�o�P攲�@/����\R�����rZʈ��l���j*lL���
�#���pU)`��#7��
��GN�ɿ�~H+���wY�o��8�6��)<�a�0G
�ԥ��)weȁ!C��YL��m�9'	 ��d���!I��l�N�˥ˤ�����Q�kIw@�3H��t�?�M��ءLϗ�S����'r����\�t|���J�
��R\�y&V��߰�����;�n�t��b���{U1‷�l��9ϟ�)I�R ��W�E� ��ma�t�t6�u�xTݨ�ל5��&ǂA� �'�۷� #R�a��^O����0�7�$S��Q�~A)/h���{=�Ub�v��r�%W���Bļ��uɗ'MnQN�:��C��g����+�<��͆Ҡ���#�w�� ���u�я�s��n���H�bۮ��[��>�ԗaI(G�c��
��h�d����H/֒Ÿq�V�Ծ����)2YIO�+�o��^��R`A��p�ڝ��\s�d�a����Pn�"��rqA��7�1�z�#���jXK�n��̦�mv�S\�B;|������1k'J(������6���^E>*b	��7r:-]��d�m�B�̋��༩	���r��6Uj%�U����)�H��V[��6��r����G.���g��êʊ�����m�Gd1���|�{Կ�})�}��`g �s�L0Z�� �cCօ4g�Y, t���[�(�st5w�	�+����4�1mNr(�O>:���hl�C����0�Z&�D��˰���Ra�4���&j�%n�jk�@*���B�N� ��ǀ�;��9B�'���}��8�/�.Y�)k�+�;n�Wt()�c	׌��	t�ߴ�Z��264��b!57�Z,e��%Ym׏Ŭ�:�s1����k�f�JL�7&���-��3��f|��)!�����ȸ��7�Ӂ�τ�����4`�s�湟�a0�A�i&T�N�'{��\!����8Bc�ÿN�#%Dm�7� ��Y�����.	c۴�$'�7���6Pz�}�o���b�֜��E���9��s3�o:9�E[d���_��E��r�����7��lC��zߛ��>��uQ�9�eA£bO����a7��R�q����gs�\�z؃���Q�5���8٘��ȗ�Yv��	��v\6Ex�R
R�J���ʋ�P�;<i��-@Z�*'2č�h C�d	�R����]�h�{dm�e��7b��*-��Ε�l�ũaJKǽye돞�FC�{���r��v���퐆��$����	������ڐ��h�O�߯�+9W��R;���y�����ߥ�)�]T��K��u2q+N�Z\�\�s�*�pPu ��m0�YB�ƞ��2{m�sk}�C� 3sS��`�:�z֗��SG�"�$�G��R�w��Mr��N'éR�09j��i�hQ�k�-��YəK�6>g�"�Of�4�k'��{+>EV��">J/@H"�$vc{Nv�I��wm�Ek��=� 6<���e�8M�k(D�;���9-v�f~G��r���'�A
�vi��qD`���Wf����myPм���y�!��:A�b&l�U"�_.��׵̛����'�ж(.�� ?��F�-�҅)��]
_��C�1��.*E�dD��M����D��P���n�v���Ѷ��:�L?��;���$��b�闫�ff�:�6�aYJ#�	,ۜ�M���)F�='�u�!F�}ʶC�]w��{|�羭�s9Z�)c��-�=Lb3%S��|�rP�mF�qw�w����`�S�R�e��f�y)��u@�<��k�'[>�u���ccV������2����[��ku����"bR�� iX�8LĔhb	����^���h��,��uB��`��Vlc5+w���!�Y��0�x^j9�ha��߲^��8	��8��}(��'�40P�HY��hi��cq�5�%b ����v�D��A|ڱ�V3wR�tSo�?��p1#MТ��`��ڬ_��Fw�	��`�ch�E>���8�8p���g�p� #��J�s.5I@4�í���F�VV��K2�2�XC�V���S� P�tQ�	���6�3��QO��B�:nk��/d��d3��c�F��=t4��L $l�QA`��7l�P�KݻH5�anԃ��s�If�t5�?̜?�Q�6�}̀���C�#������%������O�j�3����g��A�=���똴DS��bY�Rp���fH\r���?�R�r�(��) ���	W�8U�B�0�_4m/��B��|�j�Nds�zU+►z����(���i�?(�����An�j����@r�@}y �6�40����㯏���<f�Y��j���31!�����d�G � ������y��5,�Qi����V(7O�m��/��g�F��A�4:2�r�Q�U�crI��tAB�<���p/�C�G[[�!rߋ���\��DB�7�Q��b�]P�,�4��&{��8#�-�U�R�w/������@��*c�pp$��������|!~�����a�X�OD��ɮp2���bvM*��	�l;��W����~g;����c�\P����c3Z�YH6�����	5v��Z��H\��dX��I������	9�K�	%|���&]���!�� ���~cYN�ɛ`��{ �[XoK�XL��y�Q���͊��v�o,Tu����wL��XA�؀fH%�;�IWHچb��ѐ������. ����w�1�'��]�q�FW�^�"��af�&��u�����Z;�}����+)�y_$�3�R��_./�y����Y�2��!�"><�=�8��x\h�Ո؁�;^[�3�TS�T.̙�	ŵX�)�/mC�Ԯ���4B��څ5_83�sҀ�j���oΐBh�lKc|���,*xY������	���>���%���W{�N9)��kmC��&��4x���~����f��A�7t�~j<���b6�[r�mh���u��dt��4)��N�j��_Et�Rr���� ͉j$H�IX��mP���5y)�l8�'3��v��v�F��T�)u��8J�+�3��e��!����RO��z��w�Y��mY@Uk��M�򀐞����9��̃{�F�9�/1�I������<�B/����c�xc�-��ϕ���i���t3:�q^�p�W|��C�1��e���=1�:�����qx���e1�A�PV�x�GD�dZ�A��W����0O�3YD�Z�l��Y����g�-�=����vs�d�"`��z��U�����T(k��ےs_�J��w�9��B�xKG��}�\O͸8k����5���$��\���7�8!S�݁W	Qa�1�o�љ�Ѧ�L�R�cU�`E�G�gM�)-�����8c����<��U���O��^L��y}���Hf|�l�v�]�$Yʽu�P�X��gW`�ܖ9}F4��-1a���+D  �l�$���`��m�"��ZT�j{����ˣ�[��� ޴�Zգ-�-� @�ht����(��k�g�[*,n-��[ X=*q5ϧ(��W}��è-�&���^��HII#��� yPy;�Ϊ�>>�iR�"e=0����0�/�G	�2�z��?���E��"}>j��+�Dy'$4�(o��Q�ҧP�6���r��m����Ed��Î���!,X�{3M��walH���<N�+�ZT�:��z�to��Jp\+��J�p��+fa��ao���>^��/>��O!��>G>��a�9gss��e�ܷ�V���#/$(,ACXU�F2�J����<����;�Vg�Wm}Jae�����O��=ë�8���T����ܒv��!���udXBW�2�@��}􂢼d����%7��^,��j�1^)���>�Е�e�Nd�����PG��_��!��k�L�T���N�����OS"�:p� �Y���[ƫp�SĹ�����3	������^����&�������v>�V�#���%l�Y���҅���Z�����!-�E�j�C*+�0�o��`?K�I�YZ�~k�{˽��-C�#�{�:��a�[>8R;[�Bm�?;x��RX�v����E�.�"+<rR.��%�]��\^��Z�R7�:�h��p��3K��:�i�j�S�%@��8����=�.B���q��>�J�BU��(���˦q��ŏ4U3K�=���[��%+�Hl�#f��%��� �[�����!�����怯4�� �S�(6b�?�Aㇺo+>á/_:�7���v�LJ-v,h�ӡl��3�No���-G��u�Nb��=;��)a�V5D�vhNF~���ۆV��ɟ1�.��%�?��Z4�><�~��^
�#�>`�J�M�=R��a[�UT��4�r1>���}b�b��Q�@�0O����oo�斾�!�2��"�V��3�zn_���I�@��b(�\����-^/
�@`��J�X�%���k�XΠ�}��̣����K2NE�W�OY�ߺ#_)�C�_m�'`ċY�>K�����I��V��#Y���o�0'*�=�p�
q%b�q&_�b�Q�+Դ�tl���k�=s��>�`$ig�uܖ�T\�:�`���Rm��o#S�.��΋��oBĝ��[{��������(�a��|���Z��MӍ��.�" �ԏMDw��x��z����p
�����ͳY�����QTo�(I��k���U��Mu�=�������q�=�b�#aĬ@�b��7��Ϙ�4
�C��Xa[<���$,��&��D|��;#%#�"�'��v)(�i^���ӕ�/��80
�>n�:����%S�sX��
-܇K����Ј���\�V9�*�	���(��ak~�n��Di틢C�yj���/����g
Q���4�Ď4.��N���UgPN�^���J������*���p� u`qW.�������~�/���=��55���`��PV����f&r8x����e�TM��J���Ӹ��S�OمY��obN�tM���)��Q����"5����+���&���h�R�,7c曠��<f�Z������(݉�3~�7���9�>a�|��L�t�A{�,������:�9�� �&�v�{�B,�V�S7,��F��g$��rb?m��3������l��5��9�.qy��	�T�;�5�߮��+�77{�m�Hk�O6@����}�����L֡+*ǽ���e��Ü���H �;��V5��%��]����B�ϛy&��$ҢI����GV�����$1��	����Z����Tި�s�$���~��7����V*p��W)^��c���H���j!!��o� X
�Z�a6*�e�	l�Z;`w7�/���M�͟4/H���RD��6b��:.Y�n�(�`�8�T4��f�u��y=\���O��?oPƥ��q9@�]�?�`�
��U�m��c�I̲��>6�ȶK�`���֎�U��䔳��/�f�.B�|3~�+y$������$�~ٛ� n�m*�&"��/~֣r����u���U( Q����Ў��}�*�3�p1H�2F�u��A5ɸx튑�fK��X�Ra�Ui�=�<�E���`Bo07O�=g<�_��<)�/�`Y�1�))ޞ?�'�E��ƝB��r�5|;��T�=ʜ�|�Z ZD;r�*Ynߛ�)Όa�C���+�Jf�Gm�K�`;sRn��=gU���H`� �!�CM9c-���J�OU��n%F�vW��I��e��UAt��3j^c�y�J��L��SAE�-fh-�Zl����b!g=��N��P���s� &N�(�y�-
�W�Q�_3�u�0��?�f��Y\���"��2�ā����55��b`���/]W�٫Χ0�)ҥ��]{���8�e_bL�y$Ȏ^}zey?��� �1����T��N>��g���Tc���{�BEXm�t�ɽ}�1qjWn���K�@SkH���9��nZ^%F<�G�>vH�3��!!w4�>�)��2�qt�}1{�zn�Ag80�	Wv�O��f�������ŨBP�8������IQQm  Fa�L�*�v�hQ�3E6
�a]��|�s�8n�QDx0�zO�VK�
�4e��/q�]�s3ؿqϭYS״ҍ�v�8l�4�M	�=��-C>א�m١�OU��Uk �ۃ��Y��g˩�g_RgU��x�UG�<g�����'{������nCMks-�7�x>��C�U��W��pOF�t�T ��S<�{���]��o���C�X?�W���I�d��t��5��Qdʥp-f�@�l�-����]_1��??��RX�(N�����w+	F�͇���jQL��J�D����l(n��z�U���0Qy&B���Y=_l�<�(��8�ЩW�-�ܙ�鄝���o��׉hJnI�q���b=��{DO�`Њ6u���rF+��\ڒ��\!�
3�ng���ϜQ���Ό�E�q.��U��ȓ���E&Z��� �X��D�i�NB���c^f����n��\�C��w�G�j)��e#���r>��2��ۺ�Nf΀l.���x{(�r���,u|!�63imś��k#�C!��v��Ƶ�Q��j%Ai[vj�O�ل/�"?�ai�:����z}�qC���Ec�1/)����N��LB6��ى��9V�M	����H�����nu�t��CTfV@�5�h�38^�P�)�eUH𦓭
��G�4���l!}YWe�f~���x�B�e.�8k�be4�l���#��?�Ϝ�uXD��4�TU균O��s_�Búj5��5�f�|�Yt!��]l��!I|���l��l�����`C����j�SH�i�M����.�Ȅ�Mx������؎�dW%Oyq���kA߲V͒�H{?ΏF�=�r�3�$`�"$:��?Aa �ټ5�?`�� ���>�>݃?[�����@41ϛ���_���R(�/��R����g�5I�79ˬ�9h烐R%��׷� ��I�B��6���`�҈��P�����-0�ƈ�|��l����V���p0 έ�/w�ag�}���w�cE}AYP��Q._�=Je*�R%�N3xȰ�"��$����yX��6��[n]*�z���,��t�!�R\���Ź��� �J�Ull[\�O��Q���S�`M�h�-P`L�"�X��������2��έ����M�7XE�h��i\1�O����c]�s�aH�-I���r,,��a�����;���Q��?c|����1������E�������
��{,�:�
dTh��]��[J�ߢKR�P���e�ִ�$��M'G�Z����iA|?҇P��o������{,ӁUd�����7�g 훧@�m4ѓ"#�c� B�/O�O�G�ix�Hh��0W��ʷ���x���%����!_~��8IVh����ȁ�pڦ�&�#&�☬��$���)��;�+��{s(���BHs�Rac��zaPN�N+�V͖���4he��rk�k����LIx���]��|�Ƙ�������ꊊ��h#�c�-چ,�%h�cl_(�����o/D^e]R��^�*��	М��Ó�W�L�`��z��,)sC*�]�^q�Ҝ
����p]|�������{��$6�`+�c����i&�L����D�xP:���d��D�]��K7H����5��Yg봐�4��G� l-���ef�� 3`�@2����+r��/uF��}������.F����:z8�8X3��Db���+��+7��3b-P�%t�r��3PY�=�4���`�����	����d&���C3o���Z9� &]z�HXD۽��d�xN93��	*c�i���q
���67�L�pyw0<Oաs��2ym��]�8��@�Gy�?�>Ԝ�w~@��}r?��Scw�[���i�u�A��1�<U��s ~%�T�C���L̝s���v���wf��e����Z�����ُ�Q�������*�W�]x(���r�u�J^ҎoP��+\m���ѷ�ĺ����9_�V���Va�H���v���$��s(BH"��� �#����@Q�]�M��?�ko�Tj�'������U��������%���S�����\%���=����Xz<G*~�ʑ��z�fD?�Er�k��~ּ[�s�J⸈�Ï<���?-@'�T&�0iB�$B�����]�!	-/�ISZ q	�fsPݘ��Ap�$~���®���M>Rp%Ĵ��*�rh<��!��`bF���cO(@xo!��
6>:��B8�h)��|:�{�� @��1���DA�U���|K�/��H�=`Ѱ4��i�!���!5� D,]\�5a$��h�R��֖�
AuA\��Cyÿ�`c��
��Fl���ܧ��U�̊��J\`���|�D��+F������M�.�������\�'DQQ!��@!�=���Ix�*]�A߻�O�İ���>,L�)_�����1}L�B{'�W^]^�층���毬1��w��\;�2`���L̅q��{���tAu��n�G�6�s��+ZRK"�� ��j����VV�}f=���Ơ٢"_��t��׷ծqa(�P��SЊ��eB2�[7�P���P����M��;_�RL��R�p|!��-�_��^��y~����,M� u����f�Xv'�{u �T����t��ɜ�&>=x���t���`f�H��&�~�'�0��CD*\�jƳ�@�"���J��e^����ȫ����󍑜C؃���\����L�r
N���]�5�=�8�|:�3v٨ʷ, n�P�7ˤ��rQ�����S.�𲥶M(���>E�xG���9�j���x�g�K1g�r�ZI�G�4�@qoE�l��h�Z)=o�5|���pٴ�ak���ی�gX-�Uڠ\��B��� @dy�x	��>P�XeBt��]�=iŉ�tč��%m��P(mJ8��=�B���I�v.N	�&۔GtF����9O�q����;�r�;p�˥3�끓ׂ����m7���	z6 R���**���̯wGv|)b�v���'�O�c�J�֒y3�R�t������e&"y"����D��@��a�F�<�EzQ�^�̡?>U�7���Z3Ϥ�^��LqLHK�&ІA%D��=���ZLe[m�u�4M��B*C�!T����0��ҡ����
���F�^��g���V�`�S�u�
S%��o��,�0\�cz!0��L�[�w��C�- �C笊�	1��B8í8��So��'��4������ ���ڍ�V�
�C�2vסƒ���8h��F�].Z`��NI7�:cB�E��LN�]P���I��[�E:��n�(����''�?ߒ�%���O-�YީXU�l��R��:M!K�������|2�!����F�w��j���_C�mqI}�^x!o�JI�@t6��3֝�R����6�_�'��Q��&�^��1kB{��Hk �VC-�QgD�o���I�W�����&���q��=�uy\����DsN�	5�r������|�2o���"C�pw��|�؎����N�T^����.c�"ьq��u������ ;�l�!�Ř� �V+j|zz�fԱA軉�]���#m�H���N#=��w���n���)L����`HxFS
�ތ��~�<�Q��Grnf�?a��4	�.�U�� B��eZ�mmc�*��� ���P*#@.np��-���$3 5�~Qa�Ő��E�3�� �uN�j��e�/�B�k����~�ψ*��D;�P����R $[�.�:Ft
@:�dӓ՞�ct0O+���T׭���`���{gD�����&�������h��s������� |�qs����?��8 0�h[O%�tkm��>��!�	M I�2�F�wSag�6�gm��<��i�������z�Ϣ��푰ԙ^_��խ���F�^+�G���XH �aTŋ���=�_#um~�עꅄ]��N�gʁ�"�V!�$���'?�G
�'
"�:k 0ZΛ�@\`��v>�BI�%c@����e��Ǿa*" ��2?����G��g���7C�*`QQ��4���*WfPv�cI����2�?p��&4�w��0��g�	p���*Oh�F���Ha;1ww�o*����:ށ���r����Uw�$���*��j�%=.x���.ݞ���m� �9:�� �J�:��"��1L�ʰWniO�3c�F��g ��(�ܴX4�9w\|�ۈ�a��K���`���J?c��17n���$ �!�y�A+��eS5��7E���f�s3�Gj
�S	�8/!<|�x->I��\nV&d.���L�Yw��ɢ%����.޶���n���5��x�3���5������$����aa���f(��H�����5?aI�yto���F�-�	m{.�����!X�O�r͈F���I2oL�X��c��
�'�j�a�c�R�.:،�ȫI`,���o)]�����vu�q���l�.L��Ŧu�.�WwT'z@X�MW�����`K�ݭM�������8I�����>��d�	QI��0�qӨ5[�H �M��Z��O<��+�S׫�-å�IY�Ҭa�m5׍q�~Ǜ`�w[�Y)j߆��Ur$��i@�9�Iv*G%�ssC�-{��X��IdP�F������Əz�������cz���BI@��GK�H�d�&-;�xUZ[���{0��#q�1��};���w��v�M?A1��k�W���!B�$kS�;�	��B!o��43�Aq����"��R1Q���C�M-���U����.���l�k��\Al���O��~����M���}I&�7��K�eV�qPN��S��(wׂ�,��V9UH���_wk�%��e����G���&��bi�x���y��������Of�5B��7����ћ��7��E�������������6��Q���;jF�-خ^���y���d�DbsV��5������vO�����.�M!�������6��*�%���j8 >��ې����U'�V���a�6$� [O�^?�3
>^Ļwh�g�����ݑ�3� �N�y��l���/�O�.)]���⠕�p����"�27u�Qܨ�aذʅ�8f(_��0df9{U�CN�M$�k�~�v4s�U|ͺ%±�0~,?��(H�I�D������k<��.j!��r��[�!~�_Қ���\��4� �0'�>e�����4���s#��h���>_�i�2?�	gG�P�!��$���}B��@�f$��?��v_�\O��D��F&�ܤ٣$�Y��O�\���>H΋|���ǎh�w>Q��₨�,N���(�t��ju��jN�Z�Y��s�B>� �rq�*�mû>}F�J%�.��s�6�pP{���4�d�FAW�����ݴ0�@�d� ����a�u�ϧ�*�w���É��ʚ�
�$Xa�T���D�����Pj=u�s7��s�7
M�@Q:���L��I�{����EpG�RK>��7�eǬ�3��Vk�Zv�"F�mɟ"�a�7"�V��:�4�'*��Xi���D&l�]�\�Z���=��Ht�
�*��s�SB��X����Y3|�2cS�+} ��̈́�oh^TǸ���-�Ҟ��E��EXO��(5�](I�{�x �_|�l\��ރDͰ��=��M�L3m�6�fM�V�}E҃�swf꘴�)�S������`hq40%[�A�O�1��.^¡�� �G
!H�'o����d{�s'�5���i}�>3Oe�Y����	&�٨"3��������&�xĩC+�.=����(�^T���;~oo�zt������>1'�O��2��0�P5�c�.�1#?��7F�~�k�l���9V6��՜��vʽU�,�~H�?�2H�~��CQ��_
vf��/w=�N�k�.ۑ?�*����bM�:�=���j[��N?�e@��8��3W5�B��������B(�S�=<
M�-o�f��6�~� 
���ID>'��؏���"�)2�tM�x�fߘ/|R���=����x���)���z���劜�)�6>���7���\����[P%�8O�,�90���/A��9�iÛ`��z��P�AVk9E����~;V�ؾ���e �SqL�C8b
��u���i��N�y/2�m�9�@�K�5�c�����]��Y���W���RV�����-�o�����4�}�Ĩ��~�x���=L'�s�t��CA5Ԁ�a�n��Ɉ�؜p�b��a�h����ԯ8TI-����co��bT?�	���uR��͇ЈΫ��
�BcP�q�`J�A1ls5��A�P��A��z�Ba��5`sؑ�|��TG3�jw��>�f��5=�#�Z���*`~�f�w��^QgxJ��C^�_��A���-Du�7��YK"�✴���O�ND��A�7�8�U�c�PĬ��i	%��IDR{W��7D6��/�H�v%��A���%ؒ���\�Wr�B�)��+�/��_����ػmQ�bH��5n[d�~]�w-�w�Ÿ���b�d��*��˛u2  �~��`bG�K���a�Ee!$�A�)���� F�@���z���4T�[������E����E-��X����88��׍o(����@3b��털!���]�����Ĵj��ܲLK�\��@\�[�������{t�
L�<�k.�����}��:��jg�{��,�{{Q��	��:��/����=����JJ �(��d��7�{˼;�n�jÔ�O��ց��U�Ɠq�ޏ�� (�󱝴E�y��1C�7,h��I	)8�����x����D�-Ek8�bUn�Μiwb:S^�x=�_�L	��M��$M��
�jړi�Z�S���h3�*ɱR����`A�D*¸)�ξ�6�i���aYi
��&�^	����x�C||'c14$/+��"·Zo��Xg\M�d�fN�K�I.�4*�?�E���c�8O95���o*�7�6��22,Ž���ֳx��dd��t�1�d���~7���P�������NϹpp?V��F�,�Ƃ�����17��l��v��������; bN�ӈ�����wo�M1��M��f+E��7�wtm���:gd�3��&��ج���$sdud�r�LxS�-2ǜ�V
i��7�$�at�|YQk:��P����s�d/��4 ����A����$���������am.u�7�w�DRʚ~�v�W����	36�u�2�Bb�r,<m{��(1c��}�J���yb2"��T�M�'�G}@%ұ������::��j�E�f�cKG
Ȳ�k ���|#)�"L%��*�0��A}�k���U����o4�<۳Tx�r^B%�}ÕK@;А����gmn��M�tB7�R�p
MY�7JxFd@�y+j�Z0��&E�}nטH{�|�Z�n �u���$�f�R�i]}i�K<�v�v%|<2/5ls�uZ��Q�����o��A�&�^�%%] ?���$���`�4��I�p	栂S:�Y�����W����>v���q�@bŗϹ@�[��b.�#��M�!�Iڢ<�ȫ��|1���5 ��\�{e2�rڍ�6M�C������%ωE�߿I�p���0s�qp烂CъA�j���6��$
��T8��PJ���$P���M� f9 �������� ��Զ@�љ����&�+���y=���u�GU��7�(L���Yt��ٌ$�҆���b��t�@(�Q��r���%�/���h��.�p`��ː��6������ t��ŅWx����E�]ܠ�ැ�Μ�u��Q_O��e|��
�5?��2k�7'vuQR���#Ő����?��i�ΐZA������r������J�F� 6\:Q�K;��ٙ�����!@�O �h����`k1w�G�8����|� �A|��M��Ȏ�'B��uMC�ނP�ڞ�\/DL�1��{Fy6�ދ*������8q�uI1�X���Bc�-��~.T���`�r�Ĳ�}3��w0q����b M��y��̕3Sĭ���M�M�+;����g�&����ח��Mc�˒iEڨۃ�!M�}4��|)�S�������j�|%����j��mK�!��pA򴖝*�IF,%BO���"t�%���w�X^ƿ����P���>k}=U�f�ճg`�znqG�����C}��@����94�)pC��H3塕�z�X��W�w�p��z ,¨õR}y�;���T����%�ZSO����[�����[9��."�Y<e͑Kj���E߁�j�"Ȉ�Y��vQ���S��SZ�P*�� ` K~'v���h�lJT�7ٖ'���.�a�lɴm+p��p��WL�+,���R.&M��bc(�9Q�����>Ns�6;/kϔs���0��x��Ѯf������`�[��ETK�jl]!��	�3���1���]np9��~h ^����9��#s?���C&-����NA��&A��ݐ�ݾ֫^@���:�=u*��G	�,�D0�c:͡�K�:%йR�r1��3Hzmhz����{�g���$��BK=l)ΙH��vN�[Ɂ��s�U��H|�J�BCT�������R�����K����rO׸�db���v�U��x��y�A�����C�����y��y��n�~	Wu�c\�V��"��J�oU��on�,�_k?���������`x���K�ae��Gx�B�]�$�s���Z�u# iV_��l!�9�Ȼy�ܯ����gc�.ddn*�2y�&��\b2I,��L��'Vկ��4�'L7l�Ѣ�;�o�.)�&H,�W	���߭:ɕv,y7�=��*�~�ޠD,L"���7P��:�ՀT"�#�{K�_'.4��b�<I�m(O��_�)����m͟���S�P�1��|��#L�Bqs�f�����*'X�k��b��.���]/�ٳ7���������`?�V��1�"~ec�<���p%���;�lR]'���j�&�O�s��U�:�7[���^o�V�����6)k�ͫ��{�U��]�@�xH�~������(sC"Ȳ���!F�x� �Q���1vf|���gԮ��H���A�c3+�׋磛N�0Ri�������:���[���[�]���.$Вn+�һlu�� گ�a3Q�,I�E���^�=
{�x"��[�b��O�#�ͅ	����K5BFb����
��E��xZTЪX�(�4�S��e:�v3��1��T)5Tkg�H]�x#�[PfL����H0�*$��v5��0�[��W��%���s���ya̢�IQ����,�3��m]��;�f�V9i�#���" :����a�i<��鐓�]��>����`�����@&�9Y�<�ۮH�ai^��a� #����-]�Z(�&��~�0pl�]�oW�˳���MaftW��@�x�:�+b�u���t���.)F#Ox0aw�׏t���]RZx7Z覸�@a��ȓ.OK	2hB�Y�%�7���AƟS	ŗ���!Ye�s���<g�Ԃh�¯	|7-�����z�H���$�����QZ;��^��U���&25Z�#>����'k�t|	;e	�aے<	oFҖQ�)ٞ�N���p�R _Jz���v�6 �j�W�1ZK'��馢S��ܗ������-D��e}�$��� U8��\\���������/f�=tf^�@�dD��ǃ"ݺ�#��������q�d?���[KT�ӥN�^Z �)�
��	4u�S�F��^s�ԝ�:ny�Wf
��a@����}��d�սȴ�k|?�ϴ�!��
�w�@9��h��W�3�O ���]Ub��[����99��Y�ܾ՜�R~XU��Y v��� ZR����v=6U���60�
��8�x��M�s��U�J�/��,���]�Z=� �l�"q
K��sJ߱b𳕸O4F,���Ȇt�C>�e�|��N*���;2��/��)����K�6��x�Ԏ2v�譃gF݅�EзE�n�<N��8�����у��62v%�6�U|[�sn�eg�/�:�˗F��әn��Ig�����Ce��AȷEg���1�rü�\�|��@�R`U�g��J*���}�� @ۏP;�����Я�<<?�
E_�����@8��J������a31h|� &gE#m���I���=�ٲT�-���ә��/�)�.A���:�Q\O �7zr.����mv��jދjxSUcl 0���6�6�����K��Gl��f`%k��9�'�P'vUyF�ͭO,�ݮ~#�n2ޡ
�0I	yR�ƥr��l�e����"�R(�*����`�    XSQVWP�$��pQ ��  Pjh   Pj ��PL ���Y���P �RSP�ǉ���P ���X�$h �  j P��PL ���YX[����C�����	�tF���   �����t8S������<�s%�   ����   	�z	f�%��  �ڭN%��� =��� u�X_^Y[ÅR�ۅ|�b"O�ř���ㄋ~���:���x/Ed(@n��\�n�v��wݓ�NG�o�3s�t�� ������7  ��������  ���   ����^� �W�1ZK'��馢S��ܗ������-D��e}�$��� U8��\\���������/f�=tf^�@�dD��ǃ"ݺ�#��������q�d?���[KT�ӥN�^Z �)�
��	4u�S�F��^s�ԝ�:ny�Wf
��a@����}��d�սȴ�k|?�ϴ�!��
�w�@9��h��W�3�O ���]Ub��[����99��Y�ܾ՜�R~XU��Y v��� ZR����v=6U���60�
��8�x��M�s��U�J�/��,���]�Z=� �l�"q
K��sJ߱b𳕸O4F,���Ȇt�C>�e�|��N*���;2��/��)����K�6��x�Ԏ2v�譃gF݅�EзE�n�<N��8�����у��62v%�6�U|[�sn�eg�/�:�˗F��әn��Ig�����Ce��AȷEg���1�rü�\�|��@�R`U�g��J*���}�� @ۏP;�����Я�<<?�
E_�����@8��J������a31h|� &gE#m���I���=�ٲT�-���ә��/�)�.A���:�Q\O �7zr.����mv��jދjxSUcl 0���6�6�����K��Gl��f`%k��9�'�P'vUyF�ͭO,�ݮ~#�n2ޡ
�0I	yR�ƥr��l�e����"�R(�*����`�    XSQVWP�$��pQ ��  Pjh   Pj ��PL ���Y���P �RSP�ǉ���P ���X�$h �  j P��PL ���YX[����C�����	�tF���   �����t8S������<�s%�   ����   	�z	f�%��  �ڭN%��� =��� u�X_^Y[ÅR�ۅ|�b"O�ř���ㄋ~���:���x/Ed(@n��\�n�v��wݓ�NG�o�3s�t�� ������7  ��������  ���   ����^� �W�1ZK'��馢S��ܗ������-D��e}�$��� U8��\\���������/f�=tf^�@�dD��ǃ"ݺ�#��������q�d?���[KT�ӥN�^Z �)�
��	4u�S�F��^s�ԝ�:ny�Wf
��a@����}��d�սȴ�k|?�ϴ�!��
�w�@9��h��W�3�O ���]Ub��[����99��Y�ܾ՜�R~XU��Y v��� ZR����v=6U���60�
��8�x��M�s��U�J�/��,���]�Z=� �l�"q
K��sJ߱b𳕸O4F,���Ȇt�C>�e�|��N*���;2��/��)����K�6��x�Ԏ2v�譃gF݅�EзE�n�<N��8�����у��62v%�6�U|[�sn�eg�/�:�˗F��әn��Ig�����Ce��AȷEg���1�rü�\�|��@�R`U�g��J*���}�� @ۏP;�����Я�<<?�
E_�����@8��J������a31h|� &gE#m���I���=�ٲT�-���ә��/�)�.A���:�Q\O �7zr.����mv��jދjxSUcl 0���6�6�����K��Gl��f`%k��9�'�P'vUyF�ͭO,�ݮ~#�n2ޡ
�0I	yR�ƥr��l�e����"�R(�*����`�    XSQVWP�$��pQ ��  Pjh   Pj ��PL ���Y���P �RSP�ǉ���P ���X�$h �  j P��PL ���YX[����C�����	�tF���   �����t8S������<�s%�   ����   	�z	f�%��  �ڭN%��� =��� u�X_^Y[ÅR�ۅ|�b"O�ř���ㄋ~���:���x/Ed(@n��\�n�v��wݓ�NG�o�3s�t�� ������7  ��������  ���   ����^� �W�1ZK'��馢S��ܗ������-D��e}�$��� U8��\\���������/f�=tf^�@�dD��ǃ"ݺ�#��������q�d?���[KT�ӥN�^Z �)�
��	4u�S�F��^s�ԝ�:ny�Wf
��a@����}��d�սȴ�k|?�ϴ�!��
�w�@9��h��W�3�O ���]Ub��[����99��Y�ܾ՜�R~XU��Y v��� ZR����v=6U���60�
��8�x��M�s��U�J�/��,���]�Z=� �l�"q
K��sJ߱b𳕸O4F,���Ȇt�C>�e�|��N*���;2��/��)����K�6��x�Ԏ2v�譃gF݅�EзE�n�<N��8�����у��62v%�6�U|[�sn�eg�/�:�˗F��әn��Ig�����Ce��AȷEg���1�rü�\�|��@�R`U�g��J*���}�� @ۏP;�����Я�<<?�
E_�����@8��J������a31h|� &gE#m���I���=�ٲT�-���ә��/�)�.A���:�Q\O �7zr.����mv��jދjxSUcl 0���6�6�����K��Gl��f`%k��9�'�P'vUyF�ͭO,�ݮ~#�n2ޡ
�0I	yR�ƥr��l�e����"�R(�*����`�    XSQVWP�$��pQ ��  Pjh   Pj ��PL ���Y���P �RSP�ǉ���P ���X�$h �  j P��PL ���YX[����C�����	�tF���   �����t8S������<�s%�   ����   	�z	f�%��  �ڭN%��� =��� u�X_^Y[ÅR�ۅ|�b"O�ř���ㄋ~���:���x/Ed(@n��\�n�v��wݓ�NG�o�3s�t�� ������7  ��������  ���   ����^� �W�1ZK'��馢S��ܗ������-D��e}�$��� U8��\\���������/f�=tf^�@�dD��ǃ"ݺ�#��������q�d?���[KT�ӥN�^Z �)�
��	4u�S�F��^s�ԝ�:ny�Wf
��a@����}��d�սȴ�k|?�ϴ�!��
�w�@9��h��W�3�O ���]Ub��[����99��Y�ܾ՜�R~XU��Y v��� ZR����v=6U���60�
��8�x��M�s��U�J�/��,���]�Z=� �l�"q
K��sJ߱b𳕸O4F,���Ȇt�C>�e�|��N*���;2��/��)����K�6��x�Ԏ2v�譃gF݅�EзE�n�<N��8�����у��62v%�6�U|[�sn�eg�/�:�˗F��әn��Ig�����Ce��AȷEg���1�rü�\�|��@�R`U�g��J*���}�� @ۏP;�����Я�<<?�
E_�����@8��J�����