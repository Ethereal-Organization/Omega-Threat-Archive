MZ�       ��  �       @                                   �   � �	�!�L�!This program cannot be run in DOS mode.
$                                                                                                                       PE  L ^B*        � ��     t                @                      P    ��        @                        � (    � �                                                                                                          .code                              `.idata   �      t                @  �.data       �     |             @  �.rsrc    �  �     �             @  @                                                                                                                                                                                                                                                                                                                                                                                        U������UW��VS��j �P�C �u%j hxzzXhNODAhAntiTP�T�C ���t�ɐuj �X�C �����\$�f3ۋ�@<�P�T�B4�   ��APQh/o�~   TTj@�r0�r4$P���T$�XYZ�[^_]��Q��$ ��U��`3��U�M�;Ȑ�u������u�O���ϐ+��А2��B������萐s5 �����u���@����ЉD$�a��� �U����`d�0   �R�R��}�r0�   f��f�t���   �u�}�<Zw<Ar ���j �E�P�Z����5��j�u���B�ؐ@<���@x��Ð��p��}���   ����Ð�����u�������B����j �P�����9Eu���U�������E��� �Ð�D$�a��                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                  �|n@U�G��j^�Mk�]���(`�Z��'��%HiS��OU�N>�j[������~�W���V�w��#Bi��)Q���ƞ��$���Nܣ���9b��c��:Z�Q,�0�`�    [��;@ �G   �D$���   3��                                   4&�kC   �vH7B     @�@d�5    d�%    ̃����;@ �̹   �1�$�T$�1+$T$��W�����d�    ����㐹   ����;@ �݃�;@ ��.��ѐ���f� t���؃���ܓ�;@ ���f� uܓ�;@ ���f� u���a�   �E�a"���i͏^W3ҥUR^@�OMJ������(?��73]hf�99����3thc��d֗�m�R"myr��P�d���"oyz��e��Q�tQ^D��w�[����z��N� �yq�1Э�a�9x��(*A�};�q]����Z��S���7   ������   ��3����3�������@���+�ȋ�}h����K�����u�p��'�q["��kq�`����k�($�"A��(r�rqpq����(N��%��kq(����l�'��l����tq i!��q�+6/y(�I� X�(�L�دq��K�'�q�'��X(�dG��q�5�O�&+Γ���`� �����v��修�/!���0�P���c���3a����(�tQ�!h�*'V�2�	˹�"�@;��p9�@G�EML$��m^{�E�])@�=~\ύ!���w���U~��:����g�*]��:���ب����_��9.B��L�4޵�?�Y���ֈ���ð�/�Y�pΊ���Oʎ�OY� �b��jp܈$��&��j��8L�e/��vq�(Gl�~:��v��i�5�@�N�]ȅ�r��C�}�٦5���6h�'��G�X��>�(���7���4�v���T��5˘r�;3�� v��J�P@�S�P�8�J�
Arg�zd�9U���bɔ�.��Q���Ǩ�1�W��Q�H嬚����8^�q�lk��v�&�ޟô��q�qj��w)��,�/��-L>{�a�6x��,	\b���"Ws��
� �<&��^��k���܉-���}v�N�ϗu7h�ܤ13Z ��0w���%�Fw�ҧ �1����_��<(A��H�%UP#��F0�l��1㟫�3��S��7wcD�x��[QHr�3��X~�dM���y)�=��Rg�mI�L<���a��w�h+��m�o	E��m����?vw�u1\H1m��I<$�
S���0��,�\��?���A��e���dCU2�(_��6��6qa���(&�fe3>�˚��z�Nd��f�"iЉv�]��ʛV�9���
J��J),�������\(�6 /N��ܹ���s��@� ��C�u�G*��D��j���:O�*�L$��u��ݓ��/�ҫ�"s�Q*�*�kb��Mq�*=�S#nǸm����:�?rm⮟�u��;;��e{�q$��(i&��y	�,�EPZ4�qze�Ja�r�ГQC���|�Վ.T�8%|�Lǝg�J�b*���!#Y���0��HٶBxbd>�;tv���)޹� -`�j��\^4��=Fŏf�J�D�w������'����HVc����C�"V�����W5�QA!-���X��1}C��\ۏ���D�����qNLV~@},@]uf� ��ߦ�N�DJw�&�j�wbѐ�wrD]Hi��f�{���˕_i�.�%��#��1�b��;�19��Fh�
�ؖ%�k)�_H-j�	��]Sl �l_4g���U�"!���6�H�L8�ې�C���VK�1xcol-���$8T�ݬ��V
_�,��*!C��$=�)�O�7�c�G3�U��^br�?��Ubްy�����I`p�96�t��*B�R�"�gq�Qg�T�6�d�g���n^�}���I���* N>GA'�,_?���Й��*�Ɲ�T��X3��hI2����X*��b
����6�{WO{w��D�`�N�8�d�k�a�1JD�=��z�����Í����QLy���sQ��g���l�i7�:|�kN��X�rs:t��0�>t�7d
�ҭ��+�G���j�a/��o
0��Ld #����?�����C�d�G�v4�e8�SG4�1]em�,W}- �ܬ���d�Ң�D�V0f���~�`�"8�y;#A6v�*���H�`��ؖ�Φ�F��QV+��̝��Zm!^
f��1a�(Г�l�=�:?>T�Xu���s̰��c�E;O���~,�8XRr�9H'�Ngb�7���y�����L�*rYĿ]��0C�u�,ߡN�p�U���n����L�Ym��d��D�EMl�cL��z�ڸi�Jl�_&�F�}c���V�ٳ��5ȃ�C��K�
S<���IuF&���bBQ��\[�Ӈ�~�J��

]K�)�,&������T��7K�B�Uq����pk, �${jǅ^���RG��ɀA~�Ww�Ƒ���=[�ӑI��v_Ã�y��j�y���Sp���Ҽ@oU�m+��_�컆a!v/�� �7����f���2X5dv}L�OJ]����֦����Ñ�>�L}Jv���7U�A��T�����Q����w�� 1����@>Z��&$�L(�a���ȤBF��P��Fր/O�Z��� wn$��8��E�M�9d*�茳�Hb�Lz|F\ /7�'�Eq�T�ȷk(8f�����$��Vr�'�D0D�т��á�W��靽]��x�(`(8�k��B�+yш�s�x=jk��:f#����i�IL�.���ٴL)���r��~�R�� A�ń���"�C	n���$�F����O�T��]X�V���th[�sX�|�W��O-�	>�X�����{��c��[�!c��6���4n�
�9��� A��aMm4�x9 ,�����6��к�����S��D��=��Y�����#�`|v��y������
�n$�Ĥ"d	�;μ����{+��g`��1��2��J�E����H W�%6.C�p2
�!��z��P�>�gc�E��>�V-��gV�ѮX��m�ʢ�J���\�q��]�43��tNPÜe�2�M��^��r�[g�mIW��ޅ� ����ǃZ��j��٫�����{̡ىKf��+O"^x�>3� �|�#��p��s^����ԣF~�?�9�q�\�}��b_&��ͨ,v,��G[JJ$�B�RV:�a����>x��_|�g�d���1�����L�5�)8��ϑ6���M�]V:K�q�_t���[aM���R�&���P�x�M��w��Dk���5���u6Zb�d��js/��l��uoZ x�7�۔/�Q��g���M�,_XI���{܁zlL��ף�s�ӥ���A�՟*<g������֌�MI�� fK��v��*��]+od�n�p0���\��b����9I��Z�_�[o���FE�T����Skm�Q���c'�:ԤFi���xBڶ�:k7T�UFr?i&��U@�����5a����z�b7�_�2VaY�ܦC�o��f֥�(ĩ�YG&{O�~[�H.^V�)z*^;�C��3l���i5���6D_��L>u��GX��45\�@�q|Uz+��6�F��|=�6ǵ��'��c�Ҽ ئM������t�ZN�~[�����n�`i�Cc��>��NKކE�p���/@��ը�G8�� h�E�\�����^e��e�G6S<#!}��v�<)�bO�1ә�6�l�	�(�F�[���,7�!Q�/��ܟ��b�L߻�z��tTo��EW���$�v�hΝ�l9�c�L�bV��
�����c]0<"�����Y%�$;�͟���lUAϜ��R�)�߆���#F#�8�
���A|�f i��Z�lV)^��V���	֎G=�t�����������%�HQ��!�D�w�6��b� 4�5��m������1y&d6E�p�7y���N'0��}���ܫe�u�
�'��������/�v- �Y(\�����w��+I!A��b���H�%�e�ؔ`��8(zM��7����^~�M4���KMTG��k�[�'o\disu贈T f5����]�)쭺5�k \_�7�1;8���Xh_�3�y6�~F��؛Z��}\�!O��M�M���Ų߭��<��,����'_�&dr�ҧ��Yw�]D�bWc�i�<��Ń�~��7S��� G֐����L%.<��!�`Qa�u���$�����E�g�W�Xw�LQ*���9��Ύ���B�/-����j?�����o���D�b��ƍϢݍ����v�Ê�w`�k�8V��A��~��)�-���4N<��~Y@��B����}�6�d�H�>��*'Qz���X�*���Ж��w�VV���R1����p�`����0_�p�GEӞ�N!�u���\d4�⯔"[��98��@9�&�y�3���"]�m��*_�-Il4i�����Z�#�D��l܋�	�qryF<.�1!���%p.�"6��������Ǭ���jC�2X���y'��L�������[��7��8������~�py�5m�0{�?)���������jL�I\�v�9���}���hB�=�Qר5�['��v�A��qN�ᶾ���1WmO"�%��v
���#��Tϫ���I���c��ANfm!����l�FDv���5+�}b7��`�2�2����d+�M%%x���7d�w�	~x"S�m9�:!��ـX�����kv{���s�o���>Cd�L��+�kkCᅖ��H�V͔;绝A���^T3��������7�+�W��@�B�3�xKq�L��?����.����S`�>���U�Et't�2���� ������œ=�ɉ�h@��;�]���eP�Z�1Q��M�����K����j�"�_!�U|���oi*�l��%�R)%�U�'�cv�p��pfq�}�Uz�R�F;����<]�r�L39>T�!G�wSL��8ܧ��r�e~-C�j"��N2�IW�4��fyG���кJ�YDA9�͜�3��Ѩ���� �]N&n�A3��(�I0 K=��z�:�ہ֞��$�"�q9X���\��*��q�r.�=إ�_��U8�[�D}">���eF��(�����A|�<�T�$�P����ta���j!/��ˣ���2�?�Sׅ5}�Sy���z�hT�[��6'F�Ա^�J�n `�!�bⱂ��􀮁�{��@_ X���\T��3�b&�ZT�=�M0x�����"��V���q�&�ik�ض e��u��d�O��M҂�Ή'5<�[c\��	��f<��h��!wW�ImH�[\�6?C��w��"
Z3�M�k�Z	5�3��i�a\����x:pT��v=�$�j�����A�l��{%��%���eC�W\f ��	�P��펣��2�PuBkh���0 �7]^2�H��Ot
$���t;�1*�֟[D�L��h�I�Dz�-��~Aj���n6w�	�~���b=y���k�������z�j7�yN�����Ӻٚ�E�1�.�:�Eȁ�U���pͬ�Ǐ�$dfkJdf�����Sv��4 ��Ԭ�5��yf�p
��@Q�C����)b����:(�l��m8�:��*���;#�}A� ����#��)�|�SIn��!���U��*"�ھ-:P3��}��
}����+R�ltg_�
��nI��Y�����^���CJ�F @^|>�i���� @xy�v�+�r}$U:�eUZ��p�x~}Al��֚���~��("W�'�k���6��x�c]^] ]�kQYhL�#c솰���*އH�iJ���N���p���԰��A�י�,�m�˷4��l�@"�y#iT�q&(������FQ˯��dN~g���C^������ �&�z�ݬO�@y���5�����®���cG�y��G%_%>m�<�@%�ZJ�B��t��ۥ�����Ҍ���?���7m����$M��G��c�nX5��G�@G_��jŠXK���i����w���\g���i��������!������6�4��%d��/*@�H�wb��!����@�=n
4^x��)�}/_�u�ຠ�s��>�.�i���8;+�}�̆Hf@c7�V��yz�Y���4�]����7�ܕ�޷b�B��I`FJ>{B��'������ �'���Q/�'-���k]��G{�U���B���dYb��e�WR��'��~ �Q�!e���t��c�p�co6$h�G��(��S��\z�ª*Ű�F�����g�O�I���.a7r�j��hnf���3��5)<φ�V\vy;N�J<��<4eru�Cod��������^t�|W�_˫a�W6�i���/�*d��oC�Y�$����p�|R���$aM�Q��Y���|��P߶H��?-k0�jv�@�VMm��{̛o8D>܉��ٲf,�oSk=�7��~���Wxp�P�xp 6��7���I��_��Cs�Q�zdBB�n�0!��ϯ��J��sԂ?d�s��T;��)�����z���I|ܴ�$"V�&�G~ß/Y"<�Oƃ�>�|
#��d�{R������a(��#ݩZ�]
�^����8+.��:�Zչ*��n�Ї�Pm5�����Mxp1����-�����c�؎��j��PM���h�W8�0ŕ�k�/�^�����L�ۚ��8蹁 md��]�El����O�ZK}��B�fe_(�/�a���������s�t����-w4�U6G�W���f���g"��v�kʸ�l�Bh��]�;�:��K���von��q��S�F�${i.q���r��^U���ɻˣ��aɤ-O�3��kW���L��ſ6-��� ����)fU$2���>�u;Y㶲L�"�L�#
]l��g)u��ޫ�A^N�ۗʸ(f�8E��8�_������E2��u��pV���J�����#uAB!��s�d�B�e���P�R0uZK�#�FaX����S�h
�nZ1x'��yO��kUyN#��"B>����9���?�^E�m�Ud�d��$O�����ZG�U��+�
�?ޙ�kaY�{Ȕ�����­�a�Y��y�i�u��f�O*��:紅?a)Ci��>�'鉢� �]`��m�� ����ӊK�� ��hTpA.�]��z�("�ZTN�V�L�]�|����ȶ�\�������@�5���㔒��3�p��@鑏�̹���з]�P�ݼ���?�ƍ]�})�Kd��L�4t�on��պ���^�
��B�R�i����Aݩ�!V�GSjL���Z�c*ry�u��8�����?�X@�zp�� lxK�+z�tw�n�ކ�W�v;���,V֡��Q�����*akv���杪����1�1�h9�qV�E2�C|-]�z^�s��d�Ua��!�E�Q���7
:����Ť�9�haf�Yse\:ہ��ZJ�3e���p�IA�3�=M�.�I	��=��J�����9��{#��Xt.t�(���[��6F�����Uz!<���U���+"��}�
r���ƴ(��'�,kY��8��؜�I�b�k>b~N02��l�*Z'�Լԍy/V�w��34��� ���
��ؾ����q�
��d�1��P��-,�R�A5��=��-�IL%�q��ƴ%67��|��g0d:	�Ѓ
Mp*:���,7�Ζ��³1���7���W��A�OK@�%8`�11Lpِx��b2�%��/�ZS�D�����%�WED�!\E쐶��3�^�$B�3������y��h?'+xQm���B�7ė9ZLos�-6h�/��ٰwUˍ��w�y�q5��(���	92Хn�H|��:�!d�����u�;dUJ�|k���?��X���}
9���=���E�:i!b��N�OW�94�%�/�v�߫;�'ئ@ݔ���{�O�c1��M�F�G�F'��P�ፓD�G��fH���"�}��P����vp�	_(фI2��p����1�5ᪿ�d�T���k��2>F���_�*�*���}�$��0=�[𜭧k�k~{�
�F�A�>V��?A���U@��ֹ���b�@��Y���ؿ�*?����(o�`g(u?�#]n����4�m~*�`�7��ta�g[خ���6n�X ���w$�k���0^��ݐ�qk�Y��瀆�e�'�7�9ݺ�;Y���[,�<{_����.f�rt������U�
�9� ��F�� ��-q �## k-uwDm�@�F�Am�1k|���V��	uЈ����+X���ޣJ9��a���_�
=�x3
�V.�m�y��<Ue��l�����7^Jq�A��T�V��ӫ3c�X9lO��Z�/�\A!�>�h�����'�r�Z�^�P��Ea�8�B�]6Q�@��!:�i�#�O�
&�%�����K��̬��Gk�s�7��>�uMK/bɾ�.xpSz��Aw��zcc�M��xQ�:z��j4�_G�ɘ �i��?���4B��o�Q)��@�Ƀ���럟�Ā�H�[Oد���ͩ��M�MM�� i�G�f#��#A��~ۅ�1�|4��L�r
�K`��N���us���Q(�c'��d;�%�Ƥ��+���QF�@js}*���W���g%~���+ܨv�G�Й�2��w����*���ğ�O�x�b�V.�Ʈ��I���,���Hվ���>F�2�J oNߪy41�5����hV�\�a��:�2��}���H�����O��Cb\F��_��Vf8!��x�����E�����+���m�q=��)=U��L��<������~�T\��Vf�C�%T��{�rp|����{*�/"�%�� �~�`�)��M��/̩-����".��K�Ok����y��bA?����̼#��|�g�����GWa'b��0č!��qŔ<TrtPH��_�f,a�3�F��n�I���tv-�ka.ڟ<�[鸺f����X�6ڦ��<=���_��C�Є����N�{����L�2�|��eJ!d�E�%�F�kS'+���
�kym�?>6P�]%kB�7�X�!���i������Z�}m]w�|6�kG�i��*�1�V.�V�+� �,�e ��c �#4���hp?�`�g$��fo�eC�"C"9�e�5mY��P<��υ��8:"��������Ax��%�ݮ����g�\o�ehQ~�2����M{_K�JQ��`"�fd6r������!L<Zŷ��*�[�dF�A�)n�X
`��5I���,�7n���x��k��D.P����Ѻ%��w|�ww��s��m�����b�˧:�3�#s�L�����L��Ŝe�NQ�~]�&�Zgu�ѰI#��e9�"����K.�A\�;�颂ع�;�Jd��Xj/�� D����UԻn�'�yfO�ټf/�1y��BjxoG�WQ��%@��(���o����0�U˪����f�d����?��ȑ�ƷzN�;�Yv'�����}�����-"Z�iT�KP>ܔ���Sw.��;�?��@A^�����d��c����u�nw*#xh�X���Y�������Qsq���C:��!�1g���ԛm6ݍ�.	�njBs4ڡ��)
@���ᬌӽt���G�tQ`FH �O���LB@A�a.��9u�
�ޙ�H�u3m�n��X�yM��!�Q#$�=��'���L?}����7�q��9I�=���cT����\ʖCKVD,^%鈍���j^H�,�D�Kf2}�
���<xC &�J�>^L�-X�~&\��8��o�<��hOuM{D��VL�����WW޶���4&\�����o@�(�>����~�<�E�@FԚϰ�~�@��(��k�x�2�����f��N�Y�~�;w�h��S�Y��|�q�g�0n�ۜU�
9�H�8v�;^�������4p�zqʴ�
�h�1��MS��~���uJ��&���,+%p�)O;�x��חF��w�t9�@���XD]�5�i����K-�2���?�nL����]�^a�\P�H(,mW�Je�V��������s��/\�}j�xLA/�� �+(�yB�w�b�H��U���@R��A'���%���0��\���n�a�l8����e^��-.H�aD�9�3�#��*ט>�C�n���6�q�i���I�uY�C���?CW�^������*̖���Nr2������%�~䪸�0����a�9����K�`詌J?�[�]�MT�f��:²���§r�J�k#J�.���čÚ���U�X1u�ۃZϳ>�^��z�ޟ/�
_uu{�u�����(im<^��?���<T�;6ƾr�ifV�?6Lu�H��X[�(��yC- 0�����,�R�A���6"t���\~�˖;��M_�9�q�%Y�8�69���~o:t�,]��!��'�� �U@rU���|9UrF��j)Y_� qwYG��ཹS��S0�ՅWw�q�vj��p�.� �{�N��L�03�i��sW<�$Uw�|I��Y��^��K��U�������jw�Zc"��;]�ђ����V�^-A��0U�F���X�WK�53˴�*oܬSӹRYt-Y�u�՘��N��m���:(��_�G;�=�n�P��rv�~�O�� ��]J--�8�f��ܶ����n,�uRwr��+��Y;�[Id[)Z��#X�����՜�{���ɼM�ΐ����л\�p�{��IƚΒ�W���4pr��7ccBN�G0��C9��o�#�_(�y�!�l�E�s��65MZ>1��Y�pP��4��H�I�oF��/&+ޒ��e7��X��O��o!w���N�\��"���yKQ1�8�SX�3_vy�B�5C��;���-��ǰ']�FOt�h��<�=�A'�f�ɩ�+Br�b��OW'����ђX��o��e4]L)T����tb�����H�3�i���+�H���4��̋I�H����+8!��>!���E0)"�<��^���V�5d?0�(���5u�)æ ��WcW�ȰN�iS�ݡf��-}���{�dF����e����\�L)�r'H�|�	�[���U�=M�.@@:����[���k��ڒ�8�,R�n'?{�{"����+�d�-�S[�5���K�<0D�l1�xZC�
ObtJi���A�'�>W��/WڲJ�]�N�y����C=��9,MJ}u���G8cX�Iǡj�p�!=�נ��[[�����nNj�QB���L�ހ���:�.��Y�zF)f��ƙW�[�k�k�G��{1)~x�0[3kŦ�uL0e��EO+�gm�]B�p.�J|�ƽ��o�1e��]�g�n��2�\G�`�{�u�����٤���tق}�q���xn�q�<�WB�����\`O��r�"qP�z�NAUHV�M�@�Ι���p�!�������{��l�|H�aj�d����w���z�V�D����5&����e<K�0�"��*���j5�����[�Eﰘ(�l���9+Apآ ���MC�&��+N�v;����7fGt(��ү���P��{9��ɖ�}*לB�.�����������a�S:vbC��`ܛ�qw EAL%�}��+��В1��/����	�S"�����z��=��-��������yd�!�n���n_T��^`�	��ľ����]?�q�¨'oѲ��K��]}�I�����i�����(�ߛ�瞅�E^��u�ͱy��t[b���-�QU���-�ϭ�	�!�ě�;��ͪ�����nN���o�0�� ]�l4*�D��-�5�nCD,/Z[��ŭ@*
6�Y	!v���\L_c!�PstU^��|�5��"G�L�s�{R��k��'�"B�
���'~�a�%9�H%�Ó��=M�\=wA4ZQ� Z�W�|�u9f���Ct-(�:������8[$K@�������X9O����QƱ�v�����b����T+�(��,1�&Ez7P��!�c��e�|�E��j27�S��k�#�*lb����s����\	��!�=��iv��wzΣq���{/��6_b�b�,�<�7���bx�,:�1��B9��k�Fw�Y8� CJ�����{��I�M."6�x6���w^�|6��r6	�q��j:�2Nb�t����Tc:�[�O%���W@=nK��*5�uSϕ&c�U�-�-��ilY���յ8H����^�$�G�cV�O'�K@��,x�y�,���v����=����%ķ�� �>���n��?�X�� "�Z���������<�ݮ�:��nA�?��`���@	��y|˹���j�qK��C&"�<��%/w�Y(�C(`'n��Y�@s��7Q��6�R<!�=������ն��`;��b!����8v=a��om0�q4��ԄD��>bGE4^り���y/�����Qr��ZoTCp�!׫��b������9�EBT���Y�ߊ�.�	^�LU߿~<�k^X�T�FU$��a�	G v����5����Α��vN��W1�-���k3B�B��1��dQ_��3�����г8T��נ����BSX�w�yN�����|�L�1��5IM��v�O1�H��r�|:o����K?$��A�B��n ��h����D��xf�?H�"õ��9j���w�:9k-]��i���S��z����W׳ЀxA�t;oz��}�5�|lt�-vB�w��	,
wpr��'�ڢ���������*.�/��m~�4��;��5�fJ���N���f��?��z���v99���rˤ�ulƂ5�C�.ה
��&	���v�ˏ�0��P�g���t��eo�!T�z���|�Ԩ��K%������%V@-�*�-�_�8;=�oRI¼��K���:n)��!�A���f����F��_�e0�9�¹��>�(	����4y�1�r�^M
v1)������|5YM&g���}@�u�>�S	u���@�,���T]^ة�7����]캡�S�)
����]�w��B/6*��}��
���w{K��j	s׉�m,�,�C��T��̛��{Ոϒ˴�M��+O�T����i�ngR7���4M����y���iEw�/5�p	������M�zC��|@nHm�jL��N��*8N�Z)}/� &���<0�*Qf��Fj�ᑷ��E���)��S���6�N8�{�$����RT��qu�󮩛��'�m3�ȧ���6����<�osXJ"�C�&�yJ��Z�g[�nJ�r�f�?*�a~r�f+��6V�X]�gk�5��+zu���Q>;�~����	*o�;.K2��w�?P)/�Q�4��7���~Aڍ���)�?jn�?|���y��=4^�������<��ª��GU]��C��/�q਌�H��c⴨
\C���[�ǋ��u�!/v`:48J�w��}.�]#fr���{8Gw%(�
DQJa��w�-�Ľ���Y��P�א�`��r]�� ;�k\�<�i��5YB�[XS�co��^ �7����Xr;� �EA+����,aEX��@A�E�/t�ޫo�%����h�����K�偽O&��8!-�^����	`&l�5�+�{9��0�$�x���6΅��d;UJ�N&��c����5Y,ɲ;n��B�Ԧ�w�vH�$ٰ,s��`+.��J_4��Q˱U~f�s|o�`hX���5�q��.���O�a��R�YN�i6o����S��u3��jO[�K[v@�`�;�^�:���Y�@�����{�R\=`ٔ�F}��,��Gc��B1�H#$z��)h�!��B�gܻ4�$޸T�ku�Oӑv�4ߐR6���f��FZ?�ӯ9!����8�P�����i���ҴmZK�9�)�<QU��.����a��;Z�w_h6��A�K�w�݆���Q��E�\_P�6f��/����I;_��Y�՟Y"x^K|��a�KU�ޕ列��V��;�	�	\Y�n/��?k����?��{�jǂj���tV��/�rԍE�ɎpBÑô��~L�B�._�+��Ȟ�������YUE��\��#鈾� �z&�Rl%D�!F��+¢Ŭ����,T�YoNKi�S�������Њ.']E0n�i82��
�8�z4��1ׅ�3-G�`uW�^���o꺙"mO���5c2��np�o�yd3�y������Ɲ�O�`)���#��;
!��n�f�a����c���`�.}ڸc^\Y"��8Q�A��$N�"K<�t���ޙEPW�.����^�>��}H���%�$YɀW���!`���u��XlJt�@A��3�i���=Y#�����������,'�q�&��N�*������N��?0\���z��&G�H��{����kS�m���l��&eI��Xcbj�wF/��-2�UuY�CW������!�6Z�Ͷ���]���xY��	�؂��Ra��:�fAߩ@ɺ���� ��%Ŧ��1��*�����R��K|��=ҩ1��Ms�1��2�=�Dp��)��sS��OSi�N�ܢ��D���&
�%���T�-��Up��V�Yi�L�ԅ�H�;{��$[U"͟����d�3aS����|�u���f��춠��>8���܉����E1��5��w�Z�)M@�*�pZ� >,�qr?���m���ك���`Fk�Aqt�����o&fg�sGQ3��[�|��T��w�
�+0�=5�_�+����.w��M��}��}�H|�A^�s�-a�-rU��)���/�ޏű%�㷮�)�X�8 2Rɝ�>��ح�s�%~0B'f���6�Dȼ�SW|EC��o�6�q�3�KN�䥞�0�q�(j�#�-Z��<�F.�E!1��а�� �k��47���~Q�.p��j
�']D�B4&�~X~Lo�D���g�+�%߿�6A��
���m7��!��K｢P��5�	���Ubhx���d�hy�4��΍�E/�.C�,�[]W���W�^�vi�u����"�dJ��	s)�kcN�G���xaJ+��s��Ӥ��~��L�vy
,\���s�/h*�ugHi�D�$_���vӖ���i\���r�X��r�ܼc���g+��ji�S"��YlM*Q|���ڑ��;œ��KT�eR��l|�?��wb��EqQ�jn�XT�~4��"ǡm41�Ǣ��+=�
9H��O�D��|��x�����T��u�wId����GY-�'���JK�(�q�7�0�`ڶQ%��\��;��Ap�K�j����
ʢ��7��R�Cşơ���I�P�9�p֙�,�����i�s#�IcE���&e�%�-7k�wNr���#�4��ⅾ�����M`Sb����_G<��������td�d
�A�ۗ|>gN�U��ZY��ѹv!6��ƅ���8����$��p�.�kᮜ(j�6����++o�h��
�FT	O$j"��F��p�c]�[3K�R�үO����}8Q���E����Au|�_�>'=yc���-���\��Ȫ|T����N�s��s�������^��F$FK����#*�!a�X�`��S�C������/�ݓv`P�c�H���ѭ˪�UI��G)v!�;�W���h���5�6�e�p��\���tTʖg�JA�M���C��DM*8��ٽ����6J����U-�����I+͖W���P:�d!]
��x��$��6pŖ�dꈔuM�c[����J�� 0���( �5���]�j�C� �7~���u�/7�!��<�X
{"	�ؠrH��X���US�@�:���/���诐�W$��PA�}���t�]�;p���*��_]��U���������G��Df�>�"g��{5fbT�Oψ�rI��'4�&=�y Wu����2d��P���s�\a��dT��+� �" ������1i�7�JǠ�4`�T�5j���Yf��.$�M�H�M���Ɍ�d��t���$�?��\���z�v[%م��K�EN�ؖ���7T�T�Ѵ��Ӵ;�����S=�{�eY&�~/T���ѭ�"��v�d�,�m��*'���>ɻ���[N��`�ݩ�b��T���!8�#8�i"-��)�7c�A}@�6� ��������Z3Q���fGP��g.`[_3�0I\>8r�~�k�e����`�,h!c�D4�WUӶL^�+x��A݄���{�9��c=v�ł���zo�'�w�>b� ٞ�,�FFg�h�td�F���h�L��ߡ{��?�P"K�TS�/������2�w'�4�I9σQhd���@ֽ�:7=���p�q(���n���[�����Z����E�o ��J�_�Q�!A0�{'G��s���c;��	NO����*��0F�Y�h�	�`���3D�!�S&�b� �T���}�S���"
���*�"�h��o�j��,V�,���$}@B��$��痍}����hsʫ��P��9/�;�pt��m��X-a���1���nђd8����]�+	�W�tӷڒ�$��}Dk��?�������s�������eP�<��_�e	;& �e�� J�b3U¯���o��5�n�zGS6�� H��"Ч�#:+���>���i��~VuA���:4c�d��0jN��D'K�)�(&����5ٌ
Wl�E�@�<�Lb�?��K�4�;#DJ��=o��p��5�{�/�<���vi�>?m?MBf���Oj!�����U�K�D�H�3W�����1�������M���Ek^JC�6h��>���>�+����)6���sS�Ă�)<vs7s�|ɨ7�?����$K�qk�"񵶐J���t��D�
����($Q�����M殍F�D�%����n��.a	�z|lc_#]8��<�(J�P�G�P�`�8#n{�C���D^5�<r�Ba������f��eUD�y��[]yÇ�G~8V]L����B� y�6�_.�-n��7!&>*�{�$�������@y e��1^��w�Bu#h��.`�K:�?B0g-����be��~e	1���iｰ*�h�m-���v}�4M:�4�q�v0a�Đ���������"�k;�������a
��֊�	[s_�u����O8=��%s�J�7����(��T$b_`IH�2�H��J�m�EK3=�r�n�X���K|� �鑸���溋(�$�uB�x|7f��M�"��5j��~}N5�����DƚiF�B��{�{��b!~T~�g��(��T��tt����h��q!���<�v-�YMfn�ѼE�eT�
9G��a�ɋRSB�+N"}���!��2D�Q�]�XZ楙�ѷ�����6 ��|��C1�*}�=�̻{����$0i�>.F�Bb|V��2|kI����d���DF�
�uO&G4�]�XkL7 �e�4���%"�ū�:�-�4�O��>��� zה?��y�[�Y����/]TVA�x{8"�3��[�2(��NǕ]� �N���=Nn>=/k�,�3:�>k��T�*"(�3�#H�~s���T��q��<lUV�	s{��]A�an&����rgka�L�8�����q�Ҷ������O�������`��n^=�����ι�`��J%:�|�β�#h�V�'���?1�.E���n��TX9�={��Q���>%���=�w�⠳~م�_�={0(Lq,�݌����Й=��2]q��!K$�]_��.}wVb�f�̖f�6s7*������Dń@ݟ�*�d�6,������Y:�{���τ4C���A�e(I��u�z�:+-iVd��jk�R0wc�tْ16��~�����(*���Hz�8��&I���-\���m:�,��_u3�Y1��YV�*��a<�T�b)��'�@3p�.��ʐ/Ը�a{��,/F���	<�� ��s�Л�K��1�@,��Q��c�f�%y*E�y0��VyI� �>@7�v!WUZW�_�� K{�|��F~��%�z�&YFW�tNݒ��Z�|^��D����x=�%���D�0'o��ɽ�i����������;o񑗏$��w~�Φ�Xk�#	����S���D)PG�d��8:��n����a�����y��Ga,ȸ�Q���'z?)Gx�ܛ�Sv��;��E���'ĺ�]���z~�(� !���{4�z|�k�*�Q��ix����(�;d���#Kk�����h㏑,�?trˣ#~��*F6��G���wraH�c.�S>X��L���y��-svTi���jk�,�v��i{��X5	<��E@�:�ď%/5a/M��mޛ��s�C8@�Z�7ў��E����H
����F��Y Z�#S�aT�R����\,)P���Y?�&w�\x�b1���II�|�9���٫�E���$W���7����H�țe�wH>�2(?����}�G�^27y���� A�s�����h�O?B�n�B�j��m
�|��[k�
��{�b|�\{�L���o�� =�&1(S�x0w�dpz���o�{Os�[��g���N��̹�!���u?��I�K �}����]��	e�׫���p~MM�~��do�� "��N�Zt��}�����f)Z���g�c��Z4���L��d��R>PM��t�,G����3#C�ꦚ,�ƹ!�׉j��[�3��(��f��kwTZ ��FX��!��?��~v�牮w^OAg��B�Fr�Vg�}>�\`��@B��ޑ@�VP�>�dEk��^FC A�׋+��Ӊ��z���r�+���r��+�%��W��
��w����	)��e#��a��/�F���3���H�#8ߌ��rb��<|>Q5(�F���L`f��um}��@[�����Q8$:��F�aIE~�v���;`1Q�����0���~���g<�0RiW��;��"X'�r��pu;$	͜
����0�?FxI���i��'*�]�|�.CY�����f�%��2DLu�f�z5"��wK�,���]4�����(o�p`A<���<�+��	�+����iq,^�\`���������:�����}��dVTȚ�
6T�+8�g~$d�?�r�
�C+(���/]�X��C�4L���Jᗺ�\mJPs��	!�⳸'k`�.���8	�lqR�jYY���ҍ���Q��o����)�`m�rH�!]ƀ�k�!��:��MJ���b��(X���AA��V ���3��W&�+�?x�X�������#{.%u��C�Ь��?�鉙���W}�x�&'�x��*�RG%�����N���=:��7�(���e��MO*����$N��X7)�q�{��k�ӷ}t�t�#�jǖ��	s�r�ӂ;�U~\����jw��,[�x
�I���=����p�f(��� {�T��c�I&IZ�Q6Pw��E��bpO��#�┩�F�:��J�O:�NM�^k�8hk���N���>"���&�-4l���͢�w$��.�BwF�P���-a�0�i�xX�x�1���1H�,
��������w����6i�@�`?cSU"n�1o���x.!]�P2;�[��
g�tV�[)%^�q�F��ޏ��
�o±�)��i6��^�����n�Mp����v�6�}�6�.}��y6��;���¯MQg>m��2/l� �v��#/Yl󗏨����u�OB��
� q�C�A �k'8��/ٛh& $��=j�5%��;��9��L��n�S�|�G�����.�^�6e�1�p���
����d��[BX��x�UYy�@Ud��煌J����HPQg+�<@ǱU�����i��&=��~���Wq|��-��#fX1e�;b:-|_����ёAC���TL��M����@A��`rmno���:�R��Y��A<��e�9_o��D��r��z3ӟ �c�Q
��\�jŚ�ji��jМ�G�/9VW6�����v�u�G�;��[p�w�@,���|w���~���k�6�e��}6�0W��rSn���Pr[��;C�?<�͚�[d�}��P����2E5k�N����l��{�U�-:��c��p4�����_��l�-�;ne�&�;��
gO>����/&ARL�Ȯ2>�z����nA���\��L�ZD+:|A��o����	8=t���{�{Ţ-	�%OQ�Y�Z��1Ad̖�$�!7`�sS:a��9�"B�b���j�gz�y.�;��0^�+C�sX��C7�F�줞Ha�Z�pw����b.TJ�y�F���=aY0�XX�4����ȶrQ���*�Vm�I2�Ӗ2�=!wpU'*�Dv�T���ꦆ�*���?f
��ަ���6&�-��y��zB�9+��+�\��q$�jI��@�R�v��P�)�jՉ�?��H��O_0���iq;��j��$ܾ�7�=h�>Bs�	.Ks�+�.P-S�a�F_��2	(G��5�>�aѓ6Ci���vO������A�=ќh�ǘ��@�	��������������ݑ������+��N�S�X#�����e,Y-�!o�BE���\w@4=�GK#�g�Z �+T{��(�?�p8��3��P�|�*Z�H���'��ؿ�_�z�˒�?�~/ƊR�Z.%YdO�H0�nd��I� t���cw����|�&3t��^r���d�\�p���Ԉ����2�ǱW�}北w�]�L�c�F4��(+��l�@����2��:e��Os�?�Lc�`����e��6R9�	�����EC/�הN�wCP�ȵG�̀h/(�d7��-����0Ȇ5�wv��K��P�F����Xi�(Yxr�Z&.�6�1�*�U6!g2�����P����2p��y�)
JVm �EQ��y�f~��-f��~f �HU�hzL�<�GdI~7���%��s�kC�qq�Ο�\���89�?�P��sKo����g����K5�ֲ�[3�3!\ң��̋F�;[t�>e�R�2��ۻ�g��i��<�x�n.k�c�����e-��;�����S5�����ea*KPoA����hn(�ǿq]���～����D�K�아������,�7㕲�`�&���k\�����U�W�2�PӁ��G�h(>��5D��x��0Rk�����No;�)��T��x�%�դ�{���u���I�J�C,����"�׌�Ss�����|091	�b��h#���Q(R_w�ֳ}2=���R�p�CH��E���t=_���|����^R���M���RƳT���48�3�U�����i�}���;�)�){�B|��KXeӻ�J.\�t`Sp���.��D�b4Ԃ���/�9��"
 nq�^��I���m�@k�&���.��J�$1y �\�#')5���a0x��=�:3ܭ�t18����u���2鶽�p�����Vae?2�hf��
� �oz6m?R�.��s�p:nI�`������y�`n��ޤf�w��M���������S�'��e#����aV4iiϡ�X?#��t�Y��vA�]�Eh�
v��Sf��^x�Z������_|op��,�K_I+�(��Zd�sj�ԟ��� l�g$K�)@F2�2wAe鉩�y��?F�����r�b�������=I >�l���:�#��?���)5e�x�g�վ㡌��E~��G]A��Lwgu�ʛ�V�f�`��Q.LDǢL��ЧX�$���"eD�F�AP�
�hS�T��VCAU������l�O�;u#�0�lZ6iu�⻏-���4u�"�`�0A91��Ӂ�V_Ia ���7Y�?���-v�������@���)��Z�� c� �4Z���.�4/OK�q�|�������ؖF�]"vJ%nKz[��@�x5�oYb�t�Yl�.����R&xԺ��4 �1Ν��>F��ɿjf��#�82A�-�obЭȲ��ݑ��&ߞI�l�ۊE�>�Ƌ�Xȿ�� ��1���h���� �����=��aV�''�Ԋ�W��%�c��Gz��\��cA�rVT	�5�C��H`���=~�f@��������|��g�z��#���n�Ԕ��%�	�ּ)�����ȇ�*>	��f��.ና@��Β���x'홺z}Ԍ?�s���: �=*+�=э#L�� Mlr&:�?�����a9K#��}6�Bt�%(�:��~�C(#�k���Y�\�k:x�NP����� oĤ�n"��E&�d��b���|iF+s��\ؿ}"�Q�>D8������B_�t.՚��<`z��)߳��_<��]��7�gr�šZg������к���M�����3�5�g#��P�~3�Θ[�o�J�@��:)H��"��/��Z���ݯ����� �MX8�C��j�6����Z��VsD�ZU2&{�ػk�`+Ƶ"��iTYbbI����M�
{�!T�[$�˃��ӆ:b���0+t��g+j(�p�z�Lk yd�Rb����y�na~�����{
 ;\�ϟ5�S�t�W=�/�2sBw�Ss9��x]#��p���&�
�u�D�6)��IK[��Y例�<���[�wȚ�WJ6ri�oy6a�l�cv������� #�V'u��_{7I<��ҫ����Lo��B�a��L����K\X��e*�CYe��6��-��d5�� �2��E��/����4 �PY�'vƍ�P�H�;���+Ԙ$���	��چ�>0c�=�\����w� z���:X(zu+�
9��G��JF�2۽���f��ȟW�~��qW@
u��r��	
�1����B��/by1�OZ��tjӎ�K�}��bfh>���Mcs�r�8��ż��#���,��%m^������~۵�]:q2��lJ+Pn��T�>^��7Z�Z�!�<�}�6�w�^g�%s�����s��A��V!.%lK�!oeE�ha\�a�/o�{{,�/�M���V
/��==t��d��;^g��Y������_b)�uDtj\�|��k �!~���U=oe
sI��@��>�,�6�
pn�лG��(�QJ=;>�č��� w*�>���%C���}�G�L-c����m+	�P�[*���f�����Hp�#�B�Ǿ|�rѼ��J)��J�_����s#�C�ZF�A�*�S`�k�C�-���u�c���d.R�L�����u���+`��ՔiG�������Xr�!��D)@��K[�������{�M�(���W�g%OFu_�Zp>���7煚���ݱ��r��^M�:L�j���T� c8���TM}�`ѹ�r/HKO�������K��*EZG�pR�mg��$>HM�m6�d�W��kQ���r(K��>A?Kݭ�Uɋ�����%Ԩg�d�R�qs�5]�S^�K�aO� w�e������Zj�| ؉O�Pˑ���ů��&<�E}�b���n��'�HA��HQ	�������m�mX��^���}��J���/ ��ۃ��ّ��}6\��.W����Eb��NǼ�H�v��[����}9�§q�>,�����R���X��B�[�h�jO�o�^����ӕmr�cd�gD�7����K����Ҳ+w1�����C���X���j��XDw��WzV��]��3"t�����U���l��(���RL}�@��5�^ X 7=��S�f�E����EF[_��7�:�w����<���տ(�oZ��) �c�ބ|�(	BC&A��{kr,U���+� ���v�՚N��9O)u���_�&㹹5��q�N<�rh��'�A�����Bi���CaX��ę���Mi����p[V緟��N������*Wc�ɳ6���SL����+6����|��C�:i-������u"b^�h��)�,�ͫ#0=E`"��̃���Q���Fh��l�v���9�����p�%�F$r���by���U��&��6�M�M_6Y�ǀ���V�ii�r��r��:���M*��u�5����wo��s}�E�L@����:	�)c"�<�����m���@1�9�
�������`#�^�Tٝɯ���΍x�mK�dJU9�a�W�S=W�9��@M����O�]��`{A詸�2t�ʽl� s���YB��\�ay%��ԔA#"򭤵�;K0'&Р
*�ǈ��Y�!�ӏ�V%gj=F��)�1�y�QjQ=�:=��X�[`E]�m�?G5<�Y��V��f��������2���摒T����_�D�!5�Ү^��[�>.��7~㌴<i�Kw��2}T�KG~������Z��[޼F�tX���V�gX�z9~}ܿS�Ed'��h��������q0�ۖ8�!�=�C8�r�6����09�/EZl�:b���T��\D^�%0懢J�x\�.�|/��w��{RI�Nu���yH+�$������j��I�>F5�K�8��%���h[}"Y{��1�0R"��a���M�Kr�CA�:�����(>�r�GcF���w ������fS�<hӛ̈��^WR��!p9�[���LŔ:�Y��5���@M$�Ʌ�2�ܲ9NSƹg�E^�uW���v�W����\�15��0%�!#E���qp�#�d
r�P�%�=��G��]���ʺb�Z��Ec���Q>U7N�:�B�Pxt�(�a� #y<�{������(�>���ɻ�65�7=6%����q� ��z'liK�8[x8�+�c_��eG�:%9	.>@�[��-�>��S�u�7:��� G<Y@������Y�o�A���֓T�ia9�m�{E=++����c�·z�ך��7x�ċv¹�E��>��k(M��H�H)�tr}�6����Y�,�.-,�8�=W�h�(T��ʿ�c&�·|��43�����]��s������#���/p�v���-dB����kz������
�g�+j��!"F��ׯTI.-�ϼ�����rӀ�϶�ݙ��3�q�!��xR?�:��O������t�����>-���Z4)�jb���I+&��[/�?��߫�5�W��§�E��l386�Ax����(�׊;��É��Յ}�]�z����d���5�o�_S��f��.A�+���gj�ŉbt؋<����@�8Omy:�-:���s�)](W���� �Y���N�6��:>�J����j=����h갅'��P���r���;��O��u��G�pj���{�p�@�m<Ix^q���c���Hu��H٣²$Y	���`H�[�O=�s���lNu�+�v��"�l�n1�Ѹi�j������ ({��7g�1q�5�Y����`�8��0VvhtU�Ab7͚r�´e��AJ~�iT��9�
��ؽ��W�xO�G��D�iS0�@99�uP���B��%�g�;mA�Mt3����������V�1ˋb�^N���/�v���M����1��2I�)��e���&��ʼ�|4[���v�_���2�Peg�}]C��=bS@�vː��/�*�" &q�d}<jXeEi�uŀ�A�75g�]�O�Q����R$4�0�K�	7��&<�6��8�~���D��5��8��s0^c$Pt�Չk}���Ǖ܃r������`��4;	�na<�h���F�n�4�[��rV���I�ƃg읆�����o�������C��*�Fh2:\�mb�)ꈈ8,���ӭ��;~�"���Z<C�|xN&�q���X�s�R*R��-[L*v�o�N!���њ{Fb��[�SM��O ��z�>�Ĵ<�@#����I�r�O9��iE��]%l�D�|��a ��*"��^�G�&�ǆ1��ẕ|����k/���aa!T��o8^!s<~�x�
̄ŊY\�23��fv�Ӓh:Z�k���3�F�R?#nߎ��G�O8_-��<��d�'����	-�����
��s\|��U7�X�W��0�bV#�%!g�A�����k�rw%-̕���)��6��1��*4�f2��V=�*)uR��}I"�I��W�r77~�Z�=m�U���"(�/*���:��V=b^���~��d=�\�V@)q
�.�O�İz~t�_3���Z7�������2@�������uv'M��}R�l�4He���.�SV�<'U��+M���7�QE�m2��fZɉ��[3z�1��'�Nq��9|���<\bn�iΛ�B�]QS}�6Cl����9�j�}�yS��W��*}	�����Te�M\C���yHǭ貥�����fh9����9��n}��?wXT���1C��ສ�ڇg#��Z���M��˝��kV\p�=�~����lx�E�)&Vo�����>/~�c�>��1����b�fͼs8kx��SP}1���Wlr�C�0�i-*
*�h]v�~a0!k��54�#+h�0M*j\Ý<����S'Ԁ��<�Wƣ���#��_iO ��^�Y^��*�8ᕾɝ�0砀�}C�Q]F��9��尮�Vg[�,�)ZnSD3�T%��<�Oqɕc��t�qw�{e�ϖ9;�ۉ9oQ��U�o�+��g��^����/���1���:�Ơ�sf8�@��K2�0��>��r�"��êdh!�mB��A��(Zv�
n-h0w�C�Ut�^-սH�v�f���������X ��7���ԕ�����I::d͵d�:h-��a�,��Ra���vi�g��[�e)�7���ߕɉ��{T�jo���y�b����6#��\�n��H�a���O�,4vSg0�	o�V���C�q��l�	���-2����i�Y���!��g=��z�5A-�"��8�_'�vz�N�E�:�q}�[0U�8��C�^��k&�G?�P�[l��uPb���O*�^��s�<N��(���LQW����$�!��`����i�z�7��J�b�����,J��B��5٪T�����P"}���,�m{�k���d��~��S�9<ѕ /ED��oS�\E���������������'+��:�n��$����LCR�pd�ǭʱ��[���Ԓg�'>�r�a!7��ۅ����@�6�6A������)$#��/� ��;@^�6�O2X��^�v��,��/}L��s��������;�\yq��[s&����̨���l�>[d�w���]0��&��͟KV2��z��Д��X,�4�)R0�͒���J��v*�荜2,�W։�I-љ/�᫧9+��6��pk#O����N�,\���{
������7�U1��S��)��wM֦�ji��S���G{M#_��E������^�ȶ����k2�)�?��V�� E�s0��&ex��a��V�ވo��!!��~��4�j/����Tȏ�� ��B3�i?�Sh�����r���z�i��n��r�J�GX�� ƹ]q��#�m8»��4]
���u{.1��q�4���`�u���F��[���8[���|�]��·���X��?�j�x��s
0��oL�rX����ְ9����O��MI9����jʀ�_��-79l���D���XZ�jՍ_�x�"���^������pT��,ZPC��Ĵ�2���$�,�K<�Ԡɽԏ��a��NN��u5:�Xϥ�FB�4Ix!��L:Ե��[�G�����#1��3DC.J�	�LI��Je�h�V�O"�V�t����ƒS�	
	��Ct�$wM2[_4�3rp��Oek�I���e{C�\MG�,�%�� �5�e���]#)`��Q2����3��N���[J�f�P�>�kOe3)��z����]7��S	A�;m����ƻ���ͷ��Wv1@8��
��Me�<)���$R��ÿ�l�ة����h�ۏ���|y�5SW�w����'"��Ӵ�'A븊���c�:���Km1U{��D_C�����+.����1U�Ν�,�WV衝�����$k���v] �)��I�A�7�u�g"��� .;����S*T]�ed���O����ӈ���� �Pw��o�n�L+��W#�&�Yg����@�As��f��/S@"���=<�7��Բ"�,t��o��b/�Ǹc85(�h�����?��� �Z��W8���ԈnؤC�}�L�� ����q?#x�b8(�[B�@��!G�3���$��{7l�F۬�����2���� �p��9l��D��h,������	]hS1�T�=��JՔ'�1Y���v�!C��8����%k�#�	+ɛ�8���Q�@~׷�|!fI�� �ީW������ԥ����aD|�.�e���S����y�9i��8׆�*�Pw��xrVLT7�II �!���h��J�P�6sKpMt���Ɇ�:7PՀw((Y-	���|)6���vܜȎ��~��Ɣ����ϰSm/Ґ�E)���^��T�m�B��4�X�e��92���A	<6�ջ���
�M��^��R��m�.�6·���X�H��(�(p�ܧs_�\�2_�V)A��d��
c+��
�VA;����d�L�=�\G�q�,�:�`���ƚU�߽x��#Y�;��]�b�aIڏ� 5 �zr~�/d�,�n��A#���J��Iփc�m�4#�E$h����RK�#����d�C%�U��7�b���1�n��6�;��N{�16ia`��Y�dB^-NW�X�ý��D݀�/�6�?ꋄ����a��B$R�0@YH~_�g�ަ�԰o{Iwiʘ��a��ts$�a�pJ*\� �$���N������J�KLK�b��I�����ڮ[Ö���o�����o��� �4�:�'[YA>mG�����\���R���bn��&]���(<�t�UK��:��R�H0��ؙ��@a�$�����s�
���f)����@A�M�������@���MHc܂��[�v��(0(��x:�	�6��HJl��>շS�I��It��{�Z��Eq�*��+/`���NH�6��M��e���5�[��Cv���%��r�ɢ�����Xy�\竻I�(wu�R����Ԇ�}L��K���h�9ޭ���ٔ�o����,�jth�R�!�ܭ�2=�Y�X�&�t����xE�V t��
��2xquz�� �q��L������w)3ݲ���X=O9}0�)BK�ɍ�Qz�Rb�~̯P�y��j\���sH��o�M0��wb�}�ѳ�@T����E0��R%�Ɗ��O�nȺ���	�a�\w��8!�_z���'��CN��!�%C�fGm�%EX�+��T;}��ɧ0Rѹ(����Q0L6z�l$�'�ڢbg��æo9\�����$v�I0+�PY敭e,���O��Ԅ�|8"��^"��i�������V�kU��'=o�{Y�e���j�=�ip��0�L���{�VcR�z��l�_j��i	�%�
BN��j��D��?��%If��%���P�(5�M�� �������V�g`�X�j� \���C�ȁuԼ6_.ʦ`m���s�=c�z<a䵠YJ��o��d�E�>�X� �I*l����6���)La�h�t�M�a��h�E����j~��M PE}���j��JF��	�$6;� ��M�l��۠	.H�d�PJ1�6�}�{@�X��T����X�VO���+2o43�i�a��[	�W����LJ�l��cPT��h�r�i-/)��4����9j��/����x#jb��QoT�N����hڢJ�i'�(e<OgS���̯���� �6���Z ��ǆ3[���� (�s���l�:� _ϣ�E[�r���l��Q�L[U��b�x ��q�)_#���!8Z��e���Զ��G۷�H�(yc��S�P4�� �������"�`kpM�O�	��н_�0��3s=���hq��)����d2����?ͅ,7(�k��#*��wF��* ��í�����E�wJk˽A%S!�D?�ȡJ/^�v�bE�tV�a�,��Q�j���p�O����rëU;a��~C	3 R�b��PN���	�8Fd�"�[/o4IE�k&�9$�H�e�	�]�{�cMy�1@��6~;���m�����\�_�m{:��f��[� ˸O��>�[XE�dS)ܮ{U���Y5KZ;̟L�=;�M�}��L��/�,��[N�4
�T.��+L�)!�DrIf���W�/?`TU��Y2b�s�{G����/��F��5���Kc��o��
�H�� ���e�sFR�i$��8!*��h�UA����ޱ�f*ӝ���F�$���I�Ur�BD�:��Sa�3<�j��oJx 2QͿ�F;�,��%eKK�p���E�9F?}��]�,`�(ڭ~��|��Y��P��^�I�H�m���Ͽ�%�iS��2V.my���d�����ok�9)�
����5��kI�A�'�	cJpĳ,C��-e2���":��1�E��ȱ7n�Ep�,=H�oX3IS��y|I�4��{��s�!@a+�՜x�Po��?��Z�Æ����l��htù�'t�qe��,n>Bz�M���[>R�8�T�'��[�����OΑĀQɂ�Vv���7�^���C!��3b��H�L�Q���&�N�9T}De7�uv�ex�����q���{� 4�A�\�,7'�k��r���r�̾�9���,���F�?{Ip}�B�AHFSs��u��#�&{��Yq��i7EL�g��2�T�������(F�pk�� ��_�Şⶀ�2X
:-_���*�:=��*�ą/1v��A�	J�X"��{�Jb�}^��c-�$UXv(�'��F�n� �vQ��:���E�,���qA������<U�+RQX�@�x*;b��~�g%���r8��;o��K*"���ŉC�zoh�٥�j/�,1f��A����;���X�q����S2r��zw�l������!v��D��I�'���G�5>���(���,��q�%M���m��u��m'~E���Vz�*��ÛJlZdZ���	zf��J05�](�l�?�~�u���v��ZF�{�������b�u?�k��b<�e����`�0UXg�)�HWB�9� �6��[%o0��&\��p"��=�2��x���P�����$Ya��?	̲�Uu�P*Q9Q�ڏxR�p��׀�0�i�K�R���:��=��N���������iAר�����)yb���ޠ����(��w�j
"}�Z��US��U,����ViD踥���0�g�DZ�`�sz<�~r��$j}�ؖC�����M�)����?�Q+� �����
�V��}�أ	`'�����MQ:x��f7�2b��p:aUܪ��z�\���\<��`��\����lhoS�^����F7{���b��0��}���>B�����:�"8�	k�����Z8���f@�MlRH@�#� �	$��!F5{�83]}D����qȀp�� �}��8P�����&q-ex�.��]��!�W���c� ��/���q�S�KAXL�t��ʎ�,����][6��a�6&K���T�C��I�e�1ό}��<$�/�K��~�l���e����b������V���`�(d;������0<��웖�Oۭ������]�.��2kЉx\�
㺉Z������ L�n7�?r�ƸOF�j���H��~���mN��ړɚiA���$I�T�+�/��o����(�{�+J]���ǥ����`��uA�����[��ht���������/�;�\�*F�Ӈ��n�=���ĳ�]���R�F�[�?�0Q5���C���q�S�b�>f3���:0~��;��C�y��*
Y�Q��;t1��&�-e�abA���;���#�o���k��Й�*���ĵ�ݱ���e}�Ͽˠ�M5���FL|�k�wy\S�B��qI���8)x�k@�Ye=|�]�M�B��=�ec�\u6��H4��_K@x|�%��� �*�'���
&t�m��d�N�?E�Ap(>ЈR�ް���]�Q� $�bԈL�^;z�/�[�f�~�\E��`��!*e#���-���d�<ĥi1��Βr��T���r�,+Y�gSH��Xe,����V^�3���S���gj��@�n���ZUQ�c��FdyZ�8UCi|���p��eݞի��^|
��=}�c'$����5e��g�Ln�6KzG!��e��r��V�9��e(�6o�|-��{H���xT��>���?��ӣ��u*�b�J����|��Vπ'(����L�p�o9k��%p4��X��^*n�g��7��^��]=*T�m��������:"�>��$jUO�u�H-k4՞;|����J<��8�}�����]��Y�n�Qo �
��UY�S����,� �O���-eO��٤ƨ/���rl�95(P󲠕�C�c��'EھI���H2m����a��%���e�|>(75C-"��Tp��|�麬��o*���s/�C^�J̉�:	T`D{7����(λۙ��5�=\�U�"��$�����a���L�L)Z�;�G(����c��0�f�*�N#�7�T A{C;����ʎ���7�}�mnl`ӯ�o4�YLT������碫b�T�<��	�3?N�l�:S�m1���ડ'�p3z�^��"��/+��.! 3�q��!���U����0�o���g���xZ&�-�'7��/l��Ά�� Ϣ��5��f�҂�V�l�?�(�U�䙨�J�۔P�u*멃w!A[p����<�yj��i
6�����B��US�9��n��g�Ѣ+�tr�gh��2��kh�-��V��7e�������� M�䭸�=��Q3IY	�����$�"`���yZ�85"��TrS�;��j-�T3�X�	���.-�3��r�����(��O�TMo��8��c��<̱~'B~�f 5#�~�eD�jj�.R��7-g����"�5���������)ޘ	�W����Eeιu���p�#��IcǑ����i�y�Q��A۳����3���������B�E�n��碻���CT�t�V&.FT;��~���:��`��9Ap`�fk�+FH���?��@�34n��-:�j��dR9{b#��[�~��*壵'qXD���jօ`H.(�@ҥv?��ɂ����t����b-b2�&��~+���YI�8�!HK�(�P���u�HiXΐ�g���6����g|���T�؛�~�f�s����o�6��v.Y\;d�� �itž(C�j5���~�s9���y���@�-`
�o!�g��p}u��,k*��j���SoRfv�əU�]^}�(\[-�Q!�9�?���e����#��e7�!BѨ� R�J�P��m���C�%�-bz���\�e�2S�w�1M���ņ<E�Q��s�th�����G��*���F0��h�+�W��e���}Ip�>��b����X����z�'�qs}� 	���k����j\O�C�
/�����^r��|Ա�5�r���G73�� ��j^�q��h�$pL�5'4��>Ş�s��M�2�S��w���Ƭ�w�gߤ#���M9�U}f�u���2�h+*�ԣ��ך�Wӫ�8h�Qj`^Fl�_�BW�WK�|�1�m�%�%�H: ��K��cՑ'��<7��]MUv���5{~̴�����k�6��a������+?�u����.�K6����X�tح!������}B�����*?���<}Xx)�)��� �9�l�Ub7.������A꼂V��yf�l�g�(����2�E[V�>��2�[�&��J�`�C���(��{q��1{��I*\��lؘ�^|�aA�&��VX6��y.��K�À�����!f���[��:2�#��R��J�0�#H��Z��L�;�Y�(.��n���9ɹÛ�Vm�`�#��x�9��)x!C>��H�ٗG��n������[�
6Ṕ[�""
�϶�ŷ�u�y��t��@�,�o�[U�Uɸ������k��B%�QB���3 ��6��Mfi�f��� �	
�6^rbrb1�k�f�m�
�c�@�v��L�OM|���ڃ�<�z<�U�91X�#�����$(@�rtV�Sl5�$���-��	�6P�/��n�+���~<�?�`�/��`#ƾۖO�w)C�Tx ��N�zgc�� p�^E��1ǫQrW}�a�s�
S��D�p%���܀񦀘��<��m?[o�L0�=����垗��#2��*)�������+��0zs�U�v6h��G��p�h��eT�(-�����[�b���d�_N-#�d$ǫb��wZ~�� mG&2�F�W:�X�����RNOC��h�o��W�x�͙iK2���/fW=��A����wjZ���/q�E�!����|�Ù��X4To{j�f!u���s:dO.7չ�@��]�a�J�ċ�C�YЁS��C$�{F�;W�B��(����!��G�ξ���LŬ�@��B��~&ܗ�Y�<��ؕs�\!�
�	=)O��O�`e����Ĕ��J�'9|KH9V�C��̰c<v��!I��,.�Q�'"�g�I�D�y���aߝ�:����4��$���xQ�'�n�B�G�e5~��B4�Ns�:�1y���ة�x-$��ypb��"�?��*m%�3��H��s�op�Y�
�ۉ��āU��!����$�2����j���0�D䫼�H�D�`��tT"���ǖT�=��-����6��؏;J��q0_s�HTR�yRy1���m �3"�Bf�&�ɅV댩�����u�u�>�V�
q/�ޙā�3���v�y�%^á�s
~`��%�rК�����5¶�cš��`N�7��m����+��D��3�f`4����M��&���e�d� Q��PB��0.�3���q���*[�,ԇ&�$�Ӧ�Vu���"
�ΪV�ۗ
[Z�mdf�z�P�?m$��λK����JKT�����]�Xog����|h�.�����A]q��� ���tww��z�El%��Բ�C�e�?1a(��*�^<�]�w�E��.�1q$�}ǂ��D׍����(zq^io�b5��,��m� �@%�6��]j`#���.6�!�֦�ja!7�|��67'�#���g!�����BWRU85Gd/.w�%*w���<y�)e���E��E��kb���:��N<�U����ޘkl�i;����t����>`C��3��PH=�9���N1մ�F���{o��bw-���7����Z{�О.��.���O�Vt.muI�v�����5П"	�:U�)�f�p(7:��sd�	�IZ�I� |�<��D�$k��;ύ��f֔	�_x���6A7�"�\�k��
,�a>T����I+/�Ů�ǭ�b��{�9����UϢ�e|�p��YSVL/�I(u����D�F��=�=
��"����
�ۯ�U[�@R2eo�b�<�ċ_����[�1�t^�/x.=[v�� \r j��/�kE\	z�1�$����đ��r���*�x��f��Bi��'�ZJ�Z�D��[�<�T�d���Ww�v��9���L���u��-��bE�4ԾBL��Db�����4���}�N�"?�x�E��ԙ�o���E��T����׵%F���G	�c�����b���R�2�o��(�^�,M���ڼ\�`�;�8P�Q� ����[JH����W���`ϓ������� ���zk��!-T��9]*f�R�o���r�ܙ���A��3n�o7!mj�-II~�Ǜ�_3�?�S�{DV/�\�5�:���bǿ�s0Y �$.��/�"�箩���,���0S�h��-a�Y�Q�RTC�3ph�0��
���x��1���3�T���\�{�r�0B���/���l|�t19bu�ͱa�C� 6/U���41

h�d���&S��=�<�w��X*����F���z�IK��]Y���SK��hze�-�i�V�jc�^V鯲l*p��"���q���p�H�^X�8<v��?�G=��u���"�%��U�k�F�6��6z�����t��:=l�~�L��<d��5l�^�����>��m`���y�9VG��V�%k�,y,.u�v ��nw���Rh�Y���h��a�ր.��$r�p9�pYr���'&@�G���/-��u��E^-B�k�-�����ʪ�V������$p�!����.A��Z��H�ۮ�p�3ڕ�2m��,��-���i��GZiT��w�Г����&x����U΁-VN�]ڪ+�؟!�34A���f���RЂcF��s�`xMQ�}O��76pO��1��$'�j���G������!�(��Ǎ�v|�*��:%i(7��3�l��U�R<Y/2�p�Rly ��)H�b����odWR���`,O���f�Bn� �x�0�i����l!+K��/
uIo�]^a�)���K���˳����
��uR�J������~"gc�����������8�y�ϡ�׉�kc|�`��>%=�����%	l�б ���܊E�o�E*��</qp����*ޢ�J�Ɩ��� ��D´X���y��(-�H�Y|�Lx���q��1������&�plG����l�=Y�9�������:���p{Mm�S��_��f��,j Α����V�;"Ȱ����{*ƻ��*��ʰ�\p�
K^�&�[)'�ܿ'��q����'��-�HQ�q`R������nϦ1�w�X�2�+
j��}Gd�(�����
(W�L����
�XQ2��j"�?\Dr��^{-KX�O�T�I��,ޙ�dN�L	�����^�ٚ��\�Ò�ד�0��2+0͏σ}�#����[��v,�I�R������p�������L�K��f"�Z}^�Ko℘�����y�}�'5k���I!9��@ȶ������Y2��ۋ�:����V��+�nW.��J�8 ��zP2���J��:l`d�(�K�����D�|d���\�v�|�����Q��և�l�G�Vβ�G[՝���*�U���˥1��\#Dc�P�f��~��)���5�
�n
re�������WX���	W�ߑBEq �>�Ȁ��/�y;�@``���ʬN���s�jfr2�fh¤oE�c���5*��h�T��`��L8���} C�p��Ȯ���Ѽ^?>�����ʉ�wI�.��p�8+��H�,њP�������q��#���43�0~l��u/�/]�`8�K�ъ��me��������3t�>�n�A9q�S�E����6��Ut����]�ޔ��G:.+��/�i���=�5�F�-���vy�4��D\�{[؍�X��7�r��M�N�N&	KOC nɶ�:�R���ّCw�Ka遅�-�QB�"�<h��\[*v�d��ʫ �4$CD�����7���~��),�Ԣ�- L��n}���y�����
a�!e��z3��C}}�{�w��|�%��&��D��H�\O��~�s)bЗ���
�ʮ,��6s:M��9��{n.�����*���b�3�V�w�q��ϲ�!�N�����,�Μ���L x9�����;�j��B)�~3!��H�~�HY{9�̎7=_g~�)w ��Fv���drx���(E'RxZ�auP+X�� ~�oM\}�����)}�c�t�����Nm:�i��۬ܡ'�3��I^�Vq��BntiF�3+ XFBn2��gRxfm����Pt8���_d+��H�I&v%�
4���;� �-z�U�̃����ls�%`X�X�~C�"����Xr(��uL	�(����K&�~��3D�B�{�".��)ޭ��}I��ے'A*���F�_m�(�-0q��홛MW�V�1`A J�H:�׶&:ޭvƿ�z�:���
��KNJ��xF���dٮ/�s��k��xK���7��h�Q;�݇U����U�'�O��.ήQ���M.�#�?�ԭ@�`=Gg^��^o4Q�n���K=�hp%<�p��#{>.��-l�]�|Y��~o��&��C� ]cLc>���+��@t�t�1ŀ�-�tPs9�D1��>U����d���L��J20G(��IW۾¡>���9���L �S�e����Q+���Qfcᏽ�@"4�3Ҩ�K_#9[A~����bi�]��j�+Ӡ��q'��PR�}���\,9�ע+��141�������pS�{b|�k���n�+���{�0��m�-y|5��_g`�}��yz�.�B�j�,�5�ZQ�	�G[.��R�����*��F>%���6���.��$�����W.�t
QٌI���%��/�B�qT��1��>����G>i��
�|�܆Tk��4ԑ���Ҫ�V��&�E
��uS�b�����B�
��J�⊴�����ਾa�$��c�{����RAAk]�7�F;� 6ר#�� ��������*�?'����Is_�X��{k���=D��T�]# ۆ��j�v2�<���,N-'��Pu_�.�[��Tǋ���S�#�|�RD�5V�W-e�ހ� F:��>a��Gt4���=l��s)��,,LJK��73d�uc�j���?@�R,�N�&�A� F�A�.��@W��@|xQ�ʩG��ŝOo�[b�9����-N(��܁�SQ�P%_g2�\�dl����w�Ee���%�,�o�iN3İ=0�du����=f��7��_L�*�WY�f�������N���.cH�����b�E��h�Z�h�H���l�:�$(�;�e�u����wI������nrO9�=p�a��l��U���٭��(@��ׄK/n��6�W������r*�:��.eT#yya�I�e��n��gѱ���dBWHE|�湪�s�p4䚈qe�{?��'�N�k!N���@�;N�]_l����\�b.�XQ��g�=�#?qg�`\����Ni�����U���G��yl2�)d��5&Pb���J������8C�lՓ���\%"��茴�ű����R�|-�F[����w!�Ie������q�'}֬n�X��և����,�/V~~iO>�O�#_��*/�Ǎv:i��Q1#ƻ!S�KU�x'M���y�v���N���
�W{%��l3��^e�R-��=���D���$V#^�ͥ�� ��w���4�=^�V>�|Q y>TS�_-��=\S ��E!��B��-AS��8a.�  G���S�+;���`5br��XP��&��n$�L�`�<�\Iv[���X7ɂ�����eX���Pi�X�?��	�k�� ���,���^��7U#�����/�gh��y��C���Jvwv`��;eE�Hc��Q�����P_�-�)�u�>����7�� _�5���GX�N��)K�����/'s�P �6����VX�������M�������-=sr�/��/UT鼴�� �
8}�[	�3����k<]��3�B3���UJօΗ5I*$�d���[Ĺ���Z�k���Z=i�?OIv{��j֠g)��)K�i�#��6�hh�i`�O�_��o�y��j����Ff<�kb�)S��T����z�!�>��_�CP[�(~�Vʻx��w@$&C��&w���M��s�&�=ia��<����*Pl≌��n0����o�d8�IuO�M�{Cߡ����;nQ�
9�N��0��v���&��L��?њD#��Ïi�@�lp��I�R���O��Jy�$>b�A(�/b�vmX�{{0 v��9�y��j8���,���p�w�)�-u����Wa�7��/������	sj��2�Ƣ�>��ؖ��s�u�ߕ�=���.�8[�ֿ��}����n3h�:�[_OV�=����/���'Z
�A�n�����ns�WrG������;-9���n�Y�e�>�t��r9�P��)�}�6Cxv5g�E�6c��r�!���y�e�m=��,薓KzH�j���r������&�p_����ծ����SM�)�ޜ�Y��Iߋ���@8WG͉��K~p���Y'(��jcݑ�w9�{!*lG�'OM��z�DW6Faw���t�7�*V0�E��;�s�d(�-IG���>��[J7ǚ4-��n��D���[��G��Э�ME���4�����Z˃�(
=�Z6Q,L��K���#z��</��1���/G�,]`9(��5 �lv3&��C�Y��r�H���n��&����Bx��N�B�ج:�9)zD4���ۊ<�x�\3E}��LTX!�cqV0o�$��1Q7�%�`��G#�7	�e'��<��3�p�m�����A�|��mC24ļF��[9�W��]D�5r{�͘0.�]��cYl/
�Iŭ7T�G.,?՚sRp�>�I_��YN�Xd�yO�_N��^r)e�H���p�((?v�ssa;빏>���c�rw�*��E���c�$�h`����	�1w/ D��ގ=�S��h8ʔ���ez')"��)�y�>���n �c�ҁF��y�х؈Bh��?+�`���G�:X��T�	��:а��V�v��ݓv�)a�qEh ;ԛ!'��+�bܳwF��r\�0��JP��d�zb�|	� �qO�����6Z7�)Fk�����}�6��+���:�����ӊ��2�w*��B"��1�p�� f�i�$o�IƐ�n8:�f=�RLbm��lB�祦4��J�����R��=��"�#�K9���k6ܵ�
�EE[�B�n!$1^�e2�~�M������Ve!��G���<�z��(s��%�u�:�g�(�9�1Z�o������e.�v ��
sR�}4��1�Ms��hƿ���=��^"�.]d���V�������zI���.|��������o@��lJ�j��޻���=���Y�x6%f�~L�0�р����Aq�M
��x����a�E��X�
(�85��%�TE�L�z�'y-mZ_ ��vK����Ag�����f��;�B�(M�����ƻ�Ȉv�5X��T�'Q�|A}���n��	��RT��� ��ٓ���]�u7��Z-o�g��W�#,��=Zf�)�����f��k���c�N�rf'��'�������"d��F;9e:��z�`��P�E"����}3��-�ƥ�Emz�5�`�[&�S%ʪ�:T~щ�B�Q�����ӹ�.�^d�G�qG�~��e,[bAg
�Wkg'�E%'])7��c�^�z!��<;,�d5XD�k��]��^�8a+�*P�ê�@��x���;LAQ<��<O�{"� ���ʒNJ� ���$�R{�mFA{��(��ΧUdJ
�Oy̳���+���b=�����(�N������w���Ѕ�JH�7������u�gq���f�fJ|9C��Cf
GU����E��vJvm����'��e��*z����,6���A�bQ�	kiض��F�.�H���A�"��dq��"KC������=[���z�"Mgÿ�����[d����o`� �ߴ���pVH��W{���$�u%z'�x�~��6�.�X��i�����u��N�ƙ��)c���3j�O��=��-�\�k�l���yƏ�z���Z`Wa�J3�;�~>�<�����Fl0��yj8�9�k��h~*	�֧��LX�!��I��x]���j�տ�đ{0�ݜ�~��/,D��R.�uhr���aN����^};qc8�m�1�oj/����lu-�E,p�ͳ��ej�3p��ȡ��!Ή��؎Pl�!^E�j�)���A��\[7��?6ld8�3dF�aB��vC�r�E��� nG_Cw�v>1�ה����ǴD�ŭ	m���P<�x��U�|�P��a�јГ܍�����D������C��aX>du����贼'���)�s5��N�V*�!���nQEHD��o+,�M�Ƨu+N$�zڤ�89m���n���Z�})>�����<&��Y��S�̬�i����&�[�[��oJL�䯏9pDA��@�꿵�An.;�R���B�U�KyG�����-�#n$��§n�:��q:Y���9��^�� ���A�RD�bE|�{X֎����*aٱK�a
K��]nWch�J�,���)��G}��	���	�o0t>m	k�q�S�(XQ�j��*�:U+l��6>?��.�f�? �'��-e�w/p����X��0�7�S8)/t�b�j�>�\�f�q�}N����#td��4�]p�}M>2��k�Ό-x��
zJ�qY5����,��T
1�L�M��~��`�0&ڠQ��%�O�{�������o�����ø��K4x�����2��=�8ƢU �1����vLi��m ������4��ß��Z�l�?]5�5��z�� �q僸���a7J�������wI�+���&%/I�1�i��%k�XgǪCM?�i�nm�
4Z&�����/4�x���T��Aw:���kC�;G�c
Ѷ���[r�mS�nqlNH�����<��1y�soɌ2oh�o�
a�z��XA��ao�Y���}�<�<�\�b��af�%�R �b{WT\�=���F��0�ڮ�⬯�̻�&5 �u��H�:X������;r��&O⭇�K��X��~��:�$��p�Nե�2,v\[nԼ1�Ȼ$*���؞��Y1"�uŖ2B>h��;8�	-��]�K?|g�i4�ι|�h��r�B�Zc+��(-!�'N�/�'�6����/��������[	^[d�Q�`�46���yPWB��A���]�⊑ù���y���|��W�A�Bb��ƿ�L�R� T4ZzW/��т�z��w#�<�a������{+����>�u�����u-H��r�Hmܧ#��)Y=v�C�r"u�j�U�w՚�����Z�Z�gqhd��1�r	���y��CiǊ���K�Y���0��5�@�	$��v��?*�T8w����c��3��;������[sc>6�b��qKt�9ָ��*�9-��$��h���G�d'�(�c��k�`\�~�Y>}��>�T�0�95����_#AԇG^�֐�I8�U�������Z?���T�ͭ���q���˻uL]�,p�	�؞�k@#ˆ��U�rD4����Ox���ro$�&.�Å��p>Y.��7�?���o�hW�z�}�<���Hg��8B���n���l�R�b�?���QI+�|�Ňi�B�c_GB�p�4^r(0��1T��!8�2���ǪQA� �s�jI��x���.�h�h�� Bt��P5��L��7Z�@.�+o����|�r��;�|��r�����C���mA�_�4��W� ���a��Q:�rp���$J��Q-�����ӰZg#B�Ҙ����;���y�6
Ϧ�����E��J(d�?Ly@�j%�I�7?���T�0��i���:!�!	HG���"a�BNo~��d�1&�0��--8ZY��K-�{�߃�2�~w���%E�S�}�7(����,o��NZ�;V���6���P._녎�7�	~nӇ�P*͓��(o����z�����Y-U�Z���FC�X�㈉)k"P��R��Ǟv���A�l6�J��-�o�j�	ٹ����Ã�����i�y��B'��t:��Kr˿ӊ���/clI{���U���'i<���ye�W�3TXu������#p��wMpwp�Ua���=�Sѧу.馯��R����G3}k�����V�� ���邡tg4j�^���h��??V�"6�8h������(�̪do��v�жR�xbO0 H0D�,5�����2�O)j��{�f���qc
E=�=�ly��X4i�ܣ=�������¨����S��P1w�xq3УЉ�bk5_��r-�-��G�B%`>I��^�0E�CK'xo��m�p�^��Q��&�s.J�eF�Z����>��b0�<P��k��c&mG�d0W?�@�V$�P�K[_��`A�N�A�͒�"y)���ڗ���jѻ>���|��\���m��]�D����,��D�m�p�Y��$�%@��cI� ï�!������-��UV�M�|.����j>��Z�sM;iuF�}�zV�Y������(J�PTʮ}A���%Jc����n�J�ᘲ� ���X����
�%#oۍ'T���0�Z�i2���Ҥ�����
P��\�q������=�|��1��m"%��@l�+��6M�X~����z[��t^W��co�=����^Z9<�6ev(��_t,!d��F������c��Ob��vR�Z���p�g����#��5��"+Lb53�끗/Sq������9�&z�'�_�&���h��i�(�e�U�HϟP����c�Sb��k*����ɫ5��W>��ܰb��Q�0���ZAAcB��f��C�6��I�UX9�I�r�Eb1�P��;�����l[�a"F��3X��O��񦗥��d*q�A��w�(҉^񶂤6e�
�2�t���~��9�K���a��+���J��,w��+ˮ�X�M�z;��	���0�������R#5(�(&�"c�z�M�ߊ%��x28�.��$(Y�*S�i׮��Kˠ�:��K�*��Ͼ|�@n�/�������Y0d2�R���V(�$�'uV��*aT��HWY�R�rA8ڷI8x�g
�/�cG�>s�+5g������͂U��ݔN��y�g��CL2XR��(���ҊV�℈�9'�n}��ه��FO��NB�3F�wEl��`-T߻�����^\�
-˯W��6�ӕ�% 	��7��h��2a�Վ�mȰU��A��j���',�v$PnDD?�2!i4m�{���w�	$�]4�1_I�k��ݺD�<��&R��h6�:i�C�i�tZ:��n���05C��Na�_��0!�t�@�(z�.�)+�}�hg��� Ecdajk��B�>2^ ɋ&PFX	�{1<�D|ˈ�B��#�8q�%�dX�b?O��yG��(��N?x��m!�@�*��6�����0	���SG�����p�f�6����ק�?�/�ݙ0�șL�����s��tI��X���W��5����CW�^a+BoWfu�ԣF>�r����g��$�@F��K�	#��]��+��Z���b��"�R���t�4�B�834qS�~iKA����*9���"k��`���)3?�6Q~�@O�*_)�x�J��_I��2�a����7��ʶ¦���A��.BF�����d�(D�H�v���s4@\$Y�݋���A\mr����#����t��X(��J$=���M��U�|?�gHx�Z��z銔�|t�;U�λ�(�go�<�^Åk����ok��)�{�o�1CA��D?ȍ�Zzx#�R�N�P�gL��,�
�\��N]��g��(�G�X����zg�RmX-p���-nc�v�m�X'����OA{�y��&D�_�v�}��#�_�����,8N�
Ć'3R���0&�8'wn N��&�˦��2��#��<�s���Z8�SX)Z�n���jYԂ���y�ؿ�̢�й|�ux���Q���r�䋳����A>�}�5���g��؇1I@��܌bq�4�����\��;!��v�~iP+��Aݓ�?���ߤ=�L5G�4��T߃Tv��d�Ջ�㌸�Z���t�a�o�i�'.�KU)�BAT�9k5������N��<��TҊ1��@݇�m���8��̌�\ԽT�k���pL:� FSP�L*Բ�0��ȉ{�Wg/m�C+z��i��!M1W^}�[x�߻�ɯ�t�E����j�L\�1��KA�I(���i-�a��Ev�@���e���(<"�Jp!>yŢ/<:	���H6�����E�bݑ�آ�f�����E�E���ݚPWr`U���BA�,Fj�$���+�,��xtދO���*��22�)��a�z���!K���_U*�&}Z�d�����o��s`�ۯiY�2�ߏ����n�_%&Y��r���`���PsGmi.�F�;o����+�$_
ZtS�)>��h����xMi�����\�y�?���v(%��B��+@FM̴��1�5m���Av}aDZlu#j�C�C�y�)T����_�!zV\�'��LN��3�>cb��g��1�����ܕ��������yt̫&#Ş�!z
K�ڦ�:e��b�����w!C�	{���;O4��\�<�gVe�<Jݐ�EMaU���3���(ﲛ�B���fn1\rjb�N�w�W�����~�C_5�YT08!v���$n��*�-Q��2v��K���d�����*FoU줚SW=�; ����I�bK!���о��3Cz�Տ�:���ba4
�,�m��ycQ�7eF^�!�8�P���K��1�&�I��i�L��&X�D���_mck
À���	�M7���"*�f�8���]�4�a'p����"��۝u�<>�{9��#�xS�g���[�a���lW�*-��1X�z!�ل��d�����ߍ���Sм������&�hgq:���G�x"�C���W�A��$։xc����u�I&��hQ�qJ^$*��o�t����(Ft��AHk������cFI뾴����{^�UQ���*��u�f�4($�{X�P!Ët>���+�"ⵧ"o��(R.���5�!�����r� $�+��M�t��¹�`FOYLV�������w	��-���@�wa:v�|g��_���h��^Ӑ�떌54�<Ҡ�7��1��zƈ��.naLj��^���J8.!	�%V�N֨����ʸ{��@h��l����2:�#�W6�Q�R�Wq���0�> A�t��1�%�eي��,���`��]'	w2�m�F�M��J�"D�s�0^V~�-�X)9T���wT��:"Δ�]&��@�<���y��G_��VF@	��Tċ��%�.��I��G����8k��e+�-7��F��;�3*���.��(!�\ ��!w9�aƚ�%�L�U����`J�	���\�/\%�B�T�����xFN���x�!,Ӡ���9<��:��d%�%��iu-����+"Km�9XVe`P�l[�^鵐�9g��� Y�:�[5�$���gŸ��������Z���~�YP0���Np�b-?P�K$��l��,���F2:t����E��>��D��u�w²g;	q�b2N*N!�YC�V������P�ĥ�z���?��N����y(��+�q�j��B�OX<�܉���q���$���MR�?�
(��@���NSp��0���]�<o���$���Ҥ���f��|ܯ��L�s�x���Uq��ؤ���jpU���q�F3���z���힜�#-�>/� �Y��8eت�=��:eQ';��"yPB.mZ����璬�Řvq�����2���Ǭ�&�y��W�})O�/&<5S{�r��{���c�i��>fn���{�E����N>ř����KQK��ޮ�H�]wC"!��EgA����xuqf�B_E�����գ�7�9���_F@����t�Hy�.��MUN0o�5��\@�i�ߊ�
�~�1��������J��봳����:������e�]T6�ƣ�,������A�T��B����<O�Ei���u�%E�jw!~0�z��B�3�"�LXM�üjk��-^�m�l�sTG2}��0���-��wl��-�?� �&����/~�ͱ$�y���&�d���a]�V]����l�F-�~N�#�Z���`d/�,�?��%�g>�ɞ��JM12��^�0u|��š�̺�-~�$hjJs)�SD��S,��o]�i�l��9��6p��Hߥ���a*�5�j(xt&��e�,4pf�q��<r_��!]®X���vr�"�F�� b��������,'�9�*+}.OKg9�1G
������В��1�a�[��DC��5WE�L�N
�a�%��'��ž�s��z$�BV_�Q�㖅���_���f��b���y�oZ�Y뺒cV�1�zrO�,�W�mip: 0m�����C�H�T$+�ӝ���v�����6�@�JxÚUͿ���~ל^0R�N�T�N&7:��s�-hN�˼Q�k��g���µ\�x��P����^�?���w���Rq
�oӹ�G�ɤ���T���w��Ji�ͯ����_�Aȗ'�қI�ǹ��EV��Ǜ$"����5���^��ib믮Un�: �P�)�l����_a���������2��vs9���qԵÁn�Wcҁʷ�F=�_ R�.'�MK3����L��i���)�	90���v���3�7`�ޜ0g.�+z�Z�'�iǏ��������r�/�
'NA�]{��!��6OQ+T���,%�Lg����QԿ]�K��f�ou�ф�E�1 �� dr��舩��2Ղ�2��w/���n��K[��1H���m����4꒚� ݙ����m������_���4���p��F>z�FI�FU��̬#�FF�������mgv=I?�@����x@#C����&酱/=Fg׷'���K��>2|��'��ś�Fެ�	�1�bA�n�@�����1�P$����+���D��'}B'l�5��@����h��ڹ�a=Hd�{�U�JI����1�����u��y��rcf��B ����[�q,���f.n # 9�X��;vdv��c�L�{,�u���$��>���+@�s�raK&}to�
Y�Q�`�Cd�QW��"�ܿ��VI{Ar�y�?�G"Y��0�H5+��=+*ϣб sw>R��[L5p) ��IX
�U籿�.�Kc��c�{�>W]�LAg��O!��!΃�95x�P�$�q�����e��N�8�T�!�Z9�$g�v�CY�Q�L���z�T��yhc18����|Aa��f��*w��]��5��+d�mVZ�o+��L����6��"΃Q"�ʢ������E�?��e%b8�"+X�7�y�<��jJ��QA��9p�$��rq4u�!�l��i]��� ���8&܈�򃗿�u�*i�Q��x�+�1��g��m6��Lq۹'�[''LЕ��O����=������ʕc֚���%�����Ɉ�G9^�|���Heܚu�7
����������/$ }���Ѿ��8�>�p��+%�Z��^�;�aP)u�?����'$��[3u.��+{�y1L���;�<j����kX[,��̥dD���5��S�b3�� -b���c#�B�S��>(ήCOi�ד��#4�}�'N�U|p��e��ًʿ�e5��o&&ix���p���(;�䆣�[(����.�
i!C*�%�W���Q��N��]�n��+�c_ӓn�����"v,_)@u(�e��Y�,/xx�`c4�n�\�#mZP3��:��ώ�xG� H��(�9�=��}X��ʎ������.�a��+��v5�Ӂ�<�9l����P~�9�v��1hӻ�B��T�7�
4�2��w����n �u��4ed7�6���}�G�LFa�"|��{��ᴅ�[�z:a�J�:�E�ܹY�,�"lԘ S	|�0��Ƒ~�9;n�qR-T9P�i8�Z�Q{۷1��T�s��b�6��+	3�l���w����pì Qnh'Ҧ�Rt�̚���)�ݭpy�Ĺ̋��!�F����$��"5��8T#�K�[��cᎣ͢�X'�zi���^�r�V���`��Ri�9
uC�%P{�
GJ���j6�����?(!|�)��i���J9[Dr"N����dW�Xא=H˅�v��j�G������9�v��L���\b���Q���B��&c���d0�nȁ���GElT@�mU �e�g���=��ζ�u���mT��l�}�̶w�ne����r�a��i��]`��̛��ɪZ͂��L�>T�����k���$zմ��
黳��`�p/�����CsA��~�q���2�wO�������V�˨7a2a~�l��c�	!�K�u���o�q�<F��U�{� ���'������r��P�>�Q�!�(������;8l�	����KPJ"�aDg�<Ҿ2z�V��l���m����nbLn������o娀�{�� M%#/�>�X0l�:�a��i�m�*z��r�p}m�; ����KJ�Ĥ:Qm� ���V*�%Xq�Q ��b��ƅs��$-�$kJ�3L�g��C��+l�pjU�T_F]~0���q�;�x�����^������6�MesW�y��2��k����1���Z";����@w躾�R��e���㔿���d�*���u�5,���-v�6�1Ig-"󄎘�Y�'�J/�9��Ƴ�	`�j��u��(;��1�Ns�a����n���|������`�j��y��ȏǌ��+�%��a��Y���+[���v�y�u����	ۺ�nZ�F�cP�lZD�R�Cb<5�&�����0������s���{����C.�a�$��7Y��O��!j�/�Ľ��n�׏\ݒ(Q=��?!���l[�w)�-�>�c�9�-A�d�E��6�Х��O����=�`\�<�a��xD_��ю�}�9���o��*�A�1u/vd�D}�ҡ�O7C)�pyH��[L�**R=��jɑ/iJMFf�Q݋O⪴��.!W��nЍ�eaAg�{�B����p��q:q͔��'���c�ҿ��;xw=N`�K}���0�͢8NnS>��=�������,r�{�F@���'؎� �������9\!]���7�I1bvR.���L�ڣ_!i
�9�����g�?�Z�kM�q���y��#Ed��Ѱ 
H}"l��QfU��޾�Oߛ+�z�6�s|.�ƦÂ)��+���T#\�����c@��ó$��`��Cg�ѯ	��)�e��c袲o4��$��wٵ���3H�!�|Xc^��x �ߎ���[�b"->�]�Q摭�mG�z�7oɶt�~��ɣ�/��}?�C���$�iO�mIo`������3 >N�m��~�pRQXi��r?Z��"Q���zM*�f��Wz��R3���	���"�>��.�+�T��	fQ�Z��Eȝ�hI���޼���C�z]*;�rf}	�0lVV{	���Ԉ�Nn�4��~�d�����ٹ���f�t���J��+׬�~���p��J��s���Y�Lm��(�m��}�EM�װ+:����gʇ�
g�����Y\���@dP�Z�*('A��!jH���@�pL��R8}��cح,=N�"�Iv�Y7���V.\x�s㯐T���o��EZ!���)	�m:KL�9]��OkE�|�Ɨ�=v��H�Gò�4�q�V�(��q�Sr7:�`�S6���lC 3�2Wi|%k��f;�'+�ry4�4��6']g\g�3�a�tµ��|����lt���<��-�Fi�r�e?�����e��u�T��(�Tn�!	�jϨ!H���	�Ȋ�X�X�^ �����Ԏt1�{ �1k~9����y��� 2�	���	�G�=��>�s��'�S����ZI7W��J����8�f��ɖ�؞9��fv�e�ďL��P���D�tU
-�%p�	U��P=`��ADc�4� m8P���P�,<�.,���O���r4=Cz(h��Cй�3d2�
UI��J�*A�i/q���W�����F7����l�h�|�5�� ��6�L�ć�\%���S�ʃ"� ����N$*"2�u
�
>��y�,J�)b�ј���W�	R|�E0Cb$�����8]ˍ�9��Q�ɫk����v6���'Ə�?ۓ�'�n�j��>�I�;��3���6��LT1��x��k��9�㢅Q��$22�G�^,����{晍
�(���p��6t?׃�qț�����3��C�@EO�d��{%�r����D-�k��7��<�e���Gw���ۙ3�"��z����܁u�����-մ��mv��8?�=�EP0Ӑ�<��A��P �z�5uQ�U˿�9W�a\���kdz�B���n�X�?��yr�ͱ�4�R�`ۊ_�LZ����G�ւS@rv���ڕ���E�4ܰav���?4rn�{�߮�-+�>��^d�Rnڙ����GW�/�a���J�Z?�|M�ׅ�Ƽг�7��UX��EJ���1·5߇�@  &��n�yl';���L'з<v��kewzp�vx�p�8�[iDG�博��b���:t�|j�l
��+�H��?��h�׮�ߙ *�?�c������}4B"����g�>�#w� �ʈ;Z̫�G�Z�mL'�ՋW:g�K�m���=�����7�m��~'x���P	�.6��>3kު6q!�a{ޘ<�9��s^r&6=�;Ȗ�jN���n���(FZ��f_+�{�z��>��7n
�ƚ����o=s҃ma��L�^��V�~�0�l��?xj�����&�DYp)��{�:�8W �X��������Z��i�C;ӄF�Wک� B�.;3�*����.�\�oذ8�ޯ�����_���Va�)ͳZ�*'��BHR�9U���$����&�d�����O�zȇמ��b7���F�V�N��oG���=T����B~�1��t��_|���u���Kē�.�V�vMA��w��E��B9.0yvΙ��/�?���?��b
y��,/]�iXT��x�b
�'j9�cOl��vE�1"I��ݍ��I�u���X�Iv|�.6:q�E�r�Ep���箮x�q#��A�aM����Ex����S�o�ζf�S V>��~X��ᛸ�s��i;�@}D�k��|2$|
s�K�8�Iv�.|�O5E$�\�[
���e7���Ѓ�g����.��m��.���,���.�E�,˸��1H2�g";%>i�MP�Vҙ��2��Ŭ�6&��E�#^���љ�.�\�Փ;Lno�P�\�r�w��m|��R���oz�u���@�6GnSɱ� ,M1����{s�0��ih��C�̚xo+2�qM�&��w�I�޸�K�(��r�6�o�D�ln���ǥ;>qMY�����H��p���?#M�n�%E![��@��ʢ��h��Jԗ��E�k�^�B�tUɡ��]�?x��ơc��^Tv������r�C�l�d�;�۪���Kj/���{�����(r_�R+��u �0�B���t��������;��$p�����b+1F����� ג�0D `�}���寅W+`�;��,����U�?��L
��G��;0ל���U�n������/�U�5�h���NKf�ǿķ��ZPI2�"W��1�%l��;prmF͆�� �)��n�nd~a��k	-��+H�%L2��h���2��(���w�y�q�e��i�o�ƙ�z�A�mJ��Nͦ*w�^��e� rR_=�?�$���|֤;��9통�c��1-�~/D*��
ؒt��*�̱p=��Xi��9�:NeD�Vܪ�GL�,�JCj��"�Z#Al"���c��4��2��2p�t~�����!���o���(��B�ű9O�@��O����Q/��<�%	�F@������u,L���J�OM�"?�R> 	'h��T-������彳�� ���:�o�ޏ��d�ar��v�����u�	���ĝ�($�F���ek��D�)ѯߤ`r�Q���%G�X�)�t><�ڢ17�h0F⿺[gN-N��7�� �Q��'�������+y���m�ޛ�;LL�_ݭgt2;�]fG��o)��kD�>|�3��{XvW�"�;z0����c�	Ί'����~��e=1�38�v�t�Div�����]*�f-�[x �"e���Ļ���!����M>��i���K�Q�.�鐾&l{�b��N&$l�|�V�Z���;u:*��V��Q�沸}𶞤���ڧ޻oT�dF���P�p�R<k��S�&�[���5ڸ�]'-cjn=r]�b��шu�f�|��f�|`�\��C��9��1Τ������&�&Uآ��6�ln�O�e�@� �g|+���I�+��@��A �ܦ��6�L�����T?��U�d}1��G����\�Q��EW�����s�e�㨞�U�p~s��X$�:q�����7���МA�/q����g]���ц^=�l�I���a�9���F���6�t���ޠt�XB�o����,9�᭙�Ҵ�]�r��#:�Y�J��eËO�=�v��>¾��{(t����F~(�L=L
���
��w|G�����,�Y�β���O��6�ϻn��3/�����K}H�pJ%a2����N0 ����^ ���uXq�G����d����QzE ��p�`P�f���z�G<>)ȳcT#?61�|(�
v5����U�zT�6�o�،^{��s�ؓ������6�~��ݥ��&�Z��'��(�h��d{�&﬊>3%��53H�$�vA����O^%�{O�����7K�`�I9Or�g~J�&��gN���ڷ4K��	),b�;1�M'�����='���Z�ؿ��.���?�<�����&��S(�nc�����#]pe�Iss�o㖶��#��s�:N�N�u�2�>s��Hxo*��T	�%��_N�v�"�h�=���;:`��}5d@�y����td��P��F/��!C.��)���g�
f�e�/P�
'rF V�=dٽo�jF�q�4�sv
�Y��X�a�ׇ]1ti��P���M�Bt�a�nb�zY����L�{
ݿf������#�|I<�F������-p��=QdԞ��I�g�W���=z��k�n�- wLk	��Up�|�S�ً�S���Ag#d��̳܈�Na~	���A�TT�L�q%f����Ӵ��84.���3���!���ݎX��m���b/.B��ҵ@��d���$x�Ar��Ѹv�N��G�s3�Ȫ}��&SG��|�����#n�rl5V���^�$�eꤓb��g ł�#xX���
�a��&gW3kE�ҫ��=s�C�L�](5���O�X�Zy�����$�w��g�v�*ԧ��|��1��.h��������m���D�j���75`E��~�6&xS	-�^��M�G���|�K�Ŏ �"w@N���@��p��[�7�b���5x��X� �]�8�3�C�� �GY=1�R�t!݇���^x>�%�Daa���& )Y���~h�q�^�T+���h�r�4�
c�~�q	�л1l%n��n�F��k�u���G��iAZ�1����zǤ����!��#�{���[爴��ǀ̼�����,5M+�d嶸�]���>�t���ӑ���ix3��2*��Wo^��-���G1�C�0ĩ��IM���� Đ��ꩡ��v��|����TI��*bk��¯ �N^��rX�"?Ӭ�v�$�&��ל�p���-�;m:�ZF��<��V#J�UEI��l���vKa��0
V��-E����0n6�@���PTþ��Y��s$4�<Z2k�;��^2OE�-扖";^�>l��1s��NgDV��ˊp5��s<��e��Ќ�o�c�։��;&���m@4�}YQ�i�����o�t�zoOIϗ��pz��bE�(=�&�h����JK�n~�f��l�Ny�*�2TV�R	(&*�VI�晋��PF�ݫ��zw� }Stpg�]�[���j�k��������?b����'p��ԥȖ��1�$�U\%��P���G]s,;3w��i�ޭ"^�nW!=v^��l��u	y�Ƽ�CW�p��)3}	py[uO��M�L�t��<:af�l��x<s&���18|��!�2�JTє����Ea,�?�N���$�$���� ��� [��208Қ��Fh������Ż�])����
�w�ؾXh�)ǐy�S���uv)��s<T,�h��@�5�F��Ag�x�[c`�U�2%��c��\W��܂�"��O�� H��NF��fޜ�ʰe^;��6��mk>k�������Ӟ�,��=e�B�ǐ�E�׹y*H��ې�9?���n����a,�����V���/�q��t�o��ni[W<§nN_������7��.7����� -�-FǸ�Ɂ��1�ۛ�wB4^�=��9��9;h<����y(.��ڬ-$~N<{Ck��)g�r��Eb�\�UMa�>�l���GwKj��R�'��f�5��R��������y8�=q��� G�_�����قA P�?G؎�8����ܵ��bѽ�U��qj�I�L�	���6�J��e���q:x6%��GA�v��w̴$��Ű֎R���dQt������,Jk�n:D�Ӊ�Xm���_rl�X�V�o+S3"@A��ۼ%4YTc$�&pNܴ��D��K &��n	]�Զ?��Mg{gx�������oOUz�M�8"x_����4���*�42�z����m��߈S���[���p��<���p{qKD��I��)�3�X�s������>�D�5ɯI;�U���Ҥt��;#�x�VuF[es���Yx��b;#�4��� 
hR��/�qL��ؔ!%/��ߍ�^-���{Xo��?]OVl
�[�����82�K1̜�> 6h��בa+Z�bd�f��&����*;�������ߨ�	��懱*MxO�I��ꟹ�ڮW��X;��7����Gg�G'��I�*P��:�!�.����ɫ3� &c�0�e�q�dU-�Q�	��(��,�~����&�ux@{�� "��`n�:FW���q�bb��*3���+�����ϯ�����<d�ن>IL���	=L^�����7A��-b~g4�vq��9ӰҊ
�֥���E�4���??�Rb^�d�l��'oA�� �"�O�A�����Ƀ��Ć�r��dӔ���fJ�� O6caa�]�.�!.0:��*�T��:kƘ��υ�mb�5(r߈�1���%��]M�"��"2��,͐=�t�11Uϊq �N_,����>���l��2�k�Cd�!m�����2�u>� $a�2ؘ�ݗ���L�g�ʣ�AM��u��
�����ͅ�^��(4�N�[�l�r`��O!P6�m��e���z�ץ&�}8m/����G�_�o̻���E�*�e�d����Q�`m�A�kѷX�%���cެ�j�S�Z�2�Z�jʁ��rv7�|�	$���u�#�3����}Ht��XD�6��ǞQ�2���S����D��G�~�њ0�MT0��J�,&�4�zl[������%D���N_��Y_�	ɟ{�TZ��;�g����QS)_!���&��	H�2����]���<��V�&;|����J�M�E�b���ٓs�d�*��O�ܗ�d�=��ߗh�k��VxX0�l�NV&o��lZc���n��/���%2��Ż�0@:�W�6;{߮��D����v!���`�WzY@U�������$g�T����v�TS�bvB��(�I����/��"�+��ؤf�l��B��B!k_T��8;��{*o��$�H=��ݥ��kZF�8P1�C�Lo���9b�����G� �/_�<�
h��ͻ���S�=$����2��Lr�K��:(�	6t��u��u��VY��8�,6E��sVE�W��;&���kʞ6��F�Ǚ�W��u~��e��]�\A�ǸW{��%�~��WSϱ��?n��@���O8��N��f�0�X�:B"õo�yW%z����)�]�{��K!^먹�K�v��n�:F�����{�1�o�r����p^k�A	ʇP��Z��V���!b���\~��BI���G��LM����z��X`�)N�j=Πıe0@w%�GW7>��0�2��aUI±$����F3D���&��e������)O�.Lh�r��T��!����=��T�ȴ���p?S�ހ��a���{����cqף^� 8.��I)K�yҁ�g�d&*���x�̝�/�8�*�x%�����B ��p�EeE25�ƃ�)V���ȶ��t�G���h�-غ�]i"w�hG*�a��.�Z��1_�yw�`�X�
����;����f*I��Hw����Rp|��i����72o�y�u�3��P��a�����PR~w*d,n�.k�m� ��*#6�6�1a<�s�L9e��T�F���+�����"f��B�``��"t6�c5��.b ;>t��?.OȰ�5�9m���>�~b����E�</����ĩ��2Q(I��r�2U��͕���ie0�u�+�*�L�}75G��2�j/�+�GAB�O?*�}�G2������!����Nk�Z�Sn���=Pd��r�>��}����O+��ف��W�t�Ɉ?��[���n0��gl���g����=�M�m��0K�R����T>ك?O+	X����z\1+��\0ns���t�B�T`�=��$�� Xjɱ�G�w���I'��1��"�z�������C��tgX>����~��H���G:�h���+ �1�d���I%���wݎ"uR�ָ,K��?�ꄙN�ZX�����A1��J0y�!���o&�ئ ���X�P�K�(bT�VCK��;C�f���U3p����"-���)P����#X�+���2o�^� ��htW˄u���(H"��&�EQ5���-�[�py���)��c�\e�]�'J O^����5�G����C:ϣ=9c�÷yF�7B^!$��G�;��c�nB��*~��&7@�g4� �!�©IP�V�m\��	]\ע���?���/��O��ل����<�ΰ�4 �m�Sve�Y6,�>��c6�J�8b�O]���D �yl��{DeX��v����øه��*�9	��3���4��l��-�[�'�"�ѭ��hE�Z�_|��Z`*�Zkܚz������T^5֛�񛁏�t�̦���X���F�z�q�'o�n�",|)P���e�c�ފ�a2xT5.�^��y���9:�<oKY	c��g�n��qc9��B7xvo�B�}�v2���һ�ޙ���}܈�����g�$ �@5m��!J4�����@�m.�z;U>�I�*//��}K�u	��kT,���b��l�7d�
'��rt�'�,("�2��l����:�NF�i+��Q?�X�S����l��1�'��v�v��x�t�dx�& b@��c��zz*�K��8���V��ɻ��%��N�K��z�ᄟţ�n��zp�U�+��_��P���öU��csD4�՗����c$���,�����lǣ)J«�Y��]�������[1��Y�Ş�A��YUA��+���R�g�S��%n��?��XU���-vt�g�N�ݖ;�ޡ�yEle�汖L=�"�RIٞ2`i ���U,�8���47���oC�vo���S�nZq#O�� ��O!ls���X���(x"�JE/]�*����Ф�Qe�Ymĺ�Z�:s��ϓ�{�oX��/��/A��N��=�>��s��hOn�~�a�����X$���Db����-�P��_�T��&���#���/lB�0h����S<P1i�>z�q���mo\��H�]aŔ���	����'4���~������(֔}����pp.��l�w����D��nUA���������j���5DL]q�.��U�9��F0͟
�t�f���e!��;/NS��E�.�i3q:.\ʡP����u��I��0�'�;5��\m��1^
%*��
��3Zy�� d����}{%N 3�g���C�y�PZ4��ӫR�j֙^h���VI&�FG|�H�4��6 ��ғ���lx�T�Wi<��pQ�WQ4t!����U$����p����#�$L��@`��L�i�tAh.�_z����(�ݭK���VIg�Mq?H�����R�Qz��+�I[
������_�;ߖe� 7�^r��6�Ct {'���N���f�7XD��c&�JMՀ�k�I��8�5�Q��*U� ��sjD��*|�O�ZJ��7�*�Lr�ĉ��������|%���"��Pl׾t�����1wxKd����'6�M���u�i�4������dUtg#�"�ޫ(���n�]��O(��K�~�<�٠듋��[�KK��
W[<�!�r�f��kDJ[�g�y����^�%�:����R�3� 3�"�C�kdi���)~q��x%j�Emqr��'��5"ݴ\�X#	�W��	"Y�w����i<�y��뚴LI�����m�<h[�jO��S�S��6���G�ߨ)7�����*�G>��x��`ϯ�����~�xv삸e˔J��=�uO��%Yf̙����+�m�Ȟ�2�G�v�
	�S�HA �����6��F��/^c�<���Kc�BhGةw��x����|�7���/�ߡ�F��8A�|�Fܕ��ʀJ	�?N|Q��h��Z�Ă�ל�n��	Q����`�_�w1��TU%n͡~���.���W�q�0�@^�uE��ʹ&�&����~ �s����u���`@ن���=r������Q����P�A3,�f�]�A����1�a2>��F�*�+P��M9?��pY��.8���z굘b,Jy	Ԩ����n���|�A�Bt#j��3�cY�(,�iYz�ݒ��s �/ij:�[�Z�w�D�v��	>���+,����ީf��L��r��2�)(�ªp�7�Q��l��~*�����q|�&^����/��(ZwM��Pi����H~ �}���F^|���z��˟��3L�~㈙=�<���PJBH�[�Q����*�'VN�{^e1��D����aXz��
6�%[O`����Ծ�0"K*A�ہ~��F��rg*�g�S��������U�:@�<��������|Z�Dz�� }�����%/z2��ܢ�'iʷL���ξbC�)LF/6�ʠ;b�;�_�[C��l���t��+� psF��be}�@WBN�1VGS^�=�B�� /����i6��+0G��3��q���@������_/Jzt�V���.`ݢ:���3�N_����Z��s�v������e(H����vҖ�*�W�"<�z���n�TJ��v��%��A��:������kZ���@�H2�j��s+/^ ���浧�
��yF@8��J�t0p@�0%�k��%Ab�+U��(��I�#w j��OV� _nt��Ɩ��γ��t� ,Z��0|���6��FX!t<�^$���"%�>�	�Sv;�J��|d��#�7��Kg��y_�#�_ưs��՗SKI��].H���ôk$���1��3^�~�t�ع�2ݤ숢���@�CT�J{��d�h1Ɇ�}m�î+���<⑩����|]���eJH��7�'wN����O� �2,ɷE5é��ŲYݑS+�=aM�	�b�H�#��J�v�9�WXfpV�F+��f�UO�1Эԛ,�
B�O��4�:x��X;d>��O��yXeO6��.�� �Ŗ%�5!�M�I6�U:��t	�li�!�w%5$�i�W�>����ŒGCl�kN�~��4m������L�=�����Z�Y�R5/��:M
��^5�&g�� Q8�������?c�(�Ly"$c��!��NҠ�y����٤nڴ��ZH �����l[!��OrQ��-�sQ�o�u=��fT~�,K�1��C�x���jgnw��xs.�w�Xe9����(�q�3��x
M~��h�2�e(ܼ�v<��%��1����TD�ʲ�"�׉8�\/�A?yZ���1>.�+�t"ͳ�<?l�%ɸ˭��KvB�
a1*������'4`�������ֱ3��Oz���x&�ޅGKM�ez�TKsm;��h����*�:p	���-߮Tv��	��s<�\���������;	ȴ��_a�.�A�M�S�>?>i=߇��z7�Q8	![�v�0�b�@e���	⯍�[.��fm�r�cK�Z��X���n������ϳ�������f���ٚ���/��w�/#�	x9��f�1��2���x�wU�B�DtiK�E.Z�Ҽ���<eOEQ[��n�n���1�ׂ_nT��j��1r].N���:��hG|���/���)�;��ʗFR%1DǦ�����ǯ��}v�1V��?Y˲���[m:O^�mx�k�oVG��7 +�]V��sߝot2p/�j�j]�kF�\�כ�Dy3�J(�|1�C�ի}+�X1 ]��`�0ѽ�O�c3Hy�E,7�R��^�ҏ�WY��þ{��"Yc�i� ��d	qC|%�>���́�P�����%�B��+�K�n|�DtV���#@@2�vc�j꼜Z6�`M���U3�����D�h-�6r�IA7�Q3�4�\ҙRL�K N����ny�A��~4~ނ_ 5s}�y]b.Ý� �s�m��|:�m�v�zBv/'&+�D�xɾ�6�������O�Wd^c���;q��@]H��9
��Ǭ���G�S�),p���Jd��H�t�F��6hqB�9.�4$_��B5*[�G�k�{��9oWȈU�,*����N�eqa���̗�ʿ�W}�Vl#��3Da�w���$��4o��x9R�&�o}h�8���E�O���l�y��u���@h9{T�|
\T��Oc�:�EQ͡���G�´��]�|^�8�Űy1��y�܎��Zg4�G���fc�r��8��ѯTѐ{���;f4>�e�K�R�j{b���PC�f��5�孥�3�K�[�.U�4�j�{�nx
s�]�{��{�����T�p�arR�7� {�3n�UtQl LV�����(oq�lǪK'*+I�$!D�-��l1��TM�V�Z�����h��o�`��2 TgϞ�cQ�M- RF��]~�~ʨm�#r^��d���������h~b�vT����ފp� Ù֊���Z8��xɼc�Q>��8�c���1�H�@�)��}����J�-w?����2y*�����F����#Ov缊-l�c��a�̹�!����M!|pt�n!�Ke%^fOH�y�9�d�7�#5t�܄t���j*��6Rv����"wbcc�=�	�$p�������|���a�����8�Mg)�nÈM�g���Jf˲1�k�炷�j����6��=�rs4if�-�KF���XYy*�5'���b8HÚ��.eUՉV�E�g��3U]��=��sD��p�r��k6l��0�ڴ�^!	|�'��.�����ug�
('N�c�g^��q�,B�II���7���a�O+��v�P��
�#xfg��C�!T��T�h\C�[�4|2#	��[��d	�A"N!>{����ƈ�e�KV��&�D���(�����9�ֲ#{�X� M[�H�T9"|�~Z	�)n�Q$@�-Kwx���e��K���J�N�/����|GD���axC5ڤ}�
p������Rsz`� ���{�A�8-~{���ߦ�lw7V�a���N�"�g�x[�8�y'o�r�䛤�U�ɾ�ѕ���V���-��4�������*���l��Ï�{Tq%ȓNٶ�X�s����
�slOT�#{9�(�jl|�C����n�5�7���L ׻8�5��i?u�ɻ8�vʐ�d���-1�W+z�a[7cXGs�&�]a���A~��|y���}d9�����@�8��y�E
2�<g�7L�4�ʭY��M��e���4\JF�?�jp'���w�I2:x7�M�{ܖNhhxD��#Tn��x�C���*�QE�yu�1FJ�aqa΃gv��ě1�bk<Ǖ,v/��&�<=A�[�F�!ey�>����k�l�5XN����8�S��i'f�Cln��.��5���
Gf/Cz�����cDE�R�#���6^k`��V������@�mA�31�w�2î&�?���۰�]K���_�s����p��me�ZÅл@NѴ�s��X�n7.�E�ht>�q��_����b��ϑ|m~���'��+��j�Z�34�}kC�j�L��3jVШ`���?��^����o�u�9F�s�w���~P��qс��o`�j9b�נ�ƺ��=[$	��J���+3��=���W,�Q�~QM���p���G���T��Ϸ�U��7HO:�+s&Р#h�����5���F+(?Y�����C3ԋ�����9����$���_�w�;7PrŸ�4ݗ����C�+:FN�����_��Q�-��o�h�`o7,��\m�+ ��A�뵂�$��I�p��Hg'玭_O�X��|����89��;ul&����ȣ2�tK|���8��K,E�}kdɺs�o2��96Au����&�r�jX�0I/�9I{GJ��Hi<��e�zj� %��jУ&쎋�x.^:"��#����G���<PT��b��:��SS�m}��jh��t	�n�}l_F�o�.>g�;[xz5�B���~��W�Ǝ�i1�>�'�d�C�hM���=�)�E*����i� �p�|��ND2�y���~�r/��g1F#٫ajt=�F3z-�`2F��>��<Vz�U�t�۾��
FX�̙s�4�{��z�X�tI�a������`�,�/+Q��9��g8'�)�|�<y�-�Aط^q��Zw ן��v�zԤ3/�ƭ�q���CO�]iIN�#�(?�8d�b���yCK���;�;�y�,�!�h��i�/�9~���f����ʘ7�/��1B�4��3��N��^E�&ٕIn�Tg�k`�r*�R�[a�M���M�%�U@�(cb��s��F31���3������A氶���6��@#
�x4#���)�k��V���q�����1�l���L���s��+�*Ł"�s�JrVb�ò�9���",��G$P��gO:7DZza����R����57�>��	���Ƽ�'*>t�uH�*_Dw���g���|��� ȝ�*��x�ɯ��[�Ӎ�@ISv�n��M$��c#W1Ǌ!��c፶K��u�^ <�̽5Q�Q.`�H?qM�mO��B@��d�tiX����k��p�N���� K:��Z����,�%sox�I�'�Bˠ<H���jP��"P��d��@��8�.�&\1�8�	̀W&uhľ��O~ydڲ/�9���<�p�A�q���v�F���"�΂gk�_���2�EH�M�FjTwxW�q���_�_=Z��ꋧ p&�������4�3����]�0{�u`5S�d��@%P�4���h��,�B��YgT���
Vv�i����%Ki�k� `�{,���x�.����D��m��+�ք�+|�_�a�������������;�?�����h�^�J ud�X��x�_��T�'WЉ� �s*���ז�!�o~_G���=�t������:@�����R�o�D>��u�8s��)y�o"a@�	D�Ǎ�l#j�QcLP�P	+�͚�c�4 f������+���̳��:S�U��"�Ȧ\�Q�EVqt����x��^i�($��UkN��W~d�,W�)|�(��+z��A��^0.��-��*�e@�D1$,�n8�C�[�n�O�d1������A'\H\?ݣw��s}S㙕72��}�jBm�^��͈�{��`��ɪ,T���*��Ȇ��+� 5��>l��^,�!>q� `43�s\��t���	�uj�<<�H��ޖ1�B2*�k�j�&d��/�ñ�u��}/C��D���1w�>߅{�݋m�2�ӂ�����tRTM�$�
;s�S*��է�or���^6KY v�H�e��8�`���Zd|ۥ�$�r<�OG ��3���m�aouLlD��Ai�s����d��Gnm��#��.���q��"��>��XX��6$M
O�Q���l���u?�� �3muT"�Y2��O�MPc?����q�-�����Af�6e=�<#�+��a uɨ�sa�G�����x�&p�v_u:��k�"�E��1d~��
E^M�����/8N%⺠71E^H�h�Q��9�$`}'��_7kx��~�:-d(�$��1s�8O��!���%5����y�S�.�I�K[�J��O�\^�!J!j1����@(�\F>q��-Mz�AJ��PX��8ꂑ������(�n��aH�$�OĝsF�D��}6�.�˱.�j�I�h�-�p��	^"f�*O8`V�S��]��eM�f�qV���v>�(�BXZ�	������y�HO�d H��>��:^���̣L��u��翡U�*y�պUn����t�05�=�!�Cާߔ��G8�[��r\��<*�n�Y+j!k�
{��w*c~�3Rp��e�*{5y݀��=��♦'�í�X��� ��ǓÖ�=�(�^�=���*�^$;Iǁ�����-���i�{�B�`R�����3'+�/��{��@jiB����0B��n���{���[3l���0�I	���Ѹpu�<YX��4�u�Җ��q��"�&�~�o�mE�T����n	�,;�dI��V�J@�[����h�3��0��	f=oD��C
��)[	��)�����ߥ���.�-���{~?��s�E&�Ty6�/E�?,@�.ņ6��
�E;��҇���zS����]^DO�4yN�l|m��
E�W���O����c�g,�"HTXE?�o���Be���ɥʐ�,�����Q���A��wQ�����+�Ԥ�_��M��Z��z��
�rƖ��;���k}��5�s��+ 3�dO���襓Z}7��{�I�J��i�ǻQ�=@�V���!հ#���=gF2�][����D��ߐpS�P��&�ϙU~�����������P?�q���3�n�E�}��^��
��K�ŏS�9Ur>LF+�_v�/��<�n���ET{_����f!�����l9w��7�n'9�~P�gn�����Dp.d��=��N�⒍��1_��1?�W8����ky6��_��;?��<PLO0q|Y�f�r����,�@�à��E�|�Z�a�U�J~��ŏ��1��Oc��A�` f����ghO��5��_O�]�K�"A�b�oX��+z��H0�Qf��k~Ɔ����y9Z#d3?�b�������SL.�� v
|��w�k���`�M}��e��adk�6�7�f3�o�w�u�6���8 ����
���e�9�
�#Ԫ��@kA(g�` ���q�I=TM���sP�/إ�R � �-0��:��F�����8O�Y�]W�_E��Z�)
+ص�[�/�V�[V4 ���S�ʭ��Y�8$��SW����9/�d!�[u3w�S�w�X�
�����D��ٰ��{n��Q	I��0�yz�a������Q\��.dm٠?Z�J.^yA-���5������Rqϧ2�?��Uyk�sd�w1�|���2�D{�Y�I�ay3wVK�u�����I�z�l�]B%h�K�f-�{�ȍ�72���iɸ^.l|�g$S�Z;��h��a�q��.^����Y%^�������z��I19���F^�^ş�!�`0����$����Ұ��$�S�l!�ؓ2�g��,���U�
p#L{�I�=JM�AL�<B���4���5�d�Cb;���T��t��p_��y��R7�����8?������`Ч�ux?F�(g�;4e�/�N��xQ����w�������3S.�{&yh,c�J�_�](a�(rM��=�e��y����λ�Ù`Ѭ��RL�(�ET�&�`�y��~�������@ob"���n�0�m4�_�M}�{�/y�"b�Y���S`�n3�>C
��okyW���M�ܤ�U��OSH���ęܣih���s[�CC0�g���(`���OUk1]���ҧ�1.oJ��j���*�p%�OJ@cu-��P*G)4�ϓPd=�q�Q�d8� �ӫF�=[�o���ӫ0�ALn,ލ�>� 1Ɲ������^T�S^�P���X]>���%WK��r��I�Y{ۙ�M>&V�i�D��X�Elm\-� �֍c�
==�}�!`��?�u�=K�0]T���B����qpPס�V�9Ǧ�0�~��H�S�A/bx�����Z�Z��f�Y_9�N��$���N���.�M�iB	w�萟���Tw<-o��Bq�t�����p"��V����J�x�p��`�'΅^�7rdxKE+A�t�#��j�pA}�G\��PJ4�RHz^	aT��ЮV��|)pβ-.��ך���4�QֺR�̤$��ɔ����*�J�Rz܁�(�=��)��M�<�-W���5k2�"S�T@�b���=�h��D���]!�8bpg�Ue�R!e�T�W0ZA�v�6�ɱ~`m��K��J�qt����W���99��r�1|Ϣ���a�}�<��膪�8gR�>V��u�)�eA�m>p����`j�	E�������)�7�!��&`d O��a��OH��Ok����)F~Q�P�!-\`���&`�	+2+#�S�w�k�r�e��Zh5j��?=i���^AΊ�şW�;:�VlmCD�m!���
~�B>�9#4��51�zV<���:8�9pHr������7/��q�u�&[�P{�SI-�{�K��\	�z������'��r(7&��v8�h���@��DS�q[I���8����Ы�հ�нǴ^�軟�q*P�~Ǌ��,�����)̥��.�IDR(��+�-�VQr�0dH-��*�kZ2��F����z���j���8�;%�l��x�L_�z��MEx�Q!`�48<%$89L�"��#{PǗ�Z:��8l�}P�q�m���آ�-� �[����7Vg��r)�*k�:��x�,�n�۷h���b�]��j%R��Q�c�%�5�\o�C�zwu��� ���?yҷ�pZ�vYw!�w�� ��N-�Ҩ"��rl�CJm�V�hu�P����7?$��A�	YDhF��؇��|WڨO������ Z	f�Q&7;�lb<˲#�1lv�rN�iDX6�j5DdН��������4��TO�)W��LG�C9�����>�����-�d���{�9&�x^�x:g~��
��Ny��>.>��Fa��YSf�Gi �h�ȹ��,�^C`g���BԠ[z--��ۖ�ެ�rn��؈ktҼJ���4�z��!���q!��͢��������`�}'�����#N8�M��,��GN,��y��v�Z���l\�(����pw���1t�M.���H���mވ���(��ǔ�c:�1�[ �E�!�$����ej{C޻a6�����4��Z�O�Ѷ��A1dnˑWo"0W��#�Px���'���(�? �#�U/�-6_Ww�v'p��{s*x*���e�&�vC��q�e�����[wΖ�fz�G�$d�Ls���������"�����6����^�/�bl`��Ká������+�mV��"�{��DJR��m_��SN�r�py`?9d���a^B	=���ӝby�%aP$��w�����xH�q{i�3������̫�
.�s���#)�CΗ��"�������r98�+���{%��,pkf	��}T3]�SK�i��y��;��l �����6f.���>ߨں}pץ#����{MJ��GP��+*�	c	3�� ��u*�"4�|3(!���F�e:���@��[�!�a1��P-��a�e��(և�">;c1�>���aB�U
h��Z���y��4H��j��-��jب-R�!��M�G��]1MT��a}fʏWQz]�j-�*L_� l�c�i���e��a.�b��tR`8�N�`���䈆�Th�7h��#Z�Q0�P��ػb��V~��8��}6%0��������F����&�t�����=!5���g"/��Ez����;���#F�1k\鉡N�S�m�ڝ��굨�X�B[-�ȿ}�;D��������޶���Z�7j��)
l�a/���J�w�3��C������-���ytGADџ^"���RK����-��$�W������7<5��k{�Koi�'[S�{�����p�Q>T��Hxbf�E��*��/X�YD|G{�	�i�BqY펜���#D�8v=���S��ǚ� ���Zƨ
7��X�T�]�҉0P��;!��֘��e�`X�T�oHwDԠ+]�E���/E[��]H]� �0����p����o��ct���
�!8�o�Coħ���֙gU�n�X[�m����+.���I����l���e�t����[���b`�B�ݴɺ�ғ%vq9s�a��A��B�NW��x	\�
���9A�7M5@��omm&]�??B�;��ΉDI��wo֛���x��z��!��:K:�v�K��s�~��rڒ&g���.�`���>8)�g�,��_�ϻ�]�N�#J*a�}��^z`�KNs:>��ʄ6�a3�;��A�6�L^a^��w^w��p"æ 12���J���9�I�;L���JtUo�g#Rn�5w�{ʗx�-J�>�����oM��[ͩ���;�ExL��noK*�)@��]G-�`�"`BF�����a�X4�R��"���
f&R����O(w���+@��0�-�C���@E�kw����?���"1�� �@8�g��=�p�:���2��-N��)�	
���'�yX��˯K�Rd��`��y>g�|�Kk� ��L�PbݑOJy�2[��h��X8�|������K !����θ�f��~��(�yv�JG�6�6]
�*���H�QI����Z���
?sw�G���r$f?��|�^@�/�4�5�~:�(���n���3ۨ�r3��T��{�O�_e=�[�i��G�T��j|�q�'�)�O��(�����$�!�ZO�ݜ�t���D��A��iS��n>5x�g �}^{߻!&ox�,`�r">�ӥ�i�����U|�#ؐ��xmAڎ���s�s�b\'\8�Ig8����"
��R�!#_�
�w�����Dܨ?����)X��a�]^b�)�v�{�'2O/�j'Ss��?VJ��t1��I�6�x!�>l�Ү	q���^/Z�X��F,�h_k�c�1����́"���E%ɣ4��9D	��4A3!�[-��Ǜ�	8S?��5����*Z#��s䰂 ��XC��^A)6���)7�Ҋ-���#+�?�p�����������Q�XS�~%�y�7XK�t�fK���*N��W7����,k�����C��dz*<���MiH�L6���bn��"jտ3#�g}�0��HM
����݉�<F���\����}W0o�4��}����.��o�x���.�;��9��J�i\/$c}�p0�4azZ&(R�[g�Y�݆DP�p	I��e�'������",�#
\Vl��u������_�o5�ku�k~pL�>��rTt��ys��!�fX�]��.v�5�}�D>��D�mR�ZW�d�NJ�안�?�NĒ ��ث r��m��Xؑ�ixY2Z�_s�F���1�R
������),֒���'4�_�Xg����t{<>��������;7��+=��h_�ZkЏ�0�� �����������ު�i9�rq*�<�K��4A�դ�FН/��5�}�� ������*ݴYd��+wF{#��*��
�d��[�N�Q]�r-�d�6���=��&�B�N�p�Vo��R��
s��sʛ�4)3�TDQ���Ԙ��IOk[��j{x���D�ҁ���ip#��dp�<Z�ĪC�T�K����$���þ=��"��O��Vإiu%t��v�'B{��"jX[�M���I'��U�$��Q3�>��ѮT[��'��&-P��{��G�&v�l���?Bq�&v~`R�X�철�$�H2_�-����H&5��J�s,�(�y0��p�Hv��it~���X���v����v
2��Jyh��Of�%��ˬ[a���0�$�f]��kv�ˇ��@Vo���׆�;�aj2bѾ����\� j��?���lC*x��6j�`A�p~$�TW;�����ii��V���R�볺m�ATڡ�̷���:�S�U�X��*J�zC\rV[�ui�-610=��0�o��`dV���^\�`�������=��a��Q��ą�)�q�,�"f���#٦uz
��g/��j���2fz�C���,^�r]JԀ���U��N�����G��	�[JnٱF:F��
\��펇A�de7
28�\5|V;��y��n�o���
��S�}{s��UyI	B�?��Z��KU�����n�C����Ǉ�%#=|a���Uixl�3Kȝq��̀�x�m�L���-A~�
h���߶�o4��^\V�}���L�=:���ۄE�k�FB�����B%�2oNP�[�p���C�����'��^�e{KO�m�!��;�)��6Y~�� ˥╳������w�Jh]�3'5�G��-ew|qYŹp�4���ydi������=��.�PPYy4@��肻j�(�1\�3��\���q���}1�D�;��S��fo6�k�{�����G��������V��a��mT�,X���%��Hɘ\;��1�n��>�\�3W�L!���y���NX�y�!U�0Y�iv
��(��s�,�wt=ցd��{)K��;��O��#Ć�CL(;D96l~�����;��e���<�<�㰈 Mn	B�������",����Vm��_9�	��Qf���cdq�@����qZ�+ �@B����('P��\ xIF>y�<��<z����L��׃�c�B%�j��Y��)<��ó�E��ۂG:4,L�~�G��L�{���P/D��񹩧3b�p�2ZJ��-�+�����
�
&��� x��nUA�Xl��/$V*�]h�6>�CIz4���\E�᩶G���V��n�!;uēG�V�)�P����X�(+0�&W��c�F�����O�Y0ހ�|�:V5тs�9�Xn���_"���K1��#����H�\�II��R���ڂ�z�=%=�C#	�]9n��k�����(�M_�tj�k��4s+8���*�����3��P?^��J�����=��ʇga,}����ռ��Y���iQ�mo���_�XMZs#�h�ҳ�$;�J���;��	����`�Ѭ�;&�4�2�$M���p��;�#ݮh�.
����ҹj�,zD�,�Ź����� �t�����7���yg�Gh��}���)w�y�.Y��Llt��)?��_ޫT ���+��H������5�6�i,K($�p�I_��ߩ
�0��%�']�Ah�o	��|?f=��j���s��'�V�n���*q*���0X0=%�9���إ���{��:����1L������C�����UB�� 
�)'�(�p��d�X9�̄8eV�w����4:�#���Q�=~P$`�~֪P�k���1]3�8���Z�0.��fqZ�g�ys����Vpk��E�� .筓M�̯m�M2��Nɴ�Xk���g�Y�ZK)��5 �,��O�Z�<Q~ߨ�FxNv�0���R��{���+q�b,��T�eZ�4KE�B�r�:1�9	Ȧ������(-(�^�n;�ۗy<i�;�ʑ$M\�Z�G��4�]�B�P3�%L
v���2�4)}��7�ĵ������a��:א�A�7�J$����%K�B���G0j$�ɻ v	�벊�:���z�g���`)ɇ�ܝ�[M������S�̏�m����r�q���l�e�g��^�9"���n[r���j*`ܢ\~�������r����
i\�Tuc�O��9f�aإؗ7��T�����m�w8T�Y�<�n���lT�L,�θ��1|J�m�M]sk�Vq�fD�ft��ί��Ý�r8}{�u�S�`���=>Sk?(�*�>�2?%��s
;��g]�� 5��k�C:�૵I�k�YG �ⷛ��|Mg�fƹ��z��-H��/��W㯊���jnC����Tt�x1�RbS�͆?��>��������J��#~���љcTJ���o�Nʍ�*���1����m�"2���Tw�c`/]6��A��-Op�,R :�jK�i�[���	�Mþ�w!�����r/#�"$��6JM��2������;6��[µv��f�<>b/}պ�sD�g�[�A�X�E��K�R����nم �U`����lեb������Uy���V�V�[��h��W��䅝C�<�"X?nL�3Y��%�X���y�҂�Xq���Vr_e��Е:�9�"v�`�G� ��x^h��#5�e���&�y��`�ge>~̡�r�@Ұ��|LY�t�2�R�)˶���6ĵ�OG�F#��3���J�>^��Q�f����^w2��0V�>'�,_"��\y������� ,�*}�,<��������Gt+����X`���d�0^����G�ԟȹ�h��f�G��n)�-(3f�;ݦ����X�zs�)�x.�#�t�y1��X�\�xD���3�*q�q�ƍi�g�L����u�)�؊iC짤�I�zA���߇��}��ۤ�~s2��Dǰ4,��|D�6h�
��8a4��t���&a����~��S�Oq1�o��o͇�Je�LY q+"�|D^���D�kCє֘1�lʨ�Fm`�H�?Z��)`�]�z�5k���,4�3qs+m�I�sut�h�E�|��^f��{+����N%�V"���l;.�,��Ve \���CF:A�KY�~br��������v��;+��{�6x�;� :]0*zI�����.��v/�RiJ�9�U�!�K'�K�!��խ^��M���+[c�1k&�\��7����(w��z�D�<�E�r	��Q�Tjس1R��6RU�}]FY�"[$47�!��*J���,(�<��@9��Z̯S�?g
ԝ�!�
���Y��`s�i��/���=d�NZF��n�uGP� x�е�17 dw�?�(��i��3��E5���_m���y���@��6bDE������ 0�T��J�7�)�T���(�Dn�7=)��$Y��c�f��'�*f�g�P]�X���N֮�8��屿�Z�ܣ
�~@z�{mI?J=��� �X���-H�rSRw�c����"��p�,r�=�� 缸p��,G�����B�0����\٨u�m#2m&��b���ed�}p�>:���|��W*�'�8L<��5�_�t㝺@�4z3�V���� -Ud����&B���D���v�d���m�l��)Id�0�p���Ӂ�qM ���Ͳ�{���v&�q\�'��x���ޥi���қט=��|pu���	��09���@��V�/�
,��S�9�m���� �n>$tm�Y���2���fN��c4J�@a�(vFŹ��7�x$�w�9�̿�Gz@�U�X����T�"�t�;~$!<�G��Q����1ٝ�*�L��J�OqUg�~T���TQYo�j7�nS4� h�3�>`���*Ǹ�c�X��%ʊ/wx��܇Z�<��:T,�e���D㨿<�,���Qb,u���ˁ��S�]k�3I��S�Z�f�V�!y��ԄVd�B�ȏ3I�8��E2�G��,��HK�	��n�8:�kӿ<ɬ?�
h�m����&>�_���4�
���f�D�]|ۓ�u�%|��������VU�Y�xĈdUsg��k�Wǒ���_W(B�ɿ(��Z\2�Ţ���u���'�1�rTs���*����򊤦3�%{x���sd�m�'ŏ ���lCUN����$�.�\�tH=[��o�U�ϭ����!Cy��x$*D������-R>��1�H�($�
Y}Q��U�H�(��k+�&SFq��pM$?K ���b�>��]�� �.e�R3�����
��+�nxP=D���6�Q$"���A���=\��!��Ob���qI!��F�j�.An��a���Z�P�U�ۺ���mw��"�E�s7�����<�CHS�W�$XwZ�(E���N��"�4�x�0��l���[x�����V��	�����*Ân(IC�N���7K�I�;��ap�g�)l����%}����,w��4B��#Q�ۗ2�L4 3�[�
P" "q�:[a
ϻ9w�hJ!|rPhO��]�£�V����ou��e}���U��$m��!��[�{I���z��rŻ}������%��b֘FU�̘����jU͵͊����Xsv	Ȭ+Yn���b�Ç�rl�	�*NA�*�}N��	�l�����x^�;��^�P��ލJ��_�A�	�B%sUa�qa�bԓ� 7k#��ݪ�I��V&��ھ���\ŵ�8Q�A����_WI���1�{�z�o��9~�����"����¦̑u�3�7�Z��]�xFl��c�>��`�~��#�L�t1�@˘�+P)I�� {��3�U	�'D��h|/��zz�Br��TR��u�g܋:z�?���T3���!LP9�z^;cƉ�ߠ2�eq�����5�l��f�?'���8�D��T��quAp&�S�Q�����v����nyTf%E�����<���v����������,�C�d���IR���j,Rm�#�rZHƎ���y5NM$���en��G�uF��Fɮ��5^�oTp�{��-e� �����(Xj☘B�� @�u��#�8�BWp������� �y$[�)l����5Q�>A&�L7��d�O�3�/	6>2�*�F��p�/�G�~����/а����
ہ���m#R�i��e��c:D�G���ʏzw&�h�oT���;�N3+�Bh8?�i���/@䈆g~^M���=Q�ɥ6<hd�R�� ����un���<�z59�.�D3�!]�;@�mA��讍���Y+$H��m����H�?�:Po���4j��/�����y毣�����v0�ǜ�k�
�e���zU$>L??a��?VO �A��� ��B\��. �͆Fe��p�����c�(d���7|gX)�PI�B�ڝ*mm����'�ݮ��:��g�<:��>-Y1��GpṚ���Z��=��ޮ���g����&z�1�H,s��ŀG���*�`���A�t@L�gjҝ���θm^�D�d�1��#�]"<~P�k��нl� B�"��Ze$.	�a�;8��Z�h��F��v���*9�9�yc!e�p�զ�*�����M���u��i.L��%�XU���L��y���{�u�EY��i�)��� �`Z][`�^P1��`�ΫPb9v*�G��X'�u#sI�����q��Ϻ��|�~t��u�1O(�s{'���l��r��_.�$�� �ΓY=G�dBnC���1�V���w[���SF��2�*Hlϳ鼍I{�op9 ]i�|Bg��VoSy>>�~����|�qP^>�}�h����nҥ����:�a�r��ZQ���dBP�XG~ܕXn�Z�h��?C��%�H���+Ԕ�mh���hO8S�-4?���Z�w��Y��=y&��@���_���a�!�t�C���(T�Uj������Tt+uv�O�%H����V��& �V�m"Fx�#�>�Y��0���zeN+O>.��@���jk�H-]��m���x+B3�R�����u2g����B�el���j�0&�a{)G�o$�jks�NI���v�G���OD1�ô�ĽK���\NL�V�7�Au��S�����.�����bM�V���/)~�Yyg�1+�B\{N^8�z\΁�D˯�{� ^�ǐfkoj�)�ԣma�k��]	/}��[1�g����l}׈������M<��l�L*@�B���6&�*pa�b�\�AuY�3�
�<Ae�}R;��H����y[ 2%���l�"�
m!H4{��0���qg���#ލ��!��������&�AEb�œ�)��`�-ڔpV$��Γ��AC�S$vp�)���r��`�[W��$�}k��6�~�ɭ��;��)�'�[��/k8�K�~^n'���X;q�A?��-�]K�6b�xN!��X���q_��-�nI��s�bPRo�K}�t��2�':�U'��,�,[���Fp�S��N�����=��P��q�9Ŗ��u>�RN���dF|�YJ����A��א[�c"�ֻ=�/��KL��fF���?��?�u _e m��=�i�����+8����z3٤:��hĲ�YE�X� g^Y��cEo	�.%FUK�ݥۘ�+c��f2e1!S���n���L &�Q@!�v��۲�]��4o`��a���7g����٨��n.e!0]qx��[�uM�V�/F���!%^ ����A~'%���6 �Iv���r��!)Mm��0V���=��*7e}��h�"Ȯ�F�&�"FTS4ƃߜ� �.�+�gw�L�9�6��yt�,��:��c%�țQ���� &�qܿ��Tl�_��C�P�:p�X���R��~"����.5���P��'=��70q�&�ŝ\>��w�r�"l�a��+o��>��:;W�d��:U癏.A]���T����
����*��� �O�7eWH1�#6 �Bb,!m�L �9����\��/?��ueW�Aj�޷ƞ����3��1�/p��y�{�?��q���b����1�%�݆)�"S�{�W�QAx7�Ѩ��=n]����b\]l�<\�ŧRj�R��?�PQ��Ah�h�9��?�70<�����N�7�#��%�_�1y�<-a��F7�*�ˊdo%�	;\6,��{X�X���
ۧ3hwS\3v�M�M��P�Kkx�
D��fɨ�	"�}U�+��R�hiI����q�=BݓClp���u����j�N �nT����21p��7L��"*a1�t��ҠZ'�z�w��$�=U�h~�eo���]JN5%����&Yr�	J�9g����t�G�Ό?��x?w�����>q!NJS�&;�Ry��9�-}��n �LҰt��n��~3����D)�E��6U������等G�ˁ���I����ʱh0ucy��?��D�Z�nY_��aƋ96w�n��K�|@��	���C��iْ��i��`@��t:e>�������ׯ�w���(J�5���U� S�4���/������i�)!"3�nY|�f-�c�
z�m�GY�WN."�&� ����'�&���v�}?�H�mW>9�܆T/�X��>��x�\j��sI�j�6�j�Oc���Di�S�W������� �YP�ڵ���+�9ċ��ѹ�
('���L���s�c�̡�,��Q9~o5_Q+���A��a�P6�w<� /o�b��,	�|�׌L��O4�¦O]���Gx�V�l�%ƨI���ZR��l�rU^������c��J%њ�Vɥ3v9�V�׍H�m�z�62	׶��"�YLeD�%��Dyw���v�&��.���QB��v>�-�NH��"�i1?U<Xa3NT��BI��I6�H�"I���N�r�)�\�3���fu�r}H���P��1}�"0��u��<�ɹl�2!a�8=~����z��+��(�_�{~�dV�t9ht�C�gT�˿��ɰǭ|�
�(�<�R�"�[��X�[-���tB'�+.������1E`r�d��#��.Q�["�a%�V	#�� �Ĭ뗄��KZs٫#C�E�Z��*�
�����Tɮũ�OT�ܝK�Yy��ϝ�$7�N��d.c:
>�����!��i��;q2���&��;k��x��ʇ�yLK2nc<�9�? ��/M��,r'�Z��lT{�Cw�E���n(` �?��p6���|�.�x�]�oq}�d9�����ғ$#���V]ٲ;��icss��+R �Vt��� Z���݊������&�#�{��:�4� �R���C�M��E���d��v�i$�ۋ����.������B�q`Y%D(�F!Y���#٣�G���d?8�B���-%�D1<VY���k\��8�Ʀ��b�%H}�u�L��
�&B�0�M��פ���0LQ�o���Bც"`�?��8MT�L��aם�u6�a%��wn��*��t�*��qYfQ
���T��GЏZFbd|�y��lA�w�?C>1�Acp|Op^�xtd��x~G�"�5R�/��H*�fs��y�@�.�ig����|����]Q��,��n��
����c
 sw�J}�ۉ�cZ�x�Ձ��3cHP�}x�43�MH�9>�r���6��w��Mv�1L�_r8iR:��p�� �,�.��5���5,v�+g
�|��A�!����ŗ���������W,��^�B�3����&E(� ����\i(@�	���~�p��U�p���O��$Lb��z�}�PS���PrҰG�B�;6%�)�gX��<�Y_�)Y��ޥq��/�q�ל7&���M���3�i2��|k��hX$p*���׃�h7~��'o����Op�KU��1it=e
>	2��8����'(��3��!��$&�8����.J�(�5�x�U�����^F�mw��v��W�|������D��6��i�@�nE�����D�[g"� #Bw��*�8������Mp�k[�[�
KW6w��	�ܖhwR��F�l�~�!{�BJgh$�[�[N�=��&t�s(���}�L�W3n����e���_��J�8���>
s�+O�7L��|]�E��x(7�l�����Fb��vSW���#�l�Ɣ�e>��7U!��5$�]�Ë��pi'ӹsʱ�mJ&^eȏ䃙�yX�7ѓ<��o.5�������NԦ5�Ĉ>U�Lb�/�z����0;������+X��4X~�S��&��j_��}�؋I&�iW�i;i1C�*��61(��aJ#���;'$Q�o�~� �N[�����5���8y�o���� ����Qo�W���!���u��Ua+�mIЉ�.�<䋕ض���HalQ�.��qn<5�n��M��H�I�"<"�G�E p��REոs�XfWi=�:�)�X=�i�������L"Od�Gu�l��ނ4
g8K���ɢ-5��F�ĉ���Z/*#N���8�f���)ԧo^�W�|M{�J�EZM�>]�B����%R��Ѧ[lFju����B��:p�)▧�b�D�^���Yr@�@��&�XM��2�|1N*��KX8�a��|��2oL��g��E7���4~�	���CH����EECU�ʲSWqݾԉ��?
U�Vt�H�W�N��m��@��/訩$��E9Gi�`Z�o㙙^�Vx������\GۖX���]zH�X�<b^ѭ�1M����vea�5]}�0zq�^�LD-��P�:��ۄ�1�_V�/�L�����e&�+�F��~�Af9��S���E��F9�M��mF�J+)�\�0ȶO1�~� ��<��FGܠo�� �my�LV�|��pK=k������<dT-�R�{ͱVJ�&i�W�Mc-�RV���_�aQh�k�Km�
���gs���p6ob�%N��M�k<����&���F ��}���pd����V)r�ؼ�'e�|�����'b�D׎�	"���&�N���&w��̒_��8%�nH��"��c5h���1�H̚y�M!���B�g&�}�����)[X0�X��˒�	�6�Y��(Č�8�?��P��o�ڸ�q�׋��O((<��&Jtҝ:�O�-J�Ѩhs��%�$��n e�D�3Z�ډ�y��:�Y���Z���[/�<�Rxʨ�ދp�wB=��f�~u�U-+)
��'��-��z'zc���m�K��i����>#лw��^�����V��٪/&`���lk�&�PO�]��':�x��͖���ZT�k���;�[��"��t,b�
�;y_�
�{1�ؤC�Ԟ��`j7���"|G��l��ox�aq�RK��%��(c+��X�/��G�g��8�R��i��IJo��M�W�2�ѱ��pCyT�m��������6��(��>��Y�z��r��X(Ƅ�ca��[Kz�&,I�[�������U��xn^����x � ����E���z�(*�rp����pD眾�Q9��4ul���2�Z�g�Z�5�b�F}.��d?�ͨ���@�r�b|Аd�gQ�Ғ}���8�-Ɯ�2iA�W���Oz��	ѓ�,'^l�Fqʧ��RJ��v��$��J�Ū���$��ށ 9���M�ξ��nh�y�)�i�J'�#٭�N����R�����I��Ҹvu����Ӂ�X�#�4����޴�D�G-����#[Da�/�ʠ��u�G��[6�X{�����Z'j�ಢ��@1��q�S�9���ѳcف��`��%P$!.�"���+B�<��_�\S�0e��_.�{�_� nD&��&�i��#���~����0J���?����\��x-��7��Z����@�gT���(��}VI`�G��L!wF�ٔYy3i<�<6�ґ�t�!8Y`v+=��"��"��3B�;�M���=�n#i��"��3��~�3�~��)�	�U`iD�Gn�"`�..�u4 �#�(�QJ�MW��ts��}�3�0�y7?��x�H%�@u����u��̿q�b�Wy1hB�ಊ�6����|�51n��2em��x��=�.�1�2‣����!�2o:�z�
���-���,V)	4	S.���Bw�^�b�z�����M�J�� K�F�th[��S+v4���+�[77)h 2�'����<������
٠4��14�I�q)�-�
x�E�+�������F�4�J�-x��I�3i{���l����H�J����w�'BOS�-+�.6��$A�n")-bc�[w9�nZ�m�5�*�?\ue��@"D��2�?N5 ِp%km�Wy�t��B�lf�:��'M�{pa�^b�?Lh��|��"O=W|iu`��8�m�W������5c�B�C���m|��p��7b��z�cݽ��Ώ��3l�J����<p���+m�	(�U�*�-�W�x���V�}�
;RC�3�:-��%p�¡��r��a� I�8��b���Y�d_���au��`Z����گm|����`Xy�ۂ��Q��d�Q8�'��C}7�0U�Fp.iz�Ǵ^b�#X3Ǎ$ēw�S@����K�vgt����+� �3�w��!���+�{��[J?�L�ԻiY�s֗�$i�;g��y���T,��8�^|�:�?���>[W�@���ߏ݋�44���;j1l�|}���Kz�ڢ�u�廩��T�SfWZ�����H2��h��Si�X>������ܒ���&(��;��tW�r*��B��Ի�L�t���QE/$䤳`[��`t��91v�7�t�XF(�K,���M�X����2X�V�Rq�r�u�����5�\���8�	����p#�F|�C=C�)���卽��y)Xe�~~��j��e�B���LX,��C�n��	[+p�O1�B8�|��q�N�r�)?3_� }�ڣ���o�۠�i�7��O��a��*������Qb���p��Uyv��Yث�\��-�e�9�愻��~��OeY�_h��؏���F��Bi�����JYR)Ǒz͠X�ڡI�ۤ�=�{r�㪯�����-	��C�ml���4x �:F�	�mY�4C/�;����A�R�+��w�p��Om�����	�Ԥ���C�b}y�S[(X���=�f���`��ƃ�S�I߆�.G��l�g~�k��+F�=I��)+�*��;X}e׸���s��zHDl^KX����M� u˕��l�>���_���񓕺��[B}���uD���noa���KF!0�*!�ȧ4����'���?��@�ro�V��SQ�p��&z6{*�l 1\::cRb�.nZo\������J=��SN�ȵ};�J��])�! ���]-�;�.��+୸���yN��k�Nċ9���x1ɩ�̆1y<{�MQ�N�:\ݺ�谚Y�K,����\?A�}IrJ�B+�2
�s{��g<��+P۠ZqW�\T�����x5>�XQ>���H�\� �z�5��JN�y�F���x�q�;����������	k���PS�Y�T��>���俹��8����t��j� `��|�ˌ�֫C@�+��z���P1�oku|@!�B�����%.L��(��q���T��	��\��U�?�@Z�*�\`�y���PϤ�[�t��^/+�J\��GT����WP���B�z示�N
��3�4����7�0O�M6|��Nɔt���x�b2c�H	��$��-��~���A,��3�q�;����8+:n������_�*���ஔ&��+�Iw~��-k#�ӥ��̃�ZGT�q��|"Ј�)��\����={���4���\k�@�'����4��.����)ջ2���tp�9��	l��$U��O��;k��ٌ����N���|���_�r��ʬ��lv�m� k����^B���7l�����y��M�`����Y���SF��*�:����n�O�x9>Z!��a�;Bx&υ
��'��V��ԃ��o��؂iaF(���hF$W���;��`�_n��y�L��ևTF�ʠ|����\U!h�և��R|��{��:q�d}͸��m3���uh~5jC)�}܃� �åZr4���]�?�R���y�X�ť�2O�MId�_ld	�I0]id��R�EH�h"x����bR�Ų�Z0N+
��oWV�#�d�����tz��ܓA���k�'~1���Q4|�<�s�(�ƾs�W��e\��֖1��WO*yRloƶ� �����|]�ތ=�/�f �ֻmO�^iȲ>>����P��ٚ��9Mm�-�a�xn-��nK�j��W_ޝ�g�VC���I���3x���i�#rM��aw.Ȣ�g<t`�O�zNqٖ��U�� ��rǬ#���zo���O!���W1�t�@�NՌ����n��j��WT���Ѩ�_���_��MYR̦S=���+B!8@��Gl���NҠ��I�\N˙JLQl�B(o�=5��t�H�0���+Ю��ȗ8�UG�hZ{�����bօ��؏�l��C�4�h~�a��wu�O=ꌴ�m��:�j2��4Y��f��՗��}e�Kl�E�9���|M�b���W:�D�*�"�B7 ͼ�Ø�L��⤢(�L�h%T���4G�o�ܱ�9�b�6R���w&��˂|�T����ط��:�]�c��3B��Νz�oG�5�k�MS�/>�V�O�;��*"�$K��ע�,騲~է&�.��G�"����b�K�%<���(�{Z���C�\75A���ƻ�/��w�'{K,��\;L�YS�0-��;_�0i�)��k�慃�%�*%�B�Y�]K�9寮h*+��hM�zP?`Jub�J�4�ip��oH��%%�^q�[�e�]���EW��|�?'�@L��a��,M"I��r#`����$�ӧ+��>V9l֙��h���M28�̀<�T��ъpS�?߼i{sd�����@�Hz�"m�i�1�Eb[�=�k�U�7\43��*�g���t��221F�ilbT�q��'j��ؼ�����||ZB��$Y�,xͨDp���+����+���$1FK��
�6	��['�G��8�\�e�6�kض��!2��pV�E�2+��b�̄E%�(���yثr���l:<� +�S��--�˧q��fx[��W/����-6���#]j�Y�A�x�8P� ���p�����c������a�W�^���Z;��Y|�-�-��&i�)m�Ί"֮ക����IV��v2f|-��Z�H����^(\���֩z�Y	S�Mր�)��P�+]��9V��~����,���Tت5�iܨ���f�N2-�F���ċ7.��&h{��D�@�[��u��t�_3D�	��K����N"dۆ��ܔ���=�ϖ�ybl�牞쀵��N.��9��@K�d0<��$�zUZ��0/��v���$�y�MŖ��(�e�*��cw�z]o�Ͱ��u���~CG"[]V�*�8w�=Q��UjJtwV���Դ���}Ƛ��� �G��SE��쀧ۤ�1�A��6T�~P��nc�dUN�����w>A�;�O�d9k[`}�]�6�OQ>�� �Ⱥ��`� ��Jp��-՜9�n�@.��-�2��� V�G�� ]�p0���j� lR*�>c2����������?�$� �*z�7(��f��(�����o~ 2!��"Z���!��(q�`����a
�����%ki܁fۀ��|����F�tR�	���*Zr��?%QA�3f|X�`�-+�?�y�����BR��9\uẤQ˓��X��T~c����L Ko4u �52Z{�p�e�¥{���z� �@4&+_�t�;qt���_'@�x<�=8w��B� �'"(�y�W��婕�����ϼqC�=�yQ �G8�Ӓ�_�.{=3o�FU�KCb�:чɦL�j;<T��<cw�OA�p�W]��ϕ=r���=�����|q��m�T	���HU#r�u(��#kGyCm�8�%��+���^-h6����������7��>W e�z���[@B���ONG�?^wؖ�c�d�2�.ݨ����� �ӭ�o��.6=�3HBU�y���$�ש�3��W~v�W�<D
#2�?d��Dkm�J��V,
 &�Ks���Ďr�)&�&/u��v1z����Y��!�L��EO��_Š����JF���8`y�dT�r��H�!����M�6�LF�tA� `��i���j?�d}վɕ\I�:1$Tł_��e�Y��ýYo��{�����J����%�]Q�G�g���OF�NU��`�'֑�G4���Փg�ܨ�4XL+��Ӵ`�J.��{Q���Z�e����)P����t,��C�B��F"1��EV��ʔѴwt�-�E���,Č �t7�!a7�y��F��@c8�Y�
�$t�(�za�j
7i���ɩ��=b_~l�:�d5����AKʏk�Qz[U���LN��W�a�7`s�S3!u`]~Kr舛��.����� O�{/�Gu�� Zu�#��M˘xX ��y��d� �+U��L �Zp7�����r�]��#Z������&�_\��f����I��H��RT��8`@q�D[��漼I��]�X/U*q�ڹQ�ж�����+����'4��:)��w�i"�v��{m�D����*�ޓ?��hh�3���w?ɷAi.Ѳ���2Tj|�NZOW�!8d�����fƙx����ݢ����� -�	���
x#�O!k*^#�"M7�j�`�;+���ެ��}^
T{;�������Jb%6����@�%OWC�%+��|���Ɔ��\�"�\��k��l�u���;Hb��?���x�Yc�m��Q��z���'������N�o⿖4$�����l`��W���W(��3Q"�0~�W��`��IE�H��D֩�8�d�9��v#�*�0"��l��>�}�æ&iݥ��;���t+�b��V,FC^��_��u]Ca����B�����4�ژ}�XÛ���K�	�θ	3�M�x\3�,��=��d߻452I����%�=n���p�K(��|�����@l�� yg.�-L4���[Z�/�t�D+H�:`$�$x@���W�H��[p��)��%�y�i��gDt�永�`���;@�M4F��̮-(��b�e{)�!Y�\ĦX[�JD=�ͧ��k犩�Nq��97� ��j,Z�}D������2��g�v�I��v-_ЅS��ƄzW���E��,��o��FAs�j�=4����5,�!�W�>tG���>�\RQQ3X��Hh�H�j�l�_T��l�Ƭ�[�X��v��b
��4�2-[���>��j�m���28]���#��u���h��+���S�n㷻��1�[\9�S�:a��ܶ���X0Nn��L���CQ��t'��t��o�����8�@e@�,��=����6_=�xe��i��zە@��EC�|1��`J���`�u���ʪX�Z-�Caǆ
�&w�é�;����O���R��ܶ�s��Z�p�8}V[���d��d��2C��HOZ���� o;�)�h�&iȐg��s2���㆒�Y|��q����������|��t:������fJ.,m�h
��m�J�����	�0ԟ�WWߡ��Q�r�9��O����K��5���T��8�z����77	�C�����&�ꜷl���P�ؗx"I���^y��ltq1�Q�W lO 1E�-"ϔ�`˸V�6��
[����D���}L7�x���Q���5T#|���������H�+��Ix�/������wj�>P{�:�@jj5i6G�c�����˖���2����������G���,޹�-~��:���>kx����W���`� ��*0��Se�1���QZ.��笐��/�LN:P�+u�┐��}��)��R$w�,��i���4��΃&�y��F^x��WO�*��i��:�)�r>n��2���J��DИ������F>ƹ�.%H\�K-�����$h��ܵw�[z1|�M��VZ����}�a���R%C��O�f����7�Y�i��:��"z-�QE@=��*��W7D˴,�v*^&5����c����O]qk�2�;2zAR� k��φ���#��CP���36$Ta)�$�����!���v�l[[����Jt%&��t�>J�Ն���Ǫ~E�F�ؓ�OJ�-�v��qӺ�E�TԘh�e�ߡ�7� �U�_8m�DMӳ�"�z��h?H@�9D���)�Ȣ8o3�A�=v��6�h�,��=��n:��o�r�+�MQf����q�i��5��<d��:���?,/���$S�]�Dh���0ϋ�����{ ��; �E$QHh�7R�8Ȗ��	�V8^����D'���Vք�� ^Z�\v���yn�4U������:�Ф� 2�.u�g��S�)�Rx��-d"m��y��_L�sx�����Ȳ�C��T�fv�J5�Q��Ї8@����;���0jn��)����^;�U�L?��/o����́��
h��]��Hq��~�_��B�uΒ�=�u�����$�6q�n6+��6M��zM����P��5�E�h(jd�u󻧛��Cd�n�}��B1࿹��t�����g����
�G��vE������8��W��35����M7,�Fg�5ew�]:��H���UOx��Nd�x��l�����y���ѥh�T�WrF!�[&�z�S��D0�$Z�"z�6˘��k"�\uiS���i�	��`ݼ,�������b���!C�=�6@��3�v���H����&xvp$d���R.H���и�2��`��lxR,SR�y���Y�^��w ��7�����nH*�F�cL?����8�r��
4l�3��rpOؠ�X������ ����	��HdOSZЖ�	��o�<.��JuUO��+¾��b�?��2�����7�U �I��fa@Ej�0�p��1"�v�^3~��)��4RS��]m|Ke��/�~ؘş�O��Ύ���nV�����Gp�c�m�ʦ�%:�yG�1҇y=׏��}�q���o����\��GY��/��ӏz7��~�|������ʙ�ߠ�ף�F��i,# 8E�3�B(a�mly;)���uo' _��If;8in1�.O�-\  �����԰�~�<�͎�h��Ve�bU�5ffG�:L.x�1��3��������кv�0�c�- �.9L���J���N�=X�;�<�iyrI�whY�B��c��	:^������=��%��:3�p����j��j�BӸ�����R*իެ�C�3��@�Ov�V���z}�_g�H�O=��,	T��T������ ��ŠAԀy2)]��S��|������D�����������=@����;��
z�U[q(��O�+����2��u��m�̊�6��������Z�J	����r��V���%�"��y-̕��/��0dup�2�`XK*������]�����#�B���9	$G�R���܍��F9;l�&⾶�S��ƻ�{f�Y\�=ӷ�ݟ�x�'�Xj���f�k�����*j�M�Cc��j�9Ya��4 ���}�����EF
�%N�\6C�+3Օ�d*l�k�q��XHW���� �n�k믱�-���ʢ��yG���Y�-�E$0�'���v�O�YG�ɩq�:i���tM��NO'�yJ�-<��v���9F3UEo�L�>K�rZu1�6}o6G��ZY���0����J�׿�P�:��ݕ[,q�,
������9�	Ҵ��4��mAv��~S�P+%���R������iK�fG�Y7�x�����oN��+��qf��7Q ~�`w\���K�z�]c��A�&E�I�nW���3?�zɨ�6(�U��_�L]͍sǇ��ǫ�	�$�b$����1~6�:�Kع��, :&
�+L48�Y�?�0�p�'��b�m�p_�8�?|���zR��ɕ	 )9v�h8�G�9�]n�!Ri�4�����'m�=pJq�4��ޞ���7<.*YW^_���x�����3LK=E�i*(D1��T��r��2mD��ׯ��ܡKd�d�//�|�T2v�֬��� ��$�S:�F��;�;E�{���I�\���}Ǘ�G| ^�Ym�{ϓD�����,�����	�:@� � 5��
\�P��9�i�$��,�fnP�:��T�������-�,�7KB5HC�J�����Fjt�.��w� $%��fH�Ã�8���zj���H��qn���k|i�ea���Tޤ���6���F.�?gSvʙx�ΒF��0^b3Y��*�%?�-(�"���'o4���.�[K
Bw+u��%�U|~:3w�������am�#�}Ϟ+j	���Z ��\\`�mG�;b�$�1����9+{)5�L�!�D�x�Kyl�k�z�N�Y���jF������f��ne	���V����`�Xa�@��u!���bv�o�ga�֝5�놸r�o�p>`��$�^��D��[��hdP�OZ���b��3�O�2�+��i�O�Ko��h h�W���	H���`�"2*�i�<���-�5��&3��#d�p{���Ew�S��a��G��Z43�0�7���^��%9S*�yH�/�M��=�_�F#�e�_x���!ĕ�[L3]��Z:���*���X0���4T4Yۊ�&$m��|��R�$��v���g;>b/��	ɟ��@�(ʿ`|k���C-7��g�*P�u����f���O��$	I�� \ɣ}A�\I���EЎu����v�L���@JO���?�A0&��}�#��P�6�4�`"v3�߅����r	Y�H�l��?��
��g]���Zt�Ȣ,��d�38+x
*y�.��x<0��Y'�ok�������"c��d8��7`ۅa����P���7Љ�Ψ��-h���m�_	���E�j��#2PZ�>9��+��y�F�ՙx�	�W�!�M�Ny|FԲ���Y�����õp�u ��oI�^�����N<_��J��抑�beS��9�K��ڪn���³wR(������L-(JX����]�ݽp���>������њs�ƒ�6Q�wF�|�0��`j���/�*LQ,��1�ҕ�'GB��\�qc(UPm��H����!,d7_�΍�7n7���W����ѱ�1�oȺ�P���B�	�=�L�B����G�ßEB��b:��<r�L����2^N�gx��9G���;1A�^{����m�a�����_f6��ô<U�N>a���k���	\����*5%\���B�R9���0���|0���m��3B-���?P����k��pA'�a��{Q1l=���%}��s}{�Țp�kV?%��{\~�E�?'��ui�I+�ZE�Ā�'� ��Im*mҩ�M��\}��� �4�p�w.I��Y�3�L�-�}]�L�n��L�Uz���f��H~j���R�!�#15��D�32l�q2����1LYp���a
(X��g��yq쮕��7�Z&f�O�(�X4�e�"�.V�y-�%|�oǁ#Y,U�H钸��5�]�j.f�4[��E�4�y�������+6dx���Ԃr�m��Ƴl�W���S95���!�	�� ����� ���dq*yƎ5�O��u����3��w=���(f�h��A�1L����J���3$��L�s�E�s�(��3�U�xs	e��Ù�2bM^[����0L�غ#�X {;r�����p���ݲ���I� m�T�h�	XS��N¿L ��
�%9���hÜ���Wv�2���A.5�t��U�Y�O>��n����}Gj��}ڎz.-�L3�)�րt%�뇟�?a�s ���g	}�%f ����UK2�ʍKT�m��4S��8��b"�4�U�]hA1�Ro�ͰK8�4��Hy��@b�7�~��JW ��Hch��T��V�� �i��o�2����H1a�qz�0����Q�К�sڵ� 9&��i�_l� 8�����N��G�pt�:@��ް݇,���bE�+��S(���o$���
K����et�s��p>jM�>nI�a#��R(�������UIKPM�X�Ѵ�2�	6w�؈��\�.q�����7d�ⷓ�(n����b�C�5"��-�mԦ)g�ԐM��#��,"*�*w׫�B6�H��T_�Qh �ן�7�g���c����1�@�5���dr�96���O�oL��х� �^��f�响�_�aﶹښ���b��Z�WK�B�׾#4���tA��Ն��0	<ď���U;	:���8ϳc�Hg��җLASlpN�d{M�o�,t~�`��|���Ȋos��U��2��S��ޚg:�B�!1WB��Y��(�n�b�Y��9��U@;I<<�'ҽʰ]9΄�s?�Ei�N��6�"[Mr?q�I->*��x2Z��l(������{���
���fO�Á,S�S���q:c�>&�����v���O�W�(a%Ʋ-�5�LА90��\�_?���!x�O�]��^��f �y�W�a������_��&ר@6;,@ړ^�(#�m�������nE�W�I�oN"��
��r�}�d���Iԏ#p�E�L��)�f�E���!�B����(p����%��W��F�a%2s�'��eRt��L��6-���J(e��y4���Y�����%[�Ǻ�	AZu�S�d�q����R�C�Y��]e����V���1	k�I상�0�&�	����!�AA wSo�u�t�9S��V��C~8j�m��z�����-ֻ�!�̬�*嶫�2��uѣ<*J��]Q���F%�Y���m70���3镍*�ƣ)�i��]��Q��#�1�x��	!V��|��܅HN��z����D��\{�����Uo)J��2Q%G�x�л�J�.�iOE� P<��a[� XY���j���n��>��;�p~��p7t������e��t���ܩYj���=GT��1��K���n|�'
�)������*�NaF�)I��S�|�"Utk����8\~ 5���)GG�D��_N�zK�y �>��sX&���]�&�ՑL��A����I�#�ASQ��{fɀ)dX�;��+�m��ƭ�.Ǆ�X`�׾ĳ�}{�b��d�$ŀӿ6���6-�� ���s��܏����o;���F�5�@��B�A��$��|M�IYW�k߬�暭��S,�*(G�W$���ͷKa����,�6֭��"����J��4j��"e�����W=�d�}�D1S��)|d�n���@��h�o��v��w����'j_ ��I��:q��
���g%�<g�$� f�J�&@�%��]���-X��,2�t&�^(jq���F������Ƈ;���{,�~H�
���̵R_b���?����c>��',(R�:�B@B�J���K�Y�B��8G>R�(<�J���W@���F��_��(^�T44����D�I&��~�^����z������!ˀ԰�а@��6��0�Ǐ	Tc�.yO1���R��qf��7$���5B�v�6�pٌ����N�� ]S�2H�3I2��EHZ��
�v�4욤������w̥_[�[�%XP�R�\^x�۪�n����|��3k����\4٠�@ܛ�)�+	{^���-�r�d�JX�]5NW�}�����hL�K�9/�ā��Sr���{=:hh�C`�F|{���;�!dV�H��^���b��۫-h�[�����Ŷ+�8x|�ܑ_��(pP��P����D�������F�Zb�����8�>?�U}��^3<T�J���P�P�խ�7u>�h�{C�\?��t�Dʸ1���O�ڕɼdWϘ����_@0����.�rҀ��rTN :~�kq����MI�o��q�=�Q�w���|U�I�ؔ��`2
Rg�@	�脤dsM7Z�>7n� �-�^3�N�h�!ի=6X`��c'>ч���~(�V�!:+O�_����U���G��L�d�IZvKWz|A3�t ���N����Q�ﱘ/ɍI�"O�8�u�	n�$�M����Jbd]���xnp
��%M�Fz��l�[升�����"1($�;9 #A@_��E�����̥¥����� �p63�~�:��6u��Q3�?�(���6��hۚ2�O�[��`2H�T��f��(%R�hħ����b�D�r�g~�M/?r�����y��[��TXQ���
�z�b��N���P.����gƙ-� ��/�o��T��Ӧ�?�T����M���z�Aw�\6����=����D�-�ⴈ��*��a�Y۬�|֓LFGg�˙��t�'�*?�z��b��d1m_�h\�H�b���f�����r*$8q���P��{J��n�� �*���C*�?��˄s���?#�����h6���%-��� x&�f��#����S�s��]Uk��u:�)hC�˃����a��;w�:E�z���F�Q��pI��6z�����.�u?��o(�yGT����5|�oR.���m"T�����y��[�t��� lϪ�ͮ�t �>_�����RK�))��W���8&�%�����u�+��x�?a�9�8P�"���l:�S�I'撻0J�/h�'�9�F��v�Z��(:�DF0⛥�<����@"�xc#ȮUw�g ��� {8���6Fx��`�� ���h(�H��3��}�)���P�3�A]��	���{���le���Q���;Õ/ّ��Tn3��S�Η�VЄ�k��M-���{:��V~��͠�e��
�[�ћ8Aiw�t���ĕ���(|��P4�29�r�I�;��$ݖ�O%m~����Q"�J��Ӊ ȱt@�8��d8΀��/"sA3��o�q49��\�{;�]�
��h-�L�e���G=��G�s�g��:e?{���FEQ*�E|���WZn��Wo,ϕ&���q�M�IOf��6�̽&uO��!�������%0�?j|u����{(�^܌�g$M��jn=-d"�Z���e����H�~~$�D�P�Q[C���I��s��~��$�A�O�V���ܤ�Lcv�*�x�]e��H
�,:e/Mz��{�)
Cl���6����`?�*Q�ߎ���oB��LR&$�M\`e���-J�4���j�_�]�+���1&�$�r�{�\x�L���-*+��K��\[^J��v���`��_�c�^ܫ��R��2�O=w���(<ns�c����~6�cn�ޜ �;@G�k���z^i��w���'����W�b�oИ06�^`!{"0-������ArN�t�l'p?�븙����2��0�{*��@�E�D��%c [��^���*�t��KG�V!�{���c[� �.��!�!�;F�%����_�aL8��H��Y����*4|��R�
��,�K��1YV9�-�N����'$Ĵp�m�+PŁDM�4	��t����,����=h���\�V��)/���!I��RB�!���R��_�/+���d>j��%�al�V�?T��@v5c��{|��lfQ�<�?w!A	v$"/rՆ{���4��4{�ݷ�=$)���'����9�a��	�������ZF&��$~P�u�tOjsg\�?�E���}����2G��!jd�V�n����X�� @���J�id�~��d����`{�:������1zU�k��Q7R�H�	ѫ�����;i�c3L�0���dp�x�Ll�����H�D�b}k�3o����\�/F	�He����y�;���9��dNEd.�Ux��[�1or�-"�������/�2�J��N&)		-h=HqRf�Ԝ�N��;g��R��c(?����g��3���%d>H�/���j]% !nF!G��n� :��� g̴�1�gHv��W�>��gyE5�A�_P���P���ƅS����hA��}8\b��9��<�����3��2�Q����c"N��& ��ЇKb�7)o;�2Y�(u�`�R`-�\�O��j�Yj��j�,do�e�g%�Cr�4�Ki`��_��qb?lÊ���O�~y&�1#'���k{
�
���L��ړ�,Mi�P���R�AF�s5PӲ���󼌡y�@��ڎ�Ŭ7�����<��7�7�>X�'����_�����)w?��S��*'��֌m[���,/U�cdJ���c#7� �R��R^��ABT��Y�H��f�~�O�ޗoV	rC?����Di�>��>^n<t���bX�]Fub���k�1�c#l!�|�З�~�Ď�ڿ�g��R�Ø��I�$�*
2�z�b���-ʃ����`�`� #�H��t���f�@�:MG�q�/�]�!�o�̡-��|�]!�?�E1�=�~|�� z��
>d7��Շ��h�ət�{2e��kl�]T���V� "��|���*i�c�N��K7��N���"�:(g���&g�cc����}|t��G�8�pq"�"i���Ru\���y<u�{uzt ��j�򌭳�<@y��C�[�\8�s��Zo0�Z�C�0��S�
��6Q���Y�x�{$���hk^B_�xG"/�'!��Ws�����V�f[��<��'��r�A`�T��k���<(�t����%͚c�Ge&����-��������`qhԊ�GB�r�6�X����M��Nq�XsA����
3��5.�,���㪨z\W�m��n�êv���9�o0�D�Smbg0�x�8�J������[$v�pٟ��������tZ���G�����h�Gy��(�?4�ڋU���@m<\���u}��+d���wU7�H����7R6����G�'�Rj u��N����n�9+���z�*��7D�� ��i䤵@���#X��@�pTp���P�x�ΏTf�`�T����_8˞Չ�ӣ������$���#w D?�8n�L�ֽ�|4�k>��<m�d0~��Ȯ�a�r^[끅sT��zЉ�EZʁ�߮ _��C �3	�AJ|� ���ž�A黷Cv
D��1�g0I 玺��f(��E9	�n�*�HQL1l�yl3AF����Bљތ��`�.����G���=Et>���؉E���L��4����C0�6ls.��w1&uu��S	�W�d�>ˉV��P3�;��s�����A[��'U+8"���?#��K��(
�%2�i�[����pQ5߫�GHH}�������5����(� ��]���m���?�RV��vE�n̎-���W�q⑖y->�z+���\�أ�8�/延�t����+�Y�w�8RS?rKJK�LF�Ȁ/lֽ1=�:%��}��ѽ2E���m����Ա,��g��9�J��s@5������c=+��T᧙ �̒:	�C�H�u�By�5�_dv~aeF�Z`�e�2��/g㎷[B����B#IY2
b�t�L��`)<ゲ�0�fa�v�_NM_�~����e�԰@����F^�z�C�5��CC�H�I-Soq�q4����v�0�:�.�������!�e@X�h��vBC�/S��-�>/��`J#��^`hϔT�VXb)R�kl�k�HA�W HFg�+����������9O�7#��P8tX�gس���6,+�QV
��8Ǖ?l (����Ǆ����	G!��
B����n��C-��jf[ESc��+p���$�P����2��яR�$��^�ϟ����B(+�$��m[,)Am��Ohp <D��6;��ya���Lػ9���R����=w��,&���VR�*\k=$p�$���v�����	҅�2嚔�"}�i�a����:#C�s��<���/B����e�fl[�?�u\��R�cw�4`)Ȟ��M;���#s6h��3��sy��'�����%B�L���W��F�� ������|���23�����*\悵򊸔Va��dO����^��E��{�<���p�ݜ��X�B�)A|��PV��t�&����w<����Q�`�(�Р� �&�?�}�*��c/`	�뼬v/=��#�h�����[dI�E�s����ֈr�δ����Y���6�#��KDi�ŤV�^k�v���H�����R�G�}V=���_�(:j�gT n�5CY>��b��ԯ!n؅�ɍ�5�0���/i*�3���0������)��9��//��4�d����j�rl"c�FC�,�> �b;�R�r6��w�X�5�p& +c��~��f�hħ���9z!W��._I*SS�@b�,���*��㧂"�{�I�MRJS;,|;w�譍^���e�������i_���:��Zz4��e,Z�A :�#s�;���a�R�w�Dx������5��m�c��R���-U�U�dt���ɾ��r�������&�ۻ�	�����M5�a$���s�x��~���e#�3����#��0�F�m�̈́~k�H��y�Ȁ�ҎY�&ň�ѩ�K��C ��dS�۔��-?��	1v�Bb�����L;Q�C��\{6��
N�FaWs���)�R�H����q��5��e�홼	�h�C�`3�H�<ؘmc�E��쑬M�{U���[�z��(��43��X8\F�c�(���hf����}��L|� �=�����y�bqCr��6mAc���d�A��D�;7��� W�΢���P��&<�4U��>L�JC��k:�v�2�<X��?H~���{�D��4Qi�d�;2`!��Ha�ɰ �/D���f_�̍q�oĦ� ���8]��W�)/�]a]=�b*|���	�T��Y� WG���Zν�wE�|�ܡ��f����<�T�qV�i�cX 9[n+x�o$�qi�:u���oߪ�2[?Kw�t�x\\��S	_�C2:k��@2�񳃵f^����b?���+"'�+���ճ�CF�؎vgcRl��T�VM��2�<�A�b���{r-�U��{��ϘQ=�.
N �[�뵮�EEt�s�K6����u����v�q"���~χ����V?�b3���4�qN7��/�����Eg�G�ɯ�����o<krB�p[?�B9:=$E(bK����E.�6kN�΅�䜜����G�v��*���>�\��^�Ez���L(����£vx}�w��A�}o* �e��Z�~���I���1�7��F䖿�3m&N<en��t&��h�ie0X�e�&��+ o�*��k�2fY���4�R|����܅F���J�ky�Ҩ�>��9��6��s/��5>x��Yy0�^��5X2�(.2���G�/AGg+@g�/�} ��R�S,D>S����d-���ҋ+ I֘�-k}��E��Nu^h��Z";΍T��nNBs�����j3�B���S酡c$�o�o�F؄���pw��J��B��M�ye�ΨSӇ22xIaa?�����k� �\� -���W����a�i*f�ۄ`��P�l�O)3���o̬��A���|E��������0��t�Q�?��j��C�8�>��̹9^���n7'S&vK�>�m��L/��cj�|>c���6m���w���H��}0�%@�&)1�LG��7�=�9UG�U �'`��$�G���;!*�г��P�܎�:�u�lc*�?
{R���*6�� T����F�R���h^=�����5ޘ�I��!Gq7n}?�_�Z��9$�lT}N�1z�&�yѵ�����f�L"\�d�4S�d���!y�x��%W�{a��0*�|��Թ��Ĕ�SbƘئo��f��e�Q�-�&`ռ���Q�ua<N�C7m����A��:��b���L��aNFs���n�NXV�R3�H��³��qd�Y !������b��p
h�]��y��7��`%�W�{U	� N��HWd�.�x8�Q�����)���L���F5�M!�U�}����G�:A���ʪ�:!c������2x�G��[������m�X�U����͓�%�\�x�$�V���4^`��e� z[��[�Ѷ�[����QjInd.�zpo*t��`�?7��4��`�o�\��1�RyN�|��ο��7�Eș������ܺo];���3�(S�� 0��I�����!�Îo��G��yr��	y�hyJ�lL��,�Xb��Rc�}X�9��%�p~��KN; �ӑV~X��5����!��R�v0Y��-/s\��?%���o�*tW�7�72wBBi]߶�	g�� �0�氿��
�9R�@&-��{����4EU��8��q*�-�j�G��ˮ>Ʉ6��µ��<�nJ��apEk�_Y�T�q�?AQ�����.��j,6�}|�������T��$~�/���G'�]��x��@dtͺi��߇�+��fDr��yũ�t��/���rD��V\�O�`P=��"�(�E���"��9NY)>���oG��li�=h���h�7���{Gm����W�}3�K�&'w��';���}������e �c<g�/]������ZO(O�N�e�ՠ�<
��Պi��l�,�-6�C+ �U����G*e3�aq�s�Gx��	/��O	_�H���:Σ����pvP)��n�1����>�c�0MSA�&���a�"@+\j7�	��)�W�D����:�g��i�s��������S~�~w��?��2Z����p<}��Ôs�&�Aě��>�ↈ��
E{o.���<a�%?-��d x�f�,�c�0�L>���;3 �e���C�o�Z1�l�1���z�ڰ�)��i���������������Af.��X}��>��<���x���q(��pn�(7��?��;�~Vj�H�8'K��)�@r�f*̟�~|��d6(יP���=Q�����xb���m1�#��΂t�r��|�`���Y$���8x�����oW���\M4��V�CФ-\g���H��51���:�CP�17:�e���[���̸a�!���)a^H�.�{���Nз�o*�Ky����n �މ�Ѐ�՗㘀��w脝���������(h e��'�M<'�I�])����#{����?��}�;ѡ\^_M4p���blc9�#�94�JI�h1�?�^���5R�LZ0��p˂���d	©���l�3.�T@��gs�K.�j8񻿌�:O3�?��G13J����L���A+��!x[��+�3��o7��	��릤P=Q�9�G�|+�^{J��������id<��#�����M��`4�����!z��pNJS�T_�zz�غҿ0�&����n�7�⨞N�y40(i{���F�z�1A�|�E�����4ҡ��E�L�=g�s��V�b.�'Ӏ��2��L,
ո 3�_/o��`ҧ�龮	ed~\�{�q�z��{D�]M*�����RJ����x����2/�����UVt��8ZC@��膖������
�F�	����f�{1P땬�#������O�U+�������@�=�<v���s����p�F�8�؏O.�ۈ�	�2<�����L�f��1�$#>p���y��RU)�@��ǯ�<fǎIW��Ib%(^�B/�o�}�0<���˶�]1L�\�I�,�¶QM-)�7{��LzEr^�Pw��|�/9��)��x5�h:q��M�:�_�v�G�x�΁"�u�[���+V�j��"�7چ὇����n��o�,�ZS�Z��P���5�)���Q#~l��XN����G�����Q�����>��{��觋o�i �(�ޠe�U����
�5� �+a*��iyv�E�h)�EP���j{Z0���d�,�Y�d�V��^��,�8�A��*�0U���(ϐݟ��p��'O�Ϛ����U0Xa^�� �+���z��]�\+� ���9�¦�ʰYÛ�ri�4du�����dE��SR�^� �0��W"���!�]�p^���^�&���A-R��B��v��r���8~�m���N7c���ח#��5tӳ��c����ņ�ؗ���ڣoA[��� �Ho\8�K����A�{^�D���Г���1@笕q�:�nWe��9��"n��hL�:�!_�D�eU���\i��t��-^O�&:�#�󉔯�>���4�!�3��V�l�ekr�3�q%^�>�8Ppn5޲R�)eu����YR�x�-���g��ȥ��J^q����g:a��9yx�}.6��̤ٵ�gk���D�7$��F�TX	efN�l��5qKo�!��Wr����W��,Һٳ8#	�� �;ᐸ��Oq=��=0��� )�3�P@m��+�=U<A�~�h1}Ɯ�p�~A�������bT0�LW��a�{���U�5%J}G􃦍���5l��p|�����Zw����c�_����������Ȁ�̷qD�k�U�~�dw���o'3�b1D��KZ6u��Y�x%��'�*o�!���Ô���0)�	���XuGio��+�i�$<[������o�	�b�6ϊ�<���|(6�	puz֞&vŰQ��to��Ά�<�H�d�Ћ3�Tw_��7�.��
á�m҄S��cZ) ��B�b��^&[Hܧt��2I�i�� XZ�����>�q�P����0�>��e��Ss�b��no��!��oN'M���c7�y��I���bn�魭g�Z�2ǎ�F=�G��he��B��i���"u��5��׺w�շ�l@����҉�	�sad�kY��B�5��������t�=ǊN$.B���l��\4���,�=Z֮��i�-�BXǿ��C��I�gx���嫴CĤ?�y��Z!4��S�mR��蒩3X���4o�W�b@�|2�1B
k
v�����~k<�����i�ꁗ;�0=ωQM+$�R��8���<��%���rӶj�-9�M����,�����G���-�Qx5�aGn2���qUH��
��h�l��٭�CW���_Z42�3rb�|�l�T���$�7����oX�P�6p�{B�É 0i�cb�v�$LhZ�@�M�W!�\�h ���� ��D]OP��z�9�>3P����Qޯ��j+KE���!�f��ܗ�����	E�y1��p�� DjE��\�ӡ��r�m�I;�ǭ5�Έ�������Cȏ�*�J����V""���;zd��KP[Yi5"@2�l%ʿ%�b\O�|Ƴ�y[�67�5��
�'»<Cn�ntb"{������G�W55���F�+kxY�:6'D�AGeY���D/�b �YmU�p�F#�B��V�AH�>�ކ����H���ԆW
�z��-fW�wWz�4ӫEDk�ƿV�d#���J������v����H�Lt0^�Y����IaS6:�38r:JI��{5�3O��B�e�I�䷹vzhMqM�*Hզs�}�o���M���}M� $�<eLF	�h�F^K�����g�2���|��� ��|��mKaĲQ�P��,5k�d�R��1]M�ζ��-���Sz3�Z�t�~�z/�.��������T��.��8��8v��N�s	�����v�+}�Q04g�ї��'1ȍ�[CI�2���K?3oԛ��G��FƬ��8�Z�ׁ\
�$i�uwe3��]��ɍeM��ceԿN�>@���m�� *�߆R�L��jE�0F��Q���R��ؤ$t�j��.q�i�D�iȈ
=�݉�o�-���&u?&��uN������VM���ۿ8��@+��-��Hz��ݣ=�/��Ruo�F�w�й��ouY����ev�g�>`7p�@��7�^��`��V��ߓA��q��{�M���������������_ �[��#3�0n�u�rB��c�,��1�b����t~�<6��h��Z<E=ەx#s�C�(�ގ�H��=��à1����h��v�YT�qHecܴw͍�f^os0�_��cߘ��	�e�>��m,D�|]�$X�$m��դ�n��� � �^Aj�R���i ��	$w��B�噗F�5���^�#��U����-��P���<E�OY�)|�Ȝ��<��^��	�Lj?�W�_��G����0y�o��v�0�:�����2�܌��oY������z�x��͋m�C	Ku��>�
W~"�GJw�]�?i�O�ƿ�|���\S�n�	�P,�T�Ƴ�&b��B�A�p��x����ZZ���
8��N6��p-H�v^6�9�z��DX���jo�w�{�]�S�\�J�І�XH��2`��fk�	��}$b���U��ߎ	��X������ؽ�������[�]����6���#�	���4��u>�����i�q��n��L�K�,M����:��ހR�7��lP��Þ���F�m�c��އ�]0� )�Q�:� j{
�M�)��b,U����lˡ&:cF��3�%_P	�rĿ!1�ٽb��6���bl�@uu�G��%���Aǂ4��ztK���n�츲�pJ�^/WA�b8oB�J�9��ʦݺG\[.���-�]ԍq�!K��;10�%�#C��u�QS�������݊q ����;�s{���K�����	2�Р�:�:�I���'VM��V���x������H V'�п��$����]�Y�ILi���>� �^�S��8(�e�������d7g(}ߖ��C�KӢ���>�Ԩԟ�j�P]j'^��;�BW�rw�\��L7*/��Z��eU(c�P�c6��\�����q��p�9zI���e�#�;?3<�托�s˰���Nؽ�׎���"&զ�_��+y�^�Lf����F�;
<eQ��2�Ҿ�?�F�g?�|��0d&�*���}�X�4���&ܱ�Mm&�T/YR�@�UM��5��G�5�ܠ�+�G�1}��_r�Uu�VLlN���������}(PC��0oZ3�?��c��4V9&��xZȝ�1�]���5B-d�����ﺻϥ���]���* �D����?b�|�8{��l�x��7��&O>r+X��S�[9�hpu���Wӄ���*{�Y�8]��&��V�Q��F��A��Vu
B�S�-k]�1�ڒ�9��\�<��錥U�ӯ2�yn�5P3������ɟu޺�S<��.X�d�M��@V�Z;�~�s��O-�w-��;w�g���gz��:��K�Ԥ��j�p��ik��f8�lw�{S1��P��`��S��g��ڋ��d���xe(IBe9��O�Ѱp�ѴkN.C�3��Q@ߤ�{�W�F������T\`��B`�0l*'�Pq�K�9��k��A��9
hS6��r��ż�J6�Wx��>�����D5=�<ۚg g�����5���eO��<��N����}�����Gl�JMZ�����!�It|�:�l�~��SB62Q�Tc��q~��R��m��TQ��ӄ����.�^�7i��{�Le��dt���uH|��\e�3v*��tzy6d�^ʐ΍��Uw·�͕��A>�a�wn����w|���s����ۗ/*����|ԙ�{�F/W�F���������Ұ,���"g�=�r׉��d��P�eL��4�s��~Cr��״��2��@�{5��^���!�U�{᠟y㼕&��U��)ɋZ��Ǧ��ڎ�Zy�,Fi��9�1ط`ݩ�O�3jbo"�%��*���Zo�N��'�#X��#Y5��?��� ��S&�7X�,Vx��k��<�=5�|t�ׁvb�_>��u[��9�������#q��2eD��4p�w�bD�DQX�5�%Z<��/P��M���s~�/�ImsW�� ��M]R?⦒2��[IB�Q�uc�n�zZ�a�<�_W��|St�R����W�����&�� ��*�
2�sb�El�5�Q�Cb���'�"�st��o��-L�ѷ�f��%5���0�2iA2�4�'�k�\��~$_[�+�b��u�<QSlX��|�b$���'�`�Y?EV����hIG�{�ɹB%(��a��+-R�	���e\��0�,�FԎ��;�Z���&�l�]�Q��	It��z�(�X��F@*p̹>��X=Nc���T�ڣ�[�	$�Es��s/nc�a�h�{E���5:+b�Qi"U�VP��6����)�D��:�o�B����A{�r��BT��� ܲ�ep�a��&�ɳ&�E���͉`!�A���]2�iѾ���=�EE*Ev�b;"���)����lNG5퓏q^Y_�XAk�_/��G��Bl���C������^%i|E+V�[�صD <T�d���5������M��1KG$%���!ρ�l(�����r;|w��KB��)`���A�3H�!\4�ȜD,�f�+�����}i�c�{���|�:� ��6䌖��}��C��SH��}�A�T��῵�9�ז�a�v�Lp��U�M)
M�m���Y0��|�@�cK��@g�VG�=��*_�O�ϴ�b=��9�+HSz*�\0f�%D|�@_O#d\>���"���ʄ��K+~����R�U�L
���[�-l�����8�X]�kV�yû̈́��3�1�5a�4��8���~��z`�3����Ϗ�5����PY�K��^�
�|Ǻq�=(r�����r��N
W'#�*U0q`����-Φ��Y�e&l�'?��}���u%IpnfT�N�ե�ԅ��ѱ�ϟ�ڎ��q���VpH�����`���XY'No�[�Z�B0`�n��\`���t���m?5�E��NP��3
��I�
�7�����LۨI���#	[b���[6��]钱l"��İs8�G�R�07{A�U��^�zZ뫂�g4iw��f@D-��IP�TGQ`��,�)g����"��fh�0���B�-�����e%�^j��������W�{�#��K��. ���1����\��Hn��ݶ6�C��+�D�o��� �	��R��#�fw9�bću�)�mJ6ċ�"τ�D>�:H/S���ۅ��P���^��R�	B�A����f�(�l9�o�������)��JV����>ټFTZЭM6�Zg@�"zW��b���u0����ݟ6+�񸊣@��O,��Y�}�=�O5���q�VB{�@)�<���һŒQm1���-<��ٕu�z�mljħ�VZЏn~�ԣ梤[ͷ�#W�z�����1��%.��	zzXq�xӃX�̑���]yo�܇EH�P<+;YX�Q����?@]�N�d&`��$0nI�@طJ�&��4����:I9�[�V��:���C�����u�P,r���d�%���3�ŕ�>�_��H��5=i���Z��W"|t:�e�[�����5�Y�-��dU���N3��/���xuR��zΚ����K��`X��v�������e�������݋�3��`�墁:'W#��,��=�dH.�5����uy�ޚm�|SXP�=_݁]���	FU��@��ـ���`o=� ˼3��5�LZz�
ZN����������Ip�S��ф�����BA��?�w�&&e,.�c���z�85M��U����<��� c?Wo�/��&�Qn�;P�S_��PTF~�M���k�2�	?��$hN��5��L\��2�wۺ	~��a�}�:�I�,�� �ao�������x�}�1i��Y�=��c;R�&�m�����q��
�o��\��
r����҇J�+n��EE����E����.F���:~�/�M�o{`���}���h䵸�9���&o$a�x]���%C/[B�I����R��TW-)?q�ڍ�E1(-&8���f�H)�gП�<$]F�]z��������$�d�o&��U�kw+*�=;>ݩ�	����&\���Ń���u�zj��j�G�����T�/B��p:�����`��5n o���
�}sN�����B��ԓ��)�=�d2i���M�Φ��B�>L�=?L[�����B��䓚�^��/�}/t���U��_FOQ�h�`��{�X����&����	_Cݝbar�<�(���K��8dVA3�6��а�~KLl��T�2���ɛ�~�}������w�X���ݮ�a	���|�!�J�d$�Xe�} *| 9�U&����ӛ3��;�_��=��聯�l/Q�ʩ�����њ����'�GhR*Z�	++��t���g��!o��D��\�z5���c�񀺣uK��v��O�\�:eb	.@��Zc�]���ds�;)�����2 ����{�B��%[�	�N�Ѱ<�F�8`��$||O�Qa ���.I/�2�bL#�	��/�������VR��{U�2��k��UI�sHO�.�97,�G���]"����J��ұ��ļg4Ƿ�a9X��I�)�{����D� s@o~'�%T�C���/+���C�j/&6t��I���@JJ]B�;�F�qe�;~+��E,hjKV"]��vm��w�M�{���_� ?�!�R���]�]��Ȁ�މ�ڡ��u7���I�����P�#�� �Q�����P����:y���ڢ�X������SD�X����7̍�mV���m��]Z�#����-��@�Y���L���@t2/��n�`��T�f/ ���1�&������]AfNc��8����=M�l���{(m^ �wx	ǽ{b���9��!��}�joD�2B�$��rJ�Bٮ���hh�84��O���a=�	����,���,_ʲ�'��Ok@����>�j6580W��u�[�a�N�����G����5?������cQI"��=�g����H����M\}���?�{���!S��']�^�eP'm���ȱj2��D��Ц��`Y���Ͷ�V]�F�4��i�P��`r6%�0V�ʳ��4��]�%{r��C~��$�G���l�O����U�\.ߎ�D4�z���˾ɉ{��\���L�,5b�_�3>��9A�o�+m�MY"�>�?��3[=U��ŭҙ`�g4y�ʱ1W�]���2�ύ��T��*�vQ�G�)夋3����,XM��-���kQ�d��euf5�@��'E�k�m`2в:�[���x(g+�g�� t���������<pW �gzS��?'γMN6\HC�e ��E%42h���\�,2�dY��֏eє��Ҏ��w� ޑ卼� �za�Z��3\�+���ξU.�ԇ�ʜ8�<I� d��ǈIzX�e*
!(*w��L�x��uU\��N��e��ޔC�XlAYc+�]�>T�%	�W�k/���
��@ww�*I������]��I�wp�]<��9��'|�|�� �q�WF�; ԝ��_�D�=�)[?՘3C-#�J���*�PM��U;��F*���i`	��smw��'  '�� �@�7@tm&��Ɲq�@�Q�GdՄ�`��-�xd��Ű��My򇟿��|ԙ��&x�s����	�b��G�ʻf��w�Y?]����np��W�����L����y�mԖ��=+m@�`�_J��9���<\�̰��\��ahS��d��������{)� �A�|��c)�_���^/
M� `�|`����X7�ru\O��sΦoKr�07�������hZ���kJ�ʉ-%O�{c!��Mw~�ē����D��ъr���BheH�dA�&�:�R��nC�
��A��� vE3��V�̡	�q����		썠��m:�hi��
�fx�x@���4���1��]eaaQFs�"y��m2��Y���<�����lE�«�����\�(B{�"7�Øъ<�O�b4ի��^��_��tTO!�����bs�ě:n��I�*�j����d�2�r��t�!oT�%��[L�߄J2�xڀ�wu�-=����'�1O9�	W���J
ۃ����")�����y�7��y��s���㘼�͋�6s�"�ǪN���.��X9�6��U�cO[�-�rh{$��t�4�Û%$��q1wɗRY��� �Z�jxhYyD{�s��G�!�=͠�t !�pFi4k�RJ���uc0T�\��S���l�o�#ͷ�9d{#�F�{�se����#��(~!c��7of��KWZ]V�������c+�=t�G^ ��Z�$���U�E�p~��}_�G6�g,�Q�nihI�Z,j#1,8vs�n'a+��Q�K� �Ϛ���ͶD��Y��Jb=�r���6&�)���,���r����8�8�g��1����2�c^��X5M<i)7?&���zԾt؇�-�W����C�<�#�G+��FRʄ��4�.!�+!��[Q'0�0V���.����<��p|͕&k͆�@��tu#Yy�(.-�j!)���TBvG�E�$ֺIС`K,œ5)��%�] b�6?�D�O�����$��y�K���97b/�� ͡�Ƴ{%�}�hjB�n��v���N�	W���s���AH���V;�K��!���c���qf�K ���܈lvF���BMsg�+�k=ք�~"��o���sܴ�аV��e����D�7Co�by�$-ɑ���lv�����o��.��s�|ߜ�j#�x
�w��g���p�~��� ͚�=�W��.R�!����7��uw "&���ٻJ����0��0�y-R�,1�{i�Nۓ���
��}�L�	V�on:��aƁ8�5�P�T���ȢN�b��+%Z`>w��[lP�D�A�28Te6o�.5�"C���.�8m���jԕ�qj��c��$aJ[~�ݫq�㣬��El����q}���Fw~��M	���tVC�&)86��T�=c�5�4�c�g�Ί�e*|J��Q����d~w>�����V6~��� NQ�����8�dl>�S�o��._oGP��4cͧ}6�_Ռ�238Z���N���o�G"��pМ�w�cG$z��#J�ϳ>���1R3��iz�ԁ P�'9�M�AI��+�)�m��� yD��z�}=�	�b�о�������9V��"\1+��|�r����_j��vkK��h�x���Q3O�ߒ��Nn���p�F+gg��.G��,z�{������Z�bڃ���엚�I�K�+���q�g��Q$���.�L/>�s�@2��V�>%��_��}E"&�G�"��I���r���K���e�� �;2,lm����`�И�W2nԾ�a�:��+[p ���A#s��]�Y�W���@<A]E^A�s����^ᑫL��E͟�Ud��^�i㷡vO}�uEZ������9�C��?:�4S1:�=,�"��x��l�.@�7AC2_wP
�(No��{���C�+hc%��h��vq��q��@���~`U7�'+
�Rw�n݅CT�+���5=B��$¤�<�k�<�m
�(Y�׻?CFib�jgO�""ү��_y�wc�cFuyMktKʾ�-��R�eu=��8�3Κ'/�!�!U���󏄿��<�ejfv%%+�StN `�>y��R6wP.�.O,�͹ќ�c��L���$>_YMθ@�
G���_��\���� hh�t��0���|��h�
2P�(�! �d��Y�*J�N��h�?~}�W��}�d�0����Zr%tgd�F�L��5�#ޑ{���;��&�C���f�s--ѹ��ae�+M�4s��7������zg�6b'4�+J��i-<n�N�=ڈ�������Ḳ����Ne�I1��a���-M�y���M&�G}�"z�MJ��Ѥ��5Id@�:|,D)�3�4I�f�T�1�
�>��F�|�V����n���:�2Ō8��ŮSɖF�yާ>���	��:_[��ϱ�Y��ɸxɇo4��r���9�'��跸0=���n�m�5(?4� t'9��ϙ��hE:ԁ�j1O3<�Y����!B�R�a��e��7��G|x2ھ����[MwO��?��?<q�T�ɇiV�������IW"Qe��L�٨�BMXDw᭬37�J�$ �c~���$����_;�M~cn�;�`�5Z�U�Vu]������B|���A᧕��؜ �d�ئş���1����(�8g`>%�oJ�7�E�����&=�9�L^�W�3�a��M���쇉
qL������`Bcp�x��6��z|Z<
w�\P���A�[Pvu��#9�M�е�{H������ŧ � ɤ��J7�s�>j�<������M`�h ���͇�{�1�	ͺ7�m�G�/�pY�z�/|ǣ>z/�e������ʇ�}�˔��匶m��ŏ%|GQ��� �ǯ!���X�a_R�0*�J��K�4���4u��E�D������p[�:��=i�Ʒ��������a4{�[݉��AJq���De�eZ~���=�.`��=�y(��Ȉ�a�p�#�� ��� QQ,<��vrm���S<
�@������*G��NH�Ѕ##*X���05��輶oU,���҂�+���K��
@l�_f}Jx>&�k��E���27V�у�{c��䅩����G���y����W��t����e:��b�O[9�j �{hM����D �kKz���,������TV�A���~��?ᜀ6"ݧn9]�J�,V.C�p'�y~���5 ���Q5:I��8\$L�6���NLO�~%[nn����|}��OE��
��	��7�
 ��5�PǏ�x[*��)�9��z��m�X�*eZ�\��b� ��&��	��A�r-�҈��r�Rs#���˸Wa�A�,E2�9�&#�.�k��o��)mt��*���نQ�㜼���M����������ۆ!�l�S]&�%K��3By�������>�G����^����/�|�LD�F�⧮��i����0el������8q�ʾ�g�뉸6R��ȇ�$u�V�],��C5k|E۟�x8<�Nc��h�h*�=��ȒF����2@u� -��6�4ԲN���FzM�Nr��t��#��
Y�E��#�wR�'���C�*��睽z��d��	�DG������f���v�.�� �8�S:p$
 h���u,��"�)T�$&ޡ��O�o;vZ�����l��d+_�O�)�ְ�e=��֗����!��J��kBJ�ƛG�LT���P除�Z�g�	�D
��ͫ;�F��`7��֗�9��(��2��e��5�g|���ݹg �2q�ާ�/ ��������X���Д{�����ٵDJ3-�{ug��8KO C����mW��mhսVn��M)���uSio�bΧπxB�W�]��)o�A2�Dʴ�r�I7���[���*�(�j83:�t���cca2ߤe��;�s��J7b��v�<#���J��H;��XHQ='~]�>��ɮn�"����A��8��?�jWMKV̝ᇆ@�rdi�L?�?>ŝR_J�Ћe{����.B��;]��K�Z����Ι,*�*�*}�F^k"%!�CE���p���/�v���U��M[A*f�*BPN��$��R�3i�t��ض�'�u��7)<��2�-=2؞�etA�Z�e�H�5��ա捧���ie{���Td���-} _r�/6�sGVꬢ�3ۭ�������c
f�p�$O�"��l��׉xƶ����W����yw%���7��o��K
+��`�ƽ���yF�����m�-�S�	z����u4��'>����9��*���J1��ְףP�v�p�:�e�_�j�����j<R6�r� �J?1�k�1J֭#,�(O�#Hg'5��s�l01Y)��N39�A���4I��X>���YsK�N��ʱ����V*�!*�vev���Q�6�""��%��<���v��H�_�@�p�~���~��<\A�O�I�?`�/��)3�hğؗ�o���Qb�u��U/�&hK�n�$����ʅ�P'�	��
a��Ȱ~.i� j��pW���Ơ�	������Q�˶ �������[	# �m����<�Io�I$�6�rpЪ�ǙhҲ��1A�R�.��#F_v6���&�uC�$�?O��/hEr:��a�<tcr��u�YMlR�i���(u`��hg��_����"f[K���tܢT��b���ޚ�\�R*I~���5�)J�8�h���	�RS��ȀTLuZ;�ǵLF����@.�	~[CN�{���Z�n܌�������&�	c%(��,��"%�a�ڱ�'�h��WPD�X$ ����]��D��^.� ��~�x㟪�:�>(�xp���_I�Hy��q����`}#��p[Öh�z�?���0�����~{I8���`��U6|��l'����4��5�ȕ���f6�F�IV��)�#�(h��K��v��Pz�O�2"7\:����i��̆K=4Jcf0��pNNش�EQ���+1f��ie�U��H�,n�޴��U�g*$o	���+SGw/���E/��d7����۔��Q���rE�4g��9�o���~,T2,ؙ�@����넷/��݃�=*��Hص0��!���`
�,�[
��{��;�٣��D���i~�|�� P�-�&p�h�{�g��=	軄�7��%nX���Y��s��p1�\���1-s��ڦ*�,��(<��,�VV`��*Z�r��z�>r��RO��p}�S@i�k^�Wf�����ܫ�l1f�ck$�p�#�N�.�;�~�����&���/E ŷ�1��N�j�BO�$-,�Z�>�jB�8'EI:�U/}
�j�[	�3���se0ɢ
	����(qo�n�y"YeTW��ο�ӧ9[�[b+�w��cW8��z�x:��p"8x�1�j���Ф��S9��ѣG�j]v����Pq>_ݭ�T���w�8%8���VA�[��}bW,.�*�'���7ώ}tٓ\:�Y�G͚m�!���Ck�W��VLn���_O���j�=.� /h�6q���%�v+���Gq$�:1V��WO�Fw�o�6�ct��׊�Q�A�l�AQ�8+�t*����a�s�S�{�B:�.�;N�Y��^�)X\T���Y��1�}�r"�-f1Q������{Ц����Tj�4�gT��!�i��� $'RBx~4'�b}����s>��b���L���K0v����۽:2���L 	Ղ�ƁD2R�)��W�`���c%q���z����E�q�00Ǖp�;��8�f?��%\y��Uo�&i嚊�!��S��w~S��я6��vo-�g���D��/�0����m�}$��튡�r(TB�t���~��.���̊��M�8��ʅD�;��o��撙3�ry����9ąL��ea��Y�up��k;�m��K�l,5�������P
�E-��7$P�r��o-D������_���[dh�f�o���I[��U�xc7�:Ѫ7r�I+�v���I�}�:��j���	��zp9��N�(ǽ�.1{I_�{�F�x����>^�������L��9]�=�6�������f����d�:���)w%w����^�?�*S*�h��˩�A��R>cV�� �`!�j��w��Nӭ�ɜ��xҬ��E��w�+� b4�P2��!_>%4����-1|�Bze�,oA�{CM�us��*L�hS�(��p��i>�qֈ-��\��|$�$Ӡ·�#�?U�<�)�7���tn7�U^�}a.��斢�-.���B]�S��(@fY`�:H�ÕO�[�a�5̃9-�ԅ�R�������HN�z)Y!�8ul~��Ϩ,�7/1w�韹R�4��i�A��^��_ ��]J`hm~=@CH�r�� &�x�U�\�Ɯy鶢��L�7V������+��r��c�o䁟@ow�@���ۅ!`��gqn��3�b=@�uNZ��=&�tN�Y�$ɋg��N�
մ~��B\�妌�����1Kd�8cTK~�h&��Ӈ�qb� �������k,/�[�){�[Qwjł�"wWi����Y1��q&H���Pg�9Tp0��.�<N�x�/i�\��lE��)ء��^liԒԭ��I�M�=�z��j���� ��Wt�i=���ތ�ښW�����θ���x
U~7ۜ���,3�ܷ�|}W6!$���V)~���a1�̕1_�wؿ�z�je���gs���HטE$�@������I��
���J�z;��t�0��U!g���%���SM}{�"��.�] ��~�K^�Ƭ2�g�4��]��J��![�ؗYV�7����Y��RH�h[KP	�L�Hݐ� ��(Ű��c{�$��t�r�5-���uqQ�5��&�eO����=�}(�@L�q���yO����ׁv�d	[�Fe�;�܋����X�7�06���N�}޿�R�����+~��\4�V4�K�\�%��[ѭ�I|�_�Oz����R�].)�\���,TPn�F�,|B�R����~EM�h���U���A�#���NXf�!�lE[�'v�s�gPg��m*�9GJ���H�2�C�y���������2�[�yӝ�!�;N�Iֳ3pկ@?�	�f;��%�쓶�����-�. WhZ=�����N�i~vj`�2���iHh<AzU���RT��L�~�	#������P���Yf��G��19��cH�:���l 9~����O��Y��*�G�c���ɚ��.2���yL�f�J�%�̐J,K6�i�W@s͕�����!b[,�����'/�'Р��L�L�-h��oU�c��[� �0�ٻ¹f�����i#|_���R;�VĤwi�?���#��F]����V5D=� ;�A^��<|�C-� -Z}a4x|��J����%o^.V���l�;��w���܃$��B=��Q*�l�Z����z�vÂv��J�z}���O[���Lu��g���aV��EI��9��_�.��d��;=V�����H0���<������0��\�[a=�o�Om������T��bFo��
���K�h��d��1���a�����a���X�-�J���Qgn=���7�?�;��JN�?��T�q�
�s�6�5r����*�F�O�C�Gi���G��L� �#0w�'�xaBUA�y�u>�l����зKmJ���
J����@Z���.�dP�T�w:�/�LE��� ~��A'l�\:��}�3�~�> D�4{D��N�t�>5w��{����r�����GF{��Q.^N����ݕ�M�����N�}*��犈�c9n�^o��?���� j�a�t���P8{V��ۀ썸�0��\�m��A���,�Ui�g��G�܋�O���zy���O�h3{�[	Njlx<S��BAR��h����h�> .���ܯ#���j/�op���t�p8�]��MJ�/$�!'�:��'27�۷�1SʥA�mR^�R���v��H���҇RZ��F����qǐ���f��O�ο����y
9pܣ�pz��>U�_�IQ�j�l�N�gP�_(܃�*������&���ʈ7؏T��e�������@�!.TYU��Kے��BQZ$U?K�ќAl��̀�y�0*�΢L/x�S)�Q6}y*z6�Jd%�ڎ�B�ԇ�sb��C��9Q5�R����:�]��S]\�������	{&�f|����E��ܺ�]��́>@|���	��Ԣ�N�'K���x�@,�G�����B[��p�K�UHP��"�ھZջ�2,ވ�4��C�"^�Ǜy�j�\9ˎ2a��ˈ�x$C4������E� �0�[�|ԇ,��������M(^�=Si��`x)�������F�F�5��dI��7�S�/C%��֯�6�M$�j�3��P�[G�	��sj�aܲ��F���f����1M`h$�D�.�0X��U�+�2��DX�B���������"�"���hU����£[� O����R�ѥ�[�-��l��ф����F�dC�z��b���@�VO
��r�מ1���SN��r��i�"--��p0XU=f���wI��L�	���.�����W�Bǒi~tu5�aۘo�[V��[6ht��?��0u��[�)_W3|�5��-�`�H�e��u�Aw��%�����q���Go����E����`"^�)e�>Ϥ�\��!���"s�R�����h�H�ؒ��Y'��GY��W5+�\��- W�W&�O��d�!���fz;ء�7��
��������u��*\��D���gR;C$H]܍:��T�w�p+=��*{�F+����DK�@ ���)�y����b���Sy�C�g�8)�Gċ�L^���[ li�:e��%0Q�*Zϑ�)X���+�(�٦��JM5F$�|p��1�dޞb�b�
��7�����-��<��_��l(�E�pe�l=*+c�����[��9~��|Ƕ��Q�%:,ex�b�T��1)���u���J+'~�Tڱ�a�$.q��y��T�C0�$Mx�ײ�W�Xk���<���ط9+"�u�s�s�<:��d���=��yFr�GQ|�&�Js�$���1�_C٘�i�M!��4���E�k���Ս�~��_i�9왘7֬>���S�G���S�e�j�Ҙ�>@���d�I���Z�X��q bH'^��Tc�Ҧy��ZJOc�;y�9��/�dB�F��MHԠ���D�'A��x���@f;TD;�?�|A��a� ���������l������/���>�?����P��oQgl8��	Sq�dZ���-�QQ�:����r�D�@�sP��z�H�����E#>C&:|�V
��g1H�i�L�be,0�=��l��X��~�&����������13Z���=J�@V�bP�TK��)e�b#}���D�1)�u��;X�JLr�:v;�E
��� ����肢&O�[��I�U6�Uq��d�����=^�􂗘��z?�4��&��I��n���W߸
O�VzJ��3��\0V4����o�I��<Nܔ�#�-j�x���G��_.��@4�@�#���ȉps��6�A��)+��iy���e3׵� ���G���y���ab�n]��b4��<Q�m1u�#�f�vB/��I�����9�@
�E�͸)�^K0%��/o�7�ؕ�b�Z�kX�������k�w��g(�b:T]}�0�c�u6�3Y�W�Mb��5���$��
��8��Vm!EM7�#�J	�l���-�2�5�L��s	.�dG��.�vL���g�"Ʉ]tpM�����l��0�3鶉���7a>�S�+�}��G\�;�M�^��ύ����w�7s�0AX6�-ژ���s���x����p���'�B�^�ZWѶ��m�u>Ya���?ބ,�Ap����[��]-8@�V�|��\��!Rs!�iD��0�x���j�b�+�x���U��E�QJW�� ˽���	�S|m�g�+"�㾊��D��|X�!����y��|��G)� �-���}֞|�F��ի�J�_|2�0��˷썠�Qz!�+'�7Gw���'nI����6�H�  ��zwZ�_	�@x��ۉ�p:l���� Kt�D�v�M��0�9��-�^� ��}Ó^ϐI�����]�ud�]�cy�Ȋ�h�̀�Z4�;���{�&��7%Cc���7�B-����f�J�DX�T�a��3W��	���[ܜ�s��2�?��C Zc�/�sM˓����V/�z�C�i������,޸��"/�[)d}n[q������=�('�2R�FH�_K#����a ]%Sp�1�U6V�����Xx:_;J��[�k�+���&�cy�:��ziO.+_�d��GcT��˓1��RG��S9���%�@�ǖTT�p\�ako-48|�o4�[)Tg�?u{� ����~�μ���OP�Wa������f345��<���o#�45���.)���|J��e�Y�}�L=Y�|=�a@�;"�2����冻y�FՑ::$�I����=w���71�+���qg��U��_l��v.��#�&*P�Sb���+6������4���:B�_|y�`N��?dy�cP	ռ��F��Ĺs2��6J��gC�_�/U,�+��(Q�n]��8߿��BH�X���U�ʄ��{���A�Ӿ�\Q��Q���Ը�����Uw��20��b��.����6����[+?�`z��N7�)� �kC���\�7c$g��N��5z��� q!��5;����4�t������ψ(�I�n�r)m���#ֵ�Y�q {A�<`�X�/}��1���d�
�B�GJoM�K��w�UP?�¬��R�kLkz	����|�I� G�f/�R�I����vZ�0+&���!3Y`����f��?N4,�Mg_=�~�.1��2��:[L�w�5J��F
�L�=>,}�A��Ϲ�ؤ�8�"�y8?w�r��L~�ַ���r�o�Q�IW\-<_�)lq�~Af��P\��0Q�ǃ�V�$~f��3���.ߑ��3�'�T�;t�E���x������<�u�l�|�Tm�iPi�)#��tBH�w�s鲇��#��Sh�DŘr�/z�=ʟ8 ��㴄
ՌԋS>��V��ti�rZݞglfN���U~�jH���]������v��)�����qB[R޻���G:��v��86����u�$�!�L�Y�5�bߢ�duD+�>�p�za~�p�i.$g��VK�����'��8wW�|Q�0�L�	FD5�\�L,TP��$g�H��h�s��Z0���(gm3|��:&��"Z��x0�a�򴀴F2�`���U����b��\�
�fCcw��7` q�b'xR�Mߘ~ߝn�.�ܱ���i5���X1gS��H��������~ ��v2�����pq0��#>�t��z=<�h�eg�RHʪu!���f�mΓ�O�5鑟${�Q�H����@s�F�%�\��Un��?-�������H�'I �J���H�� �N��yj�E^5�8�42e!�����[c�׍쳙tг]q�6I�S���_O3�I�T"�	gX{\�t/�*/]������D�:�"���y�y[�}�ǗW��u6b�;7ad�\�Q���_��7�����r�I�`m���q�^Gd����v9�OO j2�@��O����a���+3���x��1�R+@=�x3l�6Q�-�imJ6K��Mf<}��u�%�t4�"4�G�p�C�b� �⤕��6�L���6"�/?���C"!5Ȟ �}��v����)�0����An�AiX}�2�v���1�Olp�(0����mBA�F�u�꛸�4?�bjd�?ڏů���E�sK[� x8)���03T�	j `�{�a��`J�wg6���E<am�(~�l^�|kk���qY�J�᱃sG��1刷���:��Q���i��k�k�4Iqm�u�f�7�0�I@������&���,��{TLvvx�\�p�=��`�%k�އ١XP0��d�l��ؘ}6�-/�ۙ�$ܨ�oֻ`m�x�I�0�3$���.�X�Y��C[��׻l�)N��	�-1�u+�� ��6��Ix@�+��a�=���?��&W���v 5R���Cx ��l	��|�,�rh�l��#0^����q�E
��R��oF����<��c�>ʞZ��ѐ���k0�� 굔�~�yru��0�1�t���sa5�ǿӮ=M�j�h.������T=�>�����fe�{B�U��+���1�J���ݸs�#C����6:^�5�i��%�ti��gD^(;s��z�֑?�+�!}��9-rF&P�v�i� Ǯ�3�YQ�j�9�%���F���^V�����!���g�|����p0��&�!�kˀ��%-�s����y{H�x|@�j=��~��h���6?TИl����i;�x������.��H��B��g����1�c]�iU�]�6�;W�k�KC�,�}r;����.�^�b��>�<?@V��\�7"�V�5�|h���怴�b��`d1��1�#j���1��2�[�h�`� 	[]G�ҮS���~�݉!DV$�����RJ���b�a�'�"��nz��A��4V.�1u�=qiЦ��75�8C:�>�4/;�*�18�Sߵ-�b����'���}#��娠K^�ŝR�ב�wm���?T?��?nev�#�qT2wz���*��G*�����^0H�fT��	5gn:�G;�3��$��nֺ��e&����X�0���A�5.'�U-�g�[t�/E^��eޡ5NU~�)y�-��;�$����\�K\�/w?�6��j��� 4w��
��F���lnBX���4�_��_�ԓ��g���Ӵ�&H�lN���x���&�ٳ*h2X�M��
����xX��H��Q�]f�oj�6O/�_YB�4A��tޘi��b���q�	������ˤo�x����b�~�Kŵ%s]�V���r����6�_߫�����tjG�Z�y��L��U��pJ(Bwې�de)�b` gZ #�����!�3����@u=�ż�����l��R��	�iZ��v�k�ʭ�[6�X�3�8LJ.��T=�E��ڼ���l��aR�P+�08�|��*x�(���,9%��R��:<<!�8a�z��{or�)��L^6 Ri��/�~J��|j��O���)��6��Se���y��?���O�)jGe�{=������C�5�^��`)�%O�����1]Xn�&V�{\�w�H�h�锣f/��T�H/s�.�v
B�O���XL����Ֆ����6���i�)R��=S%,�@ק��!�D�EM%�d���d�0�i[ͷy!?�����1�;2���I �-ܧ4�+��ƖK����0$!#MF �^H��6U��4ɬ-�k�۰�D��.�)f��b�4�0^Ã�A~����7��L;|&ҁw7e�^����1��_�\ZٙR%딉<��X�\:إ�����UQ�kB�`���X�xh����]�v��a��u�`,�[m�$x0u "#<�Ƴa�',Y��>��Rsc<+�p��M���tx7>�0�9�su�p�m[�l�YYz�f�t�����6y�"u| K R)�վMba\[N��d�<�CA>_��+�B������c��(Q�l�C���),~ h����� sK��H���*{�U�-�>L��C(q:MK.ڜ=iUl�]a��po�ʐp�)w�0�:Q�cdR��o~)q�\�q�$����z��`Y�Sk����Ͱ�Cs�>�8�P��Wvv�8M SKCL-�Ix%��>夢ɪ��+�����x�����mE�Z�B�B�JBAZF4D�Eg6�U�7c��Xf�<G�Ka]�6+��JF��(��ݵ$�3��� /��܎���RY[���?]]?�����N�x�HL׶r'�0ۏEx�Ҟ����AC�&�[����R	T�#Tp`y���+%b��!�����k�쎁�VP3�X���=�E��������)�Z�[����`�
<Ȼ��.�yX��S������xw��ެ)��6���^���{�]����j"��Ej�� ��D��o�o��Go����Q$�2�6b1+kR]�g_���)�8a<��A' �5�Ov�؝`d�v��6p�������Ǒ�,s[ɠm	��cr|̮�wh���W���P&Ĉ�k��"�ׅ��y	п����J�J`��t����qH��t&��8g�3�V�	JK7�Ȼ�p������M]�㹌�B�/�I�[���9m]A��N�Z�GS��h�i���DĶV��&	v�+�<�vDO�4�k��)��MO�wD�7�S�#�>�Z�#����꒓��DQ}��� ��3��H�ϛ#�5	��(áa��mE*_�
\N}��bO��d��b�1ł��z�a�W^���ֆ������;B1h�S��b��J��A*�o��:�1n��VZ����.=(�7��;���~�uУ�K
>=F�j���z��$�P���F閜+��{�
��?۵~ق ������N�c=�_N�= ��
�1�Lm��+k/ TW^��,$��z���V½�P��R�݃P����i��A@3��w�2`�w��~����=���)!n�s~"�EYͱ��Bc��Bڀ�f�
�����8nr?jJ�F�n�C(\��#l���Kv[�䲫�=CL�8(���W�[�nڒz��i[�6��^K�L�3Ql����������<vO�s� }0�@�-4]A&����G�ecn��b�Mk�+0Q����P��5"�������WT�-�֞B����F����c��9�61`���0���ǈ�"-�H*�΋m��>�1
{���#8���Q����Wy8h�bh9�����Nvrtu�-�E���?Tqe&�h�Ձ�hO���ՔJ��|k%�h�*}	���ɲ���L�V]��_^߼h�p�WD��2���"Y IZ�3hY�����H<���Ph�-`�7hUs��lS�)�M�Lrn8��6�^��F��qa ���z���*'��|��L	vheZ4eJF����3;B�eMnR�J�~�çVY��-&Q@�Q���W�F�Xr���:0���XF��it�}�^G|�B���0E,;�Y����.���:�*�ohG�|WS�4E����^�r>���(G�t�����+$��.{u+a���o�-A 3	O��nj��L�󏉢,�2x���R�BTc��2�l��� �_�oc���y��Tz�l�%��+�/m7���v ��F
�&��d�8g#=�`^�L��tR��ߒ$�T��#3�"�d2v/�v]��"���D�@��� ^Om��H�޻�biH�0�ޝ��S{`9~{�0���Q��`\�T�L^�Ӵ�sC����`XǱz�sD0j{�a y��� ̖$\!�������C:�Q@��RZ?;Z·��j~�P�0"��9rR�Cʭ�Tgh�ׅ�!:@��"��C���;�xX��Z���B u�{�[�N]��k���i����ش5�m_�ڄG����Z�09�I^�mג���/����m���#Q�GVb��m/NyT�e1V��ٝV���ΌVp�?D�F������퀧�7?օ3�)�v�z�r%*��2����
��+&���b��|�=_d�(�*��ȸ �/���^h��	�3\vhԴGvM�k����r��}��|<�#��(19>c�F���Ra)�(���8��t���k)2���?�ς�'aC����'i�I	�7���H�Ȁ�)���n��"���)Kq��FGY�W�#iM��{0>�ؚ2f?q�Q7�u����S�X���Qu��/�麇���jY[�f����*�� ����~�"��=����!2g�PrR(S��:���_����o��مi,����2G���>/#�tI�A~���ֱ��y��ǣ`-�iF�-�s��1&�C�#�9��g�&�)�-+�wb[ϸ�f]� wv��(��0��?������0ȯ���,��u�z+�MĖ��s�N�Օ>7������;��� �j�
�,{�R�ۃ}��z��R��4���Gǆ ��6#�+��)��.�������|xyh;�����ЂH�@������k�ť�i0!a��x�}O[V�~�3����\�^U���s�qh��e5��t�^�?ٳʣ@���Ϊ᳥z����*Au|(Wfɵ,�+8��`yv��br��W�	�۔+5�u��z蓻J�%�F�lz�m������X�'w��LM�:n�T�-���x��h�̚qJ̸9��h��E�c������_ڤlFKb�NbOo�p�o�(֙��nB
����Jlc�����ǌ�c�9��)��������>N��i,B�����N�+Ϫ��#�CXj��R ����@pBi帓���Ī"*+eh(|P��aI��jq�1~��0Ѵ���Z�GS�[��|Q>��W�Oi`p*Z�z�|?,k��	C��d�����<M?N���F�ј<�1�pwx������~�иz��2h��n��$��#���f8��\�yx99&z�K��t!�e=Si��_������1��n��ӏmy)��t[~���JX$��@�b�.}4l��`�y=��i�9J�����G�.4g$<xJ�EaU���Ac$m�iS �Nk���]� ���W�;� �&3�P�M��y7
��P���ߞԓn�9�+�������rv�H$�?o1ź�
N���/��+g!�t�^�Ӗ�j�?����ߢQa򺆅�t#H�����y�2xE!ӻ�M%%J�GXf��q�	$�V�6<��d���ĉdޠ�(֙پZ��}j7�Y%,4�`2��MFwm%��`b3��<M{%qn^�*�AM(���xS	ɦ� M����գ��ü6Ϩ�������������H���yA|�j��^��Z�f���K!$:ي�c��40oܞST("&r����+�ӜL��07�4�w�_�x���\G+L��*^�"�&�Z�z���-���)��hs�n2���jO�[t����Q׬$����_u��F�WzG�+~�y㰙4tȐǋ��#�����*wL���3�c�Y	���R���{x����<��zJY2�d�:��r�Pс�U�j�%uX�f�Ӈs
�eR�Q�l�������Z�u�j�� B�s�k4$�ͺ�N�0]��U!�f����#7݈�,��7*L
����V�����f�L�*KP� N/���&�<�)��%�Ly�[�/A?�X�� L΄!ϱ�C.C#j�d�ܷM4)�x�1μl��R�B2?ư<�E`����j�Yc[��{��R)!L� �4�
�\�x֭,�)W]ȏτ�3��6���;�R l�qey��߽"B�u��٧��kP����QdB���d}ju�H^�	��W��E����}�=i1J"a8U�q��]�~9&�YË7̾-��2I?~��nX�*Ń ��?��韘ד|��26'�&�)>�60�E^c7�3 Z,�ܐ��K�&�E\8��P�A��υ���$}1Х�W|C��j��I���f���=	#F��pז��b�>���/\��#���*	0�_7E{M���G<�dS �2Ĺ���|�~�ƃ���*�~��<�H9loe��S4��&r��T��r�����7ʃqos���6s�Фa�����\̮��9��4�a��(@^�����M��yn�ys���K���L�"�C�����_��Z�@1�޿' %�i��}b�IU��*�#���K�ݑ;�%,Ӡ�<d��x4���hO�'����:w����T�f��_��d�)�UU�]V��'�2
e��5�������#<*��I%~�j�A��$�a����������T���Y2�H�����kTw) w��_���̵�a<h�ծ�ƴ�4�j�(�@u����KC�|N/"o]	B��))���7Kԁ����T�c#f��V��P�7�b ��F�>�x�#?_TF�)��<��������w2���l���eJh;�w��1"�0׿�))��~e��[g�81�.�+P�`�}P�3����T;kC�dO�)��H�,���h��p8�B�I9w����
/�Hz l��V~�V)]�}�(��!<��������,�}'���9�g�T���^��ls���#p��t)��F�AN�_3@�l�~G����*����byt�""�PM�rD}�1N!ӉK�$D��豋crW��r��-pY[l<�ufT����/W�
�c��PQXiVrϞ�I���+}�]aT�#&2�qd?yB M��
�Z��3��H[!����	�p��w��vk���}~�M=h��w�o��N/�%����	�р5�ð���Zqہ��,Ba�(2nw�-Gl)t�S�"^���[)*�_^),��t>�����)����s|�>�/~�|������[yy��XX�z�w��w�8>���f���7��X!q^/������d4BX�L��3�w�a�Qö��q
'{��+�����b�.�ns�4tKqc�M��L/�0�4J��!u��Z@ԑ�y�������������?�4*�Lܜ�4�B�
�p�z��)ǟ|���:�(NyP;ɳZU�� R�	��Fc`�g&'eo�e�OO��t�7�nps����p�W��r�0"��0m35�i9+L�Ē2֗�ڠ�K��+��W9�>�>���ޑ�i�qLU}T�.Q���˧�V�uhqU���a��k���H�n�i�ug{�p���&��@��;��[e�7�����7�܀Pd�=["�V�h�� t��9F���\���|_�����'�S����£	n�5����3h��!S�K�%��ք�쥍�E!j|�cc�(� ��D��"A&胺����KR���~ �+r˻�����z��k$��������d�~?Y�1?DCۭd �`^� K�4]7�,���Wg�F�m�]@Õe��^���]��S��e�~\�$Fknݵb��:_�i{a(p�H��r�q6�N������lf�o0��Js�UUY�r��Q�0�S�ƅ��~<!��!>��>w�5���NFiUeXx���Q@���bL���ۇ����eP�.��g�s��u�f���!æ�Uh��q좱*�S¼�����Y�h�$ӗ��HNntL�Wa�LKj2=�r�K���p �#��^O�RZ��r��-�� �0'W����x���5\�=����0#��Db�S���J���v�U������<���d�`�D)пH˪Y~��1��/�<JЧ�ZT�;���"�i��׼R���+Z�|UǞ�E3��/	h+!V�ګ�I�\�;V�AG!p���i��1-G��=�:ϟ�/�}'�dQ&�����-�J����3Th�0\����� V#��p�,	��xk𾉏�Rpӹ"4�m������n��,�/���W�Xa�|�v�����*�����R�hce���W��E�S�v߰Z��]%�@B�Xch�&�3>�Ƞ�0Y}����7�k�S�<׾C�
&�v�ևMzjm�ǃ7!o��7]�e���Qx:���]u�
JT�ƚ�r

ʶ�C�\ry�����s���*������_�d��>�|����J�&�������`I5f��,-��ͳ�����y����72�6���1�wo@��O6rp�[k�f蛦�N�,٢�.�� �O�h��;�(<��D�K}.��h�F�@�28w��Q@a��NAQ7�����}��`�e�	�2�fU�'+)=|~��W���p��?l7�^�4{u���vT��i�ca�PS�y���|�|涆8s����J�j�3�Q	�,�J��,Q�K�۾��Xiz�g��IL4�kfSSH�]������f5�4�e�
ftv�~�7�T,��e)����[�kԭ���-ȍ�:&	{��qW�+��=�E����t���La�a�W����u��S�Б_�A���C�����#V�
b��µ��,�r� ֻ��;4���O��n� �WJ� ��� �6��[SP��Si����u���q������{��5/��i��{*R��?w~TֵT���Y]S�n��%��96�2T8��6��_8؂�P�?��k"����X�9��|����|d�ewc�@��]��Nk�̃��myUwp�`i!�]���PwC�%���y�E��s�*��8@+N����p����۟��X�Z ��1P�9�<��-/��'����" #�h[��]�g���L~��r������p ��^�2�_
��\W�B��5��<�kj_�pNϒ�
W���3/I[�+�	u_+|p�R��C��8m��p����X�<�E�%"����3v���9Y(T0�m@��&Ց����퍏�}���K��֒���z��Z�F�د7?�D0.�K4�.��S�^�y�H�姡A؋���]:��7W�����j�T�ۑP�$B���tK�� ��>Ӓ	��6�k +!�$���u`p�Zv��-@�0���㈫V�ް�^��o��¡�-���ͮ�v�� �#6�h7f���I:�Q� ��ς4��x�ؘ7���R"^�(��3R�u���AǍ��������wO� I�6$0&��.C��\%.K�<iܞ�&���&��[k�o7��a
�w�xV�}��!��p���5���=��+�KzIc�-� _t�M�o���dbm���f"�աs������3��H0���	���������c�?�8�1����)淒]Å
m|�X�X�2��#�9||��9��9R2�OD92P��Fʒo�0��rZ�h����%���}�6Rh�TRsοe����Ѓ\���tZ���cО	���:�U��A	+�^�@��M-�\�-�V߾y���r��!BwK]}:L9z����4�M*����,S8�Xu������w�|�����d��;S��h�JTPx:u�d7�i� ��|WޜG�2���;?��#�oȏ�7c���nk-i8W���e��3|�)<8�LutՃ�����&n�%@�PӴ�Huۻ�A��4V���V%�1�6���!�'���G2��9B�cp�M� ��F2Y=y≯×U�H��ڊ�X>���=�%�y�)���o���W$c�K�Z��QF�Ə?��op����5�%�)	�/_�L��<?���W uw�#Zt�F�a;Bl ��&���!KV�.���9ë>/!�é�
:$�e9�p�b_���ѫ����q���M���4����X�nY�1`;��c*�?hkE�r��ǜ
�fG>����0vFf�=f)��̒*���ӽ��=�7*�E�.I���3<a�<�
�,׾'���y��^����4o���פ��C��-��Y�,����?3^Js�6j$2�>������8���U��8*���d���XS���ʞd_�S��,EV��o�p2k�� �������>��v�{��-`Z�cI[��;�L��E��PE`�,��$#��G� ���Jo��d�s22|��&��*W�cP-<������>`ԩ����HZ��[�{�V�':>Y9�U��������H������"�h�h�^����5e��w�C?J\b���
 �e����z0�3��D..��Y�!NLr@	����B�6���S!_ ��w�� ���1���l��k]�#�	��,��7�ܸ.�q��9�N���m��ڮ��ݓ�%�/]WVq���RP?ݴ���jP����5z�#/�αr{�(��/���T�Q��`B�����U�^�L�
��X3�}����(�da��?�C|�kq
�s:���U�dxE��B�2D��_o?�<�m��g���Q(�J%�w�X,��t��RD-���\l���v+��ezh��5f :���8u]ڄ�4��L�kc}�M�\t� q [O�� �ATR�C
�jz���m;��Q�\Fo)\��1�F���s،��}y�0X�hT�	���\���]`9jQ蔱%:�`W���0p|l�]0�U?H�N�������X� 2Զ|�nn��>C��O�B�Z���鿴�
Ԕ�nѺXLv0<�ꕨ,�>x<}w;�tue�x9)fM$etn��BA3�L�	-����ݔ��r<�Sk�4�������i�|��Zm�3�~���*�fԦ�h��C?R��af���)]�׍xU[dюH��w]/�hA�;��t�ԣC��o D�l1B��v,�M���P�J�W|>F�ck-�j��a7�b:���שP���?[�Y���n�����Q$j8��{RO�[,r<`�VgZ���%/�;J�.弴q��NC�դ�_��װ��� $�e\���ۅ�S���B�(���r bz���훢0A���b�^GF9M	�.�w�Ue����{�9��j���$:~:T
ث�9H��;86�R���k���w��8��Ѐ�����:�
ͬOFk�L�=bhţƁ�����)-v��[-�
�l����`I������t��W��y$H�fMs�x��K}���
�{\hc�=0��C_j��qh+���Q�p|�nB�/�/k��j��4�$F����D�l�r`�,�F����fe0^��\ZD��['j,��k�M�l��g`P�5'���l	��X���U�a��Ă(l�R�Ю��"$�L�K�v��9�I
�6:B8������ޯ��U�d��t��i����A�g�ג���[�� ���ݹ,������]��` �o}��S�%������lf�X=������t�2Fϩ߷»�mӃnˮ�Bˈ{N#��H��d��!�q&&�Ν�&�1L�.F������S�t�p�0�:\����;*5��yGX*�]�i�h5Q��e�Va�� ;�L0Kj
�����;�U��!��j$�*�u�b*��C ����V[{R�0�6I��,�W�`1iI{JA)�XK�s�����d��u��[��I2:eE(�ᠶc�,M�����+���$��hw�[ic)j�*ůl4��m���-0?�+r�;dݩ����E�AT��h�f���,��!��"`��@{��#��]��y
X�����������	2��Q��Z��\�P��_jL52W�n]NN�t�ݫ�j07i��J&�/ vG��< b��l�BK�W�	�%qħ!�D�'8]������fi^�<��L?���C�1ٓ {Ui���<�=x����ڌ�?c�톉��M{P�^k��q�W��N�B�]>�9�餵&���Xb�yhM��O������Ц	�`��j�9B�DVoz/�F�Ԙ�1D�W��.K\޾���JT�7����?�w��X�:�e�u������t�
x�m�ٻ-,ہƭ�V�@nm��	Uٷ�M�B�9b �`���Ii�E5���B!��<�z�}��� B�yD1��I��h�N�'�̯�l
8*���g�+����y�����%�k�]e
)A�֧������P���{O��9��U\��;�Ϭq��ZL�#!j#1��<a�/YU]7
ؖ=]T����OD`�%����t�#�Rc6MbdKH4�j�]�ҧ!�u��z�y���j�2L�ӳ�2o[7���Ud�1�Hh��۔]/'�Ρx��J�m`.g.8e<j��$[�- p)��.�(ɇ�{z���
�:�4�}��1�����;�@�9+�
�ՈP24�����U�Im[���8�7�`�Q��dedKC��C9�Y[ 	����w����UQ��w������K�1��l�k,���M�Y�e,:����@�L�Bm#�����^�O�=��*v��_�ر�;��tu����O�[�J[Z+��B �F�_���4����j������6�ڵ�fg-�OրK��X�@�ɏ���ђ���MG%�3~i� ��Zَ�E�x3P4�Q�8�?R�0�G�>(����|}�d�9����)����\��_��d:�oV��y�zp�l� �+ѭ�a��7��f5���	�=ؔ:�?�k�T�^Mb¡���/"k��ĹhN��
CKqN�}#'�s�WH��IiCƥ��S�p!�>zMt(��V�?��I��)͘�Ž�����+����� �>���anyD7=�n��N%��'���x��N)�#0Q�&άb���N���{cI�mQ=�Dwcȱ�{G��-)C�|x�_�^��������\/;�����^GU����pZ(�c�cu�,a���k���р�JG��<�UB��ݼ��}�� ,�,�z�mr�h߽uG�*�󛇄�3p����t|?�_���ڋ��b��JC�S@Gr4|^��g�Z�Q��b�}���s��'�>�p����\��t�l��>#���%�'p<p�J�鳕��1�H��������>�:���v�e5$8�֣�6fH�� ��ۉ� ���`Jٳ�T����v�Y����!�C���l�+��vN;29_�����%{a�sGd�E�7���j�cO�w��&B���c�>����mS�⻵!^L�]���K��>�w�tG5��I����ᴥJ��^u�d���[.��/j�/���Q��r�9{-3 ��"�b����W�\�&��eh��z@�D���i�y�%��Ė��g�c;�:)�,�*�u	���_������BB���Q�}����2{d�I�@�)�p�~�Bcw�W[�u�q|���xZ����-�^L|~whwϥ�f��ÈJ���L�� Ig%*4�\=��n���&;9���B�C�g�����"xｘɄ���f@V�/��Q3�����f�!��c�\HȚتI��C���h����sj��|��?@��\�d��F-%J4��'$�DIk��:r��z�w��޾�B[媤p˰��a�H.qC�P�C_z��p7�0?���⸄
�Q���I~h�������۽2�0k��%�5A�a�:~�(;,D���G���;Sq	]�}���Uk��,�F������0@�N_� s������zY��Q�e�4+`\�wMHj$��ۊ��r��G3A�,�D����'8;`���Dݦ>d �<9) �B�Ly��͜ě�4�h��o�EJ��W���N&
ÏqhhA� ]Z���M�»ہ�����W1�jؒ�$�.ce�QXp1���Z���eh��/�ڧ��������D�o�8��s�����w<�0,�9t�$��Z`�շ����� ��Āآc'�b���"�Jl������s�w��$�`�X.�P^�;�ZR&��:|�>��Ve��\X����6rA�e�چ7hmB�" r�w9H-���aOhG"��"��#��#���Dٵ��Kn�Fڇ���)Ԡn�Ӡ���?
�t�w\Vo)���8
-�?Çs3�w��鯄��|�U�]c,S>�C�ߕM�=���-���`�ƅ�@�%�A �����{�,�>��{ ��>[��cQH�*{��#���(���5/���C�	���4��a�GYt�Tx0\G�5��s1��ձo��%��?8'��Us�g������CZ��^���J3��e3���T���Hy�P�/f1�;� ���O��CyD�Z1gGR�l�q���;zl�ݮ��]���@�r7�����$r����4� �'2cB�dۙ͹�q�
TA-�A���ؘ�p~ӽ#����x�y�j��u��<�(j5�kX�(		Xo�k��qU�Z\���g��LNoz�_�3Rޤȃ��-������
}��T��h�6��f�~M��i=r�K����y�B�(m��#�(rp�z������;��Ĩ�y�(��9����O -��Dƍ&�+TuS+wQ>7�.�O���� X\Z3o^����l_�����3Ġ"��<Zc��64�,5�w���@\�᯷�_�6'����q��� Ppk�H�.<�^ĹO�ࢪ�u�����s"z���;Z� PoZD��X����ŋ�V����"�L�\�Qf����%p������{�{�h�j� �ߔ��(�a������r�JE��T���Ry���(4��AU� ~@d��l���!��2�;Y�z����{X��NM���xo���-ył�ߵ8������W������Ž��hɎ�
M���{��v�(Z�N]��D~�E�	�/r��S��/�D�s�J@�D&��֚{�g�J�<��{��S�n+u�$��/�V l���H[Ԑ����g�^p�C{�ꁘ	�!����#~ųy3���0C3�Q0��?���I���=A����#rC�l{��I(�к�%�+i��O�͙��`�:��r��R~�����)#��J�y�.�zs=��c��x�=��{ ����W�b�zc�Ɛ��ピ�T�f���O~�����% ��@o���!W�&��Tu�rm���ݿ
�<.�q��Sy�����ta?\x��/ߤ�D���[~��̛dÒ�D� ��8K�-���t<���lf7��1�?��䪞�ɺ�;�P]�i����!X3@8[K/n��0�Ϡ�ݠ�^Q��n��"I$���g+�ř|���34�p��Y;dpG�!���n�
v�o<*ɯK�Q����a����~��>�<z�%l?LM|OU9��i73t5߼�%}��P�<���v�0�,a��o�9��,0�wI0�^�*4��=��#Z�@P���ߺ�׸��KTݨf��CE�����.h�$VQ��h�� �땫��o���	k+�ȐvN�I-�	~�qA��Ti�FQZ�3�=㍖\�H�E+��X��
�p��������7�j���H)� ��q-�Z2�jX(��e�M��0�@���֝{Z�x����V�.�$���6��3�ٖ����#�H���B�PV7�c �ty,�
��{�bY�5�sD8���%���ұ�ő�2�wR��ߖ�֧`�Z9@ɭ�����8��ע".�6B֨"Fn�B0��vw9Z(t����-�Β����G ��s��D]1G\�W�@�q�O��Mq�p��D˞2�e^�����F��	�<#�S�co�i��♖<!!n��Z��� ��Kc��WB�n$��#yô�`���X09�_���j�s�G���+�f��s�.g�5W��I��(���t�;o=O�|�Ĝ'	���Z���g~L$U"oK	BՏ	�b]?s�k�ؾ��q���Vބ�n0D���=88�Bf�Ɇ\1b������Ա�r��ά`x3$���:�'�d˳`V4V���%���c]�?rmWJ2S~�ϸ����YT ��g�V(��x�ކqlζ��T�+0n�jR��j���b�����(ֈ�Ç̡����hz����A�E-��tXx�]�-�B�HG�����<��
��j�f�V�p~���8
�#������3�nԫ��_ɠ�w ���
�x�ejh����+y+�b �O��$�3N�1:�wc�焞��={kq�7�F��!�3L�*4L�sȖ1���%�#t��� ��Nuf~cx:����NN�z���GN(��O��o�?�l���]%��嵵C��� 8|��C���_<ީ�9�^H��5|c>�G�E#�Τ��,�r�:��9y�V9H��a!�M�#֪�G�Z-��:����o:��K�ў�+*��p�fb8`t[�Je�� �����;�d4��;t���4sD6�ٟ�h<��{&�ҕnң�u{�{1�W�|�01�!o�g���68N0M�t���ns3� @Z��e�As��o������/"C޲Uw��hnZ�}{CÝz@�!�z���}i�-��>C��ӏ��)����<v���?!	��`;��>���w����r��W�@��2V[a�|[a�E��\H�}T	~X2�k�C�9J��ğ�]uZ0D�OS�}Hy��Ʋr��P���!���i`I����B�i7]!a��U	����H_>��[�9�1��\O�t^���b)I���1�T̥Xf6b&�l���9͵9���2��SAjd���7=_p������<�h �"I,��!�-�a��/'ՙ���C&cgA;��oox����z�-P�D�o[7%H�F��26����t�G��p��2�rW�i���?�(�0>� ���+mM7�v�h���E�/u�Ʃj��<i�Ei���pݝ?8YF|SG8�3̊A�M��ث���ì�[�x3����<�^�N'�,�VE�YcU[�n��͐��!�K�$��ǅ��52L�9\!���7hfIhadŦhH+��h����f�2u+�Hp7G�oY�-
p�x%Јj���U�e����:�75}:�t�4�������Qic$�WPA�>D�K�7�n�7�}'h0�H����ԣ�!"��+��R-]���������L����V���?f���� k��1]�ʍ�،�� �@����s�,�����s��WC�|�[dREᏼ�1�P��>�dAP<�^�t����vv_8ȏh����9*MK���9�~�VmS��������;L������EH�UG��62Z�D��?�|���������P��o�9'@����?�cB��qB�a��Uv�����_��f�R���U)Ytƹs�q���TW0���=�mK&L��u�grsS~4!��;x���}pؒ 
3ڽ��� kͶ�ju�����T�����B�Li뉀��������mG�N*X�DIb�a�p�� 	S�k��"��,���W��<�p�Cl�䵀�=��4L� 1�Ҕ��#ɲ%�'� � ���C\���PI��.��t������g�ل���ΒT�u�	bB(��fzۂI�лuZ>n�j�����#�� ���XA'���DҐ~^n��~1	���z]۞�e������5�ti9 9��BZ���@tJ՝0��ȹA�aU�VOd�������Oo�?�ʿ�R��M��v������ڏ{������4�ݞ���"���!�(��V%9\ϊ�s��c��D�0�����U�O
��TƤ#��D5͚ɭE��NoY���*�d����Ǜ<.�Z��_�*~C��)�ӡy���?QO�Ke��+C��0U�N�ݣ扌�H�8+��=AE�"#w�L_yȢ���UY���T�X�H��#�����e/A�(4d���fVj�HW���ĭ�[~�����c��Cj��5/�J!�V�/W(��1�آ?�F��C� xm�",�	�Z'!�U�}�
a�`v�3�b�~n�y�2b\{�U�H�`��|x��x��-�c�N_��8���I9Bp��-f�E<o����ͯd):�iۇ��IX���y$M��N����|YC-�#��j���Z����K���icH1~���)4[��Z2���[\��y�����x�Q�}A�&���u3dbp�VT�S�&��րB�݊"i9B�r���C���P����e�YNӌNU�"Iަ3y4�]���Y:�D�� d����r"�w�WK7�`�|��/�����d]=�Z[���2�w�A��4��L�	��cGz���i㰕d?�jI1����G�)"E��綻�~R�f�[A��'L�y�8[�	����YA��"��9�Ȁ�)O6c��ʣR܆Ȯ#����z���@a����"�K������*���c�V|���8�L����b5�'�m�4�xo��B�C�f�sB}�靱҄?�y�xU �B�F�a���3~qB���)��5��($��d���,D�!��r�N8�ڪ9Mn�O��CaB4vy�Npğ¨p��=alK�2/e�����9�fl�>='%@U^���Q���ș/R�w�G��7���pz�b���t�ޝ��5*��ž�U�̠�2����6��3H��%�F�Tp��n��}�t[.�T<�Q.�Ƞ�	�3�'JZ]�Y���13(�(�{��E���D�A��]C}̭j�KxA3��Q�g�|�s��3im+�������ܗ8��9zdU��Pf�Ԏ�Q�3W�8x6�Z��(P(�U}��V/Q�)���
�ri�N���]����E��4��_�m* �14�~&��3��f�]��JA��(���׈�³��"j.��3~��k�wp;qS��k}��h��j�U��V��.�'�"�5wX��cYР^q�l�!*Ϥ��{a��M}��,I�|��j���jv:c_��0-��~��O��"�v1���F@���x�!y\jq��5X,J����v�ݖ��aN&~UWe�띛ߦX�zP C?M�ݱ�,8��)�Q�sG"�Z�u�+hK9�i�SWhX� ���?�{��)(���q��Ú8��\��6�}��u(�Euh��[?7gn�s�#�4�V\aV�0�r�X�lM�g�1<a��~�K7�\���j���v����2ٗw8'f���m4?G�Ewɿ�M������Y�2,{�<���?�t�+��J�rk��1.�,lʠ�J��t./ȡ��m��]�"���[s�#����f�b(��:��kI�}���:@����H��!��@��R�]�C륊
Y9���=��oMSJ�+��	;
m)�.�n���ҟ
b/� yZ?��ff>���>^^��qlOa���K��>�������˜$;QF���NK��LAP��PJ��Z���܋��7�͜A����q(7D�Ѱ�h��o���ɜ,�OM�"Ht�,�O˜�����;�~�֫��"`d�WVRZgJ׿�#�20]�t�ZOzP2�4a��$�枓��M�i".Z��l�x��Y8��>�FC4_{w�H�u	�-�[	l?�-�(�����䣱)tgtHx��-�I\�c��6
�aT�3[�E8��2�b-{�d�G�̞
u�o�[m�YWғ$�w`2�/���iߌ���vZ-��zȞ�w'�#6>e�i!!�F�bRݱ:2P.nh9��v؜Įcea��B�V6��Ԧ�:��܋
niW;(��olG��;��81(^��:&��,REf��0� �01�?��z��Q	#y{wg!|Z�g�Y��P5�Gf����I�$cŘ~ܳf����	�����K�S��ma��y:�O6Q����M�/����\�I�����v&�c�-����4Д�K%�Z�����ei~��<sH��O&\�:��@�KpLF!W��P�y4���A_�f����5�K���`/[��1O���`��L�4�R_��M���������+��	֏��Q��n�"�\?Cѱ��L%��}����*A7)Аd;�{PY/E�Y(�2p;_C�̢{P-�a�Y����j���ȕ��i]�� q� \�d������Q5]͢�5���D��Ua/6@�R�i P�u�W��`sK���wo%�G�'��[�f�5�ΑS�a	���ґ@cb�|��NXf�p<I����ǰ�b�X叩�X�9���݀��F*�:�I8U�xT��@T�����ʱ���u8l��.dH��s�!qb�>9�S,����V�<�! ^'�Vk��������P �����Y{A�
��t!v0��X"Y��� FW#����*Ԕ�K�I�-��F�n�/��LN���H�Dק�Ϫ�+���;�'Y�v����-҉ �c`�����8��7K�U��-�����	Qm����P�����՞�:ɷ������|�$�"��v:�Q�3w��{i�
+���B7��`����U��@E��A�-1�#;�(q��f�4��g	SG;!�Qj��jL-�`�s���dM�xjRz���MW<d���[_���#�wq��y�YOe�ݪ
�PR����Z+����=����2���2�����뮚B�����e�\���-���*���;X�%}��$���xz͜.�pI�N*ȶ�Y�c�5��g�X�б����.b��:Ow,���a���"�9̀�FZ[%�d���7;�����-a8�#ȹGXl���]\G�����|ssi���"�X^��`�ئ���؋�����1x����j%^�������o���K�\���[$$�p���Ö��6����ސ�$��֦뵴^��]�6 g��	l֡��W�� fh��yֆ�R��=�[g�礼`��T&4�Q�N�j�r������������M�Ubjt�@���/�^��q��/�����xG�:B�r�]/��;�?�͓�� �버z�,���n��c)F���If}&!�6����}w%��ÏH0߲N����-�0��Ȩ�&������vW8�5�#ʷ�%����
0�uJ �L����uյ���pJic{,���`5��hܦI�Y�R�q�y;t#�2��=��T�R�/!"1f[��k��>~lfP����_�&k�B9����P�j&W�������$�Էu5`ʧ�f��kX]ޒ�8�3���\/�i���V�_�_���D;��: 2��?N�J�m"k� 9;��%�����<Rx�K�<���?��DZ=nH�Lγ>c8Q/Q����"���(~�vДGkaRx�?��V
뉁�Y�K�BA�(�� `����+��}f3aZ7vu�y�(�12�b;�R�7Y� ȗ��O���t����?sB.��� �{g�CiyB�@)�ܻh�N3x������ �}�FmLG��m��	�/�����![�N<ݕّ�y�*��ʼ�M�Lt�o�<��Ogcߕh_��uwU����!�6%M��<�����o�a�G�m?7�)�x�Ļ)#�ʞ�M�-8�8�d�/�8Cv��t&�`��|��@n\hf�5���|Ax�t[��5�S_[��d�ȇ�R�������U�"��l� �/'	ğae�eh_/����P�LIK߻[D�H�;�P�`���J硺�f9у"�<�/�r�	�8{�yK���)���ȗmִB$�dSU^biFb��`�;�2���j��I23Y/[O'��xi�D�Kz��J�l��!�����gN{v�J�p�N��!���Iq�E�j�|M>_lU��h���-D�Br��
�m9W+����3}��ҼϜ
��w5�{"��;a����!'��D}#\����[&�:���U��E�9w���ޠ����^�Dt��B��I9��n=b�¬j�T��~zF�c��ql	Ն�#B�@� ��R��TkP�]k�&�0���� ���#}��47��h���k�5���R �+Uv���.�-��E,�7P��`��(Y+*$��d�B�.��)ṅ���+��1�W$d����[zP������6cp��a�7�������hwױg�	/��t�FT#��t�U:V�/:i�G#�.nȟ���Ěx�S2�E@w@h�/J�v��iԩ���V���2y~���ԅm�=FD��7�|��#x8	AX#��	hߛ\u��\EI�o�p:A��u���`�q�y@��4���M�a�+�JVm�`-X����RE
�� ��\~�\���J���G/���LmB��X���D�����X�\}B��3ʭ�H�Kz3p-��/�nut��
1X؃L�h�XÒhn���F�����"x�Y2���c�ZF��%Hz�YHh4�T.0��ΤS�r�R9��q�Ѡ���L���n�^�F�gV�lJ-ԉ���\���[�c�w�98}�t/0���GI���^�oM�c��?W��4uG>A�7���ޟ�lw����0���Ⓢü �c��"̙A����G��Yh�t4��VA����E��[�A�s�{�i'1��T��÷' ���dy�Қ~|r2Q��|{�u���l����/pJg��1�Bϓ�(���#�<�^�iRx�������.E�#1���7�gq��?n�I��.�t��1c��J7N��z��kA�$�	v�6B�Ov����|�V�e�WA5��G�+3#%�Dp��{�%��L�N�`ſp��8�]!�.���y����beä�3����0&�C�S�����.pD��L`��i{����̡�=}�����\Ec���,x��A/��ڋyK9z�y�Q�ՙ��� ᆸ�m�C�㍠dC1Μ=J%�0nwr�QC3��k 9���c��Q����v�(�yLȁZ��&�8�{j�څ�w�IR"(�4^Ϝ�<����ul�>�R�Pu>[Lħ��CK0ΚҬ�ͅM�C���y6w󭾵»���5���c��Y�tH�6r��Մ��>��>�l�
�����`%��6hJ�'�oJ��h��z��`�K����+�TG5]{#Iλc���T��m�p;O����
v�ı���s��=�2K���q?�� |�3ܫ��c4UN��	B�S�e�2��Aa&�[ڢz(�1�����\q���Zz�h�zE�w���4A�[�����-��9��&|)��\u��򥜭���i჏� #��-�|~:��m��OQ$�lL��uD[0��G3	I�蟋��E�j�W}9iaJk�>��������yA�;l�A.7c�)���'l���Ez�(�%�Qj>ȷ��G�%�Vw{u��-c����+'G�0k��'�,]a"�7-k�^ެ{�X��M���J���v!X��GI�6�~�T0���oS�čMt�����GQ��hr ��̇���\x�-)5��J���zF��)�z# ��d�cL\
��+��Gz���G�u^��i)o-�E�)�Z::=�#���#��V����N�N����j�E�8�X���+����KឡD����,�h�/�����Q�%ꈼ�o�ٗl�Kѽ��1q�Z�k�Q?[u�G�$����〾Y$m�I��| �x~l-3�&�*�ĉFbh�̀���8�TP�/��P⇯ �!�$�� .�MhUozUq��(%v�V|�Vt3+��� n�
����
Mgzb�).�%�Rs@e�]M�kDc�f��G���iC$�Q�ϝ�@#�JrC��c1v+K�5�p�2��z�}�b��v�!!O�՛5�+S��t�HF#c����Y�	OW��r��J���ξ����p��3��m�3h�b[��,�0x� $k��#RkC� ��d�^NcГ���Q	6�R�r�&�΍�ف�.T�%Ar����a������mt�]����B|�	k�5��+y좳I/Y�F��kX�����Y���1&u*&Z���d�@@?�%�t0<F�}Z��;m���A����垍Ʀlq���ϢF�����ĆH՚��-ZXzrJmx\�*>hKh��7˅�`����O�k��"f��Ă �X?$�`��a _^���߽xM��
�J�ovg�k��$e�����y��_��	@1�a��`Ԓd���9I�Eq�	�������w������F ?�?��m�q�^�|�ă'��ĺ�f��LX2���qjU34�K�������^�)6HF9Z�E�)-��b����|Q�C)[�BP�T����J�A>ճ����|�{�IԷ(��#sy�����z߱C[<�_�ϑ�pIUxMu1�[� �n1��^�ĊK2�}]�?L����i;��C��$A��_�S�Mf�wZz�jt�	��*��jp���\�;��0������ԗ��Ǻ�-]��J-��ݷ�˺<2��̀����bg`m��In#>��z/F/&��	���q%�r˙D&����b�y�dw�5��Ĵ�7�(V �z[����疙��'ʆ/�I�ϿX��d�n�p���@` ��V7s�	<{A=��+��_�T�r�3�e�`k#���W��R%�/��~�h��:)J���R��as8�{[�g��]=�4�߃��!�2�t��e�G}�!�*���wu�`?)J���a�cf��ÿ6su"Z���:_���ndr���C#'q��Jː�(�r�����5�Ҟ�Eٸ��-ϩp�O��W�bI��b�fM�b�W-P�A|��*nR�������ﻳ�W|d�d@�[����N0m����|�U�g��d��I�<4�T�6����B���#�݃l�쀸�O4$_q	�ߍU��]`�6$E\:r��y�Y8BZ���A�S�ZW��/�R�8��R{�9��hl���:�v2��w�b\P�q~���eS���n)ɺ���{{�>�g^p�_w+�R��+ϱ�8Z���fxt�N}�qƠ�'�AV�>X2�[�7�w%=�\��,&	�K������?%��+C?2*Ta3��h�g�@B���p4+�P�+��Л����� ݎ>|O����5�t��$����2�#`�X�T��� o�XW�y�������o+���
�k��h��>f����`S��䂢;}E^��<�U�.^����e�B�eI��ߘta~tv2S�Z�|F�����x,��9�(S=��? -\�=���t�"�X�]0m��2k�0b�h����2L�G��k�n\�Od�\i��jߓ}6�;��xsԎ�3�Șڡ������eB@�c3�ZPv��P8�.'`�h�y.�R�a4῭5��5:dQ�+p|8~u���ϗ�0=!��Eeׂ�A��CX&�r�#���&�%]*�p���i#HK��9[����x~�]��f��\�B��=[�r��F��� z-Ә���ٮeP�Wp�^�]q�����d�����B��F6Um�, 8SƏ����N�o{+ɦ�r�G���pLA6��_L�x�]V�!�LV5� �~� ع�Hzv{k���N� �@Ö��[>��C��'���`0O�^���Q��e��D�I�S�C�sIx��Ɂ�A�I���植�����vm��=�0���Ek|ԅ>T�G�?5��0A������ҳ��P�@g�>x�Z�}�6����®f���7�L�v}��N5$z�zw[�·���\+�ub��z}�P���W^ِ����pі�Y��Ō��j�%��3,�!��h����`)�i��F�dG��-b}��Wļ(���辰���BW���0I�>2b�CS�k#P���θ����h�8�I0�>ts_hyJ��5�eB�[
�D���}EQcX&�W�@� �2�a99���]u��I=���IO5����J����n�$��9N�\�G3�c�7�l�o'��r�ف#��������%ȅ(4ԙ����rt� ��244���Q�����uv�o?����?��0'1��ā3��(V����ֶ����ԕs�C��E)@zt4�5����>@��9{����E��n���D�p�=����t��o�v�
�"һ�zU���,O��P�{��x<Ş�D�C��,�Sl��5����M�a�����6���Y��U%ėciD��ϥ�n1��&�1�\o��N���d�l'rV�׎T�>qyd���w��O�8��N��p�a'A�V�,^�R A��nm~���-�Jw�PZ[�OUg�V�@M?t�?�����I�a��8��q�|��y=�go"�@�Zi�A��UN�V(��Hb7�4�u�O{WB���i�]s�������=>�v��ω�zF;N:#VW���y�Z:��/��K��~��)�|��u[2N�,������h�"�ݧ�W��RX�� 1�g��j/ӱV2s� a������>�a'5�Lg��
ܯc�e]!���X�RB5*�<����~�~��:�	�����ce�>뙬��:��d�6��$��F��=6=�2�)y��TO3Lэ��AN~8����3����V8�z���=�W�po�G>��+H�~t����̛���7� jAݑ�oJHbќ���#�s'���ƀ��1d:�����v<:��/F����D�v,m}Kþԉ>����|7��3 y|��"����_+`ETYms4|;��yW��-*��H�����Pm��(�2�� �0���r\�P������4r�X�dn�S�����B*�K�1��a/&)�dw4 �%���R9�T\ʿc�!x	�=��6!�7���t�1d��!�/`el[�x�E��_�(�Z7C�n�W�(f�۷$�7#��ivPY��L��g �����3B�� ��U��ҹ'�MŁ�3�v@�γoe�����v�葓���]t��im���W��cy�~SXT��X]���D�z`�˟�#�|A��d��� ���̆F2�`0�����[�\�:�=��G�k^�Z�#�f�ʄ�\��͒������C{�'�w�J ��\<�d`���խQ���z���A��t(vs���@s�2����҉!�i͑��P�_�H�s]?���-c*���]��Z��mj���:�!>�!f��� P꒏�	���h\ۗ� ��1�zG-���H�@y,�2�`I%}C����KX ��hU˵+�|�{�Oԫ�Y@U���ď6< <P����<&"��6b�՟�g�����$������yIeԗ=�ڿ棖�bؾ6�\hE'hT�'o�Kl�N $�����@�Zs��:����hb��yN�8�,�spW]�	F.>>0�թ	�;���:��f�Z/Դw7F~x�M�Z6��J�2Ν��0"�x�Ǘ�rt������U�k�	�`��̈́��'�X����3���:� w���:fi�ϸ�W�u��^0���0�cc����sC��tm�׽.����4�y�RZV]���?���8����v��3���3"����ك��T$Q���1M�V_�-�̻R?������;����N�PnpD������4�%�]��y*i��
W:}��| ��4���Նz�F\+Z5"��ր���1uEp������W�/=WB��po&L��,�����D��d��!>��hB�'`��KӍ�lD�SY��d�����V!k;�Uc|��l?Z]�c���:�@�E�5Z�e��Wo��+�ލ��ǚ[/��0l�b�U�n�B���z��4��n�Q�dj�5qp����T.,��Ҋs�Pj#�����p�:^t՝��fc������Mz��,E|$�� ��r��vHn-����$J/<q���2����������X���&��r�\6n�)ό���^}?�N����Xo�䑣��Ͷ���8�J�V"�Ah�+֟���穓d��|������x�Y�����*<�V� �0a��3�5py�g�R̎���~�!p��1l'�
Ҩ��:���6V��̔J5��BEpݺK�ʋ���j�ۜ���1.�4����D�Tp�N���,�YH�QkY3�#�6��K�Ƕ+�p�-�͖�襽�}��#bW<T(*tRHV���"��sh��6��XZ�6=!(�k�F'�/��:�:�KS�z��zZ�h�	3\���p�2W����$�I�	�tm��
���y���t�H�P�Aq-��]=+-��h<�?�4FEߨ�L����5(��`.�Z�1�Ϗ�JD��,����"��֯���K��Y��Q�[,Du��|G�f3_���Vg�O��WN{w�>ԼX�ŏ}aK,|�ڍ��4؉n? �ء`����ga�ʊ��J2+�N���e�D;�є���+��S� ������(��|~�m�����*l�Xž�v���J�m����~W]u�u}���_��'�
����w�%AD�|@c[7�����No� ���W����H׵��1~�x+>�y�2�{�auE;���]/� (5����R=�J���4rB�Q�y����3��
.)7�C��c<^�!u4W���� ��49�]IK���+ȱ�����h��U���m �L����]~���fc����8����c��6���CC�}�|�#H�ͦh`�(8z�����1v��c��f����g���oL�7�!�"�ڶӰ����Ű�3K��z��3N4�8��-twr9�mkP�ՙu��TL�/�H��~vƷԔL��3��Eӑ��fL���P�}��ɴET�?-3���l�f|�_�ᷠ<�f���������Z�ĒB�0�L�n�H�eڧ�-P�H�z���[���U�N>\D2n��E��͟uxg��PK����P샏�K�Z��LB��P�z�Y��Iu�l���bE�>d�g�a��ٜI��Sʣ����ˉ�3+����W:�B#��r}@�c�6{L��B�y����F�P�?U���3�����Q��:�,��%���|���W0��yF�؏_"�	�5�3�"b�V�V�k�h�eΈ�D�fI��uu��,�5��ذ���Dչ�I.	G���jd��<�!ؑ��WqL��QT	g�.�X�pߩ���J$�᷎��F1��~�U���}���a)y2&��$�F\�����.
H�̮����_��f+�/m7,��,��jӥ�;�4yk�#/�������5�*��>j�y��;p�!�9<i*ŀ��lx@�l��m8fZ%�W��>6��^���uD�w�-��#{gc
25��L	�(�����ʱ����� �kXCcT�D%)ژD��	`�3;�ě����(���R�� )�ӱw�Q��fy��KB�:��X8�A:r���m�I�b ���N��{N��J�hM��E{��3c�$a��ڮ#e�12+�/�"�N����L�[���ջ�s� �Դ�]�h>L���S=q�|u���̯!7���?+ˍl���p'b���/�yaY��I��h�jH�� ����R�ϗ�i��_�C�JrW�x���Љ������h �[-Z��R(i#WL�V�0�\���!H�㝬�T�<k���/Orne��fp��R�MtWE��.�36�	��[Ԯt$�t�,��*)��M�Se�R0� %{{��(mY8�L�I��Z�0D�yuZ���c����7.�6$	�G!�?H�˂�����_@zO�f��Շ+=B���	�w��k攗��W���&r� H5�������P��W�MA��i+��j*<n�p��c�oc�4�؈xם��3�[@/�R19���w������03����m�i��'�%��E3�A_[ ;�o ^�lS��?�1ح`ÉP>Qެ�M��I�Na���]��]NK�.��X�k:�a�%�N+�	a�P&���Ñ�Ŧ�ZmD��D��x�S"B-^�/����*|Ŭ,Y���$�ã����t��)��d#�~��,W�,A��v	��M���4\�c@)?���j�����]�˽_ig��%��/��|w�ۯ*��eth�{8�Z ����_U�@��_��u�}�Җ4F��i�4��C���f��m�-8q�h�O���<����Ŷ����	�FǍ=�����T<���
���6����e���B�a�6�W��F�	����li[�e��\!eb�m)OɈkq���D�:�n�I?�>���!����.h��e�|�V{ɳ̵�O�|b@w�KC<*��ъ~w��T��5�c<8���Wk�ΦԒ��|��E��X�����ؠ��k�T����:�z�rٟ�r��h��C�%0�|�O�,�$��_e.״x���[��:�XMA�ղO�\I��
5#���5����^����KR�\7,6����9������l�ģ,��p�XƆF�۟���g�H�Êa'��B�f��K�NDM�k"�Ύ\�ߝP���e��ȤZ�0��N���dc��`�kf{T��yzנ�Q�t��u~N�7n�E��Td���q�_+�NDI��)��<Y8F���4����/�5PZs�����vX�ٺ�D�Sn��6��X}��7F!����2v0�f�c��K�O������^����AW2�ߵy0��Y�(�c��)(�Wm94xOZ�Q�"�\[���1D����Bw/��y���C<�6%⇈2�2�3�C#,oUe�E���4D�PAu*$.Uw{�@���$oZީ�:qg4hk���	,A��Z 9fgH�}yWU��qḱ����$��نTN}7_>�iA�����+�N5k�{nNG_��H[�
���G�CSh�S(��#�*������h7���	֗�tV)�Q�����{�Rܱ}w��^v:�h�C�mI͖�v��&��;�+�4MmL�;�Q��LI�K�$6gs���)���C�)���
&I��T�-Lh�zח��UҰ�F���[�ʌ8�%q9���T���*��[;U=ٕ�a3"0Z#Mpo�`���$oRSA�"�$-/G�A�Gpm�����{ ���a�ˀ������uU�I}���.e3��%
�HT�����& Y�����c��}����&���j\r8��s.Ɨ����tTg|���z��<���|G�Ȼ��L˝��dX����W�3�2��M�8�4��"|Ip�w	�[���enƍ���Rmn}�p�ό�@��X�L�\�E0���:\C�f�L�ex�ĭ������K���e�0#����2�^�@���tS	 ?�p�}_
�E��*�� ���z���h���J��<��	Q�;K�q�磥���x�eT��yK�V^�j��[0?L�ٽ�/��%�mZ.�}���֘U m���e��#\:�_�s/s��e��&�\��&�����VҊWG���σ�?lT7�y��~.�As�L��#C�r����P�9��}D��%�Xyw���'�o����l�!�~ͨ<t�
DA�Z���[� �l�����Ŕ~{��aʣ�9��ŧ���ٿ�2����� ��,4��ǩ��R��\�o$�sd�o�u�m֋�S� ��a�\�����P�U�7�y
��V��i��YHV�N�3�p��뵆��N#"h�b�S� jqĻj�M�~��%�t����nڈ��}O�/��c���O����#�
������c�e�Pqʓ�+�����AI'�VWe��Y���s!E%_ClJ��9?�q/�k����*N��D�����[t�U�v�&;�Z�%��i��M�hqs�L�i��������6
:IZ�LQ�ݘ��"N�|)�[)��¶W�ui5��B���D��a�]9\(7� �?���A��C���W���Z�Dy��;��,A9�P���->�zW�AvI�0�5]��cG?%b �%�~��%BX���
[��D�}�ހU�����Έ��0�t�rͣF?Y^K����2N���~�U~��bɝ> $�d������]5VJ0[)H*Y/.2���?��a,�j&B�ߔ9��|�ҭ��&2-m�+���ć��� ���K�A�s)���/�3����8N�����-��P�2���c�]���x�E�^�a)T��Y��J�qj��+#����6�P;i���^�'��
ǖ�P��W���zc�����^O��]|2<*��{����������O��0�>\xJ���Ș]�jW� �Sn]vQ�vE��),SLAC���/r*�<�Y��_�U\]��u�����!~4?&���磫�9b$O���r)�PV������E�h���w��	Dj ��B!έo�q�Kz:")������FFއ8xX9�� J!BlVLN?��������da���r�t)����D\���9�������+i�КH�@pL�S XN�H�����E���&�b/����������Wz*��h��+WF�|t��gz#�F�Z��#|�����4g#���ӇSY�-(O�d_��<�7	�@��=�H�֓�
A;���㹳�n�円&��'���~ q����ן�V����!�t9�Z{b��_�eָEVu��K��J!��@��O�;��!g;ư��ߊ_�=� 9��Sf��M�\��#Ü����m;A)uy���?��6���`hi�3z)f?��'�܂גUE�Гw������~�����z��:��Q����QP�{����Z��>����I��X]������F��	Fp+-�eH��,#��'�(u?��M���0�>������>��v���m#�����f\�	�>e����C��� �2hK��V'�1'Q��v
m3z��K�"�;bf_�>	 <�n�9��h;M��M�ߣ�g%���Z��b������#\n�ڻ�S�NT�&
�ԔE��.r|��b�l���mq�j�T�������M�j��Z<<k��m�u�\�ܐ��6D9P���n������Eء��i�o�>���yo=��z".w^%���+��n��,��q�&S�s���B��ɈU���;w%+���(�#�&�3�j�d%秳�@áw�����6p��.���2�ӻ{���R�|jO�h���STy����}���p��<6�m��w 7�e��&����u{��z-�ԗg;`YȀ)�!���zLJF�^���M�xn�çX
qK>��,\O/[hE!Z�\!ag%e���o�v�Z�X���Ar�������?�l�Qӿ�{�p���'�q��kZ�.�kx}�|,���d���<��[!:L�,�lEP.q	]H���8I����a�U����q?�
8��1�&��
iP�����}�꧲-�cw���Xъnju��>zՊ��De�:��M�!8T���)�
P�������Zj-��qWå�Yx�6��d���_��]�	D�5��5�V��Z�\:�VR���]?0�	r��Uα��v ���0V9SDJ���h[�ݩ�G�p�s������.�z��W�U�X&��
�<�\)���� �G���쥥����}�(5�|(E}���hEn� b@�K�=���U�+f�s�)~ԜM9���)d�@�K��a���>��;�{�t[4���h՚y��ysV�rD��;��ڪF�Qo�v�J��A�ؗN�xo�ڄȤg��jU�8�pH��}������F�f�g�fu8��j���$��hd{�b2;�j���;q|ӣS��d��a�8r���R���hF3�Nf�/4�0�g?�t`j
��&U%l���<Tr|{�N0H�H(��SXb�И��d�ɦ e�#x�[�=�Y�O�m���)ѩ/kYD1�m�_l9�/F���U�q�#�o@�E��.e�kn�Q��Eh�e#�]�?����&BS�R��i���nI1�����I3���@h����%<*�ߎ��
݆�!3�-� ���gCb"�vŧ�X��>��i�ԏW߷	�T��m�������{��tM[zrW����D�}�; �)X>!���OĕU�K*ˇ�0}�"�WGQ'I$:�ݺ��%`���l���4w�����9�+�8F�>�f<�
�/�_����ԊԸ�n�:ڐ���;o�
��u8�x�	#TgT�O�eDX�ۜ!hzސ�͗�CwtRP~�C[��`z$�p�� ���I�h��b��T�/s�v�%\}á�GtS"�pJu#�5��2�*��&��<lXo�s�rw��j#(-lC]v*b�U9�8�;+3�+'+�4�Q � �H+�u��B�W6��0'�P�F���yv*��p-�2�O��Y���!���a<�c9����.10��S)�zXaN;����M�D�$oXD�����,��<���u��3O�����pvӚ�}$8��&_�a����~׋p��@���	��V�g��6��\U��<\w���g�*�_�,C��9ɼ��Փ�= ��S��i�;}j*��ʅ硏�%�꓄Fd��O^�.nfq\�ٿJ!�:6��� �-��7ja1W�ۨK^�D`.�����nq���uD��1MmS��,�r�u�>п5n��e)�ƨ�"P���������,�[�[tOdҞ��-�I�23E2�ቨ�{���]�����?Y�����w���5K��9 ���Z��Ih�������W���9����;���@R���O�V�G�isE�"�k�4zNN8�'�K�����)�M��j��8���ʍ-o�Ac�,i�I'U
*"��#�<���}�� ����<s��nX��B�AF*D�-+ϖy��JM��/�ES��뫇,d�"P��a(
���J��{,�w�m^6�v�+�;7GR���}�a���lu����kq�Ǘ*zSV�^�V����ҝ�p��k�Ės+��YY�z�@UeM�Ὠ~1����RD�(��=�+`_�jܒa�^q��M _�I���>�+�˘�l�Ii#k�}��G�&g��19�qUO�	î��Z�� I Z��1�ʔ���`�~�qԺe�5S�	pAg�	�)���W�W��|�2<ؒᗫCH�3�2��ѯ����#W.6~����Ml����d����I�N��͸XG>�B~Q�?��)ZS-A�Uދ�{@�%�Y-�w���_A�Ki8ͽ���-�\�Tx�:�P(-��)'��Jd>	�rS)�\yS�V4r�v����߫�Ng[�>���<F5x��[�D�0�d����A#�L�D������1t݅�͂�d�Hz��N{qС�G}�����WtB���r'�Ke|��]���8���K8�7�|���*GQ���>����N�a<k}�
8��1�Y4���y�O�<T,uy��
2c9���0�#�5�����l����N�O��Q����<��k;�şa�t;{|b#OJR�^��^�ĥl〞E����:�D?��W�J�v+5��M���
:.�rV���e���~��ڱ��X#�!Ҳ�ep�aB�Vj<�B�i������iM/�ĵ+$U�ˌ�ق�P.��;�7J_�jͿ�?Դ�A_Y�;�[D2�1A֟>�����.��	G�%�(u}I�XT�}���_!���֘�H��MǸ� ~%�Έ~�l�9�\R���9����F�9�LE߃ٸ�"�7Bhפ��k��
1�s�o�t�cܖRrPV�]I��YH\���d{*Vs�)��ٗt���A��΁Ɗ�$c.춹���7`��u�	��a,�3��\.«_Ĵ��Rl{�Q���|Ur�0D	���Y=���<�s�&H�0~VD�Ӝ�]�$����m������@ّx	�X1g
��׎����xᙥ^�B�a��3�%�S�Fs�����SG��(!v�����~Dj ��b7�+m{<���Η��� ��R}��6�HfH�i�M��5��2�9v��Y�?�g�_�é�4r��^Ү�|X�s��L�����u.��=�6+������GB���H����fk��}\�ץ�� 
���� �w*pf-?�~���(�!5)ǃH&s�k��ղ0}$��v�稾Q�dѢL��ٸ=ӆD�	��6��9�AL��!G7˷���@�[G%%���6����`�\��R�(�ٱY��듎9Q��Ű}aL1˜�� |�,R̪a<^-sϮQ�"�F�����G��Ə���SW����c�c^��'�N�>[�.C��t�g�!��h)&^��9�O�����ub��Z�p�y�M#���u�d��e�Y<����T��~��c̈́�s�t�b���wb@vU��x�9��5��ݦ����i���ZꜬ�_U!�b�5��tV v��="dx�-2�w���G��+�r��֑��IF�ÓDz�]L�w�c���E���z���7�����F59�[3�uH�1�����n���VXN=z
�l2��^�ܻS�{�s쾱��J�Ǩw�t4%�"|�����D�I �`�Οv`�j���bV�ԧ1���	�T06�s;���M�`P�F�I^K䵈@���?�$|����V����>{{����Mr�u+�qD�R���icԘo:�ַ�4=�o���x q�CP1�qkmq�*7�;'��sF����k4���1uj0m�g���6J$��/=�ی�טBΧ�5ά�Iw�^m�՘�����X5?���9N�.��aG`�Enr
�S�m�_%/�eӱ��}�B�>ߴ�.�JE9��We�٬4��� jz���b�D"5=B=���+������[֋��CE/��||�'��d��y����]ח�s ]�3���c����+D�H��8�9�Tغ�������N��,�$`a�E�^�?Te��E���јG���R�8Q���t�Bn^�!�;��<����s����M��W_�xo(�Im;ӯl�bI�/�������I�5Y]R����N�S~�m+���>k�������9�.Ϥ{�����Aig$����}��С��?.C����4|uh0Qo��1,�Nz�i���$�P�U�U�c(42v�D0�T�|M*4X�Z��Қ�����c�3���I��9�[�bf ��}�i:*���]�-�"��9Ry�%�#�0?_Sc҈R������-�x��?�)j�=A]a�I�+u����j9����BZ�a�\�	e�����k�~�2�R���B���n���)�� �5�f�Ƃ�sk~O���f�XS��o�+�#9
y�0�X��o�y㎧\ ��>;ɨt<��9qG��M�b*�Nz1[��c�pq�_wCy�Mg�Q��<q*�7��11���ğ�q;��<J9�n{;�����+�t��犯�NP�·��J"�I�{��N�@OT.I�1Ai7�,�j�0��S� �g/`;t�N #�n���E��&��kԺPǴ��?�t�Z�Ut��f
�Q�0ap��"��vE���jy�F�ێ��&\"OF�7ll�n��ՄC��#�܀&�)S����?D�L�+;SA��\�
c���U�+��B�%n��tq�!Fn:$W�bşyw�{�����f���G��Ah���ދM�׻�,oF���ֆy�w#�X%K�j������Sf��g���f�� ��hʴZ�M��r� �v���B�_Y��i�?�1�T�i�蔈e �n�r���H�@�nt��1>\n`I=/��3t��`���oQ�"b�+h}x���u��{�q���W[���0��]񇅭5�]ʔˁ�ϖ~+,%��ad��{�K��l-�㓵���8�?oK�=�䲀{/����؞�I� w9DP|���'��P6P��#9�2�T m��On*�,�����з`ߦ�wё�=�$��X'�V6��t���65ފ�`�!�����z�ZS���?��NY'������� ���di��A���`'X?����:�IU0����I@��l�&�7
�4;���G�kt���|A��8���y��Qt\� Yv	(�{�*l<i%V�N�ǜh��T���sgc����M���D�v��*��7�c0*��@���g���e�[}���|K;����(�l�te�-��� �?7��:@��B�a����-��Mˈ�\��}�p֩�9��x]�>1.X��U)�gv��Y8���a*t���ۀܻ��y�UG�H����x�e�*���5:�Q&��&.�k���t%��=�c`��4V[�9L�N'?�ېTV��vīJ�y�����h	n�%�@���}���[��(3��;�S30NLA*�JHW@Z�Ԡi�QȿQ�p��!�T/�����n����g�Yv�V�n@�� ۖ�x2	��#!1G�2�o�_�_{�.�Jd�c{������g���&� Œ�����5���P�J��&�U�m����%��/&��(�t����F��;�缳����0a�\��}R|���#q�ŵWg�P�W[���B9%O�p	�\��:�|�_�Rc��r��_�?<3I/�QU��
i6�qZ'��1��Ȁ�s�`��c�|Rɯʓ���O�c[�xA���%�
7�V�{B��#T�0�vs�8���������3%0Č3�Ο����D���XF�b
V��C1��8l����$�C���NW���~N�afܢ���δS�V��V�o�ǯ�������	E��2�����h�=��Lrɡ����m���X��ypo�Xʨ4��a8R�yR�]�pKɜyЌ�L����ޮ��1Z���r�z�,1h7��fCrc� ���F+�v�m�N�&2VSQ�ىI� /�nY�
y��~�4�!��X%�"���}��OQ9�&K�sծ�r���X�_z��@�{��� ����";Ji�&�S�"�V2ǣD� ���5e�3}���Bm]�R�m{vt�X#1�=VU��� ��k�`&��oK�+�R���\��FA���Ԟ���H3�G%���cn�ng�Vf�+N���݊�g���"�3G���}=�(�f	�э{S�L9����,m�@����]�7\
��}�a��
^*Xe��G����N �?U\���x)�����8uR��lӁ�q	O=�>;�N!���檚ѱa�:t�̋�}��@uo$�Ǿ�
s�����>X����<U3�*
9���� ��ĽJ��R��U]Xx��%����\H�7��L�}���AIݚ{CYNᅒ���K{��o�&�aW	2,� n%���c�DPv�t~�ĕ����؊{��$򚇩HnA8|��Цd��[��2}qs`��e��/�㈾7!�����]*0�cq�ƙ�LM�-��u�k+�o���n6$�P��P����{�6�$�L����hb�N�2���[|��ʢkR� ������j(�]��3�����R8f+�k�R�,�5$��x���=����&6�����~w�D�ш���6,�N�l��׌���G�:5S���FUH�'Ǣ׉����h����^�	pQ̸݋,"��9�G���rb��o�a+�(r��߂QJ���ZF���LY�$*b��*-MT��"r��c��r�e?���&�bS���m��B�PSbM�6�W��v2�c
�ln&&��Z��h8�X`NM��!�tE���Ax�E��ڎ�����`�5�{���&'ێ�:#���xgXq^l20�L���!y��W+ �͡o0�o�o�����4�Y�X�or��&p����~A�_*S�=�@�K<xwTh��{>rFߣM���%���wz�;/oB=�����q͕�F��`!xV�A�c4mG�+r�s�vR_q-�Y
+�$��ߢ)��^Ӏ��v�h@�V�n�8�t��
�~'���q_qDPq7s�)$t��	�ש�LZ���lK�?۷��Т	�1�du�>DmTW�0�9-����%�������͜3a�+FKƢ|�u�(@Bz��>-q W�i�+rFzCi��f�B�"�"��S��j�VInWI�r��]�G��·��s*H���?�)r��C%Y��[N6�B���/�B� .�� &��$��Q�� ��^�86�tf �2���#���)��1�uI�R��G�ww��C�,3)(/B��b$i.�����.ܒ�W��l�:j��M=o�|����v�Kئ�A���f'�L=[g-�>m��[t��EK'[J}ҘA��D,;a-��N���:��!�+��?����Q��WR����,9"�s�ߠ�@w��3��j�	�෎�5ێ�XyG�̀s��HDc2�"b�h���Ş��6�=��Tf���pQ�&ɫK��|��7m�!�02��
h�ȭ�>�����K,ռXվX�o���e#��Qo��ל_�,NX��B�3&��������\�u^�,�o�g����}�4j�W�h[����Qr�	]�1��2��kX��5/ݹPڤ�6��s/��O`���|,�S��!��?������T�?�O��1�ОKg=s��Ѷ<��$���f�����.������)�3���Vܐ"ob��M�%c�p���u���f-�R:Ys�:�OQ&��"-�e;�)� �,�`~�)u���O��ͨ Oh(�;���C'o<&B�_�z�̈��*ŵ�G�3B8-|ħ�Q�P߶}��`��Y���'JAPDH����-�9l��e]�w�� �h5F�|l��U\EAHve��ʘw��9�# �7��)�v4�k���0�_�O��-�v+�n�F������Y�H3� ��E��:;�����Z"���B��m*�^rt�h�\╆�R�H��٬hL��m�cnFZ�P��2�Т$aw���}g�Ƚ�.oҎ!Z;�.Yh{Ia�7��ɢ(�Ź��D��f[��]����󤖇��S'R	Y������S!z�C�s��z�r����/���Ѧ��'u0����dL����ҝ�SQ}*a����i�k�����k���5���F�i�b���+�n�ݑ���Z�m%0�Ⱦl ��~iB G�0 �ލ.Tb��uX�^��Hi6phض�E���w�A�J����<H���O�� e!��VY����ӥt���ڊ�Ӂ�v |�>��L?�a�]�*��t�+�F�jҎ��B��?	rW�]�Τr�V�T=h܄���{��Ol��|4�t�(銳��+�i^�����Ɗ �x��x��D�u&�&S�&T/��kS@m/%8������c����6�%��p�h'�8n��<��c(d�I�L^��*D�W ���o\�̛�qt�#&kw��Ү��5o	�Z��{_/�]��=TM��%�;<&OF��ca�>z�g�^L�pK�������mH�h�y�O_��0�1�?5��5��&�'����A��儩�$�X.�W�chZ�ڃ皈������B���Gצy��f�B^4{{�w�ZЪ�xtp���bѠk�AfF2+-���No'��A�5Ʋp���,N�RK�d�׉����� �7�ҫ����Ŧ�̯Eq���7��/|�	[�����,��j<����L�B�f >��	��*.:2�c�X�Hxږ����~P�¤MnЃ����Գ��*��$��0�xhchz�\<CLF������JO,��H=�RR�7����rȣ�
Y���@�i2�%	e��X\ͥkO]�OrH�����eY�~�I�ڤ|��Z?�Q3�*`��Cb~Gl6�fJl���ł-�n�o9~�&�Z[R�]��Y����7�L��%��9O��6_�C��,�s�r-C Þ�Ǵc�7��.!�S�ˮ$\��|�̢��%ZN��w�����V#?Ĺ�ON@��B�D��0NW(�Ą��WmA!veY��UN��2������wh���P%�Pӧ�2T�uWY?q��Tn�9������GeU_܃�ٍ�M*C��K����d��	
D�,k�/ɌJ��8�e���l�fTl`hJ��S,��B�Dڀw����,+!OΉE8p�:�@�;a�:7o�}_U�G�F��E���2����Q����Н@Mv��2$����[
��U��٪��m��@�4�!ث�0J��ԜM@�%���{!鄌�덳TY�c߻Ho|'�m|xظ4MZ�ڬ�"�#��3Z��fE�S�"L��V��Iӱo�<����*��ߛ%���t�՟�U�;��@v��3��CW�{Dc�%�|ۮ�[��+E�[�e_3�Z�q�/ �`�-_ֳ��U�jޯ��5>0B�]ۊ����c3�e��.H����{"$P�h��Ö1�rV�?q� ֿ.��4�d�m{�s�Ǎʿ���%F�����}�<
b����6=�������1�19�XX���e��n�Ea(jSϟ��w��|��Q,�q_��v��7}Զ�����_��C�f�5�խ%�h�[���/?d:L�";m:l,�d�Au�4F�hA�!Ҳ�c�R
`|�n(`G7s�M�<��$��utf���T]/@#
r;���h\DH��lqB� �&������9�@k�6l���բ>6��l�/��-v{t�~&��>���ÃU�hfQƦu�r6����Ǘ���Uw�[���8���I�>8�/rQ0���B���T91��s��Ԣ$@g�^�w�K��=� ���˺�æ�(��dC�;�����W�V,t��A��!�u��K�>�AU%س_k�,���"Z����o�a�����A�`�g�)el�4ޅ>f���z�`�|�T���¹P���,��E�3�M�V��Ip��r���ǓU��t/��c�=`$��[�|�"MA�Xܳ{�1�����޽�vɝ�7�$��k
2\Ko6�C�����(I���@'���!�sQJU���jkS*���rz��DS��������Q}�Y�V�C���9�ۍL[�>����ұ�L|wBG�&P2��;�"� ��4"��#���'�`Q��Z���ԃ0������`N����갂��\]<n���ga���;ԉ�A��Gާ)|��.!E���ҍNڼ'�����0w�B 2$�80�փ�勲}�_�H�����*`J����PB��)���0 K�/|����T��N �p[Sa�承B'!U� @���9�)��F���4uы�a|h��"iv�;�f8������&��"�<�7i?|�V�}�p��"ѝ�b_��n�C�@�̺����(��vF8%��b�c��&��G�A�$�|o6��^��Øc��J��:"�xC ���#Mw�,l����$�mn�UV�!���];-?藸Wu�ދ&��W1FȈf�9�C��)�~�_Y"��"�}N6�4����y+C��S���.��^k����2���K �0fi����Wq�-L>c<�������Z���A2�g�q]ط�;pkj_�BT��Z�t�Z0���8�ː-\�r(�D�n͕���k��:D��u��K�?����G�[�:;�^)��~��͗��Yá������4���M���)�c�8��׻��i*�\2F.�BJ��N.�Q�>��c� �sm;P���9�Mw��X�N(pZi�u��v��N�k]�7�_����+J��wS�"�_7.9o�-�v�W�"U�S^2�z
�����yJ���c"5�����Qѣ�ߴ��i��L�jÖ�<%Wf4����*8�6�ǲ�i��9��p�W��=��m�W5�$��R� ��D�^B}�����^�1@NZ�7� ��r���%����X�j��Ҕ��EH��0Dͳ�Ё�K�����'Z&G���b���qR��i3�5:^b�)%ڊs�~�6k�3�?T���ȩ����g��<z{̀75���� im�[N��Yi���)
;���qRr���a��l���T/���s⍡ϒ+���;(�-$�/��7ɩ��$��t���$����U���P;PK�tc3��,�����;�MMn_��j�!���s�ڭ�+��M�^y�@>+_O�+��O_��@�c�׳���ĕx��P��MY7�����v�o'&��g���(~�2&c[����C_|�,�{��O�;���cH�]��J*�	XX@.6f�1� yJ���iˉ�
���h��?pN[����0���$&���X��C0O�A�G��*��� ��Y�����Hy�b��w�\��{���5|U�����gMCI>`�����b0[��ד^tg��>Q�\�̴��~1�\F�>&	bI�>�)��O ��F΍��F�@�EC:���ƻꓥG����j9yp�4{}����ːb����ԟ�ԌM|K=���Ѣ�I��HEN��o�}��G�s��t��YtB%Dkj�!ثs�aQ�
��	����1� J��y�wN����̄�24���Ұ�|�u�uY��� ����
\&�WRCr�@��J�[�3~�{�A�\��~�m�ήj+�t�".J�	�����(�c�S��'#���vW�Y��^��u�/*ΖrFg ����X�nFiԇ�]��N:g��*�}1�Hk��]�<��Grk	9��b蘝��NнM'�@s��W�J��&H�W���\vl���')&զT�8ĕ:�u7G/rB��1�	w�5�Q�&ѥ�Wȫe-f��ו�6�M �k�a4g�Ĺ���e�7���-Uy�1҆
/?�2�Ώ�.�&�y�ł��.&��~:0h�{,҂X[0�g-DB4��J�X��mz�T=�Ȗ��)�Cp��t�����v�3��J!��	��꧘�%"�q��H�L�(��3q�FUO�@=������K���h���9�&�rŊ�͆ �CE�R	��Vq�I	!���GR��"�E�p#���#̍�G�;9���\�h��
5��g"�8����Lu��gIK������:+^ͨD�Jl1���q�q�x3U5Ш9!ؖU���g0�$G q�0_E!�~o�����Hd��B0Ͷ�E�o���xΌ�����m|/��3��@wkyHa�
.��`M_�
#�/ω�d}Sh��;Z��0��h.d
+�^�]<n��ܶ�3�rD�a�r�ւK�$FK���L�?�� �:�T@	�u��Y��	1 I�m�]/��,W`�BR�O���#�֑�C�+�d��uU'��QH3`�K�wq�3�g��m@^� �A���b�`�H���I4A�"ڹG%yh�Rn�KXw9126�f���7`���1U�`7�����u�z���$��'gl�A�ǈ\�L�Re�!�Ȋ�7��T���+�F��R}�9!�ܩ�tca1�K��GC݌�vVP���V�Aok֙ �)x�O� �YM�Ǐ/���mTXW�x<t�
�А�0~���d��}��j�q�4�Z���)����b?�(>w���IaB��o��on��(ӣ�6@���y�0����^����ɔRr���ș�/B��1hF֕�RF�Nn4(bS�O_�x,�E0+sA�z�kih��4=���������:s8�[2� �����4��"L�$��R�G+��}���U�=hTl�s�+�:�(p���z�́�t^u���1�~�bL���'M҈#1r�Ҵ�FO�#���X���	G?Z��Uݾ��9����6��IK��?k�q�P)Y^�Q�׭�ƚ�kH����ڕ�a��F���L�j:u$�\ΐuJf�����<۰���"������� ;N�@�/�ak\�s3D�o�u�����NjLQI�JD����o���<��"�����n���J�9k�p`/����c��3�~E�e����5���?72[�O��	=�[�����c�����NM�լ(zbSlv��o�P-�]vi�b俊ǋ�����]���~�, ()�P���3_��i&V�vҳ���;�$��y����DS�w�^�n���kX��=(���p�=VM���@�MX�5���N^�!�w�r��X��JJ�Ck��M��Ļ?�)��YR��k1�}�}ԢxP����N�Y�eP�.USU�K�7M�lH���Yt���l����(�什ՑP�x,�;J��B�2�e�z*��`��^��Ww����������f�b���2� 8�L��.ES4]07����+�ck�s�ߤҘt�]�]�m�XyϿ8�8x���4LaP�E׷ܣ��ڒ�&5��t���~���0XB��ױB����h

�})��漉2�0�FFE��̂|{���?v��Y0�{�Qx�c�ߒ5s"M�%8#���&����1��g�l/?v�0�a���<��齍�)�J*{�I_��|j��\LFŢ�������q_��bW�9#)��60c4�Z�Iߋ�k�
��T}�\���D��9`���<f�(���Y�rn�`�H�ȣ_�����,8��2�?8���M:�
�..������n�[(`ʭc�!�rpS�ӢXk_2��%���Ge7���$B�;?�FO=���!*on�y`/���}F�]������Y^M&���'IRS��(qЗݚ�t�6�f��\�4zܒ������j;�ڸ�X�Z�tfōF�OX�-qv�_�~wX��� l�7���M�a���Z�Z!cf�W4��.�1��?L��m�JF�o/��I���g��Uo+�mb���`3+�(�w�+IZ��V��=���ξ�~Ţ��_Ū����,<`!<�FXZ�Uv��[���Ԙ:��)?�a���K��jH.���k�������ý�Uɤț��.�6|E͆_�qA����#J��^C����(��1s+�l�� *�Fퟜ�����.���Υ=���h�|�\�#مw���3`;�y�ه.���9�A�z�C�*w���o�6"���T�N����?i���ܞ[�,�<�����Y��úqgg9���#j}���T���F�:3�[���W�|�r�c:	�/�/i��������*��B_��~*�eK��~�n�Sh[�.�b_h1xރ��Of��}�A,⡵�3M�ndn����?E�)��2vQD��P>��]��i���w��̓H9��4��P��_�-@�EJ �/�='�KZ팫�mC+��Nk���y�٘�"�W�!xO{Iw�|˭��Y�N��b?܏n�mEh9�ʯ�b�
���h4��ܯ��Z�Ak�&$r�a�N��3~f�!�/kG�0�?Px�֫GD$�x6�)��'��5�#ah�-+�u���k5²堰�׬e���i{��Dd�0�c��:�|�h�*���(S��Y��M��R�76c@Ѹ(6���2!���^��x�P�1��57�5�̖~���f:e�y;5A⯣e��a��z_�g���1�$��e�LYyat�})A4[rX��'�[���cL&5p1h�C"T�� @e���[Ŭ�Oҽ���#����#�G��7(E�����!y��'3�]�ʜOͬ�2��b�G�8������D	�A>�p�)��9>b�qQ�.E����2�~?�;� q�Ĕ�6Rbޗݵ���`2����Ţ�����H�[$j�{v��q.���m��"�9|��K��\�Xi>���6Յ`�<U��O������zx���1�@y�s�ǰ��-Q;i�-t��1N�Ҽ2:Qv[��1�$�C`� �2�vc�W
B�_�[�R��AJ��\!���K`�G�}�J&�J�����2�+���J?vF�)��9u\O8@���T2�C7T�sV�8�������MIXwހb����E��B�l>����.2z�. sϵƟ0캮����m@{�i�s���ȶm4��݁�S�| A�nF�"�!h6:!�ڲ�_�Pg��B�B9�[c����۴�u�?���jD�J/֚�[l�^�Р$��,��Ƽ믡r�Q� ���?3�$Z~�z��r�x����6*����l����Eϋ-�
CZse��3�3��f�6L��=ǈz�N��o@�ؑ���Z#�G�W��2�ƥ�j���(9�y3�SGEΘbQ�x�z�S��$K\/�!e`p	�&��"f����:+�b$���.���bSU�"�%'NY<�~�ã*�_#49:�){�U#;+`���؈��8d�:��1!�<�T�Fp5i,���'�^	��a&�Ԯ q��S�B6�Վ�	�.u������B�8��iMT�m��r����U?lǫ��/�m�OW�U:/]�*c���]h�ts�����q�ONNDO] u ��ڲa\��f�fBƦlu�E!�1�>�I�]Oﾂ�2]\|�т��+e�XD����J2-�:�C�T+�ʹ���>`�h��c�;�R������Q��q=�����;�F�e��Y��M�Yj�_sM�3*ӡH�J"I��6w���:�������NO�"�����rH^(��.���ʫ�Y�����c�<{x�e��16M2�W'��؉bq�\�e��O��j-����	�0ڃ$��G�ͨ�q�c��}̘S���ӱ̽�AkW��b,�O7�z��@dh�n۹�P�Z����5�l�i�����`��m���}vM?e�gڤT*�}5����^ToE��χJK�|_|�'������4Q�'���@��IN����?PI~�}�?���1TM��� ����xФl)6�^8��e�%7�_�p�
�?�����߆��:|h �RN�����X�{"��Z�s�kI���jU�D���������J�z-1��&˯N=0o8�:��  1��:d��n�+ ��4"2�V�V��M�l��YMp��HQ8 �d0�~�-�W�V��.�TL��P�_j�G[H7n`�h�A��)�T���bk����̅�e$��?���ϯ��$�g?�&�+˒��_sq%��=i}V��¥Suvp�#�q�ɧ�-ʓ��-���r<VS��}8��).
2(vbd�qaM� ��ϴ��p�b	ɦo���7lg �ݪY�!,xv�h(�^˟��� �ʹc/r�L�L_�
cS�΢��A��UL��伨�ԕ��6���=���P���U �
K����t��I�#m��Z����J�ھW�(��gSώ|�9�z��E�|i��G��H�+�u�?Jj���K��?�q��ib��S��e֎��e"M(}職�a,��[Y�Z�m/�)�T#���}�yQ�Q�]�,C[�������Q\\��u��8�����N&�\L��h����to��`y(֚�[��Ƈ	�@�y�2L��#����A���O��$sD����!_����Z��B���`���!�����	||���6x����ݡ곧�}��F�>�0���h�av`	�j��0��������`],��y'��w�ۺ�wiV.�(W}�-�Y����*E4|�x;��"#l�9�Z=Ш��Qm��|�1��f0f<���M�?�_P�[�Y���V�ğ�FBN$A�\�(-E�yt�R�?�#�)V��Cj1[��- ���-�cc�&W�����=�����v��(�aB��zZ��u�v}���ղ��"�L�Ԅ8sM���DR�}$)�K׾�o&�!&�x\h����5u�Fik�*�=�/z黋���U1�b<N��
Q�k�G@���B�@��H��#�����g�#+�""�\�l��Xl���T�̯"
!V6Kʁ$*}������+�V�[�L��ԋ�I�߃�v����UE���^��Ц�q0��G�Z�R����������n5�Pp�HbEUQ����-�\�EE&:�y=%�J^b I_(,�1��J���ۙ{.Z3u�!*�k	�,G��p\����8�'C���#�!1.�C�
��܏����7�fƅ�ȎM���-C�$!ؓoNw�mlUB�X8��\��=hP�7[/�Y؝Ͱw���Տv��I��s�+/��#`���ڰw���X�,뇩@�, &��柰�֜��z���fN�����Tbf-܏�C�W(��ë��}����5`�1�$ɢ*�F�2��No\����45F����|&�� 6�*��R�=�a4��k3ϱ�<+x�b&�����k˜C|I=�G������J,�o�L��uW?/u�ɇ�0,��C�v�ԍhv^4�:PDa�J>j��P�;��r/(����Ͷ���:�.Q��T��P"�O��:$������@̸�S������`"Ȁ��qy@3s8��#�Y�c-�66�{Hb��vp,-'l�u�G�Zp~b�2�ٰɿ�Z�hn[���"��"������ڜ`�̐�$8�>ҽZ���-�%h�s@#���.�tL���<���ˆb�&w�ëO�9h�ʱ��W4����?=�'�xi�t[?.�u�l C�v�7%�(w��[��c>�8	�;��,�f�X��@�G�Ý7T2����ϲq!*\E%�h����t��~�ᰎI-�+���D41p/T���쫌��u``-��Au���I���<R����B~����d��3
F���Oa]�!b�H�l�LMK�j8s'X�d����繋���<wj�7��H7rZ�j=�F����7���)\Hn�&�>�9u�z�Ζ��*ν�\��s��j���;�y�yN/y˘E܆ !���Z�]�o�R6"�h�*s�]X����$����3&���4��+���"d����:gw���(���O#K��V�IFb�ȸ�S� Z;�RO1\d�t�q�Ց����4��qK�W G��}o�n������yy>�� �������˪L���,��*�f���+/��k����E�n� ���վ/w[+��-������s�
��k���9{�:#D�8���t8c{$�C�pVDh��^�Ļ�7q��׃���|#w�K�`��|uQ>4���*Ӄ&����G�R��꓉�� �G�X�(i��ā4vu|��KZ��܄N��3�v'�7���:XojBj7;�J���%�
����E��k#&dh���ӥ��������Lgi? U/#~`��"yc:���f�
��>X�@�u�,M�(� ����l����š�~Q ��>M���R��傀K8�v�����D���H�:U�O;n�t����0��h8��Ӫ����IΡ��#�I��I3��'ڄ�^�Z-��\�6Y9e�;��Dڂz�>��P�HV������&[O� �'Rzm_�P��.�֤yT��G�%N���$(���q32Z�(2�5�k��b���~� ��P��V Zև��f(#� -���98�X���>sU�rQ�������)�a��haք@�j����0�&�����q�'�:>��&����!<U=F˻���u1VZm�w��F~�T�G��FʱY������x�c��i��C��Y0�2� �ׅ��E��_"G���xr걵l��˞wN���}�7�V}�ℬ��A3V<v��u\eHu��d��NC�N|��9�*�ߠS��:K��\�g��-ƿ�����������XulG���|�4��R��|>�y��Ӄ�}Qթ&V�4���z�r��!�$F�̃�fi���N��H]?��"���5�h������^/bd
�d��������<'i��+��,��q��RZ;��7����Q��#U��k�)2�p꡽jVZV ���B_qt���:�-�PrH�+��wJ�&�oL�A�Ҫ�x�����S����KS�z�"�Wʑ-��m�~�\�i"�]�Wbz�(y6�[ �������.��J)��?$H/��+��B֑�������T��_�a+����E���"�?�y�;�_ ��U/r�G�";H��Yl��"~�܎w��N�
��\&`jI��~�����-�D1��q���Iz*��%xP�EjWg��F���(	��Y�0�1���c�s���u�@�fw� �wj�1ȵ���Ǆ�B֛�=�3��f�n��������L�~�*2�7B f�
1Q���O`d{��k{���-N�23C�a[Ҡ{����d(��7'�օJ�7���9.E�3w(��Zy�G�aw�m7j�qUug���}48pIɐ�8�{*v?�2c{"S[U	#9�%�"�l�5=��q�$�>ĕ^p�"��{AT8׎y���¸`�R�/�)�ʅC]���B�+�$��ӟ�!t��A��(|�V�ܘ�zQ��L \$KW� 5��w�%�H>�Z���~*�%�/�v�*�A��)5���Br�_�z�5�@��YJ��+�S-��[9-M1k�!\�j��Y�	nQ�,�+H�|W3,`:���}�( Ɯ�]���W�.��ȫU�V�;ӍN�f���9y�q���:l$�pY�#{�b��M����w%�X}@�.�HP)P����8�4rw�E�)Tr��S,g�'S��3������y�͢n:7���7SI3���!��yZA��C���0���D-��'���f��9���m�_��l@���}v*q��9@�^�q:�h}������#��1����, \����f�J����/�}�q�{�Þ*Vn�}���m`�iq��8�PR����d�co���kL9ޥ�#�L��tz� f3�*��
�`kc1����^�rn�f|���Q宵2�D��x��ۇ[����\�7?z�$U���3X�r�3R��7�4�����]U����mױ��䣕���7 �s�*c�&or��u��T�Ȭj�i5k_�Gs򵢶U�hs���{���T�r�ЕF6PQ�3�f�麽ۜ&
���FY��(?���eϨ6��?-�v��#�����p6w��Oހ>�j��H�0;(��d�K:��e���0X�0U���D-���߿������H��ԙp~���7�է����9���6�;ѥ�%_ZG��`3I�ޟ"�=�;�'��-���+�u���-i����NB�FB	��wn����0,2s��̃Ͻم�IKZ��M�׶�_z�w&D]r�P�i��L*�>�`�|����.W�ȣq%��b�� �ƵfΓ����0$1�����]���2-��D+�NNG\�����)f��n���_�:�l�O�D0�v,��c���+��v]��.�{i󕂜K*�l�{�5�ɱ�h
�j��Q@��H��Ъ�j��`9>�C�҄@��=�=������������Ѕ����N`W�%��r����s�r�g[�L�<�|.?�ljfK�f�?&Y���-��`�?��Ir�e|���u��"e�t���?gU�����4�}�-p2�>�n�����L�l7�NUH���v� ��'Z����6�4�p�l�A��5G�D�S��͜Y�c����=��p��2��c��p�G�w����Z�7�	qUv��8�Y��C�s�t��.a���j!Z�_���]?������	D��8P��n���k��6�+MY�����1��ٍʽr���E�ܑ���Xj$��!V�P�rv��(�g�}3d�d�S�#Yv����gM����LS�^�-� �� ���П	X��7�g�0�o��`�d���O]Dwn�۞5�/d���w ����¬w=J����N�&��A*�v�I�٩0}���JA���Y�idE���,����ֿ�ĽAXfm�ﱘ�"O}$���j���<,��;�ᴚ$��-Q־#� ��DG,T�޶Lؽ�pa��tI�O����é�1��pő^P�����
�}��O{:���n�-�Κ�Q�-zo�0���סڳ�ݷz���b
t���:�x K��(�B�o���)��K����g�߭�d�.`c��N�1��g`��-n�8��4�*���\M$C8T���\�e��!��F�`rG8 p3�{�X�S�L�*rA�!�;�#��	h*�M̴U�y^\����_~x|nɬ�D��;ԍg�f��	�׾�s�kyM�8���y���!��s[{�����aI��{��)���9���b�co^O<)?���Q�����N�/��P��A��Y�7�7��6����z�lm��L��b���k�Z�������d���P��Ruy�'���'qqP{W0?��9	t����(@���UkJ��p�k���P��ޛ���Mj\�K�r���!�%'E�l|�,��
�S������h�#��\t��!�1ؑ���e�[�j��<���B#�ɑG;Tu��
�uht�� �_��E7O�x���T�@��Wo����Qu������a��'6�r�9�gPK��,�fA�ף�1߲q�}h��}��.v1G�w퍈wno�JC�z}2���_���M5Y)�,�����s~���.���A��|����x������C-RW>�=�۩��Ln,�e����
_Co���u%Yم�j���VX�Q���w���MٲM�ƣ�^���_���K��#��W˾��am1����X�|��u�Z�/�f��F؟����R��ב�\��+t�j��[�<�w�P�<Q�E���z�u{����LRA����>U˶�j���M䅋��4ke@O�`�<s�ǃ<!���b�k���Z��;9�,'�	w�s�%̍����'��|`{���$��� �0:�+p�bn��a��������Q�~×�L�c<�^���9������VՃ٢x��ݝ�U� �C�?S���d	g��@�wQ��N#�?��,Kfp[VA�J��]%���g�08�j,��n���=��g��w�ˎI?�U.u����q�*�p�����LbUV�HU<��͔_η��`�?Gc�޶�ׄ���Zf��<�� ��qt��.nv��4�py1e!������~R���Y�5ٽ����?����1�sX˰t���
^��5��0:���dͿ
!�L�Q���8q2\W7��ecI{�,1�h�9���u�v
Lڜ�׀��}��S��	��	#O��ok�#�
f��/t�:�Ak�-���)sP����1�s̤��7�c�k���z'�z�C�˞�tzt�j�.��9D�a
���<����g���$��XD}|����#�L�_�
ug��}�y�@�xɓ��Le���&��q��h�����v�z@k%���^=<K� �ED��]b�)��O�8{>����2�³��#��� 4��.�J,�4y��nBd����Y�@b�n��z�����eɦF���$�MoP�6���F���[�C���K���r�M$" Xz�RC�Moi�ݬ;A���fwF�h����/�>����1��AH�A�v�\Ⱦ���l	�A�Z��S ͯ��~����Z��x-8oS����]�>W�4�qk��6���+휆�C�/��?��\���1���~,]��H��R���� ں%J$��g�7��_��C�K�K��mbw��w�����)���F�@@�:+����H�+xn�i[|î��dG?�it��H�i����^\�&ךk^���Q�����5� 6Ҏ�MK-\��C�Ic�U]�T��ɝ��j�Z�\��W0��R�v�=e>��H�|
�ˢ��������cNpC���9�`Y����ʹ���c�%C��G�qΡ�?�)J���!����MfQ�	dF���ߴ��s�H�v�x��촰�f���M��+��;��F�����<�j$�����1\<,17t���p�+_Z�_��,#TZZ!�>�6��O�l���*��Z �M Ϊk[�P{�7s�y��Ç����>%�Ꮋ��y�V�Ĺ��t�28�'*�����آ�b�F��ٚ�#L���ʩ��YKU��.7��*ϲ�q�@qʃ���@!m��6��N&���˶Z����j	*�J�Q�؀�B�����O�~9e�=�l�J�r�S����K�`�w���ٲ��0�Q�3hx�t��,Τ���oc��<*B�1�c!����zM�u2��'5��#�,K�۝��1v38�=�r������bVBdf���q�h~ݥa��h�w�k�b�߬��|�iQ��kFo��ƛ�K#�㭟(���A ��T���V=X@��t ��G�R&������ �x��>ɿ��
��(�d(�ɯMK
�j17��\����&zې��F��J���w���1'�>!��B���ݲ�{+��̗�'��?Hצ�0Zr.��&޶��:a��	�j�g��|���"��� �x�ٽ�h�3�z��X�u�`VQސ&2=X&�@ɔY�!+���h�}�o 
���r�f͈O���T9�|�-f��.kS�"�(�Oc�
vg��l_Ǎe0�K�0�9�	Q�<���6ؒ�������봨$~�h���*��#��Mx�"}?������J>E�QU�z�_��"Bp��s!����k���5R�cʄ#	��an\F]�y�- mN��,.�����!��i' <�&�����X뜇��c��:�wf�9�7m��*+0bk<қ��CB+ݽL�xtEȧ+�j^�#II~�]Æ2A�f���=E�]���"��\ �0�Ӱ�X�0ʄ�$���g���z��6��za�Z:h"����8:��2�y�"�V�ta����VF.�9�h�Ɲ^S�i-,A�hS���G�vv+bS��W��㖯Lk�%�z�q����g��Y.�?�Ǭ�p�}/=ˉ@��n͔㯑$ (w��h�?K�����v�GCj��՗ƃ�辒S4+Al��\��� �>�|t��]�1(��d�bò�M��-�@���R���3z�'�ӁKr�љs��U�|+�~���7�0SzP�7N\D^M�����3U��cZ��dw����N�}�ؕ�!�}Xת''0?���0��ͷ�n!�rT,����Q��%yN��z��7|�d����cc���bۡ�>]�{�E���,��T`L�������%����<Ё��*�]�T�h�ٿ&I>��A����a~v������G%�q�����ɴQ�W�&<��I0�Q=�!0)�Eg�g���<N�P�U�P��k�U%=�(%l=���o(\y��n�a2��)������21�a��E�f��:��G����4��)�-(�&X/$g�[�"��W�D<�yu�WB���"�y��f%��2����w�jG�MH+������\R�W�:^���S|m��Ɨ��%wUcK�\}v�SKe��+��Mi���__cJw=�q�0�?������ʦ�_��p�Kj&�\��l��z[7����;f��i�,�>�_��@LŇKa��
n4�z^��	W��Zt�������ɋ_E��S�|�n�:������ ���1
�@.�	C-K���P>����Rg��D��{y��E�5���DEGF��pg�@㳞�+�����f�N�[��Y,<8� $��u�k������D�LqF�r����L�꡿����ڸEL�'�8W!��c�:T� &}7Hz.��������l�(3!e�H�j�+�U�d�D�3waL>q��(�)��!1b�++"��s��u���9@��r?r�ͺ��s��2#]�N��P������o����	�G��.�����l	t�Ĵ����߼���i1
�J�N�*\vE8@S$�u^F�:���cI}W�X��I�7��vv��H�J�x%���$K��m�]�2P`���������R����p���e+H}��ۭ���N��c��M��$���q�v
i$�ـ�^���n����I��{Ӌ��JƵ�g�y+
zp%�e�	v�k��97�5�(�5�����v���#�H��w�J�$(���NK�eu�v���å�����������7)��2��D���Է��:���wM�s�c|k���8�_��뚩ZsPH풛@M�gK�Yn�l�ŭ����uT0�i��Aj�8��ʱ#�4'&��M㘏�2nQ�?@��K���;��x�ב��.,d]��(�kH��:�Q|;!��d��p�I��L���&g@����X(��\/N;�D徍aCˋ\'��k���&qM��jp��1��N���Љ=���n��SC�)��O���}�������y��[M��i'�1��Z�θ]��R��`JMS(��o�a(��P�u���m]J�sDv:Y1s(������5��z�\`hu�q���K�Q�9���eI����٢rK>@��Z�X�c�ʑ�`5�ƈ�2"mqٟ��O�����`�[}��B���9.LN4,X^���S+���e�mQ�@I�1�zd���n�7+ �GT����X�JYk�Q�(��%#
�=5�E��o�$%��(�Bg�A��gW1 +�eҍ��e�wOTDKT�_�x���k{t9�(�)C!��T��8�eV���:�:�B���fd
le]��]���m�Q=�pT�F�UG������
 W���9�J�Gd+�9w<td�Qw���*F�c�.��K��֬���ӌ�p��)�2*��ҋ�(}v��~� �A<�y����/��/�Z�7�X17W]�[���U�]�6����>\Dlk���)h,y"[�tQ�#� +]X ;�5?����D�TɅ�<�ap��_�<�D�(껜�@��:��ozE�����p���@�J��%~�^6��l0K�Z�<�E/~l�	G�,r+gC#nP �j�֓�+����X��E�>>��ȸ�}�EA�[��tIL#lv���w�H������
β�yZK+�����`���\�+�S��2�����������RHg�<��N^��>e����9�L,v.�H7��>��$�h/�l��n���U,Q���%B�.�)� �z��a'��2���(�_�a�F��Huh����CL$27��-��Bnz���Z�,t�t�9b��~_o�	���?�U1�&�I��5�a�M,���ui�X��O��sk~5j�q�3w�A*w���kS�#�J,.p"��B����u�8	}�Nr�b"�o�L���P`����m�_�H`@{������7��зv�y�3��;d���W
3k l����9�+p���-":`)!�#�eU���;��PR��P��S��Hc�3zQ�����^���*,`�O��R�ӌ��_sR=�h���Z
Z�e��7�ǯ���n�"r�Z�kq)�-N��X��{K�*�_u���-{���CxY�*�f}0�n��v�n�Ϊ�/�G@�{���i�:u�Ga��<��(�����Č�#y�ӆ.f�^����{���fӨ�PMA%��7#:� ���b4�?}@��f�I~?��d_I5�R0>:��O�[�#�n}c��,:��%���6�&)��s����T��1��n�y!<x�ʝ}^��@��H�R�IS���Μ�2�,��<�w�9)2�H���p#w4Ăv��r;�K�Zny�£�8f�Q�a��Ҳ������)v�4Mo���?Kg��.N4�"3꙯�T�@k~���x�0+����AS�`��iuR�9��gAu�����jg��<�u���	��T��/�w5���P������rm"E&8��mP81�/l����gKx,d�\3P!wv�9.�3���F�l��C���*aɖ�9As.A���		V}�/��ŀ"�h�7��bV�Y���"���i2\��G�\���g}�5!(��O ��P�o*����Ǘ��m��kPq:�З~q-J]�7���2�@-�IՉ"�˨(l���aU�U2z?:���?��vmB��Kg�YI�x����U�$�SOo?��nm�2cD���9N�7�c�wv��_y����EeMa<� �f�%����M��;��#��$��[
��Ed{E9��s!JZv�8��	��k����Y\Tq��ϛR�*�$�:���*7�����P�_樝i��\�5�������bV_7�5�H��lQjH^�;G��7@F�g�'��z,�[+�/�M�ẵ TP��ѳgV;Z��9��k����Q\_�"U@aw�5Q�i�����S��d�:����錠��
>r/a�C�=����>Ai♛�ĉ�Z�������lyB��t��N�EV]T~�qb߄܂ڏ��k	�U�sL�}�����;m�P[(c�Y����V�>�����Tp���y8Xɏ�� [[)]�}g����+�[�^�#@?��D!��4+�Y��S�=
'�=��+��y7]��ḹ�-E�~�F�����2P*� �Þ�aGã��*��=��/v0��c2�Ulj�����s� z}����Pϗ��eU�@�
��~D|UJ8�jؼ���Y\���0>X�=��qE�e�:�g� Z��+;�^<�&��T���tw@���ؘ3���[�Ǳ+�q>}����rI;	������^K]��l����ƀ��/�ߖ�՗@ �Dy���	� RiZ�W���qJ��4���O�)�4o��N5<��h�S5��J@�9
hE50M�Eo|Q�S�漐��éf��_��(��J����7O.8uv9T6�?#R���>lX����� Ґ1R��%Bۿ���4�I^s��K)2��X��>�@�A��G���/�Ԩ��䶣���o�iR�5���	�/=k��:2g���؄*'�H���� `Fk�L0<n˨+�{._�B�{�.���?��` ���O��Z��v� xaDK�a�r�����u?�4ݡ��c���E���Õ�A��eP�S[=o���&މ��lS?9�#
�G�譚�
�2̀;� �8����D<�%M�
2�5ިދ<�2�s����a	�q�E�X;\lEv�VŇ(b*X�=I�#2w���/�n����@X43ge"�pj"�A�TX��F0�z���Tf$OM�J�.��˶��m"���w������N���f�n�	�C �J��Η�'�rjNI[�v��vɒ�0FL���]��������jh�r����*Y���UI�v�������x��z�bw�'�9S#]���(��B+x�ˇ�bZ��M[�\ȇQ9��GX�Y� ��昀�.�:�G�N��l2�������\Х��}��LM�9`޺jMNhk.��َ��Z��f�65�9mr���#@s�����-��2W�P�����y$�o��,Y���h0�oH#Ɛ��SYP���@P��`)'��겔�j�smbz��V�{,K�r��!�qo�`�R�s~�>x=N-'Ap8��p<A���ҁ; ����|��C�}�:�qYRO%Ն-�B�骗̉�D��A�o��Fs��d���gKZ�/H���fnf����s��K��o��v|����(�zf��x��c-�!#�"J�`�S��?����y��������� �Aq W~&"��9�y��A3�X��1�.ͽ2�O�g�p�v~��d,�-�u���5�|>!�S�V6@=�)G�YG�s�?X�|�ނװ�Y<�<	�T����w�-jsg[q+3��5Ɩ,���;5�����)�*�qa'L���9_z� ���&�u�NVM�U� ܵ;���1�?�X�c�%��X�J�yzB��u.|����l������rz��-=T��Mj�.Aڲ	���C����wP�&���O�����Թ�L���������]�/��:�Hz7�2�=��$(Ew3)�ˈF��4"�_eb#���y'楁c������� -웜�MF�&��Vg��	H��1f��p��Z�ԩ��[��¬����F�������� 5��*w���
�N�����Hc��n�׆���+��Nk�����������MjT�s�!�(�Ι��W�H/l��\dT�����C����K���H�I;� T��,@�@���H���	}�=������d�H3���T2��0D��K���O\ߓ('��8�����Y��%�D�����>쎾��{���=��vg�t8�t��l8�?����6�{�B�<�L��鮔%,�k�X+vCG� b�`=��d)��h�����
s����t�w8�h�	9�����?E;	%_/<9�|
���uvY��|{����yE.�гkd��#&=r�������� �NI��Qjɸޮম��H:{ip�n�DNE��#a$��� ��0��2��xl��"R;���IǞ@ӑ m��;?�	0C�<��9��c%����j�@8+�O���X~*���JU~#8��Q����7�R�G$���2`3��w��l"9�ҕ�+D�ٷv<����5Re���N��wEݵ�oA
~8E�]�v�
�8��'Neg�AH��'��3�we�&����.P�.,���T=��XD�:Cψ�7��y)�EsM[�c`H��K�N�8�j���> Ե:�w�r��`���h���%c+��@pb#-�C��D�P��� �]�V��1�ͳ!��5��	P>99�G&j3����"x�$�I�QOO����'D��9z��X����t��p:M{�֎�{�l�G�tYBr�xs�dֶ�:b"�a ����r�����J· lQ�t��i�9l֘U�M����"��¯�.�.�4vdF[��1J�ݦldzYY�`�t�*m]���ބ���/�9>f��4�Hn�(��`�&Z�(N�!��)���6�d�)����c!1xbL%p�uI=_����$O3Cn��y��~����q���:��0�I��*�5cH:�o����N�����I}���h���?� �e7d��4���0=�T0����x>��z &:�;����+�q���)�u~�����<ʒ�Hv6kPQ��������b�1��6�F&�Z��XL�X�,<�����$��HbW�KҔлi��Ĉ��������,W��K*��&�5wd��ǰ�H�c%�y�o��h4����.�	�
����`�J�g^��n}�u�#Җo4)�N܅Ƅ���O�D�*	�0�����Ϩ ��ӁȞ5��έiy�׷m�G�L���zZ�H;(w��1�S��k���͌�G�g��x�<x6u��}ê�7�9>'O�9�A�γզ��w��t-�(F K��)6 m��顲�ӻ��h��ϕ%T����ˠ��K��$܃�/����ć���#�x���D�w,3=�<��Z3ĢL�}�t���:��g{�5?���2�D�]kZ���$��zyoQ�Y�qU�y�I��,x��G�9�t�@D�_�&�<C�3��Ց�{f�Cc���eT��R�8 5��|��ѻc�q���հ����aI�6�����,h{%K�%R����c�b�5�R>��oef9�4�I��ȟ%����z]!!�Q'b9@���M��,6�\��������%��N���n����d�����! �h�a���b���B��G�g� ��(fj�}����	Q��Ҳ��׌[��㷵m\���q~���ݛ4i�96%v���j��t��B��2W��%��p^��k3��,��y�ן�#\=˃��2����k�������x��C-s�]ޯ7d����X�eZ��|�!��i���[�zV����*���4m֌ԙ�j�����
�$w���)��+����t��QGD �S�v?Y��7bѧ�g3GX'Ѱ[k�t�^Tl	�[�:�ġ����+����9)�81e�#vy�����}�.�0��zt���d�Nʁ��\�櫫6��j�][^#J �Q���������N;����eHޝ�lG|tpp�k��c�o"W+�x�ʃ74h����pt�T��"�@iP�D��b^i�i|�������h�y�e�x@x;P��B^z�-t�9�c���Btb?�c�T6I�sz8Ղ�;g���p7�;��t�#�����¦���$��7r�^9uI�6u��=��Iy�RKZ'XG]G}������]�� ��>�h�q����x�d�M���5�:�!�04ɚA��Ǒ�?����{~h=J�;dV{ɦ +j�綔�[2�V_��&~����xy��Ņ
g4@t��1�j���A�&�?�
��(�L�W����Jp�v�e8j9;�zJ�	��(ǳ����Ь�dҮb&�S�o^ł,Zt(_u�[7�#HψLٹ�Ŏ�m�WRh1�Y�_�R�,h�|W��v�=<������V�e^L^UM}W��W.�Au�^l�zߨ1m�/��1x|�9�'J��0��"���V��	8+���.�z �篲a�n��TG'^�<z@'%IG�t�������}���u�.��3\���3��'��<��e��$��H"ƭ�ʮB(n8D��#�g������gٍRݰ���4��u�k�s@mo�������g~�u��n��^�4uҨ�usQٙ�ʇ�A�y-�F8/��}V�7���n)��3B�H�宋��jx��U���jbğ���XhȝMl��D�>��<y0x�N��,�+�J]C�ݟiY�gZ�j�T�WY��0�7LKP	��q{�VO�գs>2�p����w�-����Uӑ���"��jp�j-�B����W��o.����ˤwW�K�oFGM���-�ɺ4!�cZ�*�8M�32����|���e��C�Y���$������?�������c�hQ���2L��b�L�m���v����MHq�aYq����B�#��b�b�߈�m�k^����6
�j�@�0Д̥����}%��ŅTh"�BY<�/�(���b�5HJ���,l�~���R�1��c��-*M7C�~6Y�R�0Qn��=�#��/m,��ǀ��x�5 U����
��
u�S֊�G1X���18�)��(��@�+�-�Ѻ��RLF��o��K��+��g@�nq�q�k�����f������جu�S�ZY�ˬ�І�MASy���, �,�]���͉4�R�Y��c%���P���*�1Ѳv�P�����}����T���	�u+�C�mw�C���M�i��L�E��7�^g
V��iw^��H����7�@���ji�M������f�/|�3�_�c�v���)��d����:��z����T_A,�DC�:�+�}LJ_V�[�i2��{�ӕ/���k�4�y���i �2˭f�t_L%˿��I	=`�����	d�+�4���d��O���1uj�Ϗ-��P�M��^�1=<��rW$q�=ԍ�Ą��L8��I	lTi䖢��K��!q��+n ��q2/ν�ԻG�
����I|�J���KQp�R&�j����U����9��W�J��ʛ�x��t�?`R�1�?a)�qs[u���/)w���J� ����"�W *NE�a��ĽK��7���e��G=&�z-n���t:i�ø�w��fыF�Q���K^P_�G9��K�"���Xڟ�
1�\3�\fD�]+ʶ��M�\oCI3�1;2��R�^̼�����W��1�V��l�F��
7��O�,����E�"e5A{���������C��{�7�SQ`'���Y)��@����E���Q���ޯg�x�9փԓ(Y-�l �K�&�Μ�VO������G�<A��Cj��	pY�Ey�ヂ
��ev�y�s�.�؜����в�tǸx�"��.���pC���Et.N�kHϺ#߾��H�;�=���H��棾�P�r(iPl3D6���QkH���6p���We��d����?�\Ɠ`O(.:CI�|�fڏ~��ȥ����?dʏ7K]��s��8�����r-g����ӊ�=���f����R$%y�ʹxݣ�$�*��Al<��@���E���v5?�Ĝ4�B���q~�Q��u?��2��+/�� $��k�/>�ho��.�^"|K�(�Zяy�5�����&�$ H}r9�2#R���/�����S�e�K㊘]Y��Z���U5V����^�6�v9��ç��������H�N]��/��1�,��q���������嶯W��I�|]� �ٗ����'NN"3������k`�y�c���E�n�I:I��������X4Qy���fs�PH:uN�X/��z>W=�[���2��'������2v�R>g��EK���=���2O!�1۽�e�K�أ� �~}��c5��m��������|�L��,�0Q��7�#�f�$Ѱg���Xs\u�(��`��Z/���	|���OP��;�p�D/��Z������;mõ�
��2�q�x�q�M����ǴCX�O�(2,vW��7[Y�=��<џ�aXn���ZO|��K��A��.�Y*��ZG\[����,�������<d�V�!��Rd��A�T�;�z%:��|�/*��T��O���f_V�`�g%(��2'�)CR-�h�X�ƻ�¹/3sD�(�bf�V�U��!ٽ�W�3��7|����EҸ��|� =5�M߲f9g�T����0�קAXi7W�j�~�]��fc�XV��e��*����J��wd���#p`�Ap�ʺ��1n?n��*��9��g�Jc�N&��h��9[sd��w�_P;3o*��/#C�D���&|Y��ٙҗ���he�������my͋��e�P+��?Vf��	��� n)�R
	!v�6���R`�h�.ݥH����R�cV�G�}(�|�_�RV8�S8Z;���'Y����&kɯa�O����^�e-z�x���6�?@��E�po ��ܢ���.2E�..T[��;����J�!!YVhd����h�RIf>��T��T$>�7{Iԗf'^1��7�`�1,�pD��ASm9�I��=�6�_S�~���o�iCTgQ� �ȴ�<w�)�d��jQ�s�vv���`U=i36�y�C6��n �5LT�9��7�{Y[-�`ƭ-g���nV�~%���H�}����!7�Dw�Ow��[6�![:�ØJ=����_��5x�{j�ڶm,�����!>�.��$�����:H6���#����(�gE��(�K��q�G�ﻎb�;��ѭ&�hD:�"�~xj�gu�qC����c�Q�g+!ۗ����_�U�?��>]z�3y��E)2���Fy�����Q�#��N}���5�j\�/�c�^�\���KԤ�WV�i���Rn^�xX��->~�8�������8^���TQ���х��J��Z�}�E�ا��\�8��oպ��)K9���Zм�!"���)q����y^�*b%�@�N޷�ߢpѾ5U�Ug� �f��A��C���we���G2����x�g��Wr������A!�	�X�hA^�`<�Б�EꢝF��=MMȃ�Xc�Mqj���?xIP`i¿�[�d�1M�q�N�����ӆ�'&�Ƀt�5�?:¨T�_u�|�V�XfR���/�S "|8��CJ�̱՞?��=�l�x����F��P����9C����p��a;Ȍ�/��'U�ȢI��{���ɀZq�[�j�
�L�p��Ѹ?��������X��Vh<Q.J�+\�t
�n�����K�Y'ƩzN-�Y�t�hv���w���J�_�l��Y�m+�I���f�%phzLDk��}�n���Q�F����E?Q�!�	��|{�Pw���0h:cCѓsu4��_�q�Mx������ܴ����?���{HS����`�E�њ!N���;�emTT�6$�~1���vr�i���ܦ� b]e!�)�S4+3�]Y��l�`X`p���E��( B���@�7�+�g�r�s|��:G=�ݖV�`�� YE���ʺI0�7�C�ѥ��D&�|�{,Έ�ם�+����|U��%��Rk���D�d��)��9�ĸ<��¹�j2TỨ}P�*v��nAm��?"�b9���T��*n�vL4����f�,"*	����X�t�_�����G����h�Z�C���r�i��~Y�r)򜊫t1���9��"|k�r*x��JO^�V��ŗ�����k8F���iF��n����"���U#q4�*�D
����-֭Ir�&؊�q"\c��NY�,�*�)Y��� �g�")�_��E?Wœ:�w}��Rn�ٶ��\�19e�5^�p������_�L:���f
��H��Ǥ�
���J���_�>G�H7�c��ݹ_�a����*��8�u�@�hc����fO\>XYOaMi��_�@c���Ҧ�$���S�6)Z�0����Z�WdbRV�t�J��@�j`�8�:)��<�2�}ʰ,��]��̈Vŧ�Z�DY��eLg�=<��qh��Y��Y�>5��!����u�P���KA��xc���O�F8����+�.����R���W:M�n�s�,���+��T�E�S�.�b��6��2o�jL�g%�}�|R�@)u��n�b�EN��5~w�=J$��k�>q-�	���{��h��m6}����En�߲�s\h^$c��k�iX0Q�?�A���^�W��{ 3�V����f�<^�˩#�v#FT��bj���\�1�����>|m�Շ�V��J"�`R�᫬�qP�4�\!���#?�-�5���[��b�O���b"\!��c{�n��?ص�3��N߁����]!�P��/	F|_�����(���x�O��9f�꒩��UQ\Έ�Α���ؘ'�eA�y'�о�\�}v@�gc��˔뫐6S%P���&	̦���M�2�x����H��Xkm�^[��$��"6�yV����~O�+1��S��I"x�`�]�:�Of8��]9����3�P�~���gb� �*{����PD�GMTL�)e�-����J]~b�5M�� S%��~�l�9�j�a[�-n�߶]�XK�6YFE ���'[X�09m�{	�G�ݟ��v5�P�|>v���?� ��*}��
�~(Ol�=�x�dQ���6�j����x�t
r�uG�n��B�L )�0r��M8�ssO���m�[����I�`��hp>=Xn���<W��BFP���Ǟ��n�h��B~I���C[r񮾋�)[��*�-9j��Q����Y-���Sp [�D���O���YXw�C�n�S��R�F����͹�Ek��w}Y��2�X������p_�,�e�h~�^��#����@�÷�jJ�ˊ�{�[�_oxʫ���H���t�T������n9mq0��m;��©���O�>�e�>��Ҕ*�G4��5����Ro���Q�8�O%�J��a9C2YⰗЁY��VRIlO�x�씀�{y���1�c�	���M���\�'F*&�7(��%w�:�����^5�;*`c�S;����w�
E��Q���L'�6��c��	���-���g�=F1Ƌg�9�؊�����&��^e&�I�F5��s����x��D�g��&�0ֶ܎��%�q"ڄ��:<q��l#���j
ċ~�p����7�V&��%G�d�H��)�N���=&�V<�yl_͈�h�f��˹�c�qO_���d1&tr�_���>��H ���n1�v��}T������]:#�+��jJ�� *��P5b*�f�fX��X�X��U�R�w�0��;TåOG�
� l����;ʂ���
s%���+.Su���>\|��=%?t��.<:|�R5̮��9l�WMb:d�qŮpI� �N�O��9�`�Ԅ:� ��
>`2��[���LδU�B�"7�-�J��-�?�G���`�V�/�����Y�˙��qu�o�m@��7�Л?ˤ3�7��u PZ3����+ -��ύC�:���-�T�s5�璒�)0rK�Ý;��^j�*>���r ��%툍(�.~�Z��>�6�1�tAz�/|��7�X7c���a�tg-KZ�l{oO?I[W��Sڒ�R�:F��Gd�^�)���3*�v`Ә֪����{��k������X������ϩd�O#�*��I�"(�A��!riN���=~�I\<��7�v֊j~�[�+�}��M���=� ڈ��)�ަ�f�zx�B"C��"�����~�Q�~�����D%��n�:�oB%1 �Yl����!n'P~�fۥg#(����	����݂}�C[?%ݛ7ܣъ<0n�(@�9��r,H[����$E�'������ee>��G��nY���K��sBp��un?/�� c/4�Y&�	>$=Rkr��S �&���85��%�=Zʒ�&�5��1Z1��Q����.Rpգ��n]�	B����TC�<Yr�j*\qAL)(�ދ�8S�2�rP�'i����1��L�}��v��Ό�D�~��+��Ȉo6��v��+Ӱ���Z�j�P8-����'���bW?���E-�w�G�������	��ہ�4���F��a��g&�񤑥���,X3����;��Or��������hR�E��Wr��K��"��ڕ�	8T�j�Xj��A�M����2p#�$P��`�侅�5`FE�k�3$7�<����'͸��Rluϐ���v���r��j��H}�m���;n5�C�[�U������@�<7���0�n9���Ӑ���%V$���Av�dbR�������R���������e�e8�mS�z^�^��P, ���J�v��S,��,b1�k�UJ�-~FE�1����)ײUU<9�s�6ҽ!¼ � ���p¼�c:�0������~��i�*E��R;R+8u�y'�bA0�H�� ���L��N�9�w������1�z���B}J�\�tAGQ��z����M�hݯ�z`�|���6WdZ��1�K���P�u�i����@U\:C���o(C�BCH�E򼽥��ǄB��~��4��2�E������v@����6���2qƧzj���^X���wZO>��gg�4)Z��t�,�<��M�>;�x�a$>C�O�Pe�]������x����S1]�8�Dc�j��e.�9g��d����(VmƎ��*��`�K���hVs䋕��T,��N�!�~kG�%�[��k��mƟ-ي�`g��b�W51`�
J0�)��I�z�8}3:r��^����C&(vC�+��f+��Ɨ���V����X�+:���_r��D�2x�|\Q��|��,	2@�4��������ꅮ$q����-�C? �]u,�}�-��j��]T���a�x����iǲ<xQ��ѥ�M��A�	�<���q��n�KG��}IP�Z��s��K���Y+4��
�	J��)�望H_w�g�w����!�� M�{)��`�+� ��3�����׌Ī\	%~XO�k�-�	����2�:f0�&�
w�!#�a���7��wt��ݻ=G�i!0�B�W�-���>��($0�Bn����M"I?�/�����bg?�Y5��?��b�?�k��������O�*��M�hntڤH�F�$D��Og7���5��d!��H-'�����/%��N0s���tU� �j����]SĿ�hk�^��bKa��4��{���%��x��(�
#�w�m-,����PP�mQ!�R�2X6V̊���>�f]�n�|��4֝k1̆濾���K�Cf��.�	)���l:���#0�9�I�ut�I�Ӓ��Z��}Uf���\�n4w �d��zP�\yz�[E��h�M��<1A�����T�Sǔd_��Ņ��f/juq���.�Q�u����"��˻Pqf�-$�&��R���&W��~�Z�ֵ�3����'4�2	7{�
,f6��]\~S�Wd(Ţ3bc�K~���y������Nd��������푇t÷���.�M�3M�h��g�����#�5�*8/2��
ؾ6���Mc�N�L��
�U�K���t
��3k��<���;�ۋΕ�ْߡ$����J��o̕Z#�7�V�/��K�ܫ֬�3��/,T�|���pB��e&�hQJ�����`�`	�b�OGˤ}�r���Z�U�iz��|wL�#v�����^�sRZXQ���`T���i����?]�9S=�v�ji�7P���	6c4����{�������rO��%��D����1vr
�*��@�U|^ ��:Qğ^a�@"����5���Se\��874�ʵ�[���R�cw`����թW5~�,�^�X�"��a�������� �׺�����֌�n���	Z���S��oU��<S;���5�cz'�I��-�(�f�3���]57hI�A@�4F0Z=��4�پ�o�!�es���Hn�|����w�OՀdY����3�������*ߤ��y�;=h�gl�%:鏠kS�g��Z#i�q�2��[�8�^:EƘ>�]m��j��h���nK�����g%��lb�0@���z�^�`*u@_�[�t�ȒT�������N"g�.Y�[B��Y���wz^�2R��%�̬�.�Q�i�t[Y!����D�����\��j��&�9<�$T��k(�@��9�<B,d�N�c0���#7pJ�a<ҁǝ`��~�]:J(��(�*��M�^�8*J�޾�\o!O�/XxNeC5��J����Gc�jN���C��.��5��#�'r�\7�t�	��%c�b��>s-��h7߷4��Bg���H�F�+L7r%E�U|��dd�<ۇ;�w�6-2�;�Rx1��n1'����R�Z����>N��́�Jt� 7L���QY����J�0�v��Ú����W��m�s�����꛿0�Nz�iԄ�7	�3�����EΏ?��+}��x����BjB~ݮ%�ދ�L��m���|΢�/J��	�;J���'���]��_6ыU�$9�$Ä������"�?&����f�.��T{�{:��O��L#��z1*q��8�V��@̉poc�4�1TRc������K����cN�DR؛�����9[,�xZu5������$Ĭ?5�S��i>�������bƈ*@m�|\���#�{���f���\��F��f�=JUTf�������7rȋGR��Q/
�1�／ayP���Ce{�4/c�L��ص6wO�EH?=j�B�nc�z@�LK�ҁ0��	;y`,�YlLŮ��JP�BKS���j�����ѡ����aB���O=\���B�D�2Q~�q��Y$���R���Frg�� ���K�X(��_�L�C�
�����)8|7�=��<5�b6�tepd'���5���u�^��Y��<����\�D�]�*i`���E�"����Z�9��-pd�6�T>���!�G�{*�i1�����"�6yQ��=AV;S<���!X�<��<���1���x�zs��C%K�-�򡕌�x�zOa��b�,lXhyR��
G�JB�g8�a}@'PN���;�����.v�"�,��bQ��z,s��4OaP��ǻ݅*
��N,u�W�8\*\���nW=��"y�nDq'9(R�۩�W^i��H��6�������A���0N~����w��O�]B4d���x����f�?ZY��@Sk�!�a3�4��~�|����6�{���*�$K��2����(������LdW��e�V:�b���uWY:k���IK�-�����L���m�nw�ķ/�SEIO���^04�˒�C��t�T�u�bA� �rƶ�"���z7_���ٹ��|�9@Կi >���#�t8R�F��]�o|λ�?k3e��ӭ�L��ii�F�A�7U���K�^�"�N�E�@�9�&X>�)Q�KS�{0��K�l��{
�FY7�w��O݁+�}���֌n�b29v�uW��U�Y��{�cr���M1���תUA�b����n�;���ėw��G�yj�쥧��Z�-O�'�iz����d{"��On ��Zd�����K/�=���4�0���;��-���`����w��k�/-\g�l���[=<���U���T�g��̕������j�}� �%m�������VQ�[�}c���OV9��\9��F��{����˛ei�K�V�Tc�o����o-ſY��*PB���m��|�#�;��o�պh�E1t	�
I
1������T�"��؇M�_����]u�G�4Z����|���G�H��[U$Р�C)e˹z���s�|d��P\[�U�b���`�Bc�k���nQ*�16���������(���ֆa�w ��/l���A����2�/���~����>��ص��(������S�ĝ�	+�Ψ|j�nxk��KA��P}���� 9�\�F����3�<��ҿ�l�:5 ��
)�U��ڬ0]�G�v�>V�!��F�~]��pv��s���I��x3��(��p�|��]9�䄝���y������ʯ#o�W��+�7#��%��2I�T�R!��˶���C�HW!�|D�)��侯�u���Qr]<��+f��C�m�-Tm�*[wDR	�����+O���/v�v��P��v,��V�Q;"x�^�X
�ǩ�3r��r�(��� ��V  �[��{�J�Z:A�!͜X,:�	NSJ��p~���"��F����;+~͌��y�n�WbZ���Nз���5Q�9j>�4EZ.K������f�YQ�V�)�F�H-�v�d���̩�<ϥ�
���¸�0y�����6-i)L��d���t���_�z���?�Nh�`�����IeZ�+�;�W�ԐO�X��ߝuN��F_��U�&���,X��LzK� (�����d!�l�@g;{��G��Ւ��~�s`�#=]<(��$z�}�����B]�`�j0��GS3QJ�U��]�ʡ��Z���no�=0tw��1���4�c�������z�����H�&��'�"+����ጒ�U4u�R����g9����V���d;��uןb�KB���O�'*�=�S�)��S�9�wg	P��݅rSA�K�j����Go�D&v�h0�\CJ`�������^��Q01㜗L��cv�b��0Zb��V��N�3<ȧQ'O�>Ķ#OZy�ƭ��3�0�9��+�<�o���k����QL+ڢ�r�l`�`λ,��i��M	҉��Z�!��Ɔ$�Ƈͮ�p�\2Q�_�V1�7�@�bqtR�	4��� P��9ǧ=�B53�I���w���rO��y��R��v��|�F�������-н���>�mW
<������vS-=��T���.�\���nĥT���F��6��՜PQ����� T�B�"%߽3�%}d��W�&m�r�P�qr`y��{������s��ϻ+)k��*���?d-RX5{8��	�g�8��z27IPn��M�lX`c4��+�il	��x��G��UX�w���0M�'n��a��LЃ�)�	b�V����hV"�� ��"���${ѲӒ	r3������4�ɅKާ!{�X� M\��	y�`(;��%\ ���ϵuD���bW����m��gi){����Pk�y�g�1�jXs�[Z�����+^+I�f��x_�D �%���à�%���@P���W�r��&HMXߙ^�;
��Y$y6��'sˮ�ͼ	 �EaH�@tұ������T�@ȳu7���p��ِbK�^(���S�poҸ�T�9])�^%�K fW7@D�k=o��kI��jz��ꚤ��� ��F1P]��o6��=��O�ST��y��0�R�U:��0���o���j�������B8ʔ�5А�@�<���N��*�f�l�L��"�������R�NR���TǗE:�ap.��["YC[���/��|��G)�.�s"5ຉ$h�Gq1��x���dnߐ� �Ӕ���?t����
��e��̥����E��,����1��ލ�7�WR[]�)�GTZ��X§��\�,aȮhk�]:��jb�ל���������j��aN���_�?Vw�e��|eV�x��ܯ�#0׮��=�xo������@8+�n�y�iap�#^QTᨰ$�~�q��F����6�Vہ�c�-�p����^I���T�֓S�����y��C�:�#G�Dn�7��-4j��e�]�3�0A���LEH�UTm
77�9Z��b�G^۰�<�s�@5Z�I`�`Щ/Y��G-� əN^�D�;���HwOYvC�9qπM}
c7�.���y����[�f[ w��h�+�ti�EDOlx-gWa:ٸ�g��:���\FO:���K*ʕz
I��ft�襦��u�'�P�*�I�π#�QO'��J�K���̒s6v���GO��_C�����#��_ٔЮ��S�!�$H*�Ki՟�O�mqK�=v9�/����������~�dwA���D���.C�Y}������.��%}�ǔ]�ⴘ�}>�$���X�t�o0q�5�&�����ʗ��Y���/�9��G��p�c�-f�_���]X�0��e�5���f����,�*kU�C�^%�1�fmƥw���;Z����(jǿ�,j�G�}Uw�JP-N'�Ẑ~��N��Р e�ü>̞�n!�PiU,:S�O�'&���Ԥ�\�&J0t9<M0�;������Tz���y*ܲ���������'_��~>{�Ne�Cl��b��DV�c:���_,����W��[_��
G��ZP�����-(�|MST,��*~���l��X:L��k�s��%ȭ�F�eQ6`�]'Fң��s�[��X<Qvt�㖚ߤ�K1}2$�_pv�H��R�+׉����Rf�Iq�̺��v	��JV������c֨Sĕ� �c=�_��eOu���U����n(�q�s]%��%��#�j�Xw�F9pAv Uښ�J '��e���y�@���c��C�e`Z�-)+GR,����;��0��`��͂aH�� �xj36����F5t2�1�Ʒg����c�z�n��;E�=�9�[��-��4�`uӖ�>�V6�o��ħAF�ƛ!f�,����\Ns��a'�0�N���*��G,B!bI���i��@aʋ��
�,/`޹�e��y�$�� 7�?Uy�����3��� T ��G,B!bI���i��@5�wq#���0O�s6)t��NI���j2��$-5�)�O5P(w�c��a�M-3va�H`�\�n�J۷v��O���]���W]����P��i�L1��LjD��S.V�lŒ�h�������=@:Qx�v@�>z���ٮ�$_�Փ�Z����U�^#��deN`�VF30&Yٵ��.:�t�$�AθM��W7״%1�)~z�>y������jƏ�2DN�>!����1�����2b&�cW9)�Ծ,ЬM�.��7q-}��gt�v�f�������}j�/75�������&f*���|�vfW�E�<=$T���h��A5�̘��� 2
�1\Z�#���t�ο��l`����Χ\ �_�*$!�E�1(��fM��ļ�:���?�=U������9�oeX����Z��H�.�Hܾ�Abbx���� qݞ<�YNEd&G��Ŋ�R�*���r#���,-�i��Y�H5(LW@�0�u}h�9��-�.)�r�m���}��=e}֏�8'�p?��l#e��0�e��>�͏[��=�Cx� �2l��?%�����t���Q�v⭵�7oe���g��+ҡd"�|��-����s�`�r�V��fQV��4z)*)�hm�W����UY�_�r�X�X�^�@R����!��zG3�-VhnP��U����J6Ubh����7}�[R/W�q*ŀ�7ގ{s�=9��A�r�������+�t��0�+O�q%ɘ�Q�)�M��@1s�0�`6؏�Ay�%�����x�OZ����j>Wf(>�M�w�:�7nt�U�&�x�[y��3it�8\��������|�����i(���o�M�����L��f�K�T�nK|���oH���B���;�Y��R�G�w{=��	c������i(���o�M��U~&�����+QƠ�d�!���� �/��j�h��i����ݹ�c�a)��N�����o�Ղ�j�M���7a#M�
�093���6mtv0`9�_��P�Y���Za+��9��H�m��R��r7�Ҡ.]�@GA=Uf�AO"�O� �Po��g#sΤ�b^��u�C�2��l<��I`����ǀ������ʖ
 ����^��������w��^|j�a�.0�V�H����6m��g���{"	c2:ueX�L�ژ�ܵ-\�����;���Wt��O��2ӡ(������݃�<����$�-����G�O��-/z��Qˮ=�z^jy{�,�>>�vLB�w�5_8��^��һv��p��c�f�0a�V�޸+��������0�;x=Z��T� �����f��Nw0��w��ƃ���Nͮ���w��I�=�a�:��亼Ej�~�HT~��&�L̶��ꛉ\@���Ӝ��!�?�<\L�y@j��ıs�69���/"�A%�N8���7�?�Չ��'���߲��g?����k��4�g�Ȇ��b��6N�o	F�ʦ�5i��8�v��
dЌ?P�% �@ã!��𚖲ޘ�klY��q� ���J�%pa&�7l��3i.�I�p�4M�Τ�j�t&�MĮ
3DuJ�3�8�{˂=(��i؏�	dxq{+t�@wq�X���]y:�ڹ�����S�SR�6�a�K�^3��^$���-�bt�i4�G3Wه���	y �5��q��۾�o�,ߔa�缝<�J�J;���86�����A���Վ5�1�/��}92R�iW��
��祚ȿ31�vOvM�X9 D^%8C�>~0�� �����"��@t���,"n�7�GQ�� �5PN���ھ����;4���5��'�Z�n��`̓��Z���5����v��j:!ظ)v���8=�:S��yx{�N�ǯh�E��_�9 Ŷն#�@v4�]+J4gԥ��,��P�R�Z�T�T`
U��Ft.m�+��0��ц����S$��^?]u�e�b�iň�%C�I�N��"{�(��![{t�B,�^++�g����g��\�T�$�iY���)̺�-Pt免ʎ9��+���!K�� c�~<�V=�M^�ԸE��ka���?�n���Ŋ���?ю�r|/u��5p���ġ��7]JW���E0�B���n������
o��'*t(m+d;���5�:���cQ��Q:�Tk�[%��Џu<P�����<w"����E�pe�V�efen*|K��->%�V��`<���Xtj�g��Hw�Ox���(l���k2�f�k?�} +�3�L�_�nT箹�|H<�A�2�����W��o����\D��D�U��C��GeX�?��]h!�,��)y��*pAG��^�� 5�j�`9��z�}�|
d��o�ř�bǪ0|?=;�KL��s�~څJ`b0�I�ai�L�2�.7eA0Qj:,�6�I0�QxѤ�_Nj!�%u+A�O�^g��5^
���8Eۇ�/��j±h���~P�� ��=$b֮@pi��Y�e�)�/����X�=qS��D-'Zn�����gs���3Ku���HirY�E6���[@�������،hf��6�?����� ��<�`~?V����pB�� ����7o��ȇV���}��L�@u�B�E���L����_8�tm����3`��*�IJ��	�Y:�z�:�&�w����/����B#鉝�^����>����
AfJ
U�\��g�������D��	���\x�u�j��b�Ac�:Q}Jgh�C��{9�����\��G��������Z;���]U�m`YXACn��P%xX�-�d�v� �������㱇�m3��R���826��l6��~"�
��G�b䭈�h-�x�����ɬ(�e��p� E�(&I�	.��N{��i�c3�I�kZ�*o���2,HHy�H�L�=�z��(]��'"�6�q�Sp�W����L�a�2�Hs�a2���J7x��\����b58r��H���gK�.��oW�����e��F����k�$���b�Fd���p�O��Qmx�|�'
yӃ�ue����>*敉��W�n�M=!��Fci�9�����'[D�5<����k�ȂP�|L�v��
�n��V�C�[���w�ԭA�X�S�f��^���e��$�4����tޑ��*�q�ɯ�z{�BFX������lF.�%�*ߵ�)�v��59 Շ��bC ��rBT�2������V��z�˝e`�\��2��&����������p%p�U�	�:�x���3n���'�z���
Z���]*���։> ��f8&�K F ��%%;MLݾ��.�:0�5Y������lN��We�ZJ���il��Q����Q�e�×ش�����4~��]���((_�1�0�Vv� Z�~����y�i@�^{�9���e&P}r�b{��u9���z�/,�m#@��`_�g��sX�"�R	i�:�8��֎G�UH���g��z��9���)�^Q��5�>�L�Mu�u,Hks�}٧d�-��>΃�y���X�k� yۦ8���֢8}�f��B�[��;�
�\׽z��͝:�5[�>%"��;W�����M߭*"KG²Ax�E���|~�F�Xo|�x�#��Ĵ ��X�r.�0r�jx�Kl8�Z����|�b���Q����9]���%�����U���������A��<�N�"?88��l.!v����M%P"Yk1�:�q��~˶d����x�:�/��-$�����\b %(����n��à�ޭ:$�4@l7�)���,��.�*f��B�2�.�ª����֙(�������"�;�j��|�4!;7#z{1I�ǭ�t�2o�g �����U��o�����编a�1�-G>�eyn��]LϬ���u�<'یa��z{��.�.�����Nr�Hƀ��=E�!�:{ �e&��4�D���G� !>���g9\��>!�੟My��e�310|���x+D �ܠ[��>�53��m��)5-&�ɷҸ�W�n��\�O*l��;���'�a{L/����߲���%ϼ��??�^Xg0(���b�>��R���R5�VQU�1�&h��r���l�}n+Z�S�v�V� ��7��A�{51�0&�e��6[ı$����d���H`��b`]��A��4��M3�~R��'Y�Dmlr�dp��4��z$�a���x{>����@�������03ml�Lm�i�m�O���zlRo���7G2�٘i>o���H�G�'w��	d������r}��Ƌ��M�p�,�J�ʷ�&����ڮo��&�U|�lDT��c����7�a7Z!x,�C�~,к�V]R��قM���\|!ٻ��pM�@��:����� '��F]�/��Ht~�?�?��yO���
�=�Qe�gte�,r�n�9NgU1H+
��!t$Dl!�y�{(}k�(���@p�-VVc�:�}=<B�#��^���#�*����w���D�/����m�V� �d���B�h�4��d� $��4�^����}�
�:H�ٙ�����e*b��������H�Rx"�FO Ǒ
7���huRϵ�g��4�1�ˆ��:}1+y��]��-u�����h���"3F�u#�Swc�*d�M��8u��a��L�����
o崒�6a=�L��~�|k��=9iu���s����0�|��o���n�֡"��Ԥ��og��r[F+(�J?R�������U�翦9��F�a�����l����Q����r$��?1���)�&����0T�=�C���pg�[�(X=�m��۝���깋�MPCB*zMxԘ�{��Րv��fԂ��7t�Ru���Z
�{?Y������8���)�
Cj<@*)�9��}t�T��(�~�h�۰���s��1'xf��>V����A9M��($�)P�iZד�Ӵxod����v�+�[��P{�����%�
8�����܉�����W�:�bf+�F�Ħ�C#2�#Y]�F�I�`!�'�X�<�+�,}Q�-��ǵ�n���*W5���#;�S�D��:��̑\"�;�[�R�Pc С/���>���J��Ȋ!�:.�rW~D�^�ܺ?_�eI�})�58��f7�!�"k��/gmgC<�1��"�wcN�Ҏ����CWy��/q��hM�b���	�L�Y\HR��mINJ������#�CNG�Ւms�)���i��Ā=�;?��N�-/$�ƌ�֊�fR]\'��W 	b�r�;j���BOX������L��;50]*o?7�'��%o�:��!����L7���#���w�NQ�x�ť)x���m�3y��J����\�ۥW�L�|�q�_�bZtnnY"��q��a� q�c.��� G��NP,ҫ���0�C"���0��7�̘�&bE2��ŔP��>{�Ip��c�fAp/o��3�0�6s!����d�:�UC]�lAJt�!�p�Tt��+ܮ1��ա����|��r��^�'y y���50�zM��z��R���]@���;&cfʊ��Q�+#ߦ�ҁb�ݮV|Q%����`U��^��P����A �/M4�goǻK�-v���s~6H�y�2I9@��z8Ԓ�.�c�����u=mr,h�1�~�Z-�v�"��J.��S����ò~:�/'cait;"����,�P�p�/2���5�ͮk�+��2vK���?[B�}�F���3K���R,+l�8��e��[�,M�KD;���Q����'���r�4ƹKl�w�U�/֕���l�]�[2zeu��4��4֠b
<En������YD;�Yk�[����J�:�����@6u�v��N�\L���@���FF�_��5tӦr����m�|cv��o<���C߹H�1Ug"d��	�7;��/[��"�6�;��f�Ѧ��#����z�C즐�{԰���O/�@Ÿ�F��!�Z2���/����-�K�����+꣣� |Zخ�0_!��))7y��؟k]o��ڌ4E��n����7�:�X���FӦ�e�STʐ��B��4�G�z��@�w]L�i�%|��������XFqk���0�c%L�Й ~����nW2XG��?3SbKi�i�ZE����	��W��Es56�k���7@{���~�ͮ!�e~�&��5�X�!�A�	��Ld(���)!󷝌�@J|{�8�)3�{�`ާ�����V�h7au*��ϟ�7[��Xc/�A�!T�:WB-c�T7�p���v�7��	&��y�iwCMLŘ���>g�cO�
'lUM_�s���P���9p�G�4�;����hp�(�5��P\;u�?�rwigW��:=t�M4��è��I��jh���.��4F�r�+��<Чsڜ��Gy%7�̰�&�I�&]��(#'��?uFѕ���zuҲ��������1�XJ�8c�vUJ�ݎLb�$�Dy�<�$��/>��4�o���8E�z��` ���Ǆk�ǲD���-����i�"ց��*�43eƨ���s���~��r��Z�/��]9-P=S�ʒ�!y��d Ry��u-�S��~%� f��I}H��hn)�����Fց�tclk�/f1����4�{�;�O�yd��u������ɲF�E�]�J^�hd�T5S}�2Gێ��ꦟ��ae�����ʛfJ}�'<`��dڊz��q�E��d(g���)�ü�&�˰K.^VHt����-U�{�^�� X���k�Z�VC��ة�9�� TKԪ���t��CȑإV�#]�,���3w��^�܃��$���N���:��k��7���%_��|0��<�ا���c��,���?�P�`s�[�v���8G���#8�ǰ�:��q�X�(,�[V�Frh�����d>�Ѿp���rg�a��5�.Rt���,�b����Z�
�� '�e���{�������5><���{^xJ��b͑��~S�J��>h
u��;��4��p��q���9hJ���H0��s���O��l�h�@Y�H�S[�Z<>���-���1_��7V�ѭΐ;:m�,��鯢x�ZP&H�|�j�<|7x�?�������"�����`_�xϲ��2XR����,Q��ϥٵ�=##nv�[�R��N�^���u/�m ���±~����y����ʲ�%p~1{��6	�
�[��\�vq�2��s2�*Xرٙ^�T8%�X3��:)�ɓ�c3�V�l�Y'2z�NI }+�Z.��.GVu�aYt����T�|���%U����!Ǣ�a*����]"�����O�p���P3�-�Z�O9Z����f�����)m���9��m]&)4��ע�� =����ڰQ��:?�u�k���7jS[���y�EM;mӑ��
|w~���s�����lU
!��"֋;5��f�}Tָ��@�K�Փ�Gg&A�t�КܪѼEa��u�y�:p�[�(��l������
���(��k"��ּ�ל�k��t��}�{���Zq������p�{� �J5���[��}���q�З��I�]��4��K\�Y46ׯ�g��E�L�=m��~4����e1u��_��w T43�Tc��W��7����	+�wfJM╝w#��F�3�u�����76�|��l���L�k�0��**�Wxn����}�I��[��F�K]q8���Y�0A�\�^���zlxw�A�C�H��)��Y��+�i�'S���?u�;�mv�c�'41�革���S��X���0��X;n��9���s�b2Y��a��_�"���)�=�ߵj_b
>�u4�n�@�&g.Ʋ'�ᳶ��h�'�S ���͢cO��Qq��u`�x����u�2�ٺ�����+��<�R��9���F�ϛH #Zq��`v!b�0"�#��m���������2ָ�GM�C��k�`Cd�p�m��W��ٜm1̜#���q9b��Nyz&��_�鵟�|�X(;���i����)�NX�S�V�)l��(@`j@�`�AS�7	��c����Xa�� w��GE�v$���pTb~.T��T�Sdէ�|�%���۸t��hJ�	�c�՜��V/�<><�4�6kTBй�f$��X�/�R0a��*vPN5@�$�~�� ���Y����7b/ٺ+�zm2GQ^���h]�6CPNc8��+��M��n��ԓ,�ʼ��{��'(?��R�����'bԇu33�@P�����4�c-ǫ́aOҌowO�i����0Vwё��$o҉-'.i�e��/�ճHF�n>-3#.��.����5�8� ���Vx�G4��e�� U�Pklt�����J���l��H��c:��^B��,;$������vR�6�F2V�C�ˁ+�H���٧�]=� �{�B�x�űN��?���ڭ��]��/��._Ҳ3#��_+.��AK:<gH�㹭)�x�&��m$��+!K���=��Y�!&nW�!WU�
gZ�"�Ul�	�rU����)�#J*5[�-����SM�RG\7��h\�Da�T[�����Ӹ.~�*��ۺ>PL����H���ZI��<)G�'��\�Q]�{�:�1�q��bc&��B�(t*���XV'���rG݆j��q��$*،U��L�MU�5���نj ~�>�Hu���[�i�~\�4�^�`�3S��"h�P�+3G1�Z))<qH�sTyRO�y��"_O��qMd�G��o'�1?�|���e�8��E2M~w���ŨaW��[y�6�ϦB/	���L�KRJ�-��	�yDP6P�!;����!�������|�/eq��d�bt�nlJ���x��D'���tֻ�:#�^�n���k�-����Dz^��.�((^�f�0���_G؃��m[���J��q����s=�}E��4�o��O�(B�k��sMI�3��N�׼8`�2L��-'�������e�W_ s�S�C���w��R��JV�R�J�;dr��|S�c�!�:Ŏ�R���Ca��3����R򁡎�[�v�tn���Y��ŕN���{�t2q�Y�~�s��̔��&b��L��{�(��^�@ʧ*�07
h%�8�<U��a��϶�� 2�dZ��CE$�k|l#s��×}.���C�H��5�^��b�}��;�uT̀����##��e�z���>	���0G�QL ����7�t��i�1��,X�G��{�e|h
m g� k��2�Ҧ����C�4ڔ�Qj�7ȑ��|�����}-�1��Ps���%���̀v�O�q�"�)�D��1�<g!J*�l��+s�L����8�rJ��^���I�X�7�J�.Ǧ����H��Ⓨb���f�[;u�䆵ދb�U�N�O�vK�?{��E
�|������4.k�q����n�&RfI��Lݪ腪�ޙ�%e-ɌH�Q6�r�9��˵^�P�g'���x���H�D{�C�7�����s)7k�=uI�$���'݅���0$"��Io4s�[޳�6��dbz�yz����`�z�D7�3���pH��$����Ht��%��HC>e�}nJ���~h�f:�M0�(���Oq�ug��eT�+�꟬C;��`I��&Y�-P^o��k���I�.�"X�\Ic�b��<Oک}�T�������r�[~�"^�~��@������sRD����z�&�s
��J�H9�M��|>��������IA|@?;P�e�)�e���ZA ��u?8�X�O�*� �F~Q^]}���o�'����*�P�f��[��"�~jLG��!����ͱ=EimQ��a�����.�(s*�ޮ�"�6�^J{�����qP���M�3>`�}�p��y�)S0����v��� /��gX�`p�A
��R�KZ3��aA�.�3�,n-�����,G/�:��+���|2�_���s�$ykQ���=�?%gV%(�b�&`C��|/���<��U�p��O�,�ʤ+�5N���g~I<��	����(0���!O���Y��7�'$u�p f��iI���K\0���zQw?���W��,�e=0I�������<Ӿ/�o�^�Ȗ� 4.�^�:���8&����;i
b��S��T�1x��$mz�'���?�,l�o��ɠ�1���Q+E�_ف3-�R3�X5����1ϱo��1�Y���J!Ŵd���´�ƿ�8N������u-��ג�P"yǝ�قp	k��.ފ6fUn�C ��v�B�V։��	kH�ο� �8�Uv\`@z����nQH��o��+2:BL��ތ03?l]�%���Um���L�	�L�6�8�x�e�O�A�T�?\z�TuӒ���ζ$EŅ��v:��I's��w�%��[���&�  Q�HI`?+r1h㜈�����y�7�9���^��{;*V�(�*�:j�3�Q��N%  ;��nW3%��u�<}Rsȗ�G\i#�t8N�PfW344tH�7�p��P��x@Usa$�k�X2��r4��=
<�(Ήv�BN0�a$�yw�d�ls��&7����J��~=��M�Y|X���ޏF���qqp���x���5��:�2ri��[��}��Lj�e�'�.�Kk������)p����2T�y]�e��n*����OC�c��P�9TY�M���8�/�BhG�v|����^��[gq�k�R�=�ۭ� �.ӅA�H�A�+��D7F��
��1�]�R!���؀"� ��*:�lrn%������d��)@�)��C�jt(7�i�a�L�1D����D���Y�7aU���$2|ޟ�B1�'��n-M���9ux���y��R��~;�G��|���X�곅�����*��~��ǉc�ܭ�|�b~�{�։S�k3E"8����xH#���a�*���y��J�~j֗�*���8G�_HeH.�ܧ(Ex�X���@�?�4��,L*r���+�t���.����+jC��T�2���),	, ��CA�����qI%26�.��p;�6eӒ`���_����} a�l�ΗR��1ZY�\�yz��XX��dV+UO0�_���zv�2ۘVb��;�_������3��=��ܒ�
�d��Ú���Dx��pϿ�-f�l������J�j|��T\��xW�m9���#��*�2���0��_�3�����C�Q�-�1�����Đ�ab";�/<ۇ�&�z&����@[�)@/F%_��w$�]@yz0X�On��TI�� |0��v��\�22���ec�H�o�������=�T���c��a�ܷ�$
F���َV��?Ŕ�2l*<v�_�+�U7sV���a��z4��v[�8h�����_f?�����Cn��M���(83H�
?�1�VЅ+��\��Xw]|-���Ǆ�o����o�Z���\D�m��&&-:w�Ѱ8K���i�PZm�B`.��Z�-޷�z>z��	��{�Ie��^݄t�F�̂&< u.h"p��I�ʒ����r�DaD����э�J
�/G�h���gt`�i�)0yÙ�� �EɆ��(A*j-��ʽCD3*4�7�$�:v���b�ŭ3��{��<eܟ>��i�pi��,��߬�MjH��eߤ��)[��o�\�=�`��	���v����9z-��������SL�)����ts������C��^�UU#U��ho�"����RJԡX�� �����s�9Z�B4�P&^+�Y���'����8���M@�6�s/)C[��&XI"*��=0�$k��vA����)�YS��C�;�W�wpoTkR��en�"���-��&�b�Y�� ��xHi�M����Xe�L���z�?Q�?;��b?|����s�ɵ�rP�!�
�����Н��_@�E�kF<���N�QW!��b�#[�h�,b&0KJ|�D������������mL�1��o �i��q�(�In�l�0��t,۶.�J�G�
��o=��6�Y��f^�j���I�.]jVs�����R=�	͚g&kA	���t�g�j9���
�n�^������o�����5������i]�a����Z�,$+D����� �F�>c	D)���'�c�j�D%*5�(�1�
�8���p-m�����Ǖ;�H���k�J��#`#�F�JN[)�.���?�c��ug8���ˀRT��.�l��o��#p�W����0�th���:Q�����/$s�):�xiF;�҄g[N�9\��� ){-��;�_20�A�W��H�P˲�8A���y����@5��Yϰ��>rA��r[���d��o�7��X1�j���Zy�̊�Y?T���"�W!-}���M3�Ư�[�D��l�_�YL�	��Ć/�ԪtD/U���&�W(�:����������`� ��,�u�n�%���6]���*B#�8E��h�pg�J��֩�)�nX�'��.>���9z�/���$�d�{��Zi�3t8w�'ԥ���Xw4����N���u3�/;�\����AY�K������k^�JL�2�����L��J�����'����y~QէX�/�*�.վp�1Kz�y����G�C�c8�t�����[$ʪ��g�_�2�_���G�x��G8�`r���H#���sß$n��@�A@H�0��Z�S�?��JS�c$���YX��Ș�j���i��?�x��"��<G����e ���s3�iG�R˝�����<��v�x�fY9���� ��e���-d�E,)/'��|�C�\V����?O�u�.�`ѡm-��;D92�}n���j���|�%+�b��Ԯ=�K^�����P%\	�=��kU�����๪=��Y�R�6�U�?���݋<�~T��'0���?�zy	��pp�vVObb����f�;�\�� Z�NI|OǠ�^�$�S(�}���]�:�Ǵ��?f�$q:�r��*����qAM��)��{od��[1+h<4��iG�-����7��6jf�c��r���CY��#PX_u;�2�|�-W�D�k����*̎�C��k�cXl�l�d=x#*BK`�U Ϲn��Ș*�(Ok�^����y\�]{�xw-��>�L�Hz��BiY0?��s{�V����f[�����)^�"�@^��ߛ� >������nbP�hƓ����$2�~t�9H-);�Hgz�w���U�T���1 {�D�{ �dw�����:@s��3���Z�x{�k�I�YoTlI^H���ܱ���BƄ���1�|�}����\���c�U������]��i��i���1� �=l��&��q�?��p��q�/n8���4ɹ���%�����0�#ۜn�_�h��sEOwڵɑ��+�^��Yd�E�|`-�FG�^�.yf��~�Z����P��!׀A�"�=���1�[�ۆb���GY�z6T��UYj�U�iz�}ձ�����C����c�bT]"�>�vO��m"L,���<�UlQ��9m8������~"Jp;���E�jL�o�1���'w?U���W���z��N�Yt���c�;�T�_(7����Z4Ėʗ5�>D���$�[�?���sGοG&�=C5|6����)h6S���͇uײ�� A�0t�D�S�8���������ݼ��'�wW�'�����U+�����/�i�ĩ�5R�Kwl���S��u��qi��g��ē����ޥ,_G�*�D"��.i���6���u��A�*"���O3򞄫g!Vb\0Sme��s�(����x�j��S<��1:+/1F��w��]DXnĨ��&��o�j쉭b�c2_!(�z�<�
;����Z�-��/V(��d]T�_�h�|BH�Dܟ+��W�����x����<��W]���G�-��sN/k�������f��c��+����t�<�������nڹȒ�EM��&��]�*V�25�	��foc&&�u���`Ұ�:t8����ߩ>+��ߚ�m�zj���^e�q���%�h(�
�#��z�L�;w�4���ABJE}����&�s=<�Y�I<�� I�r��s;�=#�H�rhU��p۬���!���^�DlCky����ͅCD<� ���.<t ���(@��r��ӭ����r.zv]����|J2��-���d�NR\�)^D����go�e4�%:er��VS��������cu"�I��i �6�M�՘l�'�3������f0��K�1��OԤ�.���Q\.�r�	7�� 9�y}P4ݷ��:O�7~�#�r��dO�����>àR�ø]u����we��Q�Z��p�՘w|�-r�X!�s\5�@�v��'��]|��U����0QHw��zaK���2� ,hn���ג�B��NΉ��idA�1���sO��&
�9�&P����fb\��(*N`���Q"������`'�N_h���I�'B\�{z�Kq�]ޠ����|�ǣ���Yz�h˯������f�^_�ڏ�g�1��@�;&F����_�#�0�宒U��<�,��b*cY��DO{j%�^���&�u��S�f�#i	�@7 �e��1
����� ���ؔۄ���IٚE����^νO6�OYF��*�i�l�;垣.>Z��K�L��ҷs����(����J���Z���5Ǯ���T�t�uY-�65�sʫ����h"��t��ϩu�4�͕6�FY�~3Y~�L���lZ���|���V#yžB�����Ϗ
�[����x$�(��Wj�E�*{�=u���HsyN�˞��m�{�q�Qvh�b{�0i�F�+� �sf`���Ť�
�\�a�d��4_�{DcM����C�Z�@K�W w;�x�4����p��<���s���j�?��X�"dmB��3�Ӓ!ц$��A�����R��确pb�Jd�[��<p�����I2��R/�:���9+L�p�g�"ߨ�CZC	z^�!��@�%�g���xX)��G�t9]�L�jo*ڸXVL��wB�8�L�ϗ�Ш������I�&��Ɇ�~�s��iC�kɢַW'�E�ڇ��j��+,��L�PsD�{��M�	.iaڱ�6���Z��_��
x��#��<��7D�-��s��FQzKG�$���c�]��^sa�s�8C8�*j@x��~`��K���Cg)	Ƚԁ��᫣��عD�2�]q ��~����`2�1A0I���pn/��`�x�y\�SǄ/nQ�o��@0�$�=,A.#�������O�R��CGH_��'��*L���`��;Q��#�iq���+(�J?�5Y9cRJ���0���ca+B�2%o�����d���oqL��hHN���+��:R�U޲OI	Ch�rpM�x�4�HCL@�l�l�|�S� �__e/4�Z���:	�#8�2\�=���W� kÛ	�u.�%(L�cx�kY�9Es�D]9�4[��`��`��z"�c/���ˬX�i�N΅�w���/�/;�.�s@	 #�J�����h�`�V�\	}
�_�D�6; 2[ �\(�p�T�ыN�&��@J�R^��K�`�q�^F��������RC�3��"i��2X�b>X��'���t4\Yq�S51�.����Sy>��}����b�$F����WX���ֶJ:�Kk�L����k��"-���P�w>!mA��������K{J�g�CtHh��+��A.��*�%� ������8~�N�D0Uz���Yd�ѻ���6X�w��
��+��i��X���fP���X�;��",�7f��,L�M��F��*��e�3^t0\8x�]1oG-���\��#[��Q����)cЋ�2bb]��Z�)��I�΅�5K��B��/"��5�;;�rFi7ڡk\��?���~�*�����`�p3Y��$fң>������ [��vM%�vw�sc���׽uQ��f��JZ��̿1�1�w�=q8%�3�0(�iVT���}(��Өxg����R��@�t:h��z�"�p?k�n��ٺ�R.Tm�����䨩�W�p��9�����	�F����Б׮S��e*�z�0"���^����N�@��F�����ȧ_��� ��(��Z���4� ���q�>xk�d�_QN3։#¤K/��v�Cw^d;�ea��]?ø�-{�姧BN��%/�P�[�y��ħ��n(a��_9�w'S���G$Y/kصyע��uc�>��v_����]���M;n½����}�B�7�R��v��dl�0i�H����r*a�'T�޺B?�ָFh����S��������ʴ�zJ柕.C�<м��$��O�6n��"L�u*��ca����E+���a�P�
�,�W�2G������㛉�b����ikLlf4*������UM:�'S��!!�82cBM�?KF ����"�c�it�o���e����A��j�:�Ҵ?[�Q��t��Q��H�D���+���A�UD���$H������\��R�ý�ܢR�z�Uiͫ����u�zwzT:�ޤ(�ؘDg(GE>96t�CB�*��Qo��;��ē��p��3z{��,3jA:��!ւeU��Sy��D���^�Rj�;�Շ3�O��~/�x	���XD����X��"<n�3�c�eM�8{ 7E���o�#�^��"ܑC����F�o^�G�:ҍ-ĳ�iT��K��ܰ�^n@�7q��b�-+eo�-�Qչ��/fd����"���ҵ@��Pˣn��{.���Xʛ������H�,�P���9v���;ʽ�V�*� �%���3mi~��x$yVy��T�ҙ�>�!��W���׮�K,�c�sZ����#���E�gO�7��J����~�d�����*
��O���M���;�
�����3��uY�}s����eܻ*Y���mPuDރ��i�*�4��C�V�P�V�A�Zt'�]���=��r�}si����:��6n���s0[1�TRcC�p�����j���g1�����ȭ7�;�Xu��½�z�N����ܱ�Ђ�����`��<�%=���zF�L��yD]������ݤ����X{�`-�tNɰ7�V���kao�_j��T.��s=j8�,��w��b�<��߶OI����8��{�FC�!��J�K�Z���K�gB�}���G[�o�O��� a��M��@��b�K��}h&p�D��('�%o
�1¶���/�*>9;M�R�	��;�ϯb�<*��w��$J \/����!<'��s��ˠ�CN�ͻ ��L�H�-"���"�V7��%G�������wQ�q�L@��R4y� �N? ?�MLQ���0��)����3S���w~8�%��&��+��|����)�Ѡ|�]�\�)Mp�1�N�SL��g�w�J��F*�E���h�|��F��P{2���R�]rl�Y�Ώr�p �&�%�B)X���ӌ\���b��p�Nlg@O���jt�����QT���N�6�oh�����d�X'�U\��ū�����| Zɿ_�S���Sq����g�
{w3j嗟�A�J�;��֒�'��@\�d�G�?��/�:StcЉ߈o�4Y��~� �̆� �A�˶��x�k��?�ŮYm ��ND���«��TU]�XȦ���9*E� �O�s�SV�F{Ze�zTD�,�� ��'�+P"��M4�Dʁ]N/�߫k �z�f����Zp2Tx�{M�ֵ�tTb?ɡH%3h3��p�z	�T���6���z�.��3�
q9����=���'��:�ʌ"��� �V�;�Y4�q��QY��p�4�9xq��ǕNSF����-��*T�KR3i��\S��Ә�������:�HF��B�g�� � �E�Rf��B5�6��$��1>YF�
u�P	� ������w~��϶Z���C�5�� ?V7�/x:t�$����߶�A��h�����J��h^qo�}�I�#�"˫4׵�3��Ͱ���i�[a�P<�>,x�;��)�=����:�A���6ͲS�3�����k�, ��W�g�m��+a��e;Jl�����.�4��ˡi$��:FJ%Y?���ud9Y��{��������"k�Ѳ9��Cx&He����Ļ�#�P�է����^J�2h$߶�������s6�{n�F�ѱ�k��4
���i������w�	�W8���[��:��B3�K�������U�ӶoO���ŕ����9Ɇ6�!�f�oSƍr�mmWG[E��k&ĈDc	I��L� �#I�k}@���b�k:;�a����r��j�$Ʒ�:��5<��i	�~�|+h(��?�������@A+��)7;�s:�\�{)�,����AA��X��q27t�1F���*Ʋt��#c��V���E�)�F�Vỏ�"�.JB1DH�<0���;e���uT�����PJS�\�
�މE��7w��ߚ�f�d����v�J^V�<� �5;9'�V3g��4�F*R/A)���IнR���X�d����2ZP�,u)�w(�gS�e��10���""��M��h�τ���E���m�LHq�ب������p�_�z.
��-�n!]xf�f?��B�%�a؛���-[D
�K/' j"�*x5p��Ү,�3�r_��Yb*���7�"���r����z���R�;`���:@ pT(:_�^:�����jP�!1%D� ��w ��C��"=Is*Wn��瑠)�\_�'�k�o�ic���qp�[�/'�s�rU�����8|�27��3��7�"|�O����gL.F����ll���ч��\��1��7ٛ��.a����t���(`ݚ�:�}�K����}I�.���gNT�H�Z�+������[%���Z�$Gt��1���%�2BZ� �9����c��7�G���=�~f�e�&���1�F��p��=B�m)���e��2������)j.�zNhE�{��<U����AG!�v��b���:�e���h��R�(��GrCÊ� �Q���u]������� @N,�a�����7Te�K��9_M>�}���W4�i%��=����z��Pw9���:"��|:��]��0r��xQ3�� �D�_}^2`�(���;���&��?s��}-�c�ĵ���-����f�2���E1�Gg0Wv���K+1KH�~�c��)�o�nZ�n*\�{7�x�I%��w��:����4PM̹o79Uɡ(C�A��S=�0�>�wKR"TĀ�kGM��g�VQK�f��1B�)|�X���$���+�B���x1ʖD�f櫊Y�i����yM��6���H���e9k=J@v��9^�&�_���70����M�ɿZc����'��@�dPA�e��+��ej��4��E<)I�1S����RA��Q���/o�g�����J��3C���2*T<�`fn<��,
����'����D�0���4�.�T���}
p|3U����N�o(�Y���F2@�Mh�x���=q�w��
�puPP��"<�Z� IiO�1;�md��Y˩#���c2�z6��u�q U�ϩM�ţjs��Ei�D�ۜ#���g�  �@�M��qV�^�g��F����&�����zKI�E��}sH�+ܙ��K�����1��v@�6��=��TM��S$�!�q�(�%������|mZ��s��[��şɠ�{��~o�|���t>Q0���rwۈ�Ø5�}�>�E~�Q�>��HwA���0^��'g��as�Qߊte��s�L嬒&�W�+��r��2+���h�vi����u��L�Z83�g��4��웊`����%��
���PY�#�@!�����Vy�ſ���g��4!
�#�b:h��PP_��4?c��^4Hs�c4K�_�kƯ�ߖ`O̊O�$@GM�g2����n,�t�1a�'ζ2Q1���΋����k�Q��áwF���̳��w���F&-.��q�g��r����wP;6i�օ�j'�?�ݦ��'��Q�5~c5��s����@P/c�|Ҋ8��эd�8�\�=��ܷ�'���ս��:o�38@/�?v_|OY|��ڛ$�.�\=�'�V>o��@�DU�� \�Y��䑨%4�q���r��y+��Z��z��~o�9�n�v>L����IT�o�!͔bҩg��"�2{���L���Xog�Gj<qHj����c�|�Ԯ�]�PF�{��'�����/��<7\A#��T�m�藾X��\�yUi؞���r�,k��U�oL���w��gQ���'<l{l���բ��d�>;6�����dT����u�6kO�z�����{D�6�;ʆ�x��1����ՠo���izn��D[���DpV�sȣ��ߥ���S�ꟻ%n���ُ�lG@ {�s���T Vܦj�Dk		�g��R��7��1�$HV��%+X�Z���0����U�@ ȋ���un���rV�a��.�oI~0����e�n@WY,I�,s_��� <��]����a��9�^�v�o�]���b^�k��^ZB�^z&�(-E���σ{��߷S �c��0����[�Ӗ���Cb�����$���B�c��'��i�6���E��έ�B����t.p�Ͻ�F�%w<�Xx�_߆휅[�_�������1�&.��z��\6�a6��w��@��[�K'��n���gkgD/(�Y���7l��V�F�<��r�1�1F(������*�:K�n�=�=濙�� ��m����Y�,}>t�/M!��]c�{�٢z���	��.�L��HA�����N}�G4ܛw��"W��{|<���]����W���wҍ|�����[���?D8��\l�Mp�QO�¬�+k���Yn�t��f�Φ��.�pCK�ϧzO�B�l������0s��0�'L#B�������o�z��<����Ib�\x�n��d�8	�,��V�i��զ��o�J5^��֩e,d�7����Y�>������N^��0�ua�5� M�����w+,�X�H���
x���%���bO�O}�L��_(U�	�w���zdV6���ɾ���j
W�1�ǉt�.���:��g��~�����U��s�������T�˃��$��H?�`��U��0��#��'*Ѡ�:����>�,^!^�c@���B�j�A��KUC��x��)�p I�g:T�^~�ɢ�^�9*x&1�-UM��A J	��^��-=����Hc��\���.�<S�����:2M�ɇ�ǔ���:�����!�l_�q���L�2���%�#E���']Ċ��ܖ�[���`c��j�Z��|��])OԄ�X���ye�4��)m����R<'�U�c�����$�"�o�]��UG�!Ø18��W�B�f�z����K�w��q�^ğ��6 �����j��֛ƦKk��4~�~��Rݷ����G�UFz��!��"ǘR��#�l�LĞ�UrI��\�8��EY�*iWIr]�y���ڶ&ǝ�8|�B|�^k\~��g�i�჎c~�e�˂������4�]�H����	���a�̒�%�fc˭S���z�>���)GIz�K�����W%����0��\���;��۲�-���d�y�#u�w-��f���p�}�hplL�/�¯	�H�@��-?-�Fi���zDNLHY��1i0�B�|q��ߩ�~1~�lJ�� ��NΙ��[�z�;��#2{����ރ�o�CK  ͵�N#��.�����.\6�9n��*Z��U���'�j���80W<�^�.a���vD���$6׃��&� lwh_�3L�~ޔROJC8<��=O��#FOi�F:Q���Y��M��MB	H�� ;�|�%>�k��x�SJ�+7V?K��H �*��/�ѵB��I1G*Wz"fP��뭳���Ms,���iy�qY˫�ܮ�꺔?;p`ty���ID���:��@����r|N�W�����\�J(�Ĳ�@R�dJ�{�1�������L\���eR��|o>��R�,����<�7]�K��hCG��Qf���4Pe/��������	6΢m2р�](�K0�:j�E�Jf���߯q!w-����;b��p���c���L�/U+�9�Š�R1$������s ��:ms�o氎����5�&z��y�ˢv�C�DY�⛛�\ͥ�Յ|���T�ڵ�9g��j�$�z��d�"̛�A��3����9XQk_Ύ�/6ubN���L5f�ެ��I
\�юC�����9�^|���r�a5�5��l*Ҥ:n>I�h��*��g�ǗNU��Hs�BE�9�(I��%��QEcU����2H�IBY��oSN���-�,�w}��;]L�K��>xc�}q�ä�5������c��W�����֞��C�6���g`��7��.�]�8���U'���ϹZ&
C��Γ�`�����tih'
J{�$���=��	��,�<U��Up��U(��&�\��xL�h~_ssj��1���o����{���Yv@\�Ln���L˼��4j�tBm-+�7�S(�F�Aɩ����g�b[ↃN�$����,)�_lݠv��D2R~�@��[�����"m]W�0��'��Ìk����\��cq��sI��ZOj'e���N�U~82��N<ը)��-��\P��{��jwnw��\����,|d�n��P[U��R��>���L�(*��l>�z����r��Ie�7}l$.��g���1�^�	s�ʃ�
�������EEб��,k�����O��D��/�3���;k�z�v�p��S/Q	��H���[��ȟW��*8�2����Ƣz�[���Q��I���$'ĺE�D�sw��gßdm�iOm��Xo�*]���|/&X#��jX�w���	�c���ǯ:��($��烊�A�� �/�V>��GI���Əb��ߺ`¤V���I���	�Q�Y��8�;:�'�7s"ؑ'���lX��2yu���f��#��&�2|����R�������{?.E Q�;l��M��[>cZ���V&�p�g�'G��~kH��bBQD�x�v*�Y�)A%��rܼ�'2�x���+C�lڜ��ڔ������#�M?�)*�����aF�ձP�B��e�ya��>��)j�K:;�������W�_��
�<عJ�l|���Ĕ�yP�a!��|�p`�t�)f��O�|��Z��WTc���53HEq?G�`������6��$7���gB�,$��������U�����P8�|�4��,I`���Ɣ�����������O�sm�F�A ��j�L\��u:٬���������w;x��BhU��                                                                                                     �� P�             ͣ Р             �� 8�                     �� �� �� š ա � 	� � +� =� S� a� s� �� �� �� ɢ ע � �� � � #� @� Y� d� o� x� �� �� ��     ף � �� � !� -� H� U� e� y� �� �� �� Ť ۤ � � �  � +� =� N� `� n� {�     �� �� �� å ץ � � � � /� ;� X� a� l� �� �� �� �� �� �� ئ �     KERNEL32.DLL   Sleep  GetProcAddress  ExitProcess  WaitNamedPipeA  ExpandEnvironmentStringsA  GetLogicalDriveStringsW  SetEndOfFile  CreateDirectoryExA  SetThreadContext  WriteProfileSectionA  GetTempPathA  GetNamedPipeInfo  CreateWaitableTimerW  FindCloseChangeNotification  GetDiskFreeSpaceW  ClearCommError  GlobalUnWire  MapViewOfFile  CreateMailslotW  GetDiskFreeSpaceExA  GetFileTime  lstrcmpA  FillConsoleOutputCharacterA  GetSystemTimeAdjustment  LocalSize  LocalLock  SleepEx  GetFileAttributesExW  ReadConsoleOutputW  GetLongPathNameA  GetThreadSelectorEntry USER32.DLL  UnpackDDElParam  CloseWindow  TranslateAccelerator  UnloadKeyboardLayout  CharUpperW  GetUserObjectInformationW  GetKeyState  ScrollWindowEx  GetDoubleClickTime  DrawCaptionTempA  SetWindowTextW  GetPriorityClipboardFormat  GetTopWindow  RegisterSystemThread  ChangeClipboardChain  DdeCreateDataHandle  ScrollDC  CharUpperBuffA  DrawFrame  RegisterTasklist  GetClassInfoExA  UnregisterClassW  GetUpdateRgn  InsertMenuA  CallWindowProcW GDI32.DLL  SetColorSpace  StretchBlt  CopyEnhMetaFileW  GetEnhMetaFileBits  StretchDIBits  CreateDCA  GetEnhMetaFileDescriptionW  GetPolyFillMode  GetTextMetricsA  DrawEscape  CreateScalableFontResourceW  GetROP2  OffsetRgn  CreateBrushIndirect  EnumEnhMetaFile  GetObjectW  ResizePalette  ExtEscape  Ellipse  GetTextExtentPoint32W  CreatePolyPolygonRgn  GetTextExtentExPointW                                                                                                                                                                                                                                                                                �   `  �                 8  �                 P   �� �                            x  �                 �   ��                     �  (       @                                  �  �   �� �   � � ��  ��� ���   �  �   �� �   � � ��  ���                                              S�p            S�p           S�p      {0  w S�pp     � 0FS�v p     {0 �fS�vf     ���S�vf`p     {v��S�vff     w���S�vff`     ���S�vfff     k��S�vfff     ff��S�vfff   pffkfS�vfff`   pffffS�vk�f`   ffffS�vk�f`   ffffS�{k�f`   pffffS�{���`   pffffS�{���`    ffffS�x���    fffS�w���7   f`3��f�    ff`s1�`;0   pfff`ff s�   fff`ff` ;p   pfffffff   �    fffff`          Fff             w                      ���������������?�� �� ��  ��  �  ?�  ?�  �  �  �  �  �  �  �  �  �  �  �  �  �  �  a�  �� �����������                                                                                                    