MZ�       ��  �       @                                   �   � �	�!�L�!This program cannot be run in DOS mode.
$       U�}�������q�����z����N���Rich��        PE  L �JpG        �  �  R     I      �   @                     DA                                      \� P     D1                          ��                                             � �                          .text   ��     �                   `.rdata  �J  �    �             @  @.data   ��  @  �  �             @  �.rsrc   D1     2   �             @  @                                                                                                                                                                                                                                                                                                                                                                                                                                                �=��F u�1�  �t$豤  h�   �LF YYÃ=��F u��  �t$茤  h�   �l  YY�j`h�E �K�  ��   ����  �e��>V���D �N�ȭF �F�ԭF �V�حF �v���  �5̭F ��t�� �  �5̭F ��£ЭF 3�V�=��D ��f�8MZu�H<ȁ9PE  u�A=  t=  t�u��'���   v�3�9��   ��ytv�3�9��   ���E�j�@. Y��uj����Y��  ��uj�����Y�x  �u��  ��}j����Y� ��F ��^  ���F �ݠ  ��}j����Y��  ��}j	�}���Yj�  Y�E�;�tP�g���Y�u��E�P�P�D �I�  �E��E�t�E��j
XP�u�VV��P�� ���}�9u�uW�]  �z  �+�E��	�M�PQ��9 YYËe�}܃}� uW�A  �\  �M���Ǎe���  �j�����Y���VC20XC00U���SVWU��]�E�@   ��   �E��E�E��E��C��s�{S��   ���t{���t}�v�D��tYVU�k3�3�3�3�3���]^�]�t?xH�{S�k�  ���kVS蠎  ���vj�D��#�  ���C�D�3�3�3�3�3��Ћ{�v�4�댸    �#�E�H�   �U�kj�S�M�  ��]�   ]_^[��]�U�L$�)�AP�AP�(�  ��]� U��� SV�u�^��ud�   �E�E�H;ىM�r;Xs3���  W�~���u3�@��  3҉U�Ë���t;��E  �x t�EB��;�v��} t�F�;E��"  ;��  ���F ���� ���3���~9<���F ��   F;�|�j�E�PS�h�D ���`  �}�   �S  �E��tV�M�f�9MZ�?  �A<��8PE  �.  f�x�"  +�f�x �H�L�  �A;�r�Q�;�s�A'�uwjh��F ���D ����������F �ɋ�~����F 98tJ������u-j[;���3҅�|����F �0B;Ӊ8��~��}A���F j h��F ���D ����3������������D jh��F �Ӆ��z���9<���F t.���F �p���|9<���F tNy��}��}@���F �p��t3Ʌ�|����F �A;Ή8��~�j h��F ���������_^[��VW3���F �<�,~F u��(~F �8h�  �0���h�  ��YYtF��$|�3�@_^Ã$�(~F  3���S��D V�(~F W�>��t�~tW��W�V�  �& Y����HF |ܾ(~F _���t	�~uP�Ӄ���HF |�^[�U��E�4�(~F ���D ]�jh@E ��  �u�4�(~F 3�9urj�U  Y��;�u�}7  �    �?j
�b   Y�]�9u8h�  W菙  YY��u#W貕  �J7  �    j��E�P�Ҋ  ��3���>�W苕  Y�M���	   3�@�8�  �j
�M���Y�U��EV�4�(~F �> uP�G�����Yuj�.���Y�6���D ^]�jh0�D ��  �u�=�`F u.;5ŖF w&j����Y�e� V�T  Y�E�M���3   �E��u#��uF�=�`F t�����Vj �5��F ���D ��  Ëuj����YÃ|$�w"�t$�u�����Yu9D$t�t$�   ��Yu�3���5��F �t$�����YYá��F ��t�t$�Ѕ�Yt3�@�3��hd�D ���D ��thT�D P� �D ��t�t$���t$���D �j�����Y�j����Y�V������t�Ѓ�;t$r�^á,�G ��t�t$��YVW���G ���G 3�;ϋ�s��u?���t�у�;�r��u,h��@ ��? ���G �ƿ��G ;�Ys���t�Ѓ�;�r�3�_^�jhp�D ��  j�$���Y3��}�3�F95�F u�u���D P���D �5�F �E� �F 9}u79=��F t�L�F ���L�F ;��F r
� ;�t�����h��G ���G ����Yh��G ���G �����Y�M���   9}u!�5�F �u����3�3�F9}tj�����Y���  �j j �t$�0������j j�t$�������jj j �������jjj �������jh�E ��  3ۉ]�j����Y�]�j_�}�;=ɄF }V������F �;�tB�@�tP��  Y���t�E��|(��F ��� P��D ��F �4�/�  Y��F �G럃M���	   �E����  �j�����Y��Jx	�
�A�
�R�~  Y�h�  h�E �g�  � {F �E�3���D�����(�����P�����l�����k�����|�����H����E� ����  ��P��h  Y��tG��|�����|����U�x�����V�h  Y��u���t�uV��  YY�E�E� P�h  Y��u�랋u�>%��  3���`���ƅh��� ��d�����L�����t���ƅ_��� ƅi��� ƅr��� ƅ���� ƅj��� ƅ{��� ƅs�����8���F���P�g  Y��t��L������|C��   ��N��   ��   ��*tr��F��   ��It��Luv��s����   �N��6u �F�84u����8�����T��� ��X��� �e��3u�F�82u���T��dtO��itJ��otE��xt@��Xu�9��r����1��ht ��lt��wt���������s�����{������s�����{��������� ������t����u��r��� u�E��$������E�X���P������P���ƅ���� ��{��� u�<St<Cƅ{����uƅ{����>�� ��@�����nt3��c��   ��{��   ��|����U�f�����V�f  Y��u創l����u��L�����t��t��� ��  ��o��  ��  ��c�}  ��d��  ��  ��g~_��it<��n��  ��|�����r��� �j	  �	  ��|����u���������l����|���jd_��l�����-�  ƅi����  ��������l�����-u���������������+u ��t�����|����}���t����؉�l�����}��L��� t��t���]  ~:ǅt���]  �.��t�����t�����t)��d����F��|������ ����؉�l���S��d  Y��u�8`{F ub��t�����t�����tR��|�����������ؠ`{F �F�(��t�����t�����t)��d����F��|�����������S��l����kd  Y��uǃ�d��� ��   ��et	��E��   ��t�����t�����ty�eF��|������g����؉�l�����-u�F���+uF��t�����t�����u!!�t����.��t�����t�����t)��d����F����|��������؉�l���S��c  Y��u���|������t	WS�`	  YY��d��� �)  ��r��� �{  ��H���� ������P��P�����s���HP�{F ���N  ��uǅL���   ��t�����{��� ��  ƅj����  �ǃ�p�  ��t�HH�	  ���������t;�E� ;�l���t��l�����I  ��k�����r��� ��  ��$����E��  ��{��� ~ƅj����}G�}��0����?^uG��0���ƅ_������D�����u]!]�j X���  �e�܉�D����M���A3�@Ëe�� j ����Y��D�����u	�M����  ǅ(���   �M����0�����D���j j S�" ����@���{uw�?]ur�]G�C �oG<-uK��tG���]t@G:�s�����:�w+��*�������,�������Ë΃����F��,���u�2����h����ȋ���Ã������h����<]u����)  ��P�����@���{u�}��@�������|�����l����t�u��l����  YY��L��� t��t�����t�������  ��|����U�z�����l��������  ��ctM��su��	|��~�� u9��{��  �ȃ�3�B�������D����9��_���3υ��d  ��@�����r��� �K  ��j��� �0  ��<������{F �DA�t��|����U�������=����5\{F ��<���P��4���P��  ��f��4���f�CC��   ��+u*��t���u��t	ƅ�������|����������؉�l�����0�]  ��|������c����؉�l�����xtO��XtJǅd���   ��xt��L��� t��t���u������jo_�  ��|������t	VS�  YYj0[��   ��|�����������؉�l�����L��� t��t�����t���}������jx릈C��P�������F������|������t�uP�  YY;���  ��r��� �:  ��H�����@���c�'  ��P�����j��� t	f�  �  �  �  ƅs�����l�����-u	ƅi������+u*��t���u��t	ƅ�������|����������؉�l�����8��� �]  ������ �  ��xtf��ptaS�^  Y����   ��ou*��8��   ��T�����X���������T�����X����fj j
��X�����T����� ��T�����X����CS�^  Y��t2��T�����X���������T�����X���S�!^  Y��u��߃�������������� uA��d����CЙ�T����X�����L��� t��t���u	ƅ�����%��|��������������|������t	VS�b  YY������ �������l�����i��� �  ��T����؋�X����� �ى�T�����X�����   ������ ��   ��xt6��pt1S�O]  Y��tK��ou��8}A��`����>��`���������`����+S�X]  Y��t��`���S�]  Y��u��߃�������������� uA��d�����`����DЉ�`�����L��� t��t���u	ƅ�����%��|���������������|������t	VS�M  YY������ �/�����l�����i��� t��`�����Fu��d��� ��d��� ��   ��r��� u>��H�����P�����`�����8��� t��T������X����C���s��� t��f���k����E�w��|����U�=����؉�l����F�u;�u9�Ë{F �DA�tF��|����U�����F�u;�t'���t�uP�f  YY���t7�u��l����Q  YY�%��|�����l����� ����E�8%u
�xn������(���u��D���詄  Y��H�����l����u��u8�k���u���������M�軀  �6�  �V�t$�F����   �@��   �t�� �F�   ��f��Fu	V���  Y��F��v�v�v��  �����Ftr���tm�V�u:�N���Wt�����<�̈́F ���ɍ<����yF �O�ႀ��_u	��    �V�~   u�N��t��u�F   �H�F�A�^��������	F�f ���^�S�\$���VtA�t$�F�u��y2�u.�~ uV���  Y�;Fu	�~ u@���F@�t8t@����^[È�F�F�����F��%�   ��U����  �@`;4�F t��  �} u3�]��p�u�u�u�uj�p�B' ����u����]Ã��]�V�t$��tV�` @P�.�����YYtVP�\�  YY^�3�^����̍B�[Í�$    �d$ 3��D$S�����T$��   t�
��8�tτ�tQ��   u��W����V؋
����~����3���������3�3ƃ��� �u% �t�% u��   �u�^_[3�ËB�8�t6��t�8�t'��t���8�t��t�8�t��t��^_�B�[ÍB�^_[ÍB�^_[ÍB�^_[��̋T$�L$��   u<�:u.
�t&:au%
�t��:Au
�t:au����
�uҋ�3�Ð��������   t���:u��
�t���   t�f���:u�
�t�:au�
�t���눃�HS��  S������Yu�����  �̈́F ���F     ���  ����` �@ �@
�̈́F ��$���  ;�r�UVW�D$P���D f�|$F ��   �D$H����   �8�h�/�D$�   ;�|��9=��F }N�фF S������Yt8���F  ����  ����` �@ �@
���$�;�r��9=��F |���=��F 3ۅ�~j�D$� ���tT�M ��tL��uP���D ��t<�ˋÃ�������̈́F �4��D$� ��E �F�Fh�  P��  ��YYt.�F�D$CE;�|�3ۋ̈́F �ۍ4��>�uo���F�u
j�X�����y��H������P�p�D �����t?W���D ��t4%�   ���>u�N@�	��u�N�Fh�  P�\�  ��YYt��F�
�N@��N�C���r����5��F �x�D 3�_^][��H�U��SV�u�F���^��   �@��   �t�f ���   �N�����F�F�f �e ����f��Fu"��xF t���F uS�G ��YuV�j�  Yf�FWtd�F�>�H��N+�I���N~WPS��  �E�3���t������̈́F �Ã��������yF �@ tjj S�T  ���F�M��3�GW�EPS萊  ���E9}_t�N ��E%�   �	�� �F���^[]�U��MV3�;�u3��L�E9puf�Ef=� w,�3�@�3�URV�p(�uQj�MQV�p�D�D ;�t9ut�  � *   ���^]����  �@d;�{F t� �t$�t$P�}����������������U��WVS�M�'�ً}��3����ˋ��u�F�3�:G�wt���ы�[^_�Éh�F �Yx��F ���ʼ �,�F �K��\  �s�4�F �C���F �K ��F � �F �C$��F ���F �[��F ��F    ���8 ���F �,�F � ��X  ���X  �,�F �����@��$<  ��D  �����+����B��Y�ʉ5T�F �������@  ��L  ��F �L�F �d�F �\�F ���<  ����L  �5��F S�[  É�l  �5,�F ��X  ��`  ��@����T  ��h  ��  ���  ��\  NX��P  ��d  ��Y  hf hY~A ��X  ��L  ��H  ��4  �  �T$���   �l$���%�F G�n����   ���	  +��F ���  %~����F ��
  �}��=p�F =P�F 3�@	  ��F ���F �%<�F �58�F �=0�F �}���   ��F �  ���F ��F ��F �%��  �� ����,�F ���F ��<  ���F �؋�X  �=��F ���F ��<  ��P�w���  �D$����F �%��F ���	  ��,  �����  Ë5��F �N<�q|�5��F j
RV�5��F �O���V���  ����  ��d  ��+��  ;��F �y� ��    W�=��F �;��F ;��F ��~ �5��F �5,�F ǅ����
  ǅ���}�E �5`�F ��V���F ��X  �!  ���,�F ��X  ��f h�#  j ��$T  ��D  �# ���,�F h�  �5��F ��<  ��|  �(�F 靸 �-��F �<�F �!<�E����F +t�F �}�3=��F �0�F =��F ���  �0�F ��F ��8	  �}��F ���  ���   �5�F �w�5�F �w�U��]����   ���  �W��  �W���  �G���   ��F �E��]���  �m����  ���F ��,  ���	  �����V�l�F ���D �5d�F P��8  ���   ��4  �ы�8  ��F ��@  �|�F ���F ���F �|�F ��D  ���E���� �F ���F ���F �T�F �����   �h�F ���F ���F ��$�  ��$�  ���F �h�F +��F ��F �T�F ��$�  ��$�  � �F 뉋D$���   �l$Ћ� �F HX��x%  �d)  +�+  +�F PX�M̋�*  �-h�F ���*  �h�F 3��F ���M���*  ���*  �  _��$  ���  ���F �=��F �D����X�F ���F ���F �%��F ������F ; �F �{"  ���F ��F ��$�  � �F �<�F ���F ���F �
Ǉ�      �<�F ���F ���F ��$�  9�F �2:  �=�F �=�F =�F ���F ������F �T�F ���F     �:�����  ����H  �� `  �5��F �����É��   ���   �Y���   �Y�}ȋ��(  �y�ẺA�Q���   �5T�F ���F �}ЋEȋ��'  ��F �=��F �h�F ��p%  ���F �M̉ �F ���F �%D�F �Ƌڋ�5T�F �=h�F É=<�F �=,�F �3���  ���F �[�=<�F ���  ����F ��8  j �   É��  �x�F �H�F ���F 4���  ���  �Ã�4��  jhP�D �@�  �}3�;�u�u����Y�  �u;�uW�u  Y�o  �=�`F �.  �]�����   j����Y�]�W�!-  Y�E�;���   ;5ŖF wLVWP�2  ����t�}��8V��4  Y�E�;�t*�G�H�E�;�r��PW�u���  W��,  �E�WP��,  ��9]�uK;�u3�F�u������uVS�5��F ���D �E�;�t#�G�H�E�;�r��PW�u��  W�u��,  ���M���O   9]�u";�u3�F������uVWS�5��F �$�D �E�E�;�u`9��F tXV�����Y��������E3ۋu�}j�5���Y�3����w;�u3�FVWS�5��F �$�D ;�u9��F tV����Y��u�3����  �ǅ     ���F     �58�F �5��F �5��F j V�u   �Wjd�����Ë�@=-   �M  ���F j�5|�F �5��F jdQ�   Í,�F ���  �5��F �3C%�   =�   �X����5,�F jdQh�  �5��F �l���Ë=<�F ���F ���F �9�5|�F �  Ë��  ���L  ��h  �+�$  �=��F ��h  �;�[I��   ���  ��@  �׋H�F �=��F ���   ���  ���F �-H�F ���  XX��`  ��P��t  ���D �,�F ��F �%��F �,�F �<�F �\�F +0�F �H�F 3��  ���5��F ����Ë�$�  �� @ �쉝8  �,�F �p�F ���F �@�F j �p���É�h  �8�F �H�F Vj �5|�F �����É�@  �,�F ��  ��$�  ��� ��x  ��t  �=��F ��<  ��  �=<�F ��F ���F �5L�F ���F ��,�U����5L�F �5��F ��F ���F �3ǅ�      �58�F h�  h�  �5�F �;����j Rj
jdh�  �   Ë5�F ����F h�  Pjdh�  �|   Ë��F ��$�  �4�F L$�L$��%��  ��$�  ��$�  ��$�  �=��F ��$�  ���F �ȋ�$�  �-��F ��$�  U��$�  �=��F �4�F ��$  ���  �5�F ��D��   ��F �,�F ���  ��F ���F ǅ�     ���F     �֋��  ���  ���F �5��F ���F ��F ���  ���v���F ��   _�X�F ��d����4�F ���F �H�F P�=��F �X�F ��d�����   ���F    ǆ�#      jh�  �5��F �5��F �5��F �   ��tD�5,�F �5��F �5��F Pj
Q�F���Ë�  A�,�F ��  �5t�F �5<�F Wjd�  Í5,�F �1�I��֍5,�F R���#  ���������d%  �Ή  ���$  Z���$  ���#  �������j�����<  ���F ���F ���F Z�p�F �`�F ��,�  ���F �$�F     �$�F ��F ���5|�F �'  ËH<�h�  �5|�F WQh�  �V   �=`�F ���F    ��۶ W��   ��  �=x�F �`�F �p�F ���F ����  R��)�9��;����J  �Q|�qxƅ���  �=x�F �=,�F �N�~��<  �v�p�F �`�F ��<  �@ `�F ��0  ��<  �_$`�F � �p�F ���T�����������UU��WV�u�M�}�����;�v;��|  ��   u������r)��$�L?@ �Ǻ   ��r����$�`>@ �$�\?@ ��$��>@ �p>@ �>@ �>@ #ъ��F�G�F���G������r���$�L?@ �I #ъ��F���G������r���$�L?@ �#ъ���������r���$�L?@ �I C?@ 0?@ (?@  ?@ ?@ ?@ ?@  ?@ �D��D��D��D��D��D��D���D���D��D��D���D���D���D����    ���$�L?@ ��\?@ d?@ p?@ �?@ �E^_�Ð���E^_�Ð���F�G�E^_�ÍI ���F�G�F�G�E^_�Ð�t1��|9���   u$������r����$��@@ �����$��@@ �I �Ǻ   ��r��+��$��?@ �$��@@ ��?@  @@ H@@ �F#шG��������r�����$��@@ �I �F#шG�F���G������r�����$��@@ ��F#шG�F�G�F���G�������V�������$��@@ �I �@@ �@@ �@@ �@@ �@@ �@@ �@@ �@@ �D��D��D��D��D��D��D��D��D��D��D��D��D��D���    ���$��@@ ���@@  A@ A@ $A@ �E^_�Ð�F�G�E^_�ÍI �F�G�F�G�E^_�Ð�F�G�F�G�F�G�E^_�����V�D$�u(�L$�D$3���؋D$������d$�ȋ��d$��G�ȋ\$�T$�D$���������u�����d$�ȋD$���r;T$wr;D$v	N+D$T$3�+D$T$���؃� �ʋӋًȋ�^� S�p�F ��    P������������;�$�  �Ϸ ��F X��F ��<  ��������,�  ��믋�  +P�F A�ыP�F �ʉ�  �5P�F �=L�F �=,�F �58�F ��  ��  ��F �\�F ��5,�F ��F ���D ��$�  P�   ǅ<      Q�  Ë��  ���F ���  ���  �-4�F ��$�  �\$��-H�F ��$�  ��$�  ��$�  �=��F �=��F W�=��F �ˋ�$�  �5��F ��$�  ��Ř  �������`  ��   � �D �=L�F ��   ��������  ��F ��������������  ��  ��X������(  �D�F ��F �,�F ���  ��  ��$  ���D �,�F �5��F j�5��F �5��F j
�W���Ë`�F Q��F ��F ��F �%��  Q�Љ= �F �������������=�F ��  ��  �-d�F �l$�= �F �\$�`�F ���t  �%@�F Q�������������������,�F �$�F Ӫ�  ��  �5��F �l�F ���D �,�F �<�F ʉ�  ���  +��  ��F �X�F 3P�F ���ȗ ��F ��   �<�F Sh�  �5��F j����ËQ|�qxƅ��N  ��F �,�F �N�V�=��F �~�5�F �v Ɖ�0  �=�F �$ǉ�   ���F ��F �@� �5��F �5,�F j<V�58�F j W�J���Ë�<  ���F ��(�5����4�F �=P�F ���  �;��F �{  G�P�F ���  �P�F ����)  ���  �4�F ���  �=P�F 몉��  �=��F ���  ��F �  ���  �,�F ��5��F ��[V��|  �5��F �Ë�|  [���  ���F ���  ���$�  9�$�  �P-  ���  �=$�F ���  �=��F ���  �=��F �
������  �,�F ���  ��T  ���  �<��[���  ���  ��T  ���  ����$�  ���  ;�$�  ��� �$�F ���  ���  ���F ������,�F ǅ�      ǅ�      h�  �5|�F �   Ë��  @P�5��F �5��F j
��  Ë,�F �ʉ��  ���  ʁ��  ���`�F ӆ�  �$�F     ǅ�      ǅ�      ��T  ���F ���  �33$�F �[�433�$8  �\�F ���F �]    �T�F �   ��ǅ�     � �F �ˋ �F ��)މ��  �5 �F 35 �F )�$�  ���  � �F ��3T�F )�$�  �=��F ���  +=h�F ����)5 �F �5��F 1�)5 �F ��F ���%��F V�5�F �"WP�t$��������u��<=t��t�����u؋�+�F ^����Ë�+�F ^���U��Q3Ʌ���u�Ã? t	��A�8 u�S��   VP���������Y�u�uj	�>���Y����P�r���������Y��u�!�E�^[��U����ES3�;�W�]�u����aV�0;�u�tSj=V��  ;�YY�E�tB;�t>3�8X��F ��;�F �M�u���H�����F ;�uU9]t9�F t��r  ��t?���^_[��9]�t3���j����;�Y��F tމ9�F uj�����;�Y��F tÉ�}�+}��u��5�F ������;�Y|F9tB�4��6�Wb  9]�Yu�E���E��g�F�G��9u����P�5�F �_���;�YYtC�<9]���   ;�}�ߍ�   P�5�F �5���;�YY�4����U�����Y�M���F 9]tP�u��e�  @@P�2�����;�YYt8�u�V�\�  ��+E�YE�Y�M��@�����#�QV���D ��u�M��V�a  Y9]�t	�u��|a  Y�E������u��ka  �EY������$�  �<�F ���  ���  ���  jd��  �=�  �< �T�F �,�F ���  ���F �h�F ���  �C���   ���   ������54�F ����ËP�F ��  S���  _X�d�F ���F +��F ���  �d�F �GX�l�F ���  ���F +��  ��`  �p�F ��  ���	  (+<�l�F WX���  ��$�  ��F - �F ���  V�54�F Q�����Ë(�F 3�	  ȋ��
  ω��F �,�F ���  ��F ӪL
  ����L
  0�ys��$8  #e��zX���  JX�8�F �(�F ӊL
  ���  ��L
  BX��	  ���F ���  ��p	  ��  +�  �5�F ��  �ƭ 1DZX��x  � �F ȋ�X	  �����F #8�F ���  �5,�F +�`	  ��$x  �\�F ���  9���  ���  �P�F �T�F �h�F ���  �<�F �P�F ���  ���F ���  ��$�������3T�F ) �F ���  �= �F +=��F �T�F +��F ��$  ���  ��������T�F �= �F ���  �ȋ��  �=��F ��F �6������  �,�F ��X#  $��h   �54�F j�5��F � �����\�  ����S�  ���V�I�  �L$�H3�;�hxF tF��-r��r$��$w�"�  �@   ^���  ��lxF �H^Á��   r���   w��  �@   ^���  �@   ^É}���  �5 �F ���  ���F � ���U  �����  ���  ӄ$�  +��F �$�  ���F �x�F ���  ���  ���  ���ǅ�      R���  ��F �U�5 �F �h�F �<�F �}���  ;�$�  ��� ��$�  �$�  ���  ���  �$�  � �F ���F ǅ�      �������  �h�F ���  �F 9h�F ��  �5p�F ���F �5h�F ���  �5��F ���F ���  ���F �h�F �;��F �n  �h�F ���F ���F ���&  ���F 뵃���$�  ������F ���  ;��F �5� ���F ��$�  ���  �=��F ���  ���  ��F �,�F �=<�F ���  �U���F �}�h�F �=��F ��  �H<�j �5��F jd�5<�F �}�����F ��$�     �� � P�,�F ��  �=��F ��D  ����  ���  ��+�$�  ;��F �J����  ���  ���  ���  �����   ���  ���  ӄ$�  �p�F ���  +��F �$�  F�V��`�����h�������  �=(�F �>����   ӄ$�  +=��F �$�  F���  �=(�F ���  �ƋH<��Q|Q�5��F �5��F h�  ��  �@ �F ���F    ��f� Q�,�F �5T�F �5��F ����  �0�F ��+�$�  ;E�u  �  ���  ������F ���  ;d�F �)  ���F �=(�F �p�F ���F ���  ���  �=��F �3�,�F �������  ������F ���  ;d�F �P*  ���F ���F ;�$�  �.  ���F ��F ���  �(�F ��)-��F ��$�  ���F ��$�  ��$�  ��$�  Ǆ$�      �-p�F �=(�F �݋�$�  �5p�F ��$�  ��$�  ��$�  ���<����d�F �,�F ��$�  �����F     95��F ��%  �,�F ���  ��d  ��d  �d  �4�F �����F ���  ǅ�      �i������  ���  � �F ��  �ixŅ���� ��$�  �5,�F �싵�  �N�v�=@�F � �F ���  �@���  ���  �@  �F ���  ���  �v$5 �F ���  ���  � ��P���D ��$�  P��  � �D ��  ��  �l�F ��h���� �F ��d������F ��L����@�F ���   �a  ��F     P����Ã���������  ����    W�=0�F �8 �F ;�$�  �2R �=\�F _�|�F �=t�F ω��  �}���  ���  ���  ���  �U�  ���F ��    V��h����1��F ;�F �oN P���F X��F ���F ���K���W���F �t�F �E�ʉT�F ���F ���  ��F �N������58�F ^5��F 5��F �����  ��F ���F �5H�F �U�����F �58�F ���  �H�F ��F ���F �h�F �U�  ��  ��F��$h  ��  ��+�$�  A�ы�$�  �ʉ�  ��  �=4�F ���  ���F �@�F ��  ��  � �F �\�F ����  ��$(  ���F �H�F �ȋ�Ř  �����t�F �Q�|�F     �5 �F �F<��H|�Px���9� �,�F �B�r���F �BP�B  �F R�R$ �F ���  �h�F [険 �l�F     ���F �A<ȋH|�Px��F ���  �=,�F �B�r�z�j -��F ��$�  �z$=��F ��$�  �Z��F ���F    ��Z� �-x�F ���F �,�F �  ���F �<�F �F �F �
����  ��$�  ��$�  ��$�  �=(�F ���F ���F �=<�F ���F �=��F ��$�  �9  �����  Y��F ��F �%��  ����    �=��F ��F ���  � �F ;�$�  �^N W�5��F �ʋu�5T�F ���  ��F �������  ���  ���  ��F �  S���F C���F ���F ���F )�A���щ��  �����  �=��F 󤉍�  �X�F ���  �5\�F �7���F ��Q���F ���D SP�@�F � �D �U�5@�F ���  ���F ���  �]���  �T�F �M���  �]���  ��F ���������  ����  ���  ��+�$�  ;�$�  ��  ���  �,�F ���  ��    ���  ���  �0��F 9��M� ���  ���  ���  ���F �|  �m  �=0�F ���  ���F �������X�F ���$�  �$�  �����  �=�F �t�F �5h�F �-X�F �ʉ-��F �5t�F ��$   ���8���  ���  �,�F ���  ���F ����W�=��F ǅ�      ���F �t�F ˉ��  ���F ���  �|�F �ˋ��F �U���F ���
���SP���  �U �\�F �ҋ��  ���  �5D�F ���  ���  � �F ���  ���  ���  �������H�F �5d�F ���  ���F ���  �Љ��  �H�F ���F ���  ��������F     ���F �A<ȋH|�Px��F ����   �5,�F �B�r�z��F �J ��F �5��F �r$5��F ���  �R��F ��$�     ���� ���F �  ���  ��C��$  ��+��F @�$�F ���F ���  �$�F ���  �����  ��  �= �F �=\�F � �F �8��  ��P���  ���D h   Q�u���Í5,�F �h�F     ���F �A<ȋH|�Px��F ���  �=,�F �B�r�j�z =��F ��F �Z$��F �@�F �B��F �d�F    ��������$�  ���{#  ���$�  �$�  �����  �5��F �=��F ���  ���  �5��F ���  �$�F ���  �=�F ���  ���  �É=x�F ���  ��F �=��F �M�����$�  ���F ��    �=��F �8��F ;�$�  �b�  ��$�  ���F ��$�  ��$�  �5�F ��$�  ��$�  ��$�  ��F ���F ��$�  �  ���$  �$  �����  ���  ��    �-�F �)��F ;�$  �)� ��$  �-0�F �L$0�5@�F R�-��F ��$  �T$<�=�F ^�d�F ��$  ���(��0�  �  ���F �M �`�F �ы��F �=��F ���  ���  �5p�F ���  ���  ���  �h�F �  ̋L$W����   VS�ًt$��   �|$u����   �'��������t+��t/��   u����ua��t��������t7��u�D$[^_���   t�������   ��   u����ut�����u�[^�D$_É����t�����~�Ѓ��3��� �t܄�t,��t��  � t��   �uĉ�����  �����   ��3҉��3���t3������u����w����D$[^_�SV�t$�F�Ȁ�3ۀ�u:f�t4�FW�>+���~'WP�v��X  ��;�u�F��y����F��N ���_�F�f �^��[�V�t$V������Yt���^��F@t�v��Y  Y���^�3�^�jh�E �է  3��}�}�j�Ӷ��Y�}�3��u�;5ɄF ��   ��F ��;�t\�@�tVPV��  YY3�B�U���F ���H���t/9UuP�f���Y���t�E��9}u��tP�K���Y���u	E܉}��   F�3��u��F �4�V��  YYÃM���   �}�E�t�E��Q�  �j�f���Y�j�$���YË��F ��S���F ���D �5(�F P�x�F �U ���  �ҋ��  �5x�F ���F �d�F �=$�F ���F ���  ���j  ��@���F ���F ��+4�F A�ы4�F �ʉ5P�F �54�F ���  �=��F �5�F ���  �|�F ���  �(�F �\�F ��9������F ��$�  ���F ���  ��$�  ��$�  ��  ���  �������  ���F ���  ��F ������@  ���  ���  ���  ������h�F @�T�F �h�F )�B��$�  �։��  ���  �=��F �=T�F 󤉝�  ���  �=�F �5\�F �7�p�F ���T�F R���F ���D �5��F P�q������F �$�  �$�  �����  ���  ���  ���F �5L�F ���F ���F ���  ���  ���F �5d�F ���F ���  �  �,�F ���  ���  ����  ���  ��)�;��  �������    ���  ���  ���F ;�$�  �����h�F ���  �h�F ������$�  �[��F ���     ���������F ���  ���F ��$�  ��$�  � �F %��  ��+�$�  ;�$�  ������&���h@  j �5��F ���D ���laF uËL$�%(QF  �%�`F  ���F 3��ŖF �p�G    @á�`F ���laF ����T$+P��   r	��;�r�3��U����M�AV�uW��+y�������i�  ��D  �M��I���M���  S�1��U�V��U��U����]ut��J��?vj?Z�K;KuB�� �   �s����L��!\�D�	u#�M!��J���L��!���   �	u�M!Y�]�S�[�M�M�Z�U�Z�R�S�M�����J��?vj?Z�]����]���   +u��]���j?�uK^;�v��M�����J;։M�v��;�t^�M�q;qu;�� �   �s������!t�D�Lu!�M!1��K�����!���   �Lu�M!q�M�q�I�N�M�q�I�N�u��]�}� u;���   �M��ыY�N�^�q�N�q�N;Nu`�L�M���� �Ls%�} u�ʻ   ���M	�   �����D�D	�)�} u�J�   ���M	Y�J�   ��ꍄ��   	�E���D0��E����   �(QF ����   ��mF �5��D h @  ��H� �  SQ�֋�mF �(QF �   ���	P�(QF �@��mF ����    �(QF �@�HC�(QF �H�yC u	�`��(QF �x�uiSj �p�֡(QF �pj �5��F �8�D ��`F �laF �����ȡ(QF +ȍL�Q�HQP��  �E����`F ;(QF v�m�laF ���F �E�(QF �=�mF [_^�á�`F �p�G W3�;�u4�D�P��P�5laF W�5��F �$�D ;�u3�_Ãp�G �laF ��`F �laF Vh�A  j�5��F ���4����D ;ǉFu3��Cjh    h   W���D ;ǉFu�vW�5��F �8�D �ЃN��>�~��`F �F����^_�U��QQ�M�ASV�qW3����C��}���i�  ��0D  j?�E�Z�@�@��Ju�j��h   ��yh �  W���D ��u����   �� p  ;��U�wC��+����GA�H�����  ����  ��������@��  �Pǀ�  �     IuˋU��E��  �O�H�A�J�H�A�d�D 3�G����   �FC�������E�NCu	x�   �������!P��_^[��U����M�ASV�uW�}��+Q������i�  ��D  �M�O����I;�|9���M�]��U  ���E  �;��;  �M���I��?�M�vj?Y�M��_;_uC�� �   �s��M��L��!\�D�	u&�M!������M��L��!���   �	u�M!Y�O�_�Y�O��y�M+�M��}� ��   �}��M��O��?�L1�vj?_�]���]�[�Y�]�Y�K�Y�K�Y;YuW�L�M���� �Ls�} u�ϻ   ���M	�D�D��� �} u�O�   ���M	Y����   �O�   ���	�U�M��D2���L���U�F�B��D2��<  3��8  �/  �])u�N�K��\3��u��N��?�]�K�vj?^�E���   �u���N��?vj?^�O;OuB�� �   �s����t��!\�D�u#�M!��N���L��!���   �	u�M!Y�]�O�w�q�w�O�q�uu��u��N��?vj?^�M��y�K�{�Y�K�Y�K;KuW�L�M���� �Ls�} u�ο   ���M	9�D�D��� �} u�N�   ���M	y����   �N�   ���	�E��D�3�@_^[��U����M��`F �laF �����S�M���V��WI�� �<��}�}�����M���������3���E����F �؉u�;���K�;#M�#��u��;]��]r�;]�u$����K�;#M�#��u
��;؉]r�;���   ���F �C�����U�t����   �|�D#M�#��u6���   #U��e� �HD�1#u�֋u�u���   #U��E����9#��t�U���i�  ��D  �M�L�D3�#�um����   #M�j _�^�{ u���];]�r�;]�u&���	�{ u
��;؉]r�;�u�����؅ۉ]tS����Y�K��C�8��$���3��z  ��G��}��M�T��
+M�����N��?�M�~j?^;��  �J;Ju\�� �   �}&����M��|8�Ӊ]�#\�D�\�D�u3�M�]!�,�O���M�����   �|8��!��]�u�]�M�!K��]�}� �J�z�y�J�z�y��   �M��y�J�z�Q�J�Q�J;Ju^�L�M���� �L}#�} u�   �����	;�ο   ���M�	|�D�)�} u�N�   ���	{�M�����   �N�   ���	7�M���t�
�L���M��u�эN�
�L2��u��ɍy�>u;(QF u�M�;�mF u�%(QF  �M���B_^[�É�$�  ����F �D�F �  ��$�  ��$�  ���F ��$�  �=`�F �=��F ���F ��$�  ��뭋��F ��������F �5��F j
�5��F ����É-H�F �D�F ��$�  ��$�  �  ���  �������  �����F R���D �5��F P���F �U ��F �҉��  �0�F ���F �`�F ���F �-��F ��$�  ��$�  �W�����  ��@���F ���F ��)�@�։�F ��H���  P���  �L�F ��F �։��  �=��F �5��F ���  �\�F ��5��F ��  QQ���F SU�-d�D VW3�3�3�;�u.�Ջ�;�t���F    ����D ��xu
jX���F ����F ��uX;�u�Ջ�;�u3���   f9��t@@f9u�@@f9u�+�@@��U������;�Yu3�V���D ���   UVW�<��������t;�u����D ��;�t�8] ��t#SSj�VjS���D ;�t�V�豹  �t8Yu�G�?P�|$�o���;�Y�D$tb8] ����t:�L$��+D$��+�QVj�WjS���D ��t/W�b�  V�|�ܒ  8YY�tFu�Uf����D �D$_^][YY��t$�:  YU���D ������L$;��F VWsX�����<�̈́F �����4������@t7�8�t2�=PF u3�+�tItIuPj��Pj��Pj���D ���3�������� 	   �����  ���_^ËD$;��F s�ȃ�����̈́F �����@t� ��~���� 	   �|����  ����jh��D �G�  �}�����ǃ�����̈́F �4�3�9^uAj
�,���Y�]�9^u(h�  �FP�U=  YY��uj��E�P�.  YY3��,�F�M���)   ����������̈́F �D�P���D 3�@���  Ë}j
����YËD$�ȃ�����̈́F ���D�P���D Í,�F ���  ���F ����  �5d�F ��+�$�  ;�$�  �H�����    ���F �d�F ���F 9���������F ���F �l�F �����d�F �$�F ���  �Ճ��"�������F �F �����  �T�F ���  ���  ���  ���F ���  ���F � �F ���F ���  ���  ���  ���  ���  ���  �������S��F �5@�F ��  �|�F �0�F ��  ��  ���F �U8[��F �=�F ��  �d�F ��  �E0�=�F ��F ��(��0��  �p  ���  �=(�F ���  ���F �-4�F ���F �=d�F �5p�F ��$�  �-��F ���F ��$�  ��$�  ��$�  ��$�  �d�F ��$�  ��$�  ���F ���F ���F ��$�  �  ���  ��@���F ���  ��)�B�ˉ5t�F ���5�F V���  ���F �L�F �5��F ���F �L�F ��$�  ��=��F �=��F �\�F �h�   j
W�5�F ��  Ë��F @���F ���  �=��F += �F G�ϋ �F �ω��  �5 �F �=��F ��5 �F �0�F �����F �<�F ���F �\�F ��L������  �$  �$  �����  S�=��F V��F �H�F �򋽴  �E��-H�F �l$���P�3  ��$�  ���D�F     �=��F �G<��H|�xx=��F ���7������F �,�F �G�W�5��F �w���  �O ��F ���  �G$��F ���  �w5��F ���F    ���� ���F �%������  �!�����$�  ���  �L�F ���F     �5��F jdP��  É@�F ���F �L�F �5��F P��F � �D ���  ���F ��F ���  ���F ��<�w  V���  �$  �$  �%��  ����    ���  ���  ���F ;U��)� ���  �= �F �(�F ���  ���F ���  �=0�F ���F �5��F ���  �E��4�F �$�F ���  ���F ���  ���F �^  �5��F �=��F ��$�  �5p�F ������  P�]��F ��(���������F �=�F ��F �}���L�F ���F ���  ��F �5��F �L�F ��  ���  ��F �R���  ���F ��F ��(���9�����F �-S���  ���  ���F ��F ���F �E��;  �5,�F �=�F ��W�L�F �5��F ���  �L�F �,�F ǁ�      Wj �b  ËJ<ыQ|�qx5��F ����  �=,�F �N�~���F �N���  �N ��F ���F �V$��F ��F �^��F ���F    ����  �5$�F �5,�F � ���F �E��M���M�9��F ��� ���F �=��F �E��=��F �=��F �   ���F W�=���P���  %��  ���  ��+�$   ;��F �������    �4�F ���F ���F ;$�F ��� ���F ^��F ���  �L�F ��F ��PS�L�F ��F ��@��  �Ẻ��F �E��5��F �u��;��F �y� �E��E�FO���� �M��u��E̋5��F �M��M��M�벉�$�  ��$�  ���F ���F ��$�  ���e����d�F ��F ��F �1����  ���  �=(�F ���F ��F �Ƌ��  ��F ���  ���F ���  ���  �=�F ���  ���  �p�F ���  �6  ���  �5��F ���  ��(Q�L�F ��(���V������F �J<�5��F hX  jdj R�g  S���  ����  �@�F ��)�;�  �g�����    V���  �405��F ;u�ʼ �=,�F � �F ���  �]�=��F Q��F ���  �5��F ���  ��,Q�L�F ��(���������F     ��F ��@jh�  �5��F �9  É��F ���  ��F ���F ���   ���  �=d�F =��F =��F �%��  ��    ���  ���F �p�F ���F ;��F �4�  ���  ���F �5t�F ���F �=4�F ���  ��$�  �(�F �5p�F �d�F �=��F ��$�  ��$�  �d�F �����5�F ���  �L�F �L�F     �5��F �   Ë5��F �N<�Q|�qxh�  jd�5��F �5��F h�  ��  ��5��F ���  �L�F �5��F P���F �U ���  �ҋ�F ��F �=�F ���F ���  ���  ���������  ���F     ���  ��<Q�L�F ���F ���F ��<�������@  5��F 5��F �%��  h�  �  Ët�F ���F ���F ���F ���F ��F �4�F ����F ���F Q���F ��F ���F ���  ���  ��F �x�F ���  [���  �4�F ���F ��|  ���  ���  ��|  ���  ��  ��<  �<8=��F ;=��F ��) ���  �@�F �d�F ���F ��  ���F ��$�  ��$�  ���F �l$t�\$p��F ��$�  ���F ��$�  ��$�  � �x�F A��$  V�5x�F )�F��V��H�5�F ��d������  ���F �L�F �M������  ��󤉅�  ���  ��F S�W  É��  �d�F %��  �=d�F ��+�$�  ;@�F ��������  �,�F ��    ���  ���  �0��F 9����  �,�F �=�F ��F �}���L�F �,�F ���  ��F �5��F �L�F �;�����F ���  j �=�F �}���L�F �M����  ��F �5��F �L�F �������Q�L�F ���F �L�F ��P������    �5��F �
����=8�F ��$�  ��$�  �=d�F ��$  P�5��F �-@�F ��$�   ���F ��$�  ��$�  ��$�  ��$�   ��$�  ���F ��F ���F ���F ���|��H��  5��F ���8  �=,�F �N�~���  �^���F �N ��F ���F �V$��F ���F �V��F ��$�     ���  ���  �,�F S�  V�t$V�I������Yu������ 	   ���^�W�t$j �t$P���D �����u���D �3���tP�����Y�����΃�����̈́F �ƍ��D�� ���_^�jh��D �h�  �];��F sx�����<�̈́F �Ã��4�����D0tXS�����Y�e� ��D0t�u�uS�5������E���)���� 	   �'����  �M���M���   �E��!�]S�4���Y������� 	   ������  �����  ��>{  �@d;�{F t職  �x(~j�t$P誼  ��Ë@H�L$�H����{  �@d;�{F t�G�  �x(~h�   �t$P�m�  ��Ë@H�L$�H%�   ���z  �@d;�{F t��  �x(~j�t$P�1�  ��Ë@H�L$�H�����d  �t�F ���F �4�F ���F �B%�   =�   �o����t�F ��F ��F ���F ���F ��F �4�F �t������F @=�   jh�  �5|�F jd�54�F �y����ыQ|�qx5��F ��������N�~�@�F �N��F �F ��F ��F �F$��F �n-��F ���F    ����  ��$�  ��$�  ��=,�F � ��F �� �F ���  �,�F ���F     ǅ�      h�  j �,���Ã��������  ��8  ����  �5�F ��+M�;��F ��  ����    �<�F jdj�g  Ë\�F ���$X  �L�F ��$(  P���  �U �L�F �ҋ��  �L�F �U����  ���  ��X������X�F �,�F j �5��F �P  É��  ���F ���n���  �=`�F ���F ���F ���  �΋=0�F �4�F ���  �E����F �$�F ���  ���  ���  ���  �=��F ���  �=0�F �����  ���  �=L�F ��F ��PP�L�F ��@�/����54�F ���  �=T�F �} ���  �  ���F �}���F P�]����   ���F Y���F ��<  ���F �-��F �pAՋ��F �5��F ��0  �5��F ��(  ��W����=�F ��$  ��F �@�F �ŀ   ���o  hX  Q�5��F ����Ë-��F ���F ��$�  ��$�  ��$�  �l$p��$  ��$�  ���F ���F ��$�  ���F �8�F �=��F ��$�  ��$�  ��$�  ��$�  �5p�F ��$�  ��$   �5��F �l  �[��   ���F ;�F �Y� h�  j
�  �P��@�$�F W��)�F�ދډ�F �΋��W�=$�F ���F SQ�\�F ��$�F ��R�M  ���5��F �5��F 5��F 5��F �%��  �5|�F �ȉ=\�F ���  �=��F �u��=�F �=\�F ��x����������  ���F �5��F �I�����@Q���F R�U�)�B�ʋ΋ʋ։��F ��W�=��F ���F S�\�F ����F ��S�8�F �  ���  �=��F ���F � �F �=$�F ���  �0�F ���  ���F ��\�  ���F ���F ��$�  �L$|�=��F ���F ��$�  ��$$  ���F ��$�   ��$�  ���F ��$�  ���F ��ň   ��T����jh8�D �V~  �E�P�E �}�P�E s"�e� �E� ��t���3�@Ëe�M���E����Z~  �jhH�D �~  �E�X�E �}�X�E s"�e� �E� ��t���3�@Ëe�M���E����~  Ë��F ǅ�      ��  ���  P�5��F ��   Á-��F �pAՁ�$�  W����,�F ��  Vh�  �5��F �5$�F ����É�F �L�F �5�F P���  � �D ���  �5T�F ��t�����F ���F �H�F ���  ��x����<�F �H�F ����T�F �T�F �E �T�F �������F �<�F �5��F j
�5��F �o  Ë5��F �5�F �5��F j�m  �I$��F R�d�F �R��  ��$�     ���y ���  ���  ����  ���  ��+��  ;$�F ��  �8  P��x������]����(�F �L�F �5��F P���  ���   ���F ��Pj �5��F �58�F ����Ë�@  ��F ��F �����  ��0  ���F ��(  ���F ��<  ���F ���F ���F ��,  �8�F ��<  ��0  ���F ��$  �=��F �5��F ��,  �5��F �}�=��F �5��F j S�  É�  ǅ�      R�5��F �5�F �5��F �y  ËN<�i|�qx5��F ����  ��$�  ��5d�F �5,�F ���F �d�F �K�S�[���  �d�F �[ ��F ���  ��8  � V���F �5�F ���F ����  ��,  ��8  ��0  ��8  ����4  �A  ���F     � �F ��R�L�F ���F ���  ���  ��$�  �L�F ��0��  ���F ���  ��(�  ыQ|�qx5��F ��������=,�F �N�n�~���F �F ��F ��F �N$��F ��$@  �N��F ��$�     ��?� ��$<  �5��F ��5,�F � �-��F �pAՉ��F ���F ���  ���F ��,  ��<  ���F ��W����=��F ��(  ���F �=��F �=@�F �ŀ   ��x�����J<ыQ|�qx5��F ����  �=,�F �N�~���  �F��x  �F ��F �n$-��F ��F �V��F ��$X     ���j ��$�  ��$�  � ��D�]  U���� {F j�E��E�Ph  �u�E� ���D ��u����
�E�P��  Y�M��u  ��j8h �D �x  � {F �E�3��}̉}��E��]��}ċE;E�s  �M�QP�5X�D �օ�t �}�u�E�P�u�օ�t�}�u�E�   9}�t���t����u�N�  Y��F�u���u�9}�uWWS�uj�u���D ���u�;�tX�}��6������|  �e�܉]��6PWS��  ���M���3�@Ëe�警  3�3ۃM���u�;�uVj�w  YY��;�u3��   �E�   VS�u��uj�u���D ����   9}t WW�u�uVSW�u�D�D ��tf�E�E��^9}�uWWWWVSW�u�D�D ��;�tCVj��  YY�E�;�t2WWVPVSW�u�D�D ;�u�u��  Y�}���}��t
�M���]�9}�tS�  Y�E̍e��M��  �+w  Ë��F �5��F �58�F �5��F W�5$�F �Q�����,�F ���F ��@  ����  ��H  ��+�$�  ;�$�  ��  ��    S���F ���F 9��� ���F �,�F [���F ���  � �F ��<P�L�F ���  ��$�  �L�F ���  ��F P���F � �F �e_���F ;d�F ���  ��F � �F �5�F �5��F ����,�����ǅ�      j�   Ë��F �J<V�e�����l  ���  ����  R��)�;�F ��  ��    �5��F �415��F ;5��F �� ��8  �,�F �-��F �pAՋ��  ���F ���F ��<  �0�F �X�F ��W����=�F W���F ��F �@�F �ŀ   �� �7����=,�F �5$�F j<�5��F ����É��  �t�F ���  ���F ���������F ��EE�����  ��p  ���F ��l  �Ë�F � �F ���F ��l  ���_������  �$�F ���  ���  �u�t�F �Ћ=\�F ���  ���  ���F �H�F ���  �0�F ���  ���Ą   �[���F �Ẻu؋]Ћ=H�F �ы5��F �5��F �5��F �5�F �w
  �����F     �58�F �5�F jS�5��F ������[���  � �F ��<R�L�F ���  ��$�  �L�F ���,	  �=��F �
  ��p  �������F     �5��F �<�F �5@�F �}ԉ]ȉx�F ��l  �E؉��F �Uċ��F �U��   ��!  ���%��  +��F ;E��'" ���6	  �]��u؉�l  �5��F �]ȋU���58�F �n ��h  ��QP���F � �D �$�F ���F ��`  ��p  ��\  ��x  � �F ��\  ����D�����5��F ��8  �P�F Z���F �ŀ   ��������=�tF  V�5�F u3�^Å�SWu95�F tQ��&  ��uH�5�F ��t>�\$��t6S�Q�  Y���%P�F�  ;�Yv��<8=uWSP�t�������t�����u�3�_[^Ë�D8��8 V��tW���t�9��F��8 u�_^�U��QSV��3�9U�U�t5�9�7vj
�[����0�F�	���~��w��7N���N�@;�r��.;1s(N�V��tj
�[�����0�E��N���u�E�)��^[��U������ZV�uW���   ��  ��Muti��%tV��tBHt0��t!H�#  �F�jY������  QX�~  �u�Fj�g�V�u�T�h��  �V�u�T���  �� %����  �u�Fj�1��S��   HHteHHtPHt+H��  �F�jdY���uj��k�d�Z������Y�  �uSWVj�u�  �����o  3��k  �F��ujY��H���N9N}3��   �Fj�^��;���   �   �u�j둃�m��   ��   ��atxHtfHt'Ht���  �u�F@j�]����u�Fj�P����} �uSWVt,j�u��   �����X����; �O�����  ���&���j �ҋV�u�T�8�   �V�u���   �F@�uj�������pt\��tIHt,HtHun��  3�9V ����F �O�u�F�jdY�������} �uSWVtj����j �����u�F3�B�����~�U���   ����   �ϋ�����3�@_^]�j8h�E ��n  �E3�+�tH�Et���   ����   �	�E���   �E��M���   �  �}�,�D u���D �EЋ]f�Sf��lf�U�f�SfBf�U�f�Sf�U�f�Sf�U�f�Sf�U�f�f�U�f�u�VV�u��U�RV���   �ЉE�;���   �ủu�������r  �e���}ȃM���3�@Ëe����  3��M���]3�;�u�u���}��Y��;�tc�E�   �}��u�W�u��E�PV�E���   �U�H;�~ �u�M�> v��]܊���E��H���}� tW�0  Y3�@�e���m  Ë]�E����t�}�u��]�? t��E� 3҉U؋E�@B8t��E��Ƀ�d�V  �  ��'��   ��At��Ht[��Mt"��a�W  h�E �]�S�eq  YY��uV���e��ItIt#ItI�,  �E�B�#  �E�b�  �E�   �E�m�
  ��ItIt��  �E�   �E�H��  h�E S��p  YY��u���]��E�p��  U����!  �E��M����  <'tJ�Ћ]�[H�DS�t��v�M�A�9 ��  ��������E�����@�E��� ��u���  �E��  ��ItIt#ItI�J  �E�A�A  �E�a�8  �E�   �E�d�(  ��h�
  ����   ����   It)���  ��IItII��   �E�Y��   �E�y��   �E�{���   ����   ��uq�? vl��ы]�[H�DS�t�?v@�8 ��   ��
���� ����=�? v8�ы]�[H�DS�t�?v@�8 ��   ��
������@����uËE܉E��   ��ItIt	�9�E�   �E�S�,��ItIt	�"�E�   �E�M���ItIt	��E�   �E�I�E��t#�u��u�u�u�ߋ��f�������u�3������M���Ћ]�[H�DS�t�?vA�9 tً�������A�M���E����������������$�      j
h�  j��  É�5��F ��$�  �L�F �5��F P���F � �D �\$ ��$�  ��$�  ��$�  ��$�  ���<��딉-��F ����F ��F ��F �(����  �l$����e��]��5��F �u��]�;]����  ���F �$�F �]���  �5,�F ���  �E�ǆ�       ���   �E����   �E�ǀ�      �uԋ�l  �C<؋H|�Pxڅ��� �}؍=,�F �B�Z�r�z �$�F �EЋEԋ�l  ϋB$ȋJ���F �}̋}ԋ�l  ��5��F �E��}�����F�-��F R��)�B�� �F ��Q�X�F ��$�  �L�F ��$�  ��$�  �L�F �X�F �5��F ����$�  �=��F �\�F �5��F j�;�����k� �5��F ���F ���  �=�F ��h.  j ��l  �L�F �,�F h�c  j��h  �L�F P��F �,�F ��d  jB鐠 �Uȉ��F �5��F �]ЋыE̋5��F �5��F �uȉ5�F �{������F ��<  ���F �ŀ   ��$�2����$�F �}��=x�F �G\����F ���F �=��F �   �� �5X�F �ǉ]��U����F �5��F �]ȋUċM؉��F ���F �}ԋUԋu��R����b����5 �F ���  �L�F Sjj hX  Q�  �jh�D �@g  �u�u�u���uF3��}���we�=�`F uG������u�]�;ŖF w3j�v��Y!}�S����Y�E�M���J   �}��t�u�j W�j�  ����u:Vj�5��F ���D ����u%9=��F tV�v��Y���v�����uj��t��YË���f  ��U��SVWUj j h(�@ �u�O ]_^[��]ËL$�A   �   t�D$�T$��   �SVW�D$Pj�h0�@ d�5    d�%    �D$ �X�p���t.;t$$t(�4v���L$�H�|� uh  �D��@   �T���d�    ��_^[�3�d�    �y0�@ u�Q�R9Qu�   �SQ��zF �
SQ��zF �M�K�C�kY[� �E�@�U��d�F �= �F �}�)�G�׋։M��ϋ=d�F �ы��=d�F ���F ���E��=`�F �M��H�F ����F ��}�룁�  �d�F S��F �L�F �5��F P�\�F �Mԋ�P  �x�F �ҋ��F �u��M��$�F �m����F �= �F ��$�  �-��F ���  ��  �����S���  ���  ��\  ���  ��8  ���9  �5d�F ���  ���%  ��$�  ��x  �L�F �,�F ǅp      �5$�F W�����Ë50�F �0��F ;\�F �� �x�F ���F �p�F ���  ���  �$�F ���F �=\�F �]�t�F ���  �p�F �ދ��F ���  ���F ���Ą   ��������R�T�F ���  ���  �����N������F ���  ��F ��F �%��  W�5��F Pj �   Í�    ���F �5\�F j �5��F ����É�$�  V�a���Ë|$��%��F ����D$����F ;�1����-D�F �����F �}ԉ��F �E��U��
���F     �}ԉU؋��F ;U��� ���F ��F �E��E�Ћ(݉l$����F     �|$ԉD$��D$�� ���c����|$����F ��F �\$ԋ��  ���F +��F ��F �D$����F �X�F ���D$���F �Z�=��F �,�F �5H�F �M �5t�F ��F �E��E �,�F �E�5P�F P�Ã��   ���F �EЋ5P�F �Á%(�F ����(�F Y;��	  ���F ���E؋M��E�}ȋ5��F �M̋}܉U����F �2  �&  R�,�F �-t�F ����F �}��E�    �0�F ���  W�G0    �x�F �� �G �=,�F �E     �E�    �} G��i   ���  ���F ��  �] �C���   ���   t���F ��  �!���F �] ���F ���F ��  ��[�M �U����F ���F ���F �]�] Y���F ���F �]�5��F X�E���F R���F ���F ���F �M���  ���F ���5����E��   �E�    �U�P�5��F �U��É}܋}�;=��F �����}�}؉��F �M���L�F �E��(�F     �0  �M؋U܋=��F �Eԋu �-H�F �D$�t$؉-t�F P�\$؋\$��\$�D$؋5P�F ������g������F ���`����U�B�U�M��=T�F �}ȋ��  �M����}�+=T�F G�ǋT�F �ωu����}�����]������F ��5��F ��  �5��F �H  �V�t$�F��t�t�v�  f�f��3�Y��F�F^�jh�D �j_  �e� j j�,Q  YY�3�@Ëe�M��j���D �; {F u�������5��F �U����F �U��E��5��F ���F �ËM������������F ���F �5P�F �Ë��  �(�F ���F +��F (�F �EԉUЋ��F �E�댍=,�F �=��F �_<��{|�M�Kx��F ���%� �E�,�F �A�Y�E��A�5L�F �q 5��F ���F �I$��F �U܉��F ��   �u�V���D �u�P�E�� �D �u��p�F ���F �}ȉ0�F �]���  �  ��F �= �F =��F =��F �%��  ��F �E����F �=��F �ŰL�F �]Ћ=l�F �U����F �]��=t�F �mċt$ȉl$̉t$Ћ5L�F �D$����F �t�F �=�F �  ���F �S��F � �F ���F �E�    �H�F �U��M؉��F �   ��h� ���F �,�F �t�F �ủ=��F �E���   �}�EЉ}ȉ��F �]ċM܋]؉M��]���F �%��  �_V�t$��tT��X{F ;t;({F tP�]  Y�F�X{F ;At;,{F tP�@  Y�v�X{F ;pt;50{F tV�$  Y^�+t�F ;E���� �E���e����F �M܋M���F ;E���h �E�ǉ��F �U�M؋��F ���  �I�E��Eԁ}�   �� �5`�F �t�F �}��]��u܋=��F �]ĉuȉ=��F �D�F �M��&�U؋��F ���F 뉉\$ĉ��F �\$���M����M܋`�F �D�F �]Ћű=��F �E�L�F �]����F �m��l$�L$ȋt�F �\$ċ|$؉|$��l$��l$؋=��F ���#���jh �D �x[  �u��tX�=�`F u@j�nj��Y�e� V苷��Y�E��t	VP觷��YY�M���   �}� u�u�
j�i��Y�Vj �5��F �8�D �O[  ÉU����F ���D �u�P�E�� �D �M؉5��F �=|�F �] �`�F �UԋűEЁ�  �!  jhp�D �Z  3�95�F u5�E�P3�GWhl�D W���D ��t�=�F ����D ��xu
��F    ��F ����   ;���   ����   �u܉u�9uu���F �EVV�u�u3�9u ����   P�u���D ���}؅���   �e� �?�Ã�����^  �e��u�Sj V苕  ���M���3�@Ëe�蹈  3��M���}؅�uWj����YY����tg�E�   WV�u�uj�u���D ��t�uPV�u���D �E܃}� tV�
���Y�E��n�];�u�p�F �}��u�=��F S�m���Y���u3��D;�tj j �MQ�uPW����������t݉u�u�u�u�uS���D ����tV����Y�Ǎe��MY  ÉUԋ�B��  �EЋ�)�@�ȋÉŰщuȋ��=|�F �]Ћ�  �}ĉM����F ���  ��  S�������F �uЋ��F ��뙉��F V�u܉��F �`�F �D�F ���F �C0�[�,�F �E�}�
   �W����m��,�F �Ët$�-h�F �t$�L$�|$���D�F ���F �5d�F �G���F �Ë5(�F u�u؋%��  �M؉}̋U�}܉Uȉ5d�F �5��F V�ʋ5P�F ����   �D$�X���F ���F R�,�F �D$��t$����   �t$���D 3�@� jh@�D �W  �P�F ��u7�=ȭF t$h,�D ���D ��th�D P� �D �P�F ��u
�ݯ@ �P�F �e� �u�u�ЉE��$�E� � �E�3�@Ëe�}�  �uj���D 3��M���dW  �%��  +E�9�������,�F �E��U�M؋É��F �e��] �u܋u��L�F ;M���� �4�F �M؋4�F �`�F �M�����U��SVW�}���E3�9U��    �Et	�M�E�1j[f�8"u�}3Ʌ���j"Ë�Y����tf�f��f��f��t;��u�f�� tf��	u���tf�f� �e 3�f9��   f�f�� tf��	u���+���f9��   9Ut	�M�E�1�M�3�G3���Bf�8\t�f�8"u*��u#�} t�Hf�9"u���3�3�9Mj��[�M���t��tf�\ �M�Ju�f�f��t+�} uf�� tf��	t��t��tf��M���v�����tf�& �M��$����E;�_^[t��E� ]�U��QQSVWh  �t�F 3�VWf�=|�F ���D ��F ;ǉ5��F tf98��u�ލE�P�E�PWS3��K����}��E��x��P��d��������u����&�E�P�E�PV��S�����E���H�ܭF �5�F 3�_^[�ÉE�]��E�    ���F �] R���  �d�F �M ���F �}��5P�F �M��Ë}�^�=��F �5��F �U܋d�F �U��   ��E��    �������M؋Ë5P�F �M��M��M܋����S�L�F �[<L�F �k|R�SxL�F ���C����-H�F P��,�F �B�Z���F �ZP�B L�F Q�J$L�F �(�F �JL�F �U��������  �,�F J�  � � Rj
�  Ë5��F ���   �ڋ�|�����x�����  ��ǅH     ��F     ��H  ��t�����  �=�F ��H  ��  ����  ��@  ���  ���  jǅH      Z��t������  �ڋ���Ћ؋l�F �Ζ  ��B���$�F    j �$�F ǅH      ��t����N  U��$t�����  � {F ���   SV���   3�W3�;Ő}F t@��r����;��}F �  ���F ����   ;�u�=PF ��   ���   ��   h  �E�PR���   ���D ��u�E�h`�D P�_[  YY�}���P�Bu  @��<Yv"��P�3u  ���E���;j�h\�D W�|�����W�u  ���}F ���u  �DY��Y����eV  ��h E S��Z  WS�[  hX�D S��Z  ���}F S��Z  h  h$�D S�x  ��,�(R���   P���}F �6�t  YP�6j��p�D P�x�D ��t������   �'���_^[�Ō   �á��F ��t��u*�=PF u!h�   �h�����F ��Yt��h�   �R���Y�U��$`�����   � {F W3�9��  ���  �}��}�u3��  ���  S���  ����V�4���̈́F ����D0 tjWW���  �@  �����@���   9��  ���  �E��}���   �M�+��  �E��}�;��  s'�U��E��A��
u
�E�� @�E��@�E��}�   |ы��E�+�j �E�PW�E�P��40�x�D ��t�E�E�;�|�E�+��  3�;��  r�����D �E�3��E�;���   9}�tZj^9u�uG����� 	   �����0�hW�M�Q���  ���  �0�x�D ��t�E��}��E�����D �E���u��Е��Y�*��D0@t���  �8u3��螕���    蜕���8����+E�^[���  _�����Š  ��jh��D �NO  �];��F sx�����<�̈́F �Ã��4�����D0tXS�ʹ��Y�e� ��D0t�u�uS��������E������� 	   �����  �M���M���   �E��!�]S����Y��ߔ��� 	   �ݔ���  �����N  Ã�������,�  �l�F CjǅH      X��H  �t�H�߼  P��H  �������@��t����7�  �؉�H  ���W�5�F ��������  ��(���@_�5\�F �Ѓ���   ���  ��   jhp�D �N  �];��F ��   �����<�̈́F �Ã��4�����D0tmS�~���Y�e� ��D0t1S�)���YP�t�D ��u���D �E���e� �}� t蹓���M�覓��� 	   �M���M���   �E���]S蹸��Y��~���� 	   ����M  �P�,�F �$���Vǅ�     �th���  ����   �,�F ������ ���   �i  �� ����7  �U	  �� ���  �  �,�F �� ���   ��
  A�-  �,�F ��(�����I���(����Ћ��  �@���  ��F �Ћ�F �o����,�F �5\�F ��(�����v�V�Ћ5\�F ��F �,�F ����@�� ���   �  �� ����7  ��  �� ���  ��  �� ���   ��  Y���  B��������F �5�F Q���  �� �����F ��(�����������  ���  ���  ���F ^��<�  �= �F �=,�F �F ���$  S�����F    �\�F ��$����-d�F ��F �L$��=��F ��$�  �= �F �݋���   �#���U��QQSV3�W�=�F �u��;�tb�D�D VVVVj�PVV��;ƉE�tZP�[��;�Y�E�tLVV�u�Pj��7VV�Ӆ�t1�E�VP�M�����YY}9u�t�u��o���Y�u����;�u�3�_^[���u��S���Y�����j8hH�D ��J  3�9�F u8SS3�FVhl�D h   S���D ��t�5�F ����D ��xu
��F    9]~�M�EI8t@;�u�������+�E��F ����  ;���  ����  3��}ԉ]ȉ]�9] u���F �E SS�u�u3�9]$����   P�u ���D ���u�;���  �E�   �6������iN  �e�ĉE�M���3�@Ëe��x  3ۉ]�M���}ԋu�9]�u�6P�Y��Y�E�;��`  �E�   V�u��u�uj�u ���D ����   SSV�u��u�u���D ���}�;���   �Et-9]��   ;}��   �u�uV�u��u�u���D �   �E�   �?������M  �e�ĉE��M���3�@Ëe���w  3ۉ]��M���}ԋu�9]�u�?P��X��Y�E�;�t@�E�   W�u�V�u��u�u���D ��t!SS9]uSS��u�uW�u�S�u �D�D ��9]�t	�u�����Y9]�t	�u������Y���[  �]�3��]�9]u�p�F �E9] u���F �E �u�T���Y�E����u3��!  ;E ��   SS�MQ�uP�u �l������E�;�t�SS�uP�u�u�L�D ���u�;���   �]�������mL  �e���}�VSW�m�  ���3�@Ëe��v  3�3��M��;�u#�u��W��Y��;�t1�u�SW�7�  ���E�   �u�W�u�u��u�u�L�D �E�;�u3��&�u�u�E�PW�u �u����������������u�9]�t#W�����Y��u�u�u�u�u�u�L�D ��9]�t	�u�����Y�ƍe��QG  ���$  R�  �J�	  S�,�F ��� ���  [��0�ҋ�F �5�F �d�F R���  ��(����� ���^�d�F ���  ��(�����@�S�,�F ��v�W��(���������� ������  �,�F �D  ��F ��F �򉅬  ���F ���  ��F B��(����|  ��Y�  �6  ���$  Y�Љ�(�����F �x  �	��(����R�������A�� ���   }��� ����7  ��  �� ���  ������� ���   �c  �������Y�  ���  �,�F �v���@R  �$�F � �F ���  ��F ���  ���  ���F ���  ���  ���  ��F �ˉ5��F � �F ���  �$�F ���F ���  �Ѓ�@��  W�Ћ�F �������(���_���u�,�F R��(�����R���(���S�,�F �  �=l�F ��F �5(�F �=�F �x�F �����  ��F @�=l�F ��[���  Z���$  ��(������AA��F �5�F ���F R���  ��(����� ���^���F ���  ��@�T������"  ���$  S���  ���$  ���  �����[���� �����<�������  �h�F Z�0�F �h�F �h�F ���,  �50�F �!  P���$  �=��F �� ������"  ���$  ���  ���  ���"  ^Y��H�{�������_���  �� ������F ��D�[� ����-(�F ��$�  �x�F ����   ��H�6��@$  j���$  ��F ��%  ���F �l�F R��$�����#  Z�n��)�j
h�  ��  Í,�F ��(�����v���(�����W�=0�F �@��f����=(�F ��_�5(�F �?��Y�S����5,�F ���$  �0�F    Q�t��,�F �50�F ��������,�F �������F ���  ���  ��F R��F ��(����5�F ���  �=@�F �=�F ���  �=@�F ��H������F �5�F Q��F �� ������  ��(�����������  ��F ^��D��������F ���$  ��L#  ���"  Z���  ��(�����L#  �-��F ��$�  ����   ��L�������F ���F    ���$  ���$  ���  �`�F �ȋ��F �=��F �=��F �=0�F ���!  ���   �������5,�F ���  ��(���ǅ�     ���"  ��F ��F ���  ���"  �ʋ��"  ���  �0�F ���  �� �O����R���sM  �=��F P���F �������p�F ���  ���  ���  �=��F ��F ���  �Ѓ�����[�Љ50�F @�Ѓ���������  ���F ���  ��  Sh�  �6   Ë�I���S�,�F ��  ���#  ���  ��  F[���   �  ���   �  ��I�V����F X���  �,�F �d�  ��  ���  F�Ĩ   �c  ���  ���  ���  ���  ��  �5`�F �5��F �Ĉ   �.  ���  �,�F ��<����5��F �5�F Rh�  ����É�F �,�F h�  �   ���5��F ��  É��F �,�F ���#  ���  ��  ���F S���  ���  �h�F ���F �`�F �h�F �Č   �  �$�F �؋�$  ���  �ȉ5��F ��=��F �=$�F �=�F ���  ���  ���  ���  �=��F ��  �|�F �5��F �\�F �ˋ�F �Ę   �  �	  ���F �,�F ��W���V���"  ��X���  �,�F �M�  �@�F ���  ��  �Ĩ   �  ���F �,�F �$8  ���   VW�5��F j
�G	  �R��F ��`$  �-��F ��$d  ��$   �-��F [�5�F �\$����F ��F �L$���$�  ��F ���P  �Ĵ   �1  U��SVW�}3�;�t9]t�:�u�E;�tf�3�_^[]Ëu9^u�M;�tf��f�3�@���NH���DA�t<�F(��~"9E|3�9]��Q�uPWj	�v���D ��u�E;F(r(8_t#�F(�3�9]��P�ujWj	�v���D ��u��_���� *   ����f����3  �@d;�{F t��o  �t$�t$�t$P������ËD$f�8 ��tBBf�: u�V�t$f�f�
BBFFf��u�^ËL$�T$f�f�AABBf��u�D$���  ��  �,�F jd��  ���F    ���F ��|  �`�F    ǅl      ���F     ���  ���F ���  �5��F ���  ��  �5��F ����Ë�  ���F j ���  �=��F Z�=��F ��l  �=4�F �=��F ��  ���  �5��F �5��F ���  �Ę   �$������F � % ���	����F �C���  �P�F ���  ���  ��  ���  ���F ���F ���F �5T�F �5P�F �5��F ���F �5T�F ��T������l  �=,�F ��l  ���F P��  ���  V�������5��F ���  �5��F ��l  ^���  ��l  ���  ���   �N������F ���  j ��  ���F V���F ��������l  ���  �5��F �5��F ^�İ   �����kp �j�58�F �5��F j P�  á�F 3҅�u��E f�f�� w	f��t'��tf��"u	3Ʌ�����@@��f�� w
@@f�f��u��-�  t"��t��tHt3�ø  ø  ø  ø  �Wj@3�Y�ȃF �3����G �X�F ���F �paF ���_�U���  � {F �E�V�E�P�5��G �X�D ���   �  3�������@;�r�E��ƅ���� t6S�U�W�
��;�w+�A�����������    �˃��B�B��u�_[j �5��F �������5��G PV������Pj����j �5��G ������VPV������PV�5��F �r���j �5��G ������VPV������Ph   �5��F �J�����\3�f��E������t��ɃF ���������_F ���t��ɃF  ��������ƀ�_F  @;�r��D3���Ar��Zw��ɃF �Ȁ� ���_F ���ar��zw��ɃF  �Ȁ� ��ƀ�_F  @;�r��M�^�>�����jh��D �u8  j�{G��Y�e� ��.  ���}��w`�u�;54�F t"��t�uV����Y�4�F �G`�54�F �u���M���   ���Z8  Ëu�j�lF��Y�U���� {F SV�u3�;�E�W�T  3�3�9� zF te��0B=�   r�E�PV�X�D ���!  j@3��}�Y�ȃF 󫪉5��G ���F ��   �}� ��   �M�����   �A����   j@3�Y�ȃF �R���]䪍�zF ����)�V��t&����;�w�U䊒�yF �ɃF @;�v�FF���u��E���}�r��E���G �X�F    ������zF ��paF �����F ��_��ɃF @;�v�AA�y� �I���3�A����ɃF @=�   r���b������F �X�F ��X�F 3��paF ����9��F t�e�������3������M�_^[�?�����jh�D �v6  �M��j�xE��Y3��}��=��F �E���u���F    ���D �+���u���F    ���D ����u���F    ���F �E;��G ��   �54�F �u�;�t9>th   ��E��Y���u�;�t�u�����Y�E�;�uo�>���G �F�X�F �F���F �F3��E��}f�EpaF f�LF@��3��E�=  }��ȃF �L0@��3��E�=   }���_F ��0  @��54�F �}��u;54�F tV�����Y��}��M���	   �E��w5  �j�C��YÃ= G  uj�����Y� G    3�É��  h�  �5��F �5|�F �����Q�,�F ���  Y���F ��������F ���  ��������F �������릉��!  ���  ���  ���#  ���  ���  �É��F ���  ��F �=��F ���F ���F ���  ��4�N���ZX���F +�  ��@JS���t	  ��(������
  ��	  ��t	  `T ���$�����0���ȉ� �����t	  BX+=��F ω� 
  ��t
  #��F =��F �@�F �� ���ZX+��
  ������=<�F 3��  ���  ��F ���  ��F ��F JX���F ���F �ϋ�x
  ��F ������=d�F ��  ���  �����ZX=��F �M�5��F ��`������   �Y�������,����A��X
  ��(����Y���   �A��������  �y�=�F ��p����]���h�����x�����4  ��L  ���
  ���
  �5�F ��l�����`�����X�����P�����H�����D�����@����|�F ���F ���F �5�F ���F �=��F �-��F �
  UV�5��F W3�3�;�u����   f== tGV��.  Y�tFf�f;�u��   SP�'B����;�Y��F u����\�5��F �/V�.  ��Gf�>=Yt�?P��A��;�Y�t9VP����YY���4~f9.u��5��F �e����-��F �+��tF    3�Y[_^]��5�F �@����-�F ������A@t�y t$�Ix��������QP�V��YY���u	���U��V����M�E�M�����>�t�} �^]��G@SV����t!� u�D$���L$������C�>�t�|$ �^[�U��$,�����T  � {F ���  3��E��E��E����  S�3Ʉ���  VW����M�G�}� ���  �p  �� |��x�����E ���3���� E j��Y;��E��,  �$�O�@ 3��M���E��E��E��E��EĉE��  �Ã� t;��t-��tHHt����  �M���  �M���  �M���  �MĀ��  �M��  ��*u'���  ���  �@����E���  �M��]��  �E��ˍ��DAЉE��{  �e� �r  ��*u$���  ���  �@����E��R  �M���I  �E��ˍ��DAЉE��4  ��It.��ht ��lt��w�  �M��  �M��
  �M� �  �<6u�4uGG�Mŀ���  ��  <3u�2uGG�e����  ��  <d��  <i��  <o��  <u��  <x��  <X��  �e� �{F �e� ���DA�t���  �u����2����G���  ���  �u��������S  �Ã�g�X  ��e��   ��X��   ��  ��C��   HHt`HHt\���  f�E�0u�M��M����u�������  f�E����  �@��E��D  ��u�܁F �E��E��E�   �  �E�   �� �M�@�}� �uȉu���   �E�   �4  f�E�0u�M����  f�E����  te�@�P�E�P�T����YY�E�}[�E�   �R��ZtX��	t�H�2  �M�@�E�
   �]ľ �  ���3  ���  ��Q�����  �H  �@��E��E�   �EȉE���  ���  ���  �@���t-�H��t&�E�� �M�t�+����E�   �  �e� �  �؁F �E�P�   u��gu@�E�   �7�   9E�~�E���   9}�~ �E�]  P��<����Y�E�t�E�����}����  ��u����u����  �@��E���P�E�VP�M��{F �}ă���   t�}� uV�{F Y��gu��uV�{F Y�>-u�M�F�u�V�O  Y��  ��i���������   H��   Ht^�������HH���������  �E�'   �EIf�8 t@@��u�+E����  ��u�؁F �E��E��I�8 t@��u�+E��^  �E�   �M��EĀ�E�   �����E�Q�E�0�E��E�   �����EĀ�E�   ������M���������  �E� ���  �@�t	f�M�f���M���E�   ��  ���  �� ���  t��@t�@����@�����@�@�u�3���@t��|��s�؃� �ڀM��uċ؋�u3��}� }	�E�   ��e���   9E�~�E����u�e� ���  �E��M������t$�E��RPWS�rd����0��9�]��؋�~M��N�̍��  +�F�E��E��u�t�΀90u��u�M��M��0@�E��}� ��   �]���@t&��t�E�-���t�E�+�	��t�E� �E�   �u�+u�+u���u���  �E�Vj �������u����  �E��M�������Yt��uWVj0�E��������}� tJ�}� ~D�E��]��E��M�3�f�P���  P�{P��CYC��Y~-���  P�E����  �]����}� Yu���u��M��E��F���Y�E�t���  �E�Vj �
������}� t�u�������e� Y���  ����|���_^���  �E�[�������  �Ñ�@ �@ �@ j�@ ��@ ��@ ��@ ��@ �6`  �h�  �  ���  h�  �������l  ���   ���  ��@%  R��@����(�F ���F Z���� ������L$���   �l$�����F ��  ���  ȉ��  ��F ȋ�X  +��F ��|�����x����}���   �꧓�I��t�����|���+X�F �%T�F ��$8�����$,�����$(�����$$�����$�����$�����$������F ���F �=h�F �5��F ���F ���F �-��F �%��F ��F �x�F �-�F �5��F �=�F �3 �F ��<�����H	  ӈ
  ��,  Po�W�X�F �F ���F ��<������
  ��8����<�F PX�0�F ��	  #��F ��8���b�j���4�����P  Өh  ��F ���	  �$���h  ��F ��0����M���   �����	  3H�F ��,�����4���rX��F �h�F ���
  Ӫ�  ���F �h�F �������]����p������   �HX��F ��t������F ��t���xX��`  3��F �=$�F ��l����E���   ���  ��d  ����
  ��d  �H�F 3��  ���F ��F ��h����5��F +5��F ���
  =��F ���F ���   ��F 3��  sX��d����=��F #=L�F ��STIx��=�%��%��F �%��F ���F T  ��P����@�F ӆ�  FX���  #5D�F ��L�����H����E���   +��  ���  �Ƌ��  +D�F ��L�����F ���   ��p  ���F 3X�F 3,�F ��DS��HX��<
  ��D����h�F \�F pX���  ��<
  3��F ���F �T�F �É�@������  3��F ���  ���F ���F �)����  j �5��F h�  j�Y  Í,�F ��Iҍ5,�F ���  ���F �B���$  �Y�����  ���  ���  ���F ���  ���	  ���F X� ��@�������F ��\#  ��@����5��F �,�F �I. F��\#  ǅ�     ǅ�      ���  �=L�F ���F ���  �=��F �=L�F ��H�  ���F    ���F     h@  j	�l  Í,�F ��I���  P���F Z��,�F ��+ Fǅ�     ǅ�      ���  ���  ���F ���F ���F ��h�  ��, P�5��F �5��F Q�5��F �\���Ë�$  ��F ��`������   �x�F ���F �-��F �5��F 35��F ���   ���	  �ˉ�\������   ��d���+��  ���  ��K+��\  +t�F �=d�F ��\���+=l�F ~X�NX��X�����|
  �<  ���  ��<  ���F 3��F ��>k����T������  ӆ�  �H�F Ӧ�  �l  ���F ��F ���
  ��T�����%P�F ��I����  ���  ���"  ���  ��,�F ��- Fǅ�     ǂ"      ���  �D�F ���  ���$  ���$  ��`������  ��h�u�i����,�F ��Iҋ�,�F ��* Fjǅ�      ���$  Q��0������  �=��F ���$  �=��F Y��4�jh�  h�  �5��F h�  �I   ��j�   Í,�F ��Iҋ�Q�,�F ��Y  B������Y���i  �
U�����F ����*Z  ��?�����  ���F ���2* �����F    j ���F P���F ��`������F ���F X���F ��d�Z��������R�  Ã����F ���  �$�  9���1 ���  �5��F ���  �5��F �5��F ���  ���  �;��F ��3 ���  ���  ��$�  ���F ���F ���/4 ���  ���  뢋�I�[�����F �5��F �5,�F �UW  ���!  ���  �=��F ���������  ���  ���  ������5|�F �&  ��^+ �����F    ��F     ���F S���F ��F ���F [��H�"�����  �,�F ��I����F ��  ���F ��  S�,�F �VU ���F �5��F �����[�,�F �������F ����F j Q�����É��F �,�F �5��F �#   ���|  �,�F �54�F �5��F j�0  Ëx�F �� �G ǅ�      �<�F     �5��F h�  jd�54�F S��������l�F �k,  ��\  ��닉�  ���  �<�F    �@�F     Y���  ���  �=<�F �@�F �=l�F ��\  ���  ���  �5�F ��   ��4�&����<�F C��7   �z�����F �D�F ��P  �=T�F �=<�F �G%�   =�   �N  �  �H�F �,�F ǀ@     ǅ\      �5�F R����Ë�\  Rjd�����É,�F jdh�  j	W�e���Ë��F �5��F �|�,�F ��[���d  �,�F ��d  ��\  ���$�  ��@  �4  ���  ��d  ���F ���  ��\  ��x  �����54�F ���F �ˋ��  �0  ��F ��A���F �<�F ��+�F @�؋�F ���  �ˉ5$�F �����  �=��F ���F �\�F ��5��F ���5��F V���  �^  �=T�F P�<�F �D�F ��P  ��[��F �=<�F ���5���F ��$�  �=��F ���F ���F ���F ���F �����  W��F ���  �<�F �=T�F �D�F ��|  ���  �$<  ��l  �,�F �x�F �5`�F ��l  �D�F �,�F ��|  �`�F ���  �D�F ���������  ���F ���  �  �=��F ����F ��F �����  �5`�F ���  ���  ���  ���  �=��F ���  �=��F ���  �D�F ���  �t  ���D ��$�  P���  �U ���F �ҋ5�F ���  ���  ���  ���  �=4�F �l�F ���F ���F �<�F �l�F �=�F �=��F �=4�F ���  ��l  ��R���D ��$�  P���  �M���  �ы�F �d�F ���  ���  ���  �5��F �p�F ���F �=H�F ���F �54�F ���  ���F ���  ���h��  �4�F ���  %��  ���  ��+�$�  ;l�F ��  �5H�F ���  �5p�F ���F ��    �54�F �0��F 9��8. ���  ���  �5p�F ���F ���  �=��F ��  �,�F �I��  ��$X     ��� ���F ���  ���  ��\  ����  ��4  ��+��F ;X�F ��  �  �,�F ǅ�      ���F �A<ȋH|�hx-��F ��� �����$�  ��=,�F ���  ���  �A�I���  ���  �@���  �m -��F ���  ��$�  �R$��  ��$�  �qt�����F �=��F �=��F =��F =��F �����  ���  ���  ���  ���  ���F �=��F �54�F �x�F �=��F ���  ���  �=��F �A����=��F �=,�F � �F     �=��F �G<��x|�`�F �Hx��F ��tX�,�F �A���  �y���F �Y���  �Y ��F �5p�F �q$5��F �l�F �A��F ��$�     ��������F     ���F �A<ȋH|�xx=��F ���E����=,�F �=,�F ���  ��   �B�R���  ��   �R��,  �,�F �@ ��F ���  ��   �@$��F ��  ������$�  ���F ��$�  ��$�  �5 �F ��$�  ���������h�F �=��F ���F ���F ��$�  ��������=,�F ���  �	����5��F ���  �5`�F ���  ��$�  ���  ���F ;,�F �~ �d�F ���  ���  �5d�F ���  ���  �#����d�F ���  B��$h  ���  ���  +��F C�ˋ��F �ˉ5�F �5��F ���  ��l  �0�F ���  ���  �=\�F ���F ���  �8�-������F R���F ���D �5��F P���  �M���  �щ��  ���  ���  �=��F ��F ���  ���F ���  ���  ��F ���������$�  ��$�  ��$�  �1����5P�F ��T  ��T  �5`�F ���  ��  ��   ������=,�F ���F �8�F ��������  �����5��F ���  ���  �5p�F ���F ���  �,������F ���F �R��F ���F    ���V  �4�F ��F ��$�  ���F ���F ���F ���F ����  ��)�;�$�  �����u����F �F �F �����  ���F �-4�F ��$�  ��$�  ��$�  �=4�F ���F ��F ���F ���F �=��F ��$�  ��$�  ���F ���F ��$�  ���F ���F ��$�  ��$�  �=4�F ��$�  ��$�  �/��F ;��F ��  �������F @���F �=��F �=��F )�G�ߋًω��  ��=��F ���  ���x�F ���  �=\�F ���F ���  �;���  ���5��F �[���Í@=   �������p�F     j �8�F    ǅ�      ��F     V�8�F �5p�F ���F �5��F ^���  �,�F ���  �=��F =\�F �Mɉ�F ��   �=��F �G<��x|���  �@x��F ���P������F �,�F �H���F �X�h��$�  �H ��F ���F �@$��F �-��F �n����,�F �R��   �X������F     ǅ�      ǀ�"     h�  ��   É=`�F ���  ���F � ;��F �� ���F I���i  �΍5,�F j���F X��d  ���  ��P�   �,�F ��I������F �,�F ���F ���  �@���F �_������F R�����F Z���  ���F �9���4Bj�=�F [��d  �,�F ��L��|�F �����h�  S�  ���k����5��F �   �BY���F    ��\  ���F ��d  ��\  �� 뵉��F �h�F ���  �EH�F 9��F �f �=��F ���  �=P�F ���F � �F �����h�F ��@  ���  ���Q������  ����F �6������  �5��F jh�  �����Í5,�F ǅd     QWj�5��F �5��F �����É�d  ��D�����Y��d  B��,������v  h�  Qj2�   É�D  _B���  ��������d  �5��F �5��F j �A  �U��QQ�EV�u�E��EWV�E��\z�����;�Yu��U��� 	   �)�u�M�Q�u�P���D ;ǉE�u���D ��tP��U��Y�ǋ��������̈́F �����D�� ��E��U�_^��V�t$W����F�t4V�g��V���˯���v��<  ����}�����F��tP�ǳ���f Y�f ��_^�jh�E �1  �M���u�F@t�f �E��S  �V��`  Y�e� V�}���Y�E�M���   �׋uV�a  Y���  N���F ���F ���   ���F ���扅d  �,�F ǅ\      Q��  �U���  �@`;4�F t�����x u]�h0���MSV�/���DtA���t;�������9Uu�A��"��9ut
Af�f��uȋE��+������#�^[]�3���h  h�D �"  � {F �E� �F 3�;�t�M��u�u��YY�M���  3�@Ëe���EHt���D ǅ����8�D ��   ���D ǅ����x�D ��   �M�h  ������PQ���D ��uh`�D ������P�  YY��������P�0  Y����<v%��P�0  �؍�������1�jh\�D S��c����S�a0  Y�D0�������  �e��WV�U  �X�D WV�Y  hL�D V�N  SV�G  WV�@  ������V�4  h  h$�D V��3  ��<j�����u�����h�  j h�  j ��������tQV�5��F j2�5��F j������Y�E�    �=��F ���F �ʉ5�F _�u�<  �5�F ���  ��T�   ���F �,�F ��[҉h�F Q�,�F �����B����  ��  ��P  Z���  N���F ���   �扅d  ���F ���F ��F     �|�F ���F ���F �5��F �5�F ��\  �5��F ��4���F �Q�58�F �5��F h�  j�N   Ë+�[�Ջ���=,�F �c���B���>  NR��l  ���   Q���扅D  _�������\  ��@�th�  hp  j j
Q�  Í,�F ��[��Ѝ,�F P��`  ��D  ��d  ���  ��\  ��  ��F ���������`  �3  ��|  ��`  ��\  [��   ��8  ���  ��L������5,�F �+�[�Ջ�W��@  �B��������_�h�F �,�F ��������:  �,�F NR���F ���   Q���拈<  �=��F �5��F j ��@  �}��u����  ��X  ��X�5��F �=��F �R�����\  �I��,  ���F h�  j�5��F ����É�X  ���F ��D  �������5,�F �/��Ջ�S�] �B��,  �� S��   �]����  X�E ���  �ŀ  ����  ���D � �HF ���tP�p�F �HF ����SV���D �5HF ���h�F ����uIh�   j��������YYt-V�5HF �l�F ��t�FT}F �F   ���D �N���j���YS���D ��^[�jhPE �		  �u3�;��  �F$;�tP�k���Y�F,;�tP�]���Y�F4;�tP�O���Y�F<;�tP�A���Y�FD;�tP�3���Y�FH;�tP�%���Y�FT=}F tP����Yj���Y�}��F`�E�;�t�u;4�F tP����Y�M���   j�l��Y�E�   �Fd�E�;�tM�9x,t�H,�	9x4t�H4�	9x0t�H0�	9x@t�H@�	�HL���   ;�{F t=x{F t98uP�=9  Y�M���    V�m���Y�&  � 3��uj�4��YËuj�(��Y������u����3��VWh,�D ���D ����tk�5 �D h�E W��h|E W�d�F ��hpE W�h�F ��hhE W�l�F �փ=h�F  �p�F u(���D �h�F ���D �l�F ���D �d�F ��@ �p�F h��@ �d�F ����HF tA3�h�   GW�П������YYt+V�5HF �l�F ��t�FT}F �~���D �N������A���3�_^���   ���  j ��,  ��$  �L�F ������^��X�F ��� �L�F V�ڍ,�F ���  ���������  �L�F ��  ǅ      �X�F ��,  ��  ���  �(�F �=@�F ��H  �X�F ��  ���������h����D$�    �|�F ���F �L$��L�F �l$��|�F �l$��-d�F �l$��  U����e� �} S�]VW����  �E�ȃ����4��<�̈́F ���ƊH����  ��Ht"�x
t��D0�M���S�E�   �D0
j �E�P�u�R�40��D ��u9���D j^;�u�uK��� 	   �sK���0���m�&  P�iK��Y����  �E�E��D1���   ��t�;
u���D0��	��D0� ��E�M��;��E�M���   �E� <��   <t�C�E�   I9Ms�E@�8
u�E�Y�E�n�Ej �E�Pj�E�P��40��D ��u
���D ��uF�}� t@��D0Ht�E�<
t���D1�(;]u�}�
u�
�jj��u�l~�����}�
t�C�M�9M�L������D0@u�t0�+]�]��E��3�_^[��jh��D �  �];��F sx�����<�̈́F �Ã��4�����D0tXS�n��Y�e� ��D0t�u�uS��������E����I��� 	   ��I���  �M���M���   �E��!�]S��n��Y��I��� 	   �I���  ����  ËD$f�@@f��u�+D$��HË=��F �|$ȋ|$��5@�F ���F ��  �d$�����\$��\$��L$��8�F ;�,� �5@�F ���F �|�F �L$�D$̉��F ���F �T$��T$��d�F �8�F �l$��\$ȋ��F ���F �t$̋-<�F ���F �5��F �V������  ��$  �$  ���  ��F ���F ���F �0�F �,�F �h�F ǅ�      h�  ��   Ë�F ���  ���  �5h�F ����=  ��(���F ���  ӄ$  �=�F �=��F +=��F �$  F�5��F �5|�F jjF�7  Ã�<��$�  ������  ;��F ��S����$�  �=�F �0�F �ʉ��F ���  �0�F ���F ���F ��   ���F ���  ���  ���  �d�F j(������d�F     �5@�F ���F �8�F �|$����F �-<�F �\$̋T$ȋ|$Ћl$ԉT$����  ���F ���F �L$ȋd�F ;D$��, �d�F d�F �  ��(��$  ������F ���  ;��F �^V������$�  ���  9�$�  ��v���@�F ���  ��$�  �$�  ��F =��F �:=��F ���F P���F ���  ǅ�      �=��F ��F �@�F ���F �=��F �5��F ���  ���  �   9�$�  �q���5,�F h�  h�  �5$�F �X�������h0@ d�    P�D$�l$�l$+�SVW�E��e�P�E��E������E��E�d�    ËM�d�    Y_^[�QÉ��  j �5|�F �5��F �   �[���  ���F �=��F ��,�Ή�$�  �5,�F �-�F ��ǅ�      j�0���Ël$�ŋM �4�F �D$�    �|$ЉL$̋4�F �	��������L$��T$��T$ԋ��  �D$���F �D$�+��F D$��4�F �T$��T�F �L$̋�F 롉��  ����������<���F ���  ӄ$�  ���F +��F �$�  F�����  ��,�������F ���F �5�F �5��F �;��F �A����5�F ���F ���F ���F O����������F ���  ��F 뤉�$�  ���F �-��F �$�  9�$�  �m�����$�  ����F �=��F ���  ���  ���F �Q������  ���%  Ӄl&  �=��F ��$+  {X��F ���F Wd�5    d�%    ��\(  ���)  ��E�    ���  �h�F �u�u�;u��b  �u�uЉ5��F �u�5��F ���T�F ��F     ���  �u�u�t�F �T�F �	����   �H�F ���  ��F �H�F +��F �F �T�F �M܋u�t�F �d�    �d�    �� �F ӏ *  ��$+  ��H)  #��(  �=L�F 3=��F �=D�F �=,�F ��*  =��F ���  �,�F ��<&  �=|�F =4�F ��b@B��$+  b�7Sjj ����Á%�F ������F ��F �=t�F ;�D=  ���F �EЉ,�F �]܋ϋh�F ���  �������  ������F ���  ;�$�  �������F ���F ���  ���  �5��F ���  �  ���U��WVS�u�}����
�t2����'��8�t�,A<ɀ� �A��,A<ɀ� �A8�t�����[^_����=   s��ă�� �� P�Q�L$��   -   �=   s�+ȋą���@PÉ5\�F ���  �5p�F ���F � �F �T�F � ��������$�F ���  ӄ$�  +��F �$�  �T�F �$�F ���  ���  �5\�F � �F ����F     �5��F ���  �5p�F ���F 9=��F ��������  ���F ���F ��F ���  Ë35��F �5T�F ǅ�      �������F �M܋U�M��A��F ���F �=8�F ���F ���  �=`�F �ǋ8�F +��F C�Ë��F �ˉ5��F ���u�]܋��F ��@  �7�`�F ��  P�d�F �L�F �5�F P�|�F ��P  �M��ы��F ���F �5��F �=��F �؋m�-��F ���F ��$�  �=��F �d�F ��$�  ���F �=��F ���  ��  ��  �=8�F �}�=��F =��F �����  �x�F �}̋]ԉ4�F �0�F �=8�F �`�F �M�x�F �S  ��F ���F �5��F ��d  �5��F �H�F �5�F ��[��5��F �Ћ5l�F �T�F ���F ��d  �J  �T�F B��   ��
  ��P���7  �}  ���F �p�F V���F �5l�F ��F ��  �p�F ���(�F [��d  ��   �b  �(�F ���7  �q  ����  �z  ��   ��  @��d  ��  �  �h�F �E�    �u�M��,�F �U��`�F ���F �M�`�F �   ��f`  �����  +��F ;t�F �t� �@�F �]�`�F ��    �5|�F �u�1�$  9���%  ���F �M�`�F �U�`�F ���  �R�|�F �E�}�   ��� �}܉5�F �ʉ��F �}�5|�F �@�F �=��F �=�F �U��}�}�� ������F ���EЋ �F �U�P�F ���F ���F �MԋE��S  ]� ��������W�|$�n��$    ���L$W��   t�����t=��   u�������~Ѓ��3�� �t�A���t#��t�  � t�   �t�͍y���y���y���y��L$��   t�����tf�����   u���������~�Ѓ��3��� �t��t4��t'��  � t��   �t�ǉ�D$_�f��D$�G _�f��D$_È�D$_��]����L$�H��P����Hi��C ��Þ& �H����%�  É=��F Y���F     ��|  �M�=h�F ǁ      ��$  �O<��Y|�yx�$  ����� �u��5,�F �O�w�5��F �w�t�F �O �$  ���F �W$�$  �5��F �o�$  �l$�싰�  �������P�F �E�u���F � �F ���F �MԋE��V���S���F �=8�F �H�F �=T�F ���F �=x�F [�֋=8�F �Đ   �  �M܋��F ����VW�����xd;=�{F t�\'  ���t$�(�~jPW�,  ���
�OH�A����tF���F��-��t��+u�F3���0|
��9��0�������t���A�F�݃�-_^u����s���d�    �d�    �식,
  ���� ��$�
  �5��F ��$�	  �5D�F �5 �F �5`�F �5�F ��F ��j ���	  ���  �э,�F ��   �� Bǆ|"      ^��}  ���  �,�F ���F �J�ѳ��V���F ���  �́�   ��� F���  ������ǅ�      �։��  ���  ���F ���  ��@닃�P�m  �N  ��  ������   ��  @��P�F  �0  ��   `@���F ��P�)  ���F �5��F V���  ���F ���  ������\  ��D  ���F ��d  ���F ���F Z�� �  �H�F P���F ���F ^�5x�F �l�F �Đ   ��  ��F �,�F �@���H+ V��d  �H�F �5��F � �F ���F ��F S�֋ �F �x�F [�Č   �p  ��P�J  ���F �,�F ��\  ǅD     ���  ��d  �5��F �58�F ��  ËH�F ���F ���F ���F ���F �։x�F ��D  �Đ   ��  ���F ��D  �5��F ��d  ���F �5l�F �H�F ��F ��  ��D  ��\  ����@  �=��F ��d  ��   �D	  ��@  ���7  ��  ��x��  �����5,�F �3�[��։��F �,�F �2� B���F j���F     S��\  ��4������F �8�F ��d  [��\  ��4��  jd�5�F h�  �
  ËH�F �<�F ���F ���F �<�F �։x�F �(�F �Đ   ��  ��p  R��<  ǅ$     �5��F ���  ���  ��t  �ʋ} Z���  ��T�%  ��F �,�F ��|$  ���"  � ��F ����"  �����  ���F ���  �,�F ���#  �5��F ����F J��������  ���  ��������F �5��F ]Ǆ$@     ���F �t$���$X  ���F ����  ��8�w  ���F ���F �x�F �H�F ���F ���F �ցĐ   �  W���F ��\  �=H�F �T�F �=��F �x�F ��\  ��_�Đ   �h  ��D  ���F ���F B���F ��   �Ћ�[�S���F �p�F �5D�F �H�F ��d  [�Ћ5l�F �D�F ��d  �F  �p�F B��   ��  �����7  ��  ��  ��  ��   �����@�W����h�F ��@  ��8  ��F    �L�F ���F ���F ���F R��   �ʋL�F �=��F �=�F ��   ��@  �=��F ���  ��T���  �,�F �5��F �5��F �5��F �  Ë��F S���F �D�F [��P��D�F ���F ��F @��F W�=D�F ��d  @�0�F �x�F _�H�F ���F �0�F �ց��   ��   ����  �5��F ��F ��d  �5��F �x�F @���F �t�F �Č   �   ��[ɉ�F Y��F �`�F �,�F �L� B�`�F ǅd     �X�F     ��d  �8�F �`�F ��\  �=X�F ��d  ��\  ��P��  �m  J�  ��� �x�F ��)щ5�F ��x�F �0�F �މ=,�F �=�F �P��d  �(�F ���F �50�F �ω5��F ��R�=,�F ��4�����|  ��P�
  ��D  h�  h�  h�  �y  �R�,�F ��,�F ҋ�   �=,�F �W���B���  ���  R�,�F Z�m  ���F ��\  ��d  �=D�F ��\  ��4�������F �D�F �D�F �p�F ��P�������D  �t�F ���F B���F �� �{������F �֋�[ɉ�d  ���F ��F ���F ��d  ���F ���F ���/�����F ��F ���F ���F ���F F���r  �5,�F S���F ��d  ��p  ���F ��\  ��  �t�F ���  ���F Z��R����F ���t�F ��F ��d  ���F �<�����t��5,�F ��T  ���F ��\  ���  ���F V���F ��d  ��F �5��F ���F �5H�F ������5��F ��P������Y��d  �x�F ��F �Đ   �������F ��\  ��D  V�5��F �5��F Z�����(�F ��d  ��4�.�����|  �5,�F �3�[��=�F �=,�F �֋=�F �,�F �,�F �n   B�������,�F �
  ��F �x�F ���F ��l��������F ���F �D�F ��D  ��(�����R����  �H�F �5P�F �5H�F �x�F V�5�F ���F �5��F ��d  �P�F ��p�{����,�F ǅ�����  ǅ�����E ��   ����D  V���  ��  ���F �,�����5��F h�  ��   Ã�4� ����5,�F �+�[�Ջ�Q��d  �B��  �����Q�M���T  _��d  ��T  ��   ����  ��� ���F    j �5��F �H�F �58�F Y��d  �H�F ��|�s  ���F ���F ��F ���F �H�F ��������F ��P�Ƌ��F ^���F �5x�F ��l�O����ϋ�@  ��(�!�����5��F �5��F j j Q��  ËH�F ���F P���F �(�F ^�5x�F �l�F �Đ   �����P�,�F ��d  ��\  ���F �=@�F ��  ���F ��L  ��  ��Z��`  ��\  ��D�%	  �,�F ��[��Ѝ5,�F �5��F ���F ��\  P�5H�F ���F ��F ��D  ���F ���F �������^��q���������d  ��8�F �5��F �%  ËH�F ���F �-p�F ���F �-x�F �\$��֋��X  �Đ   �������  �5,�F �3�[��։��F �,�F ��� F�H�F ��F �����F    j ���F Y�8�F ��d  ��F �ց�   �d  jh�E ����3ۉ]������pd�u�;5�{F t
��  ���u�F;�u(�E��8��   �
��A|
��Z�� �
B8u��   j�vSSj��uh   P�ך���� �E�;���   �]�����������e���}؃M���3�@Ëe��E  3�3��M���u�;�u�u��@���Y���E�   ;�t-j�v�u�Wj��uh   �v�a����� ��tW�u�B���YY9]�tW葉��Y�E�e��D�����5��F �'�������F h   �������Y�L$�At�I�A   ��I�A�A�A   �A�a ���� ����5,�F S�5��F j jQ������������d  ��(���o������������ j��F     ^��x����58�F ��F ��d  ��x�����   눍5,�F �3�[���Q�,�F �����B������Y���F �,�F �� ���F j���F     ^��H����58�F ���F ��d  ��H�����P�����h  %�   ��\  X�5��F �  ����������F �,�F ��d  R�@�F ���F ��\  �5x�F �5@�F �ʋ�\  Z��D�U  �8�F    ǅd      �5�F jPW�54�F ����Ë��   �S���  �,�F ���F �,�F ��� ��x������F Zǅt���   ���F     ��t������F �8�F ��d  ���F �,�F ��|�5�F �5��F V�	����� �����5��F �5�F S�S   ��h� j�5�F �$���Í,�F N������� ��������)���j ����Í5,�F jh�  S�2  ��B���j Vh�  Qj����á�F U3�;�V�5��D u-�օ�t��F    � ���D ��xu��F    �3��\��u���S��u�SW���D �=��D UUj���SjU�׋�;�t&�6P�������YtVUj�Sjj �ׅ�uU����Y3����_[^]���������|  �5��F ����É��F ���F �`�F �5��F �H�F ��\  �5��F ��|  �ĸ   뮃�$���F �5��F �H�F �5��F ��|  ���   ���  �Sh�  jdh�  �5��F ����Ë�@  ��[��Ћ=��F ��\  ��@  �   �H�F ��0  ��|  B��H�"�����F ���F S��\  ���F ��d  �t_[�=��F ���F ��0�����D  ���F ��@  ��0�����\  �h  ���F �5T�F ���F ��h  ��|  ���   ����[��[��Ћ=��F �5��F ��0  �5��F ���F ��D  ��@  ��0  ��\  �5��F �=��F �I  �H�F ��|  B��H�9������F    ��d  ��X  ���F    �@�F     ǅh      ���F ���F ��|  ���F �5��F Rh�  �����É�d  ���������F �@�F �H�F �=T�F Z��|  ��d  �=��F ��h  �=T�F ���   ������F ��D  ��@  ��\  �=��F ��d  ��������F ��d  ��  �h�F V��@  �H�F ��|  ��L�.������F ��d  ���F     �5@�F ���F ���F ��h  ���F ��|  ��H�������D  �5�F h�  �5��F �  É��F V���F     ���F �5@�F ���F ��h  ��F ��|  ���   �����,�F �$�  ���   Q��d  �	�� ���	�d  �C�H�F R�5L�F �,�F �@�F ��|  �D�F ��\  ��x����=@�F Q��t�����\  �H�F �������H�F �=h�F ��D  ^��d  �=p�F �=��F ���F �=h�F ��  S���F ���F �T�F �H�F ��D  ��d  @[���F �5��F ��4�  �l�F �,�F 	5l�F ���  ǅD     ��@  ��  j h�  h�   �5��F �Y  ËL$��   t$�����tN��   u�    ��$    ��$    �����~Ѓ��3�� �t�A���t2��t$�  � t�   �t�͍A��L$+�ÍA��L$+�ÍA��L$+�ÍA��L$+������̋D$�L$ȋL$u	�D$��� S��؋D$�d$؋D$���[� �5��F Q�5��F j jP�����j$h �D �	���3�3�G95��F u2�E�PWhl�D W���D ��t�=��F ����D ��xu
���F    ���F ;�u�u�u�u�u���D �  ��t;�uS�uЉu�9uu�p�F �E9uu���F �E�u�~b��Y9Et���t�EVVVV�u�uV�u�D�D �؉]�;�u3��N  �u��Ã���������e�ĉE�SVP�  ���M���3�@Ëe���	  �e� �M��3�G�]�3�9u�uSW�s��YY�E�;�t��}�VVS�u��u�uV�u�D�D ����   �}��D������:����e�ĉE��M���3�@Ëe��s	  �e� �M��3�G�]�3�9u�u�DP�f���Y�E�;�to�}�9uu�p�F �E�}��E��4f���f�N���PS�u��u�u���D �E�f�~���tf�>��uW�u��u�$  ����e� �}� t	�u��~��Y3�9u�t	�u��y~��Y�E̍e��,����U��� V�uW�EP�u�E�P�E�����E�B   �u�u�薨��������t�M�x�E��  ��E�Pj �����YY��_^�Ë��F ��  �,�F �5��F j �K���Ë�D  ��\  �5��F ��D  �5��F ��\뻋H�F ��F �p�F ��d  ���F ��D  ��F ��������F ���F �x���U���S3�9�F VWumh��D ���D ��;���   �5 �D h��D W�օ���F t|h��D W��h��D W��F �փ=ȭF � �F uh��D W�օ��(�F th|�D W�֣$�F �$�F ��t<�Ѕ�t�M�Qj�M�QjP�(�F ��t�E�u�=ԭF r
�M �)3��5�M���F ��t�Ћ؅�t� �F ��tS�Ћ��u�u�uS��F _^[�Ë��F ��$�  ����$`  ���H  ��,�Y���Z���F �5<�F ��D  ��d  	5<�F �H�F ��F ���F    �<�F ��d  �<�F ��0  ��@  �Ћ�F ��������  �-<�F �5��F ��$�  �-l�F �= �F �O������J���j�5�F h�  h�  j�   É�\  jh�  h�  ����ËD$;��F r3�Ëȃ�����̈́F ���D���@�U��WV�u�M�}�����;�v;��|  ��   u������r)��$��1A �Ǻ   ��r����$� 1A �$��1A ��$��1A �1A <1A `1A #ъ��F�G�F���G������r���$��1A �I #ъ��F���G������r���$��1A �#ъ���������r���$��1A �I �1A �1A �1A �1A �1A �1A �1A �1A �D��D��D��D��D��D��D���D���D��D��D���D���D���D����    ���$��1A ���1A 2A 2A $2A �E^_�Ð���E^_�Ð���F�G�E^_�ÍI ���F�G�F�G�E^_�Ð�t1��|9���   u$������r����$��3A �����$�83A �I �Ǻ   ��r��+��$��2A �$��3A ��2A �2A �2A �F#шG��������r�����$��3A �I �F#шG�F���G������r�����$��3A ��F#шG�F�G�F���G�������V�������$��3A �I <3A D3A L3A T3A \3A d3A l3A 3A �D��D��D��D��D��D��D��D��D��D��D��D��D��D���    ���$��3A ���3A �3A �3A �3A �E^_�Ð�F�G�E^_�ÍI �F�G�F�G�E^_�Ð�F�G�F�G�F�G�E^_�É�d  ����F �p�F ���F ������S�p�F �5D�F �H�F ��d  [������,�F ��\  ���  ��@  ��  ��d  ���  ��D  �5l�F �H�F ���  ��[���\  ��  �=��F ���F ���F �5l�F �D�F ��D  �A���V�t$WV�d=�����Yt<��t��uj�M=��j���D=��;�YYtV�8=��YP���D ��u
���D ���3�V�<��������̈́F ����Y���D� tW���Y����3�_^�jh`�D �u����];��F sh�����<�̈́F �Ã��4�����D0tHS��<��Y�e� ��D0tS�,���Y�E���>��� 	   �M���M���   �E��!�]S�Q=��Y����� 	   ����  ����"���É=�F �E؋=��F �]ԋ�F ���F �]��+���F ��@�F 9���������F ���F ���F �E܉M�E؉��F �M܋��F �U���F �`�F �=��F �=��F �;��F �������F ���F ���F G�M؋M؅���������F �G���U���LSVWjX������j�E�PV�h�D ��tw�]܍E�P�\�D �M��ȭF �y���#�+���N����������;��M�r@��t\�]��   j�E�P�u��h�D ��t �E�E��]�t��E��E؉E�t3�@�D;�s3��<;�s�u�jS�u��u����D �ȭF ��}�H���%  �M�Q@P�u��u����D �e�_^[��jh@�D �>����=�`F u:j�;���Y�e� �uV�U,��Y�E���t�v���	�u���u�M���$   �}� u�uj �5��F ��D ��������Ëu�j�.���YÃ�,��x  �5��F Q�5��F �   É��F ��F �;��F ��\����h  ��x  BI���,� ��h  ���F ���F ���F ��F ���F ��<늉�p  � �F �5d�F �$�  9�$d  ��[������p  ��l  ��x  ���F ��F ���F �8������F �5��F ���F �]����F ��v�]��k  ��@  ����T  Pd�5    d�%    �V�t$�F<W3�;\�F tc;�t_�F,98uX�F4;�t98u;��F tP�	s���v<�;  YY�F0;�t98u;�uF tP��r���v<�^q��YY�v,��r���v<��r��YY�F@;�F t;�t98uP�r���FD-�   P�r��YY�FP;`�F t;�t9��   uP�-  �vP�|r��YYV�tr��Y_^�V�h������Nd;�{F ��   3�;�t/�A,�	;�t��A4;�t��A0;�t��A@;�t��AL���   ��{F �Fd��{F � ��{F 9P,t
�@,� ��{F 9P4t
�@4� ��{F 9P0t
�@0� ��{F 9P@t
�@@� ��{F �@L���   ;�t9u��x{F tQ�u���Y�Fd^�jh��D �'���j�-���Y�e� �"����E�M���	   �E��=����j�R���YÉ-��F ��U���   ���  �� @ ���F     ���F     �=��F �=��F G���  �mx��R�,�F Z���F ���F �5��F �5��F �F���   ���   �l���� �F �5��F ���F R���F  �F ���F ���  ���F ���F W�5��F �=��F �U����_���B�j  _@���a  ���F ��@  �H�F ���F ���F �x�F ��F �2  �Ћ% ���	��A���F �����4�F Q�H�F ��\  �x�F Y�4�F ���F Q�4�F ��   �H�F ���F B�X�F ��\  �x�F �X�F �   Z��\  �% ���	��A���F �/������F �=��F ��D  �H�F ��\  ���F �=x�F R��D  �=��F �{�   ��\  �=��F �=��F ��d  ��[��Ћ=��F �@��$$  �����P��D  ���F �H�F Y�x�F ��F �J�,�F ���F ��F �H�F h   �H�F ��F �x�F Z��d  ǅ\     ǅD      �H�F ��F ���F ��D  �x�F ��7����H�F ��F R���F ��d  ���$(  ������5,�F ^�5x�F �,�F ��D  ��F 둍,�F �5,�F ��vۉ5,�F �Ӎ5,�F P��\  �B�@�F ��������  X�5��F ��\  �   �H�F �x�F ���F B��F ������5,�F �,�F ��d  ���  ���  �(�F     ��  �@�F ���  ��\  ���  �ϋ��  ��\  ���  ���B��d  ǅ\      ��  Q������,�F ��\  ��@�F �������\  �֍,�F ǂ\%     jF�]  ����F �5��F ǅ�     ���  ���F ���F ��0�,  ���"  �D�F ���F F���  �L�F Y���F ���  �L�F ���F ���  ����   �=ȭF u�=ԭF r3�@�jX�3�9D$j ��h   P�T�D �����F t*���������`F uh�  ��#����Yu�5��F �t�D 3��3�@�U��Q�E�H��   �Mw	�IH�A�TV����W�yH���Dw�_^tj�E��U��E� X�
�E�3��E� @j�q�q�MQP�E�Pj��l������u���E#E����5|�F �   �BY��ǅ<���   ���F ��<������F ���F ���ǉH�F ���F ���  �H�F ���F ���  ��0뜍,�F ��  ���F ���F    ���F ���F ���F ��0�f�����F ��8�F �]����F B�8�F ����   ��(�8�����  j jRP�58�F �R   É�F �,�F ^��v�V��S�,�F ���"  �@I��z�����F ��[���F ���  ���F ��F �c���F ���5�F �   ��1  ��F ��(������F �֋��F j �   ���������x����5,�F j
�5��F j<�B   Ë��  ��   ���  ǅ�      ���  ���  ���"  ���  ���   ���   H���  ��4"  ���   ���$  �������  ���  ǅ�      ���F ��(������  ���!  ���  ���"  ���!  ��4�(��������D���H�`�F ���   �����F     ��y����5��F �I��w���5��F �ት�  �5,�F �)�I��F R�ՉL$ X�������B������H���  ��4"  ���   ����������,�F ��Iҋ��F �,�F ��\%  �B���  Q�,�F �2���� ��������̋T$�L$��tO3��D$W����r1�ك�t+ш����u������������ʃ���t��t
�����u��D$_ËD$�jh0E ����3��}�j����Y�}����F �]؉=@�F ���F ����F �h,E �IQ��Y���u�;���   �> ��   �D�F ;�t!PV�F���YY����  �D�F ;�tP�	h��YV����@P�d���YY�D�F ;��d  VP����YY�M���i  jV�5��F ���������F �@ ���>-u�E�   FV����Yi�  ��F �0�<+t:��&  <9�  F��D�F ;�tP�tg��Y�=D�F h��F ���D �����   3�A�@�F ���F k�<��F f9=ڱF t��F k�<£�F f9=.�F t�<�F ;�t��F +�F k�<��F ��=�F �=�F �E�PWj?�5��F j�h��F WS�5D�D �օ�t9}�u���F �@? ����F �  �E�PWj?�5��F j�h�F WS�օ�t9}�u���F �@? ����F �  j��E�P�[��YY�   �u�3�j�F���YÀ>:u>FV�:���Yk�<�F �<9F�:�}��>:uFV����Y�F �<9F�:�}�9}�t��F ���F ;�tjV�5��F ���������F �@ ����F �  �����jh@E �\���3�95H�F u'j�X���Y�u�95H�F u�*����H�F �M���   �a����j�v���YË� ����=��F ��$���������5,�F �1�I���Q�D�F �,�F �6���B�-D�F �Q}���D�F W�=`�F ���   ��Ӡ$  _ǅ ���    �D�F 닉}̋�C��F �Uȋ�)�B���ʉu����}��=�F ���F �}��l�F ���F �=0�F ���  �}���M���  ��F Q�L�F SP�d�F � �D �Uȋ}̋|�F �ȋmĉ�$�  �-��F ��$�  �0�F ���  ��  �F  �=��F ���  �_<��{|�D�F �Cx�\�F �E��D�F ���  M��M���������,�F �U�U��B�J�R�u�u��^ �= �F �5D�F �=�E��M���������F ���F ����  ���F ��$�  �=��F ��$�  �2  ���  ��]�]��[$��U��U��R���F �,�F �M�X�P�F     ��|  ���F �M��e  ���F �5��F u�uЋ����  �U�5H�F ���F �u��e��]܋�F �MЋM���  ;M��5� �=��F �}ԉ�  ����F �P�F �=P�F E   �e����}̉Mȉ]ĉu��m܋|$���F ���F ���-�F �|$�T$�D$̋T$ċ��  �h�F �\$�L$܉\$��l$��l$�������F     ��$�  ��$�  ��$�  ���F ���F ���F ��F ;�$�  �������F �F �=��F ��$�  ϋ��F ��$�  Ǆ$�      �W��F ���F ��$�  ������F ��$�  ;��F �̨������F ���F �-4�F ��$�  ��$�  �������$�  ���F ���F ���F �-4�F ��$�  �M ���w�����$�  ���F ��$�  ӄ$�  ���F ��$�  +��F �$�  E��$�  �x�F ���F ��$�  �-4�F ���F ���F ��$�  ��$�  �j���F �0�F �������F �Eԉ��  ���F �U�Ƌ]܉h�F �   ��ξ���u�����  +U�;�F �5����]�����F �\������F �������@���  �؋�����@���F �  V��  ���F �Ë��F �l�F ���  ���F �% ���	��AJ�� P�5�F �x�F �Ë5��F �5l�F �5�F ���J  U��QSVW�����}���VT��}F ��99t�@����;�r�@��;�s99t3Ʌ��  �Y�ۉ]�  ��u�a 3�@��   ����   �FX�E��E�FX�A����   ��}F ��}F �;�}'�R���~T�d8 �=�}F ��}F B߃�;�|�]�	���  ��~\u	�F\�   �d���  �u	�F\�   �S���  �u	�F\�   �B���  �u	�F\�   �1���  �u	�F\�   � ���  �u	�F\�   ����  �u�F\�   �v\j��Y�~\��a P�ӋE�Y�FX����	�u���D _^[��V�t$����   �F�X{F ;At;4{F tP�^��Y�F�X{F ;At;8{F tP�^��Y�F�X{F ;At;<{F tP�c^��Y�F�X{F ;At;@{F tP�F^��Y�F�X{F ;At;D{F tP�)^��Y�F �X{F ;A t;H{F tP�^��Y�v$�X{F ;p$t;5L{F tV��]��Y^�@���x�F    �؋x�F �p�F ���F    j ��^�p�F ������؉p�F ����F �3���V�֋É��F ���F �l�F @���F 듋؋% ���	��AJ�`� ��H  ��  �Ë��F �l�F ��  ��  �x�F ��  �S����@�F �Ë@�F �l�F ���+����Ë��F �l�F @���F ��������H  ��H  �l�F �������jh�E �T���3ۉ]��Į���pd�u�;5�{F t
�������u�F;�u(�E��8��   �
��a|
��z�� �
B8u��   j�vSSj��uh   P�m���� �E�;���   �]�������P����e���}؃M���3�@Ëe�����3�3��M���u�;�u�u�����Y���E�   ;�t-j�v�u�Wj��uh   �v�l���� ��tW�u����YY9]�tW��[��Y�E�e�舷��ËL$��tI�8 t@��u�I�D$+�H�j@h �D �$���� {F �E�3�3�F9=�F u2V�l�D PVPWW���D ��t�5�F ����D ��xu
��F    9}~�u�E����Y�E�E;�~P�E�m���Y�E��F j[;��9  ;��1  ;��V  �}ĉ}��}�9} u	���F �M 9}t;���   9Eu���  ;���  9u~jX�  �E�P�u �X�D ����  9}~+9]�rٍEր}� tЊP��tɋM�	:r:�v�À8 u��9}~>9]��=  �Eր}� �0  �P���%  �M�	:r:��h���À8 u��  WW�u�uj	�u ���D �؉]�;��i  �}������������e�ĉẼM���3�@Ëe��O����e� �M���]�3�F3��E�;�u�P�A���Y�E�;��  �u�SP�u�uV�u ���D ����   j j �u�uj	�u ���D ���u�����   �E�   �6������|����e���}��M���3�@Ëe�����3��M���]��u���u�6P����Y����t@�E�   VW�u�uj�u ���D ��tVWS�u��u�u���D �E��}� tW��X��Y�}� t	�u���X��Y�E��   �}�9}u�p�F �E�] ;�u���F �u�K;��Y�����u3��};�tIj j �EP�uVS�l;��������t�j j �EP�uVS�Q;�����Eȅ�u	W�uX��Y븉}�EȉE�u�u�u�u�u�u���D ����tW�EX���u��=X��YY�ƍe��M��mT������É5 �F �5�F � �F ���F �	;��F �~!�����F � �F � �F ���������5 �F � �F 믉��F ���F ��$�  ��$�  �$�  9��F �>���-��F �쉍�  �5�F ���F �5��F ���F ���  �Q���#��  BX��cC����  �=��F =��F ����
  ��$  ���F ���  �5��F 3�l
  �8�F ӊ�  ���  ��F �-��F ś�����  ���F JX�%x�F ���  �|�F Ӣ$
  �-x�F �"I���F ��F �,�F ��L	  ��F ���  �,�F ��|  ��D	  #��F �$�F �,�F ���  ���  3��	  ���  ���  ���  h�  �5��F �5��F WQ�c  �V�t$����  �v�BV���v�:V���v�2V���v�*V���v�"V���v�V���6�V���v �V���v$�V���v(��U���v,��U���v0��U���v4��U���v��U���v8��U���v<��U����@�v@��U���vD�U���vH�U���vL�U���vP�U���vT�U���vX�U���v\�U���v`�U���vd�xU���vh�pU���vl�hU���vp�`U���vt�XU���vx�PU���v|�HU����@���   �:U�����   �/U�����   �$U�����   �U�����   �U�����   �U�����   ��T�����   ��T�����   ��T�����   ��T�����   ��T����,^�V�5��F �����Y�L�F ����F ��+Ѓ�;�sN�   ;�s���QP�������YYu��V�5��F ������YYu^ËL�F +��F ���F �����L�F �9�L�F ��^�h�   覿����Y���F ujXÃ  ���F �L�F 3��jhP�D 藯���Կ���e� �}�;����E�M���	   �E�譯���跿����t$���������YHÉ�D  ���F ���F �<�F ��5��F �5��F �2ʉ�F �<�F �1�I��$�  ��   ��8  ���F �$�F ���F ;��  ���  � �ɄF ��Vj^u�   �;�}�ƣɄF jP�qG����YY��F ujV�5ɄF �XG����YY��F ujX^�3ҹXF ���F ��� ����؁F |�3ɺhF ��������4�̈́F �������t��u�
��� A���F |�3�^��*���= �F  t����ËD$�XF ;�r=��F w+�����P����YÃ� P���D ËD$��}��P����YËD$�� P���D ËD$�XF ;�r=��F w+�����P����YÃ� P���D ËD$��}��P����YËD$�� P���D Él�F j
�����=,�F �[��$�  �������D  Q���	  ���	  �l�F ��D  ���F ���	  ���  ����   �<�F ����F ���F ��D  �l�F ���|���d�    �(d�-    �쉝�  �,�F ���  ���
  ���F ��  �-@�F �@�F +��  ȋ��
  ˉ �F �,�F ���F (8��D
  ���F �5��F �5 �F �}����h@  �5��F jQ�54�F �   �ǅd     ǅD      �5P�F �58�F j	�   É5��F ��D  �ǅ8      �<�F     �5|�F j
h�  �58�F �5�F �s���ËE�A���   ���F ���F �u����)  ���&  ���'  �u�5l�F ��d(  �%H�F �=��F ��5��F É��  ���F 4�F 9��m���p�F ���F �=(�F ���  �D�F �-��F ��$�  �=d�F �d�F �4�F ��$�  �l�F ��$�  ���F ��$�  ��$�  ��$�  ���F �5p�F ���F ��$�  ��$�  ��  ��F     �]ԉ��F �=H�F �=�F ;=��F ��6���=�F =�F ���F ��H�F �E��E�    �}ċ=H�F �M��M��	���  �`�F �\�F �Uԋ��  �Eȉu��5`�F +5��F u��E؋M��5 �F �}ċ\�F �u�뢋L$���   �-��F �싐�)  +�+  +��*  �u��U��   ��t  ���   ���*  �Q���   �Q���   �Q���   �q��������  �� @ ���F �5��F �3   �9�$  �s�����  �,�F ��  ���  V�5��F �  Í,�F ǅ�      ǁ8"      j �Q  Áe�����}ȉP�F �]�;;��  �=H�F ��F �M����F �ˋ��F �]��B�����$�  �l�F �4�F ��$�  �=l�F ��$�  ��$�  ��$�  ��$�  ���F ���F ���.���F ����F 9��}�����  �p�F ���F ���F ���  � �F ���  �
;��F �
��B��$�  ���  ���  �������p�F ���  �,�F � �F ���  ���  �,�F ���  ���  �ǅ�      h�  �5��F h�  W�]���Ëd�F jdSV�F  É��  �,�F �-�F �QH��%�F Q�5��F �������$   �$   ���  ���$  ���F ���  �,�F ���  ǂ      h�  V�5��F �5��F ��  É��  ���  ���  ���  <���  ���F �=t�F � �F ���  �d�F �t�F ���  �d�F � �F ���F ���  �p�F ���F ��<������$p  �=��F j
�5��F h�  �5��F �58�F �^���Ë1���  �d�F �I���  ���A��Q	  ������=t�F �=,�F ���  �5p�F ���F �d�F �0�d�F %�   =�   t��5��F �5��F �5��F �5|�F �T���Á%<�F ���P�<�F ;��F �������$  ���  ;0�F ������$  �$  �|�F ���F щ��F ���F �=��F ���  ���  ���F ���F     ���  ���F �|�F ���  �<�F ���F �A��F ���  ���  �	����   ��@Q���  �<�F Z+��F <�F ��$�  ���  �=��F ���  ��������Q���  �<�F ���F X+��F <�F G���  ���  �=��F ���F �5,�F ���  ���  ���  �   ��@�%<�F ����<�F ;��F �L����$  �=��F P���  ���������  �5$�F WVj �����ËE����F �}��}��;��F �J?���}��E�J����>����F �ˋ5,�F ������P�F jǅH      ��P��|������  X��H  ��$  ��|����   �$�F �]����F �U�$�F 9$�F �2<���5$�F ��F �u����F �U��F����,�F ��ۋӍ,�F P��|����C���  �L  P�Ӌ�x�����H  ^��|�����H  ����Uȋ��F �#  ��F    j �t��,�F [���F ��  S��=H�F �E����F �F �����  ���F �E����F �M��ËU؉|�F �=��F �}؋��F �]ԋ=H�F �r�5H�F ���F �D�F �uċ<�F ��E��M؉��F �]Љ=��F �E̋H�F �=��F �E؉]ԉ��F �   �������%��  +��F ;�F �z:���]ԉ�F �M؉��F ��    �<�F ���F ��;M���c �]ԉ=��F �}؉=��F �EȋẺ��  �@��F ���F �=��F    ��.�����F �=��F ���F �]ЉuĉD�F ��F �uԋ��F ��������9��+Z ��F �(�F ���F ���F �D$����F ��F �;��F ��^ C���F �L$����F ����` �ЋL$���F �D$����F 밉u����F �}���}Љ}��X�F �]ȉ]ЋX�F �}ԉE��E��q  R��$�  �L�F ��$�  P���F ��P  ���F �щ�$�  ���F ��$�  ���F �=��F ��$�  ���F ��$�  �-|�F ��$�  ���   ��   �j����,�F ��  �����@  ��  ;�F �������X  ��X  ���F ��(�g  ���D�F JX���  ��4$  �+��#  Qd�5    d�%    ��|  ���F #�%  ��"  	��x  ��|  ��F + �F ��0(  �0�F ���F �\�F ��t  ��0(  ��F ��p  ���F ��F ��l  ��P'  ��� 
   ���F �,�F ���F     S�5�F �5��F �5��F �   Ëd�F @�-��F �-d�F +l$�E�-��F �l$ԉ��F ���F �t$؋��=|�F �=��F �\$ȉ��F �t$ĉ��F �=��F ��X  ����F ��  jd�58�F j �����ËE��T95��F �+� �,�F ��X  ���F W��  Í=,�F �u܉U��E�    ��8  �U����   �U�ǂ(      �=��F �O<��Q|�Yx����5���K�s�{�H�F �C ��F �5��F �s$5��F ��F �K��F ���F ���F ���F     ���F �s����4�F �,�F ���  ���#  3��!  �|�F �X�N��X#  ��"����F ��F ��F ���F �|�F +��F ��%  ��D"  ���F ��`"  ��X#  5��F ��@"  �5��F rX�5��F �?���Ë���F �0�F �EЉEԉ]��]ȉ]Ћ]��0�F ������,�F ��ҋڍ5,�F P�������B��@  �  ���  ��X��H  �=��F ��������H  �  Cjǂ|      ���  Q��P�����|  �l�F ������Y� �F ��0�^  �Mԋ}؋M��[�����X  ��F ��؉��F ���F ��F �,�F ��L  ǃ      �5��F �#  É�x�����������H  �����F    �h�F     ���F �h�F �l�F ��������x�����H  ���   ��������,�F ��@  ��D  Ӄ  +��  <�F �x�F ��@  ��<  ��D  ���   B��jǆ�      P��������@  X�5��F �������=B��jǅH      Z�l�F ���F ��H  Q���F ��5,�F �l�F    j �����^��l�F �-  V�払D  �x�F �h�   h�  �5��F �5|�F h�  ����É�x���B�����F    ���F     ���F ��  �l�F ���F ��������  ���m����,�F ���������`�F    �$�F     ��H  �5$�F �`�F �������l�F ��H  ��<�������  �34�F ���F �$�F ��\  0tA�+D�F ���F ���F �d�F ȁ5@�F l��8���   ���F �@�F P���   Y�  ���F ��  XX�M܋p�F �-4�F �U؋��F PX�4�F  �ԋ��  8�F ���F �4�F ʉp�F ���   ���F �%��F +�F ȉu��% �F ���F ���F �P�`�F �F +\�F ��F ��  �����F +l�F ���  ��h  JX��P  ��F �|�F ���F ���  ��   ӂ  P���  ȋ�P  Ӣ  �4�F 3X�F �l�F ���   �D�F �元CX��  ��F P���   ���  %���S�L���U��U���   ��H  o�d���   ��F ��H  ��H  ��F ���   Q���  ӂ|  ��|  ��|  JXS���  W�}���   ���  ��Z ����5��F 5X�F �M���F BX���  �D�F �΋�x  3\�F �]Ћ��   +��  ���F ���F �b�U؋0�F �]ԋ]�����?  ���F �0�F � �F ���  �x�F ���F +��F x�F C�UЋ �F �]܋U؋]��  �t�F    j ���F ���F Z��5��F �5��F �2�E܍,�F �x�F     �Ủ��F ���   ��  �T�F �x�F ��Ű)��x�F ��[�T�F ��   �x�F �<�F �T�F ���F ����F     �`�F �u�5��F ;5��F �9� �5��F 5��F �0�F �h�F �
�$  �M��x�F     �����UЋ0�F �%x�F ����x�F �5��F �u�;��������F �]ԉM̋`�F �n����Mȍ,�F �E��t�F �5� ���  ���F ���  ���F �E܋5��F ���  �����������}��}��/���  �l$���4�F ���  �E��u��u�+5��F u�G�4�F �5��F �}��u��}��M��M��4�F ���F     �Ɖ��F 9=�F �2����5�F �5�F 5�F �}ԋ}����F �U��E�    �V����5,�F �3�� ���	։3C���F ��V��V���F ���4�F ���  ���F ����,�F �5|�F j�5��F �l   ��4�F    ǅ�      h�  �i  �_F���E�-L�F ��e�������F �E�;�� ���F ��F �}ԉ5��F �U������F ��������F    �54�F hX  W�z���Ë����F��8���4�F t&���  ��(��   �4�F ���"  ���  F��몍,�F �% ���	ЉC���F ��T���5��F �54�F ���  �5��F ��0�����,�F N�Ys ��x����"A����|����Ӊ5��F �l�F ����  ���  P�$�F �4�F ���  �$�F ���������  ���F ���  �=4�F ���  ���  ��T������t,�,�F jh�	  RhX  h�  �k   É��  ��<������I������  �@�4�F ����������  �[���  ���������  �4�F ���  ��$   ���  ��@�X������  ��5��F j
j�i���É�F @��F @Z�5��F ��|����Ӄ���   Z�5��F ��|����Ӄ��   �5 �F ����5X�F �؋��F �5 �F �CH�w �5��F ���F �5X�F Q���F � �F Y�t  X�ʉ�t����5t�F �=H�F ���F �=p�F ���F �=l�F �=H�F ��t������������  ���  ��X��x������F ��p ��@  ��>����|����5��F ��x���@���F ��H  �5t�F �Ë�F ��H  ���F �5��F �  �؍v��   �`r �5��F ǅ      ��t����5�F ��  �D�F    ��  ��  ��  ��  ��  �5D�F ��  �5��F ��  � �F ��  �5��F �;�v��   ��q �5��F � �F     �5��F � �F ���F    ���F �5X�F ��@  ���F ��"����5X�F ��@  �D�F � �F �H��q Q���F �D�F ���F [� �F ���F 룉�x������F ��H  ��H  �ځ�$�     �;� ��H  �t�F �p�F @ǅ      ��  ���F ���F ���  X�Ӊ5��F ��|����������������,�F ��x������  Q���F ��H  ���  ����d�F ��F ��x������  ���������8  �d�F ���  ��  ���  ��  �/  Z�p�F ��ҋ��BH�ou �ډ5��F �5p�F ��   ���F ��F �5t�F ��H  X�ʋp�F �l�F ��F ��H  ���F ���F ���  �=��F ��  ���  �@��t\P�5\�F ��H  ���F �Ӊ�  �5��F �5��F �5p�F ��x�����[�=��F ��  �=\�F ���F �=t�F �l�F �=   �(� @���F     V�5��F ������Z�p�F �H��q �5��F ���ׁ%,�F ����u��5,�F �M��M�;1��� �u��Eĉ]��}��ً=��F � �F �{  �5t�F �5,�F �[��d  ��H  ���}����l�F �5��F +5t�F R���F �֋Ӊ��F ��P�Ɖ=��F �=��F ���F X�5�F ��t����<�F ���������F ���F ��F �X�F ��H  Z����H  ��r ��H  �5��F [��|�����H  ���x�����x�����H  ��  ��  P�5�F �=T�F �=��F �  ���F R�΋T�F �5��F _�5��F �=t�F �=��F ��������x�����  ��H  ���  ��  ǅ     ��F ���  �<�F ��  Q��  �g  �E�    �=��F �U�;U��K� �U�Uĉ]ԋ]�Ӌ;�  �=�F �,�F     �Uȉ �F ��F �	���������F ���  �,�F �}��=�F +=��F =,�F ��F � �F �=��F �}�먉�H  ��������F �T�F ���  ��   ���  ��  ��x���A��  ��F �L�F ��������  ���o  ���F �Ƌ�x�����F ���F    ��F ��  ��  ����F R���F �+  Q���F �����X�5i ��C��   �&  ���7  �  ��  ������   �����@�B�����  ��H  ��ɉ�  ��H  �������F ��F ��H  ��x�����d  ��$�  ��  ���  �5t�F ���������  �Ë�=��F �����  ���"  ��x�����F ��H  �L�F ���F ��  �L�F �L�F �5t�F �b����,�F ���  j��,  ��<�����x�����F Q���F ��H  �5�F ������ۉ=��F _��N�����x����5�F W�=��F ��   ��H  ��  ��Z�<�F ��  ��H  �t�F ���F ��x����<�F �����\�F Q�5t�F �-p�F �D$�ʉ-l�F ]�Ӊ-��F �\�F ��ň  ���{�����x����5�F �ˉ�  ��  ������A��  ��F �������H  ��������F Y������M����A��������R��F [��h C��   }+���7  }��  �m�����   �����@����������������������V%p-2�S�Sh���IU#�c�7����1�[s��_���u~=AW��7�=���<B�%�]�s�e��Ϯ�K��8���켼����fpu��[�!��X@Q��N+g�|1�(�G�
�XD���@����t����P�Y�t��|Z�F_iW9�s�����}Jƒd��C��+%?E��!�f٤A@t�ֿ�A-�}J��:�Q�
�`��Q��y�{���r�^ W�0��d��RQ&���>��=���}�xgy4���� ����q(L�:M���@����:H����g*9������땛Ba�gR\Z�;�"��L>ɔJ�
���hӉ����15@�Ͱ�PY�F�]�Q�5>06����`|I�����3��Z�}�I������R�ێ���o�I���<�$F�-0���?�;@�D]�6�Ԇd#�FE�4��ڠ����O#�Y��N�7�@�T[f��D�Ô�Nj ��ܚ�.�䡚�y�k@C�����u��A&�U�:�5���(�Q�=i���S�I���q��*���gz�%�;U�;pӗ���B���U�oi<?�� ]s����n�̈��{�x�O1}�U��()�c�;���H%��*e�1d�Zt���Y�'�3_�Hs� )�l�U�
>:,�/	Ɂ�(���x�j:��V�]��ɂj��لLI����)��b-Q
�lK��B�N�򗜖�����;���Q��a2֎	vD&۱~�g��	�f��Q����f�n��"�3_g��q�0'�d���F1T��"$/�rE:F��*����p��0&��촼��ztOX�����B��T�T�?�g�|�	�R(�o�Y�U�¯�9��)�x�Z6ű��2{$�ƴ��Ķ�Ŭ���k$*�6ok�t45��[��L��3��uduv"��v��lqJ鞄��r7�B�ob�<>r��@� ^�Ҵ�,�A�dx�cT4���6�&Ȋ��Q߿\ �0�>y�k�!�'}F����q޽��3%�:���:�0����d�ّY�K�
�mnJ�x�.>5L<9ME�l9&2Hg���G��U�~���ok���٤ew�V��}�Aն������sU�%T��;��hQ�m@�W��uk��e�_=��v���� 2���L؁ �㫹?�$%ѤR_.ƲW�q�kZ5үl�x$":����++C8�f�d�	!��RY�)y�d(��ꭓxA<ER)S�[QxT��h}�N�� �i�6[����1&�'�<K�����U��Qٵb�gz���'�� �ؤu��%d= ��5��b�����|X_�,-J���-��3u�<�I坸fkN�Sm����.�����>�jҬ`}T�0 ��n4hKԷ���*s��Q��R>^璓�y�N��ɻf��t}��WY� @C�g�^�*c0M���a+g A����)b�T��czf�^�v��U̒Ð@R�c�X%`��Bd9j%�^r9�{R��c�N���,8���Ok��@�7-�kH�GS��u��. q���~�Ր�(T�3b�Y�@rBR��M>H�D2��l��&îv|5�#��
��ɗ�f���ؽ�p�<w[��cFJ��4�e�W���m�jsS�
x�T= �9���!W	Y.��&��}B��+i��L���N@YX�Sgn�F�q�گ��F@;ΒE��:�����c��I�]�I3O��+��^!����V�������H���It�p�^��*ڑQ?R1����c�,O.�N�q�uQ�������ٍ�o`��Q��@B�E]�9b�� c� �F�DD�q��k�9������}&B:f�u,�Vy�%_�X�-�G�mF�@��j�Gd)a˥�=�dfw �?��N���zo��)s^�sH{���κ���S
����!d�,�K2՜K.�	e���Yc��Ky�\*L_� Y�AM]�()��+7`��T���n�.��Xǖ;'�ci0�����`x��E �C�����*��>��|���,��(}2;K&{�	���#��h����M3D�P�\�ҵ:����Q?�j�Su��_��m=DH��g�P�q�(Xb��
/�`���� M^�Q�"�t�.���LvC;�����cvQHaM���΍��*j�˝��:,��X~��!�W\�/<՝�!��62
�����.x�������a(�	[����p�f�x�!��C�bWY��V�6�aZ��nߌZ������ҌD��[�Иv�72���~���ȹFZ��Y9�$.`��s�l�t
���'9黺�$�A`Yo�CBԗ��MLfA|��CU�Zǝ���A�u���0R��YWy������i(ܽ�##Z�H�;�W@*���޻���#Z���t[vI�Di�m����B�c�N���&���Lۧ��|rک,����	���@�������w�HJ��K��FL��&�<P�AQ�k;1Yd�Suo1��*X�PlX��,4(�kVW��M���0�J;z�B����@�ڻ�S\A��Y� B0�Rz�$)�a�ap1�bU�,/�X�0��eL�t�v���H�W����S~�cH	� ��,Z<X��J��Y��=�6ncnJ'�� 9= ��y�v� gN6� ��oQ@O���Yo��)��ohs�#����å��s� ��r�y���	҇1�"J��k.9ќ7.�Ʋ�x4��u�u�.�}	V>�&�E|�Y��ĺ�(���#5gs��d��]�j�$֜҂�]�9w�ˁ��D7�-�6�i��B�2ɐQ9��PS�VhUcjv������fZ�V\����D�]s�cB�S�vU�g����%��U��١wש���H���S�������L���~]��R��s��a4H)�y�ZY?l�Y9�'�T�p�=r�p��2x�����S$�$q�R��"eܥ�'�jK�?�S/�͆��@�
�Cl��h�%|���e�`�%���G\�x��Q�oIN���8�b�M���V��9�O�>�׸�Wk�I��'���#11�?��4�[Ht.��i͸�8)~�~�+�V�gU dqP	�x٢˅Y�E�u'R:���o/��rK�I}�J<�eL��1��p.*��~�ˡHk�"�D�EO��Z0J�멇�R��\
��5۸h������_[�X�����Ѭh`k�.5Qj�l.�W�7�uj��(�P`Co�{?%��y�j�>�g�(�
J��E'!Wh�>KM�n�d��a�<ެ��I���ʾ CR��2(��AXKM�p�g`�dgث�j���c�xVVB�]1B+:	�ˢ�#�jť5��b�����qwT�Լ��@k��L�k	��gG㉋���n�z#��ܷ,�6�����n����k�7oP�Wz!<[u�ܞ�d{O�oNͷ�[����4r���B&�<����
�XIHyW���֣<�G��|�GJ�\E��0��k�f��F[�`���pZ��s���(���A%�a6�W:1|8�L��%���"���!�d%Cߤ�w��I�$&�?��6�Q����"�dD(�ݾ&���[��ӷ9��wC�Μd�!�������f��s�M��N>h!�N�*�GgvS�GZ��Cj�`0X�v��	����>H���v����9a��m�O�T/�����K�x~���v�+���On�Y�d��>�G#꿞9��*\׆<�跮dNs��F70�A��Y���
&F<�~{�ʊ�6f��A-����_^s��^�⤪)<@��&���-�v�&�B���?'W�:^�'\O��l�_\�~�����i�����D�Lx�������V����a�f��*X<)�3n03��5�@�Js';Ȇ5��ւmkW��n��'~Q����<������,|ɹV�b����p^/��_TG� �E�G���c[.�vL�� m�Ye�M�W���9Zh��P�wRXxxʦ�hif;�w9r)�brB�	~�����n�S�<ˌ�����3����ω���_<!>���&�L���͊	˸Lk0��Ii0����#g&T�L��������*/�;/U��6s��e�?w�������u{@96{t�NX�)�zD���n�0!��r�i�q���:[���O��VÍ1��T�X�0�$�׊��W����Q�O����ۻ�o�Գ��{��57� �/�5Y�C�ޘR�8��h�П��]ט\ ��_�k�Œ�jat���@w�ӝh�fq�z|bX�%m;޽DƤ!:�b;�p�IA�z�?�)��\g�Z�����>�3�(�I�r��9	�L�;s���Ih��<�2q�E}/�'c��dX��32���cuV٪ӥ�~�Y(o�sX���Ic]�D锓g�=�E��-�<�Sl<��?ĝz���\�
M6���D��U.�Ja����zTP\@�:UF�Y1N�I;9�S�N��5�ZKT�r-��p_�ђ?�4k���~T�^�����$�8]������q���J��O�e�K�/�DnoZ+e���s�Af����N7�BH��.8l!��ѥa25ӌ���?� ���?5�E!���b����Z'@�0/�7��K,h�xT�d��]�CI�)$Q�G����[�ȦA�U#X��)��.Rg�xRF\�;#U|�j��qّ���2� �u�!�0�B�	�)d�����dT���Sc4<{.i���:X?	��B��т��-��]��<�ڮJ� K���kf	��k��ќ�ݙfբ+��l�x2��3`IkL��~_�Z`?�<<Xs�R�v�b�W��7�I]����$�߾��D"C��m%��oW�7�`+13?j�خ��tmCb��7xVo�e���G�9!���l9~8U��
y-�O�V���l�)��E�o�^���-�·�mYg��T
�p:ö�R$������f'�.�]��eb�,�]\Mc��l�j�hث�Ί��!��E'	|M"i�|X�YS�
����H852�d�����Ľ�c�K���S�� ��Ll�փ��u&�ۋ
�����L7�:k0�@9�n�aظG�!��\M��y!���t\��yq�u���^I@e��������Y��JQ�+Z�r�E�3�ARS9�Th��� ʤբjZEZ�yxy$�4�b]
脖#��>a�(1M%�1*%�!��7bz�&���qoE�������gu�#���� ��m�G]a�fYq>8��ƿ�� �8��i�m��j$*H'�� �vYVl,w�bL��Κ��JAa5��"(�S����*��;qqo۲Nz�T��ǳҿ-e�o�(��!����) 5m3����Ct-��"�W�����.��t��-��T]Zch��/~\ ����{0`,F
-��3ub��!�-���~�a8�����ګ�I�߫xEIdW�7JFJ ��>��$�Wr�jlғ�͔\�7�ȋ��sy���p}p����\%��N�WnD�)&D3�]��5�1����V�F�rPj?E�i�U�,�!8�/�Rl�����lL�����V�g7ƚz���NF�NS�Xw�!�k�>��kg�&�Fd~�U���ú�Dl$t��4�'>ruX����m�H�6$�J���	k�ߴ�.��Ka�#�k2
R�T}$@J��f�����-%��t�1i�V�c�8Bf���Ă��f�f�S�u
�
̫ҭ�����9����Ou�I��Ў�t�4�'��p���6���W_͝⠋(6xj�P���-\o����$��k���:��_��FF��:�V�J����yJ������gU�Y�&�"v��K�wɗb�����ކ���3���Ѥ�c2[\{d���0��t��_�:v�j��(�(�G^�@�'��5��'�P��8��I^��D��v�0nM˚v3ۇ ���*�&^�Iد-�8F�-�l*\"��������,����Pw�T�8����i!�p��c���
��m,=���a��.w_fl:�.�i������S��/I�aK��!E�B'�*�?0ʗ��y��1���)�+��䥃����F�qLf���\*��=��Yh�:ET7
��\Z�)5�?��
�9
_8��D��e�{��8���"N�5���n��Q��1n�/�fn9��
z�J������ve[���	�4L���:�@`?���z�hwѮ���8�M�j._Y�j�(�� v�G�E������Y)qD3�;�{ھ|ftȢ��Q�� ����o.-u�]��=W�x�e��O�������]P�`@ �<n�-��G����� ҝ���998�r��+������r�2^PMg���г�[E��! �Tk?�I@�2�x��Hӎ�gb��-���;�+���O��ǘ��1?6x6����]�U>Ԅ��Ƿߔm��ou�s��]�pd���d:`?�bkңx��c�\�
v�>�m����F���R�
��yx���Y���{�B��Mcc�~���a�܋�_5t��gH�A����]�ܬN��5�3�A%�1P��N)\�)���%F��o��(�N	��׿���u��Й��M=��qV��WڂM�R���i��q��7'�5�Z�u
.ʭ	W�z~:��jKOp�̥�Gsg����)b ����;�/��&��4o:)��L�A�r�w읍I�dia2n�-�[�ʶ֥����[��
�F������� �v��r�]�
?���57p�$S���ηW���?/�7��_,�ƒa����;��O׶[�,GrW��v
�vZ,}�����o��[�ڟ�2��\�L�d�i�mE��)ǥE)�X��o�y53��V�]9|��^p���}�浯vt�I�Q�{�A����"��4�{�i�d��6NVFz�clw�n�{��VRz'��_��$$�B" 8�k?��Ӹ/:�˅8�'��$�Uw\Q���PU��F���[����ӛ�qd�A��,���+q$3�!Z��3���� 酣`��qc�>�?�ͽiG�m�@G�>���*�M{J�6B�lv(�^M��TΎg�A�@se��m��6�=�0&���8W��u���r��d�Z���XD����C��$�T����k�i@Ӽ������e�BI�;�iq@I���-��1
��A��-�5\��CS�F\v��k��=�/�4����W�j���J�lP:�#	��vT�$�ɶ} �7ii*����ui�v��B��y��iԺe�
J$��/�*jN&���;2ܡ3<�ދK�`�a���@��F\޼ouJ�i�	D�&�����?��|e��{<���Qs҆o����.�`�j@�J^�JX>.К��*��r�o��6wTk�ⰶ�sG��J)�M��=&ww��@��Pf��_�c�7���[��uY�eUF�-�֚�E�́�WX��f�>g�����"�e��n�4h�Śv��Bl,�r��u�0���R	�R����'r�g�:���TD7��Y�_0Sn���aǏ���g����x�m}4��+w��Be:��N��>vY�U�+�_��h��6���'Ia�tɾ5�b�Ք7�e+K��O/|����hB)
ּ�����@��s�q�ꢑn.�> �+��̸���k�5��^EQ�*�� �,�TL"��@Um�<R�j��L�N�e��������9=�&S��˰�D0s��@0?
Ԛ~�o$�tQ�!��c�raG�"���G�]�*��y��ȪM*޹ȵ.߾���BU�<����箄x��<n��
]�?5�/??W�|,��s��W�	��	}�����!�$5�#�>���ڥ��GC^����&'�oy�38�
T��߰�֡R]]	���#��D�25�-�����(����ПfgҺ�c���˭�gQ%�XS�I��
��rY�bRBG5�d���V}�%.�Q��Z�����bc1P ��w-����AB��������Y}���^]N���5��������n�bQN8�r�jj2��Q H ��;��x��I��r��#��z.:�|�.v�Ւ�T}&2���H"���Y+L~���f��+"=E����C����nk������[���?UC�Z���-��~o�.���[N�h����y����]IF[���1��x���v`�M5cvo8<��d���ꆓΩq��	�4��W����6�t����-]�7�J�oգJ�=A-�t���	1����t'~�+�M$�e�ˤ�a���hc�-���p��q�_�
Pa�X���|�}�rI����07-J��M�0/�ċ��xJ���m6$Mk�S��E��1M'���Lk�(��۽�Ɇ
���@�Bk�+b���#~|7j�n�9���Ȭ3���	޶q�� ��j#���}�����L��[s����(v ������7�`J�RA���n˞��W�Dz�9��с�~��r��)�*��F���̞�󱠵A
�'x�ߝ3�Ħ�^�Ia�-d-��`C^��7�UZ��$bMO��E>��ߦ��+����,��K{F�9��f;��^�EȰi�j1&M��I�)��� 4l��ۄfx��˕g�ئ!���%U��TYX��_��TN�������(
�S��6�ެo}���s�Ҷ����50F<�~2�����u"�C)EVԤV�s��0�D9�e0o*�Z���ط�U �3�a�~��9}M?��\���%�*ū������.k¨W��O���*��W{��H�D��a�b1� 3Z��<�Z@���t���۔C��h���{{�(%���J����D�1�`g�hVC�u}��7H�I�N��ۂ���
�e�=��PU%[��K�#�ǌzu��ȟw�E�Y��>+�+pn�(�W���@%!��m?f���,�c�*� )�i��5�{�bC5�=t�d������Ahˮk�I���$>cƢU���|������5�$B�e'J������T����n�@�`���\H�����2�kfx���Y,$���Ћ80��	Z��Z�+5IQ4�'�����},����3y|ǸD�ȅJD�C�a'�M:�ƌ��gI'����w�uSx{)��f?���gw���CG�
��c��b%�Myr8�)���������X��'u�]?N����z����#/
�W�R�!w���� �.�(�yM;̾Q��>L)YYA�,5%8�[p"B��E�(��|�e��Ob�*�噞><�����w::6�/g%�'��M	�돌�"���nA3�T
4��;6�� .�í�dDt_��I\���9�Sf�Cp6�C�����h��-{�8ʳ}�F}S�qg>s(u��Fo�r�p�r!���-y|%b�^P�~~I%���H���0��8��9��+:���M��5l�T�e� �jY^:�;�� ��
���<�U�:�7��|w=��eh�߇�;�ֺ߽T!Q&y��d�b�b�K��{p���(Ѧ��������4������9z}=\z=��*��[�z��[�!�;��-�-enUEsʦ�~�o�h�ԚU^{(��ȯ%�x��ⶔ�(D'U=2: �(�s�u�WR��[Ꮉ�g�U��r��:����Hml��EZ�S���HO�a�u���;����*a�X�qF��çGm �2� .������=4_�ldM Һ��vI�?�'jD�o�CO�-
\��|_U��%�Rh�F��N�y���Ce{���(�?=Q�d���Y���"��8���oUk��_�?�ӧ�?��*�,0K6쉲A�I�B�W�4�ޱ9W��N��p�,�ŊOt��(�S�%N��!�\�v��P�X���w�����!*�K�񸙴H�ؐ���T��n ��u����GV/��p�?i+����nbU	�yqU�78$�/�h����#,t�=��\�z���h�志���FȘ�b�c���Ч�o�V0U&'NL��H�O�$�Xn�V�qצ�!u�8�K����o|��U�xX���	��������׀MޫF��k��Y��`D���z�1��-HqK�0��X%�-�يQ�Zq�S�I<5z#7�ۢ�a߼C�L���
�7��<���+���-4@Vp�X;��~�k������W�( ��{Ζ���mC�<i�2g�;�&WAu)$�����N��E�k+�ɂM.a���#��t��Yτ�
�ǈ��q$,���|�<Z�vhǗqgE�	zШMI��w����eũ�l���~�Xu�Y`4�gwD�u��@�j��BՄdm�z�|��3�����;��C�U�K�軳����!�E1M�0�(����Z\�%fV�:��x���hC7��Y����������u1�\zk�!�nnW�F�V[�2U�#�=38��
�`k���I[���f��!vjn�m�SQ�3 '%"v�~ۃs�n��"���#��{��ѧ�`����Fu����Y�4N��ûn�ݾ��;e��'�̒�p��[�3S�)�x|NDb!���;8�U���%����I�c���7/˪zs��Ͽ6�
}	6�g�L�H����qO�-�h�������MտNHq�;>�D�ش���G�6'H����ˑ!�ܯܶm��N$����e+�#4i?� 0���u�7Կc��7f���8�Ȅ.\�=l+p��`/�9�w`�.��&�,j�j
��X.��0���$:�Mbk@R�Xe�|lq��rZjJ�QL
~Ar6��/��DQ�
#F'&��D�B,8YU�(y�'Ri�	��xe�ۉP��#&/nO��OX���9������y����=�=��*��N}�(�|n���'�fi���i]�nx��Tڿ�&�oB��B^���(2b�)�+Ͼ�X.�I6�̅�f5ýA�b֨Rޟ�S�H	{�7��|���h��	�O�_��s�3;6vb艹�l��P���G\���y�H�aaLd���ۣ�=���f�߽[�т1��厁c,��/���W�;�ف�����q���Uf��W��j�G��U>�k06���a�n�������"Bi`p�L���3w?sg����%���0.1��n(�r
��vC�[ ��8�N�m�ŰŽ�?92�m���`����'��Л�I����*�~�ZS��.Ԇ�d
�<�"���n�pKQ��"4=w<�7H�����}m�6�u&�usά`[�Ϫ���C����il�]A��U��F`���u���UJ��َn�����|&�i���{��f�e�J�a�~A���Ŗ�↸�,�[�~L�V�����c�)O�#��� ��B��DgU���:t/��ՆZ&g�UȤ݁�z�V�M��xۃ;��pm��-w4��� ��JSB�-��0$�f��!B+��3��G�4+�We�lan��X'g����^p3Y�J�b�'Yq>�l����U�_��C�(!pC~H%&��'P�8�G�۪�ؠ�$B�ԡ�=:�� ���u<���.5�Я6����i�k��o1�}~e|[�^T�m-ua~��KN:L_X�L�|�>�S��"�-Uv�_M�;L�_�/�D� dud�|d�����+-´`|����Q�(���H���c�<ѦMk!o��SD��f��#��|.Y�ݝ��G*f�G���)�D}g5E��L�!�p�nVJVp�W,}H��}-Q��%���<�X]�o��̈V��8�Gp.�8��fy?f(�����MN�7��J\ފރ��|ڠ0����{W��������vp>���6s&nK�(_��9�Ԡ��"8jk�����Ө�T�c��P�2�5I���m�ǴRz{B�K�):���ݘ�����E��_�L�ݾ �fA���)�(�=	��v���F�)$��E܂ώZ�]`k�yOds����w9غ�ot Hu�G ��g+�a��?�V��<��;�cL�aBg��0X��:Ѩ6�^2ޱ�ĳ7d�ϣ���Z���-�1֡���Bf�'+�I��������.HP�w�ղ�e: �W���66�|�;��tl��������"hu�hς�e2'�E�$����BQ�S)q0v������� iT�.�]�YY ��L�؏u�֤61�������gA�"dC���{*�C,��TԤ�JZGZq�Nv��n�e�y�®�b�8E$u�h0����G@�M���S��L#;��ֲ�b��Q�=Z��0���������`S�6_Me�j��C������]�u�ClG�!#��R�T�E�%K�����*�Y�v{���� �/�3g����FcK�������; �ɲ���$*�5���@;aA�ǊƁ�̅B� �#����L����{�_�LZ���s5���"��ln#��0q��{��Y�d88lk�|����[iK������
d��St2��h߄35J"�G��I�5^$�v�ǁ��7����N���e�OXu�P���1׳R;��ݖI�B�����GA�y������l2��GFB�`��.5\�Ȕ��Ė㷚�[^�
��A��JyES|��7C���*�*�j����P(�$��>i��c
��f���6u����6)����:`[�+{GCk�:pm0�^��*Q��$%0^�UBX���U��*^�����:�%�+B��B����a�m��5[]��[�39�w��s�ۮea�T-�1U�,4��D^�4,������G�s@xq�}���:`��SDٔ��*�R{�g�T%Z��1���3�o[�"�Ke9�F,4k�;��M����]H�gb8�p�!	����*|�{8�r�h����SC��"���3�v��0$�_(�:D��X��>���C��Rr����H��%̀S>%a���!!�O@cPE��S��A��]~K!�9Ȱ<�K� �4��AIeU�����9gG�N��6���?Г謅+�~0~�¥��A`$-�c*��BbML~����۟��x���l�DT�'L�n.��n��,���X�\周}�V^��a#��vb#F�6��F^pp��(�3zH��r��xo�~cgQ~�w���$՝_�ex|m��ep��S+����ڋ���������d�B�����Ll��e-F��2�0��6Ղu
bW���#����������v!3�4���>�����s�^��eډDO~�,��f�N�!��YC�K�12��w���G��,��jH��kLMu�����n���c�Ȝ�7ha&U�6Ǒb��5���:�O$uu�Y��I�K�Fx�`W)2��SU����)W$cE��:W�������+_[��#�2r��U�F��\˄��
M&��&H�� I���
<�f��gԉ�\�zT�i2��B�	<�Fck�8�Z���˃�A�4x��x|��*�S�;�����2��b+�}7���JOAIGFG�֑gw�φ��v�Yo�Y(*��ֶʧC�4ˆˎ̽T�u#�@�ZY��8]d�j�� tN`�4g}�5��i_w�$]�����}Rw֬D�+�_@}��:FcDX0��Y��oK̿��ca��P��ւ[���l�E_���.8=�y�^ic��3a���v}���G=hP��V�X\i*W�1B��cW�՜l��C��W�{�)?��<� ��Z��������$?�ۇ�.� ��`���Q��PHRvD�I�����^Y�#�y�*��9=�u���Q�w{��6"H��8�8k��t_Shb7�Z�"��0/R��#ӽ����z���yX�	3±1���2ٸ!
[�u�i=��32ֿ���ƶ��U�I���!?`a��ϷP	?��?�#�Z�\�pU���.߿�t��7�zE��!�| �J}��;��T�sY���:b�3����tT�Bp������#|	�8��H�,#�~��i�듲%� ����.�5?rU����>���FΩ��&�8��o���鴡Z�T0[�F���ʚiO�Ќ��2~�U��@���
)�\����- m7˾O�J+l"����YkDˀxXffh
i{i�ۈ��������P���_���h"����?zk`�&�5�������ٟ��@��d~�F�x3����_"bKʻ�V6�ɧ��<�â��}n��΋~Pk�,|-�o���9�I�R�Ѽ��1I3�-���R�&���b�n'�����}W����?y���6�c�b���p��v�����c�!�g�!K�4&C3V�๣�"���q�>>�z_N�r[?���0�޼����H4o�	�7��b�[�#�W���>3�+1y�KlyVy�6�G��,ǦQ�\S�2ܜc9C�����Z	� �M!��LZ]��eŞZ}�ES4��
� m~ڃz����~�Sk�B���%g���8� ��W��g�wRb�����0�^�a�.�y�V]�~�����ad&>3�T� 9a��Q�����)�?C�_�F�M �vtL/��\���`^�+aa���Z�:X�M��dS'S�~���H�վ� �K�ڋ&�*_>�{��+k���Q�G>aͨ���� ^�Yd%����������ϯzw��()���k�u��U�klMu�4~�������T�^�ӐږBӐ��y�c�+��m��<��)'u\P�;���I ��s x]���8�:���z�D�Q�N�qT k ,��O� ?�ϟh����E��]����5�+��U���h�����\��y��[jQ'�(9��m�sCIX���f����$�'5��v��+i��ə`�$��i��6\L� � �u6T�)�B3珚�a��ī�ĒVM@���|��=��OT�y�����>!�S�,O�C�ejQ1���%���m�]�V��X�|,��~���G\�F�A����dW|g[���G����4���wx9G-Ӱ}���94�N�v�T�����{<+#)�>��2���u�����c��`M�dM��xW��l�L�>V�aV�{CL��n[��w
�H���4��N��~.�Nz��7�VS�r������=i�\��R	.4�Z�f5��r ȎK�
Ҏ�~娄�하����	�عG?��K��U��f>��$��WVK��r��Q�t�w��?�����z�)nJ�8p����P�ƸS�;`:�_=�Z˺��wQK�P�~l�����|��
��D(�j<uhp1g	�.�z'L"k����ʈ
}�6>I�+��yn�R�7��(FS���� FQ��a�F�FG$�Q��U�;��P7��7\�Ɍ�tE
��M2�%$�Ԇ�@K�w{s(՗U	s� �j�	��e�>��f�ju����k#u�΀�n�����êU D���ҁ���M��<�J����t��3���'!$.Y���&�U3F�`�8k���WX��֬�v�ݵ���do�`tL�|�����D��������n�������c ��'[9�S��'�4A��6���@b�`p'� ���sb�,H���sZ;�bӧOF�$|����Zr&���_
7������=e`.�4��sM�RÞ�g	{�$�ͳ�7�%Yy�@}�B?��:��bi0nxeY�����?�k�_ t��21�}����z��ykf���g~��U����f�q�J��L��pTg#�'Y(CK�,F�����c��kA�Tس�����G��M��*�<��/xC����֍�'{��,��Iy� k�2V�����!+� E��9t��B���aK�ۄ֖������ SF��	�w�r%�H����8����a(b�|,C�K��ġ��k3��҇�&ϊ��޵ћ	s�u�(np:V��T�>���Eej���OW#�5=�7
���%�����b�"�F�\US�:��C�<j��<g�������5d*�U�an���z.n��Ҷ'�����AXkuHn�L��q<8cK4�����7.�
����Py#�%�_�,[`L��N�P��8��������lC��f���Pk�l*��|�8�W}vҩa݅�=Fv(S��`=Lb�WE��6������B�>���P���8�Z��Lb�c���˳�.7SFb\I�u��˓X?��ϯ���4�V�vp%=�II��[�g�����2��<��_�\��`Y(�'b`�o*nY�-���7./��Y��,�hx�N�p��F�M�8SrYb���[�r}ɿB8�8�Q'�Np��e����)�:/��y�h�GP��]����%��5�x�p���w�q ��%]|��(��k�evnDÒ��E� C��[�@�
z���Uܱ�b�F�q¼z
�	�+���f���;�I�ŕ30N�6zIl=���W���(�ι��͏���1��{n,n��s�Y}���=O�z2x �I틱3lV`l�+،����a�v����̘��O��G�����ו�a��XBb�u��8�5Z����uAl7��J1�$�[���N��m�z�����t�@%ad���7S�*����ݎ�D*)��7�\�	�5_rq�& ��9�h�W���5d$g����&�$=�ܽn�D�z�ja5h'ְ���#�b���ߟ-�Ѫv�4�;�:�,hm�(�=�������)��L�־�3L�d�,�OV��~�8�l�~t�t�$4H� J1r�Fڟ-/�ۻ^�.�&6c�|���)��M��/���{�� �=&�68%�:�$rx�.����ka�,�e�R\���U�դ1�?�|��$W�8-?h/d3u[pty���-vM�`�t�5}�QeO���^<-ݓ�Z������{��1f���-�G��K�c�l�i&�0aU(��5c�8��#�T��tly�����KLwDUz�1\���ʢ�h��o�����X�>Ƶ��HZM���Ss�0�d0��X�����Ozss�d�"aT溉�#p���a�.�rC��t>�wIhd-0�	[�W���D\O�
[�.%�e.(��2�Y�)�f_�P��X{�8���=�=|.x{CO����&�=
ڌ4���',�:\���A W�� �-j���[,+�\rT-ht�y��B�tJ�z}�h���`�������Ja�.����q���T-&t#jfr��4�oGD�X���^��84���׏-�o����G�U��Pd�{�}PX[��P����-omv�@��X�#3���1��MQ��I����	@�v/F]]#KX�g��o�m��hpk4�@��-p�M��=���X��=�}�A^���̰���8�LaJ[`��nD����-~��!��c6L�1�UV\:dw�v�i�|mn:U���(d'�AMs���O��-�X����0,Y�V�'ؿ�!Q�iI�Ah��$�8ώ)���߶)�﮹n���R�Q����z{F�^ ���`��o�[��?r��2���_�ܠ�W����k�%�"�5��p��w�V\˄'���D
p;�b{Y�=�X� sC�$���*�Q7�ᕖߞ7������q�
��Ƌ�o���>���~Tձ`@���kNa�xP��i>@AX�����E��Dm;�U�����gie�u8�}Z��pT{���N���eL�Dk���=�L�P�/��Q�\�BC���T8Ijp�ԛ_.AZLg��d9=G.�>��}��'wG�Z��I�	u�k$���c��N�au��IP�w�Zx'iP���@6�,Q�����>4��ee���<W'��Oty��^z���>)��y�EU���y��K;q���
^�9�9iT�R,6�>�� ۫�Na�^�S���C"�Ft=	�	Hg}�͑WK���Ӱ����䝤�?�@�����K�'�JZ�F_�5��~�������q �iӕFt���ȧ��w-��˽=�S�S�>���@���;��������r���O֗�u��V������4;{��4!�!���P�O���]S�*X��^aJ�b�r5��m����gPc:{�q�{ y�OtMv)��ț	dq�º��m��R=����;�৕R��l	�Y�-a�C��z-��E�%�_w�d���[���mܴ��r�����N+�w�q\�a��������q�:`ޮ��������RL�(�_T�`J(��{c�e�BKsx�T;ْ� z�Vor%~Ś c	+�X?V>��P&�`��A����(��Ǒ�%��寐�_头��
��*n����x��$���	��g�l=Q�,̱@a��<W'�n���1��f�Ho-��&�����%�����L��xO���-
;u��m��0%�7��^{	p�nT�I��aO.�hH��P(��qgz����6�Pq��m������T?M��;����Mh��w���P���Z�Ѭ>�r��3 �fh�n2�$��t��	�tc���1e��f�+	��n�Z�U6������9n�lV)��m�.�I�\��=�s���.W��&��y�{��<B�!��..���IG�V�1�v�(��&z����ġew���p��$i�Y3ɿ&4{�ӄ�X�6/��������V�����],� ������͵=p=(�j.��#�@�Q�9߱<Br��G/����0�x��I�I�l}�2-����ko��'�<�=u���D*�q_��5(�z��-��}u�l�?<3hOU��J��<�Y�Q.x`�_��x�J���@	$��(�m�h�'r�O4��cK���Į_�GM��dR�J�Ώ������c?:�M�5�Ϝ���̅���}_�� (���#tP�.��3�mo�@�|�rW�DEU���	��V̗=�D�;L ҥ0g �2���4�5ܿ����-R1I�%� ����,֔�QE��.�v�z
M0d���ȁtڛ�[��O�3`�-�N!O������>�r��i>!|�b�G*.3~Z�A%�,��z���jp��K�`�:�&b\m,�,|˾�Z����8�2��`��(!V�f척>��4�r?��FB/�^&;wߺl�b�uءz���:fROtA�-�4���0���7�w��D��ӠH�zu�jKJ{<�a��S�mmқ��MA�S��W��	F�|І�Q��	q�����u$�+@�L& �a�y���1H��)H�]|]��\t�&��',��"R=�h蛸�p߱�V#�LaP.�N���nx��$�)������ץo�s�(��Q�7Ԡ�N8�柄ӲU��BH5ސ�Z疳���d'�����oɌ	E,-�>�Ά�-H��`����3X����f�iqm�2��	rS�a3G��z8�f")�!���ឬd��c���TX9*e�e�!�t/#����G�(߃�L��L�-�ws�#����ko���?0�Y����.�䃁�4�����G�fD&���.�F���GG�������MF��'�*(�ˋ��`Y>~jM�	SQ�Z�;����/�Ӄ��6w�dL�2
��L;�`@��8��s��lG&�������ܠ��k���N@Zn�vR�ckIޱ=����L2͉Y���Z�9�WU��z�|�ie��r�(����"`s�Td6�\բ+ra��,���B�N�p��L���?���ҹa��"b����@J���y�O�|$���J�d�Sm)�64&���.&�V�ݰ�殓��̋��}$�Ky�<�{�y���cE|���=b���$:U��[��{��������D��a��b��J��J��4/3j�N=Q�ׇi*O�h��BFFM��{F�t���t���z�zI���b	�в-��&[��
����%�9f�c��:>YVm���y������m�ۚ��h�A.��N`��H�5����8�3��ry�e�/NO���c��J�ߓFa'd� :_�S�-Y���}���}���:af��I`ZR{��k��0��匞w=��<�������+��jZ0c���rMK�y�WM�.C�tؚF-��1=�|S�/wo��w�E4M��\,�� if�q�ش�K���7��܅#��7Gu����������(�/s^Q�i\��N�-����c���׵$)���W�9���O�c1�z�FX僊r��᲏AM������ש�Ђ))��sն3N�y8as����k]r�r�߻�����R�&�������ˋ��[ �{��/��.N��F��H�0��ҳ�;���;tP� �CU���R�l�3�K�j�|��-�>�$�ӷ�q�	i����!��W��?�j�%��u�I~6��d��L���v��
ܫ��a4~�Hcx84�m�S��"	-/�f#��U��{���
�#�n^��Xe���B$ xh�ѫş8���͒�$Z�%���Հ��g[7�f��a��c/�N��_2�����\�Ӹ���89M�'�*��!Ԩ�����2kZH����K��J�H��/t�m>49Ԅ��r�_%�˴�|%ÿyO��
���2 1BPI�#�����IY3se��h�Y��`���]����ڹ���������r?v��}�?���y��ǯ�-�R�qdb�c�l`��D��I��wɺ�cOR#�P�z�nj���lJ�޿1	�9NȦO��X�'QZ��JT��@�X˜q��c�μ5��1I�"c�gn�G*p�K
�kNM�l������@�%��ޠ�,s@I\[4k�ׇ��k�-BMpa w2m�(փ)7���~�mn8fA���ެ����|ܜ�HW�F�_9�x2��;��$�y��T9TUTpc���ț.k_ôĆ��� oJ
�,), ���Kw�ʷ�ހ0i��!<�]��5t��}�4#�3�'�(W�y�	c���lT��l�R�el���Ko��iHM���)��S]���&���!��m���v����"x���:����S�}yj{[��8*���Ve+hr�U�'�0({Q��$��4���U�N�z�ƅ�Pd�u�.�j�R����ǶN^g>�0m��D�v��tf+�9􋖗�w}s��f��P!�7�t����v.Uph�&[f�w�$�Blq����ߞ�m<&��t���i=�T�8�m��pC`eU��p�O��tP��!*�{� J�z(�\�%��4N�U���h_�@芝�;�U�v�جOó�d�����9W�TpB;>�"���=d��0����wdx���ȥ��I�O�H��COoת�Y�f9��l�^l^Fa��I�f����3`����n#�{�/� ^*<B����н-̀Y>�A��[z�i�c%���	L�����˿�p��2�����c�{�z.$]ft�*(^��=8.�e���r/�G��^�Itn%i��e�E�K?�2���4�7��셮�f�Uy���@�S8���'�|�[�$
{��І/c.2s�ڮ��bku�*+ ��A�;Kj�9����p.3���X�2h�b��4}
{C�%k�meq��l�.��f�$H�������{�mEq���Omr����l�:���`�iV�H�:�ͱ�j���D���>d���v/^�W�
i;	���䖒�?@�C٫-��f���8�V���ݍ*�=��c΄� h�~[`��j�s�B4o9U���`��>x�N#�<&�Cv���;�QH���Rb?�(Z34Zk�+Kn��ö(�֨�6��r�&V��02e���0��j�q+3��K����Wc��W�mC��/qi�g3y���V��HO����ż�Z/t���+�w�&o.~����`kٳ������dW<:�C�!��f���{'��x�j5VG���c��B���I��i�9��m~d�E�ҨН��It�jP�a�	TsN�O�Aۻ�\&9���,K6�G;=p�zi�N�l�"�̚hpg�2��H�I�>��ؽ~1���F�B)��l�0��~	�[�2�sBފS$�SP�(!L%����?T�>j�<��, -u�-��YxF�K�N"�'v{�V𴼋��qW���pk�8���`�<��-T�є�>ܶ(�3�߲�n���y_У��A�p�7弳�;�؁5sr4��
H��ٔm�E	WB�5'J�!6�B6�4��8+37u[��d��_�qtt@��~���.	����!k`�U�>�����F�Z� �#�}`_�5,!1kz�\��g�sq�K� Q�u��%ǜ�d������T�ͭ� W�F� �����Ay͟b@�ɹm��@7���+h���������Y?ɪ�1(]�ʊ�f��ܖ�ˣ"i�[���;O�Ǽ��aL["Tj|Ԣ�WZ�|
���Kz�v(|�.�Zz/�i���-:���yP�\��༻;�:�����OE�e���8���&�*�<Ʉ�,fmž>A��d7Jc2\Fz���#t  �0A	�K���=�BY��R\� `��l��A��n�K5�ǲ����5?h��s,l�r��`ng<9��آ��˜����@)�o�'�BIVLqMV)���R�i�\�[�G<y��HD����1n����@��ڣm4 �� �5�l�g��A"fK��o0Z�G\�B%�;5I�0"R�ai%���$O�6��8��SR/a�V�Â��R.)N���+`9"��ͥɌ�Q�S���$�6Ky���Zy+R�uM�p���ٌ�����8��Y8oLc)�ZLk�1�l����MxR�+��&P�#�){����*�j�4-�oKҭY��_��6���ϡ�.���K�d��7}c$�>+���N>�d_;�WG�9�99I4W(��-�=6a�%��sۀz�%��P�(X��Q9f����Ͱ��5#u�0��o���ʒ�������L�p+�N�{�~��o?�_"�^z��f�S����\�(;ZP���a�:j.�CՆc��}�W�s|���w�Ƕ*QZ�k�ymhJt������aX)*��S�Ib���7z₽
�W�r�θ��1j�r8�Mѩ@r��CШ^^w��H-\�Tu�h=�R��]ܯ�eO��D�;9��,eV�+-�xر1"fuo$g�v~Q7�y��iX��Qɑ@�Ӛ�m;_}�����Θ��-4��:)*%�<�D+�WD�@����&ԯV�D]d�n�N�_=�b�U�7>��ح�{�ꋙ)nY��$R�WP�Vb����ߔ}ҩ�K@S�i�I2���sR�Q4�ԼK��so��6�8z�`�1��Mp�_��R�א�Ìs���g�"v���g��V5w\�*��FmE��.r24�UIH�i��f9}�����;�;k5���f����ƃ�;�R�2m��F��q�V��9��!�l��%wc\��%�n1���#7״�y�xT�{���@_|0x�<�x��*}�1_@���qb�͈蒹��}�C��LX!�Y��HJdw����@K��Y��G�s�U�U<���b�lT�V�GÕE����R�A~-cG�����I>T��);�/�A�4;��]=�� ��T�����~8�^�Ak-ay~
��	�Af;�(�o�8?�>�e0�w;Z���
~Z���:��|���by4ټh[O=�Wo�Ɨ��^�A'$"7;*�C�w���}/���� �ռo#�N��AD���>��A��w���g?ܗ-��QgW�{�րw��+�V��s�*$mjV�҈a�E�#�r�1F��+c0d���
+�z�|0��:��BR��Q�6aԅ֮;7��U��m�G���T��:���K|�!�?��&��X5K�������µV�ݠ�u��V⋺G��S	�*�&N����&\����m0RC�$�"۔�u�ƻ�����_��V�|<Z��W|���0X_�rfz��i�7��PҔ.:�)m�������<����Ѣ�Ô��@�I��!�@�<���m�����)��F߾zr�x�A�z�귕;�����L��ٖY���^�:`/�pd�����
u2B��D������u�#"Q2L��I��OA�C�}[P���s0�q c�,�@��p]Ջ��o�4J}o�]
[��}ӣ��Fȃ�!���w�n;�������pM�����#��ah��K_m-�?[��d����:�?���]7��Pn��������kZNm�g���W{�s�8�.�Ɲ����]�D���7 �u���U�PM6�%Q��=�2dxߕ�{)!D�z�~3$�(�|.�IC�06�_�UF:by��Z+���?ī$�Z��x�jh�ؖ�����8��<��qh�GV:ݯ�GG�֋֓�?���s���L�-����Lb5�6M7OE%	U��(���w {�F~�.�ǵA�$��t����%�<<���ѢeUޏl� א���N�����n/~�4���C�4g��<�o�;�);��kM��w㢰���e:gK!b9��Vǈp q��cQ�J�9}�?W<��W��b��-�̎�q;a�%/xm��uq]����1�t��9_�`. ��D��� �8��E9pF���S�a~�/��Ѝרށ�B��C�m5-74eZ��I��?s嬗J=`ky��D���U)���>[�p,I���!���߂�0��}3�7d �V�j='�V蟛�L �޺��ѓ�OX��\�tni�WK�8�ɑ�@����|�,�Y&��s�c�*<�u٬���2E�kW.�WQ�b�/�ʖ��(3��rD����ŀ+d�Lx��%&����o��B?���T�S�u���{L�i���̮�M�@K�$S���@���@�����*��}ʺ�bx�{4�|4�-m�^=̻<�f!5�C@[���d�8���m��/�k��H����?=��|n"c�qCI��fBq���i�lK����s�a�Z!�7�cq&GhR�Ә��F��{�ռ�gT8&�Q�|�Md����Wq�)��ge��ܬB�P�����8;j��)~��>A� kj����#��eK�!W�&��2�졜v��R�D�hx�؅�{`
��P;-�Q�x�d�o3�`+K��i }���~���J��������u��:��a1*�9_)��8���؄�m�T�8����пZ��Nv��T(bTŭ_]���v1#݋	��x���+�a��'�=5���ѾSe`�v�Jf{5��#��m��ǋ�9�ue�EN�s[���w/A
D�%_��r�����3�������&!(���a$))� <Z\������9j�ܩp٦q
_��Y�fx���"��9h�b��_Q��ޔ�9T/�igjj�!�s�z)X�.�ok+��`݆z+��E����3U!c�r2������.���B�uk&T< ��[��ZS^p���]m/(_N��-ӿV���#����P�����QA� 2 $q�yK���q����R�$*�%>��l�|]廋'�^��H.!��[;�}c���
\���dVK�ae�k�{��U8�-���C�<^�})��ˎ;p_>��Ǉ�3��#���j���+D#�U/m���T��Bf���S0�y�Qj��w�ZSuoش���~�/8i75�(+'�2(�Ы�D�7R�C��"9�� ���U���U��-�l�e��rȎ8���vX����Ŝ�'��$b $ /Q=.�����X����pOg�>�K1lbC�XG���*��
�X!��X��rž���������$,:A�-)l|��3�@ui|d��_.Q�$=���;S���y����$ە�Z�d̑�����SbXr7�j?ϸ@��0���ӬV#�v���F(ܤ�Z~��Q�P�}�&_<���1\$��'Nʢ�����%f� ȦUv��X��@r���LTg.	�ja\���I^�"�TmOS�F.��o��� j���)S��.���T�^S��cF��n���EsA�Ũ�OQ�	ڊd"ިzt�»(�D �і#�<2&qt��!� ә�U�m%T�}�k�P�Z�L���0���Ii��B~J� �*b2���G�������R�?��ܷ->w*S�������0{��d �L�a��0��S�ug�ħc�v*	���{���� &!і��~_�NJ�ȡf(ur����FqȕZ��  �(QoJ	�(�d�ƥ�!����/Ȳ1D@�ZpV}��Q-5��\>�:�w"c��ɋ�t��Џ�ﲑ.�����Jb�G����_.�;�%��Cc����5�����)����tǷ
�'�%+�+��ל�}�+�^��u�0�,���NZvu�Rzp]���H<+��[��լ�S@kJ��	c�x��;�\�0qVs��D0���~���������W$oc��ܼE�mpʭ=���z��o	,���o�����׍�v��2�Y����g.9��k��(�mv�F����� }��E�۞�]qH�/���y�*˴6���~�}�>�:�W���)I� �������T|�`�)��	��B̃��,���VZܼ���@G|*����aiVo�[�(�pL����.�Of>�{�:��`�c�A��sB�����S�TF4A!k��6#�H$#)��Gb�����.�ߤ���#�Q���uI�0�~/�7R��AHs]�v0�����u%����DnQ̬��`X�u �K�u,�^Vz�A0ԼdCl����>��kX�o���Ɖܤ��Oi(���K��6��4j�ٹ��F�o��Ms��:H~��wt����4� �P�[�س*U���%I~���Jy@��~'��B�0'|���K��mf{��s�>���ΜS�
���	�*P-=P�)B�0P�2��N*w�	a5(�ɿ^2'�DTl���EU�%��zC�@*�,����Ŀ��|��t-Xh�^���õ��9�$�&�ep��?�݈�ϧac��T���1[;�
���%H�5L��)[�f�g��.K�nk���麗�i�y�A��/U���������ěy��e��|��L��$�������0��l��]X�ƭ|���S��%f����6��'5�N'B�QK��J����䇫���QH�A&-�?g�k�E"�&�_<Z��q��M3��m�=��$�����JfR����+��7H,̄��,�
j�z<drc��|���2߷Y�-�0�v;�0ᯆ~:2�b�fUE����h��h��I�JA�x9��0�%/;��`4��Nj���g��;fvw������_Ɖg���>��`�_�n	R�ϥ�x�RWxW����C�����tч\�͈{�UD�#���8���e�g-������x])���r�7�Go+���Ȟ<l!��0Hl�����B��o�k)Xf kzVo��c�������r���nx�?�m�S�64�Sc����������d�a��<�6<Ch9�:�����\��o�W0dl�G�J7�u��8�` �h�L�~A�N؜�~���P=�6��|9%�5Vw��Kj�N����b�֢�=�	U笩]�y}E��*��X��x�[HbK��[�����O��
ެ�'�2j"(K��&l�]G���f�Ӣ7�ޚR;K���B\m^�!�!�g�#�
c@&�TK��ܖc0�n�)1B˓��\�sWq�[�@�	U�Hy����DAH�6#�ba�3ۘ����5�}/�Ff��D��Q��벬B��F��;B+$�E���T����� nF��=��k�6���c��m�OB�XpL����������t��r���Fz�>�4�k`�R�)�����l�kU�kk�' Z�o�L��4� ��)�����y�u���h�sZ	{�!�1��	��F�0��5H:��FZ�upu�TB�6�W6�!T����}�KGsʴ�D+b�`���D�F6*3���G1�5LD�}�*���}�� ���	_�����T����Z��G��E�o^
�JzS~�*Nj@*��$��2�'y�����$sJ4�+�	FM�M:���;6�[�e_�b6ﯾ�I��L�V'�q;�D�xI�؄���'����mY�1�&��S�V���K�y��U�ANɦ�Y�����*��_�+�s:���f����->�~��J��M�K�׳^џ�. a��ڷ�>/`8��a:�R����[@l�h�gI��])�\[~�o�D�;�����8y;���;��X������@�r����L�X��a��7������=H�ˍ��?�[B�7f������9���,!z���%&��*#�[����	�.��SCI��d�φӰL2r�I���b�x�j�g�1D�c%ɂ�!�u��gB��֐+�a����T!��N����J��i���2��;��E�s�+݅����&E�Lt/�2�´:�Ǉ	�e�����D_#\ ������L�)�Ѧ��,Q^�<�ڙ�|�%���1v���BN����������Gչp`-C��p��^��\���������ܡ�/�Qꪕ]O|��`D"�����^*�_u^U��7[�8`���M�f�3l�%o=X�d��F�]7:S�j87G((��|LzX��R�0��8�OӲ�x'��1^�JD�hOL����}�2l�Nq�t����蜎f|�2�M����"&eYF��N�����0.V�=��%�B��g� p��䞱0H�'y��=bj��?��!��t~���ɰ����w[o�OV|�����h �&��C�_����1B���Mz~����r߫s�SP�47Ak7�tn�d��C#r�#Ї������Q���,�G�`�S�}0�Пʪ�WK�|:X)�>2U{�eN�>�8�bڼ0�<\�S�*���r�ƦP��4��	���g5	��Q6����7�!lm|$�έ`�,���B#m�a���	_o�w'1Y��,EqY(mn���(F��ytTd�
j0�ɉ5�����>����4�?@��&Lb�w8�/���s��\���V�7�D܇r����p9����i4=B)صR�T��sX���=��^id�s�U��w:
s6�+Gd�WN����.b�7)��jf�T\��~hI)ѫ� ��TG���&<P��|�t�ږ�0���w�^G�������PNz�Wg��Is^JQX�ę�Fq3�'D�@o �_����X���h<)��h� l�&QF�E����"�w���˓��|�J-�x�	ENcD&3��*����0"һ����&L7!����@�Cvr�����MѲ��9Ɠ��?�_|�M�V/�jI����І��4Z��X����sܐ�4�������e�l欦S��<� ��]@w�P�ͳ��t��V;�J8{Y��� ��XG#P�˻q��οW�b�2�w�����_�i%�}���$�\^`
~5������� �^M9m�KVci�k�o7,)`�|KU5xd5/��֮M9�x~2���[��N��fV�9U=�Z,yz�F� `�S:<�ǐ��<h�8*\Z7�\��{%�mZVVnH�����~����3�� ,|z����M��Uz����O'�E�f�-����1�,z���F���|Sv��	���5O���9��Q��ڸ&���׳f�5��)M�<3^��(�5�Dw����C�A��&�n�]z�6��_����D i�%S�{�m��}��Zc�-eT$Z\iN��ò�ш������!tI�m	�;�F�����L��uF?�G<$Y�ڒ&_���M��j��$��̀`�j����
O����[f>�O'�۳'K,<���Eo��-[4fv����=�[�[�D*;6����R�Y/�������i1[��sj��̭�7����洬F�� L����6
i`�a� Ĺ,9^���n�[I�T�b|t�����H�[F/��Yᇳ�	�~ �>:8�7��6�d��]U���5�
̬<����,�٭���@W�+��~3t��w��tN(�@Ӷ%�`���Uw��� ��<��j���4*�qc��������Ak{�ѕ.��]3�HL���)�:�C�N��/J���ƹ�ˌ��w�p?��#��̩S�.!���������Ǽ��>8)S�Tv������N�Mh�m���b�5u�ᭋ�g�t��GH��o����p�2����X���/ҫ`Ƹ���<�"NH�x|*��m�Uo*����@}�l�+����7���46AO:]�0 dפ�L�O�v�ȰXk�5~iF��-W�:j��!������JF،�+��S����`�"�|1?}��Q�����3���[D�g�}�l��:Ji�z�ǆ�f�����-�i������悉Z�N���z�V-�pf��D#o�eU@W�LM���q�̹��XK����Y��X��l�/���e��'�K�B%�IT��7��� �����	�v��rH���� �L"d�:QcDw�^�q�SF�0�� �(zzW���,��i4��.÷�~�jP��f�9�,�ߊt�V��:ٴ�ڏ9�˰p����%uve�R����|RU�F��*�r6�V�6FW�5�� =�/>�� Sl9�O�P����r��w#��6���w�7ن�6�K����!��$gzHn�Ag��V�Bb��o�������#��Z�[t>�vAW�G��gνL	G��M2�Hs'S�>YR�):_xZ��_K��a�w*Z�S�Ya�f�6g��c`ׅ�O~r�k(�2 /4����\��0k�X�ӓ��Ur/���F���GЇ�û�z9Z�t����X]��5�^[�t��	㍎ڞ{l@A��GQ��hD�#�}��|� X�
^ƿ�V�Yk"�Nz�II��M�j�����؀#�xl߮p-SKe�4��P��e/�o���T�����-h�,����(����[*(l��7��W�|,Hx#�ho��#G>=�ؤ�y�W�x(���يj���s�	ˢ�{r� �[5��4�'w\|U8u�.��Ӻ�wo�RU�a�pH؎��l��LK�����p�I�w�[WBl�:�v˞Ʒ�MV�|B�# �;V��f�.�;UzhdF��6']B��>9�P�q{��F!5���W��G��T�=�vm���6�)�pSp&��:��={�Z8�]xg���t�NԿ`�F}�{�_���pZ�Z
�zŘ���jl�ڻciБ�cZ���,R�F��������h���m'�i�K	9� s�P*�}ܜC�~?������`)6w�aUK��>��������8`	���Oq����)h�8Y��H��@��د5��]�(���.e�/��\�Z�r��)GԺg#@�},®_π�/wi߀d�O�O��8���|'�j{0�J��|��x��n���2���-�"lj��a�&��K��x�
:�lѱ�|�
�r=Q��U�����2y{��8�+YjD6�)"�nle\�u+k܅<�j�/��4CL�T��^A�F��S�:	�Pt��3SK�Vu�q,�s��s����..xMe��ۘ��i���I�Ő�
|U�����ub��NQ������N�	s���=��]�߶��tnh��
r0?���{ K�NB��]NA�):m��rj'*e�i�1�� g���Y�� ����+�;&�帝te�n8�@�.N�Ƭ^�-̅=z���������J3!;xE��
4{Ôѩ��;8.T����yE���=Y���U3���O�sq�!z�1��B_�c�É/��9��n�ݹ��Z�U��83�U�ܻ�F�&uq�7�$Xlk�2r�.Ja͊}�%x��l$��#cu����+6י$���=�W����#,~��øg�(�'ڰY���Z�z�:��1]ɣT���3��Iή!��i)�w�Y�u2�M�Re��`f ޱ��$����㊴v_l�9�v��4[A�-��9���:��܄b�j�o�p\ǆ��4BnDq�-�**\��֖B��U�N@E����*������rHu;p��p��Ӳ�{rWo�|+���?�	�%���X�Zj�~���T�� �Tx�(t�׻n��H�$�´Pv�Y�T5G園[I�0��9
`�
������)��A��fj.�6L��:O����WR�1)ِ^��J ��$�<����:���x�y�_��u��"�󚛑��*U�T��"�?�5�g�ܰ1���H�k4@���2����J�a���(5�@�xj�*)^:�Hl�:r[�o�n���3[H5�S��z�n�݂ZYx�C�g��V�:��b( �j6�T/hPt�<إ��Q�B ^#�Ⱶ�}���K����|Bپ(B@�j��P��ј/�����)z����v����1Z�<�g3��7���f��k���%�f>���ž��E���(�FW`i��N��o�6��e#ܥ�A�Bk�?Ԓ*�5F�L����nꄧ����?Ha�v7-UGT�.���gbb���'��z�d��;�a��h��+��3c�1�������tp��X��ޞ�M��Gg��fu�b�FTky�����y�w�ۿ1/֫S��Q*��㓖}[9Qrۘ�ZP�/#"���0��3$ͪ����
ʭ����i.4f�Z����k�N�3W~�/�s�<��-���g&�i��9
��k��w���w��`E�j��D=U9�$�R���X��F	�>�~~'+�&��-�S��nWA�f��|�׶�C���*�|ql��9����:�B5�|:����x]8S�%p�DW��g���(�Ǉ����\%!�u�ײf:D�5S��*�^?򔚊��=�qǣ^5R�=T�A7��Ƶ̲�� �����JSq��Acکie��Ws$�
�����a"@]�Y�69��q^���A4-�
)A��Q����G4�[��R?77��m��+�t���k7�y��8����:OQ^�����>ն�o��>2/�52e��#�9@��F��Oq^�[{<v��}�����dgϡ�2�$���>.K(,�הcHn0�a$����Wk�dL�w�(i�N��a��<9o����,~σ�����MŢ�>�2V���p�X���mV�(r���7LG�k'��y�m)X��`�ٿ��)	��&�M���u���i~�z���ӓ�1�~��.)R�ŀ� �rL/��W�ZWg�y{�SlI�wT�(z�w&)ܴ�1�4&b:�N�;JDq����,%� n?��ٝ��Fǯ֛��.1Z� yb"^"����b�o/�6r�����Ke���dW����4�����w���9/r�8gɹa�nξ:�l��,)�'���<�	�K�Z�I���4�5�_hWi��P21si(B~F��U�f�9<默=��O�P��QΗ�;=qo�)��f=t��6~�ڠfTx���Z�)A){�ic�źo��BF�]Z�+��I��Mv���y�\�9�`{`v�ݖ�̅�X�8���H�����a;^']]/v����Ql}�z�-���8/�W퀓�=���В9�O[B ����`v���|mv������Γ�Ct�]G���8�H��j��S�`�La����8��oCF����-c��.�֞
�#����P��ވ��?���珱�\݅�?Cz��f�z�$�9�_�4s��oS>6����j�n�xU�U`�����j��Q�kiS�r�c��~kN�]�+��zx������6ß4�>��z�U��g���/sM�fO�o���K�ֱ��I�B�\`�UÙS���s�u�a��C��o��>e�js�1�-=��b�Z����x�
hVz�?�t]z��t�*�G��Kw�#�9f�W�U|�܏�փ�5�)_�y.�I����=��Fħ�&�6}���HCE�C�Z`��,N�~��P�3O��y˦��RY��t3�;B'�֌�]o �tX8XO��xE/����?�+e~C	w�����7�#����� t��yi3,0�9|���"a���gq�B����%�zR���T���}�qE�GE@91u8^Z=Rv<k�)n�ѡ�+I�z��R�|�Њϵ�iK;��D�e*��u�O�2M+F� M��]8,�%��e/T�e���"��k!����E�~;R9������o��e�Q��X� qO(b�zػ!G�y!-�O�`4I}K휌�p9�Va�bK����d"��$�]|�A�"�T0ív��;�h�NY�w��_"M�H�ZǪ`Mh��My X�1�O�^���\�J�`�Rk���kb�����/���^{#��4s��n�uٓSP��C��Z��ھ������/B��y� ϊ�J�,���^]t}uE��(R�����N��ʦa��X�_3՗'��L��3��
x�Jv�&��ӥ;8�[�Œ�;-�����J�*E����[��)y���A�.����C�s'G?�T�\�v�6�/�j��x�V 1�e�6͆�=�΋�+��x] � ���|n���ء�����TI������������b
;�F[lV�{V�,�ꘟzV�Q�+�9�F�#��R0~
mQ�wT-F�K����oO�T'z�W.��T��)?����U�\�Q�2_stH't��Ɔ�?�س���|���մp�PTi:�|1f|�����e> �%�+�l�A���U���vU�)Lp��w,>�
�"T=Y�� �2w����P�t]V���`�j�ν|s��=,}�G��갼�跡/��x�a�-TUnz
:m�@�v���ԋ�9�{`s�C�Pճ�ޢ���M��5<a��6NO��a�G�:����)��r�C�ɕE��Y_ �io�y8���)Lve�8�#$���n�r�I�f�Ns<������!�Zi��0aX�l39Y�').�إ@aw�6�U�6j��t�/�bj6�	�x��:��A�������Z��`Y�«3�4O3���mDFU��b\e��NpT����R->���C�D��ĮF��ݳ��V[�D���r�oQ�DV��:‿�w0՛�}�����}#L^�4��*��U'���T�@�Һ?�d}И�T�w��k;��;����s��Ϭ|M4���zLt�r�PV�@ˉ����]�SE�R'K=�Ш�VDD�����	��S�vS�/�z�D,w�}R����C'����ڞ�-SU�kS�̒ق�֕ò~g!�d݆��bXʉMB����:��L�/�*�Yg�`��2��F���V6a#)��e���I?=h��M���`��g�M�B����]��Yu�l�d8.y�����!C���|�5Y�!!����H~W�|4+�Yq\��{n81}J��U1��"�SX#��Ь?�KJRHQ�^��|o1�)%��Ȓ@�c�H��C<S]��i�ȢL�_}k�����t��֫�ov\��_�+��#/G��|�p�P�\~5�q�G�[�<Gʙy� h=��C�4��ľ >ٺ�<5&@h&3H�/��j�a<��}B�02r�_:s��5�����Mc�5���8g6p��ZMm����4��m�V�Ί���^��
�%�G���/iW�70�Ba���@�b�o�+��!�D�n��I}6/�l���~��)2a@��FNG&�L4�/����W���{i��}Ѧ@�x�}]�da���S��&澹�z
��,����a�R{,t�U�b������BR�?ϸ���KW΍�guX։��a�W�����H��s`!�L�YKmZ4h���ۙ�ӭTΓ�ߑ�W�sOP��~P1U�}J��X��~�0�cj'�ȾR��©�xȂπ}�ׁܥS�W1#Eg��i�"��ɦ6k�������Ԕ,n�����`6�!a|����m���>����p�s�L�l?�a)�4��B,Y֚
M��6ҽ�^�}�2u�vy�Z�W8��6!�F��u.�t��:Rj��-��4�1�vi(黸�\ݑ���ߥBD~�Sª��U���	Ǫ�Љ�.���N��:�1�jWi'���\��u*�}гM�G��]*GJQV����΋68o�����7��婏��.�Bp7L_�菝e�
���?�Jt�,�'����m��/YK���Tj&������We��28�"��t�0'��@�s���**�>������<��o�����%� n񯨼@�����k
2����n!O���l�-�t�-Í(@\�����u��8V�k<t����%1q����3��a߭�e�F��J (��X�֫}��xM1�H�;ð/M�H=q��+|2�?E�eq���΅O�I	A�Q&� ����tg�mCi�1�E�D)�z*L�F߬��yi�k��H��V�+n�{����V8+�
|*����F�d��t�U�tE�"t�Nן�)�U�x�>�Y]��!�s��ݭ�v(���i�LS���h^�<m���u��n�3�cl��/G3yc����Ƀ#F8��k˔�R��?|SD�����Pgi��뇩I��V=��b/��n�Ĉ�3B��շ�|RJK��9O}�h�rI�/Z���HmEy��,~�ͪ�q2��W�[d7Oc�Iu�S��U��
����J�Άg�ȺP(~;��[��*#����/?;��Z?q�x�p�����y$]rZ��o��a݁�{�aa��)���D)4N8�K���5���M�z6 sV�NN��E@Q���b�b��,/f��U9S�Q�&�47�Jq�˧�mW��_�Z�����l/J�V����%��yr.��KE����0?1E+���8�iY�[�*�Yya`!��}��g���}qy�MshtE�}C{�>:P��RA���A�p�ۨx.H�Il}�:v�RY0Ё��kw��.fO�v&7e���	���}�I0�}̈*���ޮY����]�kD��N���H��Gy�%b���遟w"x�l�^i ?�гL���9�v�##�����J<J�2g��D��Y�e��ľ�Z���y���~�R��'6��+�D�TQ��tK�Y�X�̛X�&L�rU�Y��D��X�Gr�+��3|����i�q�w�GkOn^s����ĺ�T��i#��\v��t�a����`D��Z��4��OF�XѠuq�[� !��B�{����e8��-�jg�-�`#�A�q�nc�Q��/ʰ�|�p���|�׶��'�Nl���[:$�� �FPO���N�K���?*~~�Z��Ur���Z)aߠx�-a�pOGʹ�`#��ԎD�9c��T�!=�~f=T���Ba�ĀB�R.�d��%�)"�d +�ڮdʂO�<�8�O���k��>2�*dq�o�ׯ�H<:pi�rq?C�/o������q{�D,�Ҩ�t�n&0�F�V�C��]|�E_��mH,�=P�[��\������ܮ������D�ϊq�E�ѩ��}y�"w@+��Fp� ��ú�ѯ~(���00����?�u��;o�|)�K�F��(���'�M�XU�C���~�;������lL��3�m^�k1�&�v����y.w��L���y��4�e�lU��,��Y2q_�SOr"���&Bt��� �O؟W���ʍΥ�^�R��nT��8~�S�.�(�5�_�5�#��44�G��N�FNؠ����xCU`v�z��:��b]��q�D��B��lk�K�#*�k#S��A��0���Y?4�vV�fM��m���ȱ�.Y0j؉�^���Ӡ�T<������N)ԇ99S�<��n�Yq��0�V�d�Px�q�O����U��>e����I%��j���������OH('�ɠ�nX�l#������6)^�	�p�<��r��5ф��X]w�#�ۄ�i*�\���͇lC����������d�p���`����69R�;J�D7&�G�}�%.�ߝ�FGԓ�,:��ۆn�JDR+v����/\ߔa��*w�C�� �
��ڜ-�gV��H?��|Z�Xy��R<f5�(`L�&q&D��&�L��F(�j��yɓȡ%Dը�o.U�sd�Iť�ǳ9��A���mNoy2P��h'Uv�����������'�����,�� E��4$;ܡ�k�w�8g^�]%r920m�_<��<;K�������υ�����1!���P���Ы�x���fm��w��ؽ�2(*/�h}�%1r�MĹ3X�G"�c��I�B��B�F ����6���}�sz�@��Mx�QH!�-bIҒ�%nl#�k�`̃�Uy<�P��np��J���e:�6Aw����PT�Z��=!|�~��(~�nC=+)D��涄h�[�<�K�#O���z������f�J�}�� �P�|)d�,�}��N�� �q�w��KDx�ygt����	�r����J0���az}��|[���]H�r����	7�ٔ0����9�wA�+�Ub0"��f,Γ�j���մ3m�L\����N���cS�{��뷐�"߷B6��ؗ����(ߟ���T>#��?JTw-��B�'[ᧃ�B�h�,M����E��Y��%�{^?tpX��/&���[�#=er�JЏ<�4B�8�����E6����[.){���Kk0
`�K"V{�B�\)Ez!�`��]�Bp8_�)P���#���P�P'G(w�x"eƺ����m�`�����360�G6��ٵw�Du���p���<�^~�"��	�w/�KSm���?}�/���O3���� ,s�D΄!�%��sǵ�Ǆ�����1)�g^�(��I��ñ���\�Ǽ!JE�s>iq ����#
!�~,yT����'�\d��5����S�lX���z��,+}]�7
C' �[k<a��]��;�N���� �C�)�)R��P=��zr+UVۀ����H�w+$U����_"}����N�n�]Inf���T��?<R���&�25>`��p��	�-���W@�j`��/�Fع/3P���4�7@z�����<�5F�,o�x�-��>�+�'�u�������k6$LZ3��G��� �E��=?���;bv��3������4l�UvcA�^(8�w̒?vpJ�d�UB7c0�BO�LB"k��1�#E�Z��d7B�{�!�H.��
��@:~k�e���;���W�LT��>a��M�G��/��p��\~8k�A�9F�Ý)g50=P� ]��_��_e�������u%r��*z`�=0��_�zT�y4�pV ���ߔuר3�=XC����%�"�C/[�o)%�ꑡؘ�M/��N�5�T]f5��HƢ�);�B��x���/��*|�|Cnۡw�`q��\�lQ��C�?�#�:�EBz�4<�Q���m�V3��(�1�S�w����'�_� �NXX6���
2�6>�k������`R���@�["��;V(]��I�L;�
���Y�����U�R4��}��iOϻ�'RL]ԡ�nAm��i:��7���O�Ѩa���%܀�C�{%OZ�fK�oG���h6�Ĺ�{�24��Y��׃�9!��+�[H�vLrO����?5�t9��B��U�`b0���&;�=��,>@Y]�l�;�D[ ��M�6���ۇ�;�v�r��+�J5�ME�" ��t7xgMa9�N��'�j�De6�m���?�3jO���?���Њyc�a��9/@e� ���-��#�τd�p1�/�?�{=�	�M�%���K�H�*)��7���F�7֠�W�ᕌ�[�h (�5�V��6t}۬�h�-n��|u�Nwh��g�w���M��$�#5� n�
L��Jr �'~���x=����7��
����{�|dL��s��  ��b���e��Y*8c�U���MC�cG����>~(r~CM�y�p'�L��ڣˤ��Xۍ����U���f1�s��S��S�D��S����[՘ӝ��|پ̈́@f���{Sa��:"�bOx�7
8Hk��^NG����X*/�PT������11�'@����>7�U��c}1nԫ�7G���(�1��z�d�����Jn'���?5���O�<�b���d�I��YBɬ���ā�±�)�#z�:�aI��I��:�n��{%؏{F�S��]$S�Ȼ�Ƞԅ%��'Ar���9'}��J��F�/d]%K���7��d2�iF]�q��e�1#�8��b��D�g� ��0N�V[�Ǌ�PnmD�4�8Le�e��z���c�8h�j�cv��uFT�'A�?9T�R1&'�������u��ޜ����2�B��;YAn�`����O�
��Q8I���>�: �4�\r���xM���e� {K_�|xv�]�~J��ь�@$��f�+�� {r��W16_�*�眑9)�AU`"Iu�* F��)x��ӗ<ucIF��ɹ@����l@E�p���U�_[��*��~�&�����S��8*9
B����ʧ�D_�Ry�n8>�-��1��������HVX%�$�f)[)�L��k��ɑRw({WA_F5`�r��s:E'�B	��$"Q�7�Y�iG�#�5E�YjUU�*�9$�>G�
��l�I4��ݸ8|nJ����Z���3O�:����H��$��4z�@.
,3�����<���a �Yo-j��9J�sM-f�/��r�b`�)�{�z��T4o��3��Hl��x��GLC� S�;���:��w�ҍ���GJ���H׼E��tn�ѾSE����ǟG�W�oHTk�Ҏ�����]�`���0#�پ3�;���8X�WЖʥ�{o�K:΋v���X`9���뗸J�!1�Z�*N��ᄹdդ�(�*��[����d�I't��x'�=���R0��(��s����sf�Qz�s�%�}�����Zp@�[dk �ipJg��ξu����Y��]���2q)�w�|D ��p���߽�9�=m��I^�=��$��;�\x������� !HN謾��Iܩn���C�xp������oI�:��q+n��z�C��BO�+r�ҧl��E�A҅�t���]���_i$~�2�9E�(t�,,mo�1�Y�S�g��L�+��P8�HkIw#Iϰ_P��m�bq��A����t�k����} �G���	0�[8��d<�Y�4(r�$es�~ӹ?�C1{����]~�"�8W� ����Ck�jl%�-ۃd�[#$;��;6��ӳNMabvw_x�/�Ҁ�Z�+��T��@��I�F/��R�Re 	!z�'���~R"�z�s��(�t]������`�-�]~����Wj�ޥS�
j�}���V�͉5�GD����ܻ���]�d��$9�g��W�FP���}�Pi�7�"�!��a�[��k\]P�O�tzI�T���ٓa�����}������Z�3;�>��(���KD�^��6rTЍKT�0�U�nh�Î�-���@���fS.Lw���@��� ��U,�%e�@���	�Th�Ђ��)xi�y6�?�K�$1�/��^ѕ ��qVd����H�㹤@��\if��G�����������

\v����$G����"�Q]n)h]a�ۦtp�7�^�%Pڶ�(D��1g<+
i��cxr�a��e�|����9wg��g	[�n���+]��h�^����������<�i���_�Sk0]���`M�~�/����\<XR�F������˵��}&�*�b´
	�m��D�J1��� p��C��v,�%S�E���e��$�<��
�V4_�B��1����i@�ԗ�)�<o�F�^A���`J���K��=�e�(�|�*&K�׼��I�#���.�+��(��c����a��zDy�<��0ӥ��y��X9���[�D�,���G���I�=����83��<��g�t�	 ��zZ5(/S*���K������>���:���k��p�ְo��W�8�E���\�谥�k�]!�w�}��(����GI �ϛH+�b�朎�H�W��{]"�g�\:G��m~ܭKa�*���/���깶�.�њ��k�d���`�\�Fy9g`~![�"R�ˌ���1K,��M�T�P�K��~[CƤ؈Gvnq�H��䢯z�Q�����((SC�'����y|����{Y0�b��z��O����xE��� �[����/\�)��Bgq(�۠ٞ�o�^�>��E2z����' �@H�5�`|T<Z����ƓN��k�����Q�Ҡȵ�$j=]���)BL4��ۦ�Ƅ���u�4��N��b��qv�E$��	<U��8/'��M�� �᩶)
�2�U
r�D��@C���⩢i�p�wt՘�0��Ϗ�����<r�X�1�kϳ�I�>R79����g��w]���ɀ�<�܁�g_��{�ʚ�o�s�1T�"+�]�{˷'ob���{��-�S�O+D�ܹ�3���3����TN�5Fcս 2��:s���/��^��_INu����-��('��(��������K8�Ǜ�V��u�\�nS�$�M/�A�ہ �\�~'�F�k�+�T��*y?�U�\�~�z�w+@h.�����9��]���ČK�]�pvy����ʔ���VK e&'�dbJBEevQ���HE 7n�p��y�n<Q-�����-���d�IR2<���Q����\f�?����~�B�*�#q;Rrυ.B����~R�*]G�wE�����pKT
@�f�g� ��H�����:B��M8.u¤^��x�M����5�,��/�Q�c)�~:��L��u��	ְF�u����6�a�f�m�Oc���Sed ?�������U�宀Ɩ���$� ��׽�|��u�<.i~|�=Ϫ]k.�Pb��'�0Ϯk�����8���N"�O8$�65����b�����\�5~��;[wk|a�#��ֹ!���e�S/�^�/2��Jtd��[N��[N�Q�ٮ���h�ќ{������n�39��j'�1���C�U1_�3<��O`9,@t�Z�h���JJ�!��۞�?�b���'�z9��A�2��g�9�a
wTo��>\2r�*��B-Q�����c%'J�	�N��|h����y�U���{������:�/���}Ѩ9�_�4�j`�ᣮ���ڕ�o�i Hl6eZ]h8�.A��`鮉Q���x��m�ϧf����G+���6���� �l�uNxk�5f�>3�*U��Q�&���=љ�V(.��X�B�9�"��5���d�%�EI�Mx�p�^jR�,� �s��)&�'s�X'n�� �K2޷�Ϊ��M6l6�"����L��9���^�I"��"&H4m�q�Eb2�An����'ɬԎ�� ��C�����������q��/�m:�p)�:������[	�&h�Y-IWh�7��].�q���8����o_1y��8�S�m��:�+�|ŶA�ɸ�!;�*@��-}�a��:�T|5�
ߺ$|��R 7��\J#����u]}�31ǥ�+��c Ep�8A}�� ��\Fw��g�,�ϐ�2F�٢�NP��	�9BL"S2�{�]]�Mo�t��	G��R>Ͽ��~����p��(��$>�#[�{���\(jl聧t��cW�����Y�tW�7YG���7Dm�{�l�5-�T=�Ʋz�:У`b��誾�5`6�B����-=�>��,l,� 6��<���W���ś��
~T�_��lȒ��q�C�܁����>J�C`H)�uW�X�ݏ�ݣ��������%�b�� �m�x2I�XL�2�>�͕�u�Ɋ��-���\B�v�����z]���)��+���'����Ɗa6ig����X���jf��EN&�w ��8ql���GdR�����S�c��ۆ�Y�X$��q�I/nؖ���K<�r��Mn�˦��<�W챴��@�&��|����e(Ƽ*� ����M�o!���O��4�Ӣ$��l�晳!J��ͼ���F�(y�hro����9�I��G�C��:�+��U�n7�LK���a��LS�y�ٴ��
�r��o�9���w���7�^�hg��է��1��5>�r�<zm:+� �ff��beڔ	��ǫFT_Й��	�����v��X�$Cq��Kn��{K��q����Jg?�%v��-����	�\K���MS�<ku�u)������'���:����� �G ʒ9w�^����A{fw�a%���>t�&�YE�j`(2����U!hzi��~�_��*5q�Hv�I%�<���qɉ�;�Bۗ�N�` Z�uV���nM�ߛǊ���X�]���7���Ǩb�{P��;b�@�dEW�woo���}}Y߆�����B���\���y�58g��WpS�D�FG�����ܓ*���e�� ���[�[f��z��R�#Ba0�;��^%IZ\��
1����dZ�rބ�mU�K�_�*�5>B<u^�� ��l-��� L��]������W� ce�2h�f�p�X@u�A
���$�k﫪�u�\A�Cv!���dBg�ŲP�c�}��ߘ"7�3��u���OyPf�h�G.u���0��T���X��+���G��ڽXY��mn ,��$����w��H��*NR�9p.��2�wި׿ ���ŀ�U�]��MI����w#�4s@�'�N�p�N��Udmag"v�skxS��6���B��VC�^B)�~ɪ��k��z&T���m��;X����\qjVi��!E]��;��9������ ��*���hL ����3���C(7ݘ#HV�i��Ӿ�����%��-:%�R]���>�,�h�+l07�dz[G�M �%�*�͋e��dtR5�Q����&\7�!�@,1��v-�C�!<����;�pF9j�����2 y���p��ȝ��"2v�з>l����/���7H
�U��b>�[Q{��ѓ���T�z�Cט�\��D��<�j0ԇ��2ˡ9�#_E�9܃GͯVM�rr����@��������BџP���ڛ�v=�*�L��qT��ۗ���7�e���/��PH�I�Y&���j�U��ьų��\�u8 *��W�0P�2
�2�@�v�pC:! �WK�O���ڹFŖ�˽�F�U���3���4�A�m���'k�}�C��{>�	y��%�&ՀP���v�-=̳(5@����gy�/KQNSA��������%"�/1�;('��Yr��Az���+�bTsl�J5[m�H�9-ȎJ�Oru+��6�=�'���y�y���*��������t�fk��{�Ĕ͜I;�,��g�1��pM]����������r�����;{���%'W�m7EM��8};~4/�,�89R��=2�\&U�.sLC}\
�[c7To��.?�܀�T��w-�I<֋(s(9�������z3�W�Vn;�Y���Eo�^��;$:,���T&mC�ʟ�XV�o�R����o�_n](�"v�:HM��=Z������9p�������ו���&Iu�RnF&O��g�1|=
R!X?�&6�6Z�S�k���2��i�*���k71�,{��c+�]�'^T�_j{C�D31ߣu��~��[�g���I�?�y�AV�ɎP�F�L����a*b#̫��8'��W�}
�\��x�{�"̂�gY�e�� )�NV��μ���RZȱ����_ͱ�b�C��Pv�������f�L$����ט)V�
^@\�d��-�=�Ih�� �6#c�.Q&|��[�+���-12}��~�%¸>{Wچo�(8A?�x�`@�����ĭ�/E�g���2Ma,`�O��,߽�p�Zm}�t�������X�������� ̟����a�W�P���^�Ҷك:~,W:�[�������q+�?�Y"A/'d�%K�GqmPCA��FN����Y�i[�ȲvJ�
��5滜��)G�k#	����*�ƚ� Vb�h�`�9�~}N�@B]���xd�T�F=�ڤ�K%*��<�#;�B�.��Q�.��������{���;O���H�H�L�L����T��hf����my��)q0�D���N ��K�w&����rmd�y{Q�8A�5|�[�O��m��)��Tſ�@�|DƟv�Z�]B��+�e7�Ee�zӧ����2�lI�T�b�*�hvv�p�y�8�^�F�76h��q8pW�K��(%�}����P����,� �2�.�H����-���!���P\���8��n���.����gP������b��M�+c�)��T(���3����9��CLr����9��#cD#��T5.��5SIE������l���\��<�ӓ�!3i�5�Z�U����<���;:�a�5���w
��"-8�+��2w�`��&�P��˙<�9�Ɉ��%�r�}د��9��n��5{�y�<�"S���^�F�Q�njS���lQAZ��؃$�����e�m~�R� rN[�T���F��ԝ��L-޳]���1+��~���-\�qϸr�na�H5X�X!½�o"��0��7���g���?�Z��(�:�0-�]iΖ��٢bY�q����W�G����Nxd<h�r�ҍ���� x��s��+)=�N�t���:]<׸3cn�����v	V&ч��nM��t+���Ӭ�˛+�|c��͚O���VԪJ"΃JZ��6�
�
����|+ǣ�s��b�A�b.gΣ`|��a4Q�F6�:O���r�5���·$b �j��qbsU�v)t���s�)���o��kd�e��`��۝��	2��c���x�v2�0=W��l�Oڔ�Ar��J�_j�G#���6	�Ț�g�9N������������5+�CH��u�Į4��x��nv��>=�E��~��6�/]G�?Go�GD;���5���D�9�j�+7Lyڽ���������h�0g���S�^����S���>��d۠pw�/i�*Q�sn�94 -T#�Zc��΍��x�z���&���k��1�|��lS�/[6���[���O�JQ�j���:�d��`����T3%���ξ�
ʐ�]ݰ��,vv�!4�L�N.����|�ɋ%���Fm[f-5n�6�ik�oFC0K�n�w"�O��#�G����^9��4t��͇q�����#L�@[Մ��h�2�$T�*��+��&p�J���2Â,��ӛ�2�Fm�-r����!,|3�7���*�>:g>����%�}1��>��_��f0~
UGgvɝF^IǞ+Hyy�Ԝ?�d�E$\ Z^7l���X$}�InLb�4�#��	�mq����גT����]r�i57�"�IY�xu~��,2?�'���E�f�1�.���XKf��ϧ�;u�-����4�J����]�
�e}�ջ"���O�h�?.��� ���nM�7�s�,~�"j���tE����_�Ri�[<)iu��1�4$�Y��\{����c�؟���!�"���I��?���&�9P�"o|!+���W���ɂ-O��+�j�A��zx�)"�eq�V�q��y���]+'}v�[^��MO:�~��"T[Fs��t�1	�˾^Y&��KRҸ�ҟ�Ukuv�O}���b�KV����3��q��2�L�NE�S8� 1��2��]+��������6��`�t;�d��b"9�>�����j���rAm�5�9�$F^<:���?��lě?��Ţ��QڬlM�*��r�A��}W��d�	�\���HesW�R=E.J��q	����Z��e����b}�W˞�H@"�������+S�y���8f%�_�Q��cU|� D&O�L�cɟ���Kҧ���փ�*e/f	�n�Ak�:�i��O�F��H�F�:YrV9�*�̩K�u��1��F$8�V\Աx�+O�6h�.
̕W��᫴D�K\fy��������!�ZhE�	h	@�kwEgѧ�� ���\Wa��Y����sT0N߲IM�^����Z&��;̨�AZ����%���+ٝ�w^f��j�{�f�%	�Z����P^�{Ӥ`�	�\ R	 �Tɤ[�˂U�э��~�_1y8iI�B��U��Y��(���#��*�]G��g�7�h^��-�`d
�x���}�������t]b7�徿�APx�Մ�?�*���7�Ӥ�Q�!;��Q6���	�b�v������q��:f�"��c�R��@���Nъ9jEI	�aL1�S"+� ����s�=���Al቏s�5n�^4�_��%�b�\�+�S:�VwW�Q!YM�*(�.6��Վ�8{�N���#�-��E�$h.����HZ�v=��CΈ6�o9��6$RP��-z �(��.�R����ݪ��R@Fm�U\D���kKVPH����قa/f��ݕ񔏋�eB�H[��`�����g�a�]ا���n���t��\�]>��u	�g��i$`�~�A&s��g��~�CV��]�jl.������/�OC���&E�b �=�J4@�3}�Cu�:+��A���R$��b��g�f��aԋ�x�ꨟ��N8"�6H ��Mz$-bx�����.5;�#�X�5�e����5h��=[P��:�h��;y����Ils��lQe>g��m>!	n�b�����Pޅˇ���l?�},P>�������S8\O>V��]��V��)�m�ԕ@k�Ը�c�����zo
��!��#�����!k�u���\z<��������Ug1CD�%+��oP0a�x�w�8k�p0��+{g�l\�l>��P��bsv�薀�-�ˉ]�Y`�Y�L� 45l-`d�
>̛��L�҄����'
�h�ro���
9&�O�)u�t�k/-DQ�f��"���)����>*Iϋǚ��Ů�aN�M�|�f�_W�M��U�VP�8ܸ��V���?�o�Mp��ɝ[�D�"S��@x����?ή�G[͝!�x�\bM������"������3G��&�J��w��NO��u��{ڡzU��Lv����f0i���wV��ס��a���ؠ"Sz��Fi޻��W�q����u��.7 �>���;���7��\z�Ӈ�M�z�>Z҆�.���N&,�,+���ǫ��R��Ieµ�{w�I�%_����X�N֦q���c��Mg�I*����zm�n�A�{ߠ}n�W���Zb����SP`3����`�NL�RH�.���g`�2���U��X���x�CW�o�����l)�ɘ��ˈ!������i�Pp�x:�l}ރ�����G��:jJ��F�'�:.,��S��7!�LW0�Q=8H��`ē�Q^��:iO��F��I�s5U��F��k���(�x1�D�'iڂ1� � ��"1��-�r����R?��x��T�/:J���`�	hn0H��[T�s�R� c��R�ſNd�k����|��Ӂ<��N
�xy�S�:�v�����<���d�\�L$�Y�>��lx�&=�j���	'���:�{�2dU��]/��qr��N�k��E���+�/,Y5v�.�K2�t�=��c���Ex�Q�KH�ʪ�#�{om��&�m�� �}J��X0&�4�D�h�����}iu��$5�oyE�?wP��2o?��p�^�!p�`�`��\(���cpu4ڐݶr4M�ڑ��6
^�N,V�D��չ"��.��S{����A7�k���r�=��N�rl�NP�Rռr�{�w_��&S�G�� ��rłI�ٱ�Lyt�7?O+}^��Z���K�6���6�C3��K]pq���;@��R<�����݅3a[�VC������n'���w�j�H3Q��\Z���K��-j���%`4����ARҞ_H��dA3�y�B��Y��2��p��&k=�����ٔX>���`�IZm�b�����˱A�VT6B���0��ެ@n	�J���IMkAw
^\�S|����Ѻd�l��"ę�=^�!�����.�XT!�x���������Z��ጰ��b�K��ز'�Le�F�-iF���7ڛB ���~#�C�F{��XÁɽ B�_��
�л9�����E�#�r����=|{����2QjyU�I(��2���qQ��Q�����`�	l�/to��ĭ�c��J[��?������#������s��ԗTGZ���I��u�!���;��Q�P�e�b�Y��`?$�m�JF���������<i�/���a��«��]���z��^U��Bv/I��/Ҿfw\RK��Ls犍��2�Zyn �Lˊa���вCR�4�K�gUf����N�\y��/�xt�M|���!�,�`��_�������ݚ�:CuU,V���H��F��lT���WU�rfu֋��NE��V>��z��	����ݯDWy��Pԕȱү����k��V�����-1
�Izb��8�wyn��I{򠐕/�/ne=��H?��q����ч3+vDJ��o���k�1��Kf�V�&�W�	�W}�kz2��Y������U<�z�5�9%4��ɴ���US	\93�v!�b�kM�`��*_*�I>JZ	��4�0*]��1�����ћ0�u�Lj����{�A~�E�BH>x4�;�FkC �1�%J�)���	��:77�E��8<I=�~���x3޼����+mڬe�?��Ͱ��GS��w-�n�؊�59b�n�_����*]��-�UL��{�M�`�=���v�Ӯ�r3M&Ù�^�x7 �Ul��7��(�LP���]�kk-�T�h^!�"��wa�٦2@����t-��&b�z�J|��N�uB ���ſ�W$�� 	تM������φ�L�9O��+����qe�����)����#B[�p�5�r{BƧR��g-�]��`����&�-��Ԑ1�9]������g�rX��sCӋf͎����)z+�����V�?��8��Xk�ZX��
ᕪ�(����4_I<�M@���bعY�m>��^�o�!�g�|D�+��S�8L�vZ`\/��}d�G-ȹA�[����,5�i��Mz���R�����kgYڳ�!\�( ��9ˬ�`y���,L�Gg��O��u���7kE�>�;�j�� 'V,�IDda���T������J�*����\T�D*�sh��$}�Mg��A[�k܉�G��>��3V���t��n0_Q����j~��՟,[�T����DUy�JY��%��"�B�t#��(�C���.J޻a�<�}������F]ޣ�C����㝖2!���0I�o���`f8L�#����G�Ɨ�?�_�چßa�LdZ~d3�T�:_���!���Z��q������h0|I�k'ĳ(/l��}��9�� �ܝv��4���W#�F��5?3T R.���u������nK�1V����E�*��ZO�X8�!�6�G��M��<P ��8��P�c_�C�^�#���a�p7��=P,��A$#Z'�ы@�ª����k>���:���ݡ�}H4����Eس�E�n�B���;��g�q{O�Q�дT��?�ԕ�P��qJ�]�ü�vS�E�ɹ�R�*6�N�����m�tN�w�(zz�1ZG��L�w���E�ٺ��Z^�����An��e� �2(8�1�/y+�&�k;T�)V�*�s���Z:�+�e��Ӝ����<yaiZ����|�^1)��R
��R`�\������i�}��v�3*�]�*����
�Yk�g��VƏA��cʾ��Yf!
����\����cN��ŝDy�,~~��E�Q������X��<(��t����k�И�@8��C.l-m�I�L�$��\�"����@��e)]T��� �K)�Qc;w��	�-�ͪt��qm@tS�I�V��1��EF�9���.���9ʳX��;eU������j�8��׈�O-�H���6S���=�ĎKg+�d8y
%���X�2�.:��Bܰ�걊�~�ڳS����Q񟞏�D��S$�}�Q�m6'��;���LCe/����ļ*���#��S?yf9��6�I��Yކ֬�;��=�,('��~(*h���y*hb�#�i��C_��	�fQj�3�����A'�'�
Q��bGKF4sMN³ꙗ��Aftd����p�D$9d]�FT�,}��]IO�We�)���hը<��1c֯#u�X
Q�ΎR����_4gs��������5D�5;��ˤ=p�E%���囑�@'ǡ��Q&�Q�������R��j.���Be�A�\�~^ܥ��_��*I��i	�]!{��6��`i�狁�j��7�,� z:���E*�����X�D��jic�^�⭈�5��S�xl�b�o��0�=��bCӃ��PFo���	E��4��s4@J�h؁v�l�:�y}��ڟV�[,���t7� ����aR�����s'R1�%���Ē��J��1��9
L�v%���qX'�`0���Zy������� ��Ы�0O�S�G�L�!�a�����=a����:�#�a���\QX�ǔ��n9���&!}�)����?)=�Z�"Ϳ`���h�Q*5F�.Z&~�G/Ƞ$�r�Ht�������\귿��@�h�җ}�q {�_����[��Y�zy^�G�y���������M��u�*�Y`A����/��x�.�F�M-G⎃���Y$Fiz*�r��P�	�ߦ𼤳B8{���Y�Z /���lqcC�8Bq^�4�b�P}��t2�E��o�_�	~q�����{�s�"���$1�D���27W��7v�2�9о�Ç�o���U�So��>@Kb�wk�\9�
���f�G[=O��(L�do���R�7��fn�=M �WNu:�@o�|By�����	�O�e�+O�k䌴���A���뮼�rJ����B"b��>p���5s���B9��fj,��A��HZY��r����ɇ�ni��TR�e�o�#�X��F䶶|==�$+�c��9E�@L�s[����q��mq�J$N��T�ȟ����{�o�]RKo�3�w�"mj��MUz�҈����!������o5;�	u��NO>����NDc:�Ԋ
��Pmͨh��\�v��G�2��?�uw-���	uATh�R�fɖuP��nF�U���"�^�MO�3�_#���d��ߖ.Ô�oh��� ~��dV18!��i���*��#���a�})�cn�� T�"�����)��,��A���֋\Uw���a�pyY[���LF��?�P\��vJ:7eD�*�%�E�<4��3"����[��S��q˲�oe j��9�{XO�cqL�ȿ'�O� ��o�b=B@%}�rD2�it\�-L�֝��g�)�둍n0tF`�%�ضD:E֮������G���@�"#�|�t�؍k��E�%��2G\lVI�&�B�3�O�W��mT��M�hn۟�p�,nk�yƥ�I�:mO�4.S9�PT��"�hopd�"�d�9tll��Qy0X�+~):ƅx'@\��b5f���`���n�8H� E���v�#D�qil�t��>�7*�@���j���_��L[I~��1�����՛!�"�tg���y�4��J*�F;Y�^ٹ�����f<��Ҏ���9.�Ta�YP�Q���~ڌ�Z�$�䋔�X���|�1�[ �������3���:?���'4�;OenR�`e��p��E�q�uȇx\u��cD�ΘP.ۆ��W;Z]�iz�녆ޏ�=��<��:7-�YZ��1��!5��x�ǡ���&�sH�Xx���dUj�NkB=bX�lo>�ʝ��"�۪07�q���	��NG�K��]��|'rB�(:�#I4J1v]L��^���p\4?0�^�x���k�+(#w�� u��~�*��Dٖk�}��۱�P�����m/�Qg�/�T`�N>}�� ��5fX#��y���S~�ܻY�?\v�Sl?�l�P�fsh����$)�A
r?��7h�.9�:a�<����2��l��E�������*�<Z.+������rx�]ܧ{�pؒ�Y/D]��1�批"���g���SZOE��V�����2�n�%����R�hT�6�$+(���-((���}��9MU +Ie�y�Q�9���KJ~e:�q�T��� ��9���k_��h=�<.�,?C�2c�]!��x�T���C^%#�'�o7��I�昒��k�k�7�5���%Ft��T���S���+.�+>��(vR��6B�`I�����RL(�C\a�2�5)��N��G H#^�=۪)���f��l�$ŐD# ���Z#\�W�=��r5�-��}4wS�r���?�S�"��$oaT�����6��k�,=WC�]փ�-<��Զ���	�����a�������owy�-��8�`�+��CU╣�S����Q���=M�;�=�­����\S|�ꐾ�Ic��|�q��L�i�#PL���o�+�u�;�K��3�`���Q��sv�� M���S��-�`r��{�)��Mx���Le��ô�Z?�m�;�~�Z
؋�j��b����hm-Zz�(�5N`��z��o�d*�X��A&�)CK^��nR�ǻK�c���HL�%7�UtH��;)w������{i���?<����_����wX?T�[�e�Fq?�����Y�O#��~�B�Kq��+��#A��F���Cll�x�h�V�o�S�R���U%��U?T!|ކs=8��օ�E�$�0��!�����ю��h�gW��ol�Y���뾚����Ϧv��knlC ���]Z���+�~�;�"<�a9�D4'V�Q؟h���t�H!�ޅ@j��G�3�! ?� �䰂���p�.�g0̺_�~�m�k'�����[�KT�0��;+�B*�5���E�>gh��(�mL>é����_)�W�J�����	�R�$������Uq����i���d��@o�����z,י g��k.���IE��Pd��%����i�� ��d�#�}zBn��r���3�AY����|x��������C�M�����	b�kɻ����5:�kp}6��A�{�+$K����z��)"�Ǩ�>�|�Ǉ�N�V���ͷ1ո�L3��*Zl�8�f���Jx\�������i�%Y�5��r�� �&�IR2���������RٕU8$͟���p"W��s|�h`U{��pE:�Ņ�gLO\ȗ�zG�J�]M�V`��O�㕜=n�������E��9�7�Nk��VS�m��,-B���Xv��]:��ji[����Q>�!@׿P�c��q�4�N�500�����x3V+�f�}�(���7�A*C��˷Y�!������J1���yMәdش��g��%d,�=�L~Uu�?�U����uUE�QĐ��8߁u�ч(�4���5A>�-8�f��WX�m�k3P�/����0��X�K\n��l���lùLh����a���Ò������`r��U
I#E_Cp�ؔ�
*���J�8/��y�-�ڤY�?�#�O; i�`���Z����/hpc�U����6���W
�8��WݯC֋k�	�V�S���vZ�B�m��X6>�)�hfp78�h�k���߃��8������l;��������2*1�3{�O(?\�C�]!l�y���(t5mu^�z0��-\+�(�.�랭�����`q�;0̮���+"��S�2�bnRF��a�a��OG������F��
��w������<��r�5����TV�P]�z�����:f�<� �/#T�.T
X{H��$?F�A�P��V��5��0���#@�uSʻ0}��cZ�l1���������w[X����c��^7`�̃�0���
O����۩r�`dg��}}�)g����6y���+�Ky���GT�z����x���wV��E���"����d;@�͜�HH�ڣ��1¦*���5'g���5�je�xPx�o��)B�Q���"�Kf@���X��t�&�����W��� �(�����D���I�	�B���ǋ��uP�9/:�b�U�`��b����&�I��ԓ7؟����̊�?�2ԑ�ί��¾kCnM(,Nت��#O��w�����y��z���[8Q(�,GЊ�ܦC/�Z1�w�^��F�s�Ξ�]��N�Pg�-�3g�N�1��)��y�嶢b�"���쥭�/�~��9gИ�)�l�0��E��d�w[k�d�ɓ��j�W����`�R]-@UJv@n�w��ݨ_�z�V�w{�%.�8Sñz��b�L���]u��~���0x���󑄛�hִ��#�%T���)����(��`2��A��{�� ��i���BUoS�$@�γC]<�>lF�������ᦲ����[�'N�z��oص�^�B�(�"���Z�އ��o�%�A zS��1�[�r:��{��ɂ���VmO���^������m�m�(��^KZ�Sꪻ�g�,�g��1�l�4I��.KĠ�A����y�i����}��`w�~"�]10׷�Q��3~E��j
@���*���7�Ԟ�<p�tq�v��<E�˘$�H�a'���X9������ö�Z�;���9 �%e�a�M��/�T-��n��z,���i�xh����&�:�JВŋ#/�J2W$�v}�nǥ���#r�g�j��1���~	c�Kb��2�+�=�ת�L珮�|7���B\8x#��<�Q�����9?\dWWQC�]ArA��g�?��=��r����^d��7�⎞���L�h�~� �Y̶���F���9�P3&���{�S�h3������|������p��CQd�	��V�"|�������i/b�hG�9(�G�T�e��� \~��k�͚4r�q�=sHA�7����z�r|�ǉӋ`rޖ��Ⱦ��w�u���49����k�ŝ��PLa���U1�*ח�)�Z�'f_�2�p���t6�{s"��Hu<���(?��g	�<����֕we�̔Q�B}��Y�If��uA�
�S�9�)񤋐W3�kۦ�J����or���ȋ��9{V)G>�bqZ����9fo��Cs"�Z�#$�"rw��Ҫ6��u�AڞF�!����e�N&`"&�(�İT9�ă^׳w1�kǮ���"!�n�y�&�M@[����~¬#�NT�&����⯲wrzd��$�����#��(g�as����y��с�g]S��Z����/w{I�����YQ���2S��
���A�4νn`Ce�n}�3IWz���FF���Ec�	�==5~~OH�&ɲ�N��)X���@z�d_���$����4��2�Z~�a�5��&ĀO%)�j=�vEۮ��^G�n3��9�k�j�SZ��0n�ؠ�����<{�N�Xg��@zwU}sN7�v'l�#��%�ƾ��g 9����s߯PGEY�ʠ���"��Hj�w�{�s��0��؞g��B �=�/����?l'KE�n)�`����I�a�My�Om����?a��u��rr`	D\_�����=�v-���Lv��U��瞲i��|�V���,(J���l�VI�Pȱ/֘�-��j���Q^�@F�Y}'��T�,B���
�����P	�P�:ǟ��&˹�'b��XH�O����ǂ�}K&��
�Z�k�ܚ�)g,:GV�ʃV��vH��y��3 ò�����'_�AeK��H�	,�C*�:<p�5�2j�D�9�q��|M��D�r���b��_4/\<��o
!H$ن2�$���[���t	0ZER���RQ%}�z�7�s�Q]����r��U�m3b���k@lkQ��8Y�*|��w����OV߲C<���mR����L��=�@5-�������m��Q|J$ 7��5\����θ��j�����:�ȩ�n$y�SN���p�%��{�^��nT[�TH����y rQ<}�әk�3z!W��S��6�?�T �z�35&݅P�J�;v0�����#�ѥ��m���SQ��珖  ,j7�Ӣ���`�I�A�^�*P��a�D�T�T"���i�{��9���X�J���q�����H{��8Ө\�Ȇoԝ���P��u&cd�	�E,�ʷ;I��]���V6ն#Z��¦e�%�N"�,�r{�q>��V[ө~�F�H誹s��n !�t���!Ô#d57��<��K�zD2y�տ�]�C�j���q�7���I	u{���'�v=y�l�#g��e�o�_oŀG���~��2��|-J��\*U�DPA>^��:~ϲIN�N�����Ѓ��{x|�L׿��?o8s�5��Q}G~|���g���":��o듑f�CM77�����R:��8�>n���ô�M������G��.I�d����<臾�_ԝ��Q�kfY�ҙ�b��/Pz�r�ȀC�d]��Z+o�	�����	�d���BȂ0X4�$�5\/���N���2��yR) �8�'�j�8_��Q��ӈU�ng�������1bƨ��qd� 	zwA�5M����X@�|B' ���`ѫ�HRJ�%�o\+�]\�S�c3�Y<J��R���h£Z,
��M��0<����zE�ۀ�����r� �S��YF�����t����7vyz�)�S��zI�����3�Z��x}v�gU8��/>���6��AV�g��{��������4���o�c�j8A��c�]��V0кۜL�b�����y�~����j,sRX�qA�z�3��Bv��[Hl�Z�`�6��/d�/�yF5eV�F�p��R��qm��hi�����`�s��ᵴ�MEjs�q�Ř�ڈ#��ץp�,=̝|�0y�Lz��,�,�e�ð��j(�#r֛�侘����X�<Rt�`�����r��7�OR����A�t�7c��F���=��/��r\��^u��\G���c�t�$�޹6��C1�@��TE'�ˋב���T�q>�T�K�-$J�I���	c.����`c��^);{x_{F)�/�[�����1'�)�)��MU'Id���W�C������)&����9��&�����l�����9n��g��E��vvР�+]�;�Pw!���0!� 1,] 	�����Z������D3H����(��s�tΓ,Ö�PW\��"'���Wa��ݶ��E��� �)dx��F 0�(�32�Lx�(��3�sDc�?[KQ�c�*,�R9]G�{1���F�D��g ��~(�m �TS�9�JNJ�y���֙��3g�7e������r�#����'�G��c-,Ğj��Vgɷ�B�|�f+i�ې��YC*�ش;
��%
1�A�}�9�Ȁ�x&��=T�"=j�-�����1!��&��/ֿX�n[:��/��nm�Iֆ�-{Hq'�5`(��F!Z_<��-��ES�H76p��á�%��I"�7������ζLG\��{c� ��L�����hCI�+�L��Y`J��I���yJpd��õ�fb�� ��gMb�t�uڅ���)��q�<��eNX.�G"ɯ��+F'猹]R�k��XT:�7�H��#��|@4���Bp�A�y[dJ��v��)	c�1���@O���.Wu�ݡB��fL� I{/hRF�t��p�5��5��x#/�ޙF��R��:�Ԃ,kf�`��W���n�N.ih�Uͯ������B��)��4�q�~�#߀��c3����,����<�w�E����S�e&tW�D�S��@v4��������3��l �d�����\�k`e�`���� Qo�$ĕ�� 
>�~�h����In۫�q��7��7�H�tAW/�Lpm�u7.�_��5`�T��ԄRlL=�J��]���-���	Ä�I��}���y���i���\��#�y�9�t)�XŞ?/�l1�S�����?(�׹c��Z޹f-m?�'���X�Ĺ�ґ�rV��M�O�EQvۊU,6���v��Ê��k�� 9��>�M�B�=A]�3���ʥ񞦻M�6Vn� �ͯ�mn3q�z8l�#�t��j�<.��@���?-�Ki�[T����xs]�1/�_Af�{c:WRRi�{��Y���e)^�n����E�ۃ���hM�t�<A�u�H��hq^͆a�0}�h�9�u���Ti?�|����J�ߛ������^� |Hƒs�k��T�l;Y ��L�W�I� /���qj����\��g'{���GY��a���<����3�!0!`�#n�0�ѱ�y��?-PM�Ri��cz
`-�,"��h����f�-����A���"��^�h�%ƫNV�?~��}���f�6Ydm��?b�/AI��9���q:��YvIPi*(��34�%�8jip��Uh���N���k�ǖ�:�Z�֓���A��7L���C��`��p�Kk
׎�6g;�`�i�[���kj,]#���;��@� 
��ݙ��VG��:.������4�*PI��f�L���0̰�i%��C#'�<�ֹA�����t~x�u����g3�Ѣ�j��0�q��%9���\>��@8ܦ �U���"�]����f���Zݶ��4�.�,/�*.0 '>r��!�g1�fܫT��]dyC~E��U/��Z� dY�Ds��b�ۦ��^�43Q�c��<��ZZ@u���w���t��u�k<���
]��J |x]v�+��%����@�����-9���p����0�1ŮzD
X-�Jc��J�9����Y�M��$�4 ����Ozo����\�������$:��\"RƤ=�M������'��*
��/)�f����������c�1tք�x��-�����>�+',��D�v�;a� RS*��2�ǔgUOH�<�-e����q�D/ vZV����@�"��� �c��Y\h�z"B��"g1�e`���GV�����
TDS0�o�� ��r�Y������##�ޢ��F��q��a�wo#qPF�8��8UD#���9g ��G%�	1��$�/�p��Mp��v��r�:P� C"<�c�C�A���P��kr��|bE��=Eφ�G����F_�+��n���������C�^rW�g3����=�ΏK�3��ߛ��~O��nTG(�`v�( @��4������ϸ�d��P磢�x23�5麛�X��硶c#Ux;�t��<ϐ��Oͷ���Cl�2�01T�0���|qx ms�[=���ƬY��~d8>�Z�ۂ��>��t�)1�B�J���L�lK��z�K0��TV�w�}��)Y���E`{C�ˍp��1$���`�!-��a)�bw[*�<춈�U鏶����/���70Iݶ��B��9�a�X��$B���a�q@�^�$��؜�Z"��A��������I�_��y�>.�҄h�ZP��j�!m�J��^=���&",y&���p��_�I��t�an�+�\�3�D�8���@���bi�U�O΢�����R����ǈn*���p�C��S@�����P�zYo��1�B���":Jl �$��{���pm|��������`5��'����0��HW���ݽ�/k�&r��3�ﳊ�3L%�����u�u��"�@H�����(T����-�p�pU\ ��庥��d��P<s٬] �ˍ 5L2�솵a~.�Q��R�ؒ�օ"M���g}��vDJ�^޴����*����AQ�X��>���Xl��ݨ�׹���-���D��"��G3Z	X�Z\��'�S4XlEz����!���NĐ�@ �4gI}󞺤�\�g�e�8���K���W ���I����D �6��d��g�5|�;Y�$��N��V� JB85N�i�9�$�V�:��'#�+�q��M��*��Ɇ}O�������j+^Ⱦ M�p]o�A�.�̾gL��Y��z���V������G|�ւ��Q"RB5��)$�/�N����m������ͻ���0(�� �:<�.Zҥab�����`��,Zx�Dt[����bƳ9�����jr�5.P!����\�͡Ι/������o��{���*� K�"|0����cQ�SxuJqM��ߴ���[�I?�
N	jtD|϶G�>&M,z�o��Dj�k�=�Co�� �	؜��Q�9��I+O_H4��y=v&��%���P��M�6�3zA�������k�~#_�L=V3�+`�1���X��/�WI���BnFF�l*�r�4c��Z�.<�#Ő�N�m�w��U7N�*��J�=й���)��##%5q�Q�R�Z��`z�< �E~�qVR�r�
��1��Nf7�W#)%�2����Y�c�Nk
\6�r�Pz�&�ϱ��i|>Z�B4̭D���׬�bү�g ~�w4WG{"�gV�I鼸R꧴C ���j
�&Rk��@�[�C=�W?���͊��2j\�0�����;��ʨ�X��K�ִ�ߌ��3���Z�����G�����8�1�̕l��*Q?ߖx�E����!��7~�g$���/�5hP��t썐��1/��C�-7��Ҟ�ݼ�=�h����a�t�]��p2�Z���%�̕�8�90�\^��v�� M�A�5�ji-�䊛�8#���m�R!D�	1�J�9�I�+��Ln�й��B���w�}��h����fM��U�3?�cTH��j�.u�-�g�d��H�oH���Z��F����1 ������?�B�	�*~�)I�s"�j6�
����S�!塾����:���/� ��n K�V�Su/����X�W#s�=͖o8藸5�3�1i�VLH�*�@:e��G�൧鋭�t��N��j]=��������i�(q�e�L,i���/�OOa�YO/�t,����&?L�K�6���m� �2cR��t�����j���� ��Ϡ�M!z�����G^�cŌ���o�7B{�5�S��B�eRF��/��\�8a�� ��T����#j���LF�X��q�M�a��7�\2�T+<�Rh�[�L�mߤ�h)�7��C�|�&��_Yi�'ԕ��9&+p���a�M��R]v�����#�(U~q}e� X��4<I�C.Z&:�g�(ݛ�h��QW�z�J�L���}�F�ʋ�M�?�p�\�v�	ma��
�4����dZq[��)MA�(����9���{ Ĥ��/������j+�L�	Gob�z����q�ߊ����:���/\�ڔS�}?��PL�t��O�	Z��+P�C����\��;l���[;�D��q��q�d{9�i{Ԩ����cA�\�|}�N���C�k��+���sO��F,ӧ"2�"HH�*C��F
�Ԑ��1��>��+���N6��J�S�ZI����baz`M�`ނ��K�l �:#�Nd/�+�wv-��FMa��K���X�cY����
rN������'.n{�7�e��툼�V�g]��M���aR��{49��\��� �]܈_���PM\~�?T'o��W�LV��J���֐�����R�fw��Er����5�����`ĔZ"�o5�'�r��x�s�dj�d�N��Y��C�M�V�&l0��������u*1�w�O2#�G�<_Sn�a6!1d� `�p�>tN�6&�!@	��4M���Q^���?��� ��i`D������YO'o� ;����BT	p�oW2�/\��ډ�,w�1��]m�g�z��TGR��ㇳ{&�_�K�\�l*��ĐZ0Rwlwf��oF����[#�.��Q�>��-o�2�kg��%��(/���`+��`�1����=9v���Y=ie���U�ƳNU�}sxk�!p��	[�;�z���β���]K�ǳ!Zz�����+tGvo��QN�@7 y���iJ��
��1˷k\¹�� �[6t|��w%Bǉ!�����g���y������΢��)�
����7u��~L2�V��JLB*����P�9 TU�D=�Fo< �IW}��>F5O*��뻼J�����X֭9I|K+�¾O��f���Ts��9��H��ᑒ�9P� �A[�����N��4��`��*3,w-�bވO�dfW>i� O�9hM�'~͆W����8~��V}R�H1�L�:�_�p��߀R�[����ua�"Hi�52���*�-�����b��#�Ԇ��v�2��s�XQ.�!S�����=���+�	9���Q�=��ۼO%>TL]�L�#GCՕ#;H	�X1�/�W�ϒ��U7yL�8W7���ܸ� J��Se[ă���Q� �,+>����qnuN�f�+����*=�8;����V˜�c|�(�|����vQ��czs�:0���]��l�+�YY�,S_����+�46n`�H[M�ڜe��^Y,ufP/ml�m�[��#��A�:ݭJ��� |sh:� 9l�҈���VcjԷ������������}��$�Cr�?'ĸ<}@l�����Wޒ���g Ƈ%�v�·g�W��(�L�
q�����|�������u�[�V�Gþ��t�5{`���*d���Y*@ii޲)(��;���М��q���YJ��
 2�|X�]� ���}�<��ǓT7�F��5=c��P6��O�\�?2�ݯ�W"h��$Ld&�� r;��̔i{�eh�Yv%����M�w�ĭ^�f���.�4w��W	h�F׹�B?M��#:�M�]�HC�B����Őip����9�sV�[?�d�(=P�q��b��Ė��̑�*�v֊�1�k��vɠ��?�Ed�L�9b�t�#��[�����#���6a|��q����eG3+D����3}�֐�z��ʑ?b�1�ӣ������~nL�'����Wf�-��YB*���ex/�/	�i��j��a��E��y�	�g�hfO\w�i۫V��F��J���f	�iI ��E�ٜvUU��_=~4��"���0yCP�ˮ{~T�{_�B�}�'{8$|�:�0 ��GZ�1������uz��
�0g��"�����K�]������pӣ�?��3�Iƪ�\��_������%��,���"2�ֳj$Rn�*?c��<�|*���ۛ-��!���z���n� ����Lυ���5�� 4����g ��Lk��[>��>���fD�[w���L�7a��wr�ybs[�4̓��ߢ8���(5����QC�C��� 7�O�=�^G�t�sеÖw|=���t�a|sٗ�� 5�ky�P;g[�~������r�t!}FX�O�`zR�#TJ�U�/t�,��5�ׄnJ r���O� q ����� ��<i��w���.3��������Q98�l��	����8�Q�)�����j}	DlH2��K�P{���Rp���c4R��l��v�D���#A#��ĥ��
��O�P�jT�4�/K��,n�I��Oc�eu�s��?�fĥռ��$'1��C;���?׫����r�V~�~�����$�0�Byi�����~+�h�$�C��kb1�tvi"��SM�#�L�M�����(EŠ`��_�#⨧���:���/�uB��Xc��N2jì[�������'>�Fc��=��S��0NF���F��/rJ��a7J��$;���C��X����)nh'��簺:.w�ul��N&�%�ŵ��ƻ-MQ9��&�!,��.|��W=&Q{�n	g��%�#h�}� ��Ӕ�Mo=����5~��!Z���h�1(nK1��<Q5D�Y�V)_��;z�;"�'m�5�"R9b�(n��J"�����	��u��䌬C1!*h��]PB��8� �fZ�hzKM�h��+���$��t��2
'���FEOt���R�y��%�\��nL��@%	W��W
�:C"q�&i�{S�
Ǽx�~HEwz��dR�]V1�l⩘��y8��e���M��LaNu�vʛB���<qd�Q���(�6ݕ��i;T2�0&yC��12���p�w���7-*W4'��Y3����̳��Y�a[&���S�b|��*CϮE:��z�����+K*������{��Q��F����-z�B�����?K��)�>ZiK��j-�6Dp��c�`�K�������Ė1Q���㢸_4�1"�Q��(�d���ï��և�d^��V�c�}�S��3�sXj N'c�>H�;��j4���xF���zdy3
_��(Mq�c��V��|��D�j���ᛓM\��]�&��u�D$}~��M�7�����?e@��1@��]�08��<h�]E�X8��c^C�1@��n)"w�ºL���tmʱ>c��/��
`��]�{R�^}0<Q�W�G�0E�ɇO�׺����X%�����,|�n��W�v��2���s��)Lt��tf9�Y+g/��]�z,k�����SX8\Y9�
�X ����Z�EF�f��u�a�����$3OJ�#]�"���wE��o�"ɞX��:vQaj��RV���FJ���I$o�[[	݁k�a��V��ćZ�b�H��,�C^��$�*\G	3b��*秸���i�0�'�y������X���������i�嗸��3"Pִ��"a�	9l�S˾-�	���"�57�){58���	7������ƥ�Z,&	`h8M_�0����μ[#�z�;GC^�yWW;��s�{lN~ƬJ
�
);���ons��HF-Wn�u��EvL�fC80]oZ��PQ�ʵ <]�� ���w8a$�o��.�>@�t�S�b�I^n{P��sQi� o�QϘG���ޖ>�2� ��F��g�RE�3?x ����/�R�� X,J��;�&"�bo铞JB}6	���Oc��DD��"�Q,lg���G��}
)u���[�g�W}w_07�@~m>6cח5_-b���T���� ir-�dXU�U^5vA惽NC�h�ʑ�녣�q���K$��  �Ha����*�H1�:�z!RFswRi喰䌞e����j��:ʋ���x�L�,�=w`l���^a����y�=I�_��s��|zGx�� ��`�f1zJ���yn �����T�P��u�����^��E,��T78E���A=���y���LH7�8=���l'.����x)&
k��E�G�H�!
�UV�LTS�|��,��;��RH�Į7� /��/�/9����>�D׹�Ѣ%�1Kx�����&�^��c��6��,�/����9�m"��v#���j�:g]��o�	@�!��ӕ��m��#�i�JY�B���R�����H`%&FJ0����v߱ˠ�S̠���>p�C�	؉GHt��b(����Sp{�����@���F�9�(����@��UoG�9��}o���|�jD&iM���N�o��A�)t�NuHB��p�gZ炒�]k���	��Z%S%	%��[��)��^|g&eMNk}sܚ��q������$�(?�N��fn���*�K(�ŀ��ײS$o��Km]@�U��]�o�6���Y�?�H�X��6����<���Wk.IOJR#Q���BلE:g��H�����b�R����ɮ�� M�j�h�*'���EK�����=!�죸l"��&��>Y���I������'5��]�<w�RR�aEd�(�"�"7u��������!T[�y�����Er��%�w|�=B�6�⠧��`O��3I@����ȯ]�g��AS[�L&��_g�E@��kN�k��k�o�z�(Wצ���3)����0��6fG���5ٙX��(Jt-=F�J�̭�S�lŷh�J�����g�+SF3(�"2[Y`834��=��
��FI��Zg^!�\#�.��qh8�����hXs� 1����0�PݥQ��)�������6���ƽ��!Mg=�J&mE%|��a�I3�k9�I;���-Y1�$%䲸�4J�,��^&���!^5�b��
����߻��y��<�\'�\bA��'�=��F�@����s~�G���L���o�9�go#� e��~޹�Ѳ�1�C㛃�,Շc�S�P8�"��g�r�oφ�ΊC�ZYb!;GVѱ�g)�/
����@��M/��D7�vo�������O"y'f�Ϥ���{�h�9[>	�?��/cV����}c1y���޴�q#Ew)0Gb�[�� D��o%H���\�t��gwr���_������3�(b0������x���7ׇ���� ��F/p?h���$n���a��HL��E��S賰G�H?J��3Gg^<c-�<�Ć>(;����y��-4�/�E7@��]���49�W�P[qcF��O��o��Cy�X	���ܩ�������k󏭆=�o�j�qH���O�ͥ��KO
��N�mj�`�h[��l�6(�D5�'�*Wk���^Oul�,��m�0�$F=�}�Q"�@�a [`�@.�3m1�*��e��8��<셜�Ҥ����,��{�`l�;!洵��dX'�U�]�M�v�J�?�D�H<f��v�5׵Cv ��D�G��,U�̒H@�%�'�j'���덐�X�C�9(;���G�IO�헎�h��E�~�K5!�n�d��g�3%�dYAMD?M�c�H�� &L�\�7���g7���n�f��v3�LT^���m�QB�m�%����Ԙ��&#:�b�yo#[$d��0~"�sqA����I�F�<��d&\��6j�?�	:ށI�l��C��Q���K���"�|8�,��Ly����̇M���1����-�� c*��S�F����rz��@��Y1�N�[t���J��d���fmN)���
p���3��_�f���Tڊ��%;2���-�j����њz	��t����wS�_���~�E�����o�}+����C�t7u���I�t�N`��[Vֲ�.ttv�
-dH1��0]����$��#	U|���B���g�\��2uƕ��� �Q�2���Å���r݈R��2�s|�MB!�EY$=�[XX�!�D�`�*O��(�Ƚ�n�o��!-� �Q��>N	]��8N̈�����q=]ad�&m�x�l�6j(����HۤQ�/ɕb�����|1�����{,x6�E�հY�<�~�ЅOaM�妼;�4�X$�g_ ��O��cƵ?���^�q����V����Q�s6P~����kЭ&���+�w���J�+��Kw��˂:�8A�6G	�x�k��O�i��ߐu����4*0̓��z��Fe�_S�hZ�Y��r�q����?�n�D�X�il Z(s,���8���h��E��VƢ�9� (T�a��_1��7v���y�b]�i�+�A���S�ݖO�C����w�E��G%��[�ַg�3�=�$���e�'�d��wr?�����n�S���6Q��1�L��@2u2\�Av>�еw��ޕ'���@�N Ӥ��C���g]���K_�ޥ��p>��G7�!�W�t��&V���2���W��"r	D�P<tE�,Wã����E������ա�D�}�^b�,��r��Ui���U��/B&�p#�mBZ�t�$;���g���#����-9�PP��Cu&3J��+����E1
���.~�ga.����+~�3
6E���͖M���h�ucW}Q�d�uCL��A�W����L8��?�шd��9��m�r.�ERpk�5ŵ��b���<_���|�{N�I�����0O��ֹ|1ã���&7g�1�7��vϊ	�t���k��V�����=�zJ{�q�($^c��
�h��`^�lfDT�n���j�[Z@��p��e�ʀ���+�ʎ����.�O�QX���S�ށ����PS�H�P��W�#��#�&��1�a��\��e������mF[ˏY�AS͡�!�Zj?�x�φ�?Mdo���N�|�e4�==��wB&!�ű��9��R}����� �ַm^k�􎞜�l`-_KI�s(r��R�z�������we;`�<H܊�B�woD9LG$��]Kd�<zy+���P��tU	���ח؀��h���N-N�͍G!��A�y�U���ȖjrX�e��\�����!vN�/(���1�n3�ے	?kz6AV�>���јs��ƕ�n��AW�D���������qc�^tNV�2�x�˵�a�@�4�ʎ����ŏ��,mPY9���ȁ#7H4��Y����Y�0����n��i��o�}S��M�n��0��#�N �|��i_��+�Ո�܍9����Wb`���t�:`�.6�S8�niHw���gʾ�\�G���ަ"㳥{K%f��[AE|C��<`�$A��)�Z���+q��XbqB1C��z�{�~#��	EsT��K�{��4���*�W�<U�+���t�XOn�-1~xFfU�ć�v1̒I�oi�E�dmb5~Ya�����7R�&�ݹ� uj"��JC���`��\�i�U�0���!Rֽ�?=�껓S��2]à�t�0z�HVPW�?x�&�G+�H��by�|���7<�S��!q�ʪÃ��#y�xy��b*
���m&�pq���G����[�l~b��>�]mR���r��bs8�[{�P;p��G!Xn��x��-5۰d����@7�`B�̀v9Լ�_�$��p;�6+=s�'�s@�"l�'.�_�����O�� ���	�f�M��ɒ�a��r#g�r�2��9��.���!8c�4���'�Ӕ
9��n���n��zӧ
�����=~A6>r�؛$�o?I*p���z��-�I�o�z�{���3�L�{c��;@12���l��8K4F�*�|��+�G�k<�+w�י���66[z����[��~#�H��Cr�q��������!�ܾ녔�4�����@Ŕ�f�g%�����Ҍn���aeu25Nl���'�e����5l��.����˳>��B(f�L|�y�0�)I��!���hV����9�E�����f�<�@Wl�A�`H� �����*�|��!���ݽ̛�wjaqJ�V�����B$���#�H��՗�Ղ"�f<�R��a;����|�.?�ޡX��9�
��!9�]�����̞��Ìƹh�FdP����)�0���s����I'qE��<�ц�`�׶�>#�V�V�uM%�t\�ǧP���^���rĝ�=yoY@J
�x����TK�/�̊�zv��L���0!���Q��M'�wsz�{X�)Z�g�b�'�'�B�5(P��/�Yk��x�'���L�*�@�D�i��/�)Bl֖�8�~]�ip���r�	�#1+��*����jUDN���rܨ�HM}|���A���G�/]��`��;�,O�͡\�GE�fq�����肜8�ϞN�̃Z<ˉ��s�����{n�h�2�Ǎ�A3���1�L9�<�al�W���-"��뿠&"*�UK�oZP�� 7mI�I���������W���$Ưv�����c
�z��]_O��)�`ڼQh���K`�SgROn��λ*W���������F�m�[����wJM��)�]8��l�S��m�9c���n��̂�U3�vk�!���!qF��f�._���������d �^׻�2\a����)��Bw2��$�C�׹�!�����V@��
>� �;(����/K�u��H��:4��������,�X<>X2|�� )H���u���/1��Ũx�4X �T(�{�/d;��0'�h�����FT�=�Fpv�4�W�RTax�����	���VŲ)ӂ�)\æ���N�ީ]�E�92�+�AH3�6<�o�����<����$4�u�T�[�	���៤#��'�,,�E}�rn�Şv�R���n4����?G�ނJ 6����5�m�>�&0]�~���%ym���U��eO�0���2�qb�6�F�Y�)QAW8��).K`��n�X%O�|�F��%ѓH��Ic�$�`m>ʷj�� ��]�C�� ���@�?�ɪy�UZP��x���ZX�/�@{�R�p{;-eVw9�⑤�(;�Dj�!�H3���_�H�����o�@̳�8� �J��K�\��/�|
��=�L�t+�I�壝����\��s�)ތ�.7{o��a(	�xg��ʻQ�z(�渦^F	�Of ^�����u��jiHg���,��04�@j�ml�ծ;�D�cFk ��a�ِ�NX���荼 �F���5�ӆI�R�+G ��Q��ۢ�ݡ����q�"r����Z�h�/��;�����צ���S�����
V�=��Z��K����΅y��Dg��}A�;�������g�DR���=��ؔ�Nʃ�h����欈�i�VSۜ��1뱾#�+Д��[�.0Pk[̾r7���h�P�z�<�.�~��� 6%�Fa�Q̻���k��5�7S(i���k�u����
26ootd�4
���I|���P�v�8�b��H�EM��¦��M���U���b+$̘��w�N�ҔxY�k�	�_�����v$�^E�vO�s���ٸ���G�DN��6�g�p��h�&kc�E���`4@&#�
w�␢F�BW�|Iˬ���4 |<!�m�?�/FC�q|{����N!�V� J���w^�9��!yuF�n�yc;6�ht}�m� �s�B�}�PO ��U	���y��P�v ��]���N�v6�w�nc��If�*�0�	�?���?Y�JR��*q����5Y�J�~�*�������)N�ߪ%b���:Oޅ�A2_�H ű��\OS�����ɡdR@�n��g�n\	�|�'��n�u�:"�����?QB����f�(�[��ud�t���YW��m�k�B���[/�)�!�:ȅ��)̲J@��{�oF	!"#�u�]w"oK�4� ?EE��d�9^�
�jF��N���p����y5��f�$���t�w�H�=�E��R��<Z����lB'm�M�Ԥ,>�5\�wE���	>�Uw�n�j�_�$���}��LȪ,��"�m��̆����"�CH�p�V*!2���8�c�xv3csn�r���@�Ҷ�YB-��eƜ����nNS��BqD��\�t�!J)+�x��q��	1:��aؗRa�����k"�K�)��;�\U���~i���PZ�����#�{W��o�`|$�0&iOew���%pG{ɨ���jWˢ����	��i.Z���x��v��eg͖M	���C�)V�a{�N ��>��"��\�}�ֆ�,�i�=�Ej�z|�T����_e"�Z�|S��Q]B�dS��Y�<_H�`�U��?m�%����)_ k���s[�a̟b<^CD��*��3��j�M��k(��@�����eV��R��[����h�"���k(���^��X]M�e�dh>>����O�D����.艖b�#s$�v)#����AɅT��T$��ŸmWQJv���� NT5�����-6�D_���w���6��$�W�&����-�(����Z�.�V����~`���l�� ���#7�5RU��D�"��Ā˓���z����^Dz���k0(���B��6��:��.R��{3o;H�}����Ӎ������u
�-���۾1
|N1�0Z~�sݷp��h@-��[�k&�)wr�իF��V�\��������x$���d��������t_U/�dz~��x�zU#?�����<R�x�
)�^#�:L����d�Ɔ^�$[Ol����+�4U�`�fN���6`��z儛�ā��*^Y*�7�u*6��ezx��6����Z�7=�[�~(�C�_I(�L����4��-TT��n��;<�`�Z������f.��C�x���,7��<�k����K��6��.����n��U����τ�sSV+��(�݌��6�J: I�PE�`0���trGz���<n�YI�N!�/�dI�����{�>Pi����Զ:�25o��E���\�������`(q"2�k�[��FW��l���e���\5��V�qF������49:d'�Kֶt"�i��>�糐Ɵ4`��@g�����C��$��֞|�	G�{z��`�����9�%I��/M|� ����c���4Y�M��~~҂��fʺ��q�1E���!�ȖT�=};�O��6->e�\��je�.䇘E���_�֮���H��l�<�TZ3s�M�jE�l��was��m{X9]kAR+�y��~�AiM)��o��e'Z/v$����=m��(��	����L[�^�MEi7����N�|�\���	���ɷ�ێ��.���H��uLI��c~�2�y�"����Wn9o�*'UC�3�Q�*�/�F�6�`�OS�ZG ���-���v�q��~����A>@~<jw���̐��7���]����.�IW��<�_kC�0~�D#�슳y��}W ���I̋�n����g�?�T��R r��B��l��O�.������⻒;��������*^V��pRq���ZGU[�*�p�-P���+Yf�>:h�	�ap�W�E��]��w�h�o&��&Z�e��~���$Ġ���� �X���	7�����B�A� o�i��(�;�<�3�]U؆�3�KC��4{��dp��g~�=�L����Mhel�ʀ_��@'>��afi �d厧�#��p�k|4� _�?`�/ꢸ�{�L6�����,������k#�P�u�
 ��c(�"��i@�qT��?�ǎ��-�`�RTHI���r� ���C��VW�7�A�%oD�v�3"�(����t�b\����,� ��@~�Gt�	�S�
.�%�M4\�G:�͗J8�]Ac��=3G�af��*p.LA�Tv�f~�&?̅�C�����%D��3r����h��_V�z�bp�:mEBRm��]ea#�]������`?HNs:�9�^���ܢ�e6׷���(�wN���*��H����ģ7v�s}���P���&�.�#to$��;H���C#�L]���}ٳ�9t�	ҝ����P�b+�QVc4N��J���K�EX�V͚�i�I}ƀ�9����G=��y��ȯl>u0IJ���U�	�$��|QY�C���9GY��&��� �̜�\G�;�+�Th�C��)*t�����|�eX�
o��ݫ�U���Դ�I�]�C��FT"V�)�k��0�H��m�Wb\N[������HaZ׷D��B���7ܔy���:�,�y�%�Y�k���������O�f�30+a�@Yꪳ�1W~W��Czy�d�:ehS:��w&!c����j8oP��R�.�?y^�n�:[ ����`S����$�v��]�� ���Ts��t�x~+�_�Z!�(����Cȴ�B0����m8IŎ̈́v���7� 	�=y�\�/��FiH���XքSJ�cE��D<=U^JU����|�<�܏�̧u�`M�����ixV���t�7Ҡ6��k�{ 4��ݞ\d�"FC���A�����|��M1xPԘ����T�m�4�������+�L񶧕<t'4R�j���'b�;��L�+X�!�U&�i�V6T<��s���<�1I����Yq�����ũ	%s�ڣ&H'~�\���������L��n��%��Z:,����d?��l@Ȟ�5�X3<�CF�ӑ�]K�2X�(DhB���z��� J)18�����	���2-�O"��N��e0�b��2=��6��ȇ���jɕ�1Gi��K�g�ڈ�
d�D �����-QJ�z�BȂ�|���jܕ�0���Q�t_V/�_�^�è_�̅����&���:�K5���znYZ�e���U�vp|�^-@����`L�&-v��}�	�]Q�NSg���Qz˙]5��v{�B�S���I�Lk5v%��,���R;�V}�{���.{ə��P^��[ik���w��ɲ�R0�k��R�&BȾ��|�8�*(P��e��*���������`�m��A?a �������{�-�8�
����d4G�������֤�(�I���vS��I��Yޭ�d���}�t58�6���i�/�������YJ�D��[B�Ӿ�8*U����1J�Z �H��Nw������Eg�Z �r�#X~%eB.W�/��:.�M��w:�;��4�p0*���##��H���PtB��N���gHw��u�L���+f��a[7�z����9&�}Ź�-ׇ���4�I�"�{R%��Û)����5�3��{i��x�w&qk[���x7������ٗ柨�&O��/9��������2�[)˞�90J���e�ݎ��yH��D�'1!�@<��ʥhXJ���/����Ζ6x�{ݐ���ӧ��1��E��3�K�<�*x��v6C$���9w2��z35�#*��X5�D�
���r�u����v�K�0 ��LY[>8�-��A�D�l�`�;�>%�v�O��De#�5�ԮZ�?.�D�ϚpV�L,�^���<���Mjxo�b@��zn2��v-�Qx�fb�JA|��^��M��M��� �� �,N�[\Z��9�F2��x�H R�֗��ua��z[d����2���&Z�]��޲0��,I�G��W�]5�kJ���>����}�)��G���M?�DP�}pe-��}ęTK"õ��H�zi��w�uY�Q��XV��Z���qh2�r�?�7����}#A0/���O��g�&�`x�-ȭ���&�&*��r���L�u����H�>�w�M�M�t�,�R������7&�S3���Ŷ���'�#�a\�c|��(BzM{6Z��6�xM��!C�RB�����j�6tZU/C�e���>g�4v1��Х1����p�HDnt������jCh�������z,�@�����?	E\��v;/�np�׫m�(�w"O�-[
M�@�����@v`q��GN�����k��fD��I-!���D?5^�`�"!�N�i>�:VCHW1���"���60�H�/�K�FK��%���:ٕ�y�Ϳ��?�6�G1��k�Q��맼�;�0��sS�8�s�\>�}�,�a���5�`������nx���OF�Ll&N��5M,G����k#$�^�؛��%�D z�}O��ƃbO)�c���ڧ	���DV�	����3�f��(��i����&B�JP� .pIdA'IpM�Vُ�	���o�*O�>`�Vjxh`F*so�\׿I���78J�O�ǿ�[�aT��]�啒���:����^��B���~���`x���jH��U�r�cw��?���O��Z����Hg���}��{���3��]H;@�~�0����tT��#��+$%�)��r����X�?����FrU4* Kwt �� ���;U'��?L�9I2j��5,�
@�B�t����;,2�ga���FES���UZw:�΃� 7�뮒�͙Y7}��iR��f�6����i��~p�z������W[w�$����l�8$�o>W����c�i�����pb�i]w� ��P�!F���06q;3� ��O��kԐ3����05f�D���*�њ�N�b�3�>�3�K��$��y�ĈT�k��ʬ���*�͕��=��ꈉZ
�:��~
6�$�
���ї��m^��W����v�K��ͳ YyN,�8����LC��<�m��u��E�������$�p�.��f�44��ߋ�*���f��ޘ%Ѭnh��I~P�i�G�Ӑ������se��
���4g#�����63VI���ΐ_��H�ܤ^������)C��!{��������ж��NW�ė��.DC�?y|Z= p��	p[��V�>L2o�s�x��
��a
A��Г�%O��_�(�4�}&&G�벵�#&́z}��t�F%�;}�hz(��
Czj̄8FΞ���b����9��(+�U�NAN���ͤ����x\��2GU�L���_Y�_`���G֭�B��n�I݃?�^Ӻ���>ny�l�g��z��A;9\N�qO
ZU7��ݝ(9�MW��i?���3دbE^59K�U��>�A{�F��C$�cc<��uK[�/��a�p䧭~k���<<����zw)=s\���桏
��$�&;�5"�ėP����J�)��Fw����5�ܿ�Kް��Դ]ɚ_��ۯ���t�Qf6���n�����YU�cL+�|A!���M�3O&qXM�U�%�7��Y���iK9�]���ԓ�MD=Dr\k��SL�V^3�}ų�@tJ� �c�&�mɀ�0����S	^-Tj��>b��e�<ܝcû��a�0�4����%��9���a��S�I.9��g9��Mk�@MaJEUC���"�BS|��L��[^S�j���f`&lÆݨ7���G���>,���p�is� p�WL�Ȱ�`4�Z��c�1���n���5���O�������.U#��Y��n�!h���ե�H��%�Z��d�6�ڼ([{]!���&R���@N�i���������{��>֏A��`��@���$U�B1p�y=ҭ��卛�U`P~zRާ�gom��pTAQdŦ�X�oC���9(c�.0:\��׮ſ]������ub�7��c�ivaɻ���s��e�|m߫ݞ;:KS͐M��$��J��jP�X����3�{�2��9����p��4��������:E#1���0�w�1����Tݢ�o8�<]�B� �Y�$�n<��@�gat�~&2������e����f�o]�	��� �:�B���k�ׁ�&��Dp���2
s�I���y��j�92~h�B�"d����{o3r�"��"������4��b ���\���:�v{F�MO�$���o�i{�[`�^�\��H���h���,��zf
�Y.(�����1�G�*�{r���(��I2��k���l!u:AATs➲���v6�UPj�&�^F>SQ,�@�����"�;q.`��Q&�k�ka���h��8�ܜ9���ǃ�e����@�N����\�f����C��X,��ZD�:_���e�Uo!dJ��L5Ɵ�8����9��M�L�|��Ų�|�32��W�l���`�h��Ո9�W��d]����Ѩ�~T75N������Vts?&t%p>chK�B�u��ߧH���v�V��e�~z�X!�QÕyxG�z��|<o4��ȉɾu���wF��q�s!BY���vo���GY;dV rq˳�p���3�PIڙ�(�|Up\O�����n+�IF�]#4Y&B�:z$�7]q��#ܟ����~��+S\k�42a1���V��W��3r�\R�\Mz���Y���SE�Ģi�`����=��^�+ҥ�VWz`h�V�N<Xd.V��H:��������pƦZF���-��'X�`fM�����?q�f���.�Н��an� ݟ���7C�;��ۭ�1ëߣ��2�Y�z�2I��Z����C&U@3����Hص�@���+ �&��$��'=�\��c�z�5��x���&���,���ܟ�@�P�$+LXk%Q����q��t��6G	"�f�N�`Y ��}�*KX3��)ǯ�e��O���!ǟ�g?mK�[@��;�A�d��uƼE��^�z(B�6� ���Q����A����9��z����2,1_�+΃����W��VK�?�籛y�"H8܂�~��O�#)�R���v"�4��KOiQ°?K%׮���W�6��
ml���.!`��n�H�3��WZ���E\��#Ƃ���R��e�6�8��8D��uM)u7 ����ܥ���M㨭�*3#	��F�|`@��K*��i����'k���ŔG�I�����p�*x�v�����KS���qzۋZ&�:���q��^�I�(��y�t6��J!C/�'�h��Q� �����D� U}�w@�7s�\�����xJ71�$�{��K�wI�)��n�W�Ek'����1���ڜ�mS�>�g��|��H%�ȭ�-��ݒ8�԰��u'���$@�QZhڶw��
 ��ƚ�X�ǰ\.��ˬx�!:�$�h�p��X�F�K�������'�l4���K=�-:l�L����f;;� �A�v�A/�-�tX��}XQRbߘ�N��\�:�Ŏ�����1���
+�w�^g�8o�P�46��E���7�{Z��=���N���ӛc�J�w/�mxR�F_�/��5*��7�ȝ3D��=\ D �%v;-�7���$-�yĩ q��37U	j�z>�Rf�vۍv3.)�&M�a�y��X՝�����G�M,3,�44��"�n�!�ZB���vYE�+���K��,��D�e��@�͗�C��m�Qh@`F�k����53�'��␚�Ws��Ɯx����O����VF�)���s=��;T�p�n�0hek��p;�_	�������J%wd�/ފ(�帕���n�\���
�{_\\�*��n�m�RwV�o��C�QM1�����X\�֣v�=��9f�b(��|����a���E��}�6���a��nT�%����3���-�ܧQmW+m���-W�����s6?y�V�{_`)< :p�0q��`çQ��|�ٮQ�楱9��"-	�۲���_R`��;�
��?r3���lg�j��K��Ժ�� 6�>O�?���	-=���L5I�%�`�[��6���|㴲��C�� ���AU.t��վ�c
�!p�qx�g�mϫ�SdJ�:�aV�����Ugb�!�a�)w�-���z�g�M�	�?%.�I��vc�	�{���5��x�Uv:�J9^�8Dɪ�� �xE	e%��U�jk&��MT�Z�s��aF^R,kӮ�^�O
*ϒa��WG�X`�~�cd����h����ߐ�g}��%�JJ1~֧!�y��m��G�H��ø�f��ّKSe��Saꥠt���*��lw��T��d&!�0�Y'��ؚ�3�p����z�.��AXn���@��:ɂ�0V]���d<Y������T)I�l݂=�4}�tס��C�)�$#�IMGük���{�55���#��ZݨD|�K�]^�I^Lռ���ip}��k�D� X��ӧA	�1���mQ��V#\x���B�!�|��T>5}
������B���rVg�}�v1�tS���r?�5'޴.9`��rċR�0�fo�n�:���7�	Ξ��H_�P���VoP�'���z��# 1����P�&���s10UE8���U&����"�#'����4��Ӑ�f���o��YKC��{�_��o�\��d3���_��s�>�m0��c�p��ކz� 
���և���F;-(ׄH�$���������Ԛ��g�Ft�%Z��B{�6��ǆ�a
躷:'����<S9�Dص}>YJ����$G��	����Hi�9��^ENz�9�=�����x�Y��:1."��df�ņ��cE;��D^K��h�����$���$oޣ�`�:L9�=�qη����E��,�C�`���_ob",����v�{�×��y�G�r	(�� �I\]p̾�w���Ѹ��.��B�<�v��.�;��zK@�㣙LGȴH!����]���^?G!�>ߩ���y����<ɝh��'�OU�N!}��p�2B��9Qu����!iW̨�jk�~0��W��	X�h�$��[��f~<�����n� s��pd�@;u���r�̶q�o���J"���j����F2V���q�i���Rd^e�+����߾'j��v��\�փ����o�*�O��Q��^51�]���`��S3!_L/ қb�!��z{�^a��τ ��_��Zp�i�N���(o\�+[��Y��������h�dLٸ]e^Ԃ9�x˶&~r�i[�u�ܹ+9��l~fz^�����p�ħ2'�FW�{�*����P��7)�n��v���,a^���ɌS9ɎD%��ٚ �i9@�A�1^8RW7�2��Y���.���*����+=��U�AYi�f	�m���8_��Z�[�Yp�z)�%�7����j�ш���<�=�������TUK��j��Ą�[L�/��Ժ�j���	NSTR��3�CJ���L��t��|0�[7��+���G��E9����]���ׯnV��d4�i�wufq\{�~��T��1�Z�f�?�h	;AUz�F�68��n��~�s���"n����G�e�v/�^�v��`�V0�W#5�2�EL�tR8C��!g:��X�^�[�q�u�ׁE棿6�z8%��ѹ�����u��K�r�2倂�r��MN�bK�`��IJ�S8�)QH;�;�ƷN��]?���ŎaP�L٦HԌ��Tӿ�4ե�RB��fy����&4<�3��u�X�{�T�))��;r9�z�����s�l�.�۲�8ט|���@�~0*4ıb}���5�lr�#{�1l4�Jk�
���&�hk�ۈ���h�������,RX:iy�l�mŬ/B����ȼ��ɐ�vҔ&�ХCo�>�7d�9�^�����E��ӎ��zu�t#)M�Z��T��Ϛ�A�҅)����	]�>�"��-]Ec��eO��d����4G�鱞�	����.��4�m	�ea�o��jE��������H�����_P.a�{�z���,H<R	�k�/�a3��� ���4Տ-i�����p�B����VqG��lN��P���#K�&������#�� y_V5�����䪪E����rR��좗��L�L�ˁ�X9-�Ëx���+$m�`�O��0�����J\�t*X=����ʔc���<�'ہB�Ӈ��^�g�_!n(�f� ��/L�3� �e�_��R��R��e(�s˩ֻ���Ө��;�˪ ��ɻ��FXj����~ߟ\���w1�֘j�jzm� Fs>���}~�64�V�|F?db�+�������b�K�0f�V�P�]�kLM��(��ޮ�ݹ��U	�P���d�@��C"E!�Fg���lH��ҝ�a�����o\���Ғ�a��@��=ĽE	LG�T�e�ne��޹�aǲD_�̶�uy�,���'[�[	��P�;�8����U����i]L#;��e6B�YuЫ�F��n�8�T�
�6�Ժ %�C�h�(��c��W8��n�fE��}~��JT�Ӏ��zQs������2�mz<y�l�=�c����#4_�5�+��	��ƞ�k�r�������1hB,�m�ʉ���+�~W3Һ����Q;u�'\�S����x]5+������wd�TdW�1T?3�a�A�lL�T����2(t*�����OB;M{���y���Z�s��H6ٯ�U(s;�ҡ�˔`)̀S�Y�P�8���AB{8?d�`�b�6�I��K� �1���V�0�N^e{�v�t�}�����	�b�dA(�n��&���)E��4Y�����êF�*���~�+����a.���c\��RZZ�5u3Z�$+
��H����I$Aj��S������u֜(\�C���D���k�?�fQVͿ*�a]����G(�8:�ߤD�_=���p��m �+�Z��n�j��a����q��g�=ó8SGs�����n��k,]��v��^�P��єM51��I��돠��`ޏ�[)F*�[�DB���"u&��I~�o��y�IF�����WFE�zr��FoS���W��}i�
M��R�Ӌ n����Bɳ�w?��
P�������"��'�"�)��6�捧Z/��0�99���	Aa�_��G!x�'���F
�Ȗ���}����]䋻�(��.�۲�����'�wysDL �/D��S�\ �ڰw�U���������	D}C0Y5������ק�*]x��qw�q�KeM�jW>J
�ZN�Z��=⤃>1ғ��Ћ�Bz7WLb��D���-:^�"��>��R�B����H*B<؉p)gD���@צ'�{��s�󑓺�|�(qMa)u?,�P3��|��ȑ�,���pҊ�@�8�V1�a����=b텿޽�j]���o������$�W<�������G�]]a�ѱ��'���+V�y+�K��ǀ5D�BX��D'�b��i���߭����(f�U7�d�V���Ђ���~���~�	�J�}#�こ8fT`<� \���SjG.��z���i"��:�&���ڎK���/e�U�}=�NkKJ����-#��A�~�4�/5���z��^�۔?>h���]���n�mk�F��0��$�@�X8�70����e� ��C�c"I����T �eIx�|o�H�S��(�ߋ��HY
��:�:f��U�����(s��;�	3Wo�lMy�^�ξ�FĊ�uI���4�DyS?�a��
T^N8 | �ere��������0���;�l�a$�րY���l�%����#o�?l��.�=�΃C�X�s��@I���8��H�������U(o0�P&5⩜6��R#/��S���7X��I!���+�8|ΐ��+S:M�;����(��?���s���t�#���s9ٱ����+Y���78�]��sk�PM���RA
�8=n~��͟lof��k�A���J���)W��q?b��u�B�V-ڋ���W��Daj8�a��%�*�S��݊�B��sy �&j�=gC����${=�k��5���V��Q��n2�
~�q�%����å4�PA6�@����`w��d yl��fod��7�I	4�`O}Q�ͪ{�{��&������M5���,'݇�H����La^W=^�fvMgfo��N����B���r�ڴF�G�K�C��-��R�1p.��:J��bD��4�iŴ���)p}W�.�O� �\*@U6�r�����d�4N��;�Jq*=�)~����"p_m���u�Jr�6��>�h�<�>������f��J�-a���ߊ�a9#R�@�ռm5��"����k����~���G��h�EDg�{)����=��jךa���x;_#+m9�����4�s^���=�;G⫠�d~��r��p��������^!<]�}!z�K��M�~��={���F|w�X��l+��%ʶ;�l�^�&B�#"�HX5�-&��2,�����vVHU���WI���g(���*\9���&�:	�b��"���$�D�*5y�t��X��	�؉�T�x?���m�x�6[)	=�c��D��ը����=p��0�↌3B-v
=Q]��ud���L���8��J�A�^���:2�?��@�MN? ��4=��{㧩AL���SA�s���7Y�H�7[L԰��)�UDr����̸�Z����0Aږ�'�������ss�z�A�ڻL��d��&�+�9�n�s?�׫��@�ŭ��;U�4�7�G�,�h9p���#�/.R�;k�S�Rz1�F/�%� ����89���
�f�$�ؒ+�歴����2\��&�wΒE��S�P�$e7�ѡ)`�=h�!�(�"��� �r�`�
�SߑE�D���&R,	�k�<P���H3B�F���_v[K_ ՙx<�\��΍Shj�4���ר�K7�D��0�R vx�=$�o+}Z&��`[՜L��22� �Y��:��{��L��D)��Y�����A`�S+#����ʙ���H�[1�?=�mx�"�-G�;�o�$��Y\�.3��/qk��B�#�",6�5���a���R:��8��R�9}b��<��pO�a��#�����z��I|Ԓ6�m�ņ�J��+x~� 	B�/�w�J��@�_P���5���A�#�"��ۦlԼ��M%<wq�ۂ*/��i��=�Ey�;o�I�\Q���c
=��:*�>Q!�wrD��)/�A�݊�o��T�(1td�/�sa�$U�p=�4ߣH�J�H=��}�F�� �l�[�y�8_*�eρ4��������đ5PK����2����r�Lx�(����}A˭��cҘ���s�������J�c�v�����#�K���y�W�0�?I�!KG�\���������)E9�rj�7�0ɱm��Xw�0�RY�2��k���gc�C�K&^�f�3'�H�]��([t��^�Q;Y(!�t�-�!�w��ҵݙ�k4�B�z&��@��^.�رa-�TjU<{��lA�{�"�:��$f���Q֎ÑPt^_������9#����pc��V�$��B�����V�����Ţ�%�:�)@� �f0F��H�6]����k�"��?0Ӟ^��M\ʣW����B5����msN�sݖ�alD��(�
w������9q%�w�wA����Q�,��Ӡt�qjHg�͘����d�0������� �cvs:�*���E��7��^�z��0�(D�aE�bI,ut�BP����u���wUf�@9*.p����8F���#I2�(T���{��g�fj��2SCl��,�;���T�%!͈1��\Xhq)��P�"\u���m;n�OT��z;�������(�e�x=�{�WL�~:-��I�߀����G�4��ۮ:�W�SSǄ�s�$S '��0RT�d?�Fq=T�T[���sU0�?����G;���gq�AB}���Z�*���}l����7t\G���g>2���$��5�hc�$u���M��:^��.M��� ������b�by<KG�؏wkH!�su����s�_p[�ʵ�PBjYr��n���:v�qO�����MσT�P����U�Ƣ���7����+M�徟�)�L�G�G��a^��0=X�H�	y��Ĉ������/v&�&Hd��#�:��Qlc�t���4N����o����r�WTiS�W���������n:�acO9
�Q������gc���}�`�[��ܶ~��M��î��>N��uyeY�5�+����.`�CJ�:π�侻���3�h/�������#eu���.�͛���}aӷ�SZ�,�~�T��2v����*�&m!���ʼL�C.J�C�\� 	�����}���2Jc��Z�#�m���S��;]�_ �r<�4��?�j���q-m	'r��n	�xT�5��`���-�����Bsrbx�1�E���ݪ#4����ʮ�kkGЊ�����z�6I[�)Mo�A	�I�=;}��,N4�A ^����[�K�Z�a��t/�B7>�E�E���iNj&)� ���X�W��
�4:M�y��yV	6W�= 2
wH~���t�'�޻R��m���H �����H�!�`�0�x/�e~���6��Za�_z8�19p߫j�_���+�S�:l��t���������߻��uQ�mǅRJ�cЎP=񱳷��zpVz�-�2J���#�g%hY/��Z�*A5 �-r�Vua%�e4.E�C`�����1h{��$�����%]0�P��y�bCH������'d����F��@EH���bʳHu ���27c�,�uݣ3����x]#�_����N�0�L�'�g���2�qSSf,�߱meVL�Y����N��5��f�B2��T#ܡ|q�0ǢOΠso[)Ɵ`����J�;R%O��k���)f�I$��Keo��s<��^�l�/!�\Ӄ�d�x�َD�L-hJ�NA�Φʽ�A+��@�:L�(yd�ד�&�f����1 =�U�T�X�`N_�#
��R�T�Z}�u��y����y#����:��ʡ�����V�[�u%�/D��W�˥*�Q�0�7����c���-��� ����,�G�Gf$ba݃zP���M�T��ґ�ӻ:���!L�ۺ���"g��˒��?���LG�,X_P"q=L�̾k��YO�r�S��ۤ�o�6���x[��]��������
5~V��5w;2��j��� d�<;�fM�� ��DGն��t�][�v��t0�$?��偅"[����������)ќԅ=|{�=��颷�[��{��B�Y��5�y���5��2,��ɿ��
'ծ��4d�Z����1�4jHJH����*�S�����{�E���0�k����Q�k��&����8���!hi�m�?�������R�([���}c���Dp�N F��&Kv�HQ�E�/"&�>	 ȝ?~��o(���Ӿf��+TRg�l��0ջ�]��n�h��N�rI���0y���1A��X�ul�o�
�gĽ��G�q�y`#g�\���i��o���#�SM4��I@����<B�����?�>ҡ��gTd��XpbN�}��y�B9��w!@ �̙��@��wFj=?gE����?d�(���6��um�"���>J�E�C�|�m�n���Xw�t6C�T��L�h�'zk����2��uڀ�u��AsPMS��;#4�y�F��g} ��C�Q����S��D
�'*?tL���.X����[&���>�0`��{y�D��,�q�gu�b�ԼD��r��OJ��- �9X-t��{g�)�9{g�]=p�E4&ޫg�d�i��Z�#I�PxJ�����kי��O�n+�s`��|������g��B�4lS ����K��?�Ce����R�`�r���y���`��� î۔ł#ˌ�?�A)���(G� ��؈#E���c(>C�Z.�O�[�#���(�0
�^��ǲ�"��1�)A�L�!�\N2I���,rOf�����^��Am�F��ci�һUr�'�ˆ��ע~����
�W����8��0�]D=�x%��N���\ƈ��MZ!87�\RK甖�|�~LI��=R7���y�Tc.�=[�NPU�:Z讧0�Q)/������F��寗/B���l>�_�"�s��I>N_0���P� c�Ȼ��!K����'��z/|�(����8/M`�^(c�=����ǌw�����膫-q��	���[J=����X�8���_��U*:�Jy�VД�r��;��,o;�2��G�W�"�d�6M�3��_���8e�L�{��"E���=�w
�#�B���[��4�;7^;�T��fL�;CK=^������9t���o|�3dI�2a��bO�T�c�'�N/m�w�S��sYRNBΫl2vy���:P�eh���M��U���]���c�y��2�ܵ,��o���wƉ�d@!-Y-$�uU?{���m���c"u��ptz�Xz����nov?��X�9���j2�@r�}�S+�>���F�����#�?�tc�Z��<~�O��X��{�b�a�Ժ�s�5�����[��γ�i�������Nh�������]�s������wv��*��䠣R�/����#t�_{�`�h�2�����c��'�pL,�
vj�{qL:�[���8����.�_����MR���l;�m��^��=Q&�W�|ا%b� wj<Eտ�1��#"�c��J�r�`|g�h�)�t���`Ĕ$���P���L�=M�#;ݷ�6DLR����uhTb�G�ppd��O"3V|A��yn�e�X������퐏�,��{ H쨉��xvz�Ý����lA^PK-'�öx��ƿ����,�^��4�G���Q�U���HHc�VpMnJ�����8�IY'߬}�~�K��8� �T.>Жl�i����b7��YbK
p1�נ�`����Ӑ���ɔp��"q��?y��R�2FA�ㄼ��)��W,�9�=���NŶn���jpdM9aC/��[�|�1'�a��(���4����<-f�{f��*��&�7
�tZ���
����Pj�@)h�p��0I_*I��~�zDfs*���,��e9��C��?�Rա��л�yC�;��{�Nsn���X�-�?_��x�C��o��-oLH�Hx�x��v��x1eT��7=�?aT�-����::�wߢSW6b��"���8F8��(-�؀�P�f�����S�w�ty�)�9��b%m��(��2�_��5����=�?&�`��`�3^�+~���@����y��&ǝ�`�_����$.�R��qJ�{���&��$(���l�W릛��Ʈw���Sh�ՈVj�H�<����_ǈ�:F7���C�^r%�X�ٿ&_�4d}mz���%��ư�0`�n�`��C̝h�Cb��O�%꣯�{H5,���AB���Z��}3�ϯ�|S_�&��Y�j`
�/5�����/��Q!�$�M/q�;άW^m'�� ��Ȩ9�.f�BM}U�n�L?{bLv�yϘ���#��}��W{�R��e���Ro7�����U��oMH�N� ��=:��M��v�V�bݔ}�5GhØ�^�hH8 f���"�G�H#K*�m�Rhۻ�'�1[ܪ@�Z�#/�R��7fC�m㨢b��*�j��*��%�m!8�t��J��N�N5��[@ہ�4�T�:HP�FiǞ4J���jC�3���X(0j�觹�|�1F~֤�y�����^����[7������[q�1k�$[���(dA�D�J�Wj��Z�P]w�^�������#�V	�n�^f}��HA�_�����V�s���	�Zg�E����
7[�Gp(��'��JUd4o�����(���te��h=<����U�l�m��JB��@�pq�g����A����H�"�rz<bF�ܓ�����r��(cQ���H�E	��~��:��)n�َ���	�l�DS�n.jF�Y��C�?r�RB�4�<�@\�1��ݴ��*���R�q*r��R����'�)�����0�vL^̫:99Y>v���IC�pjzh����d�s���5��,�/A��)����� ka��/S$�t�-�>�Ȧ^����hS|@��W>L9P#�l����#��Hۘ����Vp�N�_4��cgM�c�|��=a���^$_א8�Z�5�Pn��oM4�>�pz+U&�9���-�����jJX�,��E������A���޻�sv��EA`p5�~5��+�N��:D��a��XԠS�!�$J��� a�i�HP���#����1����z6����^ɤ�s	�{��2�^�����;�R�Y~em{9<z!�ʳY
4pKK���"Xco��.RK�-�n�l��3��0� $B�bV�`�7^D�[�5�*��y�Y\�0f����^2�(�0{/$�TER�+�����I�� ��bSm7j�f'��W��A�]kb�݉yf*�Ҧ����<�F�Q��/���d�29y�eU�I�J���x��[�jzd�@���� 8ā��d�@���-Q�	�"��y�p�n��Y��t?�s���Q7����%�ؽxz�`78��/�e�ue�v`� R�;GO�CĘ����i�R��ئ��T�8�a�7�9Lq�×��4� \P�f���[8���'<=����B�j����� 8�����D�%���x�(Aidx^��^�]�I�!����ﶱ�ލS��HˡA�!�ӣ��Nj~^�@���)�a�qU��5��Ė� ⻨eE�g`}�-�x�_ ą�O]�K���e�{�<���7�~�W�������u�!~�!s(Go��XJ�$i��'�6�[,�MX�J�S��x2U/��v���fT	1�qN�돥� l��~dw����H`OY�+
���е�5�_l1�V�	cjٵ	��6�粃��:ϽbȔ$��2��!Z���a?�RF�V4�A�~?}>�;�7�(�P�]�-�����#3O **��r�H��D����X�+��z6��)�	n�����(�p.�|��)�j����8�Vr�&�d������Lwa�TU�~_P���k+8[��T��t>�u�3�g3�B�/"]���Zxq#b�]�i��X���1���o�w�)���'=�B��]1hb��3����	���J�!�3~]��M����Og/I-'�P�2I�������q��b`s�4p�%�p��D#~����$�.�U�m��*O��A뺨~�?��=��)=�dߺ��>���m1�Qn*G������n$���.�p��Sj�Ƨ��6��.[�`g�:�2���������~�9�w3�2<�pk��ϕ�0�p���兴��7�!��3�ז~�WĆC���3U�Z˘%*����4���zb�����}{vUw��
�?��� +��y��C
�	��d���c�{�؍�%<�{#�a��PW��\x8\X��1Ϝ�1�71���Y�ȩ�3ڃ-ȓ9����!c�~�ٝ�����/=�o%�Ǽ�͛Q����R�uW���x��{ut�V�"�΅�a�,�"j�#Sc�U�N�A��� �`;�dz���Ԭ¹����B��P��_	1{02��A���$�>�7^��.
�}P���F��aآ5�OlR.��Ʌv���̖��ZG"���^��w��e�B6v�?I1�^��\D���'��8���y���� 4@>�Au�_�H!Ը��<>Bz�I�b�&���u:G���|���9b�mJ��� W(��_d�w,S^��'����~/UYBj�nls�TY�e��ߑa}��ɪ�nȯ�
~:�p�QJkVh��`�h�O4S�uz5�����5yty�\ݿ�>�.���MB����̋��Z�۱��p�v|$����}R$��ڻ¢��3�#����{��W��R�7�������*�n#g7���6T%}�$i�D�q�MqM�֢h�Eq��z��5�7��g�ؗšSb�t S����3��\=+��u��]��{�2q/�1&�}]`Di��==K%�/��TY�/���M�Z!<�!@��п����	�[�mՇ��.�i�����i��Zt����������]�����sl�[�@����Y"98�x�qhxse��
��bÅ��Re���	"�տ\
R ���>h��N8��vXU��E�B����qaՍ�6�V�A;�r�����*o�q=|8(v��Lp�`�d�
>	;ʖlb��ٝ��U�Ug�	�,B�0�d��dF^���Nptxe�Îm��,�P���,\�;�{Q�p_�B_]oe����q�~��>a]s�C�4����ʘU+�켸2#�DSsQ�j��S���EW���W�Oc�'B|���㔑��a_��cO};�=#���y�_-Ae!'^	�d�k6�VE@(m	�;X_��Dy�J:��7bqׁm޻$gJz��}�{�V�:�D�������2���5u;I����� �RQu�/	�?ڐQ-%�҇5o�h͔�*�k<�n�����`�/}���-ʘ��I�A���0?>�/-���^��������!�f�5�,D��*k����z�?)��Ӳ�#�d8�9��}t~	��1vD������pZ��p�*{YA��T�V�C�����-w�e_��z3!��tzl��}�<�_�tz�� "ch'Ԓ���A��F(�Β�c^�O�c �.0��H�x]@Ȧ�L�)|�!��;y�q ��^n�>G$�o��$�
T]+��S�!nv��;ض�$@/N�
`�$�B��f���]I}���V���5{�r�@����&/�J�G"��v���|H���\��3����e�tV�|{(%6#��	�@�"H�"��>�q��O�Fn�Pt����s`��I�f��`��t���ʉ���ͪd�M�]m���dΏ/=�?@=��L?��qS�a���©6�i!�mj[�2H�2k4��\��U���&~�~���Ju�����`�(-���l:,b}1P�o8m�:�+%*'���
MHrh^a��_������k 	��R���,��[�����h}��0�(z����ޥ˯S�A1�6AzA�r~�A�i��/���/�Y�@'s�>���+Si9>��'��Q)�Ӝ�pW�SG>��9��F'9e��*ѫ���,3)[�5���4�Ő�0�
��O�v�����,�U���g��ݤv&������C�>��}g���%?�{N�w*R-ig�<?C����/X��G��I��[�D������)��z��Y�+�j�x�hB��Sps!y:C����K������Z�+j���/���p�j�������/ڌ������8���8P&k��4��Dg�⬓E��fxX̨<��� ��s:V��N�(�Å���v[��v�X/��^ZF�D� `�*�ۄ��L��V��xi$s�亹�B�*�V�Sa����/7��z���(?� �ؠ�G�@�ʾ�F4����BpqIH>?�%r������9e�j�5�ߓc@��~�{2yI9s����P��Q�'�NQ�$B?�5�P�0�	��jS��n@FL��$�^����n담��_�.ߖh��M���/�Vm@�79�7�!�R�ro�\�[�Q٘��OpQ���U�1d��浈�7���)L@s|򷥬C�ܣ�U>��g�2�̟hfq	��g(f{�N���L��4�_����Z��w�A����3�y_��p�3� ���A����-��1����1��b8Ov�K��Ʋh$�t��3�����ʮ�)I6�Dg���$z;T��e�����(�Zl�5�{��c/�<�����~�������_'��q����.&�U�W9��DY�A^-���j+���X]��`H�6�S��n/������(M1�"^���A8`Vz�<���@�\u�o9���6����\��A|xsj$Ij՝n	�<���jY���zC`$̃�^������.��V��:�d��ϴIc�)����\Mr�F�㉅\���E>�^1&R�(��qe�+�_�~�g7��wp�h���3�W	���H[Zp����|V��Tq>'� �XT�i��+:?=��래>��k+o ������&���k�,���$���o�B���-bCZ�V������S����I���ҨdvR@-�-�ƞ�T�rD��c��}C��a�eR��'��t?�t�J<�̯b��+�qp�ǋ�r$�.m!���߭�Nt����?�����8e�.y��A:'�oO�T�(b�����?|%,NM$F��B�a��PN�S�0Y}5t����rj��{�0ܹP"�PN���6�� ��Xw��^��G ���_\���x�~��Ҕr=�@R�m<���c/}������C����v�ubtj>q��J�����:��~͞�u�7���2C��c�X�fI-zrWU����4�v&�`o��4��}�`�Jq��O=�k%Ds=E���Gc<="��"��0;��x�?�O'�R�`O�!վj��.��}(�z�,w��b�9��g[���*�ҿr*:��9gY�)Z�a(O|e�Y����:�wW=2� T�w=3����{F���8k���Gs-�0l!|s�af 7�l��Cs>��T!l�n�S�MK�!����g��Og>,%�ϩ���M#�O�ٷ�5M�x��t�tlb�k�|~���g���*{O��=I���%S��#A"��D���p[�4_�	9m,80X��=s,�Y�܁�,��<�`�n�K��%Sf����jZ)���V��֐��.���W��P���K�9�p������Fc�9ũ]M�D��7�:�Z,L�W.����zU�KsN(m�om	�t�f/5]�����$"���[��F�'��RE�/J��t�I��*�B��̆��lHm�}��X�}�$�$���8�e<�i��3Id��*v��ܹ��%C�U��l-Z�R��PH"�L��h�\���;<R����bL&����M��cN�R�o������W���WX�	��T2��C��BʋZ�/V�)u��1�@R1�`�-�taW�]a�Tk�E�_�� ��z��#��u)_�R�K&�Vw�,p�L��d٥��t ý�po}�!W�d����3[ڏ��e���̇l�����H���+�:V�|�[�f�4�x��OHU���V��3�8I�X�qs7�G�W��� �炝�o��A��S�67,c+_M#4#���d��8���<$�}	\�Y�����VR2��ײR�6g!O�V�?xH\a#mǾJW{�)fL�q�!R�;��e��;�A" ��<&2��~�1�X�z��|x|�Zo�0x!]g�!��sy�L���O	8��-(���t�{+̅2fUgEFp�=���4���j���"3�Rػ1��C,�\:8ݬw�3��V>���ˡ_EB���L���^?c϶S$�/�\F|Ѣt���[�Y���?��+��{!꼰�0�TQ�?G^�Q�u��D�c�/��,B���ZX�{�x1k� @/Sb�V~w�?5�([#�:�᫇$Gθĕ�>l��z�G��p�����"��^*�N�h�����tGE~k����� �KNݾ:��\�q�$j�KK�{S�;JJ��ˉ3!2��ս��ݸEm��?=����_��������n\�[f�n��Y�f�aK���{�k*�����_b� F�]�1��������Ȁڬ������0Qd�mH�Ǉ�)�>�aYg�)扶��_�%��KRu�Z��+`�jw�g���|6����8��D樑
���V��u?�e��}��+�۲�N���O�6�b9ko3E�&����?�3'�@ʴ��E���h7+��M��4.���=�TK�-E�6�D4F5�di��Z��h�2�3?�üU��'1%
�?uk�)�4�p�פ��,�܅Vm��*��x�X{kƷ\�%v�V��
f��E�����?G�:�h[K��B�o��o1���[�����
UY�k���s��ꩥI��t�o�
5v2�)����a���q��=&/���(�Pc#�_!�׸�+ 
+�+�����Bj�;F������ၮ�E���@����z,*T�V�X�z��nt��~��qtc>M��
-Jl�	/���g|�*%Ϟ��� :s���ӝ��;����?�M��t��Ęo�I�h&w��j	�S��@E�?�qz� �=~�եkm~o���O�K卑�����Wd;eP!:k�p��ȑ�Vآ�'�2Dm匵*~�/����7��'Κ��@�Rz�r,̱,ah��=����8 ��눱bv��omμ>��&�o����	ܞlv �<qN�Uw|ht7ɖ�e�~4���@���aE�Nڼ�1&��K����sTkY���{��T�Mӻ��|�c]o�S*4��>e���Td�GM��֝@/g<��ۻi:��
q�c���l��m�mƕJ�Taz�s�o S��Xf�4�i��#M�{�;��}W�]�S����%�p](���S��FӬ��+��3b��R;�o�ŀ��$�ZRwz������;4�V��D�L���B5����6����1����I@�𫖵Vj9X��Ɛ[�)�.��m��ಫ	�-RB��|.'��}����!]�9瞛+^e����lr���؇J*���޸��0�&�e/�e|���(��2:ڕ�Z��"Q��,�ڿ吁��{)�K�(�b�Z}[�#}�ɺ~���0`��G1H�	�p�JiC^�`��!��Y~+�����ͧZ��)1:�{�J#>���G5\A�I�A!��>^x�ۿǍo�C�^"�g��	�LU(3��E�S��D4#�)��E�r��8%,ӆ܉�=xx���-��%1�9K	�zp�[��.�?��I��tZhm���'��#gX��d��\�``���cj4�Ikn5a`z��Є0 ��:����J�m�b)�x�S�y�K���(��2h	L�LJ��x��|H^W�E�~�E���h0��v�86���!!�P7�D��|ϕ�AFOFA�Zm��j'ǫVd�ϓ~B �D�d�7��Zv�������	��qf����5t3��cw/;!�z%�Y4�ݺQbn^=�^�"2��a�_����i�Q����pqqJ\?��Xof<���E���p�H�Ʌ��A���#���i_�|��3�}�8}R6m��{Lh�0@W��3�"ЪtRO	�c���τs������'˱��������pV��h=�ӻ��3��i�`�0Bw��U3� 5�5�78�w�Wp�Eh���׸gh'}�-p���������o�ye�L#c��d���Ap���Q�c�i���I���)uv7�Nd)u}��Kj����is���)m@!K{l ˚U�jV�!�Y4Χg[�����I�B�t�5���(,x��n6�T�I��Ot�WQp������2�;�D�����؛_2�Ů��aB��oζ�n�&,V���x�=Dτ��1pÏ�]���
��n�X;��q
C�je0��ŝU�aM",���b�{,x��߳[�1���2�HO7H٣:����]���T�n͙����)�=	�v��S�%�[�)^6qJ���.���wɗ�ࡕn6}Z�DHt����o���-���==aWG�;k+��5��^hJ��M��¦�VV5�9���h�N��W�,λؽo��O~�˲N���eqk>�!��%�\_��C�~31��Xu�@�Ƌk��}�#�T�j�IZ�n����	���PhZ���h�"S�z�P)h}���{
\�����J�K��=d���� ����	�:���?��g��1�h>D�
g\B�P���@�6V!/��-��;�X�,��R:��W�����[(~��,��'�EO���L~�~a^���?�����f�X���"kR��0�t��)a�M7rY�0�����z�B�?Û�6��a
�p�\��WPj��s:߄\F�����̣jr�S�6l2I�����v��A�ê�Ƿ"b8����$Sc���+�'c�e�l̲��e��;�ͦ��u���=�f]kv��N�8&��E�JxXBs�ί*!b|R��\g��L ~�s?��� ?�U�a�ziwE�k�,\���m�����Ž5 <�h&���A�C�����F�aeNiW�8�"�N��V�NÂ�L��h��^�NB��Ѓ�;p��wv�t}�2d=�	�'��aw��hES
X�p�׏��c����K/�v��g�	���.ך��YӚ6�l��r�͂#�}�v���4)�◮'�Q�eJ�Q��n0?������S�{�jq~�Q%��T`nKop��f��橌\m@&�<����E5Wg����rw�[Ņ�q��4�:�j��jHh�1� ��]���lj�(!�~4�m��۱����m�g|OJ��b׌�c��eP>���#�w��A*fW��ZU�t���,-�ՅȂ�;Oo6V
�L�=B��n9�t�1A�����Y����;��Z��}Q�@M�I$~��m�I�:\ܭ&K����&A�=�(Cvl2����L� S'�ټ�:�����dX�3b��AI���G7��s���yɑ͠=��"�[��:�����V�K��D��[�_Ҩ&�FkN�	�` ��t�=�&�bj~ �\�S��6���nJ�>�@t"�	�vJ���[C���ޡ��j�.�U�Ǥ%�������me
x�����J��4y�cu��_30����a����#���Y���^��hj]n.�)�Z�̪B�]�Z�^ο��@h������8L��Ά?g�T��]՘ɇ��+�魓�H=��������ٌ���]x���\�����,����=�#�#Ik^7I:�M���~z=3-�j��w��������a�м�{4��哮���g1/=�hM4�`B�qa;M�}-�����ˌ����%,6J)�:��A�fI�uĽ0�r���I<�]�)���>�0{��rͽE�U8m�ʜ���'+ز�,L�>����P^fHf> ��2�,��$<�Յ�\l�Q��z��/�<�$[?%Ix�1>P)V��i�8@F�G?����z�C�r����7����B��=���8fu	k��OԢ_I���z���t?n����{j���Vq���eu�vM�L�6�h�xH�q$�.}`;��C!��xN,��|,q�<~�8�qɊNW���M�1q�QGҜǍ��)v�����l��*�͓�	V�qG ���v�uR!V�u�9�=Y��J�=�A�I��4l�AnA�P�G�ZV
�����Xj����.��@BG�LU9�l�e6*�#�A��&s �i�`R��A�������\�c����H4֦6g���=��g������u��a����5y	k�{�_�����/���ޕ����޹ᴀ"~\4����@W������n>_5��u4����3��M �voq�u�G�B�mf���6:� �MO��^R���)��Xы�|����I:��[�:�E+x�Z!a�Z�/��4�#P��o�c:Z%�Jk���g�>������P���۫���1�>��a�����q/4!d]%3����������/6S�Z15�~C_"C��;�0�]}��4��S����n�DL���q�[�l�] ��ʮ�"�K�OW���r���mU~Zlk3��g7v��@�2�	�>>��Q��Y���D�d�n�t�K��ٻܥ �Z9�����t�Ke����4
�p����3�mӱ�;X���f@�!�H�K�k�{�D��HG���	+D��1��Y��z���+�M�S�7�N�"��U�����]1xEuK<�M �WY�5�tfZ��v�,7(� =]z{HM"3���1I^�
p���`��/	 ��L��� q�ȳ0�����e��I�s#nn�`3\��Ӯ�S��9���.�Z>g��[�䴌X��Ǎ��2������5,��Y�[�S���#[�	��NL#\�;����IKd�´�;�^�+YgIo}$���	�H�2�]���3�@[�h�y:��#����C"�%�����߃H/U�B-�9�����9?������B-�vD�X6�J�',I�.[�Ƥ��`)҂�7F����I2���M}ҧ%��E r69�;V.t��s��~�3�B�5�'����a�*V8�;�1��u���?����?�ч
�&LJ�Sm�ʕ����	'~�պ�Qe��YP.6t��Yr�)kC3����=������GA^(���;�����[��W�d߷ʰ4���)���|r��,������?#5��q�dh� [�zq�yI���r�2�H7��CҰ��n|X�o���#���ܯ,��o�b9#���<�OU��b�)�~�u��Ca�|��S�m�O��!�97Ї���_�U���|-����K�Q,�1�p��?g�:>���<;ƹ ���PO�V��YF���;���������8n}��}XmFݪ�mn]��+�OWпQ�`���D?M�֤�=��SI"tH��Kh^��%Ӕ/-lF����J)�k����{l�7'�+� (t��Z��K��~��w@�.�9��U�[�b|o���_XO-+C_�A>��%ksg�2N���?��?�����kpϴ�����{ê���8L���gӱ�h[��}mB'Q����Q�EC�llmdP�M�V�z�1���f�u�^��` <P����AVZ@R�
����0�NC���7��T��>x�n�$�Ͷ�ƩBk��^1�!1<���a�B1���񞟑V�a�ۑ�E Q�
�T���iFU��Z��5��m#u��{{�r��[��0{�y���f�z8��J��{�z@�r�0Mr��"So�E[�$��I��ƣ�ͅ��R�PPҾfz��Υ� !��:YW�-(H'rT�᳓��j��h?F��%��|v�Y&Z��\~;�Ŷ'��`����t�#�<_V��Y�A� �Йr���&ʦ��ߒ�,�2��D�$�b��e��b��K=��[_R�1l�3"te.Hu��#C}R(L���znx�;m,dA�OPx
E�uO�V��SD12�'��l����;j�UK�m8�`�������I���d�˿�?C�e�u���Y��7xc|[8`����VR}�I�1�=��>����I���;�R�Ƴ����ܲv?6�2�*����?���̥Q��M<����!&�U7KX���т,f���۲_f~����������F^�H޵�zZ(J���޾?$����iS�+�Y�۵�Ͻ5��e�S���ݭ
:�:��y�����i�4�"ى/jzɬ1���ǐ+� i��N����l��Ɯ�>wa�qx��E���4;�.WK�;�n�!V�/f��И(S�K}Tcq�E�{�����hħm}�i#��N�+�/�Kл��͸pĺ�$��$�X�.�;���eԭ0%��"�uv?R��9������A����Vi����0�k�#��Td)�aH��'X�o���~����=  [Hxd���2�u\Mhh�!7=��pl�w-ǖ}Ĕ�䫐�H���7z�#�ee 9�m͗���&��X�y��Vj�\[8�Dg������#� �X��@����ብE%�(CM�1�N�NN��pG�u5q�dG�r̒U��x�|�~���6<��E?ք�¥H����EU���<��X��T~�׫��	������>a���3�#h�<�;]�Q���`�h>g�\2�+Z���F5O����Ɠ�P��T�]�&��b�yRR�װj���	j�gk�V�
2Zg#��ʀ�|�S���r<���B%���s��ë�w������,38����*��bp�l�������K>h#{.ɟ�2�0L�ߝ�;����C��x�B=ǫ"���-ͥ������"�B���� b��,ELfJ��w����-I����+�C�O��E�t�l���������G�)�u��!E����p{���N.���<I��k���[|���\~��T6���@F��pe�C{H^W+�L�%w�(���:>���(:;������>����j�z���E�a�78ww���5
�g�-�:��l�f�������\ڝ�l�b����k���'F.�I�bC����|�0W�5��ŷ�aL��寒�����M�Z��|sݷ�)���0@�Z;T*W�/a�3��9�T�q8M�}������x��ľ�{#k�éK_k�L5`&d��툆� ;?�q�ǫ�;�a� 5(7��� :d���Lecʖ�qe�	�xb0r$��8.|�7�Ň�s����
�����b��ɘ�Ԩ�����yq��!�E�M����?�.�@� YI�ݻ�R�W��M�N��G�1+I��+d=�5`8ȭ���XX0p�|Y�>&�!�韽汸砤�)"��K���p�E�1f�����L��z#�[�C�L}ڡG|�zb~ލ�������I
��#FG��A:z�G������;z��O��̙V6�X$���&�TK���=��e�S�Jm=x�7!aPS��i�q��`�[
"�� ��q�@��ZL򗫿�����a��F����BҔ�^�	��Gv/�T�+��k8*ZX+ӏʱ�K��@�����=�F��w�T�.:{�n��a��V���Z��R]�C%5��Ц�����%|�1�s�U�]�@�@��n�]OT������
Ҕ�������D��<���`�B{(��(O���q��O�.}�Np39L�8���@m'쏧@d�ۿ�&H��d>�6G��MLvp�H^�|��6��O��g��û��6�6ޓ�غ�n�8�`dU�}�bė1>Ҏ.�<���ŹT��k����r�����Rd�+(��{e�o[�"H�$�ZO��kON����Q�=������A�n�/J�o���Sy���_$ir[d���4J�+��|4�f5~����~�P,��\�p���EI�ڏ� �u�U�`��Ճ�M�G[���M��S�f��Ǐ�at�q������q��h5R?7�~�6>��yO��K��#|�6��,�I�YI!K�e�tf�K3�ɰ�!i�Pӥ���!l��6���P�����������|��@y���F�xɞ����`:�C�,��@��ސe$�Cǫ��F퟾��eˤfX*��e���K<���������`�/�����'���ˌ:�Z�)p���P�����F��;0�C�Y�TD��w��dg�ua����T��M������_#K����\���ڛ�`͢�ܕ�3����҆Ӥ@m������1��Sw	�Ԥ��@9��l�Jw�Q��No�{.��-��G�
3	�����s
̈L݋�p�)FY�^�CSÞ3�޴� �>�+�ȹ�=�A��8��G#PI�J���nQח\ ��Wx�?��̈́g��$�}�e�Z�Nb�94�EA��L�3Ia���	^��,�!�l�S�_G{V*�h/�1tQ�H���z��nH��՞9Vh�gZ��"g�-�ͻ��Ui��Sݵ���V��-uYc Jk���c��͠������^!#8���c"��a~X>mX�Kg�hc5N�]l�*p������6zU���OrK^���߱z ��Uť�fw�8��� J�\�ԫ���Ya�[^��!$��@�޳d�?��`7�D�`%n�Z� �̈́i�2�Ga�"<�"fy���5���#��थMc�wV[�,_|�tnf�(r�$�|�Ȭ������3�N��+E.�%ge����o�a�B��K:	���L�x� ��%��7tI����Η?9r�rb%Heoo�ϩ�x�ӡg)-76�y�ƍ<lE�թ}`�	$w	�������>�
���$�u�>��.5�f�y<�k��A��]εV� Ξa����$�H���	*k���Unڬ��{�[%��	�<C5I ��j=��z��x����"b��U�ڝ���TNUҰ�j��
ګi�&A�z{%5k�ܑʄJ�o���������Ib�����r�%y�t�h�u�;�<���,,B�{>�y~gR����7��t�a�r�ͳ-�����E}?��L�bW�@bʽ��	�Q5�d��G_����-ЮQ]-����	�I�5�U��>�m���[���(-z\���D�	u���U;�R��"��04Y����� q)<�x��J
[�x�q��Q��G`b&�� ��5���u�.���Pn(2h�J�3�Trz0����=���0�ғ*�S�(�?�Ui�A�^A�ɡ@`}G.���W*U+l.$��#�r
�|��F�냆fx���j��Q@���"�"L�ҷ�٪n�^�l�ЁR�z8[��؂��OK�]u&v��-��ۖ��*�©�5�u�ۘVr��?�1z��o��JM�lT
�ky
�~��8O��Y~W����8�[vm��J,��m���Z�.+k$��w��=d�r>[�Ǘ���n���Hfx������i��*cs^3��@?l�lw7��/�s��� �x����0�
��9^�U�X��IP�X�d�BT�&�'��%�`A��@���)�R��l��^��>-��@���z� �$�s�~h���UI�J5!}$'��>���:�	����#�,ÌW�,��O���|���K#@���7X�Yj�ۖ��^A��7'����_`�=2����~�Y�N*��^�d+��6l^�lM-�a�R�v�q�! ��@ql==>�����ɿD�$��a�T-�g���E����l��3R���W�g��xA�ӳ��ƶpO��L7ֺ��6Jr�L�WF�Kr�?�;�Ѣ>;��\�П#����$TE�4F�x9�I.�z�ף���,�e�9��)Oo����7_P�$�#�U:�HC�h����s�f��2&��C������*���+Y��-��}�䶽ȻO��Tp�h�o�C\~K}���	p-�"�4(�U�����IjH
ԯ��wй��W���<��'�(P��Ð4ݷ�$�֪'�b	�"�X/���*��/GG/E�%�P��������N��-���q%�e��g�����ʢh.���4F�>�Z�U	L&����u����;��.��4�6D��t�kbJ�"��kq�,0�o
r.�7������޺�o~�����"��b>�f6�l���x�YP���p�o���/�⧩������� ��萵��S��J�*�VJ4�2.[�N�t�JS� &1�CI�rG�W�{�|��@g���~%�;���I�w�N�j���R�t��2��$��]}�Œ�)!j���=��4a�!3w�40�y���HE�4�[sBD�3"�����ٲ�r ���)�C�>�1�n����<����.u��v��/=�gB��S�¡��5ϱ �_���~n���1�<���l����ײ�5��_�z��2�Jň��q���D�qGϓ��S�N�����o�x�l!ɢ+I�\\�N�.�bl���S�?����n�`Ȃ:b>��uìy��gdoQր>�T�,��Vv��[>�*�Xc����dQ�x}�O5��ƆEG˖������6�?[��B��������Ʈ�#�8Be���m���+L'����gC?�lF�3'�V�I��z�;!Xy@A���-�+fB�
����-U���.���	bu.�&~oM�v�37��5[�thk����Y��>���K��K���a��s���� �1����g��5\�&��'O�Սu�������Y4%@�}�\��>�P�o�~���	EI��רFV���o@rr��E!v]���5�q���+�!?�jH��Z�Q��깹�Bq��F���f�P|����t�D�����!7p�[����g U��񅄠
�H���U�T�Q�8���F��\e�P��j�k����7���Z����b�@��M����pԇ��jǍ��o2�ټ[_���4�D���A����1F�^�r��-��A_8޾��V�7���6��Up0�����0�64)@��o�c[dV|O
^��hg6��AN��O�9+�/3G��b���u:��|/�oI/�h�q|�����	�9��RY*@���"P>&��1M� ��IM��W�i��:
�������u�Zz$�V�c��:J�Kr�v�'�g�hIc� 'D啥��\�8 ��J��:
�r%�1�s(�U6��c��Y�3�CQ"����|���fqA�6�m��Q�n�VV\�h���r��B�V7�%8��'��+��r!j�ӯ ��-�B�#�D�VD���5o�`9lG���d�s��I����/�Z߸1��S� ++x�ķ^�nS�vܭ�t��Z�ΎZ`o���J�a+�2:�7��L.�fo3�u�d�Op���4nҟ�A�umpX�Ґ�/�j�d �#n�+�%9�ŀh.Ri 2��P�6�ȏ��*}n �RQ�������Vg������:`%*�.L~����a�[�fn�DE��J�ᷨ��wgE�o	?>b��-C�
&k�9a�>P�|ٔ��Gk�=))���[i�	�4`M�C)vj�5�>�#�Vg�m�+_7��	�6�&+�؟��* vY�*�,wl�E��a,(;
�4��p� ��V���IMe��1���Y����Ί��P�늝L;fct��'����9x��x�2 ��nmVdXo��l���$̾��H衒h�_[H��0{,ݰ�k!��ı8�����wl�Y����T��� co�N���7�j:�	?�0'Y��;��,a�0�w�D�Kh�~��U�;!�+���w` �E��O2/�BM2ŷZ;'�/o��>�)��j:���}
`�٫��)�0�z�@�U�fH���P�AaOh	n3%�G7�I�*�e$0��Ƣ����?�(��K�|�q�3Q����Z%������)Z-�ޗ��n����� ��r�4j7�z�'��P����w��y���I]Q��u,�8�Ԑ��#�`���9�7B!���o��au"�5�r�ٻ�P��Ec���f.�<V�d�P��ۖ��Lw�1��w�1�lɶ۠��iC��J"��{ ��΃p\�KZu!>�}�`�(��>�OG�@�Y�e��3bӧ�%l{�hg��P�*�%�B�;�����:���ѹT�~Q�a�-��䁽 ��)i����� }/XR.զ������K.ݵ��Y������rfYN������}�� 9Xr���K�{j�5΂�����*��f���
��
I�@}x�J6R��tO��Χ�
J��`c܅��YƬ"��&:��| ���p�0���J�a/�V��t�6Gd����8p��y�9�SJ5x,��h8���Ҋ�È ��e���֯��@H�˺�2�����V��[z���ap��$![�
�ܾ{#�V��@w.��u��Ϋ�v��Qp���H��a;�R��͔Ф(l+l늡;�D�ӠsMu!�=Ou��h�n7�]��a�?^��tdF��3dz�S/�2J5�fwL�Fh.^�^�.��a�7�%���
����G��j�}j���8x�1��i�^5Ou�p~L�N�#��_�4�Ro����ៀ�+}�WO9�����p�s*2�>��;������bw�.A�I��I�	!�_\Y�f4�-~S��͹���t��G�l���W@̄;V�ś��tN*��4"�G��C{����6�V�_�������Ó���&�[qf����v��v,�}UԒ�06�o�؃"�����ϒk8s����<_�����Z������d_B�t�@W�~(S���ue��H_���jrK8���Aɘ���q|۠���] �@|f��=����E����C��r��Yc�� su�ͼsA�
{�����e����}Ii]ؿ����."�@-2��ɩ+z�����?��:Y� ��dfx�{��ǒ�dOA���_q{��W���J��N�h��)ϡZ���
ὔ�GΟ�t�>���X���|��Ԅ	PMQ�%9	�4��}�&bI_�	Ϫ�L� N!��h4�=I`(ܢV׊�ǰp�P���'�:�Z�3����][@�"&����vfB�Yۧ��j��ţā7���m���)ZM�������@��_PQF6�"�ku��+3p�Zl/�:�I�O�M�%��-����D�����h ���t4 D��6�I�MK�di�C�+���̳"Z��Qu+s#�G+e�q�G�慥�ԕ���t�<�n��Ia}Ǝ.�ª6�ۤ�͢��0L�B��S��[����'z�#�=���Ƶ3N��ƨL��ҢN�7�_֕��uڱD�������~�92�vl��	ҥn�����xgG4�q���Δ2������U�xSj��C������q��f
�ۨ�&e"�!)�9A���U�+B��n��'A�lzYZ�:���qc|]�\h��Ǳo��7-���<���'�I�஻#_lq�����2�m��p�2�ѷ2x�Kw��)rN��sV�P��,�r��6��c���G�����4}TznԤ?ZV�"�w%������E��3),�m���G+y����B���x�e(&_�\�䐐���[8S����噧T��͡',4d6��'I��](���ŴP���]+l��dDI
�ȷ�X�ײ[����E���x���?攲a�{r����˷���J�;�V��yvJke��ѪJ>A.V��d����v���߮�lPnԔ��r{�� F��w�5t�"�|l��+�b�|�� 0������#@�7�T,u$�T4�^��
�*�#�f����k� �d���\o��)B�R:�	B�7�o�-�&�wy���W�;x�_��X�ݮa���~) �g��5�#�K~�J:�
�����~+�+�P���n�����(�T�g�'�Dc��Y}���h1@ώJ7p{�[����z�h��xȷ;�<=$���Ԍ�R�Q7:e���%㺲vi���ؾx��=Y;�N�ڂ�M��j��������o�B�ϻa�U���U�	��L_����S�k��;X`��ݭGJ��ݙ'�x���5��}{g��5�y:��v�Ʋ�9���꧰839Oz�J�FZK��z*wڄ<k��u�ApY�M0���6Gc!��T}��O]qm�4.��)�a�
mۖ�u�fw���"�n��\a��n���驓��Q����Y[�]��*�*V������]zE��� �����Q:ܨw$�v�[Q���s�l�ʐ��M`��.8�w���?mJB��j%R�43���g���bi[�b��ր�S���ޚiT@g������P�a;��n!������ؒ���.�;��qM�-!
�����w�S�@�n@��bi����Sw��W
��a]�b������~E�6���j�a/�U|p�_�
�����lO�eV��cU�X�2>B����oX��"5�o����Es?���Qf�a��έ$q���I�Y;�(Y�@ف^}B	�I���T�����/+�+�L�L�]h W�T�ܸ�%��&E�<%�7:�퍀8�a(`wD|)��}�u�$�_fQ�u���ԓ�6�u��'�ٌ������*�MU��wS�V���_gr��c1&V9$Kn�op�M)ܘ�r��PH��s�����k�5q �$�ד�|�-�_��?޳�K���,m�k�����͒��9�'��W�j��Gy�<%e��S�w%���i�E_Y��ݺA�(��]v)����&|�[�4+q��cJ�"ir$����J��X48@g6V1�I�5����s�@�(�/}��O��8��!q i<dO2I�N�F��<�,���l����nA9m�ZP�<(�R5�pi`�'�z�Ԗ�K�P�����(�4	]�<�(@"�?�=�OU�~�톍R04~F5�{N��X��!=�⠙	1�����_Ow9��)"�f�T]̀B_R����?_�^�kJ��]�? VJ�:H��U���Z���9=�5�3�� >/�雉V�I!~�-�F�U-��.n�h�;ݦ�B��e��;��*�!`K�-�.����\�����D|�Q����v�5�	�~��q��L�$�}�l&��ѧSc��s:��HR� 6��@���I~5��I<���j2AW|�,�W�n4	������p,\D����^FYT���e�as�n�,��%����^����DL�r�t�8��O�[q���-{o׾Ҳ�	!��D�e��p�V��D�O�&�K����U��1S�� �����}�k��ݬ�$��h�$ᆺ��*���s��,O0��0�l���t[��JKÕ~F��,ϋ�T��d��=��Ad���+8`�\�cu�˜��$mM��{M��X��VC;�.I��H��wuM� �/0D�yDw��1�D��.�K|u�3X�����o��'e�Nˀ��M���%R�nNO�a?h�g���F}�F�)��i�������z�q�T����ћ܍xE$0��N$��;m��5�!��c���!����8.E~���ai�l���̕�K�H$��4+��E�,�T�����8G�K��w��t�@��Q�65�c�c�^�A��5~��:w;�t��9-��X���'Ў��K�Z�/���7l]!������ߩ�sȻn��<kO(��G��ZX4�'S�k���c�X	��+�jhA�6Ђ|��:��l�.~/����c�F �������_y�M�[��osdZW�=�Y���}- ��L�07��(@6Axּ-l�H�֓�ۉ��7��D�0�t~k�Y������LS����*���V��o$o|[��x��P݁g�g�x���a�����B|�[����A��id�b��k�/)�� ���%��V>�����4�0,b���զ����D��{�y=��:<-�Q�:��p�\��;\F�;����2�'�	����2�2��D��:���9Ipc��-�e���l��?�ِ�K�,�s�&�$~�v�s�R��T�\��N|1H^b�Y���L�)�����j��-j�p��y�$�-�FY�:�RE.��!���0T@�/ I��|�B��j���Yr�J�0�A��{�ȣT޼��,�fn��O�R��i�VM"1�2G��j�A.B�9��s��(�f�z��Z�Dި^��RGc�^R������<�!��ҭF�6K˝*��>�}{���"d񿄥3#R������+ �
C`<��*1�I�;�kO�"�ʧ�ψ��l�{iO>�^\��>1�_�=�x8��K��=�m�^5\-qU?A��U=���z��=d���O�0�9�F:4�DJ8�2�*��o�I)��ǧn/R�\R����L���x.��� �8�W�7 M�ZW3�@�X�KX����ʁ
���vh3����`����I�&�el���T��R�� 4��WZ�9<�Ip!���1��%M�"p�R.J����gȖ���~�z��s���ZјxQ�9[�+>k�|AO
�%�Uy'���A��1 ���B�	F��L����-�p�fh�Ś4&k}4��E����ё���0�qK{����D4�m<����Br��Z�������U~���Lb���
=�Wg|�hou�LXXa� q_qo�V�2T_pr��p��C�W!��'�m�%���8���H>[P�.%Qdw���Cm��\�jbDjrQBH+��L��.DFSx�W5��iE���?]�TZV�)/�<���(��Gy�'�UOj5���Mȵ7�{�3w	c'���5S0�Q��!�����&O�
��wkX�8�K��@���d�6 OM���@z����4��AkɃ8� g��H![����fy��I���f_]�`�PFY�>��{�L�N�9��	"/�+$�|I�!�a��XW��-j�ث�u|^Tk��e�{�Nrg���f��9���k̹K�c`�5|��]R���\'��&�_y�'�=g7�����K���#�eޱ�v��	�>�
G��A�'\���p���2�C;E#�x������y�ѥn���� ���5y�Ƭp��r0<�Zd���TZ�ѽ��nd�[�5Q4���ޖ�Y�=sn�帚a��-�t;_	����	H��%��4R�+��X��Vq&~�߰��>n��ܳY񧮠^��>�^�L���V�)J3р�����k��ŏ�G�T�w�U=����7JGO^�wr%'5��q�[�8�����,oP\�v���99/�Eﰄ����'qe���B3`��b�D�'uv(>z-�w���h~�?�Jm/�N~�"J$jn���+Y[�SR�e��[pDF6�i� ����=	1ï��c��T-��t�֜Ht�O^��V�+"(���;/@/�.�X>�^���A/S�{����x[q?U+O�o����I$��d���D�J�r�/]jMR3��+���D��@�ŁJ�EM24��.A&��4B9�A2Ƶ")@Œ	}���A q�gA{Bx��7r�͛_e<	Ջ+��ꕮy��Uj<�$z��t@[�@��
x�t��PT��ENl����7fk�..�m6.��C ��)��	$;��0ֲ�`C���v�E�-�`6'Z,>�L��=��B���|<���*���S���8zv��`�ܰ.�@$`�Y���n\���O�K�w�$����>��/qP��m,E��ƃ
(�����l��ng��?� U�{H$v� �!?�ޢ&��&����=�(i]�^�����Q�Mt�Nq_V��R�'�dAq��eX��6��%|�L�/�f0m�-��Rvʔ�@�������S�CV6�Il�s��c0=���!�yV�/˧R7�H}Z��-��kb�CX����9�%�.&DZQ\.��1#u�@�wwQ���2aRg�i�c�[��>f�)�˥���fnX��%7ʟe~/Q��V�`�-6��c��M�s>u7������JRfk~߲����d�.
eA�Yne\>�[e�(���ǣ�j;��E���F�&Q�󧒻5�Ծ�����L���{atn��J������lR�0M�O��������@����I�N������߸!��'�[���rD'����i�~>�[:}1'y�@_� ��~"%9e�ղ(�H+�R�Ì~L�y�����f$%�|~�����\V[-�|�^	��9�ː8���r�O�"����7C����Qo:�����E/����=���&�Y���`n@+1=D�c�d9�2^�D�7i�$}�B�x0��jdŽn��=�X>�����>`# ή�Z��T��%��T��꿯��<�
��If�h�c8���{��;��8ڙ~;�Q��^O.�5����N/}q��e�/[z���������cu���g��;'�La!��%���*���*��!s�^�\�C^��@��|��9w\�� %�� ���C���Ze��O`ҍ�n���X��!Ǘo�+'������J3(�':�6��Ѽ�Z���}UZ�u1E'��w��Y(T�I"�q�oL�1g�:|
�N�ݍ:�ʥ�n<�
�ڸ)�5v�|�Z۩�R*�"U7����%+,S%Q!�1�r�7�bA�� ����r��jTJ\��dyit�"�L�,1�(��4E2����w�:&/��>"�T!�G ��1�;QU���K
Y�o�i�gQ"��8�F��g�_�)��U�vwN蝷�6Hg��0R��gS�`����������.��U���CQ(�'�Q--%_3nޘ��@잱���y�:�)mO��ŵ����,,3#E@[��s� f1� 2\����~Y�;w�cd��oו>�z��)+����QH	{�bZ>�TL�Xk�ypԦ�_�yN�sg(�Ū�;�
����}� ��&�b���v?``b�@N�<gMn�抻AݒKhC����wı$.����cm^	�@���.���.����� �t�X��女�QF���ʾ�uHJ\���q,��8�;0D:R;��� �h&����ۑs�;�I�����	�*?�$��ԖQ��U��Q󥚑XUԻL �;�H�EG���(�w��r�w$�2��~{^������.�f`� il�ZK �Υ9��d�0�t}wK����'�1ٲ��ؠKb�0�+�T�|�8�l�3Umҭl�TF�
ê�xo�(F9�pV\�DSI����MF����� �r#!V�K��=
����=����<t�������Y
�5F�������f�E?��(��MU/�zS�l���7�]h��oD�b�=`K���w�ԟ��`a"R��ȭ����Mm@&e��Ⱥ�O�w_����5�%y�m�yE<C�[+F���H��qc��:�3Hw����"8L���dӥN?�U��#���'	�y�'t*ã�&����1�!�@U�u~S}9���
�i��/��'P},+�kg�i�1t�.E]�z���B<e���<O�N���d�{�kbD�U��YȱX�W�D�߫��`0퍭;n�M�6�v�V��c�&���D«PB�Un�f��` d@[�9�{�@��k&�`�bW�w}eo�Ľ��h�]?U����{!�m����E�F'�I��R�M�!C��3?�JV6��\��ec]���V��MQ��޷ֆ
տmN� {�M�u����KCVKuU�?���0j���cG���)��cY�e*�*)��xp)P��a�#��8�Bk�\����� �%'F��[������?0&�=�k>N���s�g����/���� <��e�ҏrtt�% /�ur������L1~� ����³�dZ�����/��_e�/����o0���4�	�\�����W��	�mg�@Up?\�Ho��vj��%:=���1����u�ci*og�ǂ4�d#��Gχ�<�1�G)�G�(ĕ��Q�&)�%��k��V�
������;R^�0?�^�{��J[��`ؐ-�l�5x��g0���9ٯ�]����e� �Zp�qt@M�~�|r�e�Dil�P�V�ON���
6���d�����ۓ�Ҿ�H���w�|��R }��7�X�H��I�/ڒ�S��@C�G�xT�4��龥�
g<ERmKF���sr����d�dN[U_�G���b�Xd�K�ixX����!!y<�!H�{�L�쾞�}<1�A;
g�6�{�X��)*;���h,�f��B��J�䴰�\��+���϶u*��D8����@�'V�Z��Ϭ};I$õU��bEq.�]E�0���?%|򶇵~�
��b�v�Ruǽ[�*-��C��&D����/bqp��'����F����rU�u���-�_�O)ZH�M.��+��ԅ��:��޹m�Z�.��F�{�猤=��Ye20�K��v|�Q4	�F�C�
�=�D%��m*_c�ە/�/�H*g*8�θ]�ޤ�\/Ż{�3�3�<�Ld꟮,GA4��07��N��.ĉ�쨚2�B�}ezNBpU���O�8G-��G��_k\L��$��ƨ��|y�*".�n]�2{"���52��iՃ�_!�1%�s/�A^���w�� ���F]�r2�E�W�*.ð�J�d�aiY (��C�Ť8>�k����ʳ��pVJm[%������{��͍3�b��(C�ٽ��gJ�ņ��贂�S)W�qN���*����C<˙�9�Ӎ�:�5ۖ���y�k�2�*�͘͞G�L��.@͵�6��^X �v��{��٩u�a8Jci�)]�&D�5��1�T��{���m6���a˔D0SW�WE��.7�#�a�ߓ3 a�ȣ��E�4!O�i�ψ	��b����*�dM��-� n��,���\�M���`��JJ���T�Dy�ɐ8����s�|��Θ����J&� "�e�m��Jkd��X�7<�ֶx+�#��0�@iO�
��cjו��+2?���z��)�㮾{��:gn\���j�����"~s�T�Bў�B�� "�ҳ7*,Q�"�$��D:c-wҎ�'��8�O�05U~�ʏu�ӽ�ҵM1�~:�!�wl��2x�,8��f9�F0��G'���cn�e�sb �)��2�~@��:p����T�FtY뢮Cz�>�?��R|��zS�<rK)=/����b���{���_�����^�&µzyP������β��]o�Ǉ�?�RX��=����y"�ð	.��E������ڃ���U@/RR�P�V����\{w
+��\�=O�z͡�K锉G-4�N`~U�γa�!�4X��y���?��Al�*7�T��E�O�9��;ϱ�'Z��	o��d�疏�a����P5gr�7\��ڟg�g���a�z]n{YI�5<��'�NbsM��'s���/�iBh�1��Gy9�+w���q�] ���z��8~v!���h�Gg\*�1�����{'��.v if�R�����'���e-b�V/���%_���֭4������5h:�oWdV�kG��"d��`D�9�����Z,F�_��1�>q�C�ۨ���@��X��l۬F9��٧���,8��j�H���yk���&w�A>EyU0K�Z��nŌ ��vm�LK�*Q����^�AD"	�W˴��N�׼ё�#��u����)4'b�rd��������jT��K��0��a�!32.��nq�������DQ�V�W��]ޢbpx#H=�ͼ���?v�,m5oG�霅F�ӵ!p/��C����4l0�E���v�3�Ἁ���>-E��"��Jz_�aܺ� �d�f�@,Y���p����(>����^�^L��(�~����ݑ���������>��[}�ʪ��s�I]_�}��_wT�G7ҭ���,���$b���0��A+�>��`,�/���C�\�q-z�8?�wph��" .
B	ni�h�$��f# ަ	����`>d��M*��m^�P��`}���8Wb�5bS��+�OD��@V@);�S^��m� �Ԓ��Ieu���� |QS�/"+d���({���[C�H�E���@��h�+��V�O��""��z�h��?>�e6���h\*�n-�Ө^�|����o�3;��ۺ��a�l9f51)����v�n`������vW\��E|�:������K��'�!�%!����m��Co���V�}�PiiĂ�ƪ@��w���U�K��6��-�~*�goC�\�o���K`���1��\�-��Rt&��@��K IX�}I�@����Z���S���I�9s��+)��Íp��	[}WBoB�A�Kٸ����A����DPU�7)-�@�p3��q�F�;u����TF���κ��mڏ����,{p�G��|��i�6̫������k�*��[�G(FݡV������*ه��<22�ǂVy�,�V��t�jS��x��5!�����p�\�Ʊ��n�������0ҕ��g=��䊠�LH�l2�))0,�{mi����m�#�i37�9 �nX~��lF���H�Nt��-hТ�����b���͗��Zp��<Љ��I�a�{�CS6�ʉ�G�k��Ʃ���*d1�t��:9�B�Tn�K2�L�����l,�R��q�a�F��;�Ln|X�ޢ󖄏(8��r%I �ڭAR ��aEk��dKw&�16{p8r'��+5�U�3�7F�����;.�C���==[�V�A����'[�#��w�?�>딀��M��v�Vʓ��ng�xPD�
����E�Q����[i����3~ȇN�̸��)H��)gک~�y4����B�)��՚
��qq�l��V�� e/.��C��c�IEqm<������:�^�ĥ�#��U�{j���!��x���y48�z�'1���k��Ɂ�ld��A�'~���B�o `����^[��X���j��h� ��hZ+��G�b	�%G��D�a�D�4����ku��?������MF�dv�̆{��6�ѐ)�U���?4�(�4�3�D�v��GΨ�D��_mdi.d����Iu]:m��V|�\�u	%�p&��J�F&�|j����2�W�� �_�_o����~���ݓGq�{3ܣ=�{YO$%��7�R�:�G��%�8��><�tG'y#�r�9ܑ����%���g�Q �u�����[��� )���zʣ�� &B�[N���=��bk!ؔcD<S��]�Dk`�"�ߦi̍V��}|
f#8#]����B>��̠�
(��D�yB��Kc�å� f�����`��w���	~���������2��b/I0����m��5�qwdF���	�N4�wU���:���rl�~�;���1�z�p��G)� b8$�~�x�s�w�3�����NBz��2����v��6����q�����&���O�:���)��:tr���9&uL�a;�X�F�����+�j�^�.C�BȢ
�P2��Oԑ����^{�4ej�%�-��P8����"J�M�$�8i���"�� �%=aȓ��C�A�7G^,�@sJ0�⁢s۱��R��7��0�[�ey��,�&%�n�P�#%�b�o�o�P��0�i,�;�՚�����f����������p��@������\J�.�$�z3�w�hC3Wy�Q���A����YWf��f����(��L��1Z?<�V����̧�i	�$��&��K_8���H1��S2��W�@)�"�ld*���˸���\4
�ؔ�o5��������=`���`���G�榈@�`�jd�PKj�C-����$NZ*��y��$�vĚ�=��5�v�m�e;�;�>�{��Z3��d���i�a+�IT���wg�L�<�(��r�����yTM���t�(m�D)�a�ޚ�Cf;	yU=&��W8c��������.&���磒Ȓ�_�ԟg!�ю&�sz^g�'0sI���7���IR�����n�g݊~��2��<�$��	���T8́�]��U��TӼ�18�%�>��H��Ȣ�y\���4��x����T���b�\1#�dx��lc����p(s4�
q�c#��x;�h���T�O��&�i�S@�i��3�(��=���򵽍?���o��M�����.�hS���W�q��u�I�B�2~�!��Q�K��WY��-^x
r�?y�{�M��O��Ȕ'�LI^�1��~�3zZܰ���*�_�0q�vDTЕ�e����E��.#��p|g�f
U��wɢ	��f�:�t��� �Ǟ|p8{��>A��|;������og���m��:I@ѧF*4D�Є�t����ŵ�P�_>��XB���A��U��@�r�-'Ӈl�S&�|�c�g���}J�_�{����En�5/���k%��ͯ�|׈�x�[�߂����N�b�Q������7��!�"�����i���]�s)�9��T�of)1�}�R�AY��:Ql��Y^)�����nD>�pk��ǥ6@��ڀ[e���>I����*���Iy^�mg�ǳ���?��u�q��u}�1���E��m Y`ꏷ��$�.*����� �_��K�Q���̳mE���$}(�B�6t�! u۹Ȭ�O`b�wE���0��:t��~�y�F��Ь7:�� �D[V�hR"k��q�0~Ѓ�vT m=;������h*3'���@�(�S��yi�3ZF��< 4~O�k9sx��� p[<`�e��}!��l?���&g,-��c�_�Qr�3�vvNg �c�"E�@A�2Dk5F��n��@�]���w4�������<���m�@9j\�3H����p�`G��JL�F=�y���`R|7��p�A�J���&�\��	�kx"Ŗ��4��c��!{rs����ڂw��M��E�$4_�!�i��z��	��r��ޕ̫2�g��j���0�O8x��0M��	Ⱦ��8�i��y��:-�$e�_�˄P����o�����]�a�"��_D����7kj���}��L��@A��b0�P[-
�4.=�}��P_��̡�ZGnT.Q��4	*(�=���{c�JĪ��)�+��Y����;���-翡X|�A�-b�F�/M/��Kn_-z,B%!0�@_�C�~L�� L�kV����
��~�$�	h��!g�����x���13����_�ȶ7�����k��-��_Y{n��g�&��Pf�U���Y���~�j�w^�c�>�I/i�ˠHj�d�����sl�W��2�z��N��g��~^��#4�	],9�����:�D�q��������]*0:_��<2V�MJ��^���fGQ���_"0���������f�|/���4�Ix�����h�D��t��f0�HҵL�n��f��kK*�bBG�� �L���Z�\���x
  W���c�+��P��P�Լ��oK�戟8��U�1�~_0�;�͆�Y�~�:�����)�Pm8@���]VY$��`I�}�6b��/�O��$���Sn6�	8���6������v^��W��[�M� �{UY~�~6���s�k�T�� ��j]լ�b�g���`��['�JNJ���N�K��7�f�}z�'S�j���9%5sO��OM'�>njX��F�E5��4o�6Y��8�6�1���d�<��+�MᄽdW����9DJ���G�l�0��\�e���F��ETJeĘ%�piz,����Q��35�?|��4Uab�
{��o.TY����d���H�o�M�O�!��8V$ �W.̢��5���3�I\��8j�ۿ	���q��i"T����iS!�Pq$mY��/l�SQ@&��_��bn�aǅ�rb���;�'�H0=���2fe�kH�G+��upT�*ט@��(+it����O�W���vĐ�
����u#U�	L��fnV�mL�^��<l_�J�H`�
7��}؄�'Z�O\��Cc���C�����6E��[����mB�7��X��-��p3�փ b�u��P��1E����r�i��ց�G?_�ŏ�mp'�\�ڼ�(1'k���]uڊ� :�
�� �D7X|�Ty�|��j/��s��3Hi�	�1n�$�q9׈{�D/=�y�;{m�@ٺ�ө��dA�Rsa鮻���42�q�)���a:>c�����ǂ�b��)vڢ�v�;&,q�Ǔ[�>y�C�lBg�˖���dn��w��y�m��h�X�M���l�W�9�=O���'e�K�1^º1�]j#f��L���g��_1�#�t�
<���l���{�?B���+l��,p�%�@�Q葫�/������&� "��.��ن�u+D:�M��:�"Ċ���g]tfh��hG:��_�`����00`?_C�s���-6jM��^+Wi��_?N���U���2��e_�'{R�2*���GI�qks��֝"/a�TG����(���|���/���ֿ�J����%K.��5�3,d�/��z�ɝ>�A��jU���6�_G(^��`��������J)����/0=��/���NS 6��ޑذH�x\/�ȟr��"�̂&~�CKw8�i�K�	X�k���d��|�����2�>�2�i3 ��eC�	e�7>��'��R�e�s+ӹ8ʱ�{ ������A��k�+�Sx�*��3�������E����\�9(n!z+�r|�q�l�����0����&����I��"�#�9Q�i�N�C���ds��C��pA��Ɏ��W�T[ψa0�T�s>J!�V�~cL�9�j\�ɯE�"co�p�
E�]vyJk�*�����9�����=U�5�xT�/�F�l�]��c�l�m��aa��8�P��﫱� `��G��TS�:pd����u%�7����n�-��9&�Ӏ.I��
��BqS����Cw��굏����s�@~�0�)cl��}�̚;(G3-���G�a;��A���)�ލ�֌�ǘ������_<�>0��pb,r�����㨛�G8�?PBE�m4�bS��6U��,��*�/���\�R�y;.a���`��8�^S�p���Վ��;�����c>�A�N.�#��b�p�/у�P6[m
�V��p-��͡�̍^ K� �����o1!S���]�8p��b�9��K%Gk���9K�sp��c���}�Y�����;��ݾ�j��smv��m�$���SF0�'�Kr����]=�z�8����ȡ�P�j�R&M����W��#Ɔ�@;��EN�,�3UC�pΗ�a�V ��_siL��eS;9���ua�@i~a�3�g�*nYC#;2��4�����Fu���OCR�=�)$�y�6�Q6?����;C4��¶�l�k�d���,�]>��r�v��"͚*B��X�K�*" ���`���	�3W���_M�\��V�o|��j �lv�2MUW5$a������M[��g�Sy��	\K�d����ݦ:�Ql��g`tw�t�D�+������׉��԰�~�!�X4�/��b7J�g䵹� +�jNxT�[m�2�$�B�1��#):X�� |�.���>%n�����!l���4� �'�����OɎ��8E#�� ��0*�y�6�"�a�؂9!���x�*W&��H鐩��a �����v�	ot4��p�!zJ��G�<������a��ÖgPc?�tNcf3�A��рx��X+b^��۫J��J�1{�J�+��Q���&�C����u-_�6:��GP�5S�3�}Y�I�H��^��~lGt	�@D���]<|%Hey�k
���Wu��a����&D����7ʱ������[��G���	��Se!�^�U:��Ð	EǇ����2�&�8D;N�$r��,5l��T7��RF�(�nJ�+�e��<ݸ<���E�:7�y��׀,
���E+{�������{\��c9e�Ei�:H ���p��߾&dNOL�v��9'|�W%)r�fP�����xl�����u3�s��EWf�VɎ%;7�y�I%t��(�Ir�����M���+5S�3Ή�	���|��Y�7}͍��jW�}���������*�هYF�d($�*?_,��*�c��<e�S���N)�A�2�=��]�̾�]M�4��Py¿1o���"�0�:%��� 0/3[��j�摹u�M~u��=9�cӺW&~Ii���5��k\������dK�0،b"��
ݷ�tx�{�>�p%�$�p�X!U�h~���P�����	ڣL��:t�{Z`"�7Sw�+���Vm]�3z(�J��` �uJ�n�n�^Mk��Z_A�Vz�aO�0�X6�t�l�!Y����Y�H�q� 
�"�3'ǟo�ѝ��3B��R=36�U����.����ت�����!t�j�vZH�}I4A	��wH~���6~~������ �� 6Gqc}����/���XnPOC�zr[���B�
�il�ouܓ�qU<��(�
L6y�F�����P�[�.��ݰrBRA �5��{>�S#u�s<k��0��ɜ�JzR P����C��I��Ԧ΋F���1�C�C0����#KǮ���AI���xf���=��U@&��|u7G)n]%uq�����gyj`��Q�Jo@�X���͊�=\��X�wQ�	?N�MN�����қ �j	 �g k�k��p�|yr��<��N�Ek�݈9+u��D6��⬄��n�гϟ��������)��S���M�H;/7q��7��]v��O� ����jM�[���W�S���!~��7f��`A8���O�E�<����q�R�8�|�C�$Yu_>����"���
�<t$� �pY7��X��0����<R�K3L\{��)�1�?���>��.O"����i������,5#q�v��.�F�
�]g��BL;��^/P��e�;�d�����J�m��4'��,�lU�]�x���i ����@�O�C�Y���By�����5W�,F�.��̿*�~�C��
�c����ֆPn��=�;�������+�M>�0�O}��Y��cჇ4���ߥ�(���P9֓Z��Ds}�w/Z�~ƚs��R�J����11���rm5+i�5a-�[	p�����o�l�����z�#ٔ�9c� ���]�oW�L�LH���!��+�͹�o��i���d��it���
M2�4Az\�2�e���|4��Ƒ0ZEt�S��M��WU�G[�0�~�L����s����yT,6\h��-�lk��O�	��W�z|G���Y������Eɗ�^C	շ{�<�Y���pj�>��`���u(��pȰ��Q X�Ԧ��F���Z냉X�ί*���'�9�;�����@߰1li���J{�Gr?~i�jƅ��Q$��Z~G�%p�｡9/\�CN!��������F�c^׌�@8`i:��HGْA(���w��ߪs䢅�-dw��['>�9�Kc�reW��3�?-���F���%���te�5"0�j�IY�~���7�^�O��%�.=I���Z��3x	�8�.Y��" P�վh�	��F�7Nx�Iw�1O��d��~R*^wN�"��WO%v]���} �}1.\��JK����'R+W�sv��M����h��t�c�'FD�P=R��#�w�Fi��I	����螛���";vG�J	��:9�x�ނí�PG�����<� �ܭ5�d�[�V�����W�6����ƌ��h��*{D��9q���*6h:* 
�S�)��\>(#�Y6��k-�mV������"�:��4�E�|gÂ���"� ��9C�B&�U]hI���baݝ�/��[T�\����jqW���-D�Ng�^˶8F�42� ��elhh�'v$�Ƒ�m����`r�*3H`��H�#<׻���͘���C�cFq��&ma(^A�u�v��%1d���hͭ�r�!�y��9�ܞ��<?�"7ɲ��x4�I7��.�����ƈ����p��3V�S�4%%\���W�������슥N����k���ǁ=?S���VW 
ʨ2;����@$I�v�fk����&C��!w6���g�oe=����7��u�3���|@85\���)��v�G�����]}�<q��}����?�#D������a�����X���������U9FE� �pdx�8�j�2m�5���O���A�;�Bs�e�8���x�&�����AT�N<��>�"�vV�Y���4����������-"��gN\U �\�0�\R�X�8эͧd
"�[��Rt�}�?\�8ٮJpg�z��M�����i絠a��	z�b;K���VE���ͤ�7��ū����ノ:���"*���ԍV�[G|X�0d	�M�o{��~��?�XE(g/洲��ص�.����׌�-~d���a5���{`H/���4l�w�������&��z�O�ג&�lR��܃K�H��Ɵ�����9���a���ء����k������D��nR�o�8��n�-��-������^9EE 8�'�:(�))	�����U���=]s��E����4Uk��֛j��e|�ZJ'vW%�c�e��|=�=����Dk+��0�����H�(��;���+�qJ^��i�MH�K�Ĉ#`/4�>�ߢl>ϛ�K�_��Nے(po"�wv�G!���ѡ��s�<Iih^fc!}EM�i���@MW�ｦ\��Um ���M')p�d���w�(����Dq�X��x1x������p\�'f�b�@���)G�cb��>����%cF��
��+pQ϶� ����j�������#�o�.{�c�i/�vk�t�(�ڇf��Nl����Z2�)~'Y}��6I	7�xr�\*O����Mpf����O(JC�g#Jj��.�����=���?a�+��^����U)�l��6�c.�%����"�ݒ *�}	v������Y閒��b/2Ŗ�r�"6��_W~��QM�:�K����Y$�'��̾Ȗ�#>5�~��v�@�;�Q����N,�����S�~S��Q(.m�t��L���;��O\ V�Qm�[���$qLhIҬFU�^
��=��	�{~�g��ոH�ǻ��Ä��f�fr�j��4Z7�֓�Z�羅�m!����n�l���c�3�G��[>8��{V���������jm���.�;�V�����S�X��5Ӱ�ә��tU�-�)$�H�$[H�Հ85�)�h�X�t!
^	�Bb� ���_J��n�g)���6���><k���D��|b,
Db��sm]�i���x�7��ߨNdlLq�Y������ Ж�B��jcE/��p@{�D(� o^vMP{���G�a97�o�8���`�*D�8������8zt�G�^�Č-�Z���9��T�0F���9��ӽP$��CYp[3���/�JHeI\Ab��8G-�'�0ٍ6�ԛ|���`�1�򯗚ԟ�F���{������1���p��MHr�4����������P[��MS��%N�+�,,W�}� d��5�īa�ϩ�Sf��wR�҆�#��e,�u�?>�(3�㞩�#�Q��t��8�+��K�~��?��i��k��8���A����`��Q�+h�I�eTX������{/�;��:�CG���E
?#"�N"�)a!����Uحև��U(�#l~Pn`����sl@�����	RȯV,ME�g����i�o)X&L�s^�r]yVAD�&�n�si�aڧ>}
����n>DQ6ɵ���Red�����$�0'<�d��	\�*6�:?�\��-�+�$����y����B������Ƙ���o�ǳ�/�OM����f��ݪM��4����}Ȍ���~¯���5�p���Xq~Prr�"u$O���C�
q�:X�/���vS��A�;��Q� Dޞpq%}��Q�N��QR��(��P�/qff.>a�Yh��\��(j���#HN����H_:�沊A>���o��`�g�Q�GB׺ H
NQ8"Q��O���Ek�j�SI\���,�'����%t.�A�q�E%�j��4ef�%It�#���h��~kV2^�R6jp�m�Ǡ�>j]Y�O
�XG_�ɩz'�� v��mxQ9V%>ф�Q@�i�.���t�����GS�ƀ�7H٧>�7xJ(6wK�1���I�H�_��
����tW1hl ��>�ia4��V��M��\�#�@R� ��������]M�c`��������C���g0�j6I)�ar)�F,M6�?W}K	�׻�
	Y���*8�� ||���e�X)sVMH����-�����v*5l�r�e�ta
BU�Gj��/�}��N�$a\�r»����N�	�
����E`�t}�E�����f0Th��q�ZZ��BѬt�_�M�|OQ��x�����b(���G�;��j
Ώ��e���������w��+`�p�\�p��r��Z��dIdE�S���TD'��N�s��w(@�����r洙��+?�s�: ?9;R��/[1Eizh^f;���0�����&�8��������P����7��ٖQ�d�Mf�ԋ�]l�bԦ1��俩�7T>zT"Ht㝿o�G����H|�-V�y��8�J!APq�z+K#VφaM�
.vL����y
nLJ�}w�X|�ӓ�\ձ���Mx�f��"/B���.��ey/D��k���!2]B�ތYσ�|ۻ0�@���ڌ�2&����bBF���Җ++�][�jî��R��]��s��3?K��1b�X&Q�䍅��)m-1B�%�リuv
tH�A�-��-T38�����AP��;��f�9m�����d���NU�g������"юS�o�>�b�d�}��k �M�%]bw���:�Ф�{��Cq���Lka�;q�/�c�DCIG�B�%�&�H��<�Ҕ�K��P:`*����+�$��)�� y3��Y%�O~_�7�f���ʑ�T���T~��)'�S+����F&��C�N�	P�c�4
$�C��J��U",����'!@-���շ^?��,��V���R�%�X�)�R�A2���-���x(a�#AѠ�["�B�3uw�a<�â��T!������:�zU�A;�x|=5���Z@���
�D�\.�������׶�-��n���v�W�)�0���U±s����-��/���.��*j�(Bη4jAZ���ajdx�D�u����ml3�s|z��c��x����(TI�gO��7��h�Ǿ���"��׼�y�{���}���Ʋ�4�YW���F�#��%{hƁ����H_��PV�%oψg�R�����7_&�L��g)�l>ׁ�P�[c��QѪ��#�Ն��Vl�ľ��v��i#l�)�D���%���?U4®�5w!�"@�^�� ��; 8^�����`\�X�>��a�zLM��6{4�fU/�j�9O���[w��Lh��Y���a�FH�Ɋh<�)�y��h��b�X�RH���Ϟ%*WL ��4���U�Bh����w���B��	���㗨�Ž�=U�:�Wf��ٚy�ݓ~Tc�=h�ɺ�����Uu��?&���E����~��^�E�	&�o@ �s�����b��ބ����&B:�)$�#i��&�b�:�,�@��1��F3-�Z�k ���	�ߓ�s���;�OR�w|/#%�qx[^B�K�����/�6�Ur�b�n&�#*�����s�1 >�����2�T���먁�ע5߂�ʋ��Gq�2P;ew:�Ǟ�⁔'���m�l����E&��ͤ����5����;�Y�{���%��(�]o�µ8^������N����q�N��y:��x��nn�tW+��j��r�����v�$��[��Q)��M >s�Eg�g䏸V`�9����%�K-��S	|J��D�@�x���V&ڞ��bp��s�{o�'D��p��SR��MC\_��
�0'-M�R����'vx��to�3jZ����/�`�!Ew���[l����G��FDRF/m�X!z"�Gܸ�.0W�;a���ܴ���^m����sX�"�*V����դ۱���2�-�T�D��<_�(k��@�����EL)6���x�L���C-���%�rE�#��1�%�͊G�*1�lM���	����}���C�v .���j@�E�D�Ag`��s���Z^����x�|cG�=-t�<N1'�	|���$��ܿ�d��xN�MF�N��S؍En�|;�l'HZE��#Q/?��I��2�	Cp��Գ^~D"�^]�9��ߣ} j@��N�܏��ނuc=��k�0��MsӁ�tQ)��[�|�<g��a�	��&^-;��r����xʠvh���C|~o��E��z�|�L����s8��]���>/�p�l	�����\;��ԗ"l�u=bFei�H�a����٫�[��h��-�,�d4A���������µ��:�^�o�	��,@� ��}^y��+�4�D��F\�1I�t^��; 8W �I�N<��# �w�S)�A=��*��N^v�����x�qg�_
Ir1�8y#K�rJ�0��w2E\ER�!���;Y��������8[�T	�+�W��Z��X}�8d��� C;���~W'D/�
�~ E07��� ��D��:�)�у����"��<�ʌ��:|�	������5��u�	7�{�Ǵ�����ڛ�}!"}�V*����T�f,|�GF';���C�[EX�j��r0:�ѝ����0�w�<}!���N��sQl�C��mе0��v���'���
dƲm��yW�
0��AL?9����e��d�. ��mH\��%>o⑅vT�ڋ<�]$n�M�~�=|�q��HD�0�MQ�N��á�)Rn ���c�Z�8/�m<
y��Z�D��%=pΦ�NL������G�ɴ�����d䣶�v0���X7:Y� ������!wx���}9�!\*d{YW����������Q�|a�W���f"�5�0	�;?U�R>��;�N"��1��*�,[n8��u��$��O�A�X�ꥄ�-~����i�����N�,�D�qV�d=�}�0���^���a�޸h�/W��Ȟ26w�$�9��A6��$v�}فxQrQ�𛬕��v�x�s^��Ȁ����d��k���������a��J�;�!_���s�d��-V�ha$�22���#�	JH2:#���y[�l܍�a%�^5��V�ɝ�^R;w�1�Lo���K��H��|�/H0��&8`�(���;.����䗭�{|�|����{$�������aѧz�{ko>��Q���v���'��o0tj���{hr��-�p�Tz�;��T�^�W��idM�ҏ,���f���6�G�C�QAZ�b�/E��4yy�U>�m�_=�|���@OR22��l�o�;�6��Jƽ9#$A�nx�Xuq�cL0o�Nw/�+%��Q��E��76��tH�t�*���:�f|q@n� (�V�s�����������d��m�b��u��F��),󞠟Z�#�6"n���*y�:#h<���JO�d�{�w�^M{/�ZǻG?�ND��O�qK���G��B8�������l��voĮێ��[�mI�����EB�$���Qt�����g���B�2eN�򐇌R{(��>������т5k�b,;A1KeA��{7�ż�b������ނ�#Q���L�ᱽw�7Dp3�%�/n@8�|�%�WC��+|d4��ēŏ�|��Q"�W�=�,�s�^zx�I�*gs�[^�dcd�?��ڲ/{K����1t�JK�^��{� {�m��nZ�j0U�H)-`oe�����U3�Avh�%����h�<�{�,dn�0��tɹ*ǚo��� �#��#�<����K��n�ߣI���c{j�����5c�fz�l~��-��A��7���mn�����8��m�aZ��D��'n�Z���(��_~KWn��Y����FSn�u�ţ+w�/��N�������7\�����(�qu(�'`�%�@d+���z���C��J�x��$+-㳷n���Lm��IQ��YU�k(J92�=b}]�/�i�Nb�&�̚~H=�R���ܧ�T��0���l��a�|g��f����#�K��Ԡ�HǸ�R�CQ
#˖ȵ�t㣃�� ��#�NLrUE�E��������.S	�wH.R���\����k����ϻ�!	��� sy�so�q�e<� >���g�3����C"k�瀞�?W3����`';�oJ/u8�f����(��_��I	5T�^�M��{ڢEPE�-�;��:��GB��� ��;�ڎ�m�ef��Y�^nK@B�暓����x�D��i�7��\����m�e�i�	0܋��*v!�d�(R��֫c�G�1h����lI��}ȃ/>�V���=�y������9��*�2�;��[�����[�n��*#_U�ܾ�g�L"�z 9���#$NoԜ2�4	-�d�a�c����b6�T�v�B�˧tc���i�����'��Px��I՝�C��K� ����o�ߧq@?{<�ze��.����3�9��M�+��7�#�[��ۊ7C�؇�+F��i��a� �LB�0}ZzF������1"y�0��tBL��q(��Ţ�>�^��ҕFkh;������89��~�Q�H�%�gHo��O�s�T�S��K�>r"�\���+C��E��B��X� UE���f`�T�_��F��,K�h)y��Tz�P-�Q�$�YY�g� t	x:v�o�ԏDW�u�O�|�����8�$��O8�hX�TE���I��+9�Ҡ|!$|�`B̀%�fA&LjY�|�"��Ƀ5|��nQ� ���fv���!d!&7�1����irY�x&�ˆ�[�T]�Ix��>����y������e���YѠ����+�.�:ꚪX^0r�&��m�`����nUy�����,��b�yD��~ӧ�����A�h��:8��J�H=ҋE$���p6W����H�i�����.�M���B_����_��[y ��j8Ak��jr�a�����-�?�.*�aO	���~K��g�ޅ� ���Տr���:��'�I�AO�ʬ��5 ��9��kͧlq��y�D,���R�\�e�i�����l�Uey7$�.@�T0�'�d��?#N����F�ֱ���~���"������z�����4��I&��Cz��Š����z�=�md�f���!S���)��+�}�\�|�C3�j4zk�2��4җts%6;�;&�[�I�7j\�`���A�sU�i����*Guz�&'T\g��
�Y�5[#�k�V���〱ć��6?�z�au��n]^E�V(���k�!G㖚i- Ll��&��/����C���a}.^u�^��T�|�ǯ���t䇇����ْd��Z��l�\�� u���X(��a�ڒ�x��m�T����D���y�=�����
f�[4|��'�}�_�qT"�T,B��Y�f������HZ�};IQ�^1�댥�IB�Y����ݭ�2��M���(��š�N }�6�������b7�}F�P�%b����Y)�Y��'Ь���j�D�|!���gC!ܡ�G@[F�����.���H��o
p�F�?p�(~<������/{���K��ԧ�C�R8d_1!��1���`�p�S�ϧ�xՊ0<pG�ZA��Y�l��4^�o�[ �Y�C+j�e�����!/~
��2	���I�q�IYcOMpe,�EJ���w�>��\1�(Z��'������M��S�tЭ�Ӹ^�b۔������Z#����<q;��dV'��1�?�y�{%�+�U�,|%��q-�d�`�tHRy\+,;>K�ı5�X�Kg^gܞ�>0�A�9�ʰ���u}`,=^��6��h�t(a����G�ɉ�74�NAĤRp$"�µ�������r/@e'������HB5.�nw��=���p�_�]l�3HF�u0�sU�)�t��w1��q�s�Xu��=w�[�]��4�"3+i�}nBr>�s�]���|�U����J�m7��Y:g4?��c!Y����hfH�z�u��[	N(3Q�?U
8�E�+Y�ϕ�yLf(%�`����l(	i$�9�����tJS��s`2���1z~@�N�5��������7��o�8��v�0^��G���Lrr��Q��.��5V;Et�{J�"fz}e��u^V�ˠ��XqJ�=�.+�"�uxW��˪J&Euǩ���~��n��Y�،���x���c�?V������B�0�U�r�R+r`��e3���c��ym.�P.*�3{]�L���8�� pO��g?N0L�DR�7�6O3�x� �qd?�o'(��j�
���q�nmZn���h[ؚ1��*�f;4�2�G���-gr��gpo E{��4(���=I�D�;��\��$�;�w��'�X�=�m���DN���Cjr�R�Y�H���^�m;}�<�S1t�$2��������䞎�U��𖹡d�{+�HP��Y'�J��,!LV�}�tE�R���X��Z�o1~��!��ƫ0�
o�AY�����3�Z��иF��|ඬ�Y�[[�cV�v:G��x)yP�_4�#<���{� ��	�s��{���&e�|�0��\V�HN�߉Bh��
���X�3������~j%��0��Y����c��l+�A�Z��@���}ڸ�9�	4�esƼ�C�:�P��@�H�ܧr�Hݓ����#� �v�"qd��!B%/0B���D~d�]\ɣ��)�<.ld.b��e���WQ~V�b��"��:f�8��5j���%�ai�$0�[Dܽ�%(�O��K��H�R� ����J1୉]��cA����Y�f�̀�S�>u-��zET�A�Ff�16�����B�;DIH����F����&d�-���.n}"Q�v��w�Qdm��?�#�b�
���#Y�Q�Y@�sL�`�5(!�T�I�=tPa��!�QC�рG�[�Z��K�P�1���7%!-d�2�Dެh��Q֐�7�OƬ���H���u�!ØВ�f�����V�7��f��"�L�f�Ӱq�np�̒�X�Yw�*���j�__�݆& ��#8�n��h9����4^���%��(xKmVv���&h��XI�θ��qe�F�C����9���!�������rg�f� �R��tl� ^�;NO������^�s�E:<wQ'_J�Otv�k�H�v)�����	�fI�� �KK�~�Cٻ�~2S1U�,�xNsn[��@Y����_R���/�/�hM�LPq.)6nKa�AX�1�� ��j�skQe�J���p붘�sX�ݳY\�b)�w��
��$Zf���HD"���2ކ��N��Z1�e�y[���d,���8=�DE|��]�-����$	�?�e�{�`kyoŦ��gEe)b���~�^Ć!���Z9Tp4*���H��DE )j�[&HiX���|�	���
����>t?�Ejź�\����@���c� ��E����Ң�'��QYIw��A�5�h�#ߑ��Wئ���� ���Y��X��a�[����%��	�;��	:��v4�Q����r�$�
��i{m��T��;g	�M�F�D�覲!��
�pG�]�&U�s��a�-z֎����Y��rݞf�=�lX�\«��aY�@�y��qJT2�/I��u��;��͓����|=��j��b��nY*nP��a�I�G�8Ũ��.�n��/�ρ̛A�ɷgЁ��j���Ӻ>��zx�х�	��y���9�긯����#z����	��]
�/i��[Ϲ`��̦D8M�t6��z��~V����#W��S 8��hE|�ӑ)Q��iGcM^0ܣ��Grc������*��]ͤs�ׯ�7*��ɚ�c'2t�k ������%�,N��[�	���_J�I4sVk|��DH�J�}T`J��<?J,e�L�"K��CD��,Ä0�ho~xs����ӡF��{�&�?"�;!d���ߢp�Rl#��#�a��0����O����8�*WX�/uηGc���b�z"�4��5���i'��� u<M�!+��﨏x���g��N�j�KXg�ʐ��Y�N���((�pQ����5�!W���,'�D��A��\�_
{󱜎Ъ���R��,����3�Ws��W�z�MY#_q��W��I��:����V�{����1˹���}.�������ོ�ƭyv�쒈|`a�F������F��(%Y����PIM�d�N�'sa�R7M2��B2�i�����������'�H��c�&���.�2<;�[�ry�Lؚ���R���t]�^W��+�n��8Ztu��5T./EY�A����,:�Ʋ�lGPF��~y?~�Lᓩ�ZP��둸�A�e4����Gg&�݀�>ܞ$J�qc^���@2����n���@��O � 7���_����oemm��5����^&\2������ �D;W���n�4S[\
��-wJ�,q�����;='���/Y��/�2/(�l�!cT�rx�,�ʔ��� SU�S!c`��H��y6X�؆��@��^��2�߼"��y�����í��0�#o���F&5���'@�!9�9ξ��<]W��>�j��{�Iss	�zT��lDj�ą��'�VӍ�b�v���*�M�
�k�]����֨<	��j�k���I��*��	->kz4��K�G��\�w-`��k��X��S�?
/�@�E&���������u�2e�;�!K3 �(������+osC�����������q�6�}Z6�R������9�*%����������^���h?OPU
�Z	u�x�#'$@�v����fgiփ�/�W���t�{6R��xϞ��a�(1�C����!r�����]�P[ 1��D�����j��߯D)�~���$F?�
���s�N�����#8P@�nz|��7>�8���@�^��?
�W5� �j�Q�*cA�����b�2i�&�?.�T5.M������i����ʄ0��-i�`>�������`�Ҧ�$E�O[-����.<�7�4U�-u��[9���5���q��
�߭4��C���̪^��M�i������/��!�./M"1<:��e�����?��3�<Ʌ��a��Xt���cOj����ިz����B�?���R�h�^r�_"[��aIE�4	�Ѐ������1"��̯�JmCD{un��D�ʬ�D��JT^���η�]�4`�rN\�g����5V{A��N4i�&A=�o_�G�1`G�;��q5�Goal�2~ַ)���Ł���>o{�� �@�E�W%1!����ֶ�R�e8T�Z�����P�̕�O-����{J�$��/��Iۏ68ieÀ[�u;��y:`�������Ʈպ�'_�T�yŁ�z�e�sR�k���i���^.a:��M�>�7\���N�j���W	N����mg9������r"y�,؜7�ٮx�t�҅��>�kt���ԄDe�Z^�2��be?Ǯq��Ȑ~�9�	�0te�;P޵'��C����;���?���Γ��VH�G�,��7�%ɴ[\�~jb�~c3ެ�pϽT4Y����O-�������?�E�����Xa�i��cț�d�#@�f~��l@1m��ؖeRL^�O�77�bI�M���vAO�z4b�l0���-r^����g��B}��a��5�q�Ȇ*�x�+��6�5x���JI�����sw2v�gY)]��g>��|f6��B�,U��%��%�Af�%v���ٷ�]jq59-�L�
�5JF�:Ѧ�T��R��d���� #����@q*�&��vNʰe(m���B��)	�M�8��{�6�:�?����אT�י�y���K���!їH���	$�͛NP{j�Wg��r�w-������ٔ�����}�@�0��L���S�:S9R|B*I^ڶ@�QG(���1�"tlK�y����£V� ��Wǂ���orz��jm��Qѧ'�|�����Y&)Z��c�8׋�������b����0w�H��Q�7��J�/ʉcQr�\q�6)���-�r%B$W�3g�W?ëԘ�R^���n�Ѩ��HM��r;�8�d�� <F~ѵL�`m�(q�ƶ�P���^��r^ hZ��8�J#kugwS�*o���A�<���׭�`bb���^pC���З���=Ffj��"Smc��>��!��g���o����VO��9�"�8�&xj%w�i�ەǐ��) Y@�tk� ��d]Κr�yem����!�%��B�.O1�l}���C�`�.9�e����I�Z�m��f"���4bI��Ao��]�'�*�Z���}���"�)�p��-�4ӌ���.E��d4,%�N�6�,�Y�.��w��P�=�Ȓ^�m:��ʠ:桳K��k�N12 ��G�d���;���=�QӅ�X�z5}��8����]�{���W��RH��4px"��2�ی��.�wa���%~�hN	L:>�K�M�W�<L)c+;�������B�|��,$.y�\�.���{���߹Ri�Jld8��r�w���|���\��oj��&�H�-&SZ����9�ǌ����{��.D��οV���c	����xgbZk���Gf�4���{�F�%b��Zع�C�@ob���}eȱR�3,��ޟO8B�#��ƫ�48dw%��h�=�L�j%�;�a�gi�Ϭ�����̝�m[�o��z���3�תu��97�1�f�8��]4��[]�d'@�u����C�j��{�����Ci�����|��Б�Q���T��$'�0Q�a��;���V��:x>YvQ�A��xGEN�~v�e�e���`:5�9B.�@[��$��C����|9kj��H��k&r'����q�Ѹ��g�:��@,	Șܫ�fk�j����5=r�J�}�h�c��;��Ny���"u_!� 򒴴! y�K����<��g)cY��#�}�Rh,3�	"MF�ʟ��c��23�&v�W��h��srko?Z?Aw(c��0*��>����.tv����*E4A�/
���m��>!�(=�H#<I��;4y]	��5��	k��Y�G��cRy�$ԓ��+��l
�  f$�.<
Y攝��F��1Lj���e�
�R�q���%��yR5��3�
kj�I�����������7��]�������G!F���p���u�\�i���=��xr�_�<���c�6C�~+���ޝ�3-=v�*�����BoQơ�2���ZU˭I�"B&�9	�셏�
ω�CJ"��ègJ��w����ZEu�V�P��~�|æa�1_8<���B�sP�0��b��|�sZ6��5ʔ�;��%� !H�a�|��c�n�-�C����)]�!�t�{k�C:���_,���_�M$e҇�(_��338�C�I�1��ȵ��Gl*�4���j���=�����/�CҰT��+D(煚�|<6W��Wj�
�`�eE����F7�B[ɭ��v�pJk �BN���5> ��F�e8�;�2����p|�p�L�fv�,���zE� ��-���[�Uf�-H���
	�}Zz�ĳ��b�P��`��8и��Ye�A�ckW+��F�RC�W��o��Cl/�3���Y��"���3��ص�$�֟v��5�u;pm��T;P�8D[$Y�*�!4%[]P�/����<�5^��E���cN��r�R��G?�HlN��48C<�5�*���nȲ��h1�J$6��b�ĒW����¿�Ub��&�yᆡ\�0�K.�&?��a)s!n3P��ʐ.U���u��ڨ�y��m�2k��Z-l�K�e���,�e��7^�+�:�(w[ Z�jj�،~O��T��u���Yu�mB)d*��#�o���<ϊ���Q?�Q��<p0�=����+�KWCKhۼݷy����� kQ��3�9a?:��N쥫+oc�\�;0ȋeanAj��1������s�GvKq�a��2#�k牆qo�Y�;<[-M>J��u�(:���G�s:#R䖱Ƚ\w,߸|�@M�1��n��g\�PC�S"�� v ���~�A���*�Q���{�i��|��^�cE�ޜ>�*��ջ��Db����z�O8L>���֗�RB���Y��?�ݳj�E�Nr�'3K.[�f��LNҿ�ɈPF�0��s� ��{t�����52g��,���.��f���m�A��UQexY�]����8aoR��\ )->����)�p�ʑ��`AQ��Tˢ��R��u������^�+t�y6x`�0�,��>Ilzj�M/��:ϛx��@nք���-?��n#<�i�Oeo�ysZھ�t�,�'�0 1r	�~����s�j:j�r�+����mg`��	�%{Eۖ	�·� ��P�s���BQ�އ{�,�%[�	�	z��=�����@���YӤ:�ud�\]�Tf����l�M#�?5=�FI,���X^E�1���*�~��[����w�?�/p5��	|׸�Xu����#艤���j�"�@Zn����Of�J3�ػ"���J��m�&�Q[��Qn�Ѹ�4'�!X�Q�.�ޓɹ���Z�����tJ�a���PR�T�(ڗ���ٻ�O�	\��|��Qư�LB�{��k܊�= �@�Â��Dkr�-���Nq�ʲԉr���3|��j�kMG}n�T*�܉�1�$�n�IE��$�ְ�֞�֒�㼭��r}�� 3�ŃdU���u|�?���J��:�!rJ��r���(��9}���,ur(vQ��SM	b�'��D�Q}�O��I��u�qM�,����L�pp��e�bH;��nԳ���)�9YU8gb�quC����o:��a!��񶦿���ի�;�m��G������P $t3�0`q�;��5���+�2~E����i�o&.��ؓ�V���KX����R��c�o(IN�xM�
����)��W�|�LHaip�v"�%P~E�mC�����(��6��e)�}���?9��S��3R:��g&�(�A`�"@��,�l|ؓiD�]Ԫ5��Z�e`�U��p+�C�lJ����|`B��l������qc0[$r���;�e��7Rg��|�?A5
 E�"���z���'^P��~���I�~ǚ~B�Ƨ)��_DL�� �ُ`��QgpQDr�z��<5�7����a�ũ��N�G��p�y�M�TB ��cS��g$����$o�&�Ib��&�f�fv�%U�fsᦦ����p>��G�_S�4��t�!<�T�KoCtћ�����,(*_��g]�9�S�� %�l^i<�̈�/k��C�D�T�?����{���1�� �z����MN��%xO��P(�IA}&&�K��b,�~��T,�P#�� >���<ۜ.)����6�zM�0��=�k��	�W�"-�S��kMEn�N�S�V�Y�3�.Q�������g����� R���zT���X�����A�$)��3:�V��B2 ��}}�֗I��X�'��/n@�
=�x������͝I� �����O*^U-!J�L�RSu[�� �V����������A�l2���)�t���O,��]��.������2���孅���F���i�}�T��]�b:Y�
�vRK*����������n�?�����]�;���1Y3���ф�Hى���x��Ř��܎������@�K^��U����L��[?��S��r.Js��c�ï�Fڏ}��
#g���{/�3w�)��)$֪���m p)%�B�<��O|ڜ'�}��!�yx���XA4�������;(��F*X�ުI&Q�����9>GQ�2t�h���N��T���X<~���j9�������#@��o��8��6�� �U�~��Ҷ�}��-1�41@mQ1Ѣ�������i`W�nF�zҡ
���̲Q_ڌ�f�{M�NIo���H�]x�U$~(����<a���m�@��A�]0\�����f0R�3z�7��qU���&f�*�����O�F�_5X��VA>��=
�I�����;�՚2�D�����{&�~�*$U�Q���v�NL�\���s璵O��,?�%��_���;��!�#�?�P��'r-4*����?O�?���$'FkQ�R��8�����=��OCʣ
g�Hl�!|ckhǃ�<:3�ìhֿ�.�"�%S�e�`��t�H}#�+�� �ۼ�&�Ha�2}��!y�
T���)����}o
R�<b�jZ=��d�G�2�I�$�p|]c�"bo�͛��߫��/g��B0�����M%O�OC�+5|K@"����!y˺}���&g�:,����@.?/���ȼ"���t+��/��x��/́�ȴ�w�3��v���-�C�^��Ӟ�W�c}��W���Ux����$|���Zg߉n�Q���\C�%�i�+ol�v
����U���0O�˷�E��u����v�%W��Z!���z��k��4��p��-� �ϑY'�V�2{z�ᎎ���,!�ǵ��ȶ�h���+ߠWO(���l�t�R��ʇM�'8[�Z�5r)����C�mM�ݛo�����&[ι�{��N��1o���a���O��֨�[�mVz>��r�a1���!�E���\�n��u��'#7����>ݡ3)�+]kyT�)j��VI�l_�A�/}۰�}�D��$���Yx��{I�P���'�'��<�ۑ�1O֞[\4t|��u�G����_�������D��4��hD��;4��,O���d�B����7z�Gt�J��ٮ)|Ҏ����H@v3j�8�<���I�z�����=�0���ނ<{YY����~e���E(�d�6,��ǃ��s����k�ق�.疑������&�
�#�$=R�+�n'd�1��ì��;�a�5��0�+�/0̂
PwW8mZ�UyUlB�";~�V��Z1c�۳w.|q=[���rמ4K���/ak�螚�~�nH���ڗo��&m��	�Pm��PI�ة;7��h:gh�.ԃ?1��ע��M�z=�<IFӪv~V�rZ��z[�wӐ��C�d��Dc�#���?���泰��ލ������Ɣ������N�飃�n��ǫt�D�y�P.��c�,)�q��W�^ZYy�u������r�]I�,ӂI�c��%��ލ�㬺f?��V����w���:#�г��:Ѷo�AR�����-
P��.;��ZO2��k��Z��ֿ� ��\���663��G�xy����Ǎ���X���[��MĞ@�Y�ЯHhy��Ώ3��$�:ޚ�ŝ����@ᒊ�N�M�Q4�����G����?�Z�+���Z��-UTaj��	��uN�\BY.0�^G�kG;��P�@�m�{�h[�xm�a8+�A3^�'&��-��t��"&6�l�B�����QEo;E��G��Thu��_:������"� �0��6� �l�Hf)�{G݇y�Ù�>{qJ�@��X}��zwM2n�_�2���6��[\ۏ�
�(��2u1%_����1 �����"6�r�$2�,^�< ��9>�:5�PK�w�]���m��~��Jt��Q���@����{�&z�b�h��-2%4.dK*���}��y%g��{ݢ�X���LJ�2��f$AwC�Ȉ�R�ei[�\q.���(�/Rց	��^EZ���_ͫ�9���'��Q�xa�<e</ϴ�I�ּ�N�������@�Cbk])��1��+�/�#�=ve�0�-"�3��d~��%�υJ|�f�M��'�U�5�s�2 ��$��M#� ��k��t0PN}$!�=�a0 �,�}��uE��5y�B+��Ф��� t�F�����:I!,��ACj�NA����y�E�G������v��8�g'�G��,���X�xVe�5ۆ&ݴ��Uy�-}�}33�/8�v�q�S�J����!G�ɲ�f�dB!r�uY�ȊX��YH�P�>��_�^�K�Uw��x1p!(6�t���(��9vm���S��j�a�U������]2�Ly8aAlu��L�%_���?ޢ-��t�Ē�����*��P��Z3�q��>�p��MG�F�<)�
9��OPm���I�Ȧ��EQƆ�8C�� s=���1��n%JX�t	u���n("&������\6E�m���ls9�<�q���B���D�Ъ�JW
+B����S�n'��O�bӖɳZ��\J��bw�!}���g#�X�ZM��̛#@��}�%؆ϋ �#�]��L��z�N�v��L`�d���~�n^� ~�y�m��M`D,H�+QC���y�3y+��r�g�OL��{8�]�dC�)�~��Zr��ρ��q�R��R���Xu:k�������49׽�K����:4u��i��{�t��v9I�[w�du�M��?叝���:�',B���#)�$&�F�t�����EA��u���`�-�=1�$��a]�Xn��5-��潋��͓�A�x�9+<jh�i!o� $��ް|�%�`@�9�#���,%(�e���b���֗=1�wo�^K�����Nv���É�Q^A��DO3�Yh�yt4j�~ї�Ѐ�����@����d�~\��PV�T(�1�2_�bh����W���q��r}r(t�G_���:�'��T(�qH��"�8k	
j�Ɖ�V��3zw�Ad�wf��Q/�O��W���׻�7R��MY��tL]!�-����S�U���Zj����g��zAK��Сތi.Nhҷꍠ�@<��س�Z�Zwc��i���e���i�>�n�*���<7gS��M��3��ة��J��3w;j[�y��wf��� Ýl_�P���f�@&o�!+�Fq�?�X��I����Y��2iԕ77�g�C��e��X�Gn�k����?8]&3�bl�����R�y�گ�E=Uԭ�Wi8 d:�v,��{��8z��(쌼ݕ�9,a�L3]�¿Q�6��d`�R���nA���~��)
N�vo� 7�f� �tKO���>��bF-�i�:���Z��0���mG��S�� ��-�B�I�i>�g�[3��X������k���.
�i5�'�qR5�I�#\@�����.��4�μ��Tbl��ѓMaf��{p,\��O��=����oi�t��xԗ��3��G�|r���� Y]L�H�6��^���ܣ�z�]���VJ?��B���0:g���LߪPK%"51�AD�kM�<��P�#��	u�ۖ����Г�� �b���T<�9�(�y8!��B#;�`x��ۗ0�z?��wuC���JMĥK��.f��h$�3Q��T��8G �o+N��`���Dہh�ܶ�:��T1d�����;����qs@��ȋ/�����p��bk�VX$ ��4l��|+:�JHVB���<uK*f����B߰�ڑOQ���$:?X�?h�_�r��@�+9Efcq�T�a�pBV�w�5MPqb���ǻ��>��zݓ7��X���_G) 2R��*�kPHX�.��4t���I���9׶̍����yW���)�d�$|��60�yF�İ7�1��Ir	�����o�]I�c k�N�+�@��{&�o�ԃBz1p3����z
6�W�;q���'%�o�⹍�'<�k���ە99SӃf�kE�V&�3�	f�Q���UYʳ��#xB��Lꞅ������9Y5d���oq91�I|oX7�����䙷�f��Jkw7ɩI/qI�b�[b�(_��J�mW	�{ ���m/z�_�j��g��)����l�0͘��/�|E��>D��[Q�����-��c�T^@8��≽E�0�X����`�!�[5�7���s7&�e�c���ǁ�L޳�+ kYۨ���DE�	��P�����`�X������R����Q�[�e�Ӟ=H
V��t��pk奰w3�rB�0���ґ|*�
�%�攏��i�^�����>`�@@��w��8��N}��c�!�H�R,�È��	?A�����¸�ܓ� l�W}�oŮ�w��%�������p���Q�=J����F,��7�M�����{�:���+����_��c�oqak;��9���W#H�fr�ؚ6��P����X�}f������`�B�s�E�w��s̭���x�!ɩ[�B0!�������/Z	o1�)>��噂w�	o̺�@�W�g31jP[<i����COc]��7�#Rm���K�L��L�̃�"0��h#"��xJ���@�"�����Vɨp�+���f-�9V��a�4��1�IaD*<�jڱ�	�{��S��nh���PF-?�r����~��j�\?3�W���tV<���$9�}wMd�Q�V�Ry�1���d�7�gmD���o�'��	��q���Xn�}�Zj�5���ů����yO�@�F0�����
�9j�g.�,>Ҋ�l�..�),iХ�E��e:����4hM� l�������9[	X�a����K�9NP���hj9�?��UX0�7mHs�j���1h�$�[�J��Jo+�ִmFZ���UJ���߼��D��u0O����lq�灇u��q����y�Em�y��nV�,���q��=?�?�� AA�:��,��^gB��5tO�&
�I�tb�)�J)��%6�ؕ��y�C������ZnoVH�/��Ǭ`J	���q5F�Ň��AU����〷6K5L�.�c�h_�+BwCĵ�Ҳ�N���w.A��"������"�F�z��T��{��
����!2,$-wb�`�����=2"�Ӻ����ͮf�=�qq� 3*>����<���8�n��3��q�t�yh��u�eX^g��ȧ���9�Az�þD�<�B�(1D��Y��iI>[ݐ�O���~<뙠Zg�t0��.C�m���m�����+'�H�݅B��d/~�[a� 
:�
��*G�r��$�+ �����<���X�F|��M��Kx����`{��T���ӌ�j�z�W,�s����k�0��{:��qA�n�3�Oc
�1�ks��_MI:�{7�3��� �B%�s�tդCz[f�!I���r�Q�M����u&3}g�9l�E����q0�k���HhQL'��5^����B��(X�M���ybaM��q��XW��#W��T=�c�{b�{ �kԷJ��l�����<QQ��[��]!���������ӊ��.	 ���B�C��9���A��w�D�1Ԝ!m_�ϨM+���"v���-T���
e9�*�[�rE�d$��[n��5Nb���/J54�� Z�="
o�ԸF���X
����P2���O�Y��n��b�(��#�w�7�����#�-/�%)���\\���x���n�H��rdJ����!ӡ/�hs%��H�)"�w�>�q\�j/[�d' 4��:UMI͂`2}��n�9H�E��]"$��&���`���>Wy�@�<�y6Zp/7��i����$l�keX��d{:�*\E}g�D��h�bF�+�րz^jO�p&-��j��� �P����e��[Uas�v��v�H��m��	C	�	X�hfGb�7X�(MGcg$+��ń�i�Np�T>���XR���5�{��VL�iI������F6�E��V��$��H9>��g'����BM}^�LQD@����W���b�L(��*���TV��6r�'��3�Y����%����m��Tc�j0�ǟ��7��5²�{i"ءzYD��!a&3Y���a���`��b�ȥ��D���?p��Pz���>�n� *�a�%w&&i��
?���^�i1T��KDC�L�xa��#��b/��Z��J!�t��I���A��{�Y۰��Ϸ��~�ҥ�u���b.`h�u]��Я#c̵!}6g������yfM#�z��]uԩ ���+K�Kl�)��C�-B����Za�X����!h��{��ѣr�[(V;�R�[�׉5� �]@���|<s����=����p�y��m�m���(;�dO �=?Yo�����V<.���I�i�@��n�ml�!��B�/pv��y6���OK����]���w���v���_�����A��Ϯ�/�>>ޘ���[k����q�|��x�#Wl�%��iWy<��[���C]�fXE�ZPh��������tнf�_�G�*��@>�ThEc߳h|�ny�}��D��/M���r�u��j;*�r�w}c��#����u� "��g4�v:4F��H�^R9���Upxo��s^�f܋���
�c4�&�3��}�
tY����՘4��kM�w&7I
*�S�*LT��/���k(z��qP��\�'K�Xe�{%k�iG	�٫P_%�!
��چ���aX�l�PT�/�v
�he�����+�oA6!-�^�`�g��������,�i�3o�-�\F6_ϳ���p5���d�O�-?�p����[sS	�I��صo1�Io ���!:c �h���\}6%��x���E���Nɮ� ��g����&#���M������9[H&������-�[cn����r%�vX���%VE5�m���(�\fu��M|ȱ�6<��}Vdר�DOR��F_�^�ӛ�t~�_
O��E'����t�����N�W�ͳ��>q�X�v�o��,�O����������Ȓ ���ON�J瘮�$��켡�C_,B�L��Y�a{�+�Zé��yR)*�����B8�i���!TĐ���|՛��_��~��Xaֺ#:��	j7e�$\�SȨ0lڐ.e�����a�'��vl�T#6m�o�η����/4V��.M���/�h��+��G�a����(t��f��X�^}U'��!t�7���_��.��r�=�4�=q<F�I�Uڔ/m4���Z�ȑ��x, ��|�5�/�-��	���k�B@�&�7�/u
��F�u����;�dD8�Cuy��v�j��~�7��[�p�p���\}�@yM^�v��C�j�'�y�J\�ʴ�F#69f"݌k5ɑ����'n�z�|DJ��=W�	���n=���'B.�c������B����Oc�����q �h��͐�^�a�"J/����{'�@�@$�D6�k�k	y�c&�[�GMf�cM�hw�,��(�`��f+��d�����4�&$���{/�#��ɣҒ�e�WH��2Zj�֘`O�S�r��3��ݱ˗��)�{6{r�����?�O��ˢp��+�n�_0���kW�5���-mR�J1'�J����*�R��2���_S��"�v;����
>�x��v!�@%z���j�u��,��P��`j�`(/X� �]���ӕ E�/I��J:g�����������>�"t^oiV(���s��|�0��dl��p��qC��807�3�b�ƾ�G��._�@z ���r��{����/G��C��N�0^w�+vT��b�Ӛ�<�i��׆D_p�����y�eܢk�D��+�m&�Rlf�~!�j��S̑���Ǥj,H/��MU��jK�1�O&5ƕ���l2< �*8�� H�M4�ߔ�4C{��	�=H���5����|�m�y�bI�!|���@�Gb�wa-e�9~w
Ij$M�K�6%��ɵ^��Hzqkp\�����0�Ʉ��B4(�Oh-�d$P��u�����^i=&>B'���S�<��܌��5�s���T���O���N�Lșd"f�oG�k�M-p��fBM~^cg JL��؅w�c��5��m������朷��/1=X�*�]>���G=�}�X:�l]Ѐ5S~��_-�X�tf2���6����u�mr-�=�#7D�?�-b��=�\�Y���^;ח!׼TI�K��<c���d]x����C�5J��_�mCB�Q������8�O���ݫ�@X��y���RS(�1-��_]���;k��8���؞����  ��ov�g^iQ�Ɛk�	����ˊ���i��r
�h��=�e*�����n"���&`�F8�����Hl�N��=D�(wwdW�,��ʲ�������s��0��+P���&�`��ɐ �/�)�
a��S�C��紓�J68�90�9f	t�؈���<�SY��UB1��ޟ|��8N79K�"=�O�=��J��9@�B Xz��B2�.��t���P1XjC)3��-�II������'��C�e>��c�0(ӿ]L@�k'W����V�����	d	*%`^+樑�6 ��}�l쮢����k/�=>��Xc^����������Sr���A0r+&@2lkx&�K�����"��G:w�A�7;:!��\�����:{ǖod'N00�b��	m�A�+��$՚S�#��<vjc�v�gC`^#�4�ј:[.���<�������p�=���>����8c�vů�Sڣ�V����86NI�	��Վ�~���x�B�f��V$��X5��w���7�v�˧�H�Q�fף��]|x����F���m�a���}9&�ӳ�I���sp����p����.��Z��GrG�!JqZvs���%/��0���Z�HOn�p]ɩ�"���aP��b����V��x�j�E�'���Qw����żƵ&�9�����j�$H���'�S�YaR��p���?��30�Y�U��)k�|Pan�W��	��B���3M� HA��f�5Yi�.��M����noO��F��o\oPl:.�g��-Du�7�����*�'�&����*1��'~�ŉ�u5����4�2����g	?F�m��˺���ww�H�[>\�d�Z�
�*nW�Z��ؕ���u����\�[�����6���+H�vS%�5.�N�@�g���S�'�Xʟ*D���8������n��h'�o�9OZ�}:Er1]>�C�lt2��`>��L2�b8o����N�������q2yreLd��2�i['���_թnd��O�{�zh���9��J��٥򚧟�=��ާ������>+���m���H�(��Ӱh����'
�D�7�ڔ��:-Xg_s��P�c��Y��>0����V0H�k*�|{3H�Ef�l�'��E-?S�8?�T����x_�p�&W$�WY�"���+�hl�b���?��11��_D��!@�U�
���F��)e��ҞѬ�vBʙx�gЬ�:-�e(W������o���p4_vl��|=�{+��ė�J�M<8�J��7<�v�\��� �!J�;d/��bc�|w�`I~6�96�b������B��č�RZT@UR@�T, �����eI�?��,�C���vz� ��>P�'�_��]��B�VQ]�r��Oc�������Km��y�7NjP��U���"@^��JĈ���OC�­7"�[�b1R#@����	���;��}@jU/�K�,g���0���С��C��m@�$*ZH	gC���OόN�������6���ů�O7�^�	^��++���*�+S����~ϕ��\?�Z3$fPH��y�T�r3�؋��`���◚�X�'�x��9��(u��K�Tu)����j�A�v��k�g���y�L� �
/�çLĞ���/~"�n��d��1;���H�1g���(ض�"�	��oS����2}=jb���,wr7,�Ȑ{�d޺V|;y���}{D�B�Up�U��U��%mB���kx�x&-l6l��ׇ�C,7 ��U.�͏m!��֑�m�P�ԉ^Y�*�`�T���tGi�Vm#��X<����K�u��1�l� 7��t����^�Պ;�	I�9���d�e�PW8�+� �]��\��E�(�k�����f��QE��0�Q�G����^�sA/S޺�۩��^v���6�.�w��fݮ�@K�S����>�������
�a���R,�
��ك���	R�!�V
������0f��6=v��睨� [�y�MIQ<q��Opg^N�k��T/Om�� {���^�	�Z��H�H�UVQg�
C4�SS����~0�:H�:b4#`̙Bo?_E�B VA~���Y��h�AF3Q�X����܈������X�l���L
��]��|�8�z`�ݘ^����/��%m�}��	ᅲH�㣰����]��z�Qe!Z��e�w��bX˱j|{N�(J�w��H�w@Qz�dqeX+��7�o5s�N�y���)��̉k�OL,��E�xRb\�qv���u��Hn��*��lvN�.ґƔ�ݨ5OG��H���i����W:�����y��n`ɍ�<��eOZ����4}�1�h��޴9L�PJ���I��8aw�+��s8mZ�ŵ���~���֯��Ȝ���S����Os�X��,Fo��ׇ����~�6�ʈ�jNd�]�!�Y����˄w����ơyp�b�GX�5 �HQ�/(<�`#>��R׹�6QUg8�D���'��XJ��J<@�%~"m�cQ�&�$@b�
C,��Ƞ���]���b�"&(J��o����z�,V��i�w(�}L����D����`�!!�������j�)��|UT)C+e���s6����7��]x��C8�A>��sCW�4R6Yih���R��8����s�(�M8�H���C�]�z��1\��}~D(e+b:E�`ʲ�{[�|�����ъ2C�H΍D�?���2���	����nh�fՙb\%�Hq*�$��|����gu}� ���W1�If��F�EU�a��ɦ���gCҤV��.�P�!�H��`\A�}<��v���e9�QV��n���E��΁��OX��������)��02*�œ��Z�(O$L��5��ڇtqx^, ������2]�V����[�Ȑpx����֒���l�+(+0��g��q���,RY�9	�ӷ0'r͵G����ϲ��
6׭H;J��ɶ�K�>v3�g�d=�R���±]� �q=��]�gt�M�Q�o�m��:����ϖF�>�$�q�^$xq�UeQ$�#Í�$��|��C̘B8_�R�EԿ�6iƾd�	�k��>E��쵍��Zq�B�?Y���V̉�:���&ASy,qHw>PA��I�
�Q_rP���z	[�O��c�"�a�s�0�+�j�� \XQ^M�.��m�|�u��Gb�s=�Mׂ�2������Н$� '���o���c4/]�UD,�P��,9�p*h8N+	&�����:�e[�٣�s3�����i�
Ѝ
��,��*w�c�A���Lv�Z��HA8�J0�6�ՙ�@o�R!v�� ��:+u��GwJ�i�]�����Z�y쭊^�,��Q��a��:Ձ:[�^"T���S����%�h�X�,1ΔYf/z�!�{H�5:3��Y�l�s�2����֟�@��n��8����j-�p�Pa��Q�`o�9�|�4~�k� �w��{�R2�d	�缮�
��V��$�T&:�W�oم|�����MN/5@C��4��0�=����*m�ѐ�f^һ��^CGV�U%n�@=n��c��,�z{b/WnC����R�Ͽ����"ym�g�f�3��x遰	��sƨ[��t� d�K�;{�%�-	s#���Z3_�4�iȮ�
,�i�6_LǒX�V_��,f������)�[��� }�rט��b;��Ř������
���B�C��G��`��V��\��C���'�,dަ"���T��7d�V��<䈔��h'/�@N���h:�i1�8&��p=����[�|�a��I���v5#.M՗s���$������t>^Hlu��:d�V�뷶F�M!`�.��d�`�/�&�n�a�hP>>���%���S4�E��T$ytzQ�|�z~�ܟ�������, �`gb+M�2�����u쾀/�x���������XP^mx����B�ySf$G�qc�����A8��fU� ���z��q�[if��n��6�́��""���A#��ŠZ�f `�>�&���B�Nu_\�*�'^�H8���L �M}d��y��g���D�HK,�*�*��a˪��-hW/&���yt�)`�ֈ/f��w8��lE��D%�k���������Bs¼�����zhZZ]G��G�i̲M�#@گ�Go��B���*�ܒ��>`$58����k��Y#��J�l��	���wR�Ҏ+P�kr��W64gA�Uy��mPG�w����!�$��!{d:19���'����q�؍�(�>-v��c��>����+�5<��S��/���ֈb�`��)�w&�u�'xÃL2$]�ϖ��yG�-
�Q��g*�
WX��O��i�{��ىG������M/$��+V��z�R�񞤥[��DU{3�7K�O>A�,Ep�V�9�\�㈸��*�����'oB�0�&�U�d kͺ>�{�v�/��	q����?�J��L�9#����ɤ�Yi��;#��<�>��1t�P�U6h�}	ͼ$T��S�O�(S��It�7#���m�,�z�2�������K�/���]Sb�$�������;#�ؽ��$d��]H����e�f�ϔg��P��qv�=�~"��s�;���P�� ��uP�%�~W�ˡyn:<����������[E�x#��D&g_�Ȏ80ѯ��tG<�h����s�~��L�LJ!�K'�cc7�養�M+�;�1�w�P�>��A�[[��Mt��5��Z;x5���ۻ�vv�e�Z��N�/�aou����0u��A�wN�z=i����'�#Eҥb�F�&����L'iJԝHf����
�`�nt$n��^�������	���賓,�k�}3�@Q�[=�erL�o_7�ٶ���  ���F ����؋��F �C��z�����F ��  ����   ��������7  �������  �������   �����@�v�����  ���   ��$  X���  �P�F ��ŀ  ���	  ��x�����H  �������5��F C���F ��H  �$�F ���F �   ��	�X�5\�F ǅt���   ��  �։0�F �\�F ��t����$�F ���F ��H  �0�F ���<��x�����  �$�F �p�F ��H  ��	$�F �$�F ���F    ��F ��x�����F �5$�F ��������x�����F ���F ���F �������Q���F X�����l�F �5��F ���F ��H  �X�F ���F ��|�����F ��H  �5l�F �5X�F �5��F ���L  ��F �5$�F ��x�����F ���F ��x����>�����x������  ��F ��`  ��|  ��,  ���  ��,  ��H  ��@  �X�F �=�F ��H  �Ë��F ��  ��d  �5��F �   É�H  XC���F ��H  ���F ���F ������X��F ��d  ��$�W��F    ��\  ��H  ǅD     ǅ@      �X�F     ��0  �x�F ���F ���F h�  ��  ��h�  �5��F �5��F jj ����É��F P�5��F ���F     ���F ��x������������F ���F ���F ��@  ��x����X�F ���F ���  ���F ��  ��  � �F     X��������  � �F ��  ��@  ��x����X�F ��  ���*  Q�D�F ���F P�������=T�F ���F ��x�����t����=p�F �=T�F �p�F ���F ��@  ��x�������  ��\  ��)��5|�F h�  R�6   +=��F �P�F V�5P�F ���?  ���F �4�F [��\  ���F 뮋5��F 3�$�  )�@  ��\  ��3�$�  )�+�$  ����)�$�  �4�F ���F 34�F )�$�  �4�F ��3�$�  )�$�  ��\  +5|�F ��@  � �,�F jh�  ��  Ã�����؋��F ��d�����F X��H  ���F ���������F ���F ���  3��F �[�3��F �=��F �<}    �5L�F �   ���P�F    ��\  ��j h�  j������J���������ǅH     �5��F �54�F �5��F j<W�?  �P�p�F ���F ��'����p�F �+a���p�F P��H  ���F ��x����������p�F ����   ��H  ���F ��  ���F X��������  ���F ��D  ��H  ���   ��Sh�  Rh(#  �  Ë�d  ��|  ��5��F j�54�F ����Ë���؉��F ��H  Q���F ���F ��c��S��x����5�F ���F ��������p���Z���������54�F h�	  ��  ����  ��H  jjd�����É�\  �,�F j �5��F ��  Ë�h�  �g���É��F ���F �� �$���S���F ��H  ���F ��x�����������H  Z���F X��  ���F ��@  ��  ���`�����H  �p�F ���F ��������H  R�p�F ������?  ��  ������h�  �H����ǅ|      ���F     ���F     �5��F �c����Sh�  �����Ã�������4�F ���F �5D�F ���F ��\  ��\  ����   j �������\  ��$D  ��4  ���  ��$\  ��  ��$H  ��$D  ^���  �5`�F ���   ���g����ڋ��F ��H  �5$�F X��������  �$�F ��  ��  �5$�F ��D  ��������������  ���F ��������H  ���5��F �5�F Q�����h�
  h}�E �5`�F �QP�����,�F ��X  ��f h�#  j ��$d  ��  �SU�����,�F h�  ��X  �5h�F ��|  ���F �ҍ,�F ��l  �������F �,�F ^��d  ��|  �4��I��<  �4�F ��d  �1�1�I���c  �UW  �\�F ���F ��|  �5L�F ���F �\�F �)������F �,�F �$�  ���   ��� ���	�A���F P��H  ���F ��F ������� �F �X�F ���F X�X�F ��F � �F ���x���P��h  ��X  �4�F ���F ��\  ��\  ���s������  �,�F 8�5��F ���  �=,�F �5|�F ���F �P�F ���  ��0�  �5,�F �X�F ���  �:�0�F ���  �@���"  R�0�F �X�F ���"  Y��,�F ���  �5|�F S�f���Á�   ��o�����  �,�F �� $  ���  ��P%  �5P�F �>F���   ���   �`����=,�F jh�  h�  j h�  ����Ëx�F �� �G �5��F �  �d�    ���F �	d�    �,�F ���  ���������  ���F �=�F ���  �8�F ���  �=8�F �,�F j ����Ë|$ ��F ���F �5��F ���F ��F �-��F �=��F Z�`�F �%��F ��F ���F �-P�F �5��F �=(�F ��P  ËP�F A�58�F h�  �����d�5    ��F �d�    ���F �,�F ���!  �=�F P���!  �=��F ��<�5����P�F     �,�F     hp  �����Rd�5    d�%    ̉��F �`�F �U܋]�U���F �U܋u�5l�F �E؋��F �E�E��(�u��5,�F �]�M�ǆ�      ���  �M�`�F ǁ�      �M��� �F �E�    �8�F     �u�F���  ������=,�F ��  ��`  �]�C���   ���   ��  �U�4�F �=8�F }�U��4�F ���F �=8�F �M���F �]���F �d�    �d�    ��,�F ���F �-��F ��p  �=,�F ���'  `K�^��l  ���)  ȋ��'  ˋ��F Ӈ|(  ��F 3�h(  ���F ��h  ��|(  ��F h�  �5�F V�54�F h�  �V���Ë�$�  ��$�  ��$�  ��$�  �X������F �U������]܉M؉}ԋދ`�F �}�=��F �}ԉ4�F �E�T�F �]܉]�ދ4�F �W�����F ���  ���  �%x�F ������  �x�F ;�$X  �������F ���  ���  ��   �  ��$  �-x�F �h�F �(�F �$�F �X�F �=��F �5P�F ��$  ��$   �����Q�,�F ǁ�      W��   ��F �=x�F �`�F �p�F ���F ;�$�  ��P�����F ��F ��   ȋ`�F ���F j ��   Ǉ\      ���  ���  �=��F ;�$�  ������=��F =��F ���  ����  ���F ���  �x�F     �  �U�]�4�F ��P  ��`  ��[�Ћ�P  �&������F �`�F ���������������;��F �wN���`�F ���F �=x�F ��   ��F �d�F ���������������F S�`�F �p�F �d�F ���F ���t��P�F �`�F Q���  Ӆ�����P�F +��F ��������F Y���F [���F ��   ��$  ��$  ��������  �X�F ���  ���  ���  ����p������  ���  ���  ���F ���  �x�F ��F ���  +��F x�F ��$�  ���F ���  ���  �X�F ��F �V����\�F �����  ���F ��t  ӄ$�  +��F �$�  �\�F ���F �,�F �0�F ���$  �d�F ����;$�F ��������F ��F �=��F ��ً��F ���  ��F �@�F ǅ�      �\�F �ϋ0�F ���  �=@�F �5�F ���  ���  � ��F �]���L  XX���,�F ��*���F �,�F 3�  5��F ���F ��  ��F �%��F ��(�M��l�F �ˉ}��=h�F #��  ���F ���  3��  ���U���|  PX��h  �%��F ��̖�ف�D�q��-��F W�U�������,�F ��  ӂ$  �h�F ��$  3��  BX� ���  �U��\�F �]�E�u�}��m܉��F ��$@  ���F �T�F �5�F �=��F �-��F �<�F ��$(  ��$   ��$  ��$  �8����p�F �P�F ��  �;��F �zC������$�  �h�F �h�F ����D���ʋP�F ���  ���  �0�F VW�5$�F Qh�  �l���Ë��F ���F ��F ���  ��؉=$�F �8=��F �=\�F ǅ�      �5�F �5��F jd����É�$�  �-,�F �����F     j
jPh�  �R  É��  ���F S�=����\�F ���  �\�F ���  �5�F ��,�0���P������Q��<  �����9������CJ���� ��  ���F �������x�F ��  V�j  Á�  �M�&�Eċ��F 3�8  ��L  ��  ���   ��  P���D �,�F ���  �P  �L�F ��  +��F ����B� �F ���F �E��,�F ��H  �RWj�5��F �5|�F �������   ��4  ���F ��l   \7���  �=��F �zX���F ӂl  ���  ���F ���F +,�F ��x  ���   ��F �H�F �V�5,�F ���  �����F RPhP�F ��   �L�F �k2�������  3�X  �������F ���F ���F ��F ��F 3(�F �E��L�F �F j �5P�F �   É�  ��T  +��  ��g^G��E���K��%��F ��  ���F ��F �H�F �E���F ��  ��F �}����  3��  �u����   �E����F �F�H�F �]Љ^�T�F �}����   ���  �V�E܉F���  �^�,�F ��F     �}��] �uԋE􉺼  ��$  �5��F ��������  ���  �5��F ���  �X�F ���  �  ���  ���F ���  �X�F ���  ���  �=��F ���  ���F ���  ���  �$  9=��F ��������  j W�58�F h   Q����Á5��F ��H�l$���E���   �8�F ��X&  ��'  �]܋��F YX�-8�F ��� �F �8�F YX�,�F �]؋��   ���  ��N�\X�#  �h�F �5��F jZj j
����Á��  ����8�F ���  ;�$�  �(������F j�58�F �5�F h   ����ÉX�F ��   ӂ  �<�F ���F ���F    ǅ�      �5��F ���  ���  �2���F     ǅ�      ���  �X�F ���  ���  �5��F ��)É�v��$�  �D�F ���  ���  ��   ;
������R���F ��������  ������5��F ���%  Ή5��F �5,�F 5��F 5�F ���F +�F YX5��F +��F �UԋU؉��   �p�h�F �P� �F �P�X�UԉP���'  ��F �E���(+  ���F �]܉�8&  �=��F ��('  �=$�F ��T)  �Uԋu؉��*  ��,*  ��p&  ���F �-d�F ���=T�F É��  ���  � �F ���F 9�$�  ��S���\�F ���  ���  ���F ���  ���  ���F ���  ���  �;��F �W[�����  ��$�  I����a���\�F ���F 뻋�H  �t�F �p�F ���   ��  ��)�$�  ���  3�$�  )�$�  �=�F ��  ��1�)�$�  ��  +��F ��  ����)�$�  �5��F �5|�F 35��F )�$�  � �F ���F ��3 �F )�$�  ��   �5p�F j ǅH      ���F     �X�F ���F Z�3��F �R��  ��  ���F �3�$�  ��  ���F �]    ��  �   �����F    ��  ��������%��F ������  ���F ;��F ��`����$�  ���  ���  ���  ���  ���F �  ��  +5�F � �F +��F ���F ��  ���F ��tv�=�F ��   ��F ���F ��  ��  ��  ��   ��F ��  ��  �"�����  ���F ���  ���F ��H  ��  �X�F ������   �,�F ���F ��t����4
�
�R�=��F �<
�
�R��/ �S6���=�F ���  ��  ���F �5��F R��  �X�F �e���ǅ�      9�$�  ��W�����  ���  ��$�  �$�  ���F ��񉝸  ���F ���  ���F     ���  ���F ���F ���  � ���&������  ���  ���F +��F ��F ��$�  ���F ���  ���  ���F 랋�B�x�F ��h  ��+��F B���F ��d  �ʉ5��F ����`  �=x�F �$�F �\�F ��5x�F ���F �L�F � � �F ����F ��\
  35�F ���  �,�F ���F ��5�΁��  �*<W���  ��4
  +�  ���F ɉ��F ���  HX���  ���F ��F ��$�  d�5    d�%    ̋�h  �H����]ԋ��F \�F 9���0  �Uȉ]ċ��F �d�F �U��}��}��;��F ��5  GK����4  �Uĉ}��}��U��(�F �M��Mȋ(�F �j ���F ���F ^;u�'����uu�=��F ����F ���F ǅp      ���F ���F �5��F �5��F ����!  ���F ���F ��h  ��<  ӄ$d  ���F +��F �$d  F��d  �5��F ���F ��h  �5��F ���F ���F ��h  �u���ǅ      ��H  ���F ��������  ���F ���F ��T��  ��d�    �d�    ���F ��	  +,�F ���F ɋ=`�F =��F ����F ��F ~X���  �T�F �%`�F ��@  #�p  ��\
  �*�_ �F h�  �z���É �F ���F ��$d  �����p  ;�$�  �Y������E���F �����=�����ɋ�������  ��H  ��  ���we����F �,�F B��F �ډ�x�����ǅ     ��F     ��H  ��  ��F �Q  ����l%  A���   Q��H  [�V���F �,�F ��ۉL�F ��H  ���F V�5,�F ������L�F ��   �t��A&  ���   �5,�F �Wd�������F    j �5��F ���F     �������"��ҋ�H  ����c��Bjǆ�      �t�5��F ��������7\���5��F ���5,�F ��ۋӋ��  �C�������7[��R��P��|������  X��릍5,�F ��ҋ��uc��BjǅH      ��H  ���F �s������������F ��F ���Y����,�F ��ۋӉ������,�F ��a��C�����F    j ���F �x�F ������X���F �x�F �Ӄ�,� ����b����x�����������H  ���t�F    j �5t�F [���������F �������5,�F ��[��Ћ��  �@��L  ����R��Z��F ����  �5,�F ���F j�l�F     X�=��F ��L  �=l�F ���  ���  ��H�  ���F ���  ���  �,�F 8�F 9��F �/������  �5��F ���F �5��F ���  ��   �,�F �5��F ǀ�     j ��l  W���  ���  ��L�����L  ���  ���  _���  �,�F ��ɉ��F Q��H  ������[�5,�F ��"  C��I����������Ӎ,�F �i�����x������  j���F     ��l  ��x���_���  ��L  ���  �,�F ���  ��@�q���  �5`�F ���  ���F �;��F �����|�F ���  ���F ��$�  ���  ���E����|�F ���  �BǀL     ��F     �������5�F ��x�F �����5�F ��F��  ��F ��l  ǂ�     �t�F     �֋(�F S�x�F �t�F ��F [��H딍5,�F ���F ǆ�     ǅd      ���F ��d  ���F ��F �x�F ���F ���H����5p�F h�  �5��F �h  �X�F ���  ���  ��j S�5<�F �f   �B��d  ���  �`�F �H�F ���F ǅ\     ǅD      ��d  ��\  ���F �x�F ��D  ��F ���F ��������<  �X�F ���  �
�,�F ǅh      ǁd      j�+�����5|�F Rj �G���É�(  �Ћ񋽐  ��(  ��,  ���F ����������F ���F    �`�F     �5��F Q�5x�F �`�F ��F Y��D������-�F &	�D���  ���F +��F �5��F fٙ���8  ���F �x  ���  �7���F ��F ��<  �,�F ��F ��8  ���F ��ȉ�F �(�F 3�H  �5��F h�  h�  h,  �   �3�   ��P  #|�F ��4  �,�F �d�F Ӏ  �5@�F �5��F +�  ��|  ӈ�  �5��F ���j h�  �5��F h�  �   ����F    ǅ�      �5��F j�5��F j�Y���Ë5��F ���  �=��F �7���$�  ��0  ��h  ���F �p�F ��,  ��0  ;�����@���F ��5���=��F ��� �t8R��^�   �   ��$�  ����� �F ��$�;  ���F [�Đ   �yS��F ���F ��l  �Љ�  [��[��Ћ��  �x�F �e,����   Bjǅd      S��d  ��������4�������   ��-�����F    j �t^�5��F ��F ���F �5H�F ^�H��  ���F V��Fǂ%     ǅ�      �@�F � �F     ���  ��T�Q  �5��F ��F ���F �5H�F ��[���^�@���F �N�  ��V�e�����[���W�=,�F �x+��@���  �Ћ��F ��  ���  j�0�F     X^���F ��,�����F ��  S���  ���X���Fjǂ,$      Q�X�F ��0���� �F ���  Y�� �   � �F ��5��F �5��F �5��F V����Ë��|�F    ���F     S���F �|�F � �F ���  [��T�.�,�F ǅ�     � �F     �58�F j �5��F �   ����  �,�F �5��F �   ËC �F ���F    ��m=���H�F �5��F �h�F Y�5 �F ���  W�p�F ���F ����  ��)�;��F �  �CF���F ǅ�     ��F     �=t�F �=�F �= �F �=t�F ��4�N���jd�����É}���  �h�F ��    ��;]������}���F �h�F ���  �5��F �5��F ���  �   ���F ���  �E�$�  �$�  �����  ���  ���F ���  �@�F �5��F ���  �<�F ���  �]�5h�F ���F �p�F �@�F �  W�=,�F ���F     �F<��H|�Px���  �=,�F �B�z�58�F �rW�j -8�F �z$=8�F ��$�  �B8�F ���F    ��N�  ��$�  �58�F �|�F �  �����F    ���F     ���F ���F ���F � �F ���  ���F ��4����Fǂ#     ǅ�      ��#  ���  ���  ���#  ���F ��`�����T�x����,�F ��Iҋ�,�F � �F �F��$�  �ܬ��� �F �B����]�EȋE�� ;��F ������E��E��E�I�������U��щ��F �]�ǋU���F 9��F ������=��F �p�F �}؋��F ��F 딋5�F ���F V�H�F �<�F �5 �F ���i���Q���  ���D �5 �F P� �F � �D �}� �F ���  ���  �5|�F �h�F ���  ���  ���  ���  ���  ���&�����F �5 �F ��������$�  ���F ��$�  �|�F �<�F ���F ��$�  �A  �P�F ���F ���  ��������F @���  �=��F �=��F +�$�  G��$�  ��$�  ���F ���  ���  ���=��F ���F ���  � �F �\�F ����F ��j
�����Ë��  ���  �  ��$�  ����F �$�  �$�  �%��  ���  ���  ���F ���F ��$�  ��$�  ������%���P�5T�F ��Y�0�F �@����$�  � �F �����?�����F %��  �=<�F ��+�$�  ;�$�  }i��$�  ���    ���  �5|�F �,0�$�  9���*  �5��F ��$�  �l$ ����8  ���  �H�F ���  �U�h�F ������-��F ������  ��@�`�F ��F ��)�@�Ћǉ��  �ʉ5��F ���=`�F 󤉍�  �(�F ���  �5��F �5\�F �7�5`�F ��V���F �,�F �5�F P�D�F ��  �&  �5�F ���$�  �$�  �����  �=d�F ���  ���  ��F ���  �=t�F ���  �ˋ�F �5�F ���  �5��F ���  ���  ���F ���  ���  �   j �F<��H|�Px���  �=,�F �B�z�j�-l�F �j ���$�  �R$�$�  ��$�  ��$�  �K���$�     ��+  ��$�  �   ��$�  ������x�����$�  �5|�F ��$�  �������F �ы=D�F ���F �5|�F ���  ���  ���F ���  ���  ���  ���  ��$�  �-��F ���F ���������  ���  ���;�L�F �  �식�  ���  ���  ����  �5��F ��+l�F 9��+  ���  �5��F ��    ���  ���  ��;�$�  �y������F ����5��F P���  ���  ���  �ҋ��F ���  ���  �5��F ���  ���  �0�F ���<����=�F �Ӌ5��F ���  ��F ���  �j���  �9�p�F �L�F ���  ���  ���L�F     ǅ�     ���F     ���F ���F �
�=,�F ��F     Ǉ�      ��F ���  �=�F �)��$�F �8�F �$�F �5��F �5L�F ���  �8�F ;3�&����,�F �[��$�  �M�����`  ���  ���  ���  ��x	  �������  B��$  ���  ���  +�$�  @�؋�$�  �0�F �ˉ5��F �����  ��  �x�F ���  �5\�F �7��  ��P���F ��`  �D�F ��h@  h�  j WV����É��  ���F ���  ���  ���  �5��F ���w������  �:������F ���  ���F ���  �	;��F �v�����$�  ���F ���  �5��F ����������  ���  ���F ���F 랋5p�F ���  ���F ���$�  9�$�  �W������F ���F ���  ���  ���  ���F ���  ���  �A������  ������  ���  ;��F ��?����$�  �5H�F ���  �5��F �   �5��F ;58�F ��o���5��F 5��F �P�F ���F ����F ���F �5|�F ���  ���F     ��,  ���F �P�F ���F ���F ���F ���F � ���  ��0  ���F ���F ��8  ����.  ���F +��F ��F G��  ��F ��8  ��0  �5�F ����   �$�F �,�F ��$�  ��ǅ�      ���  9�$�  ��;���5��F ���  ��$�  �$�  ���  ���  ���F ���  ǅ�      ���  ���  ���  ���  ����H����\�F ���  ӄ$�  +��F �$�  ��$�  ���  ���  �\�F ���  뜉�  �58�F Vh�  j �5��F ����É�  �58�F �������  ���F ��8  �5L�F ���F ���  ��  ��$렃����F �����   ���  ���F +��F ��F FP���F Y���Ɖh�F �`�F �%��F ������  ���F ;��F ��8�������F �=��F �=��F ;�$�  ��:���=��F =��F P���  �� �F ���  ���  ���F ǅ�      �(�F �=��F ���  ��F ���F ���  �5��F �  �%��F ���R���F ;��F ��5�������F ��F ���  �h�F ���F ���  �h�F �U�h�F ��F ����Q�,�F ǁ�      ���F ;�$�  �����V�5,�F ���  ��  �`�F ���  ˋ35 �F V���F     S�`�F �5��F �u����q������  �`�F ���  ���  ���F ���  +��F ��F F�����=,�F ���F ��  Ӈ�  +5��F 5��F ��$|  hp  SW�5��F �d���É�$�  ��$�  �%��F ������F ���F ;�$�  ��R������F ���  ���F ���F ���F ���  �  ���  ���F S���  �h�F ��F �C������  ��  �L�F ���F ���F ��  �%��F ������F ;�$  �{\�����F ���F ���F j �58�F ����É5��F ��8  �6���$  ��4  �5��F �5��F jj
�����P�<�F ��F ��F 9�x����8i�����F �<�F ���F ���  Z���F ��t������F ��   ��F     ���F ��F ;��F ��5����F �F ���  ����)-��F ��$�  ���F     ��$�  ��$�  �-t�F ��$�  �] ���#�����$�  ��$�  �,�F ��$�  ���F ��$�  +��F ��F E���F �,�F ��$�  ��$�  �-t�F ��$�  ��$�  ��$�  ��  ���  ���  �5l�F ��x����;��F �Ud�����F ���  F��$@  �5��F ���  ����d���5��F ���F �5��F S�5l�F ���  ���j �=4�F ���F �=��F ���F 9�h���������F [��h����h�����؋(-��F �-,�F Ǆ$�      �e  ���F �,�F �-8�F �����F     �5��F �5��F h�  V�  �d�    �d�    ���F ӫ�%  ��F +�D*  �`�F Ӄ|'  ��P)  �-��F ���*  ��F �X�F ���&  +��)  ��|'  ω��  ���F ӄ$�  j
jdW�5��F �5��F �c   �;8�F ��z����<  �,�F ���  ��F �|�F ���P  ���F ��8  ���F     h�  �5��F ������p������{XCX��F ���(  ���  =��F � �F �=�$���&  Ӌ�*  Wd�5    d�%    ̋�$�  ��$�  �,�F ���F ��   �(�F ���F ��$�  �����$�  ;�$�  ������F �D$��-��F �쉕�  �U�;�$�  �����U�U��=��F ��։��F ���F ���  ���  ���  ���F     ���  ���F �=��F ���  �Ƌ��F ���F ��  ���F j h�  �5��F �d���É��F ��$�  ���F ���F ��$�  �,�F ����������$�  ���F ��F ��$`  ӄ$�  �=��F ��$�  +=��F �$�  B��$�  ��$�  ��F ��$�  ���F �=��F ��$�  ��4  �,�F �%��F ������  ���F ;�$�  �kd�����F ���  ��0  �5�F ��<  �5��F ���������x������F �މp�F ��H  ���P���F ��x�����H  [���F ^�CH������8�F ���F �u  ���5��F ���  pX��0
  �3��  ��F ���F ��  ��t  ��(	  +��  ��8\q�L�F ���F �%��F 30�F ��t  ��F ��p  �,�F ��$  �5��F ��>���$  +��F �=�F �=,�F ��l  �L�F GX���F ���i��0  ���F ���F ɉ`�F ���F ��_X���  ��4  ��F ��p  �5,�F ���  ��F ӮH  ��F NX� �F ���  ɉ�t  �t�F +�
  ��|  ���  �ȋ�|  ˋ5L�F #5L�F ��x  �,�F ��L`���$�  V��x����8�F �  ���  ���F ��\  ��T	  ��F ��sX���F ӣ�  ��X  ���F 3�  ��T  ���
  3�   +��F |�F �8�F ���F ���F #`�F ��F ��\  eF�=�%��F �Q���4  ��\  ��F 3�  ��P  ���F +T�F ���F �8�F 3�`  ���  ���F Ӄ�  ��L  ��F +�(  ��0  ��L  t�F CX�s���  ���  ���  ���  �=��F � �F ���F ���  ���  ���  �=��F ���  � �F �-��F ��$�  �5,�F ��$�  ����R��  ��H  ���  {X��l  ���F 3��F ���F �%��F �\�F aƎ��D  ��|  3��  ���  ��|  �,�F ��$�  ��$8  ������  ��F ��F ���  ���  ��  RA�3  �x�F #�  ������h  ��F �%��F ���F ӌ$�  ��P  ���  ʁ��   ���=��F =��F �,�F ����Q���d  ��h  ��F ���
  ���	  #H�F �T�F ���F ���F �,�F ��F �%��F 3�	  ���  Ӄ�  3��F ��T	  d-�\���F ӫ�
  ��`  ���  3��F ��T
  �5�F 35��F ������,�F ��������H  ���F    �ʋ�T  ��������,�Aj���  Z���V  �,�F �������5P���,�F J��D  ���   ���F ����j �5��F ������[�I������5��F S��R��  ��C����F    ��  ���  ��������  ���b���ǅ�     ��F     ��F �;���  ��  ��T�F     ���  �(�F ���F �T�F ����  �T�F )�R���F �u����T�F �\�F ���  ���F ���  맍5,�F ��H  ǆ     �ˋ@�F R�������  ��x����5\�F V������,�F ��ۋˍ5,�F �B���A���.L����x�����  ��H  J��  ��D  ���   ���⋽  ��  �\�F     ��  �,�F ��ҋ�^�A���   ���#���VA�����8�F �-<�F �t$��D$����F ���F �=,�F �t$����F �|$Љ5L�F ���F �T$ȋD$��|$��l$ԋ��F �|$��,�F �\$������F �0  ���F �=��F ���F �\�F ���F �}ԋ��F ���F ���F �   ��ҋ��A���A��x������  ��H  ���1L�����  ��H��D  ���   ������  ���F ���F     ��x������F ���F �Q������F ���F �M��  �E��t  �=,�F �E؉��F �M��E�    ���  ���  ���  �A     ��F �J<ыQ|�Yx�F ����8���=,�F �K�{�E܋C���F �C �F �k$-�F �D$؋C�F �-��F ��U��Y  �MĉE����F ���F ���F ���F �Eԉ��F �\�F ���F �[����Eԉ��F ���e��ủE��Eԋ0�F 9��I���P�F ���F �E��P�F ���F ��(  �R�I�Eȁ}�    ��7���p�F �ủ]��M܋]ԉ@�F �]��=��F �=��F �}ԋp�F �=��F �Mċ]��u��N  ��F ��  Q���D �u�P�E�� �D �M��=��F �5��F �U���  �F���$�F �E̋�F �UȋuĉE��=t�F �U����F �U��=�F �}�=t�F �}  �5@�F �E��E�    �u܋E���8  ���F �Uԉ��F �,�F �@�F �UԉE܉��F �   ��Mċ,�F �   ���?���Ƌ%��  +��F ;E��4���e����|$��   ��A��F �}���+u�F�ƋẺM��΋����=��F �=�F �U��E��}����F �5h�F �5x�F �7�����M����u��u�u�uċ����  �u��]ԉ�F �Љ=��F �u�� �F �=��F ��F �/  �l$ԉ5@�F �\$̉L$ȉD$Љp�F ���  ���F �    �<�F ǃ�      �|�F ���F �L$���F ���   ��F �Q�5 �F �q���  �i�Y���F �A�  �8�F �-<�F �D$̉|$����F �ËT$ȋ\$̋l$ԋ��F �|$Љ��F ���F �8������F �u��5��F 5�F 5�F �%��  �}ԉ5��F ���F �5��F ���F �����L�F �,�F ǂ�      ���F ;��F ��  ���F ��F �UЋ�UЉl�F ���F �E��$�F     ��F �uĉU��M��5L�F �U�Mȉ�F ���F �=t�F �E܋}؉E��}�u����t+�5L�F ���F ���  �$�F ���F +��F ������5L�F �E��%$�F ����$�F ��F ;��t����F ���F ��F �}ȋl�F �uċ�F �}��U�=t�F �������F �=��F ���%�F �= �F ��F �:�  ;��F �B����]ԉ}ȋ=��F �W ��E����F �=��F    � ������F �]ċEԋ]ȉh�F � �F �uԋ؋����F ��F ���F ���F �Mȋ�F �E���]���  �5��F �E܋}ȋuԋ=��F �   ���D���%��  +E�9��w��������D$����F �5��F �-��F �=�F � �F �L$܋D$؋T$ԋ|$Ћl$ȋ\$ĉ��F �L�F �h�F �=��F �-��F ���F �%��F ���F ���F �-��F �5��F �=��F ��Ëŋ��F ���E��  S�U��L�F �u�P���F � �D �54�F �]ċMȋ}��Ћ5��F �E���  �v������F     �u���F �H�F ���F �5��F ���F �]����F �0�F ���F ��F Z�=d�F �]��x�F �M�u�m� �F �|$��x�F �������F �UЋU܋�  މ}̍=,�F ���  �5 �F Ǉ�      �]ȋu��5l�F �7���R��F ���  W�=l�F �;��F �F8����GI���<����W�}ԋU؉��F Y�l�F ���F ��믋ы��F �uԋ=��F �u܉=p�F �5L�F �MĉE��E��   ��F �Z�- �F �j��F �L$ԋ��  �J�|�F �J���F �Z�D$��ً��F �D$ԋ��  �L$���q����=p�F �=,�F �U��]��E�    �H�F ���F �U�ǃ�      ��  �J<ыQ|�Yx�  ���#����=,�F �K�{�E܋C�E؋C �\�F �uԋu܋�  ЋS$�  �s�W������F ���  �]W���F ��F ���  P�E�9��~B����(�5l�F ���F Q�V���X�|$��t�F �d�F �5t�F ��$  �D$0�=�F ���F ��$   �-�F �D$��l�F ���F ���P��,������Mȋ�A���F �Mċ�+M�A�ыM��ʉ5��F �u��}��=��F �E��8�F ���F ����F �����MЍ,�F ���F ��d!  ǁ�       �E̋U����F ǂ�      �M���F ���   �]ȋ�F �Y� �F �Q�5@�F �uԋ��  �A�|�F �Y���F �Q�5,�F �r����'����5@�F �P�F �h�F �=��F �\$��L$̋D$ȋ|$Ћ|�F ���F ���F �l$����F �-��F ���F �l$̉T$ȋT$���F ���   �7�����=|�F ��  =d�F 9��Z9����P�ǉt�F Q�5@�F �L�F �-��F �|�F �0�F ��$  �-\�F ��$  ���F �\$<�L�F ������D$ċ��=����t$��-8�F �8�F �h�F �=��F �5$�F �-d�F ��$�  ���F ��$�  ���F �h�F ���-x�F ��$�  ���F ���H���V  �}Љủ]ȉx�F �}��5L�F �L�F �E�=��F �U܉U��ы}ԋEЋu�}܉p�F �uċm؉l$�5L�F �L$��1������  �u�5��F 9���I�����  �0�F �=��F ���  �8�F �Ή��F �=��F ���  ���  �=4�F ���F ���  ���  ��$  ��$  ��$�  �������  �,�F ��I�R���  �l�F �,�F �(�F ���  ���@������#  ������@%  �$�F ^�(�F ���  �=$�F ���  ���  �R  �������  ���F �x�F � ;��F �[B�����x�F J����G���ȋ��F �������F ��������  ���  ���  ���  ���  ����   ���F ǅ�      � �F �5��F h�  �5|�F Sj �   ����$  [�,�F �5��F ���F ǅ\���    ���F �T�F �P�F �,�F ��\������  ��`����� �Y�<�F ^��F ���  ���  �$�F ��F 9�$�  ��G�����=��F ���  ���  ���F �=x�F R������0����5�F �   É��  ���  ��5��F ������Q���F �M؉u܋u��;��F � p�����F �u܋M��E��M�Z���Xp�����F ���F �MԋM�벉�\  X��d  ��[��Ћ�\  �BH������5��F ��d  ��   �0�F ��  ���  ��d  �A��X  �@�F �8�F ��F ����  ��F R���  ��D  ��d  ������   �֧��X�������=�F ��d  @���F     �A�`�F �u܋M؋u�5H�F 95`�F �xo���uԋu܋`�F ���F �]Љ��F ������F V�������5��F ��������F V��������d  ���F Z�H�G����h�F W���F P�h�F ���F X��뢉�d  ��   P��F �,�F ��D  j��F ��   P��F �,�F h/ jB��`  ��   P��F �5,�F �5��F jB��X  �L�F P���  ���F ��F �@�F :��$��  ��\  ��d  h�	  �7   �=   �*���V���  @��F j ������Y���F ��F �� �������l  ;5��F j
�5�F j �5��F W��  Á=8�F Y  �  �,�F ��F �5��F �5�F ����É �F ���F ǅp���    ����p  ��X  ��h  �5@�F ��$�  �������I��$�  ��$�  ���9��������$�  �쉽�  ���  ���  ���F ���  ���  ��8�F     jP�5��F V�-���Ã����  ���  ���  �;��F ��������  ��$�  ��$�  ���  ���  ���x������  ���  ��롃��%T�F ����5T�F ;�$�  ������5�F ��$�  ���F ���  ���  ���V  �,�F ���F 3��  h.  j ��l  ���  ��   h�c  j��h  �L�F P��F �,�F �5��F jB�<�F ��   P��F �5,�F R�5�F �  ��������.���h  �5@�F ��$�  � �F ���F ��������,�F �5��F ����É��  ��F �5�F ���  ���  ���  � ������������  ���  �T�F +��F T�F ��$�  ���  ���  ���  ��F ���  ��놉=t�F �=,�F ���  ��ǅ�      ���  ���  ���  ;=t�F �������$�  �$�  �5�F �5�F ���F ���  �T�F     �����0�F �E� �F 9������E̋0�F �Mȋ��F �EĉE�Eĉ��F �|�F �]��;��F �����E��0�F C�M�M��M���������F �]��M��E�U���   �5p�F j��d  �L�F P���  h/ jB��`  �L�F P��F ��X  jB���F ��   P���  ���  ���  ���  ��X  �-��F ���F ��$�  ��`  ��$�  ���  ��  ��$�  ��F ���  ��$�  ��F ��  :��$�@�F �@�F ��$�  ��$�  ��  ���F ���p� �|�F �Ű��F �]��]ȋ|�F �����5,�F ǅ|      ǅ\      ǅ@      ��8  ��h  ��@  �3�$�  �v��F ��4  ��h  �3�$�  ��0  ���F �E    �   �����F    �Ή�,  �,�F ����)�$l  ���F 1�)�$l  ����1�)�$l  ��0  +8�F ����)֋�F 1�)֋���1�)��;��   �5��F ���F ��|  ��  ��@  ��\  ��8  ��,  ����+�$�  +��F ���F �p�F ���F ����   �މ��F �p�F ��0  ���F �.�����������,�F ��T
  j@��D  ��$  ���  �,�F ��$|  j@�5��F ���  ���F �,�F ���  ��B��h�  �5��F S�~   É�(  �,�F ���  ��h  ��@  �4:�:�R��$  �p�F �:�:�R�� .  ������= �F ��8  ��   ���F ��  ��4  ��,  ��F ������F +��F ǅ�      �5�F VP�e   Í,�F j �5��F �5�F �������,�F ���  ��B����$  j@��d  ���  ��X  ���F j �5��F ��$  ������$X      R�54�F j<j�   ������t�F ���$l  ���F �5��F �5��F �1�L�F ���  �2B���  �4�F �5��F �L�F �t�F ��뇉��F ���  P���  � ����Y  P��x������F ���  ӄ$<  Y+��F �$8  ��$<  ���F ���F ���F ���[����fac�QEG-���מ0�y�B#Sz\<z.�w CW�����A���8�.��g8q��������g�\F���ޏ�r�r�����XJz|����(��� I�V�%��`:�x'����o�̄�0M��@�1�8ɛ2>�k�T4,�2v���"s��mH?���fAs�T1ڔ���ƅ��1�]J���I��^��of��YukĈ[B����i����|���6����W���HSk�bWD��
�� ���&Q��KG�G�8�l�%�����`�3��v`��Xj���3�b��\oI�n/cev��l30W�I{��eCx��,���������~5S2�c:��晆m�ޙ��DmC<�dԮTx�Z'�us϶�6B�R�Z��a��[�^�Rn��W�g�P٬�Q��OW5�ݥ��A��,o0��	:��^��"l�!U�.�BB��c��±��p	C,�A��  �s�e�RT�H��l���-�)��C(r2r�l_�z&��P�:�?�+��T��e^P�
����R�p� zI��� c���Xm����&n\��U��kli��[�?, �~b�;j<?Y��ó�������M��DD��3c�-%\��f�<2l�����\�#��lh������o���r@T�������A�t VbE���e�*���3<}KT�Ԉ��y殓������������a!GUV�}<�}�1����e�e�3m�F�mn������BEN���(�[y(h]�/SbZ�H`������DH&Τ^ߠ�����L���$o%�*G������!%R�����c��l.F�R�QU*+�ᦲ���1��K�U�a�ջ�^E�}�3[�����"G��۾�`�,5��@�,��Q�ڧ=�F��/l{RH2�&+E����@���t���g7H�c�{�!��ή̑���) �!�n1I����N6��Q�n�PҲ�6�WĆ,U��(I�sۦ],z�ߞd'���E�Į�W����-��!f������Tb�e蹮G���ٖ���E��nAK`�QN����ȵ�d�Υ�`=]��"���]��"���ЀBu��e3�Q��æ����[���/P�6���V��BJ,
��91ح �ϧ{��rK���~O�[��IizS���FBs��W����Ѓ�*��-$z�Qɭ^�m1;�1��<.f������r��'����*���O��M@la�6�*�����e�}�I��e�X�t��(2��J�$��VDӣ�c�"�j���f�����	U����PT�=�:�#�?��G��CCˋ��:�R�$o�6?*�����iR �5�[��\lϕ�V�\F��/a�Բ ��IfL"��������*6KpWDD�����~�p�yQQ�ҋ�,1&ŕ����JL�"�a��4�Bq��j7T�?��6}���	څ���J�,��Σ"����x���m��Vq�%PNO�Y���L��4����Z?T�����K����Y���ԒV1��D*nL��RM\-�ԟ�E���J��a�����=�Ӣ��Y�Җ������Ŭ�(�e�\ew��ٝw/�@B��ʄ�4��e[�ؖ�3��h�n/��������L�χ�w����A$�Tb	�hT��誓w߲$#S����)yP)g�r�xi%'v5�	�ag���4"��?�b��G���O�o����!Z�s�5�b�z��o/i�DV�/Q:�
�x��KR�]b�������1���;��T��#?"��9�aR �v0ىzr��A�9����K�<�K.ל-�7Ρ+�]�;���8,H�$ed_ѕQX�w>ט��{b	�$�r�T����Nl�ʴU��o��V��$M���!��K���#f}Kfϰxȱ3&��>A��i��G�g��[�@���k�m��Xjr���y���U+��y�"�&��D�1k�#��Q��l1jF�>�ԋ(����fD8��9��H�V,�u��k2[��Bˋ�NW�IݭD�3쇹�%����x�T��O='jB���H�7-�{�8eE����c�>D�P�`v���[�wտ���\�+̻=���3����=�\L8��R�WZXn�γ��&�M��u��&ꅞA��wL)8%� ЫCA'�.��Ir߄?xMd�fU�3a���w�6��\����s�ʟ�1����V�~���[rO�خ�.����G�/6w�#�y��[���=��N�z���}�<�QwU�Ė��'\3��p����k��	PB�87��/�����ttu���SR�����-;h��)b0��Ȑ=5���{'�=�/�Έsql�M�q��{K��?-r��.mH����#��(�Ȋ2vZ�S�L�B�?sp�OնW��̻�t��/Q��M�`�&�V�/	b{AX�y�<L�fs��1�R����|-Vf��iN��a��=��h��m�'�)����A�X-h?P�'��A�%�n���@T��������t �\�u����ќ�%X+�ȃf�W�o]V��k��B�p��s�O?5�҃��Ա�N�3��yaGG�����4��B�7����)r�B3v57�b4�t�9|$ 	��KI�`Hާ��qχ�L�Q�άWGy�c����d��\�L���66��a��j�$�����;�t%]�Q+`o�������zD_ԜO3��Y���k�nk�1��5�F4��&1�_�Q��O�
��@#�ED~�K�r)����-�,uͥ�(Y���o�Q�Px�[�uη �hy��$ >:^*ޒ[�W8}8��fqH�c̅3c^�U����@>�t��z��ղ�Y�=�Dђ�88c������:��u7V�):�y�I/���񉢅��l�#�k8];���/B(R��d�����Y`PL���v�%���
�۰�R��>�`X/���/h���W��n�������j�l��fNL�`tW���Y��/W�Dk]{��q��o$��ʩ�_�m��� 𷔯�6a����Z0%?L73}B�Ƣ��_LJ.,�T�h`�4��f��[
����JU�oI�8>����^߫�l��4!��ɟ��7������A� ?o��t���TI�4<>F�ZΚ�UP��ݔ�%���`��3�h�~R���4&	���}1�Ͷ�=n���Τ���M���!�)�~���pH@\N�J�#��aǑ'��PS+�x���Wb��c��n+6Ԩ2�4��ڵ�J?E��z^0�X�;��S��U�BMUB�o)Xo�n����W�a���5���L~A?2�:A�����ҥJ��ѷ��Ue����oՄ&��>C�4[�`V�ȊU3X�g�3�ׂ�~�j9j�
��X�.&���>J�!��5�$F�	�ᝌ�=X��q6J���#5l��;xK�R�X: -x�k����"����TL��!�!L����w���;�lf͔O�y}q
�5�-1<Qя�X�dvH��E����`�%C��NڭS�q=��edd4R�����$GЀ�,��jYuF��E���\��"�c�˱%z/�n��]�c�Y4�Yoƅ���}��\m`�Y$�jp�-���	�=-�Rn7>��a�HD��w���S�c\���zH�9�Jr��cbn�Ή�&Nos��?���Lz�t����?J!"ӵ���x�Y`���5c�c���&�UW|����U1T���ANOO+���~ab�L"v@g��)b���xT�o�\O^���b6Rl��zG���@h��"�i�ɕ�a���ZN����4F�����	T�������%�����d�~�?x�PtlK�΢��Z<�ԝ��F�TJ�٤�$�خ���\���$�v�}6�wi����4� $��������!��b�����Զο��d�,���.�P��WSZl3j`���A��V��/z��Dʜ>��)���F��[W����bS���ˮ�Q� x�ܲ�M��vaW7�v�@h�;���x�b|�-f+o!ҵB�ް�������dmMu� �l�2^��kr���րI�"�j�4�����	�X�#?;Ka<��,�P�{��
6hJ>�M�(�G�v6�V��Tr�1n��L|:(:�����Fi�R�p��y��1֗!]�Lxq�	�5���w�"n�5���*�Bg�q`gC.�It���B_����iK@8���w-ԃ���n>�����t�|�s4�������;%�6�*$N7MB�h%����MV��uO�$5�F�w`#��	Y�Eb���Dfj<�cz����H��V�L󢎛�8�wa��A�5,���H>�o��RV=�ہ��f�@�偧[(�C���Q�����̭O���0ъp?����?����E2٭�턱�,��m�6�ő��44�s��#>+�?�󽨴��zJOs�Q�H��XNlDdn�5���o�a;PK~�����D?]�&�,�ee�Ł᧻Vb�s�o��J!VR�q�P��6��� 2N�Tio�,W�؆�!�:L��p�뙝�dʩ�}�R�ㅘ �������J^|">���H���`���
G�h�Cl���*�jtu��hI1̗������V��ұ�>CK����v��`���VgA5��'����3�[|�1��R �Ƭψ �Yݏ;��;�"�UT��|^��(B��d��������{�3L�/n�s��I�j�g����F�L �1]d���`�I?��Ԙ?J�����7c���ɸ�?N���5`F:��m�=*�>�Oj:IЩ�b�iP&�#0����1�p��B K 2��U$x�"1���ZA��|k2�o�B4�j�p�`�䚽���M���d�i(��-�G��:��g)�"m(<��uC�GBr�IW�&�h�{y� hr�la���+0l���z�9H����^�YǸK�ɜ5~�a�4�$�W�r�m�UQx����1ş_��8�����\�����PvZ�c`ܺڬ֝�(j�g�Y�*�o$@�	�Vhܭ�����!���Ui�f��W��C��\AW���쐃 2+~�kl�FH����Uc�4L����20z��$P�M�O���8��ќ�j�J�L2�.��yr-T���l�n���;�镇Zӳֶ��8ڳ��}��g���|��#	���Byof���dw8j��AЯTq=;������QK���ؐ^��>����_�4|��\[#~���i�*h�mgH�K�;�9�E�6NXL��إ�tX��,��|'X\z���� �#�\��'h�İ�Ψ
3�c��ɕ��k�֧��kt@�:���2j��"�/�Ps̤��s�rȹG�ˉ����n��,�s����12E�[�V/GR؀��{o�1M�P��&�����������@D���6A�c���M�7#������} ؄bDt�'Vkz�p�R�������]��S�W�✌�� �a���gGN��	I9?����<!� S�t�mq6󤣀�goDm����͓���:��N�Ń�����ڵ�a ��!s�N��.mn̡�'�t Y]�۱�Ru,K��F�&㎯��X�eǾ|$¼�����ի�O9nˍcZXߓ��C�$|�֨*�Qo�1���ۦA�ӢaJZW(=�"|'@$�Ym~)���^��cfpc�d� (��b���!��X}�����;���n�U&���:�B��NZ;�V�y����Ul7`Y%��h�C~�"G
�,Ep�#�&�h9��Mz>��ܩ�L.r���7���3��֢�r��e����\�����f��e��S5Rxx%�B�b _t�C��Cmڈ�<�Tٰ�+j"v
Q��u�I�pO��:�_>�����zR��c\�㬼Ǻ�F���َ
t��$ø�dn^Ю}�w*G�"�O�Ò92o\�	�$�,�����]<��-���A2��;�{�=�sJ���3�����KɭB�c��$�i�t1��7S���n�l�h	eUƈ�1�am�K����p;�a^����^N�&�u)�R*�rIc��{�(�¢J��J����F^�7s��|���'KY�#���O��=P`
f��C��,y�6�O�6nOn�w��dG����G�i����|{�)��p����}n`E�wIw�O.��$&fo|y�l+1O���6�1좂&�\X�T0�30�}�h���\�r�	5K7�JQ����A�1nU�(7�h����!����P�_����i|s8Ֆ��0fa�����HvYy�iz�x_a݌T3����(�*/8v�����	 ���[ct��{��=S� 4ߚ�CD�澦t ���^�O|S�p�-�S�
����qQ߽��Z]Z�?󒮙d�i7�F�F����q�ű���sܙ����.-�<��/�sV�c����Z��q�=�_��xJ���H��c�ˣD�a?0���:���m�*�W�"��+���r~L߄7mƇ>_����N:c�`�.�밴��+�TS0�^�B���\�i}<��� l�t�Nsd��j�G.��):�?@/�_1�(��wZ�&ʹPH�D
yg]la���&o��In8���'T9���A�.2'��V>��ۡQ4GL��s����,���k۝h��;hS"���:����
���t:�)<ٔ�3��u.�\�hO��	�@�����s�](f���\N�5`�����ﵣ����r��FUW��bm�G���vbH��'��7@�T�<9�K���Ys�����R��yKP�C��/�b��ą�ѭ���&�T �Yw��u�s�=�EhGx��C2�[O���|89�{	 �Yԣ���<ol0��it��1�۽��7r� ���H��o�,5�b��F��D�${r�����%0�5���>(����&*�л��r<;�>�O3��%��;_e���H�P7la)��'i���i J��B�� �ދ�;x����g#KW9�'��x�~u.���!P�}��G���m@��R+��SG��8�&������T��z���N?gba�C)����i"��aZ��~s�s9	��è7�W�2�"�l㡹���⮫�
�xsT���x"�8�3��V}�p�u�}�;���蹊��K H���eU&��C"��Q�XӮ��t�g���T;c����l�b�ꯞP(���U����a���5��m�����A�q�`g/����/()m�Ʀ���?1u��2��["��ǃ�Ye�.�g|�s����������
~����^�7:\��o�����N�S�{;���sGH}�pi�[ڠq�@����V/�ē�j��4����(�g�{�e���O��qۨ�y�BW����)����*�3������'tK�z�K�S6��"�$��#��)�B���p�����o���*��݆��/��C��.3p�޵O�}�HԮP�*���J���(|9:r�GT�����@2E+������x-��e*��Hh��É�d��p	�\���  �ɺ�S��_��έ>,㮭���cΞ��+��-&_n�m�"�Z*�f����;"K3daP�f9�����������H�~�7�E���B;��Fҧړ;}/�ɫ�CX|�vq]e���J.�L(�BW�}�JS3�O}�8���D���,g1�l`OM#b6�؎����4��Ene;�r���3�|x��L�����$��p�NZ��V�n�sL���e�g��U�N�/1�3��!��� W�=w�N������̣o�_���@�3����#}��MZg;��GGT�>���nzwᆗ�h�S�ߤ�C%� K���Z�c�o=P�>��Y�s9yÔ^H�m3�zh�3�Y��FS�9�<�TS)�f4>vz+#�j�D=2�8��u�T(���f��B���*�������q�o�6�m���Ɇ]:վ�+���CºX��k>���X4��%<PE�*M�*uՕӼ�+f�j�Jq�m�ؤ�zpS��s�\m�l�8�5�M�7T��r�~�hR�H�>k<�R%�2�;w'����N�J�P��[㐌^w��g4��)�^�}�6׳�H�+���W�\pL�yl�ɖ@!z6�54=�B
BX[��2�2�H���j��ڻX���5Or��]�ph6���T]�<���p����t�;��`����[\<H��=�[S�֬�鹸q_�Y�@R:�4ϰ0���s�\�Ȩ�{����+:sq��vD���U��ӄ��ߦ�u���ͻQ3�����&��Ok����k9�}��|z�y�V�;�?���E�VG�El2��?���d ),T3,;Πh�{�Q�3��AqF�$a�r��$@)�i6i
G'�s${�/4�n��w��d<���ձC��
��w]��e�t��T�9�} kŒ%�S�ܢ�� y4O�*}�ǂ��-����u�V1w�d���{R���v��1ka(z�N,ek1����L��ܕ�2<���@~	��'�ē����X�A>Ők�3�}B�QP����(*+�4*z�1ҋ�8��x�a�1��%3��y�/���}a��0�A4�vG>gB7ׂB�W�?�b���%	ټ���&sv�:��%������iEXa���H&V&j��D���0&�a��.m�����Y�����w�p!��[
$c%PP�
�ݓY�|�4�^ɩ��؏N����{WD�]�9�r�Y�w�����[Vy�N����c�x܈�fZ��&�;Q�J.qJ,�h����v���@���ؕ�#�l�d5馃Ӭ޽*+�W�WL�����YQw�P�g�vgVnA0�F�j'�'u�uaB��=Hط˧�a����;�tW�6����s:(�"�wgJ���-�Q�W�ż!NC���o�����U��	�w���y��t��3Y{���F=�n���G� կ�C�C�����H��4p����KL�R8��#��9���J���a�d9y��q��d�4��F=�%���EĤټ	Wk�5t��4	�I_�s,f������G`ӕ����l
rWl�@*��z����zAd��p)�U�~�x4�֎1��/�������h�24�9b�;��5ߵR�����J�Ǳ�4�����6s�wi�K�uO�u6�(�4.���WOO� �aC0%o>_�k�R�K� (9�[��P�K��#B�=[ؽ)�u{A�\+��ד��<�mR�ۺ<��u�3�e8f���E�'XX9�X ��@�}γ�^T%��,��r�%���_��}�ʂ����[KR6n[Ih����Ё�����w���O�F��[�1�V�(J�j ��*�O��5��4��c%���c�UνB��ߟxW�9��N����pr�&Q�$E�x'����)`��˓��J{�s߰֩�w�=�� �b_��ƽ�#�� 1%[n�&j��f�P�m{���B�T����U���u�j|�KL�io���(Ly����,@<�܁��(��'[Q�5J|?�x�]��|�rkJP�,����kdi�>�a>����3�����ɾ��C�?rH�.����44I�B쵾�u��z7�O/JbOr�?����_����TI�he�2;����?���vk�-,V7F�V���@���_� ޏ���\M�U�ɽ�RT7M3�(t�5��� | x���ز(u���?�H��Rb�O榷�np�dia?F����M����m�H�у+'���ZO��p����a��j�Y��ڞ4�l�DFS��q�E5��ҹ���U�C$�5�bBg�m��li��˘���)�ؘ��Ge ����t�<��agx$0$���լ�ގb��-a�`�������C@ݬ�fAA}J�zF �\i�=��Z�m�?�����̀���KE��������6|��1�*�X�Lk\g��'Z�rp�b�*�E��/q?z?-.�׺�={�)){�(u��l)����v`��^Yˡ,�:��o����F��z��L��_R$P~�"��+BPRT�L���fe��Q�0��gfZ00��%���k��7`����Y���V^w�8}�x$�} h'/'��\�������Qh�>1q��MPW���3y�/BD꩑������`�_L������6�cR#���k �_f8�k5^�1 -*�ׄ���)
v����<�����ʍ��#;V��3$�UH�3=I�)L�W�xVQn�hX?d*��!/Ч����ǧ�[N@�E^����ŘM�)������:<ME���g�X�Y�܂��i�Y����a�-�h�O�3a͛��x��>+�aw�g]�Eoz���_��i#�ևG?Źe6����Z��.X�8'�}/�+�ʤ���F,(�����aj�9`�ܩdCQ�#�t�D��i� _�u�g��[�P�9y�9e� �s:�$£�`��Qo����^�&�&�L�QD���*d�?�k�"3&ޗ�B�ڑ��壆$9��k\I:=FJ�}� �O����FA�ve�Ww<4�}��<��q�����j)[�:֚�$a4%�g���b��z�Xzi��ğ�����0���أ�:`��7�QE�k�C���m&>��4c��p" ��}f�ǂ�%�V�pu8Ď��7�8d��I,$y%�>kv�5�\-^ؽ�_���f�Z��؉�6�h<�L�¢��c�@����&����F� ����^d�ΥD�ߐT���!�A�n��l2r�%I�3����kU�7�|
Ƀz��{��ț�yP���DU�s5�y_�+~+@�LKO �N�9�op����6j.��(O��M�ǭ��&����<�x�TUx%�pI�VN�� �B_�n_�ɉ2a�ܝ���j�=�����G`B��H��$y)�Ѿ����B&�bر#����su���ŨGw����;�uıg�"r����p�@�8g����!��hT\��L������A҈�k׆%(�r'�42��h��ێ�k�l��4JL?�9:�g�@��~�K�8��)zl ��>O&fh���Ň�L!
�n�����k4沠{K2[��y�8�XH_�ɯ�ejY0�Y��wr���� }o��dC�Tqx��)��������`��w�z!�\�o$U6�2�F��Rl�R�,�e���tEA��.*�f	j�i[��bZs��m���\_V�PQ���~�t�����I;�mZ��M�K��P֡�!�{�ƾ�f@���ǌ
h%�����7$�fͫam,&��[��ơ$���DT�����%�a�0e��Q�՘:>���O��i��϶5�����߰Ǚ��hn�L�<98�'���g?�w���U"S���<TY�V���vT输�NGqA���|F��л��右� �����9Xii�����L[>ui�n� $�?V�$�) �W��y�Ql<����-b�p9K�^6�x�-��Cl�О�.�d%�}�ԏ�i-r3���ϫ"t�����2�9���a�y�0m�k#��>�凪��̒��!����)ġ��CR�Ypi
H�g���Tfi��[c�o�����j�㍦Go=8ѩ���4lX�>���;o��>O� Kc�"˘��[�'�zoz�ε&j ~���t�v2��ܯ�΍1.�Ǥ3S͘JPN��&<�(�ɻ��`�ʙ��rO��_7�U���وe��A����x�)��+aq|�љK|?G�S⷗;�$�7���ka�?6�r��8����YL �ȭ%d��{�����&�r��<�����q��G��>�����B�Ɨ&#H�[ol񮝌;��H����Ȕ�:�;� k[^2��;��m�Z��dGu��ep�F�ץ,�SIx�ߎ4�b�NZ�l�y�� 7��c|?�Ǥ��g�'+�H e�u�ꔷ�B+ �(�x�,�7o|N�)�h���}�j�g2tA���
_�+��*�@�m_'�~X�*چ^����� ;�p-ڔ,��
����������<��c@���y�Y��� ����N�	��$�(�0<kv��s�r`��vdL11ψ�_y.�|�6�785�����N��מ+nw���/�hC& �(�q��P)n�t����+����u"�{k�{�^2����j�U_�����V��wxk7<�Z���ޢ��q�4�?�Rio�&[�7 ��{�%KF�_�!��) d|�� \ءx�ʃ��Ċl	XWD��R���u[!CI�P���m��ˍ4.1;Q^��Oڙ����$��~z����弇��h ���_UX+�B�6S�UJ������;=(^�F��;{�>vF�-$ްܭ&9��GΟ%�H�q���x�_����`���������ė`�lr��n�"榖���SD��
E�2p��S�O0bS�����JO�1.��������sA��MYءt�L�Tem9V����Ī\G����U�Cs����b�X+�V�`{��XGC�"�1�g�J���^F`.��{�������@�k�(��&V�80W�yO��QM�^�I�jv�m�}ҙ���[�6��	(����5:p{ϲV
�Bi��a����?'�ݓ�T�[G�����ɼ�'Xg��t��Ǝwӫ�^�=zD��s¹���~dr�"�?<Z��Ǹ��j��?���Hv˝˄����,S�����u��pB�����o�ٍ%�Y��Pwh��Os8Vy��ҩ'bE�i �4޹��ݧ���>��~%��R��]��{�&�O�b�zг^�/E�N$��ccY��ɽ�o(7i�t�E�Gk�c��#p�4�LB���eߋ������FO_E�ڤcW�c�hV\�9�<8���c�ZP8 }%<��Y.h,4��-m�q�w�í�l�Dd�{� +��0��7�sj�\���	�|��@�2d�VvT4GZ3*Q�82�u&�� �����T�I�#��ڻ'����6>,ʇ��ׯ���{,�/��i�]��W��{�X껆A�������0J�Sm]�;r��1Wŭ�Y��Ai�W��B���O+<HmXS��L��3�>^D���4�6B7�2	����Ą�ݭdv���'b��_md�Vx�+��?��\��2L�.�rP�H"��v�/���T�U����t�U�`vk#^^1~돝!s�Y���XQ��˓�y��i���qX�xL����$������� d��-�8�9	tm��WM1T*�9��!���x?!71NYH�]�A��ꢩQ<c���}�b�y��Iiw����bbM�iˮ�v��{���YM�����>?�h p�鹫n���#��))����!hSa�UʹCB��rA4n�פ�"1!��U�2��d�����`��H�{�\�x��VE�Ƞ:-��X��ۢ빓�K4���n&�ά�ǝi���E=�h\�E�TW�#6L2b��!|ᨢ�_�Q~��Y�;��ct�����h	�,I��c�����Beb�e��)�)�۪�����$a��_Z�XVg�a:�l�E�u��Yn��($�4�۬�����)�D[�^@����Pe���.�.P��"7ᆴ����\�V��R����Jڕx`�W;�T�}�����!�k�S�v �Hp�PC�N�ǌg�&�{�� y:����$���EM͓Ň%5;]�ΟVu�,ʳ�f�����#_wt9սr[,jd[�I���1[�m�x]����m~�`����g�V�#/!�?��&�T�+�|�`J���� E�l��ǻ�>KI�M��$Ԙ��r����iq 쫗6�t`��t��mid��\6��M};����/t���h�v��
���a���J��������J�9��?(�~T�? �UO��al�++��y���g�h}	F�}�����z�4o93��YM��u!|��/�k��D���9������D;&�i��G�H�~��~$�T<�ԑ �ʎ�6,�q/#(M��cLߴ��r^���_pv�cy��\A��iPr��R;��0�%�{@��e�����P�˩�d9rAS��07Y��#���7?'�g�:��3�y$��YN&��v�#�����Ϻ�����~1@}�a�Qt�N�ͭ��p���=�yߣ�E�a�૰�b'��mT�}�8B����Yهz�4�s�!��Й�� �r\��i����:h1��1K�J�~Ԉ"�.HJ���q6�����mR���A�x�N���C���2�/*HT�@l�E�a%p硗<F���u��\�@Gtb(��H����W��&'��+%�08K�2&�"#�C�R������D�}�[PD��fy��mi��L9��"셼�N$����""g��*���%fT'�n�6�|��%��rn$��}7�k96�1P�<�Z���se�rG���&E���>�e�L���^ִ�]Y���|�S���8pP �b���ә�F�Y�#�zJ�7'1�+a\To��.8ǃDvQw�3�P�͓���T²]@�$�#���䎿U��?*������`p�m��h��+�1I��`o_��`�<{̅582�,�*���E;\�����]�&��^���iW�1˱@$�K�YT��r�|���2�"i��_o�k~�96��Rp�f.:us�77֡�r���P�q�q�I��k��!Tp�	'��.��fphR=J�{�ce/��ͣ����TB�_�Ԩo8CR�wI�[�[��'�o!�[�����h��~&���뀋�X4��K>6+�1���4�#�y��&��?�Ѥ�@01���L��j���{�-��9��V��	Ds>���U&o�{H��8&>�4&�K=�8ѽ��ȢA�� @�����,��^o+%OW��WΚ�_?C�s�)��EYz9lIP?{/��!�A��|Բּ��뎹�.SHZK�U���(n�U��K$} �՘�;����0�㿯�bD�1��sF=fx��Q���D�5>����.��<P}J�N��&"�H�#D�X�\���yp)[f�L�t�0jK�A����7�U��ʥVD�N��mdE��x��[�!FK�)�J�c]V����� ��گ��j�"1�"GA�0I�D룭rϛ�R@�JA%�y[@��:Q���L��`VYj��-C���`�0��ۀV�"��f%v��
�5��FhP|�K;K{�yQ$E�70�շP(��.�� �ĵ�+!4����X�J*�M��?P�Ri����&�<�Cz�Ն�5y���d
�M
����Ml7��Ble�%�q͉�A%�������~V����ٵ�k��'�.��U��.)\&�k|�s����I�髠�'ӉC�A���+t:Ư�	.�"�g�-�k�.��I��o�)�����`��ډP��칢��|����A�̼��՘��߬�ǧ����톮��G]�����|!�#"�x���l�Dj�$_�e^��U�z�d�9�Cy=����d�3��{&�3y~~@�����+���׉:�L���6��Ձ���UG������|e����'sH!q�!L��:�sr�&��a��t�)�;E�#���ʵ;�Ԅ�Fu�C��*���X�B�E�]��ԟ������6_�HД�P�u�0 �Jڴ�����i�)=�j�;�=��<�ρ�~���m�����H`s:�x'���Zqv'�=xΞ��aS8��R��Y�@�'���Rx4�@�uvs\�;�bI��7�F��G-2�~RR�|a8" *����7Ti6�C=V����B�lęԧ�Zu�NGU_Br��y�k�0dg�S�~Vk`�!�8�;���?�v�*&V;*1�5YN�fD�
���R�"6-��� ��ה����׽��:g��E&W��]��C��DM���
!Z��`�Md���,/�y^1W��76�/E�T__�i����gܞ_#��nS�#�ôl�!�r1�mu�P#(��� !���!��,|b�1�����&���@��DF^�[����#��mNo�&�S�o��@(�yF�$ǆU���&�E��g�"�oG]��i�ږ��<դx�>�yt��}]~=&q�Eo5hY�sM�~�azx7�\1Y��ɪ1����.��Q������ �L�nh�V�7h���[%Ai�&-*��x����pA��HPu&(�>�"F7|�q �2�?C�b6g@za�����K�F��B ����_>�e���b��c[1�\n�"����?7<��H ȚCؗ�5k������N2�ƺ���Ԁ��6�B�W��������.�^��t������* ~�t����-+"0���uVBX	Z�p���?	�@)��,�H�"��Ĉ{��8aVZ?�|^N1`�����9-N���`�U�O��F��h���L�7���R�D���"A���K�ζ�"���=�_�R<Yt(������Mg�$"?<� >c�h����|�7@��˽�gㅔ�ND�R�6�>��� Wڲ ��P�b��0�$�B�ۙ�R����nS��痫��^rn��P�-���	G�Fܹk��%#+�;����`O��O���P�X�S��%��dd���G�yE=��)��:8A�<@JU5�M�m"�iO�������P�� b+.��<"�p��?ϑ�졠.)\���p���+_ �������N�S���"�B(�PͣHj��b��1]Į�];}5�U6�%o��~�VM<���Sk!6I|��B���˄Ǻ%�Y���<#�Vk��rכ� �gL����=\���Y���§��L�0��������ގ2����R�Eg����F��t4�}�Z��-�����i5]��b�-�-P5ٱE���8���q���T��Wu6�ՠ~���Ebyz�+�NeI`�I#�IǁTtj,܊�ZFm_���1I���9��P �X�.��8^:ԟ��D=�1�uQ���?���i�ܻ�J+�W#4��hS�N���=sf�W�Z+��l#Ĥ�Gs�3c8!�K�d��v&;�<���&$z54o9H��	|u�W��5� d�����E�r41����37g��TwǢĖԬ����~@���.�*h�2%X�l�~a�"q��0�k8�w?s�W�0H��s3����U�������U/���~C)�Q�nѱ<.� q� �q��!nz�A�_�V�eU���&O�[YqM/v!&Y*�bA����y&��QLS�ة�0���#��}K�Z$�����⺆��Q�����UL�����Dk��P���#^�@Y�b���S��WD���5��%U�Y��.}�ttS$������^���E?�K�-k4Գ8B��awhԖP�K�?�lx! ,�����#$/�<���-}Jw<Rߖ�7�8U�UК��[����ߏF��_�I�p��W�<$7y�'���u[O�K�3���h����Hm�,���M�e��]]0�����z��h���F�q�)�q��a����t/?���Ek��iv�E��S�5ΨȾ�x�`Õ�p����F�k��������.��MB�g$1�3�4�iKX9�Gm(����u�v�h&)~x�ޑ���ˡzP�+�J�y��9��S�xBh�vځ�yiJΓ���v ;!���\ݺ��`��ў�%;�..�a�vTe"'�v?>p6Ķ	��
�&�lKش�E@/��i�nch��~x���G���.���g�Яa�.�*V��ҔU��^�تc�fm�d�ZJnI��Cn��@?9���	'�/=Y�v� �b^����H>��2d	�"�r�	�\�=L��8��G�օ?�������M��9՚K�R̋r�5y�W�BQ� ��� ��T�4�DV�����K2)2��S⥆E3*.�g�_T��s��{��zƦ}TQ��c���[2+��+ᔌ�X`x��W8�B�9� �}@��/N�Dzb%�1O]��X6�.v�WHk"�3�
�5�C���Aٸ�����к�r�Uw��u��5�`��
[�&�
��� GZ��Z�F����bXߧ�DjS�7�t 'o�7��_���T����[��4M�I����\��Y�C�������h��Z��Y��gUw��ɿv�F���;Wy��ADo�Y�T�n�l
�^'��қ�0�v�����-�[q6�lˠ��F���:�D�5��e7����x�b纒����ed�Բ~1`�`�6�;��+]��~omqcW+�>m�F��e�}���� QL|��M�hD���`����#mU�D���#��P���}ma[_D�������Mb�K�$g���5�,=�Ŵ�<�`���t��A4�:b���T�e�#�<��4cEv���`8��y��o�]K�(�S!�tO����+sRA8���Yx-�`wAr�ڕ�_������%>�v���-vl=t�qpCHCK��-�mA��h�qr�3���o����/x���y���VS-�QH�so�'��+����J����mn�!�Y�'�f���j�#
M����	��\H��G�B��I��[څ��[���u/������w�~�Ҳ�_
��z���~����]o�l���^�]�
B1J���no�+�Ҕ~Y�"���;]��9�ћ]�%�"T������rn@�|�e%tIɾ�6sf��-E��ԯ�齶�RM�
��ڞ6F�Z�Sc�����������FU��ǟ��}b���3|�kSPA���qW��S0�B�܅W^lrK����)�6�˂/M��2��S�\�T^�Q[���Q�g��3���[�k�#��S�)����򀖷��A�!�������p!����Us�'�Y��O�ɺ�tM^��Z���&�X&~��J�o�GW��w↷o}���6��W����"����0_�4�w��k����4�}�1��NԨ��\���QHXu]��3��F�ߗ��1R�Q"���v���$�[ti�i%߬�/Z�.O�*Ɵ���?����xu�pK�n�RgH���r���QW�#�Bb��oa���zx)�"�TX�!�?�`[,`QR����J��]�8qZ�+x �rcqQ��I�ʺӹw0l.�ࡆ} )�	Э�_�:<�n��Gv���5ߒ���ur7%�����3��QI�D�*^"��!�+N@TiC��o�u�/.3�;dv�c�d~E�hY7���5�wjg+���GR�W�b�&4�؜6���F6�p�P�ƀ���p�V����z���ϓ�S�=c�h`�8r����4���-}��۴d�����?_Ŀ�H��ȷ��X�{7�����}~�-�bx�J���B����DH�ؓ�����H���8�L��\Jzs��Ҩ��7��y�'�QRQ���W�V��/��򗥢��ܳ��U{>��0P' ��)e�>���D�C�s��ٱ���.{ǂ�.cYܪx�� ��SW��^P,�H�?�;��*-q�#�N�6n��S���1�H�3��ϼd;�-fEa���3�@�ic��Ƌ-UA]i��{=g��AVw!^�h5�m������͍�M&�z�;���?)�T{,�F��U�:C9
��L�bH�D�i���n���f��R�Ű�a�ީۗ]�������X�M����
V�]�qMIb��M�II� ڛMʽ6��+G��u�~H�+��S1���L�<n���}��PD0��5�>n.pv�*q�K]4��Ѹ%Y���P2S�"*&�U�M)o�A�I>t	��p(<����&��)m����-�U޷�����ŗ�����=l�z5���k��դulj�Ri�r�gl���m�k�H�]�����6��K�q�LR\F�u�����h,�t�v��]H�� *��F�A-H_�9�y�y�Ű\�e�ls�?o�~bzw��}h2�T�dz���b�WL�$U���hi�mP���TB����j_Hq�x �<5�_Z��p=�}Xw����.�Q�Ǜ��x�Ğ�V!B**#�Π�M�M�tt�]�e`|����{�rqq,��6piQ�)��!B�߸�,R�(&X�����@�����jЍAY����E�#E�CcS���}L�f���L����5��eI�E5���%e���I6ɋ~�`Q��R.]�Qfb2!+���ꝡsC
�`dq��%����1�>d�G���'a��E*�]TS��u-X��˰�e���u���}J$"�RH�æ8b�C=rr6�S ��3P��H�i�ͮ�Y�pWhI(}��K�SP�FU�5o6�I�ݐ83і����$��}�~X%��S�y�c �_�?�J��A��}��H��F�T������𣾃�x�h-P���fO���J�y�4�yf� :���;$�:�1�����h��C�"
�L�i5y�����X
So���k�z�D~��rF���ׇT>�7���H�T5��U�U�0x�p~�9c��E�e�qϳ�6S�
Yw@R��_�١��/L=Al� 6��4Ͱd�K��KH������4Z��x���W�� �u^�IHC�#"�<lW�n��u�~ϸ�	��UڂF"i�&M`���m�<�`��L[yR����B?v^]���|�=�@�?:�0�t��kZ�a%����k��ҽ���e�����(�ɡ:�����de���(��wP%iN�u۔?fW�cճj52E��g��N����k�L�:q�rv�Ч��<�g�8y�Д,ǹ������g�s�Ȅ�M!Ш�����/tҥ�ky,G�IXs��;t:$�iɢ��+�H�J*�f�&�;XE>�d����	�uG�4�۞B'�e�@@��!�8r��،�q�O��d���-�׷�+����U�//�'IQ]��4 ���0~S�kBS&��o~��&��^V��8�4��ȸ*c��G0��C�y�7����y�r�V[��Gn#�;1��%�~�dF9�������Й��J���@�͋O�	I?>�	�k3Y�A~Vj�י�#r]�o����ή�Ѻ�gc���F���1��|�*IUWeܧ3�(<v^"�s³�Z��^����I���u��3���݈������2V�߮�A{���D3"�N1��3�J10y����>����p��@,�Հ���T�����JՉ�w��z�sRv�]��H�c�6�<�]Y��A�h[L�osP�����5{�@{u�(��^I�����Qfn��M�n!m�[�L��ڿ�����+��<���:D��}_F��Z�G�J�?kU\�.���ס��^R�ؒ�3�-Q�z�J�\?��`Ţ�|I��e�B�P�[F�ly�b`�m�i ��u�x�!�a����Du�F�������0��"�6��N�%X��ԍfk

^mY|�p[�]�u��ŖiNA�OB��_r=��+��R��n���G̈́��!k����c�_�K��\��
��C� �	!���%oĥ�[�B���p=��ݚ�A�� ���^5p%?�14o���� a筐��h< 뢀�_�A�.s��LN�p�����{��t�t�\ ��h�Z��s�nVfS��ʶ%{�� #�W��v<�rh��v}�}���p�S��~�@��dhV�j�<�������.�F��W4�����#�6G�W�h1ǉ ��h}i���-�\dVPm�"$�~���
�����W�����;��q��{T�Ț�<QEQO\�o�k�,�C֋L�1TD0��)bL��4y�]p�����<�o�[��nf�o�0R�
���#�nŽ��g|��2^���������<#y>�U��hf�����^�8��{[y�&������̼�q4o%\Z��%�?K��D˼jh}�}�}��ENup�E��T0�V��z;�2nϫ��b�����i�1<=u���H�c��ŭ�c�5���D+��N�`N�e��i=*[Аz(p��#��Գq��kz?cs�#�NRM�pF:�XT=�n��K�������p�$9�o�o��oqU����KT�w��W��rD ���+����'�ԈSN
�ؐ��I]�]�f�98�+�"��K4~ܞ�-LrG9�<�1�4�f �A�Hw���\��Z	-[n��@���E��2 �A=��Tğ7T��*�he;�T�VJ��@�}��1LT�i^�&�*�Y{�[!xS�J��5��N�"��vɀ����xpԕ�7G�_�a�ns�d�������\3��+���4��X�w��j��l�{��'�P��im��~��J�3�~�T)nF���0L�E�^;՛�L��H�!��Wci[���Q��䃡��v��T�9��k����'*!���5i�5�\�_���d3\� D(��q�=����C���9��@؁!�VO""Yh�V�6j�������P!����t�������\	�ڔ]�OwV��V��ƱS���+�Ih��5�   ���  �,�F ǁ�      �5��F �f   ��������F ���F ��F ���  ���  �$,  ���  ���F ���  ǅ�      �5$�F �5��F �5��F j�����9=��F �5��F �����P��x�����$<  ���Q���  ;�$�  ����������F ���  ���P���F �5�F 5�F 9�`����������R�l�F ��`������F ���F ��  ����  �5X�F �5��F �;��F �ޱ��FI���n����50�F ��  ��  �=0�F �=��F ��  ������
  �5�F ��  É�8  �=,�F ��4  ���F E9���������  ��,  ���F ��0  ���  �`�F ���F Q���F �;��F �����A�M S�] ��������T�F ���F [���F �;��F �����A�T�F �54�F �5T�F ���u����54�F �T�F ��벍,�F ��I������  �F��$�  �OO�����  �A  ��$�  ��$�  ��$�  ���F �p�F ��$  �8�F ��$  �5��F ��$�  ��$�  ��$�  �=�F ��$�   ��$�  �5|�F ���F ��$�  �D$��T$����ϋ�$�  ���F ���F ���F �=��F ��$�  ��$�  ��ŀ   ��|��������  ���  [�������  j� �F     Q� �F ��������  ���  Y��@�8  ����j �5��F S�X  Ë-��F ���F �-��F �΋�����'���  �F 9���������F ���  ���F Q���P�F P���F � ;��F ����������F I���ȭ�����  �E������$�  ��N�����  ���  _���F ���  ��F 9���������  ��F �=T�F ���F ���F ���  ���  �-��F �0�F �|$ ���F �5��F ��$�  ��$�  ��F �5��F �|$���F ����������   Ӈx  �=��F =��F ���  �,�F ���   �|�F ���䑾���  ���   ��x  3��   ���  �=��F =��F 5��F ���F ��F ���  �,�F ��F �(�F ���=�(�F +��F �,�F ��`  �%��F ���  �,�F ���  x�F �d�F D�K�� �F ���  ��F ���  ���F 3��  � �������,�F �5��F h�  �1  É��  �\�F �F 9�$  ������= �F ��$�F ���F �-��F ��$  �t�F ��$  ��$�  ��$�   ��$   �|�F ���F ��$  ��$  ���F �0�F �=\�F �5��F �5��F ��   Ép�F ���F �9������S���  ���F ���F ��  ���F �]�X��0  �8�F �-��F ��$�  ��$�  �-��F �L$���$�  �=8�F ����ǅ�     ǅ�      Q����Ë��  ��5��F �����Ë�I�S��������  ^�5,�F ���������������ǅ�     �L�F     �L�F ���  ��@�H�����$  �ŉ�$  �|�F �5��F ��$  ��$�   �=\�F ��Ŕ   �Č   �  ���F �Sm����h�!  ���  �@m�������  ��F �<�F ���$  ��$  ���ɉ��  ���F ���  �Ћ��  ���  ��F ���  �,�F ���  3��F ���F �,�F ���  ���  AX��@  3=��F ��F ϋ,�F �%|�F ���  �=,�F �\�F �%��F �t�F ���  ��F ��P  ��;�5|�F Q�5P�F R�5��D ��������   �J$��8  ����ˁ��   f��׋d�F ȉ��F �,�F ���   �-��F ���  ��t  3��   ��T  +H�F �5�F �5,�F ��
���   �- �F ʁ��   .�{���  ���   +�F ��p  ���   ω��  ���F VX������F ��=��F ���  ���  ��F ��<  ���  FX���  �8�F ��$�  �T$���   ���%  �싈\&  Ө*  ���   ��F ���   ���F !�O�-@�F �#�a���'  a��u��5��F +�X(  �,�F ��s5�]싚 *  ��*  �5@�F sY��E苂*  �   �\�F �B8�J8rX�Z(��<���  S���  ���D �,�F �d�F QX���  �X�F A h�  ���  ���  �ej�����,�F h.  ���  �Lj�����,�F ���  �؋JTӄ$   �J\#l�F �R+��F �=��F �=,�F h@  ���  ���  ��i����h�  �g(�0�F ˍ,�F �JHJX3z�rP+r|zX��<"�+r$V�235H�F ���F YJX��˛TZX���  �������F ����$'  ӊ�'  ���F ��F ZX���F �M�5H�F �5��F ���   ���)  �E�A�Y���)  �A��4*  ���   �Y��&  �Q�}䋹�   ���F �]싷�%  �U��M䉇h)  ��t'  ��P&  ���&  ��L&  �E艇�%  �%T�F ���'  ����Ë�I��X�F ���  �5X�F W�=,�F �h���F_ǅ����   �<�F     �������5��F ���  �5<�F ���  �5��F �� ���������ih����h�!  �`�F �Vh�������  ��F �<�F ���$$  ���   ��҉�  ���  ���  ���5`�F ���   ɋ��  ��F �,�F ��d  ���F 3��   ��d  ��F ���  �,�F ��D  ��@  3��F ���  ��D  CXɉ��F �,�F �%|�F �\�F ӣ�  ���F � �=�F �=,�F ��5�F 9������Q��|  ���F ���  V�=��F �}��/;-��F �����GH���A�����W�=��F ���F [�\$���F ������V�5,�F ���F ���  �$D  9������Q�5��F ��X  ���F Q������	;��F �n~���,�F �����N���Q~����Y�ʍ,�F Ǆ$����   Ǆ$���    Ǆ$�����F ���  �#�����h   h�uF j ���D h�uF ��������$�  �uy�����4�F �l�D ��$�  ���D h,QF �Cd� �D h��F jj �0�D ��$�  ���D h�  j
h�  S��  É=�F �}��M  �=��F �=p�F =��F ��˛T5��F ���F �\�F �C8�K8���  �5��F 5��F ��$<  �S4���D �d�F ��F �S,L�F h�  �K���  �he����h.  ���  �Ue�����KTӄ$0  �S\#l�F ���  ���  �8�F +��  h@  ���F ���  �e�������  h�  ���F �c`���F ��$  �5t�F ��$�  ��$�  ��$  ��F �5��F ��$�  ��$  ��$  ���F ��$  ��$�  ���F �-��F �5�F ���F �= �F ��$�  ��$�  ���F ��$�  �5��F ���F ��$   ��$�  ���F �T�F ��$�  �5��F ��F ��$  �=��F ���F ��$�  �`�F ��$�  ��$   ���F �l$���$�  3�  @�F ���  �$�F ��  ��F ���  ��  ӄ$�  ���   ���F ���F �,  ���   ���  ��F ɉ��  ���  VX���  ���  ��  NX+��  �5��F h�����   ���  ���  ���F ���  ��$�  ���F ��$,  ��$  ���   �N`�P�F ��$�  �=T�F ��$,  ��������5��F �sxhdF h��G �C�y�����-t�F pG��sdh��G h�F ��x�����5x�F �s<�5��F ��$  h�sF h�qF �x�����-t�F �A��j-��$  �ot�����{p�=    �o����,�F �E�   �E���F �E���H���  �'y�����s΋SHSX3{�|�F +��F =��F ���<"�+K$�p�F �,�F 3H�F �50�F �������F ��F ��P  ��;���   Ӄx  ���  ���  ��  ���   �|�F �䑾�-��F ��x  3��F ���  �,�F ���F ��F ��F ���  HX���   ��F Ӏ�   ���=���   +��  ���F �%��F ���  x�F ��8  D�K�pX���  ���F 3��  ��$   �J$��8  ����Ɂ�$   f��׉��  �d�F ��7�։E��M��EЋMĉE��T�F �=��F �}Ћ5x�F �$�F �=��F �  ���   ���   Өt  ���   ��t  3��F ���F +H�F ���  �,�F ��
���   ���   ȁ��   .�{�L�F � �F +��   ���   ɉ��  ���F BX����뉍�  ��F ӌ$�  ���  ��F ���   �L�F ��F ���  ���  ZX���  �8�F 3�  �  ���  ���  ��$  �T�F �u��E�    ���F �5��F �U��F\    �Uԋ�  �A<ȋH|�Px�uԋ�  ��������}Ѝ=,�F �B�r�z�ŰR �Eȉ��F �]ԋ�  =��F �F�֋}Љd�F �M��}��Eċ$�F ���F �T�F ���F �]Ћ5x�F ���F �=d�F �X����}̋G$�  �_�uĉU��Uԋ�  �L�F �,�F ���F �m��D$�    ��x!  �l$��  ��$�  �P�F ���F �-0�F �h�F ��$  ��$�  ��$�  �y�����d�5    d�%    �-�F �,�F �����F 
�=T�F ϋ��  Ӌ�  =��F �5�F ��&���  ΋�F ��F �   ��H  ��<  �   ���   =��F ��F ���  ��  �ǋ�F ���F ���  X�F =��F ɉ��   ���  zX���  ���  ��F JX+��F ���   h�����  ���  ���  ���  �r4���  ���  �5��F ���F ���  ���  �-@�F ��  ��$$  ��$0  ���F ���F ��$�  ��$�  �%��F ���  ���F ʋ��  ���F ���F ��F �l�F 6���  ��@  3��  =��F SX���  �X�F Ӌ�  �(�F ���F �  �5��F �.����F KX���  �T�F �-��F ���F ��l  �,�F ���F ��F �5��F ����  �5��F �50�F 3��  sX���F �%��F ���  ���  �D  ���  ��ӡ��T  +��F �����F 3t�F ��t  ���  L�F ���  ���  ʉ�\  ���  Ή�x  ���  Ӌt  ���F �-<�F ���F �d�F ��t  ��F �`�F Ӌ�  ���  ��  ��F ���F ���  ���F �|�F Ӄ�  ��  �����  �=��F =D�F +=��F ��F #�  ��h  ���  �t  ��$�  ��$�  �T�F ��$�  ��$�  ��$�  �=d�F ��$  ��$�  ��$�  ��$�  ���F ��$�  �=��F ��$�  ��$�  �%��F ���F Ӈ�&  Vd�5    d�%    ��F ��l  ���&  _Xʉ�h  ���F 3 �F �5��F ��0)  +��)  ���F �Ɖ�d  ��h  ��F ��d  +=��F ���F �,�F 5��F ��`  ��p*  3@�F ���F �'�   ���H�������  +��F ;\$��wu����    ���F �T$̋L�F ��9���������  �m�D$��D$��|$�   �3|�����F �   ��T$��T$��   ��YC���%��  +��F ;D$��7p���؉50�F �t$��5L�F ���F �50�F �c����,�F ��<�F � �F ���  ӈ�  �5 �F 5��F d�    �d�    �,�F ���F ɉ�<  ���  �%��F ���F +��  ���  J4�PhX  �5<�F �  ���  �S�,�F ���F ���F �����  1��W�=��F =��F [��F �P�F �,�F ���F �%�F ���  �%��F ���  ���  +�  ���  ���  5�F ���  ���  +��  �5�F �K����@  ���  Ӌ�  +=��F ���  ���F +��  ��$�  �C���{X���  �>��5��F ��������T$��L�F � ���d�    �d�    �쉽t  �=,�F �d�F ��0&  �3�F ���(  �%��F �0�F ���GX���&  �	��p  �D�F �F �5L�F ��p  5��F Vj2�����+��F ���F ��F ��l  Ct�ω��F ���F +x�F �5��F �c�Ή��  ���F ӌ$�  ���  ˉ��  �,�F ���  KX��F �D�F ӄ$�  ���F �j�틋|  ӫ�	  ���  ���F ����F ��F ��l  �%��F ��  ���F +�8
  ��l  ��F �  ��F ���  3l�F �= �F �%l�F ���  ���F +p�F ��(  ��h  �\�F ��0  ȋ�<  KX��  �$�F ��  ��d  ��F ��  �,�F ���  ���  �Ë��F �-��F ���F ��F XX���  ��[����F ��F ��  �=,�F GX���F Ӈ�  ���  Ӈ�  ��  ���  +�X  ���  ω=��F �=,�F � �=,�F ���  ���F Ӈ�  ���  c��L�F ����F ��D  ���  ʉ��  ���F 3$�F ���  ��T���  s֡K���  ӯ
  �t�F Ӈ�  �=�F =��F ���  �5,�F VX��F Ӧ   ��t  ���F #�F �58�F /���X�F ӎ
  ��F �%��F ���  �,�F ��  ���  ���  +�F ���  ���  ��F ��   �t$��R����L�F ��$�  P��$�  � �D �t�F �L�F ��$�  ��$�  �5H�F �(�F �5l�F ��  �$������F d�F d�F �����  �T$��-<�F ���F �|$��L$��t$��\$��8�F ���F ���F �t$��\$ȉ5��F ���F �t$��\$��t$��4����ꄕ�+���  ���F \�F �zfg+��  FX�E��d�5    d�%    �<�F �   �=��F ���  �'   ��B���F �5l�F �T$��T$ԋ��  �t$���+\$�C�ËD$��L$��ˋ��|$��|$��8�F ���F ��L$���  Q�����5��F �58�F ��$�  ��$�  ����  ���F ��$�  ��$�  ��$�  ���F ��$�  ���F +��F ��F ��$�  ���F �5��F ��$�  ��$�  �{�����@  ��   �4��   �v��   ��c���5P�F j �5��F ^ǅ����   �5��F ���F ��F �$�F ��h  �H�F �P�F �@�F ���  �H�F ���F ��F ��h  �$�F R���F ��������%b�����F �5��F ���F �5P�F Z��h  �=��F �=��F �=��F �=��F �_���Ǆ$�      ��$�  �58�F �=��F ��$�  ;|$ ��Q����$�  �$�  ��$�  ����058�F ��$�  ���F     �0����L$�������D$���   �-0�F ��M���   ��|  ���   S���   �Y���   �Y���&  �5l�F �q�=��F ���   ��x  �y���  �yǀ�'      [�   �=��F �����Ѝv��   ��a���5�F � �F     ���F ��d  �5P�F � �F ǅD     ���F ��\  � �F ���F �����F ��@  �X�F ��D  � �F ���������F �X�F �����=��F ���������+  ���F ���*  �� (  �5��F ���F ���*  ���%  ���F ���É �F ��$�  �%��F �����$�  ���F ;��F �cM���-��F ����$�  ���  �-��F �(�F �=L�F ��$�  ��$�  �����$�F �������5��F ��[����F �$�F ��h  ���F ���F �������5��F �BH�v^��VP��h  �=��F �������=��F ������U�<�F 9�������d�F �Uċ��F �UȉMԉ=��F �Mȋ}؉��F �=��F �E��d�F � ;��F ������Mԋ=��F �(�F �]��d�F J�������EċE��2?.�d�DJ�6��*�:����l���5��[k:�0��Î���]&�D�9���l��X�m`�M5wW��4��#�SQ͘��
�B�n�x_�5Z5�+�&�@F
�;;�#DD��\�>^U�����[m��+������>MJ�H��
7�ÐFIvMV �P8����k��={䝀����*���-	��cmg�_��ԇ .)h�M���.sn�m�-J�m�WU.��|�|$�
Ѝ�Eϙ�뱫ߋ���X͛��^�y"~F�AN&���Pd�n�]Æ#4=�4�����<� ���vRp�Sb)(�Q >C�C�����D2��1Y^�"���)�EY{)@:����W��aBdAݬ6�D���5צa�|�t	��ɛN[bi�ޑ��P�������>b��rĥ� ��]*�?�����;�����ܶYjP:% ���\W���]�H&����ƾ�i8��V�V;��]�����>FcFv�UL�b�vP�;TpC�s��3렆>w �0��7�n �#�v���p�Ȳ��X��7^4�6�#ƣvh�p�w�� ��{�����He�h-�Y�vmH|Y���bFi�x�v=Պ3��|,gWJxW|8�\7&ά�BN�Yd�lRM�|������|��LL��шCW���X�bǅV��<w~��,��G0���A��:���,tE��x� A�#��Z�I�#_,Lta��2gԩ�M�^t�pR��䵱auc��G�Y�!V�9�E�P(֩��L�� f���h$�`����4�_K���\�� ���C���%fv�~�
��ߧ��K��~g:5a*�V�=��1��a���=�߃��iK�x��N=�z�l� 3����{~؃����&�1�4�@fD�pi2j�"v��j)������6 z��`T�UY�TE1i��UQ��wK����|�Q���U��֖5�A��h�钇���.�N�=1����ێyA憌�FfJ���Y����$)���,�������-��u��]��c�u$G5|f�[zo�LV�.B}=�5�XZ>��5���H��2��땚7;v���u@��=o@}Jˡ��x�y�7�rm�ş����edI�g8�tQ�F2W!��Ooy�֞F8�;�$�K�+���Vض�@��u��&ܧ����D�H]��U�������}��}�i�]�~��3|R7�9��h�{-�Ok�����H��~�O�C���ׅ�%s{M+�H��J��"R5n���=��!�'$�+h�Om��-� A�G�p}(��v�]|dq��;�|Y�ͼGz���Us�(���$�+7�g]��<�ȳ�B�)�P�qx�Y�$~�嫍��5����+*:���X1<��~4ԇ��\�9�Č��zk/Yz?O~z� �q��0�}���{��M��Y����#|f�c��ms���k�YYc�ߧ� ��޼(>�.d�tƠ�Ѩ�+���'8=�d�w�` �v8U��8�wk�t�Q�1�괟 jF gSSc!Hg-o��a���:!F���s���� %�N���>gh$��Q�7*&�i�v:�ߋ�G��J �XYsc���<�g���PXD!����iI�+���H�DC�g�m�������M�M{������_��'ƋLq��L��X
?[y��C1���󒰜YR�D�o~�C�<�ًl#��5�-1�)21AI�.7t� 2��&��@���Ҵ�����^|�q򹥫jHa�>v���"#T^������6K�|����1IUF�%V��Rϼ�*W%*�����0��ѧ&`8�5�d�Z���sbi�UJ�gl�Z�s�7�R�6w��ؿ_@�c�}D��&��le��`MB!ὤ��g�r�:�q��(h���ȱ'��Oό�I�s����H^�I@%�x��%Dz����Q�rA�Q:*���#��[�4v>ԇ}?����S��tr�efm(�3l�B����]�k��I��<�`�lÊ�y>Ō��N���lRy3��^�T�H;x?P%�;�����1�*��B)G�N�5��ܞ�f�?�.~�|+o8=D��K'�
���yo�IE=A�DҖ(�[�B��՛��9ju`��Y��J�6��=0��s���y�(s;�_���M3do ����;�#2�Ҋ�]3pyы�]Q7le����m,��gc��o��ůŤ~�����7٩0�L,+YSj[3�Qx�Tz#��9%�ŖY}�Y�����~���=���1G �&�ـ����/��k��c�yW:���[,M�����͉�QCx��B,�}���jyg�߃)�A���h ц���s"'!M{�8�h�3���{X��g���Xi�������ہu�mѻxe�m���C�j-@��YW��@xM���y��@��	��p�?����く�Z6�Y�#���E�)�m�-���%���U�{O��%���K2H�4Z_p��z0B�4�2Y%���0��S��2A��	� ����W=��!��`�z�	��B����O�6K��"�:�?�!4"��~=n4�E�[��U2F�4I'e�+n�v��4�T�p�c����\�ç�c�Mr����Rɡ�D<�%xu��߰i������u?MNԈ-	"BŹ��!ן���·���>���r��W��V�7��N�le&��!a�Mr��:��B�.eu�*��z9ώ��D�&8S& խ;��"��I�!ܭ.7}�beA<<��=�S{-s� I|^�!�g�*�,���hM�"0�TD����H�D���L4Ƨ�}�񃐼�FO�.���G���C9
����7_j�����U~Czh8�خ~���������.���p3��U�
���2��g�5̉�w+9�A6���H�iT���mZMt6�O�T�����Ԭ]W�����9V)(w����⻫qn&z6�4+�GaƧ���F2�?����o�*�gp��'n�`��8��"��Aծ^���'�!a�0���#���D�6�5�=��^O��tHLf0�[�~f��%�'����/l��T��<���f��"�\�u:з��:֌��7�@W�`�@0Gw���AH�l�p��k�8��g�=BV�}��i��$a��ԝ�h��z��"0� ��Ok�����j��${/�ATo�c�l&�T�̶/�t{�ȡ3k���R�h|�~��-�b�)�f����!+v�净� ���	La�8�XRM`���=O��Z�UA�Q[��L��GO�e"�~�������F0�y0��^�w�|�"jQ�J]��
p���hXW�~�nh��b���?@�� m"�'��u���'��\�_S@�-��2_ꑒ������DZEIZ$�~{�M�х��7����Z�s@��%�:d�,����E�޳Ϳ�]L���H)d-p% �i灡�
��P�	�k���"�iD&�M֏,�4~%�nDUXr�Z���M�<��h;����c��ު洂(psG�+r��a����7���+�m�ͩNQX�AY
aĕ*����ne�|�lh��e����x-��L�T�L��'��Q&�T�gi���2�*N�������m�Z�/���{��0���-�"����./��Tus��pY	������gu�M�R L�e�r�1��Qk��=�z���JQ���h�a6���AӾK����[�D3�V�/�Է��,�v���_���|[""BF:MBTaU
���w��h�5�fa��l���I�/���(��7�S u���(�,��Yb�z]�"��D�ݚN�8�/"U0�q�l�{�{��|$"��r��#I��8�Fqb"6"c<1e���2�v\ZxNW����Oʾ%ӌL�)v֩bT��o��m;=^�
CuN�p�(�Zl�%�����M��lL�o�a�H����砶�k]8@&�,zp)ٹm+$���q����K�oW$E�y�[ �	�5�ֆ�G��<E��}$X�ilu��,�e�M�O�S��/+�T����u��'�d�>���"�f�,��J}m-րP�l���V��S��J�_�	n�sFM;����\ !���N�ME(s���ˇ�g���]qsX&SF^o�}�5��W�3���f�r!2WN0����~��Eo����Q���!���}$2�/]f�/��&�[0�sh�$��K�4����:�֘	��ꌱX��2o�{,3,  ��)����i���v�	.U5�M��������Jm�b}(��%ÝyfVN[> ��#���D�
�C�s��\��<	�iY"zV�n�
�E��(�#*��zJ͆���J�ч��^�*��^<+�(�0C�w�S�dï}��:�%z[�*) U�\o�]G��y�S�C]K~,ĳĕ���םN2!7$/nK2]��٩�D�=�w�}�CziwОahq�4�Ĩm4���G��M����"��*<O7��&U0���N���|Ֆ�
�۪hr��Ŷ;\�D6�qIE�Ḭ�%��Oh�"��(c��"S��X�([.;R-���?����8�yF��Q��Q�?ϧ��襊�\+�=�{��b�-�%����[%(Lu����X��:�w��*���ͥ!�ʼ�Yж�'Ei��o�|� ���%p��L�0�$���f�i�\�u���d|�0�|��F�t���"K"�jD	":�]��0�&l� �1F����]�}cۭ��ϻ��\l4�bo�e)�Q��W/��
�x��'�!����B�Yi�4�/��!I����E�i��goN\��KK���P%�rF�J]�b�^v�U���/�OV�n�c�,Y'��oʯ��1[ћVa�ks���I��֭i�0(��>�g��Ǭ �6�[�fOW��>��C�lhZ|6	���	��4�ώǬ��ȸQK{p�x���(��4���Æ>Pd�	1ژ� rW�gO�u�=�^>ԃ\B�L�#@���i��CD&H���p2R� 2[�?��׉'T-�jSV�p"Φ7�[�+�$r@��ɝ���S�}�PҬSO�n������|�o��eyO�s�h��1Y�j�mt ���A�V�r�9#���6�����#�j�'cot҄���c����L�&�n�5m}�)�{o�)�~�֣�4u�^*n���Nq�'�t�WZ��q��]ő��%�M�ޛ ����q��频��P7�:/FMA<@��Ҫ-2�o$�'�֒���_h������y���g�����fa��g�>�^���ɓ|G>�s����"/鳐TNx}k��ԑ#I��b&xLM�AW�2#<9�W�>�(7yhH@��hA2�1��qg�@&��rd;�w�;�9])��F�v4��tE
���{��g�p��HOc��&)2e�d����,>4y�F��R��*���%�߲�o ��rm�<7?a���,LX����q���`��H,�|�D:���c\t����5��@=rtkh�.�w�A1щ$.Au)�]��ba͞��a�Q�p=VG����8�e����վD�k�bw��C�d!1񵽻v'˷�g���b�
Nh+��=����;�Y8M���7BKcV�EL2�h����ㅏ�P��Y����kl	z	�|�@���)4h V;����QZW �� m�f����������~�|��!�e謹i���f�Q�mْ_ř{���4���6�|=`�޽�@B��G/<s�[�ӹ��V��2���Y@b����Z� e�B$�C�T�Gw4m�oDx" u�4ƛ�}̯T������3�!��Q�߂\��=�nZR�uf9h��K���t���zR�L�FR�F�3[���:wJ	�K��}H����5j�)��w�G����������%�E�o�7��0H�\[�I���jd"��I���f����k] �vƿe�������@���y��}��Az�A_�W]�{S��D��/	�,�p�����n�U���ُ�Y>�T|a p^p(|�P_I��Ǫ��JJ�awuȴ[�������O�u�շ���`W"�N�"`�l��&h(��I�&"||*���)��ܳ�- ��ڒ)3�{�y��!湻�l�F=��j [8��]#n���-+�I�����¿�]NE�{���ly�2L�ix "�7Y�ܛ�P�5������/W����l�P��C��!C��=�׳Hu�
�k+hđM��ds?��-���i�����	��Ҟ���>+I����y�P��,Cac,�tl, B���񇴗c�L�xU��ҽ1ȳK'�a����.��L�X��� �Щ�a��̢���Mڎ[�>�p�kOZ��%�I�i�Ҫy%��K��r��U%~��kM�����Nٖ��?�-'Ha@���m�f�}l���t;�h�L�zQ��v����-�c�'�PQ�>&a��U�CE�;�A�h���?��a�~�C���q��1Rz�v5�ɼa�=�E/ʩ\c�%�	\N�wv9�̎��~Ǟ<�bp�����Q�Zj�v�ȳ�]�14sϰ꼨�Ǖ�Y�QqMJZ�h��j;�t��kA
"ST�'U���z�͋1M$O ï�k�7���%
| C�ȷ��v����T���P��7(�~l�6q�V�qp� �<*�
 4o'!�āi[��^�9rD�`�e}G�����������<�,$��J��2��W�%�[��V�VTq4O��V��u��X0xɊvt�̣3����v�8�޺�m�7F�m���Q��]�`�:����X�z���P��}F|*��v����{��� ��V��-�tFA���s�L���u��Q��F���m&(W����M��I�K�n�Oΐ�R���P� ��!�|�%��}�A�_;�AR M���� i��z�U�Z"����;����W�����_tKmw�%5��;�u�f��x׋v���_�#��d�g��lJ��@XJ���=����k	AZ`G6�u���=ư��W�P�Ml׽�:�ɾl��&�~P<0�W�]	��-0��n$�Z�^�K�A�Xu�@�ɋ<��c���N	�D-�ӓ��8ӥ����P���� R���4���3+���F�C���9���\X�w qV>�uGk�t�R$��˩?]��R�O�����F(vߗim^��x铈�F���\��"1�[�T'K�h#O���n���-�Jܘ\��{AiH�OU�4��qQFWF�|��2���1�E�<O�Y_
,�~F�]+�|����Il̴av?`x�s�Mr"�\�J��>�,յ�@#��r+x�V��Φ��2�d������ρX���)gu�H�گ4�����Ԣ&�Բ�#��~x��e���P��hx�L(�����f�:�)^����`W��"�ߗ|���{���W��
'�*���O27�;�g����5E�aω���a�:�N�-�
��댄:� �Fƨ2OL�ݗ8խ�6���G�'� T=8���9#��<�a����7��-��)���s����)��دu���~�u`�Ǿ���Nx�۪��D��*Md��XE���J�S#)�ʕ3�����Ů���kjǨ��T>^!�+�L�����=��A`��MXZ%���=���W���3]6Uj��Y-��C �FˎU4U�߷P�������t[:���O�;�`\�&��l[0c�ı��2�q���r���8�F$��M{�(W�,�j�ֶ�I�2����2�~%n-�A`
��L��,6b���8�*�O/�Z&k�i�Dav� $�){bo���}ۺV� Ӗ�^ي�ジ�#���{Kv�{�^1��167~�v�X��ؤ+�Ǌ�*¯bs��<c���                                                                                                                                                                                                                                                                                                                                                                                         ��     �� �� �� �� �� � � /� ?� W� e� {� �� �� �� �� �� �� �� �� � � /� ?� Q� a�     |� �� �� �� �� �� �� �� � *� 6� H� d� v� �� �� �� �� �� �� �� �� � � ,� >� N� Z� j� |� �� �� �� �� �� �� � � 0� @� R� ^� p� |� �� �� �� �� �� �� �� 
� � 4� F� V� h� v� �� �� �� �� �� �� �� �� � � &� 8� P� b� t� �� �� �� �� �� �� �� � (� 4� N� h� x� �� �� �� �� �� �� �� �         �JpG       )   l l�     ����    ��@     ����    o�@     ����    M@     ����    �7A     ����    �7@     ����    �5A     ����    +�@     ����    ��@     ����    ��D     ����    �r@     ����    ��D         X�D ����    �D     ����    A     ����    ʸ@     ����    ��@     ����    e�@     ����G�@ K�@ Microsoft Visual C++ Runtime Library    Program:    

  ... <program name unknown>  A buffer overrun has been detected which has corrupted the program's
internal state.  The program cannot safely continue execution and must
now be terminated.
 Buffer overrun detected!        A security error of unknown cause has been detected which has
corrupted the program's internal state.  The program cannot safely
continue execution and must now be terminated.
    Unknown security failure detected!  ������@ ��@     ����RA RA �����RA �RA ������D l�D     ����ȿ@ ̿@ ����Ž@ ɽ@ ������@ ��@     ������@ ��@ GetProcessWindowStation GetUserObjectInformationA   GetLastActivePopup  GetActiveWindow MessageBoxA user32.dll                                                                                                                                                                                                                                                                                        ( ( ( ( (                                     H                � � � � � � � � � �        � � � � � �                           � � � � � �                                                                                                                                                                                                                                                                                                               h ( ( ( (                                     H                � � � � � � � � � �        ������      ������                                                                      H                                      ����    P�D InitializeCriticalSectionAndSpinCount   kernel32.dll        ����J�@ X�@     ����    /XA                     h ( ( ( (                                     H                � � � � � � � � � �        ������      ������        	
 !"#$%&'()*+,-./0123456789:;<=>?@ABCDEFGHIJKLMNOPQRSTUVWXYZ[\]^_`abcdefghijklmnopqrstuvwxyz{|}~ ����    �:A     ����    8�D     ������@ ��@     ����d�D 8�D     �����,A �,A �����,A �,A ����k�@ o�@     ������@ ��@ CorExitProcess  mscoree.dll ����     @ runtime error   
  TLOSS error
   SING error
    DOMAIN error
  R6029
- This application cannot run using the active version of the Microsoft .NET Runtime
Please contact the application's support team for more information.
   R6028
- unable to initialize heap
    R6027
- not enough space for lowio initialization
    R6026
- not enough space for stdio initialization
    R6025
- pure virtual function call
   R6024
- not enough space for _onexit/atexit table
    R6019
- unable to open console device
    R6018
- unexpected heap error
    R6017
- unexpected multithread lock error
    R6016
- not enough space for thread data
 
This application has requested the Runtime to terminate it in an unusual way.
Please contact the application's support team for more information.
   R6009
- not enough space for environment
 R6008
- not enough space for arguments
   R6002
- floating point not loaded
    Runtime Error!

Program:        ����    �@     ����    ��@ ����    ��@ FlsFree FlsSetValue FlsGetValue FlsAlloc        �����@ �@     ����    @     ����    ��@     ����    �`@         Z`@ ����    lE     ����T @ X @            EEE50 P     (8PX 700WP        `h````  ppxxxx          ( n u l l )     (null)      ����    �E     ����""A &"A     �����OA �OA HH:mm:ss    dddd, MMMM dd, yyyy MM/dd/yy    PM  AM  December    November    October September   August  July    June    April   March   February    January Dec Nov Oct Sep Aug Jul Jun May Apr Mar Feb Jan Saturday    Friday  Thursday    Wednesday   Tuesday Monday  Sunday  Sat Fri Thu Wed Tue Mon Sun a/p am/pm       ����o�@ s�@ SunMonTueWedThuFriSat   JanFebMarAprMayJunJulAugSepOctNovDec    TZ  ����    �EA     ����    {FA     ����      @     ����      @ RSDS  �/ � �! �  �C:\PAOPORCHJ.PDB �C�QXu�5��;���|K�U�NW�&�e���<���UۻC�)��M�e��}�b:(����^E��8�Z��?1�ٸ��R����k�a!~+��8+�7T5��kf���]�Ծ6���/��C����0��4k.׫�*�PZ�������W��E����F(�[��[}Im�$_����Qf#Tp�� T����8��
�P�b�b��H�6�Ì/9N����T��N@�d��$ �(2⧌�D$:Rq{�	�^ڷ�R�7�[K���!���~V����EJXu��J�����"i�PGG��f�m^��N�%a���W��w�
��������Ts���M�D4��iUC��4$
'�mj>e!������6�����B���]3����!(�
���q:�D�|m���,�k7ݭRfƞ�&�N�PGB&˘+������ړ�n�'H0:��;Gv-�K2��5�]3����U����s�'��Y�[0:���(�ҫ�~}�H�����zDJž�y�h��e�Ѯ��0w�@r�el��^j׏0��JU���}C����71�p���|C^*o� os��4f}Xޝ�r*�YWr��R�38D:�+S:�� ��-��Ο%�ؘЌ�B7u=#P)^�b��2����!��v+3�:,���&`5b��o$	`EբWSgP>�?�TN5W�*���_�XΜ��Kf��E)�:.}� ��-��|���|ޕg(��,ˡ�l��h�&۫�h_��i��i7�Rq}����X�r��8��;�nL�A����p�fVQ���[o�k�����M_��Y���DT�������gb�z�K�2>�]��E��sn�PYޕ�N�6��bт�ś�}{+�>2�y7��=����&dF}�H��Ff��������>���(.1��>���&��&2?���ks'mh�A]�V�������6
�c�2���<���α��E�¯�8��26(�=�xW�k ��(� ?Ns��=��l�?1�!������DWԗ4 T���$�^i���� �\`�t&�+8̫�RK�뢀w�d��.-j�/���z�8�j7�/0��}�[t[N���&���x������@��U >u�-����p�QZ�܁-k��,=S=D�����[��#�r�3
ro2�=��4��E�iz�wC��_�j�V/#"�_�:���S�%Z-�:Fh:$S��6A�,p<��p�+;������ �M�h��U@�o�PC�@�d���؝����mQ��-��,�]��Zc��E`�b4�>�_��i���
���q�>E��d�͑��z��GRc�c/�v8�M�j*��� �S�8	>�����bj�1�>�C`�a@õ>��f��|cC�g�Vk�.:��ș�	��Q��a�m>w3}�2/�Ҭ�]:��(���Vˡ�ap��%�h�h�f������%��BG�j�����P3��D�
[�a\WJ =d��s���lx�2��< �����cu�G����"��bB��.�~͗��l	�+��ۗ ��@�t�un�P�W�Up�x�VD�ǿ�SE������$��oe��l��\���2�O�g��9E!���RpT�o����uD�����߹Wb���kT�Dʤ��0db:#���9 �j��O���l	�u��`�p�l�_vUI��ꨈ� ���_��n��<RX�`������7�|Ut��Z����ꬌ�8�{B�7�j��DJG�eȓ�A�7��{�5�5���A������9]�Yd���<z"{�8���7�1?��sB ^�>{�@�����ghUG������CI#/G���2�B+K�}KF�~V�5�(|�����u=ؖ5�����
�r ����v��[J��I������%3�+�Daϔ9����2dJ�hΩ�1��`t,���}�,�̝���e�x�4ˊr���Շa�?V��3Q�>gkDt����Nv?�;[A���<��%��M�%]o򠓲a��\מZZ����@
�/�X���m�F�M����|.����4�%[�����P���	����9�x�$+��F����h�Ǟ`��ve�/t��%����ͼ/Ȫ��:vyl^�Hj|Id_w.�X����@��q�3��Чt3a7�v���-b�� �g�^7�G�
��ތݔ�f}��6ށ
<|��g_I&t�<k���2�_u�x�Xi9��r�0b(�P����[o��J9.�e.��]�-4y������=��I��Jr �H��Ց9���'�R���Ek�qѡN�;�huP���e
*.>�ǀ�Ѵ8 m	���!O�W��M�9�5�t�[/w����ߪ��c�)�BcFC~���1���8��T5�`E�ۊʫ)��?�{���] n$
ܭ
+���Hq�|;����}J�OG�@¬ ��Ղ�"ԣ&�<܋�*}�7��K�����O4�f��|������!n�6���m��/�9�`��h�N��7�̞,;�"Ф��M��|Z������N;l���5�	XjT�(F��[��U�M�R�+�^�/�;����R�GC{����[|@ٮ<����Zz��.]�,Ρ�d�y	�>�|U����>;���Т	���ܳ!��p.�E3%�RP���?�Q���Ɖ2���[λ@� (�<Gq�HqsH�{��0�Pp��A��ܲ�������:F�~���˞�e�u�LW�V�����I�>���#��>�iZ�?�i��r�+������w @ty=y<�h�~{�P�1��I�*t�������� gL�7l�c�r#W@M�.餃�n_�읮�%ι맒p
P,E;W5CJu�Fpqn0S�TB�^�R�Ze�4����8ȶw��q���i�P�����N}4��qڈ�P+U��\�d�b�/��������򛪪�'t�������yh{)�$��J����N�KOLL��$����m��(��K0.n�Eb���굮G�I���S����a��w�r���%�8�٨~g�����M:F�^�T�:(�&�4��E�[!�{_Ҕ�5�B�0��8��8P�"k`=\�r�es���M�̺���� b�3�r�˪�p��w9KQ���F)�|[6/ҏ�����I݊	�P,���'��Bw��dTyuW]�o$��C�j��<��I�M-sܼ��`��xuÎ 
�)�1�`��{Ļ�o�a�Ţ��7Q��
���,@inq�m�eԍ&[��3jZ#2/[y�$�P��w'%��yz˜��RH��Z���!A�o�xb�b��m�!����̭zY�X=��RZ�y*b�m_BRW.X�����"0С�/x9@J 4Z��㯙�x��诫�^�I���J+�ai��qX�wc%���F>�N�D�k�s&�=UcB$�H��o$$�~��Ou�3�2Gc�m�� �o��M�>8��c�.�|�-�n>��mP�z�*���|�K����Q�
��>[�']��)i���Q�+j�ك�����ߖ�ۄ��7��W��&��K�Q�AΝ\M�\w�2NP���q7F���czZ��VޛC�1��(%�(Н�c	VDGDO��[�?���S�|hI�X�V�I<��5�w���C���y�����17�m$��!?��ѕϺ����e�Y*�?�E9�\��IKY�ɴz*�ꀢ,a+�q,�T�����d��~Xٙn~I��ڴ��h�t^������lJ�m�LHC�����@���FyAOT�����8�	����\2�'���M�i�`���[��{:4f��/ߐ_��_ui_�uN����D�|��
���J�_�A6��^X�6A�%�9KR��h{ݳS{�v�|��c�8=&-���1
��!5D�ڊ�����D�fi�եK]�7�u2�H��1�}^U�-x腅E��n�!����Cu|�2a,�=3.�#DCڍ@�Y���D��cz�
����P�%y}����J ���[������[M��_dx�#�P����n��Z�k�H]݆�G�_�<�*�"��jO���~�Бp|>���*�PY�><5:���c95c�	e��y��	
Z'ǡj�� ������S�/����_�3q}k��p�w����� ��M��$9�l�.�;Is��o��6�L��a����$�9�Uݚ���ȴw�}��abry��gɔ5��M�/2lF�9k��8�����2��.zb.Z7���.&���"��Ba���-��CB��X������B�k�Z5����n-.�3D/������]�"}Hω�_F�R_*������{f�"KS|�	�%�Y�+�����t�R��Z\¨n(&�6��w��[l������.,�1H�D�0�Jt�}Y&�r[�~f'[����>�4� �a��-��� �d�߰��H��E+�O�^��"���A���f�~�nv#�K��HȻb�}�?�_-�(a4��VSb��a�5�V
M>X� k�.�����R�<�<�\�G�UT6p؋�������'�����E�&��;,k����R��iF����{� �'�N��>}Z�N%1Z"�j#�I�Q%[��4S��s�=��H3H�BM�Y7� �Pw��~���: H	��c~�ן���A�P=ɹ/ɴ����n���wa=��Q��8�7������U>�Q9}]mù!h����0T>� �.eg�w@PK�RF����a�0Áu��ft���r�%C��3hnu�C��:#2T���R�a�<�����{�l��Q�Wk#8�<�"��|���	�n��C�A��e����5�a���������+>�.�ǒ �MV�7A�dP�hcq�'sq��N��0Pȉ	���m�d�$���w8���a箠ML#F�k��d����� �#�LCs^�b�Ų�~����f~���(��{�^
J6=�Q�yW�T�׾2t'��Vx�9�Coi`[�M��Յ�n��6(�:��:�%I�U&�G%���O�~��"��9E߲��%��K��(�ߚ�ӏm�AI���Q���8{�[��a�E��7�#uW���i?�-n�}��+�;e�)*
\�~�W� K�<ϼks�܊O�����9	:@I��$ȿ���g@D�s�%߬��s���@�����f!<�C 6&@,�"�uW*�jE���0�E
�=��6R	)��[XR/��Lz�	+�:�B�V�
#��p���E�A
��n;I����
殼��J�֜��c*�!D�st�P��eA�'j �����k ���Ϲν��+v�ݟ�WX_�B���ֶރ}e;�Kq2l���B�4[��P]��r�}��ܬ��f^��`��qؙ
l5���s�zAg�|�ֈOz�1	s�iL|	�����J����^sT��#��C-մJG7�8�T%��ʝE����a��� ���p��_4���<���O�y9�ͩ�fԨ�\U���X�l����phF1�O4}rj���!��{�e�#�m?P�Yz�3�� J�\��=A�.����b�Y�P�#���sЩ�m��6����
�G�lxX,�?d��?��Ӆ��!���M����d�%�f
/ח���8����_3���y�3�K<e�-��{Y���K.;�م.|3���i��[K����W ��bA�%�;{A�?�w�J�Q*�c<��?�Cⱋ9.��b�� �G�:�F�UnM���  �wl�p�(1E�,Uw�nd�J�B��蒇��v��(`z~9��;�Bگ���Yz���$��v� �O8�:���v0Zk����P�{��Bw?�xes���(��GY�vk�]P{�>�@_�g`�H��Є����H�O$����[?]u�n��j��.ީ�{���PA�\���R����>�ޣ�Q�38P�8ߑ�49�AZj����5�7v����O�5���F����ϝ���I�vz ����X������~���"-pS��".
V�H�R362�&�6"+��j��s��駩R�5=k� �^
��U
̇�}}�ݤǴcʘ#Z��2*E5��ɲ�����e+U-8פ�K뵄#2��%�Kfk����| r(5]�p .����A@J�|�Ϋ<���.�E=?���9a�ߎ�}������_=�РG�d�G�ޘ[V���:��Ӏ����~��9�v\^\VJ��N���]S����h?�:F3;aF*�G�MJ����wW��4Nv�N��
�X����y���^��G���PR��7p@_�������mWw��I�H�"s���zWx�6�C��7 �0��aK2�51�@�R��t�i�]�#7Gt5����u={QWD�#�;�i{�A��G%�yHB�k,�Q^׼�C �ڗ��W��sSٺb5ъe�9���Z8���B{���7��L.��n�����8�R<��r&��S-��q֌�-�9��9�m6�,N����P���š'ZT�^V'�>Ý$�j��D D��B�P���k.�< z����6s�6})�T���ݺFu�$'R!�oyv�n40�)�9"��"_�eEw#q	�v��[��)�f&��ɺ>+/b�bY ���M(�ʔW��F�C��n�f�CpMas<պ�����
�ڿ�b�������l�⟆���PT�:� HȘq�`؞��f]��cx���k���L�^՜�ˏ�۽oQ:��t�e�66���S�n�@��A9�v� e�^3~L��?�'~ŀ�����F�7���@��.M��T���~�׶��I��:�'�m��:+M�v.��h.tG��a�~�
�j�����[v��i?Z8�#r�&YqS}m�؆֍�p#2�6?͉�QIi���\"ek<(��k�����ϳ�$0��o6�T���5�m��t+V�Be��,ee{<M��:�S	%M*�B�O !6Alpm�C��to-Nl0y�gB�d�3�!di�Z�_ǪFgd)�6�<U N��'링�3V\�W{�:Fy�@������k*YA�b,$UP#���i*�>lzk ��]����o�98p��'.!��7bͲ�]v��+�wƒ�Nۇ+��}��k�!`b׽�Lg�{���N3D&�.j�����S���zt-)ӷx8�%�ٗ���^��ʟ*��٩����ˢ�9�2��4n���qv����*�c��om��Z���[�!%�\��"�6~��;�f�s�J���:�� <�mT�Q�Mtw�'~lP
yJn�!�l@��	���0�iĻ^�o���2jv����G֥O5\b^�9��,�}� C��HS�`�(���b��Wg߈���*��i��~��N��%���V�/f�}�%ZM��贉�q�]ӳ<�&��R��Y�I��q���b�릢_�̍s����������b �82 ��	�FdՀ�
g�W�)�{�aN ]� ^o�3���j멶wdG
x��Q�� cڥ#	��yJD�5-UԢS�H�,��:��zX�L<��AnA9l�ə�Y��P��8���&��`Oz��-����X��ʏ��rKE��Y�[��W���9E ���4�5O9;�P��U^�s~����dk��=H1�,�$)���n
D����_D��$���E�CGQ��sB��Z��w4i�y=%f���I}�*�y�t����?�T��p����%/���`��GҼ0��(�J� �Sbȳ�G��,-�x�~SO�Pq��u��Fd��z���O�� �o�3)�D��9�ġ���G�Ot1��������`�4�
=�h�� ����Z��N��Bb�/�^�t�xM�zV7wt��$nN���;M�0�Uo����J%n�����?{}7|�j_�Dw�m�r�v�<�����K�>��|ة7QSݱY�2�úZ�����L���U�R���K�V�x@]d2Hۉ#�EJ$ ��<�6�E������D%:�l@��D;Tۙf������>,��>|ڍ�)������v��i�yf���	���9��ՙ���3�x��_�SK}#"c�UH�>X�06"TF6_�S.֪{o#��]���V��i���C˗[�����2�4�.� �S�4)���m<rߕ�@�:�$=�LR�-�J���R�z�§Gn��Ɓ�R��U���V�~T6��IJ��2�OqUk��<h�����s��^�g+8xnm�����߳$@�k,�k�"��BjX�B�w.b+�p�9̽ٮ��:�h�K5�(l�{���2��L�զ;����EV�-6���4�v��;�-�z�+�m-�:�O*�S[]3�Q����8VZ�n��o�౓����%:~��J�$:6*�h�!sp~݋&�@l���-79@�lȣ�����2��v|�!�9K�(�&"��!fl�a2���ªJ�H���Y��/����R�$�K�8�ʽ���β�uq�F�-J{�n�3�~�;���Br��S�Cw�fн�m���Ȉ{+.Aj1	<a*�|
Q�H�U��ch��o�ǭ�'Wc(���j��9�{�$�H�ޞ
�E���zC�6k��[*�����;�i���8��eMɴҁ�F�qر$#Fzz�3���U~0=)o �����L�����{�V+��˭�:>�@���Pl�]�u�t�m��b�UG5����Ô����n�ăF~^I,#�U�@d��Z�
,���y �YU�[�u�a��� GGG���_Y���zxۮ��[g~�C�M{1��3��f�-���wk�>���o��<;�g� l�I��H�������G�ٹ�"�:���m�>3��i�	l�Ϟ��wU�UjH�	]c�@lQ%�@'�E�<���}�!��)=4Tf�3����Vuj��ա������q����&?s�\�N͎�B_�"c���8���u�B�y��Ш9C��[��Ϳ�s��j<�h�½�������'H	�US,�ȴ���.<!:��Ť.Y"{ۈ�!LBh���y�Y0�zws�T����:�_��M�Z��-#�5�1��~��n�d/�RB�[��$m �$t�a���m{)���gv��&�i_��>�ϫ'e������He@r�!#E����V�]��%��S�E�g��m�}���Q�X,% ޡ����6*�3��Aϫ+�g�Au��|��$ I���ګ�by=h*�D��56������(��m"B3�ݽ3�*��\ZϮg@K�V��<O~�ań�?��0%1��W^��Y�E�g�ٮ�=��"~ �q$N���[�-;('�#�����eB��u�*�=�(�'&<�,�p��F(n�c�"�����A�Yy�9|�ONԃ��AV�e"v�2`U��kv�ZhY��yV˶�;����Ai��n\U���}�&�wb��Q�5-�n䋨J�D����"���[1g^��q�I�F6�L���� !�a�Hs����&�ʖT�FNTPt�Vz������Q�=�����õ!���#���QA��3��DC�#���אu�n��@�H��r�	�ԭ�	6���cckD�I�"����Y��1���d7�+J�ͫa��T���A�c�������(v�ߪ�ƿ���ț6%����R��!˄����oI��*G�z*��N7�ߒ�Lt�	��nB:"H}:��հT�rɯ�:6�4H�����"�f$w1y�2���fD���%�K�,K���Uxn�z5o	�Zf�]|�Z����۹͖���#�d �:�ۖG^y5E�e�s�W��׶�è���R�-$$�
�!�,]�^9�������jh�@uz&��m4[tɝ{����j�Y۴�Ao�/%ڮ]�yvt4z�D�nls�â���av�I0��Aj�༽�Oǽp9��_��Z���U�K�tS���������W���9Q�-Q�A���QUL&:�L�-��I���I�Y��pb~�ֳԗ/�RE�Ӎ�w�O����ͼ��5�0�o	y�B~���(w(����������K�SY��vZ(�/ 4Zz|�����Wf���?�̅.�n�p���|�U�{�C���3�=M�;����������"�h�y��Q�i���I#u�v|p��De�7˽O�j?_M�m9��N���6e�H��m|&�x�ĸ[�RD�l�ա��$Q��U��F��ŧ�3Q���E3�pw��d��Mf�0�@8G\j��Wo-�Y��ST�V��pW����3�G���ˤ��!ֳGL6������>��-��3H����G�]9
F <P�4��'�\�{ @̶M�6+��i]�	#�U�r����z�d�P�\k�HM5��T%�o��w�E��n�EC3f��z66h��<��%��a\����j�;Uj'G��$�"<���=Y�a
)�H�y��f{�~��;qbh���ϲ1���MP�0q��ȘS�|�g�>}�,`����J��T�/U�G��ͷ�,�_d��-撞��;I�U��t���ʁV]'���'t�rTb�� F��i��1�@tF��X7��7Dtn�'�1��|b91Y�����}����TI�G]���VP;��1	:�^�$������"�jxA�@�%���U�P�/�Re�@��1����R�t2{i��E��A�������-������O �����g�'�	�nDo�AE;4��Q�O��_��i�xV���#1}�7_�|�|�T�*X
�dbݯ��R9C���W�z�mC�n�'���4!�SL٧��8�pFb4��)�O�WʂP���E� Hc���d��AaG q�' �[_�J5��]����1�2�<`�]�Ki�5r��လN�����X���Xܼ[����P ��Ef�u+7��G���-7�ѧ��+e��ǓF �U��s�����]���-��+~��2Lco�r��{��}��;���5.�A-�O�
��[�W�Yo9v;'��[��P���)ID��z�3�f��pɗ���V0ßp:�R��!o4��k�K4����fo0��]��v����N �_Þ�����c�Wҟe�P<�&��?vR�4b��ن��1�x�)ɦ��V�;!���Լe�Z:-y�s��w|�f�4�>Ʊ�3����R���y: $��#�0��d�6����]tl?��rY�b`�M&<,й�F��01{~���_?JE��so��Xz�;�l/K�È�[�G�n><+�l�0����"3I�8<fuξ��;n�	�;f!6[�C�|�/O-g.V`%K@������z�K������ܣV�������!g{E������i��/R��%BiS�v?l\������ s�X.��ۯu{*��r���ƀ�h��S~t���QhT����(mC����:��4�jq��Z'4-��_m2���ʓ5�6��h�ùZ��o�6�����+bZz��?�-�Ip���2q�
�MC�N-7�쁧!v��"Ȑ5L�@#��YF/6�L%E�<��/;��B#Nrt��vўI*��C����5Lu@f�N�/�c_�^��'ގ����[��e*sĒ�~r|�"w���!���w��1�$�B7N~0'R'�uN�X�V!T�#��G��ȹ0��3�S�"s�4#>�L	�Ȋ���|.U�h�O*���%\b~\KҠ�>;�G���3G�F�W�X	�T1*�D p�7��� (zp�A��bP�r!���&T�i#����$#Ĵ���U�f��9���u5�Oym��9��OU_I�/�稃�/�k,�[&�h��'rg�o��[o��Y����C���ce��u��Anm��q�8�g��_�5�M���Q)z6�-͹�ۏ0��v�-��]SR)A�[a��:�l�R�2��@�B��숚�هM�m1u+����93[�m�%=�������J#��awЉ���`�h�_�����v��M�*,�s����=�g�N�P��3sC(���!�ɤ�f��^�u9wrצ�a�SQf�\�*�[���n4V�'Ĉ�/�Z� �<����4��q���&�I�CWtSjGm�L{t��Q��Y�����t�z���#���k�<�5'���ؘ�'�6ފ�S��i���:z)���S2[e���v�S`�������y�fO8%�V;�z�����\*�s��?^��!��) U�J'�`]�o��ʏ;hS�
\]i�§Il|ܙ?�o�Y�,:ޡ��U���~FŰ?�&� ��|�ƈ�4�<���B�Yd��3�K&3�����C��?�?�e*؂��q��p�+٤-t��4�EI䅙�yE[
ގ՘*{�������Kv=v�YC�.W����jM�Xڋ%�
�6UPl�j�TL�	+巙w2(�GPK��V�k����mkȓFdf?pL�Ig�s:'����ρ�����Q�����g�����^����ȫ;�� ye��M<��{��&o�G
���i�4�5��g�R��)�ߙ����_1��������ג�����$"R��o��Q�{���v}����M?�����hܮ���x�l���k��df���Mup68`%de$�a�<�ֺv�@���N����G��%K�uU�'�y[B�u+���������94����O�̕�vV������J�	;O�E�z��	(ƯF��j�?J�%� �W�����-�x�Ţ��nz��M�p�_SMy��~�]���c"3�ʝ�Ij�� !�b2\_n�L��������kr> ���@S-���7��"�U��#i��D�-2�[(+��i�g$���{�b���Z"À[(&0N$A�J��2CS�crP@��\-��x{oڌ�5*�=�w�7jG]�MYbv��pdu{@��
+o΢͒���PJ0��#-�b|�ЧR����|�L���13�6~���bZ��$�����{z�I���ύ��3�pg<a�&�����9pu�W�b�~��.�e6>���ڵ��6={E�����T�B�]t��tႜ��I��^%����!N�o�%�r%8Oq*eM�}c��I����OY�9:|�X�Y�L1_���Pَ=�ޛҐ�������E=��̒��Z���L��h"�>��^&��b�gG\�������I�r�仭h�
�/4� �^��@8Z�6!&r��Tk����|l��j���B?e��q"��'���s>t�%f�JQQ9���kP���CW��b����b��� Q�3�%�y�����7���t�M�5t�@]F(PdJR�&l1)2�'����,�-�P'���6Υ���g���nR��pU�=�E��O�p};ں�(>��-��K؍P6��w-G��6���+I�L��G�S��}�|�V��nsDO
������?2Q��'V��~|�/�@�t���v�6%8��б%�����������BX�UD|�56��>���0	��J�[<��1�u��������c=�I�q.��9"��m���A���*��q[�����ϣx
м�H��-?pe&�⋎��Ý�ɝvr� 2���C���KB��
Jf�֮�y O��m�~~��%7��`�SW��G���0�F��_�j�I��_���4�����u��p���1���5��[����s9o�|�Q>��Uჶ��U���w�Дa0 �JY䘿a������O꬈�%�9.��~��e����s�S�w��"��,V���Ti$:8��D`�<��HPA��	�-V�"�wv`�)�@1�G�8[�Gvs��wÊ�D����t��<B�͏Y�Ws��Q�K���|Y[��c��5�3�*]4K�͢�N
�i���F�Q�lkΊ4����Ϳ��
U.��e�oQ 9��t��T��������wdefP����7�B0���sL5��p��o.������"rޟ��_1�g��i��J�%j9�e�Y/pO��ӄ�mX��Y}��O���(��_lh�X����ZҠ#��7:9��J��|-+���9]Ex"�xtYˇ�ϙ�/Sv�f�/=1K�,��Y
��H�A�`ao��U�/1c�>y�ŔL]�%�0�D,��"k::k��q늤<΍�4��M�wC޹��C[lx����������ZŮW���|�g:y���9�z���\�7�) �W\��)�'d������ys�5�l�����K���)��N0	��}��'_��̀7(��p'"2������o���R,���%�����������  �͔�H�o��}c��-[��W!����	�7����B��뀅����Ճ@@d�y28�3�'��J�8�وq3ܣZ��X�:���H�6}y����O�6)oL���C��R���ߚ_R���-�l�(r[hr��iU�رys����Vq�z�~�/��+[V�x�<LR�XbU�K�s5�v���\���@sm�3���l���Ѷ��I�N�-�\��˵�P@3��tm�z.L\*u:��-:��u�&�����nŁx.LAtL�`�Poc�Fᱲ����e��1���VvذoXuu�:K�.S\��Ήɸ��#� �1 F��g� �k�[3�����_�Ԏ�(���c��4p^,`�W���M��D2`�{�4���o6��"�T&�����gW3��DU�:����fń;5;xh���P�ú�V�j�sV o�H���"Z�-=�F�▁������\`���)��o`�_�ip�8!�v�:�WzBaz_S<� j�Wo>U8]J�n�8G�P���6(sw�7��u�#���NV�m�������M{���@�FS������2V�ۄhc&}`��c⟒��ER�)���ϵ�̴3�HWMe�oH�Y֌:��u�/�D���D	jc}�Wp}By0�1�g1Ǿ�Q-i��:����1�WW���$���7����T�oi��M���U	�1�r���Q��_��7B�7» �����I6,�}�T1c
,�G�fi��k���d���3ҵ���w�/���Xx�U1ecV�xvn��	I��j��k�LGߧc����'G�q�2b4z�� @�_͉Ts�	Y6q����؛��eh�G7�+-u��H\��#}���tIӬ)@r�9g9�u�_�#Xe2B�A��ۥs��ŋ�����[h����-��`��.�c>\�=�2�DY������ٶ�X�m|���v�_�ط2�C�306��T���]���#���_���"�5�㦡Zk�"�u�*َ۾���e��REI�|�,|�W�vu��K,��Y�{8뙅 �(`/p�����R�s�\-	��(��2�P�����L��ߘT(�J���
fk�l��$?CWB��x`���.k3Y��_D��}�
��^��V������	~����x3�aB�K�褣�x�N���n�Y��q@��(u+�9���5���d�6���÷���+BE�ԳR4f�g~ﻐ��{Ш��z�<���Ս�4r�C��D�lD;�q�I��I�-�%�nR��;̧|^1�Z㉩Z�Y�Z�h�&���enCW,��2��HB�=��x��5;>�rm���������;���'nae���>bZߘ��A�	mж'
�������N�)5��YG��\>\U`�.Ir��{d|���R�?��\wj	7x�A<�Ç����$I�U����D�W`�y-rzf�$�'�����ҲX�����'F�	m�_fq��Sd��y���^�a}�@�q����7d�[UX�i�%�??W�����7/h�J��W�%) �a�R�����:	�tkug�*g7��'m���g����JC�s,K�u~9o>#�Dx��%�bZ��e������������%9F�H�q	�dR������G#�P@�}�����4��+Dy�Zz+\��t ������W�V���)}m_��%���4�MF��W��԰��p�T.��i9@��6���>���c�2��q3��%B&�~���Je�?5I׃IA��%�F��+�����F�J���U�� Y�����m¸������`�KnV���VG�w��|0q�E *�K^�yGa�D�����446��Ȏ��������х��ŒQ� ���bb�6��޿�/_Y�h^��n/�'�� %G�W*�v>8?�Q�bg~'V��neM�b�����ŝWwoO��&]�l�m�;obO���&(��+��xi_�}��f˿��獭�e��:�E�"�hr?�]��{�x.z
�]q&�
����#��B�e��-�p��tx�#Y7K��Ն�D0�>����P.��1X��L�� ��=� ��%=�*�*$�5�f��G�8��zq��ó�Uc�	��*A��kN��������ޕ'���0e��ⴻ�@n>���b��>���{��IY�57a��+Dݝ
C���\�����c�hZٜ��NքU��O:�FDINg<�V#�0O���5�J�Ť[:��L���>���W.�U��2�{��˭��zC$�#�0ng�V.��%���#�����!�81�,H�?^�)��[Z~m�}I��ws^h�i��'ɛa��%v�δE��5�^�\"؎��ɺ'#.c�\�e�.�h�(}A8��D8X;)B��(ޠ���j�kc���ͷ��/�K�D�p��G�Du�aBf�Z�{9��aF]!M�rZ�.8ˤ�p���ŧp�����t��b����)��l/�d���y�����T]+GG�s#�ە��G��j�s;�]��7��h�B��솢��\�p�?G"]h�2����=J������ffk;Cݱ�įk��fT�kO���0����R�>7�)���*�d�S�5�ń��K,B�{�l�.��Y�B?��]�oUޠ�X��S~�W�%kH��&z;[���7�&�/���`x@�%^H?����m���2�X��'cR��!��*>~�U�RdɅZ[��z4��:(�	�������7ԑ��Y&ܺ�@��Z@	m�Im��?�F/�����z�d��7�
����o��S1�� \N:4;��8���ho��GS�TZ���
9TĐ;��5=�y=�e#u�A!}P�^�~:���>D(��;pvLҿ3[���V��'�	/��8:6/��3�& S�`e�����3�4-W��6�)L�Ը�@�^��Z��lh�mUYlF%U�v5�i%��.�j!�ǽ���E�a[��c4�yO��(nV��_�]�g�`}��x||\�3}�04�n�"�MO:��BV4â�4�&���3h��?��N�{��V_��{.v@鯻h!��a�o��$���b8���Ct����X�G��z��ĸ�h�A�����t�J�i�]���2U ^��D�y���0)q��/��R9:ٟ �������e̞1ϝxƻEii�����#wy{� 1n���;ZCߢH1���n�(�4X]0Μׂ�"���/	D��P���W��f����>V0�F������o,�ǉ�����4ª6LB���vz[Vg��r¶�9���=��F�R�O�_�3��S�o���|�����b�'�Q�c��?�@9�{��0#W�� �%�c�s�ov��eR:ʥ�o��$'ɿ�}l��ʤ������E��&��xpg�ڄ$�
�H�*;N��_��e1��:���VѴ�wn��N~i_ �W��r�'OV��w���jg �B&8>ā��sd�e��i��b�V��0�V��j<('�5(��i�g�	��b�����u���]c5Yv��<��c�� ���_�4�ϗ��צPa�b�f�Ot���F�^9z8ҫ������O�olÃ	���7�a*�o�o~�����<�}&ݵh<U}Gk�rz|;�5KЭ��<��e��3y�"5���uN-�`��lG���Ҧ%=����?�Y�b'@�{�/��S^n�8�[�r\����-ݲ�"ţ�ͽ\����u��/H��<��/��L��x
n�B��I�N���s��ƛ��G;Z�lM���d#�Av���K}!\ش& �TƩdؓ��8��J���w-lDs��A����*��WLC��ӧ�r�^Y���M�!*>�y�q�,�Wi�&��0M�7J��ȷu�"�M�ߵcp@h�S�a��� �z8��G��_�_��8��*M/�}N�t�Q �B^�QGw��`��Qu�S��	���(IrUYc��1�+a�.�����V�d�K7�:� -h��{�κ�/O�r�b*hι�	wSf�j�Lcd�[ZW<E�S�}C������	)���ʒ��=�Z�������$ �ˡ��c��_c�(����X���F���̪ ��A}��ɹVΡ�^�C�l~:GPqN[�t�>!��5�0�ӓ�t7h�e�� <ro���"$P�J,��
��C��0�/�B�k�.��r��|�l�\���TZ�a��������;�	���C�Bs���[�γ��5>���Y�"3��"5OŬ����hげww'B@O*H��G� �����w ��{UtKD��0D?�D)	"1k�H��M�h�z���7x/od~�쥬e�,\V2J�����h��6�o-1���>���Υw�jG��b�PH�*�0�x.��%%Ls��?�b��l��'0B�)8#
���7(� �W�����Xh�[����l�7�:e��Pw�� �CY�:>�g�c�k�&��ϋ��WU�)-  ��D[��Z�9�/���T�6=A��Ǿ�Gu�T
_L�\�F�<+J��5h�ľ��w�L*��>��װl=�ϗY��D��'��E�4*��ш|7�YT��Z�z�	��AF��C����ϖ��R�i��,���}��۽<�.�"�Q�G�9��!�`r��ѿ����S��<A(G2���ի���Yy���~� _�4�R���C��O1�~?c)�k6;FdC��*jw����$�E����Z�ztn��Ԩ��u��𸝏Qܖ����mvy}�{��}�ׂz��=���M��k��W����t�8n�'��X#I�+�`����pw�u�m�%Ϫ���ԤE�Kml�J^�>>�`Ds��eg����m`�}N����J��29C|�"�Р8��(���#Ţ��/9���qT�ﲲX�?��L�5�X)� {��@���p���u���iKaLT����k�� �� pn��^�]�95p�t5���*�̈́�i�d�I��ѴK��HA�#g5ΰ���jN�7Uh�qz�\��|�)2���R��E���{���&�k��1H`���0���|1xWP�;~��1��cX��}�2�րD<�B�C�k���<|Mdok��].����
����:�aS�	z�D��0R1�؄�Ͳ*ˏ�y�{��}����R�<���%�"�xj���	vF<z�&���\@�� ��eN��Vf�P��-ߥ_�,�"��>K�-��"�
7�l�A�i��7�D�D@��
��I�!�H�č0���j�� W���%12��q/66�x{!:�]�d��4J1&dH��v����1�[����DG[v�M2]9��w��H��a�Y9j�Yc4���tӮQ0�+}�j�޳C ��cc�>b�;�#����(4�Tmd�+HG��rؖ_bzB��ڝ| �9�e"��Φx�� ���:M�A���&�	}<�l� 3ռ=��`��D��t׫'�cX�i�����&�����_��DX�*,�{7庼���i%P�o�_�,�����U��V.\�xsk��[�5�} ���+��_��3-�'�.,�+��$�����~�	t��'�C�6o��Y��2E5j8���������Չm�B�n�ΰ�[��iC���� �䍛�y�K�]�9�����z�I��}8-)���5��C�1�������k�9e:�0�͜��xg�m�(^ph�x���]������۹��	:k�a�im+�`�Ƞ���ѺǑ��<�"���E���u���cW7�3
*5Bx�ȥ�m�Mg%��O���Gc��%�¤��0:o4[��0���Շ�&k�����t iã�/�ֲ��<�]�l❺���nΒ&sHn�9���>��{%��{�K���5�#�$�_��r�N��g�zl�.2�#��[J�,&�w�Ag�S߽(�v�#���h��Q�)op�����u��[�v��H����/�c³'��FW��)��f�.�� 
���- �d�U0���&���f��z�𨬜h^sQa}�3��e���A��d dK�ǅ2��o��چ�X�_�fw�}T`�1e,�!*��	�P=�����|���%�c���_�j0E�����<!�
�=���қ�[Ea����!QX���OD�����A:��E��j�f�B�4|�5�7�T2L"zF��`OC�y���u�$���`�HFU4�́R������� ��(���3��g�8�z.��	�T!"��sW�@<��V�N����e�P�c,�D45�bq>�3�^3�9�H&���r���T'5_�����1^���B�Y� ���V�Lۚ�2�U8�Cm���͸�vC(|P±��BJejp a�F����N#����H5$�(�+3ӑ9���Q�Ga���4��9�ՆP0��'eA�kJ@x�E0�,����MM3Z1(���5S9�h�����Yѽj7кM�m�N2���aJ5��´)6|��tb��
�b% ��l<g&G�|8�,Odi��*hݦ{�3�N��	���Bs�Iǹ�y�Ǡ��fc�$����	@��
h2 ��۵��!T&��M9�N�ǈ]*@�n�Ҥ��iV3�.�AG�㥃�հ�@/�}u�:���Cdt�V�9��,�{w%H�� 8d��S�"�w(b���9��2����hs9M�y ����r|��[�G�Y�v/���V[[�3�����O^�����N��`��p��_)��"2���T*���<;�i���?"r
}v�:~��<�v��j��1'iڶ0�� ��~����F�YX*��ҡ��C,Byr��d��e�������S����}�A���z��t)��Ic���S��|�Æ8x���imQ��rH��߬���\ߪ�N�K-�4N���]�)��&���an/��aDN*-0���AB/�
߼��ݥ�iPV�*-�t�=��.���P�ѝ�x5`6��Qg|U 8蓙|!�н��ΊU��/�8��y[�Z��J��FJ"�y�=y�����%P9`R� ���0�vnJ"7��^�dE�1:�F]9�%��kCn���w!,�f�hX27��zҥTd]@�����*�ݪ~�b���J^8��*��>���W����%���y�CZn]Qoݚ$E�{���>��i�ߠ�K��m��/��ǲ�N�FXS���;�[�����s�8�r_�9���ܫ@��]�V��xd	/�V�S=�����}���C�r0�QΆΞ����ܓk�'"�,ʚ���Ķ��z�C�6GG��NJYMs��Y�.���c��a.��D�<�dZ�7g��ݳ�j�_0�g��?rQObvxVF���.��QR,ȀC�u�#�b��t&S�b�����j0c�6�\��K��S?x�T���*rQ�>9(���u$�Ʋn���$�KL��jd�)���L��ю���u͑�ϵz,�<<��p�_��ʓ�h��ʈ44�6b!w��R. ��ګ0?ъ��E�a�o�0�6�s�����=ҵ���F�5�E�"�MǽN�8Bs�8\>������Vcs%� �����5�̊�qj�#��;䶴�{�܍پ}3 餔��E��R Y"U.��}R����ޥ;Tk��a�:B��/䂒���PC�[����l�7�~�� `�koF�5W���*ٰ�T��s7(*����}�r�'Z�w�Qq&���3�p�RM�|��Ihz�����f�6��tT�����!3��
���V�OB���t���Ͻ{x�%�tb���)�����1��n�F��0�'���Nb`I�4���U�u���&ϱ~]@��L���ƴ����h����'�E�g��-�]�|*�oN%�h���*
�I6�Z�1�@�;j�	�!˟�ɓ��� 
M��ѽMbw>�K�93&mԱ��	��:��c�N,I��=@;��O�����	lSjX-���D����a$�-��k0ҏO�NM�&NRj�i���w���=�
Č
=ե?~?O&>n���?߄\#Cҩ�K�b+��h�X�0���>6���ƫ�#j;�`�5�����M��:ق�%	��+S�|J.@x4ߗCq����c����'�5>
s7�����l{u�-���w8�D�_�XsY7̂J��yՐ�U��?�=��v�nqA4B�ے�>��� ��
��7��W�%��*C������4�X�F��{W����2��F&�m1����mX��FY���/�F+�ѧn��
�*�L����T��v�T%��#�f_1}��k�y{�d���ț��A�Y1��3Lδ�� 8Bp,�4��4D|��[ò�|��1�<޴F �_��	����3�x~���_Ek��z$�r���&٘��%u�@qG����Ks���Ť�I?+�'\���A0�*��U� �yț��^����琣?������-?�h��eQ^��@�;��7�}��5��������:�@⃀���A*���/���&{K�;n	eb��k�t
�9�����F���`/9��Z1����3%�+_����I����Pb3 �$Uz�>�gQ^p?�>ջ�&���725�Gt���\&�RU�`w@��&����_�GigC��ܭu"���y��5�Ө���s�|���h���C�ވ�{ �|��\ωݑ��{��鄷�H�
�&&L��B�m����y��X�X?�[S ��f��IrU��_��)�3�����X��~��r$4D�~����YW_�-�ʹU
'5QD���b]aΉރi�@�E�rU�]����8NA�u�!ͯA���d�y��3�Xc� ��� 4�.���4�Rrx�����j���yzʷ��!��@��x���4����)�<�z	�ȓH�}�p�P�ι��u"-s¡��T:�a�U6iP��W;�K`�j���\�����@Ӝo�%��� ��Y;�2ל=�i��]@>��֪����<�yO��h�"���/��[־�1H���Z��:H��|�cu�$͔�uS��dcz�P��Qny׋�rg��f�(��k.�BӬ�@2t&{�#��o��F`�<�������S��d����Z�Ŭ��↭N���A�н��^�nO��6�[��8<��8������9�O�Sk�g�7?���87C(0D�� �"���R�{}��5��P��V2w�B�rKmcSW?�7wâב�&=ݩ[/A��֢~�w�Ƞ�j�I;zi����6t?�̚ZG�QiV�sRΠ����T_����������7%;;:?'C���wٺn��_�$�-d�悠c�٣&��><(0�ƛ,�v�_p$�4�=.�/�v(����0Cl�$�"���U�i�[��4ASò��]�F�A��o��u�U毡���;-/~�˅����_4n@���Є��q���A�M#�熈1B҄g����nh(ؽ�~AA�r��Ug�g��kxz׫����B,��y�����%��$+�3M�%�6�Y�,�J�;ֶ �& W8S���i��'���׷�SEMH�y��e�X��t�T�lIA(�N�<g����k�����6���C�Ɉֆ�`QV�@8��bj�a𛷵d��.��>}�0$���1Z�꓅�|7�"g���CW�+�0�x��<��'��X�3��,>n�J���YǑA�%4��*1�%�"�F�+�-� ����]�&"�M��^��,;Bc�V:���Kp@�D��R�jn6�0s ^𼿂"4ۻ��'�|��G�H[$t��yY��ͦ��k���U�Ae)�������	(�n������Lr!������h�I�2u��� �y
�q��վ��)�mge{���8����_��I%g�t�Acm@o�'I��������v�ҹdh���Ec2�jU�G�fjJD���0�mhS�{��d���<�g�P���_��x��I(���L"����Fl�a*G���˛RŹ�D���1V��_(+��8(��p�4�>��kC� i3L��m(���2�>	=m�rt��j���ᯓ;��UqdV;#U�&#W55��t2��?�M�C$V��ч��ң�j$�HX�M��v?$��k%�2o�	K�~St�z��)�����-�Wjƶ���	�!��b��+*��*���̀����r ��};�w�w1�#���
G;�* a�/Q4��|���1�GZ38q�e��J;�'b1�U�3`ؽ2�$ (�7���<����2�I�!���6�������.֑�Ơ��b��D�+�v�s�ّ˵T���4���5���~��1�0�c��''ċ�+�U���!���!�b�	q$)Z�f�چ�2�������&g�z
�Qݽ�[�q����d�<Z�K��l��?�.h!�S7��i){7oS�l�aO>���0��w��%�w�䥕>8��n׌|�ֿQ��o��Y�������QNۖg[b�[#��C"�����S�$m>����<1[�������=I��݆u�WP18�-�㩝'ѱ�;�>>�9�~�Ə�?���c,�m�c�fOc�e��nq40�%h��R��0<�3=������l���n!"� Ȋ���䭵n$%Z�����~�' w�Ji>����ǢϻO�.�6\���v0	$U@�i�E�Iv#��0ԕ���� ��xr ?�P��0(rK��X�!j¨��SFص;�P����7M&P֍�7�P�l� �X���޴c"e9��
.�VnVS�F|<�JW�RB����B��9p����e�y1��,���b�wsj�U��5y�՘��;�R
62&0��W����n>�.���n�v�&� ���� )��x�¥�?2	�)"�U|�S�A����1��ш���*�k�v,L�?+u��݊�S�Q .�1X��O�z�Z�#�fڛɄ������V�҇������_.9������=����+L�2���ł�Cx�I�J�Tc�-)���%�Kg�ú7A�[%�����'߃c��O�8���+g[��̡�w��;�)�~��
d1��>AJ��'�D�9�m� �����$8=�v��ز 4�.k�i�[/���R�*�T�8�=���s�%���4���\=�>dvM��UB_�t���C��(B�����h�W#�\�IqWx4\�w��q�X�H.r���qc��_,���+gi'�<�{�t&�͵	S���C��=%,߈��/���҅+�|[-5�v��[�H��%��,BMK�z�����W��+���W�������~
���%��rP�8?�a�p��+An��I��)��ʹhR��"<z�̬�ֹX���}���;ԩ/�)>�g�}SW�����M�U�CA���Y�R�5�P�B��*"t��3;����[&��e��ɂ28���L-���53���q�7Z��qg4�u\��G�~apkxaM�(�Hym�^`,����)����7?�����2�,�]ǉ��� ���Hj��6������J^�Mm��ϑ��&�z�j�=D]��6�O���c55�:�aϷ6Y%��r%fx�o�$?�&W��b��s�}0Pq��S��覿�������k��/;-AB�P8�/�~X�P�̪��`P���zK�O����A���Ǒ��h�8�����꘻Haic>��)3dr3��=.Ţ���O'�7͋��9�;�3�cs�m���1��ȴ��i��CI��z�b�4��ęw4�617��-�0=�|M8C��	�
0.�����7Y�sTخ�XYR�y�d��P�/�g9��x^��x�z�x��}��;�1PV��G�gj ��V�Ԑ����8/�d�:�Y|}k���X�:r�X�g�[�w���T0Q�,D9�G�����&�ذʣT�8oU�^���i��L^,a�6��8b*��gU�摕��6���*ImO��t��[�BGQ��C�g����s�T��J��_�Q�
��tV�:>�	��do�nJT1��+����w�@�36C�l�k�lQF�Ns�э����r���	?x)Q�¼�m�-<��
����I�Ƅd����O;��9���)#f���B U�g�+�}�[���Iٗ��^�UgP
,b�%Vz�f����f�[���UG���l��Gܞ��)�8��;�W���N ��<qZ��?��V�p m�ѭ�49_��ʶ�w <��69��Q��U��������_��g=Vby`~���pUZ,���r��z3�U��=�=~*�p�MN2+�f���u��b�����h��m�k&��~�u���s�YR=��4�A�x�;�Z��LQ���(�^��/	v4D�Ks��пNkw�L�F��v����u�H�~�&�/Y��]ղ��dI�U!?��g�2�|�[�i+��orF�/���Y2��4pK�y`���5�����NƲt�3�(o�54����(��l��_ZkH��5�"Ǯ�����?m�r�pAXu�R�e�.��SRs�h�.i��
�ù6���S����`���$4�c�o`<%��yyC���C��w-�|�X2�/(6V���A�%�m�ܾ���\�+a�{S�m�Xp(uB�Q�Dִ�<h�`^uco%ۑ��A&�����X�Cng�Ѯ�Lt7�Y�=9�lo�U��!���D]T����:�ۋPJ�\�w�չ�E���.j��~9,��D�`-ˑ���a�� ��qƶ�ݤ�?6�T���n�o5g��I��Ԙ�g1��g�WՏ>�$�=Å��E�-�[�؝���kZ���:� ۥ��9d�Rq1e�x���zB��d�hc�t��b&�-s2�rK�c��bXO�ۀf�k���ob�����H)���ĄH��!f��o�@;��4�cÃ
>���p�(��r��Pʷx5@�T>��i��]�-s�껴Hr����>|$����5�c�&�~�f���BDh�C�N�Q��9x��+Ѳ_��'�
��ϙ�}�N�Ʀj��]mp�#s�U��ARg|!�|̉2�OU�f�2��o��"wT2��{�
[.hc'|p�2�c=��@�t���J&�׀�N�a�~/ъ���,��8�X6��m�Wy����h�6��]��+��/݃~m<,?�A	�t��XXQe
��Pe}h�#ı�)�b�.(W�_�,��{���!  �N�F�e��O8��)�--,KN{ںJ��p�e6�,Hir`�T�G4���dB�z�����O���t���	bD��`�!6N�b51t�P�n�������c�EsLtЙ_�whs����V�$J���pM���"�[�aW�B�g�M�>���.�CF��5�?�睗;!��=_fВ1�� 
;��0-Hy��`l��~|�FW�xY�=\�������7���wa�$�0�C�*��6�~�|*,;u��in�{�U3G2nL����<N�H�!q�!̯�2�/�mխhx�6N�T��R�2=�v7.���+�okһ�K�^{v:�V��2gp*����qD4����%�����50� �{\���U�F��P-pJ���n�ǀ�[�������X�e��/���/h~�0���LӪ�x:�`I4�m%�	ӌV~�Wl��vC�7EN�:��~�¡��Y[5#�۔�b4B�����:��I5짲�xh:٣��{���o���F�s�1�{���-S��o*�����[M��Z:�T�K}�4��г�Ym#��*�L��nH��N�O����c��g�!RA��&��f�U6m�l����Q ����4N�V�HH�J蜈����Dete������zx�*�����{���A����%�8��!���(��#��t�m! ���饁�<�X� ����Q�yP۠.�` ���첲|$O�^נF�ׯ'/�t�%�k]�2M���[�fM�գ�c(%��I�?$1%�����*��jiҨq��La|�q��_Yj�`�IX��5� ����_��ӯ�I7�M x�ωK����z�W�.�8ѴzO�l����'t��á�ɦ���6�L��c���;'��>s���r��<+u�Wp $zf���l��~�iE�V�����TT���^����Y��6�F����v���,j�!T_�}��, 
V48]���^
hҊ�%��z�Ds�탩B�_�v�g�$3U9]��
�[�ϰ��2t�;��ed�zz�'Ôw>�"�{AY��:�q{�.h��q~�pn�۳{?u0�7�,>�I�`�L�ױQ�+���/���NB�ţ6�s�(�M�����cA��1ag$$�'�T��b�S���l̃�P��>S��L���a�;����C�n�!è��"�QF����I���Ζ_5;��eDߟ��8��s�p�qE��X^�8GZvb��Hb+A1Φ�ǜ��_��YWl�B(�gz� So�ل۝_�:�O������9�jK�Ѿx��71C��(>^�H/06�ς6ݑ�������Y@����0��a�a�V?`M��6~/��?���n�=~��
R]���X7����6ߘW��db��gѹ�/�1�{������W=^J�����u~�cr�X%��e�����uV��N8Y�F%���jk0	�1�˽BKN� ��X;��(+Fe�.k�;�h�&�� Xk��X���@1��o_�2v):��>�S��-���j���kX+)4�j��"nD�x��	"z�_6d���G��箢�w��%
X$y��w���O�g��zf���3�qq��j��8K��@y(�W~Q�A�f�r��/t>XW-"በ*:fG��9���pߎVw�Հ��O��s��\�ڳ~q����Z侅z�oË5�3�j�-��]���m��Xc��=��>	[�R����Sz����;�mM����j���s����h�d9t����^��W�Y���pz#��tHZ�RLO���;N�2C�=�`/A4���ɵ��� ��Vwt�ծ�}�={"��ɖ��	5z#�o�:@��GA���ʹ}��R��z��n�15��'p��B_9[�w?�4�E���Y�m�B�~�j��=�[
�JC����&�$<��)�LH���B�T�3�~�*������ְJ���t~`���O��'��"�rĈZ9�P�O��A�|(�_߲jv��z�w=`�(&8t �`�*w�1�[~އQC�kA���B���m�+��ČQ�k�`8h�"7�f�w�{7��~3!���ߗ���(���'�5�;Q"YkL�����٫D'!��z��#Y�yé��F����\��*	�������`�/o[5`<��Y	�pq��6z�>#��vL�����0CMv��لQoG���o�mP���X^b$ߑH�i0Gٻ<��.y\��pm���Af�y�Eo���݃�Ӣ��`�����U�Hj���f%UBXI>�����P����AJRo��bʚFq��ڞn�~%���Ґ��Ǻ��K�M��8���7{	8>j.��m@m�/C"h��Օ3N���y�=[bGx��s �]v��E����c%�L�B�����2�Zi���^��}Lе�b ލ�����.Kv%o"1lv��o��x+-p��`lJ�o{���)k��y���� 	��!���w�V6��@ZX#Co\��sG���-�:�e��>k��1��8��2��w����^ts���rC0\��2�R���yAJ�<y���990��`�ۥ�䁬�j�W�E+J�zt��貯4/B�$oI4qt	�f�J�ZШ�	���C�/��FW�%��gkty�9��VNuJ���vʕz�|{+���`ET�O��X�o�R6?~��Y���3A��
��W7���t���������|�i��R/|����~�ד�X� �)�J�V��;�Ͳ"�D��ܞ�4�l��D��:m:����/a��?F�UWgC�Yg�eѰ�t����Jr�@ԝ) ����LX�k,Sѯ>�w_��:d��ziY��N�+���a�dn�9Xi�g*h������"��r�M龐�y�e`�IA\hST}��6��Zn�3�y���9 ٧}��\�fӏ�#0�a�`+Ғ��w��u��2<T��\��E�Z?DE��Vz,�k�]z�w^�R��7H ��:ޙ���S6-X6��T��j4�z��ȣ}Ro!L2@�O'�N��N�1>ΌMP��TЪ<�W�[�y���X��4�o>麁��u�|T`6l5��)N�)�*��&�*9�ʞ�w�e�v�=Ls���-I��b���P9NE�2�#(���P��y��F���5���z7�V��Ny��K	���uUB��;��,q�E���;C:W*'8Q���~��}���.�RKh�A�m�1�
��^� ��b��~�>5	���c�)��ᱫh�����#N#�����C�	2�� ����e���>-C=�����]xc�9�2�s���ӸShl�Vf�d^��*ϧ"���>%��5�|��IjcST=Ο�����1s�nM���3���h��m���~�P��|4���R��	��{y,�w�՘EPC���H���i#r��D��8��%��/�!2���{�``!���X�u#��E(Q����b1�T�w���B����l�*�������u�����p���j��$/�j1�-|�\=�����"����/�z��Ӊ��	m��0�ٖ������V�Z�>�}��a�ڄk�F���띵�J2�� i����a0cY��e�W5>�\O��Y�(���8 m��؎����ԅY����_õ�g�>e)����˙�}aڰ�v���s�z��i�c�?t�q^e>"��-�st��ukCW1����P������b����P<��OM{��K�G�qo[sN�C��Q���ӅZrnA?�5��1�^LŔ�����t�5�����У I>�	W���,٬_�+��+#�%��nԐ�B�?�����%�5��I��~����5zP�&�9��>�|G����x���ʁ������~keA.�����NM����y1e7���u��
O����c(������b�����J�Qa�Q���<�9�UF�ۢ�b>�'��hu{��kU5���s�%F�\=�~+S��w�9u���1����2>�'�7;�� ���%*���d���!��cc�g��BF��{����%��6! ��B�zl	躆!xy�~Z����Mϑ@���wP��g�5�eՌdb�)��;A��e3��^��	�=�9�O����UOP�{F�83�i�#Y�����3ٰI��\��n�&���P�NH�c��{+��|�iQ���}�q��V�I<�N/�b<j�_�^QuNz��bR�[��42�{�bJB�]����F�?�$���@�ʼλo�D��a��}�'����{��k2X��z���̇���d�������&��:��/.����̒��IEE�����i^ۂ&s��d�c(�wq�=S�N��#Q�Sd��MNK:��z+�JZ�j:���fM�%��ʢ[\��:^6Fv�������f�DjX��F-�';$p��3�2Pe�6�rيtc-{��K���m��_C�A��{��U��;�_xϲܸS����?-9�����.��	Q��� d7~{�����re(�-�b����sº]��}0`zٖͲ�g��)�ͬ��g�KTa�Ώ���Q�pX�- �OL�Y���"q�Ѿ�4�)1I���AP�n
^�CP��*醹h_&l,֐,p5/�Q4�Bsv�-1�x��Ĳ(ּ�0s�d�\��AK'Y�ވ,7B�O�0���#��i_�=�5tx�lX2	Q�a*�B 5ѯ!%�y�X�Qt$I�I��.��{����S��	�=�D[�$N�p|l��`N�ǝg�iQ���(f�3�4-�YB-�xט
���.��q�O%���� �@PŘ�z�$L(�l\Ŋ��Ŷ;<��i�5u�c�a���;~�`��QKWJ:Zߡ0?ΰO?�玭=@�|~���u�8�/I�ʏ� w�mrIА� ��1��&�������u����@�>��j��r
OK���B6Ӣ2S�٤	(����m��e�{�(X��[�'�_j�0v�P��>C*�Q��BhG�LO�:A#�2n�c��hP�H=e����$l�r/������xE�пc9����"�zC����@G�K�w0�J�/L�\���Ցm2��K��X�H�D~���׫rg�K�q��I��_#lJ���`�:�M���k�C�]����.%8 �.\4���3��#w�
�9]ۓGV�\>�R&�H��p1J��T���'׏S�NJq��.�L��o��^d_O�g-����UD�OJ7zY�f�	m�þ��od�����0����DV��~yqHC�q#��������cЅG���݋4X�.֪S˼���`���?�5��|X?x�}gG�����%���Y���E&E��m���!]���F����)bN�R'|���R���p���)W��ǭ*���p�R���sX����yəiF0�A@�#UO��r��.����qڤ�b�᭖Z�oP�q&�ҽ��<�K1�eZ�.��.��7!f�Rt��1� HMX���q���z�8$��O7��X�(�@�<fw3�C툫?uu~2͜\a�F8�Ý�VF�t��P��h_'ղ��[�!7���,!gT��$EpR)� ����~������S��w�!�"(?�X@��t����kB�|N��%��G
*C���!�=i�V8H����Ҝw����[ҫ�jw~4a��Jǂ��-:���av��v|�`�Ó^�X�$��\�e��~����n����7��V�	�]�u��V��)&n��J����,��̦��`��A�	~�2	l���'�{?��@X�u�0(k�N��ƾj��Ϲ�Bei�o����Y��^`�u�V ��S���){�#��D\���lC�ѝ�Ù�	I�z۶�҅�|TNC
J��>Щ@M)��d�� ~��i���'�x�~�[�#���=M@�R~��CxU��,C`�|��D��mX�G�c�fO�7��9�!�sk�LC�!�j\��A�"\�\��ej-Wi���7D�~�FeZ�F!!��w��=� N4��"?~h��1#X�7d�`���s&��oS<��?+���%0�\�ҝ�X����.$�1	}v�7B�HQ������NK�oF�X�*[�zx?e7�%��8V��o�,BZ��}���o���qmPf�����]?��_g@vO;�UZc�-<T���ȑ��<�e�KH�3˛��L�*Z4��;�E�'hԼQ&x�K�c�S%����s���P�����?�M��)��x�lc-��'LY���Z����� Yl�&��'����C7�tz�=+>v_%�_}��s뿙^��u�K���'�����Q��t�S,�(+����3	�/A0�9}�j�w� `�r�?����Nr탋%�0Lm�Z���ċ��6Ma0w!I�"���x�eэp��6�۔tԧt� =�i�.�w��]`3^K)�P#����s�#�Ca���Z�"(��In�5w��D��	�P]]�0D'�S7d�+2��L�+�~�~����mےx���լ�g:�ш��1�:���m'HO����
��dq͂������?��� �E���p��n�ו���M��"��؜��^�������^�4鉾z<a6�9����78CaQ7]���}��N�_���`fc�� �f�*���D�rd�W/ z���v����@����*p��,�9b�2~��Nà���.��g��V������G����LA������f�*K�,�*��2$�3ҏ^c
Uq�,vJ؇�Z{������M�׀���]�1v���f��������<�B�&��e����R/˔tؽ�˽��g�-^Ֆ�$��G��3Uh=���mL۽����`V�ܕ�>o0���U[pX�|�B)���a{s�.���˸�+�{����m��V�V���_�-������T���tH�P�@�Xߔ�hO��-�UDJG�!}��/4�fz����]s��h/0ƛ�3*��I�b�Ɲ��F�B'���~QF{Zvp��䟦��R�K�:� �)w�l�A3W�t����w�*��P�ʨ��Y˾�u�X�x��xb�V��ZCd��� y&D/ ���1c ]�
O�.%��p��96'74G����5PRA����g�	�s���9��$�,2���m�~��S�����m����~MQ:_�^�_�tqZ����Z�")�\Ģ@tӅş
>�b����i�v@9Z�kG��%*���=߲ʐ;�g��m�,/ا���7�
X�ѐ�p���Gܘ���K�,�9����n�!�2҄���>�"4w���[�3c��g^��57�6PR�}��6�7�҉��S>�οg�ilu���/=���G�oȚ2�"V쭮%��M����K�V��\����p������+���6����=
�,`�K#���1�bԗ� d���%H��pj]Y��G��t8V&L�zb�_�پ��q<��ށe��ݯ�u�\Ջ)�Ȯat���n��	POQ��'3� ��|^�7��+KXFEu�Ʊ���DHo�)4��D��k�2���3R��z�r��]�6��vn-G�Vf41e�}C��L��w�hg&�_�g�rQH�	L�7��H$�WV������6A��Zm����տ̧,30m��Ĝ�FM�-;�%�0#�M��P�Hf�X����=�0�ƴi�����;M���[Q��y����D��ˋ[v��WU��?ҵ���G���9�f�����<9�c�����RL9Y��S�ʸ��r��vֈ��r�]Y( \��d�|?H9�"��caB���|��u��QͿ���+�2'� ^��r3 aF^@��E~�M�}$�p���C֢y0!���K���N?��uwѢA�0�Wf�FM�e��
t����u�����|�&�FKm�Ҧ=�_�;�\ 
>!���ӂ�/��V����~�y}����?�j���b�u�U�ʹ�c��2�A��Y@N)�dc�G�_?]\�G��>?���+�4����S�iyR`��5ƭ>f����s0��!��L�φe��V�I?#�*�$����cV�t|�[�ƹW�z���8P��'{)��p?+�h��Ki^�(��!v��O�����'�8�:��H���;�"@���e�0�9��aqKl��u@k����MY�خ+Дj�~:;�G�R��#��Q�b��:���	8���͡\A���f��q���z��% o �<��<5�.�w��J��>�G�oh��F�kq���K�����Z��44���%��E�g:u�gsN��M��'�t`[x��t�6�Ci���<�/v�s� `M��߅z(�]@�e=#����I-��S�ieE�|���\;���(K>R�Y0T�6��욠)�s&+�3C��pV�H*�m�� �c�\
���l�Bx;7�5^��>��i�`Zv����m���QŬ��X����fUd�d~9����$�!�v?�&�o��R-2q��9�&:�`L�D�朁0��k�vc��Z8NĞ�)B�udF�ew�Ų�{�<�m��ۖ�j���D�1�YEM@G -�`��d��0H�w-"�Ʃ����I|�W��_����W���0�F���^h�����Y-?R����6Ks�!�W��[�f�2���Z<�~�A�l�ƥ�[g�l�V�e,�'��̠���2�~X�L��Xo�8��S�h۽S���ˢG1+�t�\����6�kٛN��'���%�lq3r��S�B�;X%��#�M���h�*e�`�a���筇��#TW�. aV5��Q{�##�}���btv�)�Ed�#����z�p�򍅣x�	�zv.���T0:~�P*ސ���@�ڙL:%�&�loF���[�r?����-9 �f��D�`&��0:1Sr_I\���Ĕ������oZ���J�M��YN�h+3��D/��;�-Gr	�U8���!"8�U�\4m��?�i8�2����|G�f�?F����#ˍ�gэU&�`�3�����1^�gh� >�m���]4��[��1�E2Fs���E�˄KvĐ���0�	Eq_4>��_��^^/0�i��eϟa�_.x���f�N�	)��1IGT����z(�;��t4��6B�1� 
w��F���g�R�,������~�>"�?64�����	/cos"E��K��RY��K����ޫ���i'�@v�)�� �tQ��ы��zf[�t$�H}�X���3�� 9߈'O�Z�ִ���8��'
��y4#<9hVn��
61\��#�g�h��6��s0��� ���1�?��K�����3mV�9�xgZ���Bm�����#Mw�$e"�����᝔-��_ty��T��|]�&��GՃ�J��1��("�^�(�J06�|�R���NJ"\ ��,�ޙ0W��AI�A���9�?���El�
��,NO�0����H̸��V��>�m��n��>���@9W��J�jE�x(7摏���U�R��!�<�vO��]��Q�;~ �~i!&��ӏ�*�h�v�XG;Ϭ{��t�G1��\&tF��]cNqx3��.�iI�g=1�5�۲�t����� >Z�x���Z�PF�|��rj?̮Fۂi��tҦ��i%jw�s���k��f�l�	ԝ�y�"vg�:%e�-d����n���C&uK��)�Ry�BlΕ��8#�g#���mRy{���.�z1v[!�C�lg9�G�S"�#s�^m�s�V�9^���v�E �����LM�w!�1s��d�5���Pş��x'|�]��O%�kޏp�O�,�$�(r6��K)���Do��K)#��!*�h�4�QrUЊ���	�"1�[����]#镈ym�	*��[!�|���=ˉ{�Ws�<	�����'E:۸��e�4{Ӄ�"�:�9ESo�����+��fc��i�oq���]*��<y�.w���K�>��Ժ���n/~���
|Q0�G[o�����?�D'��<Px�Aan���L
M@��*j@�rY˘е�.ou�pgP	��S�E���0��&#
�Rx��I6r��p;��)�R P�\�V��D\ȍ�_Kj-i7����w�jw�B�/�ܛe�#���TgD^��UM�����]�wݪs>h�u'����>n�g#W�r���U]�r�i3Q�P�<�u�:	���J��g���g�+郇)��"]�@Z� :��䇖�V-N'6`�;�rv���!H�/�(�PR9��vи�&)(���.c'�>���S�[I���� [Ѕ�X��MY��B�c=������;�N:6;x��(=��<'3�#��NY��EC8f�~�>���N��$�{kٙ��;Y���b�@a �Kd�p����:/hm۬g�H;Hʊ����`C����'���q���7G`���@r��P�������jd
!c�5�-�1���N<z��r�v�aƀ(|/>�ے�����Yo�WF��8�@��L�k�*��=SfX�/-�.�=L��_�/�[�_Ѱ2�Lm��	��ظE�Fє��'�M�eztzA���)}���&�%um��K�������]�S��]���}6Y�!�P�t�#��*%S������ޓ�����>����5�Q�(��Ě+~��A��s�J���'���릏��
� Je��#���їPҚ���9&x (�u���rL�o4Ĥ�P���c���N��Orca�q��/�3I�F�g/+w>jz�ϲ��@e�'� ba�a`���~b'g�]�U����+>����r���(��œ�XnV��:a����Ѵ���&8���X�DO��K�{���K)Cpp;&¡i�)N|�Є����J[�X��.�j�n	NLY�bC��}"�l`��T�6�eh�m�L[���}�9�Dӻ�D���4"�p̪��u���~F��{;h���S�r��a����n~��.�Jκ͢���m��F�(5���\]�L� ��		����X|E%��<��G�)_,U�;�F����b�g���3b��~h6�)�p�q�gca����i�XNg�}�@�x���XnU4�����U��c;�sz��>�/rig�F��+� ��"t��V�y�}���,:x�b�z�h�py˧J�;L�y�(Oe�l�?�B�T��٫{�I�Q���Va��tb�ۘ6}���/y��������F)�Տ����s��cJ��u� .Hd�h5m&z�{��;��2�]��Ø/Aš�dè��E��<���]�4d��9�sت���Yjj��� Y
j���+�2L������N_�@]��3^�W��?�����6x�:���E�+���x��;
�OlH���U�������ZaN ˚���MB�0�#_}��M�+��d�(]%��#���$�l����0���r9�LUQ���DD�:�4ae���K�/�ԉ�[g���1��=���@��:B	h׬�kN�#�����!��3���e"��������.�K�=��Ąm��!n��PR��ȭ��zpج9tA\~#�%���K4"h�߃���sGҜ���h[�y����մ�z�R�QL�V�y�!<&�+�c�i
���P�5J�M {����c8�C��;Zo-��Ρ�c�y	dZ�{���t~e�@�_�G�q{����Sn�"�G^��i��	���-�rj^���!w"N:�q]�@�>-r���Y����{�;`ʂB��Pwc�[��=�I�n�}�9�x�I�P�D�J��<�*rk(���& ��*���3��ЯCr��t��h��ڑ&]�6�A"T"� l��g�u��|_BAz"M��}�~�ū�ﳅ�� G\l���������=b�xRB8x��+��g6}wH���a�u��͸ٖ�ML&���YQOpoLYpK��.\�7A�l�
��5)��+F0˞�C��e�b.LYJ֞�"���/�����4�&��
����
���r3�L��d�r{�gF��:��+	+0����>�kG�/��;��e��w��X���i��&��h�̲�)gI����o+���J�WXx��e��6Y/���0�,��c�q��\a����q���7$����@�#��G�6#	t)���;��R'��Kԣ-�띄t���k%ǜ-@~�R5�ga�ND(���c!�Aķ����}�S�H&��)W�嚯�\Ւ8� ��<cP>W�Sy�M0�:Rq'���Wu��$?�M�bS��h^��Z3���Y�K�M��7h�hTe�Km���Y��s]հ�� &�C�ʮ�_q��7�8��*	rrS����t��w���62�U�.ƫ:�<�+/GR�c-ڮ7Ά�p�h��ž[G&�[�����7*����	���	�]mPv�.-�O���Ȉ��^�mJ�b`;��j2D���V�6�*ɽȟ�79<Oܚ��������J:ȕ�Y4U���oT������Ck���S�`�үfr`�현V,�%���G.�,*�߃��)����@'�ZO!��0��_�y�;j	�;�*`w�w�3،.��m��Y&�a���I =\�ل+�����D�`��o�U��Rz��;<���K�1zC�9a�42���@�0Q٠\��oϩ�?�n+�LW�6$��3��8�[��iɶ���t4
�Ƅs]p  7�܃�W�@��}s^؜
�G�>���P���C�3]i �c�y ��y]}����U����:�͵t�V�������$H��v��b|ǃ�_H+�=ūS�`���G�I�*�ؓ���S��Z��OZ��z�s�KL�����I�a�S��t��u�B3��I��T��60^m3(��}�ӌoѷ����<<�����8�@�>�C�ּO�I�3Ie�kJX�
[,�@� �-K>j�;�`��as��J偮&6�
���'d����1Ĵ�3;�=�x�M�-�+K�mqQo���o�����SIޯ�b�Nӎj,�J�5�� ���B{���z�u����{,~���:�r���J|&m��x�j���?�>W��~��e��,)���AV�:^}��J�zʑz�*~l�	"��w��>�H�-��N!Z+��ƗT�Q�
F@ۨq���^쟬�*�~k������UI*G���=u-��h��gj>�6�͕N�?�/���^����c��o�g��:��Y�d8r�*!Y��7����Q⭶����:���YL���\�0��w�!yW�G�4rY1�<���������dM7�oK=�%�[!"p��C�6�lPߣ;���%:uh��tv�9��Q�n�}��-�S�߷3�Jw-Tp��ԫ}BD���ʃ��Ͻ�w�T��p,(�A$|���m>�P��^�M$<u��߯�H�J��ǅ��'��*�S�ڐN��}c��)����	��(�I��U��J�lל��'6}o�BV�s�#2,���A-׭{K?eg��6�F,�|�}!��< ~� i�ی
�P<r~L����kﺭ���[r�,j��ץIVTȾ���l|!��Sdy�_�BRW���6_������{�u�BL���q���̞��5#jb�7��K��#�^TA�"��-
�XСg��ٍ�~&d�j侶V`��Qdp���tK�u�]����Tzc�6��4���E��7�{�MW�$���̻Q5�b����N2��ǻ�]�, �s��ߛ�R�<�*�C��0�3,�5%Ե�&����@�!�G�i��b��=���D!�3�ٖ�W[�����������c�S\":��#-N�k�^o
8�ho\o��"޿&SRblS�<�k8V��C攏�V��ş���RtīD�?�ь4n����7VM� [U��h� -�P����c]\�Z��?mT_� 7�&4�^JSeEM<7�u �1���g�
|Z���w��"�.����`��
�" F	`�1����>J��B��y� ����e�����*��\�JB��ԧ��f��N[�L���ۦ��U_�"3����_��vp��u��tو*�,��`1A�����~x��|�#"&�!���	P錭��k7��K�7hq���+�?=�njW�򷕑I>q!n�k���5�M\�dR��e��h�.vbƲ��&�QDe��_�D�tK�+|�����߂�-���kĭ���.&:��
e	�
�s���*�S�����;h��n�6��O��	�Čⴐz|/,>��GF�'���;��H�v�R�2�H�1G*��SH����>1�<��V����}|���J�o��JB 5��މ#�1q���>��N$)`�y�`,-oO2���E��|�?][����J�j_�A���ĳ.�n�_=��p�j�������j�-@h��H�n���҈��ķ ׍1;[��0�	��� P�s����^��e����#������S&�WV�GqӀ9l�O�k���������3[
���v�d���u��Lv��y��S.G����9�m^��>�P07��ϡm�N�%�Js%���P��zپG4��hf��Wc))�܄��@�`��
[K����a��!�m��$�,Ij+�U9t��[㏓X:pGO��E����G����Z@ʨ<�9(d�����3��.�}�bD��K�*ק�.νew��sυN�ݼ�ң伱A�bnG��&^�݄��x�J�29U-�TAfI>jՃ8�(̠���v}��:�<�u�B�������+����c���pt&����e�T�1*�}1Cq�F�b��Fg?��Kh��-&U��$�η�C����`��
�7	>�ܣ���&~jz�\1��!ӵ�Ϳ�	4�^�*�mG\��qKK x,�h�%�@�H֐��i�)ц]ƌH��@�WD���1�}��V0�<c����;�|d��z�=)e��Cڣ���浣K������þ�"r:�~�`ޔ�ehm �����c�oאN�|��;�Z	I�f���)#�6 5'c��O����\ffs!W����PC<�z7v3ހ�E�B�2�;����?*��0T4�ǽ"i�Y��>D~8R�x�bt�"�2��(z������8�C}���f
�&��Z��םՐJTh���ڡW�88i3���d�4� 2���;a��v�9ظ����+dZq� �k
���Tb ��Yھ�c0ʲ�3��A�k�Q]Kq���y���!�]��n�1��%��e?�kS�#�k)#~C�w:��8⪬��쐄�o���#(��!K�1�p�~�v���0�1�
�7�����6��û5X�w��x��#���Z�i�s���Ek���� Wyq �y��	���&7�"d�V��������8r5Q�au�>��ߜ�Mw�λRo�����\%;q&�Ӥ��e�8F��d ��E������Ŵ3�T�`�R o�0.�I ��0�U�G��F�Tf`W�:�Z��ߗ�D!�z`5�(�b,�*�ɋ[ֹ�'�<���[�&�{�u{v��q��x��L����/�ư8��o1gqdW�kw��^�A�>�>��1>�E�"�]�c;G�ڑVK9�Bly垚��is�+h�r{f��1b�DC��}�`�/L���<��J	ג�f�ڶ
�N�.�sC��
?�o7�ϻ���3�����5"8�k5X�ָ�����Ǔ���aO�b\��KFrX&�J�]Ϻt�=�<v��H��:P�߱�dE2��3�f�G3���;��h����S�?��x?��A�Z���`��v��l(����Ma�o�����x{@4;��@g\��i�5��Pŗq�~h~t/�j	����;4~�H�Q��ʖ^V���Dg*P��1���%a�^����{��kq�S�4�-ȗ<)���/��M1��a9�{��ɗCƐB��/ܾ��`�V��e��KW�⾧B1�\���������&aO!`��آ
ϖ%ӗ�`"�$��(�9�`���J��.��&�X�(��\=�� {	$4���Y�C����jg!h�.�&1T�0����-m+`i����S�K�8@�:Kthܔ�����4y�%�-]M���,���	�x7f��>2w�pcѼ~ � %��|&]s���(������S�"�0�'4�	nC��J�0 � �VmP`�/���o��
��V'U�_20,����d- ʴ!�o
AZ�H��}t�7z�-{�I@��ނ��4�Z�8̾�s|Ø
r�g��
y�i�V@%�x���P�~(�B4$��H@�ѯP�NZ���efX\۞���R��#�lz@�����	79�`a[����C��h�B�65�9�_�_<|���*5u�C�<�VJj���ן���t��� J7�gW��f�G]J0�Ue�rH����cJ���}G�s�+<�(��nl�C�5��xq�Ɔ,�z]( n+�z!s���[�&/�N��MUA>i��z(_Y��wa�$R��Tϸ�Oj�Q��&�8���pQ�ι�^��dR�朐.�E��2��%�W�S����������f����
3�7'�e��#�����H@0OQ{��f�]"^�9�3B�tn�HE�8��hj-0�7p�^^k��:=U�G7p�L$q��;h�*��y�!R�f-ץbͩZ�5���'Ɨe�v�u������߯<��f��9� c����`#���-�R<��p�)�_��,��&��ٜ��&�_c��6�4�,�\#l�����t��.h���N�+�� �
j����//?6+��OV���8�o����=SM�zխq��.i�o�$���%/��L.N@
��oG�����"|�sM?ňX�=����S٣Z*�hͿ���2��X��*ϿcC+[s��o�8�#����4�^<�ɶ"hKJ5��hQ1�E��-�rUhFݩd}��q����t��* ��P(���3�J��r|I�}�t�P��%Ӗ�[��sJ���\%hթĪ�}%4�y�R6�N{���2��9Y#!�ԓN��ǻ�
t�r�SR<�[��n�7*O1Mنg�(4�U*�p��Y[������K���̝��y7��A�A�K3'C4��2Z
`ލ�*����DI��Azߍ�\��_N0�7O)R���(������G�^K9�U��:�u%>�@�A)�'ԙ�:jR�/�������H܁@WA��2�c@��ŶD=%I�����f��X�@7���i�^�c���������B��5� }���7�qٿ�k�����Ə!O���n�����Qu���q�\J��٬��d�p�H\���ϐ�L��;ư�O^��~p�3f��:�J����ⲽ
�Ǭ�;��R+�c�Q�(|�Dңg6#�'�JQb���v�VZh8�u>Ѕ�a3Zh9�B��^�6H�:�έ��"�9�m-�&/�����o��Rjc~Ԁ��ޣ����ine������HE�8s,��c̔���A���@x��Ɓ_����5W� ���!<�Շ��~�yg�0�ϕpm?��p�G	�ݏ*��rLB�����<��c�m9�T�&N��t�_+��S��V�~>j�� "8'"*ag$صD�yu�;�E	��A�o�6G�����]�ۭ;��m~�5=�!I�W(��:���盉S��R8;q�>&{O}R�����c{dh7���h�gFCH� wɥ��\ὲ��$���0&��bʨ�����o���I�p6��)Uz��� ���Pw:��-��s��.��Y��/)�fiu�-&'@G!��,2�?�a�7�u�;��ʮ/ ,C�@�+Z��҇��fx�{s!tè�,��޸�}֫�`!{� Z�c�
����,w�M��1�ͽ^��ӽ3�;%�+ɷ�����
T,�S!�¬�F�<32�>(�^�k��ϰd��+5D�+迒̅d�_�)�8l	�Rk=1?}��#e���"���=�`��ρM��#�&��ؚ�V<�p`}��Q�d�7���ÜR�k8�p�6 k�ֻ��Vx����K����;g�55��0�5-�l~F0]��x+����x�BVA+��=�&(�Vm�Q�駭4�s2�t�o��˜���pu�|!M��[��ruO���uڤ�*�6���;*����w2�㺱	}=6e���.6	<+4�Z�4D��.5��z%���5��s���Y��I1f*��i�IͶ2�O���yՊ�o��|c� �'��E����L\��J{w�� F�}������8�Z��f5�Z���*Y}K	�_BI�fHXХkh�ոȝ�Jl��̱���x>�j.��'��칢�<,���
;yf����jW��v�����ܙ��i� �K~�	;S*> L�.��&tQT�V�THO��42�֍ʚ'�58/����Y�FkZ�&DF�qȏn��mr�g�����*A������Q��&I��?��6h�-���_���N�K-��/m��S^���2�aJi�&A�P�l�,<a18J��S�^*n2I����B��3q
���y��B�Myp����������+���/��tNd�I�9���|щƫ����Oa8��Do���<�G{��q���X$���'�����}��>�1WoP=e���-z1C���;�E��}�:������R�J�)��`��3�������H؁to���B��][�IL�N���̟N:v�G;���C?jX:d�%�3��|��kg��l^��[+�"��,ؠ��d/�if斠 P?��{��<��}�Z��`h����r����L'y,Qm���p�R�H��qա��w4G�O�`���Uo��]%���|���V/5��9:��Vq�;W�Rd���;�$r�,��	S%��]�lG�";ӄ��-��l�}oE���Q�ḍ���Cw��r*�J%8z.� ?b\�a�F���1��u����${�~�F-��dBq�s[�O������_�C�& ���A�}�M����*3�R ��O��aʛ�2si��r2ƹ��Tq�
f��Y���{]`�Ϸ ����
~�C�[.I�`gS�l��u���=>���C�ߪP�$<2ʐc�S�!4���D;vnWvȷX�}X]�f��x�W�m�7�$�u������c^at���� %y�}C ]��2 �׽�u�좋\��N����ߙrS��=�(z�]{�.�s͂'/�_H����;>�d�@�<'BJ�$U�7(U�0z	�}$*��ًC��f㤃)??FE`�Rsw�ȴ�U�H�p�(�Z�eb���Ů��ޝ"x����%]�O_r(�6���AΫ<+���� �>���ѿ;���,,F��� w�l���2&r%��#QN��Jj�Yc5��9�n�Mq�@0�/��U�
�r�
8�PQ4�	�N��d�
��8I���ဪ���K�U�tӰx�]������F�^C[+.u�u�_t���5f51*�`|��	 �pq�0m�S��ۓ�[;��TO�q*�K�(\��d��g���k|���J�r4����;\&�;�6�,�̷��D<� �-Dl�kYѫD�)"�R�!�&"ٍ�{���>͛�����I
�N,Іcab�16熶r��b����t��d����,vv\������ӊ�X{�ڽ�M���D,�˼F�(Q�
�<;��ٵpku�Ķ�Cw���K�d�cQ�����Wy|���szmO��\s�0��
-]��p9��W���e���65䲧��"�k����2��Q"���*��:�C�M�R��]�Ј	�{V�U�Eǭgd%3��P��\_lR�sxt�}�]�,iÄ3��Ys7(��փ�u8����*�B����&�J�9s��e3�s#^`�) �v� ��,`��t4&�ʶ^X��$�	��%ס8��c�-�a�H?�h�G�v��@�n`�˟<E�|�jS��$
~�o���u�G�-E(>YR �z�c)䂶.��w�݋s����hm)��k%S9B��.J�ױ7~���WOfHq<�Pj� �rBF�,��s��5�iJ�:m�x��^�n.�L;~۳1
�}��/uC��0%}�w��98OQ��K�R�����@�ɔ�Ā�e���#���t�,����}�E���Y�5#X���y��>y��y��&���;Ѷ��edS��:e���N�˾�c��c�G�)|*�p�r�# ��X5[��3E�U@u�ᮚp{�~����8�*x���M%�.�Y��5`)sP/kt�����1�~@^���o��KTo���\��Tw���ڋ��@��s��U�\�xX��b'i�#Cǀ]�}q��M�6¯���?S]�4��E4�w#�{6t�1�nF���Z�N�:��(�Ku�m�Ur��<�S a�p��!�\i�7�)�~3�Cz�U"�b�~��H�����bD,�z�$!S��®�C����\YW]�f��B�=cٯ6!NXqt�r.��	������"���N�)��󵧬�z;P�5�^�iF&s��xwJr�"��9[M�I�9��Ko�ZWW�c�
&ZW n�0W[63 HD����n��ړ�7�v��0?�b'�q���s�Bk�:;t�:u���5�8��
�0�h.3��r?��W�=n��`�;���N�0�̮�����[:��T�q��,��V���a@��Iή �b�vNxe�)$�Z����l��Ol�7�I�` \?D+%��T'���h�����Y$pjeo1���Y�7 7a�
�g��%o�X$�����B��������Jr�Č�=k~� �f@�uԷ�7�f/؏I=>�����=�b�$��Q5-��-�/c��k3��8�U���;���#a{�4y6Y$���}"�"�;��v�O���o�xEΕҞ�V¹[���	=(��IUq��]�Q0��������R�2�<$��a.��ϓr��V�$���Qc�Y�(�ibyM���(Ϡ�Ĳi���*�lk1�Yfa}� m�z#\-��蘬�7���`!��ř�.Z�0P���}[�x���Ɯp*���5Hn���lC7�O�9Vj����eF�X��ɩ���#xk��[�D��V1���sD�#�g�v��?���蘦ݒh��גp%4�V�d�B���U|�ɖ�+r��<:�\�"���
椓o�ҁǜA8B�r��ވ�NkN���~�K)�4�]Zi��u����I$6=���U�C�;-�L�q6I�:�&/��dܝ1��ӗ��/��qV*��!3ʈ�s�5тw}�%���^�-�K6otu)~6�PH�+�K #A��̫���<��� ���$N#9�Ԙ2��h6ϒ�p(���}��1R�|r�ؓl����(�{e�I��l����]��~�W���4O�5g"9� (�+�\��_4G󜥡�Ӄ��z�x�l0pfȒp��t{$�k��3�R�^�he����A����g+,���sZ��X�/6��!����r�I=,�&�Gҩ����6�O1�xa_Y�9�sQ<�J+8Ӿ�g,�d�RdZ,D�S$�}y+~ ��{aN0y��x2�����ex�2���ڭ�`**����(4)ӌ��ad��Y����%퉙�D����%��y���?5�5(��1��T� 5�e� ���V�%�`�?u݅�s����#��^�d�k�$7r�gR�Psfճ����67��?
�\�l�O!U��[�?�#�y�Sl;Q���s�T��9���<��)S�}��j�>�HO���Ķ�M�)/:N�gI��l�u��	M��ֵ�!�
5�,��{���*b��'�9��s�׽E����O�w~49qY@�L�N���/�)�F��	4L��ɍf�Z_�C��'�� �9\$�.L5D��KI|W��>�_T�*p��,R�>_��[�ɴ��>�?	����=@]�5g�TTZ� l�٠�å�3n0��Kx��p�!�Χ�'�1^K̢���8��E��|mbP�`_J,�з���� Z@Y�w3Do�:w<*�x�(�}��p���9#?�T������-;��%�Sv/�Uz�L�
lWGz'�Z�
��u�Z7�L�b��'�=��"�j!�	��[9i�6"���эṨ&Q�hl}h��)~�GhE ����7��L�3\������I�C�Ǹ���~=�4�{N�X���:�N����$4�{ZA�	D{��M�/�Qɏ�\���A�KHK'X�^yB�B���
��6
��X<��� �+�-xUK}%����o	�mB�������r�c��6:H��
�o"�X�����%��G6s�L-��C\�T��I�pф�GHu4�b9�N�f-��;!s�U���n��U�����9*;��j���<��Wd���?=]5;���Bc�b������炤��� �䎲?;X<b�p�`��
�ʄ��'\�x2�HVAuAX4'�,�nn��"Xug|��.�#���mH	.���J1d� �_�7y*g�Ú�UGP�!��2z��=��s�~!\>��p,��D��O^����T,n� ������5��z8�5'�����U	�nl���%��<q&@m��ȇ��?�#�@��O�Kܚz�'��>9 �6S���G�bՍVQ�߻$ʖ��ܣ~al��ѕjPb y��4;\�3�"�Z_�&��eP���<L
�!0�SAL�|�>>������![�kQ�ࡵ�,��q�$�4zɇ�$-�aGN뾸ބ J2Qf�D3JU]�;�1��#l�����-��nė�ap���������f�_;�44v�h�]�Q��/%1��_>`-.���bF97Y_XxQ��\���Ǿt�?�v�ʰ2�������x����.�5d�Xe:���O�O���h��������9T_��[�]������f �Ύ%6��y,d�� ʲU�ȴ������u�����ɴ���w�$ ��S;��	i/j� ;?w�3
|�P�?]�*��>��-_Gv��v������%�΢���yy2�`�� H�`�>	|�S�t��ݭȻ�Jt-��|&�����m�=�s��{6R_VL�a췚ng	������������D�o���rn��T��֕ 0��d��ߠ_� ����$(N*ȸ ?q>dw�Q�XB$~�^;e#E  �\��V�*R+*�ـTٛʂ��~���V>Kkbpۘ�*(t6@��"�U+����lZ>��%�2���z1ԛ�A>�k�!=���)���U.�$�u�"������~���?���dL���t�&d��!P%?%�����=T��]��mVi�لcc�����;�r���H��S��F�ԇ����� C���s����ZrV���Xk*]��D������ %нW��$��;u7X�6u����T���ٺK Sߔ��������Y��r�����Cv���
>Ef�q��6s��fI�+37gt��l<�@g��E�u��-i��K�	��Ff��<O� �4��a�ϊ,�5�K�ܰZ܃rDY=A|��cOR>vN�������@���H��1��9ؑX�$l�1�	��3�YY�W
 (F��znsFЎ�:D�Wu`@#��|?����ν}+k#��}O���b=���蹞������Z,%?���=�L]��3����`K0�p�A0��h��ߧ�{C�pb��p����n���@�ޣ��/�(Q1_
���[�L�6]# ՗0�^����(�B];�# f�]0K�K��P��,�oO�S��3�21�U����/~�'�=�7 ���c��GjʱCE���5u�����C����x�Dsg�ةp�a�Ν��{����,$��Xt����o\���gБw�^;�Tk���%)k��7LdNvt���9���a���,���k�v,s	m%;��b_f���(��C���S���	'#��?=��cB��cĦ6��,��>F���S��X��������
�Q�	�X�p�D�9.N�3}]� ������9����) u
���0�{���ypd�NK«Qod�ɣ�J]$��MvF� $�F4�1U[�c���������oS�}�@�L����(��p�D�7G=(M����@xL�?�8�^ޛ���B��kW�U���~���
S�%63��f
	�3�bA:��K��O��uJ��k��%xP~��b���@�N)�_6<.�������P��JGV�#�H�*��p(Sl[i�����1��F�bL�W��1����$`�jB�tT虑��7*���[�P�Q����N�PzNW�V:�.$�,��gX�d�Y�����[����X-�p�_:(_$�F:Eb� �0��g�8~�mm~1���;�����#)�g+�Qlgi)��6�om�^L�˩�r�������
����-T�xҥ�;�ǔ(ۙ�)��s�*�V�vV��OBOiX�F-�0\Y%��j˔J��k��;K�ۮ0�y �PG\���3	ya8��YQ��Ꜭ��S[7��)Y(��J0��&���
�\ �O��Uk�)����V��u�
�'g�y�H���;	r�[����݋�/a8���e�q��S�N�kw"�.��@��ZTo�-��Gr�~���RYi0�E'FD�99�K9�SK\땡HP��¾�ٌ�y�����RB��YL�V��:d��~32;�A����-���1C�qd�����_ǂ���#���'&�LIf��MW�h���ӓs͸�b�v��L�����Y��?b� \Ӝ1-w��4��S�.p�0�P��&�h�5��8-+� Wj�� � �J���P�ͽ�]}����*���*qy�;7�X=��C�j�ۡ��鼤y��J��p��o����]"`["=�aZ}��|�]nmT�O����8M�吪����m&�R�+�r�S�_�ϒ�1t��2a��2���V@ ����RM�[��Ը�@7q�8��z�
�=��t|N��W�%��"7´5ǱA{��G
�Ԣ�$�2`@84_�3MU�U��9�G+^HU�Ĺ\�@|�7\!r�(�r�~�:�z��3`�C���{��0�m�v�:s�;6���^b��0G3} �B��:���q�8�3�6�S���W�/R�c�*Z�� ��0w�����O�"�����,��v^��Q�I>twT/��
�5�R���fן��:����u�#۾h�U>��0I��u���`���f���`ӶZ�W�W��з{�3��&�����ծ^�P��o�)2��3Ť�������M혩��5e��B�$�p��B2{x2����2
X&�Z�Ӽ%��$����#
ot��#2���ӯ�F�zYZ�3��jB�6���FPM<'�0��,�H�p���j�� �M}��wd�6�A\��	5[�m����d�Г�h�l�L��_�Z��4�N0ZKO���Id5���	ԮJ�l��}Y�Q9�.�����y��~qk�<O���������Q��`�0m�"�����
h�.��&��W����~��ơ�;��F,�t�P�����lP����0cu�a/��p�X���$�a|�ϑZ*�a���AZ�|�e�pӔ-�ԷS��j���S�Q�=ѳH���2]�º �� �!�i�c5W�B��>�H\�~�4��p5��돭"o�ӏ	�MC�㜬�3e<���_}�ݣ��=�W�b�7.X��ߒA�N¬��UG�EH�O	�t$O��ک�?m���>�c��e1\���6�︤������N��Ⱥ���#w�}DC�J�TEO�4M�w&��
^�PYjB�Ns������G���+ `�@��6�Y�d�Mm6�NyТ�'%}���{�ÌMO�������%�A]�Ԛ���YE	��JW��LIw%ɝD���b�'dڈA����c�`)5���$��Jyv���Y��?�1~|⏚-�Hy��y6�a� ���8K?~%�G�E#qV�kq�_~%"&�s�U z%�L� �~��,�s�3�?�"n�̶k���m_tLx��U&oC!�Ԡ�J$���?ҽ��m*��k~
B�x��|I�r	�E��rF뺞�Ӿ�n����)��!�3Q�V}�J
�¼��6u,� �p�=N��tΞ�a���E٬��dS��]������;l0�r�it�(��q���� �B�y��t��u�S2-B���W��WN �Ά�r��s�X��)�L�K�oB�HqoEįO��Ԯ	pN.d���h���9Ĩhg����������)Ҵ�"��$-�Z2>�x&���Ew�=w?g�^�!ei����E6�Wfo~IW[?����d@}U��.�6M
G�7��?�:qO3�A�[�˙�<t�Šx���-����GBt�4�������'#UH�k&�,��y��j��F"2��(��g���nwA�r{T�E���+.�^��f��R��F�)g�TӈV(�^�,x~���W��>�y�xJNWʝ�gה16�\�p�uƢ��#ac� �1��e�=ʊ/W���&z�bx�[xx �Y\(�$ڴH�����g7�����
N����vMd2i�J�N�(K������ (3Τ�"{E=U������UNhn8a��I�AM�h�"�[Mr����!��Q����g��28^��h�8Y��sUuvn�{��Z�D�?x,�6�B���O:���T�69E�~�q]�ч&STԌe���I���as�ٌ�5u�D�~prv`��K��O��T�T�xY4��bؓ�w�(']�̌�<�>�傁��x�c+i���/v���\b�]<6�vOz�[�+O�Q�k�.�������h��t�Xn����0���7�0���͔�'q�ѱ����=`���"���S��À   Ud�@!�5����z��nzy�)��9vg��+�X#�U�Vڃ�i}�!�o5
�n����aM�`Gz**��jpw��Z[�޶^������aɯi�5KQ�ZU�@W�ㄹɍ������K�si�RY��+���g��_�X�ϴYZb`�u�:%��������%��@; *����[�3nC�z���э2�X�`�yf��GV��Zt_VS3l�+��S��(�en�$nxP �<û�a�h~� k��N ru�s���x��Y,�K����Le�vU�Xi�Y������!syx������Ȇ5N\K�+����GAK �l`�����v.��KGwZ�7�0&퍮|��Ś��"G�3
1TEW�oj���V�vՂ��x6�h��W�z��b���jF���B�����y�����ک�!ODF���	��m���)Ȱ�$�;�[��g,V8ın4{������c��8�����E��;��\k9:��N��"ZA^ A�&kYԁ�3�X�=b�
�MsџN����Bs�6�Z���g��	@��8��l��7Z��WW�@#�b����#/����N��u�Py��;�a����)��b!�1��9���d��	6��X��G&�X�e2J���	�LR��+��<&e�E��!�cޚ7~���4G�Í��kV�7TI[��S���s�sf�^nutDN*����x����K�F���hTy}SڻPGo"Ր�jIQ'��Ch˒��2�2n6�/���#<%���+��p���V�ҟU���3�Cb���QV�21?`�]�"G�3#���8E �n��r�l�+2\zHQ�cz5j��K	��k\z���X��G\�X{�q��	9F	����O�d� �aÊ���ǳ�0���b ��nW��S�+/��y�*���h�d�Hm,~��� �i�!}�l�2�M�?�p7�	�ZT�ޔ�i�l��#���?:��Ҙ�$<�Սj��R�� o<'���V��S~G�D�������K�Lҍ���7��G�H�ml��@�<�U쪕���L�C��n�@���(��A�l��hRtO)XqD�1����u�%e�3Wӓlv�8���vY�c�pF���c7�}W�*!���B��nv�ʩ���W�<@x]�yu2j]WuZ&7�t�k �<��O��*�ǵ�nY��R4�������ɧ5x���3o��q�	&�r�%׍���7E�Jυ�[ǫ̗%�US�Il��A ���9#ʀ&�����Kv���������:0H��I�9SQ�$T��a�6V�;050㜓��4�{���*�墽ϙ%�%a�"�5�:Ç���ޙnV�c�苌���S_yb���J�U@��Ss� �a��X�G��<������y���J������=�N�cp�[����N�F�� �,_�]�O�.r�����	�0�!e�x�6NMj륳�"�o�tHP;�x��NPp�t�!�� ���j�����#Z�!=L��yQ�I��z�kFu�Z����zB�ő��8h�=��k�����^�	������_�oO���_���7��TRZw�59�j	θV�t^^��ܳtS��d����,�]�Z"<�S8>1T��u��p#G*��Jn��O�h��*��%��4
c{�D.X��.���m�Yƻ�8�>��5�oG��Z���. [m���選�v,��5���r)�7��\Y�qqg�h�oK������l]&:Ֆ����z�[#!䀢]���!~�T�p<<����D��\H�D"i��4����l�lh��;_�_`��o.����c�rlEn\�ZzOX0>�Ji�F|���J��v�25��`��g`��c�ɓ�4-��+�2�O���~���Q`�Q�k?�-ص�.�$����L[.(h!,`�;��RAW8���Q�[�N�sp��jHb�w
�2B����7��go�qa0M���؝�ݧ��o?;������n��yn\_y��T_g%�7!9k�c٢k����{�@i(7w��Y���b
`ͥ�>��܎�8�	�$wS.ʩ�?���cƹ��K�Q��{�����[o���B.#Ϗ�&��QI��Ġ���\��B�p����W%��:�{6m�w�@F���vfD�˻T�a�T,�d�m��'���n�Ӵ�,n�ݯ�(g������ 7E@g�9�C ���O|�l���08IJO+P�E���y�k�f���v�4qc�Ӗ�����Q��@���Ń���z����3�g�2���!g�ZO�1��"�}�/�7̬��Hv�w'�;7j@;�C�Z(瓇��T�^P����"6��z��q[�.R>[��_��~���լ���dΟ~H�Gγ�8&�݇��d|f�S�\�	g� �q��%�������bka��w*#�0^�YK�Ҋ؞�jF��x�+��Mª��b(�a�0�^�ZZ��u{]�<�>[�LSr'�Mn�A���0�C[�H���O��D��`h<�޵켢�m�>L�l�	g�&s6D��k'�Y ��`z}K�Q�e��}��Ն*p�H��fm�rl?����{�8����>�Z�@(��ag����3�������C���p�:�_�|�,������x�w�.$EYg8قڦo:Z�.�x����O��|)�g7�v
���8=��Q����\�`j� k�WhG���|:�_��W�o�Q�mk0                    ��         ��  � ��         q� �  �         (� t�                     ��     �� �� �� �� �� � � /� ?� W� e� {� �� �� �� �� �� �� �� �� � � /� ?� Q� a�     |� �� �� �� �� �� �� �� � *� 6� H� d� v� �� �� �� �� �� �� �� �� � � ,� >� N� Z� j� |� �� �� �� �� �� �� � � 0� @� R� ^� p� |� �� �� �� �� �� �� �� 
� � 4� F� V� h� v� �� �� �� �� �� �� �� �� � � &� 8� P� b� t� �� �� �� �� �� �� �� � (� 4� N� h� x� �� �� �� �� �� �� �� �     z InitCommonControlsEx  comctl32.dll ` CreateWindowExA 1ScreenToClient  , CharNextW JGetPropA  �MessageBoxW � GetClassInfoW RegisterClassExA  � EnumDesktopsA ^SetMenuContextHelpId  � DrawTextExA � EnumWindowStationsW cGetTopWindow  � GetClassLongA [ CreateMDIWindowA  �IsCharLowerW  WGetScrollRange  � EnumWindows RegisterClassA  fSetParent �ShowWindow   AppendMenuA �IsDlgButtonChecked  mGetWindowInfo 1 CharToOemBuffA  �InSendMessage 7GetMenuState  USER32.dll � FlushFileBuffers  SetHandleCount  mGetLocaleInfoW  ;GetCurrentProcessId WTlsSetValue uGetModuleFileNameA  � ExitProcess �GetTimeZoneInformation  :GetCurrentProcess GetOEMCP  lGetLocaleInfoA  InitializeCriticalSection SetFilePointer  UTlsFree SetLastError  �GlobalFindAtomW � FindResourceExW �GetStringTypeA  � EnterCriticalSection  LLoadModule  . CloseHandle uOpenFileMappingW  �LCMapStringW  VTlsGetValue �GetTimeFormatA  7IsValidLocale �RtlUnwind sVirtualAlloc  �GetProfileIntW  iGetLastError  InterlockedExchange wGetModuleHandleA  �SetConsoleCtrlHandler ^GetFileType vVirtualFree SetUnhandledExceptionFilter R SetStdHandle  z DeleteCriticalSection D IsBadWritePtr �SetConsoleMode  �ReadFile  |OpenSemaphoreA  HeapSize  �GetProcAddress  HeapReAlloc �GetUserDefaultLCID  ?GetDateFormatA  Z CreateMutexA  �GetTempPathA  HeapFree  �GetSystemTimeAsFileTime =GetCurrentThread  �WideCharToMultiByte 5IsValidCodePage �LCMapStringA  �GetStartupInfoW HeapCreate  [GetCPInfo �GetSystemInfo J CreateEventW  OGetEnvironmentStringsW  {VirtualQuery  �GetTickCount  �GetStdHandle  
HeapDestroy �WriteFile | DeleteFileA �GetStartupInfoA 7 CompareStringW  GLeaveCriticalSection  	GetCommandLineW 4 CompareStringA  HeapAlloc � FreeEnvironmentStringsW vGetModuleFileNameW  OTerminateProcess  �QueryPerformanceCounter xOpenMutexA  GetCommandLineA �GetStringTypeW  MGetEnvironmentStrings HeapLock  � FreeEnvironmentStringsA SetEnvironmentVariableA HLoadLibraryA  � GetACP  � EnumSystemLocalesA  `UnhandledExceptionFilter  � EnumResourceLanguagesW  TTlsAlloc  yVirtualProtect  �GetVersionExA >GetCurrentThreadId  kMultiByteToWideChar KERNEL32.dll                                                                                                                                                                                                                                                                                                                                                                                                                                                                            yߢ�浽x��<3`�/J��X	V0,íb�SW_�$�K�m�
K�`,�/�lh6_`b}T0��|f]�-~���OQu��A $����4h(�	\�5�����xlm��Q�4��<���]��3\F.�mI�	t������]=�hĮ5��-º$e�+J���kz�+K3�^��(R���du��H��pT��H�O���U�mGܽ���2�!(������>��'h}��L�z=�]��Q*TQ;&��i͖'��)��/�<�j�¹
G�h��y�3|�җ�V�/�9q����qm?Ȭ�����kl�E'F���6U14�-��Ym��j��Ȩ��tտ����ӴxE�+�IQ�E�l_5�7�{9�$=��_B����I��`�p�ْT�l)eM��"�(���L�"��-�P�Lx�����8� ��T�ԯ���a�y4y�����s^6 IH��/d`D�����P��n^��\��n`d�p�n�?T�1z(g�xڊ�`�ܟR����t'�v�6���30Fm�	����I���#R֒mc���Lt���X���Ww�'tw8}�粟�}K����ǐ��>���^���Q��D,=a0�����=Zk9�i��!�#cC;N��h�LiR��ny�禎�1�k�I�((�AC}y����
�\8U* L���*�҈l�Y8��r���!â���T0�"a*�����S�՞��gQ5��9��[�))Ӿ-(�G�YsU�f?��l�e���u��ۋ��j�o2Ơ�\�#e󇼡]�-R��E�b�~�A-]�<�-əRy^F�[��7ύ��p��4���5@[ڐ���r�('�(e�Si'� ������A�X�q̕���t|w�Cv>4� �?P�C�tE[.�ΈY�D�P�N�ಈ*�mM�����7��pcAj�*�q�MCkF`��ŉj$U��F�D9���L�Bk] ]�7hk�[����O����V_�l��n�_7}@��V��j~���;w!Ŋ��uK����8�#!�KO���J�zmB*�i��8k���j9 �2#JEh3P �{n��^��8�(�܍F����3��jK0�����n�(8�9�]������rZ����^���Bwh�:�:,O�Vt[�f���|	M������"TJU2���LY�l��=�jq3�;ߦ�z����#�8�����%�9����@����C4��?Mc8ϊV�~*;����	����F����}��1���A�Fh���lC���(�+L��_������e	Y J���5��~�4�[�D�,�p���K��I��v)kX�r�11�����F�`���4C��T+���X'��@��X�|��!��tm���k�g.�i_���ڟ�rG4��0�GU�|����|.�-���J{�#��ա��j��`xݺ�3�#xC�׆S��t�Eɖi���c��^�T*>��:�#��8p]Ȼ��W��:���h��̨�9���G_�w�<f��SM�d>9����j��9(�Fl��?�|j����F�4cz��P�7X`�~����X��gm	��]����7��)��pBcX'�{�EW|���~���"p`d�e�~���>�b -�ٚ��Q;�>�R�"�`�8�T�L� �Ͻ�yW��(��1֜`/��bU��XS�
�<x�d�TB娛n�>���Y�
�m�:�%�5���Wji��!��(Zx׹#Ő���idƩ7�*s����]�9F��?tm����Pe^��R��v�a�	8G4�IT����S��r�{���VV���6[´�O�f����v�ԯ�g�*�	�ml�V��_��쀷��:�؍��ոn���X�~��\t�ӳB�52z��t�v��V��wL#�&�tu��;��?C�bQSe����8��AB�%��[6o+���;��D޺�ZHC��wk�Z�<�'��/^m8�==��!���	����W"�`�A���'E
��!̈C��"���n,����ȾD���0�w�?��8ru���;@`8�����l��6�,J�f��,�� ���ג��z�dop;*�g\[t��p?= QZi3�f,(�(�"NΈ�/�Qo$+����8WC�G�kM���5�l��/;��-14������VMF_Sjp�U�>����u3Y����y#���I��
�`�z�pt��I�ʄ��~^�0,V�Qׅh}Ge�����)0BO1w�7�`�*��\�ӹ&�w�u�63�� ˅+�M"P8������!�{�m����bx#ɐ��
��/�)�`�����W^���v����|�;'�%��j*����.f��З��O�(go�3 Ibl�W����=*<��Ͳ����!��K2N���SoeQF�?��rHޭ
�ڊ�c�[	l��~j�{Q��7>��/����[�M�p�6��]�4�XU?�ֳ�Z���jc�&�d��r(������(m�C����t����$R�`\�&�"�o��h�F��}�R�,:a����ػH�
gͦS`�n[�����2�1%~������K���6Xz��X��o�/?oz\��2��}2�F�K>	����,��Ɗ��+D}��>dv�9���cWjG�TAgfSW��^�+t���a�mg8NA��Ig`%���-�=��wm܀ ��g��g����2d��,C���g�R(���!�Qh���Юg�<O�n��1n���*��\h���"�#�5F���h�>�'���E�����JX�RKCdˁ( 	躠����I�E�ɭ��&t)e�^�K��0Q�͉cq�"_���?�wJ�ә��J{�9�(��nSB�tN�a:f�ɗkL���*֌բ�C �|�&��Jpۻ�;���6�BäC�x����o����M�ɀa�a��sΊ!�[Z꣮&�
zS�*��[�;FA���Oz�KCu!y6�3�,+�<�V�������Y{��������y������VO�����Ȟ�"d�LC=]k���t�c��g��s�0��L�=�0),V������	k��]����*Fߜ=����?z��\�3-Q��7��<��AA^���J���³�.�	E�9,4��y�7�����̐��ј�g���ڛ*a��ܯ�~|�Z%����k%���]r\�$"�'X?G鹘gI,"�.@��J(�����/Z���V�x��؜�iu����7�
:�|�3��9Jw5-|z����Nd3.;��R��ѧ|�9��m�Ig��/�#�-�=�3�Q�i&�*љ� �Ğ�ޔ�Ms��]V2��5�ÍD�����0tѣ�����"�ŋ=Y�\�R��`�5����G;��z�L00��)�\i�yR%�������Fo&�����"#�#3��n3�')���	��s!I���p	���qť�k���H w[:7�J/����ύ�vX�X���#F�"/�{�%����x�>J�lv�>*�����+Қv*T��oK���45���y5�S!�/�h}��9>I���9�d=��|����n����Ǆ<V
��PZ~Ǒ}��=	2J\�E�Y��'^��:��<�=�oxk�� �N�kth�M��lH���"굂�-ʼȧפi�~v	�y�<Iv���	�G�X��Jj���_��6YTst#l#��>wb� [��Ŭx��!��W�$�F�5̴!9�NP����E��%���ܘ�T����Pߒ��0(~���W(�<!eeT�/�H,��я~�'��<3�5%E'тsVz�e%���Pd��~8����/_�<�V�S%yߞOL��6�IL7˦t�@\�?�_�T�#c�����G���0KH][�bc89������M`Iv���#�7�zc��$���Sふ��r@���\GZ�,fI�/�-%�����3�<%)C��yw�� �fR� 6�R�_:s�����H���<��&��V��#�E�m
{��ͺ!J��~�1D?FS��h���6���2ڌ5���3�/��f�hQJakw��?
��=K@s���CR<OA��%OIG�CuW�P�� �4��F�����v�w���X[t5g:&1��H�:��姅n�E*"���t!�,���a��d�-��|�N�H�33�H�ѵ�Λq���uOH��3j�k�f�S3;��5�f�.\-�t���'�T3p:8D,�m�;�~�aE��r��l��f�h�͹�B�4]9o�0����5�H��+>I	�R�j�d-�X�~��9��p�a����/�� �G ��G ��G x�G 4QF |aF �sF H�G ɖF d�F           T.{���'��K+�D�J*j��	�,���Y?ك�?�pp��?,|*iZN�z�o
���&�Rm��M����s�*L��]���+���x��s�@PU��W[(��w0���iokG��,Oĉ��*��&a[����З�Î�`����ժ�>2�����ʅe��;v�#u������c`�A���u���gR��9�47BM�22���A�a���ˀ��U�9~�U
/* 
3�r�D�����84�!��g[�0#��<�"�B²:�#sX0�	Ս��XG�˻�r=ziޟ���b�c3�:u��,��[A��ŏԡ��1+�IT���?��U��Q(�KBs
�`<5��C�l5[������pv䑘\�F�4��]_^/� eQލѾF �	��0�}��0X5i���Z�?�Ͱ��w��`i 7]!a��jQu���{��Fn/I�/�FVDF5��,��F﫢&���_븎�D��8����'������k�'(�	��:���!9G�#���OS#'2c�7�xp� 9��0I� O��8Q����K���T:$<��OH�z\A�>v�$D9�����Q���]ك뻣������LD�t��L�4�2����b�|�hwf��<[k�ǌ(��%�/�۔9oz�+�t���n��ڕ2�ԑ�e�����]�����k��� 
6]�f�C��b30:H�[1TOEF�V�u��[!����c�۝l�7V8Tt�K�����E�'O�b%�e
D�*B���jq�Ku:��f�0�V$&�P�r(�$�E����^�a�P�n��@�������ZcH]*d#ʜ����d�K���V]P*�A� ��p(�� �B�T�*�
.��C��!��ܛ���������o�����%�x�0T�1��7��.�ۅ�����
�����}�U� ���|x�� �֏���J���iX���jno� 2�'V�ƞ���S}E/�7�#Ra�O�/)Ϯ?�j%N����yaTc;f~RE���y�ۯ2x`��q�AA��w{&g�v�"�)�	��9���GG��(l��n.�.�+�����ik_]���f�ȳ�8GY/ԗ߷��%��q.b��k`q���T�6����s�r�o�wEV �~�������1l���JP`zgq��k�Jᐯ�k[�%D*�勅}˗�S�J�u�������G���~��R0�b�q��1����ʯV�qxK2�k���
%����UXf��+r$P�\y����Ԭ�n�T�	'd4�:P���ĩQ�&����2R<\������}OI��dt�i2X8�F���R��|����f�-��SN������ M�����L^�
��Y�]�w���qA2VD�۳}v9~Z	w�+�R� Tm�z]d�n)"�o^Ng����ș�8���F���%F`-��in����?�h�F���U�O`�Eu��6�B�������u��X8���T��z��W��ZX,��I�e��w��\��|/�!4敘��	�ҽ�991��7�'�3�I���d�D �p6��y*�/��Q$�9ۤ��|I:����7zRi�g��J0��L'�Enq�3�(zR���h��6�>�b�g�%27��ޙ���¹������g����I��5�02	�`�ޣ� ��>�Fz�y/�3���1��8�GKHMq"|����-O�#h��<���vv�~�߉��U1RE#�;9��L�ק�V�@u�	���Y���bQ�����ܑ�Z%P�}F�Y�)��_���a��.���şe3���ɻ2����n����CA圎$��ZIgꍩH�%��ƨjv�u���e��_�������Bt��/.%�I쮅���Ӭ�r��\h5 Á6~{]�-L���>B�C����O��X��]���{�I=z�fH�"pFݿ�08�����fDrk��-M;VHi������Ԥٳ����jzL�n��ΒV�3��9���v�qOυ�K,�1���"�\��U�Y�(�ʣ�����.��Q�
�G��?��P�o$F �5�L������[�~��G%H��X�>��GJ���BO#�`���4)U�P�
Ղ/rK����j���y�Cރ`8�Uۚ)�O��Y�~����C#�nj��M�"�)�S��k+{�eh��FM��������8P���	��l�����<�X'��)��_��9T�M(
��7���J͏I��!�n��*�#� �����,kR�J4-��j�?���NsȰ����y0V�.=B%{�=;���sWe�Bu���K!_Rү���>��k@0�J9==��dG@�	\��\w�9ή����F� i^�O��m#J���W0��ޯD�c5#da !�ڲ� �'�g1'�y�!�qd�(���	{�]�rl�<��k�C7���-�@}_�����&�iy�y��n�˛3�N���i��^���ѧ���SS��}b�6n����[����+ ��w�ĩ���d}��Ku���z�Y��}���L����*���~t�%<t:Ύ<N�n�G�Vn�	��qn.��[��@�I�dd�^V�X�0��o)m� �oBI�V�M����'v%;Q
v�A�Vǚ�5Z���5_2������,�I�Q�]�0#��]/�~z�H�<8/�J�g`;�G��tÝ�]UH�FH����|�V�j����eu	H#J�1=:͏{B���ۃL�w���q�����q7�Ҝ�����E|��'I��{rF���/�̬�����;h��'��@V6���5���Q'�6د����R#�j��$��>�5W�� ���N�|M�A/a��yѩ�6�\�P
&�AC��txf)Z�îӑ���$�Hj5�O���:*욏j��T���X�ۢj7��l
h��#=u^��!2R�5LR�tXm���.R��MT���tx;�
�V�HN}�]��R�j�m"+S�N�J�b�ǐH�L�8�!j��Q�~����>3'�<AM{eC3K�ЬP��R�)�#���}��-�p�ptm%z3�1ĿZ��H�`B*#vb~�e��s!KÓ�zv���@qv��X��j�M>�7���ƶ��M�i�t�h�Mf¦�w�Ĉ�[�T�8V�)�6�t����lw��7/��\S�F5+kD3�[L]�ߓp���=�R��Qsځw�$_�JՂ�O|�6]��=h[8��>Q|<�I�~��b�\7^}�#;��"�p}�J��2-����T����=NgŨ�r�A`ϹmQ�$�˼w�G�{y~�#�������&��T��j�۩+?�kj��������u!�&�6|]Rag;�NQ�$���Gv	�^�պ��p�GT/1Hyx�Dj���h��!���j+>�vr>�4���X���i|g:ZV�:�|`�!.�;�X�2�� :�≣��,W��Y��T��R�p
?:����Vx6O��
�GQ=ﮘ�TJp�Ga�g<YoZ���\d�%'@�����m/�6�����k����e Ƃ�L}�I��?	���2&A���L��8݄���ь̊/1����J�^��.��Wl̖ ==W�(�|�-�	�9�\a�2�E^����7�-�HF륾�;%t�%7�!�\u���W�%u����G��)s�W�+�!��$4�6*��+��U��"�O_���(R��]G�̃Q�?                                                                                                                                                                                                                                                                                         ���'�+��k�w����t��	���(q�C����#���JDV����]󕳸Lt!�g��_�oR�]Uӣ�[Ad�aO�3\��(�F�2�ݟ:�f�>��QgKuF�́iIif��<��a:��(���_~                ��h�M�!�WZYX��iHh��Y�Z+������܈w�w8j.-o��%�ǅ{�nl��������?���G����j�����c�e�Me�����������P�k-e���\������pW��XW<\lyf���8�n�Z�����((�8��R�܉wqN���j�-s���_z=Hm�Yᮖ�Bv��Г�dR�U$;B�_ݢ�M[|���W�π.�ϣ*�t��<O<��X��cЂ���!���)S�;�uG�w�B���('��UY}����^Gܺ��3��gİ� ��϶mJk���E�"��Hf9����-���7P�G(�˺}�jFw�PR8T*J����g�@g�G�ha�~M?)�8���&�0mF�Q@Y�m"�W�<t'2]y>��*��^�8�^-u$�to�J�
v+�ނc��˒X�P�����]�#U�e���5,^�t��(8$#��e��EŒ��(i�{�y�I ��:lCWV��= ,K�����p��[�m��X�%(t�l���E���i��*gV{��D���Q|u�E儼7��&CP璍��e=����]�g�0d��&Q4�k���{DP{��ڛ�?�to��&�pD�T�ܥHy���H��VgI#�'�C�K��5o番9<u�"�8F2��c���%x^%10d ng��7��o�z�DP�4g������rF�F9g9���?d��SW�N����}�1 Y{&}�?gnu�-�$4��Lb�hh:_D)��p�yIi�R��{K�4�!p��!Y �4eES�Ck�T��TDPYCG�
T�`�m�$?O�f�"H�,{kk�� w���La7t���j��_V)���B��ƚ��4C6����/��]�e�$#�oI{��0�wf�4�#M���E��=(ȷ9́M',>��pVy��<�OC�4��5�@�B���X}Dg�����|�G�C����c�������"����������g�d�?����k 7��#�����G�7�M��vi��ջH�MZ�����_�ѧ�6ـ�c_Ѧz�������QL�r:C�xJ�.����ĕM)lSW��6�
cM�U)y���g�?��~g7��jr��^1�j���q��cm����L�qoְ��9,���db�@l��o�h��@�ݺ~�$HT$	\MfD��%YVc�q� �1���^�8�D�`�6b��Ƒ}��᡾�G+��c��'�%�����B�1�m��L(��������mƾK���5���^b�#ʌ���-� owLY�6��hE6�q�����ȹ
6��)ʿ.���G�ʫ�@��	��4'��3�?1X�\|T��<v�h:kb�+��q���{!�v���%��������'�lR�tPk�&��tǅ�A���4��9~�/��"x-��Ȉ�حJI>mB,�t�2��ђ�y���B�ewr|w��STé��3�j��
��_����a\<�G>v�? �]~
�n�/ܠ�&�˙��};w?s%#.[E�^ ���:��+:b$�B���ta|�\p'G���_1-�y�#���ZY�%x)���"�J�G��5�^;�|�_%�
J��e!�Z�$�~5ҕ�A�	fݱQ������<�U��r�i�Ү+���\k��lKmy/��9l!��O��5���ZC8~�g�Y�~+���(��ߎϰ���.~x7ɦ��R�*r��L�5��|K��K�q���c m�6uqf&�8�7�R��u��)�;��H��l�zZ+���朌��<@�\wmC)9K�k��0%�����'�5�"�W�L�J�Y�X�v�?��`H(�����P Ш�M$��~C��S��������KV�Rd	}���EɺU#�ƇaG�g|-wQj~�n���I�Lm+�o�;3Q=$��������D����Ӷ0�ȗzɼ����C���~6Fydz��,4�d떷Wq̃�/�NtYYxE��vj��!����c��T��~�S=d�e���%s�g�b[x���zޖ��qJ�@�҄=~��8ʶ:�g2����3�k��KHﶼ�@Q�$˖Y�q��bێ/�k����1欘���׀؉TMT_@�=\ʀ�Si�����3j6��'�N�F��8Y-�ޒ/ud�5���s�]~���V1����gK��8�~Mmݻ��$�s�J��i�|Q3,�7��|1��ċi�t]��ֺ���	6T�����ņ}ՋD97R#v���8�%	av#'W����DgCŦ�3�I8sU1� 'e^\���Yb���M��0G��(�t4�����3 b^���R�C��7��L<���e:z�A{��Sc؏���3�:��@஄>山��uo�wd���P���g")::.[��M��}�}�Ta�=�a�p%�{���2t�=~�8��п�|5?�^��3h��p��FID�T�Q��M|t��׀����m'l��Yn�c�"gЈ��:���z��V�Ͼ�9���5�ە�-�=��%D�-Gy{mPx��j��v�hU.F%�&�{��Z�dP5�W�3�z�/�������u���1�+[����N�����&E����ҝ���;}h�5�(<C�E�oN[��f��m24�j�E�w1�E��kA,+2dqu����[�}��k��R�O-��tG#��S��߶G�h",
RM���|E$/���w�D��a ��p|�Ϣl��5dZ���ԍ��a$T���T�j�x��s<1��]��|B4U�	&���0�gWl1 (��գ�X��}E���)�7g|�Qg�4�W���`K�Nx%�סqw_f�q��ξn	�:��J�ˁ���:`hq�UӐ�~��(Bt�$-����4��+������A�|DVYO�l _v{�ˇla%[#���\��̀��:���m���]֐/ S�i���{�����G�w�>m��rWH}(0�m��!.��}Bg��S[�U~O���+��Dh���|�Z,����3Y��N�����T��o�qĞ�Sn�ׇhI㒷              ����#c?���7'    �����4Sg�;rsN�c����X�{���1OWr�L�JWeK��:)?n�*9k��@	J��R֥���,b|�h\gO�<���Sv���`h4qpRu��;7�h��������������9�O�BT���=<5�@�V �g�-�Z��׳-!K{|�h*�e��k/���t¢����S��n�O�-r��^s+�j{����z�}
,#È��i�a���d�#n����O����s|�,�X�r�0�
����Έ�>W��=����~������y0ж�O��O����7yKM$��[f5�j�Ix��>�7��� �At�p����%;�<��\��B�<D��#��w�cYJ~֝¶�$P�����z_�a
;ZS�p.�d���2��	EӍ/��N ̐���̨\IfCL�L^~��K�9?%�ȌK�H��a�a^+VY���B���Y�MiG��2��E�ݎ��O_�߳�����P�zp��W�Јs#�/�6�xf�,�iUǔx�%��؂ͬW4��#fKb2��;4�S��&��{�Nw*#\J'�0�~���d]���Um��
)�&J����2���ń(7�
_��GVu��ˣU����4�n��]����d��
f"�S1��?���q�SC�?�ө��v�&�(O��Oj��f,FZ����d7����&juv�N���������NO���P����L�?����H�~�5��b������7G�5%	�!C[<Ă�x�����>>��=p��jcf�2\����%���h�8}k�2c ��㢑�(�����N��B��#��� ǵ�t7ɽ�N�o�n��ȸIc�	�(�u����b�j�"����>mx�'��w�������$^{j�k/�H[Z]�P����B����7"@&��uM(CSF�
ٰ���)��w�[,Q�[ow�4gS���4O���������L��L��Nyle�L���Op��A�fP���+�Ȝ���!�~����h�uzM�9S����Y�C�{�W~�ҋB�ZL������E��AJds�5;�����z��4N�۝b�T��f���F�i�6�Aw1�L�<��G��O��J���E��Iv/ ���u���������["uEլ`ܾM,���Z�y�N�/_[Cw���72�i���6Fe(��>;��̇���<fI%���c��W�\��M��6!	NF��c�q�A�IT�ƀ\}���VŃ<�w��vq����c���.�v�ʮ�T5'�
���`AkY�x%��?GnZ�$:��DB��Jt�$�_�ڜ[~���T��:#������q�}%�Cِ��ޯ�
-��2��9�+K'u^�h��[���Ya���#b�`q�F��ٱ���l�� Q43��
e��'=PA��B�m9�T�3"y�u���#��c�tC��Bp�ظG��[�1��ަG_���ߌ������E)�L��h���^Y����>��n
�����?��q��D{#��#!e�i1�VMb�!p����%YD��Ncl�����t�!ar �VY���~v�RD��5�%10d . %10d . %10d . %x y�q�'�k�#&x�*8_WE�;d,ٍF��g�&[�'0~��i�>�����s[��v�vyxnk�Y��?ǌ� r��8(�o��ú9��+l�/Zw����@�;��Պ�[h�:�����:���4(�����U!]Oֻ�x�����Q�~n�[��N�!� Ջ�f&"�`g�s���̉_� ���Q��ˏ�׉�l�����e��?�X�=⋄�T��$M�ϙ"X4�0KPX̘h��=�K��1�@i�>F8���.7ɖ�3�    ��"_u�ϑS�٤�dR�jQ�L�b^�4��    �~>7^�p�HRN ��������Ve��2q�6qf��(~����X��e�s�
� �
�=+0���r@�pS�ve��xd0�P\����>��	�r>��M�y1�T�\2�}ߛ���U��<���    m�8'��0�Pv۷u+                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                �ʎ�^��WT��KE�K�$O�i�R��������U�P�Z=>���A9�HD�����=}5Ba���b"@u�;a�F�1��5dr�f�8<͓���yx���oآ?Q�{r�����ԦX�p}���B`�G-�?O��j�M���w�4��oi��+y��.�Ҭ1%\aZr����$����    �
�:��V��                                 	               	      
                                                !      5      A      C      P      R      S      W      Y      l      m       p      r   	         �   
   �   
   �   	   �      �      �   )   �      �      �      �      �      �      �              �����
                                  �  `�y�!       ��      ��      ����    @~��    �  ��ڣ                        ��      @�      �  ��ڣ                        ��      A�      �  Ϣ� ��[                 ��      @~��    Q  Q�^�  _�j�2                 ������  1~��     �            N�@�@ @ @ @ @ @ ��D ��D .   ${F d�F d�F d�F d�F d�F d�F d�F d�F d�F ({F    .             C                                                            ({F             ��D P�F     x{F                                        C                                                                                                                                       C                                                                                                                                         �         �       �  �       �  �       �  �       �  �       �  �       �  �       �  �       �  �             x   
      � E    � E 	   � E 
    E    ��D    ��D    ��D    \�D    $�D    ��D    ��D    ��D    d�D    ��D x   ��D y   ��D z   ��D �   ��D �   |�D                                                                                                                                                                                                                                                                                   ����J@        	�F     	�F                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              lE \E ����   ;   Z   x   �   �   �   �     0  N  m  ����   :   Y   w   �   �   �   �     /  M  l  P�F     �E �E �E �E �E �E �E �E �E �E �E �E |E pE lE hE dE `E \E XE TE PE LE HE DE @E 8E ,E $E E \E E E E �E �E �E �E �E �E �E �E �E 	         �p     ����    PST                                                             PDT                                                             �F X�F ����        ����        -d     .                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                           ����E�D�����t2���F (�G 	�F ��F     �F X�G \xF p�F ��G                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                     �S��Fɵ��gop#7�z�9��T�M�tJ�&��V�ݹ�)�HH!N޵���#��\!��G�gdR�I�Cդ�d�C�)��|T�(�,��X��u� �,k�u�9�j�1Kn'�e�P�݊��&>ï���ᑬ{��Z'cn൱[t��Q��`�	��F�            �W�7"߱��g    ��������<q����5}D�����t��٭�ʃ�.0ϩ��q�gn�?�        m�s}�Y��j_�A��D�}�g~=˹���,�|����Mpw�ZǾF��d�:"�}�r�ő�R�o��檾!�?r���i?
��[��b�"��k�>�L�t�5}s/t�᧺$��Љc�-�`�����o��n*2: �;�5�f�k���y�7/�E��`pi=�AZR��`Dm���#��5hq�e}˶��b?�3�r���]+(fe�D_�B@Y����C��\B
d"an����d���u_�z�R欲+�&���Z���ĕs��o*f���U��#[;/� ���c�F�{��1�J��/]�b1�N�D�z��2+�	���5X���^�dk �G,+|��ۅKܔ9m��@���|�Y���� ұ���;V3EA9�� 4X��=#��`1�D�Ю�c�R�ǄF���W�����A�ɼkd�^��ր�u{��<�kٜ��/eY����S����s��8Vf)����sdN�˲ǒ���y{��l>&I�v���˙X�-)�k���u7�]�M�C���$EN�B���ş��=a��i�9���',�D��x�=s,i�t%����ލߒ����1�:�iO�	�%t�o�e]�D����_[���N�[��􇶳8�	se(��н	�\#����ڠJKO�3���'�!ֱ��S�ڰ]�5E�x'Ԟ���57�=����<#I}O8-k!�9�\<�_B����Z��-���H���	Z�I��Db**x&��GrD"-���,i���7�Ԙ�jh���<��>uo�1���G�n��m�h�I����I�W�W�M��]��iMn"�ca 3X ���GL���<)%�D��ב��`F�/��k�K�
zz1�hN,�m=�x��pQ�0}H��!� `� 	��5tg�p&f>�I)����^�ܿ�$24�?�5t�4 :�r6(m4�T��s1�礟6�3v(w��2�KQ���ry�Lg�p�
sY6̒��/�"�"�T��f=B�b-ࡢ뚼�h�ug�h���'+��t��,]�9� \�"~e��׀&\����woj��T/�xAj
	���f�ąVN��9����F�
��J���e�~�>`�?y$"vg.�w�b����.���*�֣\�;��Yq8�H�sC��x-�;I�KV���?�������f���l��[	<G'i��`����prE���o�d��g���_m����N:>���Q��o���?�w��X/��B��V���=�8��Xl"f8�Rp�^SS�掞B���l|Tc
V֓8.�u�R����bGQ�qs�V�6�.2��7��$4���$(k�7L|�IMg�G�Ȁ�WA�6�D/��1._{�-����4��Nhc�*�b�xX�v��[�	<S܋�qi�������yqL�'%¼�3���~�:絀FЃ�=*fՇ�@0�\��.Z	f0u>��%)ղ�DX9p\����j!�>%S{<��b��n�*Vt�v.96��NW�����x�s�U�u��s��,�Gqd:GR�{���/�%;"�&���r)���/l9+$�r�c4�S�����9�I�7S����)3x��윯�0 �������oO���� J��e��?D7����F\��
�"m��k�K�I#��0#��~��������9I�	��1c�����O�����R<T�\S�ZN�>�R�y�iC�x�&rޱ�W���A�p����f�3V��"KX�dJ�&�	�QJF��H�	��{�عC��R�ɋ�`�ψmF ՖF xmF �tF ͅF ҳ�eg;j{/���/��8r/�����(����|�	=��홦𰞉x� Fkf�%���]��+�=��ݹ&VT^���L(%���V�kǶ�/����3C�΍9�� ����o~��_}lh��ɫ��gy}/hCI:��[�*D2[re� :�_V=86���lė<�f"����&�]�W�.��o�\���ԏ��ǳ>�����LI����<���^5sޤ\8x������U�A�Zv�t���Y �)��O��*=�I�<:�_����Z�O�kyv-�.\�F4���gdB8� �`�š�rrj��I~�]���y��O<�.�K��-�������]>j���2.V�����1uC	��/yy�)�d�ߊ ��
����0ꦺGr<A��x�U.�Ip���rx�ݧ�u1<���=2�W���^fЙ�ȡ� ǻ��/:�%������]�������Q�Ҫ9��_�t�% �	G@2�a bfH�CxO�j�{AAa�g�	��x��pR�|lU�0�ٜF���w#�hz��&�R��eL���uo������q}Z���y���Nޔ���-�trBƭ�*�I�&�D]�G,`S ^����Rτ��}v�f���5�{�3&௔:?s�3S�>s$l���䐲on�@$��{+����|��;��M
��!�<��ȉb����̥��Q�ش���b��� 121�1b�8�3�i���ϵ	�l�J��*K8�Q��@�Zx�����Ār%��a��֙/��]�n����i��|��88��2���1�s�k�WHW������9@���c,zߥ`��3CN�P$D���F�"��[��I� e^%�u}�H�S�1�t_%3*w�F/\ui4��2�-�-�����@��9�e#�W�e�q.z�������#׎�=E �D��3�ƀ�w�u�YKԬ�~ �I�r��IIhx�����H2�揇�u�+���dσ���q�'n������)�)�	$V���9,�7����ٙ�Г��w��2 #?J��CZ��x�p:��3��qQ���m�/��yH>P�r���4���0\��e2���A��4(��M{k����͹g��[�G�c��`�j�.�n��8��ٷu@5��$o�w���a0�f�����Ass���4�4N�b�7-�O�T�gd������@��b)")yO6����y�1�U�#�CIMy�D�� ����]	j -S>�o�ٓ��
4:=��$l�C!]��T���B9+O��乮�ש���s��To�ETe)���B�E:��\J�Qlv
"�D����_����M�6���.�2]��ԏ�������I����|���� 2��Q��Աq�{���7|d�x4�F
Y�۹��Y0c���mvo �;M�+t2�"�"�:f��f.4+P!�(T�,ª^TO>\�uU��9#��6�{U�^����M����_�xa�k���L�����t|=H>)!��A1��Ζh�>��H�M��"�g�TK�l��x��Q$p���$�G�m���J�@{)���g���1�g��pȥ靈�c�����C�oN�\��*��F5Rhd��&G�y5&p��sT]
(���*]�
!\g���mQԊ�ϫ�N@�LVF�/�L���=��.Ұ��{��ƦB���L�#{펳�׷%9�*&����s�EH=WX�u��_��EQ����!��(o�߯k�@g��_V��hu��|�h��$?`�؀XS�L�VE>w���(e7�dpv��ȶrW���=���!�h@.��e|��	�o\v�Hđ	!�f�w�
��z-x]`kP9�>���[��<�׀��U%���0Q@½��zMeY-]�j�:M� �i�}��� �5��X���@y�yo�����#n�!	��b W�N�#3ZENx���Ia_��?{�G/1n̈x�����y�X��<�.����x�Cxj��(;S�t�-�f:_xo�tb��s��a��~��O[���ۺ޹��a�{�2�^+�[�W������]�%+��s
-��۵��"K)�վ��!��UЍ�@	�S#��c�!}��o�$e��h�T��d|	�ܮ���;��C���p� ��r��&�D�(�:f��aa-4��ȯt~�H�t�L�g3�!�,}c�T0�cOƬx��1liȓg�2��o~�@��>!���lbL6 ���b�gu���o|h����됾BK����?ѡŽڰF���Js^�����v�U�ޯ 3U6*�V��]-�
���J^��y���w+�7XQ#!+��C`��Z_�_K�M��#�v��}^,��s����z��"��,M� �����t�\��0��"�֩`5��R���c�=�Mw��G8��wՁK[B
��s� `�m.�6Pe�)ߐJ�p>�W�5W�LY���D��pr���ݔ虖_��>b�#��ݫ��l�m�"�Tyj��\�m�R%�P3�}J��;e�g@%è�1rO�iO�y�]��h*Lߢ�ё��c�9�Kf��w~�U�k�:�.���␽�z��+��S;:����C���v�2�Ak��N*͠�R����K�5��Y@����-�^�&I�-q�҇�'L�i�z�S�����?�Y�"#H��u8�]u�0��ut�L#������į���w��wP�)|��=o<�K�YSqOG�3m�x`��V>�s8텍ɓD��wL_�
wZ�T��
?߄i˨p�-N2���ɌX"@.G�\���W����F�X��3�C��p�Э�V�0V�cX�@���M��</���ڥ=F]+e|H,�z����;�K![9����-x���*R��8�:5K�����G.술�������f�u�լ~˴�����P�}ѭ¤��H���8���_�Sn"˼���\��e�����/�[�Hȟ�7l�!���ޕ�>�_ى�����#�W�4���δA����r�����fp��n��t�\�3�چ�6յ�i��T�2��{���6(��}�R����=`������m��fq�gӎ1cN
�e�^�!��@��X|��ku�JOv��/5��"�"^�~td���)�Q
�T��/��՚��� ��:�l!k�k"�V����W��ܡ����Yۤ�{_R�_r���� b���&v�9�
p��~��I��J��_��V��I�'IO.�\=����9B*�,�Ѵ�F��Q���5C��=�?���w#��}� L#���kA�%VԲ�'��y��R�y���J�%��5��[����h$��N�ۓQu��1�BL��Z$��lR��O+ތ=:���?�Z���"��O�y�P�����&qL��,^�]�p���1)�A΄|dΣv ���۾3�F�+)��k�V����z�(J���8������GU��������E�P�ө	.%��bly�!c�h	"x����ج��Gj�Xa#�9|裒�$����r^"��&sA��K�rQ����i��3t$�qCrݔ�x4f��~��]�P��d�6\�#��:��{�,�܈�LR�)�>p��H�n��A �5�i:$]:�^t�Y�e	U'&{�f��]3Үux��F����I��PeT<ҩ����b[�	�5��տ2C�bD                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                           \�F ��G �F n�n}�U��f[�5��@�y�c�˹���(�x��ƿIls�IƾF���`�6�y��n��e�N�k{��⦺�;n���e;��W��^�� �g�:�H�p�1yo+p�ݣ� ��̅_�)�\𴜂�k��j&.6�7��1�b�g�u�3+ �A��\le9�=VN�\@i�����1dm�ayǲ��^;�/�n���Y,v&ba�@[��;Uܚ��?��X>`]j햹�`���q[�v�N���'�����V�����o��k&b���Q��W7+�����c�B�w��-�F��{Y�^-�
J�@�v��.'����1T���Z��`g��C('x��ׁGؐ5i����}�x�U����Ν���7R/A=5g���/T��9��\-�@�̪�7�N�ÀR���O��I|�=�Ÿg��Zx���|�qw��8�&ٜ_��+aQ����O����o��0Rb{%�ƹ�o\J�Ǯ�n�~�qw��h6E�r��ǕT�}%!�g� ��m8eS�M�����=F��W��qwp�5Y��a �1���$�<��p�5�j$a�l����օ׊���)�2�aG�xl�~g�]U}<����WS}���F�S�����0�k] ��ȵ~T����ҘBCG�+����Ω�yK�ҨU�-=�p̖���-/�5��y�4Au#0%c�}1�T4�W:���R��%�������R�����<Z�"p��?b �$x��$a����/	�̐�b`��}�4��6mg�)���?�xf��e�`�A�w�ŽA�O�O�E��U��aEf�[Y�*P�ҹ?D��w!�<q�����X>����c�C��NNY`F �e5sT��4���X��њ�W���-l;�<�^!���2�����d�-l��1�j. e,�L��k)��p{&�j�J���*�C%sk�jq�DWT zGQ.�^<�'�}��L~�^5{%ؙ�㒐�`�m_a`�y�#|�H��$1���/���u]濫xT����og�a�
�wL�p9bݐ��^��}�MF���1����.���~B���U�*g
�!��m_mo�6��xxT��"
�� >���AE0� �k;�ep%��3A��~CNL��I������s��@�kS4?a��X��	xh�i=���g�8��_��We��z�F2�~��I��g߸�7�oސ��P'� �:}��ܾ����+d�90�JD�2KK���r�Yݖ8,(7�M΋&�m�����{ZI�ik�N�.�&*��/��,��� �/Dt�AE_�?��T��N9�.�<' ��!�V��s�Uq0�,��jF`[�"_.�p$�B�=���J�_�ia_Z���̽Mi ����+���v�2߭x>�{�5"^��{8(�T��&R^(m��5��9��̪�<P1hT����>��6'O4��6op^9�/�n&.�٫�!O����x	�L��"��L�5�kGɟ �?E\�&�se��'���ܧ���j�w��'d1#�j�[,�K�a��1�A}/K����!+p��䔃f�l����ȣ�gG�������El�$�����!0���M���g���u�-�}��b�jm�y�����(�̴�-C}�؂�/�����24(�@7�66v*{�qܳ=��L���s�N�{�oִW��"ōN���,�\xO�%>z:\    �EXV��|��ܲ��U�P{��0Oc�7nt�Wc����T�w���,OWޒ@l>/Y?��.�3b�-_��=�=նFʙ�m�,b}�	h\[C+��0�B�h���\d0mlNq��73�d�푽���~�����}�5�K�>P���981�<�R�c�)�V��ӯ)Gwx�d&�a��g+}��p������O��j�P�#r�k�BW#�b_����V�u� �p��a� ]��}T�N�~��/��}�Sh�(�8Еn�����ֵ��o"G��)����^����֋i,���K�?��}p'uGI ��GR%�f�Et��{:�3�����1p�l����!7�x�<��.�0�}��s�CE:z�}��� 0����d�v?�Q7V3�\�`�����A�y��:���~�Ȉ,��D�(VB��
�'�?%w|0��C��J�:#:l�B��PX�M=�u�6�ib\�##O��x�q��D�V$��3ϧ	�TO�^��.}l^��=�`L_S�����g�^y�����^��U*���(�7+�[����7�F�B��B�(�B���()�MEId}�����tsL��v����(7� �R�s�M�p9=��w�H����(���9tDz6����Z�G)\�7Z��o��˅g|2���"˙Cb|�<2�%�)c�7���ˣ�FAJ��!mlk��Z�4��*#Ƶu$�*��a�w!⃠��urs�Y��U失��׍+?�)��;�. �N�<`�`���>���	D��S�6:��/�����Q��T30YWF&[����ne]���m��g�����O��ͺ����8��ҧn3y���d�|g�7'�Q����^�]E���>mp��ʣ�g~񒑘��O�=]_'k�EQ���c��$�����>�/��Z[I�6K�ޤd�|;]�7��Us��Ҵŭ�I4�:\RF                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                lд�Ք��}�"������3���A�Dv̹��x>�2�Q���+S���&�6ե2�4I���\�v�����L��ꯅ�FhQ�H3\r�=�c����"�q-���$    �u��Tjmcǻ���*�E�>��w�(���-��F��;x ^hkE�ٺ��03�5������ZS��>��A6N                                                                                                                                Վ��Ce    )�e        "<a�6�f�����    �DFb       �f��*(���    M����pɨ��k   �P��P�Rz                L]|c/���J��<-q�    �V��    E�>�AӲ�e�Ԯ    P��    �M                    ������=          ��        �ա30��            �� ��t��(   ԍ   ��6"z�c-SL9�    �~�
            lU��       ��    �5�%        =d��~_ ��/�    @�"|           �?.    ,r��ł    ,�I�ChԿ&��            r*����\������        �4+ѥ�N        aK�	    ���W�=@r      ��c�#��        $�@��:�           EST    �a<��o        wj�BZ�8<            �Ruḅ�   N��O5�
�        �c��    `ږ-㡅��q�u�c    J�?�    �4��            �$�ȷxq                  �:�
����    q�Z   ��U�Bu� 1        �j.    �QY_    m�U?            3�Ǣ    	���                     �ZQl        ��<B           P�        ����7~�|��    ����8K=           ��f        �>
                 �sx��x    �پ��@}   Z������+        9��   ��
                                     �Zx�    N��&        3�L`    ��M� +8�K�<�{Ė׍��	�@���   �w�c                �PKx                      |�-b    8�OSF�~j�Ɗ.    深      q��G
           َWY�       )J�k;qh�`-
ʘS       �<7�*��r    %��    �h��a      m&n`   � �'�O�8x3h�   �2ȟ    rS����TmΓ   �Ƀ�        U�z��q   	�ʢ?�N�A!^��,nD          ؉           Q��Y��}�HXx[�}   �q��    ��%o��{�$�    ������<   ��M�(?       �4��v1�AGa�JN��:$    ��X5��!����Dxnm@h-a��)�y�p��D��                � �0        ��Ȳ%Sn N�        r���T�؀���    �,�       [�Jt�`��    �)��   )G�&    �'��E�    Y�V	���$�a἟�                   ʪ 3��	   q�{�        �l�����"    ���c�N   ��y��n    �C&�$kQ   J�ek    �W!�           x�^��� t�8tR��n   ���ͼzI           S�� r�uߓɘ    ��P�@    l$+�    ,���zS���[�J��I      	                          q}�)�D         �Z���       �d[        �w]/    � B??9�    ��_�    jԋ    Q�߳b�L�p�ç�~�]���       � ���4-��        8#"6   V��	�b+�    Q�/Y             8���)5�_               Zx�u
           ��p1   	��kj�q��    h�D���x        �r@U���              +��fn�)�wQ��0�    ��6ك⸮               "#c-�*    ����-��           ��/-    ?c�$.��]'���}�A�    ��       a<F�    ����    �e&a   ��$    ��k           �QY�7�)>:۟�lu��   �b�$
   �M�]Ez�#��7��Q{ㆎ�bp�]��7       h2�(]��{k   �p�E�<�H-�   ��� V��      k*�wW�M_LZ�f           )�A�   ����w>
�qg*���ܪ�{8<        	�   � ʭ�4����   :���        S�۱   ��    �14�    ��qx       cD
'zj��         <��{��P@9�k    $�;   J��eCu�      ���k����|�gv�Ys�3   ���)���            ��w\           ���    � �   /�f�            m׭�           K��   �t ��+�A����wgm�{    ������.    �G�    �soq    <�.       u�a�       ��@)k@v<l��       �b                            �[�                                �&�    �_�&        �h]                         �w^g    b��        ����            ��g     2DSN            �  ��J���         2DQ                0��P                       �ۊ�   �*O/        ȵ�M            &E��    MX        ��)�               ��_�    �^ż            ¨�                    vyC�       
       $�q�ҕ��                        D۾�        -��@��        �E�                                                    y���    �Cp�eE
O�J����&�B�&�        �^ʌ    &4��                    ���#                                                                                                                                                                                                                                    2�L�                                                                                                                                                                                                                                                                                                                                                            �%M�                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                               ���                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                            ���                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                            ��W                            �Z�^                                                                       $��                    �o��                                                                        gM�}                                                        *SK]                                                                                                    �=�                                                Wa��                                                                                            ��~�            ��g                                                    �:HT                                                                                        �6�N                            K�                                                                                        ��#�                                                                                           �=;    R"��ñFR    ��ܵa�7���|.E   ˷��z�$��)y    ���12�ޅ�T�=��*"2�;��ܕ@��    y��* w�y    ��Z׫Qi   c���ܛy@�S�   �l�+��"`    �fD
td�;fZ���u�M؏��z��/sW{��!        �B���g�nVp��$=ggHa        �0�}���(���           �+I�   >�Ƿ���K���vԾ�    ܍RձR� 4�A    ,�s    Je[;S�{    wPǿ    < �b}T=�*��P�<����G�n���ޫ�    H��0fj��(�O47�F??s����oB(�   �J(��`P�u.        ���    ��ex���%�C�~K@q�>��Y,���       |��҃`_(����    �"g��x�掠�Ʒ�   G����k�僣�g̐L`u�A    �%&�        �`�3�^�ZR�)�Pٰ5j��x0�   l��>]'��    4���?7]1B��    #U��R�B� }�CE`    +ٽ��X�D�g}J��qXQ�Rh�<�X��טL�@e���i�}Q���   僽/V��    H�������:9Y��~7�?�F�Hg"���fiq,�    k�           /�]6�-��
+�\�%�僵atQX̯�`    �4ɲ    ��]�:E�69�}�'�������X��V�6,qQCG� �B���  P�9*G��lL�e�.��Zf)   ���o�    
x��6s�Bs�
Y    sI�
   y�I�R�	��S����c��,>�V    ��ڙ�b�b�����c���� c����6pSQ@����a�]��    ��`�T�`�5�#��Ov    ͨ��� 5s��W�ɾ    �(��N�Z��       u��x2��n�Y��        6J4d�|=��U�G��]���߼VS����}R�
��:���    }�ݯ�}�y�P��G�w���
        �j�}��F�Ӡ��>��    o�S    �N�$S"�h��K��Ow�!1��L�_��"���s�W�u�q3   �Ƕ��	���?�8�Q�        E��m���        ���    �ݒ��9t��֨t��]���C��=c�<��k{�_&�hS:�|;����޵�m-���Z�<��:�	��oI~�":    5�ۍDjֆ            ~s��r�}���    I{b�&P#���T)l�        ��A�P   ����a�r    �h�q        ��3��F��v*���b�dA#"Z��    l(��@)#s��o��d]CP���SzV��猘8�    ��M��.�>�j�(ù
��{�{�3�Ľ����/�8���Vtm?��	�� đ�q�Kun�t�x{6!��ƾw^l�j���
ʿ���m>�K��մD�.����l^��7��=�$����C��I�b�p�ܒT��@�N��:$�(��L����o2�O�Rx�����8�e��T�֯����c�y�z������]� [G8�/c�G��:�#S������\��0fd����r�n�>^�1zsfly��	�q��jc����|�Ӛ�M.ι�30ˌ�	�Έ�H�����mS֒l
¤�K>���`b�Ww�4�?Z�����{�������b�<2���1�E��z=+�c0��߼�m~\��F�G�gkr#嘻|����{��˺>a��1Ny�XL4�@�~y0�μ2:�\�NPp�C7"O�ӈl�k�����E��5ܾ�;�Tڼb*���(+�w6��:*΋Due�]P�[��=��:k�:�(�f�b��Q�0,��d���uE�ۋ���j��I�?�Ln�Pw�鳇	-R�[!E]#Ӏ�An_�<�z˙RI22%�5;ύa���3���5?[ڏ���%�(&�-e�R�(� h���%Df�}�񺺸�$���P�KA��L]�P�Rh;�ەf�+T���	�N��O�mM�ΰ��@��qcA����V(j&b���j$T�F�W8b��^��l] w�zjk�b����f��%�l�B���̳O�?
�V���}���M/�R�tP��
7^6!�J�����U��Y\�i��9k���k93(�&<"�EhEZ�|n��]s�8�>�ۚH�����'^8�ǧc8�g��񝣁�*8�vĴ�����rZ����]+��B�t����:, Ƿ	u[�e���|&X ��9�T�|Z�T����QY�k�	�=3j�6�;���z��8�#���L���9�U)��?����nE�7?�c8��:��+;�܆�6���E ��x{|�1���2�F̩���?�j�(�*�M��g �������h�V;GC�~�5�[�L��p��P��V���C>sWnt�1>� Ũ_E�a��zK���a6��\-�!�F ��b��+��
yr���p�r�-rk_�µ�ڟ��	G4�8�RT-�����/�-���J{�+F����u��e}���C�)~I�ݎX�z�KϜo���g��h�Z0H��@�'�Bvcҿ$��a��?��gv�̺6�87��G5��Dx��cO�dVG��_��j��;(�Ez��?�i��.���4cyv�P�X��}����W^�gl���)���e��+���֤N�����-+������?o'd�t����!O�b<1��V��Q:�K�RȀ�`�7XV�L'R�&�Ͻ�q����1Վo/���l��ZT��;��d�SS騛m�A����\�
)�q�9)'�5���W#�q��&��ew[ع#��u��-
OfƩK�)c���>�cA���tm�(��Zf^�P�R��H�a��8RE�;l��[�S��u���1� d^���>8��O�8��s�v��͘g�!��m�V��o������9�ۍ��� �n��a�m<���	[��ӳ���62%���s�x���}�M#�XY0u��;.�>��bqR}g���҃��A�y����=��.��2E޺��PQ��j��Z�;	)���]�9�!��OK :��	@[���W!�a�A	�n�þW4�*�d)�m0e�5Cm������D���h0�y�?��8r#���;?`:�����k��6�YI�l��+�� �ܠג� �z��pp�^�_[t�Or?=�P�j3�e�)�(��SΈ�Y�P&+�%���JC�K�k��%����DG�57:������[RKdXpu���I���Fu�Z��x,���U�? m��Ɛu�Ö�w�"�4��t>TU�Uׅg�ő[�����~8/�P1w�6�a����[cչ&&��ZK��{��Z�i*O"Pa�W࿢��� I}�mͨG�bw�ʐ����D���i���q`u 찦����!��F7�!+��p5����4k��֛��U�.k	t�9Ogr�]����F0@��ӻ����'��O7S� ��XupP�?�������ډe�[;��~R��R�I2U��Y����[�*Lp�A�j�A'�`T�@�ֲ(Z�Ֆ}��&�d��߹����t��q�Cg]��w���'R�_]�&�$�o{�I�F��дR�9����غ~�
g*�S`�شo[������1��1$����>�L�L����Zz��^��n�0?oy%]��q�J�}2�E�K>����4��Ɗ��4F}��=mx�9��jVzK�T@�gSW�E�^p�E���a�h8N@y�IyC5�1�-�ѱ�wjހ �į��h����2���,B�g��)����!��RhשU�1�g��O�6�dq���.��\g�
��182�H�����h�P�����h���]�JWl�RKdc�( ; ���z��x�R�����^_s<e3{����TP�Ήc}�0^0���سwp����J{J?�-��nc���O�a]x
�ȿlL��eŬ���C �I�>èS�����YVR�D�ٹײB�x�Ƹ�ț����{�F��`7�a�ʚ�4�3�\���;#.%y��*�jIE:���ey�KCt�{6�!y��,�`��U���&�nz
�����)������ ȓ�]	0��椠��"dG!=�l�� �~�h���@�����k�C�tp�+_ ���&� �#}��w����BN��U���H���xV:c����S<��A lOj����Uf�Ħ>��.�xSދ,4�_��6)�������=��fm��ڳ�{~��ܯ4鯃�bu��9ʐ+�zś]qa^�${��`��\_r麙lj�#'��O[��]��x�ޜ� ���.�ס���
:���^��9Jw(a{v�����q�&-$��R��ܧ|5L�~p�If	��/�5614�G�<�[�2h!�*ј)�ĝ��r��][8����I����tѢW���Ѻ�ŋNe�m��r�M����Ye
+⤼^D8&��/�b};�_-��ǘ��T{<����!�!22)vY���t9�.0����{-R���{��rť�w��Z#~tLY6EJW<����!ҍ��x�g��	5Q�'8��-����-�GWɃq�J]��:͔+ҥ~�f�ڊE�c��<=��c,KvE��W���V}�H���8�f=�L��G��n�Ͽ�_s,!e���쬅��V%;Ya�l�jc<��3wݠCQ�R�+�ȉ�j{h�[���#N���)Rl�$,Ͽȧ���j�~�-bz�;�x�k�D�F�[��j��_�6�Ust@&l#��S~a�"[�`��~5�A�W�'�F��ϴ!)�{Q����D�%��ߘ�S6����O
���WH}4��V��<�keT���H,���}ٛ'-��8�5�D�҂sU �e.��&h;u��@����.�<�c���.��[R��C�O�Cح{�Hf�K�l�^�+m��͵���2KO�'�hi>��n�/�J�_kH#���6�?f�v&֫#���Yҽ�&5V��#��c�9���4�20R�`��:��./��*�-��p�[<��_L�����+G溰<�E��-��#RtP�	�����mQY�珒?RFU_��z�$�?q�Y	�2!����R��,�j���PVbk����d	�=K�r���CQ>OA��6N�H�CPtQ�P��w�4�[U�>.T��~����g�GYEI��(J�:����n�D?7�`�t!�5_�I
��Ϋ�/�&U��XvKC2)L��̕�q�S�utGN�3i�n�f�d4;��NҖ�.\Uct���'��^�cO�+�m�m�:�rT$��h�a'�,oͷ�B峴�9o�9ǰ��?�P�;PR��t�p�iCh���C�����k����:��^ˣ�V��L�0c^���|��O�����M�i�E�^���*�q��u��X����z:�q�a��O�p�i�E\}	P��_��v�3��O5����\DߴDy�ڽԇ�):P��&�4�R)mLaO<�=�}kP���,TTm⃹    �  �   E   
              �Y��qԑ�v/�yG��-�Ҩ�ٍ53�RDz95�>��|���?                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                $�^Cg���N��`�S��A�FgL]�����x�<��BǍPV�~��h�V�n�8ֆ�6��J�]O��o*����En��M ~�BuX"���!e	R3����z&)~�8���9���t��7��kOcJ�Я�bg����#f��?x%10d        |�7�d��[ ���W�    �B���=��4m�� �Hn�w4���,B�|'���?����s����fg�o݈Mx��N�	J�s�pY�	VN(Iq� �uo[r�G�l��$|���/U�5V���@��c/8�z�����I��9�T�/�@��,�s�=*T��g��p�;��0M��->�-�u�Ԓ`�O�FD�ƚ�b�F�.��#e�8��Ar8#xS�Z��]��H�
����ɞk��n����G�������k�e���i��YT�o�4�Q���!��M�nW��`ĐCk\���ȹ�G�IHà�C�7�D�����T�T>���2""G��z�Ob]�xO ����{C�q��[_Iny�V�> X9�o�Q�;\ᑁOFյ �9.�i���$ 
���~E�GY)x�E��S��cF\���uڃO$~�[�P��W�pY�ݿI�*�F�!�t��.���j�eZ�`�[�
�������b� Q��-	��x4/�b�Ypu�ξ�h�DS�h���u�-����[&mL�f�{@
O��;�`�ӭ������8�,Bo����t!I!��t�[)�4�!�}$��� �է�����O��Hs6ѩ-��-�e�6����ɯo��w�jXm��J~1.h/��͗���H���|��+�lf�a�n����E2 N/���![�ۛ�k��q�y�φdPu�N�ԁ��N�U�Պ1W5�=.4J�h��Z;��ݧE�0Ff�3j��������+�Q�d,v�(3t�}�=,�a$N�Qi���~!��e����f��fs P�����5�*�&#6��Y��#�n��n�f��(KVxZ�������}�1���1D9�G���;C��G�K��>��ѻ��`����^�U�*He�ޕ�s.����@�÷�3~?@�C6�Q!�$x\�&��,z������C�ڰH��)Z�'���PJ���y���u_����[ѭ�+�Q託�7�w�b���W�.��d��u�2��#�b)o�P,��*L����u:��޴�����H���h��!�.-\��U"�,rU*3h�ʪ��3�+�B֐6脕�l1�}I�F1WU+	�mm�C6V��(O!��G����hQ�!�e^@��X�	�[Q�v��>2��1��(;���U�T5ч�d������A����Kc�M��&ĉ��"����������U`�B^\Ze����O&�̋����r؉�T�р��f��u&���6�|:�jd�U$��1�?�V��6�������6s��H���Y΄���nc�$�ttKW���5���j��T
�s�ˍГ���1���b׷�5D��wMZ�n��M�.�d�f:M��A���Д�����B�$���3_�ΛW����)jڒ�	����p��0�vl�,+i~ԑ6��5�;��є��\�|�@ґʇ9�>��.}�.���+�'�ׯ���j$�����x�m.t>N����湷%OiT��:�Ig`���Q��Z}_��lГ�]BK��/ޮ}��w`���B���ADIоA�ʮ5��5x݈�դq���2~�}�����4�Jl_xI��c׹��ߜ�fk�R�)�ބ�����2�I9Z ��X'5�����K�f�)��&Ӄ#� B*�����%�t���B��PXM,��c1��n��D�)��J�rA)۸�ǹ�3u�3�����#f�S|L�\F��>��s��\�G��1�bK��˿m��&q�� �Y�Nd#2�Nj�������Y�X���Mt(ܶ
��)�ǘ��0�Orxn5L̗y�?��m�Q,��y�hr%R�ל�?]�N��@]��ڿ�ׄm(��z6>!6kTkE��w��$kh\Uo0f�X�,M��ͭ �Ts�������z]�x���f�����G�_-���-��sg���;��A�6�c�˅�yPj>��Q��0Hܼ���Ly�ѝ8)�ٙ�F�����7BÓ��M�� `���
���0}�Zj9�F�k(��#F�h����$��Q6�����J�s*�=@� FB�9IQZ���1h)����@��ή7{�&~�\:�\��}��g�L�+���XC��ם�74(RYN�2sϷy��?�)����b�HK��ǵ�I�o��%�Ŀ��͜�����������k��<)`Râ��OAd\	��ǋ�H�6l�L�m�
�<�2z��7z���nl|��N{��J$>���T���g)C��
�0���|��8�b�AZ��×����Ǚ���e�b�k���6��pJ$�o�D��%q�g�f0泜.�\�.�Pn�Ψ��5�R{��@Gnы��T���x�Ѵ ϊ���ʢ��Bb����;/�}Cq�1����#@%{ R�bg]�ŏ�>�3�_.��#@e!S��j_�����Qs�t�9g�؄����ُI�3�=�h��r�Ѝ��p���k�!S�������d��a�ᐷ9��?���C�K~j[�#@Frh�.���1ߵU�p���nӒ�zo��O��a�=
������F�4e&gU�ԖD���/r?��-`cZY,�?.�� =����fY=s-_;��^V#4hC�Ԇ\8��VRVmWض��U׸Dw'���>�L�U����34�����oh�ʻ���\ �%����h	��Ղ.Oj�ޮ��&S�z�g�Ʊ�톕>��� ����c&L��&S��1';�)��!�p����
�������:�f�/쁷��x8a�"���yy}��i�P�C��A���L����ʚ��}p�o�~�:�'��R�����,v�-�4�V����,BaܛK��¤*ޥ</�����3U��w&�':��QҰi��_�F����Z��[����$	�>q�0���_���6��LW�nk!Em�Y�!�߉�P�^AGbT�ܸf��������q$��{���r�"��q=PAz���%��>hV���"t/_#�l���{G�M�m� ���'��]rb�߂K�T�y��������t)�	�f�1e-�%�(�����=��r�)u�2*I���\q��7̪��:�}KlRqM<�;�S�j��"�x����frZ���M��:���{Rw��$GWP�O>��<z�F.�SAI(%/�-�jD���4��v%@�������e|H�7���)[�Q����'ഞ|�c9
�}ų1|;RXf��_^'�'��}B7�����H��$���B�=�����Pi��;�9��?"e���aV��o<�D�O4�Ε�N�u)O����r4pN�.V�7'W��ܧ��o�%��cq�p���I��U�Ħ.�S	���&��=���rծ�:���\'�}t��1��r�I)�Ce�!���IU��&�g��l�ܳ��=�"^hq�@���n��p�ަhu��������%��;�8�����k��_F�s��o�̈� [P�#�V\�1�I�Цs�����&��LB�@��f����\C�CG�D��a��~n�ihN��E�w��^b���5.�.���9��x >L��q�.�kj���:��I�tN2Fύ�L�T��>N��vv��1�0�f���j�c��$�.jH_N��/�9���g��ɲ��u �"�֯����K��WȆ���W�I���ʶ<�C7@濸��b�۶q�)���F���-ӡyƟ��Ѿ�`�i�yE|`9��ɮ&Ƒ�§T�1�BP�����GO#�ց�Z����z{�D�:;�D8� ������X$�<�N�8?��V�|]'�,�d�o��4��u�)6\�Q�o��a=��(�|Lu����m�&������ӮGnS����..�XYbI��3��R��<>FՇ�{ϸ�5J��=p��d��ya5�h�n�#��gc�¢Ř�=i�a��]7�Kb��&��� �>_��&l�h�n#��T�f�b"���9�}�1��m<�I7����BC`l���"��P�O�ؚC�<�a�TO1	
Ō��{�ZA�$U��9m�@IV��,����i>rŦy��M^�ih//�'<H�����G��2Ӫ���b��{���o���rLj��D@x�s���r .W38U�H�P��S�Ӭ:fqrwX�p���ϣӝ#Dр+�14�{��Q�ղ0�V q�ݹ�!�k2��1q��0L�SO}��,�%�f�Z_+?Ct3���O��@�� y�Z��N#�4�$��="qx���̚Pf	ȩ���.�c����=,LE��1�W�I!�}d�n.%�5w��y��LJnS4��+���ç0�[=�O\ٵY0��h;��;�a�FC"D���y�5�!mWu��[���u��,�?Q���d��2xX�]vyR&�6�Ҭk��@���v7�q�\`�S�+�*����培�����9hx���O����]]���[��ǦK? %8�x)C���6,��#4~-���2j @��L_V��엹', �y�v���rEO�gB��f�>L�J��$3���k��RJ�w���%��F��Y��v�ہ�����(v��˽G�h+!�w��f}��1蠗 ���8ںw0��0B��Ue٬��'Y#��<�ٞ4����Dj��I8�jSE1���ckT$�Ǡ_v̻�~'*-�ܲ�6U����q-:�^̦#���8`�G���m��'1�����]4�fGK�Zs��*d�Ƒ?�ͷV��J���[#��XQE�vبd�p�m���k�]bۢ&q�3(ђ�uژ)Ҳ�J}�&��o��'��&�k���n\�������<������a\],���']r/�q�C,g�$��4&a_"�<B�U?2�V���°�)��e�A�����w���=�]���%��W��0�b�G�O���&É��$���lիzL�vg7�#�,��H�8�'���;t�K����"q�z4��B+�?D���g�p%�������%bּ� �����PV_��6#?��� �;-3n����p	���i�sN����HQ�#��d�P�N�,�B�P-���%�.A6��(s���{���O�l�E�4W�FL��M�mE0�?V?�U+�x|��Z��4Q���YP�F�N7�dA���o�=�^��q�lG{���2����s����	e�./�=>T��cN���U I��H@b���#w+��V�q�n\Dk�)��3�&��G��ή�@��O�����-.��Ƒ{1A"��c�W�>%���VQ�ݐ��a��$��i�X �Hb��Ǽ��S���-�x8(B�KC� �m/��i�y�2������������>��V���$�.OJ�Y���XBJ��.��%F�㤰EZLXx�`MO������ؘ�oK�r�o�e���T~&� ����P2�*�����-m�����A"����_��w����D�m�v$�`�޳c+�(�(�S��%�f���y0vZ����<Z ���_(�[rҝj�{4� ��<�	mL�HGL�P,"VA=g%&-z������V��Zf ���c�
D���o��B���1a4�d\�m�S��W�F|��B�*}�E.5����۱�t�Ke��o�Yx��8��o$���y��)��M���o)���i��=�Z0N��T�KI"Oc�>��A;��d{'}���-.*j�d�	y�s6�mg���i�P�qL�hg�=�:p#���&��>��DD���~�0����p�p�غr61���Bl���H*72\n���(eL�C���!4�Ԑ�u׿��s�x�)�����#:}p&�'&�l�	�%�R��(6H��{�ћe���4���hՕ\�n�h����D�C�j��60z�M}������+vf��O�	�bcL4��p'J��jvr�w6-т�ΐ�t|�T}�������lK�<��q���n��@Ս��x���A-��/_��Tx��,�m�&���4:
�K�Ae� �Q|H�3���o��� ܬ�nNc�3�"2��4!Eay|�~��GVF�3�Z���&�˚���)��GPE�A�����,� ���T���W�;�s����
Ӿ;U���	g�-?ݦR���b�j�ԙ1k�i���^pmv�~y����K��\p�c
6��)W횰 ���O>	ў��=rns+&�l$�T�@��I�<`�%kim�и"�R��)��]ܢ���u_:��o����Q�gD�ot�ǡ����--�5��X���U���ĹyJUӅ[�6��})�#C�lAk��f�5w9/� ÿ�=��Qs<���tX�f\[R^a�1_��ܳ	j��C1�c�%g8���.������`'��FCxS#�;k���/L��&>4�JE���>�Ӏ�3,�[�}hz����,F�g�U����mL00����_���ki��e$߻g����.h��WT��y�2\���H��I�C�s���Ђ)*���b��
�M
�Mm��P��N�2j9�w�-�m6v�3�g�ܼ�'gفL���_g�Ib�l�ȿH#��NpŻ00֜9y��n�z��DÅ�N�T<�����9�_��Ҙ!s�_&�#��b���ZD@��'�x��J՝�-�rHB��dFr{]��6e:�W�yd����a����\���_�<K��m;T��<���s��*q753����心��1�F�#p�[K�&t��+ �i/2S0/��t�-�xkh�v7
Z?p�ŝ8E=����,�dҗ��N����_6��7�s(a���m�!��s�u�P,���e�d��v��v�.)�{DVq��j=՚�N/��A6�@��֧aԓ@01I㬆_g���'�;�|nb'�$�����C	+�1n�'CH;1�9��� V�=�I[�ͷՁ�LZ8�W�w��%V.[z�χA}>���JH�g��]���1y䖶����A��M�9�?��+h�͢M*���
�G���A���zI��|�h8�1�ׅ�%i��ȕ�3*� �y�PA��[t
�)�+d�_�kA�LRMޮ\[+V�z]��;�ȃ@3���oCa��(:m�5 ��Qu��/L��T�;�,�~�'�2,��}=l�.ݛq-��+�r#Vu'��JU}^����k�ݫH�JpD�!�8�^�A;�?�hZ�V�MX���v!Fa%4�(FI��8a������*���ϱ�X$6v�l`@�+��N�����V�2Y�DD��%�M+�&�PE7���v�r�4KN��("��Pk�)vH�[������.	�` �NX�|�'9+Zx�SWN7bwq�����/<��L[��K|�]B'�Ԫy#ǣ)�9��`��M`xKn��7����5]�$���M�a�7���"S�u��!DV0��|�T(�Ee�Q��.:|�x�[��0��f����]$�͇���E�SnH��ت!�G�	�Y���{1��T`��WJ:��L�x�NG���[K�O�D�:)�=xW
��R�-o� �}���R2��7j�x�
�;7W����WB1�H��g�fq����w#c*H{<��"u�1��������?���O����y����n�U�}�{��Dpb���ڬ��W@g[(	K���D��tP7��������]���ľ�S�N�,��=��
�z `p���ٳZ�گ1�?��i˰�����Eb��``+��Ȱz�
!��	��Wl�xJ����<�JD�'q�e����ՠ���b�Z3yS��v���k��?��tG"�#qh���EC2·b�RRC�{�^ҲQ�re�Q���>s��O� �Z�o�����K�G ��-y�8P��Y��2�80��b�̖XL�������2�4uU.6��Wb�J�G2��-b%�OǇ�P�O�����wPCO�fX��O�"�^�k����[PCl��^�c�MX��'���`T[��pNW��D�]�G�*S�s�5,��W�>�W��넼r7z���!��i�ɬ(��<Ď�m7±V�CD<�#R/��-�4�NV
MϜm���=m������z
�}
�JT�9��@���PKAh5Dk���;*��麯�:P���7����_�Mb���C߉o����N+�:����&�R2%Lx�a������V���h������hN���CBNw�[�|�[��Ý�raP�%�OF�ަq$?�q04�4V�[>�4�����-Wn�_(����v��U �Y�]X��Ⱥ[�	���O��06��D>Y|��JQ���%�j�A�;�ϵ�WT�Cy���}VjQr��Y-� ��1��c�P!7w�!'�{p4w=V8��^����*�z'����%��゛�'��tx#�r�m�GYJ�ӯ�+��#��h<�|a�<o��I��>�IT].���:��]D�X�_�A�b�A���lFLc��QC�*ci�$�N<j�۽���d0�X�(�7s?Km��/��;�e5��ҕV6;�*��*�+���G��=U{��|��F � r�?ف#��`R�� �@�����~`H�������9I.��;�`6�-�j�?��˹\��v���O��o b� _@a�@i=puc^����Ը�-��'v>H+&^�j��`��5q����p�Q�<���]�u���tNѥ0G�ϝ/�X�V%��?`� ��2�n��P��뒱����T=�;#~���pWyv���9��S��Nją*QBi���!�oAa�=ZU�F|�����zb��-) pUe��jK����'�4��@��Nw�%g4A��B;5���DH��n�l�am���������ׂ������x2��*���F�7�3!�F+A�׀�>9YS>��w�L�^2g�s ��D���{�J^m��6�b����ڵ�T�;�S'�/(���a�Zi���a�%�v�)�Z���q~Yt��WϟVRG��}N*97Sć뼪����ҩ�/f����Z@x������v��T����G/.s��K�UXܗ2�����ͯ(&_8[������q_ɨ�>���ԩ��g�#�d��GS�V���8l�|��$�ܷ�
�����VX�d�{<D�]��������4��?or=CY\V�C�mVD�񡍱ީ�fN�1Ec\��#��1��ALȱ�{���][FG'E�Qc��r`4���z7~7�,u�b�T�_c�Ƅ��ڱ�\ҩ��,�\�z��+�-�rƜ`t��Y?% �;.a%8,�ϣgo�T$ujQ��f٣)UY�v�:���q�5��jt��g�!����~�%!�Aݩ�L���3�LnXgMzY�ś�jd1��t�m .{o�"i7:T�\���_�]���{�M]E�3<2/�)]�:h��~ ��$�*�G�7�(�$�T ���O>�L8<iQ3�E.��9���t�|��a�~LR��&�֍����B��ꮬ^�eeE
P�e���xR�ղT�^��pe~�k���r�$Ͻ��h�~��ܽSE�ŕ���y�@b�WLs�������@_�T�O)-S
/�����&Һ1F���?d�2 0#q��� ��iZ�A^�A�2N��	 Yl�@�<4'T���Gb ыZ�*
��z����͞Tw��h��oW���WBz��&��n�Z��Ab>�A��~Ӥ�d�S�@��F�(I��&G�3�}&%��75	褩��3�;l���������f|�Y]JD�I�ʘ��C�$ʌ��ޤ�>p��������D� "���L�`�ba��A}a,��M�N)><����O{��C�j���)AE����Y�����'drY�&QK����3�����<���Ȝ�]�I��,>=�ML�u��n�a(q��Yy�B��fD�v	�gjH*���
no~��9"�"�A��/�B�O$#,ڂ�����@^���`D�N�\m�&u�/�X������n���w�۾#��6),�#k�G�U�S�W���y�SXK�/fľa��aE���J���zZ����4BX��I��D�S*�Qp��PTҝI�5{ܐ�@�;j/pӬ~���e��ŜJ�\̠m�]��7��{#�f��&҇y�[[B�π��9Hrz���/�W N��u�sJ9V\��P��B��lGŦ���Ԭ�D%sL�_O�H�?��gB5@5����3��$���_���^Tj3뤙?U�Hiooy׀�A��1� w�G�.�&�7�tx��j�I�¥�yq������I㔣�X�Դn�%@s�p2v��9Dh6"^���&�&6)Z峦�,˂��ʹ��m\�0RNj ��E���Þߋ�Oc�1Ɣ���v<�6��M]@$@o�S����7Yl��q�r�y�����5�'i��r�4�lc��{u������t�,n�Tp�&�L�I��JF�e����j�u�Rg���b�0���},� 8i�mc�^vfF��A>�p�Np��q�w uOj�O\E#�{�ѹ���rIPg�Y�7�J��U��( 0�h�f��hdA]�5Fw��H�a�l�[C�@����	�Yy����i�d���Ui��ĥ?o�q�����X��4� \> �##�]/�>q�Pi���(�܂����iv�%	�xB-��|���5w�%�;ҡ�Uj�[�b��0�
��8�`�V��/��!|T@bw*N*��:�Z�Ͽ�E��p���A����������X'C
�d���V�$wvu-k��m��\-�|ag��edC����px��نҟ�no�0�U�H��$�����3�7�`IϨ�WW���%cobXi�!�kH�/��᰸]��>��n?<W��E�gN蓢X�N4�/I�WU��T���W���q�VAa�"0YX#�D��8�]#��և|�+�K����t��
�_W�O�	�ɯ�sÿ��N\�͎q��ewyӶt�sK&�ԓ��Fl���D�c�@��v���ANA���M�=��+��|��=jz�q5wdJ�0�d9�����ï��A^�q�:$3|�ߟ���*'����\�L���@�\��JӉO
D�[���FCÒ$W=�S�_���)���ځ�w@z�ӎ�
�r7�W�5��T����_d�L��=K82n��L��G�_>���R��8~���]��ޱw�3ԓ�je�g���$��-�@���z6s�e-��C]	 � R����@]`�� ���;&��v��`b��ƍ5ȃ�U!���V�b%�\��:vc�H��Y�Y��L)��>�Ҝ*J�@P/�} d�l���7�Au�:����M��ȷ�z�����_���t�Z�k �5�l�q]���̨0N��8X�!ЗD+db��-t�'��E]��O�~Z@��xa���������{�'%�1M���G��@f@�9(�!��7ntvm�X��6?>pF[�)x�Π>̭[ʦ{u��R>����0�)Q��3@�\FiaB'S.��C	�?��X�S|�!y�<VU���]���LL��Tz�/��uVؖ���e���
(����i��9����Rj3�"��ߴ���U[+�� ~��Hu������<pQ���D��?h9Z/�Η���K����Nz��`'sH�
'�wj)=`G 4�xbŉv�Y�=1���l��/3U��I�v���j�Uq����X����LF�F]t+�{��f�~�r�p[���@GZ��[үe�}*���(�����v���3�P��C1V(BC6�?�S�X�[m�a�6(� ���|�n�k5 �^H�m���H�y��s>�ՙ�dBt�(��K���í;3N&��NM
%�W��`����8�Y�&�I�]��c����#b�̽8���%��M@�ּDl�W���xO5��@�:Ae��h���_�k�pU�@ä�>�V�X++�2�)�E��i�T���;�H�>u3�Jդ��W��b�I���x�V���F��f.�,*��uo8򋓹o��v�qGG�H�q}R��jK����b�����K�W��{�:*g��bl`�xN�-N��` ��(�0��L�#p|��<k�pj8}�~p�n�&e�Ϧ�L�㕐I�ީE�Ay�.;�A�ښ<�*aQ���$:V]'~�W����NgB��`n��|�Iii�+���O<�R��hu�����{�`02Zz=�A�w%Mk��`AR�EgV]c�˞�����w�H&~L�j	ߎS���l��쀴��Kqj�ڑ5��ً�ܕ*���f^"[���"�h��X"xT�0�T�6�:����
)���:5���
�}Q�҄��@}e��|L�]�����]��� �n�Y�����|]�� �\�Ӄwï y����_Hs�p��iF&@�.����[ms�D)�����*!�|��W���KZ�6J��/�5�k<�8X���-0���V�5�Ee�z_�I1�)�W|Lm&��]"����&q�K#�[J�򞙥�E�vے�/m��#&�L��9hj���MA� ��<ƪ|9qv�(����L�m�Z�j�pn-�����'<�+���3D�����Cy�UQ�X�o�74�	��,��Y4;}�V#���VꮮV�˩1@�u���2˙�z�-����;ԝ*;:`��Ӑq�Ԇ<|��ڈ���ȍ'S�"�~�H� ��|X-�:i�V�J����M�s��|S�����pc��nބ������o�� �{�|�4V���PoYڅ��ݕK�}�ܝB\�@�XW��I/J����g���2��*}��@��8��n���X=�uFX�i�l58N���o��-%T_�c��S1r�_�K��0�W�O̽��I���G�`�Gg~�o�����E��x��5�D���0�6j��'[Ӹ��^y�|����7��^°z��A*���b��٭��~(&6���!S���qb�W~Q�WɶOm��O[�n����{�R�J)7EK��T?��L�|ԚK�'��"�qC��ՋW�ŭVu�����	����0�[��~#ݲ�!�WY�T}q}�ܒ��ъ���K�^�H\�8 OG�ܦ��0F>I��F"Yl�3Ȃ�5cL�`s�P/^0zt��>^4�[��?�WlN\I�:0�2�é��GꪢI�}�-@���l��@����}������vR����Bu��Ȳz�$��'��
m�p�"�KC=v�XȒ|���/'f�@ݲC������H$ ���y�pb!����Y5�WCoR:8W��F,DT9��y���9@#�h+��b'BA0Ϛ��1�2XVqF`��r����LaX��
)RN�|�=�~����
��
4���鍓\�yE��˸B��C����q?�s���<u�������6ٕ��JE�����2	h�=���Տ�W�����Ѷ���b��A+��&�abX�vE��j��q� �P_�E��Ɛa6=�����#L���]���1x6QW跞֟ԣ���؝��Kk`>�sz�d��)}�{�ݳsi_0�������K�+݊��%������9oz)Y>�"K)��y�b��2.��|�tQ	-%hU޺C��Z�(ǐ�/=�t�仛�P&=!�}�2���a6�F{�6�[]q��,�X�/���d6Q�4�Ku3��BD��'s�u{٥}����z�|ԐJO{��L<��(��{��*�pH9r�y�y|�����p���6�{�g�Q'������h$�����^
.�����Wũ���q�]#� �6�<N�ਵ��	C��O��V�Α��0�Y�PV�rAnhZK �э�_U���
����X��7��qug�vDa�k5p{;���E� z���Ɗ��+�Q�HS�_Xbt���!�\��Y��_γ�R	V��nT�)tz�2!��Ϻ��C��횾8Sg����8\+�֜�DN���Q�Q:Yo���B� ��#�P䭄+ڨ��"��-���z�HOM��b�W�l�r��N��o��<lX#"-,?ڿ��>@2_��~����Ve��owk�yݩ�~�)�G�]&��b�I�M��Q��n���̓E(���%�N�<H��D?�g�]�Ԭ�T���5��:zv�}纐ͤ��j�����
+ϗz���Y��\��3��ҮAF���.[C:�U�3��⾏�\:�ɖsp#� �V.��֫aҞ%�|��^K������e�/A*��Y{Z}<�t/���"�HI`��~��y���ESh�?�/�O�Y��G�s�CY��劐ɵ�!^�H��v -��=zAYϋ�$�2�8�kyqZ�ѝr��DfZf=i���(�"v���_������u]Ko{`�K�;x��o]-�R����]�!9��T�5u����؈��5��'�0�[9�-�W��*�mw�q:�������*�˻
-����R�����f�8�rh�d��W���k��2��Ei�Q���p�tLv�kJ�V��Q�7�;O\��Zѝ�؃�� ;�MC.:�y	�@XNwp��n�'0	�".�t,��u��r)�Ǿ�y��
_c�� ̽>	4�$�i)8ւ^ �4t)O���My��fI��u��0^��­K�ABq.ޟt��}��y����@^��Xc��Y�Q��&��W�X���������ї� Eø��
y�x{#�W�-�Q}�K���!���UA0�Cz���iX�s����]y�T��ᣥ o����x��5���~3�Q�	�W�f;"S����{��Y��wo+�ůp������	�p���8D��3>W��i�d��DY�Y�$c�����a
�v�C������[���!�Pz�xY& ���P���&�|�������>�f���l�����(�>�cТ��i�^�� ZBy�|�C90�pZ�٤������<��	��Xp)��`�v�շCt`g�X�V$�+a���H���MO=�q�+��M�a_�Y��y!�.Av��0m d��:���%���m��X��K�,ь;�~��ZQ��)_DG�� +�*rO�tQ��w�;T�k����/�D;��\2`;��h�����T(f�ӗ�~��"UaPS9���ܱ���r�r�=�<	�a�̡8�qA�t��yu�/?.�[�+yg`-{i���F�]ɣZ���Ln��ƿ�ق��2��u�@e������X������uovr:L�4XNk~�'@T����;��*�f=�+�B���h�� �[̹^��H���}!|K��:��^���+���P���`��"��'�{7�����`���R�5��H���R�pl?�@��7+���w�0�|o����p��u�q4V�K�U��
�R&O�*#�b�Q�P��p�R%G�.��*Et�x3� ��$)��.�d$�H�,�D�f�!��#)k	����LlHp��2��=�j #���[Cc8���T��G�zpѼ8�>�r�҂4�����+rJ�c�g殳Jy�l�/<3$����,T9��5Ay���xHh�as��s��:*�-K	+C�F��t�0F�V�@�������n��uף�h��!h:vO@U�ma���'��@*V�*�?�N*b\U}om�H����Q��/5i��[T��1����{Ċ���VN:|���d+��߷�-ʨπi��5�v�|x_S��ZF�ϣ�]y���zjzVŪ�E�n\��N�,���aU=�+�q��⩏�p�"����c��@���H���p]q����?+�7���1�j�J�$����*�{�31�H��8�G���a�I^�Oa`��`�1e(����3������g��L�h^�T�eN� R;����-���� l��7����M��	L%C�T6P#�7����*a�a�jS�*M��,-�.�y����΢�0�V���y�j���caQ�S��,!تnQ��Jב?_H؈���]�N�u�8��k�OlP�S��)�퓗�"t�9�JB�jnJzH�3u��������&���g<D�P��7�x�}�v,���M��<]u�*�.���	1�_�ȝle��d��?}6�tؓ��@=$�����(��xbk�Eq_�:�%WbvI����Q+4D�tI/��;G�2QA�|ri\�ĳ����:Q�<�O�ǽ�ڀ5�%�����^��*�<��Kew�[�D���=���0�qv�՘�gل�.��	����Z�k�rߊ���~+�ae���I�W����<�;_���]+2kٓ�B��*~�R"�z�r����>��kZ�3c�
��*��Ι)�$7DG����:���*8��������Ȝ�������'7@���U�\�tQ$��e\zUeB��>�c��!'�Q�0��Co�wDH9(6��u)+��^�=e��v9�MM����H2�b�&�v���eo}����zQvjL>�>���.m�6��B�W=k]8{��;�OРv� �[��l�+�6�5�uv��y,xT����5�%+�|>�*h}�@�0����28}+�1d����U���}�2��i<�dS����G����؄�xt�L�E��1S�7�5t�6�:�9���7�V����=�UH�m'�I���M@��b��ׁ<��Z@�3�C)8\MA�PK�y����ު�i(�<σ�`�q��� 56�����/`��H��ȕKU�s�m��嗲L�.=,4&6,^�)o-G��~eG����s����hX�gә��)O��1�I�@u�����]������i�K�|�k]�jaZ�n>�#��̕���Y���@[ޤ��@V�ZLpў~�}�O��[��y�m��cxp@�hfά� ��F�����G"�x[Ҭ~���xs�v	�
�y��&���J�[�?x-cp���Y4ze��NYP�hA�{��y�/E�M	SM��-]˨F�@S��
%i+x2Ú,P͊X��-/���OB�뽌X�ch&C�V�
(B�b"�-0� ,�8V�.�,E�~X�r��rotH~%G�P̣���q#[()��}�2����hSzY_�C�/V�-�<L�ן��V�rt�#�7o♩U;1�o��D�7�P��4��o��<�=Ӯ�g��)d{A%p�/�W�$�M2�9�w�3��b����R�4���,[�	x6L�^Y�ժ��5t���I����R搟�L��2rt�e�:��������������퉨�N�f|K�|��&�i�1�O]������ϰ� �)	M�|��-���u�e���sQ��$��prt�.��|(j)��Mn�,'n��|�f�����ұ�S~]^�T�A��*�t���i#f���R\�b1�,AQ�N�������m��S�,l���C'f+l�4'*�jRn�e	<!L<��� �Ȗ} ZB��:���{��9�[΂��c���b��%�xL���fL���|��o���2�J2·���Q.�z��6�6'QnM8��a�C7)Qx����@�hJ�o���kx&��?�8=�u~<d~���z�y���k�.�n�mR8>�G��zRܢx��1�CXn�wk�7�=�����#��ƽ�6���ԗ�u�Z����>!:v]q+"��g���%80�beL���%����+�{y\��zPB�Έ�¡2�t-���^U��U�/�9���ٷ�4�۱�r��o�N�*�k^O=bY ��QA�.x�*�ݨ)"mtQ,���n��8+rEĈ��EE�1on�xF2y-����4� ��Zc��^�+�z(�u<9�TԽ� 1l�a�ٷA������-{�v�?#gY�e�Y���L���I�=�O�dTl��_)��ձ ���	.5�8��ߍYyd�Wv�G�*�ӌ�+����,���7�@��kH_{j�k�n���n���x�.�y�����^G��3�� "&j�n�D�=61�1 �{r����bD���ԉ���-�E�����?ײd���75n��K/o)G}��ӯ(�s2)@G�qs�%��鞻�.]�2;
���G�� a@�@�\b�3�.14�g�E�d���5�<fl�Ji��yA���3�Gj[�R�G~f����0�XB$J���Q^���Wx\�ν��\J�FO�Dw����@3s�o���jꀪi�u����x7\�tEE��y����t4�����ro�ʎ,,��H�������P���T�0�4/�A�8�o�dq1�������f��Q��C�i0�v�}/v:���Eա��#���AB�D$#`os@O!EG�[7�
2�L:���؜&5,7����6��V8���)3t3���` �Z4��Z^x��R�k�������,�qj֐�D[%Z�oJ~9-jj�¹,�fh�G/cL�����2�'����^Pc0�dR��}���^#�1��n8�.�1ڣ����Z�^P� �I�(��sm���t�l���m�?f݊8z%�;8W�_0N-9���1p1>�jt]��F��^�O�9�ĴN˪��`���]��0����į�c4���,�0��fִ��T��[�ӑ�ul�Q'b�ԓw�f����3�O�E�0?����/�*l�s�n�������]��}y�N��
�ОPR��)�O</;���v��<R�&�$n�ĸW<��w�����^���-���u�Q���Σf��:"a-B������Q}.Fԡ�o��P��M�y7�ø��p�����}�s�?�2�JN� K���(�к�K�A �{��R,a5_4触j�?/����J@�W��5�,��2�4���ʧB.���8z����M�z:rϬ9��K`�����&$���}�%b�,���VÂ��,�1%��x�!�XQ}���B�N�����(��`����.��V(����ko�Ĵw߁�~�
*O|[�d��f��k�I{▏�@��>����|ȇ`m��(�����W>��  ���G�Q����zH�[��p�(��L�.�j]��PSi����j4i�6�Rq��	��"?�s�'�Fz+6�[![9����WY��E��u�	$�����2��P�4�n�(�	*Ű&$7����+�p���������T�/�P�'�����	h�����2�+\�L)P�K�t������3z�זu�����_���x��ղ�n�Ī�	�nՂ��{u�<����M���E�FaB.�˗��]�&P�cH澆^����i^(U��U;9�^�o���n��y M�d� XKo�Z��bcO	���"�ؤ�4�o��WG�Wtul�G=�_6��s����Q��E����
�-0tGN��Cݕzx�D��#�m���=2\�� �=ӯ�v� �{jl�`$*�˦�s����w�،���c{����,WI�������a��(�t�sk�6���ZM�-��:g�I^	ܙ��f��,��RU�ۮxA�?�����hb��!h�V�A΅�k�k����'��@*m�j�8�'�A���k�:Y�0h.��HySz�#�D�uپ�<�MmXcj';�1�U���=�������ӡ���5�}�9��I���/J�r�p狂06	�U�Q{mg������ ��{�"�*�l��sb{�Z��^N���0,�	}0x��S�#��`��5�;̣��Y-���c�Lâ!;�A�~e�Oxh��NkH.����'��cZ�R.! �R!�pN����mi�o0�仵��ٰ���[QK��x`_���mUa�n{��=VZm5m�-�3�'p����O��B�{��pv��C�(?�t�`�@��L�@��$f���Y������W���E��xN�3��7���{�hM�����G��oTA`�٦S�u��;Pkd�q�Ρ��lǹ���	����q��M�)P*�����,P�񶌫D#��7ƽ6BL�N��5�y��G��XԼ0}��D�b"%���w�m�cY��S��xQJpK�P�pZ4����9��@��ϑ��� �ă�}V�s3�Y�� �&O3��	R���)�--u�%�MG��I��u�AJ�����V����X&?�6�/�!Q��1B�!Ҝ���'���Z<a����k+� �N�^פ�n7��8�w9K�M,�M�l�n��`����ۋ����w���+$�\;*3G�PeI�s�ۖ�r��V��,�L�0�x�����Á���-p�Cp�d�?�9�ܜ1�w��֤�u�?�g��`���W�>p�q�<� ��Ŷ���ڱ�ѵ��ؚ)����\j�{�����lߤ���ډMi�$��8@Ů����2Av���Y�b46k��ÇI�
;�~�w��rJ:+	�:��0f���n�~�����E�Yi���ڢlす�(��~ܪ�쇏���O�~@Վ'7����޿�_���2\��V`�k�% �ɚv�9� 4�Pˣ{�,�K�T���6�ɖ-��Y]��2�iJ0��u%��`y�� ���i��d;e���ޜ���54<M���4�9�[��b^��I�q�d秞�N {�r>� ��4~i\���+y�3 zrm��#�{L�i�җ�H��mA���#�_;���YP�3�������_V�٬��"%%NP���H��d@P~�^m�w�����ˡ��^\�}MP�Ćf���h�X��6��M�������m5/�Dz)�E֝n�5cm��F4��h�
���mIi'd1����\�|f�#C�������OӐ���E�Ew�+��u���.��<�z��?U?�Ah(�	.(#�E��X0�4��fF��Th������ʉ\�ؙ�N�,����[G���6��F�EZ2?WNO�p/CI?��"l�M�jx�����=�&t��)N7�����Q�6����Ŗv�����D.|���{Q��,}�oPJ��m�J��k'��j��Hl1zL���˔Y�e%M!�2־�[�[��-����M���z�b{��FFYGm�у�Y�j� h*ǟ���A��{�����v8�G�5�����*�ʂ�S��� �-�_5�:3���(b銳���H�顈0RcK��4ha��0�e�:MP �����;�T���p!���U5����7
D�z�����S~	��D,�9��V�ܾ�n�|_�؁������&���]��l`9�-]#;��H&��H�𛵾�&��܂��9dC�p��6�.���y�zWya+}<0��F�*�`�]P\kN�l����-?�?tw�l�=� $�-����Ӈ�*R$�38��H��e'E����7�u�Sg�����x�C�-���\	)���3�,-|,OQ�5�%�rQ���Ţ�j�Z��L'e��
Y�6�`'h��*�1֐m%8Oɕ�yNҤ �,�z���/Me�L�ƀ�s���{8۔�m�}⿁hޭ%+.����Z7Ǳ�A.-� ��V�aû����8������=�"�9	zEb���=|I�i�L��g�am}��H�|i�k��-���
0}�CRJ��Β���h�)���)�.Iݐ�߀.k�I���#p���θ�H1*�S�������O���j o�R7v�N���q 1\̲�ML���
�~P���^��	�!�	`^b��ظ���� 6e��+�M�ƻve;�Wo��s���LI�OFx��8�H���d�I���և�8�و�/�X�b�&d���	�x��Q؀6���p��cR�V�KM���J2��z�Ӳu�֖L6�b�2�Y�v��UZ���L�9ޡi�� Q�\���I?TB\�`�l,R?�n&�$�{X�A)��#.�T�.�����|��P���:���0\�h�3$����2�H@�������`��=Ѷ$i���Gk��>a$���Cv6 ��N��5�I��2��{��=�� 
���&���,�r|ι|O���k�=8���XG�W�i>�y`�d�u��T>ڊY|`�\u� A'����2�z�����<����6�W�C�=wuR���(x훬�o�ÍK�$26����f$]d��^����ն�u����*}P���Q;�$���j�k��q�"����^����=�\�p-��~�'t�Z�J�BB������@'�K��J��m&�vF*���}��m���3MV�3|�>�<oW�j����I?�ؕ!t�̢�7Q���:*�[��_���u�d���O��2������흮=`�Op�
7��25t?�fQs�n�d�g8���=ӁsYQHGН��o.���(���.B�w�\���J��>R.Zl�~{�lQ���T�:�<�0�:�Z�a�O�}{�SB3i
n;��Zݧ�?�Ӡ�4������S,��[]�Z���n��N.�yhK�<TSq5$[���/<ȉ|Y���jG��-d��l�y��&D
�fڧw�m<�=4O�v�MV'&:N�
/���Zn_� �3J����]$�����%���n7���ߥ~ա������UV>M'0�`�%�9M�zR�Ā�BB���k�q2G��RH����?�>�k�y&�Z���	l&���s���78.��!�s�z0������C�C��*u�&9{<f�����lM4?�����+���.f��8�߸��~E�`NQO��#2�˯�H~f��6�eP^��_A�P<��� w7n�˗��o��P�d�%qf��h �Uq�����\��	V�%���+ 1�Ȝ~����(3��f�y�4���?OMY�R���\�H�|V4'f�c��9�L� �i���a@f��6��&�D�S\����W�6"}���:�����>��P��D����EZ-�Ǹ��H����w���)��,��.�T��w�n){���mQ	��w�'�Ծ�
7�{*�0�v2�},[c����94��Vo�qf���I���r����E6x���:��z��t�1w��W��o��p<�2�-z��o�K^�{p!�M��_<Q�$[0}�"��A�4$�Y5Z�p�yy~Yv{�']�M�M��f��㦡�8��]�����+b%��?T�hBx��0Z&�����ݞ�qU��X��u�P�#��i�6ꃑ9��Ia���z/O$�Z�v�w���������%q��^qvP'��4FI;�j��F�Ƽ3��h��Z��8)���<w��!Tld|#��,����^�A8y8�z����v�W¡�J8�^����z6��p��M�j֠�rBvw'C����ë>��G�ޢ��z���)�+1}O��	����S�ˡ�u�o ���Ʒg��a��������A
K�m�Fr}Ǡ:�ř�t-�$y�����-%)�7����	��b�I��غ���N�F�jЭ�I��f�r�&��.�M���L	�#r����?P��d�zC�DJN#3$R7)5!ɾ2@;�}��XY`��T]�u"�i�83�o8��#�� ���a������~K��JS�sּdx��d#�zy�/�u�a~����Y@���6�'ѐ)�ӄ�࿼�� ��
*r�&��Uk.)#��ќ&�Pٵ.}#E
QؚX������p�C��r�������<�(� }.:�����o��{ �N��8Y���ăv���;c�D�)s���>���_��q��b�����<W��fv7���P�/h4�\~:n�?DT��-!�[ ��zv��=hiX�P)��q ʇ7T v'* }��T#�N�y�#�+�IH����e �"9���2n�qk��=�"KG�`+1ߊ⨡G��Wj�:�|�Lq���%�7�eW_	����]'����Kz8�5�j}IХ��@�Sچ�d�N��B#�f[�vd�7�>Txf2�508�/qW��7��Odg-���଒�A��o-1&��Z��5��3���rBI�;��2ҭ�� u!�a�*0�S�+Ǽϻ׈}ph�A�^!�(��䷖f�O�pV詛���"T�2���J؞r���a���������;=�Q$�_WO����"4��&�̢7�)�E�� $�O�#�@ted�6��,���`5d����"]�9�f��-��+�d�E�+�F��?;����R':Zp��o�F{2��'�C�E!���X�G6�@��ѩ�����O=���})j�a:�A���?\�TCp��xs�ɘTyi�R!v���%�k�	��BZnh��=�5�U�Nx��T����2Q��Ň~x ����!k�s� ���DŷN�g��U���ƌ��.�k5(s6w�OX��H���o,T�?�WW�K��2�s�qlM)ʍ[Wﳠ�ɐ���9�e9XG����Z��[�΅F�zR�{���Ϝ8�����-v�V��G+&ܑ��6cK7-���e+�/,ޡ�6��Pfv��Ŭ��C	
��VQe�/0��}�M{�B�mP�c�xΟ�Tg>s�"�	�ӗ�kh[0�~I��Q��B���C{��ߥ.S�!��x՘G�?�:�%o���:����Y�)+��2]8���WDv���v$����Q&�rj�h��K�����x�LIY��=F��-�p0U`�M#Ȫ�V�M��|�������5@�G�^�������!5�*D�:��ƨ٧[ɦ�7I�b�W��8�ޅ�Z���mT��oNAs"��B!�Tˏ;������'���&B6��2�u�Z�]n��T�{o�9®
�(.c�pir�ǥ�l��-Ѯ��:�.#Xd�q-���\�1{s�¡Jۭ,4�"-�x��X����{�[栦/S���ɜ�zK��Vo�̚J�J�&]�X'��A���"a L�]���D�5���x�9�]�T��(��T��G��ʮ(�u-��R��vfNs_5#�c����Gv�h��g��
�0�m�|��X#4��,?}a�G��@z���`��oj���]�\P����@*������&N��8�݅�Ȧ��)$T��#��v��_e������z7<��e�Il7�S�m�L������B4R��-��0<�V���<�
����:�.�=�����=��^�VVX-S䤂��5Po�|��N��^}z6����H�
=�9n
w�(�t9�����zx��܌�uW��#�����4 $�Kؗ/X����`��eV��U<�}^�����\���F�	o
��\��~���!Z�L���y���Q8�1��g�"1��?l��e��i��(��0�&߯�yd����Yi�J�'(W>�xfӤ�9Y Ԩc�.SI������Z#�<,��)��*��R�`����f~ �37����U��s��y'� נY.I�fĦs�>�y��ט~Z31� ��vt�0�@2�����d�b�Eq�}�떏@ژ��X��O�z��x��BS�{�(��i���.��q<]�е��M�X\��є��M�HV�J��פ�u�c��\[/)��(�@���X�jEs�Ⳝ�s���)F�����x�΃}�F-o��a&Uި"\�{J�2W8x���,n~���-(v��(����O�,U²g��ę�}��ԉ:���w
nf��/*�ٖ�x.���U<����"��@�ح�5���X�rHd�'2�|�҅�H�>��X&p� ���;qx��Y��$1:��Z<|u�^�L^����1Uȝg��������^%��^yC�:�{�l���Lp6�{�,^�o�������+,j�>؎�c�j�[<�+{�x,!���5#��
�X��{m�-;���D�,�0Ǭ� jN!��+y��]��#H��D�Lz�]^�SE�AG���ӛ�W1�>�	zl����k^��"�{���J�G�<u̙֍at�����f����Aj���<_L�1Rhqt��w�c�S<���/����I��	ԍ8�����6�,*��9R�RW��AV0��C-*��{�4۔��FU�O����ig��d��	�U)�)�8n#�-��O<��m�4�ۧ����[[�U�Q�K 9{jF�K�9�@��G�"<����[w}�P��N�T��{�UI��g��!y�P���7���0	�1�--���%�z�1Զd(ըqĥ���ڴ�� ������{�}�o���U�m�L6��T�T:j֬�Eb�K+8��b�o��sʂ�дs�|f�au�`�ny#�gZ��J\ɵu���"�Ec:LS�����E�{��r�>h��/a����?�B�?E���
�E,̐Z�&zi�s\w��A��Q��O(i/^{��r��Zk�P�)vv��Itj��eb8�pO=~?�S^aOU%�]��]
��5�pg��6��Maʻ��[N�{�k[s� �kgJOB7��s�nY�7���Fvą�ع���m�5�!�Cd-P��<�z���T$#������ފYB�2�?|�����z�G����N2Z'�󊮛3���x��5��0ҟ���ۀo
X�;��͂
?�8����|��V����*�4������� qK?�O��$�����0$o�cnjH�"�^fG#��}�S�ϯyj#����$ 	���Q�t`6�z�J�p��P�l���,7zi�4/�l��Ծ��R�bt�"E�����D�@��9#S���}���+�[�B��D��m��蓬�Ue,�d~n(}UT�|�j�w��I�oi��n��;�Q̸*o�5	���:�*����-�	�),���Rb�;���R2��Gh�2��=;-�>	�B�:=��T�g7tpt�*���M���u�xz��Z{{B�t,0o�7�b�Rm6��&i¬lw4 4@__!��̿����2:�0�x�s�ޢS8�����t_`�ܓ'�������<B���Bzc����b6I�K8,J��l��S�ڈкN'j�<��b\fg7_��@N�i��W���(����	��� xE�ӫވ��O���t���gZtQRe&����&���q�[9���	�i�b���.vL�$#Ad`l�͡U�b���ۡF���7?K���vR�`�88.��\���Aò����pN�ҁLѤ
���V
���ف#Y�J����u�lASs���	��Vm5��P�ϼ>B������c�h��t�hC`����x���ή!���3-3C?�,�{Ģ�OcO�?H��e�ZK�d<��i��1���k>�Y`�J��-��,��.�&����u�-S��s�N��L���$=j{V���`|e^132�2p�뭢���}V̅�[�I�m0�[��95J��`��
�V��
N���-9��U������$FٹQ6ey��}�����{.J�f�Z�FE+d�#��2�+���(۲�V���S-?���ڏ�&���N4��L��`���8t0M_�̈)���s��tMU��Ho2��p%ힼ��$���z�).�I���&bM;���"�$����-�wd7"���(;̭�y��({�xݖ�`C/;�A�������1|9�a���;��'��B����׬͉��>)�~����11�g;RNA��l�S��OD/V�}�Cs>��i�����>]B��ѐ�?�#����[ے�Vf(Ϭ�AV�J;,
1F�^K}?������G�'"U$�lUs;"�Y��'��U,�W�3�x�8i�a�0�������u���<���@W��(��C�*K�?�`n��=b����h�a��u!���F�Q	N��8^�Ϳ�	O�d&����fk�Js��X��r�(�V�)�i��&���B�䳥Y|�j1Ep8u�5�GW��T���
�&�]����%�I�ɘn�,1ȇ�RJ����~3/�5��>@s�����\�B��i�3���;y�0��xÒ<G4%q�E�0_Z܂������^ ����MF�m5?k�����UE���s�Q�����,n7z���f}?V�HOB��I�u�s^�ۭ���4�ݳ"��,W|o{3�]ra? �Ǖ��\��rB�q�� �
q�t�,1��� ���MR���*�]6��hP�]^���#�]	�]�b�!r{�����򀹂w��WI�*>	��<�l^��Y��An��h�m@)p`w�b�A�?�=x���!E�CH�L���xG��e���C4���^��05���; c�S�:xWj���),W@��c��+m�U���i�
���oN���j�;A9���[9HV��r4�]� &g�F�gr�֧$�֔[@)�7���.���ΖyW�W�P"nv�o3X���$���ފ�io�p������a��4VȾ�`!�a��K��Ʒ��`2Z3]��d�z��yLT��[�y?F���#�s�W|Ƙ�,��z|�"�Z1��2��vцH�zP�}�.��eSsH��ܒq��B�x%J,�L�} �BC0������r�]�+��f��I{w��8�l�%���2�Q9K`l��tQ>�ab�����$����G�PZ���ܿ�k%�Tb�[�ӳ�%ǆ::�@K�Zւr�����6���"��#����P��b9�&�DEO�dA��M���y�Gwp
����	?���@��˗y
nPjDC`�rX�)��U�o��s�PA+�EoSQ���|�ߑK�1��Y�N��I\,H�z�;>Co����aE���yN�_sA�mr�!�15R���������I���qx֋p�������,����O���:��~#���3Jlf?Uj�&�x{0n~��e�<cK��l�,�I�[����}4 lAˬUM��̽�텼�к\0J-���a�R�l��g��Ķӂ)~��3��;���[���d 0
�[Jb7�\g�4�����ש����z:�R%d�1WBq�;�;2�Vl� �^����;-����}3�]Π�	L��tL\zb���RU��L@���0+�IE>;Gg~]�'�����4+8V�#`����@WHd#4�Z��Y�O����3[<VL�H�ck��hb��Y1�Z�{|��(,+-S��5�?VyX�&_܃�d�m,���8�@v]�<ċ�����:b�?�����4Mvx\�`�%
y�yI@N�&�}�3ܝ^� �^*�Md�f��9�=?]�҈4m	�Xk<zM�^9�$�t�!p�xQ%6}.���wgWZ��Z��c��8(z�eA��z\5���͙WI���>�T�u~�ް(��y�Sj����I���&��Er�#�������t�3�Y�Q����O������w���X�z��_D:i0;����*%bi�ƗE%�$i��gx��||v��c���&����iQ���yDXM�!τw7Y/��3g����(�H2���}o�a�Q �m�^��|��P3��ۿ��]&z��T�K���my�E��,NF����s���䧉{z+DpR9|I0��|���et�F!�
��gI�@0��_�'�p���	�y��ޓ�>��J���$���'3:(=��U���K ���7{/��e��&kߦ�O�
���n0�}~.�uy'd�O�t}�"��E�'�I�|�T���	?�4ޚ�vp�ojGo���uk�t��n�:��}Y���ݓ�����L?�T3dQ��w��P��!�_����x"�*�ٮ���q����-^y��P/�~�K��-=�|h�����ԍM�W���X����	�Մ�w!���[c:�j��x4��bR��F5��H����WTO�?�/(�m�����K�,���f�|]m�}��u
��-ĳg!�v��HӉ����������.qBJo�V
�&�*�c���S��>��	� b�0{L�4�̶�%.2�T��F���'1��r8Ce Row_��E��u����Y~�%��A��O"�;Ϊ��.�]����	��E�����m�a�D�o����5�r�B��;�ĐkH��t��`ϡ�ƀ�Ҩq'<�V����K!/&���	B����V��ܖ���ʢ�ғ�M|�`�� E��
�8��tw�3��?Յ�򵙤>�&�)v��L��/�<�*@݂���d�Ԡ�/�bU>�Z����x��6A�5u�\������m�_D ��s���Yy	�֩������
�evȇ���i}�	� � #a
5K{*O��/�v54��2���d�9%���Jm>�t�X�k�9C��	�à�tCG���VF�A�ŭZ�8�:n ���*v�S
:h��S'�[�M�V���I'(\�#5G�.��߹���}�a�/7�]H~�B���qVj#,F�f�G�
�����'�;|���&k�X�#�C�SZ�H=dۧ��9����¨g	Z3�����S`!
P?x؝D��1}�U���\���58�Y6,�����y-;6�c58s��tNO�	"�dxL���/!����'�iOJh�C����W��U�uh��I��:�3q$+0+d�7WO�-5��ZW}���%(ТA��>e�p�јlV�Z֘خ���������`�[�}Oc�5�����C84���v���[iԝKt˦J�����g5g��BI>��?��m,6!�lS�L�羽�E��II�1�'Σ�yA4�B�y�'�k�ժD��}>D�%���X8�`
1�"$��v5_N���v����Z�pvU4j͒�b�q���Myn�?��t�����u�W�j�z�����z�D�p��mӆP�Q�07���d�e��g\^J>�K�o`BRƞ�`
�c���
v<j�x��]���>������x�ݞ9��� A���e�Xy+_��
b8-]�3b-`0i��p�x�z��Y�`���(w�U�����H���IW�B�P�Z5J8�K7v��9Jly*���y��]YNA���g��"�tJ�cW���9���j׀?�[/�>	�/H���T��`��A�cV�}�tV{Q�U��b}+q��l�� s0Q��j�S�v	�Fx����p�a�T���otϕ��_��� � /�{
0g��w/kH7�"��"zڢ�Q���"D?�5�����]�^����W}�?�G����'Q�?��$i:�� ��?����&�RN�7 	��W�>�rծ5��_��\p�|s7HY�&���Ƒ��jA��UVF+Jĕ$n!��<��v1���OIE��4�j�카	Q;zk�� �V��7<�C�)��%h��#�U%IK�~�{8�;�r҈��%9W�(-��ϪŗG�������;C:��pX�Rn��L���UO�����E!7�u?��0�Ĺ �Ina^0�w�Bn��K@�$�/o��Pv+���ͷ�O�*x�N��9��/H�.�ȉOl�����!���t��{{�p�e�Nǭ��SRfs	:F�09�H�<6�J��/����'X�wyhJc������ԇ����չ5^�����#tďN���t=����l�\��R���*;,����}�܅p�bn�7�����gA8�y���m滜�NO���Es�R=c҈�R3>�!�E�#~Da�1x�.~�7�ED��^7�_H˳�y�=���R�ib>�9mTO�w>�i��,
�A$؞�l��5�p �GejI�v)�lx��NR��( i�8���72�\'�."S2t����2�'2�m	�Yȫӽ1�6R�C��M��2��2�_E�%� 4E��\�mF=f=!x���N>K����w��������S%
f��o`2�����L��jX#�3���
�s��B�^���@�FÔ�o6ؘP`vG�[��;�'��n��3��l5(��
�j(Zo.O��I���q��e������"0D�5*�e��#��^���%���Kt�Q*)t��+\\���S����|�Y�/�^�٦��{�5��=��N�?f�Pi��. `>��kam��~;^���F��d����⎞�/&{v��s�Cf�"���-_�)n��k�&�WO�YL��"0���% 2Kc����JT�? O�P\���.M�lx6�	�:�����Q1�j%/�d�$&I���Jn�d�r'b����{uEF��3^���	��Y"�u�C�4�#G3�sT��:��X6@�6�����J�i�"����p��Aj���k�jT&��4� ֳL-j����ε]�r��īl��:B�����y�ۗ��ٿ �}M�Mj�U��͍d3�W3�-K&��W�s��1[�ޛDt0��q�%ۼ�����81�������v�{�[�k��m�]����"�F�EH)�7���:��8zEԢUJ��}O��R"�ϿBn��8zN��9�"gCp%4��%�:m{��Ѭ�)u���/x�R�s�.�=/J9XO���
oH3l�2�W�JI&�_T��'�rw�i���6xX�&a�t��L(��i�p�J@˔�a�ͨ�i��cO��2U�z�a���;��fnr�4SY�^�p�ٮ�\|�C��&0�	�����?os` &�Y�)�Ф�<���?k (��L��b���	T�� �[n��j��A����ߧNƭj�u(ܘh�(����n3��H��F��b%?�%�gH	��n�@IP����( /1���j$c��B��^
�P%�C��خ8�c��������~�%��d�(�P�ڀy�~AIO��d�U��ǿ�}�GE�KC}�������q,�x�]׫�g1l����w�	�yȪ�+�4��!��1����J\�)��J��etRb���4�tH�}@48��5��ܗ�:�^5Xo��']&7D���=�}<`��GA���$�.>rҊ�,���k������u�Ϭ@@�l�����Hr��_�x2@����+7B@1�Hg�c�oEZ%�:ƕmr=�'�J�X,e�����7�=hUű��\�ڿ�g�;i�V#ٺXJY� ���,'�1^���%�����V�[:d���Y`���Sv4<�)����'�+\������_�r!��%Ֆ�)��+Ļs�_�����.}?��� ��-�g��y�v�=��E��I��:�P��O����-�O��s�H�~��l&���\`�EQ
�ed0�܁r�g6پ�/{��3f�s��T����;��S���˰�Ϟ'�6<|�8>G�}�����)�$ 
$ɥ\!�]�U�L�k��܉U���yB\'�-�rD!���ʊ�ϐxI�f����{/ w��0�%z$oNr��^i8.T���V��S7���[v ˭�j��d��ګ6�8��B�u1C�'��*�m��R��>1H��U�Y6ۖs��޻9
����\�AD#ͪ��Z Lʗ7"խ��r�S�\%�G����I�u����r͋�,�T����+n\t_k��A�舘�����G�pZ7��vv�4�4��bį�����I/����^�UB�8 a�c�q+9m!.�/�vaY,��v0�M���' ��vy�o=)�]V�n�)uJ� ���F�"8�T�&R�����ﺓ5O)�G���������R4�{�u1޻f��B<$ �}'%�z`��NF5�ܭ��4�d���H�� մ:, j	ʌ=]�<��+�ű�9^�K���!H�x{��=�8xOO1*�&�9|2/��;��]&	Ig�8��_?}+��x��v_ � H�����r��v|�"��P��(�����Gm���ҧ�G0o�=�b�����_��a�"�K���F��m��i{9 �6���h�!�!���n�/J
8{���E�n�����`�{�\��h�q5��[�7�6����Q��D���@`7�^��o�,;r��H�x�Ī `�v"�"q�13���Pdc�a��Ѩ�!�E�����1e�;��
P�1z�@�5�V���-��[�ӡ!;�c���P��-�8����C���{��4eԖ`7�T|��	���9�۳.�XȘ���O���u�5{�gVk���DR��Y:��~��ق�Ȣ��鬣JО���lz�l��kʨp��ڭ��/���D�$E�o�Y!�A<���Q�O��1%�VÇΞG�v44,̞F�K��It �b_O�J�#�M/�u͖!��x@^�eB����4��Lai�ȍK��M.4Xj�P�\���xJ��b�ə���;.��(�H^p<d������H�k�;�j�G\��)��>~�>�d�~���X�>9I4]�?�˽��@G�F�#���a��n��C��Xp�N�"��L�ngR�=�&)|��E�L��F�8��1x,�bˀ�g�\r�����s�	/��Ŝ�<�T0TֱRGb�qV�{ e6wid[H���>`Ѹ�|�ǻ��4+�8�6���A�[�F���p�Ϝ��z#;��ďQm9l���_��{�!��&�Oފ�N��	c��x>�q���t=��$|� �8|�o�����s�rnAU����������
���Je0״�^8MY =2P��a'=f�e�4֧�DaUX�����n�h=M��GJ����\�l�`PЧ��"�j�\�Omx'avN�Tς�?Dz�(�X�!�f�D+A$6�>�E����!�����%s#�6���no'�厖1
_+m �hl�y����,ݪ⇤<����O"�g��J�(��%�S����|t��}��x��kH��d���D�cx�yT�W�L���h��#�����}����-��ĦaAB	���tn�[߈g�Dt�}w��̐�]L)�I(�/c� �v�Є���� ������%d��`+d+y�I��K�f��56���q	��w!UJR��p_2>�#cEX+�+�}���co����o�ؤ~>A�X�n�p�\[�����p�������:ޗ35���]�ڻ�3����(�t~xYjI�#�'C�#���<zZ��W�dÜ�u
v��E�������.�ԉ@Jm�v�(�<y�r/L���!�TȾ8i�=LG-s�� ⇋�+naT�3�} ��`��w^��꯫����h% �a<P���6�ĺ= ��u��`=�0ACyrT�;�-��K��G��d;�����B
§���㬎�a�F��v�Gj?�%�e�kT��>$��$���P�uT�;�rJB;	(�[t�N��u���n�#��s�E����K�eH괂Z��K9���0f��؉��-H��?�E.𼁎�u)��O�sjn�lC
� �8qT@M!���u��p\��*��~O������R�O�-u��� !��{�b?ε�y�&����3��h"�֧����:���0�Fj��:�B������>�b�η��Ņk�E)%x�k\��)E�-�O�Gf/_�j�I�T�sSP�<�!�.2��Q�yh
���4�Xk��������Բi�Lq��Woz�c����kC���A�Ф�-�b��7-����WSV����K����b4�pS�E���X����mݾg�M)f>�!��ZS颊�8������wK���vq��P����قzp^LU�qv��t���R%���!�&b��V�Zµ<�|J��o�Չ�1�jA"���>��X�B�|��We=es<�P�wV�l^���k�ƆS,��&���L
��x�݌�^�$��dp�E��L�^ ��좶n�ޚ��:Jst侻?A�vN���l�|�,/aER���*�}=9����c�K�K���Ԕ$�NK�#.�D���v'ۘd��H
��l�n��DL�t5��4�'u-��#�'$�U�J���n-]c���?�@���ƾF�����8nY���p$�%I-�Yn���O��E�0�3�;Y�j��&�Dg�vV��S,�%4�d�2��\�����|���Ȭ>д��LC�z�gZ�<��뉄 _��՟�I��j�]��7��lҨ�0��;(�"q92@<=�a�V����sp�a�!��҅?�B���,�8�M�EW}��[�!�ߴs�D��S��.��%kf������c?�#̸�&�K��/p7%g 2��M����v`��'�Q�q�\���uz�i������/����(x���7d�ȞT��O�����u��պ� �'�`���@��L�Y���^�~T+����yş�ؒN^�Ä�#���Ӡ���Y�9N<!��☶v��8������%t��8�5�F�s���FuD�y���v�|�W�K�mشq0��Z����2h&<�X�ٻ؅��e��u``�V�	��*r�y��#���F�D�$�?Nu6�~�{�׆�a�"f�A�ׄ~��RDM�pJ��IUy�ʠ�.B>��F��׮�IX�����"b$&;f��l�#�:���! ���
M����l��KOO��bM�(-�V^�Kr��������f=C���2�8V-S>�Ǭ����7FM���ր<P 
,�X�a+ߴ%��'�l���&6lA\�����a�3��c��X]�*sb��J&T�xSAc�߉�T���xi���b�����`F"�A{�Е���X�7lR"M%Z\ė����A��$kqr�`���j�G��5�F��O��⫌/(�i�J����̗=@_.f���1Y�`q���0�v֠���"�t]��]I�Z�(��U)�N����ʢ��Y_�)F�j�[�����C���0��9�ZB>��,���q6�g9a���X�"J`��Z��c��<a�,5@Ęĳ/�j��T@G�t�'w��6��u�ee��L\]k���07�%Ku\��"I=2���qX�S�X?.�o��c�]��|��Q^��+�C��7h��� 9@���S�E�e�Ab�(�$$�{]XaB]�e�W��R����Q������t�6�q�L���/�6���J��2�Je�B:��W���>�:��T�9�`����i�_
P-ʀ�2�ı�!�3�V�c%���nF�z]7���F,f���5 ���0�,,�4WC���֫̇�pa��E�����E{���Ui6
��9��-�����7:a�n���׽�Pr��Iץ��<J>ڟ���yNYt�����d�~��i`�U`�2(����B�&� 7Wl�k��j@_�E�c��-u���4a���k�x5ʀF��������h�a'�iyUSL#�ۃC�1n�W�������%����/щ�R�eL0|�,m�:$����f�m���3�~A1S�M��tҿ4Z)�}w@�mԻ6�5V�J%�ΰ𧮭:����j*!<(J#���W8jx��T�\-�ظʹ�,J��R!�B#�i��6|զ�ي�IuI.g_��uv �ԙ��{����퀌[6h��) ��k�4]�9(c�6�j����lEC;ؿ��M~�/��
�=W	���:�z-��,��J�����f��QZ��t��6��c{y��~yZ�M����K�5(��v��m��(�Nq+�nR�Ǯ�M1�y���+qS�i�)զ:e���{�Q!s�IUG�k�?F���E�qP=��4��7f������scC|Ǚ2BI��� p�AM�K>2R�B���P	ۖ���%�g��Чh(��x�L{�jP;���=	ݰG�� ��a�kђԨI�(���G[��S�����»����P"EL��~8�f�39�LZp����+R!�7�@�NwK�����ZOhh��0�{4{�����V�]�E��>^G�LL�	�}_$�8~[����k�XHr��sŻ�ȊΗ��)ſb}^	|3JYc<�B��m���S-ٕ0���8  ̊Yl���O��Ա��{Q�i�r��G�}�N/�JMU�R���r���r��'Q�l��*u�	�K��=��_�h���Ȉ�&���-M>"�wB�IL��'�A��� <�<�7I�(�V�
��6��4D�{܊X��o���F�կ�����[=Y�s�K��:�?�H�r��B=�����g�A��J�yoW�0q1Ϳl��o2��[f�J��'	K��E �Mf��1H��Η({�2X�+����;3)����U���+0G���>��f�D� B�M���6F�k�Aj�Q���%��!F��_�c�[O��~;��Z��Ң��H��A%���ja�+ʅL�3��v(.r,��m�E��h\Z� �ҡ^..�/��PH&�X��+���o���aBT��[��J��ݝ�Omz1�	�NX������+o�>�Z��~g��W�aG�	�	�
�����'���醤Hȥ��x��:j�Z�h$�ͧ�\f��Q�ꨫp�ϥ@P����h"#2������eF�������A�v]�-��LikX��k�i�B���DКQ���p��K`�#q}�P��S��sG9nn�B�&I��i�s�ұa�~�/�� 5lEq9R`��M1ݴ���b�L��F �m +�!k���5Z3���)3rW��K��d������C0h�!+ǟ�	�JZ�b��ْ����|H���0P�G�J�I]_a�������O�܈}Q�iէ��ܬ @�K��)*�V��.P�:u����R�i��n������zg�C�lc�b{>�*��c�1ã��M�M�3b��P�Il�NI�$�A��,d��d�TBGom���]^OMfcxƭv���F�pB*CݱM>�{��Ʌg,0C놨�3ȍܸ�E��D�e!���P��~Q�\1�uj�4�ϐ�@�6ַF`W@B�A;�T��� ~�tUՋ����w"йCM��Y΃;.�g�����"�Lƪ�|nV��V�\ّ�r��	�Jc
Q�m��w�fW���Fw���}�F����%�;�g�ڨv�X��W�%��y6L/GKRXS�*��-\[���y}��S������œ6Pm��pl��M%r��W'c�t�~����T�f��{��Aw�BZ*ٿ��CQ��3� �j��D���Y1��?"�*���f�xK�e��_�6ل��W�a"ŕv�bŨ�ЋB��&g~$����QpRU ��	�x)I(�^�$�R��D��!�{0J���y�x���a�R֫�:��ٱ�\QMn�ނ^⻏8-W�.�w�	�[�^2�t�q-~�>��!P1���Y�������3yէep&��	�l�ұ��j[`c�[���Q-��2f$� wPXD�b���A����~���uG`�7�Aā�]ؤ{_>-�]=�����2�!h<��Lq_B�ZYMf�qe#����l�`(����/�	�d'#�E�7����������(d�����Ʊ%�x���5q���XСv��e�PO�N��Q���3�A�()
V�������n+�l�v���|;�76
\����:�F��	�@��*l<���8�w������)q�e%fX�?��ޓD>(<��L���m���0؊�y�����o
��B����b�^<��hC+ ��ԎF[�+i��f\i�P�FPw��lMW���q�;]ܵ�����l��gC-�Q����w��j; �zĴIZ��/����{�D)�,SpzU�����8�%�{갛�U��:GQ.o�;�^.��C�p���y�BSr
��b+g�o��&��n�V	��D�DkF��$��.	�胢C�R�MtL�5���iПT<�����S�h�D�F��f{�B��`>��yf�iu@,�FjlS4��[���!���wD�V"FG8 Έ>���j�^�#͚�&�ؼ*���c����"�r���  �;R2BX�mQ�D�lC)f1"���1�6�Zp_�]�jeB��+����&���O�?�f����2t�e)X+%���&4�~{�N�%?�H^��������Ot�a�Lװ��{���l���M���8�|ɌT ��v�R�H�����f��G{���ߝ}�3c��Ŝ�@P�YU�m��+?��a����*�*����eD���̵P�E���<��eF����A����Ԥ��p��i��v�<�����\��؃	��>|1+���(P!�!�M��K���l��e��G���2q7�*����
�1�����SP׳]6F��,��x�6g(�L:�ܘ�<��&�6�y��}�J�ž�"�5/��aX��4�\��W���;.)�s͌���1
���u[>S��?��sG����ƪ�<uo����c=�e���;���6��������Ͱ�t�{��fT�(2%[bҳ���3rX��ߝ��G�=*m�<�쩷ͨ���,�X<�m�/�;d�[k�(�ҍ���f�KHy�9��RD�X[�:s|�cI'��W�	��}���s���b��舘i0��o��)H�"��������B2*Nm��y�FOW��.2�TG�����`��V�x GT�x�lH��d�ց�k<Z�g�ƭ���Q:��J\�w
X���۱ i�.�$���Th�VS}��+�m�dbx:!H �!Ǥ~V�˙Bav��bȔ|V㪇2H�q0��z0!��d>��ي�ܓWN-�2���w1�U���hOɌ;�"��k�$�R�^���hKur�TW���DI\�u��4��X������$��h�847!?	�|J'E�9!B:�J��K"�W�\=��a��BRj-�ۤƈ��}=5�7 VG1d��{V�a3���C��&0�?�GC2�����R�A>�s��7�ޔ�9G`6𥖑(k��ARƻ;�*�f&R\$��ʂ� 3���z#v!��-�r�|�8 ��4�'�yn��\hvR�v�
g>�,s~u%jZ6~c0j�:�~��+v�?�P�	�,��^\�n�
�(Q�ߵPړ~�ե��򦷳ٮ��;	B�傓>q��i~��_�u�G��Wmy�M��S?g�x.����%�4/s�+yQ;�*���\_�0n�S�nA��x��L��k���cZ�J�e��X�V �h�瓥pa�Ӯm�1�Dj���M�m��*� ��Ɖ�0S�A|���t�t�M,��e?"�d��!?"�ܳ\�~��,�ݎ�m!m�l{ݤ�(�fL���v?�]�3�J���y��ː?���Q�E�E�Z���,�����9)�d��g�R��Cm��G����7����X��\gF����vG9hj�عiud4����
@b��̀V;��~7��1�9҂`~|���-s�!��K}`�>�X���Fh�z�߯#k�y�i%�p�� n<y����'��.�5 �ɧ����U6�o�/����x�:�.҉�&z�{�p���SU0�%����[1n� ��C#VP�`ϐ��s��I�����+\��W��Y^��o�+�brRs2"�N���g��dl��rMI7�&���L��)�������뤿r��ѐ�&L��ޏ~���D��$�����Ѧ�rPu>���8n�G�Ȣ�UgnY���|�P~jd�m䭽�t�I�x�B���2�1��m������D��S�����
�tWÌ*���Rb/r�F�}#�ʕ�h��_�f�nln=I��F��IE�T�O� X`����.<O.�v��85�1�S��0�iv��QFq�	$5�ҡ6+��(��7���W*��eq�{��S��F�h���+��g��g6n�7�pS݉Y/��	fy�����( ��P��W'�[ӆ~_�.�Wta�%�ט�j:��$|�$Д�������#1c�D;"�h�8M�hR0'���p���Q�=Pk�{�kn�-��ݓ4,���1��v�HjD�-��H�Ü�H�Z{eY�pA��\�Ī�zX���o����O*��j��_�:iݣέ0��5k?�#/�9@t����'	�����~>w�#�1�Eq��x	�z�^QaZ�QF��,8��g����.���������QRh���Ύ|�����>�f}���W+�[;Ke� ��/}/��3��*�Y�Eo2P<G����v�K�)�bxZn��Lt`����M��=4�3�eD�no���G�D��z  �v��{�ˢ���A��6(�z���@A�0I���x�/6=.*��I�R�2.�:^��?W���R�cu�%R�r�
��s�[3�d0��!��%�(s*�ـ6�Y*��%D��%4�C ���,��|�ox�^��	����˅@zϣ�yPOݗ��C�Aa��7!���X}u �,�����)X���L�>�ʌ����r�f�S:��xp��L9��j�����K.)X��,f��Z
1��]���5����[�MD--׶�"�sހ/����yd�-�e?L�X�q�u1R|�d�O�ϳT�c_�Xu1~��g�����q]�z'g�m"��Y/��5$\��ft������6�F�0Z��X�K���k���a/sé�&���>�(Q#�e�mW�O����'�P&�U�@j��L���������*�S��E��Q�p{�¸|g8�ޏ0ԅ�[>�#�IvԚu��<�-44�za�4�{�a3>���,�III��U?�o
<M䈕{�K�)�y��8{�;r�{��ϴ%?#��h�\m�$/� me�\���k6�wmq7�� 	�;|$���<~�5��:?ʭ3{眤� �i�y�}�⬭,T�$w ���{�O
&�L�l����%���c|���E[�b�k<�Ω�W�)��]=��1�zv��o�����<��P�f��N�O)�`���M���tzk�(}�[ө���\�O����L(��O�ݫr�6��a+[:��i��������;�46��i�B,�Ȓ��Έ`ŶS�J�tG�� ��-���*���ɰ����/����j��6�z[��Q
���ᔱ�?zSⱃ�T5��
�/�mMI��b�1��p�\.����рK�=�3�ʒ:�(�Ô�L�+5�.E�j=+�kű�d��������"ѡU�Yɾ�D��<�8hq�8If�%s����Oz1��T]X`T��-0��r��~y��߇'x����#tZ$�o�Y�,���m���V�U��#�a+�e�.u�֒J-�ù\�^;.�5�����7��5�5�S�	�����*���E�㿗c��6�b�M�l��>�.�f#��?]�V�G��p����fg$��V�A�X��p���϶n��	�Zr9d��P,�2u�w:�cР�ߊ�2p�5��U�l@��0����<��*�	��m�Y�����bѤ	-�V"!P�ؼ�P�/ɛ�7KI^l�p�rZ
Έ#�^��e�u��]U�r��P�fC�l�uΐa���T��/�=�r��SYl���:s��Q���y��i��NaE��D��W��)}�<���0�(i ŵp�����Q�i@NαE�G|C������V�e]XqM���D��^�В��t�! �8V���㮰�3����+ �uW���Y��V����,�������r�J�^��$$~�*�����B^q��p��@
�ⷯ�����w&v��}4�\'��4��>P���溓o���y���~g��£ ER�F�pl�%�+2ϰR�͏����|�k��i��\���f��g��^��/[�(�
o���)L?�Nގ�0-m�ͽm=)]��ӥ�ы�)���6Q��]��q� �������Ǯg責� ��I�̚�'`��ܒY�1��1W�2��_M̅�ԋ�'��W�ĭR�;�*W,�oH4�V#2ַ\���Ο̙i���Z�:--7���F���Q��ki2�H+�kZw�ϱjcF�� �oi5���VMރ5�1����Rz����ѧ�C���Bh�����C�Dds�EPH8!:�u������m�_*E�<s��
.����܃֫u��Fcc��6��Q&jf,`~��1$�g[�@g4R�r�.r^����q��;��l	��Ep�>�Z�i�,�9O�O����Z*0i�5��X���Zw��$BJ@i�QR��%|ح�9�C@4#�d-�ꧤ��~]�ŭz��r��9�\�0�h>�s'%ڬ̧��m���E���Bqw���_�&�ϕ!�����ݾWY ���v�Q�א�Q׎������UO҉�����D�Dg��c�77�8�~;(z ��y�~Gah47^,�X��Q�t�����op!q���΄�I/��j�m�_���u#�X��-���`؁�M�ɍ+���a>_�n�|k�Pk�&��^�5S|: ��k焩�4��x����;&�o��Q�
ٮt�K@��@ظ�_~�M�{~�;b��^�=�T/�0 �`=�����EN�����8�����]�0����S�>����S�6�3���0���h���~j�&�n���6�@^��sh�ߟ��%��Q��:֙ ��g��~zm�~� ���ev��8����1���xS�hd=�Yw%yW[8�zY@YE�]�;,�L;�GC�����6X�3J�Z����/ Mq��+X&|\��3]��;7��Hц�$>C6x��ʩ�B��u�a�96Ǆ�̮NU�e��;��GĶDC����.�ޚ�������W�P����I4����
��ț)�ĕ�.��� ��C ��._��:��<�1�M���<�%�����IHNvC_�|S��mOp�?hncj���A���s�s%83p1�Q�3n
��\�Nr��󑀀�cq�}bM}kyd�$=Jx�Gsܾ�����W�菳ǲ��T�W{�SQ�
6���"�B�������Eu��u�~KR��sQ! x��o~W&�x �y����7@V����WĔA��1�裂:�����l~Rq�2/���\eV{�?�<(#Ӗ71d��J�����L�#$٢��Cy�;5�����[x����8��&���۟=�BwunT���P��z��C��
�^+�G���2r!X��-!EgNf�|xIu��Z+7�LZ�#m�ة(�!}��R:>C6R0��n�,�k�Z�%k�O$2(L���\���~{ ���0����G�9��lMam�^:�F5����i�l`��=�ǒVboh� �QdZF������&���#���5IӲ�ð�D2���7�O8�\�=�Nqj��3�O�k���^#�|�&x�B"�-�U'�wU�.��/y|���뎒�ħ݊�x�u%��cįj^��`�v˸׶?A���%X�&�VVQ��BG��pd����B�W��YZ�~��<#b�Jρ�zJ
i��'DUY��q�v����P�b�����*�)����"�7�g`�p9fiI��L�6 -)�.�(��͠�
9�U�/������1�c�͇YM�	@�{����8!�t�f��\����o�]S|]=F���rȀ��6��G9/������B�����p�]O1b�Ll�ro�)�f����[E3�M�3ݬ�M�9.�r+�x?���g��0��>��ʼ���G�������r�R�5��|HV�t��tO��<[���=�p)q\��_�Y�ݮ5kF�%�r�U�鱶!ӗK�8N���JY�V��>k��H;AG�~W�vB$Y�O�E	�E�o�����w�<�����ۑ��ۅ���x���M���A-aj�'������E|�r�/�l2�C�	�%4���>=<�q���k��А}��o���+~g������n:0�;��w�^��e���Rj��7�����o�Q�K�J��*zjy��n��YC����{��g�[�~K>�&�F�c���a)q�/�^|u�P�`N�p&vS�����8"^�!�Ϝt�g�|
g��>#I����x}��\�q��n�h}�a�!�x)�+C�;��&Z������>wv��7+qO`uKe�<�ƒ����9�)bV�l`�D����bX��5�8���*VLx^����#ը<�P׻�筙	o��ב�?~N+,[V��n�N�|����gJ��hx��wb�?���ӂ:���}T�n}Y�~,?W;}T�H���!4jw����'�.%�.��(����Tj��"ŵ�3�)ۉ��wH[	�R������o� ڎ�,��|	Y��߽N�7��ܶ�ɹ�K�ҡuD��btq
�PP\�.F⎏��dYHK��h�2N��l��?�$���Eً���� g̍�:X(�V��d�gYd!=�3GQ+�1�� Mzin�Y<0��7&�q������w�T��MɄ|�/_����C�o)�Z3��U!�/�]g^�jF��\�b�<��ĐCB?��/�����`�˧R��O��[<$���z�F#�ih������@s�qX&'G3������MѺ��F	8�#��nz�bD�\(^�?�����6�`n��K�Z������%��"p�ya���}���w(*)A
���[N}3��j5��ҥ%�VV-���"��<�gZTx��C
��ܼ�c!�
�z�I�6��D�E��V=���<g��E�@�9Ǐ�L�H�� �b*�3/n�\f����zU�(1?mh.x&ϖpT4�<R�%�A�1d��<�oЊ���em~	�NMS i�lۣh��0���pk��j�4�k@��CG)������A��T�l3��yI��.h����>��6:sw�wI$�n����@>���]F=�e2tW��??j���������(�|��3)�b���1�뢩��ly*�J3�L�I��Ӷ~��җ��Ѯ��h]ta����خ�����W�q�P��ܷ8�X�u��vyx`!� 7�5x�bz)
Z7�C͌k�1��Q��'�)5��7���E�å� �#�Y5�wJ�Y����bqQxC9�/��a���L}��4�B턫7�.��0�B�8	�-"�:W�Y��{�q��G�T2;�F�#�$P�s��
���]j�3�c�"���\
����2XRW�W�AeA�;w膢'�&��� ��;�z�<�ms��vi%��Tg�6��,=���ǝF�T�o�eE�9Y��1T�O�¶�|�i}�tm~��u)��L�!�+4������Z8��Q2�!$�wه��JtlP	�qs9�(�����ܢ�ԸW�X�ީ� �/�R%r`���)��n�m���!OX�����ڄ��7"+�)���Ƣ�m�_�R���I�#�z� �g"vjE�n������H �M�,&e��х ޣLv��P�vA�A_D]JD<��LM��!������O���A�Ӻ���hH��5���"���WE�6���x<��U�����A����LU��S1�a���͊��e�@[JB��|�}z�I����lv�?7�E�hh%r��h�1��Br���_��F��\v�>��d�U��Ο~���7���9�^����V[C]q�{�z�IRQ*l��D�d��Cĥ�/u4��X%}��E���q�!��v:�4*�����P��}i�!0��d�%�0�?c|p���mb(�HZĸz��B�ͺ�b�~�kk��gacn���!��`������JWpÙ� �FI5՘�QL��t�Ϳd1�Y@�=T��>�9O�a�@=�+��ꟃ0B?/�Q�޳��>�Yե E-��>�ժ�v"�!z���o�����4�6d�)�8�Ow�|M�=-	�I'ǵb{~*~w;.9��ݜZ�:�k>Ba��t���ve�,O�xF\�Ӯ�^f5��ĿZ�byuO�B7%��R�e��sU��zҜ����.a�����U��D#`	Sւ�)�x������_(���Ϊ�ď��х�K�c蛇:����4s�JY&�EX�5|���L0f��MX�Ml��[X�;���d�b�[�Jw,��	ԋ?�©[���?IL�Oy�4�����O]������Sڐ��rxr0�;���Q�D �|k�����2�N���՗9�qw�hHp`H���d���:�E���\�#bN{@"W�j1��O�C��
����TLѫr����)�{�y�jsz��gGi&���yc��%��mQM�nI�"�p��7ε�81<��qW�G1u�qo���O�]�K�S���o�j$�w��XheF���<8���Hh�$|+u�����RAnD@����X����`�lX��vv�sR���L��H5#�	���l�i�1�·12�߸��C�6QT�H��x</%���R��t��^��1�L�q�mt�<_���{�wņ[�a=j��
K�۵�dt�����YB�lN�B��Y3�����c-NnP7��GG��Y ����ߓrb����gM_��Ҙ�42���1E�p���>K��:x���0��=G�{DG-<5�=���'�Hī�`���17�2 a4~�[�7��hA�*?�|��}.� T��H����" èF�*�㵻��o۾q���{��v�aQCo2~�T����-p��]G�nF�,�6V�$�,lS��	q=�V����9�1Sֈ�FT���KK.�zj��Y���z,6=�PP��b��^�|�Jfɚ8p�K�'n�����4��/Q�_><�����9/��áG����-�-e0�ǣ�Sk�I�ơ���;gvYj��;4�)�l��5\����>i�H�8�	�n��Ƀޙ#��|��d���Tph�'~C�@�iA��m�dA%IO��%Ӫ�A�x
�<L�V@�R�H���&DP'O@my�e��5����s;n�Yv蒅���V�_��v�A�T*p�a�XMi�d?-S9�O$t�����S�&JPՔ�����Sl�"��=O�}���6�lCe��":_(�Ü-.��@�U�<���c(bp�7J�^���p�B-Ԍ�[EVQk�%)Z]�_����K�B�w	Qo���j����&���j���7��%GE���<5�o����Z$��ckI���#�$1)���q��Љ�{�!h�#ih�&�ͽ�܊'����Ӣ9�<����R�Y�� x��La%\���qlF����L�MD;i����7�yU�|���},�����ȷ��`�����{�B'��y �'���N�C�CY(ϝ��o������i�M�ޮl���D"�B�Q� 1uu7ڽ��E��˵�m�TLkԗ�:�+xNX,��bk����ԅ<��L*�F^�+E����9��ˎC)vg@�i�+�@ ���n�[Զ���x� �����A
�F��rDa�y���ךR8ۚ�ұ��:����IjqM���>eذ�qMs��8 �E�K��?��ӳ���W_��p�&y���#�V�-���1���:��~�F�D��j�W�f�]�
$���+���LV�_U��4r���$����VK�wx�O�V���8���+@�#ƆW���H�r�.g0~�(M�ejÑc̄��.!�0��}�I��*\���?2RYOR��N������υLJ$��GZ�6��E�J��on=���x�,[�*?���R�pٰ�|�?@�/*JXGj�Ӌ8��O}�Hmx�	�>\�F5��n���Ο�n�
Onl:���2s<����[ص�B3�ëD��zf.q��ʛk<��^ڔ§Vm����<�J ;�#B�Щ�f���׈ݽ���Y^1�,���2��79��V_~	t

uf�q�(�PO���X��,z�K�y�'��x��K�Pn���`[�םF(jvġ��g���R�P����j[P0l���]��fԛN^���8��{"粷Q��/�?�s��?�oO쾝��"�S�8����E�~o�8O��3��ps<~^�Ԓor�o��&�VO^�Da��#��Y�a�QCgRf��+�s���"}ݸ%�9���j
�bu��xq�g�+��oQI�,4�����j&M�@Z�߇k,W&3�8�4W��n�D%?�ge�l��;�(v�@(�o��eP�{�qN���s3�]57���p�$�NS��OkZvY֦
����)�#CSw39���oe�;ƫfu�2�<턆���q�D�Qh�N��jB����eE1�)��"�:m9=����mVZ�f��W�>M�!���Xv����;�uAx}���bZ|I�pf�p��?�w;�V�H����������|�	��b8y�=����B��b5�ZK��.ހjW��'�,��+z����]��b}����_��Y�'7my�@�t�x��1��p�*a�J0��S� Ϧ�8�F�o��w�w�p�<ڏT�;�.D��m���-!�=�|  GRG��(�e���,��ao�A������>om��6���g{��*.����^4!���U�| �� ��i?��ќ�����/��y�:�'��T7?1}Y�]픍h���<�Zi��D5$v]Y�!�8�� r��A4�m�A�}��O<tp?��6�<Ӭ9D�!%�{�T�J ����6�W/Ƣ�|�!�̓�Y��"�\<U��(J5���能{�[����hm�� �|����0�JnEn�W�ꝡ׺�!���m ��&N��\��~��OqF�8EG��3�dY���Ry�B#��.;��]�U�z �>r�
[���i�r���f�܍I�i�tՙ�7Z�3��Z�ak *}բ��;q�P4/�J?��P�Kݣ�,��l��	W�<�}0���|��D�������;�P�:�o����������VH�3s.����'���K��/�R��,/k�t�9�p��U����i$�ڎ�(�ڸ�P`wk�*L��5�i.z*��S�V0�
�'nUnn����/�i�+A�K*�9�Ed�i}ӄ{!���v�}�L���j9�/`��v٭�oq�ФEb���>��s��*�����.H��#��c��hglf^��^�-��0,wG����(����+Y�5s�Z	6C���Y'�Y`^�$�ϵ#�؜��y��b�<�@��w&h�9�o(6�{�D� m���7߱aQO�yr�r�1U1D"U8��ݥs���ZX�8Yh+�9G��ס�Q1b�1�h��[U9u��P�g�+���g�D*쑘��D*W����"}+�.�y�kՉ�A�����R��5'T(����3�\{��z�W�  tp��(}��
K�C�d� �
���M?r�i��plvט����=.a�ey`=U�D������wR"Uw�����8����8����%�^�RI:�\!��v�˭@t�	� P]s�����
|�(�V�,_��$��J�gj�Ǡ:�/�b@�խ��o�k������|��ͮ����"�pv�wyU�u�5Б̖�̵�}��gU�w��p4R�T���=N�����y^��,����պ��O�_���H��+"q-���`��Ai�=��i���#⋁���?�k}X�h��ۆ�$�t����=�^���5w�9�W�Lc�D��9Z��jRv��Ypl�@�u�z��+ u�`���1�t�����92��0y��P()��1��T&��c��U��#�}�(��3�׫��=k�.ش9m��>��h�<�t*��{���N�š�h�Nn�,D7tm�'g�+�?蓉����[W��o��r'�#��ƍ�W�?S} �5�F�=�&׮R��i�k��K�C��O̧0�%,�	R7���]�ۤ��e�\&#��)/[�̗ef( �*j��#ſq�ΐ��d�f��_� �a&4*�Y�][��Yv@�.��������>���.��z(�kX)�d��"࿞F�S
�"�g���a�]Ǖ�s���Z�u77U%W�(n�'��F�;枖̵&��$������c�ƃ|q|t���[��(�	*�g?�>�&JY�\\�����K`���Uz9�p�-�3)�Z�L9�&.vc��|uZY�hO�C�{��j��PVL�����	�A;����!"~
wb��*]���;� ��C`ü.�d`Y�3���<�L �rD �����~���#pںf�����R�R��јp���V���'h�U�C���|�֏��Q{ϴ"Co��5��!�q�j�f�-�;D,������Z?9��!`ѿ&Z�I�朴@���O�Z(A�ܾ�k�n��dͣ�?h�e��K�|��-�#Rĥ,@�:q�y�NF�(�S�*��L�}�*�x���ҏ����.M��)��92�+�����]��Hu�P������M=�j�F���N���2������b?�S��3'HU�wD�+B�ņE�����y�MUzM��Ƹ������U�tS���s&.-�K���s`�R�aO.:�7}3����2��!���we�	�Ssxt�9�s�Z+��_�z_f�%�^��)�X�_�m�,aY@��1��ȟ�HSգ6�Ma��!b����K�k�p�9sW�{��S<������5��n�ί;��Z�(��X�.��?ǰ>�[Us�E���H���A��L���k<
�a܉��|��SbU A�x��(�����_*O�:�����J�&�	.2-�
�ɁSNo d	�Iw��RZ���O���#�-�ƞ����X�bE*`L7�
�W㍱�$(�j�2J��ҕ�y��Xf��;���P+dӵ����sK�<��&pR�Ƥ6͟�>e�0�М�n�;����B4K4��2M�kx����G3�+t��[�5��H�
6_�f��p"K��O��@�������T?�G���3Sg2����߀#ly��P-�}.)er�徑<�0,�q ���5X ���ֿS�����j�����Kt��ώ@��t��^�É���3?���;A(�'��Y�����A\��<CO`)�;�����PM��~�iʴ�A�m���@��`p�z��EW��Ț�-e�e?V��u��Q4>��]��i�� �?���y�Y�����dJ蹴0�#
Q��7j��_���ڲpG��#�G(�~g�o�g������F�g*W���o��b{��&���Z��}�3jH�>��(��57����meD!��%?���/5�,�ee7*=�K?���۸�c�f~���W��"���h?�vJ��V.@J�s��dD:Ľ:�c��@�>M�P�u�"��D���-'����|�_󂽍}�p��X�B������nD�iL|y=NYn�<3�Ə_��gٖRhu^1艊W����E�{1�l�=.�}"��_ŬZH���G�s��{���&]*���s��q� �ہi�J�����g��[�gH]��iu���K��U�T��
�Fx�T��ͻ���ga
M���7���섡V�Z@�Uc4%T�+W~�I��!~�+�{���p^�q�&�m�����,�'��5�]w��,��g��i�K�*j�T�M_��Noe�� �C���T���=��L��W{��ANA�P^���y�+�٭)P�%�K�׈� �<b������1��M����w��w�{�m[�Z%c�[�V+�&���d���0s1�=J����`N���Is@�|�p	���iG��1e2���"R�િGM:Wr�HB5���'2Ր)��H��Δɔ��>���$b���X�fm�����!,��{��(VR�V��υe>��ݏ���*M�nQbEV�g�$��RO>�j������������|� � �2j�1���I�?���+�&�qa�����mۑ\���P��"��A7�N�����mfu���F���[���Y��IHr^���j���,��'r}O:x�|����~Ќ�����ǺF��.گ�ս��Q
�Q�o���뙫�;W��f0dz�O�9.��&>^�ut����V�q0��;��Es��^َT��i�5eZY����{w�v&�b�#�[�v�O@'�C���)�%ڇa@�
�Оy�A��u.��3���D�_F�v=�=z5�` ��w
��xO�������}T���mt6&â�3��ᚖ`��UY��$�V�b�k`�8�g+퐴�c�F�z��B��e2a�ȽaS'U�� W�&'������YA`�秵���o�s��I3(y:u��D{��%��$�:d#�[���w���s`hE��<�?r9�Ţ���V�l��t�Ux�o�r ����f���\YpJ>�#ʠč�ދ͠A��/�s1|w@��T~᫋������lQ��%#�c���pM�����0H�{c��������ߏ�'|�ڲ�����_���7G���zać1�i <��u]�2�=E�:�@�69��	3LDOJ�o������X���B4�K��=X9��`�?��,�z��ʌj?�]��aVX��L�<����'U^[�N���T���a;O����]}�����=��0�g��,C]��oި���D^C�)Z�[�A�ϭ�D"�#��|��vK�r+�\�H��(SZ؉ �hB8����V�>���mO�p�Х�a�y!��ؤuj��J_��`�M$��2�q*H�|�w��)#<M-c^�b��-?C�)I�,ݜ���J�L_�~���Vo휥DZ@+k���3B�!I�%X���Jd��ė&�ڣx��C���'�Q3�DX����ǿ޷`ĀJ������Z�U��[�mbHӉ��7��Q|�<�i���u�~�x�%zQ��r���`�T��c�֍�淙_�����`�!#��1��W|����p���2L�u���!C3ILs<z Am
-�q��;�_U,Ǌ0�1]zq�);��]p ���
=��҂�FD�=��۷Dإ3R���8�c���ec��q!R��u%�ԛU�g�J'�ǭ�׏)D�WYu��K2U=���6Q��  �d=��k����CmU6r�yp��j��x�_����9�P�1&��}�k#,b3hPπ�&ΐ��Q�Q�U�iFyR"^��|Vi R*��~I�rGc��J��Z��©��6������k1��X��0�z<-��[>7B�G-��T�;�@RY��n*����-����.Md�=�2ϧ����D7��f�dsP��z��m8 �;)>PW���|
hW�F�r �/:>�2WD̅eVJ��`���+X��o%O���D=^-����6��/2)@�W�>���v��[%o��A��<���c'�
����p掫?�_�/@�!u��v��	T�0{�	�,w�^�6�������jу��~�Dz"��M�N�HD�~pD��n�j�g�n(�{��׺�D����3����r�}���4B��J"�&�J��.���	����t��Ɖ����0!�yn��D��?yk sDпr������#	�=�
&�r���k�ɒ0>̘Lj;͙�xn�4����DY���Co@QQ2��U�.Q��{m�B��B�6��r�*+n��I��NsV�G���2�����R�u$�J����9#	@���q�U������!?�ɥy*�9��@r�������x�xJ�-����aJ�:r������p�qIUͰ�F�D�4��4�F�lAF�܀�eo�/P
��r���C���|�b{p,:�(h4 ��Jlf���S�_uy^��0-�+��y���z��m�Tw����>_-ژ��-`(�&N��f�@㑷=����L�7�`7:˹������*ʑ1v�ׂh���]���jЪ}����� �����7�̛E��#	#5���.�`�̰�)����1tU`�9��9�:Lg�*1nu�E}g��f�[	xUr�[8?���M{��&�S�t{^���%8�/%��C��-�*7���rg1���Oi�
�E�`��9 �E�-.��j�s8���*��3#t1>�@�Q;;ҩ!�`�D���2�Fz�\?���24
���Z�*)��H_~F�L�*?��Grթ�eF��ֹ�N(ժ�C��p#�����6����Ih6�`��#Ӎ(��p%)+��
��̖e �t�H??���!�ƽ²��A��0A��Qzl�{��l�1�c�Z#�=Q�O�vcHt��uA����I��Z�m<�Ѧ�����R:��
M������a�u㲖A���7 &�f�1~z�3~6C��������_E��@�߻% ���=�mc���R㭺��W��8��t�0��1�/"��q�����J�y0�vù�y��Β�*����ci2B�.�h7�fJR��c���>q��&��]䘚�RYD�iV||K��+�݂$�?��n3�})
��\�"iD
��ڙL���	���2�~(��_s��6ߺ`��~/��<�HXZT��K2�FFcy�)u�8*)���X���#R[��\#{�x;�x#�i�f�E��s�ܪs�(=Fu����9�
��ZZ/����*ߝ��~�9-pש''�(���W�����	-f�!ﶽ���B|Y��ݑ���>ѥƛ�A�*�䦊W���4Xl�
����5��^���̏G3��v�T~�9d�`�|3�*FTm䓃%{�o�j�GU���D�L�rBAa����������K���{��7���@1��j�@q�1n��6y���W��:ǐ���K��`�?�����S�f#��c�C�� �����r%:��p 8�4K5��ʶ�r��y�J�ֶlM��a6Ӣ���SǴ9�ľWܳ$G���
�4�������\��
��+�l���xg�'逖,y/��wA�l�3)�t�T�بnP���ο%�f�II�I �"�?��Y��G魌P��-V��X�	Y6J�9]�x�{���CZh+_�E��xz ���NIS�v��rVI��"j�傿PB�N3HR�3?sa����x�FKOXgܜ`��� /&~�w�dJ$�D/Y�CS[�y�.��%*3��M`���.~;ٵ��I]^aAn��Y���+$�vQ>��#�9J��������e��R��x��Z��M=��I��;����q�k�l�f�m�k�O��`��q�_�ӈ�A��n{��I\��&~=��P[��*s�%l�T�А��=-�QUX?:&B����a��a�>(�T���!'	�D�D��p�^X_fT�0 "��q���`�z���ݻ�(������BiY����sX�Ӯ!N�aX9ʳ�-O_^ø��>�$6Uq��>�_�}�+��M�H��F';`�?���Yf��W���[�x�	�"=9��>re��L��
�ؾaa�@�6��Џ���D���E`	|Fz����!W�ژv�r6 ���k	��G%�l�HJ!L�Ki�\> �k����Ô����Q���!�h� J�	����2�B�y�7����o�������2��H_d��0

���J�y�t��t�ɏwq2��Bm\N^���)[0��VW���-��PGc ^_�>U�΄f�0еΔj��[U&�H!�LSSt��<V03m�*��=��逫�0���yhK����2�׭��D�G��Z}��?��d�fH�"&��-!P�9>nxgm�H��s�<�}kM5�
�����EߠOqʛ���|𳈧�YzQ���63��=�����c!Fl�Chŝ^�ߞ54\b��A�3(A~��H*�qw�~qV_X|F�l^
���X��d���?�*�/��">��w��x�&k8ԟ\��؛ �����>����v.I�yhI7��E%��+t:�p�Ѱf��/�6��0.�a�h���߅qC�>ǋ����ߖ�����\�1��-)��[��F���. ?���Ob� �%����HtC���0=���*��"�h��Na�, ^�<`smcESD�"woy���}ں��Wϓ-�B���|��nfD�m�^��࡚n �l���ܸIU|�~��qW[��X�k\$��j��Re쁊�Q*�ksF�@�(NĄH��Y���}�ÿv/us���V�@@T�F��r:����B7���EI����WҀظ�L�|
�p���u+���� TF_��Y�7�Y1�l�a��ߒ�x�65Dúk�LL�i�j\���<;��,By+wb}١7������t��������qyX�cvt�� �]I���K��L�A
�sè��h�(J'��!, Q���Č�?�j}�anf��EC��(�gB�Do�3��	���D�P�#����>�yxX�~}]�$�r�yp�&Z�r�D�� əu�\�ȗ0�H�c�=Ԛ��N��+�T�M[�(��cD�v`��� ��J�[����Zb��x,]�z~�v^*�a���Ko���D� �����+O��b�烝:'�Zb�ג��m�ՓG6��9XnY.�6ozRR�H��m�7lt�-L��h���Hj�D$UF��y�V�T����6]�bi���U���盜����htw*��k��R5�V񪴘w3�hsɒ��J����}S����'���(�>(�F��4�J@b/ϰx����9h�$'�ve��l�=)��w�ʛ.�j${��}>;��ek{�M,�
��S��vg���0tG�����&�&
]��}a����瞔9=ܾ��%k�"�$�
�6��d�)��}��$*��(�򑱭���2*]�3K��"�����|�Vi��[ך2%[/?�=� ��J��Z�SQ�6M��+a����m�_(�>��e��>׎[h�v�R�c��%ٲ.,�(�2��C�%�	tZ&�^�����	yl;Y6���Z���1�My$ 5K?��p!�e&-΃D��K����~O���%�o���S�\2@� 3��c�)�=+��M97�/�5X�O�hI�� �v#�����RvY���d�&yb����� `[��LWCh��@����F�ݗ�
�?Ha�	%TXXd�R���o��}��~�� G�]i�{h�Mբ5�:��v�Q;�Ľ�ְ�y櫘E��N{��cy3u�`%�S1f{҆Y5�{;6�nJ|ʻr�5}P��C�Z�ۛ���t���Z�cV+v�Q

ҫ�oW�8}2seB���᳾:���Ba>�j��
���*���([��f��,\�v6*��6��W�(�h����Bi����V�k����H�(�L"b�7r[з�w�*�%	i�.�� "�lj[�($��]<ˁ0�����I1`�����{�N�"�����&R1�j��¨��kIH���z^��fC�����\��a#Ahj�+}�QIRӀ�@�c#�����dg�	�檴	S�[r��?����:��7:'���"�ڭ���5F'��b����\���hT����D;Q�ǅQ����gJ�ʱ�e�ٿ���W��\�S��R�� ��0k����E"�s~�f�.ߝ%�j�ܾ��XD�s�O28IZIH>��L8T�ޗ�/r��5��A%yΘ�*�@N\ُ�d����Bs��ol��ɑ�j(�t�x�;�4R���]w5jn �;]��t%!l�P���\���                                                                                                                                                                                                                                                                                                                                                                                                                �,_�R��N<��O�R�t����    �               �Ǐ�˃�[����ګ)h}���S�ӃNQ�[��Վ��5E�d7 vڳ��u?)[ <ˡ�҂Ja�o�T�<�����qI��fwY3��/�B0L��4�蕪=@y�&�<RJt�n����fۦ5�W�yrʒҹ��(����F�Il�J�>۫~eb����y��n���ej�ByRD�w$�#)�H����pK
.j|����k��'��{�B
��[n�p��l�q�{FR��p&oP�j��v�߁uC̃�)-JI`�"f�3�)e�a�ĭ4ͣ���ϝSR{��;�b"t�r1m_Дrf/;�t�,T  �.]v�jRb�'H�h�����}�Җ�W�/�Auq�@Ȭ��5Ñst�M/N��>]9<�5��au��i�Ȩ� ��x������׸|I�/�MU�I�pc9�;�=�(A��cF��!��M��_�w���t��-iQ���&�,���P�	&���1=q�h���iH��t-�CB旺n��JQ%&��P'��a-NC`����$�va��}w        �T����ʑ׵yA��ˁZ��`����x�ܥP���H ��jI#��'�G�O��9s��9%10d    ��G *7�o*�~ؿUQ�4�f���p��rE�I9g8���?cܲSWuM.���|"3 Yz�~�?f�v�-�6��K��hg{`D)�jt�y�h�U����!o��!Y28eE Kk�U��SRYB��
T�|�m�#	@O�e�#H�"�z�l������`�v���o��ieV)�[�B�(ǚ���E6ф���/����e�#s�oHܯ�/0yf�X�PN���I�� *ȷ���O',����(pwz��<�?��5�?�D��9^}s�������K�G����g�������&����� ����1��f�e�?D�L�kڔ�#�ֶ���F�8�MJ�K���ٿL�Q^���������ѧ*6i��c�Ӧz����ʌg.���N�q�E�8�O���,Ĕ�+lS'��8�
b!�U)x���g�@��~g6S�jqd�^1ǋ�������c��ݰ�q������[��9+P��d�`m��0�h����ݺN�#�U$	[.hD�G&YUc�q�v3���c�8������a��Ƒ
���2��,�颇n�'�� ���;H�1����CM(�=F������l�ʾK����5�B	�]4�#�­Q�-�~n�LY���hD�7�p����s�4�
6S�̿.����G��F������4'�n5�?�Y�[lV��;�
�h�j�+��w��~!�up�-(���Z���'_kc!QJvPke���sH��A�
4�-?����H��"w�.�bs�� ڭJH�wB,�0u�2��Ֆ��B�yr|(�:VTè�3����
�Lf���ig<�?v�>Ђ]}� o�.��~G�˙�	��:�@s$�1[EB�#���h��+9�%�B���tn�(�'r'G�m��_0��y�"Ȭ�Z9�{)���"�\R����s�]R�|�^�
I��e ��Y�!$��6ҕ���	f�BT������=�U�At�i ��.��؍n��k�oy/\!���1�����5���ZB8:~�f1\�~��X*����ذ���2}�?ɦ�R>,r�@!�P�4��|K��O�q Ԇ�Dq�:yuj%2H�7/R:�u˰�;���J��[y�.�������l��E�\v�G)9�Э�4)��H��*�I���W��J�Xp[�-斓�뢰I(�}��P �)�M$��~��W�����e�KV�Vh|O��WȅZ#��[cG�fB0wQ}�p�Ҡ=��Mm+`ݬ2=R=$ˬ����ŝD����Ӷ���5j�� ��BC��~5�{dz� �3Tf떶�r�#>6�M@uYX�I��&K<�񭰃�c��T��B�S<N�e��e�%s��h�b[w���z�W��pK�@�ѵC~�8ʵ{�g1����2�l��AG
���?m�#��Y�G��a&�/�j~��ි笘L���؀�GL�_@x��Ɂ�Sh�����dm6�跊N�G��8�,��/tj��I�s�\?���U���iK����~Mx�˽�/�nv�Jz��|Q2m�7��M3����i��\���ֹ_�	5����~�f�}ՊE:7R�)�ڻ8݅�z#'1���Df�EŦ�5�J8s�0� &�c\�{ԗg������0F��(��5�ǣ�B�3 a�����C�:��z��
=���d�|�Az���Sb���75�:!�@୔>�Ⲍ�t��wD6��NT����"(*>.[���}�}�T`"?�`�r%\�z���2s�>~��7�����{�@�]�3h�� q���E�F�T�⎣�t�������lWn��X�p�c��hЈ��>������������9�J��5b�&�-�����$t�-F:{mO���i��v�g�/F%�Y'�{�>]�dO7�WW�-��/�N����Ζ���0�1[����N��U���%V���ﳟ�����h���'}D�E� R[�{F�ـEG�$}�X���0�F��\C,*3jqt����Z���j]�R�00��s�&��9�����GM*+jZM��|�G$/�5�w�K��&��t��Ӧp�<<h^�- $ے��N��ĘX�n�|  x@0]�]��F4U�0(���W�gW�8 (��أ�W�}<ߎ|5�7v��[v�>�~����_��N�,�ܥu����u����r-A��Nh�戚��[��x�Yה₣-/Fx�#_���;��+��ڐ��@G~DVX#�l ^�|�}�N�%Z����`��Є�͒���l_��aڔ3W����z�����K�{�Bq⁽rWGd00�q���%2�ӪBg��[[��O��\+��An�����^0Ð��Bv������!��Z�'�n�q���.n�H��_���[����K�B��yTG}Ű��QD���p�[�>TC�]��F�����/5����<΀�2�׳�d�o|����=�߁6z�Бl��>�;�7
P����"e�hsT�M��n�s}I���/�Ž�                n�@ �WA �XA         eYA             �  O2  A#��� e�-��s5��|�h��'t�j��*�;#.(��+���s��IBl��s;�k�uz��uh]��%�W���{�7����������;��WD'�µ��;�`���G�E>�3�����i����sC�cpڻm�8�DI��f3�-?FɣR�Ѵ.Ye���+� X��MH��zU�s��n�m�RZ��f�k�(�pz���c�� g3����wO��g����l_��\�8����L�m�ن[�@Ķ�+��S� <�!��4�U����{����W��"A\�˾�%�� f�m�ώVB�)��@�R���~uxd�Sފ��e�e03u�@�zP�Fsߜ�i8G����s@|x�d~���l1㕠N��v��\�k�ֽ�&4�ܤ��f캎�"��?��}�B<o@_W��ڡ�Uҡ-�����HR�T���e�q�,���V�)7�	�U�\U]t�j!�E���j �5lR�v=��:ԫL%o	��D�w,�q�����
9m5����57ǆ�ʭ�����S�b�3�3\l'z	�-J�A��Kw�`��L`��OR	<����I�M\��
I�3"z��{|"�![J�����1�Nb��n/�BS>����6�~�.-`ayf��l|z#Nn���#��w̨�
��GM�!ho�l�Ɓ�$2�	!�A���Q�!0�j� ƋdP��QN����$�����9n�h��ko�Ga� �)4�����k��L��6�y��F�Z܊���j�ă|�2� �ը��͉��/��MR�4��
P+%~V�}6�QNK��:q/B���ZH�l��Q2ަp�bCi�~=͝�ی�Y�5�
���ŮQ8�|	)$u]L�Cn4�)�c��9,z�̤�����g��5_�z��Lе��om��De#Ǖi��Xx�,�w϶� Sn�:E����)���9�oo�Ee^P�'�-͸�"�=���
fu��侁©��R����dZ?+���2x�}�oA�>��OG��4����s�[�\�
sʨ��'�bQ�ڴ�W���^ͬ�ͧD�%Giݪ�+�_ƹ���k#(��ril��M��ڳUQ������QDJ*��a.\ڃ�G&ļ��~�q#	�6J��SX��S��6�]D�(������B�q}c,�̓��%$�Lp��w�u��B'�$��pT`雽�3�O${s�~Bp*���R�������\)4]AR�����wՁd���YjԪbxi��k�r�/o���W�s�����,�ٲ쁥ϗD���(�U�WY�1��`z�����aӎ��`������4��By�a���5]��~+��1�N�vH�Xz�cr�W�+o�IK���0�o&���d)���U�| :�G�cMr�ò�|x�V]�PZ����M����p-�3c��B���FB�@񾘸d���CP�J���h��ϸw��#|�=K���;SG���o��}�Ts ��h�_pie�$�"�9~�O��M�6��g� �M� �m��v٩�Lr
`����;q��w�(�����H(p�+5�|Le�:^&��RnI����ޅ�j��vÕд�ɒ)���ǇYG2q��;DS-?� ]1���cR�p%�)��)�Ǫ�s�RVד�A��R�M�V�7��C��kQ�Y�abq|SV`��B��q��%�2־���4���]�b{�5V��sL;u@YJ�����T���6��o�pC!ٖ'��\��<L*��{�"����F#]�oԘ������$�J9X&չ���Lj^C��p���8@�"�b5p��r?��7��2]���+����2��e�I�r�R��[���?��a�:�e�&i`Fe0��,y��x���������~����~S�(�x�(��(
~~Hڔ�I�]�mV���=jX��B9�/h=��&%G?�x)>�@�M0_��$D�����hw���oI���D���T5.׭��ƀ�T?�?R� �^�џ�|��׸�4e4�~��F	1Ǫ��e��2w�Yt�w��p��~�x�]Z��|%���*'H��6��{�3[����g�U��l}��B�)��)�xM���hU���K����6�s�{�gÀ[<����ae#U#o<�<V[Y��k�N̹�D-C	�&��i_r����k�L�;�\w9ƈe~�%��2:.ű[�8�]�I)х���
���"2��[��k|��_aōB�lU��6�� �����]@t-�H������AcqJѷ���i��FK�;{sJ ��`�7���� �y�A��C{b
q�\f"V�����@������v0C�s]�"�M0�I��XF�m�H�˳{�!����-���}��ݧ�E+�|֜y��K��R��`]��
�����ktq
aӘoւ�L,����}g��׃�<��p�m�G��`6|�Q�Z_�NSIs�G���nM�A��~l��e\���3 �M�)Z�}��v͢1}�̎N��ލ%e�������|z��4��X��e�p'*:48Ɉ�I=�p�c�RJ�]�f� ��'(Ż����>��+������oz��&�d�3B�S1�T��wΤ�y�@8/���4� ��Y|k2��t���6d����5��(������ǥ�6.�R�;�d��;sĜ;���� �k�֪��~^�ā�f����`-���*G)�_�7���6��L�GƘ(�A"u삩�	P��������[��/E%��R�(#��pn�lH�	"�1���\%mG]x��9gX�͒n����'���"���*�4���� +�(���x�g��͝�Y�<�p��� �0��a�pS�~��ҡ����n��� x�v�&���Ρ�4�i�S
ML�WL�v�9�h�>�8x�i���}p~��l옍Ob��s�7
Ov����Ce�yⴻ�<9k�L`��Ĥ4ʏ�ħ�*�'�Ӝ���S91U��:�ۖ.1dJ^g`�rF��ê�����e��E�t���0������=�pծ`2����S����+������ܹ���J�K@���Z,��U�\H��$���B^^=͸^�l�h�
-�G��C�D���H�T�&ц��@�Bk(�(��&�Vs���n��u^���ƥ�״V�)jDXꗹ����GK���g?u����h
#�!:�r��T���ѭ�8H���:�](/ �G���Ͻ�������j��7�3�NdA�?{��C%��9�.!©�K4�+k��s�RB1E�>q~��D���E���7�4���	=r�����J�5�!]Q"Y�K1���¤@�s����`ʳ��M��,�k;�U���qL�����h7�g?ǔdwH�z��qpP�o����
!`-���71<4�b��;��o�����j��i27����$�	����~k�Ã��Y��;�+���������%H�t��$Y�+�H>e�Y�)�����y�����U���7,S��5��;���?Rܸ�?7�*�"s�0�u��}Y
� E8@%�"���H��*0�����mk9ɒ��".�~�b{ipB����I�RϮ��ٔH�i�^lP�E 0�J�S����u��8����G2壔5��W�]�8w	�����\���a�7��)%jՅ�|ℱ�w��ί��F�|C�ٻ���jޛ Xd���A8qȻ�DLե��I���ݏ�JĥW&�^}P���O��-��[@R���f��7��g1��J��i�P�6~��(��4w{D����Q�|��Q��W ڦ�?	z��nh�n8,�W����,=�i���`�g�eTX��±��\Q�p3�I�ӽb�n�EJ��d�}F�B�P}�dL^0I����W�2\�5��,v=�c`t��~��/������@6�g�@j�V�F_��L������*[�&�m-��r����Sk%Aeб9�do¸��G\�EJ�6�$������>Ԍ�M��Rϲ�ߖ:C^���Z'G���d4�K�k���0": ���u �3d�� ��K��E�
�ac��^hB�n���u���}'F�l������G��<�p}�Q�kvQ�����Zr�)�'�X(����x�.F���+FeK��Ř(h�u��Z�@T*�Ǭ�������'��2�yOx r��ϛjt�qmFa� ��3Ǜ�������OO���v)��QXk䱊W>2��9��u	5��5�#PV��UE�b�=��%27�j���ݷ�����%�vwmH��L����[�N��|BuE�NZ7�"����o�o�[ny�tB$)k�&�� v��Į��	;_�נ$5�(�c)V્�`�!����Uxr�B�nLb��jScIs2C�4"��X�����Ia��w�o�V~Y%��1�:&N�8�]�4�L�ZL�.�ݰk��v6���?i
���4Y�����Bc&if)�����C�yy�\�܂���^oW�$���	FH�	���
@kW�M�}^"�^=�����h�3bi��ܫ�k���N@���;�;w\��f���y�:�PKwfQ*�� 
IiH���x/O����Z-�6^ĒUf���~�P<ļ�Z�K"�E}w�j���=!��N�!u�e��?%�n�m�|���z�O�)x(��8���ZւP�i���lv�����
v�޷�j�RtN���﬏ZLs9 :}��|q���r� �1���_#��]�����iXur���-��`�<�����&|�<���F�K�7K��,s0^ַ�egi��p'��6�;p���s@�-��*�¢N�	���y��0�[�I���3Y1`�
��aV_=[w��C�fa�XRo^������ܫ	H"J������]`�H������@���p]���.-X�2z��C���IOJ�$�1��ꁦ���&���)���D
4�׎MsZ���k�\�Zw�%����ev�rj�m�E��o$���,�eM��0��bS�cōe�/#���㡟W$Z����,�Eax�S�B�A��K8]�¦�,Uӫ�dz�u����}�S�}�	(��=aP�kZf[;(J�� P-w���*b�! ��\x_~d7R���utM)MG�wGy��"��������o��C_aV��W��>��b��1
c9�U�Kr�&`���Gpi�� n����&����+�̝b��r������̦�tRm^8P����-�<[{r�H� u�>��"��N@���Pt����N,I�vo�k�#�!T+��\T\#1���lƠ?f���Ç� n44˙*y���2R��P0}�_ ƃ��ɜ-"�d0.0��U�gpQ�*:�D��F@�B��ix�Z�~p�Y�=$�p���q�ʉ�q�*�O��|:��<���8��P�n�nF/�џ�i��\9Z�����(�b	�_��Xȼ�z÷��Ș�d�9��-�(��	�����D�kiY�o���)��P4:��|�sB����ȟ�Zdr?�O���<�!�lnYC�X�M�Ӕ                                                                                                                                                                                                                                                                                                                                                                  0  �   d �   �  �   �0 �               �  �  ��  � ��  � ��  0 ��   ��   ��  �	 ��  H �               	  �   � �           � Ȁ         �H    S n v   w e u    M S   S h e l l   D l g       P    *  ����� Y r i .         �P    �  �  ���� R n r       @    � ? I  ����� N n l i y g t h .      �P    �   � ����        �@     � � . ����                      	  �  � $          � Ȁ    	     ��     A o h t o h e   u t t s e   v p p o e a r   s r t n h    M S   S h e l l   D l g       P    Pb $  ���� C m i i s      �P    } h � W ����         P    k H �  ����� W e l a a i   a t p w y r o h   j h d .         P    � o �  ���� W t a i a p   f t r o a          @    Z � + ����� S l n t e r   s e a e t .      �P    � $  x ����         �@     m �  ���� Y d e r e t         P    �  �  ����� O h p s v h   d e n e t   d r n   b t d r m .       P    �  e  ����� A a e e   o w w e a y v   r e e l .                      	  �   (          � Ȁ         b     H h p u   r s g o y a    M S   S h e l l   D l g        P    � � �  ���� O l n g i   e t h r u       P    ; � �  ���� H h o a i t          @    � Z   ����� D w n   t o a a   t i r t a a a .       P    � ' 7  ����� F o b t i o b w .      �P    d ! k ����                      	  H  X �          � Ȁ    	     ZX    G i c c b   n c a t e a l a    M S   S h e l l   D l g      P    l � �   ��� W s t i s      �@    �    ���         P    *�    ��� R v r s s s n t   c a e         P     � �   ��� T e i e e o a i   t e o g       �P    = � �   ��� R m o u o h h s   o a u        �P    � � [ ^  ���        �P    �  ;  ���         @    � � Z  	 ��� T l i h   r e e a n        �@    $� (  
 ���                      	     0 �           � Ȁ         �p    T r s r a n    M S   S h e l l   D l g     P    Q\ S   ��� O s m c h       @    �  �  ����� R y r t s i t   t t e e t i r u   p i t e o f e .       P    �  �  	 ��� I s i y e p a o                      	  $  4 d          � Ȁ         ��    U t h b    M S   S h e l l   D l g     P    F-   X��� A e h       @    V j z  ����� A t o e   t l l   e o n e e r a s   i p a e .      �P    d6 ! Z���        �P    � � � � [���         @    A� -  \��� N w e g h r         �P     �   ]��� S o s r h i c       @     j�  ����� O a e n i t f s   w e d s r .                    	  �	  � �          � Ȁ         @    C z i h l a o u   s l i r   m t u o    M S   S h e l l   D l g     @    � |   ,��� N m h a   e h s l n a       @     0 �  ����� G b a n e s c   e w w .         �P    � � "  .��� M m e t s      �@    l � | K /���         P    �  a  0��� L o o      �@    � a 5 K 1���         P    w  %  2��� W m d y n o a r   e e a        �P    { %  $ 3���                      	  `  p �           � Ȁ         J�     N t l t o h f u   a l a s s o b f   v h m e o    M S   S h e l l   D l g        @    � �   ����� E q i l i d t   b a i r t k e .         �P    h � �  	 ��� H n e   e n d s o o r u         �P    \ @ �  
 ��� H d n                       � �   : �   � �   � �   � �   � �               	  �  � n           K e s e n   e h n n s v l s   f e r   n d o . W E y s d   r g e a l i i w   u m c s e e c i   e t u u h e i d   e f h r o l t   n d h d   w c l w i f h e   d r i m m d   e w m u e a t l   u r o h   e h e   l r r   l o s ; F E e t s d h k   t r o e c d o g   t a m n e o o   g h e u d   i r h   d p i t w   v t m w i   a e r a i e d t   t n p i   s u t p a h o r .  O r h t e c   e f e   r h r n t p e g . A E r e   e o e f a   u t a f r m   h p t t u   s e s a w u c   a n n l e t   v v t g d   i o l t   e y t   n l e e b y g   b a o . C H r i a h y o a   k a n s t o i y   e e t n s n   s e l n   t n e s i h c t   n o u d s e   e p e o h o   t e i e   a e i a r l a h . 9 N h b   e a a a n o                                                                                               ! E m d w n   z o o h c   e i t   s m v b l e a o   e l r w v e o ; Q M n t   r o e o s o w   d r r f   e i h i h a g   i f w   u d e j t   e h w t   a a b t e n a l   t a m h e   i f t i e i f   n m e o w e   a e p   t s s t d r . : T y h t r h   s f h e g a e   c t l t n   a w m s e o a   n e c t e t s   w f t e e o s y   t i d r g e   m a t g ! Q T t e s   c e d n i a   h f u y o   a n z n f o o   e l a   t o l n r i s e   h e l s   b e t r e e   e i c   g s p   e w a d r i r u   s y s o   a i d a a m d .  D e t   a i i   r h n v w n   e n i e h a c e .  A e d w i d !  A i f a h n .                  	  R  b" �          E D i d i   t a e e   n a e n c o   a m a r s   t e e g   o o c s h n e b   l i l h s   s h y   m b w v p s   e h s s f c   e a t t l r r .  O b t f h a   h a l   t k e n w t e i . a T e e w d o   d n t l r   a l t t   r d o e r n h u   t y p   n e s t r t t n   a i i a u s   n i h m c   i o r   t i g   p t e r e s   s u o c i e w l   v e n   i u y i g o   y i v n o i e e .                                        	    $ �           H t r n e e   h s r t o o   w o i   n t r   i r i e s !  I a a h m w i   s n e u p t   a h a . I O e g t   l y i   n u e l h y u   e e o o   n s w o n t o   p a l h t   e i e a e w s i   e r a y o o o   a n n d n s   t i t w g h h r   f l d . 6 F d e e g o   l i a t e e l   t k g a n p l   a r h i n v   d l b t   h c t   r n i l h r   i u r   p l t . A U i e u i t   d r o n o   y r t b   a i b   n s r a n s l i   i e i t h n   h i e r p   e o h r n n i x   l n t h t y   t s r t .  O d f   r p t d h o l   i i y ; ; U t t   e e e   t d i   e l s n l a u   m a e e d h   t o f n n r   e h l n v o w t   i e i   d e r s b   p a d f e . & I t h i   d r t n n n   n n e y   t r m t o k e   u n g r n r y   n a s w . " R t c n g o   h s m n i g   i t r a r   e e h r u   t t k t e w b . 7 W s e m e   d t r i f   v m g a   f m p t q n e   a l t   f y r n e i n   n u t i n a   l r n y e c   i i c .                          	  �  �' $          M S u b f v   e o t e s l   d v r u r s c n   n r t   t s o y e s i   y t n s e w   e o h a r   r o u f i o   d h e r   j w i h t e m n   d h g d c a l r . 6 O s l w   r o e r s s y   e d m e   h c p a e e   o l t w a d k i   o a p d b i   a e l   v a i b o t e e .                                          	     ) �          A U o n n e   e s t d a y   w e n n p e i l   w r c   k r v c f   i e d y a   c b a t e r   i f r v s   r h o e h o   a a a d r h .  D o w   d i u p   b s s p   o b k w k o   s t e i f i t n . T T r n t t h   h e k n n n h   c e t c   y e e i n c o   n s t o n r a y   s t s e u   i r b e d a s d   e i o e h i   c e h o   y r d s w s   t e r p c a e   o w n h ! " A t e   g e c d a e n   h e a t r i n m   i v r e c k f d   m a a . - E h i m n e p h   i t t t i n a i   t a w e t e   p w t s g g l p   t b o   n c o i u y .  S r l l h u w d   s s r e y d   i o r .  N s w   m f n v s h m l   r u l n o i . b W h t g   c a l   c e r e r a e h   t c l r   o o a s e   e e u i a h i t   t n e r l a   e n u r   u r r n s i w   e t v e u   t o r n e s   n n e r p s   c o e a t b c   i n y a o e r   p h w .  R m v a   n h a   d c o n n h w   f s d i n y a m . R T d t   t t n a l m l e   p e g   f a n i y p   t s i   r e t d t i p a   y t s o   i t o   o e t o r e   a w p y i f i h   e h d a e a s   w e e i h   o s h a s . D H s i p   c a e n g i t   e y k a i r   e m n a i a t   w y n a   a i v e e d   s s e n s c c   t s f i n h   s w d t h e f l   t i c . Y R g n s   h o r   n a h u c n t   d o a h e m h   n c h o v r   r l n d p b   n h a   r s u l i h   c e p e   w s r   v g n s o e t a   a r o i e y   d n t a f r e   n a o h n . + A o h h s h d   w p i z o   a m a t   b h u   n t f   l i s a n b n   d e e r h h p .                    	  �  �. �          E C t m t a j   e e p e v   o o i f r a   r o b t i   y e a   n w e h l   a o s o l l   y s k o   e e n i s h l i   a r r p   i o i t a c . U H e t y   h t o   i w o r w c   t q t g c   e t i o v   i n a r   a t f e o   h h c s e o   f t a u s o   h i c f e   r m w m s e i   b e a a h   t e d r   a h d a t i . ( Y h s   l a e e t   d c r e a i   i e i o n w s   n a p t n w   a h a n s u n !                                           �  �               	  �   �0 P          (                �                        �  �   �� �   � � ��  ��� ���   �  �   �� �   � � ��  ���                       �    ��    �  �� p�  ��� ������ � p     p    �    �                   �����s������ ��� ��� ��� ��  ��  ��  �� ��������������������     ���������� �������� ��$�� �� ��;�� (�� /��G��	A�� <��C��V��O��	L�� C��	^�� X�� K�� W�� V�   ��, �(    �� ��  ���� �� ��%�� ���� ��+��4��3�� '�� &�� 2��=��J��<�� C�� B�� O��I��R�� H�� D�� J��g�� Y�   ��  �     ��  �� �������� �� ��+�� ��  ��	0��7�� +��1�� 9�� 9��	C�� C��K��T��G�� T�� V��Z��[�� [��	c�� O�   ��	 �    ���������� �� ����)�� ��%��(��;�� /�� 4�� .��B��S�� <��[�� H�� F�� J��Y�� b��^��p��e�� k�   �   ��     �� �� �� �� ����1�� ��!�� �� -�� 1�� 2��5�� 6��
=��H�� E�� J�� K��X��M�� T��l��n��c��`�� e�� a�   ˶ �     ���� �� �� ���� �� �� (��/��?��?�� 3�� >��	<��3�� D�� M��J�� H�� S��H�� L�� [�� c��	u�� Y�� g�� t�   ��- �     �� ���� ��(�� �� ��1��<��-�� 0�� 1�� 6�� >�� B��D��A��
U�� <��R�� O�� ^�� ]�� j�� o�� S�� c�� X��k�   ��  �     �������� ��2�� %�� +��	.��F��A��6�� 0��O�� C��L�� <�� C�� \�� P�� W��v�� `�� q��_��	k�� d����� q�   ��  �)    �� ��&��$��,�� %��	3�� #��5��=��G��>��<��H�� >��J��Z��]�� R�� e�� d��k��Y��
g�� n��z�� w��x����   ��  �     ��%��$�� $��6��2��.�� 5�� 2�� 2�� 2�� 5��Y��L�� O�� T��T�� C�� \�� g��]�� g�� c�� g��m��p��r��{�� ��   ��& �     ��
&�� ��*��3�� ,��9��-�� 2��@��L��W�� G�� H�� D��D�� P��X�� Q��b��U��|�� R�� ~��u��f����������   �� �     �� %��(��7�� ,�� 5��=�� >��K�� >��W�� O��Q��`�� G�� R��f��i�� l��W��`��|�� x�� k�� }��x����� ��� i�   ��%    �   �� '��3��0�� 5�� +��C�� B�� >�� 6�� H��R�� B��f��P�� Y��o�� W�� l��]����� f��	u�� q�� z�� x�� u�� ���}�   �   ˩    �� #�� *�� 0�� 4�� 4�� ;�� ;�� @��J�� N�� K��N��g�� V�� ]�� b��l�� e�� R��p����� k��f��l�� k�� ��� ~�� �   ��+ �'    �� 1�� *��8�� >��S�� @�� >��	I��N�� I�� N�� O�� I��	g�� `�� [��z��Y������� ��� u�� ���{��������
��� ��   ��' �     �� 1��G�� >��C��G��C�� ?�� Q�� P�� F�� H��Z�� [��`�� i�� a��|�� n����������� |��}�� ������ ������ ��   ��  �     �� :�� 5�� 5��@��U�� ?�� J��D��
E�� H��_�� Q�� V�� q�� P��	g�� ~��s����� n�� y�� ��� ��� u�� l����������   �   ��     ��E��O�� :��U�� :��W��]�� Y�� S�� V�� _�� Z�� d�� g�� c�� f��a��v�� r�� p�������� ��� ������}�� ��� ��   ˸# �     ��E�� F��]��	R��O��I�� E�� `��n�� i�� i��V��j��e�� h����� ��� f�� j�� |�� v��|��}�� ��� ������	�����   ��  �     �� B�� F��\�� Q��Z�� Y�� [��`�� [�� a��R�� v�� f��y�� u�� x�� u�� v����� ��� ������ ��� ��� ��������� ��   ��  �#    �� C�� D��O�� X��]��Z�� Y�� V��c�� q��{��������v��|�� w��h�� y�� ��� x��	��������������� ��� ��� ��   �� �     ��
B�� R�� X�� A��]�� V�� b�� T��	T�� s��m�� x��{��}�� |�� ������}�� ��� ��������� ���	��� �����������   ��	 �    �� A�� X��c�� S��
U��c��S��Z����� o��t��|�� x�� ���g�� ���r��������z����� y�� ������ ������ ��� ��   ��* �     ��H�� P�� R�� \�� b��[��l�� a�� g��y�� s�� ��� �� ~�������� ��� ��� ����� ��� ��� ��� ��������� ��� ��   ��  �(    ��c�� P�� \��o��c�� a��r�� s�� o���� ������ ��w�� ��� s�� ������ ������ z�� ��� ��� ������
��� ��� ��   ��  �$    �� U��W�� Y�� Y�� g��t��i��x��{��`����� ���v�����
���	��� ��� ��������� ��� ��������������� ��� ��   ��    �   �� e�� ]�� b�� K���� g�� i��|����� p��v����� ���{��z��x�� ��������� ��� ��� ��� ������������ ��� ��   �� �    �   ��x��	T�� _�� n�� r�� m�� _�� q��{�� ���	��� t�������������� ��� ������ ������ ��� ��� ��� ��������   �� �  �     �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   �   ��$ �) �& �  � � 	 �  � � �  �  �  �     ��  �  �$ �+ �  �  � �- � �% �) �  �  �  �" �  � �%    �                  1 �               	   1  0A                   (                                                                                                                                                                                               