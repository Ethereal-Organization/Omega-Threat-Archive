MZ�       ��  �       @                                   �   � �	�!�L�!This program cannot be run in DOS mode.
$       �,��Mr��Mr��Mr�yQ|��Mr�yE/��Mr��Ms��Mr�Rx��Mr�Ry��Mr�BKt��Mr�Rv��Mr�Rich�Mr�                PE  L �?HE        � !  �   p      �y      �                          @    $�                       P�  k   $�  (      �                   0 �                                                   �  �                           .text   R�      �                    `.rdata  �   �      �              @  @.data   �0   �       �              @  �.rsrc   �                       @  @.reloc  �   0                  @  B                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                U��QS3�9]��   9]��   9]��   9]��   VWj^Vh�  �  S��   �y  S���q  S���i  j ���`  �u�E�V�d$  �uW�[$  �uS�R$  �u�VWS��*  ��@�u�u���&  V�#  W�  S�  �u��  ���'  _^[��U��S�]V3�3�;�WtC9ut>�};�t7h�� W�`  9uYYv"�PhH� W� � �P�
`  ��F;ur�jX_^[]�U���  SV3�9u��   9u��   9u��   �u�Ya  ��Y��   wq������ Wj@3�Y���������t������hP� P��_  YCY�u��������P��_  Y3�;�Yv!�������E�PhH� V�`  ��GFF;�r�Ej^_���^[�ËT$3���tf�:MZu�J<;L$}�<PE  ujXËL$3�f�9MZu$�Q<;T$}ʁ9PE  u����t
�D$j�A@X�U����  S3�9]VW�]��)  9]�   9]�  ��   9u�	  j3�Y�}��]��f����  �u���uW�r	  �E�PW��	  W�H	  j@3�Y��5�����4���j@�Y��9�����8���󫍅8���PV�u�������4���P��8���P�54� �50� ����j3�Y��=�����<����]�f���EP��<���P��4���P������@��tLj3�Y��}�����|����u�f����<���P�E�+EP�`  �E�j@P��|���P��_  ����u�E�   �E�_^[��U��QQV3�9uW�u���   ��   VWjVjh   ��u�� ����E���   SVP�� ��;�vxV�c  ��Y��tkVj S�Cc  ���e �Ej PVS�u��� ��t?9uu:VS�����Y��Ytj VS���������t�F�W�QPS��������t�E�   S��b  Y�u��� [�E�_^��QVW�|$3�;��t$��   W�E^  ��Y��   Vh�   jVjh   �W�� �����teSUVW�� VVVjVW���� ��;�t=VVVjS�� ;�t&f�8MZu�H<;�}�<PE  u�D$   P�� S�� W�� ][�D$_^Y��t$�u���Y� U���S�]VW3�S�}��Z�����Y��   S����Y��W��   ��   VjWjh   �S�� �Ӄ���E���   WP�� ;���   WWWjW+��u��E��� ;ǉE�tjWWWjP�� ;ǉEtNWVjWjh   ��u�Ӌ����t-�}W�}�EPW�uV�$� ��t9}u�E�   V�� �u�� �u��� �u��� ��uS� � �E��E�_^[�� jX� ��  ��$   ��$�   SUVWj^�x�h3�3ۊ0�x�P�X�������x�h�����3��3��Չ9�Q����Nu���$�   �L$ �D$<�D$8@   �Hh�0�x�L$(�Hlj�L$0��Y�Ƌ׉t$X�|$\3�����`  ��\$j�މl$Y�Ƌ�3�����`  �t$�|$j�D$\ڋT$`Y3�3��`  3�3��t$0�t$(�|$4�|$,j��Y�Ƌ�3����`  �j�\$�����\$Y�Ƌ�3��D`  �L$�t$ȋD$(j�3�Y��3��F`  �|$43�T$03�ՋD$<�L$ �P@xDP�x�����y���L$8�L$ �D$<�������$,  �d$8 �D$<P   �H�P�L$p�L$�H�T$t�T$�P��$�   �L$@�H��$�   �T$D�P��$�   �L$�H �X(�h,��$�   �T$�P$��$�   �L$`�H0��$�   �T$d�P4�L$x�L$P�H8�T$|�T$T�P<��$�   �L$ �H@�@D�\$h�l$l�\$H�l$L��$�   �T$$��$�   ��$�   �L$(�D$,j��Y�Ë�3���	��^  ����3���j�D$8�T$4Y�Ë���^  �L$4jȋD$4T$P3��D$L3��Y3�����^  �L$$�D$ 3L$T3D$P�#L$L3�#D$H3�3L$$�\$3D$ �l$j����D$<�Y��� ��� ��   ��   t$(|$,���t$X�D$8��|$\��3����N^  ���3���j�D$4�T$8Y�Ë��^  �L$4jȋD$4�3�3��D$��Y3�����]  �L$�L$@�D$D�T$#L$3��\$3�#\$@�l$�#�#T$ˋ\$X���L$ �l$\�L$(�L$$�L$,�L$P�L$ �L$T�L$$�L$H�L$P�L$L�\$`�L$T�L$l$d|$X�L$`�L$t$\�L$<�D$�D$�L$d�L$@�D$@�D$�\$H�l$L�L$�D$D�|$�t$�!����L$p��$,  �T$tωH��$�   �L$@�P��$�   T$D�H��$�   _L$�P��$�   ^T$�H��$�   L$X�P��$�   T$\�H �L$`�P$�T$dˉH(�L$p�L$H�P,�T$tT$L�H0��$�   ]L$�P4��$�   [T$�H8��$�   L$�P<��$�   T$�H@�PD��  �Vh�   �\  ��V�   Y��Y^��t$�   YËD$3ɉ�@ɼ��@;�ʄ�@+����@ �6_�@(т��@0l>+�@8k�A��@@y!~�H�@g�	j�@��g��@r�n<�@$:�O��@,RQ�@4�h��@<�ك�@D��[�HH�jj �t$�,[  �t$�^\  ���U��E�} �EteV�uW��   +~H9}s�}j jj W�\  �FHW�u�D0LVP�W  ~H�FH})}��=�   u�FLPV�����fH YY�} u�_^]�U���SV�u��   ��   W+FH;��Ev+��Ej�E�j P�wZ  �~��ǃ����E������E�����}��E�E�j�E�Y�Ë���Z  j�E�Y�Ë���Z  j�E�Y�Ë��Z  �u�E���hp� V�E�������E�jPV������}����j[�]��Vj8Y�vZ  j0���VY�gZ  j(�G��VY�WZ  j �G��VY�GZ  j�G��VY�7Z  j�G��VY�'Z  �G��V���Z  �G��G���Mu�_^[���̡�� Ð���������W���������  ��t�D$��  _�h�� ��  ���G��}�L� ���� R�h�� �  ��Vh� j
�]  �w��NxF�|� h�� �  ����}����� Q�h�� �p  ��h� j
�]]  ��N����}��T$^�B�����   �$�@ h�� �   hh� �   hL� �   h,� �   h� �   h � �   h�� �|h�� �uh�� �nh�� �ghp� �`h@� �Yh0� �Rh� �Kh�� �Dh�� �=h�� �6h�� �/h|� �(hh� �!hT� �h4� �h � �h�� �h�� �z   ��j �j[  r | � � � � � � � � � � � � � � � �  	    % , ������������V�t$���t��h� PF��[  �����u�^Ð����������VW������3��G��~h� j-�[  �G��F;�|�h� j>�[  �G�L� ���� R����h� j
�w[  ��_^Ð�����L$�D$��t~�����Ð�����������VW�9����t$���    ���+����ȸ   ��;�tOr��%  �yH���@u��Յ��w�G   �7t#�   �3���;�r3ҋ���΋W�B�W;�s�_3�^ø    �w����    �G_3�^Ð��D$������������  ���Ð�����V�t$��tWV������~����~��3���    _^Ð������SUW�X����l$��U�����L$3���;�tY�|$}
�D$   ���V�3;�u�E�   ^��D$��} _][�;�~��3����EG�T���3��3����ȅ��D$^��} _][Ð�VW���������  ��t_3�^ËVB�V��}�D�    ��,  ��t��������   ��uj�����F��H�F_3�^Ë��  jP�u  ������u�F_H�F3�^ÍG�ȋЃ�+у���D$��t
WP��������FH�F��_^Ð�+�����  ��t3�Ë��  �L$�D$�V�H�ы��+���1^Ð��������VW������|$����|x�VB�V��}�D� �   ��,  ��t�������  3���~��  @�D� ��  ;�|ꋖ  R��  ����t��  GjW�v  ��  ���  �N_^Ð���SUW�H  ��� �N���3ۣ�� ;�u_]3�[ÉX��� �   �X ��� �PB�P��� �H�D�    ��� ��  ��� ��p  ��� ��x  ��� ���  ��� �X�D$;��l  =   ��a  P�}������ ����Y��� ;Éiu��� �B    ��� �X�%;�v!��� ��yG�y��� �Q��;ŉQwߋD$V;�~��� H��y@�A��5�� ���N�Ћ�+�H����F��� �   9x}�x��� �H��   ���  ��� �H��8  ��� �P��<  �5�� ��<  ;�~+�4   ��~;�~�A�+�����<  �5�� ��<  ;��9�<  }��<  �5�� ���  ��� Uh  ���   ��� ǁ   
   ��� ��  ��� ��(  ��� ǁ     ��� ��@  ��� ��$  ��� ��,  ��� ��0  ��� ��4  ��� ǁ     �  ��� ����  ��� ��  ���� ǂ�   UUUU��� ǀ�   xV4��   ��� ��=$  ��t���2�y�T|ޡ�� ^ǀ,  %   ��� ��0  ��� �P�L�H��� �A�Ё���  ;���  =   @��  ��8  ��� j��H  ��� ��L  ��� ��P  ��  ��� S���  ��� ��`  ��� ���   ��� ���   ��� ���   ��� �AH�+����A��� ���  Q������� W���  ��� ���  Q�v������ j���  ��� ���  Q�W������ j���  ��� ���  Q�8������ j���  ��� ���  Q������� j���  ��� ���  Q�������� j���  ��� ���  Q�������� j
���  ��� ���  Q������D��� j���  ��� ���  Q������� j���  ��� ���  Q�{������ j���  ��� ���  Q�\������ j���  ��� ���  Q�=������ j���  ��� ���  Q������� j���  ��� ���  Q�������� j���  ��� ���  Q�������� j���  ��� ���  Q�������� ��@���  ��� j���  Q������� j��   ��� ���  Q������� j��  ��� ���  Q�a������ ����  �(j������� ���AH�+����A�
j�k�������� _][�HI�H��� Ð���;������  j�D$P�(  ��Ð���V�����t$��t0�T$W���  3�����~�1 ���  ��A;�|�V�6  ��_^�V�t$��tV�A���V�  ��^Ð�������� jǀ      ��� ǁ�       ��� ���  P�m������ �����  ��t	P��������   ��� ��=,  �D�    |�j �]������ ����4  ��t	P�  ����� ��8  ��t	P�<�������� ��H  ��t	P�#�������� ��L  ��t	P��������� ��P  ��t	P���������� R�  �����     Ð�����D$� %   ����$�@Ð�������������L$���t�T$��}   ���%����Ð�������������V�t$��Ё�   �%���~�N�L���9 uH�������~^Ð���������SVW�����|$��O�K�Ǚ���T$���R�4�u��_^[ËǙ����|�{�ʋ�3���I��u���3��s_^[��Ð������������W�����|$���u3�_Á����V�H��VW�x�������uNVW�i�������t��^_Ð��������������SUVW�d����؋�  ����   �SB�S��}�D�    ��,  ��t�o����T$ �t$$VR���%�����   ��D$�L$������{��N��ƋL$����D$$�ƙ����|�C������Ju��C�T$$;�|)���   ��u�;�|j������C��H_^�C][��Ët$ +͋F�<�����8�D$;�|	�D$BЉV�����C��H�C_^][��Ð����������V�t$W�|$;�t]��uV������_^�SUV����W�������o�v�Ѓ�;�}�ˍ<�+�3��|$��~�͋�+΋4�0��Ju��L$�][�_^Ð��D$V�t$VP���������t5   ��^Ð��������������D$� %  ������Ð�������������QS�\$UVW�{������l$��  ���1  �D$SP����������  �t$���  �UB�U��}�D� !   ��,  ��t�r���S�l�������t
j�.��������%���Ɓ�   ��؉L$���L$ Q�f����E��H_�E^][Y�;]~���   ��t
j���������  ��uv��~7�C�;�|(��    +�@�,�    �Ћ���+�J�8�D9u�l$��~3���+�ދ΅ۉL$~���׋ˋ0���2��Iu�L$��~�<�3��L$ًL$ ��M_^][YÐ����T$��u3�Ë�ȁ�   �%���u3�Ã�u�B� =   @r�   @��   �u���S�\$U�l$V;�Wt_��} �ʋ���   ���   ������$�@;�u?����������;�/}_^][��Å�~ �u�[+ލ��t��y���J;�wrم��3�_^][Ð���������QSUVW�v�����l$��  ���`  �UB�U��}�D�    ��,  ��t�}����\$�3�����uj�8��������u	�C90u3�9\$ u
j�������|$W�;�������uS�.�������t
j����������%����؁�   ���u�L$�Q9u3ۋM�3;�~���   ��u�;�~
j��������  ����   �T$ �D$RP�����L$ ���9 th�T$�%   �3���u�L$ ���tM�_��EH^�E][Y�3���~)��    �T$�l$ @���R�m;ƋT���T)�|�l$�D$ �����0�M_^][YÐ�����������SUV�������  ����   �\$S����������   ���%�������   �����  u.��   �u�D$Pj��8�����^][ËL$Qj�%�����^][�W�|$��;�tG3���~�S�O����@;�|�W��������;�}=�GW��    C������;�|���7_^][Å�~��    �W��H�D�    u���7_^][ËD$PS������^][Ð���S�������  ����   �\$S��������u�D$Pj�_�����[ËV%����t$��W��������  3���~"U��    �[�n@����\���\$;�|�];�u"��~E��    �N��J�D�    u�>_^[�V��������;�}�VV��    C������;�|�>_^[Ð�����D$V�t$��t3����ʅ�t��3����ʅ�u��^Ð������SVW������t$�H�ƙ�����D$�X�ƙ���   ��3�����_^[#�;����Ð���Q�D$�L$U�l$W�|$UQ�   �D$   �     ��������u_]YÍU���}�E�D$�L$S�]�+�V;ݾ   ~P��L$BSQ���S�������tF�ց�  �yJ���BtK;����ƙ�������������D$$�    �΁�  �yI���Au�ƙ+T$$�����   ���^[_]YÐ������SUVW���������  ����   �VB�V��}�D� N   ��,  ��t�������   �~P�C����L$���  �QRǆ�       ��  �苆�  �Nǆ�      � ��%����Ё���  ;�0��;�)W������D$���  PSQ�,   �F��H�F_��^][�j�����F��H�F_^]3�[Ð��UV���������  ����  �l$�;�u�D$�L$PQ�`�����^]ËVB�V��}�D�    ��,  ��t�����SW�|$W��������  �D$RW�������  PW�{������  �D$(    Qj����������  R�������  Pj��������  ��3ۃ8 ~}�P���  Q���  ��PQ��  ���  ���  PRP��  ����u,jj���������  PWP�  ���  PWP�  �� ����  PUP�  �����  C;|���  ��u>�D$��u6���  ���  PQ�&������  ���  RP�������D$   �����|$���  ���  WQR������D$$WP�����F��H_�F[^]ÐV�*�������  ��t3�^ËVB�V��}�D� M   ��,  ��t�5�����   S�W�~P�������  �T$QSRǆ�       ������D$$���  PQǆ�      ��	  ���  ��R����W�W����F�� H�F��_[^Ð��������HSUVW�t�����3�9�  ��   ���  �L$`PQ��������  �\$dRS������V��B�V��}�D� T   ��,  ;�t�Z����|$dW����S���������u0���  P��������uWj����WW�*  ���N_^][��H�Wj�k���WW��)  ���  Q�x�������tӋ��  R�e�������}
j
������9�  u���N;���  ���  ���  �T$ ���  �L$��   �T$,���  ���  �L$$��  �T$4���  �L$0���  �T$D���  �L$@���  �T$P���  �L$L���  RPP�D$$�l$4�l$D�l$H�l$T�L$`�I-  ��3��3�y�   �T��D�;�u�P��GC;�t�l��D�UP�Q�������~���  UQU��,  ��Ku����|����  R��  �|$h�؋��  WP�����������������ۉ\$d�w�����\$d�F��t�Ћ��  �L$�T$QRSP������D$ ��3ۅ�~WWW�x,  �D$��C;�|��~��W�+����L�QW�U,  ���T$�\$d�D$+څ��\$dt3ۅ�~WWW�.,  �D$ ��C;�|�)D$d�D$d���_����F_H�F^][��HË��  ���  PQ�0������F;�t�Ћ��  PjP�  ����t���  WRW��+  ��9�  �s������  P���������\������  PPP�+  ��뚐������SUVW��������  ����  �VB�V��}�D�    ��,  ��t�"�����N;�t.�|$W��������|3�W�Q�P���������X  ��|$jW��  �����?  ���  �T$QR�#������  �L$PQ�����\$0S��������  R���������3  Sj��������  P����������  ���  Q���������}
j
�(�����;�u
j��������  ����   WW�B  ���  WWR���"  ���F��t�Ћ��  PjP�W  ����t���  SWWPPS�#  ����  ��u)���  P�V�������t���  PWWPPP�^#  ��뚃�tVWUW��  WWS�  �F��H�F_^][�W�$  ���  �T$QR�n%  �|$,�D$$���  WPQ����WW�Q&  �� �N_^][Ð�����h�  j�?  ����������u�D$�L$PQ�?  ��Ë�  ��t3�ËT$�D$VRP�n?  ������u
j���������^ËD$��tP�M:  YÃ�SUVW��������  ����  �VB�V��}�D� L   ��,  ��t�����F���`  =   �U  ���   ��uj�F  �D$P�������   ����t��  �\$ ��\$ ��0  ����   ��tI���   3�Q�%?  �����t/���  G;���   ��
t��t���   R��>  �����u�� ��0  3Ɋ������   �N��<w��
ty��0  ��  G;ډ�0  ��u;�  }3Ҋ��u��K;�  u;�  |j�]  ��t03���~*���   P�m>  �����t���0  G;�|����0  ��0  3�3�3���D$   �L$~D�~<w>�|�/uH��0  �; u�DA< t��L$�<-uA�D$�����L$�<+uA�L$��0  �D$K;��V  �L$ 3���N��<v��@�  ��<w^��uZ��/u&���  �|$RW�   �
���W�������3���   ��.u*���  �   P�������  �OQRU���������   ��P��@u_��p��   =�   ~=�   }-�   =�   ~=�   }-�   ��~
=�   }��L��{u�>   �f��u�?   �Z=�   tg�Q��~=�   }-�   =�   ~=�   }-�   ��w=�   ~!=�   }-�   �=�   ~=�   }-�   ;�sw�L$GWQP��������D$K;�������\$�T$��0  SRǆ0      ����S��������  P���������t���  SQS�������FH�F��_^][���j�j������F��H�F_^]3�[��Ð����������SUVW���������  ���  �VB�V��}�D� K   ��,  ��t������F����  =   ��  ���   ��uj�  �\$$3�S�l$����Sj�D$(�����;�����<   ua9Fw\���   ��u�D$(_� 0�@ �FH�F^]�   [��Ë��   Pj0�9  ���   Qj
� 9  �F��H�F_^]�   [��ËL$�D$    ���u29Fw-���   ��u	�T$(�-����   Pj-�8  ���   �l$���  �D$    QS������(  �����  ���  RS�w������  P����������   �߁���  ���ۋ�u�   ;�ǆ�       }���  ��+�PQP�y�����;�~���  ��+�PRP�`��������  ���  �~PQ���������|O���  ���  RP�l������  �F������;�~+��QWQ�
������  ���  ���  QRP��  +�����l$�~ǆ�      �|$���  Q�����L$�؃�;ˉ\$~�������H  �L$(��L$(�\$���   ��u;�  u��  ��;���  ;|$u"�~<w��u�).����   Pj.�7  ��E;�~
�0   �   ���  WQ�������  WRj ��ǆ�       �K����F����<ǆ�      w��0��:|����[|����@u8��}��A��|��4}��G��4|��>}����>u�+   �
��?u�/   ;|$}�~<w��0u���  P���������t0���   ��u	�L$(�)����   ��RP�6  ��EO��������D$����   ��(  ����   ���  �T$$QR��������  P��������ta�~<w3���   ��u�L$(E�D$   �D)�/�)������   Rj/�5  ��E�D$   �
���j�����F��H�F_��^][��Ã~@uD�Ź   �����t6�|$(���   ��u�/=����   Rj=�85  ��E�   �ř����u���|$(���   ��u�/ ��F��<v��@u���   Rj
��4  ���D$$�L$PQ�G����F��H�F_��^][���j������F��H�F_^]3�[��Ð�������QSUVW�����\$�l$�D$��M ;�~ �D$�D$ ;؋�tPU�������$�L$��L$�L$ ;��tQS���������D$�L$ 3��9�C�\$�U�i;{�l$|9��   uG�9�; uL��3�+؋�+�;|$|��v~�D$���   ��t	;x��   ����;�v3�;�s�   �)G��뾋�3�+���+�;\$|��v2�T$;Z~
���   ��u:�9��3�;�r�   +)C���ċL$ �T$��t����u_H^]�[Y�j�q�����_^][YÐ���������SUVW�D����t$�|$ ���;ȉl$�D$�L$��   �\$$;�tSV�����D$����D$��F�M �W�[3���uC��3�+��+�;|$|����   ;|$��   ���+)+�;�s3�;�v�   �G����+�3���T$ +�;l$|��v@;l$O���3�;�r+�E�ʋT$ ����ҋL$�   �	+�ʋT$ �E��붋T$$R�������_^][���j�M�����_^][��Ð�V�*�������  ��uE�VB�V��}�D�    ��,  ��t�9����D$�L$�T$PQjR�   �F��H�F^Ð������V�t$WV���������  �|$W����������  SUV�����W���������؁����W�������V�\$$��s����ȋ��D$(��@�+\$ ���D(��w{�$�K ��S|WV�������kVW�������_��SVW��������TWV��������B��S|WV�������7VW�������%��S|WV�J������VW�>�������D$��}�3   �;�t
��}�6   �];�[t";�t�D$��}�5   ��_^�j������_^Ë�SJ pJ �J �J V�z�������  ��uE�VB�V��}�D�    ��,  ��t�����D$�L$�T$PQj�R�c����F��H�F^Ð������U���SVW�����E��E;Et�MQ�n������} u�s  ��} u�UR�O������Z  �E�    �E�    �E���   ��M�U�%����E��M��9 ��   �U�B�E�M�Q�U�M��t(�]�}�u�U3�����Ń� �����Iu��]�E��}� vH�E��E�M��U�;Q|�E����    tj�G������   �M�Q�E�M����U���E���M�U���w�E�;E�|�}� vi�M��U�;Q~�E����    tj��������[�M�Q�E��Q�U��P�M�Q�UR�E�H�U��P�  ���E��M���M�U�E�뉋M�9 t�U�E�M�_^[��]�������U���SVW�b����E��E�    �E�������M��U;Ut�EP�������M��9 uJ�U�B�E�M�Q�U��M��t.�����u��}���]U3���Ջ�����Iu��]�E���O�E����E��	�M���M�}� |5�U�R�EP�M�Q�E��Q�U��P�M�Q�  ���U�J�U��뼋E�M���EP�"������E�_^[��]������UVW�h�������  ��t_^3�]ËWB�W��}�D� 
   ��,  ��t�q����l$U�g�������t
j�)������t$��u
j��������  ��t�GH�G_^3�]Ã�u�D$PU�}����G��H�G_^3�]�S�] ��   ����\$}5�\$��SVU�=��������t��   ���\$�WJ�ۉW[t��_^]ËL$QVU�
������ݐ����VW�i�������  ��t_3�^ËVB�V��}�D� X   ��,  ��t�s����L$�|$�%   ���u#�u�~O�~�I�u_3�^����_$�^@Ë��  RQ�������  PWP�q����N��I�N_^Ð����D$�L$PQ�Q��������@Ð�������VW��������  ����   �|$W�O���������   �VB�V��}�D� 1   ��,  ��t�������  SPW��������  Qj�������  ��^���3�;�[u�   P+эy��~RP�v������#��v�NPQP�������  �V����8w⋖�  �B���r�����  G�@���s�FH�F��_^�_3�^Ð�������QSVW�����؋SB�S��}�D�    ��,  ��t������D$�|$;�t
WP���������������u<�G�L��A�L$u�C�   H_�C��^[YÍT$RQj j�,  ������t ��W�L��3�A�����tWVW��������C_H�C��^[YÐ���U���0SVW������E�E�   t�  �M�9 t�U�: u�EP�%�������  �M��  �U��E�H���U�J�E�x}"�M�Q�E��D�    �M�,   t�����UR��������u�EP��������tj�P������M�Q���E�P�a  �M���   ��E���   �3щUԋU�%����E�M�������U�E�P�Z������M􃹀    t,�U�U�E�;P~j��������M�Q���E�P��  �M�9 �8  �U�B�EЋM�Q�U��E��H�M�U;U��   �}���   �E�    �	�E����E��M��9M�}J�u��M�+�I���UЋ�ދ;�]���+ڃ���U3�����ŋ,�� �� �,I��u�l]뢋M���}��GGGG���M�uЋ}�3ۋ����Ã� �� 3ۃ��� ��Iu��]�E�    �	�U����U��E�;E�}C�M�u����]�ދ;�]�ދu�+ރ�U3�����ŋ,�� �� �,I��u�l]��h  �M;M��  �}���  �E�    �	�U����U��E��9E���   �E�    �M����M��	�U܃��U܋E�;E�}P�M�M܋U��B��Q�U�P�M�M܋U��B��M�Q�U�B�M܋�R�E�H�U���P�  ���E�럋M�M��U��B�U؉��^����E�M�T��E���M�Q�U�R�E�P��������E�    �E�    �	�M����M��U�;U���   �E�E��E��M��Q�E���Q�U�P�M��Q�E���M�Q�U�B�M���R�E�H�U���P��  ���E؋M��Q�E��L�M؋U��B�U��L��E�    �E��H�U��E�L�;r&�E�   �U��B�M��U�D�+�M��Q�M��D��7����   �E�    �	�U����U��E�;E���   �E�    �E�    �	�M܃��M܋U�;U�}P�E�E܋M��Q��P�M�R�E�E܋M��Q��E�P�M�Q�E܋�Q�U�B�M���R�  ���E�럋E�E��M��Q�M؉��c����U�U�E�M���U�R�������EP�M�Q�z������U�B���M�A_^[��]��U���dSVW�����E��E���   t�j	  �M����  �U܋E��H���U��J�E��x}"�M��Q�E��D�    �M���,   t�����U;Uu
j�Y������EP�}�������u�MQ�m�������t
j�/������U�: u
j�������E���   t�M��Q���E��P�  �M���   ��U��E���   ��M��U�3U��U��E�������U�
�E�������U�
�E��M̋U��E��M�Q�UR�(������E܋�M��U����    t/�E�+E����M�;A~j�i������U��B���M��A�  �E�    �U�;U���   �}�u=�E܋H�U�r�3��6�EԋE܋H�U�r�3��6�E܋H��U�R�������R�E܋H�ŰD�����M�Q�M�;D��s3�UR�E�P���������|�M�Q�UR�E�P�X������Mԃ��M��͋UR�E�P��������}~�M;Mt%�UR�E�P�������M�9 t�U�E��M��U;Ut(�EP�������M�Q�Eԉ�}� v�M����U�
�E�M��U�
�E��H���U��J��  �}���   �E�P�M�Q�P�M�Q�x������E�U;Ut�EP�M�Q�m������U�E��M��U;Ut(�EP�������M�Q�E��}� v�M����U�
�E�M��U�
�E��H���U��J�8  �E;Et�MQ��������UR�EP�������EԋM����   �UȋE�ǀ�       �M��9 �'  �}�t�U�R�E�P�M�Q��������U�B�M��T���U�E�H�U��D���EċM܋Q�U؋E�H�M�U����U��	�E����E��M���9M���  VW�]؋u���ދS�;U�u�������u�r��u����E���;�ru;C�vOu�s�}�_^�U�+U����U��}� �  �E�    VW�M��u����}��]�ދu�+ރ�U3�����ŋ,�� +�� �,I��u��]�E�_^�E܋H�U��D�;E���   �M܋Q�E��D�    �E�    �E�    �	�M����M��U�;U�}e�E�E��M܋Q�M�I���E��U��UЋM�Q�E��M�;�v�E�    �U�B�M��U�;�s�E�   �E�E��M܋Q�MЉ�늋U����U���E܋H�U��D�+E�M܋Q�M��D��U���9U�u�}� u�E����E���M;Mt�U�B�M��U����5�����  �}�t�E�P�M�Q�U�R��������E�H�U��D���E�M�Q�E��L���MċU����U��	�E����E��M���9M���  �U܋B�M��T�;U�u�E�����M��U܋B�M��U���U��4�E�P�M�Q�U܋B�M���R�E��Q�U܋B�M��T�R�
  ���E��E��M�;sW�U�R�E��Qj �U�R�E�P��	  ���E��M�;M�r�U�;U�u�E܋H�U��E�;D��w��M����M��U�U�U�럋E�+E����E��}� ��  �E�    �E�    �	�M����M��U�;U���   �E�P�M��R�E�P�M�Q�E���Q�U�R�W	  ���E�E�E��M܋Q��;E�s3�M���M�U�U��E܋H�E�� +E���ȋU�U��E܋@���!�M�M��U܋B��+M��U�U��E܋@���T����M܋Q�E��L�;M���   �U܋B�M��D�    �E�    �E�    �	�U����U��E�;E�}X�M�M��U܋B�U�R���M��E��E��E�    �U��E�;r�E�   �M��U�+�UЋE�E��M܋Q�MЉ�뗋U����U���E܋H�U��D�+E�M܋Q�M��D��U���9U�u�}� u�E����E���M;Mt�U�B�M��U����P����E;Et�M�+M���M��U�
�E܋M���UR�z������EP�n������M;MtM�U�R�Z������}�t�EP�M�Q�U�R�0�������EP�M�Q�.������U�: t�E�M��U�
�}�t�EP�M�Q�UR��������E�M��U�
�E��Mȉ��   �U��B���M��A_^[��]��������������UV��������  ����   �VB�V��}�D�    ��,  ��t�$����l$ �D$;�ǆ�       uj�׼���F��H�F^]Ë��  S�\$W�|$PSW�����L$(��;�t;�t���  PQP�U������|$$�L$ ���  WQR������;�_[t���  UP��������Fǆ�      H�F^]Ð��������������VW�)�������  ����   ��8  �|$��tPW���������   �VB�V��}�D� P   ��,  ��t����W����������   ���  P�&�����   Q�������  ǆ@     �   ���  �H�    ���  �B�@   ��   �   ��   �W�H�����  ��   PPP���  PQ�]  ����tj�>����F��H�F_3�^Ë��  ��B���8  +ʅ���4  uj ��������8  ��8  RW�����F��H�F��4  _^�VW�ɺ������  ����   �VB�V��}�D� Q   ��,  ��t�Լ����8  ��uj蓺���F��H�F_^Ë|$�D$WP������8  PPW����W��������}��8  WQW��������@  ��tN��8  ���  ǆ�       R�QW�q�����8  ���  PPR�=������  WPǆ�      ������ �N_^Ð������������U���4SVW�¹���E�E�   t�  �M�Q���E�P�M�y}"�U�B�M��D� R   �U�,   t贻���E��  �M��U�8  �E��M�4  �U�E�P�MQ��������U�@   u8�E�P�M�Q�U�R�c������EP�M�Q�������U�B���M�A�O  �E�    �U���EЋM�MЉM��U�: ��   �E��H�M��U��B�E��E�    �	�M܃��M܋U�;U�}X�MЋu����]�ދ�e���u�+ރ�U3�����ŋ,�� �� �,I��u�]�E�D�    �� T�� �E���  �E�    �	�E܃��E܋M�;M���   �U�R�E�Qj �U�R�E��H�U܋�P��  ���E�    �E�    �	�M؃��M؋U�;U�}G�E�E؋M��Q��P�M�R�E�E؋M��Q��E�P�M�Q�U��B�M؋�R�  ���E�먋E�E܋M��Q�M�Mԋ�ыE�E܋M��I���E�    �U�U܋E��H�E��;r*�U�U܋E��H�E��+�U�U܋E��@���E�   ������M��Q�E��M���U����E���M�Q�U���R�E�P�e������M�Q�������U�R�E�P���������|�MQ�U�R�E�P��������MQ�U�R�_������E�H���U�J_^[��]�������V蚶������  ��uj�VB�V��}�D� S   ��,  ��t詸�����  �L$�T$PQRǆ�       �Y����D$���  PQ�h����F��Hǆ�      �F^Ð�U��S�E�eE�� �u�]�[]Ð����U��S�U�E�u�]�[]Ð������������`VW�D$$   �ε����3�9�  t_3�^��`ËVB�V��}�D�    ��,  ;�t�շ�����  �L$lSUPQ�"������  ��$�   RP�������  Q�������  �D$HRj��������  Pj�������  Qj�Ը�����  R蘸�����  3�P�|$d�|$H3�\$L�������4����  ��l$(�\$�|$ ����   ���  ���  ���  QRP�������  ���  ���  ���  ���  ���  ���  RPQ�������  ���  PRP�[������  ���  ���  �D$<��$@���  �D$�0  ���  ���  RUP�.������  PWP� ������  ���  QSR�������  �L$8PQP������D$\��0�����  Pu���  PR�������  PP���  ����  QP�������  ���  PRP�z������  ���  ��PUQ�������  PWP�������  ���  RSP�q������  �L$8PQP�_�����0��u���  ���  RP����������  ���  PQP���������  ���  PRP��������  ����  ���  P�����������  ���  �8���|$,u���  �H3ۉ|$0�B�)�\$<�8�  �H��ҋD���L$$�X�\$(��   ����   ����   �L���T$RSQP�����D$L���  �T$ �H�D$ RS�T��RP�}������  ��T$0�ARS�L���T��QR�]������  �L$X�؍D$@P�B�T$DQ�L��QR�9�����@���W  �l���D$<���  �@�\���|���|$,�3  �&  ����   �L���l$USQRP���������  �D$L�T$@�Q��D$$P�D��T$(SPQR�����L$T��(��3�P�D$<Pj Q�  ���  �    T$�D$<�AR�T$0�L���D��SQRP�W������  �D$t�L$$�B�QS�L��D$,QRP�2�����$�   ���(��3�3�PRPQ�7  ���Y3�SRSP�&  ��D$$S�L��3�鋎�  ЋA�T$@�D$4�T���PSR��  �L$,���D$0�ڋT��3����D$0   �   3ɉD$,�D$ �L$�L$(�D$�D$0��t+����)  �T$<SWRU�.  ���D$$���  �5  �D$,����   ��3�+���ʋ�щL$l��  �L$�    �ӉL$@ʉT$D��  �L$l�T$ Q�L$@P3���PR�  ���D$$����  �L$D�T$@QR�T$$��3�+ʋT$D�RQ�  �L$4��;��m  �   ���    �ˉD$H��L$L�M  �L$��3�+��ˉD$P���L$T�/  �D$L�L$HPQ�L$(��+��L$D�QP�"  ���D$$���  �T$T�D$P�L$RP�D$D3���RQ��  �L$4��;���   �|$$uJ�D$�L$ȁ�   ���   �T$(�D$ T$ �T$�D$(�ŉL$�L$<+�ˋ�\$<�T$�����a�L$�   �+�3��t$�L$$;�si�T$(����D$ �T$ �T$S�D$,����D$ Wj Q�T$,�D$$�	  �͋�+ȋD$<\$<���؋T$�L$,B3��ɋL$(�T$���D$,������L$��  �yI���A���  �L$R�!��������W����|$4�u�D$�D$%  �yH���@��u���  �L$xPPQ�������\$|��$�   ;�tK���  �D$tRP�������  ��$�   ���  PP���  Q���  RPQ�������  WR�j�����(���  SP�Z�����$�   ��;�][t;�t���  PQ�9������~���  OR�~�C�����_^��`Ð����������L$�D$�T$V�t$+��;�wr;�s�   ^�+��;�wr;�s�   ^�+��;�wr;�s�   ^�+��;�wr;�s�   ^�+��;�wr;�s�   ^�+��;�wr;�s�   ^�+��;�wr;�s�   ^�+��;�wr;�s�   ^�RVPQ�  ���� �T$u=   �r3�^Ð������U��� �EV�E�E��E�E�B   P�E��u�E����P�R  ���M��x�E��  ��E�Pj �  YY��^����������������W�|$�j��$    ���L$W��   t�A��t;��   u�����~Ѓ��3�� �t�A���t#��t�  � t�   �t�͍y���y���y���y��L$��   t�A��td�G��   u���������~�Ѓ��3��� �t��t4��t'��  � t��   �t�ǉ�D$_�f��D$�G _�f��D$_È�D$_�U��� �E�E�I   P�E�E��$   �E�EP�E��uP�  ���������������̋L$��   t�A��t@��   u�    �����~Ѓ��3�� �t�A���t2��t$�  � t�   �t�͍A��L$+�ÍA��L$+�ÍA��L$+�ÍA��L$+������̋D$��tD�T$VW��|$׃�t2�   t�:uRFGHt��8�uE�N�W8�u;������u�_^Ëȃ���t+�t'�N��W�8�u8�u����8�u8��    �_���^Å�tċ�8�u�Ht8�u�Ht��  � ��  � ;�u�H_^�����U��WV�u�M�}�����;�v;��x  ��   u������r)��$�u �Ǻ   ��r����$�0t �$�(u ��$��t �@t lt �t #ъ��F�G�F���G������r���$�u �I #ъ��F���G������r���$�u �#ъ�F��G��r���$�u �I u �t �t �t �t �t �t �t �D��D��D��D��D��D��D���D���D��D��D���D���D���D����    ���$�u ��(u 0u <u Pu �E^_�Ð���E^_�Ð���F�G�E^_�ÍI ���F�G�F�G�E^_�Ð�t1��|9���   u$������r����$��v �����$�`v �I �Ǻ   ��r��+��$��u �$��v ��u �u v �F#шGN��O��r�����$��v �I �F#шG�F���G������r�����$��v ��F#шG�F�G�F���G�������Z�������$��v �I dv lv tv |v �v �v �v �v �D��D��D��D��D��D��D��D��D��D��D��D��D��D���    ���$��v ���v �v �v �v �E^_�Ð�F�G�E^_�ÍI �F�G�F�G�E^_�Ð�F�G�F�G�F�G�E^_���t$�=  YËT$�L$��tG3��D$W����r-�ك�t+шGIu������������ʃ���t��t�GJu��D$_ËD$�j�t$�^   YY����������̀�@s�� s����Ë�3������3�3��̀�@s�� s����Ë�3Ҁ����3�3���5�� �t$�   YYÃ|$�w"�t$�   ��Yu9D$t�t$�V  ��Yu�3��V�t$;5X� Ww!j	�  V�  j	����  ����t�����uj^�����Vj �5< �(� _^�V�t$��t=j	�Q  V��  Y��YtVP�  j	�  ��^�j	�  YVj �5< �,� ^�������������̋D$�L$ȋL$u	�D$��� S��؋D$�d$؋D$���[� �D$����   �4� j��� �s  ��Yt<��� 3Ɋ�� %�   �-�� ��� ��� ������ �@#  ��u	�n  3��r�0� �x��)  ��� �$  �i'  �&  �  ��� �>3�;�u,9�� ~���� 9�� u�B  �$&  �+#  �	  ���uQ�#  YjX� U��S�]V�uW�}��u	�=��  �&��t��u"�|��t	WVS�Ѕ�tWVS�������u3��NWVS�������Eu��u7WPS�������t��u&WVS������u!E�} t�|��tWVS�ЉE�E_^[]� ��� ��t��u�=�� u��)  �t$�	*  h�   ��� YYát��t��h� h� ��   h� h � ��   ���j j �t$�$   ���j j�t$�   ���jj j �   ���W�   j_9=�� u�t$�@� P�<� �|$ S�\$�=�� ��� u<�p��t"�lV�q�;�r���t�Ѓ�;5ps�^h � h� �C   YYh(� h$� �2   YY��[t�   _��t$�=�� �8� _�j�%  Y�j�}  Y�V�t$;t$s���t�Ѓ���^�V�t$WV��   �NYx��D$�����V�t$�  Y��YV�  Y��_^á`Vj��^u�   �;�}�ƣ`jP�9  Y�@ ��Yu!jV�5`�   Y�@ ��Yuj����Y3ɸ�� �@ ��� ��=x� |�3ɺ� ��������4� � �������t��u�
��� A��h� |�^��B*  �=��  t�))  ËD$��� ;�r=X� w+�����P��  YÃ� P�D� ËD$��}��P��  YËD$�� P�D� ËD$��� ;�r=X� w+�����P��  YÃ� P�H� ËD$��}��P��  YËD$�� P�H� �SV�t$W�t$�����w��uj^�����3����w:;X� wj	�/  S�3  j	���  ����u+Vj�5< �(� ����u"�=��  tV�  ��Yt�Sj W�I�������_^[�3���V�t$WV������NYx
��8@��	V�)  Y��V�����Y��_^������������SV�D$�u�L$�D$3���؋D$����A�ȋ\$�T$�D$���������u�����d$�ȋD$���r;T$wr;D$vN3ҋ�^[� U��SV�u�F�^����   �@��   �t�f ���   �N$���F�F�f �e $�f��Fu"��� t��8� uS�,  ��YuV�>,  Yf�FWtg�F�>+��H��NI���N~WPS�%*  ���E�6���t�ˋ������� � ������`� �@ tjj S�)  ���F�M��j�E_WPS��)  ���E9}_t�N ��E%�   � �F���^[]�U���H  SVW�}3��G�ۉu�u�}��  �M�3���M��u�3�9U���  �� |��x�Ê��� ���3������ �����E���  �$��� �M���ỦU؉U��U�U��U��x  �Ã� t;��t-��tHHt���Y  �M��P  �M��G  �M��>  �M���5  �M��,  ��*u#�EP��  ��Y�E��  �M��؉E��  �E��ˍ��DA���U���  ��*u�EP�  ��Y�E���  �M����  ���ˍDAЉE��  ��It.��ht ��lt��w��  �M��  �M��  �M� �  �?6u�4uGG�M���}�l  �UЋ0� �U����DA�t�E�P�u��P�  ���G�}�E�P�u��P�f  ���%  �Ã�g�  ��e��   ��X��   �x  ��C��   HHtpHHtl����  f�E�0u�M��u����u�����EP�  f�E�Y�ȉM���  ��u	��� �M��E�   ����N����  f�8 ��  @@���E�   �� �M�@������;ʉ}���   �E�   ��   f�E�0u�M�f�E��EPt;�0  P������P�+)  ���E��}2�E�   �)��Zt2��	t�H��  �  ��  Y�������E�   �������E���  �EP�  ��Yt3�H��t,�E�t� ��M��E��E�   �  �e� �M�� �  ��� �E�P�   u��gu�E�   �E�ũ��E�u��H��M��@��E���P������P�E�P�� �u�����   t�}� u������P�$� Y��gu��u������P�� Y������-u�M��������}�W����Y��  ��i��   ����   H��   HtQ�������HH��   ����  �E�'   �<+����  ��u	��� �M�����N��t�8 t@��+��  �E�   �E�   �E���E�   t]�E��E�0Q�E�   �E��H�E���E�   t;�M��5�EP�  �E� Yt	f�M�f���M��E�   �#  �M�@�E�
   �E��t�EP��  Y�A�E� t!�E�@�EPt��  Y����%�  Y�����E�@�EPt�  Y���  Y3��E�@t��|��s�؃� ���ڀM���������E��u�� �}� }	�E�   ��e�����u�e� �E��E��E��M������t;�E��RPWV�E��U��'  �uċ؃�0�u�WV������9����~]ԋE��M��뵍E�+E��E��E��E�t�M��90u��u�M�@�M��0�E�}� ��   �]���@t&��t�E�-���t�E�+�	��t�E� �E�   �u�+u�+u���u�E�P�uVj �  ���E�P�E��u�u�P�2  ����t��u�E�P�uVj0��   ���}� tA�}� ~;�E�]��x�f�CP�E�PC�L%  Y��Y~2�M�Q�uP�E�P��   ����O��u���E�P�u�u��u��   ���E�t�E�P�uVj �q   ���}�G�ۉ}�����E�_^[��/� �  � l� �� �� �� s� U��M�Ix��E�����Q�u����YY����Eu��]�� ]�VW�|$��O��~!�t$V�t$�t$�������>�t��O���_^�S�\$��KVW��~&�|$�t$�WF�t$P�u������?�t��K���_^[ËD$� � �@�ËD$� ��A��Q�ËD$� � f�@��U����  �e� SV�u3�W��]����]���	  �}��}3ۃ=@� ~��jP�F&  YY��0� ���A��;�t6�M�W�E�WP�%
  YYP�
  �FFP��%  ����t�FFP��%  Y��>%��  �e� �e� �e� �e� �e� �e� 3��e� �]�]��]��E��]��^F�=@� ~��jP�%  YY��0� �ÊA����t�E��E����DCЉE��e��N>t^��*t2��FtT��It
��Lu7�E��E�~6u,�~4�Fu#�EЃe� �e� ���'�E��"��ht��lt
��wt�E���E��E���M��M��}� �O����}� �uu�E�E����E�@��EԀe� �}� u�<St
<Ct�M����E��]�3�� ��n�u�t(��ct��{t�u�E�P�  Y��u�E��v  Y�E�3�9E�t	9E���  ��o�^  �
  ��c�,  ��d��  �j  ��g~8��it��n�W  �}� �}��   �!  jd^�]��-�~  �E��z  �]썵<�����-u��<�����=������+u�}�M��E�W��  ��Y�]���}�}� t	�}�]  ~�E�]  �=@� ~jS��#  YY��0� �X����t!�E��M��t�E�F�E�W�p  ��Y�]��8D� uf�E��M��t\�E�W�M  �ؠD� �Y�]�F�=@� ~jS�[#  YY��0� �X����t!�E��M��t�E�F�E�W�  ��Y�]�뻃}� ��   ��et	��E��   �E��M��tv�eF�E�W��  ��Y��-�]�u�F���+u�E��M��u!E���E�W�  ��Y�]�=@� ~jS�"  YY��0� �X����t�E��M��t�E�F��M�WS�r  �}� YY��  �}� �M  �È& ��<���P�E��u�HP� � ���)  9E�u
�E��E�   �}� ~�E���� �  �ƃ�p��  ����   HH��  ���������t$�;E��?  �M�}� ��  �E��E�  �}� ~�E��}G�}�?^��   �Ǎx�   ��+u"�M�u�}� t�E���u�E��h  ��Y�]��0�E  �u�E��N  ��Y��x�]�t/��Xt*��x�E�   tjo^�  �u�M�S�8  YYj0[��  �u�E��	  Y�؉]�jx�π}� ~�E���� �M��j �E�j P��������}�{u�?]u	�]G�E� ��Uˊ<]t_G<-uA��t=���]t6G:�s�����:�w!����+�F�ʋ������D�BNu�2���ȊЋ��������D�뛀? �  �}�{u�}�}�u��M�W�u�u��S  YY�}� t�E��M����   �E�W�  ���Y�E�t~��j��Z�]�������L�3˅�t`�}� uR�}� tA�0� �E����DA�t�E�W��  Y�E��5@� �E�P�E�P�  f�E�f�FF��F�u��d����E��\����M�WP�  YY9u��(  �}� �  �Ẽ}�c�r  �}� �E�t	f�  �`  �  �X  �E��]��-u�E����+u"�M�u�}� t�E���u�E��  Y�؉]�}� �  �}� ��   ��xuO�=@� ~h�   S�  YY��0� �X%�   ����   �E؋U�jY�J���S�E؉U��}  ��Y�]��S�=@� ~jS��  YY��0� �X����t]��ou��8}S�E؋U�jY������j j
�u��u��	����E؉U��E�CЙE�U܃}� t�M�t$�u�E��6  ��Y�]��+����u�M�S�9  YY�}� ��   �E؋M��؃� �E��ىM���   �}� ��   ��xt?��pt:�=@� ~jS�  YY��0� �X����tv��ou
��8}l���?�<����8�=@� ~h�   S��  YY��0� �X%�   ��t7S���D  ��Y�]��E�}� �|�t�M�t$�u�E��X  ��Y�]��\����u�M�S�[  YY�}� t�߃�Fu�e� �}� ��   �}� u)�Ẽ}� t�EԋM؉�M܉H��}� �E�t�8�f�8�E��E�u�B�E�W��   ��Y�F;É]�uuU�0� ���DA�t�E�W�   Y�F;ȉuu>�M��}��u�>%uM�E�xnuD������V����0�u�M��u���M�WS�   YY��M�WP�}   �M�WS�s   ���}��u�E̅�u8E�u�����E�_^[�Ã=@� V~�t$jV�N  YY��t$�0� �p����u��߃���^ËT$�Jx	�
�A�
�R�u  YÃ|$�t�t$�t$�t  YY�V�t$W�t$�������W�  Y��Yu��_^á�� ��t�t$�Ѕ�YtjX�3��3�j 9D$h   ��P�P� ���< t�  ��u�5< �L� 3��jX�S3�94 U�-,� ~D�8 VW�=T� �ph @  h   �6��h �  j �6���vj �5< �Ճ�C;4 |�_^�58 j �5< ���5< �L� ][�V�5X� �5�� ���5�� ���5�� ���5�� ��^�VW�=\� ��� ���t+���� t#���� t���� t���� tP���6�����Y����X� |��5�� ���5�� ���5�� ���5�� ��_^�U��EV�<���  �4��� u>Wj�������Y��uj�p���Yj������> YWu
�X� �>��S���Yj�   Y_�6�D� ^]�U��E�4��� �H� ]�h@  j �5< �(� ���8 uÃ%0  �%4  j�, �$    Xá4 ���8 ��;�s�T$+P��   r����3��U����U�MSV�A��+q�Z����W���΋z�i�  K�}���D  �]�M�����M�u��j?I_�M;�v�}�L;LuH�M�� s�   ���L��!|�D�	u+�M!9�$���   ���M�L��!���   �	u�M!y�L�|�y�L�|]��y�]����O��?vj?_�M����M���   +U��M���j?�U�IZ;ʉMv�U��]����]���O;�v��;�tk�M��Q;QuH�M�� s�   ���L��!T�D�	u+�M!�$���   ���M�L��!���   �	u�M!Q�M��Q�I�J�M��Q�I�J�U��}� u	9}��   �M����I�J�M����J�Q�J�Q�J;Juc�L�� �M���Ls%�} u�   �����M	�   �����D�D	�)�} u�O�   ���M	Y�O�   ����   	8�]�E���\����   �0 ����   �( �=T� ��H� �  h @  SQ�׋( �0 �   ���	P�0 �( �@����    �0 �@�HC�0 �H�yC u	�`��0 �x�ulSj �p�ס0 �pj �5< �,� �4 �8 �����ȡ0 +ȍL�Q�HQP�  �E���4 ;0 v���8 �, ��E�0 �5( _^[��U����4 �8 SV��W�<��E�}��H����M���I�� }�����M���u��������3���u�E��, ��;߉]s�K�;#M�#��u��;]��]r�;]�uy��;؉]s�K�;#M�#��u����;�uY;]�s�{ u���]��;]�u&��;؉]s�{ u����;�u�8  �؅ۉ]tS��  Y�K��C�8�u3��  �, �C�����U�t����   �|�D#M�#��u7���   �pD#U�#u�e� �HD֋u�u���   �E�#U�����#9�t�U���3�i�  ��D  �M�L�D#�u����   j #M�_��|��G���M�T��
+M���M���N��?~j?^;��  �J;Jua�� }+�   �����M��|8�Ӊ]�#\�D�\�D�u8�]�M�!�1�O�   ���M��|8����   ��!��]�u�]�M�!K��]�J�z�}� �y�J�z�y��   �M�|���z�J�Q�J�Q�J;Jud�L�� �M})���} �Lu�   �����	;�   �����M�	|�D�/���} �Lu�N�   ���	{�M�����   �N�   ���	7�M���t�
�L���M��u�эN�
�L2��u��ɍy�>u;0 u�M�;( u�%0  �M���B_^[�á4 �$ VW3�;�u0�D�P��P�58 W�5< �d� ;�ta�$ �8 �4 �8 h�A  j���5< �4��(� ;ǉFt*jh    h   W�`� ;ǉFu�vW�5< �,� 3���N��>�~�4 �F����_^�U��Q�MSVW�q�A3ۅ�|��C����j?i�  Z��0D  �E��@�@��Ju��j��yh   h �  W�`� ��u����   �� p  ;�w<�G�H�����  ����  �@��  ��������Hǀ�  �     �H�;�vǋE��O�  j_�H�A�J�H�A�d�D ����   �FC�������E�NCu	x�   �������!P��_^[��V�����p� ����\� t:jtj������Y��Yt)V�5\� �l� ��tV�4   Y�h� �N�j�X^�3�^��|����\� ���tP�t� �\� �ËD$�@PP� �@   �VW��� �5\� ���|� ����u?jtj�2�����Y��Yt&V�5\� �l� ��tV����Y�h� �N���j� ���YW�x� ��_^á\� �����   V�t$��uP�|� ����tl�F$��tP�����Y�F(��tP����Y�F0��tP����Y�F8��tP����Y�F@��tP����Y�FD��tP�}���Y�FP=P� tP�l���YV�e���Yj �5\� �l� ^�U���HSVWh�  ������Y��uj�2���Y�5 � �      ���  ;�s�f ���f �F
� � ��$�  �ލE�P��� f�}� ��   �E����   �8�X�;�E��   ;�|��9=  }V�$� h�  �!�����Yt<�   ����  ;�s�` ���` �@
���$���  ����9=  |���=  3���~L�E�����t8��t2�uQ��� ��t#�΋������� � �����M��	���H�E�FC;�|�3ۋ � �ۃ<���4�uM���F�uj�X�
��H������P��� �����tW��� ��t%�   �>��u�N@���u
�N��N�C��|��5  ��� _^[��SVW� � ���t7���  ;�s!�_�{� tS�\� ���$�  ��$;�r��6�W����& Y����  |�_^[�S3�9hVWu�  �5�� 3��:�t<=tGV�n���Y�t���   P�y�����Y;�5�� uj	�����Y�=�� 8t9UW�4�����YE�?=t"U�D���;�Y�uj	�����YW�6�����Y��Y�8u�]�5�� ����Y��� �_^�d   [�U��QQS3�9hVWu�F  �P� h  VS��� �x�5�� ��8t���E�P�E�PSSW�M   �E��M���P��������;�uj����Y�E�P�E�P�E���PVW�   �E���H�5�� _^��� [��U��M�ESV�! �uW�}�    �E��t�7���}�8"uD�P@��"t)��t%����� t���t��F@���tՊ�F�����t�& F�8"uF@�C���t��F�@����� t���t��F@�� t	��t	��	ū�uH���t�f� �e �8 ��   ��� t��	u@��8 ��   ��t�7���}�U��E   3ۀ8\u@C���8"u,��u%3�9}t�x"�Pu����}�}3�9U�U���K��tC��t�\F�Ku���tJ�} u
�� t?��	t:�} t.��t����� t�F@���F������ t@��@�X�����t�& F�������t�' �E_^[� ]�QQ�T� SU�-�� VW3�3�3�;�u3�Ջ�;�t�T�    �(��� ��;���   �T�    �   ����   ;�u�Ջ�;���   f9��t@@f9u�@@f9u�+Ƌ=�� ��SS@SSPVSS�D$4�׋�;�t2U����;�Y�D$t#SSUP�t$$VSS�ׅ�u�t$�z���Y�\$�\$V��� ���S��uL;�u��� ��;�t<8��t
@8u�@8u�+�@��U������Y;�u3��UWV������W��� ���3�_^][YYá�� ��t��u*�=�� u!h�   �   �X� Y��t��h�   �   Y�U���  �U3ɸ�� ;t��A=� |�V����;��� �  ��� ����   ��u�=�� ��   ���   ��   ��\���h  Pj ��� ��u��\���h<� P�p���YY��\���WP��\�������@Y��<v)��\���P�x�������\�����;j�h8� W�  ����`���h� P������`���WP������`���h� P�������� ��`���P�����h  ��`���h�� P�  ��,_�&�E���� j P�6�����YP�6j���� P�$� ^��SWj3������Yj_9=`~]V�@ �������tA�@�tP��  ���YtC��|)�@ ��� P�\� �@ �4� ����@ Y�$ G;=`|�^j�����Y��_[�V�t$V�#   ��Yt���^��F@t�v��  ��Y^��3�^�SV�t$3�W�F�ȃ���u7f�t1�F�>+���~&WP�v�  ��;�u�F��t$��F��N ����F�f �_��^[�j�   Y�SVWj3�3�����3�Y95`~t�@ ����t_�@�tYPV������@ YY���H���t0�|$uP�������YtC��|$ u��tP�������Yu��@ �4�V�����YYF;5`|�j�����|$Y��t��_^[�V�t$�F����   �@��   �t
 �F�   f��Fu	V�m  Y��F��v�v�v�  ���F��to���tj�V�u7�NW���t�������<� � �ɍ<���`� �O_�ႀ��u�� �V�~   u�N��t��u�F   �H�F�A�^��������	F�f ���^�V�t$;5  s@�΋������� � ���D�t%WV��  �t$�t$V�(   V���  ����_^���  � 	   ��  �  ���^�V�t$WV�P  ���Yu�  � 	   �-�t$j �t$P��� �����u��� �3���tP�  Y�����΃����Ƌ� � ���d���D���_^�V�t$;5  s@�΋������� � ���D�t%WV��  �t$�t$V�(   V���E  ����_^��  � 	   �  �  ���^�U���  SVW3�9}�}��}�u3��f  �E���� � �E���4�����D0 tjW�u����������@���   �E9}�E��}��   �������M�+M;Ms)�M��E��	��
u�E�� @�@�ȍ�����+ʁ�   |̋�������+��E�j P������WP��40�$� ��tC�E�E�;�|�E�+E;Er�3��E�;���   9}tbj^9uuL��  � 	   ��  �0�A��� �E�ǍM�WQ�u�u�0�$� ��t�E�}�E����� �E��u�,  Y����,��D0@t�E�8������  �    �}  �8��+E�_^[����� h   ����Y�L$���At�I�A   ��I�A�A�A   �A�a �ËD$;  r3�Ëȃ������� � �D���@�U��SV��� WV��� �=�� 3�9�� tV��j�����Yj[�u�u�   Y�E��Yt
j�.���Y�V�׋E_^[]�U��E��u]Ã=��  uf�Mf��� w9j�X]ÍM�e Qj �5@� P�EjPh   �5�� ��� ��t�} t�D  � *   ���]�����������S�D$�u�L$�D$3���D$���3��P�ȋ\$�T$�D$���������u�����d$��d$�r;T$wr;D$v+D$T$+D$T$���؃� [� U��SV��� WV��� �=�� 3�9�� tV��j����Yj[�u�u�u�   ���E��t
j�����Y�V�׋E_^[]�U��SV�u3�;�t9]t�:�u�E;�tf�3�^[]�9�� u�M;�tf��f�jX��0� ���DA�tN�@� ��~*9E|/3�9]��Q�uPVj	�5�� ��� ���@� u�9Er8^u���  � *   ����3�9]��P�ujVj	�5�� ��� ���x����Ƀ=@� ~j�t$�   YYËD$�0� �A���U��Q�E�H��   w�0� �A�R��V�50� �����DV�^t�e� �M��E�j�	�e� �E�jX�M
jj j QP�E�Pj�f  ����u���E
#E��S�\$���VtA�t$�F�u��t2�u.�~ uV�e���Y�;Fu	�~ u@��F@t��8t@����^[�����F�F$��F��%�   ������������U��WV�u�M�}�����;�v;��x  ��   u������r)��$�X� �Ǻ   ��r����$�p� �$�h� ��$�� ��� �� Я #ъ��F�G�F���G������r���$�X� �I #ъ��F���G������r���$�X� �#ъ�F��G��r���$�X� �I O� <� 4� ,� $� � � � �D��D��D��D��D��D��D���D���D��D��D���D���D���D����    ���$�X� ��h� p� |� �� �E^_�Ð���E^_�Ð���F�G�E^_�ÍI ���F�G�F�G�E^_�Ð�t1��|9���   u$������r����$�� �����$��� �I �Ǻ   ��r��+��$��� �$�� �� (� P� �F#шGN��O��r�����$�� �I �F#шG�F���G������r�����$�� ��F#шG�F�G�F���G�������Z�������$�� �I �� �� �� �� ı ̱ Ա � �D��D��D��D��D��D��D��D��D��D��D��D��D��D���    ���$�� �� � � � ,� �E^_�Ð�F�G�E^_�ÍI �F�G�F�G�E^_�Ð�F�G�F�G�F�G�E^_��U���SVWj�W����u�  ��Y;�� Y�]u3��p  ���V  3Ҹ�� 9tt��0B=�� |�E�PS��� j^;��!  j@�%�  Y3�� � 9u�󫪉�� ��   �}� ��   �M�����   �A���;���   ��� @��e� j@Y3�� � �4R�������� �; ��t,�Q��t%���;�w�U����� �� @;�v�AA�9 u��E����}�r��E���    P��� ��   ���� ��� ��Y�� ��RAA�y� �G����ƀ�� @=�   r�S�   Y�� �5�� ��%��  3���� �����=\�  t�   �   �������j�#���Y��_^[�ËD$�%\�  ���u�\�    �%�� ���u�\�    �%�� ���u��� �\�    ËD$-�  t"��t��tHt3�ø  ø  ø  ø  �Wj@Y3�� � �3���� ��� ��� �� ���_�U���  �E�VP�5�� ��� ���  3��   ������@;�r�E�ƅ���� ��t7SW�U��
��;�w+ȍ�����A�    �����˃��BB�B���u�_[j �������5� �5�� P������VPj�  j �������5�� VP������VPV�5� ��  j �������5�� VP������VPh   �5� �  ��\3�������f���t��� �������� � ���t���  �������〠 �  @AA;�r��I3��   ��Ar��Zw��� �Ȁ� �� � ���ar��zw���  �Ȁ� ���� �  @;�r�^�Ã=h uj�����Y�h   �S3�9`� VWuBh�� ��� ��;�tg�5�� hx� W�օ��`� tPhh� W��hT� W�d� �֣h� �d� ��t�Ћ؅�t�h� ��tS�Ћ��t$�t$�t$S�`� _^[�3����������������̋L$W��tzVS�ًt$��   �|$u��uo�!�F�GIt%��t)��   u����uQ��t�F�G��t/Ku�D$[^_���   t�GI��   ��   u����ul�GKu�[^�D$_É��It�����~�Ѓ��3��� �tބ�t,��t��  � t��   �uƉ�����  �����   ��3҉��3�It
3����Iu���u��D$[^_�V�t$W����F@t�f �V����V�   V�����������_^�V�t$W����F�t4V�f���V���H	  �v�`  ����}�����F��tP�����f Y�f ��_^�S�\$;  VWsr�����<� � �Ã��4�����D0tRS��  �Y�D0t)S�  YP��� ��u
��� ���3���t��  �0��  � 	   ���S��  Y����  � 	   ���_^[�V�t$;5  s@�΋������� � ���D�t%WV�U  �t$�t$V�(   V���  ����_^��_  � 	   �]  �  ���^�U����e� �} S�]VW����  �E�ȃ����4��� � �<� � ��ƊH����  ��Ht�@<
t�M���S�E�   �D0
�E�j P��uR�40�� ��u9��� j^;�u�  � 	   �  �0���m�$  P�%  Y����  ��U�U��L0�D0����   ��t	�;
u�$���E�M��E�;��M���   �E� <��   <t�C�E�   I9Ms�E@�8
u�E�^�C�E�s�E�j P�E�E�jP��40�� ��u
��� ��uG�}� tA��D0Ht�E�<
t��C�D1�);]u�}�
u�
�jj��u��������}�
t�C�M�9M�G������t0��@u�+]�]��E��3�_^[��V�v   �L$3����� ;t"��F=8� |��r"��$w�B   �    ^��5   ���� ^�Á��   r���   w�   �    ^��   �    ^��\�������S�����ËL$V;  WsX�����<� � �����4������@t7�8�t2�=�� u3�+�tItIuPj��Pj��Pj���� ��0�3������� 	   �����  ���_^ËD$;  s�ȃ������� � �D���t� ��?���� 	   �=����  ���ËD$S�ȃ���VW�4� � �� � �<�����~ u#j�����~ Yu�FP�X� �Fj�^���Y��D8P�D� _^[ËD$�ȃ������� � �D�P�H� �j�`���Y�U��j�h�� h�� d�    Pd�%    ��SVW�e衘� 3�;�u>�E�Pj^Vh�� V��� ��t����E�PVh�� VS��� ����   jX��� ��u$�E;�u��� �u�u�u�uP��� �   ����   9]u��� �ESS�u�u�E �����@P�u��� �E�;�tc�]��< �ǃ�$���  �e��u�WSV�0������jXËe�3�3��M��;�t)�u�V�u�uj�u��� ;�t�uPV�u��� �3��e̋M�d�    _^[��U��j�h�� h�� d�    Pd�%    ��SVW�e�3�9=�� uFWWj[Sh�� �   VW��� ��t��� �"WWSh�� VW��� ���"  ���    9}~�u�u�  YY�E��� ��u�u�u�u�u�u�u��� ��   ����   9} u��� �E WW�u�u�E$�����@P�u ��� �؉]�;���   �}����$��y  �e�ĉE܃M���jXËe�3��}܃M���]�9}�tfS�u��u�uj�u ��� ��tMWWS�u��u�u��� ���u�;�t2�Et@9}��   ;u�u�uS�u��u�u��� ����   3��eȋM�d�    _^[���E�   �6��$���  �e�܉]��M���jXËe�3�3ۃM���u�;�t�VS�u��u��u�u��� ��t�9}WWuWW��u�uVSh   �u ��� ��;��q������l����T$�D$��V�J�t�8 t@��I��u�8 ^u+D$Ë��V�t$;5  s8�΋������� � ���D�tWV����V�(   V��� �������_^������� 	   �����  ���^�V�t$WV�3������Yt<��t��uj����j������Y;�YtV����YP�� ��u
��� ���3�V�j����ƃ���Y�� � ���d� ��tW�����Y����3�_^�V�t$�F��t�t�v�϶��f�f��3�Y��F�F^�̋T$�L$��   u<�:u.
�t&:au%
�t��:Au
�t:au����
�uҋ�3�Ð���@Ë���   t�B:u�A
�t���   t�f���:u�
�t�:au�
�t����������������U��V3�PPPPPPPP�U�I �
�tB�$��u����A�
�tF�$s���� ^����U��WVS�M�&�ً}��3����ˋ��u�F�3�:G�wtII�ы�[^_����������U��V3�PPPPPPPP�U�I �
�tB�$��u�
�t
F�$s�F��� ^����U��SVWUj j h�� �u�X  ]_^[��]ËL$�A   �   t�D$�T$��   �SVW�D$Pj�h�� d�5    d�%    �D$ �X�p���t.;t$$t(�4v���L$�H�|� uh  �D��@   �T���d�    ��_^[�3�d�    �y�� u�Q�R9Qu�   �SQ�P� �
SQ�P� �M�K�C�kY[� ��VC20XC00U���SVWU��]�E�@   ��   �E��E�E��E��C��s�{���ta�v�|� tEVU�k�T�]^�]�t3x<�{S�������kVS��������vj�D��a������C�T��{�v�4�롸    ��   �U�kj�S������]�   ]_^[��]�U�L$�)�AP�AP�y�����]� ����Q=   �L$r��   -   �=   s�+ȋą���@P��U��WVS�u�}�x� �x u;����
�t.�F�'G8�t�,A<ɀ� �A��,A<ɀ� �A8�t������x���� �=��  j ����� j�W����$   ��   3ې
�t'�F�G8�t�PS�8  �؃��.  ��8�t�������X�u	���� �
j�g�������[^_��U��WVS�M���   �u�}�x� �x uN�A�Z� �I �&
�t!
�tFG8�r8�w�8�r8�w�8�uIu�3�8���   �������   ���   ���� �=��  j ����� ��j�g����$   ��3�3ۋ����t#�tFGQPS�G   �؃��=   ��Y;�u	Iu�3�;�t	�����r��X�u	���� ���j�h������ˋ�[^_��U��Q�=��  SVWu�E��A��   ��Z��   �� �   �]�   j;�^}%95@� ~VS�'���YY�
�0� �X#ƅ�u���e�0� �������DJ�t�e
 j�E�]	X�	�e	 �]��Vj �M�jQP�EPW�5�� ������� ��t�;�u�E���E��M����_^[�����̍B�[Í�$    �d$ 3��D$S�����T$��   t�
B8�tф�tQ��   u��W����V؋
����~����3���������3�3ƃ��� �u% �t�% u��   �u�^_[3�ËB�8�t6��t�8�t'��t���8�t��t�8�t��t��^_�B�[ÍB�^_[ÍB�^_[ÍB�^_[��%��                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                               <�  H�  V�  b�  p�  ~�  ��  ��  ��  ��  ��  ��  ��  �  �  "�  6�  J�  b�  z�  ��  ��  ��  ��  ��  ��  ��  �  �  &�  0�  @�  N�  ^�  p�  ��  ��  ��  ��  ��  ��   �  �  2�  D�  \�  t�  ��  ��  ��  ��  ��  ��  ��  ��  �  �  &�  6�      "�(ט/�B�e�#�D7q/;M������ۉ��۵�8�H�[�V9����Y�O���?��m��^�B���ؾopE[����N��1$����}Uo�{�t]�r��;��ހ5�%�ܛ�&i�t���J��i���%O8�G��Ռ�Ɲ�e��w̡$u+Yo,�-��n��tJ��A�ܩ�\�S�ڈ�v��f�RQ>�2�-m�1�?!���'����Y��=���%�
�G���o��Qc�pn
g))�/�F�
�'&�&\8!.�*�Z�m,M߳��8S�c��Ts
e��w<�
jv��G.�;5��,r�d�L�迢0B�Kf�����p�K�0�T�Ql�R�����eU$��* qW�5��ѻ2p�j��Ҹ��S�AQl7���LwH'�H�ᵼ�4cZ�ų9ˊA�J��Ns�cwOʜ[�����o.h���]t`/Coc�xr��xȄ�9dǌ(c#����齂��lP�yƲ����+Sr��xqƜa&��>'���!Ǹ������}��x�n�O}��or�g���Ȣ�}c
����?G5q�}#�w�(�$�@{��2���
��<L��gC�B>˾��L*~e��)Y���:�o�_XGJ�Dl�                                                                                                                                      EEE50 P     (8PX 700WP        `h````  ppxxxx          ( n u l l )     (null)  runtime error   
  TLOSS error
   SING error
    DOMAIN error
  R6028
- unable to initialize heap
    R6027
- not enough space for lowio initialization
    R6026
- not enough space for stdio initialization
    R6025
- pure virtual function call
   R6024
- not enough space for _onexit/atexit table
    R6019
- unable to open console device
    R6018
- unexpected heap error
    R6017
- unexpected multithread lock error
    R6016
- not enough space for thread data
 
abnormal program termination
    R6009
- not enough space for environment
 R6008
- not enough space for arguments
   R6002
- floating point not loaded
    Microsoft Visual C++ Runtime Library    

  Runtime Error!

Program:    ... <program name unknown>  GetLastActivePopup  GetActiveWindow MessageBoxA user32.dll          ����� �     ����E� I� ������ �� H:mm:ss dddd, MMMM dd, yyyy M/d/yy  PM  AM  December    November    October September   August  July    June    April   March   February    January Dec Nov Oct Sep Aug Jul Jun May Apr Mar Feb Jan Saturday    Friday  Thursday    Wednesday   Tuesday Monday  Sunday  Sat Fri Thu Wed Tue Mon Sun SunMonTueWedThuFriSat   JanFebMarAprMayJunJulAugSepOctNovDec    L�          ��   �                      <�  H�  V�  b�  p�  ~�  ��  ��  ��  ��  ��  ��  ��  �  �  "�  6�  J�  b�  z�  ��  ��  ��  ��  ��  ��  ��  �  �  &�  0�  @�  N�  ^�  p�  ��  ��  ��  ��  ��  ��   �  �  2�  D�  \�  t�  ��  ��  ��  ��  ��  ��  ��  ��  �  �  &�  6�      �lstrlenA  . CloseHandle �ReadFile  [GetFileSize M CreateFileA eUnmapViewOfFile ^MapViewOfFile N CreateFileMappingA  = CopyFileA �WriteFile KERNEL32.dll  HeapAlloc HeapFree  GetCommandLineA �GetVersion  � ExitProcess QTerminateProcess  :GetCurrentProcess � EnterCriticalSection  GLeaveCriticalSection  
HeapDestroy HeapCreate  xVirtualFree InitializeCriticalSection z DeleteCriticalSection uVirtualAlloc  HeapReAlloc >GetCurrentThreadId  YTlsSetValue VTlsAlloc  WTlsFree SetLastError  XTlsGetValue iGetLastError  SetHandleCount  �GetStdHandle  ^GetFileType �GetStartupInfoA uGetModuleFileNameA  � FreeEnvironmentStringsA � FreeEnvironmentStringsW �WideCharToMultiByte MGetEnvironmentStrings OGetEnvironmentStringsW  SetFilePointer  InterlockedDecrement  "InterlockedIncrement  kMultiByteToWideChar � GetCPInfo � GetACP  �GetOEMCP  �GetProcAddress  HLoadLibraryA  � FlushFileBuffers  ,SetStdHandle  �GetStringTypeA  �GetStringTypeW  :LCMapStringA  ;LCMapStringW  �RtlUnwind                   �?HE    ��           x�  ��  ��  �  �  ��  ��     CdnSign.dll Csn_SplitSgnFile Csn_VerifySgnFile                                                                                                                                                                                                                                                                                                                                                  �{ �         �|                 D� <�     10001   CA5F136A67C6B50ABB0BE8FAC9A2B4B3C4F15731A5E63E42CAD3193C7FAE0E167133D2B9E174E5A90D7DA2DC4FA5B2F68921AC5725261C2F45D9C25A63204FBC3631798984A3403D6B64A54A6617AD753EE573AFEEB108A72F340546F32BF41469FE9DD10C87DC5DD0F65FAD95182A01EAA8B563588ED78176362ED014CB18E9    %02X    0   ���u��ڌ��(�?�wy���r������P(�I ��3��ĵC:��)��&T^��[�K�	�� �� �� �� |� p� h� `� X� P� H� @� 8� 0� (�  � � � �  � �� �� �� �� �� �� �� �� �� �� �� �� �� �� �� x� p� h� `� X� P� H� @� 8� �� 0� (�  � � � �  � �� �� �� �� �� �� �� �� �� �� �� �� �� �� �� �� |� t� l� d� X� L� H� @� 8� 0� (�  � � �  � �� �� �� �� �� �� �� �� �� �� �� t� h� \� P� D� 4� (�  � �  � �� �� �� �� �� �� �� �� �� �� p� d� X� L� 8� �� (� � � �� �� �� �� �� �� �� �� �� p� `� P� @� 0� $� � � �� �� �� set_io_buffer_size  big_to_bytes    bytes_to_big    strong_bigrand  prepare_basis   mul2_brick  ebrick2_init    ecurve2_mult2   ecurve2_multn   ecurve2_mult    ecurve2_multi_add   ecurve2_sub epoint2_negate  ecurve2_add epoint2_comp    epoint2_get epoint2_norm    epoint2_set epoint2_init    ecurve2_init    ecurve_multi_add    epoint_negate   nres_dotprod    nres_multi_inverse  epoint_norm mul_brick   ebrick_init ecurve_multn    powmodn nres_powmodn    set_user_function   pow_brick   brick_init  lucas   nres_lucas  nxsafeprime trial_division  ecurve_sub  ecurve_mult2    nres_premult    sqroot  nres_sqroot nres_powmod2    epoint_get  epoint_set  epoint_init ecurve_mult ecurve_add  ecurve_init nres_negate nres_modsub nres_modadd fmodulo remain  divisible   nres_powltr nres_moddiv nres_powmod nres_modmult    redc    nres    prepare_monty   powmod2 cinstr  cotstr  instr   otstr   crt crt_init    fft_mult    powltr  gprime  flop    facosh  fcosh   fasinh  fsinh   fatanh  ftanh   facos   fcos    fasin   fsin    fatan   ftan    fpowf   flog    fexp    fpi froot   fpower  expint  logb2   build   sftbit  frand   ftrunc  fincr   fpmul   frecip  fconv   fcomp   fsub    fadd    fdiv    fmul    mround  mr_shift    dconv   fpack   xgcd    mirsys  subtract    add putdig  multi_inverse   mad mirvar  isprime nxprime bigrand bigdig  powmod  power   nroot   cotnum  cinnum  cbase   egcd    fdsize  subdiv  premult decr    incr    divide  multiply    normalise   jack    otnum   innum   your program    Unable to control Floating-point rounding
  Specified basis is NOT irreducible
 Specified double length type isn't double length
   Number Base must be power of 2
 Exponent too big
   No modulus defined
 Illegal modulus 
   MIRACL not initialised - no call to mirsys()
   I/O buffer overflow
    Flash to double conversion failure
 Log of a non-positive number
   Numbers too big
    Flash overflow
 Integer operation attempted on Flash number
    Attempt to take illegal root
   Raising integer to negative power
  Even root of a negative number
 Out of space
   Illegal parameter usage
    Illegal number base
    Input format error
 Internal result is negative
    Overflow - Number too big
  Division by zero attempted
 Number base too big for representation
               called from   ??? 
MIRACL error from routine          �z     `     `                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                      \� L�  	-]   ]          ��                              �             8�             �                                                                                                                         �  �������� 
                                     ��    �� 	   p� 
   L�     �    ��    ��    ��    h�    @�    �    ��    �� x   �� y   �� z   x� �   t� �   d� � � � � � � :� :�                     ( ( ( ( (                                     H                � � � � � � � � � �        � � � � � �                           � � � � � �                                                                                                                                                                                                                                                                                                    .            �         �       �  �       �  �       �  �       �  �       �  �       �  �       �  �       �  �             x   
       �  `�y�!       ��      ��      ����    @~��    �  ��ڣ                        ��      @�      �  ��ڣ                        ��      A�      �  Ϣ� ��[                 ��      @~��    Q  Q�^�  _�j�2                 ������  1~��                                     	               	      
                                                !      5      A      C      P      R      S      W      Y      l      m       p      r   	         �   
   �   
   �   	   �      �      �   )   �      �      �      �      �      �      �           C   C                                                                                                                                   C                                                                                                                                                �            h�     �� �� �� �� �� �� �� �� �� �� �� �� �� �� �� |� x� t� p� l� h� d� `� \� X� T� L� @� 8� 0� p� (�  � � � � �� �� �� �� �� �� ��     .       � � � � � � � � � �  �             �p     ����PST                                                             PDT                                                             l� ��     ����            ����        ����   ;   Z   x   �   �   �   �     0  N  m  ����   :   Y   w   �   �   �   �     /  M  l                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                          �                  0  �                 H   `  d                  d4   V S _ V E R S I O N _ I N F O     ���               ?                       �   S t r i n g F i l e I n f o   �   0 8 0 4 0 4 b 0       C o m m e n t s   ,   C o m p a n y N a m e     C N N I C   Z   F i l e D e s c r i p t i o n     C N N I C   F i l e   V e r i f y   M o d u l e     6   F i l e V e r s i o n     1 ,   0 ,   0 ,   3     0   I n t e r n a l N a m e   C d n S i g n   N   L e g a l C o p y r i g h t   C o p y r i g h t   C N N I C   2 0 0 6     4   L e g a l T r a d e m a r k s     C N N I C   @   O r i g i n a l F i l e n a m e   C d n S i g n . d l l   0   P r i v a t e B u i l d   1 . 1 . 0 . 3   0   P r o d u c t N a m e     C d n S i g n   :   P r o d u c t V e r s i o n   1 ,   0 ,   0 ,   3          S p e c i a l B u i l d   D    V a r F i l e I n f o     $    T r a n s l a t i o n     �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                               �   �0�0�0s1�1�2�2�3�3�344w4�4�4�4�4�4�4?5U5q5�5�5�5�5�5�5�599�<�=�=�=�= >>/>7>D>n>s>}>�>�>�>�>�>�>�>�>�>�>�>�>�>�>�>�>?
????&?-?@?D?H?L?P?T?X?\?`?d?h?l?p?t?x?|?�?�?�?�?�?�?�?�?�?�?�?      �   
00*0I3U3g3t3�3�3�3�3�3�3�3�3 444*4E4V4n4�4�4�4�4�4�455(535?5O5Z5f5r5}5�5�5�5�5�5�5�566+6T6b6n66�6�6�6�6�6�6�6�6�6	77(7:7G7Y7f7x7�7�7�7�7�7�7�7�788#858B8T8a8s8�8�8�8�8�8�8�8�8�89)9I9X9�9�9::6:T:p:�:�:�:�:�: @     O:;;;;   p  �   4 4'4/44484<4e4�4�4�4�4�4�4�4�4�4�4555 5$5�5�5�5�5�5�5�5�56=6D6H6L6P6T6X6\6`6�6�6�6�6�6�78>8D8�8�8�8�8�89999"9:9?9I9c9q9y99�9�90:K:Z:v:~:�:�:�:�:�:�:�:	;;; ;9;A;F;R;W;t;z;�;<<<)<=<C<Q<Z<k<�<�<�<�<�<�<�<==B=p=�=�=�=�>�>,?9?�?�? �  T   011�1�2<3]3t3�3�6�6�6�6�6�6�6�6�7�7h8�8K:_:�:�:�:�:`;t;�;�;=>1>�>?L?`?   �    0%0K0b0(1�1�1L2y2�2�2�2�2�2�2�2�2�2�23
333 3(30383D3I3U3]3e3m3�3�3�3�3�3�3�3�3444+41484A4H4P4V4a4i4�6�6�6�6�6�6 777-7@7K7Q7V7\7i7�7�7�7�7�7�7�7�78�8�:�:�:�:�:�:�:�:�:�:�:;;;7;H;N;a;�;s<{<�<�<�<�<�<�<�<�<�<= =&=7=N=X=q=�=�=�=>!>C>W>�>�>�>�>�>??;?e?s?�?�?�?�?�? �  �   00M0]0�0�0�0�0�0�0�0�0K1R1�1�1�2�23323>3N3�3�3�3.4@4O4a4�4�4�4�4�4�4�485L5j5v5�5�5�5�5�5�5666,686�6�67T7f7�78f8y8�8�8"9>9Q9�9e:�:�:�:);q;�;�;�;�;�;�; <2<8<�<�<�<�<]=x=�=�=�=�=�=�=�=>7>F>H?`?g?o?t?x?|?�?�?�?�?�?�?�?�?   �  <   000R0X0\0`0d0�0�0�0�0�0 11!1K1}1�1�1�1�1�1�1�1�1�1�1�1�1�1b2~2�2�2�2�2�2�23343:3[3e3p3u3}3�3�3�3�3�3�3�3444#4-434v4�4�4�4�4�4�45#5A5R5e5z5�5�5�5�5�5�566606>6G6M6Y6^6h6o6w6}6�6�6�6�6R8b8�8�8�8�8p9w9�9�9�:�:+;8;];�;�;�;�;&<:<t<{<�<�<�<�<�<�<=&=-=?=G=W=h={=�=�=	>>;>@>_>l>y>�>�>�>�>�>�>�>?n?�?�? �  @   0D0�0�01'1C1�2)3�3�3�3�465<5J5�5�5$6*686�6�6�677P7N8 �     �7�7�7�7�7�7 �  D  0000040�1�1�1�1�1�1�1�1�1�1�1�1�1�1�1�1�1�1�1�1�1�1�1�1�1�1�1 22222222 2$2(2,2024282<2@2D2H2L2P2T2X2\2`2d2h2l2p2t2x2|2�2�2�2�2�2�2�2�2�2�2�2�2�2�2�2�2�2�2�2�2�2�2�2�2�2�2�2�2�2�2�2�2 33333333 3$3(3,3034383<3@3D3H3L3P3T3X3\3`3d3h3l3p3t3x3|3�3�3�3�3�3�3�3�3�3�3�3�3�3�3�3�3�3�3�3�3�<�< =�?�?�?�?�?�?   �  �   �0�0�0�0�0�0�0�0�0�0�0�0�0�0�011111 1$1(1,10141`7h7l7p7t7x7|7�7�7�7�7�7�7�7�7�7�7�7�7�7�7�7�7�7�7�7�7�7�7�7�7�7�7�7�7�7�7�7�7 88888 8$8(8,8084888<8@8D8P8�8�8                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                          ���/���3���%�m�KBwA���K��M��}��^n	W�~p �əSj�(.���T�參��
4�l|Q�Тcg��8TQެ� �-�[�L��5��K{v�w��T�`%���)�Xb^�g�wF�wF�wF�wF�wF�wF�wF�wF�wF�wF�wF�wF�wF�wF�wF�wF�wF�wF�wF�wF�wF�wF�wF�wF�wF�wF�wF�wF�wF�wF�wF�wF�wF�wF�wF�wF�wF�wF�wF�wF�wF�wF�wF�wF�wF�wF�wF�wF�wF�wF�wF�wF�wF�wF�wF�wF�wF�wF�wF�wF�wF�wF�wF�wF�wF�wF�wF�wF�wF�wF�wF�wF�wF�wF�wF�wF�wF�wF�wF�wF�wF�wF�wF�wF�wF�wF�wF�wF�wF�wF�wF�wF�wF�wF�wF�wF�wF�wF�wF�wF�wF�wF�wF�wF�wF�wF�wF�wF�wF�wF�wF�wF�wF�wF�wF�wF�wF�wF�wF�wF�wF�wF�wF�wF�wF�wF�wF�wF�wF�wF�wF�wF�wF�wF�wF�wF�wF�wF�wF�wF�wF�wF�wF�wF�wF�wF�wF�wF�wF�wF�wF�wF�wF�wF�wF�wF�wF�wF�wF�wF�wF�wF�wF�wF�wF�wF�wF�wF�wF�wF�wF�wF�wF�wF�wF�wF�wF�wF�wF�wF�wF�wF�wF�wF�wF�wF�wF�wF�wF�wF�wF�wF�wF�wF�wF�wF�wF�wF�wF�wF�wF�wF�wF�wF�wF�wF�wF�wF