MZ�       ��  �       @                                   �   � �	�!�L�!This program cannot be run in DOS mode.
$       �J%ߍ+K��+K��+K��+J��+K�wR��+K�w��+K�WW��+K�wv��+K�Rich�+K�                PE  L ��H        �  �                     �   �             �     �                                �  (                              4   0                                                (                           .text   �                          h.rdata  �                        @  H.data         �                  @  �INIT      �  �  �                 �.reloc  B      �                  @  B                                                                                                                �L$�a 2��  3�� �jhP �r  �  ��u�F`�H�M�H�M��^<�xK�" uq�e� j_WWS� WW�}�W� �M���� 9Pw�  ��>�� �%����"���� �   "��3���E� � �E�3�@Ëe�}܃M���u�������#E�F�~2ҋ��  ����   � �\ D e v i c e \ R E S S D T     error   \ ? ? \ R E S S D T D O S   S� V�t$WjY�  �~8�h� � W�Fp ��h j j j"Wj V� ����}h� �k   Y���h �  V��WV� _^[� �h� d�    Pd�%    �D$�l$�l$+�SVW�E��e�P�E��E������E�ËM�d�    Y_^[�Q��% �%                        �  �      "  :  F  X  ~                  ��H       2   \  \      ����� � RSDS�o5�#@����TD��   D:\RESSDT\i386\RESSDT.pdb                                                                                                                                                                                                                                                   �          p                         �  �      "  :  F  X  ~      �IofCompleteRequest  EKeServiceDescriptorTable  5ProbeForRead  6ProbeForWrite AIoCreateSymbolicLink  0 DbgPrint  8IoCreateDevice  RtlInitUnicodeString  ntoskrnl.exe  h_except_handler3                                                                                                                    4   33Q3]3h3�3#414;4@4H4O4_4j4y4~4�4�4�4�4T5X5                                                                            