MZ�       ��  �       @                                   �   � �	�!�L�!This program cannot be run in DOS mode.
$       {m1b?_1?_1?_1�"1._1�21__1?^1E_1�18_1�11_1�-1:_1�%1>_1�'1>_1Rich?_1                PE  L �ܪE        � !  �   �      �`      �                          �    ��                        � 8   d�                            �                                                                                    .text    �     �     PEC2�N      `  �.rsrc       �     �                 �.reloc      �     �              @  �                                                                                                                                                                                                                                                                                                                                                                                                                                        �<     �<      *�����Y��!�=�`XW��A<�!���|.��iqlɪFS:u���\��H��!ݟwy��9[&�j�y;�|`!�q�Xpڂl>�Y}�y"ڹ<�!wƋ'V����r�Dhi�W�:x��������`?"#Ĕ�I��~(���?��"��HpYrȈ�d������)����â����Ӄ�[%s��ʹ��Y��s+	�Q�_��_nl�O?K�oZOy��W� ��-���(�|�`-���_2��M�?x`�"�K��� <Y8_�#�Ǧ�y�n��$m�t��`YP��2:
�<\7��^:b����9���n�w���c%<�c,yV����Wv_ȑI#r��QVC�I �^VI�lH�mAP��O�ǿ!�6)�%l8���}+�nix����C��;`���Br4���i�iҲ��SԷR[@��m/0�X �c'���Ju ^���͵����̄�P����2�(�:�a#�w�w�oH�x�/�MI1�g����FR�:tn%E#W��p�l��ٱ-�!�7�|�)�w&�0��*�-U^Md��v�8@���zӓ��> ���S�5-QRV����p���j���#o���fl��"8��~�[��ν���B�ĠX��.����Xu߬%���v�bH%��?}Б��I��Vd��� ����JT�Mw���L�K_���Z��-aVo��4�w�`G{n�<��N$C�	������m���r�	Cl~��[`@��C��uJs�Xރ�b����
�X�s�UO��ՒO V�+����z�6c2�����z&�����R)Y��O�į<c}N�J�ńS6����+�H�|g���[f�o4b j`f��YCӖ��F��K�o�I"v�gx "�Xt���r�LI���������������ZO��{P��cY	3���"qy��
�D+D�[�Tȥ��KE^���}���:А��}�G,>jP�Nh��S2"���v�S� tA�S�z&ۯ.�)�9��B�	�y���AP�<iuɛ�f�G�J�{^W�4���:1_��i*7�J�l`��ge:F��w*Q��Ih��dAׇr���ՠ?�6�`��C+�Eլ䘹m97�1�_���K��n�X1��/��˦3��S��g���6/=���:^�y 8Qg�����@��2�F�CSi��V�����Y~2+����q���2��<)��cV1�).�W��c�ѻу�t��(�j����eq0����rڬÿ+�Z���L��ةJ�i*�tH�_��99��.��n�b6ᢆ��h�Z>T���J��rVV҉�[�G�nm^!͙vD�;Ba��y-+��YB�>�X� ���]�L��$�<�6��
���n`��Z�a��T_�⅘� yH�M��9V
P�����s����q)t�*��5����Z%�2�!C� �9�o����U�^��	�T7��1g�9/Ԁ�^�T��.y".�a�D.c����{
M�<t�� �Xr�J;{�B����b�cm������KF;�5�y ��߄/�&\>:&�Xd�5�o�9rH�<���1�$L>U����8���}��6uw�_�À��m���uZ�C�6�o�<b9g�$�JQ�؂���5M�3[&[!��W�!Y�Rx=��H'^,�ׄA4wL���(���)s�%.dI�r�4#"�"3�L�x=p�ھ� ��B�ɂ�nBZA�R0�HL[. ��K�Z@4�ْe5q��(�Ş�ѯ��0j�� x�$�`��~4�@��h�f����{�NH�ܯ+���>Mep~r��<ϴ�@�Mӓ8���q�M��I��{毶�a�[{�l��]�z�p�� ��.���ވb�i���#�U8le_ ��LE10	��5�_��|�vs�̠�;|w�X�ep�!��]�O����h��-��)齼j{?����=�)m�m��6�G��+-��d� ��B��k~dY�<d��p�̂\�N3���%������Wà������/��c��gx�L���F�[��!u� I���
��o}��f59^7EӬ��n�|VbP�YY��#����d�Y��9f�a��"�|:�ۡv��o>��eZ:iߒ���Mp!fK�V���/����E�H�?y�O��)�V��l��b��5�1['�0P8��3�x;ph�Fv�_���?��cN8K̅A���+*8�>-��dד�䪂���΍b"��)I�~���[��Udb􆠑2]!]��q!c~:ch��P�D_P�鼖9�Օ@��AR�;X�\���`N���c�oRT�>e�z��A;���d�*{���R$��+��E�U	#r���f� &��r�#g���8,����y(�e<@_#!�r���tt�Dc�Zr>��T������b��h�]@}R_�eh�m s���	���(&^���/�g)w�ǁh���/z��^���I ��X�[7�nAG�r80޴���)�� ����b��JJ~H�V+��L1}>ҳ7�n��.�?g�(%d��Z4���2���XN� '(5��~����I��$hi,/��>��5Q	�����덬,��I�c�ͱU�(�J\�W���e2(��0�рI�$`�V�ruP�!�����P��vպ������jT�i/)J�;ug0?���U��8��w'�\��v���Wh��Gi��
���Ѭ��K�f�}�(7Z,�J���@���P���wgF[w���/H��W��\z�ۇ�2YiA�[�;�svc54vJ>�������e#8�H��4���^��P�O�6�V�(E��g��~����<���4F�by�3���K���qH4��]F��'�I�B�ֳ�����M�hX�%���%r~خm�k�t���O�����C5�X���ķ��+	\���[�v!�����l�����S��A%��ʆ�f�|���Eu�'OE]s[kh�/s��4���j:/�_��CLaK�o%�x� u9u���y��N��{���G��*�6��Ʊ�gE<SOB5�� ����O�ra���
���w����Hp,�t(8e�'��C^�����B�����X���:G!�XC�3�I>4D �S{���k���8�YW�uR���~k���xh�Oۢ*l����_��ɴH�έ���O����D��t�|bG�ۧx/���Ks��U[,���E��������a>a@TbSq-����I���K�_����Qu����3����c��_�����G\o�T��~�N��,bYy UB6p�Y@�]��x�WjR�:o���E�\�<B0;э�ό���8�x������~����+0��%Bxr�r���t���w��,��[�4
F�~�hR��6SMc#גدtwϙ�YM���(�[J���k�>-/B�J�����oP�N��F������ ��5����Im���W�u�)�N<���p���G��)cʾhxԞ�,��S����ґV�a#)��D�ʗ�	�t��w��K����~7��|&K=J�u�gQغ���F��}��m��;����<ޗ�7ć����=ހu46�R!���������<
˞nO0%�%�`�:Q��h �x�J����˙�E�V;B�ֻI��
�a�Cf|1���#|^ �c�E�n��M��t��t��6ۆ�w��Z���4z�Mm�~�X��Ԋf��D��ƕ	b�9�G��W|���f{���7�ZIn?��V��FC�����׽L߇.ɳ���Lfֈ���k]�A��5o���
�Be�����HW�Ug�NY�GK��������	��ǥ�JO^��5ipN�� �c��F��Z8���-տB�$�U���P�o���	�5Q=���6�%7lH��~�H`S̅R�-\M�NR�i���e�4J͸�(��饬B|ʊ�����l�K���H\5�w�Mp Z�x1��,�;�O��57��󣨶q���X��
/�h^�������h<���+@BV���8�R�D��������'��X������T�Iߎ���k��UXDe�$(��AK��:�.�Y/]Yd�����2���c�>��v��u�2G?<"p�o�$R�����*>��?��@S=�Ḇ��B�k����n�	��@��e�P��w%���L&�*�C��;�y�/���m7�j�t���_=���1F;f�P�h�Q�����VD�օ��m��!�Ҳ�$�'\�
�[Z�}����p��)����+�6]��.kߏ���ڧ)�)67�Fh��_ɪ�Ó_e�&=�9Ry �z1��8X �3ﭔ3�� 9WSa=rc9V�m�Q��X�4�W�vNO2O���pIJD~B�Q��ek��2Z��z�@2�G�ݱ��4�� )+��T��8tyT��<�P�r��SC���\�#�<(��.�JLI�K�U���I���  �,���.L�£X۝�cۊU�đog5]�]�/c���"��&��}����euJ孍>Xzz62˿���$��͜f4Ёc�9>\�v�39�M,`$W�%�<������(#����%&'���^�V-��)��Q�X=	��n8�n4b�.r�� �=�VJP��^�����l.-~��ᔜ�d���ɷH<C�ם�hŵ^�PjL�c��S���u{n��@�rc�d��d�ku;� �ާ
꓃}5e^��)����#��,4�j�C�+Vѓ��ԲtJ����x� �[�����gf�����\��~�`eht�lp+�����k���l����bۄM��斛G�N�n����B����N��[z��_��V�5����*�."+����%Ĥ!� �4HDR�3�+z/
ǭ�e���i���A�$O�@7��c
.�{qn�^�������;�Hn�2�Gx��h4���Ha��Yu#loL%C�X�^�#l��l��VV��VI��=���YLKE�����!�/����)&���!XY�Yz<7j���p9��#8���ʟJ�Y)��~�����Ӯ�����P�q��K�)��Cy��#h\�c�ZA�	��J�eT�2i�����+e�D�dHޚ������6LP2�����S��Th93�ǵ7�H�@������gGv�K�C:����p9��9��|��v\�*��0���T�h��2^j����>��������2�4j[r�}z��ɐ� ������S������jO��,����0p��/�7�MxY)،�zz��z�܊��/�l&K�>�Fݣ� +{~\�Tjf�1U�U�io8��~/�eθ�Z-~RS�?���?�'`�`��+#��$�/#_eI�X`�3p��<�p���l��6��M���+�[!��v�WT�'H[N��󄐁�ԥ��x����� �vQ�I�)��;k��լ��h�,�n:�З�< �n���S�b��O8�b3D?�DX��'�2	��UH:��nJ�,�Z��Bĉ�x�2��{�L�,�Z��� G��ߣ�B�@�{�`G�k2��ԣ(Xo�l�o]~�K�,A�:���j�#c�9��PDD�景i����g��=�y�$�YwL�l��O��#b\��㽃s�fEj=$F���I���\/>�/PW�.F�G=��D��;�*����O��!�B�2*xspB�Y����	%��9w���-J1`Z6�DTc��/����a�d��DO�8�2`.��:��x�o�[U� _t��t�H ��nx�'�-q��s:��U�l�
kc���*��QG,C|4�t�͏��@���E�h=�&�Ӕ}�v��s禤��ߕycLI�ACRr���*��N�#�������?d��f��+�}Έ�Z�������?�SU5�R�np��F�f���(R
���*I�X�XۇfX1DOL�����6�K4$�����#Aua��q�pz�'W��XO�����P�)Ud(#��GJ��x339F.��[��#Q=�G�c:������oJ8G�'l���H�s2P<�O�3�OM�Rt���)[N�?�����Q�o��ŰT���K��l��х&S6Qv�eF�s��t����l�/�Z�a��,����NY�P	@؍��-�v'�@�N��F$�Ԃ��?��gἲ����Ӹ���T$s�B��D_����7-	`suc;����kX���q,&�-�7S�o�+gdCsK�y��N�[h�{t���pP�@�V|�[��"�=�V4MJ؟��(�`��˪pƈa�YA<����ړ�A�K�NN�]�-(�4AYf�a*d�����c-��l�u&[��6ф�1~R�����n�x�yz#S,���T=w��k���?�ĳJTY-���8�1���%�۱K��(�"3���05�cr!�
�#2������!h*�9�3/-*����:����cO\_=W�� |Ҋ��m��o@:�&T ��ށ���||!�wB�Z�w�T��R���(�ம�5�_�M��z6�ٽd���h��r���Åd�f��Wq��BPD������i�,4����x2�о�F0�I9���CL�N�Jf�ԁY���������>˳]�PRt~�ڳK�����+sQ���%�Y��#��nst(;��%��*ʳ�U��9�&�9/��y��Ŭ��=�7HS��!��i}�7�a�*�2]��C�I�
�lF+L�@LY��C촲A؝�q����=S������À>#�g?O�"S�'~��L��-�{X�^Y  ��ʼ�����<��9�`��juʯ2�2Zc`�n����d�ӋQ�ɳM��j�8)��'G/Hw�d���"�r��`ʨT ��dUXX��jf�:e�cT3��t�p�X�3�S��_�a�`q<���P-=S��*|w�6�o���b<���l��,����2)C$�f2�$�}�y힦�R����=M"^K� ������rn�+����$9�f����i���e�o`��~N�PѲR������������ߌHV�\�|�L��g!���=����Ed��x�\y��p��z/�|�Ϡ�����E��L6��O$q�ʻ<d|W2���UA����m���	������}��:B�TS�	T��e*y�N�Z��2G(����(��%��i������S`ӍKg�7ocnM^ m__�l`�,D����`d���l�>`�l-���l^x+�*Q��w�]..���A���_�~�|�jQ�H]a/�[�$��P�n��a��;��A?+j��$�������-/1�f�i��%�[����v��~h`���1R-�����c��%;I����aF#��U�K�R���w�0��H���9���MIw��g��ܰ�"vɶ㼹Gj��o��h�����"tˏ��"~]@y�)�$9zTSf'5n�X�w腰R������=�W�M�p���9)/��X��G���l�@?wM_fGE�j?+��@2��_Svg�C�Lb�x��3FaE-nYkaX�/�	E$�������S:����Ԯ��Y^�I�E�LR-�)�˛!O9�B,�*@}�_�VG�,�f�0!�5�.��p^����������X(d�FdN�BJ�.v:3^�d�����}�����<0Li�ɵR? ��H�K`y��$���u"a~u)�"��uf��'��_�q��Hvv�`j�����W�LJ�b]��&a���K��2�`ϭ��Z���Y��m�������1��1���p�u�[
�u���@<~��e�z'q�~� LQ�M9͡]��"�&��ʣ��*�	�ܲ��I���N]�D��+�v��]��G8��;5O2���LQd4�b�n��zy�#�W'�9gb�7K����~�񴻠C��J��"=��	�xH��Gj�{I�ȯ��p���<{+�n|�W$|ͨM��>+|幕py���^q��w����/�@�e���],�~�ȭ���jV�C��d�u�U3Q^����4{;�
��=n6#��2[f����r������w��H�%+�>u���pR([�13��A�$
�J&�"���U�]�G�=���P5��k��1���ϥ��s?�%�Џ& �<x��C~n�	Lj�JbI��2U;�.s��q�l{�<�����6Y,���A��!�h�ῗ�<��6VYT;��H�@�C���U��S��8H�%�.�]���b��-R#Xq
�L�>��]���4����Yd���-a�B�A�Pl V�V������+�E��g�u�FT|��^�?���l�V���5]�&���h�d(]C�bC	荲�~����
�n� �&�M�X�ަ�%�xQg��*SM��P���K����g��_�M"d$N_�l}�Q�D�%�����L���$��eMAn�J�s���ʧZ�X��?�H�۳�{�2X��0m�^;�$��kO�1D�o�<3�n�4:�Șn\MC�1�_<���*~h<d�k���<ˢJ�e�4ۋ��VtĦ��ؤ�ű�VMN3Փ�Y�K$<���n,�5t���?�9kc�<"�{�H�S��#W �멭�`��a\�8�����c*��>�F�tW���?D��<��P.ik� ����4�P��:�n:�/\Ϋ4�M��3�N�u�DY�W������D=��ڝ�Y�cݚ14���x�h8g>O0�U�}_R\=�u4"R���<��y�� ��Tw���^�ȫ1os��x ��#��s&{�5�o^ʋ
�fBg��p�&��.t����G��0O�tj�J��t5nz�q����]���	��0m}������2��a#���z�uWS��N�jK!9�ATq@%����p����Մ�>�9��i����T�2�^y����ɞUv��mF�O�}�.Ƭ3�}�oj�G+,�:4/
�!��H�r�����_������X�c4>����j;$S��$[���S�y�_+���si~$���@+l�1Z�;W�I�NeP7A9��ܗ׸2�6�{(.�>J����#��=\���?At���h�v�ui�����-���VM�l*Ks��	UA%Sއ��^��C"IU�uĪU#��]���ʥC����6�2h�9W�?x��<��z��".�¸�	L�A4	�5�;GRO�5�C�x���`� g��ld�a1����)�eY���o�<:��Ί���	~fc� '�7ѷ����9��r
���u�uE�CW��g��ը&��I��q4?$UZ��љu�
��r&E�N��B�v�_S,D������{l3�'�|��\+�vt�k�HR���tΘ�<AL��t�e�@��a;	�Y!��W4���EU8�	��;��8X�7�F�P˦O��U������D���f��P?�u3��B���O��[��k���/}9��JK��Q�µ8�� ����+����(��c�KvW��se��	�0�v���h1�����W�(u���%f#����Y)�O����\�o/�J7��';!$Q�d�Q�m�t���ya�*�́`��7^��`�BF<� ��G0�L �v��S��&�c�x�Q�g_���b�~�ֶ˽������)+IE�m��u%	�Y�dt����R8r!k�� Wg���:�V�ctK��iE��E�x/���ěR�\?��@���#3��I����t��Y;i�i��!|<f��e���X���D����#�σaq�]�$2�D��&�N�|u��O���M�GV R?٧-9��"`��ʨ�'�H&�:;(��v��|
�sཤJv�Cv���R���w��BO.�_rlp�lYy���K%n�d?'���m��[ynd[ze�l��ќ��wΚϡ�H��P��d���f9x�]�ϔ��*�57�8u��-�^��#P�Ud���?��j6]�0�îן ���������}�Z,��l�ؗEX�8���� �"X|˓�&'��ǏDI�|`l�@�Z�v�w���BJa�G1��ϴjo5�����0��d����|�-zp�?5�O��A"��D��
�VU�ى���O[Q�:e�f���8%^�ʛ�mGT��A�I�to9�IIE�[���<�W��mȩ�̇C_��8C�>�]��8F��O;%�ØDMǉ�Sv�*ѹ�ĕLm��D�~M8�%Y"/�9�pTfz<�ϸ�3w�ŁөGְC7'��W�mҲ��gT>��5��k'W�������ا'�-�l�{PW���'��mz]#��>���b���Z�9Xf�-ޓ?����{hs:?����^-W���_q)���5��m�⁖�r�ޣ�l�~�3d "^%�D%x�7L54\�DȄ/��2�����y�XPa�$я�eA�C��dO���u�x.���E�$��e!F����ý	�p�m��}���?��X6��,�#�#���X|o�A��^A���k��ggC�TO�?�/��o܄0@y�a0z��;E��)�����+bN���t�Z��FuInDV^���ѵ� �>��Ho�У�:�m�-'�9����'���Y*nh����s]��!.w���l�}`_ߒ&�q��}���Y��k��a�@�>5����mX��:Q���Tv�
i��S��=n4�_h�tG�ԃ1&�����3+#�U���/�;���3��<��Z���AE��IN	[�7�Ó����� ��g�ڻ+�Y����
;�V��`���р[��%�\�ވ��p��u�'�k;�^zilw��f?aætk\��nٱS�>+�����Lb%19r��Ή�U��_A����Zj �5��D����V�u�1�0�U�GF:�k�h�(}��Ä�zRlCW�/���T�\&�-9���
���$Hs�7��`̱I�A���J���>zj|0�eì6s� a�8/D����q%:�ܜ%Π�A+޸�����%���Srץ9�$��>�r6��Ĥ��_���[�}^y�Շ�ZN+��%����I�>r�"!s�	�Z�����=)}��C�R�yV�=	L��s�O:5�(�U׌a�<D&3�r�ݮ�%�W~˺l��ޑ�VH>m�V��v*��4�K��[�ZN�Jui�����kg�	wX`Y�Ո��}L��(���z���F��p|�l7�CJ�h��t��2�� T;%�z����ނ�Mm�A��V���ku~��r����|aI��q������3X��Rs����.���/��=��.B���<M�����2�I�����2��d�E�^yt�i���C�J���RR�QZʙ�o^Z�j���Xz���S�F�s�^]��Hh>\��2����s�bx_cl������WC�Ǆ<'�F�7�Y��xO�o<��l�du�2��*�V�,FG)9#(�>��6�����lM,y[��>L���#.CR�������;+8����d`<Ʌ��-�B+���5H*$�o>f�#.�d^��t��[ז'��.ݠ�͢�g�.�#���W��8�r�|Gפc��658���an��pl��J���
�2�a�wr�/'���dj��17�TFk��	��#;-Ԣ_��b��O*��!6ʏ po�0�]TBUj��9Y���(MS��*U��x���&��
�w�\C�7�1$�L1J���������(���Y9�e��b����Y�2c;���C;ؼ
M2�	.5�������ؼ��;zp������Aƙ	�|�.��*(��	H%)68�t�1*YG#�\�tf�*"x�'��Kv:���9"3�M�p��3 NG2䤷]�0a��r�l�F�m4�'��r��_Y��D�@k�������i-�)�N������>b޾H$�c�ޑ=�r����d��z���e"s|"`B �"���#3�z��{��Z0�R(���Ou�#��
8E�a��m8�L�8Q�'�1� 7�ӱE�7d��4�%��ֆ��.�#����7bY������b�5�7e�tԂ�w�zZ���ט
΍)L�5�@�d����1Q��I���3�2��ۅ�t�̟�R��@�&���s(\:��X�̟���T��fC~�	 {�d��~;]A��9�0m̠ǹ�?�&��[*�5��Obk/%&�)��"�QA�ĺ)���Ӫ��+f&j�G�Iӵ��3F��������N$܆bԴ��Y��m0OZ|���4yqQF��6>�wǵ.�؃,���n�G��:�Y4-z�h�="z��l��r�8�"l+'��
�xF�x{�$����펛�Y=�3��/��\�4��z�?Hp̺���(6�y�ec�8ݔ�քt+p\8�sB�Ԁ��lu���D�Ĵ����	�هn
k�玠�I (p	u�8�X7#�׌�i��!(8x�
f�d}��������RM����D&�!} lԬ��d
8��!j�$�G��n.��J��}=:#	r���Rt�V��˼��R
��t���� Tݜ��#畓DQF(�,�q)z�����>���8�!Y53��;̇!�Y�0�󪸴�Z�U�BV�_>Ӹ\+���٪��)Ik� q2_��l��K�׃Z�@��d��������?e���ۂ�.�)�t
	�.�#��qϝ�`��n��ٹ�z<���&�wG�h������"v-�2��S��!���.�Ʒ�)�Z���E�a~�@��Y`��P�M	BW����V�?`�����5�G���7G!���&*��RT������P���XW�2��,�D����&��43W�
�Փ�/�*�Ad� M��A1�Ϩ�5�̬�<,��H����62�AC	�7;�k~����L`HI�'(���#�uXA�sW�9�4k���9�2L�:�z�{z��0�^Y�3՗S��T�Ǆ�v7_�O�,,C�l���
 ճ����gܚ%ޤly�K����t��M>j#k�m�:F�Ẋ�d��Uk�ƞ�큹j�sAt�$L�����珵��1'hډ?W�>�g��$XQ)ly��&Uo�@��؃��PZN��9��L��l˘+��@H�7 ��U��S4\1��9b���গ���Y#`#�H�XDu��eC�/��:�D<�_��@N`t^5:�6$���_#QN��
�#=�m�÷f\�TU��Z��W+�[z� b<gZq�9�D��	��u?�m:D�����A�����!	�����!��O �0�	fP�.�# �e��+xnZ�b,����� +\��멛)�S�uL�lC�|��ޑ�
��+�x��y��2�޶�Z!Y��VrJ�.�?$q�E�t��]��V�t�ض�x�	Hko4��<Ь�~~�R����ƒ�m-������P�^q��&�	:Yl�Ecn�=��kYN"�-e:<��6����g���!�>v�$.�2��mֱi�h]���0��P���ݬ8E�Q������rwU��,�Z���Ē���00k�t��~�4f�?������A2o�Q��IIn�ĩ{k/�|	ޓ~�	lҚ�n�%p��Ĩ#1�TNA!MrҸ�G�l��%(���;u0���z'i�Zf>*0�r�K�$F�~$�ńؽ]�(�1�t·�y� ��2��CPsx.�t;�bN6��������Ԇ�D!�t�{�~��4��,d �{OS�|-�ݦ�#��j��{�m��EY'�2��
�=1]��;�^�W1d�C5�(S�~��8���a��A��a�P����30p  B�KNc�2d��|ʲ̎��l�&�ъ}2�oO�]է
�:�5��ލ]�#x�2웢�N�.���ϱ�5�ȑ��Fc2㒝��N�{u��R���I�8r��sΌ�+����c�m^���tYD��_�̙�p���\R��_�j����+�#k��T����)_Y��$!�:�8�@݃�x�<ɳ$b]z���.�z�Ÿ��a����i��Ke��Z�UT�MU�J�����t�b������h�R�_�;ሷy�Z�K�o5)0�w��*[:q��l�Ptʊ�ۗ+ҟ��s������=�S]�w�i
��z����7_PU<$��r�$VC�L����~Ĩ)"���x���1����$�p;r_��pbHּU�U��`\�ʈ�o�����An�`zrQ�@�F��*��c���5��G�ʏe8@ 4���-����"jWڅ9W��_�J���d�pG��^SLj��_�"�O���O��<��M�UV<t�*��m���t��]M+s��lb�	��
��ۀzY$*ǵ��,��ey��Q�n�#��g�%��SKRaƍp@:K�r��z;K��O*I-EGB�'�s���(;�aw/�M%�.j �?@�e�����6�R��m����'{(��P�;C����^�}�N�^�P&È�܏�%e+&a��q��I�0X�����h���������(s'7�`�Ƨ*cf_�lq��#%v8v�V�ӟ�E�wY�"�KwX�A���-z���M��"9��$�wbAe�A_�W��]H��v��r�I`]>(A��K��K/�V�m����.WUEk�ۢ;��kݔ�M��Ts�	���yl,������������h͙Ǔ1�������l��W��lZi�4|/��nsC���p�I#wr'�ߢ��ה�,| ������pv��)����HS���L�Crv/�����JQ,�6��(/G�n΀���nǲ�1'6�4#����E��d�~*���V$�DN%#��b�[�j�f=�GM�����r��^Υӝ]�>9���ZgS%��K^�%�loA{¡�����ˊZθO�/�_���&���xs�Y�����n�k�EWzITo���Z��Y���=Y4�R�%;�(�u���Tn��+Fy>�\��ІD�Yc��7��g�%VEq��Q.��s�Pc/���!:��*�@s���8tܽ��Ǿ�I]�%{�5�=B�e ��}�=��!T���RB���4�8�$jLUl"5j4z"�W�"&�i�s�rHކH ��	Fs�-�>
qͅ/e��o�"֧������F��R&��2ūak�;�+ˡ�i�Rg�#Ng����&�w�_���9���l%��O�)�Od{�eL�pu��]ݕ
#1C7��.-�6�e��|>W�G�<��e{<&()�=�TMc�=4T�Ih\�.��m���Y.!��������6K��Q@�����X|-��߿b�,�*���c>mYe�*�:���tַG8�bF"zh��h�z8[�y6hd�8Gc����eE9f�nNE��N$��m�DPY,9�����Q��Z!�쟜����M}�}��HN��W�YQ��φ����b�G�͏��ЁX�Õ7�K����Fe����>0�䢓<O��
�~������䳾y��>j}�]R��q�t���R(�8�;�#Z"g�3��2m��)��1J�Z^�U+vO�D�x�@|'d!�bn�F`�eKi ��9�)�	�ۿ�'`$?�j����H$כ[�2��c'��c��v5�B�kj�H	�u؋������FG	RIX�j����N�}Ͷi7ܥ_@����S�p�������v��VI2�%;a`��w�����؂�*���M7�#�8�UB���˴ɸ��	��i)mMi��l��U���������>˨��j���b��
ח�q���Жf`��7�N@�:VGS��ߘ��5�"����ktA����k�H�jk�����U��EG��f.DEq��\��X�S\�3HAk\��[�rY4|�M�z�H�r��;N��[7���qW1�M�����~�0i��<+X�i����S}L�`z���ԣ��{��(���Gղx	�����:�(�VX��>h&F��!��ᠢ� �48�$|>(����ر5|t]	^���ذ�G�jR?×|\��#4�O݄q��!�-��7�R�0�>��	ڸsj��+���y������W���(NX|�ioj}J�����3Gšc���泶������Fϖ�Ar:����>�s�e�k���l�i�`M�e6�sl��z�$���^��83$w�	�Ղ�!�j@4�����������������D�����pO8y���"�����#<c��N�U���n_7��v��P�b1�NJV��N4�Ƴmg�*oT0+1;Xƺhp��������a�Vm�^�f|�p��^��uJx����
������~�LH�-�N5�bK&�bZ맓�����wuo� +���,"�t�����,�s_b;" ^�і4�F����x̃Jj�	*{�N2Yx��%��9[w	�ꗴ��'ֆ2����D�o
y�
M�>�k�T=mS<��Xɞ�Դk+]��{�*"B݁Mf%���A�/����YBR����P�s��'wV��D�ۜrM�n��Rxg.�|��ŷ�Gc~ӛ�a��a���o�+l������n1g\U[���֤�2����b��U�,�ۀlA�r����V��M���Q�LÈ��a�*.@�����2�i{�5=�`h���x@�[���3�d��)n�񻸯�ۖix�zM{��3鄍�VrΙ��cp�u�5hܽL�Y��r�F lph�����x��o��&b|��]t��Д���WDu�B��(	n(�0j���W��a�_�g�⃚��)�ҽJ�.������[͍*϶~�´��Ĵ�s8��;+��^X�N�y�#�Q����~�4K3�R� �=&yj���` �a߹��N+�Tō�_��똓��1�]'�a�q>f�r��Տ�8�7���4�u���WU1L�;߫��j�z�fԷ&F�Ck�tuc��ؙ��≇I�a��0����v:h�9W�Dh�o�f>��ɐ/�цC/%��VJpǊ�#N��@����\�o~f-�2���}'�i�-=!���Q��fG�.X#ӝ�������Ȃ�Y{�Hq6-L����O��l^$$�Z�,>���Vܾ$���C�X$ŀe*�\�[��wl��nhwwXWk`m3Gg>d?�_B�>펒/��(;ITK�k�X3w�w�cg=k6��+�|�VrE흱q(�T||��l�~�F�$a-��z
{r����'2��|�p�m��� �u�]�8��u"|��PTz�?y��Fϒ<�g��7����O����xPݑ�$z7�_"H�-��09�i�1K��X
�R�|�����E��zO�Y֍f)ra��Ќ\'���LB�q�c�8a�rȀa��̡�[ﰰ6`����ʭ�RfE�I(V����Gi���̔2�0�
����-�r���O��R&�
rfhp��̅��[R0��RǄ�:��xwhjɌ)�;��8��1~lRb:�_P`܋�p�H����	���p�7�J�͸��%8��3��\���� ~�MH�/;�<�3#��F�=]�a����%S:! G��K���69�����[�5N�'!\+K�KkT��*_��ǲs�ݞ"���x|�ձ��@Z�^@�I+�;]6T�֠{���X����J�"''*%�@���cz����z�	nqM���,�H�Q{� ��@�|X�y =%��K,71h��L���UpW�A�&�f��6��#)��r2�<�}����U �l:����������m~)�Uʁ�I�q��e=w��D��ɹYlxC�~g3ѓ�Լ�cQ;!�r��]�AAm��Pbƒ�lb �/j	� �R@s�O�z2W� U>���
�r˹"C���=��AKګ
�Ɓ{Hyc�wJc>����{_�9����5͊6�2��C�1o���o�����O���9k k�+O]ݬ=4�����؍��y~�8*�YkfA(�S���ĳ9�nL�=�
𑱫q�I3s����6�����N�| Z��E����C�-�Gi�H����K���z���l8�}����v�V�#�0��u�&?����J�ݸ�t#�\�=	'A��=�G�~s�	�-�0�AP��������\�c�N����hv=����B�F<,�D��_:H���oD�����' ߚ��g|*s>�l�(����w�l��ښ� ������5Z1�X�"զ@�nqj݌=��r�ƥ��5�q�yO�9����K�2�#;T��%x̣���d
#ס7؋�Q�L�}�x��ٝ�ٲ����ݯ��w8$�%JOP�6�;�tpu��9� ���WbT�Ih�1.��Up�Qoѱ6�C2����)R�9`'I#���k1NSL���(�]mFk� _8��cu�cw�3\��`��nV)^]�+ÎO���)8
u���e����=�pH�g�v"��2�<��o�@��n�[��6j���u���u]{��ͦ���#��=��#l ?�(J���B�Ѿ��	`Z�����[���,�o�h�d����3R%j-n0��	.,�]�W��PU^TU�a���iڞmv�!.̏&Q'�fY��P�w8�������f�2��1��1��b�A7rcFu����莣3�ez}�\�� P4"�xn�Z�A��ፉ�{�	o���-�ިF���%"�8L��zG�<iU\�C��: �����8�x�gݑ������j_'5:-y�u��S}j6P%$��l�)K�{g��`G��ߐ��4�5���BVјm1��M�G��	�]�K~!�֒��B���[mw��92�������A�Hm�M����5�����V�Jo[������o��Y�Y}��,hjiTL�${!�����%��1���~�g(;~9y��QaF#���(,����Fg��q�o�SZ[/M�H��a�,l2��O"���Kjv�6�$t��If`��8�*��/M�O�4�-$vheA�Έh�-����������QƏX/ _@����m ѭPz�+SQ�Qs�~7��·�*������7"_��Żas���j�~�4󆾀�,�� 8������ʓ<#�1B��n�b�����T����g_8C�~�+/��Ԝ#��E�t����'�p�.w�an�=E/JE,/�\ˍZ�d8�#ߴ\�4p�Q�~�T�7j{G�EB��_��tI����"(�4�,�֌�p�A�j!�.ޫ�EO�)�R?���~�,(K ���3��;d�� ٸ�&�Z��z�E���oq�}U1Hp6�xw[��)�*	f� �fD��"H���(�lGB�~:987�QKؙ/�I��N���M�:է+�֚HO�6
;��\$���w�u\>�pY�[�U��o5g�U]� zC�_�"�l�S_ >`�?˚P\�����Ǖ�xҰ�A@��R�j��������n)�=>�07b�rZ���%�|>i=������p�5���4��.ㄜ�j%}��p4p-���q�:=61
\��V#692g�t��)��xNY�$����ם�s����]�Ȼ�G.�K�9$Z�F��# �5�([�;ly	���=���1��a��m9܋]���($�yp��4�J�Kמ87��5|ɊS�u�8���7=�5�>��U��_�<��Y#Y����VRKs�i�f�o����-�3��<����d����z"n"y���f#�6@K��U�3ҁ	�f��\���r �愄�1M�x�oE�<�uWfd<j���{Ʋ�q��5�����e�1U��VV�@ �㕁�'�\�Ku��=� 6r��ٛב��fN>��
*���~��/�!)Cl����\�]o)����N_!��%R<�_5�}��}4L���ZO����O�ڿ%U�i��O�ď���w�F�sl)��o�X�|�R}u�JX���P �w�5���ц���F�2 ��Q����W�!^	�e*3�=�e���6~
���ЖXL�&Rg���KV'KPݳ����
<�a��JC�Z6�X��56����_�R���=�����8�`�d�7���6������bWH�T�dm#l���N6&��0O�m&ḁ�'&s~-|��m�'觔��D��9==��[]Gז��];p>���&N��6�	��j��lH���^?����������1%v؉]���v���w�4d��UbқU��A�r���Б��R��s��ߜ���|<�c�����\��8�p���$0y%`�}c�l4G��������	���?��rt�c͇���R�:���S�8+�!�����l�#�)��r�9�i�5&
��7/����W_W0��seC�[:��m��MP��Y�݅�L������ ;Sx�n7�4�P�jR�_@�Ecղg4%<��tJ'�jA#~
E���[�dN���z΀���`��ZxR��ɻ��?!#�d+/`RDj/ӸL�Pd�5    d�%    3��PECompact2 N��(��F�>�5끹��l+�
�U<}G���-Ar��r��:��UL��;�ΚYهCKmgU%h�C�����AW��*� =��=��K[G��ǖ !a���ԣ��x��Σ{�{�TY�M/��6��(�9:��Yc$OMў��jڗyX��-�}��h�>��jKUt�����;��Υ��I]ι��@��`o��?��#d335Y����,�����4N�����
����"�*�Ɓt��e�����OrT�59s^]�)��͈3BAj*g�Z<�a�<hO�H#�S^�D%R�y�zh�\-d�e&�Z�S�6_���>�i䓅�"3��u`�1
m����I�X����iS��/��3F���mX���'7A�j(V�y��a�kl���P�a��G��%^�@�M�ڴ��j�zF�L���A'�wX���1�zbm����/���}�4�B�)��B���5/UL����2G*�� fG��$���{z�Lԥ��a��*�[ݟ�<ɷ�RԞ��7���)�����!�Cp-D %���Ps�gpRz�n�L�)0WV�v� *�M����� %P�c�}�F�Jϣ��>r��$$�hC6�t����θ�9Eo
ñ&伽ཿ��U�ʡ�bh/Rd�0�H��F�Hq%+`���gY����]WnҊ���鋔`��,DZ
�>ݎ����dhiW��KҲbH���B���|������4hxCQ�ky�����tp�3�j�#��>^��/t�Z&k����4�t��\N�����J��F��]��IU�+��坪�v�lGhp�@$�u� �N�!V��c!h�*�kD!g��Ȳn���_=�:娿���K��T<�f��������3�S�Q��N� �Ȑ�H��p9�o���Hu�M� ��( +\�'RL�d�/��b7Jߋ�yl�/��[��l��V|�?9�2��P�@y�F!��&��4Lm�g,J�s���%}8�rS����4�!Rh����U����J$�B@#T"rcp �6$9�Y�DJ��j��nhv�/I���(^���`�-�yv�u�4�e%z<!n3���5�s�3}g�o��JJ���M����.��o�Ph
毗6��3��-o��M0L�de���S��KBՇ7dث���t�<�پ+�8�5� �c#�Huǵ&(;�_�˶��68�c��O�IC�we����!&�xr���P40=̎Ք�+gȗsWW%�����L�۱�%��#�ܪ��Mh>L>�k�g��)+7�(�,[k5g��c��+P.�"Fw\��W�i�փң�˦l�)���R���-Vm+ތs��_�ރ�v��E�7���܍�U;=ݲ�Z�9�EaEP�S�����3�W�����s�-�%+���W_i_0Jzx�Ĭ���,�_[|"u�#�[[��+��jٞާ<S�t���=���
I�
���֕��q)�n_��G��b
$��0�]й1�L�,�|l�����O "[vG����.����7�יĝ�G\�����_�J�Gd�ӟ���>% %�Y7f��v�\�?�ԅa���D��6B�J7�K!��O�P'/-��*�[+��p�kAd)o�@YB]�6�l�V<'5�+>�8�_)�!���ܬ�V� Un*�l$�ّ�C��q	�i�+q;�M��wP�Ž�EK��-A��x2�n��Y�3�Bw�>Vx��D=��y����>K�Ŧ2�8�:2|f��$L�!�^y�Z�:�����2��jCI�@���_,;U���|ϰ���E����}[��O����+�� ��r&%n�N�a�H5�Z��b'䅧����0aY��>��2h%�{�	ë ��&��Pd`�2�4�JA�BI7g��ld�$���0�p��J�X�}�JǏ����\�8�9ޮ�hY(�0X�!���8h���
\'S)�5���NWHaUf6�c���͑Ȯ��9��fhG�F���u%�j���Ȉ��l͠PfwLb�4� 5�c�u	�ϋ�ҙ�N<��������B�4jo��|�}t4�%VD�68��=���c�������\%���|� Lb�՛�g����+��o7�Ҋ��dP�{w��V� B�]���E�W���	�,jt��vS�	�$�����5d�a�(;Pg�H�QJ8f�	؁Hb��n[�����ᬸ�%��L
EU�U�BB~�K�T���n��x/� d��v��9>�_,�ɸ����h+;>�K�"<�Ć�GJ��z�(�E��bZ��7����e��Wírb==�U !�. _��'�y7eI����B�X~���#x�Q����"�9f�EN�l<���}o�1��ؾ?��M��d�k�57��k�+�t�ya�����4�h2�O��m��y�1q¯��Z) $鍇��nF�S#�G�iS>��+����l~����&+k0ó���E��	"%P�6�{��̕��i8b�_�$gv��2�e#���j������[	R�D`"�qZqʅҹ�X��_��q�ò�D.�v�f�zIG�|Xm��jm)
o��N�8�6�p	�˷n����z)��]V߰��%���
kf�9q·����W���N �O��+Zy�b~�1�� [��|:�2�&1,����e����4�}YH=^�j4�,d�<���@w��-�z�;}�xn�L<o����a��\6M�%�L�q�1|iG" jܴ=����pܐ9�G�Z�����.,�"��EK���o��CXa�s�8�5��CN�B[Rx�E��
Y`�����Lӆ�(�V�캉�h����Y��q=)�:�s
�l�&�M���ٹ?/]f�c<���|�9��o� b�Z�:�V����ka8Kv?��ӼMl9rˀ�r��42�z#�i�K�����S56����?���`�.�xl��T�j��JT|�&<��x7~Y}t�KF<��U����:�Ճ)k�[���M��������pNF��}=��00�ڟt��H+K��V�P^�&ll[e�+��;�������U$�B�},�'?n�v����F�v���J������p�Q��^��C��Q!�F5�j�k��}'��@m�0��P�>�r��u.����j��K�U�w��"������
���^��AM�҇���B�9�(K�5e��d�L'=����a`K�|E��L��O��m��No��-H�-5E�).&�Y�d#A��WԮ��K�ޯ��;��&�; �"!`����i$�O�!�E�\x&��{����3��Zv�)R�p�L�^m�)�l �������:�������%K�c��kK�W½W.Z�����%y�塇I�AA��Գ[^}�_c��cZ���z� �n�Xǚ���� �r2�'6�3��뢄ٖHd���,J�]���W��=���%�cWt?kF:��nY]�~<5Cb���([�8O7������3dQ�􇳝s�q�F=���� %�s�k����/�ay������5���\1+譇���JL8�JZ
�M64w��Ѿ�zƻ�@��>�F���=���i#%��&��e����b��e�J
��fm�{I}ːv���Ӡ�")h�UC��p�f�����.6\�,�?�D0���{��������d�#m�{�w�e�x>\�4�Q�
�/4��E��c*`73�ޞ�45�Fo�hlf�\�ƪ2�(.���|��җ��)�e�q�m��/zw�! K�����(@ܦ��C�t�%`)�H)|m���Jv?@Ā��Ya2]��U�u|~�ʢ�&��S�~���Cf�4�jFz�T�mĜ�Ԍ]��Q��jY�A2�4 ��k�$���Y��5dB�~*Q����������%����s���L�� -C��>�N��lN�*Ԁ.,��Z����V�FU�u�z��T��VL�˔�|���v&,�s|�f��F��Cfr�K@�Gc�+J�4�t;��fK�`��T���2��M3�?�O���YT^�*Uv�W$��"�8��}[�=8���7�5���
�by�|���}7WH#�g�W����W�g�L��	�7\�xFMُ^�$�Z�x�(�@�t:~��N�/�q��r$���~�;k��jy8�O��n]�fHR΋�Y�(�S$����aڠI��Ӆ^���Nq��6�)��e����NC7��E8"^y/LPӍ~N��uW�4O��.Q�3{YV���Ʉ�|�V���z��$Q+@;N�Q� ��`c?���a��Yi�'�9�����o4q��� �K@]���2Z�$߹�Vr�\���1A��|xb�R�Τ��%��qq�Ep�-'��D��'�[���~��&�1P�6D(`��6c΢ak /%Ý��t�q�䮐}��f��f�,�B߆{W5"�Be<�{��y��I{K�v�ҷf��N�@�=���-'j��=m.���$��������y(u������acJ ռ'���\h�>���H�|�vr<@\!��q�tY��(�.R�ѥ4�(7˅p�6<���?��G&:ҡ�^�!v�Tz=�"����k�kO���%�g4��}��!��'6\�i�e�ל+U�ā��n&�4�d����q�O��PUΧ�N��C�)�A+6�I�:^b��!t5jY��%?@�~���}n��a��3Yh�u։��YG�U��!��?>����1YA4�����@�<����u��R%������´�ᛦ���W����!ֲ�1�wA�\M�J[۵|&%��l�4_��-;��!��7X�Q�ۀu���B}n+z�5�n$q��b6c��z�����Kp߉��ǽ�/�[ڨ� ���������*�lm�n)lϘЩ���Y ���=�Ӗn�"����Xgt��f/3gL�s(�� +�f��t��uF@?	c$���L�_�&�l�4�z�xA���e��0�\�n�|��ו�8�dw��v��Hz��@J�6H���d���˜�Tgf"�8e��X5z�v5�S9���K ��@V����2*d]�B�f���r*s���
Y�n"����)J�<��s&R|��d{��8Q�m�Y6��l���nCK�",���H�ټ�v��C���J�?!��.ٽoDI�S�_��Pݣ�]�ʊ��X�)/��v.��gMXq��y�}�ܻ�e�v^kC�7����LΡ7&�3�%��9(�e_�|�l�z��L�=����9`�-���:*&7��?�1t ]���XP��w�!���X�Q���'��r���ҝ�$%sa����u ����_])��b���~M�Z���IL�#!ZS���g�nS�Gh�.o��I��w�D�ĵȔwg�W�_�O���k��C�2m-w#��~)#��H�<b�zU��I�{B��a �w�AD�/��"|s;D�:����ߞ���$�C�A�3����|#�ʵ����*[V�o��2���KƓy�3��
��.�����j�3�"/��vE �sO�}��a�T�U`$~>�]���y�]��'f�29G�*�������q�A6�������[�[���+�K�:
'u.��I�	Ő��^.�b�O��?D���V���}+Y�}���;��9鰈Ws=��=�� |{�	�N52���"�<h���Y#u8���@��m�cY���Sk�
�2���Hk��:����T/f[>{w��HLI�,�E���_m������9Ny�`ؙ}�WL�aoẁ���x�T�s�>Paﻟ+��3	�ٷx�^3OM�/."�$�ġUh�9�����W�t��~��l��!� )Y�L;�*u���$�D������7s���keҒ�mW�1� �Iq7�<|i�c)�j|�*�*��;��zF �G��J=oC2�nP�i����IFz��Slrx��B<]���ҙš���+�	�E�F��KIO�7U,j���U5r���/�W�U
M%�0���ʊS]h�l����)�� @D+���ct�o�1�'A,m��?L�`�|ͺ� f���Hl�>s����O{Pנ�*.��+~��	X#��$�*&Fw��f*�+;��V������p�@xچZ�sb,lh��?�\�{��*<=.���g�1K?��R�BƁ�7�.�e. ;�`�������o��
����FK��P�:�i�B�H(z=�,�is/c1����2f���Ye�P�f�����6�Z�K�6�+�^����?ק���@P:��w%XU����0Oh�tm�I�Q�?a���8�l4����J����hH�2��nL����ÿFߎ<�l�b
��w�BmP�<47�@Dx���d&�o썺�j��-@�$_ш�M/=v���)��i1_���N;�&��.pc���μ�75��K�g�=�� �yn�L	g��b�ʊ�=�~=I�e�r�&�9"j�22�/�ڛp��m�U� ��g�Q��T݄5���X��4f(/��w��H4� a���67O�����\�S�{���3��.�{��MJ���]UО6��Ks���S똌ѥMhd.�~�U8��������a��I�" <lV���t]��}�%vZC�%���0���^<?aB��g���R~�1:���+J&���߅�[�C�f��rv`��w&We�6l��X�O�	��6c��>�ܤ���|��������Vu��[�A�7@���gCJy�m(D���H���x�KF�$�`���Fl�q�|���r�{�1Ʉ~�ي\x$ G73?#"t��oĭ�n�dϼ?��D�����˧H%,�5&Zx(���9Z5�"J�x�"H{��{��)���GQ�"��*G�tƃп֙��%/Z�$�Et��	�D����י� �WGs�Fs��ݬ�7iS���*�fK./LQJ9��_i���C�g�zaϮ�Й�5��OpQN���M�0�K���N����`�H$ǞK��H�dX�.' �a��g���-5���2��i,�&~��;�f4��3A��	���/�������t��yj&�w�^ �	na��T<������xH�B��ؤ�����z�ߓ����/x���/#�5�)��0�BXD���&���OmCE~@Z�<vtHۍ ��c.�#��["�v	pA!~|E�������Pb���0�?UM'q��(�e��Sυ{q��������ܭ��w"� x훞ۇ� �q���A"�f�@gv9饍6��!-�������(���Nu�=Υ{�u����P;�	��Bc�UMa_(�y@��\�ft��0�y��~��tލ�:qE׋��= 䙴>��F�r�Ƞ�����T�[3�0C��.q^�%�'�9���1t�V릲0s��k���T��e��C ��j�|)#���|Q�a��
שWl���,�#��v%8��a��)x�^fe���ۏ���f/,3��"1{�+N6ʇ.�[�0�	�2�k���H�O�p� ~rG}h����͐aЗf�V��f����'Pi����|�E�U�NXA��ٙ�Ұ���D]�2�cu]��"Wd�YȀ/{��6Y��il��:��j�l'{nW��7��b����ǷHZ����Ýj\��[���c�;��`4����}h�<%���åi��R��N�m�%�)��	/	VB��6�U������!�E+8�I�X
�G=��p �L'�1s��O2*]�����Q���D���v�A ���Wmt�����H#����!һ���Mz�Z^��q��U?��;+͚�#�z;=�\e1X�X��w�B'��|=��ݾ��:0;��<t���v3Ў��a#|eh�H��kz����8��Ю�UP�����:��´C���	!��ʑ��G��R�M|���Ø�9��gg9 .S+���J*�6�>

��{G�)ƕ�{Y��7�/_0��/��2P��@,�Y���V0n��@G=L�6�z.06�̫��V��5v_�V��{��i�i�U���I���V��
8}O�يP��$���x�ro6�hFW��dɾzi�N�cw�gP�*ae(o�>�k�N8�jD�fxk�Nm{����j0�S�[ }l:=�.w�4
��$�F��H�Ű�U�Viݪ�l��|�(�P�Aj��p�D俁��=���A7��L{"�y�|8h�VM�I��~R{t��@����2%���ܘ���=����O�U �MA���YK�����y%��8��%�x:m�Մ�9]/)2���a����QG�'Z�3�*Y�����tGQ;u������_��'��G�,�]�N��j莝�Z��FP^�{�Z�#� t�F���� mJ����*:�	��V��	��*�"�%Y-�m�ӛl�H�B�cs��H'����\_��c�	��2JRS���b"���	U1��\3�@Vc�*�xt�j{M`!n">���>�7/�|�	��S���&Gͥ��J���ZK�Vpy��E��ST�v"o&�$�3N�!&��/Mvƽ;��U�𵴺/�@��V��� ��2�^$�a�����@�A�1�}�iW��3uD�N�y���"7�����:�&�C�7��pH���Anq|'�����	�fC�_Y����s�8S��X�Z��UJ�W�r����"��Rc4H�Y�tm�����&G��N�����_�/�pԋ�ɩqԩ�S���=����HT���⚱;��I9G�"�G�Q��4�L>�&�@%P��V7MUf�\{9|���n5�?�$�8{�����6�2�`Bü��g#��U�4����K�VD�#wʄ� ��Omfüƈ��:F����".$s���B�1�������@Ԋ�PQ؎�A-���g�sD������ڒg�HXw��֊V�4y=�W���6b��Rl��\�c��'wTK��� "�zW8���n�y����y$�|$�QZ�̸I՛?�\2)���Tr�Kf��G�kRKt��&/~��_K�w��3F�5]r|��@� (���-�#W�3��J1
�O�"ڲ���wA�S��Y�����}�?c��J\��_o��/V��~�6ۮ>���1��y�^N��e�.�&���=m]*zZo�i#$.����Z�w�{�`�Ԛ[IEa�1(��� A���-�q6(��]��spb�]���&��g���T@��}�l��Y��9���a|@?��/-�u��Zv����� �|n]>?k��~W�e2�k:�,Q�G�N���z��BځO�)[n ��n�c���RH�J��5����(�S�v�NnhL�03ܢ%ȿ�= )���ӯ'^4�/��a��=*�"lc�?�*�{�3X��VUT��l@�AӢܭ�;6 �1,VbD�?B��0�+����WI�O�Xm�ϱ������]ފ~�4��Ѹ�=W{O�A�ua�F}此k�XPp1���;�QCHLH�9�[�>M�ێ"\��3�iK��u(���L�S������o�\ޠ�����'��L���S���a0�B����vk��K�W��,"�D[���/�MӺ�WM7��T��O�|x�����6�v��>���a�@}��!���91>��d�ߑG�h{@�<���Ln�n�k�Q����N���&�gu�(M�ϧ|�qOZ�"뢷�	s���%�AY?͐�X�`�Ɛ��8w����Q'U���uM�c7+�|�ڝu����4�YTr�����^��TV���v�S����2��Gߗ�&�AN�u6V��g������~"�2�1}�=��])�	3~G�ݧ�Y��t	��x����y7��v� żaZ!��!�k�I\$���"|�U���t��@2U�^��b��H&��Zt�I9��=�.�c���K1t%�Ѫ�u�tK�7��S��7�����XT�Ea�]2�n|VZIg�u��	�UAѽs��4��ڌd�&��I��Dm2�"��[�O�R_K6~�e*�a&�9�﮸��~S[��Z-���N������1�/z�o0�����V��$��E~���<k�RL�!N ����ÕS� b�V%�v+@���B9A���062�lO�
y:��������Fx ~sX%͚�Z!���:hgZG�1V�KV̓��;���������0Lzw6��;�Ѹ���5�4S|<��s�n�"#��Gr�)c�����eJ1,1c��9�1sT�m�M��FL]��
��=���7�C�}1�}P:+IT����o��p����Fi�y�
#r�1֐[R�8�#�=�ю
.}�Ӥ{ɶ\Op(�-)�f&`s�]ٔ�D3�T����̨2zv�OR��Ϋ�,Œ��^�O��3<�?��ϥZʅt)�*b9����\�+O9֟w��c=��hb���NP2Ajp�;��<m���,�䚿.�t�6p
���GqL��$�z�����)0��6v �/�K5,�ӭ��z�U�ZG
d�.C5�;$L	���i'T$�Hn>GB|�d�T�AV�G_��т���M�H3��g�:��9CG�x�`D[��M6��O<W����l����`v��G�՗���t`N`��Ӿy�@j�JӼ�˕P�M�<=<MB�H%�3M�OP�d	]U+�!��uU�\?��:p>��p`���-x��RC �)���fo��J��1ds�딍ߝ�'����w##�[S3�ɥFV �����i�iƬ��Y	uT��;w��v�z�
�Og׾^��.��l��j�A/,wNk�V������73g�k�����V�Ù�r&��^�W1��8r�յ�z2\<M���2Âjݨ���@��y�L�\���Q�}t������5�����d>Pl(��R+Ӎ����z�������e%c�F�-��gs��<�����?N&�΅uEv�������m�����t��������2*��|�f�	��G�M�7���]���hΫ�'�W�43W�ʠ�)�u*�򀇓��Ë���T�:2��r�E>Y�>̞Y)�6K����;��!�)%��Uk�[���l�G��Yb"�\�z����f
��e�8W�L��c¬� !a�{��p�WM]�Nx��?h&��"��K��)U^c<��	��_	�c�҆O��wF�.v�w����&ۅUu��&�2��(�5zP&��J�{04�ƩH�H�����ms=>�c�uT�ƛ�0\?�Ǌ�d�&�/��+�)r a���Dڗ��j�;,��[0��n�8h�5(�&�5��,���]^��Q���`Us�>m U�N�.�j X	���EEE��g�lb��>m���~"��\Ś�ӴF�:{�D8y��Y��0*�vD[0~\<Y�f��Rq���:�7؄��t�5�+���p�Ch�z���1���H�h/�n
�#R�����mk�
��}���KbC���$�i"��ڼ�	��K��K&�'vu$��-t�I �R��!�-��ϙ܏��yփMǈ9�{U|�����2@ԕ��0�q����Rʢ��kK��db��LVz�~C)����O%�?�H��Ѧ�q�����A̍-�[C�ר_U%�Ab�}��}��^R4�O�CJ�տ�����1=4o6��{2�V�mʡ���RUY
p��ׇ/�u�SX���R?湘�mS&������Dvt9b�$��`\+R��y����8�"�O��8�u�3gs���8(�C�${h3B���^��	p�e1DR�uY��hמ��|5��[m/�4��\�0G�M.��ST�0��Il�R"Ҙ��Z��5�����Om��\7br�֍�����K�Qw���2���`O���Y�RG6.q�D=LB$���1D7��A� �f�3�W��Ms6�o 㫗���B���.�9���k�0T[�����q�bP�$Aʆ_�}�� 
SZ��;�;�O�7�ZT8��D9@�]�H^��!�b��m���@�D�䈥��O&{J�8�c�8K�墲��Ȉ�d4��D��K+o�71R���_�L�?�^�ܳ��$]-+&o�!n�״e'�.@�1�t�ϟ�T�M�4p-}O��l��ʎ&����)�N��	aN���a��
7,Xr�6�y����]#j���X "�d����^�g���vr��(D��u��y�=h�w��u#�A�G�|w"*('��P,���
����Ja7���_�f� E9�xxOڣ5J����P-�O��?!TFHv��궉�,���K�*���=��T�s��lA��=4[ر�=菵�m���Y��(��"De�*ip�Zji������:���H�2�)��4�	�F��w_�*�;��I��2�{C�@#K�����Ȉ�#�X�x;�i��D�{�0����{x�\��l_�: nr�^�b�~�:�ïy�W갊�͒V�UW�Z���-�a��v�1S�n�����d!���{F9#����"�m{XL�V����K���*Ffz���P�8�])���X��3�.�O�����GӇ��vm�v a*l_^;��le��b�� ��\k.A�z�F;1BMg����Ƙ�@���/ ���^��b��N��y�>;w�	�O���>��<��d]� ��7j���E��C�G}�����u��*���T�#��l�N�@t0��-�Z�x���Q�A�g��{B�ф�qG�i�� ȋ�R�u�WI�i�)��d�F6,�s1E/r�Ւ~�| ���7������F��8n�"G��BJ�KRuÓ�З܂{�	ТJe8,�m�^�c����d4^�
;I�8Jڜ��kb���8������Q�SG�]_i=��,�x!��y}��<���35���$���`��S_5�D�4��g[j�U��R��f����q��U����
�ڎ��[��{����;uMH�S�e*�c��?��v[�=��t��$�.�~��=�'{�*L�h{g#գ��gA*�"3aU��Qt"�&T����s]3�Tf=�`+�1w���8��F�oS��V�ަ�gbXڋ�Uv�3���I��7tt�tg\��4�,f�b�M��	����Z�5{�U7�_M�цǍd�&���o�?�鵀f����ծqg����� �6�� �8 �_�,AGz�ܧ0�1�=ǻKh�.��֊6�}��S����j[α	ļ��oD���-�v�H���(༜C�xS;j���#�]��!)�s�/��}݊ � ��������$��'���=D�do���\��c!�H�'~�3gZv:�\O[�%4Q�H�a�0>^�i�F$I5��n�'�}�S�kmQ4.�|G9�@��r)� �3PFĴ��:f3�S��l!�~�����9d���vm����:��ܪc:�#�Gb�������D 6ɜ#_��6�C��I:1������i��U0�,�@{]r�f�Bh�ʭi���יb���Ɨi ������z�a�a�N��8��&,^n�m�9� �vY���Fi��.8��������)1�~j���dG��k���JΡ���?YK��xѧ9xG�M�|�����?�녈k�U�1�]�D������Ͼ������ <�ס�ט����p��O��?�2y��̯��b��.;���"=&�N�Tw2BZ��ޗ$,T��+��[;�]u��h�Sj�����Ogfak�O��uM��G%k��]^,|SCZ:~Y�;��s����##�i-0;A&C@������{�����.iu_�M�_nWܯ�e��ϴq=���_@h�Yn��Al�n�j�b��җ�p��ɜ�B��Jt=`N������z��_����Dz�u:�@�%�"4�@Z������ �}6Lw����Nz����W<~_�'���~�d5�3Sb�O�'&�t]l;�E~ub}o}��o�U�x�5Wfd>�;���4��*�5ќ�t�D��M��.7)�-�,�����8��u��b7�b1�z����QL��8�JNP��!B-p���ԝÐ��\�Ҍj�A��4YD�M��?u��[v�� �.�2憳GYb���['H
���}��5E�ب�Lsbm��r{=]��vq��,��-wñ�������	B��Hը�%��O��.�*�n�����.&a���+�NX2��YF�)������T��~��]Ն��f�KP�Y	O�Ā �C�9�U�`Tq�����tP��կ
ZW4k�;w��,~�`������{`H�y���?�q�6�l�ݴ�����>�Q�'�gٽ�~@�pL�MQƞ���K+_v�������Z�IvXH��*tPl!	�����{B7��X���=�R>W/+/�D�#?}9���{x���A4"�l+��+�P�(��=zwC�5s8�$ar�kf-sh��/X��T�H�KxC@;�y�$yES�up��j����?P]�"Izd�ܦGf��Yk�S*���Ĭ�B/���
	bv(�(�_u��Sl�O���E"���i��*~d!����G��S�I`n�#��هLYR�ϊ�a���������FÚ0\�2;����	NH��k��P���P<���x��m��HbLx��y{6�ʄ��
1������P"�7��Ξ42�,���}�������G��ӷ%�����qE2>��	��&I���
*�����ڴ�����U����<ѳ��Ꮈ,�lﳥu*�^um��{(��z
�<�{��ϻ�I�)��[2�Q������4�8٠���S��h���^0xOu������ee��	�`j4떎�^h�]��-�陽��\(Umo����_u�Ę��0�4�ck�2u���{y,���j��@U��Y�Y��
j�+z��`Ic3��UZW9����H7������R�L��X�pT���O��W�qNۘ���k�����Q��i�`�v�l�+���z�>�Q�cIAN$��vY �:���=�Ik�[�l��~i��e�����D��L�����Y�	�c�E\������ͤ"i�Vb(.�* TQ��ԤI�˕0?�%B�")y�l&`�������zՃ.mT��l��C�fX�����N�MF�/��G�� �� �����}�yy?��4bα��jzbJ�m�/���퉿=x��kKD�0c7�
]6��
^Z�R��|8�0�������gݪK�X��Ň��Ʃ���w�pf����}�������4��1�ebwE� ȋ�m�f��D��g �����-)~��*�P�3��ۤ���vg���|,ޓ~���߭yx\�4�g
K�b�}:xh�G�)����O��-J	�R�|�n˼"�9,�%A�B�����+Td��-�c����}���P8I![�$��ST�Mݔ��\w��P��;������K'-�тs�Jf�                                                                                               �ܪE    b"          6� 2� 0�   :� �  input Ġ Ԡ � ��       �    $�     @�     ������ @� T�     ����� T� \�     ����� \�                     kernel32.dll      LoadLibraryA    GetProcAddress      VirtualAlloc    VirtualFree   WS2_32.dll  ADVAPI32.dll      SetSecurityDescriptorDacl  2�]�ҡ�� ��2km��ձ���#����7Ri,A�H�0�
U��r�u4<E9H�3�BS�XV���g��W��@�E�8ȸt�X�NO�U�x���`6��]��u��}c�&��tY�eq���M7j*P���Z�}� ����AoJd�u�M��?�����]��f� U�#����=@��<�sf(��͂0���]�F�E�x���N����9u�<��8ƾT�+c�0��7�hu�
}�#� jY*MԠ���ݖ���
�B�ip�h\� ����T�M=6��@>�+(�c�1,��e{�u����gn�"ؤ�]u�����u	xs��3�ب҅��1X���a)H+ƋGv�0��؉�Ttg���x�s��Sa�dz��$ub6��s�����n
�i!g|�����I$ݹ�y|	|e�=��2�
m��t	�Qk`�����ɜ�-Ǵ�������$In�#
DCy��j�N���$�2�}H���E�S���ȓ��Q�ۤb�
l^���0_'V�ЈË��9U�V�Wy�����աB�&�(1��H�s��6���X�Ubs=D^*ºV�/u)3����Hq���L	�jM����������im)��+�:g�]���i&A�Jx!`�L��@n2�z�Js#���D��2�UI��ub��k�vtQYSI����F�������U����U��D%)�.
�1m3�1D���2;��D�b�`
Qaq&�q�%�k(�eb��bh���2A/17_Ҏj]���"��?�ܘ���<�C@��4����;|b�.���6F�H\��:���R�	+����,j�z�eg��mF��rjxY�����9�>���y�#�$��С.���i��h$� �u���s@H�p������?�����,`��}����a@p��
��C��~;���9�qr)�
��uЍ���B
���"�gG�2}�O���M��ڹ����h�B��Jf���n	�|?�R }�C��&t2���Hp�+�μ2��ÒAK����7u�M;������E_^� ��[����cV(�� FW�j	Y�u�<_|phKF�����p}}��9��X�d
����� �Pj��QW� ����Q����p��VQ����܄r��QFVON�A�WAP�Gm�Q`
@�8D���Ll].�)��)4A��$�#>��#	 Y���00b�yM$���l穣2J��­���<���fג���8܅!SWVĝ ]���T�����F���;+�y{�XV�v���!�2��@��{H&tsD����#ӃG�{@Q��ߞXDr/4o�Z�x	Q�:%�0�N,��Kj@�ʒQF{�)!��V��%r���6���(2�GM4����I��C�:9`nt{��*W�6�[DTu�E��-0��W�tR����Q�3�1P1@�W�&�����A�R�?�TЖ1j��D3�S@1���7�"%uC�QK@p�����7��F�%R��W�5j�E��&�v-�F�]^_[�b��N��[��A?��	�Q���D�\VW(~�r�X�BvtR�~��P!֓%�E�Z���L��a�uś���HZ��G3�G;�_;�tY�w8H�Ry��+�������dV�?W�	�O%�f�\�C?��ņ����h�������O�����:�uXRvI|���vRs�f���[��#8)��!���<T	CQ<��0J<&t
�D��.P�����F��u}�Z�y$v*x�l�
��6��;�}4prF���U�,���t�����u*:v�I9�����!����sA��^Y��Ft75;*U0���L����;5Q�7\�f�vR�� ��bY�I�1W5�Z�F��U?}MN���C�Xl�tM�Ls1}(Kd��������"�{���{RP���ʄ%�Z�f;2�=2���
u���#��(��,	0�QRHV�ܤ�d�T�)���}�nAH+��6J��^� �|KR�f�H,�RI�WK!��!��Q�v�X�@td��Fu)g6������Z�Ð�;}�u
���<�@��b0M-ss�}+ԜI�^��N�E�@�-�-@��N��)�haI�&9\(��t$�DC�QN�h�~3��!{�PWQS���HF���@��N�p�msvrb�2��tE�K�[��![�F"���X@��9�҃OӑK����N��BNc$�w��JA�U����������n��>~¸tDR��8�	%�j��Z�A��fσQ@��G"iZh�loM����R,��묝#�V��D�Uo{\�*0+����;MHf
A��6�ak�'mK*�^�@< �H�|��'����`s�2Q�vP�@%�8	B����,���Y���M�#e	2�8xC"�TR%%��]cAp�lic:aton er�n|)�� �u��.The��<vcd�%s5�l��n�t�b_va6�i�d�SDL�BG5f�d,7al z3W�*bN�n��|us�32M�y=ag�BoxAw��1xtf��[�	�"[DGS�Agkpn6lwExitP&���C���Ha<nd~�Ozp�XG�tzM��lM��Virt��A�c�����	���+Ҧ�q'$�I�	RI�w� `�t$$�|$(���3ۤ��m   s�3��d   s3��[   s#�A��O   �s�u?����M   +�u�B   �(���tM���H����,   = }  s
��s��wAA��ųV��+��^��u�F��3�A�����������r��+|$(�|$a� d� �  L	  }� H� L�    @� D� �� ��Y �A�T$�R���+ʉJ�3�øxV4d�    ��USQWVR�� �SR��j@h   �sj �Kʋ��Z��PR�3�C �K �C�K�KʍCPWV��ZXC��R���F���+��V�K�N�׉�� ���KZ��h �  j W���Z^_Y[]��                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                 `     �0   �    @=M=                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                        