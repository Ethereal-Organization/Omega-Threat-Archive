MZ�       ��  �       @                                   �   � �	�!�L�!This program cannot be run in DOS mode.
$       ���si��si��si�ld��si�Rich�si�                        PE  L I��F        �   �  �     �     �   @                    �*    '�                               � <    � 4�                                                                                                                  �     �                 @  �.rsrc   4�  �  �                 @  �.idata      �     �             @  �Themida  @%  �  `  � .DLL        @  �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                �D.w�h;'X��k&��Ti b)IgI�^�I\W#��3g_7�W3'+� VZ d3���{�u�0LO�7��˄ӗcX'��7#����_ü�3G&3�[UZ�dǬ���Ǆ���c��[XG�ܫz��8x�O�PI_��K3�&w�_ [&���E�IG]�a?�z�� ,���'��YT�_�FӮ�M�f��K=�i��nG{E��4k]Y]#�� W@+V�Tk{k�7I�0w�������d K�K�����(��Ϣ_՟�K�_�_�R5W���Y)�ðm6x�Ub�M8���@&"_�1��[����د�+xK�e�`��5,�y�<�/��}ldL 8�\���B�,�1K�={c��7I�?1U�4A@ DLN��C��c���	B��j.?����+UFלx!ڟ@�/P
/�)?�]��^b��7��Xb���ID0C�Ek��M�+#���;��+��u��_8�Zg�Q�T����h�� ��X�g@k��}h(�LOt�� �%K�I�T'�߷�S�O)�	D�6a ǏI,�NxSsO��k��}��G
'���g���#�/xB'QC3ҷ<��H�T7q��;s�[X���
�Å��Orvx�v�{�� @@�OS����E��O�f�;GSW��dw�%oh���S��@s��<��}��oh����#\��p`ۺO��gOЙ���yL��߆/�9�Y݈����w�x�PSƏ�~P�7`$O�t����mO#��/)�c��s�2c#nZ�H�M�)P<'�r���+,P�]K�N����0���y/Zۇ��07�d�Oc�4��}ӊ6�ۛ���7dSO{�Z�i^0���,/���XGh�՟ [V���[ا[��,�'0�8<'�i��#h\�A���E�!�/$@(�K��у�P�߲��	���K���gk���X��s��{PȘĽ�����d� �̢s��X�B�ݻؕ~t�϶c5T' �n�4�+�+��E���,�Ad<,O�6�@�ܨ�f�4����?Ǌ]���݋wo
���b'X�K"�n�V>]�%kPƼZ�'��
�Bu�8��AIw�	\���S��z�'vj�[{5$tnK�b�n��j#Q�t�����n�(�B���^�<�AW�қ�F`*u��G���G�o�8��tM�x�XUw�M��A[sYLy,	�g�8�ܦ�"��R��"n"�@2E���~�Z��L'�/�� �P=��%W�P���P]3��Ãѧ�[�ħ���Tc��W?I��8T17���=��� ��cX��@i;4�uW���d\���	g��{�`iO���ñL�h����kĨv�w� �L�~�F�+E�0�Z�Tt���g]>��|C ��~P�G�\�@ '�J <�a��͐$#Xu����;d�-<��1>�r���I�E�LW�O�W^O"^oO߇$�]�z#���#l����~�^�O7(�+�;�y��s�F�BY�߃�#���$ly9]	(xt7�p�Rb\"L�WE��^���=�_�x�L�?,�0x;@r�E�5"�w�/HEw�64$#�b�L�wO�4��÷�d�;�cӻlG���/LW�_�Hd�K ���O'�طdW�g̋(P���'T{H��W�w� �d��E��`�8(�����8���wE�K�e��'��C��@��� �l�!kOw� �h�m���g��㍵̰�N��EjG��o�3��}[8�0���k�otg��X�?,[C�;E���G��[��W�ۃKOt�(f	��&.���D��L�cx4�oY5m(ʷ2�h�A! �Q5 �g��:�8|.��i�
O+5�5���P+ �X�,�C������[8e{WY];@��"Hd/_�O�v�';W�,��,	40!g�-,c����x��˒/ɍ8#4��o?۴��%7���D[�`���[@37}A_>�K��4��������W�Sde�S�K;6~�T_�-I�k��H5��R#��%�^� jI�A/7駸��VX׫G���K�L���#�OW/Q߰L�5�gVH�� E��������⸳�(�e��&d� �e�:�]F���n8�N��Uv;�����e��� \c{qfV�|�+8�XJW$!W�����O�.���sK���N��q$�W�g���Y $���c?a���I�;��"[`�Wg�HmS�ۊ7�0g���t/4��Ww��D�Ut�=ӝ)@ǲ��_J�lgS5;�n-���o�n��̯�-�P��dw((��`���J�d'�JI��	u�Y�mCh�5G`��SC�%��CvF�I������?�����ouO(�1+{�X|Y\x� wy�C�Ls0����Z��i5�H��p�e�h�1����[��7�D=:���s(*56�e�d�t��*�opOd�Cy3SW���� 8�x>�.�;_,h׋Ks+_wj	�?"K�(cv�׀��Hk�4Hoh�VK�l��[.4�%9��/���#D���hl�7WY3H������ ��J{KvfL�^p|'k�{i�ܧy\�@�ڵ
��#���?��������0���p��' ��7	��0hԏ�;��Lg\�hk��i���1�\�c�}'o�@�OA�sW�\3(V�H�����F��쏛+�pnp������dg�j�59=�E @�#oZ��[(��X�����xX��C��Ӽ��=����Þ��0p� �gcj+*�0\g}�v��H-�h����(�P3� � �gp< �EU�d 믽|� ���SQ���\���^��(���O�K��5{ �E����Tm���c�[��?�㷍T� �U�@\��u�g(x�óu�W(��{�m���/gJ��O?|���hc\�Xx�ড়ug |nu#���G�c��Z_رu;⚒L/��)i���� كg��~���σ\B�`�, �l#�S.@�e� &��'t!�XY�^��A�=u�t���K�y+0�P���pP;QW'�J�T�����L�)�'�����{Uio�I=��7�#{V����+\!6� ��#��#�&ܟ$LA?uO���OWA����'�1�ŭ`�k����6H���5���q��F� �'H �����`��Oo'4�+}H�t��H����Lr�W}��c��V��I@[�xo}�[�{�%���*o棘�ק9�;p	gFL�+�Q�6�SK�o�;(�k�G�;�.�WY�/��헍�0{!���˔^��&�^*�W��3��Ζ��4��y�9l'$G.�6��;�L�k"�7�[�Fd�HZ���3~7Z�0�Wl��E�M���4'f3`T����?�q���u,kiy��-�+6S�lI9t��{�T��ȥCP_�]�fw�,"a�x��x���k���(��n�|/�۔�#O��[^�f'� ��V�7��`K�+�y�|;3 ����Tc� %��$7s�;��_�㖥OP(_�]�fo�`��ᑳ�t#3 ��ӑT;�,%��%��c���(��W��O@c�E�9��igK�3��f:\�����1�/7A�[O�;��˃�d��O��[^�f��Փ�f�G��`[�S_x��烂��(��W��g@�[c�;��'|�[�P��O��[^�f����V�'��`;�Xy�|3����{T#�%��%��O�fÜϗ_�T��x�CP(_�]wfs�X ��� ��]^T��|Ǿ�?Px���:�򫅏�#o����]:ܼ෼��+eH/��3G�x2��ˏ���AS,/E�;��{�c��h�GP_�]gfO�(��V�c�e��gW�dP�,{����s:`���$��%��3�f����?�#<H�_�;S��_Ⲩ��V�[?��`��g��\tS3 ���[Tg�H'܈��瓂�(�W�؛A,4�;��?|'3ې�O�[^�f�Ĥ��fo�T��wW�SH�{�t�f�r��;�#*H�_�;)(��᧧�q�W�[}�/G��s��9�CVz��j��y�TEM�F�L�T��{EGLYޟ�&tJ*�۬c�������(�����bM 4�;���c�� d�W9����}'��� ,�9T�G�}���#�K�pƙ_��j��{��$ho�Z�4_%��DT/���`���l�W+��_p�h˔5.oY��?��_�|T]T���w�YׅL�9ć��}3�Ąt�( �7L[H�X����<3X'�T�4��T���T� ��3�<>�(�rg2+���U����\�5�V�-%��|��EG c�Ly��UOw0\����X���<7X#�T�}��w������[\F~X�؃@����|�(x�8��80�r�)H_F���vcLr�>�D�������|Lׇ7Q��I� 8k�Wct߸L����cL'[\�X�)��X����d��W}o5�U�x��� ��L����üu���"�B_�SE���;���i V;	�gE_�����l��Vj�1�KF�V�_�7��w�j���%)��� �u]��H<U�&#�PC�ìU�Ȧ?��$��RH[�jsڤd��4��W논�H�l;����'㏤&PA�5s;�BU���\{��j(@�5dӢ5;�������_m/	\y$T3p�6c��؏ F@%�A<�b8�;�j��W@�e�'�_�����?5�9��:�G@�C�^,��%���#��Ⱦd9��-�	8g���72���!�G}}��Up��&�O�'h3.�o�?�LŢc�Ms�M�5Mde�$��Z~?��_+=Y�O�=[7�����4��	��[Od��^G
Jm.�D�'$.0��Y�ðꇷ<f�FxmC�T�?���߾,K�B'C@�7}+gf�B~;X �L��c4N�Wg#K�Y��xw�S?-0��H���G�0_HH�':�S�Z�b�B/Q7�M@+tk��,��sX�`�7���7.=ȩ�xќ5ݝ��7 ���@'��='���ё����rT�E��#���Ķ�'�w��
|��hO � ?-W�� ��#�@#IH�#:�>,
xhf?�7���ӀvQ߻�%�-�@H�$@ �,S�=W��?�O�����_=��%/��	�'|Ѵ'�Op��Q�e$h�S���DS� �G��;�?�R�C^�K���	|W�M�[n�����J����$@8���ӣ��s���.��X�t滛�� d�˗�e�����\�/pmKZ�1�CoX��'O�&��Os��f��3��5�߸i8_}�5khns], �L�)"T\�b�{K�_�'�I� 8g��0U;H�+�\e?[p�X�����!xy�� �cl���>������#{�����+��S���%��_���hZ�{s1��Ŀ��0����xL!(Z��Sh��EO\cx\"+�u0���H�oR�'%�0���౗;� �. �;0�H#U�%+��cv_cT��X٣<�h?[ ���Xc�C<�h�]�h(�L�)�eӿ�^S���Ϸ���˔��#8��\gc�dKx�ܨ�5�ќ�	nWg��:*�HT�p�\ #�F�9�����cTH�Or����Y�'���{3����'�bX?�&O�08�2R/��Xa��[��o �5ƻZ�[�[.�)G��Gz'X� c�:�T�{6'x�(L�I�W>ε[w�c�4�xLc�-_{0�L�)�g�]�P ]'��=��(hLS��V{9��b���e����d=e(ke
�r�k3���|�ǚ5�c �Wƿ'7y�+L�@���a���/� |��W�\� U�;0��Tm��([A`9LƗ� {��������}�+�?� a9��3�eӊ��?�� ��d `�#3�Ul��軷��:X�T�'���g�z�0�L'�tUg;���������;Pt�#��Pv���9�{h�W	I{1gF��T�[�K;ҥ\���`O�cT<OJ�(pL�;x����S�>%\��Y=S�3�L��s^\`(�e� ԛUX� ?�GC��`��O��M�7w�c>�C'��;a�s*f f�싛��T���Ep��պC1;�J,T�k3ܯ+e�K�u���[��X�||W7��}l�� ܚ�{,���ߛ(�L��O���L��5"ٹ8�K���ZU.J<��8�+�j�A��g���m�'K�IL;@�3��ķ(u��l��g��d�\0�C�e�Dy+,�T3��6w��� �ԃ)�Tr�'���� ���~`�'��s�Kc�N� h�3)Hg_(��g!���KK�&�¾j�5�'T��k^�kpt�o�F���K��04H�����|ޗ'P�rY����x[�+�����@eh��7$)�`�vۃS'z*K�|<K7\����c��	W�5��K?ct�ȩ�����cne�v<^����a'��?����>�y�� s�d�g����;�G��fL�^�l�/�k�N�;@t�d��)�-\Jt?���BG�cDk�:x��я�+>�v;*]?HYc� kǠ�U��G�8{(�`�GWA�h<[7�8�Afcd3��"nc��E�B[��Z�e&S� g_?Ժ'���+FX���V}��~������8���T:h���v��B {�j��e�[�BY*�� /Z��WeF[�X����� #��Kebu���c<DkVs�?�F��8h����`Z«�lk����)x�ۇ��Y�ā%O~(�|� 0DL>Dl���M a+tn�����%�`UOBt5�Tןs�������~�OuK�k:��7Tu� ��(�G�g�M�(G)�Ӂ�;R�Y{85�_n\\��d'��W&
�O�S2�[`k�n�k�;��+���k6���6�(�_߷���@HF�g�JT�V�+�?����V#��f� W�+F�3�p��%y��'�s�M?D�{���Ud�+f�����Qdg�)�q2f�I��ס;(My�|K��Pd7_f���̃�8�G@0M+���!�l��W��x��㪸�+~t�,,$X\�ro�c R_æ̢C�����>�l�"K!#��%��FP��wQ���
iXWs ��l��؏�H��os�K�H�}s�)�fw���G97z�Gm��_dA8w�G�J��w�G hXBTT7,x�MxL�G��"�w�U�e�[��]��K31��G�[7$�=��/�s;�c��JS�����(8�Y��'t��7�f��9��Kgx��:��ׄ�38��g5��;�;��6m��/(�W��G�6���r�3�seS%0�D��޵M��9�Y�/L�[$Z9�)|�_J<d���3)`�7�htSc/v�f���p��W�D�3C�79��gX�;)hgS[�ܫߗ �ԏ=�kG]c^A�%T~�X�0�d��z`�gI��]iB��]
'�S�XD�e��}7�0ghW!%Y�8���Yzo�GPA���3��}���GW���&�K�g��I;�",�;�K� �ns²�_�'��g7�n%�0a�VGUOc��ޛC){5+������16�֨_I3t�GgE���Js
���BW9��4��F�5�&\�H4H��;�k����Ѹ>�:DS���|�jEM|Á_Օ~��-�<X�g�3j�?�L%��V�t�ǚ~ ��uT��*���e��dv� Vߚ��tSr�n5&���It��$�AC��Z�ԋ�xa�4�A�zV��}hc%�׸0��������Y$|"*qo@-o	 �[��o ���8�+"��3�{�2}W ��3I��Gk�����ϝ��a��r��9>k��&%=�f��֊mcC|avHI��/�UP�A��f9P�������+��g?k���dy^/��cJc�z��1�I�=�h���Y_�&3ޭ_��oa��� �^�+|D�60�;x��nug%�.GWyx G�#FK�}�/�895 $�� �Ѩ\W:� ��?���&�Lh�8���>Ӷ�,�����L���p#N��hE��\�UX�S�!��3�G�Z`G�|<��{8���ߟ��"��[�G�I88s)/��;�)5M�nf7�|:�c!c�HK����򜐵��"���kqG�k�����P.)8	Kd�D ѧU�[[*���O�*�������[���cŗ݈���Kc�[ 
���:��ٟ��X��8�>>�o�e�+�L0%�XX�U*a�7�g�'XJ�{�g�İ��c�����3'E�c��_���\�/7��f�v��<��g�S�b�?�X��]�6+��m8�����!�	�r���S�G�%�h87u.0p-��*FX ����?�b���K�LU�Hc?��_�_�L�g�T�9H$�sKw��ojX[�K��8{���"�W��]/7KE�7SE�P�DV��3�ռ,��4,��
o��̳/��cX}w$0�KyI_����{PcD�d���qGTi`�8"�d����(X�;3-�8�+"�ķ�~�X��l#=�k�6�O����jɗ|���7+C:��K&A�E�#7�8�)�OjY��#8��HD��4ICbK_��^GQ�PpB��#[ɼ#.�;�J�� B�5���Ф�'�BV5#LQ��Fi;d��A��oA��%�v%��8l�v0��K����WhK�߈~���pXec��f`����ml��� 4SH H75��+ �D����Oے�_�`ۼˠ�f�����k�?���mi��mH/;���wZc�_P�\'�$we��e	T�d���j�k~���u��g�
�8��y.��^�6���lg�ӂ�{����6IoWX��F͙����q�0�R[co|���T�x��Peh�7������߲b'T�ڎ|�\E+fE���Q��}�Г��Y����@�����2�ڎ�v�8�A�N�h<ա����:f�[�{�^V�ܚ]�7��>FL(������۸�H�?\l��yv����"�\x5`L�"�df�[�{_��� l�x�߼7�f�� �OY���o����<�i��6Xj�7P��z'�u5qKT�<����B&6������R��_k�Oq+�k���4�K-ȦZ[�{���OH��{g\' $�{\/|gI��Q�M�%056�Y�8�&��K7{W��X�?J�b��1R{3!D���0w[|�(w2H<]�g�G4SN\��UÔ�L����"��B�߷=K4+H��s�'���#��8�����@f_�T�73;�$$gx��\f�	_�B�(�C��<�FXs٩AъQ[�_�f5�l�O��v5s�r@��#�6���q��K�O���@��`����Y�3#�gݱ)X�7t����l�Q�#[q7b�TV�>��_|�6ۜ����"³[]u�[3������fr�'=���@�������Q����)9<_7H�]��o�.fB������o;���8#�y,�å+��g4~;��m�Ӿ��sX'8||� �p#wb[8[8y�wyg8�4�X���[�P���=w-;���#�.��<�@�R�'��K&�ך99�`H�/�+���3�?o����y�K^�O<kV!8�����z9���oK,�^�\.g��{W,_��S��O�jۿ�c�<Z-�H��CXb?�#_Wk֏�C��s�$�g]��[��gś�:`'�
u��X��{�$������{,�^�״���aQD�[�^�f7[d{�u`n?Gر���K_��C�p�6Pe�__�d�W_�à�fg��g��ںX_�_[�׶?�Q�+��[<[<y�w�yk<����_(�[T|s1#��,{*C��aO�cmR9�=���M��X��Q���[[����K�:[@K�/�����_=e� x���[H��|Awh��h�TE8kX�A�(����<�=,��B�v�̻gX#8�{Kӆ�̛ܰ׻K�7�Y,5�P�]?Y�<h�W�a�mOO�k��8�������0|@˫��Sc���Q���a�:��3<%�3{?�
U��x��� %ó,�K�c���@�빬�Kd�Ŀڴ�ka\S�j\�!yK@����kH%3g@f�	���c��cŗ�:d'�D)C��Ww_�fw,�T�9�%r�'B(�3�{�S;���G*x�Fm��7kcqm,g�_�x{Aydw�x�A���%{l��c)0����D�K�x_��[���6�W�;[.b�~	Qg�_W�ӱ3��[=��d�@#��	���xwB��pE_��G�0zP�;�:�n8��K*�YW�5�yi<Ɋ!/Z�@�{�����O��#Qh�d�ɦpǘ���oW[]�ˏ�.�JkI���k���2�a�A�rj�tP�0�H���Q��Xj<�-c⎟�=����g���ī���!�]#�c�c]u�]� cȏy'��l(i˫��Q�7iq#.a�iS�E�b�[{L�]�˿�Xb���c�Z��<���Q���I��7�^س��K���!�)9�9��h�;�fEehwlȔ��YD��lKW�d�6.�L"A��?�#,�(���/|c@���:��;8o��v�$�W>4;�$��,dF��fqW{F(0�3;�� �<�8�GI8�ZD�SɨX%�%���B�:��Ӆ�qs����CB?��/@KG�:�Wd_G�Yg��c�0a3ja�3'wr&���=��hF��(���\�=RXm+�k&�;K7�W��N�l��3���=���]���`�m��|�?+m����lb;"���_X�7�{T+	�� ~�3kG�:��sO��`%�����˧�<�w����6W����8�f�1Mx���l���E�L��Ⱥ'2�(���H��笹k��q�[�:����D���P���P�X��Q���\�g�D�傳)d�:w�#����ȳے�T�<$t7a"K�{��K s�/S�=�ai���`��Kx�£��F%^G�u�nC��c7��M\W�D��{˘�?��TQG�ιv�/2���#xTC|��@u��K<J��Q��4�c��6��m{>'�fb��-YZ&���v&[C���	J�C�c����,ɹ�����[c���G�Pf�P̌v'��E�\��[_�2!������?5�Ze,"J�Mq}h{`�D�?8~QxoS�k
���v.��+W�"��{|����LG��V�Ԥ1cq?��%c����<�������u:�>�L��_����\ �4�O[+:��D+zo�^3U�T��K�WzphWZ�F?H>Ӱ�fW}oO�WE�:9t�HF�2�UA�JG�9Om[�Z�K��G�g\|�%i��pg%���&[#e��x
yW �M��KB*����ޡ5��M3,�{	P�c��@ $p��3�xg���(���{��q/Z�S���y$��+X댡 W�[	�s��k�#t��Z����r�u��qg�,䫼ϴ|�终1���[���}�8Kӛv�;߉'HZ�Y���>���<��O���`�A����м�E~��@�SL(�>cO���n�H�y�guN'P���0�R'�̗�o�����ib��[xwPyw3x�PE���fcZ�Sх&j5?������ wK|�%���6�����v�O|�?+vȜ�.��=�G��#~������cL�@Q��H\�B���4��L_��#�����3P��{�/o�-�Į��[���S?�$��\�ph�8p4�"�_��BW��C�ׇWO��v@T0|+���4�[��_��Oez���\-#���%�%��8��Hw%�^���}�;3����ۛ�&�@%g�=z��L�|c<�\'�%�U9M���/x,�'�u�(���
��KA�}�ym/��<T�|��f���t VzO�8�{T[	H�j�2-@t����ei#�ϸ�u+|��c\#]'�%�U:L`����5�: ��9%�3!{Ud!܋3^{"ó =�ӓfօŻ�+���0OV(�5�p����qW,?�p�Ɉ;|�+Do�d�n�Mb3��Ww;|�-;U��<S�����'<�Y�҉l�hs]�G��K#|�B���c�H�;\D�����kXw7S{Nӟ+Guc��S|v�<��c|�U_��o[;��c8���Ϛo��E�GkY�<�'T����됇f����}D����SX+X���i���Tc��}[��.�ݗ`s�����^�ܦ?����&�KK7�l�݁/��/ü��cD�\'�$��4 ���1_~tc1ߓwpZ^)Dg@�E�-��8���ʙ�NG#�f�Z��Ӣ��X�5�8S�$h��v[�_2ܷ���g���Y�D��%۸��'<�vW�]��ó��u��(�W��'�-�
�L�bC��u[:+Xf�ޥd�߉��d�۔����6��������7d�F>��ڙD�t�XV/Z�d��$Mg�ǥS\`�a�XS
Wx�\y w+|��!*K�i�g��(XI8[Z�c�j��x���wC|ʊ<����@�����O]+$��Od�̘=q\��P�0 �+�:W[g�K*��:A�J���-i�q77��_8���ު׷�\6�g�[]H�+��d4LhH�}]�3w\�V(`5�I����{J�`�����X���"�Hf;[h|�U>Z�S �ڞ`�?6K,��/�g�Zt�ߧls�K�{�'��S�-�&F�- ���#{Ρ[z7�8K�D܇#�T�O�/�]�Q���W�Ǡ#8�k�ǣ,clH�K�d?u� Q�c?V0k`�(�G��8i�\������<TK߄h%ϳ.\��!d��_�Y����3��߻�]���d��'HWa�:�W�dsa�w���T���_{�c����_~�K{����1��ǩ1����P�]��7L!~@׭a^J�O�z<5^7�#�v��Jt���{���_�H�U�R`A��8fO���3;ϗ+N�̘@��S��́-�<�DSc/�������j�%�Dߤ6�51�(0H<K|&S��pOT���X[�_�_��2���c��{��K7kY}c���G���(�������C�,wW|�M*C�CI-]X'L+z]��Qh���`�|G>G�d��[�S��,�d'��?�T�L_�W��+�D�8q��G�Pw{|��$��k���߅�q����㷂���[jh�W�dcf�_}�(<�뗁SW�Ggݜ_��h2l$[��[K7�W��R*�@��_7a����>��H�N:�/��8��x��>�E�RDQ5�@���&?�O{'Έ@0JJ��d��@EW�������i�0I3�a\9Xa�����[�Z�+���/_Ȳ�d�����o@�^)��Gw��`g��0��'���=w`e�u(� �x�W�LA�OJ~��Հ��#0��[�SDK~��c�^��!;�Ӡ� I �U[O5c%G�lDc�l���#LS�#PS�#T��#V��A ��� ��� �{ �z/O?�O�;P$�$�E_�kǁ�;�9�����dh���d�i�M{(12e�~珐fV�� *�C;�3jG��V���1#����� �<!av��t�On�\�8�img�L�j@����,�^�:���N�̀��O�@���#��2�⮡{��,ͿcX'8|NӳʣC�A��oSK��3_���c�U�`g�43V�6���-�ST����{����eg R_o���(���0SV'��"���@[r�������+�v�OP_V ,�Kb�)�{?{T;�g�Y��?�)���}�:oWKe��v����І4GE.{�84ܵk�w��r@5]s�[���e<d�H����}h�c ���h_D]�o��K"�r}�{5`�>�Y[��,O�g@��G4:P�3P���O�jwJ~���b`��(N���Ի� zڠn�``hk��N�� ���K�5I��~E����8c��0�P/%�?G��u&ص���(��� �}�B���9���LKn?����]|��5�G�'Ohd8|Yuׇ�_B�V�ٱ��?��d�"S���1b�1�']�pd�bk��������q"�kE���'~�7i�\�`�7����/�Sp���V�d�6;ͨ���ZA�*<��yd�h_h]𓸯L(G\ytw�|��%�LaApB<��w�|+�i$��_<�FI/e7�tg1�K��wm&�D�m��{`5�[�+���s1pV^����c��K7�W��Z��4 ��KD��GrU:˓���T�%h�Y�>���a,/�H�`k���f;�/Tzd������|A� ��J�:�ԯ��_��w��8 s�OI��Z�&t�N���d��Ca� c�f�3D4�]���s�� ���gq��0G��8J���z��r#����-�l_#��_�za���eo�,��gE��蠕��iX�z�Kc��pL4��ME,v�v�l�Ʈ��+x��F�,��J8���1?�)����/�X�=�������>�c��<a�e��d7�!�ԕ�3�d	���mo<I�x|\wm���6��XX��m�o��#���#��tc�>ZG����E��'�?7&�7@+��,� �u�P����=�\�� ��M�vdY$'a�p���\�t��8a�mI�G�����؉�iK{�tz.)Zb���H�m�i�@�<wQA��?�G�H�;�Fo���z}�t? J��Z�$S�wP���x�i���rh�'yןU{=(l60u7��������h�Dp�E�K�3-��IS\�rd\$��u�Wc9$�p��#�
`��֌�7�c���k0����l�m\��}�LDU�O�m��d��,�> ��.u�;=�����`^se#e����I���}#s�)���k��M����ߏB ��B�q�8����}/eW2�:�k�����!ro|j�%�]�Ii�1�g�@>���?e*ΔW���{`��e��5�py�X�A:B�l���.��*\NB�-��!%���9�@;cfM1 c�TW�ۼ4�+����h�@%1 Z�>)0j���N�=a���>k�?U����a#3����?�|ͻKW��"x^������b�#/Ǔs;���gg�y�����ሒ�q��Fed�<}\,�|b凭D���߷1��e��Ay�!�cI�
�(��!|�o�6ĸ8�$)Ig�7��*�>��kHM�4w	 ߴ=4���T�:� �Pd1����
hB;�SD� �A�:'�DH�::̵t9�[��Qw>�eu?#�]��5���7C;��+��h8I��h[��+�6�y��A�:r�Jy{eP�%������5IZGIy�`�;[W����b�{(CSm;�5�/��0<�M\�]�Qޗ�Q}L�M��N�g{!���L�T"z��]A���X+
�5-c+f?h� ����_���h�s��?!AW�j���u�w�]�7\g�>��K��{`mm��o�����Xbk�dP-�m�ZAkɻ��y3J��po
$n�K��gi�kE�����`oG؁X]&��M|�R�9�ל]�G��G �A�|\?d�f돫+=��� ��!B��Kek�[!�O.�Uk�h*�� ��#N��H�C��[xQ��3@g�si�Y8* 8)���x�"XG���h�_THs��fS���?�˼9?5I �9���㖲4��y��HyL����g�{�,�=P�9���哗gfk�;�W��c��.�+/���ض��V��;\�G�u�CV1��;�qI��kUm���d��!ƥ4p���y�Sd�����u�~Q��&`���E D��Z&5[�!�?Gc	/�3����Н��8�3Ҏ��D �r�#�4'�@�'[y,q�{��D����G�!w+�DvQ�8d�7�(�ж*t�����<M��<���05k��F��W�v0�v�@�n����n��)c���C�OE��N�����rñ��t�17�릸d~�3�}<C���A��b%]3[����R��L�ǳ�C���7(�MK��\ Ck�����P��@��{�X�����{�����!.�8�)����GS���6>���ۇ|倶�_x_�~|�%o�Ì�͞��4�?d��`��K���K�S����1��z#l~ku��dp-Z<˷��#;G׀X���g�'c��:@�#O(���և�����<�'�T_��L*�7���\'`*8y�+d��_��w;���ČC�B��L�=3�WH��W�Ż�.��+�h/�{��@�듁SS�`�)J���ȝ@�s:|�_O��`0�4�Hc��6%�� _(��q.��8����+❇S�k��˳ic6��H�]𿸛9jԽ����ٔg��f�Z��s�l��;*|(�����]�ˏ��b�!?���9�����P��5j���`H�g8��VZ��#σ+fgh�ns�z��[c���fo����7�V	�d������������Z�An�_�]�f�[�{i���\y�G���%ש��LZC�
w�%�O"j4{,��*�{g㚳��{��xVG�pd�^a�:0��#D%�3;��)�����0<[�8l� �#NM8G��-�#WC͔������NW�v�[
����_�oY뛰�8��Wa]��~�[&��GR�8���h�Xm�ե�;k���V��߼�X[p�X���!�HS4;#�o�G%h���+7[�C�*��'���[ͫfi�ac��8��-�kr�v�mۨ�7+EUy����u�&�ز�+ 觠r)+��b6D�>j(\Pf�I ��-@��2��7���A@J#=o+�W7�c%��}��0��l�� lV��GO���`d�ga|��*�΢g�Y��bj<�<�s�_�������^�/c[y�#�W�ˏK3a�;�CMh�"�C�_B��f��unZ�P�Urc�e܈�$�eC�H`�J#}c�F�*B�x�?��)�r4d)c嗩�o�wo� o3+���.�v�4�r��乐�P�J̆sәq =���uB�"#��q6���s�:F��o�)�� tG���`��\�րd���o�oX��J��w�6;]�=���`�+�]�9�ni������g�`��Ci\�� ��,T�4��=��+X_�+�{f|1[�-J)$<g���U�+�E���������p��@Kؓ\5HoKD'��Z���4ŋ��9��`m�8r���N�g'7#%��7L�Y��Y<�t����_�-3�G�Sv��VoX9.�+��G��e�IS���f�huWJ�bA�UX9
�A��(�<�[/�ϓ9��g�݈���V.
����C��K&D��C{�	�*���2��an���\?"�t}[%��Y9H�!������2ܰ�˫*�����e���i�Dcd�ʤi+i�����a�w|l�ُ�K ��g���8{XkP������kn���i�[( �h��5\U!t����*��7j D�7V���ātO�M	$�}XGC6�d�o�Zae	���l/��#"�(,�&�ڂv�k��Q�V�aM$(�(C%YFi$e�'��т�I�.��E鈃cu�r���ӱu�����IP\'����ׂ�ؐ��*f,��8����w�/CU�c�[Y<�?D&�-�GA^�U���8��_�S8�x����!n��A>Ev�C��~����nX�+�Z�& %�;&�����Wu��l�;�b+�@ �r]<q@)@SѼ��8e%�A#'�*����|��l�K����~�KysF�cV#�)�F�.��G����G��C��n ���9{� �(����'3��H
�2�5Ku{�����\U��m�U�r�;�X�ZqNk������ft=��>n8��M��Ĝש1�KTm��i������@�Z[������#��H+?����+��q�'l�`qy�fg�����bQ��J��e�d�37�w�&���O���(��d/���_|�#;��g��q/1 
ܷ�����Y�L��a0{89�+�E���av���~�d��yȃ�QhHn�寔i��+���2�^yNo�nJ`;X_K�:eYI��R��������!�?<�@V0C�Gx�:���qYSΚ�L<�S��sqQhɔ!'�3?��Z&���q^��V�c���T��]h8�q�;ou3^Dͱ-�[\�	Q��D*�L��A�p'm)[w3r��	"z`B�Q�q�!�qe��6��bUbW�g�EY����_`�%%�b�=@?_7A�v(���Yt�&*�y,k�×v�S�^��ْA�L�+jAl�Sp/��>���:�����'Ɖ�|�3����`T�d��fg=y]^#f��-�{_���qx�����K�Uɵh�5#�~�k��%�*��J�S=+�1�_s�ug��g�q��#g\�j�՚?4�(\� �kCaﴇ1&���B�����`��K@��6�j�35=�#D�DBW)>�D���o?~�_$���B��	�>-�k8�|�l/�^��?M�Ȱz��[ii�G�[��� 2F�u}u�mN�"nܨH/[�I&��y_�G<_��EG�Fso�@��vk]?�(�%dR��&��[8�y�Hk�{���3[ѻ���'����z�t���F��a��S=��c�����>���!�( s3^��;C��Muph�_@�D�aK�n���k�����]S7{W�L�.3��qWdY�lE#��猈�9sxO}���[���~"Q�$��I��{�_P�l�'�6Co�v}�(rAm]�ЩL��\@ ��ۋ�o,e~D.ϭ������|cu��H%x��3�@+��W�֗�^�8���co(%03;�"�lY?@p�2{���xc��/�4xU��m�Agh�x@U�#�d�G3�b*͒�i5�j���8�σ��r��R`��y�{A{J#���q�#��9'���yőD,�����3(,X����:X2!?G3^y����@Tkߔx%n��9�?�7��_+aÖ��^��e��c\�Λ_���n
܊D�jW4>c]�@���},�wQu�t[�G9j(�r7[֥X�i�Ķ�RU�V�X�<���@|�I��G����ip���:KIB����`ۣZ%O˓vhk�E���gL���bESKBk�-#Ha'1�]O�GA��}a��IwvQMH� c�]�[m��7
�q�?���ڑp:X%��#���|1���4^������?����9�Ue��M�&.��1��D��� k���k�L/y�-��H�HS�S�����\j��r��G>��5�g �$'8�E̊L��J�}t���PjI��'&��J��2,�z|�왕�c(3R���ܿL�p�{WmE=P<������/@uHR���\�ChK�D����S�/rA��3���Cd� �<���=/��l�8$�y_*o;X)G�����
�&57h7U��esՉ��� ���,�w�vh�AK��"����kR���sBh�c7 �(��Id����G0�����C��Eso�KI��'{I"��"sF���W��G��w!�B��&�Y̋���:ݳD%�����\P��H`{3����<NBX�=j�~)pP�F�o]�DBG�D��i�ֹ�ӳ�$X T[����O��*�6�9 J,���T��.D5)�q|��7w6S�kU�	�a�/7Q��cÿ�{ ��TK,�l�IAG[�����J��3[T�B�Q�o!k��}o>N���n|4ٱ'��E�$�)%p%y=���%8%�Tx*��JYke"�⍎z�N4�bO19K��@4^�I�0k�5�w1��<D@��u���Z(Uٕ�N-�Wx%��|��.�Y�YE����х:��'\DWz�M��k��{���G�|����%pZZ�	���`X�N�А�k�t(�{�Ѯa�Y|VW���`4m��!b�_��5d8��8��_����i�=q8�ո��/�d�4_
GG��:�Jt�p<kaXo�5*/��:7<���޷G�J��|����'���B��;��+���{{����_�, �#�WI�n%���3�רTp�0]'-k33��3T�D�$]SJ�6��Mڣ�G�)O��]�u[HwWW�5�|L�Cl�X�a�^��9,�'���KQ�O�� +�.�� �~�q�^_3�n��i����)���3�Sb�u��)�g�c�Lâx�W_�U�W9�O�{�I_q";�^(�}K%���7:�o�o�HЗ yG7ֻk56k�d��w�$};��d`g7�`��rR9����<c�S�g@'��"d��"͋"o���{�C���e��MY�O�<��׬=�����<�[�t�Xf`7J_d�%m�4`�OP�!x��a9��8>o;m��;��k\�P��M?��$_�eD
���;�3@!5�$��8y��8��6T�*�WxVv�]��T_�Zd%󨄌�9�=������`psV�i��ģ���� �`�����'�{�9������w�x?�̏3 E���KW'�ޛ�=F}�xIk�I��
EY$�ȓJ�3<+�+aWG�ju�6��?���FdDX^����g)��)�x_@�]��_d {�s�{D@7�|��,!�ʝԖ�߹{��	�q��[���c��E *}Ls.���Y�]f�]�{�A|#����/�O�* J���"i��rw�czU�'{�Ht]���+��14?��0���#~�4jڃgq�j�e[?C�e�(�'����e�G�#��Y@u�*�O�4S�l�s⨼��Z+��GHG�,�d�NH�hޟ���Ӟ�X�hK�S�����O���'W��mo���I�}lV��0�p-5�	��|�HK�W��(��]-�U�����㨸^��q��K�`�UO!�-����'VYV�<���?w-)[�W�YKT\M�Qu+Y�l�ȇЈ0��f\ߛ�$�4�I�F[�#@AnB`�e/<=��N`���XJ���-����X'��`�B��Jۏ�h���>��3�.��g.��S�}�N���]��h"Bԋ	�wYH;�)J�/ا̳���(ȭt0S61�_���J3=GkOK3��˪j� �Z/g��_4�����Hx�%޳��L�)��
�H�(�&�	j�G)�l�O_?���7�0P'B�T��gou���+/�h^#W�b%�C0.&|E9%�n�i ��4����!�����F;���Tfpnک�U�y�k6�m�2&w�u�١G;��'W�Fh7yO�\	dQt�-F��4���-G��7��"+��`�Ȃ9��Cs�]+��w&���T�8j��nDoe����9L��#-H�'l�3� �����U��sx�ˡ�G�#�Ў�I��ղNI"��c\~Mѷ��K+���.�+Di����(ʩ݉�2��� �@�b�jږ�_ `ه�oԳeE��0�J��F)tm�;";LN�3*w��ޓ���>��R���O���@E�u.���>��ٷ��s̸�Mh{�8(!.uP��i!3���OLS�!�ޫ��PB���Q�'����]�/I[��QN5G}݆5uB\Ro�+�ރ�d�,^63j��A�N�">ͤ����]5��+	J��I���I�qf�(`�<��[9���Z?�v@�υR�J�['Iܿ��{A��m)�Z�j�s��z�˃�:̷ #gc=7M�Jo�{'�O�$�+{��;[c0�kB�p
��$@�r�P�t{�	#�[WRHE�2p`��΂��(�P��+�Hk#a_�h�6��Y�c�K��h��A{�Y
�F�T�J�j�'.�@@�g=�ZT~�7b���%�dQ@�`9Ah|�0����V+(���r���q�ͭ��ޤ|�ޕ������y 9���(�8VyȀ�7��F��l��"�7� /^�?���A-0��&@忆�eWo��c����D\��8�7-��leg�P�0����.� �O�F���+VCv�n�Hx{���#�k[LVQH��ǈ�b	�|�9�,qE8�E�mg���$@��Mc�DI��ξ���R����9` ��h2TVwK�iZ�������۳,��.K�LbgeCMd%u�=���s/�2�~O�_=�6|�!PI!�xR�3}���[�"_oPc�_�m+����(�I�)_s"�'�&ӳ5=��md�����̝@���8w�^���`W]T���'�@c4\���ۉ������;hs,�Sֈ�K�|���D. `(��9+X()�#�'�*�[�S��&�؇k��/����@��uD�&�TI7���A���j0XT!���K�fe�7N�<t��s�os�BԌI��(V���T�Xf3�M�~�>�I��{B7/�&���j$����d;�8-�,IO���6سA�_I���_ߩ�M��۬Yw��#f��H)Q�f8��	�߇ �BP�7CD��z��"r�n:�fp�����3?"/�& 5E��s�i�/��H�_-��-��7���U��-�������8s�u�_s�2�Dq(���"�󙜇߉g��DQ���/>��{�P�'+��{����֏L��M�]�h;�&K��������\ٖ�~N��o#%���N�虇��Y�����w݃�!i!�u�j�z��VYY�m�H_�����
Qg��$Oji��8�oaƂ-���(ا�W���M c(���)B�4.�����Cc�cG+ �>�Y$�l��+>y*f���5�G1�l��{S? �ClO��XRF@:D�[�L=0�r�{$�7tC2Bf����s�W+A~c���N��f"[t�xc��u�����NY��8X���m�9<��.�p���;�M-�o4"p���Sd+]8-oDyApZ(:G)Y%*ܛYң#�ir�9u7X��و��������5
�	�u];p�,8��e��9՛9<`Y�f�79�=$g��?9��ô�7�5׉{C��S�K"37�(��)W��tR�?�B��O5w�P1�[C;�X2R;<�R>-K\١�r�'mS}8�s�s���ܷ\c�PBр�gH��>{#u�S{�H)Wxd�AS��/�Om>��i����,�i�D�E����w7�$�2Yqe}(Z���b=�7E�|��$�2��|��39���S@߃���Qs�������Dڞa��I�\�nX��ru<����{�>I0h��7agD=�qk���s�{�P��6�A�q{�*���F$N[RO�X�&�\�][X���=I,$S��7�xo==/b`�a3n�4�3Ĝ�G㔳}�5��Pd�wUhBZ�/�B��Ny�]7cqW��`���7���V���TAԝ��6��u8\����0%cA`]@���'������Q�_��{P�O@8�'~UG���0��'Y�4�S"1���/_���Q��Ї�\��z��#�(�c���{��؀

s!S)�_�`�;����ߖu�7�c���:sfu>_���q�+�rB�{	hн\՛�X�� ��hgg%��x�%ZZ5(\`oZTf+ ��'yD��Pȉ�%խ��7k�u�LL-��f)_�X�R�f;M�,75��G�_�|�z����e�/oz��Ͷ�#-9D.dX�O����4�#a�̪�+�M@R�28�s-xe���I��"S\cꀗՓ�K�,�W��L9[��-�|�P���rZ�Z��@���#rW�ˇ:�0�w&KG��義 b�!��㊑�YiYR��YF(�n-��b8E���un#ڹEV�N�J$,�~��+���^���'V�@)	�v�]4N�5����"@ħ.�KD����]S8��G���IT���E[�s��9v���kGa_�(8�C�q_?�hWGwY ���u��wI�{�X�-��������w7�yC��'���Zթx�Ֆ���d,x�zH�Ctd7�?ɹ��%��{�S�Ӫ3�M�O>��OfO��c�.��KT`�^�F�f��?��JNF�Q<;[ k�6"�+�ۉ6ogRɈ�;O�LO���u�,T2�<����zHu�,�3'����C���g^�éyGh����]'YJ�P�\-�#Dx*T	��c�(`���н�YO�T��F�W���9^��ې��
��b��.���q&����L �Y�"
���!g*1��'�y���a9�Mb���}Hū�uH@/�#k�����'2_���؍�I2�-b��Y,D �A���˨{��<O�S���K3��qk���;��chG��(K�O/�N���"�E�:!%UTS!���4�4_�G�w��ه&���b �x�9�^���!��?A�KG������T��qr����#�[^�xxUW��ZZ9U���/: i��߉�뛈NPJ�L喩���(�`�y�el��)���[9�>ska�b@�p���e��a+���t������&@�.$0�@��@j\d�FW��OA{k[a[�U���������w��hؐz��ɦ��?Dٛ'4����l: ���"*hH���᪜t�@�n����Yo�*%�Z��
#�+��@KO�3_��T�Ǿ�Oݟ����Fb�	��"���G��H�7'�P2��LC��,7��|7��r�2�X=��_>�/�]���E/�a�'ڜ��g?���bCc
3rRl�e+Sv
7(��1��Wd=S��+�Ӄ%v#�o5t����Cb]�'ܜ��4)�>=s�{h�,,���`�몝��!�@�#�<*��� z���Q#��A��a+ںk8z���I�p��^����H"E��,N�/:��t�>�XC3Ѓ�/��gQ��{�Bs�T���S�H�NH�C�'�fҰ;w�F
�n7Ф���bI�t-�C��1��Hs��'@y�tH��_��T�_q�_�6µŖ��3�\��C���4cH_<?���|����Lv88t�;�le�9�WW�;�P@�_�5dܓ�pXh*��g��g+�sv����-R+�Y�C�$`2���ǫ ����f����$u�'�\T&9n8�( Ҳ�� ���Q�(Y�j��[��v�ԅ?�����)�QH����]^cF�;��;�'ט��j�c�=dֳSR�Q�}3]�ûxJ�]R�]���h9v8@f����K����l8tH!��~�t;U��C<ؽ���3qc�h���gE���
�7	@6�Xas3�f�|�J(�K�[���hw��>pga��K�߇�CS%�oIP',ƇvU��~/:����;�u�U[{�3����r��l����2|�Ƭ��.g��"XKl �Lo��;9�F��d,V�?�S�J0O;K_r?N��,��+J #4�@�y\l��F?l�\��9�S�L�(邐&�^���>�}��g�X�Ӿ&�j�F2�+'ᜧ@�lPw�v�\_O'�|�NR�μ1��#`�y,����
,��H��#XM�Si�+ ]��x�w�P�g8��a���I�LÑ����/HP���K�M�M�X�asL7k#ʖ�N.CP�"w�䖊�B��T|��I���4=Ѕ��jc�����(�#�D9H������'��j��
��������#x�ӓ�a��&PjD��bt��E���\�!��M�&�����#z$:Mq�X�39'�zB�qs�l��T]\t5w�Hܚ�U>Pg������Ct~櫨�;�gx�3�|��K�hfE��u�E��ѧ�@:{HlCydtc+���j������0��i�1�����?_?��֯��hh��I/��@#�E�3^��kp��W�}:���D��EkK�{=�����	��kox--�a���נ�Guih�݌��W�s�)AZ���Rd����=�I�ˉ'��
�t�F�B�rH�����q �@�T	lf��`]#�۵�>b:��E:���Rx���	��+��f���SR	C�ȓS�Q&`(S�|8�(���y�-I6��mJ�-(m�1�8�Mz��<Y�"�>:j�B�d�ϛ|���fJ�S2v�!	l��F��CA7�U�2�@����8�30	7�y8��|RK��Q��V�y�P쿶*�H����ө���ө�Ӊ�f}ko%����7ķ�I�E!5vܩ�S���M�[T�p���=χ�S���e�{컱��d�n���*r�����@<�`�><��7�h�b�y�"��-`�-�����FR�ܠ�&�k��N���fn?^�<%��	?Gl|[*��)"X�@��c�F����,�f5�/��9��BZ|�����&9��i�hu�>bWr�����WIqQi�70��e+%#d�'MGۊņ��(5X5h-��
+Τ��<�b�'���cG�W8!�V8'�"q?�PY '4	'�«[���G���?��o��Q~Ǭ~��6w˳�oLj`�I't�g,��ca��EH[��W�1�{�W6u����k��Cq�^�O��k[��k�&S�j�'fՃb�
m�O�4��7���~)�O��8��#.������a�!��I%_�tU��+��kx�
���}����{g�Ub��@M!>#�b\�첼�o����c�Yd��;�K�0�>|��'�H��m_:I������<���@ |�7C=W�?�q�A:w[QH"�8��B*�E��0�A���O�:u�'*����;��dC�'����L3ܰ� �\����AO bz�/g�$./g��,%��Ի\�V{|��7�Р��K�VY �9Ti�8�&����t�9)���c�|�Ps\����?wa����'a��4o�d��i|�m�q�HEr�� D-�-��7Zp��^��DJãϖ�`���X0
��z�UF�ue��$��N���O��c���hoW���'�E��:�\ I�o����\�0h^�#N�k�Ϙ�̟Н��P�[<�s1Q�U�0h9w��st�v�I_�c�㈛��KYw�GF��#qY�bΜv�"�g���޿g�8'�v��Ւ8.�?4\�qǣ+;': r>��%=���� V���E���5���I�*�8.�b'1*�}Y��< Q�3d(|@�*pI�+�Vlpm�9�I)�͂W�n}���Êh��SW���j�<��G�M���T�O��}�J@Rl� La�~����<�o���*A{��|���k%��@V[ݫ��n��P��;�� ������︉�u��U�~)��Q�Bw������lU�Ϭk���=���?ĔYj�q�O���76,K�)��ud�q�Ec:M�8^A*>����:c��v���%	c�Qر� Z��b����7�1/�HR'�\��o=koA_���5k�{��^P	0��e�������sdE�@����X��T���f�;�k�W�a�D�����y��NE�Yy��?�xZw�
�y�e�����~?M�ܢd���Jk��Ka1(�����S�҄�e"�z��=�M���3��Ņ 語����U�-�9��y}�^�>"T+ng?�?+�C��	��D'|?;�G�؋Ld���ye����,��|��B��	���/N�t!�k�H=�
Ek�0<`�H\R�+KtK/	�=Ht�"h}�pS۩�T(�Y;��Sp,�8���%�4m�j�U4�҅�gNR�tF��h���� x�.?�Z�:O9�-�v,v~r+F�S�6:E�dP�Gu@��b�k�3���u,�Q�_�.+������g+��R��6�$���ka����J���H��uk���z�W$r�I��)N�WS�
g���l�d������BިU�q�=�#u�G!\a)�KPT#x<h�_���K��3C�T���yH��-"�3%57C_f�x%����s�DS����<�7��O̜���٩�U��i��'����w:'}M
u�DD��t !GV���-�۞��Qq ;��]�SD�h�%OxV2�ݐA[��𺋏`[#�?���2�U}�������!;�]��?v�⻪�æS�[X'O�(h_	L �Y�u�T�fD0e�Qb���܇D`�u��<`0�ٰ�X+CX��R�+-��	Ź,N�Q�A�`�X�X2OW� W��-��H�L�H$��UDQ/K{���;�C!�L�`]����c�2�c�3�0��S��s�0f��<0�Y����9q}	.!I�/����;$Jx����O���������58��"��B�w{��<R;X���2��n��% SI���^sq�ˑ�)_jz�_=���+�<pܚh��f�ޗ����PXFr��6��H %82eg9\�?i��g ���A�qO�-E��_p|}G���}?kO����2K�!jAJ��F�Ň*�i�Qg3�S7�g���TF�aI��L�T߿"LC�A/�w,S��Ԭ3Gw��#�7!�l����{�]'���� B@v�KVNw0b,o	o�Y�e<�|����xY�Q[[�[�%?�Ga���ʠ�!1(�����\���]S�E�#�=A@K����c
-{3(DW[P��a[�O��m�Z���8�Md|�F|��e{�A h<|���,�d�):����;��S�p�"�;!�u�d�� C�E� p����?4�	���aq��<��6�c?��9�U��Kծ�$6,�Q!u��ca�71S$y��x�6<fR������s1���#Rh��n-c#��#�w}{ �L��d���j��l�� ȋ���o�r��-�uW���K?�Iӷt����]���_�J+�6�\�=7Us��Wq�;��5NCc���!2a-ߊ$t���c���B?L��,;�D|X'��=�g����I�a"���:�<S���Y���d��3m�3���ͳUuLaG�+�κ|�. '�H��T�?{<|7���(_x�NE5�0C_fTpIf�U�O���ǹ�S}�+;C,(_𯼒S	 W�{,KT�?O�z^�d���2{#q�W2�_��3j&�ӡ`�UW��\�K�(��(0�E\M7�^^Ʉ^��b$�Gb:��S<��K����L"�S���x���d�i߸h1n�Y�c�8h"�4hЂ ��-\�*Sp��� �as��k�M$z�?��]�7���(�������<�R���kt:',�E�Hٹ4�i kޯHʀ:b��p�XE�3zd�-���!����~^;��f�'�#�E�$�l��bw���5�H�d��O���0Xua�-#�����"�/"�R�abHP�VZ���Zr�3d��%�� �F�P_��$`A��(�N^��i_h�cg4yT�tz�3��F�28Xt���N�On�+f_��	T�h]���J�3xj��O[AoGV4K�So�ْ$)a}Ffqy�`"��m�r1!�q� ���k��n�����L?X�ȉ��j-�*.��!��؉��E%�?�}<4+��?��K�?���fY4�i�T� #��q�Bee"*3���M�&��7]�'��L7�xPX�pQ�0�>g���X�&�׿�#��.��@�ߧ6yײ��5��%'Y3�U��O�]aO�ڋk���?+�vQ���g�;X��k����K������ M�XJ�ʰ4sӂ���ͩd�U��a���uޅ��ز�������(T����ߵ���F�"����;g� ���w��vc#l�Ђk�$CH�'�<��_,�g��7��/m�+AiP�^;S̂����E�@��u�V7J�&�Ri�z�7,^�R��-�ar�6����^,�|�K<<D�����������DQ%^�۴K�3gl%SR�j�d�p8�DS�%����`q@f�V)�\��ć�I �h�_w��Y�,�/��N�7�ω�+�;��@��^�C�]����BT��G�O 4E^�����u��[����nHP9 �`�B7p��id��dK�#h5g
Q��c�:먽�������+£�|j�:��@\| N;L1��/��#��g:<O:��<���3�3���Wy{�y��ٕ͠wS�=�敼 �pxT�3����f�h���2x_o��� 6w�`��U4EY.���Յ&���ɰi7b�P�+�(3WM��������RF��{a�\l��k}wI��ի9K�YQ�y��f-�"6�G���6<�\��N�E�j�Hn`����CjF��[��Y����5�t��;mG÷��5E��`oxo��N2]�)$���� ��fkE��s'�68@NvX�%
�'���[�!&��,Z�S�"��K\�%�A��~K_0Hf�4���>�
^��|�OQcFW�˥�Z��NG�G?����w�MS�M��%cR(��b�{: ?ۜ�ljB��@;O/:��.+�MjS�>.�;�d��&M��XF>��9L�;�`�@�X�>��6��*8OSuK�}ʗ�y'@U��ڂ���2�`#��e|�F1m�'�GA�+W�TЗA{b�3�'�NG}F@�n�2 $���ql�)��[��g���
K���e��a�?�U���+A`q��cA�1>�a�����:���߅�)M�#-�Rǿ�z���2�a�/ ��F�n�CӃ�G��:$R���UW[���(�k6��l�
50ɢ��b�%��ǫ�B���U����%�&�xĦ���U!�vL��k4l�5�R��Ur����L���^'���+SA7��p�>��e3���~�g������i�qfn��v^�a,��q�5��F���RL?bݢ�7��^��A�gx�֎v��<�mu���jF?S�G�w�h"D	j�E��V�w}�G�s_R�f[ި�k�fO�Z���#�ip㧛M,ˤT�Ơ�Q+�?��K�7�.,����\�'\�
�0���&'�-A��u���c۷��r}<5w�<�ك�AZ�4�#�ܽ&h���Gdp��_��9�=���;��\��r[���V�ۨⷡQX�'i���ES,�k�EE7��:��:�.*��~S���	dH]Cs�Ը������U
���1?�Q��*��Yb\P�z�M[;:�UC@�F��EX���
I�Ϳ��s�L�3E*�Da)�����ϻC�@̀�8%��"R� �|tG?����2+���u���3 ��k�KM���+�ڎ���<D\�D-��� ��9_�~5(���cTWy�c�  ���c�狓�������� A4�|D�\���9�Qy������𵕇VOS3d�[<��+8�8��X�1K��HTE���O0WSZ0�[<�7��'8��й�"u�_%ͨ�]O3��@:���}��������[u��;�F�hk��>d,��[�3LO�n����7O [����"�e�j�O�7Mh�l�#�/�UH�X���r9=�S�-�]8�w�_ɀ���gL�#��ߔj���z�)��zO�ic�=�ԫ��hh���$�$7�Y�r�l#�����{7t��Ԧ�'� �\1Xg�+x��7�!�n������`�Az@�5mhO�kc�׸#�۝'$����?8�B*�@H[7�O�P~�	��l�[ �3�8M?�#4�_z��{)�������0���i��4\���e���bO(��iO�c', �!�\R�?LU��<��i�X�^��@�R~r�S�7�[*o̾8���铕�E�?�-�+��2	:��QՇ�H�u�d�/�����q��uy�f���C�?�p�8�!$��b}� � ��;�_����h�	�gM���k4|V�?�`Xj%UaZ��j�VWό��`�K�*hK�0��8�A�0��5K/Je���_����	�Y�����/U���}����xHq�I7����;��3@�4�	�@�v�[,_��(f����]��:��nd/����|��3^�F6�s��`��Z�����;�M�l)�X��R/:ӼfLL���V�X�F3/��6���*�1�ݍ7�|�z��ⓚw�Q���MH8���X�� @�9(�#������O�.�z��SW�D�9�d9Y�O�R2_qH�[�2)���xL�7�_U�$m��K�`������d��7���9�Mc�ۙ���+�I�EIc�"9k��������1��2az3=H�J��Er�	P#cG�*�su��8-g�k"-�� �/ry}�����R��0��`SU�;�;�Q�G0��E�@jT���
�<��Z�,���a�8�<���n �S,i�a�h,dt�XL㓱.@�C��'&��iSF]�,�;�����w[��Jۄye9kx>��b_���a9��4?dg!���@y�/ulr�5,Pp��{�ϝ�$��Z8KAQR��T���#x���r� �-��	K���	l%{�T���F#��۬[�3gQf~{?8����C�0@>�R�O?�6��؆]t3M���eo��9T� �H�D�1MCc��=��c"��c��9��K�^'��c��NR#�R(> ���1�З�Fӡb�_���O7�*�~��ϣ%�i�{����N+�{�-�=C���/�8P^s�ጶo'��w�V9��C���S�]��W���Lymԝ���% ��H�X���<�wS>F{�[��S"J��2W	J���j!���P����P+Z|@RS���$`��,�а'$.,�Cn���(q��4�-�0�#�!��-��Bu����;���ε��+5D��%N�hO0��I���od����3:b:�w�A��ƿkM�T�v�V�G��0��\�a,g)��F$z���^���x�#�;������P�/���v�$a���(��M5��g#M�&�F�a��WpÉV���I�
�eW��N�N<}��J�]o�j����[�5�WG8&��5�='��>Ͼ�*��<%�@��~6E�� �� �5ݵKy�Wp��0Ҥ�^E,Z���%���E���wM�Qi�Z��TLy��S��J�D�3ɰ�Q��J�sNK&��k��/��B�`�I��j=�e/��u�`,F2�s�h^p��(�~1a�.�8�?ȡ�,!^��c���'L��#���>ܲ��-�{�,�Kr����X�����ԡ�`К`w� kƬn�/.�&6`�2�*tw�@�n�5�L�M�{H���:�K(E�{7s�̀VZ��b��'��?���2��@bw��UgH��҉W����㸼��vN�a�Q�yE&_	��h�����}��[H{�"���>g;������}������v##}��G��2zN�jT[��Fk� @ Th���RN���V$V�u����z�G��x�N������5��Y_��JW�VO�5I�5���'�U�����/�N�e=��J�_]�� _���Ѕt�Ve�����xƉn���'C���9�ۯS�T��(��7��w�8+ �;cy�%��?T:f�WC�Rث�<���'6��0�#������72_S`7n��� �;`coJ�yV�fG�J�u���O���V�{ȾF7�v!�{�|��Wt�n$@���~!m�����SWP��~�nķ$*B|�GG@?��S� �7~���Tƀ0�Ş+@�� >(��\-������ ��y ���@��?��ƿ��w�u���.J��>�um�^�5jfj�pI*1���w�`"�!��.ʒN:������a>/� ,h�j�X�b�b�u$5|*r�+ޫ*K��)<Ȟ��`q�PW]*DDq8�B`�9�\�!C�oX�;1ָ3�Y,g�;'8�#h��D(�T�TQuN��]�"
�Wŵ����2��.=&���4;����lg���ԀRK��0�8�T�Ý�ӝu�G����˗��P���&o�?gKJ���.����ڵAE�{@�au�(�9�hB�V'�>��Ol��^Ԍ�D�6�;_K�K-��U��
�Gc��]@a�_2�@�/0�9be@��I� tr�%�뇦��D�t�O�E�r�3F(���SH����́o;�M{Kj���(��@u��7a==���\�9�+?�۹�t�����
n�/<�kƽE�X��h4�?�_�M+�����r�ϩ'�H��8��C�ɛ�O�)RR�X�a�L�x�'�Xly��� Hw�^����7u�GY�kw����-L熍���,�S~^D5�4	�
n7X��4H7�P�=#<8�w?��/�����  3ؿ}������񧄒b�ѳ熀c 333�VO;���.R��V�qU��J�^]��9WL�?x$�����I��Z���w���x 섷���!5���GN"kd��Q���w���
#����c׆!]J%Ƈ����+h���G���_�Y���ۨ虒6D��h�XZ�p|��+%/{e������RR���#P�ڛ��S�!d��w%]*Q���m�J��A�W�K"���@@�s�[�srGr���pb���Q�Q#}�
�h#rB��u�Vq}�}$���B��i;�uT��F�l�,[G�P
qFe0:��H�Ԡ�����é��������jj�V�~���,�Xޗ{>�����4�-��O��"������O��
D{�}�L+L��圸/�J�}��"!!��:������2��:E�l�Er��M[�Z$���NљX���bpzG��Vy%��ǰ�lr�j��M��]SN��_0u&U�%�x)-h��SJ����Ǆ1�\A��L�'��Cwn�&M��wc8���P\c �*,8Dm2�y'��#�?�uA٫v����?W��z�;�7=��a��z�FZ#���M{�'J�����-ɒJ�Afi��V�m\�_�D|�}/L=s���{7��g|�낢���mK#��Yg�����݂��U� �Qq��G������R�]%�eW���'�a�kC�q�sug{�ñu����;��Zs��S'��Brk��@��VL�S<Z ~���w����k��K	��@�]a�(�K�����ia��A.܎�k�@�v�mr͋�w�aG���M��[͝4��c}y�!vџP$�Z ���n�U�y��:���f\�M����S����ޥ�U8�#A��C�*��;x�'nt�l�S��
nT�S!W�z��3(X?'Otv ���L�v|��r�NI�~�qW:[ 
G%��SE�dLK
,�I�o��B�8�#�
<�zKf!c���E,�+�%��F>�r��W�9��+[�M�)�d0�gg��$������v�����[�,9`��k!ؼh�o,!@U�M!��C�ƁQ���R��ZO
[{>7�~ЇZ�`���5��c�xn@9^�68׏R��Y��Q!5_�Bz�HW>�.g[��2�>A��e�̒�t�u���>R|G�ifi9N��6�X�gPˏ?fR���D8:�M�?)�}l�<���7o�#�7},;����k�	�@Nc{�]\��!	���ͮ�A�h_����^Q��8��a��.�̐�l���I"7�X'���{ ��i�'�s��zķ�J"��X߄agD{p'n�׃�<l�����Ny�¥����h�Z�9߬�b�^W��?0jW}�L"F���;�h�c�#�/}#�q!�'2HR���{`�9Lc'���t�n4�0J�@����(�Z0��[�|S�(2�'��=OjQ�њ*���W��ἲ1�"gSD7wۃD�Hr�t����N�P<� ���=��F{sGpțV�((GT�λ��+����т�{Ӛ՛?DL;����u#s�{�+aL����������VS�5���J���}<�e9��#�LF�<G������Z�uZ�ʈ�~��;��{�3\��IMo�?�V�MK��O
�	�'�cdr(��TX�_�)8f@G]�< ��~5�}a�ׇx����� q�f����hW��{�Fi�u���e�4?(�:r�8�e�1�b�)�����-Q��?`�"x�x+8�"���#�x7xp�&EV�;��r�Io�M��V�㛈Q"��;Ow�&x�#-\��7��A/t��Ϡ�A��X���=��Y�_��=���v�ě2���:��+�YI�&�W����vgظ��ڧ%�37oa�j���>2�Q����r��k3�F�����Y%��G<���ˌ�l���IJ����$�&�n��q�B;�uܐ�1w_�|W�|7�/a�"�d(��	�s�Pd�\��A]�U$I�7#qx�[2�zP$�\9n�G��8�V��& yދ���k4��E�F����'9ȃ��}�ѫ�׋���k4��E�F��d�e��Fd�Z��G&Ø-p;� ��$��ڒ��G��� y$d�;�Z4w|�z7��w���v�׸�cm��Kj��Q���b7��_���v�נ{cU�xKR��y�5R�Ұ�}_�9��n0W׮nϸn��Jb�M���:�lJ�:�I_�q(�W�����_�s@� iU�����I�Lc;x�C�Xe#[8wX;W�D94؋���e�[��X���{<�`[w;��,YP�Re�.�	$��k���*��{���R� &k����n4�
i&`�����g����0^Ӈ���e��N��Ҵ���
kx�)eD��K(T�����J9���ߡ��e~_g�TmG�y�{�7D/LPX�'F��� ������"`�Lw��<�V�����x�Hi�w.&���.�X�x5׳�։�}X�1���S^����� �Gq�>;�"aWD@�*�II:�����#A�ᆺr�a�+����݇ؒ�<v�G�gE��y���	@jڗ�X�*=^�����OP��U:H���9�����j��g?	�����fL���B*Qi��0��Y�����7"�Es@+����;�\_G�0�m�[����~q`��G���5����i�{��̢��H���k�'aBo'QB9����o�(�U3��(|��A��E���sl�$xxcV���k�Y�6���m��#�~�I����e�c%����+��x�U�,:q׫4�wD�oK�[gTv��>d;�[�)�yx�|j\�+P���s�4�sh�ښOC`��Xg*"����Rqi]�]_�c�[�a��F(f��X�.�aןCT���<:ݟ(��?�����wh=`�;Wǆ2�
����`S���Y\u�6��@v�:��c��[�y9Gh���hЎ����D��;�@�d���f�]fӷ����WLAD������3��C��?����D�d��f��g��q�7��e� ��o6?���C����x#�2ZG�s��o��_�x�c1�.C�ۄ���BV���0G�({��P����o�5��n��j���I(H���4~�vwx��r_C)S���J�^�|�YO��h����R���I�Z�D�O�����i$e�+��8l�C�3ԅ�Wɱ�K��9������Z;�?��{0�W4OS������d������󑅾÷�<X*1�MÍ|���p�F-�^�j/���[D���c1�ݡ�sy*Et"����kǄ8}�Gj�Gaso}7�?���3V[ '��&C�L-T{�&6j���{��pp�E�0�#]t����S�O��v�6`�$��t{;)�E����?n�'��3@h����͇7�CG�S]}����_�;V�>���z�'Ԃs�HW�W�F5X�Y��0,r=�b7�������&Ϟ�i�WSe
Y�]f1]��"W��$wW�->g�-0?�A�/=����P���u��*@p4x%��,#֘�i�U�����J�a��|�k [+WEr��IvJ+z<�1��0��[L��t���0%R�'�AZ06��;د�	I�u��[����m�MEX��򔹋�B��L��&]�8>��j�
7����GZ�#_��:l
�.�X�����6P�{��|�	D�����o���O�jn/��\`��y��'�n|��-qϛ#�F��t>"�,N��!���M^})
A�0wSC�D\��	A�c:�-� E7�EM�
���v�"�?Q���fsQ_��I`�6����9���g��L'�<e[[n+(Zq���*A�o/��^�(f_ּ���_��{�roÂk�Kwp�Re���E`Yl�T��)��x>���Gcc䋠AS/�Os'vk���E�χ������M_�t�l����83��y�aP�Xઇ4Dwlo�h�A�f��d�Sۭ����&�0��S<$��N�k���:H�s�H������
$��r�k<�d{�% �r�g�ߋg��k	E|k5|��ǰ�]Y�5 K}�+f��wz�f/�� �T��9s,���1pԨ{ng� o d�SX�R�7/�i�w��"�ǝq����ˉ��EW��+\\IvY��,MhJ����p��5XD~(<h7S�0"��O8��A���52�yګ�A��(���-q�4=\`L5����?�ݟ���f����D�-�|�"6�� F�yY�ɗ_Є���L���*I�����:D� ��.��N"c�=R�f
��gНcj<��EzF7�@�U�{xX��߱�H΅�;�~���r�+EL�_0C����(p����;#O��*.-���d��h�R~p�ߣ��֞�J!k�x�M��Mڶ�艩V�$0+��.H��r��+�@P��]�񱗚#���n���B0��j:Ek�U+Y���N]=_��3�E�~@��IF���,ٸ��	�s&'��T/�l�^)���գ����D�D�3�*�$�0�[�:u(��4cL�RF�D�B7�uw��1Q���Y��k��_c���t\�'귢��c+�C!��G��!&�`�&_T!7��@��p�%3�z�1:����-f'�RK��֯u���.P U~o�����?,G��siS}'.�5{��?�>�����7��)�&�d$ �e����\�K�J�s���<e�8(�(D&P	�Ƨ^��f0�3o�2+Eb2��ɻ��ӗ�N�'��Td<�w���GDI����(Ї��O�1�W��}���(�p�<��36|E��4�2�3[�a�f�7��_��5�����#��*Z�q���$yh_;�.�KEg�8(��!{�y`_`���].[x
����=��o��.f���C'=�'%��R�w�-��_a�c�c�2ҫ��KW�R��E����[t�XG_F����!!����;�h��'#O��e������N�t����7�q�|�I+;�CO4��{�y��: ��LA#�<�w���oMj�g�Tv �_��dLÉ@�=��Eq:f��SfW�)M��s4q�n�3�dX�{�~z�o֯���mP�(P�C��Ew˅�*��#&�34�l#��N�;>^��=��d�1p����m=���KN�Ea�J��͸�K/��f��ӣ�C|���l�tٯI��'��w����DJ���rr���\�9ԗ4f������-�f���"����3��|��^v���?Z�K�`R�o�W^�!BvZF
y�����O�ȝ��p	�bN��=��g�*Fx�S�2$��,Wt,y��y��\(1\��FP�XC���Ƈײ��23�<n�� �8�wd��k����;_M�몣���C���;����/FXe�zo�H�)@�0X_���n�5;:̹ǣ����@��Nw݇^B;��CZ1y���_�U Ć&EU��_�мG�y�������I�G��u��?��D��+�<��w�gሣH�DӲ���Q�?U3��M�)Oc�G���`�_I�]��0LPD��W��R�0NPh�	�X )�����ɪ@U��v�{���W�M�(�����������t7<�[x����`S|{gwİ]]�Jz�x�+���<K����t�ą��oZ�{�5N��_Ϭ�5`��\Ww?��s4���+Wת�a�~&(we�^�n�fe����]W������U(��>ELiY��)
;&Mu��/R�㲏u�ґo)'N�Wrܟ���7c܁A���>D�:0�P�T|�:P��e���R����t�!���"O�C�ߚ�4�d��$�/S����%O/���W>(2�Q�a�q��143��/a��<O����ie!�۸ Z��y��?~=FM\��j5]��u^0�]��u�3���d%�g�R���?��u��S7��`�ȅ��G�I�k7��)P��A���p�Fa�>��Ň�S;��I*�Ev�^5�?x�X= ��p}bQ�7{ŦMt=%�T����Ji�)��z�+�W"��OM���dHH�T���%W���e+��Vn�C'�'ŀ����8^�W����WW����\L�ܐJ�8�d���B�w���ՠ�"��AIt��C�ݘ��C_�S�B��»7ߑ6�W.�{p�OUz7���DG���y@��%�#A��_��D��5$5=Z��$�E���J?���KU�U�vK�/�Ļ�{-GS@Zc^���<��<�1����1\Ӟ��H�W��U����V�Y�c�~N�n�2dZ��=T+\���Q9�1��f�ͮ#qP��
e�[�c�:0*;��;:���%M�5�M��3�5'2���(���9̉�T�Ϧ���)�2��5-bp�3F�??�1���3j_�)'{��;�㚰q�r�I[ل�\��	:`(m��y��-`��*�Y��W4K���F޴*!�}F�v��?�S+k?���@�x%	�� �IEsH�t���^�R[��[��Y���<a�L�q�i��V�����&TRL/:�s��On$;�wE��E���O�Q�E*Q>�������
�N��1�-����� 0�0��ޅ�P�����\o&	#�T%�(,r���<sY��O� ��.M[����ւ?H���3y�,�
\hDH35S(^��V���i�,B9�ZO�3X�P��
d�KF[~%V�h����{�>���t�E������V*") ;�Qd:�l2d�}�w������U�G���L�#�?���.%���
/��$⹜%��D >��H�xu�H�Y��L �ns[Ȭ)ԼX7dM�c6��-#^���i�1SW�/��<�U����%`�i����k�4�QJj�i�e�`/��F����D̪��k)�Y��e��'�@h��h�"A9Nߞ�3.
Fi�0��o��0��ؓ�!O�M�����hK	=�߻�C�WjU���a�R��s�k�<I	� N�XK� �_ӮƸ.�џ푍 �w;�r���;,�X[�*�qZs�_{�C��5��,K���RXǍ���.B%�":VUe�Y�^���/:3��Ե��r�ߛWq��z-�RA���2!k�..�e_�sKr�[��hM*�YIp�3=F�%8�s��H�l���ߵ�'p�e�O���F�cI�i��҆�G�ѥ)��5Td'�
�/^�6�`�%�jݓ���$'����^�(�{�a��.q��f�HE�f
�3X���*��TLff��
&-���d>���� ��7bZ�'P܎;<4�o�kx���A>��Ї��½�&8Pc_g��_X�&-tA7�����<4ΕC����a���8��3/'';F�3�7*�~�*XG��;ۡ(g�c��k�d���U�z�ES�͕��I��a�7�c*�L!{��b�0�G�U�����A+B��(}S��Վ�	e��_�?�YO��+�'?�Q��
���h8B�gگY��c.H#��o��R��)=s�р��%�<
�_�ȸUK�<���,+���6nS��S�.�̓D�{�{Vf=�#��R85�0�wtz;[wFAIcd��ؓ�TG9h��a���	�њK�[��ZU0g��M�(�3��!7C�#T���[?��0��f	ߎs��p{�K��;eoW�SU�N�<��F�������E�{�h����0��ڧ��`�o�$_�FN�3�����\�luό�^��
�UgH�F��U�Um�53G����_�m�IH�X�+�z���sLAm<�W��3��E�R�S>��\F��X_}�	-5�63+G=�'��]�\�(�K�"=W�O�����D�I�r��_�+���3?���GC5(nx�(9�U�_^!�#_(ϻ��3�b�]`;�u�S�������|�hf�Rqw�{U7{�r��1?@7U�_��_>Ay�w�=�!3�CFZfAe(플BX��a(Dk��r٦�Y���\����`M��|�&'`�o�[����]?�	m7�>�D�u�P��*HW�6�$D:`=�?���^���Dch�����Ǣ�aSX�5�՘���5�S͈�3=*I2�z{3��S�p�i�DW������+��D�s�4N�p@.�dD7cRh��=+���>=s%[�+��2�,3J;F�'̭)�`-T���c4�D���/�4�;��Cg�Ey7W�	'�4�%���EU���pX`Mלt�y&�.h;`�(}��^)a��QB����7�=/a�'��̧)�g�_�ԗD�G^{����f`+]M.|^��Nl�G�$>�d/�:�-q_�2)aQCs��D���/��?�D5�_����x��@��E^�*�[��8��0���wO��;<�cG:�(|���R6z������k�0�����[���4���э��w�<�a��`X����4{�k�f�3���[D�Dlb�D��DZ)�{�~�I0j��p%+�~�h:���݅�D�3� $��Jg��:ac�*-0g!եNŋ�s-3�6��8m|:!��,@
�>�A�]�LB��A�Hn��[��:�bk⨄����+�j�+�N��5>�KS^��wk��DU�0��=AN��\3jv�`�\�Zs��0�����w8s��BF�9��YC��Z�"C�)�*��Y<΅�߀�G�?3T�G*c�NԻ��JJ���8e���_;��P�׼ߗ],:��;g����-.�]��j{�)TwM�SR >��b��_X18H�5���N8[��+fT,\�"��Y� W�_G {�c�ŶO�_#���~8a���_]�;�z82!U��ƨT!qۣ���C��~I|&cO�6Ui��&�����Ι^��_����3�8���:���?RW/����`���oB���&��Σ�A�5�S��s��d����3AC��;�'?I*S�!�`?�f_C�oT�w�������̃|c�'g?NH�����4��=%hsf]:��|��\|I0���p���G�e]od)?ܢ	�Q����<H���� �,��4���{���i�4�@SJy�'��/s��t�B�"��)����؃ _��g@�XS�]��WZR`9$������TE��s�DTx�������@߶�iD��`]���N��H+��OӜ�د��ȟ1����yc�a��7~x�	c�Ǣ��7���[r���9���� ���U��.���@��bsZ�˧h�E�36X�����g�*1T/��Á90�Ew56ߗ����
���`����\O���[��3�6��k�b�D?|!�@���^汘���ZlH'��mh���T��n��&ͣ,>ͷ2m+�
���ZR�U��CCSa�E�Mޚo��d��qE��] ���?8
o��.Y��$���R�ߌ���33�(k}��:���i�N�1�0��M�S�w,��A����;vY�l��jX���%Q��&��A:�7:x�)!�We��Q��G�ȍ�Y�Yiv��mj��W��"_�z8���R�����q��u$3q��4����?���p�9R�bo�l֬ff����i�V��ǿ�nIBdx�	�P�썍�@e���7��$ԃ�X�OW��m��ߟ��&���KIL�1M��{�Z;��Ų��Z��A�/+��}��#���V��ܺV)0@x�QB�W� H	�K���3[9^E�r>0"��Kwj�2�%G��]�N�O�C�ʏT&+�e��nx�_ڃlvp2Vh]�;#�u��$nE���6ާ=SuR�2�D�iQ��uږ4t��2O��"�V���&K!X��J�����z�0�����!�&W��\+�N�2S7z�-3�2�XgH6�ീ�ot@ qx	/�M�vs�'D�]��i��Dp�F�꒳�v����ˢ�Мy<�+�-س�<tH�S�ևC���O�٬Q�Ģ�_��{	T��.��;B��Kl���瓾#�0�1C,�	���Os)b��O/#4�82�wI%�ͮ���ɮq��'ё���>_�:a�+й4���rMU���?�6c�{�p/:��
$�#�-Nc6���b�oMCD�oHyRS��d:��^�� �~i�Cdpӑ�؝㗱3z s94=.��!���lMޖ��)1P������5�v*��ay�5D�Q�[�ېE����|�Y�Â�'��RR���_~�[L�� �˯�����lh,=�{�Қ{�s{�DY��a8�B��ou�m��#�<���k�^>[����-r6��`��:���5�FvV�S&'��D+O��3�F����H>/.?��_e�e��.���|7�a�k���l�w�дVu�v�U��I����-�8'�gew��#P�c���Y'"�d���򃔺�+�.2 (���	$�Ѭ�R�@1H�'֫���6[Wj�ֺ���ku{�
���:�M[�[_O/֦E�E,��������Rs�-�{�Jп���m
�*���7����U3�__I���'�P�&��.Y绦i�T��7U�W��p_A
E����3��x�� p�\������R���?�Ϲ1����ܯ��]Y|�]WlS5k���B���R�	7^�`�%L>����bc�"2�B�_��s2��AK^��u�g��kAT9B���> UvP�7e<����"�Rم�.u�N����^s�q�/��x�>(5A0d}[p�e�u`E5I���lAh
T̐�������7�0�&�]-OW��~�=�$^B>7	�Ք;���)hBc
=<�k}\��^�3e�፭�[����e-)O;!��̨�],�DuX׬9���%?<�^>n�����B�X J	�2#+y�gW���̂�tOE���dӇ�y�p�.+[���b��ea�a����Ii����x�x7q"n�'�HQ8�?�6K��"�.~��'&��h�
�[A�Y�J��wŦ�+Ny�_fn�c��b��l1�:G����8�+�c|�]s�v���=9�z���A�>3��q:_E�k-��6+^9y�7���� �G3E��&��/ ��S�:ܲ�8�S���eQE&QM���E�\��ͅ���M�Ζ��ݩ��M���k/`�,�`Ro�H �x< y�j�.�\�"X��ӫ6��{z���;EP�u6�Z0��S�Y��_ҝ\��]�g�������!܀k��7��g�H�83���U�A�X�����50fL�?�K��S���6`/֣�r�5��
$r+��&L(��;T��nv�߄F�vD����,w@k�m�tL�����J�"����#�狠J䃀�ƃ��'�0� �\ w8;E�����] �ڋD��FH8T�QTС�0�c��`/�]�~���`�}�<L7Sq���Z�`_�8�~9P��RT�7���)�M�\����P�*9���� ;���W-�Xiqo%|YEj�!𻑡�:�ǫ0��6���Qҟ�=�O]^Oƈ�+��0u��AK�߾�\E�$=D��ąT?��`�4��UY��3���h��X��˙��x�+�q�7y��'8y���gº���"�}v4��=Q�<Ҵ�p���j�1^H:��yZ�)�o���mVXnH�h�N�V��Os~�߉I�,��Aάl=d.�E�6��) y|P�a���
��(���_�ҋП�p����ml��"QH�:��J�h�S��Ņ;��3�b7�͌E�K~��_4�~r:DW�̨6��
a���a�8G��C�oF#�1
q˪�.����B�`��>���J���Ҿ�n��i�'�����A0V�M9��M��u� U������Hظ��g ?B[�s�g2U����f���A��J�=繡�cix�Lu�],��D�S` (O�;, :2I���")��5�k�b��f�v�\{K3E0���q�+��:����}p�#��ɘ}$(�`�;xRC�$�3[V�u4�V8��K�e6;VW�HS�:��@��
&�
ۄ8,��2�I�k"�sԭ9�k[h�W�X�#(UF�N����țW+�r�y�?K�/�YA��]O/��.W�}2ns+�(YkAvsf�\�"��G��}�n�(7�C��~�v/��w�v~g�V�z�馮���nQ�7x�E��~�p.��P��7w
�Cgay7Wj+��/kY�ɥ�Z���+|ӓ8iT���s�~�աq�jh`G�X��`|��(��w�[T+�~Z����\f'���s�G}��+X^X�踎��ZC����@W�\����Ϫ'�'m �~�v��Ux>(���ǯ뷿Md��1)�\W�3EQ#A�X�G�'����ޭ���Sq�5�ӧ�O��#�۴���]�(��bd(8Kd8;c+�L� L� L� �L�5r �?�嚞�'����ۣ�yjY�Z��̻���n<֢3�W�O�Q=�t]��8�-��#��b�}���<��O����y��l�ZoT�	�'��Jٖd�ތ�'����f��3a!*զ�W�*)V��Wk��������[n�2�w�G�G���J�������)D 8�#�8U�;�ӿ�A �U�;��S�he3[8wl���2ܬ� ȇ��}���{���[8w��VU�e�ۅ��8�3�HU;(��eӧ�9 �U�;��c�x�������P}w$��c����`O!T�ݼ_�CO}L����s�H7�g�OFl8�Qԅ�q�3�$[2�z*��S�1t-�WR4TZ���\�M��r�2i)3�Ĕ����$��o���	�C�]�>�s�ʄ�u��t�|��R�]��(��CAyd�WpP%qW���5DD	�{X���o�|���|8Y�=z�I8��I�T�"h_�|\(> �SY�{�e�-�O���N�E�;X4Mg�$8E휄f�98b�8z�8��I@T�"p_x|e(� �SY?{e�-7��h����=y�:߾��C��k3&7�@�c���E_A�;45n�Zd' �q0<K����t8q�rz�A8#�sI{T�"�_�|t(t �SY&�{�F�(��������L�[�~���k�]����8)�| 4�z�],뎝6�P�z8����~�S)��IOT%�#Z�dq'3%L8! ��:6��s�87�|4���]:���6�^��9�%���a��#@�b|��''c[A|�L8w���:D�Ld�8E"���_|�@k�0�K$��y�z��8K(�||1T�f(ON� � �R<��7o�~	�+��K9QY���u�����T���[To|�6�xX����8��ɟW�#��{yӃ��4C��P�i���<�~�Oa}��"��Q�=x�qc�^��u�,,���ч�ï�����,�Z�C ��P�[M�#m눵̐4H#��5�?*�1_����e{��9�hÚl���[���K�;u��+�4���S���Aآ@����u��˂4��7*z�;��6�dk.�IITkr1�S|�%?�+�W�.Γ1�u-�\��+WW����U��ﴌ]Z�|	{>z㟇��'S?@b��j�P�x7�0s&�3�a��T���}�^B��s6�3�a��b���!�7Pd��f�\#����d��A��3���W�\#{�${j�G��}�цjE�$,8#���]	u�K.���Z��5;��$؟A$�8�8W�[x��`h[�$�$fE�'���W�9�E��PK���ۑt��AW�;�LC�-S�������7X�?�8PV�Pݐ=_ܜ�P���ܨ�̓+cT�B��f��a�>��eU+;�G�8G)���<g�{|W�(qŀW�`�F�����T3?ce�R��s'a�ccSYdfC�8�uS;�G�8E=((`�;X���#7]So�C�S$%�����k�_����eK��!*a�'���	�ܫ���St�5�ӞȽ���͢�]�~��3�nH��U�j�ٙ�p��q�~�N?e�>�U���>d�%�#Um���M*�Wz	trs��b��i��U�	p3k`>�@�l�� OB4XR{O�t9�}bQ��]c�Ε�%.�ņ'�< �0�fvp]BH+��/F?Õnp�3�d2rsa<��a�Z��у}}6�>��a7G[�����A;XJ	w���Ν�j�n�B�]�؀Ui L��ٚ{�(��Z<(�k\\|�o9���{�KVc�h�_�]��&������g�l�9�>���w"���]>L��0��Psu�Xg+��#Q-�������e:�h$}�_O ��V��f�Ad��l�W��� <��4e[,wX7_������K��Ipv�>��(����N�m"���9��p�f�Y���p���XC��:�̰K�����[H�XKg�+<G\�ġF�Z�Se�.�	$�K�آ�aiΓv<�߲�s 2N�����!����uͱ}�>�؏��(E�
�u6q�E���"ȳE#d��"N�ER��	#Z_E�qT�"r�Emq��"�E�q�"����q�8"��"�q-Y"5�.�q�Ey'�FqHE�
�u6q�E���"ȳE#d��"N�ER��	#Z_E�qT�"r�Emq��"�����B�`�qE���"ȳE#d��"N�ER��	#Z_E�qT�"r�Emq��"�E�q�"�3Tp�7 $��*J���:c�����m�p��\G��@M�,����3b�M��Щw�)�<��tE��*Ɣ�Ȫb�WꝹk�@ʹ��B
�	K�'��9���f���1��Z0fl"��E�t͕����π�T����P� �;�v0*�(�8j'�e���W~5�@�+������ҫg>-X�n�C����d�#OL��k�3K���Mȋ����X��b�`;�� rp1A�G6+�U#�RF*Ƚ��%��T`+����Y:v�����Ng����0���1K{;|�&�����R���X�@�KQ#�4f��_=�~\7��G��C��ր`�{g��TW!8�����'$97�Js���(X��T\No�ibA�������}��E�X2K�K����Ө��m-�"��EW�a!GEn��
��I\���_u��wy�D\3�}��7�*0`�#g�2�»W̍뫦�d��{�G�q�!�?�X��$#?��왡4��g$�,	R�R`%M�Q}�M�,�F�[�����R�� ������H���W�`}n���g��H�����\�=E�m�ealmB��69v�R�U�'�.�� SxGp�cj'�X��$S��~^a%�fQ5���dU��+Q����a-"�Dt�[s%�
��R%*#bkq B7T񹇉P��t��*5P��v
��������x���FG >5�ccҡ�X=/��pHW�a=��>��b;^3\��2�2����@��~��@���GMy ���D@�\qGO�yCOl��S-1R��|e�$<KaUV��8����
����yyuX9U~R�v�y��_�ߗNB=�����I�����D��{�Wu�B�|�f����#���Q`�,C�������P�@F�0�g1�qm|�W��4o�&��I.G��K�H2���8�}G|r�R6j�!�O%̘�S�jV��h��d"5A��as^�U>��v�h**W3��e���3,��@I�w~�8T{2du���!'R�@.P>5I�4�x��*а�y;��%���==I!h;��1�e��4A[eN�\5�v��X@NW�nw-c�z�M[vt���1�@Mq
�Q�DAW���D[X+#j�~De�@e�_(���+�'
v�> tvD�����+��c1&k+��!O��aS=K<��NM,YS%GBJ-r|�&�H7�c`��9��C���ƾ]O��FH�ey1��ț9�*�[HZ��;p�rs�t���D�Q�w`0~�t'�&b6v^6��6���k�`��츋�_Z�d�*�.8wc�@�+������K����c۾���?��&H^ t\NBO� �_êDY�_���}��2]�v�y
������J�Y����+#,y!\��]��4�y~��	<5�`��֬��ٕ�+c³�^jY\}jWG��H_X�hh�8~�z�t���dJ�x@�6\�SHV�׽��^-(�u�$���H�+�3 ���Is�PmPz�u��YN�I�P�q�`��|+�C�rk``��$_Qc�q�+�}/ॺY\+F��R���X^كU%A����&��8\	DE��ks��D!2�-"1<�q3G^o�y;4�G�2�j5W;g��U�@�y:�9'��?;��?�j���$P�9�q���W)PA��W?�N-m��b�GH������#��8�l!-)��'	*��W��#�`�sy�o~��("�B
�Z(�QY�3�S��ƼWD�*~V�Gc�:��
�L�q�;��^h` Ѱ�,����a������������٭x}X�w�o�O�:�8����5�'�_���%����V�D�e f�v��i/�]�4�\v�y�v�.A~%e-do����#c���<9DBZ��.d�"����d%Z�����9���ٳcAN] ��2���m \��Z�8$s.�dl�[������u�[�c#_���s�s��J7[',���,�,�6)���@�B?O�4���M�L`J8L��bg�a�}Ǌ!�-I[ �{?t�E���x�h��.�/�|��OMU�yJ���{�2�H%@�M��1�a�eTf�Ck��� _��|�k�8'��y	xI���[Eʩ�*J�WG% Tk-���1v���:�w�O�Y<~�r���X�=$8	���	�aN��[�k��iӍQq�)�ipEu�x�e��_�x��Y���lm�E�r�@���r;)����^�Qn�ɼ5���K�o�~���e^EhN�V�FiI6D�wr	s��oټkh�Ǉ� Zw/z�n��T��DV��(¦a%zڴ����B��?�M��4"7{E͟�D:ʦG�
�DU��0�Wр��C���wR�5Ӝd�t��΋�1�U1�����=��4K�lv6*7�
���sغ^�51��b�
�H�Y���1�T�3��� ����}��o����Cc�K��@���w-`E��E���D��<��(b��.HIQZ��"/�S�L����G^a��FX��r�ǳ)\r�C��~��q<�Z�l� �jF�	����'q9c̛$ �S�rx���B�6:����1�mC��p�Y��k\��*Λ��tn���>I!b:w��Ύ����Y
#���F֜��5��"(��R8nyR�=�c���j��a�"R�jF(5��[s��`Y�Z��L��]#q����!ܕb���hYA\Wqj�ZX��\��da���~����c�,�xNE�׍uvM
Ii��� Zkʯ)��<���l��� �nҦr3��S8�0_�O-E�@�p ��7ؿ�a�ֿn!j!������r0g���b�7S~��Pgv�k��x�� ��b��iduO}��-k�Vnۛ�R�>�^��R�D�[g��<���&YǞ6-�v�A<}�7~��:1�3����?ވ1}d��F#_ߐ�*�u�#*@�3�SWrJlv�n�W�q{���ᡗq�����E���զ��H%�p|���l�7C�)ݍ&������^��*$i-�i�(� O�Ͱ\O�#��{s.�؂�G���Z; ��׀�����u���8��i�a�	8�I�����bƊ����j�p��=7τ]��������]T���r�P�l�7��uVh�dn����l�����z�V�u��U/_�+�"5���!���M|����t���wl�H�Dq���.�3g�)$���Y�+�*�n�Mu?ۨ�oҐ�s��]$�W'�sˀI�<.S���C>cF�{8j�c%̀T��[�`j,�K�K3�N�!�Rqˇ�Tx@�R�l�^'���u8(+"G�5�/«�M���C�%���\�?"��I��][^���L�������7���]�*}jDtn�7��]��I�8�����-��;=��jI���h,��V|�(r�C&&BB�Z�K��Z
�뤃d8�7P��K��J�x�L��R�,�9P_��Y���h�������V���+���G��pDKrL���΂��a��NkE��_T8��-$�@���?�.+X���X��q�o������T)��'0�(n�Pw���K���W�̺�@m��f����7%�U�v^*��
`�F>D?k��#�}�"�W��a2�X�����Sq*�����]��#H�䃦��Y(`���M��=V�>T�K-����9'B)���Rq�6���߿�������H�AQJ�9��@R�I��35``�ӫd ���b�Z61WB�%��4V=�sd�|o��ԧ��[���=�1d7^�����[�e�!T��W�_�%�@Υ=6{��k-�C�Iـ�K �)�>}�9_�	B
*�=�`�3sR��0ևZ��2�GEAF�?�%����"���p8���p�|�p�⟮���tKx�q�{ߠcd4�)�ůR��c"��5D��:�)�{�)\RӍ��U�����`#N�f(C��<q����G`_:(ԝm�N�:_�<���4�De������KIF�)��^�`�)^��9ɀ_�ː^3�Y� ���#y��Y^����A�d�!�v�8}��8	T�Q8L=*9�|uV�^o����0J����W�����Ɓ�8�@0x1o��h"5������I�>�5o��"Ai@x�$		�����q"C�$�cN��ҳ�[ Q"�G�3}XνpTă���E4)<O�l�u��JD�� r�.��8,W��4O�b���r�E��s�:{�����o�{6IBұk�YsE�n��2S��I!�oG��N���<b��(�Skt ��"?�����x
<��/VVT�ܓk[w;[���'��ȁkX�5`S�<<g�I873����0^�`��V��.��V��KO;c3wX;� ��y�'.+�z ���j�[lo�'�8�����f��X$=_����u�TO�<h.E�G�$�.��������Ң��m�mk;?
F?��_a��'F��"�j�uS=4'x����Z��I(g�#e?�0�S�ڥ5//�B�.��i&f��8�T!~S5�Ķk@5��p!�Y`�F�s���7u�kO�<�� ��v�׸�c`��-=��s�	�AX������b�	E?'�W�g��%'�!�VP�<;���O��	F�h�|9JA\���}/`�#��G|�I�@�f�L d,����YE��K~8S{c�y�C`��K��y��ZB\QM�3gm�3���u>/��>2,�w�^x��T�M��>�����g��J�bd�2ѫ�tN���\W�%`]q�B/��I����`�;fM�-4c�M"�c������N���y����=F�]ZN�5�t���P1ME|F0��E8�ͮV�-�(U�.,K4>!$�[E2��ă{$U��Y��A�]�l���&I7N�N�;*�7�'�:�n�$(�%������v�]b��:�,�8�/�+�<OB"�\d?���Xj��YbQ'<J����tn�=��%(��W�`=�/&#*�]�8�`Y1j��J7���ys@� �4��c��'�M�Iu� /@  (9��ғ'�+/�rF.*`Ƹ�J#|u�0@ز�y�4_m. #�?r(K��t@+"fgU�%�D�a�&I�G+�앮p���)��:*�у�1T@Mc�ob����r�k�M�TT�-o�ON���-��^E���1DU���HT�N69�'LWqRi$�B�_
3�3}������O4�JR	 �3lG?%*K�.,��
߀�����UT9T�Q*�E������L�7�!i�)zb�+Sv�Uy�M�{��ka i��b��o�`�ꇥ�f D!�m�7܌�5L�!��x��O�ֶ�B�[��;;�bD�~0v*Q�EГx�A�_|]�4lG�H+��k����?{]�
qT:C_|�I$r�\� d_��C���0am��^b��G?6Y��,��j+��>��':��0/	�w�1�jEH�<9�I^{��Wh����'�b���]��&?[�<Ych<��K�\�b"�����mSa_�>�3l����e����9�}��?����.�ک���{�U���5�(�1�5>3��o:f���!�1`oD������#�W�6H@.���\2��%��~�e�l?ny0�4��%�Sss���4؄@XT �B);S��:�Yj.���x��<x8�ȟ˹D�,-b}����</}t�[M9׸�_��B.d���T��a抷���[ 3+!�K�6�$`�ML��H<���)��XhV�Y��&҇��0���N,k�2aE>��8ad ҕ����ܥh��遞h�E����-R@q��壍6�sW�oх��1b3{k�_k�����g�� !��;<W8A�F��W�~�l��D���1|6X�F������@pb`��eKs���"�C�c�E{�@MyQnl��&8t/#��-g+w86&�Th�l�cz����;��S���@�Yěd�ӏ./.J��Kۿ��.O�i����H6 UG�kLV=s�=o�C�Q@VU	 ��`�N�@��&�!O��L2@��a�@�.�����M�0k�nb+`�x�Q&@x@���[����e�^�fS�8�n�/·3�X�94=~�� khOGj�Bnr�)ˇ�e����MA96f;���^S��/�v`G�+�#��Ho����0��P'D����-����\��'�C\��D����Q���$���:7ie�d���a��Ԃo�57�#EC(��'�`�F�^r�;�t?-/��m��Y�GuE�E�����-�j�hBqv*ul-�f- 
���N��Se�$�r�p ��s#�?G��`f���P6��o�MSWnc��<�H"���;s�#�WQ��8�{��! ���QLEYcRa-��=���`�(|�Y�/�I��
7��IDn^��RCYUD"��+�X�}9p��$'�=��[Coe/�3 �qЃQLdi�@��@���R+�L�r���9�E!��Str$M�0���K��рv� 3z�0�R-�z�?LM��Mx�f����Q���'I[�s�[f���[8mr��eG.Wfw��/����Q��w�3c�y3��Z���1�I8{�2auk��XUIKo�ٍԱ&`d��E����x1$��`!�O��k�0l��!j�c��8I��6%{Xu�gкW7<_:�/I�E������"��᮰Ve����_�N}F8��2D{w�Z3K��w�dt)d�|�x� �q��vl+�u�ʎ�a_�:y>�pp�-!y�y�y�=��: ��E�,��6^�4�'iL~�F?kߕ �Vq���-Bw�Yxl����;�B�ܕs674>5�b\��NAr���WF�8`Z�D�E�jc�@/[��o6W0u��E������H����͉�hx!��`��ᖠ{���\i.�y3,����^��R$�bkW}��|t%��T�\�=KY�#�Cq�����U+�dH��m�L�I�?�˔KʹCb$�����c��b�r�-���4Y�۩@��;�L�S����~�����ۃ���M����-9D��)$W��Q�Ka�Gj��.i�^l�%��
Z��Ȝ���1�
�&N� _4�r:ye�,-y��X��\ M'��O��a�R��A<�KOC��h�����D�!X��_s��@k���B/*Rj��Z3�je�z8FE֥WG�����U���4���#�
V5]$⭏Y�*��~Sz�@��I�9����j�A�̇p �W�#%��`�?b��މoRnI��gN�����ep`�n�����"�"3x~�`/��J��"�A�Z~ވoa<L�Nǚ C�NR�6�PDx1˕��8)D;�N�Ӂ0��;g|���R����W3z�Z�$Z���k6rl�[ �34�$,a�Qrv�r���)���A��*@ٸ}䰫i�!������d61��0d��9����څCh7�}B�*t�����f�d�{k���1 �27�n�Z]�^�<�qI��B��/N}O\S�����/�!a�o����Ί���
2C�vS	1�p(_	Y0��~0��/w�4x�()M�M1�$�$�[���Ph Tj�!5d���K�a�ѣ��y��>�C-�pn�=F5P����dx�$�U2�NU5'y�c3Й�}L1�Ϗ�8�{	:�8�=�kdQ�h���0n�Yh�	ZR{.d�����3�E�����T�1���*������/SUW��1�d'��h\U?��0\�� �f�oY��f`�7K4D-A~�*�w�m'~t�*0H�L��;��26D���Z�����뇀�հ!��5z��8d�Y.�:�ŝ�T�Y�dQ�����s��!�v�� |(RO�óL�Xi�����TX٘�����������0�^�o:/Ӓ�US��Gx�_6N��by|	�x��R�I�� 8���>��f�f�sd}�=e� ST�}�8>N�\�1�8b�`	or]�䡡��+���γ����HL.J�N��s_w���$�dp��H�i*���x�ۖ��_�\��'J���[{^i�L�eYp����\����f6��*�7�����v�#�Ô�Ow�r'�h0���Y�j1|�DU�fSpJQqnO�V������륾o���A�tb�T|�o���B���Af�n��:|4*͛�������� �W?��y|�x���iM�i����dW9���aF���c*��xWs�)-����ȍ�
q�nY����Jh�yDO�!�y��<H�)��Z�ƋZ��E�{�}�Fѱu)j�Մ�T�>��ӳ�
D�0W����ބ�_F<�_rɨGk���5���&Z�w����!I	�bUH�3s]A;��u���P��ڧ����*a�{�{	g.�m�3��T5���͝�=+�����=��E�1��BSU�zFQ>v:��{8�Ug!g?�>���@�YT��zV�c�_�b���)��D�Dy@.;OM��2�߀?5�Z�C��3��eÝ`8����F�����|
f��۪/=[���8�h}�iq�S}ҥY��eh,�m7/�?�K��#Eً=�B��qv ��t$E[$�8�<��K����33��}�%��]
��K�u\�z~�E'eE�dT��]� �_�[���e���k���w��C���_9K@+]L �����w3��9U��S�B��Cw�+�m�{���|�����,���v���<g����/ ��r�h���㻻uaږ����U���bS�h{���lpcCah��L�'�E�D�<�AQh/9cD4�|��@>p�2}�.3���9����Ҁ��@|�+V�_�g�~a�Lh��,�b�ӳ־_]'B9�G�^��J�J��
\;����}����X�;��W$�br�\8A��d�!�ED[hj��H���=��yM�EN��k����-��"��8iLdjE���yi��u��(lD��1,mX�ڠK�R��z	ӄaI���N`�!�x[vozm�-�T��f�?6��%�U�#*Fňq���7��V+
�R���z�"�\H�QY7��pH%7�І"�N�V[#Htb�6�{Z��З%?%����"8�DYvcND
j�?���'S9�Qf�'!�ƺ�vj���s2�da�|9}�rzo�SxI��^�Np�ܢ�G��}$�.�-�,�%%�o���Jju�cn0��#�?v �F�L���������9�9�J�/����	X/Q�9J�Dn#��(���Od��x���ir�_S!��q�#�t��-$H�L+�m���/b��_��rq�B<Z������*x		�f��d�#�V*����D�����)ƀ,�Dɏ�+XƊ��2�W��'����ZL%�ɤ�����(�K����L�F��/���2|߷un�)7�0C�8,����L�5�u�^xe7�O��x�
lb���4��b���� ۜ��z0�����j�[/�9��8�FN��	���.�/>�s��ެ����y�o�^	K�1�9�"�1g��;���4�Gs�*������iJ+s�	Z!��\�hC�a��ʕ����U_.b�;�w��K��	w]�L��ͤ��,�ǞFY�j�)���SFN*������_�x�+��W4RE�/O�Q�۞�6��Wx� !2u`�RcWB�3��Q����>��ҷ�����d��9���<���/��f�|�d��0�OI��*qW3�=LkuSx�@.��L�.��W��9�xWf��A=.��K�f�?���T2t�q&Y��^����Up��y�;Ͳ��7~��DXM}3���8��ݙc(w������r͐�N��ޭa�����E#q��y��>����l�Xsm,QΘW�7�1�,���a��2���.��*���vt��&��!�R�O����Ei��k%^j�
_k���e�(Eg�bIo��&=�<l-j�D�-KSm��a%�j��H����80Aޝ�j��8�So��;���~?�>r�6�������Q�1�0��f�Qf�̜�.�4������}%�ﭰ������<H�5H����-"O�\|n�/$<D-�#�W19�Dͦq�V�1n+�mwdO��.�a �\g������>V���L�X���]<ȩ���G��Y2>D3 �2��q��,�s��%+	�sdE��`�iVח�6�3�Ӌ�@�Tk�D�q��e/��K�:g�u�G/y
g/�f��}��2RBm*â���'�	,XAM�[��Q� ����+Y��X3CH:��S���d&�F�隲�(�P4�(�x�1�Pq��bWp%����+�����Y�E�rg2�DF��&�Ѕy*U��
�G�Q]o���"�eZ1��$��Z�jZ^
V��F�EBV��'#^{4/S|��G��A��! �N�Q�B�|�q6��:_�}2�WE�]�X��q��CO�	S6�������l��S��6� ����IP.�#[�U6�38�z�<mw߸��#HL��U�:�.D`e��8�O�dT����<�`��{H�)$g�_�ʿ #�s���4��gS���{���ͯ@��Gx�B�$�0�7lD�O|���ߗC/~����'�Ks��"T�����-���r㟏-�7P���H�5(���=t
t�����S���l�[/׼b�bh}�pS�M�EWl��������)�1�˕O!�ߐ(6�}��Q�ao�C_;��K��MH��jcE�=';�)IKHYGPG�T����'\�K�eSH[I��?��o_-����?�����x�ۄ^jpdQ#��\��A��S�����ǻi�!g�����bl���>!�%0,cI�'����X#eS�<��oHH�g�<�}죀z�TW��#����[��{��'�Z��-�Qᜯ-�T��g� �y�9_8���3̩k$I�C�I�)���C��L�a�>\o y��KK�uS�g�k�9G�;t�_�;O�O� �̛)�g{_��[9p�;s}���E������=e������`���b��F��"E_|F����ߒ���=��Ս��g�  D����                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                            I��F     � ��  �   `  �   H  �   0  �    I��F         �  �    I��F         �  �    I��F      1u    �2u  �  �3u  �  �    I��F      e    �    I��F        0      I��F          @      I��F          P      I��F          `      I��F          p      I��F        �  � �  �      �� 0   �      �� (  �      �� �  �      �� 0  �      � 0� �       C U S T O M   �$B's"v#z(U`Bw0l"j#kԿ(c<%$�!���)$+&(' �-$!�,M$a�#�DW�L�I�@�KCJ�qDVd5HQt߄"!��q$�}v�iL Bo���,-g('UeC;uP�iA+P)F�k��HY7Er�wABR�"p#U9����1�9Us�,�Vj���#'<�MQ��29	4/`�6[We4�I���V�G]��37jc7UB�h	/�[��0M�N���b=5�=P�95��l��Y�m+���@5,q!g��j$��&�-�"m'6�.��&�-"'�6c.$�-�R�#Oi5�>*x�]-�>�gG)+ū,��"h)/$�Y�!e��e&�a$"�*.�Z1�g!�e�'J�$ժ�"vU+�'"R�4X-�$g4`+.b5Z�>U�>ͭ�?O9��"+�?5�+��-٪$�fږ�#�	Z$�:�c"�--Z$�!�e&�"]:ގ$wj�Ӌ�y���\&�*"ŗ5,Z"؍�e��e��5��r��?�h�&��4��e0��59+:V�ő&,��$i%/qMLVUWJB�DH8F9KXQ�G@�P[DL#ajv�HJ+A@( /au`$i$�� v��5�/"�%'.$P �-��c�7a6�̝02)|�!9��ذ$(6+[�!�v�-�"��M-t�(���k��Ck�=5�1���5IY/59�,�0�!&:�9Q@]�0;"$��ɯ#�m�E9ADQ�<"y�-�4+��ee�9WV�F<�C�P�ŝ3U@IJF����1 [Yg�z$��4��ߥA(,)m5�JUa7��37*1m4�!"a0#� 7&InCv�@�,2�VQa.B�C7,m�/ 6�b��*d��5�-eJ!�,97mc�w{aK��t����a�Ǭ�6!?,��my�Q��4a��<�,��<+,�o7Om_�$651,'�7C4A,aI�i7��m]���a�׭!1�779�C�,q<AC,Wm�����,�<��,��a�ӭ'0�<d��,�,�<O�,ma��v��,�aᑬ�6��T_ �>q4�,}6�<�5�,c�${�4�Y]�,�a����7[ U	'Km�am����`��$'�KIa=��7�Kuh�U�,�9a]h�u�7��-5E3o,U�m��1a#���7��mɝ2a7�<�9p�ɦ`)6#8*�]c)��u..j�m�+ �d��P1#e5)�-�0�,42x�`&�a�s���@�5���*��5%� )=��Y+�$�O$������&��o.1��e��>�e�ػ4M�.�a��E2��P*�;��1��4Q�Qu�P�O5���U͞A��7�{�5�n�͟N����.�!���dtQ) am/�b���U�?g�!}Ο�;t�qyb�`�u1��(}��ͱ�s�e���vy3�r8Y�1��i�� �j�k9!���2}��ae-���"�z{~�Υ��"Ӯq!j��ǌ"��-�d��T=�i|st�f_kc\�{��Ӣ+���_�Ssa|�æ��M5l.b��4>	@�3�c���?dٱ��Dt�Q7ښ��O�f�=�H</kh�J"QLC\rfKA�RfIDV�3=苴-�	�^�7!�iP!�q�%��`��4�m��*���5��:���V&JFNb@�WDI�u��U57Q\X]B��hvrlk�fSn���61%nFMH�5L�DI�CQ��v�f��I	�S>�VL?�5�I�)�8d�o;�-�1-5a=�4,ؤj�,Am!�1�_� lm 6@װgn�K�$�3�mB��C��at�#���Q�4��'C�'P+n�7]���b��F-� {Pń9@�:�8h`� ��<���l6Me��_iWϭZ���9��졮y��Q6#�$$\�5�s������GnE�f�rv�)�vLy����^��s�t"k�r�B@�iQ��\MH#�?��׋��6�sp~��!��*Ԭcmy�i�YdJ[k��3��x{~�ã� E�}vj�E�/���ّ�k �)�6�gu9]�e5u�4}�1�+��>9�3���x�*VDt-�5�d��hqԆka}(�.!�0����Cڠ<��H?�C�$Q6�@*sB�{�Evvr�#x02:{y �͇t��e�`��[ u��͵7	f7��.`"-?�݅U�u�1�~�-�Ia�e�3\��7�$��/1�' {e=��|c1m7*u��Q1X9fg�uo�=([:rpN������qf�[�fEY�xz�=�T)�)P'����E����9E:M9�&g�4 �Jg9A�ͣM'�ru�)���`sO��}�|�V�t�fl�����@{*�+NOZ1�X��1u��L&s�A�-`͟,s��*��$:.�5�,x7�)5�o����Kl)4
1���V�T��')-�7�I7+�1@[=1��l_�-a����,P7������Ӧ�/>�:��D-�,ݵ���H�A?ܵ�5Ea�u��u�W�yX�Ec���h�)`�#Ť�'�!�#ݨ�)u( ���<!62*�
f�h�1ٍ��d*���fs���m��-ܐeQ7�X�7����i��U�uM�(̈́��nd��f<$?S�aT�8�?3M���O����c�`FDY)��h���U�s�H���OA�	�M#�|񐤠րD��iM�t�iD�!c�^�Kc�qf-y��I��Rx�x6Ԛu�4�)��6�L&t6N�u�a��� ���E���!��4uD��r�� ���$ M�2�62�!7%�baQ,wc��4��9�TbԴ���Q�ݗ�;��',!5E(��4,�i�}}�Am-�i)Y�-�!��c9�gMϩ�[+P]m.#r*��u��VX��G)<YT+�[��cf&�j��3-[*M
�%&+gj�@Y��?�dxk��h):ux�id��l�o=�|�l�Wx�Of}h��A[s��E?w{wVe�#�#�45��+u��z���v7L�AExc��:�/�c�c5O|�,փ�zd�doAh��`�a���kz�&�]~n-db' ��QA5�}��l���(1|��x�qlK�s��u!�=�����e	��'P����e�k#i�h������=0��Y"'gh��G���Qv���P�O��7�e�F8�p;x��Q/}ӂh`��V3~7��&)���,]*����*�OE�sY|�[#!�>���e���$.x�O,kYQ�F�ˠ��a��@��FQy�7���/𥏟�d#��Y,Pg"��8a=Q-u���v<�p�{,4-�2��)n"�qOh��b	p~�/��~��-�
0���e��,��e*��m���w�x�q�O<@s�T����j�0Ѳ%��>�c��4It(mn%�s<r�xX�1�Q �*?P�Io���W;-�'d�"b���:1;��:�o{�ip��;b�:,$��V?���$!>4*�-�)�dWʮi��ם�*V#do'�W߅�O/�\�)�|��?)*��DR2�+��*>'�����!te/�c��z�=���r����Ʊ!"�e1��WdbS�?54�Qw%$���|���K7�X��p?ib&/1vAj��1+Gjc	 x�]$���1 >�uN��v,�)Ctj=�S.������P>����m��&	Mh����u�0���*�oe<�������2�7-��&p>����)�-��g���?����w#���&d.9$g#���}��M"-�5"5e��a�mu)ift25"q��}��y�GE�=A���-�"XՀ�/��t��1M�0��0�N"�ҍ���Q3r ����U1|����T�n���4�&!)$A��,i�IA/���`�����Bm�Ra�"�K���լ�m+8��)���?�LB4 �K�a5tO=�
�7n����c`1�15=�����,�-�n?R�or��7&!�gqD��f���f�fZ�)�)�f���f�f�f�*��U�,�1�ǆ7����U�u���)��)��)U�)m�)�)�)5�)�f�*�kI�#U5Q]ZY���A�oA/���¨Ù0�m�#���A��<�)���-��@�4��1z��$ �-Åmsw�5!��l����O�*+;�g�k��C-?	���Y8d?Um}�u��u2]a�7�C=���y��A�*�P&�c�X�_�e�`vڱ$�Z�ei�(��f��ݣ��5ni�N4r���u��o,�r�S�5c��Ig�9��(vt1]��}��X���m͐�YU��rʵ]�l������	=&(֎O)[!|5Cя�3�g E��!#���-�#1))�`5�*�vp/����=����w��?�(��="@��(*���)9}]x~��v�=����`�fb#d��@���ud,���'�k!��N51�McJd�Ea���sjml��5���iy�{iOn5g=�[9#)'��7�y�d�\�hjLܪ�l"s-A%{��(=g6Q0�d�r�;��u�4ow)��=�=g�4���M-u5�֬$SQ����:���ݙ a���r��nd�'-��u�Ck<]s"T��5]z�k�R+WP-]�nr$�� M]e�Wd�=��	5m�X�)��,��N���t�x󐲅��\�B!פ��	C�ϻ���7I5�V��7b�SVU�s9>*�.>��g�A33��eZx�*����A��w)+�(�M�g3�� ����1��q�Pu����4�o�g���`�t!�|�m_�e�%��ӷ�V�A(�ns&.���>��*>�(�\C���@})��X�_��|�.�>�m����#/T�н�^̧�	�-E5j���.�15�}M����;�5iV��Pd�]��J���fg]�X�Uu+T��.�p�/́�a����^��<`t��	�w���q;Ԯ�5�ti��A�}u)@�1WX}3�8�-A��Y��v�m� "ojT����eV2S��d�:-~_X���X)lg�dix5L������ǅ,=��5�j!���"�6�s�c�t|u�! ��� ZU	,QM=Td�b	t+��z#C� �*U$�=�b31eQ&�k}&dig��e59$�k��v)w����R5�td1&�)��[��Vkt�6$��9 Y
�ɕI-r��mU�n�);�Cq�=f1g�*��/�k7. U?��ѾP�c��/C���wo+�{\,7�6d�[붎�pwg�FUQCa!�7vM�q�|�49���7�e�a�acK��Gڵ��� /cu0�8Q.f�i4�}?t�l�Y
�� eP� Z�_��W+j�Ry\����l�='�#�pgdy�\�-�]jR2¶�#��I	��C%A/*�����ϸ[7g�sC ��C�c/���6�Ʀm+6���WC,��#�Q��٬��.-t��mU���8��Q#���&�,�Me~5�(�Q�iz!iQ
�
���#%��$P<t�=��͔�-ڍ9����P�Rtz�g�[!S����sf-�6�b��,Tr�����z,��*�����!&����H�n"<i�9��b���A���	����,v�Ar�tYj`�����3O}s�����z1�dtq�o!{�u g$2zΘ�ڣ�����qO�/��58���~,� �`*������Ω~�����O��0�o�n�ao�y���Ko)A.�e����5ud��35���?=53�*����f�S=�-8|s� �+{਍��6�$�)me4]�NoVD�y��N����w �\��$�d�Ӕr+�7ҷO\G4�/r��"��UAV�G�S����A�6�|�*���X6���_!#z�=j�s(�h�籃4u����/P�zE��̢4��o��'�g'Ά\ìk~ ���}	W	Ej��um������?&/r(�f{U�F1�J.w�e6�^�j�g���9�n��P��7u�$�;�����
�5R����4+5P1�t$Pu)�)5'��!��;�9G|���y�͖��n�\-�D����]��gY-陧M0�G�_��;F�J6��5ݘ�u����e�d-ӏ��Yv!�:��~�1�Q��5�2f#��l�a�{^���$�F"��mn|N���8s7-UK	̀d�-/�c�95�݆Q7����s�����i��Lt�y\Au�_����OT�uQ(��Iɜ�#�<�?�灼+�G�n��kS�ub��c�n��L��^�0�.�5���a��4�0��\�X��V�i)y�����;횒=�7�9��Zh�	 /�|�m�-��lѣ퐟e��,���a���Zj�I4y�w.U9fQ�]TY.6��W���+�R�A�W�<�9��b�XXg&�k	{ �r6�,q9���rC��/s`�ϧo��f�[U=��P6�C���e/Gar�W��<[3`Uv�mP2G6	��/=+�E	,r�z�g4r6G�FD�)}���L�g$�ի&��?5�����8"�k�f��t)$F��n5-�H5�K5QZ�~7N^m��4J��-f4��|�4Te�\eU�<x�5b�{,�-�#���Wʴ,�5VDaL�e�de�;�t�)i,���5I-���B,Yi5�＂���X=�,[��7��a&Z)����l-� e�7�,:��4�e=�I�t,ݬ�,i7���7��i�,��0r�t2��le�ev�$�o'H�z��u�<tG~,c�!�y5��CAP,C*�,�na���,A���)�,oe��e�_e��$J�&�5�wj�|,F �G`4y#ntG�4��#�,C,a���,�,�6,84�$Ή'��a��)�4��,�����a�ʭiԶ�=��`�m���<�,ͭJp4CYls�]<�IfL,��<�\Ga-�v�K4�&�,Q���$:�ma�e	�<Z,���4&�'Lue'A),3m�D5���\-��o)g��#�,a� w�E5��5F��,TL\w=e}��tF!u!��!.�)9,$w��q���,�)P��,���4lr��<��,p��'!��mњ�aO�[7��c��qM�p�ݥ��]Ҽ�]@4�&�5P�5�lt, n&�5�i54u5�j5��4Jcs`�qv�5�d4�Y/�a/SՍW-�!g4rTѲÑ ����M!�m=m�٢!���a���AMCM4W,`YM�o,q�{1�M	,evM+4=,��McՌG�,!��M��lJ�,ThM͑�d�,�BMc�A�,�vKM��T��,��M�CIdS,`XM�q�t{,@�HM-�	�A,vM�
�a|Mĳ�+4-���-ϴJ	��Wjql�M8[�@-x!��%P	=�m��m!r�g��"�m��Ң.pi=��\��9��m==��m���,�<	ܤ �Fv�<NU��f+ĳ�o3�`��6!��4/$},X���B�4��muJ����Q��Y�<F<�g9H��حFW�-��!�T�L<���`�#�,6��3T�'���Ё5V�0k���H4G�䐱��$�!|י���-T�׵U#
��ԇ�tPv��U�5�"h ��4�$յM%����~��+�4�%�z	�A%��N`>59��-'�6���Ge�U�'��&m����W��k�E�@�=�g��n�0t($��7�5kD��E!�)�,��<�,4��9""$'&&! /��b��t���b���������j��/���z�!aM�f$�5a��s�N|�cl'}��b.X1 s��b���I�sCgAw�s��`�:Ua�;��3�5{�:X��?��� �f�gΟY�CsV?�U�Bs�40~�l�h>#3ue�g�Wj9�mOA_+�~��@�cz"l�h٨�Ex�tMI��X�C��u&�u��2w:�c;`����AQ�f��)� ���u��i+�jv��gj�	Q'0-���-��2��'�Q}sK?�0�C�f����*p�^��$)w�V���m�&.�P�8�X&�V�f�;��1l������'�m��+��&ˁ�^�)�P=�~{��̧X�O=�S����'`���x��Ŵ7�j��r��pd�'ь
I�� �|� sW-�K�N7�t/7��w{Ǭ5s���A�O�݊�t�Y�y$f7*�4;�m��-�"�05��1�⁹���r�`/§��b��W��v�o)��Y]�O!��-5$�#v�;I�@�ْn`1�0(
)�
�?�����M�:�Q�	����q�Q���=��0��ɳ`a�Y�t$�-ͽ��֚��Q�3HO;��17=�k���D�Y2`�<@�G�#����L���T1}��w!>���ֵ�����E����4�1�{�w�H��"v���3dJ�|��I�Y,x�*��o0�.j�9!��#�lN�n����Q9 �]q6Ͷs�@n���+�w�ꩦW�}Q��V")C�XA0FGb*��|�,� (J�{���Λ�Yԯ��9�k3r]t��J��9����B<�1!���v�f�z�g=�Ǿ��q�M�2��7'D���Z����Q���-e�I�CZ?98�Ң�כ�)#�}L+��,fe����;f̨!>'�":��.�d.���q�ǁ���:ĭ�(2�h��9�b	�TO���%�# SE��>Z6\���|}��>\N��m_��O��t�}:|�wH�����FGA�i>��j�!�)Z�^.�$4�)%G�I?
�1[�h2q��x�fܓa]38<Q	#qH�H�"D�{��A�考��t#m9-e=��e��� Q��.�P`ف��v���`�"G�W�j���A� �Y�~�w�w��gt;DD�>��g!2C|Ceg�e���=$��e8�^R��G}�d�!����5g?�4?F�u#5mtI�}r��*=�Y�Ii��7�<��a�U��S�	4�5?`]�{��R�q��'�4�����[{W:ZZdz渺9(����eۣ�����'(Y �	Z;����$O'�2����w	��FU�Y}%A��-po/J��0��1��o�=t.)��-/@�?�'�Ε�J�|L7�vٻ�)�U���Z�6";M�@���o�E4� �-;!�U���1�%� ����o,~����3Җ�3�Q&v���Ap�֙_�h�=��	4'�����=!	r?�dr���Lp�`!�+78�X������P&�(��DO�~O u�&�j��<�b�Ee��e�v3uM�v�̐�w�ty�Su �*�إM�~��an�(��d�u�J�����[�P⸮8/�)����O"��1O�Bδ'[i�:�@�/X��:gL�)Fqc�p-i p��҅��!�a� �VA
��� �+��]�m?C1�u�i�PlH�tpM�o��P��fP'3��K2z֦7��Q�8l����	=��1:�5&O$�{3n��y5���c��x��ߥ䬮7Q2�=4C;y=��)�P
�z�E6���
�l��9��&�d��@Y.u*�`Q2�}#�g�gO8H�dAI�F9�M���u	L�)-�'�UZIs�G�d7�i{�> rpU���Y�dQr���tАa55�Jfd��@vO�s1��:����!_n-#3���L	Y|��lkdSh�tg��#=��q9))�u1�Qe�M�2���J0SGs���w�E 5����M����d4M6��v���oU��Q����m�^�͓_�!�{�,emo��^F��n�!$Zc�r��e.,[mQc�D�3����5��?�I���ߑ�z���cP��o�"�/�QȎ5�g4��/���2�n� &��p��2�(M��!��nF�-'�rQ=*�G}po�FP��W0li?o)��w�k݆�d���5��6/	Q�J�1���dQQ"
�v�H��B|��>�u�������2���J�o`[G����D� �	��&�7��/��XN�YE�x��-
��!��Dm�Yj,}ku�7�͆nT}k�/��}������а�� Ne�w"�����6�����f�R�7S��)��~R�a2�X5ҹ���Zy��z�x�k����7s���,t�|�6�l|�S#���8�7tM��J5�0�R�A�W{�=A�8��	�(����#L����&�<����(�;|9?�A�C�d5��:���m}����#/o��a�,�zy��q��4��5�"o���8׷.��Y+ѨX�A�5���{��o��ց��q7.��a�P���)�kc,k��\=����!uo.ۮS},SD
+�N��-�;��)4{�!�vA8n��� 84��o�+X��T]�5��c�3vͷ�(t��y�T5	����ǻ����[vyy	 A�c�d4�{r���2��[�(|VYQ��)3�Z�br 'Bٲt��sP���7��N�ҾJ��Ew�d"_�,�L}7 � @��9����X�^CS�6A${�V* ޚ�Z �p�%z��Y���gc��לh#�튪a�6w3�,,͎?"��_e95����2*���\���%��9Xq>5�@�54�<z���+$MFQWISJU]�%fivlay^d�gTSRTc��f�/��Ƙ-g��XylKUFWQv@�S0#e/���#̴�/��8�. YR�Q)pi�;��䘂^m�0�
�.�Dئ���#3|�
�[]~�����1����#-M7�{��e���t\!&��N��%�d-P��_$�O/}���֬��!��Q"�<��Z�4m-��b)\�$�(��`\j� �ȸt�4��-ϛ)�K��Pu?���:qܰ6�7��w�6 �Sa!��46)�i�Ta�cwa�^�0���_|�c��� �
:`��A��ҵ��4�Q(t1�D;lmw�� ���]Ϩ !��L;�%)Θ�t&u�U82l�<.�#��7n���K$S�j'��7�w�~uƎu��r��췛'׋����a���¥��vr���۲�?��5n��gv$�5���=�}M'��ށ������F�d�A��M�`|�̝�HӰ*�2o���|��]�o-��(͘bf	��q�={�<ꙍ6'�"95����&+�F�̈?r�F�G�:�.�25vW�9�j5��E?����j�m�?��7!-�A�}�#�+50�pr'=@�o�5��06 8�'�~�M���ĝn��2�]�h�Paϫ:uFP}K�!k2w=�nOwM�Alt2�̘v��?�+^5e���4k.�vb���l���#�7 ���r(-A�t�}E,����ua<A6ٛ�o�ŕ�w����Vt??�|}9�g�^V��7�Ҧ�̓3.����u}Mq�u /j�'���И-�����kt�Ԍ;�m�����)���/��c��˦J)�5{��Z�B?Y�V���c̙>��xbmAaKW�4�+�
`}�4]7�ZG�����$� }z�(�bV�F2`��m<�`�q��2��6���`�`������[�F�:�ñ�)�0q��G1&��,+wusuE��A�&�����5�l�7 �կ���)5-���5$̶�@��F�&���)��u��Ք�-��)��:Í;Ua��,��`2w96M�Abe!u<�M)�l�� ��ݒj�5�A1)�Q �Urm"k=��04$e!���I�g4+�>�e��-eC5�_�u���5���4�Lx���'�mPp@6)���֢l�Po��>��ׁ
O�4�$Fu��6`5���?̨8yI���4��.���M��ur�;�ms�6�O�]�#�A`��[��Q)�t�T���?�B0���{XnD�L��.�I�JW�5P�]$d=H2%��'�K=Hg�'��4q"�o[�	-����^Ae9�}�I��.M�nW<a"sf�V��͗+$>��G�$1g���$F���)��~��yd���N��y�uN2���Fd�=dj�fgM�/��^�Ѡ�yd��%�$R�:_����f�ĠGd�3U���濽~����d�	��fZE�/�W�PF4��PvWQoOy+U�]��-�g]�;�0}�:I5��#�4n�g33T��U��|���X�JM�O&�ح�T^��Z�|�	��a�!�f5��"1R)��[��\���y;Z\�"��K0�45��]�X��6$crMH^�)�&�r��V44i*Q�b(i>��BA�� M�O�9.�#sA�1�x���n�5���w��0�0UNe!��scש�u[J�8�.M����0&e|N�0 �]����'V/� ��	u��H�)�M�(;l�Y��PᎮ25A7j�Xt�1c��M__�dnuM�?��c|.k�K/��da ����By/
~����΄QM`�������P1���׈�E]aH>���Y��7�P.&��m5�Gob��H�0g�)tM�`��J�W��I_n.���wM����%��oQ��$"P�!�������R�	�}�.*�s/яe)��t�nβO��w�nP�k!VVq-m�q�lQs��k[*�n!��-g��#�Y�-����%�X�^!�.)��m�Q��*���z���S�sf!�ӵ���=%��Qk,�5?P7F��U��G�v��V���=ҰW7��8��6�7~i�ZCi�k��S���2�跩C��<y���1�Byl$1c/b}Yl�l4Ԝ�io7�r�H��/�k�*���?c8�Fk\�w��am��!ng�1����~�z�&��LUuQ8efN�g�����*��f��<@�07L~/����g���.�F���Vg�0�� �?/m��)� Ӭ=�[7��KUz;�>��Zqw�"6t��:�1!��MD �!���,�4��$3$8$��'��G�,.L!8m
�g{'�:!R�+j�}" i4b@Q�JFPH�K~�KBI2f��p��SAkR5�l�kjGO�F�f7w�BL���W��7JG�1�l$����I5DmS9q!�c�[�-o54���,�"ݭS���7zUm���,"��G�X3�i�?�RF�����qO�t3���'fQ,IcWD&0rJ�Nzf�C�s�ݢ�&�4�-�'E�5�o���g��������X0�5���ʸ�g�&y����f�J��%�#Vy=��K�x3�4����*�[����4ϻR$�G�rD�+�F=T�om�<:$-f7u��r��_h���Ց����5���wO�6(� ��b�V�vI5r���K�e���U-!� '�Y k���75�@��$��5A��]���5��Ѐ&��œTi���q�)l}�5E/�����{�E��J0/5�2b1�6�):Z#+Q�1��k-)�!ݥ�/	���U�<����e'�޾7��?tլ�%s�5���|��ز.nTe-�;l�-��4'{�ϲ��b�\k8ɥ����
e�ru�/ٮ�RD�5#R`"�}h��+s�iG��>	�q`'�A��a;QK��y6����Qe����Ͳ���43�[t'�Rf�[e/lQ0��4��۩��,ǝc8Z�v�����]�>�z�G��9���ޤRQZ�Zo�8��A�@4�w��y��Ӵ�$��M;��-���j��`;[C'�sP5�?˼��*����Z�e��1�Ŭ#}��s�Z)/T!��7�i��N.����5)�E��X6�r`�7��J�T{��'rqE!�n�~.��,Yx[&M��/Sw�m�%�Q^��#�7�y�(V&���ѷXi�2�L$�V�3u�G:=�XQi��H��P��^UQF���,*9
V��FO'�5xn6� �ܽ&O)z7��b� �Φ��/*���]]�%��R!P+Mw��2��4���"h���Pz,�fl�6�j{a��,"���mb-�Z���E��,t=���b��7����3қ7�6m?
s��v����1P(�Y��sv�?��ΨI(�3�f:�\�{�����-0#��,޲1֧�K�����R6�oc
�����E(*$;!+/��,m��V
'ZC�~��}҂�h��k9�k��z�(�#��,���w#�iSRl�kܴ-ل]���Q��sZ�R���G��h�n�-�]�B<���'4�޵�Q���ι����F�1g{,t��a,$� r1u�(���H���@=����d�0'���=��4�Ӏ�U����-�Sf-�&3a�νC�Y�g�3�1t�OW�A�!>|�<b��uvl�h�l�4h�r�A	�`��
Z�-�>: A�4! �'	�bI8

E����s�C=S����-�e�d&�n�g7e�[ �j�?Pm�塶��J|+l Q>1��G�!�3�H��=f�1�΀3t����*v=�w��@�5݂�V+n3��G:��c;u��loege�K'���7l5g{��w�g>,oo�7'Cc�6c:�Ϛ��/�C�<XՎ&���o��w���h�V*�hё�׋��0�ë` QQ�.p���<w��g1Q4=�O �I������Q�8q#dI��h�u�?�*`I�� �Ԫy�u+��?��[U���H��l;)��ݸO��Ё�d�|y��m��$:c�n�*#��ѓ��Ye��-+�8`&,X"h� ���"]�w#|V����J>�n����5#!-1=�- ����#oM�[��/����E�%eX'Z��o	�� YLP�[t��}��P/����p�C�۴_d�,y�ڰa&D-�R0�,���,ö�17V"�BkW���4da�8�w1j$�v��h�)ب{e�1���\*��K1Rm�o� ��v�[1��+_q�PAE\h�j�e�S���$1[5��u��*�1����EP#mO��/�;�OaV��D�		Ί���������ur�����&fV *�'��nX�}�n��R,H�V!w��R����k5kK��^���&�1QO]$f_VnI�7\���7}̳���gU�����U�-��eìP��ԝq)*��=XE���V,&�b�48�ic�b��*�@$����.x�SV	�m-��h�`٦2a!1��6W���l�f.�S
�in��e&��hi�ݒ�R��h��-��F���)S@n���}�#��fC��n	�W&��p�����^F4`ʠ_=�h��P���)�n[��;p	"n$���epX�"PA8Xcu�9F=p)�7,�,�s��FOg1HN/CۿC�묩a6ϤY;�MѨ}$���m������*!nP�Y��3�����TPi�o�.x'fP,an�5��X[~@l�<Y��c�yp�H)|h�6Pn�&�"5�SGD��p�7�c�&������GUP-�Y��Gu�����k	��<��7�=�CU�`4�R�����r#_P����x?�L�����?�Y�e�������-�P#�Jc���o3�b�=@ 79�������J5�n���=�Ar��t�Os`?��p
\p�5@��%�$k9��ʞ��I�� ι�x�a�t����|��H�T�7�6���&P7�YXd�]��;-���B��?��q�t-6�j��;���8�p���h���ڵ����N$gqz���rP�q}�<�5��3[&��Q7�u$�>sZ90eycR�����l�wKn��~8����E�t���=M�5Mzu��~�!X�6͝���'��s��X�c�I��/�3��5��sauu�d�/�{����\��T��^a �t4���Wj��Q���n�#5D +CsP�#�ړn�l��Z�5�t�Y:n��A��o�(u-m,	��b o �vP�2Y�h�'b!-5�ѯ`.��1�r��+r
j��S�� G:�k]�Ȩ��w�c��>���N��r3,��G�欛�J~`!w�ZW �~5�#ᮤ��g�/r��.�"��(�&����52�t�#,e�r~��7w���3� �A9�S�vN�`*�CR��]"��eQw���P�x<�C8X5�&z�S�-Z}.Qf!�P
[ �+"�a5�-o�����4EP�=]�Λhv�e,���($�"�'���ݿ�Ф�����4|&�Z+Q�)�/Y�/.$[�΁"e�GZ�'**p���j�7�9s" ����uf�t���(f���P�7Py6��{Q~P,(d�k�'�.2[g��<p����v��+���)uA�}�f�f*�l�(�1O��J�)�tX&_S��1�#�h5h��C�q�7p�7QTw"30��174
/a(`�׮�Efx��Qm�$�1����������P���K�Q�
�U?N憖Pp��A�� ]s9�����fQ���5?���*�m����sY �13�}�eF'�u����O��+��46}Z/P�ܼl?/͢��0�杧RY�ӫ�0��q'�)�ZiQ�ܴİX�ic���� 0�7���*f�\�0��ge/΍�4p`�a��غ�DN���3O'+���!���d��V�w&���E��x�L@�P"�Ip���9��:���4͵U�N�Z]�m�,h��9a�B�=��t��I��yѮtW�a>.��G�3C,�6ү �k�j�k�����-���n�C�ҷ!��/ep���7Q+�^�g�6��-#A�U�
έ`ƍm��& �r�H�dGb)?gE��!�H5�Th'Pr�5�R��D�!M�lu�1���4(�����o�e�O]5Q�s��!ݠ��1��`��k�Mf��|�o'9�j0����<g.�a�;5�i�¡���!��m�ap=�?�qn���Z�Z�3u����Nn�7�7�/�!�D���*����� M'(�Ϧ�?���hЯ1�k0�hgJ.Prr?�:��z��!٦��4Ĩ�d���<�
l|�7���[ �-����a���*�ݭ-�S�l�|Q�l�Tb�T���L3��O���~L�k�CeՒBG���A�9� B�W���R��?O�11�0n�{�t�1(�2m'���,v&7�)>�`�K�yMKb6��R�0�v4��� w�0=͒������/@C��(�p!`5q,��e�|� �h�%بp5wM��cezt��Szו/�Yi7��D��Aa<)i�z3�#��_�j3έv#��_�!P1|ֱ����A�x=V'�ro�K�[g1���w�����]�[qre�({fv]�h�#¼�#qe(�wmU��;e`$�MmkS��T�4��O"�Vo!���*Ͷ���^�c��u�q䝁%�Q8[1�߅Z)C.&P#�	QT� ��T
S����&�u��/��1�ᲄ�Q��<ej�n�Ѥ]|d]9���_���.΂�|r`��� X5P<�nTMR� u��	�z����G�XQ_�Ec�n9rY{��H3_�����l �Qy�0Q3_�C5n|r��{�t�H�Ng��p` q�m��#�Q,�&��!�����J���qr P � ��l��������@��ڝ"Q+��:�*�p��ʦ"MH7
�����=.=Z�;���3O��w̔$z�,~)��/u'	5�lR�<�.N��,��1��k�;	r�̢�O'�1��)�:����fv�p>M�����/��_�1��9 �.7��P�Ǆm�Վ�}x
][�?ܽ-�]M�
|(nAݚ)I�Po7�)�X(N��v;"���͏�^e���h-�9`�e�ڬ{!Qp�-Z�,�X?��,���ersv7�ՖF ������E_�P4�=aIX��
j��K'�N�OҤ1��F��Q��<$ީ
�K1�Θ�X�.�TI7-~ͽ �975o�7?�s3�-ZT���_�Ê-��eX�fg!���w�n��V�<K��u̦^1�"�fԘ?\P �-���bx�qY���zۭ�*�4E���f�Y&a]�Y EY�fW'�Ξ�gM�N'T��lK�-����]�@������ ���YS������a4a�ʎ\m~�E^zk${�~b�n����+,�v7�e=rQ3F���
̿�K��$����7���qو!�d�1�l����^��������3�׵�� ����m�i.�D �Q<��ė�)-',OAN�P,�|q�!$�
KIn5l���,�5���_^�P�����j�!���<�s��>��_�M9��Hn���Cu��M$��gP/�/G_����M�1�: �3��M�o ��6�w�T_P��7���14�0��,F1rs?����Q��x�H�-D_߾�m_[�J�k~5�l�3��Ͱ�4A�aYh5)�ـ&�o��}�9{���A��\nH�u��!�9�P�\�� TI.���p2��ַ$��M9��'���K6Ɨte�Ųߏ���e$��B�Q
\�UҜ�`.u&���t���lw�yȥ3 밫���[Qf���l��8=h4�]kb;�YTv�/�W��[ x=ŉ��,�$P#yՁ6r��9fH�޴�+Jh���{���R�!c9,ltuv�[��;�e�Ι����lo5!,m�w����&h�S�Z�k�>��f�^!3T�z 0GR��ɮ�j��5�3�OM?��6a��Q2��'1Μ[�C̷v�n�"7�S�\�2�e)��f7!Ω���R:n�bo�Q&K,�u��ST��&�R� {W�bk!�K��M�G)��5�٧r�aj��E s���-M)#���.-l�P:�g~���R�4�q�',j�0c�e�.v'Ie3���y,~Έ��Ԛ��&aGr\v��Cǋ��Q�(�m�Ğa֡ �:�]���rg9{�s�~ܝ��,i��p3Q��8��?� �%��s9��3�g$Ѥ#��68����k;e��'X��ac�0y�7��Z
X	q{)^���N|�����pm1L�SZ&=�{�|�n�'�8�p�ue-�Al������Z Yf�Qz=��n���G,�QR0|��(�/Z�v��4{�����6�\�o��^��Xᘁۃ�!3M�6���5� O3j�;A�g#Pa$��F��i�cQ���ib}o������`�%�xݷ6��[�'dͳŅsˁ�4E�j1]�sdw�0������'�W7C��"t��uY�bw0�j���G�Θ����!��������z��{��A&)̰ɞ��=���l�+���v�:�Q3P�w� _X)�/)[۴�,�C��8�u�Vg ��>����)�:�搷���s�D1�UK�IuQu:�Wo�s�- sCd���&+�"/w
�����.7������g��S�Lx�J�-� m�T��ΰ�R=�.��~= ��i2ί����w�{�ܝ)��Z1���{9ܗ�n1A�}���B_C�5Cu (��lĠ���,���5駺I�+Fl�(�1@��z�{B�\r��^�#�r�[�� M�D�t�G������թT�����&Q�<D�|�?��M�Qip�7�gr�de3(��
�^V�lM6Mt�D�T�פᛊ�dN�$΋���[j�rLF�,�uW1��L�-�bu,*��C�O�=�ͳ�z�&�xGM9�5��Vl�;C���<e~���U��V }wf�*��r&uo����Mi��J��|
P�O�6l�g�
C2�>��g�����74�\�A/��+i��Z'lOͩ�`�}|��q�a+�47�,,zr{����*L��Ǖ�X��6v-���+k�`�w��}�ݵXї�-d�m�-���U��?=MM����쁹���k ���u����<�_5|������5$
۟!�hсy�h;�pQ�}��¾m=nѿ�J�
���ۤ�*��X�Hٶ�5;.�����D/M����c6E�C���=�j���	4��{*��n��O�Hvj#�%_kp�)]������.�v��p#��$
�p�XV8�j��6 `pT��O�v�[���"5,QmPR
%WЩ�!.����Ѓ�5��L�^������k��/lR�Bv�.��Zk��]]�44Y�wm�{�}�P��Ѳ�2��T��UI��7jM�j"
��B�2���Y(�Q6lR6Fn����1��Pz����
0� G��1dN�02�l����O=�6�M�O @V՛V�LvL�O�2�4l�1cd1N��~���T�Z�A�{�{��"�&�Ǣ�ԕ���]���*,u��F�f04��
9���O/|X�9�MEn֎�aM�$�`�.3+>���C��]e	�I�f�u#]eqaM�ou�W�z����J�!ͨ{�����>n�"�Q�k������yh�W��jɣ^k���|P8��OJ-2��0��U��o+��YS�Gw9�i�CF8��-&�fC0P��r�:�����-�{�8A��Gga1X*;=!��ce[EP���,>߶,aͺ�TQ�I}_ܥΌ���4yy��#M~����tu�Ol���M��A �YCe��#˥���� ���8���$P�[�u>��������k� ��9e���q9��fC��36���E�O!
Y{	L�ʗ1���(��,<�m
�{Ɨ�X��E!3C�/���
˕�y�[m�l��c-�lۏoHq��(��b{O�W�<���ajY��P<�/a�oC�-g��f���m�����������h@٤�S� �|X�LB�i"�ۈ&a�x��J��6���t#���{1�u�7=T�4�Æ?��<N=��������՟,p��Pgsv���8�9�yA�l��o�51����/�b��~��!�S"U땭�`�܀�$7 ��6���.�I�N/^@хE�r�-�x�^��eR��d	��\P[x��`�I�[/<v��WF=��tGA'��WG
�#�v�:ӹ|E�P��8⽑"/�2o���cv넴*Dg�jW�v��g����-��PI�lr��	d���D/ـ4��Z=�y+�s�G3�i�i�m���q`{`�O�
�S�o����l#���{�Z(�9?�z*��\�o��'��f����p!'�f"��(���*j��1s*�����}2Vs�;�M�m7D�?OS��M��<m5q��4�~L=��s�AF�)�]jʧY�	�u��ϰ4~el8_�43J�\@� {���](c˽b� �9A �)�`f�������v����[��bJϣLҔ�qi�5[N������Qj[<�lrUg��5�+��o鐨�ů(����m�Pm�R��TfA�L���f�U��h�F1�����5D�q��zE�hq��4GPR�.خ!�3�ZVf����P�v����Ek�
PK
�/��b|�~>?XͩJgx!/pw���Cm-�rCX��&B/"��6)P
����R��5�[��z��&�B�P�[���^�Ғ�'[I�؎�c[4!k|�1�Ӽ�,$5�X'�{Y�}<oi�Ѿ2e=���5[��u��{͒�>=[K9�������!B�g�l�li%u�0r�"_��կ�EXX4�Zc1���╷���
�
&�®;���NJ(4�&� � a�i�gr5C�Ė�=�f��٭ h��̑� �-4�s<�4�zvV����e��e�|�� ��FE��uѷ���ơ��s����β-u��d�݉�b$�}y���S�Y���6P]��3$��u����:ե���o,�]��ӹeQb�A-���k��b� �=��ap�z"�`�$N�D��z0 u4c�G�I�&ί��E��C�y"8�z�&l'�Q)�-E��� ��`ѧ��e�pҬ� �f�y�of���ծh���5���jb�Y�`*W00�̭݄�\���H,���V���%��Q-<t �7uk}�����G,�\yc�t��T�n�'�`�
/�=�7j.��tueK�z�Jn��7� tr��n3��G_�n5�3��B^�hw0.Kg��iȦ��a��u1b�S$�77el4--7�x��s�v�t����|�R-N�u�A���mQ�RBm��A�0Hw���6k�D�_]��g1i�4�o�3�<XP
�A��(�xj��-}��ư��w�d�	�(�0V�h��g���������I�q��G1����\oz��{c�a	�)Q/1����&Py?6mL�=;ڕI3N��fk{o��ozj��k}7�����x�:�ǒ
�`Q*3"�0��{�C!1�Wx�X�wɸ����d��q���Ȃ����Ɲ/U[�-v�����1w[`;����]��#��2�eU�)J�0�����Uu�.�9M���#]�t�k�48(�	�	IB�j/�`IR��
e�م�1�N�{aD�08�1�Xu����r�n&�eE����"��4����1LX�1i�e`��D/nX/;�a���1X�15;�mm��i�]T/ X/3�Z�UG��4o�==�e� 4�X�(5�� ��Y���|����l����ÀAa(UYu�`�њ��(�lY]Z��<���dirPETky ��cm�
��|S�d�
_.��R,���X��e��t�7/�"�ƥj��~���J��b�945�͚��c��D(�3�j���~�����0���A�b#��ڼ���2�(4*E)uuy>�['["~!����˨?2-vy�!Q�)����3-�$U�Cҡ,�Ξ�$z�,E�5I��M~�`��&��rju��r�՛||���.�gs�������.T0�A�tį���GA��sX_P�yh� �k���a�k	�w�Sh��*�o�u#gȠ-��(�/&�6,/5P,�w��f�+��.g�����G����4�
��pr�,^u��AԘ)s<�m���պSL)##�i���K�f|`y�Q�n{��x���$O9��L�@`u�<-45�+�1��$Mu�苀��x�\��*�qr�o!*��G�g4!�c���`���P�'*�����C��e�}-@f[���i�F�:6� ���y�l�F�)X�:��C��K�L�p��ka��--4�z��l�Moխm�om��J�#�܀�n���h�͘QX�zQ?�a&k3ÛGp��Ӡoe��=���;aP	oEr����0���3���oi�uӻ�y�Y� �af
c2�����G��ca�'E��q�ix�d��T:�&x5����AϭѾԎ.��i����5����إ�V��a)��R��n�������L2e/.e�/ja��B<umh�?[T�-A�cma��͝�=��km�tK,P x1^��$=`��a�)Ԭ�-�<�з��@]4-&��Q:p�������
�xDO�4�	t����v�dz���z����
���yq����~
á��yG�H��o���#Q��VD~���"�c�D���YջOt
-�p,�P���A.�\�6����'�=s�z�}���rK�(~7���k��)P᩠
اj�(�6��,�"�� $���'������L�h:1�Ē2��j�3��5��[7Nӭo�s!^nA&�yDRO��6�[�Zȶ��'9D���Cf{��-Q͵��C�5�<�X�#�'�$�QB�������.=�k�&����'h��P��{ҍ�$^`�G���`9_ �m=�A*?#ͮL��#
���*����`�,*���<#	�1�P��1��P���[L�6��d�-3~�����	l	�3e������ |�,[��U3e�,Z��� `�Ch��(`���$���!��$�p���;�� �no���
����Bm+�-A�B���c-j�����l QL�T(Ql�,U ��>|n��U�#�
le�d�E7#�Oe,��;5�G�ck�V�D�ӈpV!2��5���-�}����
z|`���3���AY�;ɶ �Ϡ�&1met5o���Pu�KUJ9#�-2!MեRͧ,�7�{:셆R�\
�5���m:��S''?5��Z�wiv�n��^���#�Qo�4:��drrpxE[�Qm�Z��7o !"ء.k��ⷤeP�w8�L͏��oU���UR�f3Q�U�s͏MC(;l�<�O�ivBYd��1'2�I7��!�7 DpѸ/�:q1�HA?+5 e=Ϯ�M�~5<��6��7(Q)�pL�6�GL�/?�5�R\���!�7�.GC�vt��/[l�Q������ ���.[>P��$�Q?m^!}!�4�S��P<rT�%�c�ur�C� �îx)��vl�C�YV7ۮ��.�5'|�@�M7.���H�j��s�'x��7G<�ٗ�����|At.+(4)-.�g/,5-}L# m!"9M�2� �����.A��r�j5=�#��
T*�.s��,a���u�+X�z�3?!V�q-i9�a�MyAY��ZO���8o4�SdsM:s�)|-�gYnu��ZL���2�A7��\�k�UVm��eV���Q��n�M�u��W�T$��T�)�)Y��dcH�j���S�Qe�pf�8�$1QkO/M�������8Qal�"`�� h���1;^G=����
�ۘva,07{��a8a@�񰺴�Y��<������jg�_~��K���0�*�M��h*�Y�l��50�0 ���&-5���4)9���w���w�Z��!�8v�]��ړ�f1�^�omZ����/3����{2��x`a;B=����u'1�����M���11����P5�'Ӓ�[��9A-D'©���>c���81��Ս�l$g���j谢�R��c$b�����>�@$�[�!�$b;��.�늃K�>�f	W��,�>-R��P��c�M��*�=Qml���or�-*��a��|��P�x'+,`���|5/7���c��/R�0794=Mi�p�zr�΄�MmI�wS*�I1�GY>]0�Y,<F�j ��X;��t����7�a@#�߾�{ٽČ�Qm��ut͉�y�|>o���,Mq��ۛ�ur�:iv��7�g��xYA��"��Z�)E>Z�P�w(-b'_�T(�2�4c�o�O'pv��6a#>���0���$��e<Q)٨��u	��];LB]�\��h.��n�x�xN�t1�}�w���P������MYR���Y핎 aa�2��m�Ym�:�����>�l��˦��/��L()[aBxR)��	���Y�)��(X93��߀�7��8�Pj碡��YǮhE?�k	ӆ4�'w1�ɲh�9�aZ fi��2gG��<O��3[�����uF	y��!��)�+#�zA	A��>��RN:)uaN�ql�@m����Qo)�g� <0M������&y"Jm$�U �<���/���@1��A;r�vn�o@L0��+�X�7�����x}S�\o��vw�f� �-�0`���@00$�� ^��#�Z�z��)%@v��t�/5��A�0�`�nj�П�3�w�g�`1�w,;,�ru�`cA�unt4)im�b�Y�wA�h�c�.{���;��<�n��Ae��CU7}�f�)��1'~�|�^���}�s�'������3�y�0{�z��͇�|���\d�r`G��zclj��j�,�1�GZE9rQ>'�=9�1���,d�73�o��r�i���x�$���O���5����ǌ���uwwrp����Q8n��Z���<�l@7�Ά��R|��w��Z-;�m�c��l95v*.�[5���_�5���k/c�	s|#l�\
�ў��@޹�s�f*�x�H�J*�us���a3��Y��|�������v���}�
[]�|�����	�ͽ��-4�#i�	�$?:�>61�sl�\��i������8���\,]�_�sP���{�r�vp�
��&�3���|Mg�^�i�q�	m����l�m���ylh0�K��k�\�<b�?�RF�h��4�>�����r���Ԣ݀CP��f�5�5}�z��&�?V(�e���)
�co��d�+���JӀ�M!k HG�n�fM<(}���NBN	m��yņ5w�q�6i7���3i���QǍ���@c���0��1�}�G�-@ĵ!v=}���Y�K��F;aA�$W.�E�m2��e��-PIfsO'ӕ~����QG~߽u���zC�
b?l�mj5��l�[V�
h��2�� C��F|-�>��e��)`�aPP.����lӄ�5&[>,���c.���or�?�O(���܎ �M�u-�|ȅ?͡�u����!zsvߖq��F{��N.͛s�L�o�6�T�MEv1�)$8�2�����˾�G�*vz�G�G�srV�gPZT���1M 9A_u�3Q�Mlm���5u07P!���[��[�>cF�qgE�Ig�1�!Y0�N굍����I�T([ׅ�rQqdS5�h�jCs�pl�o������-c5)6e15�+���+�h-��cij��  Q)��͟��X7�pZ�rp��ҡd�nca���ŭO#=A=#9-	&�#UA w6��A��N��m��U�9Po-R�Q=���S9Ж(�����Ѕ��{G����.���tn-	R[,' M$�禬NؤD�|�a5��A�}`P=�ZU�}_��Rw�c��Qޏ}Ѕw�o7+����P/�\��W���ۿYr1!����b"+5>Y2�-=���$P4rc���mU$�k����u�O <\�5��5��*�s苖@!MB�-���	��gY=PaZ7Q.u��-1�Z�!B[k���n�Ͳzo�$�O"|�gۋ$�fn�(�E?u���[��!
|h=�Ak9-BA5]�]U��H��#[UnA)c1�Ǟ�xk�Q5���x�3���8���,mi��N9�م��7�7)	����8R���Jn�A�@�1R(�5!��R�l����P�$7q��ͱ#GE	�kɽ1-�mکX���D�,�F�ެSS��`�P" s� �S>��k#!�%���`f#�W����=�)Q�����΁���me���i�u1��������s1CUc�tD<)rO�Gm#�]�Vܵ�ru7twO��9�?c�z��렰�ف6�a��[M@qJl;de�����7=��S!t�)��o\��p�Kd�Jk�{�{�d�!�xَ�"m!5|�t[gD*�1��a)dM� =Zh*�3�3K�o913��Q�B|�Me?�U�a�7�7,�*����ݖ����Dk�<�]u
i��]�wR3<g]cS���4�|�1�
�g��O*��C�d��crޘ��]0 �MqM�{�L�~sOl5�M�j �Zr@��Y�'r�xnp\��q�t���a�_f�W1�g$J��4�O�?66�1���5�6p�A�=�OlbE��PG�r-��(Q�.>}v0�I����"��
Q	��lw�M�Tb6�>
3{�#-M'����+��>lfǘC�x~``���?���ħ11���Z-,1��Ib|g���m5���qn�MrT.��\7�|�Ԥ�nvnP���$4A!�͠Ȧ�p?Ee�+��\��557W5�U+��dtFͫ��D`Q0	v�+6r�7/�'P�Z!�b
�>p���(�8�}u�r)`q�S 
d��,�s�\t��y�5�u�Q�n����V��k>�#�o3���ll��7E� d���_� Q>O�r��w �$=k.��vr��đ���t	�o�<��ux��7)MCJU|�A�Uy�[9�D(��1c�l��e�"}�}��9��E�o(�6a=Fh21�GeP��ͬc�e	��<�0HvX=�@�t <�e���PQ�^�o��L{� �d,"�G<�tm��	c�6?��h�c���BbT)c	[�)S3?{���b[7	W�.�pJu4	@�|��8O��O��J�#��F��f�a;٬�e+�U9�}lZ.Hk��w!��u�۩L��T	��E"�Vk6%��1����7eȔW��*��}�uu$��,�2��½���w�A�b9t*|�1j�=�pw��u�6�l�>��:@�P$O&to��@N�`�z�Xe���JGP�h� X�IG�f�1{�.� 5Z_r.3�Q����~sXx��f���o��.B)L�]M���;�M�#�ZŰ�֥�+�
�+n�G;��p�2�w��t3iS�8���j�'�!&f����hS/�V��������GPP�=�C,}mP�XK��b�~���	�em>~A��U"�tWh����;�x�#�4U�7u}fy��h�a���rP.2���ke(�q�#0y]��`�F"�6*��͍~�DQ[��� '�y�땱7.M�^� �!�Su#�x �P"��+ �ϫ	�'$Pb�Ztu�@e�uO)����>��7�]����#��s�]��5 HQ��o�d�J$�g�F{���w8�t�c�����1g�7�7���t��� �cP�v۲�7�ݮ���d�r��SL8�zI�u'7Qi�a]4��<u�4�g�g�;�^T$��-)bT�!$Gi<�3�x�`Ũ��5Q�� ��������J�\�wu��N�:kq֡tS�i�Y�srkLxO��>sw;���~����!��|Q}罥ow��^Ao���[��d�m�z�o��@(��!1x5��.���o��ɂe(��#񻦱�2/tvdmrgo�<Y,�� `��7#S /P-=T�:P<OڒO�4�Kcћ��N�Ƭ��z�]���`R���4yht/Fi�3g�\�)�a�6'Q��������`"��w��Ψ5P��o�dO��7��u�[����6έ�����-P7�eQ.O����sxdJ��`߯'}{�w�cM�˱wg7���5?n(h�5���δc�]q��խ⼧ eΏ�փZ1mX=s��#R7Q`+=W /
S��"3kQ�w4$��5a6Se�0�e=�e��d-a�Pࡊ�ƍ�����.���h�ѭႼҽ�E���Xi1r �A�`-a�s��͊j���t�+9(9���n���"�F�݈�Or�,s�/7�� �Q ��Α�<��}�m���X����-��7�C�i��*�6͎$!lI��N�}[�et�3�iQm��V��v��	Q�)Q�'9MEr�6K���w���YL�}Xv�/�P���XL6P�� �����P��Ē6%� �~Y-;u��ї�V�HD!PL��>̀-<�ԡ��iy���R�����#.n{�q�#�(���#	�n�^��彬y�9�s��SK�9̂V�����Y0-�1�V�/p�"a���~�=�Ηm"�1�f=��ο"a�	��=��w�"� �6=1\B�4W�*��P/�l1�q/��W/1�/�a�W(�1v=/e5�W���/߻a�XWt�y1��/_mzW`�W1��/i�dW�0�1�0
�?�rkn��.1-=�|po�6�1��ae/3�m� ��(mC-�n#�c�G'����Q>��
Q5t��{j�x�'ނ��g�>�³ C� ��Z���b�j�Q�q�a�������^���1�~)]A9X+YkY��M�Y�)@"$"'Pӈo��]���uSU��Gw9Y�N�@)3\�4i*����$���rQG�)�[/��V '�7���$�m�36���?$[7a߲V`t��T��d�E��$
��Pn*�|�� l'R�.w9R6�׊iwVF��s>���Z�f��SQ(�fP�	7���Q��47֬��U���]���|@�ǲSK~��٠��0zj	�o�*�r�����e�P���cr��1f�v�mo�"�ei�?%'d]!��l�Pʨ n�5h��(�\�\8�[����4@T������r���]1�%.������".6
��U76���r�v6̈́.�o��w���cQ0��*�'��e�n�SK�\=����'�� zj�/�nk.�/���:�
iG�&5����j�@C-8)N�%���!QEt/$Pi��+�Z��Cto���|u!�����Z٤��>ڣ�!?�&���\\�^�l�a,P4��NV�R�#Δ�l��~�g�է�z
�aO5��A ӑ7�l�eQ��{���=Ni�5�-X��- �l0*� ��[��ĕ�uw����zt��*��Wqɑ�^Oe�
����M�����MB�/��H/;�<�j1�ʛ��P+j�*l�w��eWu��6��ne�1�?���7$sM��Z0����{�)�THwX�U���$o�ՠ�������� p"��[�T����>���,5�c��q��^�|�V����tI�Afs3��껶fi?�)qLqho�	3Q*2n+��(P�C�@9M��}��WwS&Q������7�xQY�+r �ő�N�Y#�(����㥆m�Z����<�Mu�1O3�VFq#utQ'��Gΐ����z4� K���=J)&u��{I�Q�o6���>�]mU>V�O�E0=�>Y�cQp#Q�)�缳���U�5�l�*�I�c n�:�1�԰w$�n9G)b�1x�[��eE�Q����[sW�iS�lU
kI�����/�!r�'��1��#y�	�<Q*�]~v-��H�-P<I�s,QwM}r��M*���&1Qxl�o���{Ԓނ�*��B�e�z��a��H  v�?ɼ71�VXqw��1�hM5p�mfΈq���umY[N�ph���,X�����Lt˷�������Pp$��$ �Yw6_�w�ϼCwK�y�L��>�`�N10�	6�u��m���`)i�]�{��Y�[�6Xܟ�f집|�<�,��rv����2y�$�63"O�A�.�79F<	=�9`#�S�@7͋Ùɨke��c��t�9��o���
P����H����s
��!��˟�E S� hA=�f/�[��b���!�pB����>D{(�PH�^�F��)�� f9`��*O]e����koa&���7vr'7�0X�*;]J~�<S�
ŧ#jv��Ҫ=n=�i�8�bU���?�.�pL!rL8���I��)	>�CU��E��Q��~�H� 1Z�qZS�s�-7�]�F/c4���z�w����j��r�Lx�֮��V���$��8'9�o���Y�lw���|t��EDn��1VY��'�� ��${��Qz�ʁ |�,0�|w�n����?�ƅ�)���fd��Du�9�0�_��t�VE��B0��ԍ&nY6ӧ}0t�aE�/uFY�� ���8�QP���C������I�٠ #�)������Qg5_�� p�$h�b��"g3Zz����n���ms}:��g��k�P˦h5O<n��2QEˬ|)�e�t���/z�����/Fr�{mr;�E��\Q����P�2��wz+fyO1�qt�7}�*�A'���Gn�A��An�U�(�"W/�R9i�33'QŤ��k*��ڸ1����c�����n��(�=�P��x���e��Qm�+uM�o"����2�6͟+�R��u�5PS	�r{9�"��x �eI-�m��.�y9O	O�뽐�̷)ɔz�a�1�ue�b.�*�(G���z�/P�-asɵC�7�8�r�ϦP|-`�U����CX,��NA�7��G���6Q�[-O�'�t5���-�!=Q?km���\ya89
{�[���2���ɰ+���F�$�'.�o�-��@Q�1�[�}O�ku����9��6ם�;c��w#L�s����5iQ։-�K���n�H( �d�51�g>��Lʧ���\l�o����a�5�)M��
�U�;��t��3٘T���;1{xd��[44�a�)�r��m�`!��ZA���y��X4k��Qia�- 	�1yy��{z�{!�����7 ��* 7�۬: lqx�B�69�P��}Z9����,۲'HmrEަ�P*B4/5�)��Hĩ	�x7O'�k�d7 bP?��9��`�$�N���'ڴ9��$�d�+�-[Őep!�Nz�62d�T��|X��Um��w�u�7pm��=9��wvP=,m�K�Q��X�_lg|�#Ջ��A8�-͞��a�ͩe����31aŮe��QL,��?	��8t�dD,�'�N�4`��uL`���(Lg?�Sxf��.`�v(J'��DaVQ�u��9�v�*�m�4] �p7�w��d<#J'�{��y�@���1�����o�5:1�)L:k�����up�����2��&��Z�X-'O0�e�*� �ɀ�/{5W01gZ��i Ƅoůgjws�1��V�|<���qkll�����E���Q-�a�ۖ�]��{����.e�@�/m�g*�F��1X)�g}x�R�$ 0��h��A&�JZ�N5M�<=L1s�L�B�O9�7�Go9��q�Qp YF�j篵7&El�̸5�'�-�m;P6T'M��-Ѻ^M�y8/.�]�e$�
x-��-U!��tx�QZ��-j����S[G��=���e�g�n("�T��^ D��}I�9]�;I�t�խ�4�Y��r�c�x*2��0�z�E�7ފ*����#����nuur�d,�Re��A���3�u� 53��kcC�^n�@^,(��	nzg�pf�A(�i_��A���# �ߤ�M�ҭ�$�P\�l�
Q=���8�c�n�dZ�f�[���3^XM�cɳ���!����
-�f��O���l���`�j�c�����՟���B;�C�z4ǹJ����pѩ����m�}mQ)nL�������D؇^d�OV�x5`p���/�Hd���s��naֱ����e1O5|�R�|��z��E��g�~�XVN\�-��g��-�s���}��63n�%�5Oe�+��͓k��VMd޹Y!�'�����6�a"���׻0P9P��,��F}�,�س�L���n��7X�����y�A��:�P��y�5���~����*ykr�]��P4�0�`h6U�	P �w]��ߚ�_n�篝v<M�f��K��)����eN��4�n)�J���X~	'W��&�L�sɰ{{��z7!�"�b�aK�9A�[k/M�ir��\tl�n�� \�r2��7*	��[2��s�8�w�#i���W$[d��:-nQ���L�,k��(�Y����"[S!|��Ț{�׷9	�`,Ec�z[���}�z�q-	���#��$f�X���í=�v�&�8j�u�ﺮGP$��(�Ae[u�RX-Vno�"�p��X��V:��)�nzJ�ިU�Y
hY��O&��5��6��9��}�F�S�\09�-ѣ9oձh�l�"��vnzbc��"ew��$e��(�'P2麱�4΂��V�
�����/!P>�8�e/�a5�&S�0<΢Fw�^a�� ���("�7=5-Rtu�R�Bx�( �<[��	,�7�>d��üQl���������a�Q?�7��[�*Ob�b���1���t���ː�
�8]���.X���p$lP	Mb"w�N�b�����`{�`+ˆ�6P��
s��Q}Vh3��?�H/(*:��S~H	��N^�_?Y*Z��Md�K�Pnj��5��Q�ku���f|Y�N����``Y�!Jɔ��s��ّ����:s����~w�lz��!�s��ɐ�*�6��Mb��3�t{�b#�ifc��?���c�67$�c�d��|q35����ķ7R����5�b���R�m���8��7C���E�)!f#b�{@-΃@u=޻63!w�=���ӹ ��3~�;0vﷂ�{�����.Pe��|�X�]��!JA�����r��,P+s[�]��u b$�0{�Łt����+���]#�? 1>�� ��(".autvY�Gΐ��f�]�#�9�Pz��1.�����f��k���+}є��E�s���v$Mԥ)�{q�G���Dv���x�t[����Z��W�"X45^���z��ҽ���ǭ��7s$�V1rZ�u�u� i�"
�n�6�^Ԕ����IE�FU�-<:	&1)E=>z�&KEF��1])��u�d $EN9]�58�m��~���٠��u]��k�57�/\#��"u
���|!�?W��񀮚Q"t&��K�(1�W���J36��?ᷟ��6m׳;x5�[=*��9&�_�8S b��;��8�L=�s]&�U��H�o#�-���h�7y'��)�����v��]�&�u1�[u�\��}������#F�E���A)�'���"��[�I�<e��k@!)}�#1t��.���.�Ũc�/s�b�)�5,��I1��{�ǟ�,(yx�=��l�A2�d����UT�3�'�3�/9�H6M�������e0Q>���eO+t�`D5�4��A[��s����`j�P2����^�現Q<Pg�Z�R�Ts��{	�&Z2��K����x�.m�-i'<v���@O
�i,�wo6dnַ#�p��`�lǫ3��4o,Y��|u18�����`5-0��v��J�D`���L
���k�<�ou��������74��\�͛l���g����S1�ru}��A�O�3�grMuGv�c-t�K�-÷^��ղT��v�oP㨮(�/�z�ӯr�퀻��ydQ.�i�̺_�����"g�*9
�	��t@� ��u�2�L��YF�a]�+�U��*�����X�r�� yڊ|J��cٹ��b�~�z�v�۰7v�D_�s��6P�� ��Z`%��J��|n�N�gBh�tĢ"O���<O��u�Qo,�U�h�["�7eH(	�K��д�"l���J&��]�eE��e9�Ѡ��(�Ź��wI��wtm�����I��Q�<4Uk����N=P�g�1\ue�U���!M� ۗՑ-�f�OTά��0X�s��&"�jq��N�p5��.�n[���?u��m~{�1��{7�ҍjz�hy`$�^�3t1��3�,���+�O��~�7���AN�@�ɮ�@h�lR-�1�v)=�2x���[L<��Yl,���`��;�
7�}t�`+
W
v36�1hj!d!P/��t&���61[Ǽ���{5h���d�=�5Qjw�wl|1D��Y���{I��#��<�,�di�<�����H���g5R����nԭ�xɳ�<��P�Hs5I��3��Z�~m�Z���L	;ig���j��?%>��'� ���l"k!�.����[��(� ��-�գoq�!&yQ`aɘhIX��J��`�c������.�?��#g2	[d� ��33��OG"uRC`Yf;Y��w!+m�z���xMu ~p�j������ظ�{Cx�w����qe� �� 1�o��m#-A)�<Q)Y�f]M�U�IAim<A)}�fqu�!��a�eA<)�f	��A9=�¥<!,5ȴ��7+9o��1��9�&59���9q݅�&r;Uv#w��9�"4�h=��W�9�-4u�W�@�#Uŕ�$�)$�.�.qe��1���(�c4Rw+1��5�1a��i*�ai������$��jfn+AI+`wkOi(K#pv;�)PJv@.+das@ulE=ji`�psq+0ba<����%��K�m"@DUcW|��Mn)d&JF�=�b�QuW�1�VM3��'I�QWF�\Kd�)3 �v)?�
g/4=D��$l�g�Ar�L�@Iu�'��҄fMD�qJ*hPIQ�g\�ir%�$i��Sc�@F�Iv�|�O���0�/fPW��qM)�Wl�	}(`;��Y�������Z�1H�h��B�w�`��q�GNfJPG[�$����1��;F'�Qi�(�`ϗ�iٴ�h�A�s�cL-kDuHi\��K���p_�iaJwP=ֽ��i�G��U\Jtiq�Y�w�2�f{c0���Vs�ϼ��l�&Yd�Y�G@P�Vo�tP6�۱MW��7�t!j��`2_�;C 3`�A�UV��[��u��SNKA3�	/�`^=!�W=�i��UCL������Nw��@�ao��M5t�#!�S5�iT_�iYs�a��:$uJA�\��XfN��$�Ӄk�}� h'pK�1�37��Ӝ��$\n��(�>oed��B�pp7f�S50`]��瀞�\6Q���`Cl7hw��$��;���:QaI<l�H k|.5��4�w��qn]p�U�7��vO14�	l��\V�cF��UgZ|H�p�)zgqJ���u���S�ԧ�O�f�Bu�m��MAl0䅐:3�[��(�b��i�'�U��QC�=��/L_�af1˗�5��|vk�SM�TK,&6�m�p�9y���Um;���"}{'>mm�?�E�E��MToet�!)0T	qA	ǐMR�~6R�!֪wC�xd��f:\�6n�\gn(�8g9��m�4Yl��]O�/OG�sJ�!��e�KR.����f��,g���;��n'�FP�ϸ���3���lE�v���7�$jC�V�bUG��TP��(�tC��m8:�a�wB	P�g�aa��+C�U���J*�l{Hawa5�B�#) ����8@�}�s5jQ�AtS��mJ���yG�y �s�7Po�27�OJc|�d+��8�L�>�h�f/67/jU�5�;q� �oz/PHAt}��gs�a~;idϴ�Z6� 8c�64f��/|cVءo$ve:!t;D��+Ҭ�y^�1LF�Y�1�Y��m�!+��Y�R}Uo[��A"]4��f7	3U��a̾1D��ho�0��_�9�G$vvP�jMBa\)7��k�d1$΍}o0�I��4!3-L�4�[�z��&M]�,�б�9� '!p�9�1M�2.M��}���)9�$���^$}U �w<�&6�o4ˮ����&��C�� IA 1� ��dD� ;��@,G	A�u|i<}bV�g)�hoꖩwXH�J�s��m`ϛ=auW�@i<Fo�I3^������;�1G$�Y�1))�'!G�bE7-�����&W�-X.$�zd{]�a�}1sf|U� V�!ai�55)�Py�?b�qY���2!�D�=����]y�	y%^ I})� �g,,�!�X�ԁ����oR.r�:d��Q�|�{(Δ�1I5��i�A�-PW�9u&IvA��HD�;�{U�.��0Bam4�7�} q\U��<e�`?+yo��W�hL�F�m���=}�	�F,<qJgG�]M��,g��y��<G-y���o�)�%Em`ilu)ҴHUI]��aAf�#B�%}L�����/�`w�Wjk�\��n�C�vq70d�?LH� fmhxM̓�-�D%w@C�&alvu�d|��/=[�'��V{)c$����`9�KW6-���-Ke1� n)�,�#�1!�=���ߨ�q�'=�&�5��<�� z�1=I�-,�N'�$¹ή7v�7$iC#�jm���E�!]���6���Ua�+�4M$��UM4mW/om`�=�|')���o�s�$"���=�]1�e�=m4<Em?�]a�W��4V��7Q�mP��S-&aR�]7�mu�٤M7!
� a�#��7-�a�,-Ŵ�ݠ�m�g5! �j�7e=},!�}�,=TM*�][f�׽:��ٝ������*��[- �=*�[f�m:�}�M��]�ܽ*�[f���:���͢��5-#�=���=��A
ed�^`A��yw�5�uS]�eW)���Q9G��q�"-U��S*5����M�!_M�e*5٭��լ"Ue���!�-ɪ-�&U���y�9m�f����	���9i\ �[U}ݧ��'�-��5��UDo5G"MU1���*5iK1f�\]E�dM!"�W�o2u�i�l�g�M�,9�P^���` ��}c�'�5,n��}�R$^�5�U��5V49���u�������5t�Ͽ�35M�(eɾ�0-��5���#wC5���+�5辪�/`�Tatm���5�)�b"����5�)�5�5]�h�u��5$�.�is�bU!@���L4V��7rˁ�v�n��X<3HK�SױkA��U�{M\;AP��g�0��QV�� nD��J��A\~Ie�r�BM�@w��US�+K� ��R~�ǝn���=C�9M�]�T��V�A9n�����m�P�M$|�q�}CDtBhnH�7-�D�@�A�Jg�@iKMR�@5=J~��F���x�/�M�Ǆ�M��U�	}�Q�G�Bc�!hvcq'�+�,��zwR��� !@z<�޾'O��a�QA,�i	��,ѴE1}'�*����g5��9�5��-�5G!!�	�E�}"$�,+5!45�)ĭ8��eNp���5Yo���Mo}�]`�q�=�-aej��!}�^xY��!c	;t�1"A�<��ϑa��!V��,��1!2i�.�����"A�91{ �}�oA"\m75݌k}S	,K�A�9�So �ceo5[��\E�,Y5���oAA'�=��0!AQឝ$��/|]9��a�w��ZI�eio��y�kA y�i-�t��rA�A$���;$���e�=Q%/)E�\ma~�]}ۃs�=�����=bA���W�	$4�׵�:Ѳ��U[�im=�$8,�=)5��&��	��\�VQnA�2R�GMr'��!�N	vp�N�4�"]y��-i <9,��d	#�/�-9l�%i,�cI��۟1�ֱ�5TY�J�<<�e|q�d�Y�� -�&=Y�l�D񂹲� �-�!��<MYy�-��q��4�j�7)"�--�l ��}e$��0���=�m9|�ia���l	�yvy-aE-ig �5A!�Ex��U,c�v�Ui��5�1#��Q���!�ݘ�5e4]b�#�Q	�Rf����|�AU��l����d�24�a/�`S@�c�	/"?�K�+��EgP��9�c�x7h39��&+-M۵1qfu����cpa;��F$�6dGJPQ��1xs�c1u�(�w@HZ=��lu�=(�~�`!2�q!� ���|9{rom/��vԠ@Qm"�AI_=�.$R�zoDb/1j2�	=XcYuW��/�Q�2=�>,�#?}31���2���V��F@]�sA��y�B8+�m,�iSa�Kr1}8dF[UQVq��$��W@TP��arI���a񦢰A	��#A�]��K5=rh	��y�@$�Ѿ AHD]iL���G�Y#�ai�+юW�~��ӽ7��g��m=�ټ�m��q�1�k PHG@W1d����FWLnUБ8=��(
v�A@je,b�vY�m1w'��"x�Ԡq/
j1;l{�	��7�f�lIu/PU�\�}���l��1d�t�a�Q�5�G��+qJ�4�64��L�a�w���_e�dߴ���z�13}��4p;u�v��+'j�GI���m!B�i-^�ls׀W��e,T嗥���A�ɲed�"�ՀW��%E)ő�CB��=-1�c���u��� 5D�V�zILS�*'��67-�U�(�|�}�WV�Ue,�*w�9�O!=�f/H�Q�4i�-+�1�jG��2P�lK��LAP������E7g�lȾu�v PU]���r}v���~���t�7j��ChQ1Ww\�.��1�6PA�,=q�/��Wgk-�w'�ZF���v�/=!M94pK���d	#ouu�Ѹ�_�wR��w��w@M�	�r�0�WU�`��ռ9�,��50୙����/G]�� r��IAg��<�iݾf�mԁ}�aHdoI�~\��mw'������M=/� �gM�h`Bٟ}xS�-6C�����eM��!���v�K��p�1�35wi9�Z�3�7مf��<�,&�Rq��G���c�w��Q*0-q��j/D�M�o���5'�~�Nb/A 4��!n5�r�����gv����u�+gPC#�vU����տUhB�y,!�2�U?9c�4�ws�SMP��RK��� ��Z��R	�P���3u m=YY�CxP�g}���Q��/��� �v��i�lc�K}�շa��>9Aq�,NBg�&/�/ґE��[��w�oA�/��,/Q���# '8�h�f��ՔrU)�Lk��j�] E)�bߖ7��{1U?�o��M�A��	�a��U���<��*I@��?�;1��]�U1��paL �;�P�G
��-����?�3g�:]�7j[���l�D�v;�Io;,Ӎ&�9d��c�u��R��a�r�WA��7[G3F@�5�=���B]P�N�a�a��H����]�����Η�	�ǵn��S� ,O�Vna�;�B`�+��6��lC�_ʗ
/B�f�H4��� ��lVc�r9�_k�H:O�yw�]hL�gV���{@;��N��WR܈�a7S�3"��g7`GÑr=j���CJ�<���k�VH2��ULCZ��sk����`��7Z��PLH�S+��+ef�9A1j/A�R/K��P9?�9���Iys eb�]���DZކ�}�M�DQo�^>ML;��k��_���3��I6����/'mU�?Fa���A��rB�C�);�^c���'��t:����/I\Q@=
9O���9�IK�����T9|!P/�U��1���a�W��o����|9i~WA�	�n`�:S�}}���g	�
�}�J��\:kER�rQP��N�ٌq�33��`��\�:@uC5�~R�4���0=��<2r(�jm�7�HCĒ�Qot/hۑ��,���ڌ���Z�v���~�;v~DCi���K�օ��pR���:�tW�C�j��<�S'�����/��nF�I<���.d��o����p`	��V}�R�񠝂�wJ1�Bk01%�f<| ��_5�K��I\K�EG�Mo�Ԋ pbR�I4�h�d�R�d;Z�h�ǁ�d�{��b�k�hw:` r;laAV�ک�����A	NcB�tH;�o�I��@0�kL�L7b>˅���SM���w �M�V�+���g�o/$
5w��Ջ�V�h�)H����ِ����K�ڗ^��ه>��\���(���@�f��,3A�H��"vjzn`5udilRs���Ա���i��P��g���-��v�m�@�7��9y�B7��V�<9��P�V�`v���>�\DYt��w	2H���9�<��kۏ��wjRA=��o�k1@�X�R�в�?�`OC�U�r�s��?"���	W��i!H�T)�S��GRf���t)�C�Jlg�w	�3�zWIV�9V	3s��s�kFf8�xC���ġ_F?5e3-Ī��c5̶4'���4)W�-4.Ƴ-�u�I1N3lT��"2�e�e��9Ѧ5u$J�df��5N&B�l]�S]Wz�=i<!���U9o���1=1)�i74a�s��ݘ�A�1-41$[S]g'�a/!$���$w&3q]&�a9�;e15�]!.	f!be��e	 ��� AmE�9y��#�<#)��:d1mQU�Um"���-5[��a-	�u�"� u,��e�/A	m��	y����g�aE�,� �.].Am)<7�b�A)	i�s.�M](��u�(Aa9'\'1���]a+	q�+)
�m:
�����*�}XD*��t��,1���}K0)��05m�y<]5)�L�m�-1�54�En	E4�����	p�	�7|Aw7<7�r�T���6yM�I�6��K�t=��U���O7E�u�m���1�)��1.I�1��a�2�u50�U<0)��~qe1m�3�mQ��3Auo��u1��\y8gy23i]i�=Ao�m�h��]g=�Y<%2~�L��Ĉb�n�c#�\�u��M!7-�v�ͭ�d,g�fF�C'`,acb��/ 1!e�M����!�9��a�ِCA�	�J�I����������!�-�Aq�G��-Aa,�m���!i�Y�a���]�,��!Q��,e �D,�$'��M�mW���l!	�m
}ZI�,1M�1&��Am)L�}eh)m�q�)�M�Y�,��3q���a�)V=4l1��l���mr'B�!)�F�otq@o�&�q)I&�anY��n-I!��5�D�i��i�i��1�q0�h�@hI=!	���#�m�m]#Akk-T�k#��	'!��ew�?uc�Yž]<viI ���6Ո��y�I�1ץ� ���Yaq���'��m�U�<&>[�7�;f!J� f�� K��ʹ��#�7)�T)"��a�*�-�ʹA�,�7���T'�����ܛj "�J\�A!�%��I�-o�F89,Yi�%|u�1���ݴ)2=W�M� @)�Y$(,�j�L0)��t�m�\�)'��ZQ��*Z�&IK,*!��)}c��i,�g�`)Ckt�7A;fk#Atxf��tA"Iw��m�\w)-��qQ��*q�,�p�5)-�p</>�7;f.G1(,!��c)�;�a���;�(�2m���<+>W��m�\)*��Q�!,�5�5�2m�m�<4>�7M;f7Axf��A6Ie��m�\e)1��dQ��*d�0�g�5=/�g<3>f�2�\f)2��aQ�U*a�=�`���`<`c��c�c?�b�a!f.�bA>Im��m\m)9��lQ�a*l�8�o�E�o;`i�Yi�c:�h�a���h��H2m���H<>5�L,��~e���Q�5)�5����2m���<>��7q;`�a�/,.)m(�+*a54�7761m0�32a=<�?7>9m8�;:a�7aE �Y�,�a�ݭ1#�C	Am,EmY���a�խ)"�c!Aa,ymY���a�-��9-�E�,Y���a�խ5,�c�Ai,Um���9�����{-x�\-����4�
��!���,U��K-��,5!���zE�m
�^���Q,u�]7�,��Yr��{�$Q+-���TU�-4=R@]b*,�1���݁5@2��df5T{��n�5��-5j5�#C�'MUT�5w7^35���-�_�+�|51^5�^5~�!a�'��н)��'Ocr]5���75Ỿ�5�5� !5M^�UI�bN$�cګ�,*�"��!a*լ�:�}ڨa�t$����!X
Wa�غ�lW#�it-�S���K�y�Z�9�&A`q7bi#3@flH�+Ek\ڪ�hUFaWV�,C��W3(��;+UAk;ڮ�apV�U�qr��5�NAN[�II�i� ѽ/��յ��}�C8Uk(ھ���
vTKi�n�\j<5}B
\itB���\�IM��1#��,Mأ90/e)�u���7$PUq�A�AH�;Vba����D��7pB5<�_�cfk��m��d��j����s��I����?�H�u��j/��!�i	+~���#�o�^���yO	5�tݗMjl�`�v�@1,�w��G�$Xy�С,!�޿̮���=ѝ!$d3�)GX �pc�	-H������-C�<�u_��!771����(�$��a9���-8.��d��S��}��+y̘�a	��{�y5�k@hc�-B�	��Fxg2&�y�!MI���j��'Y9o9=4N�gl����ew8��lMe��U�kZP�^�gE�" T�)E��i���d|Tx� �X�^5m���� ����!�i<)!�m�sf�n���i�Ee��+���z�a�it)颈:��I#8���	�����1u�PrE)y\�1�vE��=�έ�5�w�IT�`K�oo��o�A̰-9g�M�D\�mA`AQaM�Y�Wq;)�S_������P��Kmv��qqw�:w�{��������?w`�.u�
���1�wrbYMEr1:��q�v	�˓�D�iU��4�l�m���`5�rB!Ii1P����L*�Q��Y\��9��wS�U���I�G���H+��:M�WAkIU/G��rBw�Yw�Q;?��1Qvs��'�G�;�}�9\M�GvN�-g�0��U� '05v.o٣�u��$ِ�;A���Y����Ӊ�W�	L�k=� ]��1���?�k�yAxo����������5��g\V�'�G8{��/@!N�Q8�AcR�}�E�y�~��	W�g9�HG@	�Q{� 1ͱ�ߺa6<�[�?�������V�p�xi��Om�M\鲷�u�iAw���!;c�C-��a�=qaK����<Sт/�)����^�Q�a7;���	�a�Dh� aWU�;�n����4��u?\p�a+�$��7���������7}V1�M�CB ��Ayq����� ]����WMD�_��oO���-��D�{�g�S)ʰ;L��m��jO���Owg��9�)�r�73�M�F�!����屋��i�C@w�G�0�A 7�al���L�	�,Q�Si���P�sq�K���]��rU�*��0Qev\}�q�$w����A�G�o]\gx�3�O�R�M��ۉqL/M�2{Umb���wU�5�j�9�C8y�G�#=UEI��u���B'g�Ui���m̀<2�����-z��aL��{n�i�9�_��3�U kV�	�	�=M����
�A1a{L\/�M�@W)-`�Aκk���,$<�1�_,E75A�rAa�d8� �W�;vG�MdG�@Y	�?��� �BQg�����+m5Ո�J�$ao���GkGq��	���qm�׌AVg�q�g�e+�U	T�TY�@�'�k�3i�jLG]A�{�J����AL�G�	~E[���,���\��Yn���K�g獭;Lk}���{3����Rh�3.q{��A|RLi����t@_�B	�d�3S�������W�i�;�����`MaD�;�:.a�x�K�뵶����1d[��-B��H��f�	IO�@��p��� ���b/u6W�G�Dkut�ї��LH�7R�wyё�L�	;ji-�N���)}	͗PT'�j����bm�m��vn��_w��Cc�jL;�L1g�QwwDS��H�hdI-�G�VcͰ.�<�8M՜?�b͆:�d��vc�y�{4�g�v���ͷi3�k9x�ǅь[�=��/Ri�N��AG(\�H+�L�As|K~n�����],UY�1鈷�u�?��4z�)\I�=A�_Wԕ@v�cz۝<` u u�	���WM�`Am��GH��.�;}���Ӱ?��w�gmP7��Uz_a�Q��?���VOG�9t�n�у_�j�m	�>�]�oX�K3\���2�Mq<�巇��WA���1��	o��o���#�ӑ�O�o��AO���im��\���74W[W�Qb3�t�� ;g-u�=�U�H�M$P3��ͷ��A�܇�j[��[7N�Qp�ś-�k�s~7��]�C�W�aL�)��x<�dwSMv�,{�tX��R�C����tC]O��3��/w�3��c}�v�ד�Cs����C�	����k�5AK����m��"��n���u{�3-��
�-�$��5�#$-9~�D8M��;���:��������������ĺºӺ٢#4bB��o�u�������(6�=��ڢ��e�a�m�i�u�51�=�9����	��d�o�u�s�{�M�Jܳ܁ܝ�����������֫qk��b*hj��)Q�S`]�_�Y�[�[�9ec�k8v�|;E��:���������������κԺۢibwB������������$C�����Ď̒Ԙ���'WQbSv]D_CYH[X[�[�9����8���;ߢ'*bFBN���!(��S�����OT�5i�W�Q�9�8a�k;z��:����������κ׺ܝ9"�+80�>; �
:�f�l�J��������պӢdmjbsBx�A�N�W�\¥¢«²�������������������""�b�B�����*1���'qC\Z����~]k�����&5��lw�ę���wWCQ�S�������,WxQTS�]�t8��������������sW�Q�"`���b�B����������޶t�z�]�[����;���Ս����2ڦ""��G�X׉l�L953�	8�7gj/u�r�{�@�I�V�_���9��2�%����������� )�6�?���Y
[[[ahn��'��
j%*flo#I�R���������������������������������"!-b)L��>����e�a�m�iL�q�}�y�E�A�I�U�Q�}[Y[�[�[�[�[�[�[�h�������������������ź��ͺɷ�j���+!l-���*�1j=�9�*���	�����e�a�m�i�u�q�}�y�E�A�M�I�U�Q�]�Y�������������l��ܝ����������������������������������!�-�Ey5�1�=�9�����O�'*G�a�m�u�q�}�y�E�A�M�I�U�Q�]�Y�������������k�����Lq�������A��������������-�)�5�1�=�9����	�����E�a�m�i�u�q�}�y��[A[M[I[U[Q[][�[�[�[�[�[�[�h�������������������j)��ł+������������"!-b)B5�1�=����	����e�a�m�u�q�}�y�E�M�I�U�Q�]�Yֱֵֹֽ֥֭֡֩օց֍։֑֕֝֙������������������������������ޤ!�-�)�5�1�=�9����	�����e�a�m�i�u�q�}�y�E�A�M�I�U�Q�]�YܥܡܭܩܵQ�مفٍىٕٝٙ�������闃[�[�[�x�������~�WQ-S)]5_1Y=[9[[[[	[m�[�'e�a�m�u�q�}�y�E�A�M�U�Q�]�Y���*�����������������������������������dg�����ޤ!�-�)�5�1�=�9����	�D����e�a�m�i�u�q�}�y�E�A�M�U�Q�]�Yܥܡܭ��Q�ܱܹܽ܅܁܍܉ܕܑܝܙQ����������	�:ź��ͺɺպѺݺٝ9!�-8)�5;1�=:���	����e�a�m�i�u�q�}�y�E�A�M�I�U�Qj���������������������������������������������+!k-�)�5*1j=�9�d5�	1 "3e�a�m�i�u�q�}�y�E�A�M�U�Q�]�Y¥¡­©µ±½¹���c�ّٕٝ����������������������������������H�jWQ-S)]5_=Y9[[[�'*��m�i�u�q�}�y�E�A�M�I�U�]�Y���D�ܱܹܽ܅܁܍������������� �"�������������"!-b)B5�1�=�9����	�����e�;m�i�u�q�}�y�E�A�M�I�U�Q�]�Y٥١٭٩ٵٱٽٹمفٍىّٕٝٙ����q:��������źͺɺպѺݶ٦{!�-�)�5�Uw[�[�[�[�[�[�[�[��W!Q-S)]5_1Y=[9[[[[	[[[[[eka*Yi�u�q�}�y�E�M�I�U�Q�]�Y���"[��:�		WiLJ��h"��a$Օ4 "HBR�X��������^��*0���	{;F�Lsc6=+�`kJ����]U|�	+#*k�
�*jn�z�ӷ�͒L�����+h�W��]:�:آ"2:b Bd�l�k�mBL�1��_���u*��g�W7Lj�ħ72lc������{����B�����.%��74��f�oS*G�wd/QW�͑�i_�9��Sd3>n�� Y�;��|�wk�mDa�ܢܨܶA�وٚ��	*-��J6�w�*�����ƉaE!$,y���b�B�Ä6;�Մ�����*�;AB��������"2�v�O��9����8���!1?��lɥգѶݹيٞ�����: nt�$Wq�;��^��7M�k��io|TA�M+���x���{"F�+U3�ѱ�0�!+Ofd\�Z�����UYQ�J�!L�D���#W�Q�9�⢯��d�@�HI���Uh�=�>�)K��&Ug{�����wDg$A:�aɧըѻ݊ٛ��������Q[�[�l�_���ע�����'#�/�>@m�'oj�������[�Ei�W�9;�_Y�[�6-c�ޕD\�#9�l���Q��O������)���fg���<��U_~�%�[4������,nOĭ�Kŗ�2�
�c�HɪճѺ�#��:��ȶ�k�kb�$/}�S]on�*������E�dWB{S+�/lg��< �*�$�+Y�, �a�-k�NЂ�t����*�b"�lF+O�CF�#h)�}�+��n�D�#69��qb~�A�����9p�QSL]�_�~�*���oDo\Ie��yc8N ������������?	"�^���m&>G���+8ԛEN�[Ѡ݋�C[�z�&�&0���u�|�Ɉ�:��˶(�%8��U�YL[�[�k�*�������w�TU]k�*y����g8	��O\� ����������+Q{Stnr,��D��ܒ������a�A$n0,_`DKw�{�_	�+"k��o*xlFdߦܒܘ���������1h�
o�-W����[�o�;���LK�hA߳с�����\�n��� "�GbTJ�7�������+՛QST{�*�����"bw@H���%9*�g���La��0i
 Qoj�o�)�Ɯ����sm7+����pĮ̴�M�K	���kY�[�[��*O�����e? W6m>mj*}l�Mc�h�u~�o:[����������ה�[�[�h��,V�dͿ� �aqj�*���&ĕ<��e cdsJ�^i+?k{�VM�ĭA��!2&�bU���97h���7'sC8>8�7O�e�ِ��[�n/(���@	� [���a��k�+	�k��*��,�U�[�nd��y��������������h|�R�
��ǳ���q��'ݏ�Y�@KVԷ D�h�s�xY	
P��������Ч�~L�IK �"G����������?!]+;��@j����D�eFͮ���C@|����Q;³�A�W�;m�!��=�*���z��W�n�?��[k*�o*]jZ�������������͡)B�/ �E% W2QSjoD�����k�u{2�*��+?�

�Jˌ�D��d�_��Ā�-WQ9g�v8�N;T�^1�����	WtQ�9 ��djbxBB�S������k�p�� �D��	� &G]d�h�H���� .D-mQ!��$�6<�,�e}B�Q�s����g}(<��J�PĶ
,ٗdm�ߢ�G���
+�-n*�9���{�:G�P���׺.r7�� ��R�t]_{	NٺY�����>a
��b�r{�2U�5�֋֘��������a� 4 "�]��ե��#m$��-9.�:�M��!r�x	U�| ��������W)Q6Sk�)Dy�:����]��SY3\�K�*�lƦ��y�bk�q�x����FU#|���n�*I����rGl�Rc ��!l2 �D�"�f�^Հю�������m��qalC��W�w[j�,'��%�� ��������6��}�sg6ϧ{�s� �mn�M�Q�]0��
�4=�]+�"O�-9������Y̧��Ų1ո��S�j15 9�o,HV��r$sAGBO[*�B1.';"��7#,�m$�($"'��;&6����+�)#w-?ZT �qB�/$� ��6�|o�7|*� &��+�;�9/'�j3GȻ���'/r�!5XL%:�R�uH+yS�O��-*)'�,�1%6����͂�%�⾨��:�v/s�(�~aٿ�	��&8#&p�/63"s@WLvBKq�P�}�Vn'20�.6+/+	l�F��m<��HА���U��\ֻS=FwJ�Q�%kjildg�/q|�f6`u�a�"FOA�;2(G�C)&:ƹ?�*���示hQe&��]��'�%��MY	R�9%�#��.�4(%r�v�P��Z%��,~�̵R�%)��>���%ӭ��� �%X}5VO]�T;0�����{�!�GY4��T���
��"1 ��发ho%���s�["�I���b�O�$���,�U�h']W�6�&d�4����%̥�^��щ\��*�TE��6%@��	�$�%�G�4��ђ�1���N-�`�%���Z �+W!�łY,3�+1f���h�"��%5I}�/��%���!U�X%D���.T��%�CGg�������A-�S���B�,B0%�4��%f��c}��P�'�� �1EH��:��5 |�;�٠�4.�>��/�D4*-" 6-���!��������Dȑ�9��b���4{Lt/ZG�#%��ڭ�c�l*�������]%���F`j�*.K���,�8�J�(tE j8Z�q%��	g�.ɨ"�{ړ��Ƴ�Z6lg%f���$s%�����Z%�}��@��%�]���bgM%~Xؐ'$&��]HE%޼z�L��^%UG;atS�%0�Q'�l�%?y��T-%Ӫ�Ő�ͮ%�n�V�m,����"0��&�� s#�%k�b��rc�Y%��� %�ǚeb��H%S���*��Z%[�ܰ%0��1���%�pdUc	[�,��,*�&��y�5\C�K�:���87�� �@TM�'��D`Sχ��Ԭ�7���Ƴ=F�7�;�C;=[�uPGS�>M�id����,*"��!���$x��s/cafR<'SVV2�F)
}UȀ?���Gfuv�A3U�&~��]i	����qa�m(a��O�l��Q�����������1�S.t,e�6'�v���4�(-�/r	�M^���75+B.	�AKH�;9b710�zpf��#r�f.�zD�cq�]F-'Z-ő%���A��0%��H^dj/�%JT�=v�!��M��%l7���@�%v1�!�_��U%H��閊%�}Y��N %B���R� �}�%҈.<��%�U��JyjX�*%w`�0�@�% ��I�$+. 6��٫%_G� �?�9w���i��k}%�^�,s�%M�g`��9����p�	��j%�Ѷ�&:^�&0�ݏu:QHG�6���%9+V�#e�%���T�C%��q�.BY"ݢ\���/�t�%�W٣x��%o+�}Dh�%�A�6�{�$�Hi3�"A�)� �-����86!'�*�..;*�S�y�V�+��ե�[�5%^���f�M�%��K�.�	�Fl�ͺ.'����]!��̺�1�+3)��3�"��g(/C�a>;����%
:��MQ�U9V
I<�#��&��-�qѺiuQ�_MtD�K��HYV��C�[	ɇ�Q	Pj+�\�FK��/��~O���m�ox� �}�>u�Lo?a��]��/��V$	N����ck���o�s/̇��`Ԓ�t�����Ise��/�r��)��l�DU�d<hK��ی�P��t;��
 1/�މtU@\[B7�� T~>jZ�I�w�VP��C�A	f` qdlk�z;YR����a�ffih��Ck���C/h+�	/)kOb�m`�-jc2U�j���Ju�:���=�i^S(pgo`1�oj>/skWbkJ�j9u���>MT�����F���8��9jww�/���o�Jm�u����}�?�9� �GHpK�.3/���fm:/�K�Q�[tk�u<u�t�fp��?���j�q	@r�EY��qy/yv [�wf��atpp��i	B�_�vsg��j�sa�h�bd���G1�͵�PZa�hi`O��j�#�e��q��'o��rnz��v�,
�a�/�]m�����JHM+����dFʰA`D��{Pɧ�C.H?G>tJ�a���!�$���G��==I�����C�Ҋ4'�{LY".E�m$�`�"�Y#-s� @'g39�E� G��[s 035j9�o?0�Vc����qX��F�SQA�\{�$3�ϸ>�-=D˂"ݻ���i�\p�%Qy� ��"I��^c��_�%T#m07@�x"�t����1%]���.��+xm��:�/v�e�+�6H%b�mi%W���[�a%J����Ʊ9���%���W9�%�&K��F^%]a���ޡ$���"�֧!+����P�e��`(�~�e���m<��&||��9	+.n\R�:o+!7E5�g�7�T9%3��^��/��O
})$y��Z�]�vٟS,���OkLjHQԩOS}G3L�ȵ!U%/�]gY�%��ur��~%i�ׁ�n$���L����:%�V�򖼀%�°ڎ�X%Fت�Mvuh&$���E��[l%"	�'��_��'��&��r�.�%U</��z"�eL�RJ�9����+F��Ӥ�����gy9�v��&#���u%����ÖS%i;r�F�%4u��f
6�y(&b>����v/_�,)hѡ���AO�]6%C�/Y:�n�%^G�ܛ�*�}�%/�M0�%=
��Py��&�D�!�ݩ�C%i����r�%�	]1xgk�Z=�'ҳ�9��$���m�;A���Z�o����o��]�|=��.x(D��/?. *��;�)!����y}�:��� �cY��p����%B�:�3΀�%Rb���$��\�%��K/`�Q#$�F��m|4Uwz%�I(H������*��7#EA��%��p&�[B%��a*�=_
$��yV�@�Ȝ%��cT�+}�%��H[1Qx�%��bF�;����A��d.۪�$g:t�ϲ�$���%                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                             ]� k�     ��                 P�  �             y� �                     KERNEL32.dll   CreateFileA   ExitProcess COMCTL32.dll   InitCommonControls                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                      7%(�r# �l rA     �    `�tX�    XC   �8�ua�5�    X% ���3�f�Zf��4f9u�P<л�D  ��g9t-   �ڋ���� ǹZ� ��
���W �Z�E PQ�   �    X-&   ��  � ���Ha�  �B��H��u����BOw-
�@ ��_/�B!�H�Q��i��l�Z-
�@ �b�Ó=/W�@Pe�y��D��l�Z-
�@ ��_/�B!`�t$$�|$(����F�G�   �u�F�s��u�F�sO3��u�F���   �u�F���u�F���u�F���u�F��tW+��_�G�   뛸   �u�F���u�F�r�+û   u(�   �u�F���u�F�r�V��+��^�O���H���F��   �u�F���u�F�r�= }  s=   rAV��+��^������w��V��+��^������F3���t����V��+��^�   �����+|$(�|$a� �?O �8�2R����5��+���G�`�����`
u�Ժ�K����Themi8daF��3��B��S�}d�\#�Restar�Aqpz.|x�
�Zj��)"�B������"�����~�4q�X��.�����`p�]� �2����a%�	#��+��� I�t���i���pD$q>�& jE�`�)h�t�zP�
%K�
��
��W�U�
�����Z��@3�	��E�@��}���t $����C�c�6�at&��F��|��IDҍE��]ǅDJP�
 �ÈA�����]u�'(��d�u�����[��7Tx���K;u���GF$JbF��B�a����_��E��M����F�>�@��6�4�}�>�m��L��J�e�����(3ۊ0���r
�
9w���&"ag
f����
��Ar
Fw$�!]����}1r���vv�d�&��v���;U
��x�����88�*p��5 �GIu��q"wj�����v���6��Qe�o�w;�&���Y�� _6>��,�v��� ����Uy�v|ɣ]R���g��a�����b��`4�9N[0vhQ=|�v;aFlu	.��H��e��W����7�GS��@)�q������+�w"4���3u ��?wv
g�03A쉌����@�E��`Pb� R�M%����ͫZ�V��
^�����D؊���#�(C�ykR�!Zr�h�t�E�!BR��NM�i ��]�5�7��Z��ȹ��j1�M �b���Î��\���s�&����<,H�.9�a�O�v.w�X���<oJ� `b��՚��qF1*@��${��+tH0�Yg��0�S,�
��w��Q>a�� �IJ�3��|������oQY������ t����#D��{� ��r�z� �uگRo,���P y(hn�b*R�T1����{�6��1hD�@ i�eR���]H�ࠇ1�;:09��& �u!\)n���a"� �<�:�C)��~�3�1H�����
�� ��_���\U)�t�<@I룴����6xC0h��&�P� ;��zJ#>�Cs!���jG嘤��(��K*࣐>���:�x�σ +g������ ����|ؐ��
�̰�x^� +�FE�rBj�2���Zo��̤����^��适�
���D�|X� �2�P~����0t�H7�
�9�S PO?�(�C���H
.�z��2Q��@�Xy�)��� ��~�gs%��ԧ��~j Q8E�
G
�k�0�+x�`�i]d�<��z��@�� H�0�@r(�n �p�ݡ�� 3��O��>��� P���a�i��� �V�<�?�>�@�<�đ�Fr,� "1���-H�+v��b7N�p�D��#���!\@ � ґv�ZX��p���� ��e�ߜQ��GDq��D�ì��AVC�,�)����{�� ^�y2���� �d5��찐GS�M�� Px��@B�X1 �[4C��9s� Kf�J�� 䥘��?5U	�
�T	I$��0� =��(���U|� *C���5v�r&y���uê���`����XG��l�P
ԯ����b�x �y���֭B�i�|�P`��̐� C�ڥ�x~"�+\Ӱ��IM �?�ہ` �i@"]du��k�#I�j �}cK�X���QM�P���e ��UK�� �Q�Y��������g�V0������w4ǅ`�L��{@Pj7 -�q�Z�W�0��){�Q��	�9{3�j��լ��>Ł�(�� GA�@�$����@x� �������4�(&��xd2��� �H��e1�^Q�� <�(96�J���>[	4�|I�\�Fw)����(m9��@te�����L@��� ��:�7@����֙��;��RJ{<��.6��������	��@�@26K���h�R�T��C�� E*��kCycZ)z{'��A�T��p����Ǣ$��C4qb�@y#�[��w�/�7�c�Q�)��)������D�d\М��ƈ������s�w�r+�Ix)�S� ԿI�<W�oL�$����AD(P�, lA`Iz�u���;���(�� K��`�(X��W?N�m���GR{�@$@<�]Ϡ�IU� �(�jJ����lW��������]e�b���t�+$���/��&j��&LF�R"�x��ꧬ���)�a��� �0f�� 0g*��X��A��Zs� n~(��w�)!�G�[�'�,���)y����b;D�ԭ�����i\����� [�0o��G ��;��-���A@��饴U��	>� {�0����@���)���������D"���7�Q�W%0�T�O.�@0�S:\��y ��J;�A��$���`	:��G�)��L���pbߢ��{������i �^!gT$L�?'�yq����� �g5�����XT\�w,4�|���Í>����[$fR`|���"�+���P����Tz�P_(��� �c�$ɢ$��l����r#�Sӫ�̸e^�ي�hh�n��)Fp�� �cbO�@� �9&M�ȋ�9��Ȝ!E��[1�A���t��yX����D��f�w)�%��I$�j� �Ł	�N� B��B$b�R� ��'V�z� ����Mi0 ��{���`	�e'�8 �;= P�O�֮��D�|@@�z`���:C *��&9� �Ϗ-)��⣔X�	�V��<���M@1��8�G�|��8��>g��l��"����@V L��ƪC�<�p䁩�r ���z���&q.|@�Sm' ��N�� ��F��9���~����g*xN|���@qy m"���d� 8��s��8P� �@�{`�I��G0 �=|���E Πa�����sr� (����oX�<b���֜C�DBvrF��N"� ��,$Lq �O<���+����{��@a���A�&��`̿L��%r��#�q�}�XXh���8�����`w���3�����>t�j�C�0D��Js�| �&;�@���0�J� v�u˜xKc�8L�ؖ����j)���vK��]�����	![�P��H�A�ˌ@NC����6o0�myJ�W���GY	�n �@������Q�����q���UsEP��f��N1ՐA�K�M�H�	x%�W�rܪ��Lv/3���YG`\�s`�H�3a-H�4H�J�t��AI$��ds@v�(�#(� �K���e7q�J2�)d�Pxb��c��U_@����Q��0*��d�X�Y(.��!��~�!6����vzIPu���2�#����n
9OtﴰS��PD��@P�0����v���O�H�ڞ<Qq�`�Ȯ��㊡�H�L�">�����	�+�ܛ����|�qQ� �A����F���h$�����Z. C!m# Bt�M[�	��4�}E�"${ ���/ ���f� H�ظ��t� �B=l�L�s
z�F�ȁ�DV�u�����3�m��A���X]�$���yK�h(�G���2IX�KС1�q��uКpIx��\��DZZ@��oy	9�q� d��1��t\4���1V<���i�Y��.��U J�4�T��:vj����t�q��4 '�uy��,Ht�����Vʨ�)s@Á3ɭ��Ő���T�a�T{���okƚ�v q��A�=�=�f.��E�p <s��a���u��B� �H�[7��0&����M���P�c|8@e��>lL��`�`�.�x�w#K� 0AD�� =0�F@�C. {T���O��q�� ��-U_8�0v@;.�AI��r_� ���c֮|����i`[�= D��&.�3@ �/gq_�����#U����Dhk$]���ZԦ|�����b+�>v� �2-��C�@S�<d� (ꮁ��	� �Uc`��&��>J�@ jiR@�� (ۻw��#� �,`Wf�>:|1 BJ�D�U i^�<K�]�&�m8)�uؚ/muX�p�(� w����iP [+��8��= 324�Cej;L߀`�OԸ|����&M�<�2��046�@EgsM F�f��ỳ��Y  '�8v�0C �3��:g_ �M�e�y,�s��~>h� >.uT�Hu� ީ-۳*���P �7D���/� 2@�>qj� �`�X�m� x�+V # �54��0� ��JhrN� X�(��.� �,��_ ! ��3�@2� I>�Mfk`� d�c��w��
��i@=��14�3F��B8�� X���^ø
�_sv4U��U�f�_�p�^���סt蠇Us�+�D�	�tDj�l�,�2�	mi��}I���v�,��xB�Z�������
T� `|�H��� ��Y�>�]0C�xN:���E^G�bW+��� (����F��Ԁ� 'WrGy�� ����`�����.T��� I6�`�J�ؤ! �A6�}=�������w�������h���@#�%� `X�(`�AK��dP��lF�y��Ǜ
p� 퐆�ZJ��L��&�pfK��` ��{�UȨ�s �O� Ŏ�(x��قpw@����E��\R YF�;n��Qì���N����n����3pR�HQ�t�.�Ey�����A[@�rf����w�\c�!��Ky<�s ��O�t���j�� }o&�U�Bp�t�0V�1)�� ��;��@ L�уwl��{�F������NJ�����\$�!��N�{<���㭗@�[W�yKؾ)T ���BH �#�UJ��E Y��Hu��	�t�c� !+�	do7SPt)�� ��w�^�-� �I�����`	q��x8���`�l�$>#4�(�Ϗ�"̙����<M@�L?�H��v��x�Z�F%�p�t��M��f���J8V��@ՌX�%��H�A�$�܀tF�	s��8B���\P�L�9 ���eEa�H`����Ј�o2kL�!�ɗ�!%xh�8���OC�rc0�0�T�M�lEB�n0\�x"o�*ZV� %�� ���� #�<��n�},�P<���@,a�=��1��uk��;�	�8t��H�G�0�w E��$���j ��0ӂq�݈ �����S8 ܇�h���q�$|)(�t����T����\� 4ɛg�9#P�,0%�z�Lŀ�\�%��t0��b4*1�S���	� �J�2�$�����	�t��!1�	wd�T�X�0�vț��i��I�0�N��F�"� ��N��Z	�SB���a ���&?��(�����W������@msUt,����0��? ���w�П. ��f}�W]uF�������H���C6�F0"� �;6K�u- H��i��1�|�ڗ	���/zP?O�w�lcj����ap@����(�`���f��.N� �ɩ��>0������ޮ;q�_>���Q&�wLAs��R�tD�$C.� V�|[�� U�D��h��;u0.�I�|�I(Ȑ�HE[Vs��		�t��0�	�)- ,�CG~�#��Ο��τs .�	· V���Iw5lf�qh��d�`�!���^OS�)�E܃o���1��,E��7���Zd��� ?��֖�H[¡Z�wa���Xu�$.�s�ﮨ� �R'�k��\C�#��NE��b� ��N�@�(=��.k� ����ݥ��cx�񥰢,Q�t��7�+�8f���ٰ�����HMD�ȯ� �}�l=4@
谊��!AvI0� A�^�Rq�QY�2��t�����ND��Ć@��N�р<Ø�p�w��F��{��&��U\(M�Ӏ(���b Ɍ��K vѫ�.�nl	>"�xd(�P͠���:i|b�E�����rt�� 	K���{5 �[XST�3<�f�u��{�%��h� ���SQ��X�"��g����}���������D�0P���}�ꓰ�d���	�tLǈ�-�	�vR���݄��\�����!�ґ���XY��p�� �M?r��l]`��**��?$��Kԙ�L�j��� 0-1�E@e? #8 ��#z�C9��8��oV���F;����_A�ۮD�3���ŀ�u��`�p�׉J�2������׌D^�ܮ�B#�k��T_�F�.�te�G��g�&��I�A��_� ��w�m�����|��yX��[����} �,��In~;� ���p0�9���(ຒ� ]mF�@n��&��‥NK��X�� NIt3Jpb=L�`�����Q�[�<�S�\0M� ��Թ6@��pT�|��k��� �*/���S�ΐ���46�l ���I��E�r@�0�\D�t�]�I@�����H=쀔�$l �`�cZgj���ͅ@��i���ӌ�0��K�P���^�V�u�_aJ��K`�]�G�����d�W4 ˠ�����z� P��:M���F�z6�He���>6������o0u�K�x�<�.ܤ^F� q��$b���f���\�$�Y�����$DPH��})W ��_�����*[V'1pt&O��A�T\�,�!(���	�t�� X,�	N4�� �l�E��p�(jxX�"�:[M@- ����1�0Ƹ�A���ߊ �EGh ��gA�i��u�B�0J6�h����B6Λ� ��
�t������@.��L�H�QL�y�L��������?��t0������?\Y@�=��7� >8e@_+A� �l-T؇ɽ\P9` ��So� �j����(D'{;�ŕ)�%��CN�.�#Zi	qI���(�а��4MN�UJ�\M *8��=�\�[u@�=h�<���?T* �a����3S�����L8�;�:̰�l�DČE6�@8�=6�%
�Acu��v=�Kl�6k���<�� �ŹU-��Rװ�u���|���|��~���4 Is?�V�O� �F��U&~Z\
�ۤ^ׄ��Q-�v (�}����K��[�$�_:
�,�:��<9�`�O<Rq�`��gpD�`�� ����?��&�� �kI��]��rU�pH���D��8�}	�HQ��V��l".�� �i-�G��XE�� �S�� �8�����ЃG�x�|T����x��#�Ѩ����q�PZ�I<=0����߈`��ݮ�}z�Y5� t��	a+{1��)B������D6�C8��<��l�&� �J��ːP���%+s�T^ ��x��'� ��0y*�SL�Ms �)"�t�l$�^�²����x˦���H6�X�ă�@6��!����Z��Md��:V:P#� ��+j�.i0X����� X������@Ȇ�2��-���w
��%�������U���>��ж��Q�`,�j���H�s`e�HR��� ��|�X��Pq��/T�"��F2(��/��B�N ���J�`R���DHPA� ��\��AU��)401��$����d�Dy\_B���,`�ĩ��\��ĝ��(a�8�v%h���]`�'��ʖ���(	�_qQ4�X��7�{Ř�`
b {R������z ��� ��hT�A��,�E � ��V�+u;�F�DB������// #�<��"|{@\��Hy��T[O����+�d���E�qyB9*҉%G~`I�qX�J/H#�g�m�]0\\eW�������^�P|��Q��]���I@��&�O�m r��;��Kw�֘є�~Ĭ�툷��4���xS ���(0��Ξ�E�������*VB)���١�M t�r�d��$d j�Q�-[��(���"�`��D�o����%u��y�	@ka��|�]�ZW ą2� A���m��,���)���(� ���K_Vuc=��L�9o0`K��|�)Ŝ�`]۫ ��1����
Eyr�\ĶC�q�I[S�s� |�.����l�_�dC�t���Ni�Y"p�	��]Ҵ'��8���غ��_�n0p�HL��� |�Sָ#��NG��#����N'���o���xO;;d#� P��Ӧ-�hu0���.�����W��@�kV�v3��B̴�Ҭ�J((� ��xR�v�\�O�$� ��>*�"@�������@���_�0�ޠ�ٺ<t���	�(����XT���Ù&q`����,	��zH ,�Ct,��dA��Z� 1l=H�E�CKhv8@�u���S�d!L3\"�	��%�d4g|�|!s�� q��i9�ѓ�Ӌ(�a�Z��.QL
8��	���V���+PW�_� ���Sz�6:&�r���Q-wIVn��J�L�A��X �� J���K���}�J��d���0a>�I���7�x�PєHIQlt`�����?\?@�ĞUS�aP� Z���%2� ���� �x$Ur�tF^?|����[L����Te��`k6 ��Q.�\y0-��"�1� �/$����r�GH�[ �ϗ\Q��;��z� 3�,ǟx��:R��/�A�*L�1�o �^����ӂ x�������;�����Z��y(����v���c0��3 ��´�f��ӄ��A�,���||��3�6?~�Lo� �v�N\�Á:hN�H�s0!�~���H:L#� ��Z:�K�\o��={��b��MJ�tW�K��[�4�Ceu,�� ���� �ZL�m�%Pj ��V��@ ��K%��`J�(E�F��|C�q�HVtF���i��bp��w������\^F ��V��hT^�I �}��vMؔ�^F��sN��1f�=��85 M��8[�&�,;��(�8�a� ���z��,�J�^F�?�~G�`s����l��!G�8Fp=w��t�\�G�A�)H�����=�� Y%)b��� �"���s�Z|���LȌ��l|$QC;5q�TR�L�p@c m�j�ʱt� 0	��pI�*�0Lo�q$.Rh&��D%U5J� ���t0!>yH�����NI�[�,ط=�N���ph\G ��R� y���m�Tќ��U;k�	Ew		ᨌ3�0r� +Dw��3�z��?S��m������ 0lE�-VtUy<H�rA��'�$�\�(�@����K@P.�7A	�`q!�f�p@D��Ⱥp ��.YCئ9�xO�����h����4�A�n �۰�1����J��Hȥ���} ϔ'-�����( �	n0,�d8g����B��t,ttF]8[����H5X�v�;ݨuT�C��������[�;�#b
�����'�.h@ׯZ����M��1oYI��ͨ+,�sX�J��ɇ����d H���wUzs �)0trB��0��Yv(�@0.����! �E����>���>V�<���<����I伿 R���>�ی��(�y8��D^`��Gz���k3�̠�(�s� �~l^�N��Ƀ�$�ΐ��vt>�a�ٔ =N�2VS��2 ht������h����A�+����!h x0��Es��^Fa �\4�,����@H��.�wВ.��:��D\u�+��`%��{ K΁��Z��Hۈ��B-���T�р$�u� ��by0��D��L�T4�t(p�H/�y �j$*Ld~FZm0X�X�H�$�L\�K������D i�}X�� |���L�i�i"8DR^����nkHa�/�ݗ���U��k~E���L � ��1kJpOE �1�/�h0qK^V˼�s0p$7� a�D�ဩr�H�ݠ�� G��(0-u0�Z?
���%�`�i�tb�P;��V��l/p!`��i D�@��e���(ڡ��0:4�>�"�^��y1p�(��$O ��]͐ @�ߝ�D�������l(����	g��!��DG�ѓ� �zU[j>$�r�wXe��@�L�P��~d^FZ&g�/� �s�ɛ$���g+�!�S�����s	t��R� �}pL�7�z`�(�VM\�#�.� Q7�8�R2�仈P�H,H̝+�,�'�7Q���p����JF����Xx����� �-�_.��J��8�;� hي\� ��Q.�y�M+�(��١��K��*��|�'�����ଚ]qH�t �R����x���-E@��lU V����O�|P;�D@Ay��_D �n�qZ zS3���y(�h� �B:/<�b ����X��T��-���@�ф��+�[y�Y�x�x�%��q,��0H�v(P�Y8y�3	�Tx����A�KL��-8d�_� @� Ŕ� \kq��S��,? �"3T�� ��Sw�vP:(�"�m�l%�t$�I@�N.�	Q���\p���^tx�)����|Fb N9��I�3�(q�Z�!�ٕ�� �q�wH��8�Z��R�s�>9Ҍ0�%r��`�����v��̠�,b�/VH���_�N�R�f�ꂦ�1]t�[�=� k�X��-ìE��\�\as�Qud`; ŬF�nV�E˞��4��q�p��pZ�Ό��ѨK wx[�ZO���CЅp��(`��P��JV����O	��|�E�lmu(�*�`t��� �r���8]�H�9L`~@e5xV�t� �� `�s
P�l@��t�O@}M���O���<��\�3Mp8��\�`�\ϐ/��Y�|HRЁ� �����6?Z��&� ����@�����XZ>�~�5�B��?8��w�;��r��th��m0�8�����s�+����,}H� ��C��>�����$F@����qng��Mu0 Ȧ(UPQ���o��,%�	�v�	���A��p�vL	Џ���X3��"�g�7�A�� �/@�	��d�	�ś�<�x>;�#[���Ԃ� ;8��GTZ"��=cIA�ܟ �t��8���`�ϓx�����:���'X�B�H��t0��(ٞ� h�/�������͢�p"H���up<-��{%ą���ҍ�12/;D#� ������;t�yQ�!�ӂ���W����uv�(���(&���^!s�O�f����/������\����Ƞ9���h���!U�t�O�P/N~>#� �!���s��@ �XBh��J ĥ�v%�4�����"��V4��cC��a�|��$D�8��g`D:�#�v��Ĕ���� ��3S�p �w{�`��i?�\b�Ƀ߂x)�.� �d��dw$�콘L�0���3�Lx�؄������X�� >Y�����_��|�����y �b���Zq'\�^��E>��R���AT;O5K��L�'����>+�������L���; ��\|��'9ir�����.
�(�}w=�n~ �f/������X'��.�Hu%E\�cҰ�qp��@�lM����S�C��Ly]`���@�����\�쇌�:�y�\��X�~�HJ��$��`�<�H��Y��0,���� p�4/���! #Y�&9� �%�\�(ح�h���b9pi��vF��š��/4'�z��V�^!s����A��^�!?H �]�P t���_Ԑ��i1 �{�I�( ��HL����lUw�_��%�P������-/�@�W=_ "\ܯ�C{�	%�� �?��%����WV� ,��Ϝ�S�'(�zI���q�l$^�tF�r>����4l��h�ۤP�[��Lȏ�%.�M�]�ar���t�!��V,����|T�H�����ZU*@<)�D����_�G�B�;f%�R�Do���B`��p�0�wd��Z�h?����S!ǧ�-����9��L@׶�_`��.0L�tF� ^z#�� $q���V	��s� ( ���Hzh �Q1h�K���; X�vCV�I<`�E�����:�,K�|�@fC��ɀBw��;��`k��}04�����E@���8�߈�H/ьJ����k*�a|0 �/��`���@+�v-(m�f\�C����[ʌ@���XlP��4��ȫ05y���p(q�yˣ��4S��B �,�!@��� Զ�yK�F��4�ܺ�0�����H���5�ne ��1���;�t[���V��pJ� ��v�N��^ I�2�`lzTw v����c���5�_FӴ��=n:�D�bk���ˍ��2� dw4��J�M�r���`}��1���G@�n���(�E���H�T��40*�~V0TT$�j3��8���#%[@J�|;M��x��G�΂$���<�爄%*��G��#�l���q���c2أ�Y�G]�ZCt��CGE�B���Zth��Q��D��H�Tl�`%tp\�|�Y���Ͱ�`"YqH��X�(�,|� �D"��t���I�P���c ��-�N�M��G�C}�� t�<��"�E��˘�$YNX�kt�DS��G>��l�,u�o���PDK���lS�X��I�ш �H
�`PL��t(�K� n�:M�.�<P`Y��(��v����H����`Y"u�:�r_�E��C5�	aEO���� �H�x �
`1,!	����YxP�G�
!Xg���Hq�����2z���m>�0`~YR��8e PV,�KG����N������Y�r2�.�����j�_�t�GlC�ֱ��HC�(|X�tq��r�T��$cČ7Xf�;��4� ��G�x�B@t�=�`#V���A�{Z}�z�T�*�Y��A�>y�	0��<B���XX��6HW`�]$V�w���u����tKoC`�� Z���H�(4,
W����,�N�G�����,�tj9�4c�Y\��K�C�y�^zp���Y��^�(�,t%"��r� ^��L@�({,tw�8�2SY������G,t�lp�n��`���x�B;:W��PE��B5�*8	��츟b������@��@�@�|�(�K�Hl��s\0h8@�dt�t����C,~�S�Gi�YeH)W `��	$t�*4e�f��|�`�\� P�6�Y�8S�u�#`t(O�`(�h��d�X� ]��<R���e�@,�s�]"�j��Ǔ_N!�ޙL��H(�g�B�u/*���$Yl8�f��,@�TH��0�Y�H3�'�m�A�s l���n��SHk`[{���T�
�G���İ�sl�"�LplN8P�BXt`dCS�����Hek�p~�Qa0��A�Ԟ����2]m�c��D�� �G$�a�>� �~�r�	��<�`F^ [�Z�XO�cY����P�,	u�`��v��P��"[�$N��HM���Hdo4P4܎�����c�Yx��:� �f�,l�$15؅�T='���s]kL�`z���LP�Z(b���8�� �G[�� ��t$È4��E��`p�DbP=��@��Y!�N�^`&Y���)�Y=��ݏp�y�
�0�u� �G�{_��)t}�!��x���a��	�
0Y�G.XW�)g� t<�4@L�~`PȨ��,=�N3�Y$�Hh��`"Bt#ΰX����;�T<�(�,�d$�����&�
EO�v��[��2�<P�D��@�I��sH#�B�D`�t$�'��Y����q�^Y@ǒ�� {@�F�P�9wZ\0 nS/t=�ְ� �,���^;e� �J��n u�T0~��& ��<C=�dG��n8���	�/���L��� �~j�w��`�$�R{HotIN�0J40Lm���@�g~Z� \�|8��3/9�v �t�Hkm�'�� )���r� �N�j�>	\�k�|[�XL 	��o�/ ��� ��y� Nv�e���� ��/]�~� 5)�Ʒۂ� �$�P<�Q0`Լ�W�t�,^� O���Ɵ z�yش;+ ��n�"	C x��^Տ��� �Ƅ�ʦO�X��G��@{��|�lb,
��@�9���~���6���,��: ������� oQ�Rݥ� ��t��9� q}��a  ��r���ʤv��d���[>�� x����� l�~���� ;���+c� �l��E�k h��b��<09��v�kil h��o�1g� �/-u��< >��@M��h;�)EpSjԠZ��l��*�}?-� 
�w��M \J	qO��,>5� �p�)Z 3��Դ�u��.��)��� �=0�^;�\��w����؜I�G���� ���o�� ��Q��� J�[���L_��@�E#�e ���~w�� p0��s��� ю���@� �N��&�� F�c�/"���r@�K`U �q�/Ǣ �՛WG��gN�{���6�x��_S� ��	�Y� ]}P�u�QÇH����4|(̮F5�-S�G� ���<,�$ �DɤK�Ob&nۄ;���B�	� �M���� �C~�t[Pw  {����I� ���ڏ����D`w��.�H��4CX�l ,�6c���;r� ��mP�L�� �~V/z�����]�D��p�N��t� d����/T �ɗQے�� ��@�&u�i ]���[ �:�hǀ 4pX����M�����ȓ8R�B2@�p	�� ~7Q����|j?��[N~�TDwy �]�1��� �̀�pS ���uoDF#�*P�@��v��� ^h{<�K�P ��c�n]�J�Y ������u�`��L�l�	������XV�= 㫄��^����7 �k� �3M�����v>{� ����%o��	
N�j t/�� �H����� ͣN�A� ��x	�S�0 ��I�o뤎 4�u�|z��fwЯ: � �n�9|��l G�)��r���}1x�yH��Aoπ�� ig�����1 ŇhY�P�� uM<�w�� ۨ���>6����2���߾� }nQ��H;v \F��Zkew:�z ��n�ן �|�EG�i�7N���K��v�8U ݟ�T� t���z5B��ȏ� V���,��KR�s�����o��x�����'�  )C�4W�-M�_���!64iøOt� �g�fH|w:�r� �v[���� �L��荴"��ܠb[��<%2�M �,��7 ������C |��n0�J�;�ۀ�6�s9�LUH�'q�0� w\�{]�7x C�A�|ޅ`���=O�w0\W�6�}�cG�Eqz F|!+�*�� �k(�������=ν �����G`<+�C�-K� ���X�W#�k������`��,�S$���E�[��]z�?� ��5�������L��:}ws�:�[����>�l����Po|Vt ��G��J� ��K�v�Q �/�w$ �sI���5�v��,D����3 (��:�® ��\g�=H� ,��WH� �\Ř���[�@�֝��?l��]k�����z
/ �@{���|�Ywy'P�� ij���_a�tZR2���� VK��MQ�L ��G��0א� k5�D�C�t\�� 2ɊZ ��P�=�{v�:i��l� Ăy�IJ �^�$�`� ���0x+ 4�	�l�ghո�ͺ���SLY�H��9n�s} &��%�tC�� l����)�Y�� �x��	1��f������~�� mW�od�� �܌C����3FA���0vh;O���`s�BD ^���N]�� ރ�ܪ��2 ��<l_��O�� ��6*x\� >}RQ{z� se���2ǎ \��[~ڵ,!EPL�`����� ��gG���$<`� z�ͮ� ���8i� ��GF�UA�}(�ͼ �Lۈ/[9� i��G>]�j�L����e��E �\@� �V�Ȝ� 1�[\�{� ƎҒ����*]7�χ���l���EȄ8w�O� (�H�<�\��m����q]p�����S9����.�5��چw�� I����^ �NE�x �	O�k��9;��8]� ��ݺ8�B ��7dm�� ��Okݢ�)�  c�ќ�H �.lwoey2,��J(�{�t ��D�u^�� �/��gLCq �$�K��# 
!v�Sp �C�7 ��s��v��v(S ?�|�Gs !�`��8�3_$�:������/�lJ�Px�� �E��Ƭ�� �3��V( b·f7�Hw� �sx����S��cU����?s '
w�j}� @+h�:�v ��H�k\� Cwᨔ��c�zjW��4�}����wlm
)rf�� �t��:��"��3�̧-�+{:C $|U`'� �蔭��_<9�
��ٮX.�� J3[�`� 4>��&#&�u ��3�7��H6 F}\޳т��d����0jG'y� �@��<��:13 Ag�5�� �n�4M�S q��F������[�J��H��۹�Q��4lny T+F�������D�L#� �ٽ���� �]�:I9x �`��w� P�D�������=���'��&h� X	[-�i.e>���Ѐ�wM������EG�v ��4Е�HU��}�X��,� IZ!YV�� 40��z;�:'* 2�E��P��3 �|�� B����֤ =��r��3�Y��x���/I�&(��� ����{L��&[y� x���� �K�m��̞/�ߤ��u�&�}� p~��� ��UK,� .u�nW��w\Nl���Ov/� ��^#���3�`ᡣtAT��k�8� ���X ���#%�y�zl@0��J:��-_�r��
�%x�О�]ȋ`�ِF�G� /S7g v��oh�~��˼RI>`��l�N���������� �+��pl'�A��`�@\o{�\) ��Y-I&�`�w�>�� +u�_� �
�{��z� SI�y�r�* ��_�iu�ѧ�{lUаt7M��_sS���� y�l	T�� �<��D�, Xo���� �s���/�p ��t���� �k�&�;�� |+
�l�!N�j"��2�� ����P��8:�>�E�f 0�
�s9��  S��%B �ء�Dnj� �g7�RӮ ��������y  �\�?m FcحSМD �@.&��x uH��\� �����'����� ��.�^� ���n��S�R I�� ~��9L�s� ��*�Vd|���9�O Gկ����:�_I ��.H�J�u8Zp�<��4{���`�d�0� [OI���=+�À����& ��ޓ	��, �8����RH x���\| �밐��� 8�y�0�����Ԁ&�{ �@%�q'�牢�d(����AxI}����� ��O�S�#~{ܨ��j�[ 3Y�qdL*~N��^��Ř��N�Z ��j$t�<�����Sw�b �yQ���ka \l�"��� *�����V� �:|��L �Cpk9ه< 4��E#�_�}�  TonB1��lc�tp�w��r����扆 x{����J k�/�7��y Nu�1�s� P^�\ԲS ���ú�{� U
��[��7 1���mb <v��\#� ��������)ތ�}�5�I��,z0� �Y�kf>�� -�}��DN�� )t�slh# Εe�xmH�������Ф�#�iS@+�K�|8 t���c��fI�sT��@���l��y; �Ci��ub D�6(fP 0K:���cF �b�/w�p ����<��;d��Ѕ�: '��{�ѩ� }�d��Dp ;Q(﹒���X�wL9���� �Kr�`I�� v/{7}�c 8omK�9:JZ �Q~C�� �(�g�� ��:���3,�D&m�"$� ����q��GB�\C g�nZ�� �:���H���9� jRnvOPJs� ��a,m: 5ﴷ�[�p �;�Y�'��5PL�B2����6��u����C mU@��H�& �9u��aF|; ����f6�ܦ��n�(t� R��]v;�� 2�DդQ�Ge��#�$�À�0ĸx� {l�9M��|= ��|/f��� X�-ǥ�A �s��M�[^�aH�I�0�s���`Ќ0zp WIۈ��K� wA)k�F\U\ D��4 I´ާ�!< ��K%Za�xƂ ٖ���m���/lE@b�J=\><� pG���W (�;L�nI��ȗc꽟�7@M�>�t@�P���3�q4������	�/� L�������C& �%o�s�a ��N:M��<�3~�ߔ���ض� b���6�#?eՀ9^Ww�� �jР3�� �gP
{$^ ���W[�� �Q��V`��t� ŧFH�t� �}��Ma�, -�Z�� $ �^דԒ�\"��� � ��|���4 ����z] Hq��A�Z��UΥ�v�W��/�0�W�['�����o1���x�
0=W �C-6��s{ 鮯.s�Q&��g<Sw�/W��{H��&it������ Y:���l=8��|���
���m�p���c̶ ]&�H��V ��u�5 v���|	�g W(� C��IVH n�\Gw�Ky$��A���ܜ��O w�F�Tq� #�� ���� k��o'~�n��ch���9�� �6quSGK� v��5�+ z�����4t�� K<�u=�	��]�k�����"tf��Z���k B(��yu� �\��U �sk�~�y����i`�� 1��R�bX� �n@,#w�� 5D�E��В�|| %��K���؄� u;t�6ޣi��"[��@���� Љ.��N� ќ�\�)> e�[�U�� �|�T�Kv� �t����ƾ� ���y�!:����e]���C���3R��O ���5� �@0gC�`�MO�N��/���TWŗ �u@>�VS�$� �B�mq� �+�hW����'�G���g.p�� vK�s@��� ��c�?� IC�4�-M�8����,�����I X4ߙ��C���8�`���L' ��hӵ8� �bǶ�~=�ո� \<-���S6�L�/�Zy� �uVtՓK hx��|�cryS �u��k�J �]��4�
� ����S N����� ���/� ���,����1�z�>5jKrL4�� +��! D����/֋u7�eȒ�I�L�,���xt�R�~� �<�J�G\s �,���E���>����C0�~ v��p4(�� D�ut/�-P��� N�o�)�<; �&a��'��� �5 ��e��9wm�@��ò¨<뵛��;b�y
�*t� /��H�= �OE��h3� K�m��, �O].��l� aI�H��� �M�3�� ���CoQ*� &ڏ|T�1 �Z�H��|� ��ЅUhx� ��LEzV�p�'	�As�\<� ���{��� �%�Jh�� M�s�eR ��FDk�jwV��B���Y��� �Eqm�k��oor�T(,h��n?�@$�9��#��PԐZ ����W[ ��&_���y �'�s��\ X�O^��� �<u�����M�����o�b�kerL׿��� ߟ�.*Ǿ �Iu���>� +AcD�y(T�&A�|�k�t��ڐ�-d �;Q�lB%�ЬK�|�� <����I�� �����t95���ݰC���S�L�&s7x 56=U��ht�>��0��y4�[8 v�Zd����U KD��2���@Mp�St	H��� Z��fo�[�QĨ��p#�?������� Ge��v��ʂ@��Wd� ��ɼ{���� �	���H ��vf�Z �0����{ 9/ՙx� ��&�'�kM ލ��Q�j 	�5hS��� ����VՖr�� ���~� �_�+ն�,�;�U �0n>8i�ɟ�=�Жx� ����!�Sa p��=��J�tk6�|׀�{��A�i�0�`�o��������cX _�QH��*� ��з�/�{�v� F��w � ;כԴ�+l�0�h���u$y�vL �t����B�\���J�+kX`���>� �#�\t�zvP&����� '�᭻�1M �}h!�B� �e�AY� �Z�,|<� ���\��tk �0��� )��rJe�B ������ ��$=W3] �,�Z�x	�t_� ���R~�O1z6 F<9�. ��K�lxP	�" ��4��Yb� �����[��v� �����y�d'�����(�� �,4	u>� o��V��8@�Έ� 	H%�t��<Q$�a� �.0z� M6���G~�B�d�l���� 
��\W� +f�,�q� �m[�g��:/������ ��� ��1��- OJ����{ >����4Z�qu f��g*� �^<PWR�yZ�n�� ������ �
=�� ]T��M�O�[o��LP��.r ��Q�SG{0`?f/# ���t�^�� ��	��D� ̙,~�Y_�ސ5�ϵ@�e��v�$�t����FWn9�u��T �qɢPU ��/��f[ C2�Z�= \��@LXOaUΣm��!��� ��C��G�;Ǳ�0� �Q� �%: j�BJk�� ���]�, �����Ȥ ������`0�� �5����?Tׇv�+0 ��_� �Y)�%��� {�ep+� :̮.5�wI}\F9����Hz�*� �w�M/\� K�lsD�< ]�tZ(�Y� N��[�FEx �{rIg4 ��Q��t� D��+	�� Hu?�8�� ��^��}C a�w�(cۋ �%W�D]�� 
�烙����� ��G}3Qi$T@� ��^����9�y���N ��mx�3s 䁞��X�\D�X� 0)��V�H�8���� ʵ���B��3 lĦ#�U�"��@$��,xv�O=c!��ę\91Z�{�Pru�>S|z& ������� �$��>�? ���Ki\�� ��I�k��?r����CZ Hm��_X� q~�0�ٸ:��j�sA��Ӣі`��Ԯ ��Y�s���W�*u2F���H {����x ��C6��h�
ȁ�����A�����(A�|�p����Wt�d���py����#g�5���� �b����/_	�v�� �.�A1����X7�,� �0�4�G'��k� ur}��Y�� �J���S� ��V�k� Oݷ�y�Cx 6FՍ�D5��J��g���\� #X1s|p�	�܅@gAP���F4 *�rpi�S� �y���+� ��w���A��|$�0�q+S��?G�"@��� 7M3�-���K� 5C�%0� �L>���c x)t�?"�7;`�������6.-�+(	��dU2�'>
�648������s	��j����<�'� ��kn�{ٳ8��;�$w �ﮬ7G�$�]�0��hw/ ��SN�*?c��`m���3J�Gi�L�սF8� �����;����K�
� |טL/��9 �W�f>=* �_uӑ32� 7ր����� �Z�N|�� LE�$��"� �TO���� sٌ��"� tW/�ڈ+n3� �8B� ԔMߴL��	��/)F �0{ ����N��� C)���M�Ν[�o�<�~JP��M�X�� �r�'Q�y����EU� �v|�m	 S�<�z�w[ 14K��QR� ���?�*� A+jo!�9�� �V����� ��xNײ )L�7g�t� ���s; ���+�>q� 2j������� M�,� �����
��� ��M|rp�cv�R\
iaZ���H� �w����r K�q�h�� �[ܺ�p�k$�l��afB߉ %�@�<j|� ��K�r�l(u�z
��r� ���0�|�<;/�������y ����'�S\�ؔ;⽉ U�]l��C ?��q���v,��� |�z���)���s4��͇u�S� ���?��L U7��uJ�� �3,=���������~�;��\� O*�T"�y?�x�z
?�1[�����0���5 ���v�ڹ?� 8��EWz_ ��yu��J}m ��pj��a ��˓��C/ 򻫋My6 �����ႝ��7����� �v` +��mo� �n
$HI )8L^f� : w����c��y��*��B� �"2���x �����Ь� p%"0�A� �{,HP� W=l���8��<�%s� �K�=2�� �G��ׇx� Q꼀0^ �9Syo��D ���x*6�� C�;Ĕ)�m .R��|_� ' ���$� C���uX��?\�v� �Az��c�}��� �o,א4���tU������� J����c?��D�IwZ����z��k�g s�w#�-�� �Ͼ�"	��oqwK��r��� �LjF�p���{���%�� ��ԟaI �k|�1��L�� J�s�ȷ� ��M�N} @����Z���;w�i�@/�N&����QV� ����;M ���t��#K� ���,
��g�Xa 2� <Ӏsq�| Z��ωݮ� P:��;��F���+7'� 	���|���`� �2�E۠� Q6���_{��x�:�b ��I� 'Ss(��� ���6ˉ�e U�t�@�� bQ�4 �5�� �h�u� b��m:� ��^��2� �Rn��ܭ �,��GTq� �
^6�tN��� 9�k_��� 3�Fѫ�^�T��;�U��fO`|�\ v ��'��,���c��t o\q AP�9ͤZ9!����?���F 4|*�ϭ�<;8��]�kSt ��b�a
���U]-1��}$C[� 
 �&� ���"k f[�5�&J ^�n;���< ���m�p ��#��� ��9YK�,P�v�䑦 ֙)w��&>?�� ��������IIr���JS o��
�~��l ^�3�x�9� ��|v* �W�Kk� 	���(%�� �"ӂ>�=�G���OK�S� ���R;̔� ^���|w �]�AM_.��@��I�{ �iO1� b��e�4 �&ֺ�U*P�� ��H�QM=S��"�@��+� _��I{0p� �,Q��vs ص�I!��� r�W���é �ZCS&=��#cG�u�� ����p+ K^��#�� E�aѰP;$ Q��84�v h��5� �M��Ǖ;� ��#��}� Q9���B5��7�Ž?�1ZHY� |��\ry =ԋ�-% �2�#��: ��4�
�;�؅���ؿ���x ��}�-́5 Bq�R�+� ���쏙��q�`j��W�>P��-p� e��cy:�O��)�q`�Ӳ [8i��>�	��'OkP�qJ.���c:I�ԥ��5 S����Q )N��@�g� X��pO����i�R������x��&.{w����dK��ɱ�y�3�YȐ�� h�x��;S \`�k}��� � HF�r� �0!^�W7 4�#~R$� �-V�jA� �!������{ ��D�� �i)`4onE	� }��&^ 0��+��X�� #�1�|c �qx��"D 脜w}ۇ��q��`lOp�� '���,�; ��^�y#�$�s�)�� K�Y`��ɸ S#�Mc ���:�p� <�Yޛ��*��q�N�kϸ rIK� ��wa�7 S븲� �~P� ��y��� ��|����� t��X'�� ���m�K �-�8L��qI��~ {��~�7 8�h�.�� ț]Z�����0�����d[m�O�A;T�@8�|7a!�_�ó�ť n �-�G�V8��NR@�MZ� ��sہ��� ��lNѴ� ��x��� �/��~0  ��ڑ�IG� 1VK=k�P��딠 !y����x� �#]⑹} >[�q����Z�*��0b� �y{�>� ���P�"��$�@�OǅTP�8zM�x�i>�� "�'=�� K�lq� $�<)��{�Q��b�'�Юa �A�Ӽ��v H��{f�@ ����竕 ]4!��k��S�v��xG�`��)� ��+�ם �jP��Ӡ��J�|��~"�(^� �P.'�E�Z9�x0�X$_ U�q}�H��������;��M��IY� :B�U�� 	 
=���!H [�c���� �"��#/� �=yM��E �k�c�K�F ��h�9t�$\�l>И� ��2
e�8� ՠ�o[T9�h�@�z�@ t���U3� A����?X�f)�i����z%����� �r�ѕ����J��`����,��H1	���!��2�����XNZ��[�����R �Ĉٴ% �2=Y3<1W� �_!��Kk=�H�h]� 
�F�)�����`BO ��(��T�N �r�I���������x|�B� 9v��b�_�ʊ��:�Hy<�@o\XQ�>�C�72ڲ��dI�O��ķ\���S�T� �Y�W炱 C�Q���	 �H�,�����  ��0X�] �%;�� Z�B^)��6 �����z/ �a(�R�� ��ר���0���"�(� �U&�á�An���[N Ӏ�Z&(v ��z� ��J ��+!�P�R0�ʾ
��Md ���t� ���pȸK ۀ���� -�m�* ��C�O�� 3�H�!���&12��D:�����h �x
�b��vI�A��V���	�0�P�[~b ]��*�4&>�5���y��FpĖ�l �-$���> f��#�$P��<U������� �5/Ԟ�(�x� �����\�4 =S��!�O�. b�J�Q�&�C  fU�� m�{��sS �w#Uן? ��4�*C��'�[qϾ��?Ⴠ0����� �AL�|V%K$��f� ��U*� ~�R�' ���3����2ԟ�B ­ܸ D�Ջ[ 1�h4M��^��� �ڰI �����0 ��1��Z  ��8He ��̘º V.^�H/�L؈ R�(3���� ��\f�uD��0�Z`��&`� ��$ƨ����q�&�䀉+��O��b�� $O�h�"��F��	&� �
� ��� �p��P�F N�g�A$= �~�D�� 	���;3�[_�|�`z �:)��8�p�q	 lRI%� q�o�؂�� \�Ð�� ���% C�u`��?���G^ ����j �����|:�f@K&Ni�PR��S����0H�L� H����8 2�P��� -�;��_�s� I	@��֞ #��'�<�v:\�" ����V�$�Z���N [��T#��B�J
��S	 �)��/V&U��c ��5a B��1��8 �-{��* ����X��<}� 3�&�E��r���&f�� ��Y^"� �L5��,�� _�O�
!�R��3�l� ���oQ0�n��W�y? )����$� �!pm��0�q`�MY�� C�2��� ��?��QHs�&Ұ���	� �hN2�xD��P��P _��s���w�:΀�4�Z��s�tı ��fH S��D�u�����x��[��. �S���qe� ��?o|p�X�� d�M�~ r��/����� ���q�:V	i� _
�8p����1�/����s' <�h2.����i��}�˾���Q� �Ht?�] �5k^F��� bZ��	� �0���N� �ɢ��� B(��	Ó���+Ѩ�v� ��g� ��	t:�Cv��	�� B��V>�f��$���~y� ��V�����#�P���>� ��jF��� ��c��Q ��� �sD$�6~������̔� ��ph'��z
�b 2��na~P; �.0��-ܕO	���P hSc]$�� ���tæK�L�P+�aH䠩� �
��(� ��`��0W��/ ��?P ���v�K@�iYZ�-�`�V�N����� C���s� ��h\/����ā5��� r� �	�Nt
8)� M6I�[�, n1��#.q�a�!�����^� ��Q��Y7-��`��Ǧ�����2� I0�N���7 @�
���0��������v�?����� 咍a�\  �fjHk$�cB�q�	��/!s���� y��hM�흩�80� �"=�	�J	�+܀[�|P ���Q��x FUS���= ��P`�#��$ �� �Z�SP��q	��Y�� A`+�8' 
�~!��K C����k&E -*%y �Z�FC\R��~� 1�h������.��@���¬� ��O�`7/E:��#�@Θ�)�gӘ�3V\�\WB#Հ�G�y a	�b��o��-1 �B<5��� 9��!	�hn=YÐ)�� �J��g� ��,0��!v�q���s�K t�|�7���<%܀��/x� �V-O�P?[(��R��u�e��^�D�!�����R �A'�� � hVȵ�1]�p��Q! �Ԉy�	 �L �r�$� ��%B]�:��/Z� ���!H9��P�:J?z #��"
� e�>��h� 4�W�ly` ��2�A��(g��%u�v��Cr�����9��e��2����`�hN �=-?Xp��������Z���!�^�@�}) �j�1�ulp� �ω��N��z �Sɮ0�� ȢR��M��9�!����Q�Y� ��{��� �� ��[0�W~�.`�� ,� e�� �7�:�p #�_�N<��2O�� ~��CM S�؉|�	 �[��� A:2��R� N��0hZ���Q�@ȹ{b* ��@R�~���<8N��3�b�a��.ƙ�柼 $0�\(˦ 7�x�����^H�Ä�y2R Ӻ0|;@�~9��%�$�� �]��x�� 1G�Tt \�d��%� ��_��� {'6EL�Ox- ǅ�}�� �n��r�r *��)^� A\>X�K�&�.�`
d��- Q՗+�w�`~�%^�/ j#l�G� Rh0 |=�� 6+��- <M�'��7���&Q
L 5bXI12؃�� �m{�% 金��b� ����4�� =��R�bx ���>P�|�OY��3v~ϣ雐	j+�=[� X����� �g�G�! cV8U��X�~� ���3u������,�<������ 6�!��ܺ�{	 ������pX� ����c ���.WR�-C��d�@Z��X�]1�@+Y� x�&G A6 ~�0N"�c 	���1�� ��p��2� �Yi]^hU �1:��G� ���Rº X����� �(.@�E_!��^40X� 1�)�X ��h�^qK�v� �*�Y!٠���%L_� ��� �OK�Đ5.0�>� �~� -�hE��M,!��`�b�`N��� X[��Q"�S
Ի'�`F� �t�4�`H 3(�e� �-@���)�}_ /���K���z����F�0� ��T����Z����E�k� /iz4}Q� �9+�u�� ��fL��� އ�h��	 �����S |�&�(���NV��
I Z'P�Y���:������;��z�M�3�W KY	�jf \+�%qn�� �b��1�Q �0ك���</��L()��R x�	��� qe������?s�r���Lb�@u ���_	��^���O�9������pv> ���F<���n����A� 7"Q\y�� �@��b���pj ��MJ%,,7> �V�7���� @ �!ͳ�� ��|�~ T�	�a���:�\� �&\|@V �TY^�� �R����hv;�FkĮ$*�
�L: &����4ҵEp�~�|� B+�S� )W֨Ia�� 8?&�6F$U�@h�[�8��ğ;���|�
JG��� P��2��"b��~ ��!h �݄��\ ����֠��  �Q��!��]B�����������JZ��Y��&4Dw��2�~P�Q�ke����z	 ���ǆ��] Y!�)�ҭ�� `�n0�R����H1��L�fhR��^#C��6�P� \dc�0��=�?�]���R�� [�
�KyU{�H��?� ������#H�XV���U�.(� �-Je�� '�_�`!ے �����8 ~�9�!�� ��ZX+ ��'�"L ������pB���0� �˗��1�&0,� �	�D�O ��x����v��R8�X�W,�� �(��S�� 	�
 ��L8 (�Z� [8�~� b�$��v: @�W�a�� �r/�4Ѝ� ���8iR ������h �p|�f����� ��驽L]�� R�DV��^ 	��Ȅߵ �N@嫣�? ��[U�����A��"� /�g�(ub�8`�>L�] )��c/W�h`�Q�^�U���u���X@�,]! ˱�e/E�� O�>Ţ�|cu��1g�6��)��> �<����q� 2�|����p (�d!���acR���p�� ^	2_ 0"� �L:-�� �3���1��? w�nZ*��� s�8�
y�x��u ��� 9� �#�� TV��@)C%8�`�U N��t*�=��� �%W3y ���窄M�H��a�	0��Yo,��� J\˫t�?�BW�Z��a�0 � �V����=��[�_'l�����R���-:�*�m�a�@u ���n	y� 8Ť���X��K��bк�J Z�R-VC�q �j��Q�����`���tk!��1� o}){�Ff:?� �4ԹZd�HS�P�� �0%��k�	���� �� ^Б�c.s�H�A���_��@��YWń ��}����� �]��P�� �D�BR�� fs�U��J	���̀�Q�� ���B@9� ��=[%�� ސ�a	�"��/�(�_t� �D�0ש��
�A�4�O@U8:�. �f	{�� X�;36�R��d@�>�0f01�(g@� �83�]�) ڇ�#^ϗ��1�I
��D ���c���oH��)@� ��*�hiP
 	�D�X�/JQ1�h�ȇ�H
_�� ��:���.��� V]�c^; !�Ϡ_*�h&�sI��� 6�=��!�� "�[��M�{/v.`x�U�n �=�ʸ� h���ٗY� �\1�8�n��K�����y� �w�[�~� ���g��\  �@�K� ����k�8� Wn��rByy�`\� X�Av$� Z���)* @��GK0��"�j~� �)�"��X�_��/�y��E9�	 ,��#M� Ý�
�R ~Y�-2��*  �c�t� ڧ}#ZY�� ҂��Q7 ����(�4�	1ݻA�� �Lf�&P�� ��l�a�q �>P��fm� OƵI	�8��;S�� L�y�(�s(����� ��1�K�V+ ͻ��&S $[��_P0�� �����l![�K�1� *Nǲ��UQ ����	��;`� N��<
v������%E����/�� ;��!( �%���r�J�����[n�3N { A�W�(�b���}9 ��� Hs��рI��V��i��w�;�J���靶@g��R>Uv����(�� ���@"�w gNë�szO�����Wj 	�wSbD� ˀ����;���-S��(�ٝd�`�� ��yY�pؼ 0h��5�Z g��6�� �3���:�� N^�	����x�ȃ�� R�
�3}�YX��2	��e\��S �����M� �Ha3��y	��0�J̚� �a;�	���b.h}��� �@�R�	 "���]��g ��@�c����� 3CQ��́ �
լڭaXg��>�m�Y� }�sI^��� �(�����2[�F�UI����!0U. (Έ�����< ���e�A ����݊�Y�0�XRt E-����N��kP�J����A B�2�%�	� |v\3�8!���`�P%����� �"p�h�IL���!��$��.%t�X�ظ<o+�_�p1��� `�C<Ox ��N�wB�
�8��9v ��Տ�V�"�Ч�Y ���s]� ������ �Y��2I�� �߉e�׸9h  F�T!��" �~�J ج�?�O�,ɪ� Viܟg��;�TY/�"`��v� �- .��B�M�~ ��P�4�恠��? �5[��K��XL� |������ �� �-�	X0� K.��+�' �/�Qr|�H]�%���(C�9
�@�ي� ����h���e ���Y��	�Q�iE`z� ����|�� !�Y$HZ�^6WA�+�� E�G1VI�\c�#Lỳ0� (�YP)�T  �,g��i��K��� ����x	���� ��h���Ⱥ �23�x0�PM�r� �R��1�� Zth(\� �y�r�1�Q���H���Y� �rX6`x &8��y��1���2Z6��4����R �e�|��1�>�ZQ�ҽ��^ ��S�K� ����%��L@Nʨ�ܒ� �Eä� �.��-��	 �^PXv�Đ ��|؉� ��D{32��dSE���� �:��.G Ph'K}��� �u(��݁ ��Y��� ]���o%s�	�q���e��� �K��s�{q�# z�~v. :��^Ľ� ��io�v�b��ɽZ`�� ��']�-q�2 �	z�� �+�3j�@�1�Ƌ؟�� sμBZ�	 ����8`j�2�I�,�i����Z"B��1��n�fC�<<��	�#��-��/"�lԡC �@��R�������0" ���	T�|� Lo���ww� $��ݦ��H� K�a�XTb @.[��%vM��ϻ��
Rh�������� Qb��l�O� �]�S3	������� I�?vp���x ���Ls� tJY��X�
��M��u�/ST �[�&�! ��_��Y��Fn� ���Q e-���! ��Ծ�� ��%#`�� ���3�V��M(�
Wv� F�1�:#��a�h� �����\�N���`C�^ \�ǵ�H G8-����� _��[5�!.�di�;�  c���>��[Y90@iK?�0�F�nHz ��:S	�$e�v P
� �k �')Vo�z p�f���4� y��(�p��r�[M  �v!iW*� ���P���� {��aC�n ��:ճ+��B���R��W@d0 �
����>�*�D#�X�;�Ӏ1���A 2�.K��-���q1�[h �uc�	��?Pa�J�]C��(�k�x]��IX�$|� ����d��Hs�'YR�.�B� -��a9V {'k?� r:��cB���� �`�s߈� O��4�o� v�1�_�$S�@�!ڹ�؀[	uk h�<�n�C~R �z�T*?�� m�����Fʦ\�Ɏj��ޱ �[��(�^ �h61�\�}� �'���� ���j�J�Xp�r h/XZO��ѕ�ɕ?
 ëqv�"� ӂCȡ��R �0ѾO�`)Z�~@��# �>���P��ֹ����.j� �'�;k�L2}������ ��ɺ�)u �;"�-�~ E�D���!��p^."_/� 	r���ޜ X+(��� P���L-,� |m��RO� �%�	��oI��B R�����Z�
�����U��wQ|h�s<��@^+I �2�6�J= %��fh� KQ��0 {����&C�  U�Bz� �\r���  E����6I� �5]��������Sh
�(����݀ â �Wb�[���PTXq��Z��� :]\7���w:�@ ��gY*�$�լ S9�>N�qq �*͘`0F�~��]-a)S���0�[������% 1�X����� �}ze�4Za �2�+T��	; � ���4�n ��D�ꇠ ��q�;1��j`H�0�V����.�O��f��iv�<-P����tq�j��� �=` )���H�L,�|�B���.�� /�"V�[' R2�)��* 7�hVk&�g�,��@�-�x� :�!�KHa�RȂ�����p/|W���,� ���;[9� ߉�Z��� _��y@�R ol�kQg?�` Z�6�DEh(O���%�)A,{�c ���$��� 	p�� ��b��P��-N�����9.1� z^V��<.> ���-Мd��Y }j$2� 6B���� �rb��G��@�S�KP`��H O����Z+�u��rR@��� �(Ɛ���� �*)G��da  Jޢ�{�� /���P� tS���� ��)�>�/+�0?L�l�� ��B��.�� g	Gf�w�xC JF"X�h�t�y� ���zK1� Q�@/�N �S�]w��L3�ʀ��� 8!��_@ s#�h�u�� �膳���U
� ���\� �E�"����'�Ld�U���vH�'.��+u��p%�� n�"��=5  �@(Ӌ0 �£X� Y�����۰ ��/O
�� ��������h�z& #Z���N��!	a�^�t�B�x Q��oY@ �21��� dZ�eAR U/�t]��ڰD-l���1vg| [{�.B�n ��%	�V ���N�K��t� }E��� [y� �a��Q́ &�#x��	��T��0� ;�O����	a�~ KC�� �-o�{*�3�Z�P�[Qa���7 g��AI�>Wj���)�b�B4L�D+�Y I�;�M
&�J _a(�V��k������K�)>��Z_ ���>[h�B��Qd��`�lp /2�۠ | �L����X ��)��i��w�:���� a��z�����e����(ψ J Ž��0��������tf^����0I�	S~uY <�1(� �Z��`^� �!���� ľ1W�f>� i�JC�� ,bqE�ž�
�Pm�� @�oW' �l�����ب�����9S x/ұѽ$ ��E_D��8Y��!��(���  �`-�I �R��X���d���ź K�:��S/  �y4I�$vT ��� 	1lՕz)�-���3L �/g5��P \��>�/��O ,N�Y.�� �\l��R$�� �{���r! Z�8��1�)�X����C��+ k���p� �a;�H|�����/�[�´�G ���<S�� �mq��� c�Ϙ�Y���d_X{� �( ���� o�����}� /
���u@&��-���_�ZR�>+�Ľ�(����,� 9a��}{��v7 �#�\h�� ޕKQ�j�	�S+(1d�|0_!Yh�4jȚ� �D��n# � ����z[�) �mS]���X�*.ؐ�=@'�ɤՊ�1�m�/���h' R�vk�JM �5��XhY]����Nx���v���hQ8y�:� �2�S�� �ڇ+��N���Ta� ��)P ���7SיC$�@{E�94 R�8�QK�Xtp 
��:0D�N�B�XЂ �u�V@Q0 Թ,�~�K I��ı \^W���%�'�� �{I�.�� �i_�� �%WUq# ���:]+ �)��ϵx}VL0K qmi�2Ĉ�4R��09x�'D��ѿp� �;O���+
n���1� OT9�:� !����� ����� V�>a��k �	�)�� ��R��" �W���I	+����. ���/A� ,m��� dc�s&p�X� 19��5 D��pA�i �ZCn��� ��ٲ�� i
߃�� ��%X� FZ�{�t9) ��M�}I� �4 �E�ml( ��_0�  ���yX�¥ #ͱ�����,�$� GK��*� b�E\����.D�N� ���0�N \4������[@�v t��R(� �ׁ�o0� S�P���= �.m	�5 oD�ρ� i��8j���pԈ[�`�\�	�)^ �`��Xb� ����,� ��F݄� �a^8������0M׾��})�%�� ^�d�
��s ߈��%���\2�Z*��ʖ����[D����b��=}�$20R�rd ��[��0e��{�s��qu����!`��J=�� ���K	XP(��� �6 i��!��5��"�R�o e��� ��2�!�� �4����h�B*��ٳ$�#X��֠�Е��1�Z�ࢧT ��0�� �FG`ݳ�y�P���L� i*Jx�(�� �%#�q+3� �bS���� �a���i ״��� �\�[c��~Q|� O��3�|[a���u;#]�' ���+��c Xy����q
��U2��lP� ��$�����K�%{@�Z�� �0 ��q��U�Eh�c@̱~'�� Df��,�B��cWA+��2�,U� ���nz �]�1 &3	 ����� ��INK��#r�	���� �b��h T��(��lE ��!Z�?�?M��_�d6A 
!h$�WN��4�@3�+zL� b�S%�[� �1�R��� �j{�e�x B���`� )��U�z� ���$�_� )=�ɣ8 &���B!��� ܨ��:�� %|��!�� �{
Yw�8rFp��	��/m�`a&����
_ �r��#9� 0�Q� &I ����(� x�[ ��LR�SQ@Ź�s� �	��u� fR�����? )&���Z�f> �_ ��S�M����	I�3 ����(&A���4���+  ���G<9gp�UE! �8����^ ����k�� XV��w�� 0�h�F� ��_�$ �aR���/[�����2�� ��k*h[ ��<���� H�p]?�G ��LoP ڇ_W�� �sX[�^� &���3! �*�C��[ ��8Rc�� �����_7���' #�P6�R/������ʀ�Ԃ VQΕ	�����@�R� c��G�4�� �0 �X��>� �L9xO^�I��Q���v�A~0�a��5����_�LwV� �)�Ya0����_��o���l ����,#ٓ�	�N�L��Y ��vm�� ?_�O�� 4pE+*���AX�1�%`�C �Ns���4 �aĐMPX� °��[k$ ��\1�?�� ��pr�w ����Np�l �$�8`�_*�Q�Ø�P �%��+�\�	�o ���y �z�hP`� �'��EZ��\� �.Ġ�� �+Px|���W�/�'�� �9���:	�;�>7&�5 �1�>�o��C�W	�఩`�(�~� ǘKY����ɠ��Q2�HW�o:�c�6�	x+���Q��?q4 x� Y�u��;R� �V�2��v� >	���� ���/Ȏ� �hg)� +�PUR�� ����a;h p4P�Ͼ� �0�5|+?[�ȸ@�oֽI�� %Y�詡��$�_ ��!�	�^ ���� ?�� ��6 �[�a1�/�=�8 T���h;iFa��Z� ��j�P�$ �y��f]� c/�H��k3�_�v� � ]�ѷ}A�� U9�F�' R@ĺ�J\O?u��������yq0���	@���00��� ,��7!�0U���ͮ�B�y�\ !�-%$�I 'S���tG b�!��� �2��YQ �(�?�-;K��ɻ�"\��
�]J �0����g5N���} �3��\й ���h�Ĉ~�p�~2�#[� Q�&�=݀�=� �o��I� kP��S��T�;��#N߈�1K�RW��L�T�@�S�0˸��$  ��_bC]A ���R�Z���C	�j���� º�^����.aH;�u��[Q� �N�C���E��L��'\��ޘ0�"�_���\������(0�� �� ��O�t	݊wʷހ ��"��r�� *׹�kR2+�h�'����[�A"�����R�V 
����T �`�4q��O$�p: D�V� q�`m�u^�摀�H�U  �v4��P �k�SB � ��� \��4�@i�	_���2V��� ��� p����<������*	q3�.W 8�髨�� ����ZW�%�����#E' ��i�B�H ��q1�Ux� ǽP7�Z]iɠ��'@� p���h=K% ���rZ��_� �+��D#� N�!L�1?� �[}(	��ޙB�r��H� ��J�]*�L�  X�3� ��=�ҹ!�?��kh�	���\�~Sn���`�� +��p���� ̓�@��7 �\��� �I�W� �Uh�ԨO	�0 ��WV/kv c?N�n�j md2	�h�T�X_%����B�
 ��[����~� �.V��
��HLt��>� ����p�  �)�]S�� �'�i�`�@���҅�G^_kpo��{~�'�f@!�?�> �.���N 47���� @�_hKO������'�e�#��<�􃉵QA/�!z����x�� (��T ���"�N �7pR�
� �	�hCP�� �}���q[��ǀ�U0�Q�'� ����(�"�1�]	�Z��S� Gv���&8s_i�+��b�vW|�A��.рQs�z�a<��)ńoX����\ 1�v(ҽV�JZ�q6? ���n�%��/ZEJP�[���]�2� Q���Lu�d��} ���P)�0 ��f�Tʔ �-8��F `;��_�5���$"3wN��Tn�*z'� �aA��I"G:�(���4�.r�: )�� �Ҵ�	Y� ��3��� �C���_A� K�퇃���<���~ �O%F���� �M��I#"�/)�PE��������`Ba� v*P��W� �隈�ӹ��X��=[�������A}~�4t@OPI˞.D	> �X.FJ� %�O/[V@�8n�x��_��9�lJ�v�8i�	VW� �Y�� ��ͬ_�' cx���l��@-���� t<G�z0�� �!��P�: �����]��G���e��d3�nM�O��*X@ &mK~a�Xk�@�!t(b� ���W��a䀝i�B���`�>cŎ57c�����.�o �����~ mИ����I;Pb�ߺ�j�@�kN�� �1��w����ɀ�V�'�< Y�B�0�Nl�{ �R��K�H�A``�,�1�@h�7�|� �S�����.l�� �xp�� %���(ㅬ 1��(@�Ԥ���Ò����0�C��"- �hu�e[�� ���ѝ���x�� �^�z�6�`�Q���5 =A��kü\�A ����_�vG-1���Q [:RvE
�� ��	W�ۂ5 ��쫐T%���O$@��>�� B�(��R�r I�'sP��&���F	���5��n 1р�S	Z#胓!C��;� �x�R�� ��4�� _J��%
zRV� �l` �F�Ͽj�����g`��d ��󘦠D��1�
��Yh ��$�,d�0�]7����h ?bo1;�VZ �:X�:'Q���7�y� �����L@ !	]2�P�:e4��;�_ӵ���p\� �W�ϸ	}� �����
E|� 0��v�������/ׂe P@�؝�V �5��%����N+Ԍ�P:�� ^- �P�A9 �2�C�lۥ>�D� ��A��o� �O�!���Ҟ1�0�d +bؽ���`l:���2�k�!���݀�	�u�<�π$���z���r7`��� 
�fˋ<~� *h���� ����Q�� mA�2�	"?�H覿��0٩ x�n&b=�-�_ F���Dq� � lP����֥ �|B�S�5��g���@� Z(П���E� O��wa9[ ���)� $\Z��2@OҠbް� Q�0�Ӊ�`f��%�KC�Y�@Ֆ50���@�KA 镈?��� <�H-���A ���+J
 �O1�g"�@��dN�����/�`,��1�g}�s��f mp��Q� �ΠY���! I՟�w���d����\NR�J�P��q�rD�QT �Y.��>m��[4���
�t~	s< HS���ٰ� �h ��%� ��}�W
� ��C݉�(8�O P�*���� 2
�\D��b vcu�H< �#��� �	1�z�(�m�v@��s<� ����G�u �� �x fA���S�J _7��ܒ���H\(�Ȅ��e@�[�P�����
��O�(0�U ٢G���؀� ;�xS��� f{?���O:832����	���Y�[��K�t" �����Bf��u��@_%S ����z�Z� �a�h�	�� "�\]�O���c�*��� �P��B\� �cd ,*�� 	�S�]u(�K۰���L�%:� J@��j��� Rh`E0Ҁ Ǟ��n2� � �c*;� Ҽ�e��d�	��@ Xn �/pZ��� `�.�	�Q �g�&5 a"z� ��ȍc�~����`�$��8]�H���2� YD��V&TZp�NQ�ߢ��a�p�V�([�"��ݜ^=+��!��� �(�'�r�6�E���O��X@�����$�� ���>+�� (�|[�!� ��ZAu+n݌�(uD���� _�l�
2 �P�u�L*$��;(���y�0I <�[�i� h-�̏+��	 ,T���7� [k�z_�1�F�`LvB ����Ӥ �P0͸45K�`> ��� ��W�4.�)ۚ�+��r������x�A#���U� r���h r|3`�qo�E����Ip�b ��"&����O��-���=�N  ��*n�$ ��aJ���� �0�� 韕��� �q�d�k�ܾ��T]����! �%�CQ"/x�'w5 `�I�
%�&+ ��bx��~ u����^ 2�:�+�M_����`��X�o�n���� 3)Y	#�h`�(򞹊��F �[I�ۇ��/��������0�� E�
��@� ���`x��� t�&��g h�MJB�� [����j	(���<��d X���v�Q����;��R��ɸ�P
� iĠ�?���U/*�ӏЄ���Y�i�ǰs+AR�:��ن� n1��|~w�9� o3�Z Q�P�{� A�d�o �� R\/h(t>�PgD� [R�A+~b��|\�(`��� �¢Ri���`GW�GM�����($�����F ��r�� ��� Y����@ �S#Ɲ�� �JQ�X� �^{�A�1� ����� Z��W6 *�!.�V$ -8���)�l"]���`]�\ ��f�( �sR-'�� V�"U�3 �bXq��� 
	 �a�� !p�.����聕��z�>㷦4� 3%�*�w Z��$X�͒ �IJ����)��Mc�iBqL�p�� ����� if����a��P%�,)� R	W��� iX8���� ��A�Y!9���R@�.i�pT ��Y���� X�0�Z&�]��VTDCJˀS ���IY ���01�<�����0�O(�R���� ��?�O0 �!`��%��� �3ua	 1��.�����( G���Vk R%}h�� ��\C��B��L S���	 ����919K�B�r�� � 0�C��Xi��&�;n�p/� ZАu�_h &�d� ��)ͤ3 [/�R���>� ����F@�@$)�HA� �+��*���o�K�k��� ��waz�s&��/ߒ�C4��p�e+`��oUi0 '�T}p ������@��-) ��V� ���z� � ��R�ٺ�p* #��v��~rq� �B��U@2 X���N� �^�/���J 	����09�� 
�S�Ĩ,���v�[� �B^����	�P�?� _:J��FZ(N�����<�i��w����9_�	`�\�� 1ʃ�dy�8�| ����O_ �}ϳ��C )ſF�i�l ��1������ �X*ʉ �
���	 ^�[��r@ŋ�p�p������� �(W���v YlF�$!�t�~��U��v�������	Y (��M~-���� �mr�� V�b�4x���L���J�]���NY`��'� Q�h>�du��� BI�,�ɽ� <�
Y"�����]ka,$R����-�1�m�� �{T<���XⓁ����C� (��B��` o�Z��ri^:�������
��  �4	����a�ځT� O�$����Ug>Ph�; L��-�A@0�@�
I�<��_�� ��XS�� ��45��0}�=�� s� N�� P��qdAQ�ey��v�T.
�%��pM l������IS0���*V�����O�#�9� '`H�{k�RQ ���� ��0�� 5.��9N�_-Ò'������ +��X�xQf 3"1�Sk �hH\� ��Q^�5��]�½� �Х�"I��	�1� �_?�� -�`��f 5��D8���� b����\�X m���}�N��K��D㼘ƴl�I�/}$��@ !ɺ�lV���20��!� >��]� %�}?��-�!���4H oj�����<p}�x�� ��sP��$'��d f[Q?��Z� �:�g�$� �V1��Π0�����`��n�� $�/�K>��R"��b Z���Wtj��  �*ۿG	]�Y_ ���-+ްP1��z�`\� U)âf
���,���	� ^R��9�� ��f���q:IH���^�[ ��L�"�� jxd��:���V �aP�<�o!�ͿpJ��V(ؾ�C.��xJ�� 1��m�]cK��^�u?�hb�� �m�C�\�y ��g^�vZv
 Uũ9�m�$c��4Ǽ�3�P����b���p�&U������L��� �0�@��Y �Zh1�b8��9��`�� ������W��� ���ǆӎ�z� ��41�/;��H Q5���p� �����n�֎D� �P�:�z� �h%{]�� ��O�. -��/��`� '��ER�I��
�[k`�Ϸ ����T@	�2�� �z���`Plʹ{��GQ���am} _��� ̬EZ*�! j��}8xK�d�1�0�S 	� ����_ ��=+�����3 @qL��f!� �F��<i� ܶ»b�n� ',�+@X� ő�y9� ݸ)�5��� 2I	�YW�48k�?V�.�J��>��� \��� ��[(v�&��� �᮴��=x+ �B�ڗ � ҋ)�IX�f��ip� H�N	  CEI�DW��7����p�un d%=f�} <�P ��S�<��=8O��z��Ԕ(D��"G��a4��j9����'� �Z:��Q�0ü�@H�e� �'�G�����;yM��*K ^���e�H ��.��	3�> =�� � �;�Ҿ1 LQP.%�� *�z:������G��V�P�s X�r#&�$ 3w�N� ���.S��y� �4�KgJ�!�֬D)����W QGB
Ϡ���^��*�U�jʽ�@s��;Bg ���f�"� �:-�Ao�u��r�X������� ��
� `�!�HXsO������\�� �0�-����Z��)�j��'�̘�.1�� Z����ᾘ��]Wt� p)�-��  GA��
M��< �Z�F2 !O#�:N
����P�?+� �[��k> )�`�༉ P����KSY%�i�W ���!��W�W��� �	>B��� ��-ֱ�F� �M�#s� �X-�wQ� �d}���fX�	 �F%r- ��Lwn(D _�Y�W��>	��� �G��c ��HT��(
 �eo�hD�����Z��" �Q��5��G )>Y�1�kv�"����Ѐ�� ����j˫L�1M@�*�G���p�� U��XW�vD '���fK��O�� s��! X���h �T�����o��� W(�]��-* �A�_h� ��pJϝ� ����l ��F�*��0��(��o�ju{��Ӯd�� �� 	�D��{5_@�P � �r��+!��$�~�X ex���UIr�Cҏ�+2��� ����S� Ŕp�ސ���w	h�D��^�<3�鳐�W ��bB�#xp� 1�!�_��kGU��Ai�H`_��%$ 
�B�)�,�b��\w�Y�C�qU�� �Z��J�^� %`_��� �����+�PMaRˀ/���  ���[:(�$Y@��ث2 ��}�)+k� �[��V�J�!L@�誆x� �Ш�0� G¤	���Ѱ%_�l�*���$�Y�n�c@�G;�R��N� �X0� U!�u������
� :�*�=� vC^-�� ��ٽ,UҠ�z�P�] �>˘�䖁 �Op���by �<WL2@u�?O������gp�@eBi7� �O;<n -y��i�� ok^#/PL��)� �Y1E�` ��4��컃 ]Z��as(� j	 Y�d ��!)Z�� ��08��ݛ ���n�|� cWP�ȕQ>V���JZ7�c� ��5��j ������ o톉(	͋��R@�1O�<p� ��^���H���[QW>���`��������R�ɖS�͐��Y V�0��b�_���[�ނא� W�H�	4_  K*�\�,k9��A��$�� ��Jk�V"�����(� )�Ѐ-�	Q  k�I|�Ӹ ���bA �y��+�� ��'�����)�2p�c��~V ؘ�	Ѥu ��=�-<�� �@[p�� o3��ub���p 4�_S� �cVY&2F� ���:��� ��/]g�Axn@��"�` �]�(<^W �ٔ!/�s�$D�@H-�Wrq 5z�!�� :�L����jI1vv �,9f��$�� ȭ<:�	 ��I��` ������d ��}	�������0���a 
��������.;� ��=�* �чڽ���� ۈ��ᰑ�?J��� 0���ϻ Gm���[�w�F$�k. �� ߫`�h&'����!ބЃ	 ҕ� )�0��I�,�#��� 1-���3y�:���&ET`D	  F�b�˕�D�HȀ�EҸ� �
�NP����� ���`�<����;�؝8 ������'�&JhY��"�.0H0� �U�`-Ι JK�o��^V S�	]�r� �/���Qg�>>�1�@+�%�W��m���	`��> ΀��kYTWbR) !u'��|�a`�����X� �1eJ- ̬=���) ���%��ynp���,�F �5��!=��6)͵��\�, ƜwJ�� ��i��\	��"��-�K�� :�϶�a� �I�æc���{J?�S�yd��O��9Q��u�
���� ��.�}( c�y�ÛU	 �R'|�[ T#���� W���+�' U�Yhd�\�, Io"@� 볹�0�� �?�1�M�H�_%��$ ˅�X��J%�3)��`����N�� =��k�h~_Q ��*!N����4G���-8�B1;��?�� 4�#'
�q� C+T	1�zO R�\u׽l N���+�D�q h���"�wn�'!�*�`� Z>����@�_K	���wX h�lɞo� �W9��"\\� �ܙX�y� r�%�&4 !�s�|w?� ����� �aNh�z~,&��: �"���� ��\�ˤ?�ЮQ`�M��T tO�ոg� �@�Hјc #�%>�� �Zʭ_	3�` "� ����>����+ t�}��8 e��K6��@XZ������f�� ��F�� ��@N����!�pb�И�_L�y��:@�(�5��{xM��-�s;)� �aO1��ϱ�|tn
�OZUQ���B� ���0a�� {����`Y ��%1}�ʐ>
� su�6� �q��H8� �����# �	�Z+�H勸k'F��u��=i��B��h ڹ˲)I \ĊEL� W� w��2�sQ hy��1m� YI�{��N�<n�cJ``�0�v� *4+�IGHw� X���N-É���ם��Y
 �hqbp1W{|� 2������|X��H%��e�d���/}� �?5��9���}��X�+ �DIV>ލlĐ%J�� � ��(9�u& �'���-�� 8i>���� �蜓����@;��,c���5Ks��iX�/	 �ө�PW� �5=�~pu� �j؀0%/X`TW F
��� ��h�S� t�!_ˠ�� Y&	�U;ّ<Z�˂b�@ �(=ρ���q�`L�H>q ��pv�% �Q0�K70Hݪ�I���>cp���!p@�^-i p/5n�� E��K-�L o&Ŗ (0ڙp��*��,J{���� �P;����z ���� �
	[Y2�u)�P�� �p�Ĩ0n��h(%����5 �#SP���_�NA	0��'�]|�B@�`�Z)���L����%�_# �sO�} H"� �k�� ��<��S�� ��[\�C �`~1��e ���WEY-�� G,~�o����$� ��2R� u!��cG~j ��8᭽6;S� �
�R�O _������[�f����� �JL�tZP ��H�K�b: ��}�J�g�(�N��7u���Њ����K�J0� �
�"�/�@�+� n�ϑ�Z $��^w��K 캰��kI� tL��Z˕ud ���X��!�*�](�AБ�� ���2��;��#�\!�|����&�`��mK��k��8X_q ��n�� �2-0B���� ����2 ��Av�dV �h)C���%. ��҃��	 ���F?�K �M&
� �� �����Z� �o�1	��G[�1�$�`�d X�'k"�� v��ZKb��u�/!c�8���~�,WUT]���2 g���n XC���D� �R��h�- M�x�[؂� ��.�7� �Fc�hPH ��������O��0��\.4� &*�/h@�����P�y�����uY h�:�V�XH <�K�3��~`��\�Ժ� ��.��q� j(� �o' +�zh.!�l a�6M��vP 8�Y�@� ��ߕ7�a�A?!�}���- �[P�� KX��תB ���R�� �/���a�) �&Vx�-X ��kNq �` ^�ѽ�~�= 1�3�[ (�hV�2{ڠ��Q�� 1�0o��N��-/�q��� ����$o�w���
Y��t�� ��"��� �ٍOb%+�a0��Gi:j�1�@�����(�\���a��n���7NupF?[G@��.M �O�e�^�� P׀�}�- ��޶�7 �ɟЋ���w��\�9��|���� ����l�, ����� #ى����	)�@�΀��2��s �9$��p ������L�� ��b),���yW	�ܐ x�3P
��rh�#�N��] [ ��$(����T� ��HS
�8�k�s�y��t�U"�m�a�x諒L�ű.X����6 �;m���	�^� ���U +н?�	�]��00Q�ӹ @�є�)b0�@I��# <�{~���� �J1�k� ��5)�|­ �@}J*O��LV�W ����k���n
���5�Z�� u�MW�I�����J0�j��\�-u *�?�,�V�� l+�	�W��zn|�x�] _��'0;s Z�����^H�� �h0�C).�@D�G���(�Z�k�ԇ	������ �X���Qe �~����k� =^/.�� -�
�d��� 8u�R��N�� ��2�Y  ����Ke� ,V��Z����CӉ�P3�/8�R���?�� it_*�E^ �/O���� ��ז������=9K�n �p P�f���W/H����0	Sw ɕ���=������������Z-�� �L���r�8D���M?��P1� ���Ϊ� �f%)�}�� !�d[T-�l./Q� ' ���@L2����F��1E|�̈p���� <0���;��f�PK��C�d0���5V_8�$!��*�`�c1-r�0�5d "2Y@e� ��M�~��� ��t��0 ��hE;	� ^�ҟQHo
�?�+`��h �Y˧!��=}^��H�� �UBЌ(N��	���א��7� ��ߔ\� �-|�N�h� �r�{~�� Z�)5/	$e��8 �S�f�� �E"��?n� �8}6��� ��KB�/���"�3����h	�.\��8����R�͎�-�+h� ��zJk@��Pa�h*U�������b�Xɵ{ �!�8?��* �1���ZƝ`pw�p� �-����(�� �]e�'Y�T|`p�
B��>-��kzi �'��������,��@%���:0� �|�2 � �C��VT^� 0����e �o[(�Y� �h5g����1 ��(�T��xKY��/ȹ�� �h_�Fu� |�[���� <�1�tRO ݨ�a��#z��j �|	Ӿ�Mg��]��� �^	��� s>��й�K,	]�����!�v����� �s-�jɳ ���[��	�9� -�*�)��;�ǀ@z��0d
��R�^��}� �M�">�� ���!��C�#� /������=;� .���X�(e��{��1�  �Ƞ���% \���g)�� ��X��5>�* ^��B?�L; �uk])+;ֶ��-��^���̀� _f���7��� Ǹ� �K�}�\�D� =��� ����ۅi� ���%MXӬ ��H�Z�� 仄���^� S�d���x��8&��	
�~|Rӝ�3`��V0 �t�o�%*x~�2̴�0͈z �(X �1� 6��
�7h<�d���u�nŀ�v	���
�>����5 �@�:ʁ �~�
�$�� ϰƈŠ�zw	�G���� Q ˈ�� �#���� �������H7ɠ�]� �EF�| ����H� b�C�,�� aT�J1��� �P'0X�� 6� ��A�H� [ɔ@ׅx�T��Z�	*�[�Q)w�� �ܵ.�� �_pH������[���Xl�hu@j@�� �؉0�� ��T��:�d^|!����B "M)8�Q �/��-�y�k|���ȶ� A3�}2,c �닣{� �@&h�6��	�� ���S� 9k��ݡ?q�
�� 7fG�9{� J����� Q�y��P�2[Ġ@� z� �I�)[ "�:}H�J`�з1� ��8Y3/!� PA�j����	�9玀�3�� Eu4�R�� _�ڃ��H �/�t�b� �_�*��� ��ϱ���G���.�� !�߸u�*� Ɗpn� X�2���� �q��SŃ��R.��1౳,��Զ�� T��.�Ć Qq( �Zؗ�/�f ��&#�x-9�Q����S2A�@KL� ;̼�%W�N ���������a�S��Q���@֝ �A}��+ ��ˋ/ �`�������V���̀Z �� ��w>��v�����k�v�x �0ο��� ����*� e�z(���,B!�!��)�_��� �N�� �^��l�~� �2�{
� ��|[#���:@,��� 	��J[� ����<� �����Z�z� K�B˜R l��%� 2��J_��w� ]Xl4�Ƃ �q��W�n�`�]��e_�/�@X� �)�Y��4' ÖP�!p� v�>`KJ �§0�hw��C�A ��e� ��h�#	�Q��Xn�_���b�1>~Z�'���E %�u��I��H4-�����9	x��U���q!/`n̺ /��0�L����B��@�X�?���P�D� �_��{[�� w�2��c�� ���R�Q�~ 	 ����_��
���*���H�� 󔳀4��D鄉`&��y� ��L��L� �>�N+��B���.� [$�����C��j���` 
�tX*� �ޟ:\b(u 	�Y� � U�존�`��k*,:G��*|0����]�ۘ�� �4�F�-�y� �x&�B� �AP���>� ��T����Ä�ؠ
r��B�"�s� $� ��>*�!�� �;��:�E�������&�� �|HŅ,� �\s�x�p g��ް���0P�[�ӻ��\�� R(ٺ�HD ��J�£! �%���� i8���.[4�� �^��Y���{�l3�'c�0��W�A����)�x� ���\�cd
 �s����阽 áxHh�f &3ӚS��$ �"V���A� �!F@���	[����
��*��}��  �PU ��T�Q1� ��#t����Ӡ$J(�ϷI(�� ��-ku$zSO̲�	�=��#�[�,x�0�Y� �0@�Z��Q8h2:;���Pn�@�}� +d�����W A��%�)�h �����;$�^�� ]c@/Q���T���Y+�� 3�vV����������o܊�T�1D0��k���e9�h �&q��Hb �W`�BN�[ȯ�&�rb� f����.��n	 !��� �ֽ�?E8� �s�y�� �0� ���˦�`�YW �Lc^�� ���;0"�g ��E`��A �{�56� 3)#��������`Ƀ�U�$I�|�^_ �����h�م(/ X��TZ���fڠ� �\��h�L �fQA�� s�,��=� ��&��J	 ��_QD�� ��%ہK ���݄ '��4d�"� E �x�ס� j��J��� �����F3��@1�����W f�#�������%Z�J1A ��\a�og������	�����`�3
O� (���h�9 �⤈�4c�v( ����0� ����Di).��� ��S���Tr�J��c� $'��V�� 1|\՜ek����� �S����+�p� �	�V��[sp� ӬQJ���		�#�pȕ�x`A �h_8�r*蘑t�G@q�J� ��0	�X
�{�/R��B�L �����}�� E��^� @��%�����k_�g�������-�!0�X`�� ���~��x!���.2nȽ	� *�
��8���� �L� !�;��H.�8� R��'�� �g�!)1�o���R �8�sK��� ��'��(�\ #�R׍�Hc�L�	��X֠�� ,3�U���/�x�ĵp�� [��)�iU�v�L���3t� �� �|�2�� ��I�Y~�H,��0
�`x�� �!ho+�8� E^�M�ZX�X�WC�- ��c�*��T�������U0�i� 
3�ߣ� mKB�Qx5�2؀�SP� 9� �=��0�_X����@Lp# K�t�UQ{� P.h�)�� ���e'Tu��| S�ߘ��׷ q�Y��]Q #<�Z���b�`�^ '|��� 2�)@EK� :����U�� h�a�/�� ����	� ��KwF$ :R�d,����� ��~����T+�G��fK�9 R��I�U�8;Ԁ�5���[���Ґ� 	 ��V�-������w��Z0����
� �πH�@�� ��j�X�b �K�Sс�MD � !6\BH;"0 S��_/�� |ؐJ�1�>��~� L�T�	�]����V�S�W��� vb'"]�?w�i	�L��յH ���-D�"q.iQ�J	�Ю���]{ ^�.t�u��#� �\[Gz� �@���� �XQ0�� W��s �Y�I��}�Ph��!ъKx�^�B�~�${�t� ����r�>Q� �p����C�$��`K���/�×t�����RǠՐ� ��x��o��1f��X@�-+)?�i��Y�xA�5`d���p>���W2�P׸[��<�Z���:����9 >uʁ7��0�2N��J(��Q\��;��CB��r !^#�%�(� V'*�Q՟�$}�q到��T�� 3�fXw Y �s&+S� �1�]043��"& �����@�<�8�vtެK��W ſ@���ϷK���.����@a{�z".\Z�VDO )Ѯ(�z�l+Bտc0�� �%�"���5�����y�%x H_OQ,) }�Ұ$^9���Sq@eh�T�`� G̃�u7���K�{/=W�.ŭ �չ��SVr��E-@���x:�)��(�ǀNY��]�/B�rP�_��X��ưmL�5S�/�^ �����t��J �ړ�_tH�� n�y1S�� l��ZQ ��[���|����Kd/��.��
��x�	��)�_�Y̴����� RU���`��H��{O^��s�M�ot�0Xv��H@˘�;� 5���[! �D�M����
]�`�T��v3 vI����gkA^���@�h0��%�)�_�~U�� 6@}���� Ihqa/�x�U��	�'��[������@-��� B���m� �=���Y!�<� ���@��(ؿ��Q���À�K	݂ uwC��q=�~� �!Q ߃���(�q޿���Д		�T�\ W8���3�F��f� RZ5����1��� �3�_�  ]�&����|y��v} �H�J��b ��� <2+ �\������ �B� �)���P��LY�O ?�� &E4ue`9 �*�R�%��vS�F��.����y,�� ��V	��u` �^2���0����k`<b��IF���2 ��	7hc}Q ���(� �XN�p���i6��ߥ� ;����� ��DYz��LT( ���N� ߉юSt=����*3�): � ]�ֹ�ܝ��H�ʽ�� ��ӫ��, �[��Y] ��Uj��-�8�p���Ӕi. F,�
�V x{���K�� /S��f�� ����2 1x��ӊ_I���!~[&л�j�"1�; �]�'d?� �0@��Y�)���<�I�	�� �J��HW|zw ��
���� �Y�y�A~P([��ڀ0�1 �	X'�� ��˧PF�����Z����:� ��:��d�� 2�-�A�:r� ^vtW%u�Sh���5@� �*+��� �<�bV j�wf� �پ��I^�V4(;�# P�0A&B�$, � �+؀����3�{2��$ r�^�+0��ⴹ�s ����р�&8�� +���� k��	1���Ь+U�� j�)�.]0h ��c0�i�` �����3� >dX�Ψ�� ����@ xK#�	� (!~�Q�3�L ݜ&SÒ� ����\�� Z*]��3 ��9�.(�  K�zW'Y� U���1��� �[���L�F �cg�G��U Y0�d��@rXŉR�������	����]�� �}_q�� r���[F�� �E�>Dx�9�� #\|�_5 Q4)«��X� ��A]=
 sF��N�<���Vv�Oc��:�	 ��qY)�?� u1�+,H�[ ����\� hz�4�����< V�ǮPO�� �0�	%� N�@t)�����@eL�]� �b��x��?�� �A`� ��ƨ�P�� ��hr�� )y��R�	�k�!�A���M?�e �j�J�z��Z��x��t �G���� v'���5_3 �,�  ��ߋ 
���aLV� цT��O�  �)��,���_�
^���`� �g� ��J�}� ����/��yh�\���ʈb��~#E� ���+Vf�� 3��j�p�{� �±�0V� �L�Gu� ��b7	�;�� :�P`���@�Q��A'��ob���t~ ���
_�e? 1΢�ĆӀ�� ؜���A�n8�^��l�#�� f��a��=p� �@8��,	 �$���w �K�i��,�T츴� 麒;�� ��I�M��8�r _��� >YU�}�P&�< ��fW�|0��zX+���@�J�ds���y��'Aj N��7�T�c����%p� ú0^1[Ѥ����w)* �zS/�� �������8���X�����,[ �fXQ_F��Y�$�`�k]�|�@�QTKY0I��נr ��
3:ҁ��ʄ&Y� �R���@�PfDbk�?� #�o� LYd<�� Z�{��> �7�w���� ��A�O� PB��x}N�L��� {hlWc9v��xA�I�X� ZUT���� =�H4�� �7���� �D���/UN�5��� � ��ǝ�$	S ]�(�N ����B� �����:� �
,C��S� �	�1̇���FXn���y���г�Y W�SP)�"J ��,�EH�8_��Z{�Y �L!q?�p��.� X�P��� �ʁnY1� �+�Q��zJf��ݦ[M�H�EH��X8 B+TJ���m`/r]�2��=[\��T�IW>���� �^��y UQ���q5	��P r@G ����Ӱ� �w0Rً*���% ᰚBtC s��ơ�Y /�<\�鬐�� fk���xh� Н�6��
8�� G ���Q� 2�̀�yk �[x��! ���?_i��&nD� I��MsQ01�w@�%X	� O�ACdY �/��Α[p��cG���ܖP� iB͸O7 !�=��)��]/1��Ah�T :�S;�NW#(�����*���ɂ��}����= �����m�C	z�;ˆ�1H+& ���p��! �� "��E��)$oA0� ��_�hi� �Q!y� Zb��� 1~z���[=_�?�� 0�U��/� �a$��]�W ����D�Bv�V �p�[� �� �1�0a�@�@.)�/>�� �+��X;� �)}����>
��	\��: ��3�����-t4�@��ï]c��	W��� _Cܧ�X��¿��J��� -؞��` !���^|#��H� v���[/zK����Z3�D��p,�[�S*���� 4�9�BQ�DX�����  �(2N�'�[w� eP^���, ��-��� �� ��" |�U)�� ����VR� ֥�	05�t� ���>�����^ 	����4 J�*)�<]��	l0�! �^�@�����J� ��� � I��0�RjZ����J�za ({�I�S�0��� ]��?LB ��V�i'n}��3���������D0�<j��h T��Q��� ;��>���� �(�)p�W
���$�S�� ����B���d]���?���CK� w�`��W���n� ��)�^up. 쵠1��� r��%t	k� ��i~�mܻ }[-�G`|s� @Z1�I��0K��yH�% ��9.�|;� :�Z�OVC �P����;�x�(�hn/Y}��F�Q@|���H���H�b�R�&FW�a�U����!�*�� Z���� .��,���a[��(�`6� �A����]8� �dh2H� ���K���C>��Vh3à��x ���%]���y  '!ū�����~
�ą��̐ ��h۷�/ �?.���$Y��# h�Te 
���!� A��PT 2Ћi��� ��h(%��&z�& ��1M< �O�*߉ !��\94�AKb��]�
�ܲ�	ю`�k >�+,�w� �JM��ڈ���@e0� X�!�S�xc �:h��*-�L�` e
��1�z�pcE���H��_�}e<�� o�|U�� ��`��e�&|)p�]�6N��kŁ�G�`���Rh�,*�^�!ȿ_���� ׁ3�*	H�� ���P饿 |��I�S �kb�{$ ]�W?N"� ��O���z�� ����� ��>L �Z �h�B1w��� �%v��2��<>-�n� ���5h A$J�Y�.X #����?@ �㚓)� >O%bR}ȱ�Ϻ���� �܇-u1� �*<�"� C�[W��<S~���Z!X�� '�"TguN����1��9j&��� �X(� ��B��-c�l% �r'ߔ) �۽��jn4[
��1�/� �l�xJ� ��%r�H�_ʶ���t��Ѧ���ȑj ��`����Ʌ 8Y�" ����L�
�u \h�KX�H��-[透1ȹ�ew��	�؆���� �UT+�:]� �^�j��� ���W h�3�p-� �dN\�]�@�� �r�T)�� � NW���YHL^ 8E����� ���� |��
���� �.��XJ�t%��xs�^�e����' I�|�r`3�� ���{��m ���#݈�L$
��&X �~2"�6\�zA�ؿeM̝ (�}P��A ��J�?� ��ٴD�� ���XB� ��U�N�������]����-�ж�S�� v"�FJӥt� cy�<�t!] �鷶
D� ,���"���HQ���P����ǉ��6�	�\ ,��I�D��;���K�t,���#Z�[�7��W�y��JR� ���]Ze@� %�*\�-��3UN��K@��7�,R��> �\  (B�W�+�u �)}��qc{@f��h�? Q<�]�4 Ƃ��չ ���R�\v� e�'�ِ�(Ⱦɤ��`z& �>����^� ����[�hOE�}@PX ��:SN�L��=^��d��_�,�з&8 �
� �P�NY��� �eo���:���۴� �r���p5 _4��@
�� 1l��0n �u���{����ǻr
�U ^�%����� ��/�F�`� @3� =P냈�i�à��� �9]d�w%�8р��zظ�g1@	6�O��`�v�)Y h р�Z�� (V	ϒ��9�Q���3��Y ҙ4JI@;�Z�!����� ���v�/6j3N ��)�%hf?'�@�܁/� ��M2���.G����@h�s��J���B�����u ~5�( à`1�#ȉ<��I�ͅO������
 �D��/�l �{	����\>:t��`�[-)|� ���ob�� hu��ޢC� L<�-8w�> �� �iR� �L�؀�f ���.ɏ~� �P������Pt`{D�Ʒ �\(�h� >�+B"�SP�wz������DE%)�]�'+�r�c`���0]� Ѯ,�<y �e?u=�҂�qI� ��Y�z7�- �����g_����W��$�	@Ӻ�sI *���R-�8@X��8��O�( o���\P� ��9��� ��ɑ/�{ �� 3�_ ��b]!�\t� 2�`i�Wg�Z߀p��'����� �#+V ��Ku� ������^ 1�nR�t� ,���E�=@�  �e�!�� �ɭ+���� ��ܑE�pN1M� �[�@�- �0�v�>s� �U��q��R�[C����� ����K�� -�\����������3� ��TYt|A� �H���*i �	��߀ nY3�!��/��(�z��@h��C ���f4Z5���������D <0��W /��y�)� _3��p�5	�K����8���A
�� ��	��d: ���}hq� '�f�lZ� `��[�*�� Ք������w�ֿ`_��2��q�X`�;$�&� �2��S ����[h� ؝�p�,�{�� ��A����LŽ ����aݰ[]6:Z���*��� BY�. Q҉ gqp�H� ����$\1� K(�U& �v\b��X��J�p!��듺 ��̀�� ���A- e� �h��<���v U��]�:ur� }��� �nG�"�
 fUzoxZ���� ���_c�Ɉ�`A�N�� �%�1�Vz�(�� ~
Q�� ���la�:bL���謵�� 5y��lT� =�a;�� y�V��.� ϷB�-}� v��K�L� �Q@�MAԧ ���(�� |	�[ø� �0┍BZ�x�y �A��� n�cӇ�Y^!˴=���v H)�EW�' ��_�^,�� �~��0 �p���#�|+&�4� ?�˺��,� ʵ����� #�(��� �6��>Q�j ����r � V`�(q�� X��%�A\l��<�透Pd2� �Ze�5[�JL�QhFO2���p�����@�%* ������ ROp�ᘎ``y8�1˗� -�U�e&�c ��N���� >@f�~_��) Ƃ�NZ� �8[�؋�ԆoA1}#��=�@ O��W���^	� ���-'x� �����3{ Q�~LY6 �ш�j�<�|= ��H�������� �;�)Ɓ� �X$!� ��H8
+�� ����`�Ox�$Ϟ� �	� ���CA�>^��gP�h-�Y���� �d��p�k ��+����?X �f�����%���,dZ���AF:��	u��YB�E ��|�.�f I3�U@�j c�>�dp`? %��6��5D>�Xs,`~L�� �d��0�>s��g ��_�����&	�� (����^=0=����D�!
�c,�@+V�(���a`���0ߧH��~h<Z�8�� ����[�G,	_6 2`�� ���\�(l ��xg�C~���Oj�� �a����h7�#�B�o���&!øah�`v;. �ۭt���8yC�������h����R'��D� ǿ��,�!E �+����45@�},� � ��
&���/ )#]��@U �ʗzp�� 'w	��`&F�?�� Hi ���1�` �lC��Lڢ &sB�O}��Y������ �0_��% �G+���- ��Ҁ�}u_�,�K�9���� qQU#�:D3Z�K2����u`fL���+*І  �y�k� )��[�S;��>2 _�E��z �u��S\�� �ݛi�"� �Tؖ]I( խFɧ|�xx ^�ϨZ� {���,�a D�5�V�g_X0w!v��p�J����8��s���U��@�l�[,���bc�=�p�� |�K)�T?�� Fw�f3 �05!� ʐ���� ��q����U�~�����P�ʆb�c}�@o �-z��'��  �H�+/ h�-�_�I�tm�	����U��� ơ�@��Å�
,�2 �VwK�> ��^�k� �r��P�m ߋ3[)�}�eAl;u� �=6/v�!I �{��&a� ,0���ׂBQ�� �U��IpL��6%s�� C1���5Z�ǀ�����lf]�`P� Z� e��Q���[ ��ܙ�� �IĶ����o� �)�GP�# �z�/>�¤ }�� �X�� �_��" �%��@�) �*�ZS� N��:!�� }���P"�T��]@U�`(�P���:�(D � ��U+ �iP��#o5�7 �'�b_ *�^���ˀ��� �_/��	 ����.���A�<�,��z m�e~
Y�� �,Q�d8� �]��+[� �%��(�^� )4i�b�DV �h}�N� ��̮�f� 5�BC�� *��9a��X�s H�4)��-��y�P��� '���+ s$	�`G �K���� WĴ�ۋ �q�_eb0`ո��D�� �F�J�� �<��BY^� �d*�-�,�K�8�+���k#��0P4�&� ��Z)���{�_Q�i!�,�� Jk��+ ������;� 0*���v��o�WӤ�R���!�m�p�	�e.'�*`�5 "%>�@�� P�'�y�� F���W1� 	T_ �f���9���[�W�PH�� `E!1���� �	O���G B0��b1�&S�\ ���NX~�	�R �Z�$ܤ� ��br� ��)��E�xt��o#�V� ?���	~w� ��^�C@?3� ���0� G���V�&tA| ��W�� �/|vb(�w	�{��!@�1�+ �s�S��8~����� � a��d��h [.��TR���3�AƓy��q���� �(!h�= �dK��Z� �PT(�`>,zMJ8ǇZ1��X�a�'�g�P��^���u� +��	�� ���0�� ���B��J`	轀V� µ��^: ��X �h A���|� ٞ�u��(��/��p8Q 0b1��Y�! �6���	ɨ ى���S=��F <N��5�}١�	2w�ro�#��h��� ��Q(�ޢ �}!nS��h�6C)0��qa��R�pt� 1	���`H~ k���f2 3IP��\�x  È	�SetP���E����%�o���� �(���~ ��S��b�H� 5����^=���\R��H�" ��`-]�  7�����O�C v�\� D](��[Sk�Y냀�hùP=^r 3K9�� �T� ֝ |;���� ��[��oA� �h
& {� _�VJ�� ���(�R ��Q�5�T� ���K�JX<�ଡ଼�� W�=$�#!�_���s�NSL�~� �X/��� ¥]��\a ��+�;Y���p�b}���' �12�Y�nՐz�_��;V
����-й� �jQ@���vZ }[���1 ¦�ug� À����&M�� ��3�(� *Lֵ��O x�-T]Yq��� i?��_L SwK��ϲw8 �h<�(��0��Ȩ%�e���?a-��x�i����~W�ǜ�
���� *_8�˙��ͻ ƺP#��j %	���3A�@�a�{�� m�B��� �V�����r�W0ٮmN �Z̢� _��Ł�>:/F �K� }� �]a�.��Q; ��(����I*�~�W�@��p ��^��}�쥐[ rvX��Ag<}� �+�WT�x�y�	�2
��� �t�%�:�8 ��A�(��h �;����Q �>�E�Y� `�m@��  �x1Y ���W	������7? !�>I� @��]�1 X�� �$c�R0��)ן���U�����1� �[��W�jv %�o�Us�Ǥ��ʋ��☭ ��GQ' �� Ah$#K�[Xq������ 0�-�w��? Hˆ�� s�AR0���෉����Ϻ�]>`Jг>�������\�}��1�� ��S����*�x����l��[$��a .�IN�<� i�7P'��V ��z����O �tM�`�\�T ��*� �B����1�?3��[� 	��@d�:U���n�.�Zg`G��} +�>�^)p���Y!�
��(,P�=	�8 ��o-� �ֺw*� �H>�5Qi �X�<�AD �ZO#�� /�֕~? 9C���`d�\�E��l��Q T��Y%+���i�Ac��" /�� y�ګp��`��>t������)�A8�1[G��!�����X8i_|��-S h�5���� ���7^/ ?
�U �&�)�����%]� .�W�E��kss 5/���- C<x�c 1��� �KX!G� �Z��h�2^�  �%H�B��E�И��`t�q ��SX՝� ���	���W���q,������xH �~[� .� �w�E� �Py�,Q[靤�X��sP ��
_Q� �K�t:�Ğ 嫵��.��� ���!M���n ��C��� ��:	Yt���@SBػn&l�l �h���K������� ��ASW[_� �}��1ӵ ;��S��R=�� [#Z��j7s Y�AP^�@���(�UAF��\d%�0)��B�`�>�l�0�Y� �fb.1�s���y��N�� z5���Ud ��ȱ� [YL#:'�P�=��������������x� �KY�H�|� ��/&��!ـ������
ndtѨ��  L�Դ4��_	�Z"ʂ |�@����8?��	K�f ���@N�}� *ҧ�%tb;_e�����`j��S 3%��-�@l�h	?W� �=��B�|Q �[�0�� ^�Y3�Z� s���V�N�	�"�R G亙 ����N�[�X������ �0�y�W� �*���X� &�$x�� U�J�cy�!�o����)C� �������� ��T�k�8��; H�XS�� ����V���\�� ��/#O0� �ʢVK&�:��>� X��Ґ  �fKؼe����n�r ������X�}@ �=�u,!� ��r����/��
"ǐ�@�dQ$Y� ?b|��Z� 8��Ih���v?z��_3��ʨ� +�Tb�V:S��-��Q�� ��a	T��
��l �w����5e_�īU��� c,3���sq���Lo��J@QWp����ry���.�8��B���� ���T* �]�s	�� �u�zx�J��G# �ʿ�0ZY�ph�HW� �&�B�s:t� �.�ea��Z 9� b)�� h%��	Q� ���Ol΄ �1�"����_������ �i��Xu���� @�3�h�	� ��,IU���n���Q�=��E@ �g^� !o��:�Ma �`F@�-���P���s�X� ��ov���!���A��S$��`���X�����e(]��~"�r%�0��r� 9P�'1���� lF��%�J 5Ö��ր �P�Ҥ��� (�X�{�6 zZR�2ؓ� %�v�Ϝ�� "�����0EV�1�U�)�;�\
��� K�?����L�: ~�B!�v M"Z�®Y wdebñ���Fl� a*B��:���ZwN �!< �T/��)�L�� �ы���W�� 0�z���S ��*�KR� bw���uq�%z<��y�\ h:B_�E�$���(��[����>�-܅D��SU�}a ��6� ���t��m0n�͸�E��t��p�/  �T�ֿ,K�ǹ5��� +�b�ԃ�� ��ۜ� �P\��i� G�9�0A� �Ԙ�=�jD�@�vP�S�l �����I�[�`*��L�� @Sɻ #�uPT����\��� ̃쑀�z��v�� ��	 � X��<�@� ���kT� ͋BP�V t�0���k����g!ŝ���`߰> '�W��� 6�~3e�L�F�E:��\9���`�' ��Z1Y��=�V %�����Sp( ����[�����O��@M�~�P���0ؽ�c 1��Z?u �����K��0 �Y6Qf�h =�%jE�z 	�RU�<YИ�Z3����%��F�4 �? e3��� ��7��D�1�!�#��{�R���9�|띕e>A�K�D� 1ӌ:-��� "�o��ZS �J��r� ')�s��I ��>���{���(��-P ��%]����[��3 �c��E�����?=\� �,c�8� ����_P� 4�`$��ʳ|ZY��W� �K�0 ho(�T�a;�\ 2`α�z� �51����:�k�d���� �g�� ��LXL�"�Q��sp� �6���K O���:� �L}1�=� ���\��  38?�D��W 4��ڴ�[ �_�a�M�*��K!�. zБ%�� �=�]	�������0�b7�Ø��QZ ��Nō�����X_�߭[��+_����P�k T�<�`��H�S@��y�&��W�Z-�{�[�0Ho���R ����YPa}� ��/�	W� ���&�!�L���� |Y%(�u&��� E
^b ������S�W 7�$��� `��(ݝS��[ ^.��Q�8 TK���~ ΃��B ͉ ���^G��p�.Ѡ�X� "����`r;��k���J	Y<�7p�9fץ^�0	 ����\+*� ~[u�A{ ��'��	�6 K����!�]�#πL4g�U ��q/�Cؑ @�A���+�
8���w] !��j ���y�#a�v��г�2�(� ������� !��>_� �x�*�\���L��z�O  �����q �h;lqz(��G�����b�H��
�h�� \$��)M >�
}�՝Q �`����h��Y��Z��	a�}�7� ���
�_;?���hzK�� �~�'W  �)�\�/���� 0�f[���� �ւ葌�\B� �!��	y�H\�X�bJw�a��� ��Ŋ��DѪ�(�]�v� � `��ͩ� �4&�R)	��״�Zu��`�%��� ��{^
�r�U��a;8�(� �'�����
 Y*���!=.ihT�AWl7p�� ���hQa- V0r���*N "A�Z� � x�jYٝ����� �hlD��� ����-���~�G c�/J� ,��[as�? ڀ�`�4����ʚ�< �(;��z�=�_��Ǳ��6� �j��Oh�_��5��b �K��!Q  �~���@>�u�� ^�+�jy- 	�V��[�N EY��` <�\%
�6� 5��R�{_-#�n~`��r�=Y ���$-� ��E>+A�8�k�w$^P�~��/��|-A���0f� K�&�u�� Ll� |= P
�W�R�����J���������N�@	ڐ �%3)�_rY \ޘ�[R���  ���bG%K��;��� �f��t^!�[��� h7���	v������ɸp�P �W(��� �K#΀��!`	��_QUv 4����� �ج6��1v�ȅ��HCB0h_� y�z�XR. b�[�J!�)G><�XQ� 0�S� ��sb���>� �VK�D�� )�!����`A��_k� �t��/�@r8��@�1��'��x;K��J��q ���b� ��`-������@�,UQ B�/����  *�bY0�XHʌ ��[�G �Av��f(!���p���J 1�}~��/q��N+@ٹ �X�t��.b�)19��q�j�X% \��QZY ��Ȃ��}�	�@"e[�`��~�� ZS�� ��!6�TY �����kC ǆP��+ 9�>�L n}��#� ��\(� ��ѺR��p� �_2�P� �d���s(.3�v,�K@9�p W�̌T�� ��ѿ"D) ��M��1 A�j�Q0L�P ��UN ��̄< ��`�0J� �I	f>��\�~ '%��� (��Y�-h�ϛ=ڀ|��H h
��zb -���s� A*`��w��hX�D����:� ."�	,5�2�]�`�� ����Q}BI9"��&Z��` V@P��M� )�u.v��Z�D�f�� � �":��uƐ ɶ��� �w�K�f� ��^	��� �����J ��(=BXŘ7(�7� W��SȆ0�� %�ր�#��O����I� ���%����k00#�� ��G��;^����,P �c	4遝X��$W� ��)ip�_��}��p�� {�� �: @�8J�� ���[ �K�zĔL %/�}5J� �<\�� x��/�0 �Y+��Pp6���}Q ��:�vR~ �A���m/+�� ��D�R�� �x_]�P� �K�{�Cu �L-J�Y� �|���V� '�c_ ��}�O��@0>Y� ��Z��LP�ag�,:���@;!y��?�%��k�����7 L�P���� ��"]��Mo7f� A'U��� �x��0p3� �e$�����	I��u�� ��j��^�>�� ��0
z� �\F�$�m��X/9�Q0XS ��d̅}� ��	��Ƿ�`��!�*Aq �����)�s� X
�JY��w?!�Ȥ� ��*PY�I[ #�Ba �� �8��GP�� /�>V� �-�\9���~ �Y�	L}�Q%���d�b���@y��) �8k�� �3+��1Ё���H S��h 8�_���(���nZ0z�� �3����Q �["���:��p����$���S�}(������ �Y*�d�^� 1U�?IL�׸q*��8ӹ 
[H�@�Z ��}c��� p%g�ߗ�� ����	� ���B�!�o�t-�l�z� P���
��3 A~���f �E@	i����^� ��_�� \/X[ 3 ^��D���{* ѥR���� ����6* ��o�@�� �
S���2 �|b��P� V0�1�3��������) Q�"�&����`� ��JW�	 �:5
�HN �#�r(���z�8��SF�1�K ���t�n3 �,����0���P�ʵ��$ВX ϰ�ݺ��lrx�Āґ`�� ��)�^�Á�� ]�$R�Z�8�̇��DMN J��� �����& ����%� ��Xp[��)�(� ��0���d,���1W%�E`���F�t�Pl�1�䠋��ݵ� 'h�BHv>_�� �P1���F ���M�0���2����R� ��g&(!��I��»\�� A�	VX &���'s}�Q �n��_�L )�L:'�/{n����[�"��g�/��ݨ֠�!p?1�\���Q �'D��6 X�$�l: �dYS�� �W��qNj(�m� ��hZ^ 6��V�R  �BY?&� �_1� � ]��h�+��>@������ �s� (Q ����G$=y ?��}��� H.Y(�3	� 1p� '\�j G��;*ޒ��� �z��,��  0e�N ��&)�3aw�˧�`�5+�S@�F�� u2��w� �H�*�JspK�P"�í2����:�H{Cs�# �1�X��t��e)��3�] *��(:�/��<H�0���&��X=�fA��*$�_t/ ?,4Ǆh� e�@Ws��] ��;TBoi��)�ᇉ%��I N؍��!X��3�
 	ѿ�f٢ _!��P��� g�df :�}�%ȉ 50ܗ !��{�� �xv��[����	�*(�U�z� ]?��.�o�	����� ����1�un
�9_�~�� �	�U��/�u�|�o_@��;�g� �T ��`&� �tÇXQV ���lؚ �h'8�J� �s�+N� "�Vi��~�	] dO��K�� /R¯� �M骚@� dP�v�V� {T^:��r\'
�~�c��˶� �����< #j��sh4 �1�ů�� ����IS�H������V)��tB��c
0 d���s��� ��Ne]� ����,�R �: ��� �f{�~�>[@G:� ��1� _P���T�H� �ar�{' ���C��� �R�&�>øJ��ف!�hWn�)u���]Y \[�9�o������ ��'�zX��>�� �U��¿W_?��$��y +�e!�Y.E�l�@f�} <�A/�����0 pҁ�`�CV þ��LQX4��Nq=����V�p�L.����K ��F��y ��j�8lJ ��
�c[ ��ٻw 02�/�� ���P�L� S�D�Y ��{�"vFX׀#�wN $�	�C� ������:�) ��.�� �X��S��)�fQ>��՛. RpI�!N ӌM+J�� fL|-`�4��� ���?���� �� %	���jMߠ����F|
���S��� ���o@k0 �;��ڣg �şH	��D��%j�h ��.fݢ >�_��̓
 ]0��|M'� !C����W(ݘ� �#�Ӟ/ _,�|^S�~� 곓�� ��m�X��G ������ K0�@F4 ��J���(�V� e@���� �t 9T�� �)݂��a�(g4�0�9\��Q��8+W; �(��F% ���fh#� 4�Ꙁ��� (� ���~� �X�V��9�1�J���r D�,���s����+��<$ �k�A
F� ��!� �	��PW�X�2 ��@`�	�3 �J�-��b( 1�,%�8 ����{�6<�G�p*};� ,3��0��)J��ho%V3b�Q
��~����Ik4 ^���_���u ��.aʋ�#��@�
� [����~� ��%G�\q �㮛��^�h�|� ��`��(x� ��̀�
�T������V�od/��\��u��pB�:�� 9ʨ�jw+���u΍o�y ҉���± �nhk Hޛ !
�"��v�CqTh������<Ƀ�1��� 0;�ht�p� ��'������������p� ~�܈Â�К t�� ��{w�2�m8�� ^���Z"� l���0���Na�A.���X�� hy!�x� ���+k� xz ŋ�/L �#h���4�{N �����,1 �5�����h6�*d�Q��N�`q��	 "�Z�~����d����@��Au�=hr>UE"�z7�	��ӊ;^���L �J�& 8�P��@� R�y�#�OJ ��8.� �����9��}b�_E����
|� KA!�^���: ��i.u�<�{}���h	��XpD {hzF=}5Li� 4
+�Pbf �N���o��]�!)���� ��%�̢P;Y�'@+D�h� �K�&�X;,Q�[���/� w�����a���"%`���S��T���`M&�,� �� ���:�� 	MQ���7$�r���`
\)� !�0�>��ED{��3)���;���	/�� ����=PN]��H�> �4��� ���_(��5e���Y�?RO����Vh�~���j𲘡Bf :1� ���L�9$��6�l-� @�y� ���<?��0��t ��P_�J� X��H� ���̷~!	�u�w%&���|Ɓ
˻0��=	� �N���8�� #�1��Qk ���+��5r- �*����X�� I[S���B!� �JpU�������� ����D�� ���A�� i�N{�?	.����0��%��� �E���e=�k耝���b":�$���s� &S���W��� K�
u�! k����#�'T�7ZD���	 C�)���< ���6��1� �r[� .��^	 2�C��[�h��� ������� �%:��$�Ԁ"��]s@��R��*S� o@�D �>�#�&	��d��-�P�O� N��y�� �ܥ��C�{ ���sЀ� a/_3ޅ�  �ﶕ4]Q �iP{(%�X�'[��@I��X�Ց�d������% �(�Q�O ��3J1�� s����C��+!�Dw�{��X3�{� Z��|�	�� ��SË� <���yH
�Q ,ZNB$X� �'�w (��vPG��I��H�%]�8� �XB�S���&�.�0�� ��b�]�ڽ ���v>4�J��Nt�~��h��n_�`5�/ �A�S��? *e���b�� %[�X�P �߉p��Z��� ���Y܀���׵�%	�rk���h�Q� �������4� @	�����  )���׀� �����5V�/� f� I>D̿* 	�)� ̟VA� ��em̚x `}����'Ds/ 	�X�Ӫ�}���W8�P�O�
��?�� -G1����������s> 3���o  "����._� ��C	�� Gz��V����\R������ !�&)ъZ +�\���O ��z1�!��A ���-@�( �Ü�� ��}�?�0P��y �'����9t ޵��#�� |�N�8hȹ�2ܠRM� ���O_&� Z����Mzfj���v �6�^IQ|��x���2ߋ�X	�P���4#��腾��/��2�S `QN�b��_6�'(��p���@S鱠�� ҵء��.�� ȕq�& `�:O;��8Z4з��m0��%6`|�v�3�<P]��� 0H��l� ]+��5�}L�� /���J��38	���V� jE LZ}���� �1H��R )WYX�� ��]jd��  �`�hH�� B�ձ,�d��AF�'RU }��]Jawy �@1��N�D��O��]��� kw�͠Z�%�.QP���8=�蜐�� ��Qv7>e-�V���I@	��\�� ��K��@����`�)�\���)�-[ ���!�5Sc ���	��3 2�[*�^�(P���dN �	=3�o2�x�8��+����4�}�����Ȁ/\��%� ��iIX�0m�p��V�hŶ �����k�j,�B| �&����_�@)`��� �齇[ �/�v�Q��\d���6XPZ����b���h�2 _
�,�1� �ő�c�P-������ ��R�!W� ���Z: ާT�b�S'<�ɩ�%}r� �ŭ0�\� �����p� ��*�P��� -�K���2�J������. S��H;(A�8�� ��!�S� Зn8{E@ZĀR��G g�C	W[�;X]�Zh�1 �-�yG U��T> �Q(�+�������^�A�nڨ�>�
�R �Q�\�#=�tW(������P��*�87� �Q0Л!�2"�Y�<�H $Q�%A� �D�Ĳ� ]'~|�( w/��v��?� c!�C�1�>Ӛ�$�0�D ��g&���8���ª��1 �����5�u�q �F&(�  ����Ƴ�Z"�J@>P��A���r@��S�B%nO.�0q$~�u� �����! ��Z_� t�5��� 	�h�S�?����~%��R����07��
JŔ�!V� ���+�K���~� ����6��b��9(��x���hϩ��ze@��i/� ��Ey�B� l��xD��e� Q��	�� \h����`���r:��XS�Q����r- 0fI�Z� �K݆T���8����"�5F� �����a��z����lP  椴X��J �1�#Ղ�z�\� ���0 �%�
	y��� Z��`���� H���t߫�Y��-_\ /|S��U��h��@���}�g��i�S�*�װ�V�M�2^���,�� pZ�aj�� JC��Fz��P�B���X � pR/غΎ_��J ?���y�v����޹�CB��A	�!`�� $?�1(��̘,
���OǺ< 8� �J׳QZ���b��Rz��-P��b �*���� �	�蠹�� ��_��$` ^-Vl =��;�h1I t��z(��[� Z��F�0� ��3d�x	>���V�cX�2" �ˬx!x��Pey 3�
9 Z�v@���\��L� �J�8�V,"��(�Z营o�D�6 �}�<^�xl���c�"o#���X�����_[��'��A �9�c� e��!#+� Y�:�LWP�kR���	V\����*�K� ��1M�i� ���O�-�` �h%�\��}� KcH��*�&�(�I�.
�= 	�d����'��V���A� "?uz���-�!��G�� �4�u�w0jz�g`��#S��K�<�	��� ��"�`s1�y���+˨!* f'�L � ��,���2B �ۃ���V �;�	��_Ĉ\�3Pm��&9�� @��2 �Ҿ�����eN� �p@�?[���K���49�� O���ػ; fYNR�4�� 3惷-t�8��Ha  ȶB�X
 ���J-� ���,t���[���X hZ/0~���p��o2`ZCq'�D@�\� '�`�Y� _��RP�� U�����vC)��M��#����!� �X�/�Đ]$�� 髄��� [N�����9dh�:A� \сY��H��% P(��� �7X<��� ��4��l��'R�*�K�X��d]�Q0� 1��^{ȏW>K�d�*�� j��/z� �!�n�Y[� *#'_
�4�{v� ���k���t�1���Y!ۋ�+�N��q=v1 Q;�A�M���� �_y?��� ���c��?����5�mf� �ӪS7��wv���]f��.��p�� 	��9h@H4 ��~a) � ���Kh ����*�/t�&�H��	M��S� �U�b�,�A�
�n�a�Q��Ir$^� ���ˊ ��-~)H�� �.U2ӽ` ��!�kOj �'��� \������Z ������ �BO���D��2	��M���%?pP�
ƥSdH$2�=`"��1�Zp� *������	��6 ��K�� ��Y�1��u��>큀��<�/Ba 1��e���� g�	ʖ;��G_x~���=�`N >g��h�Z.|u ��qTj� :�
U-1�u%��W��f��« ˿gw���+ �WO�f�� %E{�8
	� S��G29�G�{�P��� e�G��]�h Ӎ�^?$I�.�vg��[ ���@A�:�0�����J��2��
\ bo����� ��,�	��h���a��(`u�B��I���gO[���w qMG��ه( �ڍ&P��B ����z���5���&�t� ����� �!�X"�P T�ث���ㄜ������6 ��g{
�� G��~��� :Z�0��] �볍���p�JĶ����9�"�S��A)v�jd��(���Xbi��DͼG� �	��_� .��,�(\� ��w�B�	�O�иG�H+9w�3����y�/��<�" ���a�o �`���5 ^$r�z����������� E�2�� ��U��� ��(��R? ����V09�D7�S�!_� ��+2�\ F���&	��S^E���$?�*1
*�Zhc9���| C��r.�-�� �[�L �A��@-�`4�@�Q��3	u��j�P�ğ�!h�_`�0(� I�5�.�O	��Zo��ie�� �(��±� H/�tYZU>���_�!��� �����`� ��}h%�O�8�_@ʺZ�1q�a*����X�`]Q /���r ��Z_od=ፀ9��N��
 ��X�� w�]S�g� ������ �.��h)�
 ���U��3��[�lȸ����KSĈ�aX�k:����q�Cr��	���[����-��{��Wh�T� ݉�a�ɡ�!�;�z[k $ ѷ�� �ܓ�	~�P����y޲����gSU ɹ@�9R�� {��[X�� J}%��� ��;��'	 ��#7Q�Hx�.  ���\Ĵ �L�� ��pAR����<L�6K<�u�� k��.�XU�t�~����w�<�	 �xF"�*5% ���IH�� #^j�����@08��� ؼv���{H�� �^U��, h ��+�C/,N2 0�rt �	�H��j ��(�5�� f��l
{ ���Q�^: ��bB��H �Ƒ�u��FY������ J� #�V���� �B��HQ� =�!"��� ��$k�X� ��h�|�d�  �W�%�-��Asӯv��� ��j�)�3s�� 	��Y�1�'�t�PW@�Q
H ��&�rKu ��h;+� ��OڹB �[�S}Hx�'�e����)� %���G'����u��@p@�~��Ѿꘅf<1�-�vf 8� 0��� ��է�\-J���fs�� r)罞�B*���`�/@y�0�E��fT�l�^����1����ιN���GO�W �T���{�
@I�,	�� �QV?%f� )Z�2�x�~�H9O��y� ����&� �'BQ���J %q���hm�זo� �@ ż �ٹ?�h���T���2��/�5DH)Gt'6(���$W^.��� s[�O  ja��*X� W:��!|_2�H0GÑ��A� Y;��Kq� �߂�eL���1d��0�OSe������ �,�d�5̕�	���n	% ���+q4�C��*�X��R��� 1�Z�`$� ^�@h�Xdk �T� K�A �&[��{G���+��y�0� ����7� hnW͉�� �8HN(�78�� �X!ʁ�qT ��D�P���L��� 5��PK�@(	0� �z�ω ���L�X� ?1$z�؆ 
}���R' �/S��F�1�����n9��)�	�Xf���D� �`M�Ӡ�@�S\�~y�������� 
Q��؈ ϰj��%� �w$K`�D H>"�N�� �ЊX�a �.�P�2 �����U��i08Aq) -�.YԮ�G!P˿p�� ����#x �O���0 J끫��%~ `}��h4�� ���
ÈC !�[83( ��N��1��˂QH0aL ��<��1�P ،�TZ�L H�&�u_4 �F���O�� J @�h&(T���d�g	��;���y��`S) ��$i(�p� 4x=��� W�M>ڠ� kH":#ؙ~ �-h�� ��J"�Y؁�\rj�|@⹐� �8t��
���@.�\���h��S ��N �7^��9�� A�R�� �8�Z���,���?�o
�u'f��hc �Ϙ��X^ � yK��.,��, )�@� �Y�v>��s &�[�4c5R �b����?>�N���J h/FW��j�X&�9�̂t�R2��K ��,�	��~IP#ƀ-�9��� ��	���p
 ���BY[f ���&*4L� ,��R�`�u �������;K�`�5�m ���2�QI���ӿM��y�-���>�х�Qi	�cρ H%R��ä ���hK{�-�n �p�! 8�d/��'��I�@�t^Ħ�����߈#;� *�h�]�?� m���9�� �,����ݶ E�����`��YS��a~V��[2��P� 귮��h. C$li]d�� �|k�0j[v6x+b���
U:����u	Fk �C���E� U�uc+��� '��bh{���e� #��+� �cI�l�*:bm0`�fR (϶�W:
�?����_ ��jX+��>�0���h��� ����:�x:"� .���Y� K��� �R�,�� �h�W7y ���X�J0B9�����K����x~O����� ��(����snjG��h�_lQ\��`+#~�y"?C� �����_�0H(��|�0�-PU��a�b �P���1 ��If��+�rz }4pP��/^ N�s�Uٳ ���]*�� �!�1-+� ���P�ȲsL�fZc� ؈[,X}� ��@�$Mx� �����9� 	�]���j� /P�ZR��f �H��ɤ� ��Ҁ�Av46��� ��fF>-" �B�� %�X�8��m ������.s�p�Q�^|� �?�+�! gӫ�H�� �Y���,z��]�.� ��=� �ArE/
B�]!\P��;��3DI�@�Q	��G>ྀN�8�}�m�耹Q(� k���D3
�e �*#�� ���tS-Ŷ�u����5��ͯ�zM�E����1'�y��V �h-X"����������F���hpV� ���_�5�@&��M�B������*X��; ��(� D����<] ��?#��0 K����-� �Qe�j�� U#A�BL0s�o���!�;ր�
W�| )Ã�5V ��%�C� ־����' ]��>��?&8 �	1p�I�0����ٿ���� &����Ě���%y`a�' J
��q�!�C��47�� �J(�� �y�xN�Ԫ�;+���g4��M,�<I (�thaU����:�,�-Q�F� E�X���?{��o F�%�	��� �6R�+�8 }�'��ٍ� P��D"�1 r�e�W�  M�_�7%O �X�sK�F��
�/� ��Vi�̍C ��T��B7�V�}�_ ���B{ �����0��������^� 3�" ���*�hY��2p;1 �l�X�.��o�N�Ԃ k!�1z# q/J��*$�O[�\V{���1�P �����UNB�������� H�Ž#}�� 	K��^y
 ���pX�xg�����h� *��H��� ��Ek+�� ���\��v�z�v��_J�A�s �	h��|�� ]P��%��Z �$Dz�B�K?��U� �MJ,���WT_�[G0_��/2%���?�(A�0�	�S��Q��:��� ���Mrz� ��Ȥ��� �W�2� �a��?��L��;�)����� ^��N%� �?���n02`@:V1��)���[�D	]h�5���l�)P��v���p1�R��� ��%���
���/�7�g�d "��jB�.£ �a������<�3�Q��X�m�i �/- l��R	 ����\� ]Y�P�� �Di�����3�^f)`�� ���05��� ��{F.�4 S�� �r1��N(�:@����I^dW ��h�%[H �"-��U��( 'h�O� ���&��_S��WR��@�p��� ��?��c<[ʀٻ���?_)�eҁ��M ��q�������U`8��P�-�A�)�(�ʠ������jb3��`�By� H5���~ �p����qw�i �D�J�@�G X��Z��W [й���P� �dY�+Z�|�T�~^���D_l)q�1���Ҭ# S�~JB����*���c=���@��8�� V�ҰZPS �ʞ���� (raq����%���2>�뗪�#B�㨱; � �Y��0 @�R��� ���]�Ju U��8� .���7�� z�Q���?��BC�f��0k� XP��-h�� Vb�_D(w�X�:�	�G �s_��� ]��.� ���[�����>��N?�@��(} �߽�'+R� 0��Ih%6� q}o#	� �@�Wi� �-���� %L�������=( inN�_1 � R9�!� ���b$^�� O�w�aͰ}� eNZ
�D�) ���Ɂ �h �/�-� ��0W%�#�r` ZVQ���P� ��z�: ��8I��h �T½���X��?��#@�Xg� k�(M���.�� �0���>XY 'և�C�U�EWV����%T ����N� .6t-J	GO �L��[�a? �1M
�� �/�S5(Cn �����& �A	
�u!� �3*4�Z:��-lr�/�o��� H�Yh$�( `#�[Jw� �	�k W ��L�^T�" (Q��/�� r@�̗�O�#x�`Pд��8(^�����	~"�\[I����o  ���m� �I\�[50���@ȿ��%���#�2щ�0�`mg aP!�W~ �{1�� ��T��� ��¥ˠ�����`� �Z h1!;�\4ω�	tI�)�3�.%�|K@��x� q�!�=
H+P �����	u������.n�0�����9�Y ��ݤ��<����Â]��׮ �X���O���y�_@
\�:�� ���%t�	� �<���� ����Kj:*X�@�,� ��U#�/[ P݀A���� �T�a��j�
�q��5`y94�!@�I��� X�%��Hp����h������"� ,��ePt U&�EH� �\A�`�w� nh�I1�� [������$� �Q��j,: 	mB* ʴ?P(�gKr jB�r�h�p 1�(�c�!ݒ� �$d�pW �z��1",׿�x[���h��Wq;$���֟eZ�[K�� �]�=�� N��Ƚ-��Ve��`��� �-
p���8��0y��'��`�� 
�H;c� �O�Kd� �x1V# }�A.�l���� U��] �;' �L�X��� �VZ�N-��W(ؿ0�*� ���m�&�B �1�	�:XZM��j�� �0T�%:�������w�t .��`<�� uL� �[|�I_�W� Ä� Βf��'�$�3 WoK��2 ����h'�E ۓ�kg����J 3�q��W��F�s:�	ͶD��� �� ��J'M8�>7�W�q���:aT]��Ԁ5s~���B�R��tL8��0��(� ?�BwUZg{/�t�@���F%�	�rUv� |�k�w�<_ ��W &��Hb��[ ��w�� z�Xh�%*�O d�p�3/��1�h(@���: �̦��+�]S"�{!���k ���d�[$)� ��F��* EIW�0�� h�H�D� ��	��Fё�� "ݐ��Nv ��~����	�R�����_t L
8 b����x\	X^&g��D ����O`�Y80� �ߊ�^%w�����3��t����H����Xx�/ʀV�p� ;��	[��#/��` �ߨ�� R�9\*ݔ�gD��G�b��g 4	� �f�� 0�a�P �:Dv!�� _hOy����'}If �[��h�O"���B�CK�A]~W�y���n �L�sYZ5�SU ��+�3C��8ʸO!!*�;@��^k ����&v�:Xb��͡��{( :���3� n�	�F$��u[@��"�q��Q�'�<��0� �a��^A�h @P̓Ô�� W��_/���p g�y��K���>������i���!%P� �^���  ����(Q� ���0�)�L/�$�^P��+2�Rd���� ڽ�E���'�@�3�[Y����&X� րp����9��h�mդ �*��! �f`�����/��&z�  �PT�f����9� ���]'B�� �u��|{  ��8���@���D�+��S �\������ V�%�������@l]= J�����H� �S�b� �Q���(���-��@eUso}���\ ��%�'��e *#���`�H��E �c\���� ���pg�C����	@�a�|4 0%��_6 e���1	�� ���no]/ ;�����	 -X���w z�&�(ǥZM !��J��h ,to�+{� �N�� �,�i@y1� ����KZ�lEL�����0 u�3�Y�� �^?�L��� ���3K�Sqa 熽 l����rR����f� s�"���n �J�`\� ��)��<,Y�bp	0��P�H�� 2T(�� �$h�;���7 ˽mK�H��Q �Dd��[�U ܽ P��L�� �v������� ʰ;��� �ˉ3��P1�vtp �Ӂ��aRZ��*�ų��l� �w��U	��kÀu��I3 `�=���0�(� 	�)�X9���q�(R�93�h��L-�?�;��w�JѪ1����e� 	 ��;�� t>�W�S� �J$�|�*g����'���ߌy ��L��D� N�!q
�|< �S�P+�2p���(�X��� ��n�Q�3���}��@��=, �؈�!Z�6u��h;`� �|W����)�΀�L�Y@��
�����C�	� ��0�� ��p�f~[ �W��1��X� �{V�� �KU�/�z��� ^��)t��H/1�\ 0�'_ ��~T�� �{)�(U� ���ޱx �k2��p� �)����� ��B�`֥�M 
^��� ����a��p :�H[2Z�yt4?�1�*�v%������_ZV\ (*>���(J��Є��	����X `@31�� t�hR� Ӛ�A[��5 \NS�;%�} �~��� E�S���DA�)o' !W� �\��2{�y�����h�+�D� R�!�u�z	 �L`,���0��G��#s� �o�B8�� 
Ʋ&�?ُ �%����� �u�׹(�= a�鲛*w\�4|9P� �˗�.� �	��eH�R�� #�$d�X��
ǃp1�K��������b�� Ve�onY� �LX�'3��[��x���VU ��;��p��QE ��@-+Z��(���R�;�X��	�mX���  _L"��	�t4�(���@Г��� W[P�aY�� f1?Nwΰ��S 3��I��u�$�� �x�0�= 7`��w<�\� Ԁ�#?�ӀK���ܭP � �m�z
 �L�4h�p� �*��8+1@� ��>y���x V��I�H]���p�e�%���^0��i��L/�)�懺�BW@@ɟ�|Y�K�$ Ayz�lhW ��,2֨��/��@i�܎�X(܀��91�O^!e���%2�w9�/��b>{@��O���9[�
�h? !�k;R\�4���J�7Ay
;��ש�61��b�� Q���~� K�S�k���h>#,7��O����Y�,* ��i��� �
Ys�0 �\�;˾ȋ�8�>����?� U�`����� m���n��:�� ?�}0k R��.���� w��?b��# ���E�N��� n?>�1�r H"�.R� l���8%� z|H��\�o �� <!� �1��^	R �uhQ����S&TY��@�� ��A��\�� y3��@�\��	��d ��� a�2�����\=���;��x>BMz� *����m�6\�� ���<9!�$Н�u@� ǀ ��/D3��S $��K<��0�)�[ ��������,7$� �	e��U= ߜ�@
�)�[u� /@ƀ�RT��4凃���1wo���� �n ���N�#�_3��eU�0!�{W<@�K ��Q^� �쮣����S�ʔ@��8B��_G��� !�Ť��m�. T�_(Șa Q,O�3�~�s� ��N7�h�@a!^ہ���n �����RM�(��H�� ��m��� Gr!��ĩ�P�X�� 0�^*�/��9,��9 �@B��� H�(ˌ� �	'���:�D �3uX)��Q ��$�P_ ��/��r) *���]�L.�0�[�l����j�A�$pnĴ)����� ��`��� 0����(R�9�� �޵�%~�� 5�&J�m h��=�ъ :,| _��C j�bt[��� �h��1�� �5-ߔj�c�zK�	3��� ������. �0_�T&�\� ��YM��2��,��*� F��y%t����T��V���QH�O���=�� x'�����љ�:�k� �Gn�� ��ѱNð� qv#s�_Y�>R㐘�d�J� �"���z��P����2��X���+�O K��r� ]� LBFJ��� �KpjH*l �
@��1� ��ۺ��^IK
�ý�H W�9[��T �>�U�͏���Vd �[��TX��^i��ЕK� *!��+�H �n�>9y<�������Ic ϗ�$���������"� ��	��0/���G�W����s Z���T��!��/��~ �\1���fh�,JQ��e�-�� )����ݣ'`{� :0��� Z]�X��?����:�1�h�i�:�;���� ���s�l ��J���� ����[e��S��01�Т: D��wh��e�}U�� P��C
<�^ �f��Ռ��P �(���!fQ@u6'-��P� ��T� ��I%y�l⥽��u�i����!n��^&_�z �)��/� D�%
�q�xj���a#<y4R���Z��> ��G�� *O�g�.C �I-Tf2���c1_�[~)�AW��?��(�LC�J����`��N M�k� �� �҃���)ק@���������a�2� Xɹ,�B�k ^��P�쐸y>�:� �(C[Zh�`S���	���%��m�.Vl������ ��� ��gK�l� ���e����	�@Y �'�^���tJ�X�|���vOuYh#>K�����ؗ �0�}T�� �	]���!�;j����U��Z��8p�� �$�:�2� 0
ֵ���Ux���)}�2�ZRQ����0y 
�S(ݳ���4��@�
 )���3�R A���{;-ى]��'�`h� rUSP��@��^�h�N9 �!�	�m�< w� �g�� Q�h�BdZ���$@�� �t*bR�����-��^�j�2�C���!9������_p|��� �e�.���ȋ3  �f����? ��J;U�� ��_�2�8 �÷�Ltk�> =��پ��1��2e^�h����X+���m�t�gW\ <�� ʽ=X���Ȝ� �M���� !�a��(Ȥ ��%�����R������g ��8+��PT �A#`BV�RQ����}�7���k��	�N�+W �x������E%��'T�R� �.���� �fkq�	���`� @=
�U� ��v�O	�( #�?@�� W�]��N� ��������90n�
 ����� ��'A+R�x  w�_��>� 4��k�\\� ��(���� W��Z2*�㽡�D  ��( ��7]#b �,��[U�D*:��R0迶$. S�!�Z�,	P����5)�� ��XB~�#�I?t!P�UV���/XS8Q<C��"�� �V��HN�  U�Æ\��~�K��鈝�� �[��(��3H� ��!�Z��J�%�e
�R3��b��+���(�ZH[ J�� ��4Ջ£X ć����~-q�਒� ;�+K��� 	�jc�4�%���M�V����ˋ��Aq0 J���]� � �\�.$b� �-t)��� 0��	ٸm<���M}����E~� :$1����HH) %"�F ��$���ƚ|�G�����%� ������q �z1�;E ����0 	X]w�����Y�e ���1y�U� ��R$BT������������� h�뙼)�X�g$�K�
~�7 �	b1����.�����?�:K�����'�:�b9]���z�쨐s�O� �&Gl �Q(��߀ ��h�{���]���,~q� ��bEހ��v���`>��c@��26  ��l�I���17=���YXs`������ѐ'��Y(�
 �f/F�n3�	���@��\1���v���!p���/�8���q��@�,�q �5�SB��, V�*c�G N��aO�h 3�|p'�� q��$��<�(�k�7 i_^�X �S%�\�x ��4 ��~�Q�	p	W.�@o�X 3�F�2�VA9z�\� 	L�
��0�a�.(��?���I��C� 78�\-�J���뀜�I2�����1� ��
��� 𕿢�c  wժݺ��>�� u���D� �e�A�5KPq��� o�LX� 8.�O�p�� 6q*n�֟ H�C�>Ȫ� 4+�I�!;��<@ ��{� ����Y� � ϓ���i/�`w��pD�*ˀ'q� ��$��G ��u&�<� ��[1�Ɨ`���t����{��
#����w~ �����_��q`{�iX/s�v� ^��`Ո�Z��~��`�v�-=�d���)�� B8�	��x��t@!���,��(�N���%��P�1� �!�0� �R�X���i�`� � ׽���j��1bx`�� �6C�g�q,E��9���/�Q
 %�z���ZO �u�!�|P2�-��ɦ ^�g�a� �	��[�_U�$����^ �q��j*� WN����;�� 06F�i��\H&I+�G�8W�8� ��_�1w 	^h5>�t���*��?�A� M�n�w �3�>P� Ϝ�ֶ� ���*�n� �ނRm 	+�*l! @Z�[G�]�.�C�+�0�Sa �4���&% �sѵP���bmbl�\8�q��u j��T$��.ї ��b5� Z��Q�t��;��og�Y9 NЭ}��JC ���1�D� ��.�X�I&0��z�o� ��ͱ� ��`�� �&c ܯ�{a���>�
 ����h�� ��,���T��ˇ�0D�+���O!�'[aB0O���ܓ� �]�GXy�� p�/Y�� 0��|��P���J�#���:���y+�!��J �~��	� Q�U���ki�%�b��ԭ��Y���4�������УB �XbAu�Ō��\_j�WD�� J -�
΁PS$8~���[<� ��x7 P"��ݤ V%Qbh�Uw�|] @yzCER�� )&:�!���L�K ݂�}�� (�P��v� a0�,�� �G���;�;
� �`�u �+��_b �r����  ��tj��: �U�G��[ ȕvk�\_���#@�S���u| ��˅�;��� (.�
��� ��W	� ��r� ���IU�*VK�����n,��2�wL:��� �j�� ֓]\�/ ���`�(� KY1�������@�{�� ������ P���?��3( XrN��8�^ 2��[RLf� S��� b;������}Z�z��58�>J�����i�;���2@��y�| �J!���L}�����@�( �[0%� ޙ '�sh��� aŅ(j�<x��i �L, �[-.w$�
 np*����1	Äbm@��ݔ �6���� (����!?�w� S+���Ml� -$�W1�) n������ S`67H�� o��.�IG�.�Wh h����	 �S���'tz���� ����!c �:�Ѻb� "��ҹ�� �P��Qѷ�a ��2ø'g@���Ь~N�W����+��� U_ j]�? bEYd�@3[ 1W�2ܸv%���*���]P��`J�V~� �z[���� �������,{� -����� @2�Y �z(��� �Ku��ppU B��!������������7��&��[�@{S(�mM�� NEP1������aY/�w�e��� �*� �� Y��G�U��9/� ����M�����e �n�[ �)ѕ�`�{� a�(AQ�:D�ބ
��� .U> �,'� 	}�9�JҀ�� ���[� ��F�� �	�YH:�<�� s��D]vX �{hg��7��n�� ػǘ�W ��P��t����\��@��R���?�m���-`c ^	��}8�f�D �V��u�i>^�H� �M"A�\ b���H[ �|u�(	� OR�0�͐�%aE����r����Bh�	>�̀k�L��^������� ��I(�� �tP�@�_��X�K��� �t��� V	Ej_N-�v���� #�Z ���0ق �9�UT�o�HR�?n�u� ��)���$Z�G �� a�q�~��~��f!��@�si  Uہ���� �x;B}�A� ^*��" 7y��� 5����z�����J
��+�b��\Y�� 9�B+"� U������� h8�q�� 	W�ʹ�� �2S-B�� �]$3�Ri�x����
�����h�r ��a��W�3.�#�S�8���� ��5�0,X h%R���> �|�π ���J��;��@*� �tQ+�����}|��(�~Z �K����p. �_�v%�Z >NOw�[������@��h*L�л�b�� ��V ̾i���% t��Z�*>߀�ۭ;[��B�������� �"/�\vo 5Bz�0t�pg �e�IH� w�/���� J_+�$�	�x�1��F�0�j!�6�U"i�� ���ȝQ�a �X|9����Z��03@Ũ��� \2�!aXd9^�������~"�-D�&7� ���_�fprW�G*������%��i���a<��}j �����&�� ���h3{\�6�uH��g�o�@R���%	���D�H1���,��� �pZɿe ��vh8Du[�Vf��
��@��_!ð ,�W�(Z2���R`~@!�u���k{�wۘ�=N�qV��Е������p |bL� ��RP�x�( %��w"�L{ 	R *���h�G��LsX�o T[�Q�b.SW��@�'�!��C
m��5� ���}�� $��	�U&+[�	�� P�w�*���@ģ�� YB�#�� �R�1Sk��~J el��ϡ 4�-��� ��J��R3�;x������ N-�8�X����� *Z�h �#�-���' �+^�2�?���� ��0
���� ;�G"S� �Ļ��XK +������Q� �p�5�;�Ȼ&��T�(<��	�`�݀7!�*
q�, �����wA ��z���ø D(�P�� cZ���������O��D `�Q���0 ���z��� �P�qb/x} �0�f3* ��R_�8�6N��� �*[" �Z�KV����/W]�o�H���t *�
�[���}x 	R��u0$ш�X;N��[� k\O�"�=D�	8D��2�]ܾ��	T �g_ �b��F/�A ��xL
Ⱥ ���	�D��|�dØ�L� �V��Y���>#����5. ��8B��^��O6`�@5�. ��s�L��\�� 3)0�Y!�d ���(�b?�W���Y%
/���D^�����R�lwx���;���,S�� T�oG�D�!� m|� ��ğO_��o�����V��Xg��G4 �=���Z� ��0;nG ���@� -�9��"�.�r� C3��%� 1p�ׂ��9�	� �iH҅�@���� Ma��]�( ��\u�	�c??�D1�&�� x����# ��	<S�|� bZU�m[����N�������<�DS��h5�� Q��!� ����(���nKۀ�� �E<pB 0���DI�:j���	9���W`�hΔ�-s>�� =X�[)�� R	��Hn�C�,=e�pI���z+��z��[��C� �S�T�Q f!�˲� ���h�� '��5��� �1�&ow_��+�@�颒�~	r��A�|�� FW Pз� ����a�u� ��+W�tP �-�R���H�5�`�� ��~l΃#� ��.2B��XU�(\׽ ��N����䤅`~�J].�� p���9o�� t@�ڒ ��>�e�!�� �O@�Q�s� �<�����Ȏ�3]����V�O����x"�X�� �T�nh%1����\���&- |⾁M0�P�ڸ������ V"�Ŕ�{� 16�����=� )Z[9���ɉ �('~� ��}�2�H [�iP �*� @�C���� 3�t���&�["��#ɸJA��xI�ai1س�}��Ͱ������7�s '�:K� ��[���g ���%6�up' ]$��� 	���M���`�AU h��������F9����41~��Z%��� 2'V�@ �[��ah~-i�y��!���`.�����ޠ27p��+�KY�� C�!ʽu�hQ����ǀ�6��W�F���ATv��_2�_ۨ�
���� Wt�/"� \��F�J ���P�s�t �Mف�_ �뼨� ߈ �]y�L��A �ܿ�K�c ��(0�n� ��
.�=��FgA�T �#� ��/�_��0�t �L�kp){� +�A���\ '
����%�� �B������ '����/�� S�s8�N��U.�Z�)쥲]��N[�@����y 2�h�	WG��@ t�A�~+�1"��/�S�z�����!� &"��<-_?0� Kͬ����VHIB�L�-��]��C ���%�h �'k�BÈ ���0j�$� ��+p/�b{�5�]�@ d	?��G��h�o}��̆���+�Z^��W�|c�� �"�Y	����!�]9����� � ������"��w��O��������� �J:��(�* I�Sv83�c ��1Jř��0�h@�4y'2�z, �3�Q��L_w 2}�c�-EC �㺮i��$�)� ʢ[S#��ܵ ��1h��<���-\)�4�N��$������/ �L��%l���8R��\ 1	����� A
ֹ�� �3��?: �آ4���� B|���w ��ݞ��n �}8�[vY�K���F�@%>�`2�D#��5� ���HB�	P(�w�^�̲4 �/���k�v ��Z��� ̲&(ɿ�<�`���c*-@��. � ��>I�_1���Ё!�@���F/��Av[~ ��a� %с�-��{zCl�Y�
S��\Op.��! `k�K�� N����L� ��Z �Jp�����2���^(���Qs�U�� ���n��[1 ��Ə)�� ��O�&�@j�zP�" �h���� ��[X��\r �W]��� Hxd|28Ծn����^!t{ �J`�X���(~�A��). �G�d��O �|/�-zq�	�@�G�����Sa�	�ט���I�^ U��:D*� �AIx�� 	ۉ���<<+w ĵ~3�τ0X7V*v% m���ε�:  ^������ZP n&�� �����($�~%�� NO53�)z��/~�N� gҴ�	�h�s q���tH �0.�XF���r�� �^��ܑ�<.	���8��p��J����y�����. R��]h Z
`�� ʷ4��� ���J����/hE]�M?^&� ��Z��{���f���=Kځ!(��I��L�� ݏ����u�� _��؈rC����4,»�'�	� ��SB�_3 ����Wg� �U{@=0�	G	�� ݷ]HYZ� 9�U�
=1� Ř�y+ �V ��@�� 4�J���=	?�� fE���^�I�B;�'-�ǎ(H�jfh�s��d���6�ߚ `B�1 E/���hZ�s@5��J	3�QR�^��� �2߉}�6	 ���q�����&Z �� @A�']^�� �$���MV�X�_ �@'SI OL���_J��h�V��/W �&��Dq�À�	��;�#C��( @#�0�x+ �p�4M2� ��C�SP�h �d���Ź �F'X!@�0��S��_�� ��-�V "W�#!�Y kR'�]i��`�
�#��=W��\S��/�� px��	�s�<;��?� ��"R=\��;�Y
��� �+R �X#�P0�J
j/�_>���i�H ����?]LÄ����#����0� �����, ��yڗ�'�]0��H���ܔ	�
PKC�,�� ;��&+ W�tq��B ����]�	 z�}q�i� N#2�M1^� {�@��ub �a���� �Ĉ��t�	}籓yX魈����S1��o�Y� �vu$�B��w��0�v5X�f�r���^!� Z� �W�0�ͼ� fw'� ^�:h�e�o �ƒ>ND/ ���h�0 ����r�  �^��	�+�� �5��z���͡b0��;���w�� \�h.�׹ Dr� 4�U@�  �mx�_�� 
�	�v���XK�.�� <��w�;W؀[��c<��-(�t��.���� 
m}8*W��/ V���x�� JU�����r� [<(.!^�� l�Z�*]J �ha�'�y R�<Fze| 2�Ժ����y&(�	z� �aW%^\&@y5�� ߎ�4�J��� /�X�g ��̭�i	�\������L ��g�� ��B�
� �'HpD�� �F��P�� 
��	.� ��E��t1 ��	<Ĩ� K�2�#W dP~
� i�_n�w ��8-�֜`W鴪����0R�Ʉ��� ������ 7A麈9� Py��C�+$�1B� �۸-� ��@R*� U��P>ЇW �0����1�L����I��F+�P�V^� ��D���	�X} �i��� ���yf�� a��	��Mմ�� �W\RI
�(�����c�W��� ���g1����bu����B�]�9��	��+ 꿆�x���_^[ �Y�� c��O�*� b9m�g�":^W ��,�!u.9��:��@V�9�� /�L�4 ����S	� �ٯ�ѼA=�� .4",��l>� �
h>9�� ��5�`�� J�2�`�v pB��Cs���� �#��O0� v��V��p� �2XY.ht;&�����4W�n ���
�� ����?��[b�0 �^��ZF�\��J@̠�H֕^i|$� S�'x�d0aO	�j˾�� ���� �&!�B�Ar%�������p}x �3�0��e����4)�݉ �づ�Z����Գ� Y"��X	�*��^o����� �P4�8�0� 	��&GR� �[UWtZ� �{�!'�|$(��C�M�����#� +�y��� �R���~l
ڸL�PdN���_�) �S���� ��Ap�Y͜H��#v�/� 0��ߪ�_�;��fN! �YR��:� �#�k�¨XT]�!�S �Qu�?r����)�1 �W*�T�s���3 �?)�ո_g �Wi~�|P؍֠+� �;v%5O���r!��ă� t(a���-h������ @щ�8` �VZ��=� Ah^�������W��+�L�;��] �)'0�� ������X�9��޾� ��P��m\�@��h����'�ap�ȸf��c�u` J��XVN[�ȓMUD@��� ����� �,��\ h��'��� �H�V�� �� .(�� ?�N���� ��1���z
�� $k�A�	��� ��S)�R[ (J֤3 �|h 1S�b�:�q W���{�� �L�s_[ ��
e<� k����!� ��z\������% �|+���� ~��h��wwY `1���;�w! ]���ib���U 	���#Q1��!h��/�e� H�M'<6�� vOx��_� ���Af���S�aT��K� �-� | q͡���J >L�4�%�;!�
��H�ޮ ���n �?.!ےI�� `�0�z ݁��/@�.� d_u1~�	���!�[0ŀ �h�:o&��� �
B�G� ��l��t+�Q K�,_P�Z �m߅aRo �{�� QG��E`ݝ�,��t�9S3ҳ���'@Q�� :��7�� �
�y������`��!�C$12� j��qZ� P��aɽ3Ww�TU �l	��:�ؤ��eg,�@�c Z��%�� �y�8ܒ� &e�[�I�  �w���ç ��'�v�<�{ 2�]�� ��������kI��D��1�'! �PV��c�a\��O� �����2�R A��L?���jQ��a����~��4������/!��A1\ (�� �B_�6�
3�����@^a�U�� �2b��Y&�P) N����. ����l;��O ��� Wa:���e& (���!�P �\/�ɉWZ���� '���L�~�_I�ur Bc�5��� S�TY��� D��ش	Z� ���5  ������ l�;i�X�� p��SA��� ��:RW��)���� ��l8� �_�O�aB� K�e�N)�7���{w�1� �Zi��Z�� h���_8�  ��C=q�\"�b ��]i�l��9����\���?`��,ޱ:�& )�\�][���@��f��������V	R�s^P�J� "\�Bg�@� ��v��P5wv\xB k!�'��"�_z�X(Q�o�� �S�+ u� m�B �
�[Y ���)t���� ���W�*�m�n�`�x)+�o��㯘5�� CN�"*�{ ���ˇ� Z/�g��3��<؀e[�x�� 7�c(H�$-�@@k�{&���R�< ��ߐ� ZS(�ܲ�� R��6�� �h^W�%L� �4������5��j���h��b�����@C��]ʨ�} `�8E:* u!Y�� , 
a�p�j't� ���[�l @�%�/Q� G�tU�D�� (ً՚N  �Z��H�?F, ��c��� �z���]Q�=���5�~�x/� K��L�jP4�AD�{2�!K�ȡ F:ڧ�_���-E ݤ
(�� 2p�^��bY��Ƚ�PՅ�	 v��I�� �J�(�\�ah�&��0�R� �U���� ~��.��8� ������ 3�۠�R"J�({n ��&��}� �!��1	�(9�_ ��`Xh:�1�  A�R	� ѽC_$�����QXִ�p�:H8^��)���X 2����� 4�h8�BK� ��H�3='�p�<���� �"��=�l��|>9�OG�d0�� �L��R�7 �@��'J�!.��� g�r\�� D�K����0�<ڃ�_F��
ZꜲ� �.�G0�y�PeS	��*�W 9G�>l2� �H!X�� �:]����;C  ���9Ŷ տ��1���$z3����� S���ʸr ��(�  ����:WiL�Pn' ����*! �����ﬖ��֯`�"�	�eB�]�@��Č|^ �[1�v�%�C���L�� ������c|l	 �ouj�X �6^馔�0�E�b	�?�0 @�e 6���Z_��xH� .��2� K�A��R� ��������y�����; &d��� \"�[�
^1d�8 Z*�R���
 �$�/x�|>a�n����� -����(��'1�m�~` �-5b�� ����ΔR� Z��^�|� �Y*��ޘ� ���,�R��e�
��X� ��(�^�A�� �/�������ip���:�AL`�,�=�0�׌�py�{+��1��2�[�J
�S����0ڠn���?����@��U Q��1��e ��Љ�C�>�Y�I%a���� ��ū�]Tu$ �	l�
\�n��@���1 ���D�W�o������,"�I�[��7��f]���Ȉ֬v���!�(���/� ;}�N��F� \���H�o ��-��P��z� ����X# � HL+	���F ����/3�P%� eh.�W� �E����*8v� 3ǳ"� �	:��/z=�Q��࠺���B��\���G~�(F��HĴ �����z� U��y�D� �(5!�\h s �3��/ �|�qÄ 1h��=��R �0��B`[ D�p�b�< a�'8]hq^|!�ɶfu�`�i Z�]��I|� �Ũ�h�E &�}N�FL<	������;,]S FT�h�H{� |`�<�@�su K���!8cP�� N�Z���6��� �	!��r} w��$�Ý�	�)��g6���&�HM � Ј��9�� *%x���D �n螹.�5���$�� ���a�
� Z5v:�\PQö}p'���3����" }���R�- 	�*
�Lk�y~��J�pGj �����0 �^���XN8 ��t:�ɰ��޶�p��W ��3X/1�<\�� ������_u	��q({Ք�] ��� ����
p0R�^Z�� �ŰOh J ����͸�=2/
!uP� o"}j ��)���]q��0K�1}�?����[T r�M��� D;ʄ��e>�	�Z"�2�� ���A�hx
�IH"� %�8���&n0 @�!L�� ����r� d͘Nn�v� ��}����. ��ނ�� w\�bL- d��!�(���n�v��G��@�
��^�#�' ObQ�_B��ʰ!���t|�^� ��T{�(W�:+�k'��o~�����	9�P���敀��`�9�y�DV�E� :�8���! �aB
>� ʌ6�^ƅ Y��-� �?o]�)��uE����s�ɸ�%� � �ȸ�p� o�y���m ���M_ �`�x0�I�k����-X���H[���u�(fh�=�ـ����O ��Ss�K0 ��ʗ%�B+�&������ Wpu(I� Q�$ �bJ) ��Pʮ�' �p��꿥 ���	*�8���5Tz��� �0�.X�4��q� �/ �r j���W �9��NY =�i��q��hP0햑$� T�`��� 4	y�~E�{L��rQu ���d��e8����_�8��p��s��~�F�� ��ݢ�,>�� �!� �Ƕ����'�. �H4��) �ל0�� 1"u͞���p��vXPLLQ:ι[��n�P�Y�� R��!��hW�`��_ C�ۜ�?� ���� ˸���/�x�� ������ W!S^��*�r� ,�R� �KY ���_�����s����!��m �)���?% �޸p����M� �{	(�ݖ �"�h�HG;��
�2�����m~F�pX Y��
��>� �� ��,� �Q��F΄?� OҾ��T�B���b" �x	��� X1��8�h� a"�#?sEf	Ћ� ��l��^��JR?��� �_� �b|���W �0���w ������ :�p��t��
P��{��N� ��[��d1q��䘷���P/[.-=XL�H��% �lz[i��Z��� KL	8f8� ������ � �O�i� l�蹋Su�&gZ Q��	 ��\��_����!� ��*^� �"����]Zh�e�P9�a! ���R�,�{� q4h+Mf�^�[k��������G
�	uy�n��W{� � ���[ ְ	��EnP�@��0te=� Х����0�%	�Cp��#� Q6��T�
 �x�$�� �A�4���K��:��Bж���Y�����~��J���10hx�r�����(�� ÕvӉ�l� �Q�1��,�L �5���> ��H��|P��){�\�N ��	3�m ��֡'w� �-�1A{Z�(�h� ��Q�����2�����&�5�G��W�i0.#��(^��ɵ��2�ǿ��!� �l<���/�3� (����d )Ĳ�My&xa�p�� ���%w�� �l@0����� y�,�%� �K��3� ���kA hP>U�׽��y 'cR�%�r ̂Z{�(�� K��!"�7/ �DXt�������\C}@����P'p������m �<�}8 ��+`P� ����_|�9R� 
�w��N��&� �.�]:� <���� =�v�A�r jӀ��[� J%��?�� ^}�f)�z.�C �!V�� 46	빍� �]�b�� 錇�� �y |R�7	'_ ��%u�;�� �FL�41L������	�sa���_M���o �gs�J, ����:@w� �bǐ��"�� '0���� ��^��\h-kDTP��Cܘ��l��R� pf�"�L�J  �&%�i�� 	.�N@�vl��O�V3p�a 1�u���� +�Ѷ�=� �ˮ ��H�c���'S���;��[��ZP	� ��k�\^�~ ,�W&M����i>@1�� ��	�����k�\����|�����C��\� �0O �G��;B� K���,@ �ŋ�0� ȉ_��� �P��|����`@d��,'}, �3�E!� ;\�hd, N�ߜ��-�	���#��SߖHl3 �5���~+���(�`��q��i�񴃂��[R �D*���� ��%��|� N?���� �`i}
U�b ��h{^� �_qM��� @i�h6��&+�Ä�.��� 3�Q2��y^uO��=��Z�� (�VT��C�2 0u&�\>6K?
�������D��(�`���@��%!�DV�z����u?�Y �����3� ̹�-��L l)�#�Hn8h'�s1�� 8 4��2�\hQ�U� ��V� �@1� ��+� �t#-�P� ��_�Fh,�e3k@I��;�-l/�d� *� �<2�!o���Ł-+@������d���`дPU���r+BC���
 /��-��(��33��`���%n�XI�>w�� :��,͝?�������$0�^�x���[��* �\-�htS $�)� � �_�em�r�	|�[ۘ��\��ܻ.�@�- ��"s/~��#�P S��wL��Ѐ <(�*i�s���h�UFK�+� W��jޔ`���_�,i��ǘ�)� �.�9: �D��A�&�;��R �9x���ڏ��`I��* �0�Z�h �[~��w �y������ ����L0/�8'�b�e����ր/�- Y^���-<�`Q�Z�����'�,��A �?/�j� �>�װ|�>N� �O	�{]J�����.��Zi��Ub.� ��	��Sp �_Ɂw깒��G�ؖ0�� '�q��? 	o�]pEJ�!Q�� ��`�0���E� 0�	� ��%<v�� ��
����I�1��0O�|m �Zq�}��L���ȿ�2:��p'`���PT��X�8��O&	mÉ',��<9�?�+��S�Q1��k�� �n?���j �W��`� �^Ҽ�[	] �~�b��,�{L�3�fn.�(�#� Z�mWR�cS �ￊd��&���< ��!^�q�����q� ]���wz� ��S@7�D ��R��E,g� ��r���P�����9 �� ][X�Ȟv'�
d`��z� �,0�cZ�� � ���C-�hP;�Gc�-�Po �f��lջ�����;�$8�� ����s 5R���� �B	a�@�#�$�*-� Z[
u�b ��@���w���0���^� �4���+ �A]�d~'���X� ���j�P�8 s�NK% z�J��~�� o�)���'<!ځ��/��K|P� 2��r �1�t��? e�	����wΟ9PUM���X ����� �o�B� ����=0� п���h���p�W��n�y��Z@���N��R�p|�� .Q'	�%2t5��i^��Z x"���-� Q(P�2N	;I������!� ��ӭ��fʪ����V ����yi�r uG�b��}F�j ����S 9��@V�>�� ��1> �� `���hLD��(����漯Z �Ip��{� /��!'���&��D+��P� �(����!Ь^���8� L�f)�%?
ڸ΀b#*٣ս ��!Ř�w� "0�Z_� ͺ����X����]�DȳZ� �8��JE�, .e�{Q�+ �
����|��E� ���</Z�����E�.�qق���W��'���G���Y�@�� Tk��/t � #!�Q	�D���;���3��5z� �X�ؓ��M h8YZ�r�\P�p�("f��=%�a�n��� [`Õ��uO�	v�^�|鉼@���DLTa���h0|4�I N_`���%� 6R�jׄ" �a� �T?/���� �H�x_�y���.`^C�� �󘃔�9b~�P��cj�� ��Z �� �jn�D/Y�5��
���3�H�yK� I�ƀ�R(� S��$�K� t��\�40-�� �� �C�t$R" ۺ��p�}�8�Z �!�0�HY �������� ~���r��v�������2�`h��я� ��Ze	�Q! �O0ν
S �?�*�	�� �\�%G�l�< z��f{� T\�a�� �Q
���9 �>�[Z��� ���3K� ,��(����Ї� �Yދ�b ��|��>�x �\�����b W�B&� ��H<�R�2�X��@� Φ�>�)��	�'�� f��. �b��A :�\�ȃ�s_S��E��3��� 0�@-��hA����X�0' ���|Mi)ruN ��J���_* �d����� ��̂�. �ݫ��9�
�� ��?��\Ib���f�`���7	�|x1��'p]��=���}N�&R�݀�F;� ��0/m6��PR���)�f9��i ��z-p�� d�&��P ~]���C� HxW.��b(��� �UZ+�]�����jO� ��k�f �G�Eb|� <��`��h l�m�� A����8z饄tN$3 ���\Eh �
� ]�� �*�̻i� ��!�x4l��u
��� �i#�� e�4]�{�  ��[��u��*�g2��~͈��ـ���-� ��vZ��{��"��஺�� X'�|�R� ht9�5���XW��r �b��0� ����:�d� ��e�# �V���D��]�i�@a�*�[����Q �yo��u��+���#�Y�S��Il��^�&T�� }VA� �=mj	�_t TY ޱ��19�. �z�ĩ��p� W���� 1�_ �¹ Tֱ>�`3� 0�[�!� �i�F�l�� �n��h*>+ �J��P�� ���O�=�Kd ��f���zH �,-��[(Շ����XZ� �:�l�zq� "��>?.BX- ��$��	�z�P���,�'[Gb��@���:} �^x�>�㐅��hs58A�@������ 0�ncؼ�V 	���9H �@Y0'�X���=G� �.���y>
��]ZN�������� �(X62�>���PS��/� Z[�"
�� ݙ�k9�� %��'�3�� ��냾�) ;+�,�̨� L��9� �{@��	�v��Y�7���0�#�\ ���ހ� u�oY�Q-�����	����p�1=��?�7�e�����k�겕��g�m�Hv���	��� Q9�� �h\1 �q��K�� �`��(0ղu�R�c}��2 ��5Z8&w2 J��Q�V��  	u��y� �^�/�z�Y|��Ex����iB`�'�;C��Oq4r�i~��n���nޟ��xְ�7���	>_h�P�)�����2 ��I�z��U �����P�� fY>�|r� W�Ϋ ����/�\�[ ���q�v� ���S��Q u)�o��,y0�飐O`�_��`6����,������Kً k� h:2LD� �
��� ��U��JT� �=6� �,	���wP[���-N���&;�l���3Fe�<�,�hpbI�=�r2�� ́��d� Z�b��`� M�]pOΨ��"��
� ��.U-b_� K݁Vú o#�"	��u
���{0:�S� �0�~����
������_�� �?*px�� ��s�kĚ N��j�O��7�Zn�����D	P��HU鼀���K �hk��;��.D ����V0�?	������AL�F �.��:��/�ϨZ�[��=x��� �q`��@ S+'�QD��q0 ��`n�V
� �^�Af)�z СH`:� �9��h���Yp��X)��V�������(�0�@����f?&�����o�lvXh��-@��ܪ���#�m wd���/bM �o��
XZ �� �f�/ �5PF�%*� �&6`���W1{�Qݻ� �����?J&0����_X����@���� ^�b�w����]�����7 �]z�K+� ��	J�e��[� �T3�% )��R"}{Y ��4^$��wZ�1`� ����ֲ(`�퐬̞�P��b�<!�`pѷ� ����������)�|Z*8^� ��t�� U�RI�Z �Y#�� �$��D"�
���_U 3�	P�0V�� �A��JZ��\Hr �� 2��}?~I l��J�� �����Eɮ�p� ;�*vD�' hХ��� ��Յ�!����T͟��W�h �Dd-O��W �:$�@�� !�2
�. 9ٵV�X}jJ� W#� N|�1E�7{�wj8��&Z)�9 \;�^'�� ���*�R� Q��1uE�AY��PO���� �@�V'3�� �aED*T� ������ �P�A��S ��섖��� %�f�2��Z��ga�.�>^ ��f(�Ұ �%QKF���	��h�B���ρ����
اx� �23j `�f
& 01���]�$�ˊ��� Z���� ��h��M` wΉ�Y�B� ��݅�D���)��~����@Z� �̖� �.
����9U9�`��R��X }�K�e��� �	��\O�� �o+�3��. � ;N�\ $�CU�Q�"	�Ipv-�f�(Y�������B�� `a�W� �썃!� 2��	�hS JȪ�N��  G�dLŜh "�I������{ �*��^��NW��>���� h�^9Q�g}�\���  �`~��;$��� ��V[^ ����r� ����a�9�?�6U%d ��ɫ��t#�� D-�^h���_�%p�5☔ ��S�g� �X[�=I` p�RZ�T9� �D�6��S �\�&� H��8 ��9 %�A��p� ��D����f��Z��!���UŲ�ɮ؆P ��)	|$_]rV2���wc	 7ğ�A�HM� �i<�x�k ��p�( u�N�� ��_��-? ���NA;-��g h!+0� _��3��)ׯ�],�Ue���\ S�k�кV	T^�|��F�bR@:+�ܚ ;����VPM�_�˽!���p �W��[_Hq� �/�`"5d�) ŐJ��
�܃Y��� ��'K1b��� +������u ��D��O�g �\�	�U�[J�o5@��{@L�� �k��
d����7 "��<P�@��8M��,3B�-L��Jj��	�Q��E�h��\K��aS2���% �b.�:���
9	^"� �̒��� ����9<Y�+�i�� *�[�}D� �a��ǂR�,����� o��Xx1�
z5˽ .���d7`��g5 ZQG��;�L�� P���3[��ܳ`~	�h	cQ��?���@��
�q ���ò4_\ cAXQR�� b���W| wD�4 ̄� ����O�tz"���$�� S%V��2�u v����,'� ���Y|�Z� N�(���Xc.�P�� (�0�
Y$P � 'H�c��"��� b�*� ZfⰀT�} 2�l��Q�LAt ]8b'@�%^B���5� "��XKH�_1�7H �}	���p�� \3�W�i8��Hm�Έ뻦 ���R�XD� �rYһ!/�i|S 8;�]�$f�T�{�XS��|z �뙔���1� ����WF�9E�0��6\�� v<	��� T����<
8���f��O�6 ]KW�-�� Iݐ��4X��`��e���� �>��g˾�vƿ��^2�����EN�����<+ �
��M݄� 5	�4@=SQ00[0x��=k� /��&n	�����3
���� �K�� \*j�|����.^o�`�VU �pq�0�}�<X�H��ؐ5� �K��a�Zq ���� ��@ �h�v=�; "�-�`Y� 0��!Z� �h��	��H3s�� Y1�� �m�HU2�Z�݅X��@��<d� 0�.n��_�T����� ��0��he� ��,��9/�L'� �鏆� �w�.�tr�U��Ԩ�W� yG	O����Q��@c�N��� fâ �@����ڵ y��0mr�� .��f	 
΂�C�  -�24�	�!�n��[� ]����w�,��y (�h�R��E� �o��A�(�Z@]J���ި �qc
W^y|y� au��J��X �GL��	�}��I72���! De�[C� �_�(wȘ �O���KX YfS0��V ���#�2� j�}
^�� ���5�QB�@�\��%� u��]�U� bOQ#+�T L���\��x �q�2��+� e��Ex 
��[U� T]�f�J� �	+�|E�y���h���W�^T�%
 kS��.�z�o����|� N�5����)$Ug| qƪ2�f �@Ģ/RUvy; �_ME>? DG���Cv
�	we� (�`���u�E�u��`ս9LՀ��	��P �`�J�'W;��G�I�Uy� `>��m�2 ow��a��0�X�����/ ���Vn �؂"+�@< �e��ú�$�2� 1�ɨ�u��X��=���D
H	C�3�]e�R!���Qi���
�( ����Z'���5�����D�� �o��$��k�^΢q@�>" ���Ht���y���NV\W �[�Y�(� �lR@�?6J 	�:j/o g#�U��n �h8d- Z�~�1ʻ &��t���K��y��0���]��:҆@IQ"�� ���`�z� @y+x�&�) ژG������t ��R'7ט{ Hr�h��/ =�"6��.xY ����^ ���1��� �|_&�~ ,W�s��� dS��r�HQH a�F7Tv� 5���D�?������ͩ��R ���DX ��-��� ^�wl�<�,r�P 1��&�
�;��� �׺�-:�C �b�$.4� ��}#J��/ �y���O�C 7[j\'J �F�����>c@�I6�k� v��8#�� ��0�C�  r��N�b`Y>� ������ �0���-!��c+퀮�� ��n0jFk� �Q݂��l� �p�h]U� ޢ ��8c� �Ox��qL/ �HN�b�B��y�u�(�k+ ��]�cLQ� 50�h��� ZaN3��1@���X'Zŵ���P� �H��	�:傀�hR4�A ��/��v���d�Da+���) ��^k�Y��(���>z�m�� lsÀ�e ��"�	�߃^|���E�y a;����p��V�R]v@b���  �:�p�� !��_�) �/�\�`�
o�^�ؘ�����`� /��|�8iu7���,@�\ �w��Ӄ�S���%�	�.�nt �Io�f����3���Ȅ:�� ��@M�r ����&�<؉@�i��_V�E�0����%�[ Ba}~@rtO �H3� ��
�Q�!���|�������E* �1�[!������Kj?Հ�%�POF� ������1 �D��]�ɭ=l� g���?� �Yi��� )	�0�?_- ӛ(��� �ŭ�V3O ��]1�F� !Ҡ����W붌0���X  �Z�UT� ���^a�/� :���Q�']n��a ��b`���%� �2��� �芤��� Sv�a� �0 �LR�Z����?F�7s6��a� �b�R ��`P�
 ^�-�_4�w @�!�¬�� ��h�};#WѺ ��,�g ��P�����{��$��g��P/�� 
���E�� �^݌ ǉt 
O�鯄R� �������2 ��BX��8�)�L��c�� ���R���%���G_�"`|��i�� �z�{�&!T� �+�s �Q��� P/�u�� ���S�`�tN p!� O�� ���7	Y~�u�0�e @R0)���=� ����_�&�N���10Pڱx��>2`Ҿ�)�7��p�Ѩ�} ��fP\۱0ȕ���Āh���(����� <S�4�� �[��f +�X�ٽ�"᫅��ϠdZe[�Ũ�t�a3� 6_�Xk��7��\5S �b�v �n��x, Z ^����0� �d&B� �+�;z�������R�q� �S�+�L�r� �K١1h ��;X.&IU�� A�@��' �	����.En]\��h+ ^id�����xI��@�ځ�0���(����	lR��g�M��L'�X���
ŗ��6`�1�#�Z��5�������	��X! 
�?�h�Ee���p( �n�F\th�� A�-T�� �#�&Ç�h �r�P���� Nμ�`
�h ��P��E����%\3���4-�	~� �29?�y���� � Q/,��>*=������b� nǞ@�0 �f^��Z��h$��i�yٸ� ��@�)� �^Y&y�9��<� b|��1�V��� g��	� PZ��^ �&������P� ��'�A��|��J,☘�Yy��<�3�mBA`�T��}�=	�h.i��Y��q�?��Pk��l80L0֏�ؐ@��  ����X�[ȓA����h�{� *ՠ���Ǻ0�b���k�r �\� Zɜ��Pp� �{�#� ,��z�  �T�:�2��P}���ϐ�+Ż �g��%z<����[W���Cp� �h���� 'a{<�X �2��>��� ��3��
�{^.)�C����	0�W�"O��cr�ꕒ �|)Y�����(��.IkL� o2��h� �!�unK= @�L���]3�S�D��vR� V
}�p� @jQS'��y �/���8� <-xs@�0X���(p�}p�7� �S����) �}�îﾫ �R sO��U�_ɛ��{ �C��	��� <}8��@q h-�S� L��_� 8�� �X���*��}?�� �2� �ۑ<Rf�൚�M�V�	����� �ݖ���YO ��E*̴�([���L ���{ J�BkR�� U�g�	F�z8���>% �&=)�����@�� ?Q��03����LA�����%N EޮX��z�>��!�a`�Ӊ� ��Kp���!�&�+ <|�-:� 0O7�� 	r1K3�,��; 9߸�� ��u�i-�t� �ް)%3�� �� ƨ� �����
2 r��_�xb 	ɲ�BX&�HQL�k����� L����>I ޏRw��� p
��&> ����o]"�	XԜ��?R�qC��>��@�: 3
+��*� J�C�V!� �-���G�&,ɴB� ��rY�/8�آ�-�b3����E"�ā��k�	��(�w���� g� �Y�E�� [�Ŝ��� �\D"�
�@S�� ���PN.�&�D�D��^8 0#�m�5���� N������ %��ϲ�X ��T?��J 17��<_[���!�� '�X�eg��v�$�A��ژ[� Z�U� u4X*CP�� �����$���,�2ȕ[j ��U�1�mH�?�7u��2`n�v �0H��c� �s(�Nf ��ݰ?�H�Ջ��3� ����`m-.U� �����I~�B������� ݬ���h�a #	������J�������մ!�X��߀pQ�� *���{��~��݀����f�2����dۀ�1��� *(��� ��J���$~�m �h�)�*�o ��̿�H ���]�SQ��vs  )_�� 0�c��� V��]4�[�N�:�*��� ��Xf�
h�r�a�N�~�!�C ��4�z���� ^���)ع ��XB���w���I��:� �t�L�
P	���� ��Z 1��OJY� 5��_k�t� �S[��4 �|���:���T�;���L8wZe2���j�� ��>E ,��*�����pJU�� ����\�O ��a�R�+7�P �d'�� �\�^�@7�	�e� j�:%��t� ����_�Lr�H� �p��� R����	S"M�� ��М� '��GwS��ń�U���z���s�}��o^ D.���_�I��P :�V�� 9����� _$����� G!ф~� %]`x��X�߮D �����2(���=�?�7�#�C Y��h��F ڐ�+�X`���� �@�����9ȇ�F�p�� �C�Y�����j���=k���ca��=~Y #�@�&��> ��H03�15<�	_�/�v ��[ȁ�W ��:�!=���K]��\�� n�O�� M8U|D�Q&o��_�P
0<��1��%���9� �z������ R�Q�k�3� �x�{KE� _�1H	��b �e��w(�V -ݾ٧������?s� ���Hk-���� ��N�p�Y�� X��q�`� ; �
�񢽐�lcԀ�3�v,��P ���^'��1 [����0�/P� ��}�� N���;�'<| �+��~����v��z?�6:! �J��0�Q��Y� � �R��r ���}�� ��ً	�`t��
 �_X��P+qb �R�@H�Q�?$Z��(�X
��+t �^V	�y� A��b4O�.x%��W?z��Y�� ��K!	<�\��+�ǵ��p� ������3>� &�l�� ����f	� YIxC�' `\���.��	)�`�v�Z�����H_"吚�	� ��K�
��P��� Ȱ�Įi�J� � ������e�t�@NX�O�8�+4�����`�3-ħ y��zX�I e/�1��� �B��w�.� �ZM��%� NnDlY�	]����L� ʨ.,:- `'���� Z��+��R M����e��@0-�}��P� ��o����
�����( 4�L�')�ZXΒ�*}�ᤃH#�� ���VK F	cO� ���R�ؠ 4�Z�� B�3�kxN��EUY��tʘ�������@ �%9u���{x� �H�g5M +�,fA�?�~����WC�Q��k�����@%U�8� CFg�	YW~o�*������=�ag�+O.�)� ȉ!�2�=V; =İ3�������B��T7`2��%p�ހZi^"w� �A9�kvt� �C[ߺ'��yҐ��z�r�� �| ޿�n�� p�J���� 6��g�qw�/{~�`�$ꈸ� �a�[S: #��	��
 ��D�*����T �����B��\{ǀ��>�!���(O 	c	iC ݏ�:���>��e�<�%_ 4��Zv�0q�ITh�ǁ_`�� ��X׻�vSr���?� ��ֿFBP�˶/#fx� ������&FW"��vj�� ���!�� ��]a#�� �Vj���� �lO��-�t�K־�z>���HqJpXۭr����4@�\U��H�Q���S}_�"�`��A�mXo�$�� �!��w� ^XFa�Z�$ �	9�� ��E�Ñ{����@�)n��]��b ���S�P=���k+_�e�}l��,	%u�-h�������$����`U�̑e ��7�X�� ��2�b�	0�1�K���������0��#�q-��(��h� ���G$� ����>CP����Y�"�_�N�8��F\�	y�K�yVW7< �b3�A�� ��ȝ�5'h�)t���N 0�9����E	���[� �h�Z���� >�Ʃ{ UD�v��x	�1KՉ1�ɀ���ν9�U l��y�f, !لR@E)���1�"��� vq��� 8Z)�e,�,�E ������ �C��~�u<Y� ���u>���L`�M��^if��0�y��ɍ B!���#<�d3��0�����>��X��% ���R0� �^�2���5�`��\#� h�v���}���1 f'�����Y {�2��r��Z^�*�
���m�o��V>���D8$�$%� S��Cb� mG��
* ڒFU"a� 2��l��� w�����>v� ���D��u	`w���x&i�=\* �� � ��n��� �[hs��8�P�NT�d ����(��1AD	�#h�T�_� ��М�� �������V�D�w�`�#�^� �+)Sz��� M	�
=1 �L�v�_.�P����U���-<�뀀]��'�~��V����Us��u �P�腴%�kO
����ZM^ /E��B��Y>��I-0Ξ��J�����/���hL[4 �RHK�r ������ ��P%����������:����\���N��.!�)�{��;�C��80*��� ��c��ق �Y��B� Ƣ����� �u�ecR� ��tP�(?-  ���l�=0[ ���I�?�� �wH( � ����9��k��,W"�^ ��K�(��� *_������LҖ���k��� �։�^ �( L�<��a����o��+Y��f�Q�H��	�B޲�^�P����0 �x�A *�` �4����=�����I�S�p�� ��	��o!O�+L�p�?��������d@P<{=�Ā���!���O�� �ւ��r���@(NJ�1 ��-g	�b��P�n�0:f?R�8�J��\ #��3e�� Q՝��
 ����IɓC�� ����� k /�!�3[?
���`�N�_��G ��!�|�XQ��1" �_�$[YBPW�^N��'�
 ��\ �P/�&>�L)�%�t��y�b2N��n���z���~�߄+��� @Q��������ǘ�\� H�`V���v M��T�z 5��%�" �UVB��ݥ �^�_�]��|i,�Et�:�@ ��8���[`3^���ı�� ����1݀ Ƭ��;Zv�r7 FA:k�� ��wj�����\���s('� �@����
 E��;�b�'�Y�U RO����[������ �]�	�h`> ���&RS� �q=�~ ��Q"�RB�	+4��eJ�����L P�@���D� z0�Y1\ ��	 �� �
@������}VC�0����c�02x� �뿲1��`�Ԁ'�9 �)��I��[B�ܡ����9 �0�`�� Y*�[�=kS\�C Q��r�(� �%�Rrl �F
]��d�P38���O@��0� ;�X��`.� k��n�y ϰ,Ru�; ���ͺ*:{%\�����.���g��e �rsP�.��d���� ��ES<�� D�ҁ��� �1��;�(s� ��]9@Z ��[Pb�����r�o s7��&j��^�O!+ ��R) �Q����1 O��$��:���2�+>� N �A�fz�p� (]����IP����^�1YX� �׃����,�F�,N P��;� ���ƞ���g���S��V��.X�@��Luِ3 ���� �h�_�\% vgt:�&� ����@1� ���\A� �����  �-�Ԃ� �.j�U���� ��E\G�O���9 cs�&&k���
 ��}x� ��!�b�j ����{2�@��S� _�{e0}� �Y]¹|� �g��)�(>�X�%n���R{>&� ^�����	&b��� �M��4S Z��)���^��/�x���� (���r���R�\ ǡq� ��t�u!�*����	�<:� ������� QWj�@���Ҷ����0�\��(��Z��=|,�GG����v���y�./.p^�% ��Z*��\� �h2c�g �<��6� �֨) �(�L�� �$���+T ;I����޸�������Ư4l��;0ǀ֌��� �%!��� ������ �~�%PׂsX �z�,?�:�X���I��t@��#� �(��'�v�Q ��|�\��u/l��m�� �8z@� �h�_�Ao�>�E/����	�K��� �ZY��<+c`����	����&�,(�`�]Ƚ����tw�`� ؑ"܈��R h}L0�� |� S	W� �x�%�U�+���d|Ș '�/;E�8j�J��"�Sp� ���V�$� K����� {�E�-]��N�� >���M� �q*F0��=S�ϼ� [ �w�`N/?�҃��JX(�2=�h�zF��׵~Ix����ӯ��k��p� ���)��	 pZ���� m�ׁ˵Y#�y�� 6���؀/3�ж%@�l~<V ��aMb	� ,�v���T �'�|���韇U�0K���c���=S 
��D�b� �L��gB^�6[�R�%`����b�S� 4�;W�n������j�,� �$�Q���	����3v	�R}��%Y[���/ Xt(��P<Í�!L��2�D� o��Ǔ@Q�:����Z�_�`-~��o�[A�(�/xǘ�� �
H�eQGX��u��<P-�Nw����}��<_�;�0��e� �Z��3�H-�zH�F ��E������&^���/�F����{� �̟�ӕR F~2	�t �9�\�� v�{J@0 x�/�i�� �S1
!�.8� Ӏ��Z* �V���d�\	�=b Z��H�e� �q�i�U %}�y�.����� �H5K�� ��Bn�*ʃ.E���j�� ��~G4�v%�x	�f���a ��.�s�_( ��/1�~\ ��#@X� �,!�m� �T�%xL\ j�"�dJ��ψ�ɀ�	��T��V�˲��]�� w��|(�E�&+��� ������K
�$!�`��ctInX`��\z��lP�����)Y��R����˥�U�S)�� �D���N�#o���y ���A�7� zQVD�8�� D�SU0: h�6Ϗ��w�	ܠ�4��Œ0#�X�m=�_Z!��Lk�f�v$X� 	�W�u� �|Չ�h c����E� [�:BӮx C8�t�fc/܀��� ����@ �2 �N��|?_]ݓy���e���@����� ���X�`�$F6n� QKD�����sO��'>�B�R傮=Uq;�����7P<�	$� �gX��  w�ꟑ��&�PI	U�_���: ��p
u�� @��[(XZ�<�t�S= �ęG���K�a ���b)Ȅ� �D��� :�ц̀� 0��fX@r� C��R� �Q��k��� ���&9
�~�92��0���h�ė�y���pM�� ���O`����?�� ]80ؤR� �Nk�� 2X��}WȲ �_��^L:#r� ��3�I��[ :�@�6� �J���1S�T��B�3`�X ��A��ԙ����_g �Q�? �� �h���P,s�\�za������ h��b+ ��l� Q$��]~vC����#%X=�d
 ���^ (�����Ɍ �'�_�� �`�s����я�U����#� ����?$h� k�ɒ�~g�,��[�� >�˳���� E  �
���&\� C;QOH�^� /��3tZ��f�� HA�V� ���aD�2�3F�h� ������?��@�a9�`ِ	 0�.��N
�fY�-2���S��1_�	������9 ,l;�)Z �t��P2� �RDM�`'�H�Ñ��%ȠT������nz��
���0� pH��[�zt/ V��՜�� a0�� ����$������\�v�%�BK hkݩ���{�Z[�8�*Ph#�pbUJ�H�(˗ �t��'�	 ݋�c:Y������\?#=�D���0�� �H�_|bd�!�0��׀ �X�'�x B�H_P�F� ���J�`W�_>i%�l������ �S��J��Y ��<�/�nh 4d��~�Ao���98HE ]��(׹ ��K�
����F&��.�2���[�< �H�]���� ��8�>[
^b�'�����0 �:YC����w!�	�Z`I� 0�1ڿ�2����s�"�u!��5� �1�X��0 ���vD�H� ��^��W�} 
�	Y�k�v8�?bx 1˩�UfNXJc ��H�u( RŽ<��� ��b{[�	�z�}���@��� �pR'���9�� T��S> �%?�`��z�x�_�� b��H:�o� �R���%$J��R�}	�X�Z�d�� (ZUA�h�e�%;]y`R,�r{ iXh-���P[�F*�Ǖ�-^��4sN� Y��� >ü�h� �"�G�r�R�@�L	�� �H�!�A� �u?��=�,*�_)��M�/�����:^� ��VO�	�TZCt��K�Y��a �P?��Ou� �C�1鴝w� s�"S�Y\ d)�Mv� �[1�+�X ��ક�� N��	!�^R n0y$&V�? �{��a�r �u;�Q΅l >���^g= `�Z�&� h[�Ě�����
�Z	2�G�`���uR��^-� p�W�b��w ,��@��� ��0�L�S�3b�!�U˽>dm�1�F`x�|��lZ���� ��F.9�$ ���!� X Jڬg�Z �*���pO ����xHJ� R�s3߮����2p���S���s�;��<��$�#��-�`�ݰt� �NP��� �[o�L�C ���Y!��[��v*ր�K�B ���RQT� w�P��H	�[����?_"bN�@��A�{gp� #[Y
O��0=��ݒ������2�J�]� ʳ/�L@Q �)�
�:� �8���X�g �஖/�	vU��-����� ��A �\:� �2�Wqi zB�X��� ����q +���'UK
����)R�;r�= ����cu��Q�?�� 3��[�� h�g���^�Qy��Ȣ@�->S<� ^)F5k �� � �o@]�&��	��2���A;j� ���\��U� ��tYZ�#J��0ӯp��8�;&r�J �@q�)� ��\Yh� �2U��)f �-����P 3Nխ F�9Cw)] ��/k|ז� ��	GY �;�(� ���Mj����&�n	�LH� A�`-Z[>�V�����nU�`q�J	� C�Ns�1E�.�:� 钋� 2Tb�g^;�� �V�W�. ��������Y]�HZ� �i��J�8A� l��$�P2�@�S��`�R� ���`���\��I� :�U��p�G8@
���� �wQ�� &������1 ��[H��V :� KW��� �P����&�� Z���FG�Q�{%�R^ f�g��J�8 �e끂�wD�@ �Ҭ0Jh> �6�ђ���~V Ծ�-���. �;q�4bw"�ɨ@(�1�%��~���by8���g 2�q�a�@ tV�^]�|D x%[	���� �,l�\-� NK#�e! �|�y�ɻ�s���@ðb�"�� F����]��?���SxF�� �Ͷ.�h� q�#���Y�@n��]�x1�Q��g�Y�~�%�m�A�+ qԎ,�$0�UX9r]D�*Nݣ�! ��Fܡ�x�%1ڃ�C��v� o�ߊ�$� �M�f.5��ņ�� ���+��W o�vh�h� E��r����~5R����"���Z 'Q�]�5,�� �L\x0���C�ɺ���B*:±le�@�W ��(q�v4� 96�ڴ0� Q!���b `?��"}����#빦$N��	,�Y �� T\ ������ }'���F��� #
݁��&pT ��)��XZ��J(A�Вo Ԛ�04��n '�aU]� �����h��Q���ɇ���� ���ή�k  @ˋ\Z<fS��
� ��;�� 	!�o�VpE \P�mK��z�w^?�H�#���� ')
D�na L�-���� ;����(��X � o�/vx �Yh�DFõ �jш�8�	%P�����2���ߞ@�RpV�Ħ�[���	� ß�1�0�a�p�� 5e��� ����Q" �F�%�s~q�8�ZQ�,�(�<�߀��̶�,��+'�B5��9\[ �	6!��e�@h�7�� d�f)���� {����� �0 `YD� �,�/R[� ������������1>NX�� h�,��� V�����O������� �P[�X+�� !ف�6����ߗ�C��P�$�Yp' �(�]��~ 2�zЩ����5�-Su��sa _���2�!�
	��. j#�Q� %�25H�p "]�ISO� ,�%0Y�- J��X	�� \��]b� �8Unߵ�# �;,\�&�9���Y�<" 0���G|�ȗ�d& J��[�v0.��C;�d�Y��C �Pmb��
�d�A�0g  *Q��	�|O@�̒\oa �đ��*�b :�f1Z��� ��GBt ��_F
 �TIw�cWv! �䉇����x�r �N�؍�`~ ��1o�� �i])�� M�` �� ���0Q;S��>JU\U]��b �M�j	 ���fE�J$�-Z���+�S�,1��pˬ.d' {��� ��Lh�TF� jH<Y#�e�����\�y�  �� ?UR�� |� P���!Xl'��%�����|� )Ӯ��*Z @��d^$� ����z.�#��@�N���J[p���< I��a���+8� �.!�`����$�P �Q��O>�%�ܳ�)�xA (���*�>� ��� ��W-�qRh��> �l�֕z� �)9�%���C �1�	lYK h�����	G�_ d�WS� �$��r�� &���{��!�H��h1B��� �9�m]��.�& s�Z�� �ς�V*� �uج&"�2.^� 7���H�����c�� �.ZX� ų��z�	 K���~� ��:�TC4 Y٨�����C��� %��Q�� �`�l�)���� ��J�D'�i���B]��=�;V5�1�� ������9X ���P�"� B���U�:����<��s	�]#��Y$3�5�{���p��yy�  ]P��b�� �p�d�rkX6s8 "�Q��� �;�Iu� % �F<��q9��kIt��ţ���(��c��S�}B���q �I��MO�" �K��A�B� �2ԡ�3 ӻ�1�) ��{�5�� >�'%-ĝ��|� w�(4B	�aï ��Y]Q ���c(! H�{$�U	���L J��(� �%���������y�R�� ���K�}�:(�<��= ��TJ"�W ���!� 0��t��K� (�G�ȅ +��/\Z� 	ֆ���� N���l�~ �[���H�i��A"�� ������� M[�S����B U�� ���*�L4;�B�g��- 0J�1�r
� |���b�� ��R��}������\ؔ =���R"��F����QV���0�Y(*:�a9� ��-�	 �Z�e{��|�=IA9l��z �B�	�X4 �m��[�=N^�]gi��}��ϸ ���-WDc�P����� | O��C ��h�[}� t���#�;�p�$�}�	* ��Ԡ�e_� O�4����* ����ݱ 3�6�@0� �΢��P� �!�7��R\IJ�K��� Ê��YH@:�� �85xJ� D�¬�X 	�:����}�	�Y���`qj��^� �0�c]��8 ��F7�� �����ɘ��� p�b�"�K � ���f	� �aj(�n���YO����O: �
��Q�Z bY��m��.��� �E* ��-��ST f ��F����E��ݦ��+ r`��P# �X5�%� ��8@x> ߺ���&��D�\R���}����üI�( D%
ِ�(�zX �1"��+ �f�z	 � (��\�
) �@�����0 �/���͸j�`b �[�̸�<�>'�Ph�.� F�ͽ[dW����D��@֋���ˀ��7	�(��o�+���C0 ���JK�a �Lh1ͪ� /���o }(?��CE��>�u�����p���%�z}	 E����5b�{vy�"�_��j �?�Y+�1 �0�@�_-� ��K�ڏ�آ ��q	�r�_�A�� 3�&� Y)>���8? ����JA��K� <�>������o`0�XQ j������ "��� +=�]>�� ^�ƃv��� �y؇��?�Q �e��E�. �!�1vjB�QTY����֏���_) x�pbJ�a
p��P!��%��0�}�u%��XJ -�N��G�5륀�LoZ�$%�7�B}_ t�Ў�CyQk����!�̴�-����&�C�F��R��	��2���'�����b�i�o�P�� 0?��� N��(�6[l�]�٬�h	 )E��Z�'w �J��!�˙�$v�`��Η���Pf�] n����2 ��'��� 򂰚:5�" ��I�ZB����D���	�z�����0�,�K� ��i�4�	 �wr� �%Q�x�������0]�P*���Z��G�z�̕a �IX��K �T]�C�q?� J��26�RL�UP�0����2�0D��PV�wtR� �7�dW9� 3+�� b �(��y�	���l �1��� ��x:����� &���@� �aT-�V �
�F��I?�� 4R��d, 蘛W����P�E�V�_ ��S�h|߬ ��w��k �~Rbv��MX��G���?%�p调^��#� !z*�S� �p4�=��=�j��}�,{ ��N��( )	�[�PL��P�to�J )�4N[��8��?wd@���� �Ү�,�=;Ú���B��& ^��� ��Kw���o d�c��YQ� }�^n�V� #3U�;r� ʺo�vb���j�����xwi@�>�ˁ\�+������7���A�`�n�	z�@��7X�~� Ru����wD=�	 �{g�G��K\�޳��� RC�	�Q�� �s9���.& 04�^���`���ZNcP����B����h�n�t`bډa� U)�(/����������;O�3� 	��KF2[ ���PH 	�_��188, K���Z�� `%��/�hH�#�Fg��p��� 2'���% �=�+���$�c��MgHB	�� ����[Z�� A��;��j!��	�X@1� �R]h��#}Z��� ����ԝ�i�?q���x.P���z���ry
o0� [�< ���k�N� ������K ��0cҸ'	j �����f h��P/Q;���Î���ps~8� hF:,��+�Q�DPOx� �3ޑ��×'���Y �52�=�� F�[^�̓ -umP\�� _>�vZ� (�
%fX� ��h�P;�aH�������  v��H�2�� �R	�;t�����N�c 0Ҋ�H��[�/!�1�  �ZX>%��}a���ПR HP}�^�s /0�+��� Zl����/ ���cs�� (5n�� �	�a�!&x J'QCch�LW�U��s �I �{}]� �f1�Xk h�Eb�'W`�A]���?;5��*���O��t~ òX!� @�
����:1��h��[  �YV��&.�]�~�p����U��S��
�p ��u�Q!�U"�A�+�1w�,<]�	���Qc��ɀ�`à;��� �D�1���� �j��.��:P~R�Z?�+���H� �+�Y�x8�i�< ��y-1$ X 9U�� PZ��]�����)���K0"�l�엾�p��@�[���O� �j-�CJ�	� ���&�Q��W�`��	 �^�t,�.�~� ���*؈ �@�Z(T���- 
�鶬C�� �$Y����ø� �
����t0 &)�8�;� �.����" [Ѡ����������2(� Qa� |F~5��(_��UnP��J 8��Ze�s�N������p� ��[ʐ3N���@ (�L ��hfr�� ���'6W� �
��߽ J{�(���� �0���	�'��(%<��h!9��0��#��� �'��p	�j�>@h+;�� η\�b�,��	.G	ƀ?�F$� ��[J�� ��! ����KU 5H#�Z�8A�ñ!��I���3�w����r��.�r ����I K�MQ��0 �g�_�Jv:�tnR%��\�� PTX����f7�_@��-[ Q�r
3ϝ� w�I�g� !C�o��� qp�w_I�e!�� �)�h %�D�>�f]�w��*`�	8�ݜ���@6 �t�PR�� ��iC�Zc&�k �P���1����W�� D�Z� �+��a*@�\I��6�S�`:��I�{��0���g �B��z�β 'yZ�� ��a�� :�����F�P֨r- �Ŵ��m�.��� ��̸9 �1�B�	�Y ����t0|�����	R��`��cHI( 2Z���<�F ����8U
}5����X*=�1 ��a(G/X����@9��|��Ȫd��z %@��
���ce��`kȰ-_ ��Uu��D ��2�yd� S�n[a�3 :�N�����mA���{�*����\�2
 �v��, ;�̙�N��u9@s !ؔ�i^c� ��,C�~ �ؐ����� �Ej-:���.Q����V o�_h���xv QS��(���}� �D��Tf��G��j�}� �|_���� rP��q�� ���^QAi8�B KCP'���X��	õ�|�l�ُ *y3_�ΰ�>��˶�M� 9���� �_
�[d� �qԺ��T� �1*��J �U�t >]Oպ��n ,������q���A�0�Q��1mzZ������
p��i������z�jC�C������N� ��a�V�.% ���j��0\� �K�UX�>�h�vO�  3Kۮ��N�#� 
����;�!&�IfhT���B/ ��D��W7 �r	�[#� �<;���K� Q��8� %Ye�W�q�	 ���_1��'����&W��0 �p~R3�� ����Ѹ{ ��[;]O ��e��֢� 1����XY.)л r~�E�	Q!��s�5W��%�s@��� ��)�G$ ,2�<V3 پ�fѻ�u �����l& �_�P!͸ 1�"�(�i �A��'� ܙ��q�m�8��[���O��`��K�J�>w��k6�=\߁�0���,c�$@»d����� ~���N�n�ݟ�('��hO�-	Ǳ�k�.��"
��� ށ��@�)�� B�0h7J% $������ ^�A�8z� ��0�1� 4���Z�R�����F0�X�>����� q%p���1�]\0��<�� Ւ�Ѷ������́� ��?
|  ]BN��I=A7 x�Qd�n��� �)�~��F b¼_N����6X fS!��y�), �p7 ��ܝl  ��/�3?
Z��Aw?��J�7��n��I U��ȵ�OШ����4 ��\ST8_MѲ� �-���G(�b 	ƀ�k�&� ��u$N��/��R�_���x�( �:,��QP�90& ��	�l��,�
"� �w}<#= ���͜X� r��ʷ��] ��wV�S ��m4�\�ʤ��|ppX�0 �e�*�S8���.f��,~2� -^����;��C�M��)�� ��3��! VG��W���_�M�琻�ǎ*[s%���#��3� ��~��P,��u mC�� ?HO�+B� ^�_J3k 0�fP?���2,숯 �%R�[ �0|wM^�	 ��ۅ����������S 1�����2 tʇ@�� ݐV>ɜJ�-�1���h+�x�b�]��-B�3	��!�� ��� ��=�'���m�n �cB��� yj'���( �\���-#H����,�|����0�"�5 `^M��ZS2����Ӏ��h� �
�X�� ���[�>�Қ ���ib� jɋ��f�0�,  �PQ�=��9(H�'r0��[� 7iP��� ����z���p $*K�ٖ��qvE�� �#/��<���$�����Ə� ��0���S ���ϻ P�� �1�[L��܅ǻ}�ͷL �cGf��� :������o �JA���' +�h$?I� "Z�1��l�� 5����m� |���*�?�E�s�3Z̶�	b  �~P�)L��������}E  �P͡�@SO ��B�XQ*M ��"�_ơ|� �.N)�wTD� �9*�Q��%}0��1aHk}x!X����>�<�i�$"�+��͒�1�����?0 �M
��G��9�W�C��9�1���L����P�H�@��{$����}� ��K	݃�� ����= ����NK���.*�4F:Z�$�<�+�ؾ\�% �' �w��	 �XpUYZ�N �\�"i�� ��.�� �(*�%�-}hѝP A1B�{��u0�
\�(s8��<�, �V#���q ����= �Z�L� �?X��5�B��2�Fo��} ��~bS� �p��� �E����Z *�)} �Re6P� ���o�m�iO�b�'�pQ���_��7����
��(� tωr��a�^ �ҕ���%v>I`��L9� ���˼Zd��)vW���w�V�g!��fh IK��8�
uEa����� �Q"'�V�@� ���8c�;N ����JZ�}� /��!��l�A�+���5q(���{�a��R�4 ��Z!��> �VY^�� �x�k�[ !� �~`9��C �B(�W� tK@Z�X�ś�Єخ ���Iy$ �`�Z<�m}�.�3 ����f��݂P���H� {���.Վ �ro/�=�� < ��ĵУ�+�f 3�^t �,�	�SU Q��=5ʆ�����*�$h�1,�o.� �+���\�0���H 
(�B��u.� �5j��� �4�,hl-�=��k'  �� ��B��1��`���\x}
Z[�Ϯ���?� 2�P���� �i�ׁ)��
o�FS&`�c�}����Z�䊒 h��H-�N�@ �;�*:�26ń���ıKH c�D�%���$������ ��KXF ի�*ܿ�$;3������� �dk��Y�@�\S3�	 V�? ���%\��ő��`ϻ� �E�h�i ���n+�X �^���� �x���A" ��aJ��v;^C|�����e��~����0��;�8+��$b��� |�6�0J(� U��L�ɾHZ�`\xn��;^ ���AOk�c���	��B;��N" �}��S (ሐ�,ɗ�;�� "R�&X+g�(���3�T9D�@����;~�@�� �V1�ۼ&,P�mԎ�� ������ ��ت�0�X4� ����@x(p��W%є���{ ��f)�̵��/������|� �2��l�K|�?������ ��$�������0��?]��ُD��/�e0Z`�G����w 1�]�IY� ���Ύ��K�S�s�𢲖�ȃ8P�^ 21Ffa� �`�A�{�L��p`(Q��s.fYs ����N�E_Ó҃3�]h�^���!��;���8�
�������U� ��T��)b\ 2[Y�uw�$+��U���S` )��=���� 폅YD43+&��` <�WT�I �����}��{ N7��l�?.æ�^�Љ� Ɇ!:�LB �� +�V�}�p�A�; �o�q�;� �1����@#��5z&��� Y�m }%���)8� �r1� �>�] [جp�f��wG%
5�ڄl ���7���)w����a�s ��\h�I 	��k}������u� ���Cr' ��g�c� 
O�<�"	�\�U��0R&0� �lN=!~ �����'2 �1h@TNi� (հ]%w �fB����1�-�މ�U�wF��P �t��0K�_�\9
�u��rz+ 6��Qa&*�N����vPְ� _����"�� `����� ^��lr��t} 1�Oq��<[��o���(҇ �ڭy�T��Vˀ��f�X^%���·
b� $�EԘ�( �3���l,�p�@��-�Z �lad% ��82����b0��Ǿ Kf�=Q"��� �ӛ���������,/�T�sZpEp� l�^	��{	,�ߊݡ ����h~�+�W�2� �K����E
��t��3 �-!n�@{� ��T��.\QU@ rP |���� �͗�hcCes' �AX�	��.��; M�{�$ �B���R� ��E�K 0 ��6_O
� ��|��2W���}S���Ps��zo� � ͻ�+��"�@8�JM���^���SL�ͅ�H= �� �4f-�~�9��S�k@ޏ`,�� >�/�U@Ɋ5*� P��`]T�1 �^��hj �e�u�7a�Ƿ�l2�җj ]R�:���� +��_47�)������V��@ ����$n �H]�XU, &)d�-p�q� Z��h�}* �����$3I�	��`e7�Y 2��ԏ�`�
�� ��L��W�9O^�����WX�y l�Țk��=i�����QY� � .a�^ �/Pୀ�&ZX���㼲 C�h�13.� �Y
����v ^�%�՘ ���
ʄvfy �S��pԿ�8� P�RG�������p� 4&�ͱ��� �J��(} �^ר�` �SAB+����0����6���G F5����)8`�a��j ��*�g��D���7h��#r���P9��M�� 	�[%d� P
��p��� ��Fe�!� 4�xL%��� ��=�1g �*Y����D�N��K�}��UE���X �����,:ޮ�A!�X����(��[�}~x��7��j�n�YB�=8'��T��E��; n�� ��7��xX��.�`0�~�	E���|$�Uu ��u�ip�O�T���w�%�o "��f��ϲ V
�ͮ(���t�v U0ÿw;�2�T����m�, NJ��ؗ�]��!ٓ�0Z\ �:Y��l; �jc�?1�5�,�'p'*h�i`�	�`҉ "ٿ?9�a\E� !�F:���[ �<����0�=��&P�P ��� <v
 ��1�."�� �ڈP�� ������ � ���ˈ�	� ���ߡ� �Yx��� C$R�W ��0h*8
�J������g2_�d��ȡ( �0���� ^�
�]����O���p f�Q�U��p� "0����� ��7�A� ��5Uk��� ��'!��7��q{� �_�a� ��
��,� ��`ʹ?oSW+m��͎� �QAv���OK��8�k��+*^���I� �d��m� (�� 	���� <Q��[/}���
'"� �:��M�q ����/�#��?��ļ' 0���/U� �5����P�v���1 :����o� -�UB��x�+ \¢�]�m�̾�`һ`����|��0��$eX���q�� ������(9��k�e\��%�� S���Q��;�j��L��4	1�Zu �0/�( �5����B �h^W۾������� �&�=q7 S�4�1��3 gU�����7 Y[2~�� -w�5N.�� ��X�#n���Z��u2+� p�[Q15�Y `=�V�8^y�`�� �W!�j1&�F��{E�o ��R�O� �X-h/�x� !�,��ͦ�;̶ �	Dpw�Z���Uq����P@���X� �_��/�v �RQ�*3K0��\������.��z1� ��R�?~,��" ��&n% \j'�h�0a��	�` -��2��r
�X� �Q�\긮��U9W&Ц���u���d<@ ů��,�� ���!R�q ��ZPՙ�� `]а��� *	E݂�� ���Xvӗ�� �
9b��;U�AҒ�c.�ܝQ ���#�!)���Z�6� GL�1�/�*� K�!��8| �̲���h ��,�DN�r�!� �v�p�� G���'��<<���� �%�B�h �[�`W)�,��� ����]� ���V`*�h8�^�Ƀ-�����qd \�8�F�{� ��=��> ƀ�J�ԟR_�-�� ���/�B�|� ��:yd!� ݁�<����B���[}� ��i/�_� ��H����+:>� ^���AL������� 2�S�	��� �/�&ף�[_�`'-x=����s%o� * �1����&70� n"\��~� tVD� {*UƼ����'��B���:�|0[ � 븙� E�]��	��t���5�� G '�mw Fi��� �n���� �2O~.|y �Ch�k�L��  ıx�� �8
�&(� ��fw��� }��#�R�O��Wa MO�#:�� � Z�����80-����a����[ �%��@	 ���DZ��X<
����� �S�{�-��x=� �KC�4 ��v{��n�x(����ԉ�]\����&	����#g��� ��h&+4	�_��,�� ��azR�S 	��~1)�� ނ�W��VH �"��3<� q1�lj�?�Á�d8�J�3��(�}ÞM��	ڝ��,\�hL� �e� EM�l��	 (���0�?��1���z3�2mҪ��������)}b ����J-�|� 0#K'|�u< ��,�}�� _!Oȿl� +d؄�s�C0�^�jXL=Y��H�h{I����!�V��%� ~Z���t���}OGe�	U�o/�Ld����� 離��t� E���v ���z��n����MųҁQ*aA�Z�)+�|TY2��;���<� �y$���(���@@"߷^M��-`�h�/� �����ap �"� ��Z Kc���{�:��<Y���k>ϖ���@��]H���G:�`��[0�\�]��x�k�@ԘR� ��A��W��=�{ �ƈ�m�>0���2܁�. �k�� V�T���W� �	�Q���xgʁڼ�e+ �Z��a�"R �.�S~2M>ut\@���+��%L����� �\^���zJ ��e���� X6)�&s �j�9t'h	@ A��;+��"a��Kl ��D�� f�~"�0 �|O��R
�?�g����j�\h�3S�1�y���V
�'��9���U��d���S� i]v� �D��TY�r�=��蟣�Gݳ������ `��J�!#� Y;��.�1HSx�,���(:��X�N�Gn�{z��gY���KB Y}6?��{>�I-=a��Z X����� �m�DQp�NA0�|�� ���ɾ� �> C)�<�Rn�4�p��_pNf ��m��>�?��c��ĺ��B@JUH2�Fn�N�k�z  �ah �ђ�o�<'�}�wP��$ ���gU�[ W:�w�r0�?�T B��- ����K��%� ����Nѐ �O���0q )�	P�([ ���F�� ��	b�����Y� �l۷q�2��w���0L�W�M����9����7�k�3@ ѽ�� �}+"��^�V[ �r���)� ��x�� "	�P�\�� Nh��Ky��J���|p ޟ[<V e� ��N�~�P"˒
/��w�����X���!V�H�	u -L�P?�T	 Z�O*��i� �r.~"/\8���J�50�T�;� �(<�.�� A����t��w�H�*�@�ӯ���G�"��� �FD@�R� �`4�� X�t��[:����/Oph��I�p�KH��M�?Y�_�����h^ �t3�/� ����������W ���+� _��g�H� 빪�8] 2Ψܒ��?j� ���C� o2W��[�Z�4� V�\�h ��w9�~f&�u/7��yv�h������ ��+��' �Б���=��DU��1�� ����! �)��� �EU
��d< �;�x-	�8 �W�N}�A �_"t��G ��|�C}� (����.��H�� �m��w���%� ��A��;��+� d�Z���
[����LO-�S!������" ��Lӂ�� ~	J�ʟ� �%�i����{� �݅d����>IXW�T���h .փb�I SeJ2ۄ(�?��&�� ��KL�� P8`(�h Ht��[�O�|�ֺ����X��K�� 5�WZt�A: �do�&�K!���L1a��z���;��Y�2�K  Z��b��
 N����H U�(����p��� b^	[V��� J@O�q0� �c��ʓ ,�	�
]��h� Z��N�  ��_]�� R\P�2�^ ��Hh�F���֚�92� �ZfQ���q6���	�Phr~I��$�� ��[1,!�V���h-���y1 ���f� }l
B�N�� O&�J%�:^@�+�mWG7>�� ��l��a� �uƁ�Q� �0�;�i  ��"��[� }~0����p� 
�a��R  ,��� �h�WV+��=��2�#�_��ۧP骮08 U�m(R}1 O��k��0~��]��
��NF�0�E a�>�ƌ��]�ԃ�6��8[� �zQ�X�^ ��P�椻 a@M�
�2~.�R� �y�(5�oh� 'sѿI ��������x ����3 Y���h<�x� ���Z����f����u V7uK*�
ز�����Z�u� �� �P.	�y��� �Xh/�g� ���+��%���X�p�� S �]qg#�� �8ޕ�&�)s���Y�`8D �V��A%)}� ًpj(� �O�l�T ��˂�2u�;�J ��8]��� + �XP��0 Hʽ3�{�}� @���(��0 #�b���& H��5D��~ �����O  ��ü	2 ��X��W;L$ �0¥��I A/���P ^-���Tq �����Z ��@_�#�S �-�3n���H�c=΀��@�0ѐ
,�(>�|)�r X#��	�� p��\���P��k_Z(����\�� ��Bݷ[
Q�H��)	Ȉ�Y/N����W���f��*�	ڴ�����#h�9��N�8
��q�.�Y�X �L�E�p���O�P b� y �<����� z!�
�hR �t$��^\��}(`��! ���-��/ ۅ���� *�����(�$ �u�D�:��0�=�� 61�Q*���r�t��q �]�f���
(Nٟ�O2��WPI-D�j l�還�r� ��b�{�" �V��N��ij*�bf|�^	�� de��4� ���[�z��YZ�@��1�� �	ha��+ ���k��C� fN���
�x ELQO��&'�>� �	l0�e2.{[��@�a�� (���Z=��p�CKšp�Aa�,FG�Q�-t�@�:ʾ �J�^ t�f)�B�t����h`5/}2 OJ�Ci��� 
��M�l���y����
����@i�"���" P����W\��� �Ȓ9\O ��	KDYi�U �)�-�� ���$�k� ��W�:-7��0)�U�f��t_ AU�z���0[xlX�BՆ�@C�@-��Q����� �yhbU
K� �d��2 ��j�)z�6 Bl�]����:��v��"*��W�=K���p�� �k/��[��賀P��+!�@�	Zʁa@�%���18��K�� ��G��� �y��	� )3��/[W��QiX���Ff�{� �8�+3L� ����> *�aC�֪�̱R�Z��g��X�j B>o	e���S
���i$�Q9� ����r� w ��9�� h�(]'�S��� ��� �� ����w� m�4_
�}����ŀ�К� �k�NJ*�� 6X�[��n���@�$wK% �j7��!@ ��]hI�,P��� �����	 -q�H5�� ��N��!�* �8��wQ� ��\U��K�-ϱ}`C%�
\ b'��}�� *ho�(��/v"� j���
����s�AT� a�XF� J�C
�P�拵�}`���� ��@��R}�{1�� �y=��օ��/�T`� '�Y� B͡/�I� �9�C韷 @b�!$(�� I��\	Q��g��X� �������Z� C�z�%m d��	G�$2��� Җ��� �N�aj�1 ���G�<:$ ���� �,�fj�> �}���R3�T*����:�9P� �(h� �!��*��w�PC�C.�6���Y���т ?��P M1�Y �� ��W��+ �h��_�O 9O�@Ѥ[�A�
�~���I0	��Kd��ܾ�+ ��Ss�n��^ �_(ދXsQw��b E.
o3�Z�U��������V 0����^� ��]!���n�@�I��p� �X�V���%G�[�yOM�� XP�+� ����$R8�� Q0��3� ��I
�y )$'克V�Th�� �\ �G� R�� �|'u�d��z��Ԉ�*�Ƈ_�(CO�>��J$\@i �/�	"H u|@L�$�-��ʋ��������ǅ `���q���8�\�,`' ��������&�? ��=) �^�L��J �}�%tI�� 	!��0�&��I�%���Z� kK�鸟S��q��{	+op!�']���Y �������@ [g�5}B ��鍽��X ��6%���` L�鱿 �'�W�}� �X�1t o����* G��	]�%�� D_�� ��8�	\ �˕d�0�{�h��O�I�k ]������ %0Mw���w� ��R��� e��!^�A ���]X����@t�.2N) `DZ�'�;|�$N�� ��W�P ���|#�K����Y0�� R��ʺ~cHa���
`e\/�y��`�� ��u^h" * ��� ����}]���_�b4�[ n��)�`�R.|5> �Qא�� F�=P���bA��"��a"�Y�[)�r� �HS �@�j_��>�����-t� � �����]�� �<�_> 0���t�\o�x�^@��f�� ��6���5 ��ب�Ov ��U�X]݊#i
��D~�l�L�����������S��OЯ���en蘴�`���x(@���=S��Ýhհ��k� A�c�Z	��"Y v=@݋80��X��G�� ����^�-@V�,�ҦD K!����\� �ޛR�� �p��C�w Ϩ�6�F7� V(
��X?= �����_�2�= |By�4-�	 r�%��zz�T�։&��4�x��0�u���Y ��8��� ����ݔ���6 ���+;�1OwX�2���U��� AB�S*�f��74�PqpW��섕���0�' �X�[�SY sp��#�f���  ��ZhY�J`��r��B�	������ Y��8�� ��' �%���?��}�Xq�\ٰl10h:yb�w�ا~���� V�'>�� f[ �Y�9*s; @�J��ܞ)�PK��-��Zo ��¸���<�Y!�e�\��5 �`"��N�LK� ����\ `��^��X���R����S�~}�����J- �w֩`} ��ge��x �YK-W�%���C�I),�|[ �*�d:� Z�?�C�':�ǀt��<�z� n�P���� 3�
�և���T S;z7	�?��(�_���!�����r ���L C�@�<��#�៳ �޳Q|�P����~|8 	 ���SB�º�li�� ���z�-�u����n��/])�0��S J��i#���, �t/�|<�� �RͺD�P l��ް�F� ��̐�%B@#?4�pۡ��.]�g1�Z� ���W�pX hUa+���	:�R���;��,��'-�����_�	��ԂiH��.K ��g��0 cw����-[l@���+L�u��� 1 �� ��U�ȿ �J���*� \P��ޫ�.8� 
�X0�!{� h@~K��R �O:�Y� 	�A\��Q��� ��9�X�.q�� (�gS ^�"jK��$B� 
���%��@��0j�`�t���� |�*�	�W �g3��%@��2}' �����
� ����\�{ӱ�!p�tPp�
 N϶�2��
�E���	�D1uLş+re}���sd�$��L��)� *�]���� ���逧�X��U�	�%�WKN�^r�X��(�� ��k����8�����zĠ� (˽2u{�/sF�!�3*���N �ϻ!$6�8AY �[#�a�����������=�.�$�`7�; �q���(����� H\�Z��� �d�R*#�x[?+������X~�p; m��!�	
� ��ʶE. �W��Qۺ �he��0�� _ ���o*t������;K�8R����p����&�S�5`{ݛ� _@+U��[]	' �Z �z�� kRs�/>� G]5�K�\\-� ��N�C�� _$��K&+	Ѱ���qX]� �1�t�0�� ��ܲ� ��U�P��):u"���\� �bW�4��7��\n� W��A��(����Pn .�0�LKV;W� �4�Y�ν ����� q�&��e+H�$@I����`Zb@�5+�L���}�Xd�^��" �UNq����J0Q0��)����� �d��Ɨ�󩿒�u� Xs�v�Y,|�� �g�%�����,� J��
�0�[���U�� �S�b0�o ���G3�!�ȹ ��W�� "�]�Θ�� �Q8�*� � �AO�y܀ �[0�?�h��Àv��>�4j`�~��Z���h�e�� <�W�[� !�0��a#�?G���9�D� _Q����~[�� dr�U�&�q� ��[���x�=4]��@wU�  Ka6��n �=��S�� ��c�^	� p0[��Y, *ֵ��� 8w	����֑ ���<4�������W  ��A��8q ������I <�1���Xb 0�(ɶ�$�t sf3���� �S��:QP ��ǈڰ[��G�Z ��J�µ��-���	� 
����Q ¹W4< ����`	}���ݗp�%W�z�~̏ ����H U_�u�h�*%� ɓ3)�P�� X���F��� 0�_�۰vC��Ɓu�ߺ;c���!���� ����K�.hOZ ���� 8? �y�� V�ʒ/L+O ΂CY�:Xh<4�I�Q]s��+ =���JK� ���|� ��@�j�� ��� �Ĉ�^j��1 Ɛ���	#�8��x�u ��3��	���_`w��T�
�����@"�Z �%���� ��0X��ݱ ��#��'�<�ۀ���`� �/� Y�_���:�����T�����W@ 0ԉ���\�8��Y�`�� ���ҿnߝVg@	8�s�{���bq�� ��R�� ��� @) bN�y�	���dދÀ �����-&���'_ B:�P�꾜 !�L��� ���1sx� 2�_!��8 �N1h���0�F|� ���J
�}@hZ��� �ݻ"�$:*g �X ���� ��7�(�B" ���! ��A��z-}%�HP&4��l *x�-�@|Q �I��;�� ��	T��' ���v!(���� `�` .1��eo;���(�	 Ɨ[���Ht�;� �l��� ��	�
1���o`��# ����p����( �d
�ڍ� 3O$��['����.�>���f=Z�z�P R��c�A� ��~��G��B��h��,�>DN i�S*ӻ9�z| )�d��E�<
�a��?�ΐ��!O�`w,��g����Ll �|\F�S.�, ;[�� ��a�k�)�8R� ����n/� 
�g4� � $(��	*� ��.������ �k�:�J�B�ty2�� ��]�\dW�������t� n`���� �Z6�!���\�1@�D w[N
�89���}��� bP��R)
��3R?�x10F{�$����I} Ξ�v��kŖTGS�ܦ�0(� [��F/.�� ����;P �5���%~�AU�V�� �����& ��vU�O�>�S z�:{�� ݏ��[��w� �ز��3 L�Sh�A �D��P	e��X��p-���V6D� ����� F��؀�J!"G�����Z[){�4B@	^�n�s <���o L8]� ۴�̻Ns'�����, �H��J�!҆Ì7���^��[@�7L
�.Ho ��0j�" ��ŻZ� ��S����z �$��'w�sq��~Kb��� H��)	 �e'?&B�*�߂��_�y`)t&���( �C���S|�Z�v,ˇ /��!L�D�p0��CN��WHϸ	�"�F �/�M��Rոa�{�G�GP�y?X 5[�Űp�x� ��h;oc�r ��K����
 ���9�%�_ D(��	����?d��. ����͗�V����Zw1N��_ �Y�QR�������Z ��$��¬2�� GY��^1��8�a ��$Q�9�JLu� �����i� ֧ݖ�' `�/��d�0�Z4���/���tH$�a� ���u�� �}�ÓU�+�$%	���]� .����Ř� )Do���� ˜��p:[��~���� ���h%u�p� ��nV���Yi�H�_�p��R=ŀ�,�'� ��I��m ���@ג�. ��5�~�K"_��߫��P��� =����^&�����Zu�@7�ǽb}D�| ���h EsIl���#��= 	鰮 YX�<�P��=W�����2G �	Y�b� ��KM}�zA�����]�t���~�xhb؟� k/�5�*u�`���p�p�� �F����8�XK n��h�� ��v@����8�^S��!�i 1$*�R�B Dd)���!WA.����v,7�V;��� !� ?D� [W��p�� o>�w�'^2����FR�� ����ڇ O�M��2�B�W�IHJ�*�>��^ ��GL�P[���&gQ���; �c ���`P� ����� �4�2܄����Q�H* ��U���=�ٓX� 9���3� *d��-O��=���/��߳R���Hڿ�EI�p!�� ��|�G�u� �k�J�� �R��ް�s ƒ)	�S2� UM�,D0;\9���\iKs �H�&�} 9`��+�.�b�:�z�� 5��l���}~�KЇ��0�%�>� ������X$r�����,�V�Śa�G�s �X_�{��� ���	� ��P񮸔 lQY�:e)� �_�>/�� �%�W�9�x[ D��4��S\k����Jq��]��0��{�� �[֗�� h0�>+��Ŗ� "��Ұ {	��tL ���r�b Z�@X�� 1Ç�Q�0�{� t�� I�:^ .]�Y�zN ��/_ER������ ����C	38"��|�Z_ �^�ON x-]u��&$�
i 6T^��.+'lc�BR`�]�X�S%�p�(�r�@� �.)�ԔXaL�>�g ���`�X�k����ؔ�YB�J��z@��- �s�\�� �4d�S��E`�
�ƥ� 1�Y�J�I ]��3 ��A暬 Qh�e�*�� ��C��FN���;��1+ ��.������*�j�VQ.�� �@q<��� $R�`�� h�gH.��� ��	���|� {����tB�)Rg ��[� �U?���� ��ɛ0 �z�<�Z@����*��T��B} �)�p�� �yD�f�[ �А�}�� �n�"<x��sP�Նp� �fRP�5���� ��	J��X� Tj�ȱ��;_���W+�߉��k|�g�i ��u �m�*��_"$�	� +/r
\<\�Y@%)�H���l����$ ��['\��ߋ"~z�0�!, ȃ#Ɛ�|�R(V�8��P�'�����Y�d[ ����> �� 0H"4.Z	 ,�'y�-T�h�~���%�L���v� ��.F�\��$�: ��{�	� ���ǱI|<����8
R�ڀ<S#�� u�k���9	 P�$�V�� Yq��y� H<.��:�.L2� dߩ��Q��$e���#��0�Z�H}�@�c��� ʠ�'�� �9�YW�(h.��� ��6�<$�����@��p/X?\ 6�5QA� ���G��� �U!M�\y<3�^�	p� �i �����Х�� ��BV��C	_<w0��N��Ƙљ���� ۅ!(�U�7 ~_���+������ �Q3��� ���7�Jr�Ob��l� %ɴ�؅� k����T|�8 �ifS�� _e���� �`%$�����8!����������,N7?t	F 
P"̸>���� � ���?�$Z� ��
A���vs* 4blIV� �o	���s *�Z^��p%�Q��i0�FYSR�l� �ZQ��(� �遟�����? ��Ƴ$0���5h�����k >�f���Ը ;�$��Mh����ٸ�8u N�dV�w=Ĝ P�_m4�  U�%�' <�
�7>b� ��`Th��# 	6vL����ٴ���YI6	O��iyR�2 ��&e��<���ϟP̠0Bk;���r���z��O��/�R� 湫�SAa9.(J���[+�����xm�~����:k��� �%Gs@���9��h/>C�-��q)@Ӂ�_ Gл��L� �"�W��-��VI	h���($�D{ �_�> ~),r�� ����B�;�Q�
���>��a����*� lL�i��ܕ%x[��H�-<KZ��� 5zh�k
�� ��/_,��\Z �Fε�7 KX�f;4�l��P����~�?� ��� o�aTX[T���~���`0M��. ���@������,� w� ������O�������� *�^J0(��S��?*�.����� 	�]CQ��! ��w�2�' F����������*�.3� �Y��[92Z$2 ;В!�
�{0\��R (�|�@.J���Z! 3�W� y#��P���%�����S߈. ��bN�^X	��`ؖ���*�O ����� �/9�I�z����f0�E_|S����2J ȩ���	B���( ?Q����� ��k%��|�������H~;P��S(ɍ4�9� �<���	� ?Yt�'�l�4=����� ��P��X>l +��[�� v�Q�h�����ԃA�`�K 0�?�^�)��Ȑ��*zb�������l�  �Sutf
B(��� ���%����\9]R�	iJ 4�@� �S�pM�*&�Z�����B�1��Q_h 7��>[�	L 
U�\�j ��P�/�� �X�^��-�n���f�1�> a0�G�ZX +�������� p�`x�/�샀5��
�d��N��@� �1j��2�A ��f�.�C %㥯k!Y �m�	�����-_(�h�A�� gK�� �e/0!N<�T��s��P) Y젥��� �
�@ˉؽ;�� $[�)��� �!	��tE��/�0gP ��K	
�� 4���~U �R�\QI�H� �D
 ��"�!@�5��D<�Pt ����! ø��(�  /��$i�8Z�������*̈@'�Q����bj�������	o�z�8Kn�0��UT �v#��/� �4	���\��,-�߰24�R�����V�qU���!`�� "?�u'�: �,�$��0?ዀ�s�&γd "i����A $�O�q� j�Dc� rb��5�� "���Հ���N=�'>�r� �[QU�� ���z\R ��[��Xm _ȷ������ >Z����+���P*�t�R<3�&D𸈳} �S��~_�| ����)� 0�	�+� �=��O� ��BK�ŀ ����N��w� �R�����{�Lk���-�X�b� Z���: �1<`�f��yդ�� ��-�|����\la/�R ���n���� �+��Cr%�P� ����}Q8Ћ�z Jͨ��2 �+��OX���0~ ���k�^ �"@w�	��r��lg%�	]�L$�B�6D	�����a�I 1gx�%�+�8y� �^����5�{]q���\�'���ہ���v�ξ�� Y�@F
<�N���� c�H�h*�� ��)����^`�T�y/ c���w �RzQp7�� �1	@��,:��ڳj`�[r� ��XV-�q F/_�����=݉���A�G���Htd`��� vl* �	�w�`XN|�C��#�-�d�y������h)Ua�����*m �%}���H@����{�-�WV��0�vf@����� C���(	� �9�@%͢� qk��y^�� ��>�c� ��a��;��&"P ���䝄 �)���Q��5B]�����-���!�.u h$0� �6�[�(c�~ �x���% \��E,J� �!����(]XY^�+a`�I (�е o��2�V�� �W}q�&� �w@���� ����4*� �:6�$�N ]�DG���� ��Lb˺ sq"�&� �,X�Zu�ː��l�v	>�3�9�y������^����"��,��� ��_^�� �̨����- GD��� ��P���(�鳂�����Q 	���%6@yaj�* 3�" �;-��B�] b\_v��M� ��[calJ�� �����1�b�a=�� !�(pD� ȈX�81Z� m���� 	�Q��u> )��Z"�Y��&! ��|K��� +�N��˴��W�� ����� \���~5� ���$_X/�8(Ř����JpVZ �v�u�$n�= �Y��!y ��a@��lh(���P;�>�|�t�\ �0$*D%^�H�L �<S-�����r� P�p��B���H��&ƀ "��\���	.m�q�� K�ZŮ	 (�zxN�� 鑥��}�.���<���	]�f�I� ʈ� ZsL% (���8n� KC�?�
�S �-��A) �hw̪F[\��J��#�C��X�
�eH��jEi�h?k�1�
�2�`X��@��� ,��:��ZA��} ��a|~�� �D؉��&�!鹁qf���PB� :���?�p 0�W-
�;����>���L~�?���H��VO$�P6 �`(��	X������ ¿8B��$A� Y5�� �D�%��s� �-{��/?� �;��o]��w�K� �Z�n�o �����pWy������� |P+踠�� ~R���ò  ��'�]�! ���k��,  �V�P3� �"��\W�9 �#�wN/j� y�_�F+� O�V>ckL 6�aHQ1�;�� =ϋ)� Y�+H2�� ��Z���T85���Nq EY1�Z� ;RV�v�L�鶲p�[D3�=�@`����G?��2<W���� ��kj+�( 7d �S��T�o��1�Z���Ԑ�[h 6/U���4K��qE�[Z�n�	�(ב ����L�2 Z񤻁'ô?BJ �{��p.�� ���|� r#c��^'� ,�:P��<� �
�m�>�gzq 1��L�� ��Q	^馏 y[��~z� ��-{����	;�0���� !�� �� 'Q�>�Z\� dY���f�v ^O���R���� a���_� pL�]
w sx�&#�
 Zl|��n_3 ��'a��4�� iX��"J�� r�O͡�'w� < ���I$hx_ ������� ��+bT?񀤛_r�|��F �^��t�� ��E��� ��g֗MZ�) �[Q
���� �	sY��<�� �`[9��Y#������`�a�5 KE0���� �^s�B� "�P� Ÿ}'�$)� ��w�t�Ё	�@-]��dAD	X��u�}S��H U�����&I`� ���tC 2ƶ��S�� |D�0�� ��J�+- ��S�2�, ��iD.�r ������6 �W���PCt���y_���\~�f��� �V�ϱw�;鷎�r맖Ɓ�H7��y ��^��8;_����0"�z H��� �;�\]Z�� 7����W ҿ��$A�<�@
_!�Ӆ �ݡ�Q�� SZ]Bܲ 	Cӫ
��Z������ ��V�S�� xQX�J�� ������Hm$��1� ��%٥9K�{��(��` L[���i WE�߀o_ 
ѽX�H0A ,R�� Q	 �Y���_����Jx ���j�������`�d�i )���	� �ZT�|�
U(JR����3�Z@M2NǞ ���)���h|A y ��|�'�0�x��/裐@H� ��C�� �%�fL- q�_z`�C<XJcP=� ^��AF TY�+��� a@��sp� 1�)����� D��xt-� �1�Q+� �����v0s\��6@� %b`)�A[ 	z���]5�V:�h2) �x{'1�sS-X���+`�� ���b�1���[��Ӭ0�z �W!�H+�x� ����]�� ��o���Q�q���L S��3 �(݃$��� u0�Ca)� !�,n/�h?���Â���O
}� �ntL_� ����K��bP��֮ U։�>�! ��UZ�1 rX3�0�sb ՘����. t� �'hӁ}�� �M���(I��� �@d�� ���h�#� UKâ�\k ȇ��)� XY��� (2��T�Rv�`������m�pQ�d���G�@B tٷ��� ���VI h�`��%� vT��2� ~R� ��Z
��. ʿ�$�	�w|� (��܋h�.E3� +Ɲ�2 �T4P!�  V΋�U� ���1���\9 ����J� �	Rut.F ���Ҳ8$
������j�D�I ������Ÿ�q� �<��� elvL�%�� ��@�0�h-�i���z� ���9ǀ� ��[ �/�r ���y!%�� X�,��"<X ]�RB���� #�_W��X�\���&�(��� �7U[G�`X,)�> �������	O���� !� ���{��;_�@� �ڊ?��X A1	��n� ��ҫ�@� d���[ -j��P�#ʠ0oh/�q��Y�$�_�(��*�;w: ��$`�!3#���Z1�� � ^f�w� �:\9 1����x0� SB��t��� :�"
��X�����W�~'<��M�q e� �/%��Tw� xA��V$�� �O�������� H�gtZ«)Q� \�%��� ���f�q�����H t�� w����2��U��� F�� ���`�� ���� �W�qA	n� �^_Q��� ��
���0ٗ |^b��T�k y�F�7�܁�L+�^x���CR����4�z�b�<�S��Ӑ��Rp� �s%�����?E������:�� 8
[�-�+� 4�_�М�"�{��V���䠞 QS����m$*\� t��!T?I�N0��� )�hk[f���`��	�� E��'�- �U��щt�y��1 ���:�[0BW�y'dT ��\�K	�� <�th� �Z��K ��^ ��|����@�o�f��涠���{ %�'O���ix� q�-� I����^��d���5��f0sS~Iw`�v�����X� 08�'�|�B ��`�3�R>� ��
������Q���0�N��t��������J �(σ��� ,���O[� .�٢gs�b 꽐��� d��m�h���q
 H��[�� ��fh���'�TiC��8 �=��"w� BJY����l�z�ً`Ԁ��=��FG ڶl0��1�2������h &)Va�z :�~v�| 1�9ʝ�x��` �z]�_�U������ݞ����p9S�< �0O�B�� U�x/��X�0��  ��3� �V�&��� �ӹ�`e� R�����n?�W�Dݾ��i��v^����-ǲ�s ���`��A ��2 #�����Z�8�`�y��Wl��� �����R%���>@���>�h�7*퍱���'�9(
�Y�ہ�] 1�z��!�,Xm�-�� /�l���> ��h{f [2����8>X�"�`ѴƋ )YZ퐱_� �*ݘ'�M.�O R����Aw��n@�*�{ ���@XZ��`^P�be��t�v 	�x宋��m;P>�H`� ��hj��� ��/��� ����^p&����Y��$S(�@K ഇ+X��,L��ӳ� ��S`+q������� �4!����A��˝ܸRŠ�����#� \S���P/����@����-���M���~� @� ��!	���	1\� ZW��+�*[�� gd�3׹�� �0�S�����fHU- v���O��} �^Q��T�b��t��K�?`�P ��\v;�� r��_@*K ���QP�� �0��
�
Ż�� Ӏ0[�� Z��L_2R ����XV�a е �q�� ���N戤� 2�zW;�VPµ/�_P����@���R> L��J0Y ��6pח�i @�D�\��}����`L)(�� ��W��b&
!��C��� �3���%4^I��*�H%�\ 9��3�M ��c�!���uu �\�I:�"W >�%��A^t|?D↮��LdM��}������<��?hv_ ��쌍b>>�} 0�[^�u�l{��!�W8�ݼ�����:^
�<����ާ�����u�BPR ��z	`�� fT&')� 9 �靚 �/��1�� q�4$�|�7�N :�Q�?i����0x� �8��K^E �Rj�P#�@��F�$v� g��R0 �V; �O�� ���>��&��u:D1��H����� (�k���� :	u�j���5p�%��h��G ��@�<XB�$O��]�Q ����<!�� y��i��4>� r���s <���ǁ �9�U+�!� ��颲L�Hzt:��~��R�e*�
 -�	 w���S� �UV�Cuy���^ 4[��x "N�	�.��@UT<(� � 0�� �X��o�.*�4]�,
�@�J��#}L��P��R�= ��o@�� \h�p�]�b!�؀���Z�v� �;��(�[% 0�fZ�h�u'�#�銕 �5�_	��^JP�ښ/'� ���햢$[ �AZ3�{*\�� ��S>.E�Ā�p�W�?��	�1�㨸�v�vd\� �8������\�AT� � vG�O� �.A�4� 0Ə$�'W��h :������ 
��23�A�>4S�Z짡)� 5���K� �'�	D��: �.�WE�+X��~ ���� Q����8�. ��ڟ	�)J]�a����� #Y�0��!� 3ڋ�*2�(؄/K�a
� $�U�k� ���51�~�;(�hmqذ� �<k�yi�-����N����ߨ�� 挋����� ��(N��@=*@��� 1���b �	���*[�G��@��X��':oe �p���S� �W	�y�� �Jȑ��'�)�C �3���J 1D�� ��R���a V��v,fS���@����R�̀�*�� �Z��[� {�\��Ԑ_ �}2��6<� W�`�1X ��.�[JO� ���1�\ ��yK����RSQ*��J� d0�� �+&�YN� ځ�R�S Ǣ	��:`P'��ކ ���$�! �3�-�S�e}5" �^d� B�\_� �'�WV�� ��Ǿ�[� 7�1.L��9 u��PQ��xf WγIY,V1 ����J� AG:�&b���h�,PC��`�(O U
�N(�� n������ �+ޫ�P� h}r��J�{�o"<��̰PB��2�_�zmI' ^�%�E��*���\���d���_Rݞ.��H� 	!ɻ)N3� +��yֈ� ���� |5&��j�u ��	����w� �_{�r[��p ��T�Q�� ����o.�ݰ� }���<�l ��!/�S�V	 �A��t'�N,�_- �O����;Ũ�U�b:2w)L� \*"�Q�9 �s�nÉ+ �B���X0\����� v��
�� "ϩ8�R��4y�I %���{	��nh��FfP����E ���I\ ��!�)�[ �,��w1�� +�^�z��?��B�: �Ͻ	�x� �y��k�L ���'3U ��1	�]S;��sP�O��� '�@н|\��/�d7��:��[{ Ix�_��> ;u��N��ڶ���h*j�����f�嫆����`��� v�t��B������hP 6��"�{� I��q�\s �B{��%�� e,�5n���ub@�W+ U���(Z` �:����� B����#� ��2*Xd^� �� �H! E��>� ��d�]�+ ^�X�
�,\B� ��\}�@ Y0>����s �H�� �_�
g��{Q (�^ �P3� �-���G	H ��W0�T��O����N^���Xp啛��na3�-	ԟ. �0K�1��� �SB��6 Wd& 5���K*� \�����JّP��������p�Ž�� �2�=��� �@"�-( /*#��)a�|☺���`׬ԗ��'x�!��]N�h�\I��Q�;N�|btv��� �!��g� A����{ �%D�J��r��D]�, ܚ )똖�Е�1���Yd�V���� ��X�g7<B����	�~�Z0�h��p�� �E�C�V� ��[�Ċ�� 
���|�� ��r4l�S8 �)�A�V�,իv ��^�4KS���· ���=� ��<Ac\ ��p�� �� KW�`�"�X !��I+�4��@P���n\ k�h�+o q��`�U#�?���J ��йX bH���=r�� ��1W �����b'� �U���������!��/�.w ��cQ%~-?t��8D���.ƞ� ����2t@G��  �]L����� ��%[��� Y�&٬��� �G-j��\� ��u�yY� �Iͨ�� ��Z`㸕@ MR�7 W�� tX�랺� �̿�7��1�&0!u LU �����@�L* ���f�&��= ���y�� ^���l� X��Ѭ�:>���%C<��M j�`1�)� _[�P�Y	sE ٰB�q�� IÚ�U3� ����[Ը ���<� LN��+�� [R�=�.�_F��ͬ���ȗ��PD���4� $(x V� ^����ZH��w%,� T���4�#�����d�O����	�5���d o�c��U) ���ʿEu��0b"���6�� �g���dmp= 	ŇψØ� E���Z! 0�o�d� ����$a��H 2�B�� װ� @Q�i"�0�2F��@pZ h<^/�Dؠ���Pl��:�j�B���tО �C4��b�$>Y�(��� ���ɐ�K` ����4<�0)n3�	G@�o� �Ç�{w� �ap��� 
��P*��� .�i��?� , ��%�������K�{�� ��[B3�h pX��C�/a���m_Կe���k��8�p�� ��&2�n� ]`���� P�L�Q�8"m ���.5� �@S3��h_��NL| ��� �b�\�� �h-�� Ve�ݒE �^0�!r�|Z��)P]Ȱ=+��U�SԡY�_�� ��3�鐟��s����%	��/�$y }�&���ӣ�	��ܸ@�h�_�� ���K� X��k�1=��Z�( ����M2��~}�
9`�&�B,$�d� R�aQv�	h(@зн��^��!4`�W ����'~� �٭����P0�]~�`�
�3�ؤ�ʀ��$ �����/  �������=ED���)Z�G e�	wL1�>r#�K�P���Y[��B2��Ш{�  �Ka� L��+�1�Y��.���c	p�f g��k7I݂ j�n���< 9�J��>_��;#׬�@�1}�
�"�)������t� &p�h�Ց�y4(��� x�$����Q�Y�A�@Dy�n=�����Bc�s�nSV B�~:�/3[ dX�*M�� �Ҩ;��� viFՅ�� e����xc �W*Z�|�%�2N5 TY��) џ�qd�08��{��}Qk KX���-� � *ʟ�� ���w0� X�8�%�P<�������>2ɀ�^�'�\- ��#�V� ���H�T�p8�N \
�R��&[�`�MN ���zAq��� �+�s݀��ZR��$1��l4��_������i2sFxN���j�k�f� :�V���.Dq���ѷ��C#� LT2ω =� A�\� f�7VN� ��R��� W��j.���1�n������ PX�,Wy: a���%i �Knϴx� d1[��O�fs��U� ��d�	@H ��f-�(� �*�\ù�B�`����� �����3�@�ŏ@��N�i; #��X�� ����|
�C�S�_q(`�����1 U���*v� �|�ft��(�� PYN���� R�/Bv��	 �w���\+� .�eN���{`;��S������H�@&6�Iv~�A��(ȳ1{ p0�o8��q� �����^� [���Co�. _���0��� 1;�"�5�tj ��)�d{�N�(z� %[����U� ��=��)ľ	K%p +��( �3�`��R� wI���&ZY��k_db����H��%�ࣃ��{ K3��x�� L�(��� H���c�� �>�9@�S: ��?K5�Y ��q��T[F �7*<S�� WM�P�(\� �[�X^Z谦 UH.�l)o ��� � �B�U�� X�5�]��"Ӵ!��.2�>	�Zp�#��J-��LX��� �Q)������݀G�>h� t*��-�qΈ�?]{���^yBp���Y�ۀH?=�P.�n �ϷK�Bh �)|Z~��3 �����	�E�ѕ@;�5��q�����Y����}rvu R�XC�j� ��I�Fp�h.3�� �1;��'N�W�,��� ��O�n�� ���=
1 �#�]��z%I���7w<�1��p:#�W� +��K�1 �J��Ɔ�ˍ ���0 �T�K�
�<����� r*^Ӹ��В� ʗ%]�9D��:����� A@���\C� ���Xʙ� 
��=_(ȬcN�0�׸�.���^T�_�Y���� cB
Qf���8 E����:�����-�\�� �6��%Ŀ�=�d���{B �XiU�_"�ꊪ����sG��`��*
����w�7C��:�my�`��!�[�� �R��S�� � �h���\� �n#��я Q*���λJ&W+	ˎ�n�6�Ї�� f�3�>2 ��dKBrZ	 ��/^�� ����N��Y_����� 9yP���
��]_�Q"?�}���P�ݢ ���5qj� ��D�G  �CW��h}kN�r����zb�Wg RS���8 �ǃ��;&	� �!˲6r' �
���T��XT 5�!��t�] '-�V�+a�� ��O ZR��}3t�	,U�0��.�� �6!f�L��� 1�Y��<y!
�� ��J[� ���R����n/�;��x� 9z}�\RP�ؖ : ��s| ��t�YK� F�un ^�:�[ �HZ��g����������� P�=�#)I���j��ڒ�X���_�UOH�ԉ=
 ���IK /�ET%� �|�+��`���03 �d��t(pݾ (e�W� F^P'�X l_����� �WF� �	%vP0��(r���D �$��@� P#�/�8�� .̹6'��K to�fI����ɕէ� ��	��%�o�6 W�)� (̿Q�%<B��-c�y�pO ��
�����pa!��<���I�Ř�	��T����a ۸� O�^ ���|��T� @�`�zU2&���bL�{�%�� �A���h �a�_\�� S����>� ȗ��Z%� ~�O��X��� R��ؔ�s& $Ah{co!��/�� �} [���#j qBO��Q��S������
�3%�셓~@����t�)`��� nh�̖`w3W׵$#�|Jk���@�@?,K� �&�WJ�s� �;�|.
�� ��"��}�=E&?���.F��6ZP��*����隌 4�q؝��s> �H�	h&5�� R��Y������Z����AR ñX<7� �O�?PpL �	[�R�S ]K����o������� Ec	��]x 4�|l���btX�C �PQ7Y�� �)(k��'X�� ���?X� ��s�}�� 8B�tL� ��n�{ ����whT	~� p�d� �<�Ѱ�&�m�.W!�z���c����~_� �)��� K�����Q��] W�%L ��Ճ���<�(!�ˀO� �P�&�` �U��R'�� �I�* ]$Sǁ&�� @�Z��'#� �irw�\�h�^J� �/�}�-2�öy� ��1���3�� <�zt�%YJA�`��
�&p`���Y�h�~X@2�7��K���	��0]J&` �i���C(� �|Zz]�� y��r��K ��o��T�M&���.������]����`l�� D�S �b�|�L dI�Εw�� ����3K� �.�}��� `�Q)J��� ��u�0�� ���@��� ��Zu�G�� +�r��@���o YR��9� [=E�0K� 	3�_YI����� c��ʈ��
���"�Ļ8�d*�3��-Z+ Y�P��� s'	ѽh �q��`�� �tN��7� ����%� ��1n�i ���	 �`M�l@;BHv# h"$g	�- �Ўyd�� %,{0«K ˙��U�ل 5H3-w} ����dĊ 0������ ��!£�K8 �,F�p%� �
1���`y� 	P����B� �o��WX�1 3?�h; ����A\i�mg����ԋ e��Eֱ  �W諔�� �b.�qO� ��k���,���� @[�o�v79V>M������ ������y^S鋺@���CL��9�6^_�N1�{� �(�h��W Z�o��be �!�@���� RC����{ ށ�|M�� ~[ݹ)�� ������"��!1�?���Zn�=C k~MV�\ �[A6� K���.f�  d�-��"�% ī�Ѻ	� }=��rt���S�3�� � �'����&U���S���^ ���c�2 Ǣ�J�8� ��0��@�!�I�p׽rY 
��k�� �i0��w��"��@Ӝ�� �BTt]� ��&��d����1��ْD��50X
 ��8�b ��/���� ����I S�\�� ����� �� /�S�X_U� ��'���	 �L�!�C ��~�J��� ��4W�� ��X�(����cp��V> *�%1�ט��'�\���0/ �\���% ����-'�K V�p�8 GW��s�^���)z ڥp+[?1�����E�	� �j��\(�� �V���� �F��R^+ PV�;�B�� D��yZ��Rf�0��`! �v��ؾ��Ca�Cf?��_��= ��5����#��%]�^� �U�Ev�0M �i�����K ��eZѯ �j�g���v�,��~�t�*���#�_2����P X����چ������/�2 �ef�zh\ K��(߿�+^�9-�M3� )�1�C ���{�,��@��P�� ��c��C��Y�dpX-)���� ��х�\ 4	H2���-]�tO��Ζ@OI(� ']���}N���+@�O:� Œ �~�m�� ����{�k���N-��A��K w_�Qė� l1ճ}*��@���RS�� �E�Jt���< �ma�k���� ��*j�� bAH�/5�����8�I�"J ��i���z���sg����� pe�}� Ҏ��!��;����DZ��A*H�	�0�!� � �C��P�|kJ��� |���'�X% ���v�+� �BU��	_��3�ԗ4 �=Z0 ,�%i�z3 �1� !��� ���[��	 D���m��qH�� �)����SY[����
+�l�
{���D��������3�.�K� �M��	���0�Z����$� ��?�gx� z��!AZu/�qY+G�� d�kB'^X� iQ�<O	R<�"�D62��l��[�=��F��N1��< A�@hX?� B(CW�x�u ��J)�M�i ���S�1� o�)2�tD �$��?�	0 �h����) P��Tu�;O[���/��4�$ �h	��^q�~���`��闺�Z����_� M����
���G;���� 9O�%y� ���~s�^]䄿 �4Q�� 	��)V�i��XХ *0�Y���K�&�� ����!� ��;�ԅ�И& G4��p�^ �1Ѵ��X;%� l����� ]"ڇ�1 Pu�/>�^��̸� I���6� Нh*�gr ��oA��� ��܂�� u5�	�� ���쵁�+��0�]ʨ�	� ��
Y�h� (���w#C ��\���� �ixR*bn�	՘��LK�O�)]za~���V u0pq������Ƌ�	 "��`/� ���t���� )�S	W�hf (����� $G��P� ��R ����(܀��{����}|���J/�O�+�{��Ɋ�4L`Kt�� V��q0�� /P��X�� 5���_+� ����z�3��a�|�P�_ N���Xn�;HU /��e!�� t�S���1 z����Ł=yBpu�'ґ�1 *	1�`��w &���3Z�n�LA. 8� �]�����m�:����-e<����	x���@s��[��zs��Y �9kf�� <B��`�
� ?hX���=�� ��ހ 3J%�P�k�������,���{(�� N���V�/��ȡQH0v�@��\f� a��m�3z�( �����q� *��ѻ 	 �1��T� �`��Z( ��1�U�Hbi V�Zv�iM���h�&0�9��}����� S��Yݧ �h�[� �1�W�^�� vs�}�a��UT]�V�v+� Q��b,��S����G� �?]d�i�� �N[�Ҙ��=����ZS��Ș �gJ�A| ���� �G�^��d )�������5@�Z��9p�V 3��U'}�8 �-��غn� [���c,�
	5}� D�GS��������J��� z�QS�4 ;���hZѤ��K@��+��y�Q"C��7�^�!�T��Xf�- 1��_�	��0��ĥb�B�uq� ��kGT ����K�� �
Z �.7��L�\� � (g�)�	 �{/�o�� 1�)+�; �_�|o�^:�(k���uX� s&�,|� (���}{� eƮC[^� @U$��I(�i���}b�Ҡ@���r�1�HWS0 C�Z�A��������u��y �*�b{%#� �L
�(����`��/� ��wl28�� @�-�N=[ \ ��e��*�H#�م����Y��须� ^� ���0�|�/=�s�[���`~)Y{�	���>� ��� _��EtL�wN8�@z�w�
X� �c�:����&����ӭ���ez���ŧ& �ܿ5� 웴D߰� ���%�`� �]k�~ ���7�[ `����������R^e� ��W�D 2 ��*���k���ց��}�) ���D1�Ļ6:���`����	 �e��>�1\h����*��kt�s����A�C���i�Ҽ���, f?1X�{��� ��h$�Tɒ3ث�P����Q�& Kxb������FXo��H�ȭP �	>���J������ ��t��������VU\x�JF�� T���b:����X�7
L2B�,/C�Z=�!�����J�{�a&�0��y� ���Ӏ���z@�21
}\�o��0���.���Xн	 ����Y;�= ?���B�� 6��z9a*�:!��PFğB��s� ��5�/ �
�ZX� �$9���0���!�R� |�%�`\� #�D;��@ �q"�(j�� 
�P?�X ��_�2݃� ��E�0Æ��ɦ\ �W['h V�!o��J;uB?Y�А Q*��I �]N�� �Z�8�匼� 4hQ7�*�p ��.sN�1 H3�;�K�� R|J<��D �1u�M� ��]�e"�� ��E��M4' dy���  ����Κ��)k�^�fP�_�����h�0b� 6YZN��/ %��	_1���}���<K�����E͎.�� �T�� ���� J�?S*͝ p�NʯhY� .�nK�d4 O��B�U�1��-󚀨�]� �h���t[�pi CK)Ё�Ͻ H,��IB� λ�<Ґ|>h����d� ��o��(
 ��P�8�� N��C�`��	�A0r1 �a#/� �R
��_� uW��F�0� ��5��>���vKP���?(Ov	w|ȫ��0]�: �H��n
� ����t \ѧ��!�a �Z� ��) �i+����:�{�ї=�� �^( ��� ݋7�� �`FSP� ��Ky����� �/AB�bͣ;*L ,ʬZ�?������.hJ k�?�I�� �K�'.	���!�<U ���k +��?|�'�\ �h��߭/N �[�븺  O��0#�X.�X9t�M��nԒ�.� ���%� Xj�`;�6^ �ߒ��?��� �L0���q 2��
�	6hrS�D���xu �$Vχ�o �/�g�i� ޱ��VmX�� .1j/~���O;n����N������\v���H �#�,駚� h!�a � 0j��46� �B��d-Z)J�\* ������ �+����	 �|�eW� �La-l"7� N�%X��10�������U��g{��5�f<��� =1m�8j��� 0W��_�u- �EP(N�������S���� �O��# �J�XB�ɵ� �6"� @V}����� '��
��>����,�@�<�ՀDv��iP�۝f�,0���y��&B+� d�^���. =�!�f/������� ��Z�z}&����R�~n�v X�9����� U-�8�] �!L(�e_��� @VS�:�� ���u!���#pb�YaJ�����i@*�	��ǀ��"� )�ЇG�:J* �Q%"��i ��G�5Y� -��<�� d� ,�\�J��[ ƹ���I]�H�;�f	�鵗G�>����\#� &V��� v�����='O� ���YĻ [X�`پ\ �$'��b3� ��u#�	���=�  �PW&b\ $<N
�Z% ���_xtiM Wy(�jb� �J
�	)�T�c]ۊ���� Q��P-��r wbl�h\ �NT%0� (�� ��,w$�B��ц�ZM���Y�<�~\�y.�4 �:�w�3 �-��g!� XLAr;�($��X w�S��	�2�� _�����pd I��{0�%���l�V����T�Q �L���8�] �)ĺ�W-	`��B��1^+�!h`^$ F��߽��8`1oJ�N�~D� l�� e�>��M0��0�� -�(�^�� �;fZ�R�b�@��X �	�)��� }��>,�|4���`q��O���X� e�$�I�3x�� K��U�H N\�7���L�0 ���0�ȿ �Pҙ[�Xh �4"�UH� �ὸ?��-{} ���w��P|V�Dϵ @��˞�X� B��:�����~��q©*�  ����k�n�.2�'~�ǐ��}O{� �h�B��%Nf�����RU �IX�o�?Z �s �h]��#}���ф�,�J��� 9Ľ%1 �Xv4�!t�M��g�X�� _����*�W[� � Ѹ_� DfZٮ"Ҹ8[�� Pimx9.�����ݸk�� ���EK���j	��-��� ���� ���J���|���-�pT��C��^��5�=�� �Ob�\��@�� �	R3�� [�� �$� ��]H��t�.BG�� �!���O�`�f�p[@�Vh�:]� ���� ����_:� ����H\?* �X��TvO +a���
d� 1���ޠ� Y	��)� G7V%��Q XYSH��� q;	1؇� ���<J׮� �/�!"�1� ���ʵ��	(�z�2\�B� ��H���[LZ$ ���lO�5G����4`�h� ��8+��֕v��BB{h� �U��09��H��tp�ַ� �J�������P�p���j��<����M� �q%�����j_ҏ8�`����}H$�>� a� /��[��L���]G �_���e�� �DP���B�ށ�cH��` ��L�&#� ��Z^0(�@ Y!eɮ�V ��{��F��y�6��U�� ����=��h���p�s�����Q`�����ǘ�����1��Y?��}02"Ͻ�ae�m� ���(�Y�� �����5/[���,�#Oۢ������5� ����0_ L���U(� ��)|�
�ۨh�#Z����N��t�?��@>3Xؙ& }��
��\�x	_�����p ��W��vV<`iJ�"������w�TK�S� c��8j �.:i%���*���2�D�7E] ��X��
'� �x�4?Ȉ� �|��0lA] ��P��;��?(���y��� ���b;� ��U�"oH
�c���'� ?s�R��Qն���\*:�PÞ?�� ��r/ � ��_^�
�@��0�r�1�@�� �(���� �̶�A9R ��T��/�� DI��36 �����X �fSP`Q�����`ޘZ ��<�M��"��! �Ʊ�Xn�d����c�y� �@���9	
�Ī����B�9�A�X?���,ӭap͢�0��ݚ��w�' &T���o| ����	S� �q���١����P��	Q!�}y��61� ���^C��-K��" F� �VT^�K�a83 dq0<� ZO`�h�z� S�ӽ6Yx  ��7<C ;�U��= ������ @��CNqO� BFR�<`g� :1Y��Q‸	 �8���;Ġ�����0�J��O	 �@(�� t�2�'PNl�1�`���?�8�@�	p\ ��6Z��[ �"�_�`nj ��>�O�7��ű�p(�uD~�ңP+�*	� R��U��- ����;:�� z�D�xr��j�;��7�͊�[�1M�t@��k�{����� ��"�5)��N��iJ� ���BD�p�N���� ,��)�e` ��Y���o��hqM�y&- 	s�U\@ J*_ɴ��" �<X
p:�^q�=5�������a�\�+@�dNŗ��	y:�ͨ^�K ��w&H�\��zyF
�^SJ���@gȇ���Al �CZ�
 0,k��S� i���=;�Q e5�9�uj�uP�p@u �����Xt !"�V��BpG� �1q�R�W�r
�E������.!����]� �yS�� �����q`�P�,�� ����e��T ���-��� ��nN�#��gd�����:��O�����XV���T���F� {�jZ��qR�� ����!��f��� ��W:�h��u�`�>~���!��]�� �w�̸+��u'��tB Y(��� /D��:�%V��	\ ����=�tY �4�������7MS�� n�h.kw� J`$B������HTO:A��p\>�b9����+�K �����S��MA5>��� ��%��X2N�)aB�} ��*��X� H�G��� �dP�ݦ$ �*�lՕޏXB� �b��um ��(
_�&�� ��gZ�% =����J� �ArR��>�.AW�������U0 x�ß��W�l�cNv��"n䯒��X��a0��E�e���,�P�v� ;)��*��� �p�Ş�	{� m����HQА'ؠZ� :�g��h ��cK��V u���HI�O ��_�' G�\(�|z�T? e��Q�܀�@��!�  �XR�G j-
���ӉWE� �1�� 9�[R�*> �\�ret�B�T�U��� �1�ɥ`- |K��aU� �O��8�����k vΈ�51�3 �HL[ϼa�!� ��N/�7 �P�X'��<� ʹv��N݈�1�p; Hˋ�'m 0Ψ��Z�4@�w�;}Q !���=�� ���nT �-�'��-Z$`�h ����B,v� ����(� 	[����
Z1� �֌&�?�Ā!����^ ����n�����o �
֣�y �Z����	0# ��_X� 1��l���  :�JR�V�X)���� � /��?��0:��G0�� H����4u ғ��݌0 ���6� >�)�߇�}�L�� ;blE��o �ZH-&2h�/�"F�^�	�Uf �u���r�a�'�����[� �9�q	�j� ������vW �����h�PR���MܵY�>#� ���_V9(�1D�S��	�0W�p����*���rֲ� '��P��%�m��3�\�y�K��R��<�Ĉ�[U��R���A�Z~�ɖ�u7<�R Px������P���:$�����B`0m�� �)�_�= Y��U	�� �`Lوp� �3�Y[�� ��C/y�sK �%�h]>�b ��\Z}	��� W��͆�u{=� '_�]D ܼ��Z��U��%�up`�8n� )�X�'/ A�볕@r�t5 ���C��Y���I� �! -�uc��| �}�S�N0G���� gPL�=K��  #|�`��?:�
�
���Xq ��W8 �>S��(� V��)��� �	�^��"`%�_ ���x2�-�w"��Y��p+ <)�dOĕ8-� Q"ع�k~ ���2 �'�n��� ��.:Z� s�򒱶� ��y�"$, �)�YS�� ���T�>�f� ��t%�� ��)��2 �U�-�Y(� XVQ�:� z^����mB>e ���Pl�Q � �f	�(��x_�P��Y L ����.� g�9hI�c� ���b@3�KS�>n������ L�wA��\wh ����}jO� �׎�P��[ �l��0?� ���J�Ik<�� в/W@؁ 5�2㥍����E)�����?t>p���` 1lEo�� wO�7����� �	$r�1v�th.� 	 {^��\>` ����&�vU�,�J� y ��P����k^�z� ��*X:���mfZ
�B��0"�9� ����.���Yi��U�0'#����Y�LD�` ��M��� v�1�, ~Ah���;\��+�U�6v@$<�y� H�� �[J'@�AOE��~�g@���]=�&�&� Y�pA� D~�E*�0%���\��R� �I��г[Z ��\�&(�� HR�@�2�\-��F������1L�"3ڀ��7� ����%�� �F��� ����H?� ]O{��� ��(���J �=.�^���k�>�@X����nY��$`�m�@�1�� V�ւف� �Y�W�� �0��'���$�nl ���Ơ:&��H	x� A�6(r^ �-iFa�X�s� �h/�yx� �.+2�E�����]��=� �_��jQ~ �k�`	�-�GE
.��^?�KL���0]6
P�����(�1�a�l��"�A��>	k [!u3 |�
ʽY" ��X�&�n�  �LSd-�}%��V����K�/邏 ��p��5Y*.;�M �y��w �F��^8�R� T 5C��xU�`)as� z*�p�& WQ���5� ������ưZ �}-x(h�K��I"~Ȋu� �J�(��8�G"��cu	��|�v �rբ��y�2#!�"��H���ѱ璨 W�K�0T_�ɐ-��@:{�N��3�m��� S�1Ҳ50�{. q�z��J�� !�v1�c��+���`�X��  ���'��pszg��D�Z;� 9r5�+��2#����Đ _�uW5�� a:b�Un sJzш6�$$>�Y �|e�)Y[���z�L�_� �?�� ƨ�(��� �W0u�$�z�Z�[���% (��/���\�q�A�Xu:�`��g�@�ո&ArE��{��M��s� �P�X���p>�޺F���
Q� ��?���Ȇ�1����� ��ڀ�v	f P�CXp���-G�����
 �6���L� �2�`�.P� ?�J��L��,s��W��Gܕ8 �;w�K.S�MEa��H@�υ��K@+�J{�XR� ����	� �p�w� "���*�� 01���[q >𷻿�f?�_,@m
� V(�楘r]h"�����eX �J�ob���H'ch��6@N �[Ϩ�(I�i�"7�;A߀�j�K��]� �D	�� ��,Jy�HKA*�r��u�X� ']�	o� �.@l�:���ݺ8� �����{Q��8W@O�/l^�}�hQLA����M�# �_tb�� ���>,'� ������� M0^�J�� ��X�`Դ� h%�}Qb< v5���3~�Rձ.\ >��u�� 4��HNa�a�&�W?��'�V��� ��Q�L�� ���՞To �ńe�(�����2/����!��_ ��M�bh�=]�}B��@�Fi% /����q�2 ��W�+ ����:.��v$9� ]TCP�N �
�����x�c�H�_ ��^�vn'8 ��X���� �|0�\
� P���S� �yc��\ �R"�i1���`3
��?���+��%�q������1Y�B0nx������,��  ��vW� U���B� xu�� �`'�oe���<���c��� ��ZQ�|�ɢ�^���h�/� �K���� H뀈;_ T���h�� ݉��3'� �B;�S�4x �� ^2_���/a������� l�+�0 �#�[���� �OӊXEH��l���$R _b�Չ<w �� �^�,� `�L���h $�Y�b��~x/ �
	������M�J������ ��4�N��[0n�`+'�C(��#�{�}x�&�IS���]� �{Q�q����U	`߷��)߄����� �dS��� w �v���|ł��w;s�h.X���<O P~^�9p��2�;y*�B�%�v���< W�hp� ���0)�_� ���n\� �1���{��?����IL�	�Є�=��/�:�0,:��93Q����V �������� �|��x�� H]lQ�k� �&�iv�(� ��-�@����{�2ʀ�dO�,�9�X��1L�� ��I@с��T��5Rn-".�p����� e/qĀW�  ~P�b�'�w�#I����. [��WYnA�� t�X��8 ��0�PV�i��	�Z���� �Ih=�8y+8³���u"�3��$-* ���� ��d��\��02]!���I�w-�i�	��	� ��׆� �14v耼�㋒��0gx J��_�a{ 5;d���� �PNϳ�	 �]���! nE)���\W������� �	������vI /p9f0� _�X�-Y�
$�+ ��ԋb �T�	(�! [3׻<��� ~���o�n~� �K_L��0X� �\yh� -�۾�)��a���]g �칀TJf�4{ �����X�q�q����[����h^* 1���D ����ƹ4�* z� ?��J�<��ԟГ 	�VZ��C� �%[P��da �&\2ᄋ�߻�& �!W�g������]�/ V=�f�7�����r!�] ��^ �0�˦�u8��Hp +�ZbY.Dp� �/X�|IE�� �P'1�n �3r����	>b�uѬ��"� �2��OS� �PU�g�� 1.� �X[\�k s����u� ��d9�
� "�CHv1K�� ��� ��0�$�E�`� ���K>yY�<���@���W�a½n*��:,�ʐ��ZUS3 ���4�XH� �9��w� ����al}��= ����~�% oR�A�T��.��_�h��w ����o jz���l�^ Z*�����Q�0��XIN �!��ﱕX��\*�0X�� ��W���� F� E�Zy ���	� ��� �Z# �鎬�n� ����p��y� �~��0s��a�p����x�[�8�r�- (�����Y ��{��A�� ��䳗X� ��[��P���n����b Z�3J' ^�T��� ��U=��c?�Zⸯ���D �L����0T���$�]�ҽ  �!1r�H?>���aU�B�� 7T8��3sż�iX��nko��b�*�պ ܟ'�� ��N��	� ��
��.ɂ?�M��)�� F	�3�RG�� ���̓_�߰���'� R>�o�)��`5�� 2hL�-�z���`��# �`,�E�� f���.*�y8F�L��N� ������S� 0�b*�V� 	Q�c�x� t0��
� �z��f�Ï�e	�\��(� 3�-���PZXI�����d&��j ��=������ �^EU �̫2j��� /,�	��)Dx3� Ӳ��ARQ��0\P�= ;�9�5[�7 b�Z`�n������ :e�=�η��X�R{C� ��0���NX��R�2} �V��!K ͯ�v�/hg[Ѱ.��(�� ���R�[p Ơפ��$ ��(ۉ�{� ���t�9��󗵁���ە�� �DW�.�P� z�Y��� U��8��D� X�z �J !ʻ��쾄 )���������A�����[�� 7/ox��b �~���Ȭ� %A-�q�� ǣ�_DK/�� E ��* �����^� $b��	� \Q����=��$����<2� ]��0@U" ��_�$� �}Z�0J��;�x_�)z��8ՊԶ�8�t��cFj�m1�� ")��~8���������� ���V� �T�,�� �=�)^I� ��$����]�� �>[��% !���8, �1�'��"I ���6�7�>�����������V�$���C��hJU��� �W_�+�� �=\�� 
��4L�.#%� t�?)0 QoH��� }�����/f
Y����à�M��_�`z&�I;�6Y� ���+��J �I�x�� �F2G�z�9*���xM�� y
ضXVE ӾAw�D�% ,BΚO"�\ a;W1@<i 0׫+��� �_"��N�u6�|g`���� ��I]�{!m���@���T���}� ���)��y"������4� 
�=������N����(��' Tt�A�/
:�9a�J�i�	V�ܤ���^�� H�5�Lԇ��� �2Ҙiq�� +��o�rS�� c��e����0ܷ����wY�� ���TD
Ɯ�e0Ϋ����@d�1;>���o�[h]< �u.L��� ��������_*�� ���$�� T��"�3Ð /	�\���� Y�Z�� T!8�yP��\��;��% )���|��}��B�Q�F p�)�N^� >����}��hP�')�d� ݺ �V��� &	۰��n:� ����8 ����x�Ƞs+�.�A��ׁ��@��}( fu���� �.y2� ە��e�	xD%�Lԥp���Y�����ڹ,1�
 �{�(� '�����3� \��,���H[��-��]0�Wq!9��2ca� >��ZLSg U��-�`ٓ 
��@ ƹ�b�Y;  �3�}�r �9�4fL�z�`>��p� O]��_��a���>#ʴ�Ҁ �]ӗT^�K2��B\:� �p1��>U�ν��B���겂`�G?��@[Q����z�ZYȄ g"ʺd)�S�r$�Y\ �Oy�E0� 	@ ���� _lQ�ʝy�d�A@��&4b v�V}��9�0 �����_ ^����y�;����7 S6U.�� ��z>Z�9����ܜ2 Y�� �[t!����Q�0��e�>�hp��*�	8;�z�L���  ����� �5
��U �P�|�[��T�/�U\='� Q�%©ynD6̰
�R���%w��ʽ:pYIp�כ�@
�'��_�0�������`�]T` ��Jҫ�6��ԉb���DV� NYk ���~�Kp�/6�$	 ?%��]� P��'hv�Sz�<�-�0�}��>� �IW	�<�ƝY������ 8Fz"|���R��2?�s� �X�!�^0���'� �DT���B sV��v���]|����h�TO	 Ҭ%�� Y����a~ ���Z��p, !�A+�hq�/}� �0�~�3�r'V ����4��e� ��	���]S�7٭`X Z(�N������{� �-�enR��� ��K���� {�Z���� ����� ����
3 ��@[�� {W�\VZp� �!�_��w� �@Y�Ľ��)0/1�6ʱ +�X�t� �H�5J��o ���8/RdV1� 	�`K�����_n� bc����2i \��f(�ٹ OrE���� �ƇF��u�1��E���K�C�"̀}F��� h$iZlg��`�XI�:����	��� ��t܄ ��� � �0!��_�� �����Q�  �h��R%T Z��X���a2(��/�F ܉�ݸ�bs �I'ghU&� ��D�{?�~ ��-@�U�+ >��6(�� �, �	��\�Y .�X7`�^\� w�W���r� !�]�{I� ������.v;9�ŀST��Q=+�,k�Fw<�%	�V9 �_�� �ą�(� 	;�}ѩ�<Q�ֹqa؀���a�`�*� �QV��9��x��P��U� �[��!��8�� ���_M_֬� ��O���P 
K��7���xp�Xӯ R*�� ���"�	h'=�
�`�5��:��:w ���`=<1��"� ���2�_��C��'��� �l�	����e@�jJU[� .�S����8����W�& N���X����ÃUT+�݀��Q ��\��?Uf8�A�:5���������ePJ��mV@$�\��$!RA�^�I4/ ��Ĉ��X1��d|�/ ��������*� A7�żh�'a��o��7 ���8Z� PnKYj� ���y��&V�3@kr0���'M������5 8 ��)7�� ѳ{]A�
� *�8	�� �Uk!���� B]�hM�f��Z "�P9���� /'}�֞p�¿@����ZH|]��c
n� ����B�� ^��:�&w �N���/ܐ��5+�� F0�`�k��� 	��CP� 1��ŮJQ S�A��T ͐'P^/�&�� �Ζ!ý b`�g�s�
 ���i��Y� ��õQs,�{��&D ��e�Z��H�Q������ 5����q ���xa"�n ���\�3 ʋ*(�ď� ��ZY:h�J ɻ -��� �L�^���q�k �J�B��Ä��@���� ��A�!�� ��8�x��L�PA�� �h;���� Zq��_p^��)����^J�- ��jDW�O� �	� �!@� �>ѱ㌊>��$UH)H��bA�G��� D�wȸ�� ��h�U� E�d[n�a_ �:c(�HwΞaR��?p�?.s���Q�'�	 ��Á%f�� {�y�k� �hl� t��YQ	���Z ^��`]*�)������ �8�WS	��9�_��^� ��i��7N�B�@ȧ� ��~���%�vFn� ap�h7���V��N�! u���n0�;)� � �W�� ��|/%���H���Ʒ h�IW~O��X@G.�KB�w"U���� ���r8�� ���	�N U��=)�� ]`�,*TiY^� ��B9"���1}�I�Qu� �F|�D��"�Sf�9�����H��1��4�yh�`̡@rBV���@4�P�����Ȕ� /}	��D{��  �s�)ժ�T�}@%ȹ�m	�c/0 #v��_� 5��s�>��^@�x���>� H�,(�X�^��0�cx� I_��ՠS�[g���Sb� �"�P-�� 5[0�^��XI�LՊ�໗Sv,�2��̶%�� ���@�R� 'q��>��&���������?� ��i�<3E����zH[�&�"
���\J٢�2~`,�|�ݓ�%*�h�-Ma�ô����;�� ���I>��;�[ ��?�-1 y<��ԯ&	��X��;֟
� ��S��r��~�RP~ �O$���;Ѕ�	(՘ 0�_���K[
�b�����u�n� ��/؈�K!�A$�� 0IQ� �o�㖄k�T��FA��`> @CY�U4��x R�0�� ��:P�� �H��J�B�e�F��W����� `� {[$�����$�a�� ��/	���� �j-l�Q�H'� w�Zu�v+ ���R���8�� (��@�c	R �<u���;@H�� !��Y�o}`bx���� kg���Å ��S�T�L opHC�K� <�����0�%�	C�΂_�mJL]R��ڢ�h���+�B�%Ay���> ���@��I ��?)5�Q� �sK\3��+�D�y��M�z A���+� !�͢���ؖ�B���n ӦZ�� w�y�KIh� |AxT���/ �eٮ�=G �"��r6���p[:�� ���w|%\��X��؉��o(n]��)�S{�"'a��/��M���m�+���Q{_���d�$0�� �ys���m@^��]C���1
 �Z��N i�D!��;�p�#��߀�����7��=���� U|^�����q� ��	Wf߫' V�
�"�� �.	��U� �-�p�LC����.^�Qz�
F�B� é��V� ��+[`�����p �OԐ<ɸ G��V)����0�1��ҫ �keA�h�P�d��?�+� �v&�� �I�"�(�y~�� -A�d��j ��р�e\U	�V��c� �_~����� ��/" 3.��8�0��#� �~ ����Z ���R_��� ���4�\" &��KWM# O�=a1p�9�-�R$ ����( �.����� �b�x"�O�P%��J��� ����U��%��݃� f�$��� 	�Xh�)��
"}ƃ���؋����bQhF�w`��� �S��C�� ��� �E��k�X�� S�;G����Ch�r���RK��݁���Q2� �!��;$���>"� ����� �I�O�S�5����#%��v/ �����S( ��UDK>� �|��� �P�O@N�>�%pH-��=�2B$�j?�ZX_[�a `1�t�{Nnؓ'��J��� ���Y�]Vߗ���V����� 
�%�*C~ ��!Ѐ2 �� �s��U �t~��� ����v�� Ir�Z�m����`{ ��]0Y�-2xe���`���d�� ,�h�M� +�Rź< H��ue% �0��F� �Ԣ:��� f1T��	lt �?��3G� ]ʨf�� g-}(� ���S�p] ވ�R*� P0���3`� F1w$Nc� �g�]s� �H=�@� �*W�'�U� �mN���!/$J ��X �V �A�{h6 *���sR� ������ �0�GJ��OqV����h �W��K�2 E]TS�M ��W_�;B��*p�"��G��� z���~�L[&,�=o`�(uNV��Z ��ck��-h"�`�2�V؆z����Xt&� ���W�����E��>�ؠ�<���i�B`�� �!�NXљ�&��s)�*�ZQ�?6�z ���3�!� y�8�-w������X*��v/�� ��fR=����� m)�2�Z�-� ����Ⱥ�Q!N��W ����tP��n�~��m�(L-�>�ѐ���� j_�bN�q ����l��A�(��\. ���am�U* �#�^�Fh� �w�`�م �3��8/�H��0�Ƅ��?Z �j@��U� �
)Bp� �%�X��߳$H�V�K��"U� ��1��xn �*�W� �K�.�z ��H��[)I �U`!� Z	º(�߀�[�HMO.���Т�tx�Xٶ�YVю�D, �fU~��\tPL��I/kc��������% RY�A/�5@ ��m!� ���R��DW�,w lk��ƞ Ch��F{I �H���Yv<�� 	���:� �.����f�'�!~�X�� �� ��[�� i3T~;I�( G��+�Z� ���,�W D�/�^�'�9)N��� �$�����ʹ�� h�u	��Cw���� -���xY .�$��I����^T1�	 �h� ����Q�/�K�i0 &�T8�a��M���v 	Ue�b# �_��'5�� �0�8���\|e�����o�� 4��1��: �Y'\�
����������P�!R	�D���� ���E���) �&h����b� �*Z�ї��has��� <���i����ͽ0 ������� 6t�&z� 	3�~��
� �]���.���?�����3 ��*���ٗX�,1�_H`u�� �3��@W .%����ayN o{DҒh_`C������,�K�D�+���[�V T:	�`�d�x�`ģ/ ��Ơ�� ��E�Fg }�SՈf���u� 2�[  ��l��6� ���ߋN� 4��6�K��: ����<S� �ށή�v� �j���� �;R��#Ǣ�@��*<ρLjt �^o�ׇ ����h}"� �Q�-�U\dq� ������4(��p! 6f)�\�� $	WYr� ݈�ˉvR�?�	 �d1%���� h<���)� �-Z���# /�,��?� u��i��e 8�f!��� aA=j��g�?��������6"�=� ��� � ;��?���V cb(����E �����$�� ����A0-���H �� 	�^��_ayo�}qx ���3t ���	���"���@u��
� �*'�:� �A^n@�K�_ ��dP�$� ���)�l/�9XR� �+S�c`<�h�R�~����~]-��)'��ːf jZ�������u�M_� �]�h�f�YCk���`�� �	�E���h ��}/&�D�@��! ���Z�� (6�шI���A'�>��T�G��h�� d<=�1��� �W�-c��L^	�}�Uy� Pk�Π�� ]M
�`SAe ���=+�� �0��)t�	k�˱��Jί ����_G�!� �n*�S^=����4�DF �.I�C�o�	�Q�p]�� q=h��`��x� �+ \�*�� �yH�k 5��K�Y��Z�ب  Q��!�h� X�a�� b��V��ý c|��w�x �0[���Pǀ��lE�w�z
�%�����x�� �J��G��1 �p��`R� �ѿ�|�٤������ $- �?�/����q��� �
7e�� %��� �����z�` �\h~R� �|��0:���,nh{М���!�8� 0�J���1 �˶�Y( ���2޺`Z��t�dN_�˴`w�=��HsE>#�26�U�R�ho¢� ��[���Y|��/��ֺh���pظ8�[��b� {�ۡh(;B ǑW����i`^�x�q��T��-��u�� ��8^�9 �����'3V~�pt �$,����~7y��Qb"�LCV���_�@`�#! ��1�K�� ���r]٫�Y���/�� �� �G��hA �1M�@+�� �[��"Z� ��;�%� Y����(S ��P�3�t T��lX�� �L�?���(1����/�Pj�� �d����%
;�0�ʨA�k�׀*�x ���\����	n�M��e\����SX�[�� � s|��!�\�pP^
���� v�`T"��(+'גp��apk� #�Ì! J ߣ�A�.�;��� w8�C��͵B���aNV|Xʮ��`R�,� �k��3�+B�\_�T�) �Xm=n�5��N� �O�R��	 =���[��cV�w����͞{������ ��Uҩ&�� ���0�<Q Tʘ�C1U|�^"`�e�V f\���R@�h M�e�i �"��ɟU%B�L�A�]1� U���(X Z���u�n�
 ���:��JL�Z	�l��ڤ A}<�h�KV #2)�b� ��W�@�R  Lݡ��'�	��@�qJ}���l��Ԋ Н\y��F �S+:���1� ���$�� '��"xZ_ �m��M��  ���3�X��~�h�!B]���+�/R
Tk�Z���2�4�>��H�s �g��� �@u) ��Q��l30
P�X� 	M݁0� �:�`��r �	�W�.y�Ŝh 1��]�� ����� �|�3X��*r� �N	���_R�C^6�%����E'���騞puJ  �-��N� #���.��^ 4�̲�:�q(��bW�J�La�S �;^�˽| G���F � ��
�,n�r U���RD�� 	L� @d�, ��2�V���� iH���
�9]�E��\�X��90��.'� �����(9l
�ா� х3�zh�~�>�逎OX�j ոm1���&P�� Z0V�:K;�( �鴄��) ��d�h� WmAt��ֻ DЈ��@y�\�] ���'z	U�� ,�}Q�K_����Տ��I��� K���APx� Mb�Q~� ��I���4 A��&��	�H)΀��;Ϳ�ɋ  ���$� _�-BԓP��I­��&���i�Z;�:�P�-Hu� 2ʭ��e&M$��j@��h0� r#��N�S��@7���* �,�
ZU��  �R��Y�G�3�!�fq �D'�	����� ��[_Ob�J�p)���-0ZTh�dc/H�� �W��g�Rx)�	�_��p�g�ǥ���[���<��b���l@̈� BA���n�&[�<�X���ʓ愨�Q� 	��߳`�B ~���L[	���'��Rq�[��B
�)A~� �[��+��8Q7� �٢X�x	���� ��n��V�y&�� Q���8�R:�T�cZ�0�#��=�=���Q����_�� ��[e<�	 �h9RA�nz�l����Y�{'�d�pR	"-�@��F�N�<�h� 3|AZؕ2��(X@� Ź�p�� ���d�� f��,��O�57�����aG��W>�E� ����� D|�רhO� �A�;���P��=�Q��7%��WO@�?@�+��	����|� �w-?v� �]Q�h�=Y���q� �v�b\�ɐ �4l��W� �c܋P� �r6��K`�`9�T�VLw@ob(�� �U� �
� wd#.���� ���SU`o[	e/`����QS�`��@��
� ����o+ ^�5(�)g 
��h��� ��^�	�� �9�S�׻.sHڃ�Ԃ� ����"�%;� �bpo� (��N-�Xfu�	h&`�� ��J�� ��^_!� #�8���� s`���]!���%݇����l~{���.#ÿ���
͜E� �c��0 M����R�q�����/��F���� -GR~�o�@b!��J`�����X�m � ����"���� ����: ��*[<�J2 ��+��ydZց*�, "3�E�Yh gw+��ʄ ���Ձ�C �£ٸ鲪 ����$� ���/o?�1(Ma0r� ]Ҧ�X��8�� ��	�0��Jl&��Z�C �ɴ���% _y��fS(ڳ�i+���zM ��u����# �Z����dN�Г`�]+ !��h�� �0:^p
� l�Bv�fL���h���b�-(���,���ȋ1_ U���@`8	�y��������� ����
�aMG�p�N� #ށ��Q?���U��� _�r����u� �^�����}n �]�@�C� 3׈�8���P
-�N���H��Z +�� �U ��h��9Zt�v� ��P.�`鎼�;�H���
���a>
�5�� ��$� סO���	8}�����X�'�9:�U���hB L75Խ`y �(�].�Ȑq %1>��DZP}��2�v�s
�� ^hmu/L� A�$vE&� bf�
���� д�G�$ ܾ @h�#� ���nE�� �"��=�]W�� m����;P0 �Rw�V#� ���18$��� ����ŵ �0C�x��)k��+�� ��1!��p`t8 L% ��M���. ��q8)N�:���(J0�r�;���֢)��i�ӟX p���Gٜ��mTn�'w\���� �גںDf �p���X�!�u��&]P����ϫ����d3O��#�S�<r�p� ��C�K|	 p1+[�� /h�Q��� ��>(�-)��� �M!�� �Z��J� �v���
��W��A�|=#�p�����'��� �S�_�a��-4�٤.�R$ ��2��F�� P�k*^e Z]Nl% �~ �;�
�Q5A��* �1J��¸�:�� s��6UYp)�	@3� W����X L��' [Y�by�^�ʬ�*�_�܁� v� �BG�����/��JЂA��B�cQ��]v�7���IW)�1��oP!�.�H[n�h�_�� �^��� ���p�d�%��i!1V}�`p� �����^�� �O�od~h8�A�Ynǁ�ڮ�� ����*N��8�t����:�N<X�
`�� ��V��W��T�����~�ƀ:N��! �D^��vh T��'�g ��P��	�����! B�a�sp| �̐��� ҋ3
��a �ק�0 �mgIRe/ڗ@3v��� ��4�G��;�=�@`ǘq��wR�A���>� �|E�M P�Z��lp ��%@�V��[��� {1�� �\ �#� 3'���;��� Z���7��g��@�A��.�EO��P�`{`��U>B��0��*%���J�Z91#�?���G�oa��t ��׊A �z�,�+�c�5�؉ @�$]����в�v`h3:W*袑t %�\�=� �/��# �����2 I�{�9�, ���kaT� ��$�� �t�����L �>��xgb ���@k�O� ���8�	�L��M�*��p�@��E�� �aR|��\�� LK��ж���Π�RW(��:�b��s���}�D�� \�=��V��xhMY�d���@b�^|t� G����خ��@C�+���@U!�Y(�)����`
�F����@N��'&� 1����Z�/r��a ����T��HX ��P�L[7)혖�� �2���W��:�3�%${�v�Y��xN �8��%�;@s�\�0� G!ʚ.��.�)��w�;����!ӫ0���^ �Ux'
�p�>A	�pP \(�*��^ �)��|�m ��r*��I� RX��˘�v���X�� !�\�gXo�B+�U ��1.?� 
��y����CDЪp� FK��,��� }��x�y �`��؋2����@X� ��&$�D( Ac.#�G� �0*C�ΰ�xJ{� ��<}�d�	�O� ��.(� z6�j��*� ��A�� +S����e�<\u 0���>k� r��RИN[���6�1�+�,}# ���i9P )�`�%Ӊ��Y�|\y ���<m9V໸
�h�麋x�`i�Yhf}�.U��� b�!	ܵV &<���y* `�Q0��
�@,z�|�' `Հ� �� ��\�1����Q�St
�P@�ߐ� 9�UT�A� �M`3aϫ_h({��3�0�U����� ���f �&�s��H�Z 5^��3�> ,F?QX+�Jz)'��`������l���� /]�5� `��"(ì>I� Og6k�o�	�b����f����?��A h�i���K� �-"%0b� /�3��[�� ��C-ZXD�'�p���u �8F��1\Zr�L�Y� �A% �/�� �H��>��a������� ��`�J��V 'Y�B�S P0�U\���o�Яް )��$__w������Bമp�� �KzڛJ ͦ(1'	������D��B��]E�\�T�J����@+�*;��(Ɠ�@T[֌ ���%+��s 8�^�i�کY߀�p�%)�� 
/x��1 �� �\0�{ �l������&�p;_rpr3 �%�x+�� P"��]��	��h��
!ro�� �����"��?�ɳ� �@���n�X��;�HV �><�� N���AEF�:�0`a�Y��	���uZ@��c%��йOʁ�)�&� �0�~RY*̳�� �
�^ �ʽ��e}� f�~td/�� �&���%��@���tk2��r�)�	Ő���N��̾��p^�@�L� �+��� ��_�U
 ��O��x#�k��@ߦ�Q U��*�2�w�����"	p�Ơ�ϲt�@�`f )�h��3� ����[0� )Oؿl}�8 �H�n�U����p��J[H�� �F�%�S�\W�g. �[!�G�j��Q�P��� ���{3	� fQd
�_��pm&�< [�O�� ����]�� �O�}�/ ¡�YS���+1�-����`XW 2���I�# 
��c}�q���.�9���*��x��:�y� ��x� �W�� 
_G� ���� ؙ���8�n_ad��{�� �:j�Dw3 1�A��/� �����Ɣ SazqǸ����	��CN�1�?���&����� �4�,�<��� n���� �)Щ�����N��XGF0� 0���fY2 ���K�������P��w��+��h ʿ)��d ��s��� �<0�r�
� �%��Rk- ��I@���Ov�h�(W��P�rp�&A� �+oDu��Xl��靤��p�	� W� �U�R� �r�;�?p������ȀU�&�	��_� ��J���hX�/�Q�$��=0	� �<
��`�A�>��Y t��z�ý ��(]�7 ���b��1� ���	 ������ 0PȖQ~�df\�] �1�nD ��x�"J� ]<L	�� ���{.����}E�X�R�` �ua�xhl"�60���:�Қ�f2��* � ��30���h�q���웂ƈ�>f�;� ��5���< 9#8���{	�"Vrb������2�V�)$^	� "�ш�,3)G���0� g@d��b^� 9��J,u�p����W :(��� 	|i��B� ���1�P�V�	�TUZ�f�� _9�e���!=�Q��N	�Ä�W�5��dT�� �p4X1r�M=�N� ���A�h U<(H,OB��p �n�h�� Z M��2�	:�򸀊ֈ �ZwB�@��Xb�,���� ��>Y]�� [��(��S O�tZ���
���w��̀��h�I�1���u?,�ߠ�|�	���1]��P���� w�z+�-�#����0�� �$	�A# �1+�EW���c�Z4����1�;��Adb|�ث�`��>�`�ʟ�~�K ���s��h�Z�.< �� �+�\a� �z48����g bV�~9�� �^�HA&	R���Qބ	���N��f�����hby�%~���^`!�鐽��{f	�ӡ1TP+��#�@���� ����c&D V+ؾ��H~�<�/<����@Y�O�N ��S�|ͽ~ Ǿ	�]�D��P
eh8J�b� ��#��W?<�7��	^�^%� �>� ����Ӫ� %����p�  '*���� ���#�ci KV_^��' D���b�� �C�����F>}B @��R\�����`��|� �����y!�V�α�� �2��M)a %�W�	��'"T2 ;���%b
�\D��(��h����v1�S0i�D\�U��I �w�/v� ��K��<^�� �%B����ر USP�y[������0�9/��X?��p���*��P��4� ��(j��)��� ��
P萰� *��]|�`+	�ZQH��W�L���%���A�� �Q
��>�<��>S�	ջ6� I��_���,�N%����ȃ� ��3��k([*`[h� 7
P������n` 钿�HȒ��$ ��WH �j�T�� `nVP�� !d+��]Q��@�A���@�� T\$hgR�� 'w��"��� 4쳢  wd�.#v� �Q���h>HTc  �]+� ����/O �R��
��  ��?���0 ��a$��s�u�E���hq/ yI��Q��L �i�� �Rs�	�����] !�����\�3[W ��}w�8Zh�|��'P-�� ��{���R ��@C��6��T&0z��f� ����_�(zZ]�	0�%�����#�u g��(����z%�o�t�)��� �����[R ���^�ں�?�u)%��ȕh,z�9 ,�*k�� �1-�V�� ]Bex�[X�(cR.�Y`vTA�@U]��l �d�� R� P��!p�sX#��'���T��S =�8�[YՀ ��Q ��]��� ��/��Z�' ������;<d�kh�:�1u" s+�|��� 	��� QP ��m�
-s��,ظ5" �3)��7@M�LP�u/Z<�; 3���.�2S���� �
�R� ,%4���� �?��1��O�
� Q	G1;yu�!�9�Zf� (2�������_ P��s݇�= ������r��(���O����6�������~�G` ��Z���p�$ ��_��� z3^����� �"�X{� � �ȸ: ���!��.��u�dO�g��3�|f M����	� �v�=H���Γ�xȂ>ڭ�^�tl�$�P�( `U�oQ ��%@�ӸH 7�-,e=��G&Y�Ȕ���u�U :8� 5.���0)LQ�`�<Z�w ���:�����"R1����|���V� �J���0�f���d��t� =��Þue�[�ѱP�x�� %�&_��� ��I���=du�6��%� ��$_�^ �<bkV��w��C?�Ŗ S\�(ԗ  �P���؀ N�S���5� b`-+߃� �d�6���.L ���h@� �\�'f� �!�EzS�� ���_C p�!�Q�� vfS�Y/��� 
��9֝%$0�Ǣ�^u� e�/h[����_f ��V�^��B��	�`0�A ���[�=����-�8�h}�;����Y��!��+ ����  ����S��9a�<�	Ǟ��.��-A�P���j%�^ �@�3�� �2�S��� р�C�|�r� ��ܠ��ۈ����27�(d &!���� )������ �ƺ�����~^ &�a�K�O>� ���l�ue������ �\�#"�(� 1G�R�d�Y	�����~��A�	�A�5�j� fY7�by@%�&��eЃ��O_0(�Wዀ�ԉ8�� G+� w^"S*Ȼ�V���_,� ��~�� &�+���BZ _���3��=] ����[% �X�V!L��J@uܖ�� 1#��ztN:��J����,�
��*���\ ��� c�4�,$�0 ��W.���B��� �=��� ����P>\� N��B.�]��L�$�&� q��3�h�|�˔T���@���-�O��������Y	��%�$��)� J[�>��]�v� !�KD��N��j_@��8�R� �U3�Y�� y���@�	#�ZX�Uh�i�ξ��P��U���@z��Bh���O��ı� NT�.B1�	)a]��Y~� �/�v���	#��2�o`@/|�-�&��a�ɴ`��� B���]Y� 1�["_���c3
& ]��p*�J� ڇ#�y9�P z"3�,�
]ʘQ� Wu�'�P��3 !�1b
���� #P��9�Wp"�^ ����J� >Z[�4�@�����t�a��{�
�����r��v`�p�����5[Q�(u@�>t~�LM ��&�'����h� ��u�⟑��=� V2��b �J�LĒ
��'�?Z��Х��X�s� �N�0�^#� �A�RexS ��o	�Z}� V$\{Q3�����j��}��� `N*�F��D"��@�� ږ��u�F )��	�] "�_�|�<�b��}T�;����� $)7.������mM	��� M�*�HL�컀�Q��] J��k�� ����K �0@��HPG.�s�<����0X��� ��v҂��=]��2�R�Ⱥ Ot������������J  z��,B� ��T6P �%����� �vad�]��?� ���	�i�w�,�k��^ ��
��H�s� :*ZKsx�
-� � �Z ���ђ�T��ƅ=C�%���	�tXh�ȑ8� �/ ��_S �8� 
�ްB [0��|�U�{ɂ�P� �[X��� ����V� ́Gm$+*��g@PQ���L Z�?\��!���q�0�;B�g] J� �%=Y ����RT� �	wQ����ʯ��)��� ��NH�5&(8�@�eoj��U �Q�u���{�0�aZ"(� 1��pGƌ�5�'�Z�XYs ���$�l� �)^��2 �Z3�a�� X/��V��  �u�L� �P��#Z�b�� ��=�l������}�0�# �!5B%.�� H��-�Z 剦؞�"�pa �0�[��WL��� h�a3�	�L�� �[�D������OJ� �L��� 0�ɪ��[����G�=)��P�T�&
L�X�{s�G��h�Je!h��� fNPR�G�� ��0"(�{�2��g��RC�� br.��~� @P���J$��:����Л�/5�u#�/-F<MH �
Hc[ ��?ۉU� :�,���` �֏�E@
 ����!��� rZA�k��3<a,�)�1th�b� 
��x	#�v>�{ � ߅�n K�%)���/S����P��� f��h@c� ��0�ZS��A�C� C��V�3��� |�"���L[L �'��:F`��)� ��,��( L�ߔ8i@�n�Z��� �^&�Sa��N[,�T� �y�I�$p4 Ղ
��R��ǃ���Ƥ���A��`�@  �1����� {����K����a؆� �l�Q�}�q� )��'�XqY *S�Q� �
�}�������WI��u@@	�\_� %����� ��������:�eǼ�	R��8�\�Y1P� o.�� NI�a4޲\f]�*��� 9<x̓� Z+^T�\8�\�� ���P ^կ�gQ�@0�h�R��O��7 �rp�VY�(^�滗�v- �0*R]� zн��i�k ��͢��3 �D��h�i *+׭^"�= &'�Q�BP	~�]� A��_ ��WX�*/� �R�ҹ	��S�hL@����8��� ����QG��{Eq��0��P�� ��W�`*� �۽4M�� � �П�|�q�d[��/(H���؛? �3��
܀�0�0��fyZ �=X�-?! ���	8��� ��~�ar h�5���.��d�a�7Q��:@�Hг�p���`s��D��Y��o��bW��] *���Y�1� {?�Ä� �)�o�'j}I ��G_X!� �׉V��� �bG2k��"LY-�<��	�Z��*�� :��r͜s�V�O�� ��;_^�E;L ��K��v>��W�w���'��	�,1U ������N ���&S_�� a��i)J~�	����l��Z��C:  ������R ��[���� �X3�x�y 턓mb�� 	"�k��*�P�gs<��}' G6�.�&� 	 ��wq���X��x% �bspi�� ][�h7}�*�q��'�١	���)����d�� ��Of,� 
��(�$���1�������6�8��^�#�U��(o���_�Q���.���%mc���J��'� ��+"ω� ������\y ����/� �rI �=E���u bA�`[G � �_JI]C���c�V��@�����\я��*V�X _ĵQq�;�<u���cf��k�_ȫ�N���\� ���h�>� s-����~K5|DQ	��l
 E���}�x �d�K�p ƅ�e�Bg@ Q-'>6�L5�| ������ kc��	~�X� P(�*���> R��鋠z ��	W�#!��(_��������0��M ,��by)�8v\�Q�R��V ؕ#�W�� �<?1'2�$ �Z_��/� Q��rU�BP����o��� ��
�\�2>�����_�b[� @��=��3�P��� 5�8��/�6J�l�{� B�����Y����[���_4�E���&�`W�07V����:y� !�	;�4S(�� y/�d���;8� �	�Q0� ���#��m�ր̰X���O!�0�0� J��h��u ��'�.!�y�#�fh�;��Z�Sm~��Q�(K��̖H[&L? &WN� ��ϐ ��v�&�%p<+ 32��Y³ [B-
��� ����,��m �U+� �0�	���p���l���T��60�!)�z�A�u ���~'��H �-:�R�n ��	c[� ��m�x� ��/�'(���� CYh��G$�N
�0� >I�! �B��^P� 2fS�Z��� �[�5�
}-���X ~���(RQ|��� ����g�r�kĠЭP	� ��^T
ǴuD �@�	V#� �,?�^-�j��P����y �R�:���� ��Ʌ2�C�4����3 �}�dс ��0�(�QY �jB�Z����.�%��[+�8��y �BVʕ��݅0������X��y ���Ӹ��� 3��	.A @0��z�^ 9�`W*N��#T"2-؀uc ����� (!�����T���sa�Q���h �aC�Z%� 0V��|5i������.����� �1��*'� 0�@�b�5�t�ـT�� �`�X��S }0��-(�vu�~��t��<
髏/W�) ÄB�Y� �E 1�0� ��νj��{]H1�	?��t�8��u�p@m #@����� X1��F"����/����f���A�l�O�p� ���Ī��z ���q�x� �t�� �� k	:]�ql� =SW�ʿP 
���/�xQ��h�&� I}1Z�!JY�/��v+�B1_�� ��$�A ��^j͋`D� ����ZI ��w��� L��,�-` 8(֘OZoF���P�������(0�1 �L
�ӌD$ k��H/K��h 	���QBa �U� r1M� G(ҹ>���$C�\� �(���Y� ٍ��ƽ��i|  ;EMV ���1�^�\���F�� \o����� �PQ,��a� �+�.D-���>���	:H� )���B�
�Dj����65N�=�r �"H-c� ��Y�Wh�b ]*)�VS��0	�灀ϖg>���H�Ҁ � �k���(� �+0���	뇄W>�]R� ���%`�}_ ��*��lP��:��Xp�x �r�T6��3 ����τ W���\ >0�:��-/ 3��j�	��uh���Z�[� �a���0�� H���� sA:��X�{�����&�pj= �\/�r���l��l�𮗥� \�Ed�P� h����ZD��*��_�		��EU��.��B�Ya7x0CwH*���+D�8B �����H"� ���)�� �]��_$�W �	vo&�.��6V��s�n��Ő�hI �g�	tE �_����"���q .��.�B ~bQ5�� �u�^�]�Sy w�庎P�  I�O_�A� ?qk��܏ 3�P1/�Y ��K����%���(��-r�s1�����
 k�=+#P"�� �e0�� �^�̝`��\�@,���0���;�x�X3���P���  ��a����<�� ����  E*��OC�U���j2� Hk�l��|	 Q��?�>�`��)O%Y �Z���dn� �2�R_��4@@�&�V� �P�75lz! Չ�+��� _�Q���� 8;�P@�LFu�,��� �h�'T �a�.�n��pH���� $�%�<c������Tg u\U�z��0��~*�a�P�T��X#Ãnr��f�u� 5R�'дL����!��@/~� �����'S #]��	)� ,��� wP����ݣŶ�K���,��%ft ����BPy� ��p��N��.��KB�����z��(��P 	���R> zk,M�P m"�V� 2׀c��� e�z��A ]
ޑjDv ����0�� ���T'���3)2`�Y �霼�	-�qن$��~�= Ѐ�ö�� J
��Z�\ 5Q�/�Ե�����LH����U`�[sK g2�W鷩 �d���`� ��h�_c�n |b$�Q� u���۶��K���J�p�Wcq?� 7�I*���~S�P݄��yP3N������
hm�� �?�/X �[-0�	� ݇<�j�h"!�T�iC_;v $d8"�����ac�1I?�� ���yڢ� ]:6W��f�|;� 0ծ<��aXG� ��`p5J� ��lid* ��g�5t��1�`P�^ �(��B>E !�4LP� �H3�'��2(��a�����ŀ������\۝ ��-# !��,�LN�:S��s�\�ZY\" 1k��0� P/B��q� E����{=��X �Tb��V� j/��ؔ�Q&#	@(� cX��vĺ `�!�_)���A Q�v�w�9O �����/�`�:��)�= %�A�RwZ,6 ��	��a �N�!� ��i,]�I==n��yke�_�"���H�z�0��w�B�}�Yu&��h��FjH譌�>���ߵ@�FiŦh ���Ws	��2S �+����� !�Q��պ ���y7-����
/�qh�5ްx l�>!N �nMY�[�)��@��9n� K�k��� I��mjJ���⹚��*�>\��h%�x�@��X^�Q ��*J���< ��������$�, ʸ�%�� 1��:�[u�|�E����`Z!��wS	�K�iW�F����~J&�>B�qݢ�w�Q�; 4ۿg���O �e��
(�� �5 �&�q�"���Sɣ������e���`e� +��R��-� �S�]��$ E�OIX߮p ��#� R¸�_���  �[�=� bv���n{2:�] zH���1���(	�Y�>�l؁BW����12��� �4<a{� Y9w�G�\:��ˊ@ѳi������ۀ=Ȅ�w;� #�`O�t͸ a�� b��� ����� �h#Y	O0QGa� � �k oS�%�E2�!ag��D���c�.	K4� ������ ��;ɻ�cg�p02�@ZS���T:�怟�|��� UfL	�?, �_܈1�� �X9σ�b)����怬}�0 h'��ޠX�� �;��X� ����a�x	 BA�+��%�� ����Ċ �vR�U^Z�?6)�4 o���bå�CлpP�L����k�)� ��T&�!�0�A�x ^HXޅ�W K������ n������ ���[9�So �_�1��� �Y�qv�� <|�L�� N(�߃hv} Q)��
	�� SE�����5Ko���
{3 >O���@����'���� P�.�� �ܼ��!�Xp���`���=~� wq�@��h���c?�H��% ߴ����iq�/���+��ye޼�*���t���@�(��&��,� ���k�M�`��\����"�@ň��� r$j�_ PR2����h���MJL;'[������)�zQ ��Ӌ�� ��	�XRiY ����?� �P�H,T(� L��X Ư ��F^�� z�p=�ў� \�
�kPU������+ ��Z��)��  ��U��/�d���C�Ev��p#�4I�k.R��0����@�91 �^�I��� -7y��� �V�K�W��T���Q�UH1�=�����]�0 �XB��(��%<"s��#' �����` v���3�u nh� �m �����O��"��Ys }��	� �}L����u ��c1~)�N ��P�/�-\�%�b�	0i�=���f����X-w�#�Zh	N໘{ �T�s�ަ� O�tJy�P�� +eU#�3� ���Ð�� �x�0
��ʵZ[�\������$ ���������/�����0�J:`Q ?�,�zӿ���2���*` uS�7Yn��P����	��؟R�} h���O?%!��H_�Q�����D�&T��S)��`��!`9u��]3�h�o�s�<^-���_A���� �z�(�e{ �3�
�p�5 ��)�8� f����y��bӾ�vиE� X��pk
 ��ӯ2�\ b;��� cOH�h ~��Yp�,��� �Ɇ�c�0�b'��$0�� *�/�H3Ld� �_
�q�	 �BU���������VP�	;�O^����X�z{�]��� �[H�b �8g��6+o��
T�^�� ;�q���-J�<�o	�!��t���_���V�&���꾇* P��9��� $E#��U h߈���a ��2�X�� �{f%����\?�� �	#!o��^0Zʹ\���1 ���3�!�� ����/��XPR ��U��� ���G�mW~�I]h(�H<��:�`>"Oϸ ���̜uNE���Kå��\h�B bX"� ��_+��1`� ZR
���� �ʫP/� h�+��� W����_����*΁�z��� 1"`?�/� ���&�A� ���{��� /��Xλb @��l�])IO��fd���j R��D-+�x� Z���=��;��Ib~&�p�� �?�� ]���BQN�Y~���T.Z0��f	�3p��+�	(�@ �$��>�����D� Pō)L�a �]01˵Q� ��OM� �b�5�LcZ \�Yz��H��'1��T|ԍL�sD�0��9�_ ^�bE U���X�/)���� �A���.K �G�'����{�󨶕�?�q�}�z��R ��]�w(�� [�Vݗt�|� �}�v��/�an���:;z�����k�'p@C@�߱��� �}���9��&� �_g� !�^2�Ֆ�8%#��� ���u�.� ���G 9�o�)� ���42�� ��$Z�Y� 鰡X:a_	fʃ��,yIg \�v�	�D�	�}:i�σ�>d� �oNשyx 4�_S��� ʀW��� "	F�H6{ 10��X�RU������M 	�mF|��' &d�Y
_P�Ahk��<@ �3�	���+�\W 6�Dn� �e��QҸ�?:՗�[ ��]�� ��^��)�X� 8h�Y�� ��!��nX�:9� �R��%;� Ű-`�_ �mQ�i%���P$�� ƿXBZ ŀ�\��Q 2չ+�HG ��9V��<�1��#��*��	�t�,�J;�!�����/QU��1@ �:�����d܀?Y�1_" �mP��
 R������;� C���t� ���V0� �3��� °��`О�,'� �g�b99% K"΂�;wٔES���a	� ��'U�г�� J�����tm����
���ڀQ���|}�sP �����VR;� ���(�� ���#
�8 1�!�W���� p5�e �Z�a@�H3� <}^!��8&�ާ�p�) q�?�'� (���%�~dX�	 �����9g����P�v�^���
~�g��0T��hӁ�z�� &0I�Y�MX���± pu%�W	��(��-@lV�
��� �Y�5�䂸� ޽��a �~& ]��H!��F�� �~ő��_D��@��}��$��T���� �������?!Հ�qk��� ��*�Ϯ,w�� ���	��� ����aPv#�c�y$�_� ��hH��� �����\��$�� )�d�S V[�� ^���*G|`�3�g?zt���`�n;� �'��@H C��N��Ld%!�D���[YҀ���� ��-[ Q| �	1�h �}YN� =6�.��f��<� \�5X?���w�� �g�����Q�ʖ0C /��!�0�Y L�ra~�� ����@ �,��	�� [-�`�>O 1t;�:�x�.� -b��}R3	��,\�k0"��u��>�3x?����")D�R8�lJb� �����>(��w�i� �1�N �� t�^�K]��i�2���`/w ���-sQ��� PW���ē '
۱q�8*�/	�ɏ�����ܦ�%Lؚp�O�N;m� Dr�*������%=����RZ_�� �N([��{)�\ ���8o�O]����/�� @��Q��*� C�V��}�� �^/�RYv�`�R�j�� �bi|!�Wp|� ?(���l Jyb��z8 
�2Z��q\ NDmtf! ����ʿ pk=_R� � ��I|w�`Z���i<� fh�KR��� ��H�4J�� ������ <S�)��� ٫.7��t{C>�\���׃���/ YQ��h�E �(���ZX� 0��)� ���P��.9�1�qAԱ0�^ �
�m<#+z|�!Á�P2� ���~0���{�vQ� $��q�� �_���h �����~ 	�Q}�n�(�w��p= 8��Б��1변`z�hgS �$��#y<a�)b��~��:- ��HjhJ[ ��?����_�x�4B ���J�8� B1�鲯�� 	�_��WY���}�������S\X�� f�FтL�� @�yN���~p�d +�[�" ��Pw���<C!���n��1 Z�+��� '3���� ���s̛����� �T}�h���3�:a�p�& K��-�1,R  ��i�� p?uD�a� n �)��� �R1#�B[9=3 O��y�߫C���0@�-��P6�@y|	����R<�* J��Y��]n�������� 4w�$RV�o ��;+X��� ��8�>� |S"��l��
-K�0`��r )'�]H@3��+�?W�@���k�t��L�i�b����ؑ �Y��A��V�)S�q�7bJz���@�����1�h������_p�>�@ak��] "b����6�\�]�rj>�I`�� G��JQ�	/ D���S� �]ݼ��� R��\� H�#K��) �;�ꡌ�* ���i��V -#�]/�����nP@�Sj����e�+�x�(�>򀁹ly,\��3P����N_��
D	i��F��|� *�
�h�%� ��鐣���C)A��Ш�cͧ ��&/$�h��!o q=}���%��|��q 1�� Wui	?�z �nhE?�% TDB#Ң ���� J�ͬ��� ��Xy�� ��`t	Ÿ;�P�� ���]�x'ט� T(Ai��} |fq�LMnD!FY��:��� �_��-��<���@�w�C�T��ȃ騢�>[��*���?� ���k�� .�2�[Z�o �E�
��"ص�M���O@V�<�|��7 �&��LB;� _!I�P.� (�+�1���~�*��`GҕPC�Y�y� ��	>����]�0 ��Qo ��h3�,�:$Y /���(� ×�'E\�%`#���_�] �˦�ݳ5� �Hc�X[W ��/�)( ���;_̦~<V\�h�0�S �-��[��>��+��� s�!ųHh�逹�<�[ ��2��K� _Ų����� �T
u�.?�=��?�L| j�(�B �����^X0� �o*�L:���.2��/ �c�e�L Y����+� Q��W��z� ˅�X�̰bPL�� �]�/ �l��	QA@�� ژ��i���	����h�e� X�%G L�5�x/�� ��K� Z �O��
�/=�'�8��,^J�ܒA꿠���y/���*� ȀëYw�,�	뇭<�u� ��� '�� �_a�S(x������IC� >�#P�K%� S����T� �!�D�$ _� o{�y YB��7"�� ׋F��!ʘ�O��.�A��`�c��,������A��@W�hx��� �2!�0�Y��lbp���Q u�U��X�
��%փx� /���;AP*	�d?� �f��O�|�ß@�
� B��3b�w ��(L�K��& �B�E�>�R�֦5O�2 ��]o\�(P� �$������p�X�o����@�R �x[�d\�� �6
� ����?�} �0�!`��G X��Th& N��x�
$�J� �%�f��	��h��vYd Gup��<���jљ1�:��R]W/�Ӏ�C�U���O۪0�P$� ���yq" ���m*_j���� ��� 靵�h[M 1^i6�� �� �����7���ઉA ��Q ���V>�������~(�BD ��F@��2�,�+\��	X���p� R)��t��}$���W #E[Եd�� "�	�YU����Qn�2܋ĉ��) |��} �E��Ļ�A�FpK��3� Q�#Z� � �S	Չ� ��8��F�|�s9ag����D^� p�s�m�8�� �'䓗b�KxJ(�9�������-i8|n �u�e�[�W�
��p��7 ��q� ��Ý�jS���Xt YP�+�g DX�H�r���aI���#[ ^H�Ps� �0�hS��u_ !���+�i� 1[��?�<Q��pЂ_|� �
��Y��xM�%�~��L�,�@��H� ߨ�3��������f�Y��	�>\+���n�3�Ծ {I���qu K�@J> ���5% W�ibU� �Z3�R`�W���׉@�� ��@�_Sa��Zn �+[�Q ��V�{�_M4�����yH�+ �?���4 �A�;-� }���F��^4`Y
�WC �����\ ��%�H����-���N��� 1��XI0�� ��Ky�ǳ�������P��x!����^��"'Ք o �fY�h ci�tQ6�+ 򨅱�����k3 ��s��-��zhS�r����m �~��>wr[ ��^���hU �6!�ҥ+x �&Y�?[� �,�G
cfL)X�� X#�W ��M˙D�� 5�B�@� º`_(�� ݄� )���{� ������j&@������8[��X�`��~�� {�ғW_���In��Zv� Ӥ�a�$�� �k�*��Y� |79E@8
�?�� ^t�_G�� Ig�*�� 1�Z��	U��� q��ST��8�'��0]��� ╀V����m9�����H�M���� �Q�� ���ݘ1	0����7� ��>z��1(��� ����"���f-����SN\��`uE=� ������R��ޮ�����!��읞���E �չz��,ꠈ��|� ¶�醵���Qp� ��ek�� :��N���[}��`/� S�\�T� �ͭ������ �:�W@$*c� D�J��s_��	�@�< �L�r['� q M�4-VX���P`�v�A�(�8��C���!���BH����}���d� \JrK�T���� �6�
� (��W-0�"�S ���%��4 ��(�
��F { ���6 1��rC�k*h>@��3/� �,;a�
�_`���u`9}�.^/x������p�=_���@�- !�F��D	�����1}Y�n�&W�t��b'���
��ؘ�.�BY4��p�� "c�/ѭW0 5#����K�f�Q��)�������@8� ±LUY}@1 �hoK��=JZ�`��!��b��Y� ���J� ���n�N �����>l �� ��Ǉ �
ޖqe�=�t� �ع�����+�:" X�D�?rQKH���Pk�`�O 0�~^��<���'���3 ִ�)� e?��P�gG��\��Z�p@  �{F���V X^���~��	v����0>(8՗ h�N�Q �&/k��7 �h�j��]��P����q )%�u�m� ��.��k�Zh^�H��;gQ��v ���w���y����V�b��� � ��c���&˿� ���%'0s� ���2�^ �9��"��#!.�]�� �[��7�� ��<�3Z� DR ���>���0A��D� ����� �A��)y���g�������"ݪ ��1� ˟87�R?! Ӌ�F	EGh��J+�@��/0 :�m��l�p ��=>�g�@ ��F1��] ���Ë(u+v� G�Ɇ��2��gT��@W8�4	 �1�� c��2���V��]^�A@�)U@��ɧ�v ��9�Z�O]� 0Y<�?1� �/���h�����A1��0 O�����u �X���?�^	�R�� �lf6�~.�=�1�8*��z ��@́"� ��e�
I����o~	���[1%E)���� >@� (����/V|>��{����� ��5��q�o/�Qs��pS J��7t�l Ç�e�"�����h��@ވĠ�0 �U��E��'�� S�3��Y ��p)�X/��`x ��W� 8�H�޾� �t�CX1��� 3!}Hu�W�*���| >��-	DH� ��$��6 �Rpŉɺ�s�2�H^ ��F<-U� ��@v�� !�X��.9Y��ٴԫ�� �Ұ�%�U?�><Հ�q�~06���	 ��Xw0-�,?$	JA��{ y+þ ����̶�~�����@P�i��`����3 &�Cr(\	 �
�_*�� �������KQ�; �B�� �T����� �Ё��5j��0���*�9R������A��r�Z|I	%�stPr��Y� ���J�V. ���L¶"\H�0 GB�y��,�F ��ƖL�@�.݅; ^�h�=��OAC�W!��:ay+ϰE��8�� �\(ឬ�Lp� �.�JB�\�n �RhG',� ��;�_>� iw��4�"��!�<u5 �I�LZ �$8Q��� ��@ mR/3�T�n �fª�L<y� �]�N�Un�&V�#h��� ���,���$�� �;�)� �	�{��[��1 �h�~YJ�����) ;�| Z�����'F\��?,V��v?�� l�.oP:�Y}�?�}!ב�
�0�&� �2�E�;  H����vP� �I9���5 2�d�`
�C ��]R��  ��/�� jZ!��@i4�[�5�)`t '�Ge�=�}L|��� 8���� ��Ƨ�� +c��Y_�)�nz� �h`%������z��QW3��b��XnH�������@��~� �/w,�.�L�b�y鋐G�5��S��Pf��0� ����Z- ��1��u���%�^��Ĩ�� d��R� �>�,��q���06�<�Ý�s����! �K ��C1 ˓�}9�h '>�t&3: ��\��Z� Dr]	���X�1��lS�ԁ�	[`d��\Y; ��.� %�&�_d ��B��� 2W�EL�� ���(B���r;�"�.� :0� Dj-`A͵� �pIJcG+ 2��_�& Z��jϪ� <�B)f�
�C �(�^X�D� ���E��Z� �:�w�I�՟�@	��R�@�����|�=m���I(�S��*���4��)͂# ����SL*� �R��>� ��
1�˰� ������L ��^�ް���\@��֚ �a��n�� �{I|���wE��c'( �P $ �}��.����4~��ȿs�-�`[Y�p) �n�y�-WQu	3�RxG �H��q��� ��GK$���i��P �_�� �U �~f�O��?�� ��u|��>w�yL X�(и8�	_���k�� J������?�hD ����.s �"N��5 ٺ?�	� ��W�.(�� �\ q/т��7 �ĉWP�OZ �vu Ϸ J��(�z�D ���9pf{_ >���Έ �)L�E'B�� jr�s��}�]����Ѐ��j��k@����;|ʀ����Z~DQ+�����A����Y b^-"�Hl� �� ����$]��/�Ǯ ��ڵ����,b-e�%�z��z��O_�ܴ��
0Ā�!�F1�����Bg �A�@��� �S\��T,G� ��� ��(�l�Q�qX@�F�P� BAa@��]��\�P�W ���aO"� ��*p�� � x\!
ޯ� Գ��q�+� /��
h*zt�V���2Mө <'W 3���"� V6�� )�_�/�u� �m!��u�e� �Օ��o��b
J�X�%=�&� �Ϙf ���
WM�:���*����թ��^�( �z6 ��Ǭ��� D\��J(�� ��^A�M �D۪�Su m꼨��'��޹�n�zj ��Y��f�~V�� 1_�O��� ���טC��;�X ��t��� lx8N�_u� 	�`؊�� �
�E��: �O��� }/Kp���� (e)2��-	t{8�1ȯ�
�� ���� ������� ���*�
�� �?��o. ��� }2Rb�Aw� Q���.з ��Ԇ���| �nS�`?0zq�&�%/�G�^�y��� �.�DLHO9�d�Y�`%U	I_�pG�� n1�hM� P@u���	 -]���I�1������%2h,_D 6��`e(�՚�UY���P���υ� S�gB��bp��[���_�;� ����u��P � ���hv ��
�q�B�<!�n(FP% �c����2X;�!�������LU�	2�@9�p A�
��� �C����! ���L��uA�Vn��!XtCQ��@��J� ?�\"��`z }�fy�W�R��'^� 1�D����}�� p �=�� ��	\@� �:O�Y� '�4D/徐 ��
_�C��l@6�0�Ҝ�}e ��k5�����ہ�;dP��.��	1)�<��-���wI�0G^����5 ���·[t2&��������  �s4)w� C�7c���� �@=o�t��� ��h8�3Q
 ؃����\|q Z1���� ��wo� ܉�)�j�����پm"��]��~�2W./�"�� ��@!�� M���I۬� �j��?�ϯ�n �u����i,	H:�,�L���W� eM�I�	�,��� Y��t% �W�X P����z`wuu9 p�"*�-� G�i@��[ �F�yP�V GB����~6 �0p����: ]��P� ���>b�F�pQ)�@0��&��Z.��t�@ ���ٵ �_�.}`����� 9�Wr�ɶ Z��Ϣ�� :?�)�hVj]}�~�?f��!�T���w�@�,�� ��3�A��U�;?%؏q��8<� 
!��$���a�J�� |w�lZ��(L��T�����z� �h�W� �����^�� Hk���R>$�<tQ7��Z��P��մ q����p&&�}? �_YA
� J;��"&�a �R.�Y'	 ^���[���  ���X�4 ;`��*�$ j����� ����JY>w[; ����j �m8��N&�� 1�S�� O�B�ˢ( �rC��8J�{� �tP)h�r I����C� ���s^�:o(@H�� F~&�\�8�+���(�ྤ� ���� $���18���N h�^L��x� Q ��
��1ͳ"�@�n �{�N�Y 
h�t���� G�0��IR�;�$>K1�
�k9�� Buf� v�q��	� �ޒL��� ���]���> �;[I�N��&��Ű�v )�Esw!� ��_qW@� �����h/ �
ŝЯ( �	 Ƀ,�� 7D񮁌�O�� H�A���	 �h�J�[��̠���2�~�rFpW�1 ���yZ ��#CM� Nq,�)*� ���G�
 ω��^U��� i�_A1�,�Y�B+ 5}0$�!�:�����'1� ���:��L H&����s� PK�$d~* �����H�L �mD�������i�`p��\u�@)���:*q� �+�R�� �J�\=
�� ��Y%d�x  	��|�� h\f��K��](��$%�*����3�=�{��2����� ��Y
Oғ|� �v!���//�pd�O���J!�6u _{3��	X}�Lu ��D���b��w�E"	�ԍ/�� R�*�@��n �X;F$V ���U�?� ���xw���~� Kn�2UV ���� 1��KW&�<J��S��-��2���˺*~� ���8�[&�� >�P�l���,��\ ��NA5uk���3�g�K@�$�Ę����@�ՀRS�2�2�g [� �]���U (�:֕�Q-s,��4��n�~�� I�|�_�WzBq�X�� �{����� �Z�x�� �i�l��%{��+ٖ���	E��p��[�m��~L�A�B� ���r�2 ��IM.$�� ��(h%9S� ʒ���G���']�~��� ��C哼�� �l5['+� }�I���b %���~�� �H��#@ �WK�x��V�� 
1�Z�)f�r �!���H�@A��=� �t�V�� �g#Ɖ� ����i� `�@>)�*� ��擴lT9Aw &})k�ec1���D�� }�Zکj�������M����W)�w΀Y]SJ �ۆ>�e� �^���A ��n�'� T)ߋѻ@���@��Agk8�i�1ո��0� $0�_	�/ j�]��� Sp2X�;'� ����^��I G�R�3�!�S��,��'�N	H�z dwXɣ�� (�;��� ^�Y�˗ м-
�t&���/�� `������"S��V`�* Ѻ9��,O#�?�:��Ѐq �!�XYI��1 �ļ�x&�� ��f�[9��� U��#_�/ ����2 d�'[H��������y:��ݴk�0�U <��mhx� �bA	�|]:�6�'�� I�F;�B� ��H� P��ѯ� $��6���|�1��QU�p��� ��ZT,m�h�U�ψ]��<�
�ߺ( ���TW!�_
���%P�}�:�Wą	ZV��`�0��_ �_@�K(�V>�3 e��^ 0�q�h�|{��%k��F�}G�- �dx�B&paH � �hL�'�@���z!K���~% �u�k( Z������.�j7�Y ���O������*@�W� V�)
��� TZ�y��R �':��/0�S4��xj�A{ �6�� �Љ��Y� �����-�鵟P���H^:��4å�>/ ���
Zw� T~=�%�z &1�!b�� W�{�~��� ��ڪ� 	X�c��AI �¤Pux%N ��(=ؐ����ž�� �� �� ZYg�����ȅ�����?��� %���P<� p�l�W� ���8���������Z^O� ����/�@H P�	����� ��½`v � afC�Az0� ]��	�G#�w?T:P��$�SK�~���� �^Y��'@� ��
֗��>��| I�3b���Xf�h����0�ᾢ�d�
���_3�!�+��b�(�ٝS�X��#-N�Q&MԾ ��`�Z[�������%�^����U�� Ph�ef�E	� �yA\� Z)#?��1 ���(r�Şw ��0����R[� e�� X������� ;�p���)� �Q��T��8%X�� ��f��� ��^��0�L �*�韁��/ '��r��v��N ��ùJ�| ��4��� ����p�� :��T	�.��^I�;H� �Q�ŭ���_�w��� 8���n o�)59 y}6 h>d_��R� }�N��<��=�h``Ow�w��ܾѸ���\h �&Q�M1|L� ��V5�S +���LULon �Bw	�� ���<�� T���֖ �ذI}F VE�5?h�H ��z$D>Z]�U%l�2��(�������� ����k��� ?�}z���{ 
�bf[�$X̖ G^c�� }���+�k r�HN�%�A ��}�P� �-�+ x��̈�b�3�$�� �q%�*�8H�c D[Ӥ�� ���(@ 8�0�Bu�  \��q�V��>���R����EԄz2 �,�_��0F�|� �� �`�� �pX
�-0 Y�&���Ȼ��� +�[( �-�9�q� ���
� (�pN#� �I�O�a�0 ��E龻 �.�@��(��^+aӺ�̂� #�e>f8U ���*	��>�Z�7hP.հ� R�	%*'� �/���I"H?��S}eł�� ��B��R�ԣ��E�$���๋��X9\Y���[�W� �7�>V��� H�U���� Z���auX�C 2��%H�vRK��a�˰L+�6�)-�p ��P��ܹ>��	F���� (�0~}��w9=����w`�Q�N T��M�Ob��bA�Q@t���� ��?�%�fh@l}w�dPD�� ���uZ�-T@BɅ�#}t\g��@�VP�]p���*�X ��� ���Z��Hb<ЛבI�>�$�� �'%�]�E� ��pOZ��� ����ė��=W�	!;�h|�~?� 0	�Yu� �\*��� �+�]�V�:f�� ��k'3��p���,h`�C� �L4�`���2�'-�@�.y? �3_�$O Q�Y"��� E׌�b� 9}��Q�	z� ^(��G�[h}?�C��� ��1� ů ��g,��' �[)@{Y� ��zT�1J�=�u 	R�B� ��M���� A�K�OB���o����r�h^��� �þGv�?���5N"��'��_��[ �0��`\� ,!�|F
tC�Z���;�pq�*�`��Ͽ�B  Ǫ5��K(�ޝq��0K[WD@���.�Nf�� �"J��Dx �A���e�0,�)��" �Z�PU��E�w���" �{��L5
�|E����>�	ȵ�� ��= ��9N�Ð��䯋 YZD��9�+e�f��/�KT�a��h���@�6��| ��I���� �K��@E�W=�ŀaG3&z{ ��h�l����o��9�r���3��� $��p�pG �S��Q�7  #_\Kd�g �u��BI~*��mH�^�^�A@1�xP�_ 9�����GQ�����+ ȅ��/��7N
DS�	�8l"Ɯ��^���@ �i�2�Y ��!�0ޥ<�����F��g:�[_�l��Q bS1���� o��	��fU '/�����a	�����6�Ey �)I���	1 N�A��� pD�^)�� ;�/� ��`����s(��0�K	��}�p�v���6|���d�jV�8)�_��*w`/�:�/��� ;�1�B�O���@�G,�;ʀ*���Kp�� �@�[��hV _�ǐt�� �H���$��W�+ݩ�`� LY ��[�����N�/ E��]��D �����H��.Q1s&��L��4:��'��|��� N��_ �0��nv��Q� -�fH�G< ��Z(�|, �$�2�P�*!ы0������5�%N>�0�@#� 1��hD� 
2̺)!��?�ay������:�>
_z�� ��'�( ��4��N�/��T�8���	)�S c�UDW�� �EOq��%� eL;�Bx�H�� ��/� �X��^�� 
� �%<�v�䳨����)��٩���e�:�Ǽ� �h*?4$� ѽ�&S���'��Ԁ0m��cx	!���P	�� '(נ~YbO	G��RQ�s��h�<NJK W�H��� �%�o	l̀ 7^U����
�ե�Y�~E���@�_> 'MZ����v� ����# Ðw:V1[v��0Q逢��� ڤc�bR(�_���׀��A�	 ��nQF5��JB�" �E�,�� �S����N 0�%��@Ľ �J^ԇ� Nݾ��+d� .U�{��4��v�)s@��P ���zw*�p� �,��!�XAD�8�J�cW��K�[ # ������U� �
�z�+��%��T� 3nY4�� ��l aF�R��Xo��
��@U%v� œ����' \䧢��4�M���:���r��� '[0��E� f�.�k��eX��1�G�T� ���S��
 ��}���| ��찈��� ⢊V	�')0?g^�p$U�/m+�`�V �_5%�Nv 0���+�*T� ����0 'I�A�� �+`��՚Pt����OZ�?A>Af9���P�˦�W<p�Y. N�D�Z�� �~`=�K w�*��^ 2�VX�rS ���؆[H������u��"�틸�ҁQI	��3.MZR*�}y�, 0�Ј�/�g�9���N�)������@� �W�O0n&Xk�M9 �!%թgu���s�v� �m��:� ���gl�3�� �!���8�(������&�� 	�[h��1� �*5�
� }��]��� ���Q�ʹL�� r��wIU�c�Pك���+�� �Z0hF�D&�.�>����U`U֯ ��a����np�\Wx ��b~� 2@X���6�����3� K�d�X1�;�ER��kS�ʉ�� �b��7 1����� �!���	` h�H�����l,� �0J����r��%q �R"���:��@���2%YX�x ��\ᒺ&/ �--u%^� ͻ[����w�5�蘸3�?/��8�v� x$ ����D�
�I5�~�3� @&�'�q�) �`�S������5�	ڋ�Y� e���� �����1��#�����Y�؅8c����@N���X(X����Q�j����`p� �H� ��I �^�PN���$n �+���!� ����P p6�����_��م�  �.O�O �A�r�='~ ��X�/� p��u��D���J[0�w��aH1��`UN Ӯ�>u_v�I.
V�Qa �lD ���>c ����q=��o8%ð�, �C�H2�� �`
Խ�E0 ϯB}V�� x�-T^� bU N��� ݁Tྤ]�v� U#[�|�Rc ��	v
��� G��U�$� ������R зt4z�@�~^����p�bE�{ �벮�\ü!���R��3�� �����}#������u��8;�H��>�$J���[���c��1�� (ӂ��~ ��M�	�J� j�3*D��q��������hTt ǘCZ�8�v��@����%CRLީz+� �� �n�߱�>u��L 8�GN�" ��k�i�A�S~��JϞ��	 �qˆ�j 3����$-7D��1
 �������(R��ن���\(�� �X!ݶ�:Z�� �>���H�a ����
�4} F��1XXN�ݵS�'�ӟ��t  �JW����* Y����Lu 8	��
�� �5[�^u G뀆���J�����P��� ���Ҷ�3>(. )�Q��_� ��׳fY�e?�нA�턁wdx0 Ni�ޮ�_�\~e4�����B��D��	u ӑi]yEZ �vfO�0 ���U��?å� ;�A�: Ѩ��*.y Gf�� F��9��+ ��½�n��� I�7s�iy�� ]�f�|h ?AV�O/W 쐍����� 0�Q��j�w���S����'� �NҪ@��� ���s�� ��&�7À.�Mk�h�3Z���	 � �%7V��� gR�S��9,`���P>���1����� �,����&�{���.�N��(P�O��)��|� �}�9��@�����{�[ �}hbAudkC�������{�#�
hG��RF`�� �M���K�tV�`I� �@xG$��� �z�����"'*x@���h���I�kw���t�3А�� "�LS�h	H�� F;V�B�2~��O-"<	�$u暝`�ތ ��2����� ��W�h�#F��� ���U%
 ���B#�}T �&�S��*��gӈ��� [Z�鏤��XY�΄3���� �$�	��A c�/�
����(�h,؛-� )��aJ*H�� D@/��  #���9� �JD���
 �T����?>@[0'�P �Lv��	�W Ƽ&o�Z
� T�p�0_{��z�0��X �s@�:*@���I�	"�K S�3���Q���x �P�*�r(�@+���Րv�W��k�gw�~���8>�U� �' �/�� 1��	BP #�w�Q)�$ 1�|X �4���x� �c��pK� ��Agal!8� :� ��
��n=�����V ��rt
� C� ^��$6�����H���3:"�N�\��ۥ��$>���' �e �ܓ���C@)
<�Q 3%(�1�;<-� {�֡ f�^qJ�}�-P��A� ��M1��� x�/�&� (�)�Z��{_ �a��'P1~H�e 嬗إ�I .@2��� {�����> �p �$�yS b	�BUL� ���/�8F���ez�����x ���L�� , ����	_ �=!�\)� o�X
釕�|0��+?��.���4��W ��u�D���(�非�\��o� ���	оW@ #����4D���p��N׸K �	0��{�idY�R��Q_h�S����C�� �&��� Xژ�GS��U��@�� ��f:<�l T�ك�q.W�>H�����C �B���� ��86[�_.%�� �/#(� fU��,h1��ҁ .��U"p #�]�(�� �/��� U��F0�� �Z]����=��1�Y����
5�-�ۧ���A��Z{p乆/�^� 8��)� �L~1-G !>/�b�e 
�xR+�-��؝ꑠ�1�����a�TD ����h!�}2 ���z����-�у����tUPh�^�J p�7����n ���	)�V*($�� Pt����� �dJ��>�*��k��w���� 0�3OC� ��ș��� �ZW�$�� ���z��!ӊjQ������ S���ሸ. 'jw��V�6��� (i�v �l��: W��[�;���/)��9� ,�C�B�3 �[�뺌� �_i�Q-K9����Rz���% ����&�� ���}:)�	 O��Q��� �C�H��J� ��|�Gf����� ].�� ����)~� �Z��1��`;*� 0��� 
 �[�ǰc;���9j/�p07��2)���_��J� ��R�c ��)0M�wS U��] r hZ+ə C��
��\ �I�6�� �SZ��ER��w�,� }�n�� df�,s��� ��lW9@� ��\��H�2�S��%1�� ��O��x (��h�2u ��:B���� P�	ظ�i ��%G�^ 5�N
U�� ��f��-4��P@O��jbv9�`���sC;,� -^a)�� �㠽U�d���p���G?���)/(��^ S؈�i����!�#�{���0��� hKir�:R�pXTӐ@v1`���;�{� �!�� L�Y�P	  �W���1�� ����Ng@  ��� ���آ�b� ������z ��e����
-Uv` �ql�;���P�@X�IW �`x�v, ђ�)�?��}'�Ty���E}G ����*_��~L�`��x�c �7��[�0|�VS� ����� �(�̾1� !ڼ;���U�s�) o�X ��ͅ���_�M ��1v_ں�X��L@���}`X3�鰙O�A��,�E?��f&�[ZLP� �@/�N��� ���)�S� �a��z�� �� _�X, �7%3ʔ� ��G�霑;�.�$U�u�h� �'/�z��AX� x�7��	,Q
����0�Ș �Jѩ��_ H%'Tw L ?����	p`�'�bS ֻ���#� |�30���� �V ��;<Z a\Xd�h&�9o( �򿀐�� �_�/;��=\R� ��IT��� "[�4e�y �~���&� �w�P���[ ��K�I����:A"B܎# so�V�� ����	����Z������6� ��!���_�2Q�pa H,�� E���^J;�� �Z��!� @7U��DJ ���4Xe� ����&
 [��S!��� W��/��H+�@����� I1]Z�4�����P���,/��0s� ƙ*3ǫ9	�AP� q��	�� z(m9��t S�����|հH ̅�G�fƲ�Q�؆݄����pJ A�nk�� �9u��PZ h�U�%M&	 +����9�����`�U��n���r%�����U\�X�')�	�`��� �8"�C4 ��!7�� ���1�^g�9��������T ��ZQ( ��cY61B:�2����	�n9ԕ�%)�{����	� �#ƃ���Ȱ��Lj��� �><���42�����-��~}�p��� *�H���[|�PC ႄ��:�$,�\���Z���1 ��Y_���[ ��Q,X-h4�I���q J��i��'Vs � 󟠫�Y�_�J��Xa ;�-e8 R��~���("�0�J0��}�v@Q�p+2� � ������[�n;� �Q��u�P���)-���L{^ �c}X́ 2���Z�o \! ��w�,0 ���]�'[%b�(�`���� ��f[0Ok �#��S�_���pz� ��� ֵ�Z���s^ �:��B�� �mH���k ���y>afh ��\9Ł�%� ;��" Y(�� �~ ���ZrP R[L��+,@_� ۠���  X��1P ��p���� "� ه����1��ܸExD�Q Ɏ�c�-@�Е.�!��O��`9�� ѿ��v�����I�] �h'{l �m�^,5�\heCԐZ i�j��&� ��"})� �.3��g�����S���{�F3[�B�R� �ZXYU1 �����T V'Ĩ
�&n�M��Xp�Ѫ �]�"	PU�  ����
��8��Q�ҫ��X��H(=s0V �|���� �ON�ƅ C�'�bzz� ��IXf`�FݵT�����[ ���	�u�]E���@8 U0�1�s����1�ݯT�A&�D���;y�l�� �-+�v* ����J9�C�  5.��W ܟ�12�� /�d��� �p�.�h~���i�� a�oP�ȹ ���?�%� ��!x�,�W	_@�"+��0 eg�툸 �1.(�[t����^@���|7��~� U��öhz @���P^�= ƺ4��hn�X�`����[�D�阮 qPV
RW)� w��1#�=��%�^��X"'�Z~�D���=�P�q� iy��	 ���S+�> 0w���A� fZ��� �t~Y K�r&�]h.�� -`��V �aF
����Z�q8��Ÿ��� �5&�OoW�� (X����Kw�wC xW�?R�Nb P�Ի,i
 k��vKś;�	�np ߿��5�^9���,���+�����u�{���!G \�� FO���h���&	[E  ��T�R���+J f� �tK��� \n���`�� �f	�&\Qc �O��#��2ذ cL�w�0\�29� h�;�΢�jB�1�6�Z� ��Q#�����P�`���O ��xHID��y��������?sT�ցZ%Ơ h@AR�� �3��n�$ �J{	�� ؕN�P�= dԝ�ȋ:�,Ѧ����.�/8�YL� W�����8Ț���J�蟄| _�M�'7Du�>� F�ZR,� !=N5o���ڲ�,��}^�X��@!����7��<�`C��Li ߡG��/�=���>F�� M�����9�����>k�A�`���@ʍ�(<��� S>_�� ]��?�\� ��/�y3� ��)h�A�f_�S�N@-�$ � �Z3�Ը�p��}S0H� ��y~R�: b��7!�0�]>�Z���(�
w�%�N��R�O�q@�1�(�W �������A��K�*�� ,XP�y��$o2�@+�� �X�����@���1�� � �,�#� S���p@-��T[���a  �o�U�%� HȾ&�z��,	b� q=�G�� .�12�^ �x�O� � �A���nJ�>H;�&�$�	 ��!.P��;=���Y K�3Q�����_�M<-@ ^�DՁ�d� �$+�I/P �oUv�D> ��O1�u �Jީ��� kϘ���U?��=I��T��}��	̶ҟX7�>A�� D �5���J��p��� ��bȫ�2����+
�`� (��.��Z �d�2��W��@ѿL&< ��J�1`_� ���|	�{j>���[��0� <�Y�h� � �m�NO�ȿ 2��U�~�3 ��$@P��=�8s����l��и�g �Y%�J+� �	�8�E� 'Ь,W?�� 
����� @ҋ͵��� �QA���>�ϧ���i�W hA
w��� +�p��g���� Y�ڍ�uTp/ Z��X��x�� �㽁�5o�v�X� ~+��¨�
UeyP� � 7wS\�ɼ��<n�I�� q%�!�� H(->��ň��/2W@.'���X�� �n��I �C%ks�.�c 9����mS&�L��V��<�� `jy�?�1 Z]�vdk"�i�^����{�Sz� �Ʈ��)�� ^h�X5z+�B�h/�N��?�j-Е�� DK5���;T����P{>B��vN	�?�} �:��w �׃�]yx �2��=�#G@	eZ������ܲ��nE���
@�T�� d��;EZ�	�aʶ���(܈q� $A�z�a9@�h}�b; �g�L����zu�`�0�!� ޣt�q�* �RZ�zw _8�P!KҫN���I��� ���+��`���<pq ؁�Q0̹#�3߰1�=�M���Y�ն�� ��v��\=��2鐨݌� �Ruy�Q����Ī��P;6v	���a������ ��5�bP
㰝��͋-h* }��ݓ�� �K�:UQi���+3`��v| �A�2�]��k!s���C�0 ���(�-P�vh �G�i#�� !�����R� �x0�������X��O -�*��F: ��hX�� �@� �-1� H[�$��+ �P��>�(��:C���i� ���' ,_�Zp	�	�K��)J��8��x��р$�nWZtH����. �i}�s�" >����BH� z!�y'tx:@\�.��^	�����p��� �[����� #�i��� V��d�"y�'8�D %���w3vxc �[s���tv�L��<��(���F������ �� 	w��� ��i/�V��`N� %](��� �ě�"f[  �X�ha� ��^
�;ٲ�繽�%����)_ �wС����m+��pb PR��yr }�z�&ڵ ��
Jax� /�S���&���:h�bY
(�_!��H ��a����S ��'�=p��U	�OeW`����/x𾖷� �1�^�* ����q[�s��O����ah��к�D	��Y$��KQ����N�f�����X�o*� {]�D�
�� ؚ�RU2���OZ�>,�y�:б�:0�k|	�3ꀶ��F�
��yX��	�� C�A�� �1�h���9N�AF յ�%1|�a�/�\�e`H	��I#��@@��� U"ҽ� ����]S�6�:�_[+�9u JL��忢 �Q�n�D��,Y�t "�_1� �Q'�	�mx ��VD�� �[�@bu z�/p4�� }BxUt;�	(
��s�~�%N��B��y:�@ �[$XZWP���~��\ �4ws<,��2�
}�q�ϫ�'�8  �����t\#�R ���0{�$ �Y��c � _�ۻ���
�h�\� xD[��e��蝯���@wg< Zşx�� �\A)Y] ?� Fpg�0 ����r���S�U�����[ (����'�� B@�?Jq0���ؼ��<�2��/.9�� ��Pon1�����U�������y_P�� -�Bf]��+��GБ[�ma� "���,:��{ 7�p�� �`?X��� ���'W�}  �J[��Q�L�� 0kPX�B� �@g!՗]�SPWl@��� 
2�����q^�3���n ���_����t���by�(�hZQ<�π	��%�� �]����{a�U%�o�� ?blh3)�� Q�@*���e\R����Ð =1���� ��
���b� 0�!�A�]��_ ��fP�W��R ډ��=�1 �O[W#��Q�	̊�p���@���#�+� � ������ ���� t~�P� � �c���0� 7�9��� D1E*ܑ� ��0�3J��	��(�� ��@q�2?H�;Ȣ�@狭 ]�R �w^����
�[�� �_|����Z� �Yb�� ~6K^���LP/ oc���- �hw�O>$\� 
*i�l.�% ��0S�� �F���&;. ��D+>�L�� Z5(� �����=����1�恨5�B�V�~��;�܀(�PG2g �[ĶR�� �Z�{��/ �~!� N�� ˶��(�R d�p����A B+2ZU@���$�_X�z�n��t�eP!0�1������
+����:�Gu|	���s
��~�� vN�(�	��Sg��G�L��^!ø�ھ`m��v�#� !lW'O�M���;�(b�J 首�$n� :�h^*�� ��k�� �/�b�B�N������
 9@�w��B�8Һ�ZQj���rH� �I���� �_�E.�[�!^x@t� � a���h�:M�����	� ��]�J�W��P�7�AH)�R!�O#a��`Z\�O,Y� Ϋ�8SG�� 0�\�h�3� ��q��$s� ��p!Q?���*� �g1� ]�����L2 ��>��+�AJ�s��ژ��S5} �j�`B) ��-p@��<�#K� ih����� ����<z����+ �S�aMF�� J�ǚ��&�Ok ��X(� \���DT�� q�j�Q� ��\�� 3겍l'� z�M��� Dn��<�� �:�Yĵ��l9f�����T��g[��`Q|�.+��pSQ3�� 
�I˥�X$8.8?Ǉ������Y	'�HA
1> :��Dc�8JZ2�`��σ	W\�р���	�� G̦���1\��t00D �� =QŜ}D A�h�GH#� �%����9f�_*�"����� I�0���c� &���4Q ��*�u��_hd�5p�>
nװ����h|SBb��)��˄ &��/4� ��a"�� ��^��> j���
]�PJ� ����}�HD�!���ˤ�I`�bNz'��3 ZW��/��xI�LDP��m�������RY&Nʡ8��Z��2ɏ��P*�D% ��JƠ��.:Mb��˺�� Y�3s�>� �GB_jDl��~W 2��O� mՄ��8��@#X�@�>�� _�n�o�8h���%� ��k��E�5��m`e~=Ѣ�C.���,g�V K້5�;lہ �)�}	L�#��:U�i��
�H�N!E'0�G
�:b��������� d����,EoͶ��3`��� �Y�K��N|�Vz�cQp�� ;��8������s��/��rc�Р�[l�� n@h(�t� �;���S=I@�| ����� *��P� �:��h� �N�Fi�I G�O��g� %ʄ����w9�c	�`p� ��+Թ���:� �/����1�
	-�� ��C���*���ҏ����̅��б�F R���Xi�9�~ T"0�.� �-��!�L1G�_�:@Dq� �^��@(�X��ࢃP�� ��Z�|ϗ �mFΰ�� �V �ċ\�i�����0� ʦNX�q �h/G+ٲ���T |M��� �p2�Q��v� t���Z���j=����{�:-�v8����/�:�C����x,���K�B  ʇ��|Z>\ r��
h�X;�����1b{ �\�EŮ ���vdW� 끼`DXU �6Q����L,a�ˠ閶@��Y��}�f�	���`�� ��H �P�| �x���@��A��{�Pɞwg�%��K �a	 ���� �滘��Y�w�X
���%�9f�N���\#9��3��&h5;���P�y��	 ��SAL! ]h��c@� �J���� ���1���� �2�� X+��<)�>�.���޼� ��h�k�\� s�;A��zg��u����\� @�Ƌ2��a '��Z0�� �$��|(�[9�D� l	�>Q���*�����p� ��_Z�b .XY��v�	*؅����gh?8�����Yx  �+��`X WQ"�3B� �t�<��RDw	t� .Z�P�8" )�X����o�F3}ؘ? vl�zIW`]�e�x �\P�TY�A@i@�(� �"�-�k� �,Ֆ�_ $dw��Yh>~p�^��o���M{\�ȭ1� �S�ƻ?�0gM��/~ Z�+���^� �2V�`�)�]�c�BZ�av�p5` 0�UH� #� �+ɽaC�cIp�Y��=���E�޾`�K_A
e�R�C���X�����j���w�� D|��$��6 ���1�^� �Q
�![ U+~��`��	_TA[���d� ��C�56 �E���'��� ����� *Z�>@��� ���'�BĤ _�����p0H2� �^*�zQ�� �&����fxJh6����O��� }���&\�� �Dڈ.���}�c���]� ��u�DPf���g&ʆ��^ ��`�Ӡ�Vv�B��j\a@�/��9�KU� ��_C �-��h�� `@����&�����D�ݲ�[( ����#�
\�ivX HYV�Խ�F�!��W����������v�� �h3-���}���`� E'}�%!����x5 ��>�nt� N{�!hJ�q|� �)����[�7�D�N] �R�1��S�wE%�`&���2� �+�����$?l� -u3��B�?�Q���U�`:�ź��������y	 �W��(��e O�@��h$GT= J��k� !�>A�#�j%�v�n �5�0\
���Q��I�t��&�� '�q.�w���� ����_�Vߑ���o������G�`ؿ�� �"�y+�$R�a �X��.�����)��Jft' �b���  �~ݭ)��B�Pj��V�< �-��s ��A���� ����I�] �%�۟)��,
U>� h�f��� �����x
R 1�����`��XG�)D�X����V� ,K���_ܨ� ��[�nA~o �a �)C�Z:���!��D��콻 ��PA�� �Y`�X0x�J��I>_�@g[��h>�H��zK���2Z �Q�<�
\w�ٛ �K�2(�d�4�
3�  ��S����}� aj�O�m��|@b���7��@����0^R鐡)*�M� �̳��h�tY��U Dy.���&��� [��A��U �EC�]�d��a0*Y�t�$��o �	�|� �*�T� ���3�u M��j/�����,BʀۗU^ �P��nF� ɼ��3�k *��[!�X?{�(i�'� �`�*z�� .pl3�H�~ �:_(���.i�� P���{N��C^�:��.h�1#	`bSW �-��<���R ��q�� ��QG��C*� ��rׁz�� *���DQ�A���]�yM� J��t^��f��AG�0�/ �O�P� ��Q��R�	�U��'g>��݂h���b� ���r�F+' �$�́�/ daÿ� ��OK���C ܠ�XS���s� {�.Y�� R(�ͼ��[��T���
�.��IO'E`�[ b��Y�K8Z� 8�?@ ������VE �EF� ��~�R�-53���y��m e�Nu��\}vo,1� ���hW\V�Á�`��Z,�z�� 
��/��� K�������h��P˃� _8�@�!�X ��v��	� ��T��m��\A@�^e<$� O�(;�Y ��q�+�kr Z�ݺ)Р-L�=��4��b�qV<�E����1��� �C�]�� ����6	� X��\��k��p�$2�_ 
@�K- .�|��x* %Z��5�� JE���� �2Y	�b� ���(��sK/��z 
�9��3p ��[K_I � S�D�� ��0Z��g@/� �M��R8�A ��K��(�J��iֈ��V�� #�������|��^� :9�Q�v -��0�� /�D�W�RS ����� c�-��I`�:¿=Yx��W#/�3 r�[E�*�^1��4̀��N/ �E� ��� ����O�� :������}7 �P�W��u�?F�ϝ�� ]���Ȉ?\����y����W Y!�_�-� �>��Q$���%]"����l�0��2W5ր̻_=�B���/#�X �Sa�덠|�+�r�����J��n�~ ��A`n�~� \����N����� F��X��!�[���S�����(
��9�2�v[Z�͘�h  N�YS֗
M��%W8����� �h.(�d� �"�%PH�  ���X�$��[,)�!�������W���[h �lU"T#����v��8H��kc��p��Yu� �Tmt@��%�	��pwYC��3��'A� ���� ��-8�m����!��B&,	ի a5�� �@�t�2	�~�:���`����w��W�3��[+�=m���׆�Y��#�h N,��'
��\�K���[�N�) Q-R�x��.�@)�N��8��-�%<�M���k��� ���O�q �Whv+�3 �����D�1��)�� �Ke��I�� 8<HF0 ��/�#��<�� J�o�m]� �\�,�u�� ��ৗ�L8�Hp�ֵ�l ϋ1� �/�|bg�|���8���<A Jrm.P��~o狶 ,*W@�'+��g�p�9�Ps�� �Z�z�> U��_�H��1 ����'< 0��)�G;?şήn#.+����� ��H�v��y j���ͻ.v� -`ҁ� z���.6�]��ǫ�7������V�ٹ�� T!|`}"�#Y4Q�r��g0G- N%C�?�Z��k�pU] ޷)ؐ�G ȓف�K	g��^@�|��z_�C Y/�i��V7�s��P�S� �$�:
�j �{e�[p�h 2�mE�X�}LJ9 1����qp !N��t- V ����2` ��r{>�f$�6���/�Ģ�w[H- W�3J���Z<�(�����f������\S�a2`@"q%t�,3�$/�ӕ���7���_��.��7��� 2H��Yܝ��0�Z���By )�(�w���L�3 ��ڀG `T�kZSp�_P"ϸ��y�& ���5آIa ���~��O Ċ��� �!܁ �~/�U �]�FbB� Pӑq� ���S���@m0���8�� �;Ī!��� �J�T����3&)����j;�����:ހ�/��'� ��,�t% �<������ (��/���U �
���u>׀X}�R�p ;�\�˺���pk>à��r�����
)�����a�t���X��YPU?@t��A���V���m���x1 ��I0�W���1� ���Nt B\�VP���<�*	�E��wcOpV�Fph�3=A���Z@���� �~�a����7�p ��[W�%�� ����� b�=��B0h ͈��O��x. �(��$j�'_xY�E�(��t� �@��_ w|O�"��	 �:�!���� ��H�i ����1� D;�'�{�` �)�rK�* ��!�.�����, F(LZz@#	�x� S��-���: Y,� �fv1 ���$�;�� �)n��/q� �l��R�~�������-( � R)�U� z�@ū�J�QP�09�WE�Bg������H�%W����< 
�}��_��;,S �z;����P���n�\���+`1M �%2ۄ�Vv�K\�� �p�6�� ���P����,��� 3��t ����z ��O��T �E���|D���ݰ��$V�� ��di ��!�Q*��{[�N\��X�;^�9>$� = 똈� ��s�yĐ1 �
����� 3��&N� �zQd�Vk� �KwS�x^�O� �� �? `�ZI^�����ϧU�"�� �_�%G8�4� z!��Z8`�@����a2 &	ы���9z  ��W��!_� �H� ��,$�6a "K���	� �!�d�İʽ�2���� V���^�@��w� aD�{T�� P��W2֮pX����G�����Q��Ȥ�u'}����d<�;����� s�Z�,(t��� 
KΙ�*�� P�:D�� ]u����\ ��_B�%Z70�q��X 3��yS�u `�&װ�{	kO瀘�L���%�fX
8������ ������	-p=��〛y��%M����� ��x��	 ��%7�� �w�?!���Lۘ o ]�'Ţ^� b��xr�� 0�Q2����0R� �սH��f� �u���/ 't�բ��})��� �
h �M���/+ N��!�[*� ��h{�G� ؁T0X`� a�$��	 92��d�
�,�����<k�X ʡj4��2�Ýְ��3o>�:�����<m���DN� ��A��"� S�L��*jB��� |�т�Qp 2	����x� []̷�'� ���~��Q ���A�
 a�R� �ߘ� *���'h�麬@�P^��7{�z� �h'
}qO� ����S<��s�� �2U����N��5-h��Y@t`/� ���޽TI�`z�3� �g�1�� ���)/�| ���"�b ;��l�2 Gs���� ��.�(�h �z�:Jؼ� ��S�淕"\	�(u�%��y ^���g��~p'!D�]�p�� -��"�8� �ܾ(�<V��� �"���[�;����qb�3�|^�ǏȐp��# �
L��, e�`;�sY� "P��A����[�N�F��&o�L �A�+��%QWn��@�Y�uٟp��ݤwЇ�) ª��}>!�-�g���e��s�c�O���`̒R��+�PƏ� �T@�Ͻ�s_ ���S�� ��]pvB�� ��w����+ 1� �� �;�� �-d��'&q �1��@�)��V���K���@��:���֦ùt��\�97G'pe �*�w� ���^8c3���& /�@�h�D K4 QT��( ��?%�NtF 'w��]D�( ����T
; *�FZ#�Y kP/C���� 1�V���������\ PR�9��Z�sX��X�f }'�]� OR��j������Yh*���/�b,@���X� �	uh�P^M��j�T�Ψ�ۋ Su��be��;��j �U��! a陀d�Ϳ�E� *5eŻ��[ P��U��� t$h7;�(����) ��e��� ��y���i�zO/P+�Kp`� ��=��f6	�q�8���d�Q��=P%���8�,��o��S� T�Z�
X�) '����Q_t ֌T���� Y(���:���1��?
�x��f�S�9�� \_�v�Ӑ �-��B��?e! ̄��� G�N����j=�7��^Ʀ�Q �����!��V���2�1H�� ���+�`��^����v����� ����~&sD ����3*�@ xP[�i+W w�q�;�C�b� :Y1�X`S.j5Ur����� � �*���e�ʰS�P ׸;�O��`px@)_ �7$�� *d��W��� ����Ν Y�k�3/A��#�����{^b x�+��ql�
� f��,�\\GE�͉_d+Z�F@@�	�;����R���,� *:�ֿ�W� f�I1K�k�2 �R����@^ ���f�-�����#�0�@V`�� \�[K
��S 	���,�� ��iֵ�; �@X�	� OQ��8�J�qȼ!�)"�;8D�ޝ
IvU	�Ҭ������}#�< ����)� 5}]�/�F !LXi"<���$C��Ѝ�^9�y��qj+L  �Y��R�/@���9��\ k���<@ �!��j'a���h�0_�́F��
 ��	Ry�� ���{�	��L��؉�%�� �M��|$	�& W �2�SU +�V�(ݾ' �@�[�� ~�#��gK 7�Rb]�(������-��q&���8Hr8I ߎ%��� ���26� ����<�N �wtP ���x�-�� J$~o�� �|g(��P ˞���v�r�(�~� �B�@��� (�Jž�� �0�4�9��:�1���< �J��$�} ���
�~�[ �X��\� /_eF�w 1��d������P��l�'�S] �GZ���>�_�j�V(������/O���� ��Z���$!��6�yb ^ۂ�Y�� r�ڐH&�[ �ى�Z}D��2����n�'�Y�j� ���h-������]، w�r��	�g�x�`��L'���� M���g�� �I�����7,��TX�@acݫ+���ȁ� �쭁 u�`��J�� %x �~��x����|[ ���o��[hu:.1��?��lP �K��Am t(\��&�� fhs��� Ԋ	֛�D�:��~ �GV1�o��c ]p
 �$���e�wy��W �R��3��1�X. +�!h�KL �Q���J�` ��Y/�B #@SQw�HX��_����O �(g�z@ & WT0�e�R��o u��h��>8�f ���3Ӏ* ����� ��u!��� �1#�]� ����Uc��~� �ō(E�J ��K߽U�� �@�P�a:Z?� ��n_�� ����:��  i�>��(�� G+�h�� ��B����&I`	�Y@���2�J�{�|����,C^�����
�����u؁�x=>� ���Qo ֹRWV�� �pL���� ��ϟ ������`I �0�W��:k��]�4��q\ ��p��d� ��*^P�a� ����Ir� Ո���	�(���Q��P��K���� ��8Bn� �\Ux� �~%��0��3[�YW# �R'/1rh������F��T+
�1�� �}U�/ ��@b$3d	�[��)�!��� �^��h �pG��q�� b�u^�tZ����H�o-?`W| ���>�� (�
����9V�P��\ ۲��Ja�(�^��B�b x�f	d�O�i�P��� E�0�̘&;�Y� UyeR���Mf �@H 5d�	sZ�n���`Y"�\��$F�Z���^o! ��be�3� ��qH��0� �E�.�8,1 QYU�А� `#��N��c�څ�~��q� �T�l��-� )U��?J���>_��B,� yu/�&G �8'"�w�z ��,��k��&��� W|����v� D.�h�@��E��	��2Q�Ɂ���)� P�_�n�� Tմ����	OSI� �T��9��h�k�|�1����#*� =������f �&ă	_�A�̀���q� ������A y0k�w���H���� �-C�)x} ,�!Y��� �5�1{�/�@k�*����x�y�9��f� k��X��S�3�s���� �����5u߸� �-	��=
��w�S���V!��H� ���ZM^Y}���qO�3 ��L�d;�� zM�ax�O�{�̞�)�pz�2�<�"�� X9�̈:V�RS�,T�$�a�� ���[���3 �5VUT�k P�����[�u�ܵ˄��VI(L�~ ��� D18����� {lR	�Y�m0�-�9�
(\�� x���2 ���^zߘ q� E��+َ��WD t�RO!�q| 3�E��>� �ہaq2: ��h6�
	�+��\�)��! ;Ż�T��e�r����"��M LܔSR+� ��G~��I� �����]1� *�`L�K V�X�� d���{�	0�c}ZI̸�>�5�Q��@�Ӊ �A�b94�>>RłpNKP��0� �i]�8� 񐯥��A� 1
ﬣ"��&` �L�鬼% �`azӜ@S*�V�7e �=Ndv
�� �`��nV�t@��@�2� �N���K� �`D!7Շ� Ú�O�0j �btJAXWs� �B!	��� {V��G�(r� �.��s[4 )����6� ��QW�zy !ʤ1u	: ���PX� /��)&Z
u�z�+�|�[��P�Q' ���`� ������%_�#�C-b�>�� U�d���<A" �@4� :�j/�Z&`oG~�X��z����!K���^���@�`\PQ�[��r8� �^[R�1 ĉ��>���$�5�-] �/���> �������H� 3�1�.&�#�%�'��p#u e��{U����jn-� 1O}>�� /i�0��P��!l� ��͆�"�I��}h ��Y�RK�8S�~ ������|� �>�
��7��4E͇����Z�
���Ҥ��%{ ���㚫 }Tډ)�l�z ye��[���HҪ �Y�z�]��� ��0	N��jQf� � �k�"��]TSH�pw������ j~b\� ��	�݆�H3$ �0��N�˻F@��]
ɺ ��I1 +N�ѬH��!�����C�k T_S|�l��Gw�wO�uǠQ� W����o� ň������ �P��V�u ��a�T �Q_�ߨ^� �맵��2���=	�
�a��$:���5QP�my
���X (� �2� H@�)�v -�董=K
�b�	�hr������u %��9�&��`�?��F7$��N�vb���� q�W�� ��P=��� U�'�(�t�� �@0�cA�H <~��hY:�;0�@��J ��~%SI� XM�+!:�[� �r�;��] J���C ��!1��T|�� �2lb]��+����� ���9P.��5�W��c+ !�i��l�����P���d�~ ׿�
��F&1�� ���z[��t) ����'�. �s� �
^׃	���Ηv%������/ ��1�Q���D ��{���<mӀ��w��%��,��f
H1��3�W��� h�wj$����~	�����=�� ��h�C�wZ�l��$���t ��+����& ��7�-��| ���o	 wYt�b7��Ь-��0����X� �B)%�^ Z(*Ӓ�� +YK�`T� �Ў�S^ ����2� �4	>���s|���!ѰV(� ��Hh� |��X�K ��ꭸ��yL�@~ ��bi�|�����'���� V��AU* ý��з� )���� C�4�W$2��I���M��J �ĸ�%[ F.�t��u g$��� ��Qõ8 ���W٬�� p쪠�"�[|YtF�r ��E��P����D(�|�� �~��� ބq� v8T�.4z��W�>(6 �r@h����PD �u�� ��I����j�R�:։���W ��HAn ��/��[wst#��� �����F'Q$>�`�7 �Upa� �XĹBK�r*WT�i ��: �̗�'� Ѿ�4Z��:*� _-�`n�� �:J�R�F} i��`� W�IU���� v`���xy	��Ƈn��\1v��?X�'���V ��W*ɱ�n;�!-�m/�Khs,yw b �}ɳ�#�9 ��Y�!���S��.���:��eڀ�N�D_ g��aJ��>��P�����o�x3��W �r%ыA
�	k��UPP����� �5� ,������t��	)���Z�v�7}$ !ob�
��\p� 1ڃ��[�< U�h��Z"�R�����G q�wg3rRo�;���a� ҟ��`�D �1�
��( �z$#ѝ ���:�.[ ���BZh/� J�L�G�] ��wH�<( �:˸� A�|�k��dX�� ��@�Z/������5r6�� �� һP�
�GJD�O��n������"��k�d%+�\O�x� ƃ'�rLl.}�C'; 	�S� �c�,�"���=�#���?\`Q�x�`� 2#����� ߀���d- �psK[�3	iH�C��}��懲 ����)�	�`�lG��?��2[�޵�:\�� ��QU�\Ka	�r����%�X�O �s����@(@���	 Z!�*���~� ��R �ݐPy� �_0sX��S3��������0 Ƌ]@L��i�`�LST�y <��C��c8ٕӀ4��� 5W �i /)TQa�v�	 ����j BT), ��v� :1	�Zp��� ��O���n�X��q {>�mK^��W,���� )V:ʍZ��@�R���0L !J���@<Ѯ< �ȳН� �(���d�V��<�%k��>/"��_\��	A� �k���m�:�`i}ȩ�ِEdj@;���?SH8�=� �0�T��� �l-�Mi ;ɗ+�_ ���˷��C�\5u���p=��Z�41����<h�� ��򨔮���?�0ЙxK @Ɍ'/-p��`P�O+ 4.Ƀgh:f3���0|����`{b�]�顒$�+�	�ڵW��m���uH���G�%���R�����{a O��;����[а�n� ���\� 왬Pl[�oD�6#�.8� ���0�[��d����a7 ��~�W��Z0��?� �U�u�� /�����e�:� b�=�a' ��0�IO� ���_�| t�3
Z�����ɭB�斩�@K*�u(XWw����}� ��HJn�+� �j�D?�$�L� L,%W� �^~���@� S��.�K"<����� ��_���6 �p'�<����
� 3�c�;�� b���]`� ���D����):�i�\h���q����T
`�Kب�� ,�; ?
 �W!�Y_zx�t �1&��60��:� ��\ ��>�ݥkP"w����r�2}`����l�_@ �h��-E� ��\^[��~Z �a3ϻ�P� (�L�J� ���҂�# �
�J�>j,�� �����p�c� <ϲI�� �>3��� �Kꊚ�= �j����� 	�A��/4 ���{@��且���!)bİ�8 � 3�fZS�D ��0P��Yv ���k��� ��ĵ\�s�� a�ewԨ� �4��V�DH�� ���8!O����Gu��`� �X������\b� ����{_ %��1� ;��wX܍� ��3^0�� *�j�ַ}v� �yx	)�8sqK���z�~�� ��p���Ա oe�W�kLuJ��KN������	������@�� �ɺY��� ��u��8�Ȏ���'h�Э�� �P���9 �k��D�/ ����Ӳw (�\�Z�@P�[���Ո�%������t@��� J�2��� �BG0v��� 勻: >�Q9驀܄}*�W;�>��!�_�p��s0;/+ ����S�w �n��0 1'��wP ��؃��TPۥ0<Rt�:�O��n ���a�՟? C��QP�&2� !�5�&����J([ڮ2�3��Y?�&� �EL�̊ 4e('�\_�� ������ �;	�n\�� n[��F�J��"���hnH�� ��r!'�3 ���д�v�?1�z"���� '�yL���� w6h��%?0� 珸1+
�� �[��� &b���z�M9�-�J�,%���,{ �(�t�CZ��&��BM �A}�� ��G��K� ������� �XjЏdY���c�� �+Ux�4����0�P=�� <"J��%�}���&�?��1؋*�� \�U��-g {!����2�a]Ph��p� �ӝ>��*$�U2'�
X��Zh�51ߗ�����|�� ��{�N» q�(�ng	� [�T|� �N��G��-�� �5,�e�@ x������`* �8'A�\0;NM=>�`�`(�X ^�3�|{���}��UT<�[��.D�� !���5*�c H@V�2�%d [����5P~� =�p��j W��g[�� O����1X�I2�u?v��K�l&�)���% �����j ��1�oi: �@u��&�� 0���?Q ��O2:� H �)�Y!� �锝í����rI	 �S  ��~M�N �m�.��� �ʲ�=�n:- ½�b ��wZ2���G�c�����D�W)؎�i ����nO� �ײ���1��W������ ��~�� ]�)(1�' L&N�
�� P��>��H�?0�衒�R����O p��^� Qy��I$�� ,���Ӷ �Y�TQn
� @0�R Ƥ	G,b�@�P9sFy �3(XZ[W�;�� ��Py�� ��Q��� mB:�O��B]& d�WZ��_ P��;����m !�� �Z3H�=�=����#C ��S��b� ����Y� �����9%o ���a80�nc��YS��o�)Lõ�� �RE����h�*4Mb<ظ�� k���3j>:� *��a��(:�9ӡ�kb �@!Z
�nD �o�5� ��g>(�Xh���`"/ 
�V�|i���@S"���� ��ĝ�4 �!�ۋ���x�	�N������	�Z� ���Ō ��y��e�� �8	��kc���(�� L2�X�
�'��s�ǸPg| hw	$��^� zQ!���  ��U^�`�Kڀ�; � h�mJ�� Ƹ�,� ���S�� ����[�/� y�?"�R�>�� \H�-��&�;�$� ��Nb��,�@ ��������	�����L|�$�6/P0� kfS���B� 0�I\ �y% H��ȁ)�]+���T���I %�(#��� �ȿ���h �Z6$��N��R�@�0��X��O>o�4�]F*�P2Ή����A�_~�� `�2�Ȋ���H��
�ؾ'�ܞ� �ЬD߿Ȑ[K� ^��\����� RhJ�e' i
̂�[	��0XEu�+�<K��	���; "��1�.� �žh<y A�P
���0 �����%s o�K���Ú7�ǉ!�X�n� ���V�[� ӈ����bhP?��S-!�V8�(Z���� ��� 	݇�w�� =��>��?o ���g�
�d��`4|/�W �9Ⱥ�(�|Kє���\�� Q
�+��0��_����U�� ��X2\�&s� ���%ױ�Rk��⃽c��>�O�8�Z)� �C��$4`�j�ɵ� �3�m�K� ��;���+�\@���0�Y�i!�P�5 ��:���P8m��Dh Y{�@ ,���� ��ST��[� C`��y�� �	�ҕ� �(�@{�`^���՜���E=���O� 8�3�P`c��)rR�G��VKPl �@+!��ݩ�CŨ]�0h%�"e�u� ��C�}�* ٽ�g �] dq��# ��:)� ^��x	� 2����`���� E�
%�� �WB���� �A��z�k ��X��� y�O�} �r=fh� VP(����� �@K��*1�  {��J������u����. 5�'�KA�LL�ͺ�B�<��I h;���b5 \��1��` �̖�E��!����X0rh �d���݉� �K���y� ���!�a� ��Y���'(�^� ����.�� R�Ȍw^8�i��	�G�_� ���~喈>ʸ J�݄>��`\��\ ��[�Zp�ǃ��X� �/َG4�	��Q��h�çJ������)���v-���X���R0I ��ٸ��u���@�RV���d�5 ���_���&z�
,r�1�j�$��Z �!D~8&� n��	1� �y�5����|��qf��	�\d����.�] �{u���� ���	��< L�B��h
�o��ù*�Ȏ� QFns}>�ο!J
B��X |m���+ �d�B�.� g��=گk ^��;��{v��JW�By��w qd�|�1��׉�)���?5����z�@�y� �,M&A	3�W��V����Hf=!�t��?  �-Z�}gR� �_B��aC�� �(U �-	!F� ���'�}� ��;bC]>��N �lqK��� Sh/N�1
Ӹ��>%�@�p�� ��O��u��%0�`�>| ���XA
�Hىz��8�� 更�^ ��Fd�<Q� W"�?��� ��jJF,1;�v�R�ƚ�-QP�ty0�;>����@p	�qZ{� �����-�r` �h�(R3Z��M9ؚ�� ���K�f	}�E�����o h�%��� @�QW(޿�}��@B$�1�t�;�,�s��� �����^M ��"wjh �X�D�! �S�4U���B�~��$[��u �J����\�r�9	��������GM/��ղv u�����L> x���3� �jKY�G� {�@���5	�]�� ҃�h ���<�>"Ȁl�O���a�6�H�/�D�%�0E��] �:+M�rJ� ��h�}�� ���n�s�Hi 0׹d�<����,� �_��� �/�HW%�\�,��8K�5 =����!� \��a< �V/�3e�!�` E?�=��� �.���OX��'�Q��	*��N)�p��/
� ��1U;�� S�E�}:� �`�#�o' a����Vʦ[���4<��- 
Ձ;hze) �_�T����� �sm�w�'	��^��-e`0=� `��/�O���� ����^1� ߮�&�"� S�!P�'��wN ��-�^��v(%� W̎�G �I���l�
�8m���$�O�%� ����F���Y�FK�t����܀)�# �hp��� ����ف:$�5�W�j�`��8L� ��O�� )+칵�e(��J�� )% #��dGϑ ��>u	�� 1c[0�Q���-�a�5��� �x�ZU2�W �k聟��ɘ� �������v�XQ��qLb�����@��SN� ��|��Ѐ��h���tB:��K&�0�< 
�ĳ"����	� ���fMq� ��ɖ  �zA�>蛅2��ᵇ��� _���LI�1� ���s]��j�XP=Ѻ��й^� 7Z1�|!���@����O�j?�7Q �����z�l��@�'\u(\��{YÎ� �2*��P�� ��}.겯� )���0V����4 >ݺ$h�lB���p*o~vQ��`+�X�P��@ 3IV��U_ �%���"(���2$��w�������	� �2�9�$>&L�?P�I Y��}j�� h����N�5e���F�>		� ��@"� ]3�QU	� Y,R�<�O 0�+D����bX=�� /��YAg�3�}�6a�Z� \d�j����h������鼷 ���q�c;��� �
��qH 'X�(���� @O\p�z< �LN�^��\?�x �HS5ʻ� 1�s%��� ��w��J� �c�+�`-) �u�C���~ lˁ�� ��՝2o ҹЂ�^WR ��ֈ � \J�?�M� �(����w� ����}� :��<��0R;�m�@6��c p:�`��� ;���[�� +R�k�� L�O	衅 
0�h�UF���>��΋ ����B} `R���|'� �h{b�%��7����\= �-��A�� ��M:������ʍ�=��_	K��R� ����A7|Ű�\�� P����� �.Ջ�	0����V�Z�X� �Y=)hF:_����a�	������H��Q ��o���� ~([�X�� 	�hcA� ČL�1�m ��*�(�IK �U����	,�-D����n ��W/6� R��3���M YT��nx ĴH�,`S 	�҉
�� �Ż�X��� ��B����o�Ā�;I����!w��9"�����Uz�^]��Ƿ��)��"*���`&�9D,�d1Ё�X�� ?����x*��1 ��\� S�ݻ�� nI���Qw�C����P� �F�1�C)X� R23�D�� i/zF�
 ��:a�G� �~���z5' �r�E�}7P Mf	b��\�p曈�n� %�-�hl5�_$�!]��*��>W��+� ��� ��S�� �[�8�0 ��������&V*� 沟ц` ��/������ЭpH{%R����� $L�;	�� ����A��h9P����0 ��8��  �
�fS�R��WM����K �|���wq�I @!ٕ$�� �1J��t�8 ����Q^ h���1�иj �I#�3�)�Y���� �<%�F^(� �3�`æ �[1�_X] �9^���J �B����� ��ps2?��Z��3A��!� ��70bzX� ��_hsV�=�؀�&Sr�%1c;!�)P�0�K�-@��şz� b/ �a�*)Z �[���H��^�%_B`�� 1YZS��&U����������(�u��@*��	H�}[ ��,��0+�\�8A����@ ��M�L��4 Q���P��`]�������� D��H!=�	="XJhɞ�@����cz �!��R������t?�xIpO)���p�0F(�\��9��J@� aY(�Vr �`O2ތ� RWn0���	_��8S` �����v��c:⒀�s\P� ��i��'U
$FXÝ�Z��l���\(���*� d���r�1 ���<h4ڙvH ���RL+>�a (�6lp� �|��2�-\��� �g\(M �v��ێ� I�t+���� @
�Ő�$­	������w��ѳ 5Z�_� }� &�t��mvt��FTh���� sH�� �[ #�k@��0�h+���j�X�Np�c^>�U�U� Sm�O�����瀾��ٌ Z�/��x=�;����`[� �P��@��4�~�@���h/�iY� �3��Ƚ�`z�����}�	�f�� ��D��e������ �F�� ����.) @�R`<�	 �\|5Y�� �*�P �u� z��H�	2}O�[�^�BoĖ
L% �/�39 7hL�)ŉt ���Q1�tW ���P.ɥ�� ,B�����f�	ۂ ���z:�j�@|����0��X�?���Z��� �T���B'<�j�M+�Լ���sn( ������ �Y�J*V��f
���/�%X���H�S �˕�&� �3�J�b4��)�`�v�@� 0�_\�D8݉w�@�P�� �mUH�e(���	t�;����ń7�/�Ќj\TDt)A Kc�2 �,�_�	}� է
��: 2��'.�� �h�$�!-( ��/2��  횕�i���@*.��>��`�Q�מ��� !�f�V ]�\J1ٽ ��[h�@� q��8*Ut%���� F��X�."T$ U��; �?�J��\�$F:� ��H�� s ݋� p�?ڗ�<�1K���w�- )�|+�� }҃ǳ��i�:�=��pNQ �;91� �8�#�Q 4��tU�� �Z飳�Cd��38���[���_ @�K�f��q0 ��dVm
X ����q���s�k_�M�X��w��S���y ¥hBXI�>���"�W���!� ���	�^� 0`�]8�/ iE�U�̳�	��!���
�� <�"�H� i����&Q'}9C`�W� � �7�d�� ����� ��w~�D� B��PAm3�0)H]��������K��+� &��Q ��0�� i���eF<���y��0
� ?���F �% �y����������9 !P�SQX �.,��%?g ��(�"�	/�8V@ȡ��i ut��������Y�ڒ<�܃�î��].XX! >Y+�� I��L^r� ["�� -��\�I�� db�%�*� �2R�V���W ޟ� Bpw�V- �H]�Ȝ� `PR�T�x ��:�vB	*�wq�(p��E �pP��kH_	��B7 ��Q��}�� 1�d5�" P�(9���	 i��ZX�h *r/_\��A���)p�o��0�4�AȂr Q��׼Za$ ͎j}�NA ���`	3�v ����Eu�n �U��� �� A/?���\ L��[�>� <��!XWz?a��h͐8	���u� ڝL�[ ��	�����3���:�I� ?����b� �0т��� �S��CŴ9� ��\�����zҠ�>� ���L��( �mO\;� "���!� 2�Z��ūv�b.���1� r�%<�X hc����{�?p��!�:�������L.S�� ��-�� ��~�����Yt���o�`j���r-���ދM8�p�_��<�5*Ʌ?�`��l ��=\/ ƀU ���31�윿��c=�++Q����>w� bf��3୵X�J2�` ���*q� ���� \0h�Z@�# �z��d��XQf lOr�>L�M8��h ��Z�� V���o;+�ln��u ��ZED ����+�a� ��B��y2�8���	�`�ߒ ف;�'�Ƥ ��Eւ��3X�����m�hq�sR�T���	��
 ��F@	���?kU �l-:�� ���h�Q3�)�IpP	�\� h�}�z�V� ��D�$W����2��x�[� ��/�W�- =3�p�.yQ �+<!#�� ��A���-
�D�	0���ִJ �A� �� �Lʸ'�� (�x�@oh� �ڮ����u�+����x�p���`; �=��I�M����V���A \�	�^*F� �k�KՂ 7,YU����H����h`>�%;� u����� )�N�D�� 3	J�2��y��K���v~�p�H��,hSk^ђ��ɓ� t�0�R#� �`8��Z� �{��S ���A!�p%�_�y����o�P {����~�K�ݎ�0���� �u�
 �T ��[]�L� M�'H���XBG��;��:�
�˸[�
?�� ȦV3��MU�x�@P�N �����ў
ܐ�O1��GQ�H�� �-2�y�j |����� �ڲ� �t!��;8��A�@�j�^HS>~ ����F/^����80x� ���Հ�F^ �`�8�K;���zR%�\�}p�5��� �qZĦ�P�L 3���qr M�-V�tp�p<�e�)@'80� ݗ�d�!� B�h�L�'I ����-� Y���=	�(}r /�<��+ �-,`W��L ���(��K��k�w�/cqxO ZP��`�ە�>Թ��+��p��J� XM�A԰� �1+�W���	Lh�/ f�]��! ��{��( d���	 :� X�����" �Q�o� �钔���� �d~V��	���'�,���s ���2�)�����'n��[0� ��I��t� K
ŌO�%[�ɢA`�� Ө�bѝf� ��p�� �~�H�` �Ѐh�4��֑oώ�gۗ�@a��k+��0��)����;3��^\��+ N��5pv�ː�$�ɴ�!� �1(�Z�,�9)m�@c�9�7� ��y��� x+�R��Z �Q�ӧ i��^�X� �[!ȿV� �Y��'|w� F���]��� ��ZS��B��߀���;-��L	2"����@�~�#��l�Xp��C µ
�� �%6��7o �kp֕T��0‬z:�B+뫧�ὖ !\ �<W�y:�� � ZNf���x�	�h%0�k��AS���F ��BM1	
����]%+� �8���� F���Ȏ\�^սNa��mT	Q�5���@��X �u����%!�\� t7��[�z�_�]d�� C閵a�Z ;����e������ �Ұ�PqU "ܫ���`
�S�Дû���%�pi����*�4K���XVa����
 ���kO�� ?o�S�*�;�&uJ���2� 	�w�G� ��7�lv� ���Q�߫X�{ �#c&�	� ��A�*�X ek�����8��])�����@:� ���/Al.�Zo�6��)� �1^�� Y���|�b,�8 u2E�� �@�3�J	,�_�k����)� ��3�H,U_;$ Ĩ��g�� �@+�>�� 2 �0���S]����"Ҕu�ڇB�?��� $R�xH�k�� p��C��Fu �_��h�� 6IT�դ� �r���� V��\!� �Qy�xc" ܨ�?@ ӽhGiv�. 	d^E'� ��J�h}�  �a��� �/@f_#�!<Ә�KZ�.X�+ >А��I�� ���t���K ��H OJ X�؝$0�>hA��$F� �D݀O ������3��)�.�⋰\�/q� �t_�1�S�ɀ�n �@ ����
#�|�P�߂����x@�g� ���$8\� ��Ϻ��|] ��"0�a� nہ��f��(� u��� z�Y�͝� h-S%: <�nk�X��}�B�
�� �qT���P�Hе ���h'q1N ���n ����	 Y�\/�� D�E�{�� iI6-��r �/
#��y
�����F����	�h�~� ���z�% aS���1-�_x�$ �R���`' U@�͚\�~�BP��Y� З�0�C ��Q��:�� ^	�Y�a�w���WR����d �.��T�&�� N�-p躌�v�� YC��� �����י?��	]Yop!9QɁ�e8��V�z|�� ZFY�E8��@7�V�>\R� ��2�* �Z�Y�% ��h;@ �ۑ| ��_;�� �"��<�� �v�VI�A@)������|� ^C�o~>ea�����K �Q�5���O �:�]��� g�PV�R�HI�u����}�`H�� (�P�'B ��5K��* �����=1������)�4� 3^��K���� ���&0�� ҂��]��%ޝ,}`Z�
b(\w�y �����3��n[!�X��h�V��p�y! ����¢ h��ZAj�� (a)�5 Þ�3�/ h��pn�I��6�{�\�P#L����@� ����}5 �
P�( �Rݽ\�� �����]$~ &�/�0�. ��V1B�[UQ� ��y�i� v]��ud {�� �N
�Wu�]�:�\��/q���ڦ� 83�Y� s�o�(�1��� _�=����: I*��-P2J ܰ�ʟ3 �Ž	��\ V>T�F`�vN %_S՘l��XZ� K�� ��zRr� �^��!��_ �E�(-CIڜ�	��Z���	��ř tj�������zY1�0�\� Tp�e_@{ ���ƀ	bs0 ZH��W�^Q�J�R�0<�� ��VZ�a8��`�*�P[�% !��Y(��� �	eP���R������s��_J� �a�R��
ܬ������"���u̥ 0��2���d	�_������%�{ ��;�)����N�Ǿ����*�7������@��j `�t�Q�� >A�2�V$n�.'�t 1�Y�S����"� dr	�Q[0�Bǃ�-���p� ���/v�l$� ���*f.0!���3�G�9 /��f��鳲����9�S�^Ј����vU":pX��; �.���\ ~"���>� ����'YPS���U��Z&�@�[d���?�h�gq �Q�:���~����{�[ �&Xw�SbZU^ ndj� �<����<8��Ee�x� F'2� "�I�H�[$�0��C� �� ?�d*5T��� ����g�f x佁���K p�^nD0�5��8v���Z�KU���z20� �:3'��" �%��Q8(�Z����#�� A�����.�?Y �����,O;��a�_@9�� �[�DL�B��	����$�8�����œ	(� 
3�=�@ �Yh%�*R�Jǿ� ��!� �:�U���a �"�X��R �D��Q��* �f'[~�-���)	-�V���0�� 
z4�jS J�Ӓn#~�LIW��Z�u�� &�r����� pVL�H�0 
fP�#�}W �S�l�	B �Jţ�o�� ��R��� �h]��[V0 `�l����S<�'�B>��d��i�v��F �hITC �<��}\���G\�� �q�z��{X�Yde�p���)+ �ʩ�	��#1Ҩ���L g&k�3�Z �5(`)�$�h1�
�� ?W���_ &�N�/�H.��1�2����������k���xP�bo q���D��� ����;ah�'��Wt%LB� A,�$?([ ������ 隆W��A&�_�	͵ �j�a ���+��<�
��9��\�%-VЌ=�� k&��U ��Qt�I	t'm� ��X�&�p-�Z�_�л c���Tg� �#s��p� l	�$�*0� P;� ���_�37~�`�1 �� �G�! ��W�'��P�% ��=!�t��w���5�]*� ��Qo� � O%��-*u� dk4�C�� O�0� �Z�"��E��/��������)]�P:��Z�� Y�ꄏ Р�ao� G�Ah��������0(�@�� sm�!��0ځ �Dl ���w �Xz-��t=>p�!����<̄i���Ar:�w1���v.Xx� ���X/�D!�n�`3�r �zx�Ԁ�;��)��p�� ̈�V�R>� ��1�) �^�HS��� 7��ê���!����@]� ��&^��p��)H3fZh�u��Q� ��A;+���@L�D�19G� m�
]�Z�2t� ���S�A ��b�$YW hp#�6�@ QF����2&ֱ9 :��� ����m��(P5�=���X_�s ��$� � �Ճ�t
���"�ȴܒ ſI)���
�Z�X[�O �b\���9!���[����U?�� ub/����>���[���Y���@����`��S��[����H� %��*�� d����ޒ! �w�&�3 h�f�n�) �_1�&�� �ҩ'�%R =��kQ
}E�\v �+�	�0nՀ���K C�*�BO�v� �I�u���� 6B��0�� <%�^�-��ޫ	��U��i�]����L�Q ��pr%F �!����|O |�(ԣ?�[�Z̚��R���i0�
���4��ۯ0�)P� ��|<ˈ�2 ��B0Ժ!i�!����)��s�v����� ��G\��0<�� ���Ǝ��8 ��_�4 �C
<x���B����Z� �����#��܁ˉN���` �u�Ɏ:� 2E5*���, Jӻ!�R/ ������� �F�'%�4m��#/
`l�՚��z w9j� �1J B눵�<�\��������g4@���q��2 ���R�@�t0 ���Ϳq*��A�$� �%��teW �ș�K��� ����D� �(:^b�8?���w���;�	�͝��a�jYp/K�5�Q@��?�� !PF���{�va��o`\ W��V�H�� /ok$e� �[��"�W�ȿv�݉���m}���pA�^%N	g��)Ѡ�f���;#�����*$���^���6 ( �R1�������T� �
�Y��a c(Ã�x, P鳎
���^Xy@���4��;!�?� ����<
  1��~ Y	��|V2 �U�'�;�uN%��� �J�D�rp�f��E�������P֗#}(	���;��@U�l R���/��\ �z�����	�v���~2%��Z�0�и� d�a>5�z�_w� �ġ��ìo����~��)���� ����� �o� ��� �Z0�S8Q�;���L�	Cѵ���� 4S��N
�6u?<��a 8}&\z�R�#�fB%+ �b�^�'� 	��_�u� �z�%�� xO���p o\��	�bD<V �$��U �:>�3�`8 'Iߐ=z�͉k˕��&�! ��[i�;1�ml�3w�H(��;� �OCs	��Y��� ��x�Z�z&������ ���.ј@�!3�ٝ״ RX���� �<w���s xo��b���T���:����Rh�NO ��,��_��#�R�J�' ��q,"���=k�h-.������'�ϰ��i��ή���!��_��ϙ@�?K�TX��L�^	��\���z{J��^LpgeU��qdJ!���K\���N���j���_�. �@�����*��?�0Q�@SV �F[ϜXӮ�����Z�o9'� 8�������~9@<1�".�[R? h�@B�ʷ�_�Sn� C+����xr)�:�`N �6pF�. ��-z�~땐�E���_� �a�5��� ����'�|� ����hy~>K�� G�s9�5 汪��R�� ����~C\h>�m ��]�� ������ (��:�cEr` Ɨ��1 ȷ0.���}X� ��rW�u� i�+����� ��2De� S�����g�?�À�*�d�� � Vo	hOJ ������� ��B��Q�J�p�D`_��� ���p�Ð� Buി�_	N 8Ra
�D ��$+�f��F��%���1 O�cԐ� #u$�L- Tk���3�ǈf����`�I� �2�WR��: ��	�!�1:���L��D�Sp%����W��_@�O)����[B ʙ;�b�(� }B����� qV�P\��% �I�(���b� 
��: �p�DZ�{����C�]�`�0	� ��H�O��*h�@�� �ъ�	�S  �;�����Z�%��4	�I r��t'� �}�y�n) ����W0�Y�<_{��o ���e�^q��,�~1�/�� Q�f��` �>����������	=�������p�}�?�pǪg@����k�6 �$�cdh�> �̮�����H�3ʀZ�� ��OM�@ �����W�� ǕԴ&��� ��
wfI/5 _J�y,	?K�|> uh��{ 0ƽ�¸ �?����Ĭ �B`� ��ޒ⁻n��5k_A�H@w-���m��Z�j�(e��,�B[�����X�� ��I*���	a靳!:?�~� ��Z�=�^��u� ���2XR} ��L|?�5 �h�9gMs ��="՚�f^k�� 
�B�/1J �(��n%:0]r� 3*�[�;� �Y}�<!�d��8@������nj�`�R�� ��	>lL%) �U���Ӛ?��0,6�D
���������9/y� �����[�\=� t0�:�-G�'�@��^CJ��t}p���`ˊ�� ��@|��� ��dk� 	�?ٕ� �����ZE��ad@�go�] O����f)�r���� ������+ �����y (h8��J)�>:� <PK��b �o������v;�����j9^1���E�02��� lC�_�k ���%x�j �rgK���2 LT ��P�� |�����3)Ȩ YRQ�õ	��vk ��ʂ ��`�J/0 � �S�F��� P�lK�5ځ ���R�బ*�v�@Q�i�;z��0��' m���lM %���W;�6�ǟ� O����9]� v�R��S� t�/�?��� )��$|׻ ��_&���� � ��P���*� ���(�� �%�[����\�' �< 0� S#����y�� 3��$�	) �(��dq�����ə�`�  ��V��� �)=S��� �AU�D�� 禰p8�V%���ˡ� D��\ ��i���^�EG���Q�iS�1�BJ�Yà��_�� 뼹����~ �{��W��� $	Zh�[�m ��y���&S" A��/ʘ�&!�> �N�H�P2���@�e ���M�Sp\�����#�[��`ir��}X� ��]Q�% ���h�J l�q�	�]zy cp1N\��,UD��Z�����_=�;��9���Z �=�&�0sB
��~� `k���6LK��X ��p�b &�)=��	 0�UϽ ̾�T���& �߸8���CtP �5�� )���n�8��	.�ݶ� ��[�/�� �|'�ˑ� �Z
ƈ���(��G��n�2�\Z &$'���Ds��@�@F� ���-�Sd
⾂�����)��0� ��f=7ZH	���S��& p�"�)�h����uM ^O��b�\�� �E�~�%� $H؋+�\OQP.�4���� �
j�d�� ���,�_�a���hex�{��� SIV"&��	��CU�^���> `� 1�	�� ����JQ2 �R
��D� *�c��_��	�
u����`v�:mF������h'Ox� _w(�0\AM=Y	�S��VU ��*<�)�=������O�*����,�h&c��"� ���`�A�� ��r��=�
�Z��jD B�����S �s�^��(���0��aLY �15�.����&��^	�? P���DJ�e��к����> ��CSV��� ��O��3.�L�F �J���4��bn�/��0�&�JD�_ �%�T�k� ���*�,!�À��$ Z����u� ů
]�@-  ���L�J� ��V��K� 	���Z� d�Ǜ#��$ <V��x� ޗ�)>�m(��``�o!q TwQ'�����f�_�> MX%��� �-s��3� VT^��c��P��t�Xx� ��!a�� �T�+�i %�7	��"\��W�Uk�&��) �}c�J��� �SO�eE��7Ī˻��1!?�[���	Ik���3 �]����L ��Q��U~b��	�_���Z��`n��`X "����W�Ю���`i��� �X'���/��A� vv��� �+���^� 1ABp�D�� h՟��;y� P���)�p�vZ d�}��8��U�` a���jeGɸg�%��X����'���u},��1�^� WA��h�� �g����8� @l��/� ��-���< S���P� d0�	��K ص�s���xi�נ�H7�P@ ��^2��K8Cf�,� ��="� RUٳ��kP	�)#��߫���'P����?<�16�(?�۠���2 ��ƀ��Z ����U�*��D�xR��@ �J¯Y��.��h<��0K=,��^�������D�E�;΁`+Y �����ܦ�QW ����^M�h�~� 1	�)T_L ke�U�P� 5�t���;� ��\����[ ��X���V ���Z	F�{��c@�-�Ч^��$5��e��g�����LO� ��� /���Z�%<��P��0/o��� �]���N� g���b�@h Pt�����P��9����`�T�p�Q L�j�-�� �1Zv&? ���{���p��\S -��aV�� 
��Z вz�h� �8A����L;X �9���M �#,(��ft�3D���o �bd�} ���� ��h<}Ǭ �br�^WF��޵��Z��%u��  ���~�C �#@7�� k�PS�6OA'�`Tj�v �?�JǓ�( ��B3��� O ��-*����caH+������
��,���L\�㘡c-�U��� Gu@�����2俜{̡�_���U��;�� &x�hkyP� �J�:W��̤���
%R��0~��A� �!�	m8� 1����P� �=�����U8 ��3��.������7]�\��I}z���u0;�R!>�w��Ѓ� Z��: �7�x�� S��W�[_V>p��^�d�YM��H�Xx,��/	$��W�_`sL�p� +�����P3�*A ��(�I�2�	�_sV i�����\�J *�3���8�1 ���d�� ]�w�E�5h� ��@�_���� �k�v� ���D�If;�p�'�X&8s� ��� Ϫ)&M�7 a�^�.u ,)�� n���$� @����W� �P�ҡX/� ������� +���J	^�X�u�r� �t� �J��3.�z~� ӈ��Qv`RW��@ڐ	�?�� ��' ��p��KSW��`��0�� �ty�{r-	�:��1�>�?� f)��"y�,�AbX d{S;��\��p��� ����� T�2��Z# �*���
/���r|��� �~'���>ÀP �՗f� 2aЉ߬�W��sQ�v� ��ׄ0ƃ�� �b|��� #"�@����!� ļ4�� V|Ho �)K/��h^<%�p�`�T�+�ID�1&0���`��~K �o)]��p I���XR� ��o�^!� B@ׅ�P��D�G`3 �!���b A�� ZL����|Q	 ����XEј�-uN�&j�Pݜ��K��@�-Ոe �U�AS�|�<B.�Mc��K��� ���P?�	�`Y7� ��Z�Lq 錉�J�DB >c��M0��`���� ��I$�.� 0���q,1 *@"�\W�9S�����	�� ֏3B˒����πt� �Jt�T�� �%�-�^� ���$1� �i	
��иK�wȃ��P�� XTh�z��+�� YV�_���~��&N-���9
i %�(;p�I��l�,[	���ݒ�b��� @K�[���d �&P�ǩr� q�!Y���0�GP[ Z��� (p_%2�U� ��-�d5 �����W�j#��������������Ǐs� �����(�S ��u`�Bq[ �s�A�)Gy �I��� ^�6��
d� S�$����.��  �ͽ5 T���:�� _�!rLӯ�v�-f�>��`;�ׇ�t�i���� �/G���� 3�J�&�H#i{>��Xn >\2fR"	݊��@�����t�f���nv0c��	�!�P, �{'ލ���J��$�����:H5|8&*�� #�!N���X�1 ~9��� h f[Γ�k`�e� �\��n�C�B���xtD!�k ��0Q����>�� �/¬����%@춞�&�̀0C��
( �S�]���ˡ�^��TSXh1b VK��
�� ����R�r }�]�<^4�\3� ��C����(ҹPc���`Oٲ�ȔT1��<
��-���R�� �#���) 2b8	Ѣ\"q����� �ABPx� ޹_d�� �����^���`����ئ!J���%-��. �8I�>B4t ��K�O��S3N��pJ��M�{ ����#�ݞN��PS(��-$ !�[>3e� h`wi�똸 � �.fW���d���!������; ^�> �	� )�g�L<X�H_�0����l� 857<(� 4�^qrA�iH��]P����X���	�R�� �1H� ?�j�_Z�0�RT`�V�ڼQ�Ĺ#� ��ɶ�:� Duņ�V@ ����r* k���y���ŀ�� ���j\9%��~�;�����1�M����>RX|P =��t5���� 6O��sL"��f�.����zW��  ��uJ+��U��,�!-�Z��� ��8� �a����(�,{u 1��$>,�Җ�W|��2 �"�}�&� �9ዅ
�X ��k~�#/@�R0���2��UK�Iz�l� �)J�{��/�O� 3�����M��G"ǡ�:�R���&� /������� >(����\��;n�ʕ[6AJQ|Ҡ9��0�u�E�| ��R���� U���� O��گX�E0��
� ;�,�?:!Ww�7y0�&� Z)�	�,�b ��\P��� BR+�V�O� oTA���~ �h�U��I	%$-G��\�C(��:,����N`�W&')����� i�! A0\� <2x�B7;"� �����g>���K{�d _��.B{ ���(��1S۬Ά��F Q��HW3��& Ή��b7hi(���2�� G�_�L	�KY�& �>�� ^]���F+K �ͧ�<�1� �	����HX.�� D�\� ��#�� 0^�6�v�C ��iz�H�W �{h,q k=���+� �*5�1� �I#f��r &�N�3�R�/�h�����b��2񊀌�<	�;�S���J��0ua��@�7 S2�(�� �XU����i�����J^�=`�t\d�& �.v`�09�Q ��[�� ��W�Z�� {<�*�B� J��'�_ڢ Y��4��� �[S���	���v�H�
+ ���Ј�Z;�s���È'� u���? |]�sN�@��$S� �.�� �_a �[V���:�����	�b �w�ڴ�%E �/iv�&,q� ��������#Zq�O���c$� ���R@K� �����;�~}� ����'��/0,� vl�^� 8��Oܒݐ�A�z�=�b��X�h�Q���, zB�˿/� ��o	� ���8Y�� �2�&��p ��hk�1d���@��o �� �!\ˆV ��R�]_�� �Eת�\�$ �Q"�(+��w2���� ���@� P������ �	gQ`\�6 �<ׄ� W��ޑ	�0��� xjM C ��D>���q����ֲo`�Z �)yJ�p ��������+���� ��͐�{���m��TX�%�9F�1�5�� m_�K�q[���D%�-�v���c� �ڐ�\� ��3����~� �k[��X?P�� VUδv�n`	<�楀�c�E ���.�0��`���V�[��.3�˻���=S- ��_x��� �y�a�<=Q(�J�H�PW��� �+R̹��� K4�&��X!�p��C�����F��8�i^	� ���'�Uğm1���k �j��T�ʡ �v��b� }|���C��b��S]d Z��°)� �7�ב� ���G�� ��!$�y`0A� {
�w� ]@[	�x1.|�E �u�a� ;_XH�������@: �+�郗^< ����*�G�}( /��| �̸y�� ����=��� 5�%�t! fX�AF� ����`����s�B��U� ��#���?��!����[� B��S���_����{�p4L5t|�Ê 2ŮE�U� �W!�To� �^���F(@�h�K!�#� ��V���H,�  �$? ���\	���ɛ��e,`>d v�Q���; 1�{���� �`���0�f[%��p�� 	1���� �X�W '�� �fZG0(� ����^AU��:�4�B�9 ��)2.����/���|��[��G�T� �0tbDƃ6 $����^_��� �:Hew ���� ��d8�� �\Ag����l��w��~=XRPĮ%���rg �﬎S0�q. ��u���� �����]���Y��1ݰԫ 8�ǜ���i na�D��� �����`� �*������i��,o� �ฮL8�W��_ށ�� 7�2xX�ɸ;�����PGq�F�z� <�����/� Lt�&_ɋQ ��~#��� �P.��2`6*S��Ź�K��/������J��1��R谠��%�#m 4�h���D_����� �(��b_wa��K�+ '@Nt�S 6��
w���: �;��������܉�xD�Ā�2W��j���\Z�08*���d_ ,$N� ��{���� \�b�s�:���q <�Z�z�H]� @fU�u �_)��B�.� ��>�1� �ֿ��`�;�		���CP���,��2&i{ H�< R�8�[������5dʛ�3�0�}��  ��V��K�r���X`[��j�J���L	� OD;la� H������K`�#;�!��2� ��}/�� ��T�	h� ��0�pڷ{⇀��A��4 �h-%`��]�#\R�,�{9������؋� ���QYVo8�X�� ��Ф�� ��U��e`Xk+ u��ƤH�E �H�2�� )��!��,YQ B�]y� h���[� ԥ#�/�1U�' ],���hHu� Q�Y%����=ꉀ�{d�X' [�\�>���� $ކ͖��{R h�`E�2v�s4� 	����XO ���	
D�yO �'�Kw�b�)���oa��;_�΅�ɖ #
��QS� ��KW�c� 9� �
_ھ iӁ�L*� ���
�R 6�u4����v� Z1��;�t���EJ�*�rb >�)wV��' ?g
��zq(�;;�� Q��_@�G ׽�3 ��]�r!у���� ؿ�@��<�M�r�	��Qv.�O� ����� �7�;�Ek] \�V��LC�%�`.Hƈ�u��l	����vW��)(���� ����-k �n��b�
gm�aO�� �0h���I���܍� q�/�,e� �\���Պ 4���0�|9u�,���W�Ŀ
� H���$��b »B7Pe4� +��*��0�r�K-��,�!o�y�� ���d�w< �G��p�# IW�o���a�?� �ٻ[�!iÍ- U+�'8�~�"�w�#]�����8���1
��kZ����d!h�r��ij C�>���x� ��X	�˯_yЋ G�-Z
� �vT��z:�[��eO����� �^h�J}$���]�u ����V#� 5�.W1zDͫ�����uI��;Z�Ͳ�h[��]�� =�;? ぢ�}����� ��Qt�U� P�@2~� ����F�Q �z��1!���_~bl��^� ̿vo���I�N����lsd�- #֡1)�X��*&��D 4"� �V�~���	ȝ�ti|��u%}��R�8cEb �0��j��, J �m(9Q P+�XY�� ��h�� � ��å�^@V�U�apj�=�12�Y[@f_R�F�L��#��)����2�ک�Xw� ��M	�P?0�L����,�z�X{� 1��O�� ��vf����	H���pq�� �fC&!�� X��gl�� �)M
1�� �Y����w*(��/	�i ��.�J4�\�� u3U�P�p	 �]0�1���Q4�hN�	�+�9%@��x�F��ϔ�G �P_P�8�T	QUBB d^-2���� �@�]��K�v� �3��R�� �����1� ���-@��D p�M��5��<�� N��3iX ,AH��s�? %���K�m����oT��� �u�`
�[H2v �P�® �����{�Q��D	�t�:�Ee�7��� �����uZL��}`��� ���w� I� �2h��Z�k �7��O�CX���o`T��%��@�g�'賸�I�e���p�Z<ψ �'��L� �9bQ�( ܂�*��f S��VX�� JK�1�Ɍ ��*�Z0#��q ��.� ��o�RE�� ��p{9[$�0��b�ȳ�	[=^��@ .h�Jo��� �3���<.@��"y2x� ��a�)�`� 3AP�Ҹ �h[��� �����̥� �1��ܓ� "��)ha�O0�����G�r �ˁ�Bx;Y���Q�/��1� �
�9� �k��^"� �������  ���,\��Q�ł�`I/{S��N��1���M� J׳.٪�n ��e�����@�� ��]�� � Y���Ʈ�=�H?v�}wW:Ȁ5���`R �G�K�u_�&�!+ *��� ����U�7 _VH�W3[�{<&��	]!�  �-d;#�� Pp1����	�鵛���E��2��m�X@vR� <|镫�1 �0��(�L�x4 ���u%W�� ������ @�	hX��3���2 ӄ�LM| �S�^�Ĺ��W�� �h	�����|3 _�G�����N��R�@7�Z��Ȅ� hJ��>;A�� BH����v	��ٿ�j����¦[ ��F�d�Q W����a����V=��{/:�*)�Q��T��=K��Ҳ`G n��O�V ��1s#� ��j+��![���h��P� �b��$�Y�Q	V3�\sI �柅pe� ��[�ɀ �%s�	yg>��!-`͢+ �Ҍ}�&�<�B�R0���  ��ָmS�	��`��
�Z����ѐN�� tXA�hL2z ��/�_��\8P ��{�h �|�[��A �釯3�9 -N�+�~A 
��R��W�	u�1��|KҊ�S K��z- ��ӝt/ !xj�k#��ݫ-��2USȤq�жNİ�:DC	\"W�k� F��Yh�;��dpV�Q!�X��Y�� �V�zb�Z�H �J�� ���f�_4� �{��0�^! �.���r� 	o$�Wf p4�ը�� �8�	w��.D�^oh��"G���˒�#�5 r�Ǘ��' �}Dʹ�E#�3� gZ`�Y�	���X�Hg�=h� ���9� �OlD��� �R��*u�4�F�	�� m�7�����P� ;(�8X �[b��HW �Kq��*�����0�� ����B���ǒ�ܛ �Y�h� 
+���` �%�|����!ҋqD{�7(��q h&uEY]#"�p<@҆��`p�Uu�9�g��v u=�aPWz,'��O`�� 鑴ז� .����h� %�:$(�/rB׺*�@���+�3��8t��$� ʻ/����P)���牮B��qr` �5�n� �����R� %�E�:��At� �`
1*TZ� ���E	 (�~��"w���EZ�u���gW�=� �pJ��# w�҇�mc kte���
G\H� /_���? ;����� �e��A �׶���(}� Ӈ�V'D�@ 3��1���[��@2sZ���?�����$���� ¹L�N�w �^������PC �)�hPH b���]z9�$9�;p@�ςY)� @P0�-�� U!���� �u�)�� ��z���D�ь�8�@�^ �"
Y�G�� V�4�ݪ0] �Q��+콩,̌" �� ��p%V�{�#��@10� �5��1 �{���7 +C��c *�{�/Q�`��\ $�R��_r.�(;�� ��= 	�����uL @}���F�^ �R�p�4� ��|.3
� ���Y�o	� \X���2�� u�
}:<[_���+=�%��bD@@����7 ��Tc#�� �y
�9�h�{����2�U\�I��!���� ?������ :"5^�� �P��0�h (A�s�JR �- �ؚ_���TO3J@�DLa %O���=P���S��ձ 6��V��?� ����7�KH ����]Y�Zx�>�������퍒�נ9~)��/�f�Q �#����;U������ 3d�X1D/,�T� '�0�� ��B���� ���cϨ���r,�S�K1(j���` ��� � ��>A��� h_��N�� uIDB�f�H k���:S \UKɮEۯ ��ك޽	[����&W�K�� !�(�R��� �Q� >�� �Ä�Ĉ%� MW�O:8� ��wn�ı(�����Z0�� '��PJ��N;��� v��_g��.@`� TӒZ�Jh� K��ȄUw����̓��.���  ���%&@T��X���hW�	�`�Q"o:`l���Jt��r� �͉B�w]��m��؀� l���?�u  #���	�� .�|�͸�`�12�h�M!X�A<F43w �ե"��?0D����Q,�� �J�\�6 �Y�(�� �^[��R>3��B��Xh Dp��?k����%��R�(�܍��p�)X������.��� ��1�Y��*='��PE Ao�c!D�PNr-�����\/�#����	� Y���FX�� y���V 3�\P��#H��K��X�!��� R����� e\h�[� ��Jپ�: I��v����� �";1���e��:��� �h �W'� ���%�-�� 2	�^����	�c' ���,
����� � P"���F��jw��/bv� ~�o�]Rhtq �𠛲��������.�!�@S�[ ��Q��]v �����+E� j��1	���Q�Z�s�\�6��S�X�E�	�c<`%  �h*{S%��������E0ݬ ��ڵ���� f��N�e���L.� �h� O���2��G����/������ȶn�b�g�X�&�
�� 6����	�#�0 ��)}\���+Wx��� ��|M��	w��, &��3t!��U�>����J�-Y��k��� �Q+�T1*x���{�t� p��^7@鈕���w������� 
��-fw2 u�}%v���& 	jO��Ը!s��;��yL g��V��|��i��@��� a���0�"}�����zf8� ��ޕ�� ��`A�� +h-NQ� ���C ��� ��	���@ ��oA�1�D [��{º�� ��W2�&� �ྂ]^:�� ~x��R�� ��󛇁�Q H�, �G܀� ��0 �E�Z_��X�1�x�xF~U )�]���v,��ǎ��Bq�� �	�J�a2�4b�AU�����G�q�ek�! �@�Z�K�� j��n��	� ��Y�/��$��H�&,� ˰����ȝ\�����=?[	�y� �`��|��!� �3���X�(��f�yl���R��:p�Q�k ��K������vu� ���(�nX&�& ��*�� �O�l-݌ R:���ؐ��n���1xB*����%P _-��^���� ��2�	�p N��_��\ s�5@� ��`x�&�85 qU��� �4�����������pʹ\�_���] {t�o� ��Y��� HҾs&R �bC�a;�	�"���-7da��]�_
�z �.�ob�S �� �_��x1�^��`�� 3U_�� ˉݸE}� ��AuG3� ~O�$EUV a�+(��or��D��� ��^!_ �]u� ��BZ+�U9>�� /�t��, �7���j��� �R�؃��X��;`8�w !ۉ���ޤb���P�0�U ��)8¹+mv� 0��2��Zi�`-��x8y����Â`XP }*�=E�� �Ŝ0�th,~.I �@�!� �D�;�i� Pn�"�| x�K+HD?� ��	����# �D��N Y�v-P�`$ t�+и�x�0C e�-$�M �H�b9� p��f��]1 �_$(�`# ��7q�,��X	�[���W0� �<�2�� פ��r�� O ���쿽��,G[�����>�����I-LY�󈻀s�Q0�U��-��8�c R��me ��Z����  �c�����$����`��&s G ��_�Oq� L��V��� &'+�㑠�(�� ��毊���
3?�� u)^�� �0�����Ԏ�BIp��O��(���� ��-+�|�� T��5�:	��e�:=>iF	"8��1%} \��g�1�X ��-I+q aL��V�G5 ��[�f�� ]<W���m |׈�l7���� �BhR������#Z`zP��>��^��X�� dY`�)� �90]�� �1M<c��~����#�� ���{��z�|��ج
�݉1O@Q�����_������o ���lK��Xu��p����>%��L�� �`F�� ��N\�  ���ꉨ w��h�:����+�Q�I� '��֥�#?Ɓ�$�²����npr��uw�@��(I����A�� ���z&n�� {��i,�yPC�R Q�1o�E��� 7�	�;�� &�����B���uP&)} A?��R�� <~��ny�Pp�K��x.F �փ�	X Z�L=����� 5~\k��1n�Lʧ������ ������v�>	 �1�uR 3�g�-�V � ]Ji\� ��DGYE�� ���zR�9A n�p��� Xwmx����� >u��/p7|� �܉��`�Yʙ 2�F9O�|��� �(��Re�&���,���1�[í�Ȝ��-�@nZ��8Jx'��]��� ��ô4�b� e�u��K�f��	���s�+�_����l ,	�
}�@ !W�4O��`^�ڽ����PR6�z #J�=�Äf ��VTz� �A�ds� �i�?��	�P/�ךp��� �y�_3��; m�.?d���@�_�r�� �A7[8 ��x�@�����,`���B������%@�v� ��5��>ug�#Y��`8�C�kp-�`c� �_�^�݋��8 ,���6���]!���и��� C*��� <[�q�G�	 s��FH�� Np�^`� YP�WI ۿqa�6	1� ��0lP������̍x�hcD�y��}bŧ3 ���Ahs|��PЂ����?��� 	�[�x�>;����]��s`sQ ��hK��� ?뽀�g��@$ ����_�q���G�P��/� @\���� F)�h�7 ���o�C� ��KI|�1@�Z����i#�޷!ʠY0$�h e,��(������݀��U� �V(�?	 *�Tf������.8����l P�ӪFۺ u/���%�X�~��S���L��9�$}�t ��J�� ���\���pR�ɺJ��k׭ ��N�]YOV �dW�����ʸp�-!� ^Ǎ�H�o �����K�B=��/�ړ$` �n	2��h�(߰Z^�����ӕ|� �-i{�a?� T�u��� e�Yɫ� �/��j�� ,��a�(�B�t��_o} �^��j� ��X�N�,� 3�.����� ��y�[�< N�8�	C/� T.S�΍� �P�+�vB;�`�h�H �w�5�[��8*�� n!��D� �v�������Y(��R��?&򏐼0��u�� *�TN�"� �@#c{��eU�D�ܖ7 �Q)$>� ��h��K, �-��2���9��o�eA �]�67��� ��ܮd'�΀�j���e�H"`��ޘ6����OE����H�瀚�/�6�h�X�pѕ8Q�s 	�[ ��)�V��W��f��հ 6��Z��� �%��\z� ���U��W�ja�� �h�D|/����S��:� H��@�U�� >a�3�uv� �hF+�* ����3p� �;T!��R� `W-)�
�� ���@��W|.���J�� ��}�{x�$ 7a���� ���B
�|� P�w$R/ �x�Sz �	�V� &�'ِ>-} �#����[R�Q��pb���� �:��hX �R� �� V�����' }����� ����,���2m�a���	�_ f�(�0��VkA9*o��S���A�
l�!� �UX��L�� ����g� tE�1�(�� ��N���C ��_�)I1�H*��(�a�	���0 ���K*z� �?���F ^ lZ-��� +#�����b ًPI����<�+�҈��%�,X{ ��1To�\�Tcn�hG�0軙wNK��rv�����%� F�5_?����YT2��] ,��s�E @h*K$P� ��8k�� b�W:�_��.��~���y��W ��@�ɉ��_ ~�a$��'y��� >�t�[ �%�}|��\i�s �?D�F�)���ܝ�М��I�� wڹ�,��� _6�� �!&�)�S ���-���� ��M�U���[
ޘ�"�� �W܋ `�Z��\L" �ē���I> �O �y�v��W����\��<���6�~��> �����G ��A��C���(� ��꺀J�� 0��u��>% ��N�(:(P�� Z{�k	�� xR�i��.$@HO �g�� Ї��
�i� ��Z迚D	ht0:�� ��pL��3*�Y�� $[h�tu���#)G�MH� �;1(]�7� id�z�� KN��p� ���~�� ��Z��2�� 绨��ʬ�,���"�� �U��&�$ ]��I!��.fˣ
����[�?�� D��a�cX��� ��x;o H����0�X)  ̣�_! u��[�zG )Ӻ����` r�TDK���Y���ຉ(P%[�<`��/��^�o�ΐm�� W�4������fpz ��BX!�%��ش c+f	 �_s"��q �2����ú4� / %�R= ]��%���� ����N��H@ L�~�-�Ή��n �$ ��/tK'X|	+i����@���
�_㌮���Ч�^ ��[����<B���2�. �
��r�P�"1�@J�G 04 �gJ�l RV�w8�����k���,N�����@o����Lgd V���#PJ
�1���;`����T�=��)��@�ﶉ�Z�ט��#^
�h�'�2�J��Y����8��@�ɟ�%q�Z�9��/�_������ \�i����;����!��)���� *֐>f�-��x@ 1�0��e�*� ��rR�Lܮp #�P1��X M4O��a� o̊!z�Q �gj���pӋ*�X�+_<	���p�:[1��?�;��Q�� � ���Z�Q�y��`��v
	��u P�v� ��٧>�=�T*3��y�N���>��V� ����%_���2h
v\�"�P��Ȁ[ 7��u�Bz WA��t�� �d��p�Ҁ ��*/�z�+�vO���A�� .�[��r��3��!� �B�� ��V+�7. �Apfh	����к�D� �:�hw(Y�- nt.1�ï� q����� ��
���>&� ��$�ݒ	䓰� X��\!�>
8rt^	���@5�6����"�W� ��<�����L�. t1χ�P���ʙ�%����X��{Q��/L�t� �R��%�
UO�e�A(���[� ���Uf�&�*@��� ���
�( 8�	%+u�����KR�b��w��� ��j��n� ��x�b ������*��(���lz1� ���AV�X�$^ ��(� �hn4W��m�V�^���Oؐ� ��7��� U�+�	(� }ʊה7��{�k���� �$�2�]� ��M^�@��H�'���xg ��Uw�b  �6�X�O(F �	S����{��k�+�@��=5��������p�����U��p�Z�.�� ��L��<>�q����j&�G�@P��� !�C��	�S� �@1��'���U���t)<� L���3e��� �a�g�X �PU��E �j"��3� ��g���Y�@��h :���� ;@�a�(`� nI�7��� 2�?P�O ��H����(c�kK�����[� 6#�\�� L�1!�J}0BY���%X���L|Ss�T[�`� �W0X2���VG�hr��`�� n�R�O��E���La�B����`�.Z���#�&2��� و�[��}��
 �@31�� �HIyK�u��~����1D&��[#��x�+�( 2�IrV�W������ ������@��0%y��� с��5 �1�B���U�2�[�ń�g��\��)%!�L�,z�  ��Ҥn/��� �̚��
~ =����:! M��έl�+� �,�0[�� p�G�V�g��Q��n�0u��9_�?�� ��ˀ��C�3إx[�����5Ϻ�eg�PB2D~�$��r J�;h� V�� H֋�9�a�Y{��A �0�!��2y��G�� �` �\���"� ���!�4k�-(�7@�H��B� \c�2m�� *ѭ��:��� ����_�.�"	�V��mp�s �|��T Z�`[�a��-�>���:�v؀@Ow�5$� H�A�� �q=���5,{���`cj1Ձ��:ܳ� 5�&�� �<��'`�"��и^�/�^�	)`�#ǖ �b1�Y&\%I6��S�� ��Ὗ����A�� ea TtO�z� �3�SQՍ
� 0�}�Y		+ @�^-v ��E&�9?� zt\��ŨJY���P��^w����ό"�Z���͋�L� 0��xj��b� VwB��>��5DWI0�xP��3 �_�"R���HY� ��>��'��;ә��Ϫ (�8�e^�O$��r�� c֮�
� f 1�XQ�-�� q�����L � D�Q0�?�� ��ڣ��Ø�� �h�p<\�� �����% ��w��Sul�?���?�"��I���C��� z�T�D��=��v�����:溻	 bл�1Z)�@�QX�`� ��+�4����BS@v˝`�6��GR�V(ۻ �E	�^� ��-�3��Q/����Ȉ�B Y�RW=��� m���`���
�3�%�u��,au ��dr1X�8����w>���z�gȟ������V�f� �v�](�R`�C��}niN��r�� �Q �Ah�I.�k�eg���!pl����^b��`&R�-�Zr� ���\�n�7@J!�- �X� ]�x���Wy�2�M;�̟X�@���i*� ��(����4��������SV�b�u%w��&
K!��gԉt �{�'���O��R� `MB�����h�)����s����q~j� v���� mKd|��hLT'	�Z��Ҵ� �,
�K1i 3���k�����? �.(��`y" '���>�� 4�B�R���||� 1;`΀�{( ^K� �3 ���͐�w� ��P!�A�/ �Z0�[���Ё�Ie����ǰ7�W dH	�ِ�@~�5��;�;lmH9 ����i��� ����-V*��t ��H�'%f� ��-X�	�,��< MޅQB� ��ʏ�a/�]-��B)��:<�^ �J��Q͍ i�O�j�1, 8��G�c# �^�ᄩ����������� �7#�h4YJ~�l���E�`�����  �)� ��m�
*�B����V.���d�0�;���z��	Sa���G��N>�-��U�-^ּ��>�����L��Z��_��Ҧ|, �.�HC ��Iͧ��n ٴ��8�� ��/��K%���`��3 "���yh�; N9|��,�a�pǒ�� �7߽_ @�M����.��P�q��~$U��hja���!z�wN ����ƭO��1��w��/� Z�ƹ%�Q ���G���L��-)ҽ ��YhE�5 (���W
���s�� � P*�G�� ��}����R�є�V�� �����p� ��TceG�P ���|�	hd(Ѡ�KF��X0� a�
#ջ� �"�C��XM%�P�^�ɼ�� s�/BL�q	u[ 9���+�`�(�FK
�m_��v@��� �PA��0.� �L�1E )�w/� �n��y� �9XA&D�rs	f��_�����L�
���� _�{���� ����[ ��\R�� ]�� N���A[�@�Y� {`܃�m� ��?�)�Q�d� ���{�1 �SX�3��� ��[�� c
!�Zp��hM�����)L�=K�p�Ԃ��V�'{�$����1�X�-�:ɐ�@g� _G��푄 �����3�� S/E�k����B'I�.�Q� *��Z��F ]��
��ʓ E�_8�[�)�a����a��x�y�)� u%V�� �Z�C,A�1�=;[�9��F�ʀ���4�� ����0��K ���"ȉ��!RO�&]�&	�� ���� #�[��=S �)b*����� GVfӾ ,YF|� ^���r L�n3ʁ��q"G���� ?���d@���/�6 ��� �xZ�4� �����P�* ��?�� � �@��^\�y k�VpCa�s���B	!�2
Ѝ5 ����,n0 �_\�e[��@@�h8�dJ ������s� _�Mf������Drن�G	�[�K� ��i1C.�Mt b)uAf�k�^ �Pn��Ov6 x���!�>�:� ;Z�+;�u�z�@0Ӹ�Hq �5�E*V�@�S��K A�HX�c�<�ļfQS��������@�� K���� �$.��� ��S��,pTV/t�0�B -N�:�1� �8}!J�;| �,�#� �G"Kd������P�P�IHs ד��K0 ���r`�� k!��,��Z X���u_Y� p͕}��` �w䗅�h��A��1:љ�� �!��oP��}2$��<�~.�\�e �mW��T� 	x���_��� c1�e���(����� _�j�k�r� \t/�h% b�a���~ �0����1# sЀ��V�/ ۾"�(�aW ���ҡ�hw�Q��`˓%���� 0Y��_�'* Zu�b��iИ�~� �~";�Y� E\���q0� @HQ3�.KPn���	@��+�-^����v�2�P���"�� ������^?o���)� �5,Z� pB"��0'� Ёꙷ�4�g���լ�2���C����ؘ�-�TpCm_ b����, �-iU�YI X>C���g�>ZR��v�B�]|s�õ�%�X�� �B��߄M0 �hs18�` �����f� �:��b&��܂a�,?�}���F&uL yn���"��~��?��	�8]p���! �XS�滾� Q0�K	���.Pǐ��o� �|+�c�������E (���R "-��CZY8h[�J�]<.� �8�4R �ش�[_��<ų��{� ��i�.^@M�n ��m��� p��2�4B a�(d�)�/,�v S�[H�6 \~���uDe 8�FC<�p� c���	 �U)��� ���8R�^'��6�e�b��w�F�5 >��'��K�jR}����� ;����0� k7{�R�X�� F�\B�19�|�H�������
���cH��1� K'�~A(_  }U0���< �8E�!Q� w$-�V\�N��ـ4�k�0��������~ ?)�g`��Q��R�p5�A(�� �
;���� �{|���H�*�I8������y�9{� 5�G~�� q���ͯ(H��?��	���H]��Et% d�M��- S��p�r� 3�V)���\l	H��>��f65�!�X_� :t���ZU����I0���TɸG�XV�'�d}� �x��P-��BO�3� ���!��82w ��-�a ��?���]z� (�^y�veQ:�I����@�� H���(`U~z P7�Zh�K�N���� C��km� ���{�]h�D�!����0�1�Y`�T2}� �%��[{8"HUt � ،
^9�� '%*rS��|h�ҋN}Ж�![�S&���?���hw�����B$&�.���4�� ��: O���A� 2��]� hawi)�$�3O�ut�� �� �z	<��B� ,��+�*7 ���X�� ��2�S_�H~��,�F��N?��i@0Ø ���y3���[�m��>������F�H� �� X�~� |���/�:W���	��4�1����2�!�Y+�`�=��nG �Db$ �/����h �#����� D�	�[X ���/{����S���2Q�����	����q)x�Z��R� V+�U"�r���`�4~QF �B�Ȇ*Ɖ��)����Y� �x��yv 1�	�^l ˝�u���>�' b!��L ]�;W��x�� `���
�Z(|� �!oL�*� P��'� YZ�Mh��ط"���a�P2 Ǉ�Р��� G�f�ě�C.Y$����%,�9�d{�4`A�ҙ �˸3^G �ބ����}n���1
0*�(���?�� ��Z�ہ��� �s��hew�� F2G �H�( ����o�� �})^B�]� XJ��d=��+?_��-�RW
 �Q��XA��Y�� ��VO �}��^�� ǿ�@��P �z���Y*�0�@�a�Ȁ�o� ����x �="�Y S�N�$L� ���[@�Q?R���|CE�������H�A 3�0�N���q����죻 O3�f�1���X B��Ƒ]y���P\'�q� `α���m 8+�2�\d ���[0n( BP��"���
2�	� �S}[��= -�!�wE> ���Qtbe �$���� ρ��E o"&�l$��)?��-~�Zq �C��x�+ ���! "k\i�U>���n� ԈI��<0��ѷ���v��X�%��|��e� ��HT�
��A ��-W�U� F5L���аR�
���	�<C(��#����}���4�p|H� Nٹ>�ufS��m���� @ ��A%8	 �9���������B!���wfW �L}*X�� ��u��k� ���{��o� ��2�h��� bC��ё-���_;�p�l%�^!���?�������\��  zQ>�/K�:��9���Ү���v ��b������
f�� ��g�"ˇ\�z r�R�ʁ .0Հ�=�0џ1���}gn�sZ��!�N Ǥ�+1�OL���� ���lH_�(d�N`��F&1� ;^��� iP ѵ��ǽ����h@�S)��<s�!'�4���N�`�.BSJ��j	 ��i�D��< �s�/~�9�w �	��X��K� 3[��Q#� ��o� ����P\��Ÿ�+�HQ�P:�X)�[����x�É+�3�ZX� �e#��� �p����` 8aCM�{$��  �JT��� �ǪO0�C� ^�LN@=�� oVӸ'��(e�Yj0��dw���*�<�'!����
� ��Z��1��_`�'ib?�~� �zC��� ׁc#`��- 
����� ��D�1dr�� �����iHx �L���!M �UO��8K' �ƻTa� ����3�Cv�p����`N� )�fh�9w��� �4#Ձ ��o�
�� V�Ҝ`�����`�ƾ ��j�� *K7�ٺ|� �¸+�?�f{ z�o�-���v0K��� @����Y� �N��Qw #?�`UYC��� ��o�� ��=k�3	
�c�dw��u� .l��/� 㵢��h ��0p��z� ��>)�]� ɕ��ƈ��g��� h2Y��w q��K����0�� �� :� ���.�v��©د�Ľ\��L�v{�<@�$R?P#�@��'�� ���*p��_	���W ա&^�6u� 骆�[�KR ���)� ��3B+�A#�q��7��L��0����	˲�>Ԝ�=ۀ�� �R[ D{��ײo� �����_��h��o���
 8��/[ �������1�`�j��� ��n��V���v ��4fӏ� �z[h�1�L�$ I�u8�� �Z��'�!Y �-��f�O���� ��BX�Q� ���%h��&C1��^�f��;
�P�� y� Ԩ��D�� �3(҆	s y�u?۸I$ �|�'�v ����c����y �E��^ o�~�� V��Nf�͏xk?+�r ���YWǕ�9�< Ic�2S( 캜+��b��w֠@�?���~����C�	� ��F%�� w23W��\V ��h�K �l�e� � dS*�'� 3��%G�� ?1�	S���=��� ݶ,�J���	� �&]�a�\�<&�} 1u�5gR0\� )�(�'��.�{o �_�����'�ӈ����� �8�X	�P `�2�� fI��0Q3�;���~�@��k��_�����-_��H�3`>���ҫ�� ����2 �E�����+�� (�3���@#�P�_ � ��Q ��h�	��%F��M ��)�A2����:���a� يQ�G�twX>�� ����c�� �fZ(�����
剰$R����"�@ �'UP�[`4W����\���N��ٶ�%�?Lpࡰ �]	0��Z ��K�
}LX`,YP�'����q> ���ۀ�;�N(�LV��Ts�/�uC�Z�	�6�h�s�$�a�=�I� �5���b����F��(��≍ȩ*�%pZ��9;� F[�^a�������g@X� �	��>
Uh 9+�0���)�^��%k�{ ��d�U��8 �H`�2Y ��h�c��	Q�� 
��	UE�@%}jdb(K�]��1 ��:��+�� ���0�O �f� '>P �(�C��� 0�*���R9 �j��o��°q ��[���p{�~$ �-��|� QT��Y� /=�*�	#� �@��(\_?Lw����=��NP <HA�$V(1��%�Z�.����6�_��#�h�� �aU�-��@X�:o}��#�sX0A�.kҺ�7 �V��b�c	�^�� ���N ��Pވ�}� f���;ہ ���M�<�` F	�;���� ���8�QH� $W�N���<�1������oS������; 0mӵ�R� �:�
P-��?���ml %0�~
*� `����-�� '��b�2
 ,�P\�[-�!�����5_�G �t�� DLiUm\o	��@b��x9� ��#��
 �4�z�7 �!/ �(��J �@��SY 	��R�0#�p�=��
X�)THܩ�'"��ܺK �0.�^��?�O��!��@��?���
����-� ���QP,'� ���Z�@) ��qa!�^?J0?��i 5Nk�'}tK
 n�-ע7E�&��ԂC�R8��
��km[�WŴ#��"���@ ���{P���R�� (59| �Qc��2N���vO�3� C�娴J�N����\0��|`�[~+.Z&� H%~�i91D X��VS���j0@d	1	�Ȅ>Հ���Q$ @!P��
���'1��<����_�����} �a㺰W�5 ��hU�(�T>�	 ]���_>� ��´Ļ$� `�/P�� �.�C~o0 1�Q�]�� ��4M��#�<S-�U���� &%Fsa8�S
"��t�=(�[�c�{:��1��0y��d��QA��! �C�3��%[��V�K�M�T�(��0͆��e�hP B�W������!����UtC����'A�X ����h�� �vr� Xk_3s�� �+��cn� �̠����T2����J0��ӈ�b��`n�� r���:�� �K�H�P ��b|NB >�L-I�~K�MG�k���� �eJ������3 *�zSK�� ��xV�&��"(d}���_�Y' �Ӹ�!�� �����U(%�P@�q1��^s� ��
��� �H�%�n �	)̓�� ��*ؑ�����Կ ���� wz�]hg ��q�� ��S���0\�� �mh�%�����!�3��H �lk��	�����@��3p ��4 �����"��������x�������y�����.� ��:���� +Uֻ5� ���b�s�� ����� �� 4�$H���(؈0��u��j� !� �_�5��4)����e�S��1�\`�� %����Y� 8��!\� s��iN�X� �_��x-B} w���;��\$�T� a���� ��^)� v� Ϣ�#�Y6� �!�-b.a l��� �Z�`	� ��#��o����G�	� ���I���~J���
� �t�_�!]{* +���2� Ȁh%c�� -�N�r�~�S~�T^��< *�:���PhB�%.(�� +�A��!��@��X[{�{S�8�!��"� ����)^�� ��t�[b� 2�Q}TD�o (�1���� �R���� �!�_�O 2?]T�d��šǎ>s�1�:�.��/�P��� �J��D� A�S��� ����< P(Ƹ8/� �H5,D\�Z	����~�&  R�a[�*��X�|�eC��,� ���⠮� [�0�W�� �.2 X�9��*�H�R�;� ���Ji� ��C����3����� ���2o,x R$fQOF� ����1�� ���s[_���� ,Q���٘ 2�����o� v���:��� �Sf!ڐ�dZހ#�+� ��](��r �������iԠ��p�: X0��� �<I�����ӊ����� �\���O� �����(�X� ���'0��^��U2�]���z�,(�o?\��� �-���O �J[�`�h5 E�k��� Y*��.� �>��<0�k��;�� ��Y� 7�1�!� Rݶ��)��	b��\��fP�08�"�����Sܳ7��:{��� ߆Y �d) ��\;	�ŏ�T^������	u͠�]�~ ��>h(�ր�5�z�
�T*��90W ��@)1��E,�;.���{_���j��� �L��* F�с��Q�� B�V �_�N ��9��b 1���@�˰���Y���%� _��bj��t� ���K�� �@l SR��N�zr �	�^�� Z�����X�����`��%EK��`� �e���z��	��� r��<��͸�����q V�:�@�;4K�J�3_�[ }H��P�� �e����"��t��@�⮅�� A�飊,-��� @���Z#ˤ���R �Ȳ� �$c 5������ n���!Ȼ� �l�~�D%8:�=� '¶�P�� ���_U��� W�2�9�h �!����[ �S�1��f��X���oDJ§���\��� y��� ��3=��� �§�K�} n���
��O��ஞ-A� �HT~��� �&�2�\֔���~�紝���0���^v@	� ��`���O0 ���(5�9uf&~ �&I}� �ؿ춝 ��,�Z�h �9o/	�R��:�{�u�� O�DbqB	Y4�@�+�U ����� ʆ�8f�, 	���# �n�O���� ��P�KU ��/���	h=�]���_ � ��� ���1�>ꀀ��C4�_g&��� �&Ԇ?� i`p�k�F _o���� ^��4XZQ�8, �Ο�Ab��� 1ƾ�9� �3J*�Y� -�O	bl�� ��/��\�N�E�@�� )���a*��Z7LF`���� �)^A�KE ���J([��~D\�n �4Q�޹WČ
��	�O���� �( �Q%�@	2w� �r�Oֺ5 �]�_��y��� ���U�`�m4�O��gP�l�(�����wc��� : ]�ü{�� 
��0E�Cu�/�+d5T�~��Z8�
���� @�~%K �a��V��f~�?� 2�Y��O��oq_��l�N������L��/��q��Yz	\�B"Vǥ�����=�%�=��]�� g&H0��՘	�� ��49$f���O����!@��} L-C�;щy|Q un�~���T��`a1���ZJ��i�8 ڰ���{�8� �ї����K���=� i�-�ӆ.�� �	z����a |�}U��Ÿ1.1� :��GH�V�hmU����R_������� Z���� �?./�e���w��h�xN9�3�!Ő�&tU���rp�L_VXY��`P&�^� t˽ZzW�,�M� N�j�
��9	ʁ��^��(h	-�>f�@����T C0�_�v�㲺 RxO*"I �}b%W�P �F	�!.X�� 0�g_
� '���.n���0�}� �$�%��� �Xt�"�� N��#�Z� �]��� ��n�$�q ���k�
h	�Y�a ��PJ r���X "�Y�h��( ^�	Q��$��5Sn=�2���\3� E�1ڙK;�4N`P܁S�u�X��8} \h��tIV5�	����>�� �@L]��,��0�S(Н�6.�R~�X>��a��W:1��Q��h�L [2ր���H�W ��� 1]sE X���K��:"!�����t �A�ve�%� �\c�� ZIAƫ�v��� ?��n[� Z����R&�
  9�hv*�!O�����0�>W)�a׀!6z��h ���$(�} �pv�\O�� iV��@�s͔����\;� 9������24}~�|�A�@^�F��� [�Hk�� ����o��� i�ـ&XR ���|��?`C�w�L�R  㮷�Y�/?�� M�g	�$ �`��0�� 3�¸q ���C���W��T+�_���� �Ղ�֡�H�z ?��G��' �ɑ���* �è��0U �d]�۠�� s�jM�Y,�8
� 5�$ps��7����� 0��Ց�@Q�B$n?`��1 �]��؃�� �������s� ��Z�-� |��� /H��f!� �nBZ0 *^�aԱz��,C� #��"�
TZ��� �^:�?� {D&WK� �z�Q���� ��y��p�? ��]8M��Z �P�G� ��d���Լ_ ��%���Z=1 �UT�E�� \)�:���Qv���@�� E`�	,���&8p<���( ��#�!�� �맶�>��[�a8x�W�u{^��i�[�`�`=W� T"��qM ���y� *�@>�^ ����� oz�	�J!��ނ*� ���K����r� З�}�H�����>��$�Ǉ���c )����0 �đ��f�p� � �S���y� �F��>������~��7Pd��/�8����&+��$[� ]��Z� ���1r?��� ���ˠ��� WQ���pN �񋂉��j5~�l?��2 ��z�e�B �k1�ab��Y�=��]|'���� bTӎ{0SE(N�Z,֠�9��� ���sPzD �Kɢ��� !����Xh_�^�f������Fw ��X)Ғ �:�����E�u����C��*�A|k�� �� !�iDft`a~MvY�\�� �!�ҕ~�H��;�:J 6����&� 2Z�pX}B ���~�*� <�-���&�1 ��������g�+�.���`ᣍf=� �Z��0	� 
�[��h� �zB'�~}a ��n�u�3i ����N W|-p�H �;#O�ٌ �t?�"�� ��X�O�� +��{ԝ�C ��Tx��ٟ �~�� ����UE����\�.���%?�� m��� �^�4���])	��` �9 BlW��]^� �Jf��/�R �-Z�=�� [V���3��H�� ��\PQ� S��(���	��Աݿ Dc��8LqK �`�Q�� �g�)6{W\�Aqv+`�1h����TR� *����P����@+͝�8�5���ɠ�U� �L|�P~ȿ8_�!����ɗ }�9z ���S�Z� f�A�36�/ꐀF1Z	� eٰ/��%�z? ���my� �-Q~�	8% �R�gj�U�h i�*���e����l
� �4aʹX� zr�`C ���k�2[ 0I���t�p���=�� ��S���b *���f)� A؅1мD S��n�Ӑx "b�_N�HeR�Zu�r��� 
���?�����F�9P�0\� a����J�R�����@�鵈 ��?	��~ +Y"n�'�uU \hW���; � LA�	R���֋��~��W���^ P�*��� 40H���E� ��A�U�<	 Z�)V�� [���dO�.Z ��W8-#x� ��β��j\eR��� �:�� �f�	YR�EB9��M��2� ]��*��v �(M��� G�B��� +^��e�D3����Y� �t�$Z�	�ox�����Mh0�J�/0 � >��A�� \���� ��wJ����4�$o�m�+[��@���S� D����'4 ���آ . g�X���"��/J 1�_!��)����3b�踔�1}[�^S+ۉN��\� �ū$�9b ���.��"� 72�{帬�9$) Y�hI=�A�R`���t !�[�Z��8q���� ���[
�ʒS�� ��=,j��䮽���/@� �W�����ӻ�����?�A���'Zh�H F
Ž�$�<�-� �+uP m��'�8 ҃�>c騫 �-)�U�� �}1R� ���*��� �VY�!H� ��"^h+����K���� F�Z_�"E0$V`� �seS� a�7ޭ���?(! fy1�@�+6�B3�O�`/���� Q
��h��^pj�z6 ���R V1��/�= �Ĝ�ذk�y|��h������� ��vNf	 �`̀�o�n������[��X\q �6���W Gw�e�?a��`	� Z&�6�?�,Ef @6~ P�pN� ���d � `����:QL�E �Yz��U }���9k'�]��1h�6�����ڭ��p�~za�E� �� �GXt� �[�c@�(��� �ݺ�N��	#���[ ����qkǵ8�Y ��h$3+ ibܔ"	1�t5���hUyE �%�o<���f&ޢl���g]� �� H	0�_�����^��8��J�O�. +��un��`X2���] �!�Q��w�N
�(���c�b �e<?t1�P�9 L�3e[�>��}0�o�� ؾ�v9�) ��"���d x����X�1 FpI��4� j�ځ�[e�{�B'�`�)�-�0����.� ٧{��J����h�ؗ�Pt�&�l��Z�n �)�[��h ��*�V��\k� �-�W�R[�y)GE����Z�� i1������O^)��8(�_ ��K�0�2� �';�a��~��YZU��dc] I��E�v�  ���*� \�<'�u )��OK�� �p��9����n_@+	� A���T�� 0�,�b��	��1������� ����T O�@0��5�f�-��S�y����~�}Q�v��@��aW+�Cj0���?<��3h�'�p�Q ���ƹK� �+�	�/���N�o�!�#�� n�.�ۃ Ѵ?	$�wlL! ���0ֺ yK#���2�L\���'E@̲U醘����_���ѧ ���4B!��S ��J�b��P ���	7 �D�)� PV��aS�0 z��$^� ��&�Ej�[�z	 ���Iqb `��%�
��^�:]�<�y ї1�0�xb��]a�� �D��E\C*;��\' �JH� ��d63� ̳�X �h sQ���T�f���)��nIi� �#}{eKW<�$v5 ��u� :쿲P��C.�0� �U !�&fk� �$BK�� (�>���w������z��?�&��@���)� wD��`$ ������� %w�8�lI /�,r -sC ⒉�Y: W�X��f
 �L�/�| �8��� �2�@���,�Y s*��`� ݁��eX������H�h��� �R�Y��g ��+ ����r����^]��	��uw���N�x����_��^
��R�ѽ�H ǹ��B�� ?���pk�H( RFh��!��TX-�4��1�V �q��gY�tHI���a�;~�4����S�8��^K����ȕ�ࡅj;言D ��I)$[�	����Kx_� U���pa|�O3 \��vD%�0�Q�'02�*��}r��B	\���6��J��x5'�`�QT�*�p?�~ [ �8UN� (�r�݈� ����+�`�sF�h�p��� ��^Y��0x�}� Ɖ�"��,� �|����<`O@���N�<8Zs �-�gj%_�$�)�|w���ck��2� 
�Y�I߂@ �l0�C��s#�! P�%˧��� ^�Q� , J����� ���	P
 ]qɅf� 1Y�(�!^��<C����?� �[h�;�>������qN �+0S�HG� V#������ �;^��	���}g���q4�� K|��.�P�d�������Z��t�mD�1+$ٮ�OŹ���u( �;���������a����TR����>� ���\��  �ڧ��dXt<0��I���+�N(�@0��,Ҟ�DP�͸;�-�3ǁ�� Q��+�O��X
� !0n��)x� $�L�i] �:~��/\Ip̎
��ߕ���J�A� ��/�ِ[ ,��j�$\@	��cpE��N� ���}�L����g��kn� �Z�"�����Q�����0 f}���) �| �~= R����FLd��� 8b�t	*)#�:4��_ �߿�+�� E���K)O�=��h�|��Q zC���.E�] ��� ı-(�K��LN�" ��X���� \� �b�h �՘��^J �HF�Q��L ��5���� %9We�N� (}G�d
,X�m@���ZV �	�ި� ������ɯ�&�M��')� ;ň�����&�X�BQ�� *��a��Z�
)�Y�@i.�0�#���~� �HVC ��X�b� 8�y��+R �����'� ʷL�� ��l[��h $�|`�q١�Q%��}	 ��Y�>����� DB0���#c���p�� ����4~ xn�;D�1 ��@6,PA %l�E��/����v���O���Z9��g=����*�hnؘ�U�'!��" ����K���Y����P�^ fXg��IZ����-�v�t $
��[���� 3Br�<�6��& � �D��1 �b��+.�%��{����) �PKzh� ˃	X�@�%��?���9)��t��d�j� ;!��8@ɧDo�"��]�|I /���&�1_�4�� ��]$�< �F ��k�x �d[��s�.��p��a 3
�Αj�} �@�hJ�� ����W)�u ��~㆕Tt\�t ��*�� Wu��n�N}|� ���h�;�� !�o�X4�c,�Y�  ��	J��� ���W0 �P6�1o�� �]V����$�� `�R'u ���Ų� ��\US38 �Q(��k ���*�SP �4����(쒷��0 =�.���>3�U �K������@�\��H�E [)�`�:fh�|��#���K��^�/ �����J� &��M�\< X-�*�1�:�Z H�]�˄Y�� ��F��ؘ ����� ~�[�7�3��X8 �C �,FH#W� �(!Ȉ\[� ��O��a� ��(�c2N����[ ������rJ^����*����=���d�I �j�+ t����; �X K�0,'�vv `p��� ��}�r=� WFu�t~�Z�����H�V�� ��dhNj\+E������s ���C� ����$�^��Q�Q���]N �	��59��� �)�'���O Y� /����#Š$x�G���j<�XА� ����t�ݗ �)*�.�� �u�	�:� ��^b� ����X�5�(�� N�E70��&	G6 2�Νq� ֽ�(� 	�_�Uy �B�P�a� ��ܶK< ��L=�����N�� !��V �>���� �P%+�|� xh^�ZȎFO�'�p��Qo�b���-�)ABu`w��8��K���� ��^R�T��|��"	�S�������Ib9� )ź���;1Q �J[�	� sqB%��I� ���u�Z, (����::�́�5�[�t!j 
�WT� _�~���q�� �O2��!�"��ٜwB ���p��7m �`�D'�z���)���� K����V����H%��W�9\� u�B�k��� xT�|X�� ~�0t�R  ߵp
;۽� �~��]�P X��Z�	� �^MB�EPѰ�@͑O�g����� �½y�T] �(ۆ�I��Z	�Ա�
�WDP�� ���#٭� l��j����^ �:_ �РS �KᨺO�� ������� B����� &bAJ��c�' �j#�u�� s�a��� 1��X�8�Z���0S�~[+Π�&��L %�ף& '�Fhm�� �7\�ê� �Ww"�tQ�
ξD ����� ���0��X �2/���׍t� �*>�����Uf��W�?�� h�*c}�	�b���0�Q2�yn R�(�~Z �<��K���ɈD���м�ݐy |���_( ú�	���s� B�ö�����q�c�l�jΗ �&�������Op��
��� �[�9a@��h��20Z�D�~Q5 ������-� �C%����0��2
t�;�Bi�V� ����s�� ���b�v #�u��I� �N<�{���9�?��� +�(3�X�:����QC`E��G�� �
"^��~I������+�U� ��*��fR 0�@Q��� ����tr* � wP�n� g�{!1�o�a	]���� 'd���E^9���@/ ��a�x� +J� ��� y���HV� 3���:")�}���k�l��/vJ��P`� ������w����JA�ǹ�p�Z0���؉� 6�o��5�v�Hh��#�p��4r�7KCQ1¹��9^@T� �'aO�k�J ��!��\�$�C4�r����* �[�V��
W �3,��t��	)޻��X���h8�UT�z� p).��\;C��z���H7 �%�2�Q�>���(_ƂF�'�*q{A���.ĸ3 s(f�5a `��%�'� ���p��qOЇo�B:���� ��_��ec ը�A�%�2 U�ʸ�9Y֯�]#�J��R�� 2���	ف3 MT[S� .� �<��HR "��Ÿ @K����y��� ukL�q.� �-������J�:���N��4�+�_�j ��(U�Ҟ �<B��� �JǇ�P;+ � X��R���(,���pjF /�0��-�_�S�	����7 j�
���� p��T�XQ ����*�k
Y�����ow� ��p�� ���R��� h���1e �'��9�z�� �|�)�GH ^�b$c�����V� �s��#� P2ɸ��� ���t��  ̀�s�ëy���S�w��0D�$R0d� _h脝ܰ �	��\�[ ��`@�Ly��A�� � �N������ �*�T�X�� ��t"	�]( �� >P����32��``[T 
�p��_� +�*�ʀ�� �	�m&�� �h_�Kx3Ź�@A���v 7����0�I�e����rn< 1�/h��4Kq� �Q�>�+^� �5�!�B� ?iQlK� h'@C��o�� ��$u}B&�P@�� �y�HU�>zה�� �+h�� ���<4?%xA1���p<{w����a_��,/ ���� G����;�Qs��� �2�V����ka��I	Q����V�h�jd� A��Tѝ�0U(N�%��]�} ���p� SPN�W��&�<M )�_aR5���+�Ii�ɉ3�h���x����`�TQ�� w���Y�-����Uv��*8�:�b�� ���1�"@`]��!�2� _y*	VF�|����@�u� ��"�_�- 'T�B!DAP�k��@c���-M �d
%�L�� �q��'>s�h4��V ���|R�� �@�XhL Uø� �l���� �1*BGΐz ����P�, _DF�Z�bN �r7�}� +¾��%�A ��`�zw7 ^3��F�& �"Y�� Sp���8h� ���x �6����w[ �f#�H}� J�!�4E���6���vbq0��$���e�K�օ����<�� ހ��� b���R�%�/"�a �*�?^Y����m�A�N0� ��U�&��~����\���n� MO���� �FYf��v, ����%>/�S�
`������I@؋�5>
� �� �~�XJ �v�?��. ���(��-J ��h�����n�x%���y� �vLp�P '}�0�u�� ��3
Z��X�� ���#��e���� ��0�� �Y�D�� '��
o��< �!R��"��@����9U�j'*�_�R�ri�ƐT�O#�H '�+�.��. ��vK�h|��U'����� �pPeq��₾�m^\�� V���'� �t1�(��,̬� ��Z�,���tK�YhX-I��*>���\#���vPr2���/.�N4�q~����"2�
�0(�[��W��w����!-�^�&����	�`� �}<= (й$Ȉ ԉϠ�;	� _ܓ��$2�hu-����V�����
���.�6�
�+�f�	��O p����\2K �#���Z9��������|����� �WA�n�0½��S��h �dJߦ� 1�Y��Λ:^��E��h�5 �L�BT��M� oP`�� }����Iz� �K]J��� )��0��� 	-"ͣ�!� ���0� q/�ae���� ����_!� 28�]%΋B W�MS���1��lX��	�%���zǣ/�� 	̓� T�#8�� �)tmPV�* hj�3?C� ���-��� �>�:�o~A!����� �=�k	�Q�� �9�� �K6�!ʽ������5�"�R�'��h�} �,#��1� ��&��4 <�-����:�ځ���������6�?$0��`�r��� ���&ژ\	 ��(��r��5O�� f�y�� �r^A�s� �7��]��%�{ @��l3 ہ��r� nӜ�EUѽ��Dg���y��< >�F7��V|�����	���RK���O ��vU�f��� ���xp%� `�U�6�� �O	���]�=�.�� \l%�� q�g��`� ���]�h+ YL�����_��[���b��E� }�y�����m��_ �1K� �x����YZ��]��p�$9h2�R�%������[�B��\S~��� ��b�� �q[ =���an��@��� EF���?� eyٲO���u� ���
�\� �HN$�I��� *�Q��o�� �=Ӓ�[ߨtO�h -�Gq��� �����3h\b�R�`� V	t<`  *������Z��+��]� X��% !4���/ �F<&��j T0�� V�h�tW\ ^�(��ۇ ���4	�� ����,Z(2��o���P �A���� �.�X��+`iS����Y/  �T�a��P� �L��O����W�0*��Η|fb����--��wo ħ��O���'d� �$���X��Q�o���!g 	1�D�%�bJ�W�`2  <�O���+�9R- ������9	*�	.�����O nG�Ј���]F	%߬�
��(� >1��w ��^���W ��;��?_O��+��5�n� ��h�R ����FL� �	H������Qha�ٵx` R
�$�r �0oSKF}� ��?����.A�� ob���_QI �>H!��ȩu�u�v�����!�8�[W0�(��0B� �S��߹��*�8(�_`��Z�S�1�&��0�| �/-F�s ���J�?8 �'�~��	�TA�ޠt"� ��p�IZ����'���9���4�g�jR���_T� �ถh1Yf��_����� ���p|Е>�s�w�Y �X��o�>��j%ܨp� ,[Z�g�d	 �=f!�U  �W�ٿw�,�O_@~��W�  �U��?�=#�}���0ʈ��0�� �)�PY� ^�]�i� �s�,J�5 ��b{�p �h�E2>S$wq� y���i���A0��@��� �Y�K��O� �c�A�m E�.D_�Z�� V��$�S�� ����@p �
w8��h�<Npk��@��b p˝�U6�va��o��L�@� g�hi� �_�n1w`�B���0�Ǘ� yÅ��Z��:�! _�4H��� )k y���-	o� ?*�|�x��H�:`J�A� ��i�� �}�gBH5�̀��֛ W�Sk����&��� �Y�{�� _r�HS�/�]���!`(\[ �M8���� 2
)�ZS� ɿ��� j����� �cq���2���H��VZ��BoƦ�B�� $����=�^�.���X�n �t�ҁ��p>�Ȭ��m) ���[�ƌ �V"վ�/��w ���3��� ׺lu�@� 0߷����� 
��XP��� �;]+ʆ QF2�U\Z� qv֖�+� �ה�k��1 Ҍ�(SfR� {K
��E� ӹ�� �����[�yZ�&�.r� R:����&�� n2����3ƚ�� �9��{� ���hO^M�� '��ua| � ���J �*@�	�Q=�ĺ���-p [�.��TFvE �
'	�g�2<� �N��G���1� ���h�s$ #�D�<� �v���{��!�-��`>��pN�_�M@4�J 5�̇#�,a���	 "p�� ���7Ps� o�O
@~A�x� ��sKB׿��C`L��N,� `dǻ���� ��u�:�� <�[=�-�$ /ʢ����9!����%9���`Liڒ���4� �2]�R~\�K.�� �ք`�=�!�$��OBz��v�^���Vz��� ��n����T ��^e��_( ��w9���� �z#�Xh;j��-UB�]��p7v�w� ���I٫�� ��;�G� \�J�]aV *��TW�z^ j�D��'���!n�ۉ8��Z� g���∐v ����;�LY��V�n� ��&P# �tA��-� �Y���ˠ6?(� X.
DN?����4֑��j&�� 0S��H�� 1�h�(˖� �-����"� ��'��5 2,���Z ��[	Ϲ*���ha������`�3Y�������PA�����41�7\���� T���|Þ >��+Oe?� �Y��)�6.����� o>�� ҽ��(&��	 K��Q;g �گ5v�@� �R)к �
?	��3��*" ���;��p ��
�(/N!� �ϐ� D��j�8Ã ��0د������2P^�� �S)�P�� �?��Wl� 0�\)�(�� � �p
 �Z=�|��S V�s�%�� ^�LޫK� �����>� �����Uo�@�ɫ��&�J $!Gx\	��(W����8ň�\v�����K>O� B��5���	�����$" �Z�,�+�R C��_ֿ ���б� ������i g��f�����0�u�)��BV�� [^	N�� i�z����( �\�{��y� ��6
�ſ� �k�A��K`X�� *j<G)�[ Y}����2I�F�]b���u�q��G����ͩ_��V�16�`��z��^�)@Ҝ �0Ӫd� 
���� �OQW�6"[.�� !���Ў2 ��$M���{h |��p�>� �b5ρ� �
o����#:��Z��yW���(�杀a�� -��,�K9߱�X� _	��"5 �hY�A�f w[O��!�n��r��3� �:��HEy`2��#�a�����U ih�P��� �.H���� 9˷�7�� 8p�_� ��+B�^ �"@�YQ
 F����]x~ �t&J�'� �)M��G :7o�(�R�ؐ� �rp�q F
�B򏸘� 4?G(�X 2n� ��!t�7��S����@�L� 	�3��Nî��-���h^�(�@0�a`Y�sV0d ArI��� ��(4� ��ҁ�ף ��e�9ڸ�w	 Q�����$�Ys�l ���Q�pk� �P��Lb�r U/`��B	�+����j�/A1�ZךY� x!�3�]' �%�?�	 /��8� �F4��2<�����3�
�č�/�t� A���| ���
�� )�Ë �.{P�Q����$\�k S�~"A�?��`Gό7��+ڡ��@����F���-"�WL� �q���>ԐP8�@ �z
�t�� �ļk��5�Qh �)�� ��&�Xb`h-���p2� ]�A���^ �Y��
��*�zJ�����"� �c����  1/��� �<CY���������d�}�ۃ��X 
4�Wipl 2�)Ѹ��� Z��:re�/�K����2V*��?R��I� 8�u����� ���N��ҩ �r�%�X���	w c�+�� ��|����[ �w͞$3 �RS���6 ^��E�qu�h��_:�� �UT��3V=N� 5�� � �޵�!-���P(9�t� [/XR!��U% a�e�,�V_ B�偘 H�d��Ac �U���!�P��� 
aWY��i.M| T�X� �(��A Z��Bzd� _�*'|>� �ے��� ;y�p���� J1�@X�9 �m�"�L �|_���� 3{����'� TQPh�\@ H���-�7 5�W9�<1;!���4X� Z���5 ]��ÕQ�� D:�m#� �]����;ס��W�n�� ٿ�HX>���|i ��5y�&@��Ѐ��t�Q -��jXZ�� ���t��e�$� �4y�� !2��Ţ �@	ɕ�u� �Z��
�����I�vDb�4�ZO��P� *���ʤ� �JR�xz�! ��P_�q5 ��{H��� 㜩U.� r��O1�ߐ �S���M ���$1?� �3�
�60>P$f1�I�,��#X� 	�q�]�{� �$!Z*Ϗ;;���v ����v�	�Tݐ sd�j� _b�]ޱ�� ��-W0� ���
� �V־	  ܪ����y'8N� �Tǿ�A��) �U@��cg� 7���' ����]� �~AUL<�q�
��}!b��e�@^> c��ui�
 �?�;�� :�]��B��<�� ��!'�Zu �%�2� 
ސ|a�� �*[�o�w��h�l^�И�� �!鶆f�<��Y�/~�� ����u�������������䂍���_�5� 
 0�Zh ��*�I 1������ q`��[ �W �P�af	F\�" ��)��`>»���w�}M��q �k_)WU�����.� Z��R" ��t��-j ��OQ�f:)�+؎R- P���XB� r�^��Q���	�:J �����\0 ��'�<�( PY�H�^��)g����� ��	#��q H2��Ss �1{�>o��8%OA��$J��d	�<�O`}z`H_� ����H7%�8@ӝ��!��`jEO ���� _+�bX� �@�����p�� �fS0��� N�Έ٫q�w���X�,.��B ���ق�dETlIs���� )��y}�#� V�ά�� l�Z��$;�.�Ƞ 9�&\h�`��ҿ�p^� x<P�������8��vX�1	�Q �[P��>Va?���� ���i
��@����h Lbc��T ��k�P��p��v������X���AI� �� �oB�G|�w t���) ����z��ٽ��'	R��W�?���!��AԶ �4�Sz���: �������]_���� ��\كb��3B� 1_f�)
�ʹ�\Yu� ����i���Z�`Wu �"GQĿ�� ����|OV$����X �[�H�a/�Y`�:�
ZW�c�S�����1"� �% M�J�Ȑ*�QA�D��a��F�	J�2��t�8 ���_1���0 ҄� ed��2�i�>1�^ǂ��J� �0�S
��*�Z �Ra���>�V���O��R�� ��� %	�p�U> �=�J��h� 9���X�� U������92݀��<�0��n� ��޵G�u-�) 7ô�� :�b7 /p�U ;�R�&�� ��?t~ ���]J� #UyϘïiH� kh�2? �����Q-����� U%/� b���TZ�鰉Q����@o�-r�� �L��H�C)Ͱw�h�0����%Vv���H0 �!~�-hj ��	p,�`: ��*��0,�wF �)�hSH�<����u
R�� ������� ��b+#�t ��X�דCH\Њ �࿞b; ��a*Ӂ- 0�G+͈M 3	ɌĚ_ ��b���[ ��F��XR )���}'���hMӀ �_�d ^����P��<*L��)$�] |S�P��	&���e k��R ��@ A�Z�?�� a0{��"� �GR �	� ��1� ��/��ע� ��y?�W* ����>����_<����[�x�V4�
�Õf�� d�e	K)b� c��%�oׂ� ��[��J
� �O~r>|%'_��Z�9��� �]� o2 ����c
���/�[ʭ��� ���^�"�7 �	�+�� �ڐw��?�P�|Sd�N�"��9ࠀ���զ�[���)���(��#�0�T�����U� �7��-��� �X��z�@��\r �p�ض X��=6`���ǜ�����!�/ �si`,�#��V�ɨ�� ��Y�>� P�c���À� �[<�
�h��	1���m�E�װ�����Fzl ��L6wSX(j �ԋ��0|X]K ��D��� ��$2ѩ�x�� ���?�X� �R��� }@�ã���(��[��Rڎ C	�J@|� P����_Z �jB���;; ��{K���_k�M��;,gΈ �+�K3�cN�?A_�ho�d'����%\N�# _́����J ��Rrb��0_�����	 �Z`f���� >�<�K�@ i/Aڹ�S ����� ��!b��  �3L��.z?��6l�4ǁ���ɉ���_��~�$�� 1+[� �X�xfZS0 ݝ^�k� �\�؀��hX)@ f��A,
+�6[���K9���ȳ�j�s\�hVi ��悡	a b^�!v0��j �1�	�W�;� �+�R�8�� 鷒��a "N-v�� �c\d�&X! ��_z��L,�?��R1٘� _|��!;� ߃�O��� �4iڨ��� �ZY
���� ��	��j�X�1���{h pV����: ��◬d�3��Ti~�v�%� X��N� Y���<-p����h�"� 
�R��D B���`O1���9���G�� �V 7�# F��y��C�Ѡ�p5� �v�P��� _\�}��`� ȗ�n��.��"���ՒtI ��p�� �P����R����$�X��]�P( T��-�j� h���$V l ��^�D� �_��L[� �ho^l{�?���
� ���_ N�J�/UKa��� 8B�[��^&���h`�.��L� �.�t� ^é�����&�� <�Q��A8������x� ��L�r�b� ����.f!��v
�|����LMX�/�������v2a��� �0��[��챶�	Z}�uC=�S������ ��Q�2j�Yk��A�«� �3P٭�� ��U~&2zZ ����r[  ��+U�j �ѻ�C�s� ��
E��k ����j�f|;L&H{ Ai{�?넘� ���M��.ՓV��}^��D�$=����h��1� �PO�`M�� �' �U�ƚS������!��A� *�k�]��.�C�� ��zat� �@#��� N��q`� ��0����X�*+ �	-��mDp1���̯�]{�&�� ���0o�E�I���Q���|ԓ �S:��V� �����y Z���J��\ ����!�~��2�� ��we˦M:_y�ԝx�	����"�� G�{ XY��, �
_��Ư��u��S����@� < �����b? �|�(��Z1�I�O�ȩ� �J��g�_�8�0�H�xr �fX  ڀ�*�V���` �)͇���/��hX0�-v� I[��|9� ��`T�Y �0��$���=(��0����]�%�u��s �D	���� �Y��l�& �7B�qU���|A s!9?��~ O�c�y@]j���"[�>�,韀�0�m �=I	�x D�ܐE�1 Ĭ��pȷ [ۺZ��P�Ζ���)_��G� R(貞������ F�S�
�u�  I}x˳U f>�ӷ�!��ƀ1��%�/��K���N a�"��Y� ^�<�!I{� n�r�N��49t�k���"� ������� �U2۽� b��(�T5 ��~���! �:���"� �5�Q0f ��I�&����b@D�0��$Z ���Ü���E�����_��	�� �W�B�����p<��%}�7�̕v�<*[���� ���X(��� �\��{� �Q���� �-�� Cu$D�b�3, �u��}2@ �L�&�� ��ݟ����12�W��* �0c��'��f��
� F��:qՉ����;U�����j`��/�	^ e�1�+.�Z�t� ����:B~ .�X{}>n���1� oT�NgO`>9��ck#�Y DX^�%S]�?`���}	���� ����@����S��l�X�ҠKeg �AE�b�Z�:�Ā­���Ǟ��?�O����<� 	�v��� �oO���� q� 0��#Mݭe�W��wn�y맳���# Z�Qd(���3 �1)��lNY E�b��Vݑ9�iL??��\:��(_ϼ
��2[�t#�H ��Kܢp� P0��� �B�Ӏ���t �]����	�/ޔ�?), 3�G���� ��	�`C�ZW�Bs��hv�S/��U��K �A�2*�� ��Z��� >�V�0 ����yz�ju� �ǀ�2� �`h"q(� ��A��F[ ����O/0� a:�R��vf���Z��P�g`��X �AU	� ��i�f{$:(� ȢP�� ��>���- �x4���~P��	_��y� ��Oa�\D$���p{����x* h�tl��(HQz Hz�S&��p1�I��n ԙj=N %�r���� 騲^� e-EU���� h�]��A$?�����D��{ �9�Q<%�� �\�����x!�Cy �"��K �d�\VaJ ��TY�+�]>���%Bzf	.1�:�-|��9�t����4�u	�� �� o�c�)ˈ �'Y%��u �\@�hK�\(� }:�<�[ �dk���N�����è9 4��4�h�6 �_�H��M ADX
p�( ܺ	3;��Z�l�D��Ǘ��M>
��݀ ��[��JK W����h �o��`�s{8b��a�*/�E����� l�X>�k� v-��;|$D�#����}���$����0�⠎���� �q[	��� nU�y��Y�X�� D?-�u �D���x]�b"3\�=�w*P�;�G��.�? 
��o���&�! �	ݾCʽ� �2j]�	�CЙ�. �>��F!
vs� � SR�h�[7#���B, ���T�Y ��JZS(�sa�@ho�.��" �����%k�)&8���g� e������U y���R*� ��9�7� f�v�i��RK?�
��kᘘ �C�4%���y������( �d�)�DZ8уc���H�8� 3eS�M$�+ /��*��( ۸�: �� -�
T�LC�I�BZ+����� ���Y� ���'�е�vD �v	�� @A�0"(� ���sV� �� �)$б��8@6�_�=X�3�JڮTNxA ���(��:���؝Yu�O�9/���р1LNp"�pYF�Z /U-�Q	C;ҏ̳ F�3�XB ���x)�� V��[�Sީ �	IqUe ,)|��� v�[��� VP�<��(� 8{�^Ƽ��p=hl�'~�d�\ ��b�K�^Θ�� ��&�R��<q/�������."�i~��xI�+�����O��=ËX ���:B��A4��� P� ��`\���q�� D-�7#ׄ4 ��nF2:t& XZOߧ�šU��� ���%�a{+�'�`�v,	�8�y`V� $�����P� �h/�Z�VÅ�[����"D�0�q� �E=�N�n v����� ���>[Y�xsm@1䒹*X# %�|@E�� c�kW /h �1���܌� .��^��# ��+�aZ�4>Fn�`�@0��x�EX�	� �-nMD2 ���/��q��1 �]*��>-i�8������m#K� O��z%�h� Tۗ�DB��Z�%3�E�	 ��v&˧_ ��8�T �f}�d�V���- ��0��:k c(��A� /�B�.h �N)�j��� z�x���� ���^ݱ�o *�#T! �c�Ί�GQ�b���$ ��q� 4߃
H ׀�Ij��"'������� ])�鮠����l�@u�x�f h@B�֖�
��^P�0�� k��_���Q/<}p���� ,�#e�(��� h�6��.��� ��V5[�� ��χI� �������+�΃��b\d �Q���wA? t1А�'���F �e4�ȴ��P 6�[��^,� �yD!W��}>A< ��\(� �	S��T8�c��[���]�飾}Xm� A�{PSV�' �P����� 9������ 7n�#�rk ��(S�g �8�M0�� #,o=��� ���a�C����<8W��-����;����h� 2&���۴ ���N\�g� h�i+!�_��%�^=���U� ��'R2� �A��bj�� Vf12���>�� їKk�������q�� �Z��j	���w�Ƚ��;�� ����l&[:�8��v�g¿(�� R%Xh̶� ������ �)��X�;J �f���%ԻY�p �;��-��F�afS�U�/���?]�v 0� nc���%��_U@��� �
����� �����g��X0n~@\�9�� ���<6� �Ժ�_ݨ� �qF��"=�C>u ��~30�5�y݉�����]8�(ƀ̘@�_&��1����b����T�����H�� �=!��Bv�{���P�� 4wl�
������~�r�	�F���S�����J���;�O��:}�`0�F �P߽x9I�V�L� 4qπO�X9PȂ Iک�Na .u�@��r �4bh��� Z [Ϻ!�� ����<R �B�_T��4=Q����Ne����	Y8������{�d]�`��! �"J��X h��3�ULN4��>���������@;�*�Z ��Q�:SP�\ ���!�n Б)'���ِ ����qC �X��u�	H�1a +U�.G� �*�0n! �1���͐ ���6���� O�-�B8_ #YA:���� *&"7'b� �3(~�� e�_��0�
a�}��9� d���<v_b ��\+ٚ4/	�Cce�i�� �Ѱ�.D (�X+� y�na���s� �D@%��s� �SWu0H���|@��Z�a���<�@��'S e��\aB��ܼ ��~Ҿ� ���;P" �]����V ���_S�e 0��Μ��:h���	�}ilL�� ;��p�� ��9^-"\�f �G]B���K����u^1 ��-ⵂ�� F �X�	�5�������/ "��p�@��1XH��U��N J�n9P�/��t�AA��VizH� �L� 	 ݈ϋ0�� ���\��� � V���R �����������w1l e�i� a �	��w��= ������� �"R�: v�&{���>�t����*� �m�A�� ��X/��b F��kt]�K��6M^��F�O�n�@�p���=J�� ǉ2�|������J�_�L-@n��\�[����2@�!�n�<[�,�*�ZRq^���T!��G_7�-���S ń�4G�&~�� �R3)���� 1^ѻ� ���+QW�r .b
�DM�0 ��;aS	��6�� �@I��t��[����Y1<'ڀ�2Z���b������+� � 5����$:��	�� s�b��&�8 Z�h/m���_|������ �S����Qrw��̐1����ZYP���CM&/��r0 �͕��{�����������29 ����Đ,0ȅh��ƾ�O�������Qp���� �Ux+� �	׺�t/ �1u�Pb� `%�N��&X��'���ݬ E�#��	�]�+ �%h�,�) ҉��}��� �?�CԾ� ���!g��Ր� �@�1�� ��Hj"ۓ�X�`�� ���,4a�p"��'0 ����hj �ɜ,���"�}�{�� �ﮢx	h �_�<7v'�0�* �Z1���@\(� Ö�Qe� k�F�>�� ��[�Z�5� ���W�m �e�24�(胫�:�|��� �N{��!u� ��2Ւ@� V� �����\� �A���"S� l�v-dW6����7�8�w� %������ ��6��� H5���4 \ �����`����2����	�8 *�{�u��}_;р��Q�V -��C� ����)�0 :�k��� 'e��*� �ź�U	X{� 	�NW�l��3���ѹA���x Ӻ�W�����Z%�`���B2ؠ,	3	ސ�Ӏ���U�>�W��K`h��� 7�$��E�� �*p��` mg �P �T��?Y� 7�m���Z ���_� �Lxyë�� h�~�&Y[��̥ /�>�f'2�u� an��
��� ��h�gE�L�` n-)��� {	xB��]���� 6�Ż���H%@�� Wˉ �Q1�Z��d ���%��]+ ��fi|�B �A5�k���� ~`ҽr: �DOf*%�G_���j��<� �� n�ͻ*R�� ����O���ꥢ%��� �^�u�r� |���=�s �z/$	�h\^� c��C0 ���z�o� �8%����Z�d4�f�ޠ�!� ������ Z�?P�A	���S�^Q�0� !��n*�� ��)�UY]�o��-����H1W�� >�@�#� _"jx� � ��J�w�{� �Lcvn�"2 ���G�%��r� �����å ��n��B[@AhR����P ���ȿ��0�3�Kh1�n�9뒀]�������X�&
�p�z ��`���(��X�h#`�y� u`��m�9�_x�<��B ��_ˬ����]�������b	� 9KPTXy# ӻ�;����K��vn0@�#��S�処�pD�����_�'<�/9
u;��V���W� ʥ�[�0� 2^b��6� 3�(���v ���w�/ %�3d$P�R���@ZV��|o1�� �`EW�B����	s]��x�.d ��X�+���2N�;
�0+ ]����B� Z!�T�c�� �h빻@H�L��4���#a �����RS+��������*<J ���-�� |h�x���yu �J��/V�Q��:��P$Еy� ���I_�# 	����� x\��Kf��u���D�4X�
v� _�䀅�� .���^�%9SpW Q�t��v�e �j	��� F��ƌ'�k�a��4 E�?+E��8�(��dF=�@��K�� �b)���ar 0���x�:� �>��Ұ�` OMI ���� iU�R��] ُ�Ha��v) ��
�>���eJ#��A| �18�*� �.D� �'_[`F�2�;)�����^{�v� *��,��y� ��u%X �bh��' ���)C`�� �\�{;�c ����H:+$ �ŗV퀄P ��DG��1 ����כ<� (����� �p3�GZ�x�F�����P� 3�(���6WUH �/i�1P��� �K��wAO%���e���� �	pǗ߸� �N\�~��_&��莩 �K��^�4� �����0���¡�	*��v ��b�:j1V@=�����z��]�� �eP^��&(�:�� �
�@i��) B}�⡽Wj l%ߔh�� 25�Qw@; ��Ye'	��h�������>y9 �
�5� '산#`1hYJ}�3�����6$)	�yh�I�!?��/�5��� ��n�֟�H����Jp���.�G� ���_�� ��O��e�� `���Z�	���l �	"��W������P ���L��K�� _����� : ��	�Z x�w�����s@> �<�,� ˈ�Y� �Вٕע� �G#�t�iH݅�2�	Q����� ��.X U(����]|� :���� \	�UE����T+����{L� �ɉ|*܎	�
� 0.o� h�l�@*� �8� a~'��G� 	��p��!���H]� 1�.�O/ n��$�� �&��hy ���
�_��a�:��� 쾗��Do��0�@�2� Sp�$�%>�<��� ~���9�!�K���Ȁ�?l� ����[� b/� ^f%]���^�� ���P*�5 ��Z��0� �!�_��q� T�͵E: �����4��$���:�ۡ3���@oy�E��=�7޸��� �ϴI[���'k�.�{���W 	�SL(�3н� ��]@ )_ �%N�WLC�g�z����9U�	��Q^0��X}�[ ��RD,�(H*���qA���W3א�P�����g����UG���V 6vR5zw�d�P�, Y�NC�O� {��A��yZY�!��.�p�/�,��%������r��| �dP+��&���t[��2���`�Ĉ3-}�	Z�r� ʹ\���� �����;1 @��i،u={��-ݔ�p/E ~0�	�Q�� *Z!�YA k�}D��e��]�M{7n�ź� ��"�1�Iم5 2�X�o 
�/7��%H����gK cY�-^* �L���'�:Ȱ }�^�N� ���1�fhC��9�g0�Yd�pX 2�S�ٻ�Z �0��)�	�RlϿ�!-Y�H��hI�
3�����\! ÅXQW� z?5���0;�~� fRQ��?� �7y��� ��!�0���1�@p,
}H��E /��j���˚�� ��(� ��4�� ��IR8f�yn���v�s�h �Jg�a�0��5 ^`7�"��c�dW�-��y� H�>�=��7@����\d�@�1� &PQU ��xH>�֡M���������a	� T���R9����24�	�!�z����ց�+�H��_�yF��؉��v� d���9�U� �S
���% Xt�����K�h.
�I�
c<~��9�ue�� w��@?�
 Q�0q�˻� *�hc��&(��N	�V �U��� `�:P��@c,���ȀO� ����߆�8� X �U2�Q~�K�a�SJ$'�
 �w2@? �/�Y.� b�A�)ŕ ~�XWU_� ���N�Z� @i�b���� �|V=��� @9!��L }&�t
�� I�6�[��,�i� �����j 
�h��0 �\�DY�K Bfw����	8�0 ZՆ� >�K�� ��"���45�H �0h�	�	S�u�8�3V�ˀ�f S�s���H��P �\�K�!)ݼ��&8�.w�P�*���1��%���2�L�Z* b> �BcX`�����O�Rq�T,��c`
谻( �������1 E+v^a���G%�����Ÿ�;�ݓ ��Q�� �kL7�0��XJ. @�{��`z �!�&�q �^ ��� ¤t�sU*� ��p<M�� ]@n߇���:9Y��?��� R���� W���s�ט��	x��<<�� � �ƊN��V;�`� ����!9{J���kr����3!A� Q��]��߾ {�,;Lo* >)a����: uQ�\/	g <�PU���[��s�~� �����O ��4/�=��٪�(��0���~�J Ւ��Yn� ��	hi$Qͮ �U�L� RX��h[u� ��U�(��� z;]ה ����~� �o���X$� ��)�9p�3Za/8�� �b�T�$	�0����'Ր�4��)( �B�h���M������ ��$!��@�"O� �������3���~�J�&D�%�M͠� K�ޅ�3�xr) ]'#R~qi�r�>�� D����	��h<@Hc��9�fpk ���b��J(�`�1)Y-
 �<�m6 ��l���n �����hP���.�Y� �?�0�� ��a'_Lu� �k@,~o���� c��i ����P��{ e�&�
�$�� J԰��K�u T24��������k��EWw ���pLRq>
0  ��Z2�P �	&z�5#�(*L��?\� T�Y�x�� �O��$f:2j�J�o�p~ ��3��Ut: �J��l_X(���P�+� ׄA)���w �#�D3�QE�;�A���]S+IG[XD���Ƞ�.g� W��	_~ �o���.O8� ��H�!�JY���L��?t*���	�[0����J h)
 �>��#\�(Y+� `������ b�/�V�} �Ŏ,�1ܖ �_T�V�	����W�ɶ 6סh7%	9|��V΀]���g	@�� ��a� �TXOy�\H �m���+���$H* ��>� �fY�M� ������� ���`8�QV Y^�!RH��.9ǰ��y�q ��)~I8_ �����Q&� {���a�%T!��@�_~0�u<��r P�d[n��� ��{V|�� �=P��*Y� !
��� ��n�G" ���0�蕐��t� O����i�X��R�ZYq� 3�_֚�� �Ԏ�;�N�z)+�岌`H: 40
콵��xx.�!	%נ��l �A��@� �}[/ʼ�c �tw,!�A��^� ~J]��.� $N`�� -���7� tBo���V �%U�R��8 �)_-,.� ��1�5�� �	{j�� ��Q,X�� ���� 
�1�^.+�� ��L�b��#�[	2���(�0� �/;A§ͨ.��[�, �=n�� �:����� O����~ �WK+��	 N�ͯ8��>^ ��gn	 j�1틮��~��)��S�(Ui�<���Ҁ�0^
ՈcL�1X�Sxs ��N�� �����_�� �������xQf'!���� @[��yH� n���ch1� z�!�bOpe YUP��Q� ��Vd-�c0�)�&�d~ HB�%�w�� 	�*������ )�_5�U�#PT��Q� ��_sd	 ꂧ
��b� �a"��1 A�ݿ>�<� (��,��3	���`0Ⱳ(�9f�Wz����F Ek��9j �^�7�
������C��VX�" ܎mH��꫅����l �%\f��?� Z`	��'(� Ҹ)��i� ^���A]� ���	� 9#� �J2�0��hTf�K�A�� �&I՗�b ��.j�tx�X��Q`�L��} �-��I>�/�����U��::{���I,�^\�D@x���� �ѭ� �O�֜(� -�ʄ�l�/����. �Bd��� ̌Y>�� J�`�%���$L3� �K��}� �x��2�	 �eW�Z�*� l�$u�_	�R� N�)�P ZpHX��g A�j�k�+���  �h0z��'_pW+��KitL �[!��� ZI���g> ������ ���/+�w8�O��A���:/��� �uj�oA��W ��hZI
 ��",������� ��.�j�� �5*�ǚ �����KyUl�� �1� ��$��ph ��o��"�\�$_A xS/�o������N��v O׵�ŀ�P~��V].٪:�� _��>~�\r*��-3Xp��[2�{O�'p�4���&�� x�鼝��%sy��۸� ��������c�� �"��� �H�/(y ��d�j�{�R��P`��a s��#��W�$+?> ��el ��huy#�Z�(���bXG�� ��*P��5c ��ߴ�	���'�@�2�x &ZI�	\���@5��$���� ��d ���wE e�W�U�# �L+$�i�� �QN����Y^hk� q��N&�	<����#
��}�	y�����L�]� �K
�~�����w�)}`��	�
� cjQ^��?� B�@c(;H�1)����z:�< 0֑�d
k�\���Z�P�h .�S��XD�*�k����U�{�ū�����x g��ߔ � v��Ї
8�X�������	T���ya���S4��\��P�_�Qa2� �V�8�1 �D�f��O<��܋<��!�XA���a��+_���Pp�J�`9ƀ ՝�7�X����  "�����Q����� ���w ��w ��Y��u��eB ��
z� ���)Ml b��TSPV �kz�Y�X�^� ��w��L?T���P� 3�=��s� �����Н ��=;� -�:���)�%G�``�� �R	��5� �*��S�� QJ�̲3�W pr��,^��\�����2�-�b�8���2���R P\��Z��K��&���<��E %)��mJ��XBi �!@�|�O �len~���> ��� �S���I�2 )d�$���U� �'��Ը�q�5��*S䌻�s��P
 �1��b䕨?���f� ������ �#꼻x����Vu�s D� ���v��P6�R �)�� _Ҳ@�[� J��r)�W%�à�A"Ή:�k�C�X��+�ޗ���!�� ۅ������ ���ʻ�H 42��	�80r�Ƚ�� (�_��`��[-N����L�e9 
 ��I�Z �Np�JP�|���=��Xږ �(��rms��t F8$�?�� dO��u� ��4��1�ءX�(��:�S�<W�����ٿ\��1B@��S��,\�� ����E ����	��3%h�p�L��% ��`�I	r?�;��B/� ��Am� _�NE���JȈ��H���-98�Խؿ8 $J�<.@%CQ�Rж�9�}��X(�ZY�� �VU/2�� ���+�G{�?���0���5\ $P�O'A� !Fk��N�� �ɚ���1�(OǊ䠼B�^ �z%l��-�:gvR��$�� �6�%���u� ���*��� ��Lg%�� �:���M=�+�5>��0T��j����<2��� �����Ju� Q;�b ^��� �!�� M�6Q~ �Z5�q�!�Y0������O��	�~+��Qb �A�H3�&pR�	�Ȏ��o1FŃ��/�I��%�$���Р Ɋ	X0�Z ֥h�l�%u�ڃi��\��.=����6Yʰ� g2	Ó��:�� v�Ѹ'P�9h�_�Faa�� �� :�	y�� Zz���~_-� PN�?�����;�@��`	$ �_� � �I-2�`h�jL�P���:��1 ��Tl�� Y�"�!ߨ� ��[�ƺ$ �5L/W�6Q �ӹT2��Z<�� \-�eY �_���������8J��� ��/��y�;`���f[�����Z�u��z�KH
 0�]� �d�_�m �w���q�Z8�r PFU8���$`VH�@�k)� p�����` ��%ܼP8Ġ���Pv��B ��-;1��p�|v�3�W� �-�D�A��:Hu��0=X \�gQhL k{1Iq����$3-����te���� D�[>� ��Rzi& ��,��wE� �L��x�S!��tW��Q B�V#��̄ ��^ �����$� :�0h��@�(S���!�Nx�2פ.' czǭ�ZN��)���!�� ��nR��8e �/�Y�� FI�S���� ƍ撴�\2DHE /q�~K0���`v?�ف�-�j��m��Z����ă����G��!D�� =��	���Ղ��y����� 0�!_�-� v�P*Ҹ�@:&��� �Rw	�$�x�WP�� 6V�()�� *N�F�����u1��>Ӄ�@�i+ �N�5��� I�BF�% �	��Ї;Q1���f��(��X4���D���U�i[ �SR����D���>7���0P�P�(���RTq�p�`� �΂KJ+] �C�%�/8�>s ��V�A�<��Ȁ
�h� r.(�B��8zG,T� jZ� �\%	��|����!� _��( 2�-[:�� ���&jDmd 
�>]�H�v��(?=�?I�!����$ ��<�t�w{X3� ��+��O$ ^�
%����� e����Z��E`G��( �� �
��Q����1�(`��	����o�h�' �.*��/�[ �J��#@� T}��N9ڪ�b��S�ɞ,��'��`�� �UI4]�?�p= )�Q�`A�� �0��|:an�&�>��� ���]~d� D�;�	hs#�mͰ9S
�O��� ��)+o�cL��/�9(� �ؑ�� �ru��� /L��~� �������.��/���8�\'ݏ r7����Oj �8�U�D ��}�εz�� ~�*�X +��
h�8 �&��o)Ck 	�D����=p���8�b�@�h� J.�N�C
|� ����9�� GzS��� 5�h(k Ĉ�'W��1rG�Ϡ� ��{5 �0�
�|p M�]A�G	XR�`� �t'\� ��W��|�*��- ��x��V����@Q
���>�#(�� ���O��y?BtW�@�$���P�����<~_���X�7�!k�G���-pZ;�䀆�jh@O b�13�>Ԣ���M `���|b�+ 9�f}[� a�<{tOwJ h�2�V
���	W/�o�#�иX��/�T� ���;�;_� �}�*�� �l~kx݋ ��h�: ��·�{ 	 rKxҵ ���,��f ��<	uQ�I�"�}@�#ً�UyY�):�� �̢��	�^� 7u�� 
1�Y��U�]����_��S��h�zڹU�� {��!� ��v2��	� �e�g �P&����"� 5�q a}��K �&�x�Q k�'��2��;�� )��L��J$� �&�B\Z��p�
� �U���Ӗ.����t �K�v�ȧ`�!�gX ͻ� C�~�D���������bv� 6��a��G(��!��\Q�� UP��/
�V(�{�`��@ ���!�R �e��ZF �ݤ��u�*&��J-����cX�<��f �[���	>� �
�SQ� �K��u�Wn�� &T�	� 9�G-'\�WD�5j�#J ���,��o� e������=�X �Zɼ��v�%����CP��϶�0��	� ,���m�s �S1��vB2f�����Y:��d�INa{�� 	�*�;� �Z��-%�~�' �;�E
��V��=�100c +��)��-�u�&���I1 xB�>rP� �+8p�K BQ�sy5�n U�^�� �_9�b	� ��2�%��� /Vv_�?�途���|S��,�7X�Hm� p�)ȞërgP¸;���
ɿ��H *�"_:� )~��^0� Q�Oc���\*� �VT�7vz `{'%�@����+>��� ���'�� We�%��k����!�Z}4c5F/H���:�e,���YV@j��� �X��S9L\)�hg"#��}�V$���@�[��0OT�����` ����Ι�)Y]p�Ҟ���� "�2�(w��#��e0
`��@���B�\ M��o쎃�� ������f� �ޠd�	� 6F1@&� ���A� ��y$T�J "�B� �S���^��z� �~����I3;*�B��(�%hfܬ	ԅE�T��� ���u?,  ��`Z�[$�� 
^6� F�|ed�s�	���0�����(r����� �[�����S�� ��'w�d/ ��	��[ ��3e��\�� `��h8 ,p����0�!�� �S��3�V �
� <�[�7� ���0�#�\��%_����� n3��^����/�\�`��B ��׌H��F pN� � Zh�3/~8�����9��t% ���'	�� ���Oy�$X� ��E<��h ��1�m�� C�R���� �A��/rU ���{hl�]0:�v�
:�R�Y!�` �_���� ;�nX8#� �Ro����> ��6�z$�U��e �Vh/F8��S�8� {z���3�1�]l���B 	���.� ��H��1�?��v �Q��P]� ���r>���� �/�K� 5P�h��|�0���
�:] 2�U���� ����D:���w'R��*Z9� @g�/�z�N ����1[� !@��*�H� է�/�S?% ]��V�-\2 �"ZѼ+ Y��S�,_H� ٽji��G ͯP3︛ �u�)�H�q������f [ Ћ�� ��w��� Z1ͺ�x�. ��Q�>� ���f�ѕa�^~� ��u��j= �X$G,v�w� Z��u[�� �z�?�S ߶�2�I���.��m��r� q��J'� |.b)��� �����` ���!з	����`���?�4��, (����g�Ĉ��O�鐋�+�r� �R���*��
ۀ��/'� ����$��@ �^�Ԡ�$�d�B]�Ǚy�����\P �/�@e�: �Ǖ�O_� g�aӭ�! ��\1�jA؀�`������ߵM!�?h-�֗f����� ���d�	�+ 
r�����Y�	���k�� �2�a��u@n����r�k ��L �.�(p�ǡ��`�̺ �X#��<�S�2��}` q(�[+��;E��~��|��[�� �"	�� )��e�_�U �pV������P��0&�_�;̓'Z�/�v�p�Ɇ ǉb�	�� �t�ױ�c ��hVr��,��M
9��*?�8� �@w��� *�����Z ��2�%�� "��	]��c_$ j\Z�� �Hk&	��*�y0a� O�R'�W K�p�%� �b�_�^�� �1'��n�!p|a�p?  �Q<"�$w;e��R�̶�XP;�H�sd��UP��J4�;�Ո�Z��8���+T�V� ŭ�p���?� gyi��/ W���I�� )�D�_�� Ľ��n��A=g�	e�� ���x�>�]%U�][��gi�t����.�S�(�q ��Q�	0��H�@X
	h�v"� l��ԑO;(x b�W"x �uoL��O��G�`���R�,������&�`J��u0keq���E[w	 ��r�ػ� �RP�g��� ���Sf)� U0�b�F%� K��e�r����\'
 9�IUqv� �A��^��H _'��g�S�L�x�̎�� ��W��߆�G'݀}�1�t �ifw<= �p���-9��7�V��)� Qu�	��A�� _��ɜ8� ���*Xߓ 䕠�4	��� ��;&�Ew N����,,R<g
�΍��.  �IkN8�h�w?)g����j��@ �G��Ub�$W�. h[5�a<�Qpi�_��v�3� w�ȧ��8 Ƒ�9�+� �`^k�� ;]��z"� @��D���~*�����B�S �>h�	؝w ��k�n[� x:
�3��� ��֫G� �K��Љ�W�!�\��0T�$x��'�Zː�����H/ OdJ�.���c>�S�! �� 8f��缾�H¸@�UӋ���� T�p�� �u����0��n (�P�N�`i�f $610�Y` u��S-�rB CתV��\��
Bf	�� ��,S����q ��? 	_���&0 K1���%�� �+R�4�t���ypH_�)��� 9��ڹ���/���^r �[�+�� `�X��0 �_k�{�� ˀ�K
�^�@,�� �;���P 0��Y>t� ^+�f[�����B���� � �7�w�9u��H�c �)� Y+�W�݅������ ���
��LK�1` kՁ3:�qD��'� d��LC��^�3�v��[W �����_�Z��&�2�W�`��^ ɟU���۷{���E}��x+M� �b��銐 ��Qɉ�� )׋rU��� "n��xh.� S�'�=��]U� �N��v <pQ���} ~�K���x�B���390�+�����#�|Z� �2�IЫ� P�={/�y<DՀb[��!0( �#��i3�C�%Bch�V� Y��,گ*$X���퐹��HB� �@$0� �����Jx �C����� ���h�dI 2��^�tz� ��,���� ��3�g� �~cv��� �(������� ��T!�_{�j"�&\�;�<�(��*���|��Sz	��3�� �g�c�:�U �#�Wt�y S?`_R�6T=疀@�0N��� ��]��z� �����\	�t�FJc �� �GQ���f} |�H��	�@��&�!����� i��?�,����{[��!�_����^�� t2�����4�@���� ��K�pS.��� �X+��U ����?��"Q��+�X-��Y���~^�H@ x���N�CP�G�Ak@�U �.��x�o�� H	�ִ��J	*���u 0��� ˃�U� [(֋���r@�� , �aXW��/�� ǝD	��F� �Űc�a$-Z��U*�l ���=���/Ȼ����0H%�����"=u΁`������p��� ���0�U�O,$8`1�@pZ	�G� �PRl 2������ #�J�|�3[E��t+;�5 �Yz�Nu8�B��� =�Z�޲L���KE���꤀"Z���R��|����� َP�ɓ4�{w�@��p� ��Dh����R�3 ͠���� �Y���	�[0��.5e�s N��3۵[A�P ���a�� �	w�N��$L�eu���z�Ӆ���{� 3�C���� ���S�, ̘V0�T ^�Wr��Y���I�?�v��d½h`�,e���I����S��H\ �|Va\q;t�+�_2��߬ 	��(} )�1�Y�D�߯@��X���m�\�I��g�%����?��e ҊH������*	���� �@gZU�� z��`�
 �]�B���7 *�n�v����JUA�e�z��X-�^�?�#ν�W�`��� ��v�6�� S!�w�i:K s�h|V	 r���An;���3�В�� (J\�%�	U<T�� ��؏�� �[���~W	�(,]�p�XR3E�Z���/���1�@���J��u䐿ps�p3��1�Z�#��� t���S~� ��U�"�F �LP��w
� ���j_� o�%;�݁f9�Q�d}�l��N��3�B*���8 "�`�Z�<�耿��L��z��a�&�Y@�`�<����Z��c`�/ O�( �4��Xhi .)�-��_+R�pW0�. !���#	9�^��\� �mK���� �/)E�d��ɢ�O0@��i����}k��0i{>M	��Z�7���&l�� )�L��� �S��!�_ �bٹ���rV���6�?��O��Z�Cb�A% �Ɉ�B�|� ����Q%�� @��̉L [������� ��'#��� h�2J$�� ��8W\�� �Ϗ
� ��V3й� �#�-���@ ��Q(��x�'a@�����R�J����C�q��s%����� 'M
�w�� s��V�YX�s k��< �F�	�>c
󼴨�� �]���*FUP�#� ��"� ^��0C�r ���P��}� �U!�~ ����%˝� ��t��'�t�?���*���"6�W�w�@� ����*��
i9�R� � b!��䂷 ������ I��:82� S��uAJ ���6��K�&sZB�+�W`��(�Q -䞗	0���ֺ�b�`��t?���<� Y�� Q3�J�- tZ�	վ {����� .%��Iɋ� )�wLu�
N������T �,��hB!���Q+��4��&�o�/vT������UR�YP�xW��`��Q`PK�[j) �.ԩ�Ӹ{ �SU
��j~C�f )�]�ɠ�^�±\@��?fh�`�)Z� ׈��>P� ʷك�(��!�j��]��GJ<�=�褈	�� :��(X�'� Y%dĮ�A�

�[`� ��a,W� ��&�@�: �_|��ND0\�"�h��\�� 9�YM�  `ta����< cp+/�� ���F�k1 A����*� -!{l�݀�)�hK����R0�G'��o�g�Q  ��)��4� ��Ct0� ���(2�@� � ���	 �\���hSW ̲��e3t �;^ �؉xz�i�s	���Z�%X��� zp!I��>�LHGl O��ԡo �ʱ~/yJ ��Y���\WB;`R�%0�  �=�����!+�@ \�w��YD� ��1���a �d�Zx	�\�� ,^&�J���9P-�s����.�H�� � �"���b1��)W���_ ������s	��j��Z��A ��~����9�؀�,0�Z@ 5�K�Xd$��;�)��!� ܂�.}� �f����s�-9�2`��]@z) *z��X+ ���.�����1�*���b 6T��W�A�>聒�2�;4g���+`Q��-������]� �K��!�k�=�/����h ^�<d�
�0J��$��AR��+��v|Q�p�]��rX ��8uR�Q��B�'N�]@ �y���1�������qMcO���	 ��~>-\lX h�tN���. 	��H"݈�*섀��Z �� �h�J����=��_ �3
Z�� U�#���� 9عME�/�rL���@��j?<�����-�����h��"�����V�{a�05q�:	���hA�i���p{ �G��ӈ \$��Y�X3 %pR�� ��7�@v �3Z (�V�k� J����C]��	�f�0�> �#'[F�N �-hU��~GX�	�\1�;��ȯ�� ���B�ژ`�] �L�I�� ���[�B1��%�v�aP*����C�m0�/�[ DpJV����:�h�e�1�2�t 3��R�; �#�[�(�� �^��_���N���z��U� m�!���1��
"�l��E��X����M����5���� �1��9:E_$�h|0~n �藉z_ �X}�`(D�9�����L���#2� �:B�!�� �z�5��p���פ{���젌	~�;���E�k�쉇 �Lս��;� SƩ���&��QIxO�e�b�%> �>��j" �gus`B� ���*!/�k� ,0�B޸ Mi\<@R)�?P� ���!q� �J +�p� �/��B�]�ډ0�\�x;�7�} G/Y��� ~�<��S� �Y޲�׺� �h�;�u{���6� }L>Z � `��1�+���� +�Cy�Y ��(�̼�� U`���A} T¶_V����S/ ڐ��� L~I�[�$� �,������\KN� ����P�� �l���� _Q�yK�# �^ǥw�[j _=/c���  q�0+�n� ��.gZ��ŋ�$Q@�>��E��/���H���3��7� T�	������ hl\�a0�U��{	����It��LA�	�R�H��� �������R�9� �F�)� �[�ܓ�$�S v��/y >d:�Կ� ^�&��� $+�6< *���߾!:�A��ݯF`�� �p�3 � �X���R �z	�Wmv 6�"��^	UՏz��"�\�s3� ��s�(�������.��� }�dF���&n0� l]�����> х�&j�8�g �ZK���H�u �H_��9Z� ���	�=?T�>����bP���s� �E��T��,&ռ� <�x�	�I�w}���0� 'Ap a\-��qN���ހ`� XZhk�|��E��(� &�#e���bHͥp\��4'���S���c�e ]�-
3^� \	(��SI���p���s�W-��BN� ��/u���b�� @p�2�U�c^	�w��)� �.(���� $HV�^'_���0萟W2@���T �g���#S=r� E���W �m����o 왼c/��=� "�V{��>�S 
ֻ���y 1 �[�� �@e!���u8�^����<\ (ѻ�L����©pX�<D �U(���:A��	��H ��\��h�3
�����\W� ��!Y�w� 赗���xs� wН��'(� y���\2J߫���ϔH SM�p��&2�J'�����`�]� �?K��?	�� ��)��' 1�ym�|� ��>Z���	�J���D*pa������B��ԝҾ@����� �NTy-E[A ��.��s�ꦙ	�w� ��3�� ���	wQ ������������p�.($�\_%��� h*I�]	"��� ���t�� �^.�!�� q�~�6�J̩��¯��8 (�<U�F�o'�� �#�P��l����'�XК� MZBI��� Tz�⸵9XhZ�(Y��}kЮ"���1� ���
 �x��%N �h2TUt� $�3�\����+;�����n'�װCW �9bU�$+�����hn I�%!�[��]-*�A������ 7���U?\� V�Ҟ���92����$(� �k8=ҏ^ ��U�b������ �J��\aB 'TA +� t䐻`Y�� [���Ux� ���@$�� �-B�Ҁ�� �TtK1�o
������
ē�;�=Yh�L��B� ��˙��o�(����{A���v�[9�	 �~s�(�W H��@nv���[��`��W ����D��X��(&ز�%�K��k`E�* �Z0 �Q�9H�J���x��c�a �]*ԁ��):���B �E �����;�=���=�	�\>�����2�ׅj� �@�,�x� ��SGĩ��q[�����+�Y�m�N��̀�R�,3�`��9[�  ϯ���N�� X��儉�] ���>.�sdMLjU�SyD�<-� ��QV��xX���7��� $�^��H� A2_�vyN<� ���V���\? $ĸ����P�_��u@�=H�] ȻS��/��W �(����x�?�U ����;	OD��@���Rv,�YH@� 5�� �3�B 1����O	\�� ���> ��4��DW|��]�R��5p��<���d.ѿ�u 2�X��;� Z%���t�`_r�)�(Z�LJ� �rR�| ��S���H� �z
#� ������~� ��j@��' NRs��Ҹz��� �� Y�ˈX͸Y.[m�	����І0ks,��?T ��s��	����x���;���Z@��/k }B�]\��� ��3���1r֘�����ft�B��N���Q
_8l��/څK�C*�, �7�O�lP �t����� � S"�[e����?�Y{ �J���+N� طk��u� ���&�� �\��9E�0����L� P��� z8��>4� 	�lC)Ә�` H�ʊr� J;7�ý� �.FRH�� +���c� J1)4�������~��T��e� �r�A�o0�/(+� ~[¡C�ab
�'����/���������7�H"e��JKN8;R|�N k^�[���` qj�b$F����aA��� �!-�|*T ,	��1 ��Yr�.B������	���U.��]0L��x_ �J��9�PI@��i3� ��	��tp.��V S��KE�ÀP��["�X��S�(�{͆!|�}\Կ fZ���T
hy/0������p�� �����H� )�"���  �R0��� ���� �}�[�PU �h-pg�.J�� ���z�`���}����Cr� ?��ຼP N��,OA�� ���v�� ;�8��JU� ��ds���W��֩ #��ZzĢ� ���d] {�s$K� �!��9`W &)·�����Y �{y�[�� zU�$ q�3e�+� �U���� �^`|�L��	�(C��K��H:cB�&M�'U�f Y�]\��׀�5����� ��(�z�OhD�xJR� �t��!�o�گ/d*��xQ �B����� ��/Ư# �S��WĆ>1�����@���0���H �w|���7�5 &���]�>� -��y��dZ��y ��%���0 ��X+c��$��,� 2��	.w��s�� {�; DLT��_t�A� �/�- N�.�0����\^h,�* ��;�'� �ؘ4�`�� ��L�m} �M)U`�0 [�����᠒��=󥀁����9�b ��P+�Q��oq�7��� ���e� ���Dc��b�p��n&$L�y�U����~� 7���&x ��,�b� k�"�0ߩ KG���_ q����ME\�1A��u f�C<�i ]g)1Z��\2r �����(i������h� ^ %X��� �A��FE� ��\]�o"ºd���^����42S����`���ڣ ���R��\�� ��
�/Mgzv:�bn�� !]�0_�s`  ��xj��J �@�aT��3�X}���נ �?��xf�<������.�^2�¤I@B��`w� ��Ƕ��� xVZYU�� hN%��1��x. ��F_��0�q��QS@3G���IW�	2�w  A�1�0� b�K�����P���"�����Z>0�E2� ��y�M�-J^��q{���/ �T�-0h� ��#���֍ ��Y{�C�L;��@���,�z"�����N	�W�� b�;��X �ȗ�3���hpZ�`����� K�Dz ���̈R�5H�'YĀu.� Q�/����WZ�)��+�(�~��<�.�� �Z�}*v ���V����]����$����^ ¼YӬ�wr>1� ����	}hu�[��Z0� X*�fhYs /�˸x�,$�% ��+Oݫ <���j� ��J�a' �;��Ѿ	{n� �`$� �ꈒs'\� V�|���� o��)B� ��Y[,�5a��3r�I�W��T�B�7x_ a�$ē~S� �`�T�����$ �w�sm+ �������Ch�5
����9���$��k ,�A�{/���ާ$� �s��"`L1Հ���AH��6����@-���7(u !�+��Pl �tܥ�_  �[�� "#�;�}� ����)ũ ɃhE=0��91S�ݻV` |��7- �P��0�d� J�?���X�/��P��(����@��v��1��3ǋ���|YO��Ȁ�)��v�8�I�� W+ʿ�) |�#a_�! ����
�V�� 2<�� ������ ^��f�;�E �P�h?�� $���cN}5 UC��.�g {xȟ�2����4|�.��*�t�� �!f.�@�h rm��]��Jd��	���.����񫋽�w���V0�wV E�(�݊��t#�1���-�� ��Ԩ�	��~P�҉���̼����Z�K1?�Y�QPz'�~���a��h��_1���l	���� �Q�8i�J�s, �AGP1�; �g��7 :�9��\� (�]�N�� ɚ����B ��!X �����Z��E[(��l�o�4�З1�\���������P�N[�qȜpA� \�Y��o(��O��� h�;
&8����7 �/�@x� �1��K\�����Y��^Ef���_믐ᨉA �#�*�� �YR��h� �k�P,V ��	��y� ��Ձ٨��EOؾ eS�J�� $��2_x ���*
�� UX��ȵ�� �Z� t@�� h�aN��$ȍ] FO�5�������Ӄ�x��J��(�X�΂�\P��M w8�r�%��9ɀ�+��� �;��b )"Y��>ZO��������S- P�7Kݥ_��# �W��� �S���U� z�w��4�'���Z#�Y �h�}��I����	�0�*�q 1�Y��/ �HUm4RwT	��)�-D�� WK��u���:���[�� �d��X�� ��w/�� �^!���5� {��n���$q� [X'V��`�#�I]����m /���� -� %��L;�pG���`B�}X ��cHI�%xݟ��`L X���G� xE:���( �S�����,p<�Ҁ�d ����ʲ	W8���� ?@	#� �!���� T8�h�tv	wA�Nׂ�<"h���Un�,�8�V �.�A�%@�K	 ]����0 �Bd����$�nx�0�bY�l�ظ\����*@�|p\ ��х�+���W�"!Y�����. �w9���~; �F1��ѫ 
U����uY;A�N�*�H/!r.�� Zp�N� JQ���1q�K���Ȱ�D ���X?�����a�c @�n9�U Ŵ��庨 �X�GM]�B ���!� ����`�E���?�� ��$��0N�B �Z@ �)����\���<��	��LZ 7���Y�S +�Tu,�ң����`�_8K� �p&J��� `���0���� �;a��x� /�>�נC�.'�� D�(@˪ L<-��bd "[Xj� �κ'k�� ���NW�=pU| ��Y� ��R<J��A�L O	�Ȕ��[8�P�)���~M� *����� +�E��@�:z� �h�q� H�0�s�P:�W��a�x� ��H���\ �DƝ
_}� QW��� ���(�U 'ʱ�aY���.��pF�)$�V�P �E���zr��Lҗ��_���`p���%���Z �h�g��>.�(�U HdN�h �A�nO�8�G ݁�Wi ���l�� �o����A 6W���;�d|�%���^� ��_�*J����H�u/�; �t"�\�$ ������X٣ �W�{S �[���D+�� )8�^�i� Av�j�Ӆ�����A��Sp� ���!N�Hb zo. 
Mh���K {��(̫� Ƶ�"t0�K���h�S� 
���G%1�|Jk	��9m��YW��~� K��B�,�\��fՑ����R�� 0tK�vP�p_ �ڱ��I��-f�2]���� ķ�Aj�9� $T͗1��. +��3
���L�>��0����1G��� ���{풨 X��(�"Q=np 31o ��� Շ�����y:���+��.dv� ���c��A=]��Ɏ)����(R>����Ao�@����["�ݻ zKHCrbU\@�>�L3!�Q+����\�� �~^� yh�L?��Y ���3B'W �z�q=���R�G���(�'! ��Na^��z-x� �4J�@( �OCE�)ʫ ��ݵj�1Ԩ���t`�g 0.Sb�D� %�evFa�]:�Q>s����-
� q���'�j %{����Y� D�w9��� ���0	S�� }5��� �I�s� H\���U�s܇Q�;@:�|��� �1���b� ���u������� �E�X� �q���% �	��1k. ��~�\� V�Gh��s&���B�`o�@� 	�[�� ��Y(�k f�h�Pm�#��9 W�V+� �N�Q;���,0�Y�b@V{5�@�P� � �q	�R(?�Uѡ@0�಻ T_Ҩ�w
�^Z����$���[�Q>���I�5S0 �Y�ޏ�![L��}=�-L�����@Fh\B �b�S�R#`���k`X���(� HX��y ����LJ�	�� ����^�a��,���y���� 鄊��_�-yp 3��'��� �W�o�r��� 9]̅��
�)�Vʫ  �z��x�`�u�9%��@O"�`�sL�� ��m� ZR��Xb,�����A�n �T�@��P �( ʲJ�4��]`����9 �T1���Q� n(�A���!|�	�}	 ��By5 ���S��' ��~�`iAPρ: 1Z���/T�@y=D���p ��W�u7� �E$Ba) 3�G�J� ۽��&~4F^��"� ����6� BQ$�'\Փ���� 5�Co�j� �=˩��G
�)퀺st %������@!ׅ�-	�_��� o[>rPf ������]� ��ί� v��[6� �'+�Hn����"�{�P�`��2�<c�+��� ����X(� Z�:[�~� ���<3ҿ �gj�D��\X�ڪ@��h eA	�͜b� W��C��� X��j��� B�3א�e f8�x��_H۬o�˨��0� �m�:��� = �w��YV���?�T�(X����O���*� /8�Q�!�R �DV��H�� �<���� ʇf��N\� ��|�1��j�I���O`xb_� ���Z[��M ��@p��� A���H#�/�(b��K@��E �-Y#���z Lnp,.�V �i�/hEJ^ JR���	 ]Q�Dx� ���|g -�A�T�� Ju�LB�!�0�r4�+հ7L���*} �z�K �I��A�> �f7�X��v9n����ӸH� �2��p�*� ������:�uT�`��Dy���$��C�@~��j>� �����$ ҸYv ��.�pn���G0x K��ٔ\l ���
��^��Q�&��j ��}|	�� ��p�-(�V ������ ���Oz�$!�("�>��`�	� ����_�
���Y����� ʊXf R	�� ��B�@�
�`��f�5�x� �K2�� �\����� �`��	hx8x �o���� ����c#�O.+K �(�� u�MI,[����U� ;)��i��w? MҾ,H@} C�xO�FI� NM��D��2��%�� � �) �WJ�� ��Պ�
� -�OF�~	 ��z�ti� (����
�s\P��S��i ���͸�� @�HQ� e8^b�t
 ���Q��J�砀dY3Ƹ� "�Ɂ�{�r ���R��f0Zߘ&�y �p�,\P����ڈ9 ��%3��+�IS4 ~oCr��~$�8R;+]�-��s�	��� �9����y� ��][��i ��Yr`�^ v�Ǌ��H �D'��1E�tj ����?��'�9c���� |Q��-�4&??������0Ʒhr�+�f�U�G�4��������p�k �M���Y�N�����o��� �
����* �P��Q<��-���bΉ�L鲝����� N1�
���� �ߏ�5Q��ۗW����P��Z�P�" �`�DI�H� �+�$�Ȣ ,@� �[�� \��h�*� �3����
�νK���]� %	O�2� �����i�� �S��Y��\��� ����R! ;����x� FNZ�w)�e
%mR���3���'0�\��4C�~���ͱ=+���03���
@f���� O ��M�:�Z��N����n��� (y0u ���3��,/ �F�~�bk R�tB:])j� ��֕VT ��X*����� ݴ}wZ%� $��Ǆ�� P�L>3=�� ���AW�; [��T_��� �Z����">�t�4,���Ѐ �P"��� .�i)�]F�&ln��k!��Wp �KQ~��
 q�����1��҃}�	�� �F�[M�� 12�Y�9� �"��>�hADO
��E�S|�W��� ����2)}�	�]����Z��˗@ 0�8�db� �C���[�%!���q�o0�����	*@� ?�^͂�(�_h�&̀��Ow ��#]h� ��x�J�� �?�n@�(Z Ӿ!�1؍ ��8���d	 �x��\, 2y�@�`�Q� ���{K�,�2 �`���xt��P/ �ն� ��L�  ��t*
���ӆ���_�� �~C��x� +�꽊��LQG ��D�	{� �;�7��!�.�&�`g< e	��wԳ � �B#��xL� ը��Lv �y���� �$^����:] �fܴ�J �Z���p�/�0x[-I@u�� ��Qi/�鳨	���� ):�LH%��������q�1i,;w�1������ �0�v�'�Q�Y�����p�) 9d���G:��X� �o��)��3��M��S ��_�{�B P�)�Q�U���8b(��h M�'	��Q�����+������` d�2��� B�P �� ��1�Lx��9�쀫/;t�� Z�.��j;	>&�� ��V��  �X�\�;	��f{��x`N��#�~�0��/ �3Oۻ) z��@N޺�����1n��N~�W^2� �a".�R�1 z�/���� ؿ�MJ[�E��Үz��K'�C@��� �2��O�����] � d}���)� �H��v\ �� ['lW�a-�y� �\YQ�;��X@�B(� [��H��Y�; �?Z�&^] �=(�\Ui �3���� E�:��)��� Z�껎/� �a�$1�S%9=*����׳�.���� `��7on2 ��Ah|��(���
S���� ^}��]�: ���y�Oɮ ���89�K �D�P�(� ò�+� ��u?)ۄ��K�� ,ђDƨ�� ��*�F/��r�}���@弅 ��q�Pަ b>��I���^�� {�+;A��(|� ~��&
_V<��,gV ��ɢ�m b����x^��ו@(���t ���pxr�Z ��ݺ��9�%��W+3�� 7>��5.�� h(Ȝ� �š�|?� �ێG5T� )*�ʧU㒏0�Q�#� �d�	�XH 2���-�G �����<U��!J��r�] -xD��{E c�7�Q, ����P@� ߟ�?��S �	ԙ�� 0�_���� ��Y���3 zѸh}��	I��v�5�	@xY3pL+��d�z )A��KŞ�] �َ{� �2�R��źXs2 �����&� ,�CSR�u$cJ��l� �1�+�%� ���K~P ���o@'W�6��`YC���Aau
Ke�15@F��fw�Ř��� ��ߐp����	L�=��Oh������P�Ha?�/ ��C��PA-��� &�H��D���j~ȱ	X鿜 �%�Q? ����-�:���&'��h $�W���q�� ��y\��
��0�� ���nX Y�/57~[	]�K��Wb ��HXZ-�<<��>���h���'� �gL�	��<_���� �0���N ꪘhT��0�%��j�0\6�}>� $!���%" �BV���Wr���wn��T|�`�� ��	�)Z�w1W(�c��� h�l��X�S��Ā�s��%	��E�&�A��@O;�vI "^��i̜�l	Y �R�}� fhI#����	q���ph���:��� ���x� >RN���0 պÆŢ� �K:�NI ����$�́����"+�@�� PB6 ��E��-��Z@��iH8בp?�
� ��F65�����A�[./ ��7��� �,�;`�� ��J�4�� �!��'�t� 1��(�*��4S��#�ޠ� O�@�h� ����FJ� "���(W^՛z@���"��C�4�`A
 }r�����	��t�����Q �k.�+�� FXA��{� -�ө�0�X �2��V �d�?)��Oh�A8U���p�� ���	R �y4������J {��!�� �u��t �� w�2#r%��:���`u���� 'E��� �]0�� \	+���x� �:�aW�I�/#sp�Y �7�a(fS������- �$���`� ��x��WR ��⥒o,��;�N9 	���v ��+�9��0��"�]$�� �T��~ \�^�����鋼�pP#�>��ʉ(�0[�	V�4 �*���/[x�k�F����C� #�P��:�|���?�ղ� '��3RV�I���n�Ĉ�] ���ȥ�Q
 ��2�<�yu�9� j� ��^���$�;)��RL�]!����@�+�P�n�q��*=p 1�R�	c ���\�)� ����4��������|@8	p����� ��7���w@Ň�1� ���-0�v�`3���m������ z=WIS �9"���v� [������x ��_Y����k���h `~R� ��#,H9�� JV�.��v1����b���H��N �t��¡� �d0c�;!�O���?���PFɌXT��_�H��ڀq���S�0�yAZ�ȁ��X.3:� �@O���F7�z|b@�� V>&G\� R���K�" �v~������ȏ� �,�7������(�1�*�֟ ;�t'T � �W��hyX v�+�Vܬ�0��(�[z�������p�� w���7(D���-��\�&q _JI�i �|O*�4�9�Z�����d "f'�WE�+��䶀tR�OU�!�8 �����|��j�����0���_ 	��%��� P�}����?B� �FO@��� �P.�� � X�$Ui�� (�kY
� @\Q�� �ɤu�m� ��@���hj ��ϗz�-��@	Y9�� ��a�5U �猆�$) -���_�R���*�X��-|A�� �!;��� /)Hx魷 �(� օ2�X�qn���&�	>��P��b����Ƿtp�W� A��c��k� �Y�^	�` ��\�h >�'
�dM =���~�Ĕ|P�8 �S5/h�� ѥ�Q���S A�;��@�� $��,2�^ \)��� %����(� ���Ȼ�� �\]�E�j��� ��V+� �po]��� ��$0�TR,�Pg 4m�� :��h�H, ��%���' Dꐼ4"�$ �$!b�]h�Jỏ4�*� F�ѝ�-K� q�"�\�, ��c1	hQ	�(:B��+��А2 *�oK � ]4�����^Z��GB�U�`q�> ��r�� ��]`z�� � }"�\��,4��`1*ċ0�Y�&�J�Vֿ�1��: �^��"� �Lv)\�� ��*�PK� gC�	�z��� _�uI]���Z�k�{�� ���`G)<�,�'�_�Ï� �/z	�^}�Է�`�<� ���vX�K �q`� ��ٗ��0�)�+l�(��[ Q��S�� �Y�Υ�i�8�* �U�W
����ɂ ���m��� H�/�i� Us�� |�	�M_#h �+�1�� ��]�>e��p��W`P,�dBh�{��. ����M�� A�Դ�� �w8���� fQ�p�&� ��������@q\� �(��� !�0�3�O )�8���=U mR��,�;�z� [�A�]�`�\�7� ��!�	� ��Y�T@"^��נm��	�@�2�C9�X�l �1-+�� �t�n
�.ȈfV�Q���a�M�� co����z ر(N��# �PX1F{�� �;���� R��N��� ݨ���I Xw��%��� K,ً��v �_�� � f��ы3�� 㚵^�� �%�v:bB���x�?��� !����:^� ���}�5�������Sމ�|�B2�1�C���F�ƕ���1(XS��V����ExO ����]a C�j��7� ���k��� L�KP��Vi%p� �ܒ9~�z;$ 	�G�HD �t�8��g 	��˅' ��$6F&Q� 4A{�* P��RQ h$lgk\f �4E&�j9�	�K�@ eꁀB�h 7���B_���{��A��j ����	(�ܔB���Z[�:<��|�'W��tM���� sh�TY����K��/�o��ؽ T�X��Lx���$A���Ut� @���\�5 r����* ������/g�:i|(� �����b�:#��D�.�0F �
!�_�;' ��ژOU� �4o�$H8H.� ������V��س���_ 홪0$o,�hE�T��[�`�:ʪˤyS���V�DG���K�8� �J���-_�{!�׸���J���Q��� �I0K	� h&�5ז�� �)�[�;� պG��, ��[�U� whSʒ{�:�&��`*���u_�"Óp^��/�h-�S�`�b�R�'3[�� d���۪ (ƀå�i���p������������b�A�c�'�+�,�< �e]�&�շ��=��gZ� &>oJ��(���� n���c�� h���&�a�@0[\ ��1��_ ��<� N� ���u� �#�h�VvS濨9��z� ����� �fC<��8ʌ 3�ņ�?������Yv��MK�������>ѻ�&�P��cU K��[���Q1���Y�	 -�N��(S� ��Jж�d]$i�_�_�r�P� �{��C �b<K� �h;S��i�� �1����t ~/��Z�!=�wRAĲ���`����O3�1Wg�@��� `�B���A ���/���N �������H�t��b2�l�&�#0 ����RV ;���#� ���{�!Oc �%1V��]� iWe���!P��u� �zRZ��Q�N���2ސ v$��
"� ���]90�/YG��C`'�ײ �T�@�) YX��
�hd�iK�Pt�~�����Z�� �`�r޺�@^h%:F���� N>�υ�B�X�me1!�(�U� %bZ�����wB4؜� /�	Z`������@]���e �*�{�+H�C�ٞ�$�@x�� �KY[p� �60:</�U �Dn
_��� ���"g�� �U��a�� �݇�'�����/�JD�	�����qp^��� !Lё�h�� �Ŷ�< &Y)Հ��1��$�L�	!����:�1p�ʗ�=P� ��K��;�1��d��@y� �B�ر��D'���T_X����4d 2��)\�2���^�� ��	���_.VUr�&z�� ����5(X���kW-@�:� 1��?��]� �h��гJ �M�y>�� )�U��8sj @��w���9%�H�� �L�i�� Һ�S|_ʽ +{��'\R �����I%� �����`~  W/��X� �"
���.(�"4�@�P�� ]�@����^ X�(��N_� M@�=��òr� �R�oB�]y�?�7# ���� |= ���
�g) �<2�$X >������ۑ]
f� �Pt�( ��-0�Ր !���#/�`��=e�T Ya���+�b�� /gv��8�r@	�J*�E�$�P �ʉ}p����f�c�� (��������$��6���Mp� ���8��z$(�A��j�_��! л&O�-Z ~�%usz/���3+�E) 럿S��f1[����X�  �q@��� �8����{��LAD��p�[��� Q�N�g� д��c�8'�x~�W�m ��\�(��� ��)ٿ�R �	*V��D ��X ��Y��y[!�π:U@.��v���3 ���e	z [���a � h{w��)N�	���� �K��
 .P��fZ  ��;�B��/ 1тb��Ul �V�ٹ |�*0� m�s���/�V(�\? Dz�,0ے  ���QŹ �Vu�� ���X�vtY�P� �Rq�$�| 0E�Q��  ��Z^*�F1� `�R��� 0h�6qE� *�K���-x�%��t�$�� �Tb3�Wf^'�&�|���S	�s�UY%;P��C <�x�k� uv�"�=tN�� '7	0��+���ڽ���Š�V
[�X�G 'Y|���h�Jq_ �����ܸ	��� 
��D�������� &UBW L~$� 3�hG�����J�"�\v� �%�	�a b1��T�;�V�� X#�)���o	�"&���1�Q ��M�$[2 �@����- ܗ�Y�lh�� x����K���� \��iEI�	5�w_0�e� =c\��q�L2ZB��@�6$
 �'d���>8�1E��* wNu� �k0^�;�YZ@��VS";'Ё�w^ 0����� ��g��(u�� t	�V4�T�� �� �e�
�� �C�D��:� Q!Ֆ�Yh�]+����O /��^��(x�R!b�o���]� l-���(ʺ �\ �|� ��on�_: �����w� 	k�>$�� �
|!D��.;����TI��/U ������gv� 
�Q�/!>:)� k�-�n� p͊�x� %\���0B ��1�l��)G������w� ��_�� P%,�g�yJ�	����@ � '+�vj�o��	׶�\e�?�
�\� ��dz� �U��0��!ʀHǷ01�p ��D�"3 �V��'�� ���´h?o ����V_X#]� ��4g����`��� Y8��:��\,~ ��#!�	g�� UE}8l�� �\����_� �F-~�2�a �h�Bw� �ϰEJ#� �Z��	F}` �o [M3� �>�w�EG���vP0� ��9gK� ꓽ��� �j)U�( �}R��� �A	�`��
��1� �p�	��z �6���0� ��H��� ��%~�OL	����ֽ���ƫ� 7�v 뀑C��$_|��u%3���z����t�b:"���ı�:���M�RX} ��n��p���/��ЀК=&#Ѱ ���(Z��No�s�AV�%& �p ��d��\��	 [û��%.�h 㩖�cL1B��"�Q��k�=� H\]*Ъ (�1_�B�h$�K�iؠ�(׋˸�JZ羨 _9�4�N W	i���/hH��f��$��	%��X/ꔻ�Lܚ� P {�]Y�'�+��GU<*��C�e�	xb4;�H~Nr� ��A��W)x�z���
� 2�=��Ѭ  o)�X|Z��v�/���G(� ^��&�N� ���X�� ��� %�ʩ �lW��F _��>	O X������tp���$�1��h�6�8��Ď 7P?�_a�	~� w(X`� �S��|# &�PI\럡*�.����?��p�NĈ�,]e0��  ��R|�'Q����Z_�b���D �[pQ \(�����'�XA)za���$ =�a��k����}��2�/� U,��ѻD�W��4� �q��a?%�L�@8���&����f_��+� �$����*��1��H!�ֿ,) �nN�5� 0�c�	7�����K�uXC-�_<����N|���T� ^��0ų >X���VB����M�5xH�G�^X��J�~qh�݈'���� ���� `���hP/ "��1uI� $؁�� H
��u���_0�#� �~R�y�h YK�pW(0��K <���7�r u��M�J'�����q\���3�`���I�Ȁ(���r ��)Ŋ����f,�� �����p�a@5�v'
�w={��U�JG ��҉��	ڨB� ��'� /�Q��\*��Z��(��^�&�@����Sm�xҪ �|[!��9 ];�Ѡ~�{ @*ʆ8�)������*.�� �	��0�� ]�ߚ��T������鄔w�3��$؇���U� Ͻk��+�����\u���Q� '�G��% ���,)�<��,�d?���X�����U����`��PYl�*j ���32F�0H��*��p�v�Z �V �[R�� �^��~˭ $�8&/��� �Ǡ�Z0�� P�ى��� ��k��(�J�N �<��e ���Y��(!x� ׊�B���; _A�ڙ�+�bPU��������>�)��I?�� 8+��%�p� O>��(��� Ԑh*�xK]��CϨ9�J ���<� �LQW�4�� ��`	ֆx� �$[�h9: �2f�_����� � E%o ��<a	�8� �V�?J[�~ �/�8��5 p붛ĲI �:$��'� ����`��h�yuć K�%����&��� ���-V&x�g�"b1,�`� 
<� a�	W��Ŗ����k��h� ��!�����2���2Z�`QVݴ���g�!�s�& Q(1��T� z0�߂#+��`x��Ot��! �_�'-�q 3@V�ʨ]�5�1�@��=R�̓X�vL�*. ��UQ2�A �[d:������ 
��VO��Qؿ�|�H� �TD��w1vXS8�@� ��u␎D i뢀	3�� څ��� �y������!6>�`Gį@�.�N��v!����J�K f#L�d��w=��\ғ8 � #
�s�)� I|U�̈́ށH�j� @�Gg�0��:|�K ל���R� ���(Z �~�EB�qU�S`��@��_ m������ ��Ds�� Sd)��� ٜ،p�R.f1��s '_�%@�&ŧ�G�,��Fu ����&���D�Z��Y�����������9���]�[�>	��ח�95�� �Ɯ|����\{K��msҨ�'5 @3
�w�����gH:���#Q`Ò: ��d����?�  �k���� ��l���62	@�$��� �_��o���5a�W��`p�[� TI�J(� �U3Ƚ�c�ե/�R �*E�;�� Zy�x:�\& m���7��� �,�(���n�`���O����f≅Q�8���} �Jk�c:X��(^�`�ϝ� ��G2h�� ����$���.ȺD�=� ��Z�*> K��q�Pu�{� ����#_ ���"Y�$�5������`˸� ��S[���;�/�ߔi����@�"x��1&5�Ib� �X�t��3 ΂JÕw�� Oi���W`E 0�¹��� !А�Z�%5 ���� ��_�絁�ét� -�⚘ mX3�������R�Ӻ�b(���U��)Ш泿 ~+���K�� ��)�E�  C�:� H�R-"�� 4����v�8�쾸 ���s��� ��yI;��������<0��H]It
�-*�xuB��d�����1E pd��~	��nႆg U �SCA_9���
V3�� � C㟉8����q�3�<�һ����w� X�	8�A ��Ȯ�^��  L1"� V�w���Q. R��dF�_ �1��\�� 2jkI'�/� ��P6?�a�~�9�#�1�����U�Kb��sq?@gO��� H�
D"!�:1<z�&�г@8?�*�w�@��>8
���S �*�q|� Q����Ɓ �XU�6l ��0����,�A0 �J@�(�_#P�Os �j����*� ��J�㯞 @��΀� ��%�X*�� O{� �S� �K���2� �_��h
t� થ*� 12�/Uͬ Xi��[�
��Ш'HrR ��vɌn � �!��T ±����R� e�A������U��M����2ǉ�T*�Z�.����E���8؅ �����
0 ��P���� �	�#�Y( ń�uS��PF��^��MU� �&b���	 *���蘧� ��9�!�dU��k���>H�o ��b;F=
�9'	O��-8�Ệ ��He�$Y�3� ��-[鋿Pc��}Z YG�J��'3BT� ?2^�`��������(�@ ��^�"� S������,?���{�@��T�AϦ���J�yV� R��*�+> �F����� �¦
)�� ����hBZ+  �Q�����eς�IR�%���`Y[��A��0�_���\�3� A�8.-Ȧ; �YH���J��� c����=�;����W���vw/ uw��X ����k���	�>�I�r�� �Ah�X��~�<�U4ԧ��&?�� QO��L� Y��ܙ�q �4��P� �DM�1�Lu�QB��P$��G �)x�4�� �|#ϰo3�sZ<@}NY�� ��P�'�A� h@�}��� �&״��F Ȋ��	�(:AQ��箇R�z /
����uHX� 	��U s�f��� �{���5Bm�� �GM�_�̺I�U޽C�:�� �K��D�� �\��d;��C��K��]�j� �Z[�CQ0�&�	��S��|>�P���D���� k�m����V1վ��(�s���`���
�1�RT���S d��0Ng'� ���� � P��j�}B�Si �宱z vr�<-�[��
�t�:����i��)��h0c}{ ��>�����Hj� �0�,q)�麊�3L��b�} �K�	- 8�)��=/ ��+��|1w Hɯ�rjT@��hb�^�*��|�1
��X� �}�I��<d8K� ��E: �6$ -�\ 	ab?�%p U�y�>���Y��J��@��h]�4� �%�+���[��6  H�	ŵt� jk*S���3����L�}&�I� M6��� X�2K�d,�$�.��M����  ����&( ������� �?�Z�A�uo �DP��^\����O@ 4��],
�� X��!�� ��6���� s��^N��
_*��K]���`+ �R[�&��p��.�!�oG�Xv� Mݧ�������@CP1�(Z ����N�Լ��H���S�Զ��U��������<����m��v' �ў��~y�(R��ld��u �W���3� ~.�D1��@/�,%��x0Lhk\ȡ�iE���$౵~ =��dR .|,�� �����=�m��b�Z
x��� y���u ̫FZ����� ِ;3ށ��� ��ϡݥ� H�\���3� �&ZW���S�L�	��@��[ʗu����; ��B|��c���1��s��่� [�j�/Q޶�$>� ��c�!�:��[h�4�%�"@���� B��ub�}�f�R(`W�/_l �N�-� 5q�z����*��2���1��4��}p����I� �ٷtWk� �
ޝ`N�K���0��� �f-��; 1>!�' `4� 2(H�dSX&8 �� ���	0�{K����*�H���o�Y ����������( ���0��) ��J��@�� "���?`�������!���� �� ���g}e��t2��� ��3�f��!���w]�� `�R�%z(U ������� ������ ��_S�2���; ��^Z� @���#����L��/X�P�y �8�ȓ@i O�~N�/�� Q_	$�]qs�( �v���� �%̤� �/���B !�l�"��@Zk��
>�l�N�@�Wp�s iIղ�]��[�9FP�W> �n��J0!�X���hAbQ���c쀼�V:� ��0 � �/��D���XA# ���ʬ ��=
�ﳋ(e8� �Y�P���|V #�TjŁ��0�K Q8�h_� O7���� �@0�I�Z8e�. � �c��3� Q+�k�p ������� �"�Q�� �D����z��N�^b�w�AI� @'S�����i�ApL�>�1� NK�� ���öC� r(
�� t�`qA���0�RE��7\p���~�Jz25LV�?Ȁ�А�-�9]���{�x�����9	R�q��ȧ��^ P���X���鷗�g0h�t� P��N��IS �}x�����	�J�����N[h (	���C�% �������} q�^+�[�|��xT¬�P�� Z���^c� ��f�M-�&���>�� �]
�Q)�U�!b(d�x�X�b�,���	0�� �ӊ:fЂ�.��s�"� �XOG��NIqJx 5wu�� �4��� +�b�^�<X|�(-.�!����B�r i7�Ӭ%�� z,P��B���|��_� �a
 0���y	� Y�4���J����F3���`��itI/ �S�	{�&q����+�s<���`�UGƏ� @�&�ZfzJ ܡkW�� �	v_��� �1�LXI; ��A��� ���8�h N�c{���< p�+�?%f 4#��	Mw� ����� ^h���M?[x��\PTX�R
?��2c@S�(�-�'��I�p �o�a�9�D��(p���$�x��p�D�%�!��� _a��(�^�q��.�*� 1AەEd!+ >��C�)� 1g�w 6}\��0� Z��h�K �X��U���� \��,�Q��0u6�7���d����_��t��'@��1����� �~/�-xy@%��\ �ƣX�� K����!q\z�g�M�P�B�)ʂ*ɀ�+��� ~����VS�G��y�? ��0�_� QӋ3ae ��ԤX@f\V0#TZ^�֗�?���H�n� �<�v� x3*�o$� ��E��ע RW8!�	���+��_� K3��¿��H\��S�����K"�q��j ���-: +�	�ڈ Á���"}m &B��A�� �k�0^�*o ��Ġw�,_��6�sk žH	��������t ���K�E�ᅥ��������N�@*V ��3Y.�t �<�2�X �֩	0�We [�g�� ]�hΠ� ��eL��� #��G���w=�I�]��[
�`DV���� ��\�h1)^��mvM�̦� ٧0͐�<���H(A,T] �V +�!��^AҰ��0�(Q ���-R� sid+y�_��:��k���̏�� 1 �'}@u ��V�&w��д����*�� J����HN %w�PS�Z���<Yp �[�0t�� h8H?��� �Lp�JX�" Y	U��A���2i�[{�'�� ��-��b�W x~27�(R_�F%Ps���Q�� yH�d�6�-�oI %n�� �> ��� ���ҭ@x~� �%ش ��s)J��( =�б'1� ��ZRN��� ^����_qz@��Tг�Q�� ?� ��'{%� �hq+� a�@C-�� [H�����>��<0 �2Z��X��������W�U �bؼ�0���P� ������l<���p�D �"��-K�a����� R��%\�� I��n�	pF�� �&�'ܗOɠ�|�R*�a���!�LP��8�	���R� �K1G;>���7# `���'� P��JV�f
n����@q�W��m!�`hKI^5H˃@���0�o��z��g� ��r�>��Ÿ�	�?H �́� ��!\� �1�� �	�hd�BX,J9�LF1�{�� `���Ȑ )*�1<�- ,Zv7X]"��Qѹ��oԲ�� *^�����rK:Z����u���� �H>L��hS w�%��߰Zl��v�̀D�;A�� B4�����Ÿ� ��.?��oLǌ	;gA ����}�Y���Z�u ��RpcI- s>"�t@\Wt2 �d)1^ ��M�'� �&���Z Y1�~��.�9' �J(D�-
�7���)�YG���s�_����VT^�<�J�v���H��Q�������b�<3� O��	]�����`���ܟd *ꉲx%)�pCO�� `j]+ M��ȭ�Q�����к�����TW ��S�ػQ#X0���&�.nՠ7�|�E@��s���,�hm �b�^ B�{f��p ���	�~�<V������؆�JT�R�x��80tVB ��x^�)�m_�쉨TߒA @@��!:I�"<Ea� �S �#�P =�B$UZ�X1w �@�(ÿ� �əK�?�Vp�:3耀��i�^��  R�b$�C:����0��v0!��Е� �3ûeHRq/�S@�ۋ
?ѯ#�h�[ x�6����$���AY{�L ��I)/�9 
���U� ���Y�\P��h.g7���e��$ X�6�^= �4�7�
NW �;p/�A$�J<���|��bz� 1��y��P��K�� h���}�� v �ǧOA �?t�_VU��X��2�6�����P�^,�6?[���59 �&������Z>`_�p�0��@��~�XYyD3"����Z�Gm��L� ��
	�Q0L׹w �I��u�1 �,�
hY� �����^ #R�!�f	� ��������'�_��1���N �z�"�� ܜ[� � �04�9ٴ} 	T_[B��  ���Q'�� �Z��T��� �R�L3/[ ��K��H�F���P����)� �3>���ү V��0�Ǌp If�4�2� ع�8�'^� �����%� f�`�_���r�@h1���^��+�Hf ��R��A�9W����uB�p �]U(你 Q�	�{D������� ��CL|+�[v������ tB�m�؏�>` y��,~| ��9����3�Ϊ�� ����p�N^	����n��(�,��� [�?^Wp��t��d�J��5v����%�>t� e,X�#�2���ۃ	��� a����@����Q�P��p�F n���$N03 ���c�� ��P
Ÿ^���~eU�WZ �	N�L ��,=�" ��ݷ1����C|��ہ���("��?拥��5I<-�� ����(_��@��5� �Q˃�t+��[��7�� ������X�� ��RҺr&�� ���� P0ѸM!%�1Ů_m��Z��O�ʔ��D�7��o�$r3 ���hD���tB�s��U�0�ػ�� ��;�� �f RX�tb�� �Ք��ۙ9 �ֱ� Y� �Ё�P�� !�XZ�E0��*�6k�;��i�y+� ��*�L� 0��	� ��H3P� ��^w��� ��|���/≀��#�ư �6�2���9߀m�wZXu� ��	E�다 ���ŶZ}y &[X��P�\��	�Bڧk�h �?n4�� �ǻ$�r� ����|�( 	h�b��d ��U�_�� �x��-K|P/����y ���(ȡ� Yk�npZ�"�@� y���N� BXh�|�F �t�ݮ�Cq��$�`��6 �cˡ�#p��-(�]1�/��K�!���J ��*߻ ���9�/B�x?� z�4C�, ���8 [ �'л�O�� L�9��B�� �=��\��u�6�1��z� �R
,��!��� �f�� Ø$��'�� ^b����PI�� ���hN0$�:\�1�#����V �,��K����q�Ai
A�+�@��~� �" �� �e2�.1�U ��:��dM>��� �L �X���\�C} <���v_�vZL�� c�O�:�� ,���`�Z��	�N�����S���Z.��ň�������ݑ�%v�m!�z}G ?����h����` l_��U*��?
Қ@Vaބ�� c�Ϙ��>�1�������%�y��ӵ�� �X!\�Q-_ HP�^4 8X�%0� W�!�wP���XK�}�^$y�3�}~ -�p�Q�������	c� j�`�[( V �K��� ����sBG�p}w����?�� ��P��Z ��z1X��  ��Լ�d��>��Q�� ��'`&��~@c�B�q� �e.��X� 74Y�)(�O+��ˁ���j�	��׻�&�0CK� �
	�o�-��A M.�� e ��h^\�� ������� Ӿrd�� ��t��kH �@%�EP* �>4ǆ�)- ��_�^�u�������VC� �>�0m�.,�LT$ ����d� � (����`$P��X0�UW��#���CD�] a����) ��?�x^ ZD��1>- j��!�:�
 ��a�R � 8�F�3�^ W�]Y! 蝢ʶ=� �
��m�;E(ɐ3�p�P ހ@߽�ڒ � Թ};� ��L^Ь��j�4 ���}m�_� YX�L� 	&����%�ꤒ���?3�-2 �� �A����ܵ ���ůȖX�\��0hP�R Y[4��Q�'g����]�� ��%b�u �a�qL�� v6������2�O ��$�Ύ. ,��FXa4 ��K��S'Lg�x�'U�i�{��߀sF�d E�ܮDx� � z̺	��d��։ B�|���W���3��~ !tʘ/?� �@���[ hK<!�"���)�U(��0��\x�,��$�#�� �ǈ��}� fY(���b�0�w�p�- �Jc}��&3 �2�����	�hHj��_�SAe�&�g>�L�� ���]~� 	�S\�R ����G���� +��z�Р� h�T��N$�a| �*	�R�eز�^���� �|K��sZ�x�k;��| uo��7��y����	�,?���Yp��h J�A����B7"��T��nx� �s���F�' ���A�� d�H�|�3�ڎ�)!�	R�p{� D���]�b3��ݍL���°�_���R ��N@`[�(��� ����?� �/�_���* ��Q�D��L ���9�^Y 1ЀǸ��+ۃ��h�R(o�5ʅ��[�m�%�\��;�4��ג�`�X(���=�ʤ �D�/���<����Z��k�@?S���Ю �B���]\�� ��_� h�f�@�K�?�#��}3+�&���$Z`�JD�qG+����' 8l��3� �H�k�	Y� D �Ձ�� �=M�C�Q� r]oq�1��w�#H�$_�����v�=�MN�@�� ��X��= 	�vd ���0$ ¯&�_ ��(J���@�{�����\u| #�&�� �A���@$n{`��H+( M�'�O�Bz� A�S;e-��:�Ջ2K�.�t�Y�q.�M(�����yҘ���Z��`�1	�W�ع0[��M ��I�+ ��@�ܥk�� nt���0Ś<N �u3
���) *�×�	�dͮ��Qi@Ɯ��aHD���Ĉ��A����4��	�̩/��n����O�x^E hWQ9 ȧ|齬= R/)��WB�U�;o���� $�Ysa9� ;�*��A� ��vg'�� ]ǲa�V����R���r��: !�Z� �5��z�}�>�X*�Lf�+��k����`
��n� ~_i�@�Z�Y EO4]�)�ť�5��<~�%���;Q�X߻F�7�����P˔��Ȼ��j���$R^;�G �8y�N����[���%P� 0·U|<�� r�݄Xǫ �ӕ��=��]���2���@�\��!Ͱ��� �8� /�9*���� 5�2��>�%/ �O���4 .�<������E 	�Z���kt�����A� }��
�Y"O �Q�I+~�q� ��P��)�|#�y�r�,��e;�����)"��4����Z�����Ց � `'}�%~� ����K��Y �CV���* ��]
3�\ )�	@4�y�Ι�i°��o `�~���Mv S� �d+�0���q� Q�؂7�W� �?	�Z.�� 3Y*�߱(� k��>�- P��Ԛ�Lh�1 ���J� �'�}`S�W ��RU�� ��)Q'C�� ��H]�F������8�� ��Paʸ�	�q����D ��)X���\ h@��N�� #[��utO��	H��D6L���(�LZ� �O�`�� q����,�����``� ����K1��n��۳6ZC t�h��qr��� e�0_��m� ���f�\k ���C�H�X "m��	Q��z��`��东 ��[��շT鱣f@��h% �ry�}��s� B#�^�5 �Z� ,*�Q -��_%��inKZ��QD[ ���@��1 ;I�Ъ�$Z	G`���0�� ���T����tV ��oP��U %*���f�+ �Q�й�_ʕ�`8�K��ڑ��5���`ϰ���<<���!�.D:����� f=�eK �����0`�� �����[U� wӯ�� d ���P�f� 0?�j��W���Հ��_*� 
���qׅ� ��4���P-��B WL����X}�"��zA�o��J �l>��?� ����-�� |�/՚�j�v@ ��_~#��0�\h:tP��r �p��yw ��Q2��(, �.f��#� ��o"7�5�� � �S�QP�� �!ـ ��[���c�u8m �b'����n�A }i�x�İ� j.CL�� X��'�O�*f֖���a�!Ԉ� �	b�h�� ��� .� �m=���+� ��O3��qD *�X0ҵ!)zuQ`�.���U�2 hc~��J�� ��3�P" �Y+Es�5_ ��Ƿ)�q� �]�/�� ���A I�Ϋ�!��(����$~���%���.S0t�� �/�j��(U@� �Z�D;�\� ����4/�� Q��*�|N 9V�Sx�� �+���}P �EɃaL%4Y��,�P�p0� ���+�n/ ���r�� �����(� �4��sX '�^\�K	��%�q���j�x�L���_	��:�}�� ��	#��
֧������ D\��?�_� ��%y���,�#(�� Z��~�.n� JĒ���� $����K��!����s� �e�N�	����'Jԣ��� �Q�S�� �V��Z�aJ ���D5�" Ы����� `�1�h-9��Ϳ���$zK�L��ط�����`�6 �)�`l�'5 	�8T �ğ��k���჏�.Za;P� n]�W�0� �lq'
�� ���Aٔ+�����h	.� ��Bw�t�`ˋ3@�X 4��6�I� �Ն5�x*�?	� ��:� ���[�� dF��TV��*�@����Zvy ��-����%V{�:���`| 4����� R �'�x��	3@w"�����F�@d-�R��0TU�F�;`fXh�\� ��ͫ*����C_p��� ,M��LI�^;G�8/��v[��ր�M�Bu�O6����� hk3��ģ	<� ��%&�A���B���X?��T�U�X�Q��趖_!��,c{���� d��*��wTy�� �����o?�2u���� $P�,H�tZ�O_�څ}B� ����҉ ��j�4��p�$ QbV!�|� � \�(��� .�BK�� ia��hv�!\�� ���� ��ŉح{�;M��:>Ψ��9��`�!pJR�/`�d��G [Y0iP�(� ����fT���夀MIyo ���Q�J��+��S$ �n �T�
�	� -�Gl�  �U����� Z�<�nWP�
��}�R� IO	�*!3� +��ZPYSE��r��풵���W|n	+��Loړ� $	�
�YW?����զ� �=1����?Hʝ�T� g�ڟn� $�^�B3(h�*�����٠ 0�M�~�q� 	�z�b� 8�g����� �O�a�X �>�fR�v/ ��������;f���0��Ӯ �RW�@t8�ZXG3�N�L�X��غM 7(��! �f)��� ����/��� �ǿ���!��8�1�/Vε ��JU����wy �f9�&�'_� ʪ�� Z�����P���ώ�ʴ�kg' �ښ����^QX���� �Ǳ6`��� ��
S��� )�\UP��^�҅O��� o����J5 ����9qhj�Bfh: �=_���T �	���������C ��� �-7�\"�? ʒ/��� ��,Tr�W8���j{�=�'�;~(K��[�N��� M���|X D��K�_*u�c�Z (r:�u ���� ��^��/ ���W*�Ű��Q)���V� ����;� :��r�b ]1�%��yO ZB��e-<�W�Ʉo���� ��N�)��<�0\�I��	މi�,C����� bp4$"��<B ����j�~ �f��X�* �ᜋ��!��] #
���3�ݶZ��0Hp�R=Q�KY��B�� %�X@�] �	����'� Z1�Q� �>� ,�9�k��!�!�؉Iq� ;)��p+�&N���l�}� /8B�� eX��G� �0���_1�  �&֘
� ��p���3��z� I�)�^'0��FDdu�,�u]=̝���.�bR�Z��X>!��J�-<�޻G���;��p�ԟ��:�<�����>-P�d0�Z��_�}@Q� �@��ZQ�YP'��	�̴ R!�q���� _��ɐ.�Q!�3����N%P`������d� ����6_ ��c��>�&ȝ� w�`t���Ca.� d��BH��q@%.h�v5 o/�{0��������w��(�=	 �W�2 ��p@� 4HV�Z�j�! ��d2��	 P�w��(9����RՀ_m�� $fkq�T ���A�L�G�_�����>� ԛ�@�N7 ��,�QJ1�Àa�L��Ҁ ��XrY +�P�������N�����G�][<î��,��`�qx �	�W��;
K��Gy��l���]~�KV��^1�����SOO���p:}�	�� \��'� �l_���T
��A� �{]� '�_h���&�e`�V�ߓ�4�E vZp�J⺌ R�*��b� �5	h��� zc@Hџ� U8k�=���ȿ���˶� ~��	Zx �$�0�X� �^YfR��ʶ?�*� �<��+�F�� 4���Һ ����N^q� �0�� W�r]c�\ ���b�'���^�R�* �q_ǭ�`�� ���;1�>p� /!	�S�X`L���n�D��	^.?�3 A/���@�$���7Q!� wl��>�� O����	�� �l�b�&y[/#���±�C� ��hbH�1�v������K +����! �d������ 1��Q ��A�%q��)�; ��@Ѐ�Z�X�y�ɴ�2T������ `P=���cG�04��b�6��yH��@�� ݝ`0tO�R-I_^R�� S��hN�
��@��n���_���s� -���p�h��R��;& vGE�� d0�U���^{)����$a�W ��1N��0h&`�T޹!��Q� 

�/��9B�,�@��`��7��0��' =����D8� 	���� MP�W1ˁ �|���:�@���� ������ \]QeK�f `Y��򠰿 �������(��}����V�Ԃ�_w���'��=�[��Y� Ɓ��P�ӆ�h �dJ�3(
����G�^�/�!T\�2��C� ;V��^t ����\�* ��h�#8 �Z����ߟ� Ŷ�8]0� Z��¿5� �R|<�ݘ��Cp���
_ (w�ad�� ���	�� P�)��<�:�.��S ��hp� P��{��'\��G$7 S��g� +��O�At<�W�8��<� N��s�ڔ��-�)�S�pzN
�H �ia�� {·�v ��L��:(� ��݅ruK��xN�S?%E �/��e�<&�� g
Э��].��A�0z���Q ����1�� Yؙ`i 6L������8ğ$���N�	�a1I�T�(� 
�Z�����	Ƕ�.�`;�V L���S� �3����KU{� �khmc9��pi�vF��@ �a(�\� /���2 �cC�)x�>�� ��=/1�� �z�H��d� �g�-2*� ���_W�N?�j�wL�A�h�� i�g1PWz�����jG� �ː��[gY8�PS ��_����L�0��Ȁ0�$�3� �*Z� X�n��Ҽ� �dD��LW� O� E41 ^����s?Ҫ���@Y/��"��【Px2�?�K��0���,�J@�1뀠%�u��m��(���[x8���|zf �lC�b �+�m��r�@����Ͳ��)�����X 7�	{���A^���1옱�3���N@O�&h{.� R��?���� ��V0=�T� {$Ҥ+�]
t>�<� �K�� +^z0�R- h�H���N �`�+��g #�f�� �	1��� Ȋ�8I~�N ��(R�����[@�V/3�L !�E�1 �A�(�	, �����a =��>�D�� p�j�Z�o 
�ඹ�N  �h+t�� ���:����H� ���>��'�x� �@v�L���B"��Ṇ�p�fZbN���~� y�q��TS� B!G;�aИ ^�E���� ����Ya��?k=.zG���Iu)� 7��ϋ^=0�X�������eƮ*��` :�(��r�� �+2�!�K	|J}��(������$��ȇ��x@\S��� Q-�UPl h�j��/�~ 
'��<߼�I��KO� ���S$T�� �Lh�7>G�~!�� y��¯�<�����	�Uep�Y��4|�F�lB"���Ǉ)��	zK 8�a_ �,g��Zt���]�V� )���@� qG�%)/Hro �21�;��N D�S��m� ࠪ' �yr M0+���&_��~�u©�1�� 4�
�Z�� (r�/fc�9 �ل�s�� X%y��!�= � �S	)�qd�� n��~^��l @��K�<��/��&����Y���F�<�� ����ʧ 	U�d�L�y� ��K�0]��ހZu�;Vh-KP+	��H����� (_<E N��CvQ�� +�U'�y@�\���W� !�@� ��^�b��>�+�(z��`U���XW\) ~����.�����hK��� +[�G�(�Ύ�����f���� 3q�A� ��o9��>s� �RZf��>2�� '�]"ܻ� �c��Y�>1݂)>��p����6 n����h ��S�]�)&
�� ����% *�3؉�A�X?�O��si w��z�.� $It�b��_ q�	��\W&�
��n�P�@�J���gҀ��@6X�d �Q��Z ��ւ< ��k�KE� n8���SLZ+ _0��]�n��j�*�! (8��õ��@�߀#P�Q �[	�y�T�ɫ���w ?̇CI� ��8�@���	��`�!��A, �y"@-�8 ��p�O��	�!ŀ�[%�&Z��� n�����] ���#uh� ,��Z3��>�[�Y"� �մ��o�~�5�;��G Vތ-��oX�	��;Υ! ܁�#�Y+�;�	I^��t� 䨗Y|X! ��e��-6��PL ��ΐ� ���G�0�x ��o@{�j�&h� ��(��� C�[��ʩ H+)	V�}^������0( ]�����@w<�O��W���\�Pz��������Ym�9Z�d ���	acS �O@n�1� �/�ZX�?g���B ���K�'�& 2>v�A�>��ͨ ���PU� �d�@<� �sML՞48H�� z�Y!����ҳ�/`�j� ]aqX��& ��:���h�@ 5�~O+���� ���^�JP��%&�X��<@�-H  ݙ�?�� �`h�R�?���*~���% ���	�U�L,���b\��p�U���&��HO3� �Y�y���,r~� HɈ�ڨ (�iؗU03&�� 4���� �V�"�ф� ������\HcE�`��X�- (�ѣQ��w�.1�� ���b�_ �`�8| ������)���5�0* ��-�e+ �`#Uo:�3/�>ǐ�I����<����� �ȼ��P�� [�v\�ۂ ��ޞ�5���_� 	keի/ypJ� ��ә�S� ��Z�	�У� X�Ky �h/_�����B��[�� ��p�h�l� -q9��w ��	��\P.,� ��"�h�J�ǅ����4 ni>Z�f� �_�b`��P N����9�{8�� 1*�謖 G�(�����g�]Ѐ���2� h�.0F�>q��K�� �b� 8Yh%,��i ��yQ|`ݖ�#}��o
� ��2��Z���I� $r�M�t��=
���P�F` BU���n�.[�a>'����`�0�����J�=?�rەA�2]`�K ���: � %�iZ� ��$��5M9��@-&�bVe��y��1���\ XK?�M�O�l����	���No 䐷�.�Z	Ԟ����1lh�����+ b����� 1�h�ZD� ���*�a�x�� �3�[�� ��z>��O `�Q.@}�$ͭ� ����*�4ӫ���/�!&Y����}��j�Sл�K%������U} ^m[���x +�P��L'_t� X0��kA 7`�C(#��\-�����V�0� �aQ��iA)�K:�z���l����-:��Xc�@��O�t>�v$�[��p w�S'����%�� �(-1�� _��C�R LpkFK� ����aL"�Y7�(?�� �j�G � ��HC�5��&�d�s��P K�U��+� ['Ȃ
� � /	��p ����4Ĉ߬`*�Z)��h�R�#� ����1r >��*[vg K�� ������ č��#Õ���T���P ���@�#�!�z���t�n�X�� ("�E����I���3 ��0ݠ�Z�+h5\^�t�� /ˑv��! �
�]���#��i�q���P���p��� �~WX(� �+�O�{ �.h4� �~g��Q��dO �_����	7̯8u �x�$h �r�"��Ć ��a�W>�,����JI(�Q� �*�m��j����ܙ�pu�@����8^�1H`�@��	q��@#���� �^L<��1��	�K�� �w� �tGS�d��~:�����\��ǰ7�0 ��(�KR 1Y&�P9Ls�~0?���*��AhZę"��a6{<��� D�X:5�� �%_�N� �g���+rK hC�O[��; �1��!�%=�*?,
�5���:N�0��. `ˀs�F�� ʸK�=V; �c����� e���� �O4�u��@q� P5��ى!�� e��#r�P��<t���_f�  �SU�(F����!ۼj�N A L�FO�$�k+��*w�� �Yp�r�8(��� \���[� 4�	�̘��U�]8� ^5����W�ݿcm-p�g @��R\(������Wo�n 5	 �R��`��1�ڂ"��a�
 ��.����.��GyN�����V���k��`8- Xs�/�
� T.[ x�Y��z	���F�� h���_�*ҹR�1+�� ��e B�J�b %<#�q�x�	���� T��]$ T Y���|W{&�vz����ہ8JG2��@ֆ��� �淓.�I�`�����e����W��%���ZP ��B��F� �g�H%ak\/�κ�*1С&�� (��'% ����n� �EK��9rs� ��� �ư ���A�{�,��Z;���	�� �ԯ-⫅����d �P�TX���N�`�4[`� �����Єr�>)� Փ��^A ��6���O� �S@ѡ�m|	�!��#�9�+� q�����n� �~��*| ��B�IK �7?V8��� �b��HQ��.l���0������>�����-��R
�B0��[�q 	1��D�� �ēS���dQ�j��s���Yz��4� l��^�3�p�X Zh����� ��&c1�2 ���Z��a  ��@�hU� �!*+��7�-d_��Q� ��#?���^�<���λae�y��j��� �F�tJ��z �SVR`� �՟.뒬 ��v�%3L� Ё�Sd����Bn�U�� �Ƽ	��� 'P��i�y p��l����W�� �n�_/F�H��I^��
�����@��p ��t#��u
 1A���:���!H�'�T�i 3���0�XA����`f� Q�B��'P�]>NA��/S()Y ���\Z� D}Ep ���?����d�%!���	��m���� �8���C�w� Eh�]�S*� ��#�Z_X� z�P3Ü�H�? ��+��p,D�H��	�Q�z�f�̒R�� �,��_�)C0 �S�R{ 4���N�# `�0&̓�� _�bZ����߀���ԓ� *�)cф��LX� ����� P�	�W5�Lw� !Uz@|�-���+����Y�5vJ`^6� �,m�V��[ 	�^鴿�~ka��?�J�� �BY���2>Uڻ�ߚ4�'��s�;Kc9�r �'��bH� ����2� 
[��8�	r ���O��� Q��y/�� >�%~Т� K �U0�� �p�?)듭 ���:Q�� 1F+�k���� ;`��#֋3���+��j@�'����^hX=1"�H 9����
� *�!���"�^n$D��� �	I��.|V� �/� `:����]��*��Y�0X�K 1[b��Q� ����f�	ULu� ߼;� �'�����\� ����6�R%�Y���☒C�U��y�� �&W��b!�pJ�� cU�� ��R�A����u�1��}�� ��fa	� �P7�=�0?�� 5����.' �~�o��&�J��h� �颩���\��r ۖ�@�A kB����} �*�1��<�O������`�Ϛ�n>`Bh| <b�DL�?�� IUQ��iv�%  ��j�A��\_��,l �Z����+��;߁��^��xL "�H1��� eܡ@���[����: Nށ�h9D ���l0�� ����I��H^�[�;~) �M��b*��_SU���w�\]~ �ӡW:�� ؗ�4��R� C��h2�L ��]g�N~�b�~���� �͞
!�R�<ޫ��'��0q �	����?��|� �j�9�2! ^Ѿ'��-�Q����t̀/ M]$��� "H�J�N� ��W�]ue��B�^9 �gTi�}� #O�Ԇa�_;�Z�/�M �0�Y)�X]s �2A�U|6 ���H=� h�S:�AZ��� ��e��T���P��O8 I�徭�n��NG ��) Z׭O	f��;�}y>��q�+��, ģ�p����C d�P�-s� �>�̐zI ���%_Y2D|6 x����E��X; ��ǧ���ėe�@�/��� �!��c�4������$ ͌X�P�:4 �qw�j^ %G�eW��� g�2O�E�� ���S���		�(��cׁ1�82ˀUEd\��h��C����3�`� >"��OG8�-@@5�� Js�r�9l��'E����ٓ(��#͸��X��[����`(�k��i��"𲪀 
�S Ʊ�2��٧rOP�a�]�� �ް~� k���{�<LJ�Q���]p�� 0���@��8 �A��{��� *0��L�'��Ձ2�ᒆ ��ߗwT'Q ����a8� �j˴k C��Y�/b ��	�U< �$�NqŔ} 鷭��I���"�v���$y���us�)��7��|% � �f��Xe)%��*��ӈ� Z͔UP��$S��p�-��P�� ����w�z���z�;�����	�2Y-��@Jըo�# ��R�L>� ���d�ڝw HP�JD���[/�2�0b��uļ�ޡ�"�#��TX��$�}� �Q�(Z҈�&�-� B܅���D�|� ��M��nhK���'�IHΆ eC��,K�[%�����T�`��\1U ���B��� ��F�.�A��� 2u�:\�R�M�j�J����$���@�K�w^h_"��@)� ��C��6�� �#��&��$ ��@�hO֩ ���E�2Z �3Q��� b�-�#%Y:�_�|��A`q���{���lԕوb)� ���x��v9�JP��%���@3(5� 1
�i�W /���8 p���N�h\ qi3A� �%]��� {�T�	�oʐh���S3 �U����e�v�=0� �N�V��;P)�t�OB��>_ެ ��S8�K&��4 $�(pwB ����12 ��!��}v`J��ҁ W�y�$�� ����Q�D��:^��S����K� ���'�QJ ��Z� ��h�8ɺ /�0ofp %�hRe�9�VIt����� �ȸ��S�+V��x���� ۻ���Uƣ���yW� ����e�i�F\t`2&�] �	�!��h ڟ���y���<������9�� ���.��L��\�h'1ш��� vW���(BE��dᨏ@�TW �M��� |��R[-� �$�4��\� j`��� ���* 	��=�AD�n0����6㥰��#������?"��߁��(�z o�-��%<�`"��Y� |��X_�� �� ���QV
 �L1����^�%vd0��7  G�ҕr�)�/��P� QDW�X�z� S�7��h� &��0�P� m��^X� t�툂O��M�� �pd� �ɤ19�Bv���0�� �h����3��GR��>�MʀC�듖 �ȯ8�, YPZ�z�� �B�pE�k�q�����	; 4�1�)�*�b\�@�v5�����.
 	�VhIQ ���P�f= ��?	V��� ��L(�8� ^�@���aW�o��V���`{� K���U�*̍�/�p=wւ�1Ë*�AJEC�� ��P�崨	��T���.^"�OV���L �; .�W�� 3oK;�	Y��F�E  l��.=$5�u/� jU��% ��v��Bo(�$��s����|cJ ��TZ�YL��d ��� K������|j��%7��(���`��K������x�aՔ�N���q� ,�*'. L�=)[ë Bj���� ���0�n��� ����|L �[���X� ���	�Uz4 =�]Z�`$}o� �^��� \P��?C ��3���۫5�n��\ż �f
魠�x �^�́m��.�i� ɝD���ܺ�}S�>��]\"��8԰Z|. �V�(�e�� *��C]B[��!n�⇨�@���^ @0ðĺ �eK���HO~"���z�X��&�H��@q�� PR���Z  ��i��� ]˺^+����V ��8_Q  ��=B�}��n� �>��(8 ��;� ���`OP���?�'K� ����J��ˠ8�g0u XO΋���{�������Z@g�-��
K�7	2 ��[�C5 ��*`��p� R���V�J�>������A��8�����Q-��h� ���"�g X��Z��P�͇�U*����?=:z|J�c���h  ,�!@��X���o�� �Pa%H�2_)�G]����� �0	�g+�� ;�ET'��- G�h���� "�L��1�� �H(R
Q������o��� ����z�Z�� ��V�īD3 ��_�Xk, 8jݻ*��)'��޸� ��f$����v��Z� �B~��H
����Ww�^���- $��{� ���H�w�Y,*���(i� �zF/?dS}�h�=	���?Q[@�%��	�uT �Ȫ�r y=�\	��P$pS�B��ws�~�0X� ��A͵8 L
뽡�^o 	�u��*/>R�3��2N��^̈�%B��� c����.�&� �sN����� H	�O��C ��˹ &!�]���� �VK3�r�}�{#v��Q%c���{��}d��@�lR.:	� �o���p ��+5��� ȉ�!ف� �����[B���8���5y� j-݄�ն\<Z�,����� �K:W�y> �_�@ ��j8��.R�J �?�+� EBMu^��� �I�� �� v�0L�[�K�� b�V� �Gdu��� � �$_�iY�F�T�� 9�h�2�J���`�+(* �i�NP�� ���U��� �h$V�� ��P�!� �8{�gK�f?�= �S��RLM�X^�vt( fg���U䰌��^L�G $ �5)�i h{�H�x� �k�A�&C��p.�)h�x t���b3�� !s��j� � /���d	=�΀�c�YC�# ���1�P�����w� �B�.�d���L2@ �p_�G�I0�!���[�p�Q�+��p���f ���k��� "'�D��$P���x0 �&��� ��ё��. ��'+ʦAm �x�J�O��4��w�T�� �.p���� /B\@ҽ9�=���K8�0J� ?�P���� Ţ������ }s�ۨw��~B��������� �J�}R' �][n����E��M �G藷�q"�'��u�	^�Ț�	%��~�e7I��/��������* W���)頩����� �P�h� �Z��6/�	���`����Yk� �BIW@~! z�
C��\��us}�������@%�Ե�A��5��"�>;� x���&Y�����/� � ����!� [Sh�D�`����^
��!��S� ��E��z �X@�ؒ �~�㵛z�[��@�A(� �^j��?�_��� �sˉ�>
 ���V1�� F[�ʰ�K���r�� ���G�	� �AkU!�{�F��;�rI;�-����V���6P��w����] 8����O��X{�2Ӌ��Y�X��w ��^[�� �0�ڶ�%�cű�A�*�� 4�IO9Q� �e
	oZT� A���%=�V��� M���݀{2X�[f���{\�# J���SX ��5G3�=�^���S��:��C
��| �K���I� 4�kF%Ť g����-Ad �"�E�t����xk�bh� _e -1�R
 �˺��K]Y ��� `\�p��g /��u@� k�P#�� ��%1��o� )�^�a��� �&W��� P���1H�� T�]���5� ahz�U2t�  �
��uF� ;��݁�+ �t�3i�Q �@��U
�� ��|9��{�P�q��=1#QA���"� OU%sՈ� Z8oK쩡,�� �?���� n�0ר�	P��X< � 3��h-r��F��V�!T3�j�`b� 
+�&~>!_ �2%�X�� c���L�*�ې7�=�I��o �� ��H;C= /Rl�^� n��棢c��q� ��
�_���H`�L�b�Y T���-�� y���� �^$Pd?� �!/��%� �� ��8^U �Y�z��I �����*" :��[�}��Xg� W�-�@XH�,�d�C O0ܓ�Q�� ���B4jr@�� \�R#���Z �K��ʻ�X��P��u�uW(�	� x�^Q� �?�վ�v�-@_���	Vn�	è�p1 �H������h� �]tY� ��!>j��:�@��	f�v��e����# )�[��I��� r:P%��� ȹy���U� �$N�<�� 5�B�.����J���0�ZYp9�x���-�]a� �0� �+�~�5'1����kH�����@�	'V�\�1`���#N��g��� 4�;� �@܀'��� �_!���t� ����+�$� ��1:�� N��g5=����]����%�b��G��!�t� Q
(�5.�>�� ߅�]�)[?� _|�a���8�C<��� ���r b�
���� ��E���z 9�LF� �� ��Ԑh�t��1����vI�� ��$#1! �����}O z���L���Ka� �n���� J�(��� ��b��^- ax|s�@�X�x �!�5�9���ވR7�[�+�� �A.��%�� :�uT���H��;����y('� ��H@�R��EUq��X �N��	Z�uPU_�T � ���� ������ r)	R��3�`�< 7�r�]@�_�%�����-0 	�X�8�h�9_,����1��flؒ� gW���N ��X+' ���x�!�r ����D� b�_ ��J�z��C\� �ht�m�.����bW��� ��Y��4��� ��`WtP�=���0�V`��(^ #��o�.�6 �ˁ����n�����pC9/`�T1o�,~�Y|+7�ց��ch�� �ɖ��X�Q$ ����&e�T<
�ʰ�S�a�>y� =B�W�w&�P s���ŘD��bn1 ���, ^�=j؉�z� 	t�EPY�" 8�'�*� ������O 	��`EW��� �c��� Dm.�>'����<@yy �[AB)
� ��\K	h� ����Ѻj/ D2}�0�p 6�K�Q��g�Ӵ�O��M �<Y	w+ C���`��$�� G2ї�� %���K�. ��WUf��ǘ)]; �=���](� ����On�=w����Ma P�-�� � ������\�� %X�f��<Lv� �P�cg$ h%����b  �FaP����j����B��e(E�W��Mܰ բB��P �?R+ں� m����'�� ��]	W��O��GJ�ܠb�
�,��K�Xio���\(���}8��˓�@�
IZ�� �����0��®���`�� �U(�V�; �>���3� 1��c�!M�\G�(B0� �$/�-�!ӽ�K�ɪ`~�(�� ��S�1i�`��� �� ���>$1J-̫� X�2*� p��7�a� `Ɯ'�W� �_���y6 �$)��� �X�*<�=󽀻2�0=�` �:ñ��xS�����	�D
Ha��� J���v%���B�lL��0>0b ������«`�@NF�q� �a�ʼz% -���#� _O���^�� LK�]~�	���`D&��f� �Iqw�!� �(�%�� � �_�kʁ�Y`vd��. �P���� ���6TÂ @�['�_+ �ڄ�ݖ���6� R!x�*N Hص��	3� ��U.p��g �'/����, ���!�Z�
�h���\��I=��|dAy��� �L,7���� �"�]� ���R�2`^ ZKS�[ƈ�޸,� �1�����d��� ���P��2 S?_(p���a�h頨.��o�u �%b�wT�@��3 t���r��� af'�c��3��_��(n�+M����)�3��/����B ��^P�U&� @7'(�W�g �Z諬� ,��f�hn5ĕ�B�K"�� ���@��r$�F,*g�x�0È'� \�qA���$0 �i�� �%�p �3�Qͨ &��;�����"ř�}�X(�=��:L�>M �D�/q�= N�y���:U� bD�1�_ �`��=�/z� {W\�������X������j� �ǜ ��Tp�i ��0�Q�%� ���}�,���u \D�7��@ V�'�0�� �ܿ	�ԡS Ϸp!�� � ���H�b�x �D@�錉 ЅS�����h��n� ���b�= ����)�! Q�P������V�Cr�J�|% ��(3�� �x��B�t;]p�6N��\4�=� �3�R� ����O�_ ЬB�)鐺;�k\�~,^�G hR>�Y. �Ѹt��4�:8����C��$n�Ъk�rN�����K ����)E ��(I	�ܩ�1Պ �rQ
��-��#Dm����8��ZM���� �����k8/,Ws>
��]�f�$�L���|o� ˰� M� ��&�0��J�D���i֭��? �=b�6 �ށ��m�| N����4 �f�'��.Eo�:�П�8��\��BuH'~@��X (��]�� 4�� br� ���S�	�lܣB<P �O$����&#X��Y [�a}ڽ+� Pw^
�!�AL� =���1��ųa������ �N&F��� �
���܉6 _��ҽ�:	� W�ۤzr�h�K?@�$'U�0���Aj��^ �-�!�:�� la�Z��(�+� �-��D�0�|������1�V�X���� ��5��*� vt�X�n��?������>�t��h� 0���W�J,��Hu�&� O��}"�|�P����!���͟��{��� �����J�k�: {$�� %ՃQ! x6 d	[LNX�q؝�G��:H� �	�(�w 믤,���2�\ �0�Z�S�� ���C�� ���gAQ a�1�}^.<� j6@���� ��zپ��~5���@Ho��Nx�eb��h�@��:.�@�	v�RK� �W�5  ,&ZLڰ�)%��XJ�$h�K���T��pH� �O)�{�9 7��
ͺ� p�4��B�0(Q�DI���C �	:l^߯ !��{� ��6B��$�uT\NС98�Ӹ� b�+w� �����*� fpK�� �uP��> a�5���� �J�([�9}�L�����`�˗O� �yeƴݺX s~�Q�T�8�Խ`��}� ���V�4O� !�Y^���� +}�խ) 1�/%��C�+��!� �{��/1����2@V(���B�)��p�]=��tʍ�
U�1 *����� !.�/}�Y ]0�(�h�d��z/D��R�:�� �t���,P�K=���_����` q���Z& ��W��T_�������>0V�\�: ��8̈�銀�1�Q�58� N��|�� ��Q ����r@A1��V�����Ź�Py�Ɓ ζH��治 2���!C�� `j�\�N� ܬ���Z �����h� �]�G-5~�S� �)o ]�w�u(� �nfhg�J��� ���.
��� oU��lP ��i~���p-E�=`K�`7��(L%�0t*���|�`�q� ���B�UTW
���K@�����C ,�sV���@�)�%��+� �2ݹt�Zf �ԁ-:<M`[�'Ȼ�+9O���8A[ �����˚ :�h�CW� ���b��� ��!�P��������i�\ tVZ��n#N ��
����� ��X��.�@��[!���k+ �����c����FYX@l;x� g�Ʋ��� �(I.'>� �����&�
�D�@� I�����1����h_��~#��gE`p���(H�!2Y������K��$���Z�R1�/E�[�� +�6����Ͳ���J�d .KQ�0zPh?�T���J~�"�>ɺ̡0x����9 �bwAmu�MU����a x+���鋰 	d�R MKbLE� @~�XӀr���1�����f tZK��z��n�.?�����0:-=%�:���k�m��� 4������� ��<��o� ��7���N ����[��+ Zאp��LY�%��G@���\�]�+� �w? �N"���p �!���M� ��/Gb� ?h�\#�� �._B�, (������ -.�G���)������������.�?�o H{��	0U���/� �� �H���) A���2�$ wF��x�^��L9��z����,��(+��H YuG�� ��CPV�� �^��M�� �2
B���� iHeÕ[6� ^X�:3�7�}* ��#����@@�"��I���U����� =�t��-p �_�!Y)q� ��OS�=$fQ�0?|�[h�6�҈]�.��
�&����k�)��	 ��XU�P /\�|�� ��J�?o���3�T>��Gd���X<W̓����#��J��a y�@�] ��1�l�~[ ��k��!K��oE��: 	�SWQzx� �F4��� ����
� I(N�b�� �gD��Z� ��ƶ�O_=������'� \0��dK��2 /�Y���
 �_��	o݄ gh�{菈�Q�n�j/����ik '~O\�x{ p	�js�>c�Z��޶� `uX�(�����y�0��Q�����>�n��c�L �DZ!�f1 ���2ǰ�Ii;
��SpW(BR� *�_	� �0�IY�� -�t/��� 3w���C��~Lӽ䰑,�<� d�K�E �;ϻ��#�3� �*�	)Zwr2F����M� ��<��� �y`�V�*N I�T��F��;��k��� ��P�Q	\���F~����Ӆ�� ��a@�So� �����]� m:�p/ż� ��h�a�P�� �W�FU^�o���"x��D��vW`1l�\� v�t�"�� л��eZ+� 5�(켋HD�0 Y
�Z�8��^+�%�b���~7 �Q�j�^�&��  ��e�> ���,<˞ Ag��h� 
1N��J� �^��7 �؈@�w�s� џ�g
��vf���zFW�Ӄ	�k��V1�������A��l������\2� ���%�� �a�-�E����E(�äO� ��zs� \X�h	�DS vIz8� �C���lt~j ������� ���['�� M��	]� ���)�� ����'G?���Y� �k��q ��W�'�!�~i �>�h��0돢`+��� K����\�|� �}��仐,�� �]P��d��$����3a�R�.�F��| v����� ���y�K���qQ_��\h� �)��̽�'�xո�{9� n-(���� ��W@ш ]�[3�� ���zy ����G�D�VO�� B@��� AX�4J����S}i��#�"��w ��Ps�� ���[�@.�q�(� �Y�!
�� �ŋ�� �x�1�� �[��^��.�E��z���Q���G��7������ Nͯ�KSI=	� 4���׀� ���,�{ �v%��PX]gL4c[�I��~ v��Vd�� ���g��vh E'#��)� ^,���?� ���Ks��� b�wF�-	����"��;� ӧ����}K��b�_�	���u q9�� ���SY:؇� ��q��� ��dh5²H��	�@��j�0�/p����O ��^C�J�R [��Y��P$����叜� X&,���4�� �(�h�.v$��!{X��p�'C�@ ��P��v���	B��t@����q��V1}& 	J�7L2��x0~� (�E��,� O�k���S�����0���VR�>0v�  �^�/P�A��.�0@5f�� y떃���x#	zϞ�� ac��X��;�<3�է 0N�v�(&�ԑȫ �Z�`� ���t�Br�3y�f% �'����� Ph�I�4 /3T�)��p�@�@&^�bD�qV P�s�*�E T��gj-V ^kPc��d�� '�����R�T�X���J��Q�]�, �h�c���%y� �-��ˤ�� ݀�1�]!% �_t7XEҔ lU|? �	Z�� !�Q(�`V�S��" ���kOT� ��+	��4 �i
�,�O �[0��;t�m����|�O�x���3�1=���b���� uē��rx� 1��O��=<\<B��l���;k0�!غ�� a�{�� �~0hgX "�١z* ����Li�)�0�A��5��z� �NV���1 �vXQ+��׮S(��h�@: .� �K����*`�c' _� p�&U �Q�]�B� D+��N��� �b8��F� J�q�P&�K�}��,h�%�	 0�\��� �-��C 	�K���H ����Y� ��q��T	Q h&���.�` )�[�?俁%ȗB�@���H��QА]�����W�+��/� ���.ap ��ʕ� =/)џ�&� �O�� �� �U^P�\>J?� Α����D�x ke�@! �]hQ^a��o뤟┌���?^V- #Ϻ�s3� ��Hj� )��N�_.�>�^���[u��,��� ���� U���I��tw�%B�|�K�:& z ��o! -�1�WG# ��s��L�˓ �ڝh� Kع�Gu �~�ǝX- �,
*$�� x���� U�����P8db�R�a@m��*����J�\ݠ1!�Z� f) �R�P��� On�3@�� � ��%�7�_ެ� sd��P+ �wq��b� �h�)�Z #���fv�/ ��:2��9�!�����
���t$���P6I,8�d��9)�U�]��}엻
���~ qA0�) �J_k���n���A����	h� 	�{�m���-�^�`Q /�Cr�j D,�z�ށ'�#�7���� �%�j�� �4���=S��TX���{ ?6p�y|�� J����� �A�5��3U ���x�iZW��h``� _����>� �����Y���l�ڽ�	;]�(m֑4�_ ��,�#Z�`Kϙᐄ2(<�y���������! r��(�\w` ܫI<����5�*� G,'	�:�г�̒�S�% ɸ�i������T��f��Z*�5�{w� ��U�$�� ���MP(� ,S�	�`X�oݧ')�\� Rw��P��x��Z,�01�)� `�Ԑ�'S�� -�,���5���8@���f�E]�� ��uloq#���O��� ��e���R�D��$h�ˀ�꤯	��3 �ZQ `���^�uZ���. &<����#͹1�� ƈ�V�� d;����	!�{���uA~� [�*��|? S,�d�Q���uLr�1Y�O�>�X��Ġ�,��� ��W4��wL�y�B E�	���^ �C}� ���
J� eS����d?����@�#��0,ي
qn��L���UN� [)�h� /s�r�J �05?�!� �"�_��)]$$�X �j���� s&-lZ3� �B+W�ֈ ���i�KuC�������G�	 �-��I�>k� Cd�1
P� ��$	q�O;󱀀�WZ�� _'(�z���\RQ骮0�& 
�5gy���� ���.ؿ\k�|b�04� Q��h( ��pRU~3 Z� ���|�:�]��U�T< �=�'�Kw10��������  �.W! ͿM�@����� �����t�u�=�����Ź��5 �Ȝ�PWE� ld0���|���߇�II�+%����� ���k������]�㋀���� 8%�q�M���
�N��p:��|�!�>�L�C1���a {C]�=���4)� *�^2��� ;,?��y�P
�静�����u-nv0���V�2 (�0X(H� �A�ו�� S�/0W�[
��j����x dB���_� ��Z�J�3 �B��u���a�n����Z�/�_�@��㿀�-� �I�\� ω�fO u�`%�l�t��_�� F�M ?ư���$�(�1ծ���}P�"�Wn�� PS�.%K�=7� ��ZNX �a�*�> �ɷ�W�� [��}1��e�� �f�V޵#]v��x�k^�" �W��'�8��J�*�& �4�.2�o�`=���S0$�T���H��� ���We����v��Y�
�@���}��[>��-����� �;e�#�c�����@���!� ��� ,YzM �D�	[@(� ����÷``����|-0�!�*�JM�SO	·��h�T �/r��D ��� �vA!:�V���+��p���@Y�NM.Tԟ[�Cf����=/ Ó�T��i) �	���� �'�B8�hw*�
C�m�(� �'^��d� ��sP�-,Q��㥀����<w� �p��2Ϗ  Y���� l�D<3@T' ��հ��� �B�SV fؓ]K�� �`|Rk B�-���� �C�'�;} J*��H���  ��]9�X a[��ZH�`�O�N*�� �f�8{�L����5*��� �� ҈ L��ֽ��H�- ��@�_A �2��{t�oC �$�	w� ���Z��N:( ������ 8E�K��� ����h1J ��- �� �X�R	�L dv�+^V�<�8��:��.� Q���� �a' ��,v���#�lI� 蚉N��U0̽�	
�] �*���� u�B-�����c��ǧ�28V�Kp l�=%�<�; ��ۂwkt N�U��o��A# �@X�%�`q '�yW��� w��M`�X UQ�{�� �� �;���=�g`)����h3��ʑ0?�#X _p�AUB�}tGY��; )�����W� �}�|{�@q0(�pI �$�.��#1�X�[n�eM� �T g�σ�� ׺��BM ��Խ/�� _{h�!, � ��	��E\\� �1�n��-X=Ch�J��� rQ��Z�� ��4�5�N�
 �]��!�_���2P`D�����]� ;�%�Ɓ����@l�� �q�^{ ���*�_ �%��|;�r c$���ZX �g�+��S>f��" ����[&�-�i`�2�"�D�L� @��] �#�"`0�����2�@1]5ȩ/a��$.�y�nF/�z4�R�� Qf�aG �A,(��� ��P�JѼ���ற/�:	�x -�:Cl �OTB��1Pӌ� P�i���h �ߠ�"���	Yeo{ D(cH_��Sk�i�'8tr Nf�R(� *�d�CX=_IB�t-���[�ύ���� & IA��|P� Z��+2� �Qz���S� | '��w� Df\���? ��J�1)������g�#N�j�7���^ v«�)r�y�V��ٸ<�"����ȑv�(?7 9&��� Y�\�KX ���0�*��/�| �&�	��o]�5���Mh�4�
"� ��z� ?����{��\
����� ���.S� ��$����>�؂���������ST�w i�
��.�lh��/�o�� v��u� ���[Z�bD ��֮^�1q ��U̻'+ ��� �HZf����\��!� hCow#���_�� ���� aZ�R/����rAD����U3 ߶�I���ꭿJ�l���� �7Dݤ��֙	�H_i�� �E:,�~.���؈��� @%��)� ���[�N �1g
�*��v�,�|�Կ� ��^J�hL8�Y���+�`3��0�Ӱ���ٓIt�pM D�1���N����*ʢH�K��i�Ē)9���PQ��%�@��C��Y��	��?�� �R� 0��7�D�p ����`+ ��Ɵ|'�eD0邪���.��� H(��� /)�P�m� K�qN��i S����������CH��jX �3%Q��� Z� ]��� tV�0�BG X�{��� N�bu[V� ��`��F\�� ���S=�~b���c�
X;����r��@�1�-�7V�'��؜iC ���Do���`[���" q��٬ YP�� ���&���-%�V��2�Q� �b���cw��� W(�&��` �1����;�P wϊ���� E�����& %qW�b��v� |��`�� �$�S��:�@� �Z�& ��(,��C |�^;a�SM�*���$>8B������6 ���vŎ� ���1�� ���`�aK{�� 
ߋL[��!G�q�T��8�����	~�+W5�ϓ�'Y�g�)��( �4t	Tʌ�� h�H�ab��w Ci���=�	 :��qJ2�wc����o�iu>h[>� V��R �-��C1N�< �^�cؾ�ϐ �3�� ��2~�VN�����&�����׀�"�2� ���]#ɁX� ��n� � ~�	�P�w"HKa 鯩H��1^�@%����.�hpp��5S�rn�s�� `gf2�v��E�1���@�^��q �.�_���{��4�CF �@�d�,�vDʮ������
�_��4`�m��� ���z�ͬn T��,���s )���7'�>�� �S�g�qI PK��3k.������ A��� �CS"1��0L*� ��P��	R � U2��< ���O���b����L��&6 �� K���'�5 ������9�]y �6!��G�z �"�Z���@t)Pˀ��M� Xz�hT.� '%���9� -+���k�Tv �\S#һ�d�(^�"0<:����hm6 
�o����a P3��d��`A�+�� $V�%�[� O��B'��f�N���	���h�<R� `���� ͧ֎��[ŏbS�9 �pQ4<��0 �]�k��L�6H
��+��O ?��{�&(� �P�iD) � �%��Mw�PϾ�T0�txT/��,
�a�z? :1�2� ^��(6��|������{]\�l �� E��A 8��]"�w���z��vn0���G��w��E���-�s� ,�(�<��V��K0�� T�X�\ 
ڴWߝ�?�;!r � ��[*s�$��5 _��j���A�%��#��F *�	@|�c QP-X�s�<� ����f �1'����X�F�ӡP`�0o}� �4��/�a 5��f?�� @�V�� N�1�
�� ���fl.I� �X�O�K� c���b�;�+�L�@���~Uar[�@ÁM� m����� ��(ه��? \��2QUJ ��O�rm- ��z �A[}@ ~m�c� h28(��������`}�
_x���6���0�5 P�}R��T� A�*+�p� 4�	S�y  �_�n�B��2��q�'� �����{�� Xs%���� bfCN���à�  ��r(- �3�
� ��	E��  9���$J��Ӹ�]e ������� �s,0�[ ����YRP�i�ZX@�I3W��^�ĸ�u:	�hɀ?��p �lkJZs� ��M0 � [N�1�� _~��	�� |�c�9% ����	W ���Nc�$�:� [��X�^ 闂\i�� �D˴��Z9�y�s��#�p�3
 ���R�ES8D�� �Yh<��% !�\�� �0�.���� A���Gn��� ���B2D� ;���\ J����ˀ�w� -sopn	�P�6TI�x0l����W�k+T _I���4 O���h�o��N���`�Ђ`��e��� K| ��h><��o�5(����2D�}��� *�[K,���4	��@rʥx}�YҀbU�CS�+�0�)����C�3�f��Y( �R��p�| >����� !���M��t���_�^��� |�	���
 ��E��y [H��^���{��R��Y�P )4 ���`E��e��c�j��4� �����/�p� %X��������	U�&�0`��g��@�W#߿�C%4��t�-r� G�fi	 O�)ذgQ� $��H%�EK��@TY��P1͸<����%��x�}A��Ltۀ��u��O��$
��%y���r	�W[yi �R�� � ����n>v3@�
�(��� <�S2�7U �.�;Y�ö�'�"��� 2�b1�� �{	�[׏� ��w�� ���3��.���q�!�0H�+��1���ַ�  ����r ������9�/��.(�5O ���H���k '�e����[ ��L��N� 0/��q�B;_	-������^9���9��8 [ ϶�:�믑� ҙ��� h�1�}ɍ/k�A򯥂@�Q0\�` F�S��;��L��+��@��3<� ��	
�uyc\�"MIcR̀n � *�k��2��$ \S�D?rɎ� �@���x����X� �X�5�N������)��` �t�Ͱ����R��H_v �� ��0�D�����X��$ꃆ <�a P���]K)I�  B������ ç,�A&R �1�H�/����ƪ	���� �ӫ��L_cpK��Y0�X"����e���0 �]S�^�E�XMA�Q ���� ��Ⱥ �0���p��ք��� �<�U�5�/ �|�
V���8'P��h%U5D;��} Z�!�� @hMRi*�����P/ Ѓ���bA�Z��p�����b��=@Q� A��^;$�	�g4��`�L0�^�����N`<d\ h�b���� �+T
/�oIA�0����b`]�DB�j=�h�#�֞��[1�����������LIB$�oy���� �����V	�+��a%���(Jٯ�q��,{-�����b�
  �hau� ����Q�%��t@"݋(� լ�
�:�%��gd�~� �=�#~� %�P�<ʐd��ſVA:`-���9�_}ѹ�U�;p ��ɷ��Ր� �_J<힉� ^9��� ���*~� �w�ϕ���� ȞL����� \�����U+wHLk� )�8���Y�# '�xo���l��+G�9 �d�T'V%� �8���_� �d׳��*�/[��Ψ��� �����+�o	�P����� ��Z[QF��\�� �� ���x� �"�!:�	X��ű���|  ��5Q��/��Y,� ��HFx U��=������`.N�I��62 ӱ9R-(�[��q�	��Z.p,� H�U"� �т;��7� ��S��	>Z� +�ʲ!f'��@�F�ټ�p�D �����l|'��c�?���f s���a��|��c��-�<9����C��� �fX(�L�� 1�hU�o��p��-�bY�`&s?A��^)�p�� 2�&��� _r�%
��� �!�� �k ���]1	�� �8u9e\:- �*���� �$�ȃ�� w�Q���8H'�#�`� ��w���� 	��Y}H +��12j� iQW�<� ˅P���� ���!�j�~�9�� ��|�n�p����+�3,�K/@d�Ʊ�	� -k���h [g� ��B x
}F"HT �|I���܁ #+�8O�<ٸ��xP!��V �'>�vװb^��\p�\�@�!Q ��a8��r ���*�R ��f�j�O�`;�*� ����W�����~B����@�W�����5���3 �hjk���J��� Ex�/���kN��":��8e �}i�d� ��q� ^��WP� b���S� 91z�i K� !L
�o�v �/~�d>� ��C��3���� �����J�S :,���߰ww R�dz'Ɂr �hoK�l���A���2~*��CW�r
��Q��a��Xz[ �̱T���U�PO�@��і�%~t&����� �� �h�Q�~�*�)Aa|��{=[���3���o@R�'?O���~r`2e}�R��`D� �/�J��A0$�Z�K.�p5�Ԭ�$M��e�@�G� ���j�c�� @R(�麐 �LA��9-boV`��� �����E���4�c��d b9*p�� �Dh��	�X�E0� �e� .]�1��eoT7z upP+ J&�,) #����}D(@���S#� �^���;`��q	�n �d i���M��� m�������;�e%�lf��W uF�X��  U���	�p�tXk� 1ۂ�@5� ���b�#�Hq N�!� �: ��9R�� cP�$�� ��
X��- q�� I�&byl+��-���±�A`U�Xd��D�y`[�	�� �r�	S��w{��݋3�n �쮕��np� ?�b\ _��!��U|� �+*4e�w�&�GI���� Z���<B�`�g �� 	F���1�� ��YQ��=ź��� MreT ���`�U�w ���x',W �n-X�( �u����! �Z@	<�1� ��)��? ��N���h�"f�|` Y�����)����n�� ��PU"`�\�}]�O�a�~�)�L� ��\���K��@�&���ŗ�瑒 ����*��3<P"@}i	\�� �Q_�1��;B� 0 �3���	/�WC���T� $�
��<�Y�_ �S��^�3�� ���=7� ��<��B81�<����OF�º���Q?�H���0y~�X h6/&����[����0q\7h ��ʩ"%-)�z pɿa� {���P�����}����x� �'*��.0��,�W�}a�� �;���^��3�4�ض�V h�#��� �%�U�� ��K�ٗ�� ���-6��S8��Q��'f<c �:h��� �]�@�&	� ��I�L� ��}oS�( �hst3F�۹Kv�W�Y M��� *h��$�/�� �v�@���^�D��Q�(�T��F���-!�񼉋� }�%h �^�e50��! �@���,�S9q���b�`��� ������O��. �T	�?D��z f0�笣�2 �$@�-\� �wу� ZP��O�U����X!��G >���L��H���h�; ��.�!�
� �)�:�u�@���b� w�	��H<  ��/�Ą5�S� OL��2��ӂ���`q��v�P�z�\�� S�q;��,���	��Q(�� ��0�?� ~�7-V�\ ��y?�k�p� ��r9�C	 ��v�0���������u7���K@�U@ʾ�� ���X(�^]����|����<�=嗿���%v:��� ���R�j�(��`g!�������h8	�����^��;�[��~�G�V�� R)�2� ���\g���`��vAC����B4<8&� �2���@.% '���X�u� ��\i�f 3a ����) Շ�$i8%x	�"�9;@�� �:���}! ��*��r���/�k_����9�a��I�O� ���Bi%PG �Ӥ 7 ��|"��H �S(�'u�az?��d	��/\- �#"�����V@����� �t��Q#�(�1� �_Ph�Z �4"��؜�[�(�C��ˊ��� �P��W��$��r�C�� d�^k � `g(ǲ'�$�s� �BD�^�������Jz� ����7�;� ���%k 	�W�$� ��u���x�x� ��%�8� �[�,�Pj.�S� -����  �m�� ���P��#k�u�*�g��,	 fZ�U�{[ �׷R�P�c0�D_�3�XY���[h��/]��<O�6 �; ,!�� qϟ�V2� o�aپ#- �(��1��Y[ �gh)J l��p��HMߒ 9�	�{�@�r��"u �w�P�� �})�NQ�� '�w�@�����a��p(�l�9�W 徿��B �a֠h���� �\
�	��Y ���@�Bw j�_��r �i��J SPU�F�xf �����&|� ����9�R���Ӻ��H�z���)@�������P���SaY�����	a^-�H�0`(Xb`� ���~�6_M ޳2��U� �1��� @��!y� ������] ڴJ�C �I��n���8�`X�� ����R�d n�%���) x�6X^�s� 7f1�K� ܮ���uSa*ȍ}����-�Yw.���`�Z1 ���V���q30���";J�^�P9� R3<	 � ���+�A '1�Y,�O�^�U��y%� ����4�0���f 	�'��`��� �
^��G�_*(f�qB L�1v�>#�:���|
M��2�> \Rx��Wo�v��80�	�(��?�g�j�Bc1ʸ$�k��X2 xӝW�H�.�~�	�[!���A��|0 �@��� e�"4�TR �=/K� +��Y�JP����m Ҁ4� K���
��  �0*����fĪ/s�@Y�I ��%_a�*��p�B�`���U EG�&�.� 2���x�� �$��L(`@ J1YǟX���G�A�I�ۂ�У��YR�.��։q�*0�"� ԭ��� ����~��u��|M8�-� x5�aN��h U]��K��JDp?sÐ���a�`�F ��(�Cά� g*vō uT�K ǭ�j�Y �W$(�Z�]�X�x=�� ���DTK -��0X��L�) �hθ{@ �R1ݺ�b- ����D~4���� �^ ��B���Q2��$�#�V ����
�� �A{�f$h �@�֊� � *A�y|��x� �N!�� I�P)�Xe ��@��W� �Y�-܄�^} V'ǋ;,jYX �u~?$� 	��_�<����h&F�츐�!PE%���01���W�`�P���NY�$�`+� ����b� w<�3��?����*I-�%�g ���O�P ��6�����S )��]� ���k�,
 	�Y�b��|��3��{P @��h�q ��۽�Jʉ ��(�$_e 	7)Y���9H�(�Z�1��Uz 4�Ӫ�fT]��p����s  ���,���|�(��?����4��� d�«]X��>� �À�!� ���߶%�s����t � ��JS�9	3�X e�y�9��`!��, i��7v�<�� �y����l ��h���I ��2��k 1��+H�>�H ͣ�ć	� ��|�!`��Oʨ )� �� t&:@��� W�Y�/� 7	� m#2! �GhFk� ��M�N�� `��bP��T�#_X��M��� \(�S�% ø�
+{ �Ϸ�tf	[�6�@i�ⱉjʙP��.(�� 
1����� ��h� @:0J����}� &<۩z%�uE{a-���(����b�]�����{W �@-0��?|� Sb�̨�B �Ȁиf��[X��K�Am ���8�N-<�z��@'�<���� �H�T-���7��bGS
� ��[) �*>�^�i0 ����6g�, P���ڱe\�"����|@�W� ��9-2��V�] �� j	v�Y:�p�$/��8 H��Tf�tOg���0.��w Z���Ѫ�}\ Vb�>�r P1
���%  0УSI�	 ɻ�_�?[� �^)1�K��0H�"!\@�i�(	u� ��꽪���C08��� E�� 1�� .�ē��� -sxoLY U^vH�u]�(N��>�� B�;@�p �J2)һ�7���,�?�����kM����D ��p9(�z �y6i��� E@*�;hk �e���l �4@I	`��<�� �-�#3��;g��� С�L+���^��<B��� ���6 ߰�d���h�p�n� o��xI�� ���SR-)� �4�/��I�� ��E�[����#�}K 0�����_� ���h��� �T�����,�1�*�R�'�H w��饏 ^��p]!� )���~Gj 
�Ŗ���sU ɒ��H: � 怓V�r `R{���n��(� �#g�B ����^��2 ��(&��� >֮aR�� Q�.�x�~��p ���;�����7��#�_ �U��:�����3 ؀XR 2͟�~KɊ�� �k]Qn�+� �`G�^P� X� �-
� !0��v@��L�hIV.�c� *�)�YO|$ 1���^��l ���-+	��=LN���Ӻ⇎��+�׫ؐ�	�sDY* ����:�W��9\*Ė> ��!AZ��ٽ���[2�� �J���8 ��u%3��~�P �������y j,뿻���E1���A�J .��z ��<��ny�
7�@"p��V {����I�	ȼ� "�Yhi��A�U@���  R�[��Z����<� w���l�( ��[��v� ,�M^�GN�w;�j�X2�ٵ^`��	�͋���y�l���h�t~�� ���'RP������|&HÔ �x�bO}rF3޻�"���[�E�]�^�pԽQ ���1�X)�U���h�[$ =�`+n�Q� �<��^�, ����� ��'���-X[�O��Im��j ����� ^���[�գ��Va
�;�`'��b;hݽ*���V����}8~_�`�B�`���Ɉ`p\��(h�ӵ~�Z����҃�������@hU����[��� Q!L�0+� `2��O�� ����{�� fh%rKb�U|� ����3 ׋(X���"�9���W�� �x3]*� "z�+�c%���
PV �)r2�X��w쓝T��-� < �Ѕ �, 2i��F�;R �K�$T0�} L]'	�_� Q��+���2 P���X`���T	�8��7 9H��X�sK�|����pr	\ h�V&��$:o��4]��3 ��{8�  �-��|b�X�]��X���� %g���7W�� 8��d� �Y!����kp��<�3* �Z�ȯ�:�hS��$�@���[��m�n��!�/ �T~B��5 ��Q�w�y� ^FH@�	(��!k+�Zo/�x<\"w�%s2�������r ��}�iP��p� )��]J���3��� ��^�&�>p��p���<+Y��������_D ���{� ��)J��ҫu��¢�?��j�A1�]�x� ��*��( 3[% WjZP �S
@�_� ���k�� h)�G>�,	¿ `�ƺ �Y0���qu[ ֗:��n� ���?HB� �
�r��� ���~g� �XJ\�%� �޳R�,��Z�Q}� =
 z1-�\^U ��滰<�3�P�`xEk�	������J��� f��Y� K���� ���l� ����G�!� �����F(�SY���3 )��y�@^�� �R��j���P@�%��2 ��H0�,��_1b��| X�+w��a �
��`��bA S���� ��@��0	�s���
Q�� h����A�1�w������r���(� �^�`� �h *�v�L�� m���śM� >�}0�^��t.�� �j�@��\�FX�Kŏ �%����V1 �:!q �= �YI�[U��Q|p� �_�{J �B��W� ��oF<��=�i��@+@�Q��<�K�ÀaY�	} ���5j`�� �S2�O��f )�]�[J� (
�͹�	 w}�f�����%�K��Ǎ �~��,]�h�@����wc �iJ�+���n���) �0>��:�/}�>�d0�V�6b~�,� _?x\N�L���Y@��J}� k�����h Ks�b�c� �	�z� �m�1� �H���� �@	���Wy����!�7J� �������;�Z�� �p*3� �J[�D5޲�!�/��_�ZG \(b��4h�r% ���J� XP'�/� �E���J ��f��Ɖ#� �
���CP�KO��� WĻ���T ���[ 5�z�V����n��q jl^�Q%�o���S �� x�0�LY )ݟ��� Z����>�x �0y��Y� �P=����(oh� -*���1�$���P�5� b�u�VUe `��D�L]����ؠ���ɀ���ݞ����)	`b��ܔ0 ̋
�[ �VJG�� >�Y�	���Ơ�y�j,+/���`�� 6�L��� ���q�]~���&2b��p!� �o�.n�Mr�����z��+ (�h/��, 4}��%L:��I�̈�U ��O��@�:��]��r �'���k�z��^? ;� J	e;�� ��6�?< K_7���� D�(�V�N n<h+�7�%�c����x3&Z� ��`g�R��P����4I��1��녿��)ɘھ ƻ4iF�P 2��Q��a<� �Jɬ� ]>�� Q��s�` �m���Xh�S|�`�fB I�ɇ��* �t!��bҠ��] N�����
�
/��i:�� N�`�)} Y;���_��e Y�|�)$ �Pb⸛�1UG���*� ��A�zٔ/���0���Z x$]_;.w� 'QU���1�H�	�B>x ���0���e�&J0�,"&b�� yߖB��=����X�����P �1H�~� @o��%��_��^�Y0l�nJmA��h"r� ��-�t��yQ������{�Y��_�X3�J� -��	�z& �W�пY���{��T'îfhJ���;� � ��!	�|q���v%���*�����+���Z�l�x:�o@Byݎ�� �����qN��` $�4AtWR	?
�5���$@�h� %��պ˞[ ��0��RZ ����oK� "B@�,�L�� �H3�� �̹ϐ�� ����o��7�A��@�� ���黨X u����� JV��Rw{v B���ޤ �oD�t�C�ҰQ&���� 1ڸHɨ[b?�%�_/���tX "o#���  T�_����
串�� ��-� hi~���� �/e���� kH����z�� [
�Y�t��,	��@A!�Л����� x��.�� a�W�qo?Z��� �:ьR|p ��U�MX��"�?��j���*@er� �R�5��� ����*�>��`x�^J� �h1�CH� $��[ ����� ����%H !,���e ��UPy ��a��?��<Z�(Xÿ��Q* ׹��	��9�[�����a�� D' �@(1� �f%Eo���7@���� Q ��^΂{��-���Ä4��� 91k*�8�^\� ���$� ������1�0�� ��f~5-�d)�g�i |�O�5�k�sb�7Y0MK{����{�j���'!��N1@�:i%�Q�/R���U�?�S1��r�zN	�����P�+��Jo8 ^E���9���R�'�����[���U��v{�T����`J� F����ɡ=��& ��F� ~���g� �hk����� |�ۣ^�!ظ�t�N)����`n� �S���ܲ9�1 Y@䝽�P5�>�D@�厒z�0�%`�l���h�৺��	�f�ܑr� ,~���8�j .�+O�FR�2��:_Tp��p��X�)!��b �1��Y�;��Sr������ A�Z�H�� �t�l�������p? �Wy�K���#��eN����H9���j�Ń��� ����A  #��*�� .�!9�e�Q�z �0O
Vf�P�������������R�� w � P`�Z%0�� f����_1q� y�N��P� 5=� ��� H�QJ�̞ �iV�t�� �r�
�B��� �\: �1�Y5�xz�}:S�����^ ;Z'�A�, 0���=b�t�-ܰ@�h�n:u e����$'��T�@k)�� 4�
2�ha b�Ȯ��` w�k���  [΋�x� ���i��ݹ &(:�F ���8�b _~볘�2 �˵uW @�tj#9�S�2	� ��#��� ���(�;%AP��[���҈���L �<h8�5[�g�Kw�G'� U��7}�� �푢�� cH��]�'�;��0�)�fwƣ������ ���}�#��`��O ����;�[*�� W�/���U >���9
�� �{�m���� �2�K`U�
 ����}E��gN���)�\\��W@
Ϲ�Q �0^­�h 9܆-Wm%>� s{���TXh�M�����n�X��� 7��¸Z
�:�%�ܰE�sN}vL'� ��C��� �g�A`o�X ��>�3U� �0� �H��N]��P"��O3�A�Bϐ��� �`�3ζb��]Pə�������$��q 0���/Ė�.�5"�;���p��,E��D�����	 K��o����St���X 1���ò|T ��P�u��� �	�s�/xs���P���f�~�%|�B�[�� !�{�-��w� @،�?H89�XݾԝS u�]kN�`{��Ķwz�	�J
Q �`�C��.'>�1� ��'��א�V�PT�Z��S�o� G6-z	 �hc=�j�s�a ��o��� ��<@ɷ% u��B0 \���
�6 ���1h+� p�V���wXXj#;��#	WC��L��V� ��Ql�/������̟Xr� ��^(��>*׀�� �Hb`&Z Jw�)� ���M�P�;K!B�< R ��F� ���	 �U��)� ZJdش(ş�AT@Ҁ�EL W��_���Z�~ ��W<�e��Q�#��0H
��i�����>H������)�g����y'QZx��� %�󜮰�Y �B�h��^>`�X�X� e'�J�)� ����px��Q�c��B& ��$���� �)P���&�� ��� ف% �Ovդ�� �Q�cY[���������B� �x^k�}L `h<v/�is���D �S�0�����	��q]���9X��O�8 �Z@A�� I-���t�x mX\}z� !����w ��0ɺ2*d E�����FJ�̀��K>OE�e���*�� ���80��9%�yqv�����2{	��Y[��3���Z.� ���S�2�N�_ ��^� ��%:�&� �ɠ���`��e̒��J� �]p|��y ���� XA�$��/ t���( ׵Vh`�����)����yZ���~�Xk;p�L8� U1��֕V�|�Z��2��yS �8�3]"N�DXt~�`$T��: ���N��_� ���Q�� �K'�`�� �d����j� ����I�� ,(�4\y�� ��Yc ᤠB(�h}%��@�'0Q6C!nu\��� ��7�W�H	\�� (�TmI� �%�����e�[���0(^�@�Tn� v�_)���� �\�`	�sc ��߄��u��d �t]+3��"@ O���Y���tz�؝� ���A!�� ���6� w 2���@ �I`�.Q�:�y ��S�7>3o� r� �P(2����L ��/� ֻu �y���M�� 0������?�[ �rp��� Rҿ���O L�|����:n5[����}�W	)�F��b�']� ����[Ӝ� V�S/�ߞu$%HX ��n  |�^j,�u ��鼾�$ 5~ ��%��9>	��a����� <E�,%��K��B�h#H\ k�� �z)���"��@�� � ����� �^�S�� $]��/�n ���>�? �u�k�|% ͻ�ڥvb?�K<���� @�� �c-���B�u�^����̀zYH�[,hP� )M�1� sW����`�b��5�;�������eP ʳ�X�& ����jf� �� YI��."� a�#�n�d���j�a~'�S�; e�� �g Y���G�0 /�q��'z���	rxD`j�\�S�M�����X� �
�P�(��;ۋ�	�d�|� !��(�R���%�Y�
� ������P����B ꨛ&��s)	WG�@��� S�|r��# ���:�9���;��{�*��{���C����?(��� ��'�ӗ�?dRO�+���# �����&~=�L� ��4��f ꊜ�UT]\ vx��i��X����]�� s�,��	)� ��+�J5\�`��H �0(�� )�:�쾴y��%"0X��`�\�⒱p�  �!�-�I JB�<�� UC˷X:�q^ ��"I�4.���1���zg �I��v�_$�ōQ��ɣ09��#��h�ޔ���qp _���[�!9,b: >���/��@�ZvJ���b�� � �9-H ��
���K(�WY�_� ��cg�X[�I\:P���t�s� 3L�K�I�H��1�����@�+�R �������O����!
�C����� �^���e V�9ϓ@� Ž��ݼ
	ZXY��*}�� �]V���n� �	�FC��� ��Qv0�U  �JX��٘g Q���u2�� �%/G�F XV�(Û����۰�.� 9������[� �\*w�� �7���U�%Jz���F��0G� �P���̀�vg �)ÝB8a �[�>0܀ <N��Z��$ gB!�]�P��/�F. ��}�����Sw� ���{�� 	w���M�(�@� Ar)�$zX �l?�yb��@���	[� Ȩ���2H$�h@��P� �8�Nr� ��M��ۯ~\�����p�b� �AQ�1���Z��b!�ɳE ���SB����{�'�\Z�a����0c��� � �K�׮%s և���Q �VY~��L�c M8z����j������]� �T�s�$��^ I��Y( b��M~�� ��h�#$�Q'\�� �ȊZ� ��� W�� O���
3�\�*�%;���0��ۇ,d/�p����� �:m���$;"PQ�����8ߖU.%@�� ����`L2_�x� �3^p�㷠� )¸`��<1�&Tc ���J�� ӻ��/�@ �����K�� �2��O&�eI� $��� ��	���'�����@KpO�u �F���")��3�@1�\Z� f�}���eɬ������ R��0O��=��^���%�o=�b�� ��e��v^�ϸ_c���D ����'��[=�q�}���^  ~�dH>���-�3�8RAQ�ñ �4:��\� ��'%��w�R���>�0� E&��� �lV��'�2�? &�s�p� �[�V0�'��v_h��G�.��6c��3��XW�,m���ļU [�ݦ��J ��h�y �M:P(z� �?OY�\2w�;-1��9{V �j���*�����<ӠQ"�4X� Z�d��u �_���l� �L�"E\ ía��+ B���<��2�(�� ����� �Z���W� �'�
����R���А�5!г*��R�1��وr���]; J�&=7 �ϒ/܇�� ���|�k �A$=I4]\�}P#�u_������ �`j()ƀ� JB����.�<�*Y jS�ھ �[�zBһ\�  �b+0�x �N�)z��� ,��2�C�F'y0�+���΀��G� hs�jk�3lZN�\`� ]	��B�� {��;З[S�� Q�i��O�T�%!��4�=wy�@�PǠ�
���L��� @,��b���q� |�ag�)� ���_� ��+��Y%��)ڰ��@ ;X2��� ؛�8�I < oԟ���1�|b A�;�
� ���&��=a��K�%�����ʀ�!R��� ���v�J����c� ��B��M&��[o�:�W�'�l QJ3�P��|� ȳk��0��:i����W \��;*K�� ,���Ӕ�L�)=U�-���������Q�G����*	�>�L 8wܲ� 
A�_��P0�QF���w�>CN �)�n�1 ��ׂkb� u�4�h�T�8 ��$�& 3�^ei� �R���� P݂�%}n �Wٺ�� �*��	 � �B!�(�_: a;��uC?�y` �~���]�r�x_��G� ,FS
	� u =]h3͝p| ��2��^m_�Ȁ+��A�\He?2q�_��ou ����O�zr! ���Xꇍ �ź6(�Q� !N>KJ��¨����A�Nrr��Xn�+����Qx[ �x�Y�1�� ��p��-/h������p�F �y(� ��a��� `<V��$�*�;\.f� ��C�u�nA�"i����O�À��Kv<���������  >f[���Z ���ͬ�	��b| �dˑB�'u0�{9��>��оr�y���t\�@��!8� D�Q�R�%��:��r�`?\ (��[$��y	� ً�Ņ���Oa�6m\�^3,q5�B� �bl�FR�� -�)��f �r���Q�o �^�pk��� �/�N�w�[�1]Wa����;�����S� y��1G@ "�
��!-�hС�!�W�Ś�� "��*Y5���� ĞZuX7��} j�ahB6�% "��'�q�	��/) ���~�w� ݉Dl]����Q܃D�[���� V�I?�*
 &������� �w�dv�� ����� ���[���~�`.�#� � -��m;�u� ��P���� i0�
\�a �h��_��< �'�>�	8�iJ���� ��� ��M����X�m<�� Ѻ��l<U E���^K/� �:��V�	 �|I�h�K��@�Y��� U�L� �� f(Ϙ�t�Km�8 [_���. ͌�N�1�&� �9.� Ph��Qï?G�� @ڽ	���tu� �2�,�lL�p"\C�P��	������l`a C�H��� N�̌��x� $Pc�i��~ y4p�KBW ��?ǻ��) ��$ϮA�dzi`�D�� ���b�E@ ���&��;�� ��\	�#� �UV ���DʌKH����� I
��3��n����R��z uި�( �Z��P���=��,1 � A�|�O�@,����?
�CI�� Yw�<���� W)6!u-� �S��� X�T��Y2 ��$S�4%, ���
����1 �_�T$�MրTx[� ��L^	�:� �Q�`e��BQ3�ܯ�IJ���5u�^ �̪��� �=C�
�� ���!�?��%�/� �8;��� 4r_�	�YXN�rq�2��t{��<�f�r�׸pmzR� ��hEJ?�%�:� '��P�R� �T���}n �Qh5�H �@��Ӥ� �T�B�Xu~ �Zƪ���+;	�2���������Ή~ �,|0;��_�	%���/ ��:�|; �#Ǻ��� d_��bL*L�� ��|X��M ��:�Ļ�p�`���y�8 �@�o`6)� ,	�Ά-�"��@?Uʃ�n 7�P��f	 ��e1�B� ���@P�q��# U����'�!�Y�mf� +�Z�'td��3���L>( m1|�2�N�q�f��L� J���_+9w�QFs �V �/{S���)�T�1տ����y�D�a�0���� ���� t.1*�+�	�#�y ~Q0��@ �΢(�-�~?�5ǃ���>������ƀZ1ͻ;U����؃�9[����w�B� -.����w��
�!�+w� p0��4�� Y��KʪN� 	�
��B b���<�/�� ��R0X� H-��  �)�>���,�%��:(�O� `�����/ x�F	�N�� �u�#|G� �����0Z9h��x%~���X�v:��|\· �8�y�C��B_{D�oX�:��� ����� y�B�حh%3�#��E[L ��"͋� �s����0 �a�kS�9���T���D\׹ }�ӎ�ψ gYh��A!y~?|�� �C���^��x u-�3�� �1$
0O0��� ��:[���� !�f����oKU�� �h7ZB��|-����(�
/�3���0��mhI;<`�OC�B�X��ɯ ���@�l7������� ���R�W,��  iʷqY �px���$ <PJ��b� 1�W���[�
������d���	 /�+7�N�qh�: k�^���uU �.*+�|]�gG�>��� V��ٸ� �x��� ~�Ȉ��2������չ��6��2�n��� ��m��TP 1��L*�\�O�~�� +=Hݽ�N� ���K���I?Y_`��m����� ��M2}�,�_l K=k@�1 �XN��ޣ�!����^# D ��qЕ1��L٧ K\��a��	E��཮�	uc���Z� S��qեd iXCk��2ӈ Ζ@�� �{i�tUs� ,����2� �We"r�@�!㋸��U����	rg�R ��B�t�H�K�\u� �%3
��t.��F �P �� i
S�� 3I��0ͳ ���`\J��WU!Ȭu�G��K O�(X{�\ Ra��j���M��O��[5G��� �"N�b��mp^I�/~f"1���;��� �J�	$#~ovu �eR�]��A �f:�-sj�,d= X��@<T� ��5QE	���,`��h�L��R :�]�$6 ����BX��M�� d���O�@���N3� �� ��[!�Xwr �l�U����Ek �*���h�� 5b̩�%�� V��f��� ( ���'��pg���#	�O�y� ~j��oQ�� }���"� ����P�� _1u�iRW� �"�ٲ�� ��Z��b���)�(����Ԩ���"�,��4%�X��
Z����L$tH��67��Bf_�] ��@ � ��-��\��������	^ �sq̻_�{���;�����sX�g�� �Q �%Tq J��&D� �~�A1®0��P+��![���(����U}� �I0��B ���?��Q�	 �h�K|b� mT!�:�^��*���hf P�N���� (X�@0��?��| ��P�^� 2�Wb/�= �������� 1� ԟ� �D�+�<�A#;��`Xd �J�[� |�:^�,���x���z��� ���XZ��X[ �L	�ީB��A5�{���! ����"h� x݇d�EB ��}�i� Ã@�X�Z ��1�uOg�>��S=,� �2̸�i�� 8�r[���k �& �)]�U N/�ui�;���y.������� +�ل���� '靥��+�����CM� ;���a/�� �@�h��� �����<>ո��ַv�pq�h8��L�\�>;@�f�Y�a��̻i�-�� ]��\�t �1�:3)� �0����P��	�S(�pY��� $���" M$��� l��v�J�:C򀽣1�� �a�����_��@�T]� H��3K&� 2�n��W
Y��)��w�B\��V�� �-�0<ue �ӿ�G��.����z�&[�Z;�h'4�V�I7,��$��� ���ɺD5� *��R�bT���_������ ���S8�Z4��Į0ϬU�:N������ �%��- ���|�	��`�Q���ͧ[����������"[����Y) �]��H ��'Uw�� �Q\n�p0W��F��������Z�% 9R P�X��L�H hO��w��I � {��� ��ϭ>|�7 �Ɩ����b �p*!�� ���`��'�� ��u~�� e��S��h 9�H�cb�� 2�ٰ��:)��$0��@�.�_���i@b� �N�%(��u� xX�E\������$������E�E	VP��y=��}^�2pZJ��k�� ȸ���$� �%�V�	�5@��0 ��[��>���Ͳ���i��� ź�dKP&���kت�`�8XLS	}��l/�P�i� \J�xv ]���F��~�_�Y�����>����
��ۥ �!�4������2Ӄ>_�߀���f��L��� ��ɳj �P�X��
f}�+� o���1*\ư ���ҿ%)�[@Is� �� �]�1�h� '�}~�k��� � �,-h�'Iz���/D$��� ��� !�W��m�cp��X��sB=� �g`�^f� �>5h@� ½�}	U�f �XV��H� K����2� �\`�
�H�u�� ���V�����Qg�!G��p;� U��@��_�����ʪ0;����ϖ[��P�� ݸ�+�� {k��!*��O��ډ�
H�(��X���4�,������eA ��n�U������}�1�) �]ݥa�u z斞 ��0焈��S�	�x �^�� �ɒ�� �L�Y��R ���&)x	� bz��"� ��e^�{� �DX�_�N�����5�Y9[p��H���`�bU��Vw��H�(�/%���Z]~cY�  >	p͝qXL� ̇Q� Җ%F�� �Y�L��� ��ɨ�� 	�h�Xd��%�C���"���l ��>�Qp�J{���(D=�����I�y�-
 �!��%^�T���z�H���+_S@� � I��d���' E�6�nZ!i���h� {L����M� �e\���.HL�]^O߫O�Cjb؈,&�06���D�����ĵZ��j��ӫ �y��[��{I�VF�0 ��@��rc� ����9�)-%���qP� ;��=�_� p؏V[) �so ���	T�E���)DՎ��X�l 9�X��Z�	�@-�#T%!�_n ja�p [��/�������;�Q�O�%�ſ�57 �;*���\ �^��Ͱ�6�H�-ɸ���I���M?P�T)��D�-"%n�p"�r� *i�e�h� ��8(�KS�zk�B%`�b TQ(ة�� ��d�� &^���R� ��V�3�� �<�⻣m�Ṳ �2�S*� X[%�_A&F�k ��� ���(�bə@1!	���T�N�ʶ�Ȩx�Y<���[��B��� t'ⱙV�q7����U�;���Tăf���Lb, �l!a�ɑI|�n���pR�9 �$�Z��0�	< ��l��\ h����Ow���\�%���� Qh��1  ��Fi�oS !�\Η ��խچ�x������$ r6*�봁� �{��ѥ�?6,"�
pJ��X�_�n� ��W$ �� �馭� X�(⮆�����P���[$R+* ���v�\�yL� �k�bw�� ��
���0&��- ������ �����K� gV}
y%��?�I���w����\C ��d�%	�1ғt��.\�F�T�����L��2p� �� YZv���� ��������h���j�!��~��$�m� �]�.�DN& ݕ"�/�{�^�pe�XҸ� `~����_ )��0g�� yX����5� �@���h�� AbX �8	���]us�_�% ��n�MpH ��uJ����d� ���fm8�,��� ����{^� ���e%�( 5����>����ԇ']! �1����� ���#=�I����c�=�3�����T �ѦÕи��6B�4�X9�.�ਤ�� O6��+�/(��C��'�����LP0P�Y%,#�e ��.B��X��hP,N�@ �#�:t�  �3K���c �P���G �!ҹ ��K�n��� [�Bb��Q$RL& �:*�� /�c4;� IP�ֻY� �
��z� �H��� ���;[��� h�+)O�F������`G�ps �����n��	��
���3�p ׳įH�~ ��XR�Ӝ� �	��CZW���п��e<т��_bu���(� )Ó��2:�}ʯ�_�H� ��?I��p ̺^5�E ���)�:b3 pB��4_� X�Z�[�?HdjPv�Y�z�,��װ ���)*�Y ǋ���w-g��t[��0I�������!�h�[A'�� ̇=�KO<��J]�A�����.dsK=`�C�Sx���u�}@�-�)!�p�����Q	A�� ��c[�" Y����������M�p[ �Z1����� $^ ���Oc�7�!�]wRX�� NV�M%���� @�`�
 1Չ�.3���e U����N��� [���u���h�O0�6�#ΠH4K ��9�+��} O�
]㥉h {|�g� �� �Ӱ8�� ֝p�9�*� ���8TB7 ��vLZN _�-� C�O3�ؠ�1� io�a�x�9}_��J�k�h� pQ� O�r�� �x�7�S� ��F���P 	��b��M �1�����̛�Fw�t}�	[������Q%
����0�h��iX0�;��"~0@��8 ��L����� T�#-	�|Ip ����ϐ <�&� �h��LSj  �9��B 
C�JW�����Ϡ���n	�Q��I�FL!O���u� ,�U�� �XV�0��J �K ����� q
\���3�2`�� 	���]%ib8!;L-w �[�A�,Y(E Ļc<R���a��g�po_����n�萂� *8-��[(�k�R0�鮟��?�E$8� �R�7�0������N�&���]�e ^��݀�4\��=� 1��j6�b�T������� �[�J� ��#ѝD����]�D�! ���MQ���z��,�'��]�� ������ sE{ҳv��dr_ `��"�� *���J���`������=DL>�1�@��-�g�=L R��q�Av���Ю �Z�Ui�S}(��w�a3�0 �1�
�S \���/x|_ H�J��e1$Y��  ��V2� M$՜�4ػ �1�!�a ���
��)� ЇH�	��1�]��%�` ��b.��U�����N�����`�
 @��U5�M� �P1��=��[��V-X^|���ɸ�^�E�f����Г'��Ѽ y���koX >�5jb Bfڵ$3�" ����F� ���Z�k�19�ܙ 4�͗a�Y {0(�ô�
~)�$���BM:��/�'�,>ȉz���  ל���;w�?� ͻ�xd�|"�T��Y/��ŋ 	'��v֣� �M�8���:� YJ5�@��p� ����� ��m��$ζ,,7 n(�P� �Ҹ,�	X�� &�f��$ �)L�, � 0�Y�A� �K>V+����u3���ZS ����)� R���������͋t'0a@���8�C��F%	����w��*n}{4&�@3yU #���8YB u��J/[:��s �O�f���� �n��� .�Xy��Y# �Qh]�
�(� � �A����K �U��C�L2�˘�Q���_ �+�S�0�� �P��U�t#x, ���2��r�ҹ`p�
�HZX���!"0;1����d5�8�^ �������L�  (��l� ���[3�@���C1�@:t� ���% �M�XT� �]�h���I @�(JTH�
� ���A20�:����K_�	 9n�h��L�x �횪0� �Y)�P���yX :�U�䮩> ����Eoe� �V�	��� ���w�$^ �l����nR�j�[��w�;w� _��si�O���= Є�6�R��!�Iy&p�� �E�W�B`q ���K �h1 �����n��� �[��W�� Ğ�L�4��TR@4O �dЪ쌖:�z?>��!р��Q� ܨ�Y�'�A `�(�[� ��ha/�G ���Ֆ C�N�v:J �KH��#" 5[y�l4��Xր��Z���KS��d ���p��\��E ����0�K�Q��/��f����~� �
3��(�� ބr@n��_ h�&�H�W$I����' ���>a�A $#�^i��4 ���EH��.	F9^�"�ӌ �e��dt (�����83 ���#��?\Ν�+�W{ 
�����u��1�������#���+�m��Ђ G���!�YR������e�h7[�J0�BY� ��;�`#� �1������_��XN ��o��SP ֟T���w	 P�J�� �����V_P����9xJ¨ ��kW�H�^ p	�\�iw�� ٶ�O	��@�6.��J+ ��z��ྈ>�1����޶���0Y3�[ )�R����i�"��00-  ��5Q+K ڠۣadZw�@ E��\�� 7��hJw� ��`��הo�� ÷�-�rV,� ���J1X� ģ@� �S ���?B�[A� ne�{� �NU�a3 ���͟* (�1�Z0� �<S�h� � �wJ}�HLK@����>�d� �:)-tvuh�Z ���NJ�* f��{!� K��Y�Z��[�C&��	��h��4ۀ2�R����=lU�u@�� �d�� B��e��6_ ���V� �2���	�� �f�1b�  ��tPC- �^��A= ��������O�F�� x'2��+~�u0 v�ހ�h �[��&,�� !�1��b �͖��ʐ��5�T��`�l ����Z�3�5~�����| �Z�����*�t� P\?��B���Lnp,y �@���: ��$�;.���� +��ܖJu̥$Q�0�[ꊁ� i��lu� �n��QA"� |�)������H)� �.��� ^Z霱��E ��+� C���-�;���� �� ���^ �����8� �t�S��� �?���L	L���c��" � ��zs[� �r��,�Q�9p YO����  �븳��ئy��� ɇ}��.�� ޚ� D� ��jN�eʧx #���5xX�� �Y�`�����i�5�l��ȸ	�} x��h��?2� jI��w��&0�� l
����BU�`v,��/ >;�o�&t �p���*��4�Mu ��ߥ� %��f�[�k;�Ȁv���;Iɕ��� Z� �h�V ī�Ӡ�	 ��W�H� {,X��Z[ ��e����d �*0��a�(P �Z�ь�X�6�@wU���cD���ᠢ� ��Zh.?c b ���	�x������z -��/~� ���2 1"J���} э,j%��� 	������O ��N�X�V V�� �. ��a�����
�F�H ���ׁ��4 �>K�x� c,��n�Y�����`R�����$ f�����Q(֗@�� �kt�~� &�Z�Y�E��ɿ�{Ҁ��6��+M%���@;�L���.�@� c	�(}K�� ��h�1�O~ z��E�	 ���� }! ���9d LbO��l�& ��^��	� )��b(� W��pU�� �MQ���"�F '�pH$ق��V���^���]���0�W!ۨ�	���f��I��c� gt��>���"o.� `)ji��_�E����Q��L�� /3���8�	���
f X%��� �wbz�� /!�	8F �]\��� �^�$P�����"�.(@�`�/G ���t��Ca	���� YT��� ��$*�8 � 2'
�3P�������]X���'��
 =O�2���#-�V�+̩� f����x���� �0��X� Z�!v�� �hd3Ц4 A��n��� �M-���	4;���St�!_�2��֙.�)�cK����@��q �<�� �ܟ����0?�k !���� ��1��̀p ��T��[��X�{ݐ��0Y��vJ���VH��y@�a
�r�>�	�]E�ć|��4� ����Q���m X�)@rC�H �=e���0 ���b�A ���`g� T�մ��5u �*�d&� �.�v2ˁ �I8C�� �h��sڸ� >ى�80  �Š:Y1K;�� [z��c@������ZP�u8C,�X� �y/&�5]��@�s�J�y�H ��+���'��3���u[X�R��I����:��'a {��*I��Z%����,@,� ۈ*�d� [V���_�?x��/����RP�O�h��'Mt�CB`�2�5WA�O�/�H�R�4���8Z� Y�%��Ks��:��� �yT� ^!Ŵ�� �d��qSah �O(��P�0	�H�` ؿaN�ߚ8����ɵ��G� ]��ƍ5� ��o/��^� �Or���	�k���� ��[#� ���|�G, ��B��Q�;=X��Z�+�K���	@��� � D`�A�r*a��J7��� 2��盧]�4 �����j�,����b�v�	N U:�]c�S$AB�y�kJ�"�U b;Z��� ���1�j SBzl`�#� (!�� U[ _�C���O� ��Z�<�� ��A�/!�t[di�Ҫ�@W;�@| YL|	h�6z�\�1�`>�-&�(�W�Z0G= � |������ `8~���hK a� 엞��u�5ew�Ƞ��� �cC�N�� �Ѽ[! l�4�?�C/��
��t g5:��&[K �!'^hr=��(Q_S �k5���U� ������b G���"�Vj �_;&��^6�� |Z�l
(�_���V@���ǋ)� V�+�0%�O��*`	� �����Q ������Ðn�i̴	<�f��7
	�� '�����R�M&���� ����kT� ���K$aV�	/\c' ��wdɲȐ@��@���=���3� G���/4o� ����0� 
�>�\�O ��K��TX� ����	J�d� g����_(�!.��+ h	�ʒ�����n3����u� ��ؚ�[��k=� Q���!4�
��@Z��e% C��}� B1ͬ��z ��pnA�h g4� J��M i��^p�� ��a�T �B���8��y���U��� ����% ����1 ��E�)���u�z�� �U� ;�#�1]��$=�T� �H�t��\� �0ӯ���5
�U���~���|��.�� ��j'1 +Y4�ϣ�`�	u�,þ���� ]+��T_��Uo�'���� �D��$�� J�����
��ϼ � [u/� Pr����=)L�<V\� �2�1�j�0�	���� x]���� (	�W�����8��͢ �rU1�R�[SP�"?XC��0�� aҲJQ��]/%T� "����� ��7���<v-���c��$� �tA�N�d�{[ 0�Z��2�y@ � �Pm�)K�G��(Z"�[�  a�幒�z�s� ��
�/�%�At( ����!�� s͸�\�9�P�r1��2� t\Q�,�Jw� 7�V| ۹�kaT�	 �cԬ�,J� �@��*��P�6� ��,g&��: ����� �.�!��S�p� _�W��� ��2ดtH�; �����$��\ ��J�)����N�5� �ٟ�Zy {������̄N ���A� �a�o� 2���*�C�-m;�&/�1 ��_��
�X�`����� �h���!�?	X��@݉z�z/��;�]X-?� ����% |��XS���0u�����Ha 3� ���'�WE�	�o���QU��g�M��%h� ����аL�	_��Cp3��'����B�y? ~ ��� N��)�{�e\�q �hg 2�sa&�>uM�\�Up�T��R�% � �K�� i[��JZd ��|��R� �p�D]�LZ:J�@��#�� ���N�@� �x�;��X ��>B���3Xi�X� ��v�X$ϝ�	�倻�.�� "��@���� ؒ���jY� ޼�a O�@�P� �^ܒ5��k�
����%� *y����� & ���A����'X����JP�>� @#T�H\�*|E1��-P�|.'�d� ��X�|[ � `M�K�;0�LD��j�Jŝ.��Ap%W ��a�p�e|{:����b�� ��Yw��l�}�B����?p��S��b
詵���v_(�*�8�N?��<fS�-�R~\X��k*�@o�B� �(�	�_���<kw! ��h6P� ܕ)q֘��:����p�o�� S��m�Tg���9��`$z(�8w ���ߨ�� 2���z5��"��p��=�gب ��&�1� Y��!�H GX��/��V �9�З���=�
�[3�zŰ�eX�	 ��q���X��@���>� h]w��3�;����N� ���Y����Ŋ�L�8? Q�/�sR� (�}Z���u��c̀a�K �V���x��I/�A ��N��ِ,� ��96�� >����8 �Q��73ʠ���/��t�����C ���m���?fZ�����(�� �#��ƺ��	~=w���D����P!< *c�1�y��fL�� �Jȝ5a��������[?R�-$�( �Y	�] ����^��'U���Q�bN<�� r�C"�
_ �]�yPv ����W	,��t h��+�v��!���� ��עJ��0 f�%D��� Kt<���2>W Q
b�����ᓡ+�E�;J��f[h�0]� U� �� �:X�#J��;�S,� �	���z -�~�9������fA�\S12��b�Z'���� ����>�Ѵ�˝V�&�9��F���d ��0���Z$:U%	˨����  ���Y	�W	��~ �0�z$  �
��]B9� 6��!�����z� ��ILA0��<+�q�� *� l���� ������(� 	�Շ��I ��t�u h�=�M� �-v���*Z�X`����` �e�l��$ ������p
�!�+��Ea( ��zkA��RV;�b��s0X" �����x�(��aHS�  YP�K�͢I<u0�ҿ���"�	��$���kh� @)��-AB���� ��DΧNZ ��!�\����F���q�<��D��@��g G��,�q� �)È�h�+X�b ��{-eR� y4Y��a�.� HG� ����d=y��� �Wvv�o� �P��'��t�����*� ��#\e���Pئ�{/��0:�ܔ �X��c� ���(�>3�� =�+ fY-qI� DS)�T�z���,���0�
�f��@A6V+� ��}q&lԭ a�C��dfQ�������X� �r_�"�Y�K�0����� F�'�q����_�v���8Z\!� ��P"��:�{��� ���ٓ� 
h`6ӽK���_����A� !�`kTe[< ݬ	��z0�R+ ���r��� W"�D�b�vF(� +����CA ���Մ3�'��� �a�I, w���(�K �H`��1qJ �d_��S���T1��[� �u";!���L-B�e��&R/��H$*�Z @�P}L �9�����=�Щ���>>�"z;2) Z���ڕPS�L|��_� @��Ra�" �A<�+����X�iM��^�yh� �p|�� F�UGd �e�'-+n 5yᒾ0	 �|��/��q����@QU��@�?� Ǟ���� ,�X�_�o�a	\j@� ��0SQs ؤ���} -)�\�� B�'�
�!. О~���o�(���G�|�BA�<N��� �hD'}:w]Sg��θ� z�����~/ �{�
�&��� � }K��6��N ���#D��y'LL% @����* ��5I�N��t� 6��Ý� _�c�Q1.� �#��C��( �$\2�8�f����3���U0� � ���$�3 ?��A���R=�� l^���� S��ߘ�av��H3� �o[��:w�sڃ��3� O#���^}	xW��К���؟� �'��Tv�. 0
y^в (��	%}e��ɏ� ����C�M 	܃��2V`��������91	�YXu��}}t�� �] �+�
�L�̂9���@��'�0=H�LJP���%��R����<`�z O��'�U�`Hē� a�SfǎP���� m��^�t� ���_c�5� !U�]ha\G0�E��{������o32 =Wg	� �&e��� ^ф2��]�9�%��E�o�0�� �)ȫ�! N�;C[� t���h{� �.����Ԉ ���5^��b�a��ȁ�7HPl ����4�? ���H���� Ɲꈡx� �h�\/��t ��vq	���@��zK�`��Z��� �����u �a��\��Oup h�=��1� 	������ ��*�B�`ю{�� ?����s)H �W@S��m0 ����XGq� ~��-�B OUv�!˶ /��#�t?� 0D���� �k9���5 {`��p�? ��u0��e'�f�%(��I�hP�5� ��R���-. �ܐ2 ]1��}Es�^��� V�Z�0;� QT�J��4���5�Yv�� �$���*Nq  �Z��hSK e1��E�� �#+x�� ��`���MO �[���'�� Y(B+��D�E�0b@g�#� �h$("��L+,`�&@�>��]��hN ��iF��a)ATX3�<�pɀ�?�@n�[-�� ؓi��U�V b3��	OZ E��e�x��$�0�1�1_ )�2�p+( ��^��
W� �d���kz~0:Բ�}X&$� �C��� ��N���� ����q�{� ��� Q�0	�(�Àȵ�C S���_��O��Th�� ��L��\?�ݓ�+ bZ��
 �_�)�	�X�"H�K�̦� *����x2 ��:��lj�P �5YL$�D� P��i�� ���
���=� W-��߲ _i�5m;ɨ?�&)����e^
��y� Y��%�{��&gh�J�ͩ�@T5� �΋<� �"ˑ6
n �	��u��� \�H9�h� ��P;6� &�_�7�H�� N[`��/Sh�}^�Z�1 ��nr@��  �	�<g'\��퍜q>.0�(��	 2�� \��LԳ�wO�Ӏ��b� �_���E�9�y�<f-��C� �MP����, oNXa�� q�5l� ��,�f�d E ْ�[U	uy�b��Q�D��Hi ��X��k� ;��� =�B�޸T� U�\������P����� Rf��r�X�Z5���³�zLx =�H�1	� \3����pu P
��l4��a���_��P.h�)���8;�[ w���(t�%0��?�����K[��� ���m$� 	(��;L
�^E�0���-% Ag�l�m ��E���0��� �u�~�) �۱������R(�_&�@����������QU� �i]�\�Xb,=�� �OP�� 1�0f
�.��� �eva	 ��0��oI; ���W!�� �wxAN��& '�\���X ok�B#@.v}c�RC1��;,n��(����r�)�7���GӦ *�JY\z� 7Tw
��� �~V���P �g�x��v( ����=�Հ�D�r�¸ ���7�>�3W(\��)�2�_��<A�t�{�!� [��Ԙ%s�P`ib� �.u9��o�G �A�E�4 @�6W]�����'�.� ����� ]�ᓜ�ϝ �uM�Pm� Z���5�� �"��^f�3 Xh	Y�Do$U"L �`�8{��� �Uǽ� ���1�y)��3	P��]� &!���:�eτ����B�� ���G�	�� �A�Qq>�1�� �u��JH ��T3�O�$�� ��<Z/�\�g��WU���	%��$����h� �p;����� ���8a�����韲��k A�1�0e�$s��ང�� ���"z
=���\��v ��BCy�2�xHP���ρ�/�K��`ޙ�Jگ�����{���� 	�WS�Yi �qM$�� ���GPH�7KT�,��ƿfh�y�|<��� <Y�E#  ���:Fy�(�f%u� �^��z�����+����/��( Y�&n[�8��;� �VS*�s5�'���� ���V�!�l>����Yto �k�'ݞ<�$W���ȸO���4g���,`� �������<��-���K�� \h sM<�����'/�"�V��@˧� _l�uh; ����ىy*��H� /\�Fչ���
�`�RDP9П��_�S ����xs Q ��W���=.��I��*<f)���!�3� ����X�h��F�)��i������ �(ڒ �-�)�� O��Y>H� �Bn�׌���+/�(��:�@&c�ݲ}�� A�C�)�w* ~�1�<#��/ �E�J��� )�k"�fW� 
?��j���c.��>��_ '=R�`�n�o�} D�-�XqQ2{� LYy3��{|@�� u��+�_ (���H�U3�Rb%@\(�tf����H<�-b��7�Pc� �QݹI%�2G��n�'O�yx �Z� �5_o%�� �yP���-� ݢ}��@~��yԀ��dB �Yo�̅1w���M )L��� ����Ꮏ y��P ��8Nz��R@!�E���<
В^��:�H+\�,� ����J�s�=�� ��x��p��S�d����	�&��� �
�&*�]�bt����^.�! ���@�s' ��bjy�"�� 	hFB��� @�8���\" c�RuY-/X M��#蒘�Ѝw� �	(��}�r� �O���$��� [5��_e �Yj����ʧ�ȣU	��� � Ћ2��� �Cs��U��9/��]�� ��1͡ �Zx�{�Y a�
�0g�^�( ް�W� �e�FE�H &��Ѓ� �
@��b �4U0�Y�%ʢ<��)������8t*/��^_��@5Ȣ����|�?���3�{����U*��"�2`])�Zȴ-ѕ� �Md� a��=�	��{���vSR+��s"��%�� !k�=?7� �Ÿ�X�� UlD��) !�A�J;�� *�g�[��R.	\B�؈��%>� �cE� :�-|;��	/�_�����@7�2�c�6 �
�����|���YYD )�V��� 4^�f�: o�h�� G�	�s�;$��,� 3
Jq��lQ/9���^��ڞ�;�ĠR�w+�=ť��AGS񅀺_�?W�w� ����hG����� �x�(慠���g��4��2`SZ+�m}�L,'��<(A 9����G�$��n�5Wa�P?����[� #�\��TV�ct�G��	v~ ��3��[�U�T�~��|- �`���Jy� '	��^�@ �h�H��]S���p�� ш;�1�	 Y�jT�P[~ �#d���� �0�!���r� ��j�n� ��$S	����T�d�V Z��B��� ����hoj� D,�)��r� =���^�%���
> �#���
T%�|� )'�X��Hz9	;�_&�췀�Q�����ᴟ� ��2�Q�i 1/�e*�>���_�8)�zU�� ����׹r �H'#� �>�4�� �%yEF*Հr���5�?� �LR�^X z� qpI�]\�(�����` P-�@�H��������t�8Gy_�QQvX/�YHrd�¾� I����
� #�=�`���H�Z҃���48@����@�ͶW� �鑽�)��t  ��X�# $�'+�i8p�3�Q�Ċ�0Ex/ V���`�� a��u�B �_���!��>�:�"�0۬ ���1	W� �N`k��n5��A`����$C:� �#�_��e V��O�I��?�v �:h�Bu�~ ��n�?|' L��.�]�� �#��R�� {�L+` �] �����Y@ ��_eW �Q�j�9\��������OIf� �ڗ�y0� �\rX�Zw(��m ����[- �e�{��!���J�X�o@�1� 	�w��>�P :2��� "��گ�V �|pz�/�	x�) �$^� >�dQ�K� ��ʵ��ϑ��dk������� g��oW\X��������,��� 1�~ns��v :�!�-� 麾���j����w�cXQe�+� -A�?̫� DC�.�| ��i�<l�J:�U 1�>2Z�� ��۸�ٸ� �	�!݃ `Z����f P�ۓ���] �{,�4�`$9Y�����#]F�b�
 �{~�ظn�� �Rl��#X� $)��� ��D��un ��Ġ��JR��g#t*㹊��� ��Z�5l� 	�}�i�1�{���������V!�_��-�� ��,��M �ý�F]s��@��Z������R} KV��.�%C"ܝ�!���1 ��c?Ч-� �$�^�,� p;+�K�[ Pʀ#��% 5��2MWq� �� �Pa�� �o��D��� ��{��p�0 �`P_��� -Y���E�{� ��P�&: 4	5�X�(/
@�-]\L1��%����p�Fn��X��g	�W�a ��KSx Y�f!ú-� ��h�n �7�ʹEd 1��$��ϸ�u������[<� ��Zਅ�X�r�S��q�8j���� �(�V)��퐘���� ����r�8��e��P`��q� B�u@D(� �3��%�;V� c�8К� �,3�Ф�_ �`�Q��]� �9Zh}���8�(�ѥ	���ΨK�'��Ҡ߇� ���M�\� I)�[�'��Y��ܥ�W&8�. Av0�� �)Ȣ�P� �ʞ$�� �Y���C  �Nشy�� �L�?w�p� �����e�� ������4 /ͧ"%�It �eB�=l-7 ��L,���3/�W�`�L+h�� ���Kt@B��� Uq9�� %x�fn�� �-P{X�]CHm���n�() �\ X�w> ���:����`���/ [�XՊ. ���U������fa�*��/�xj��H����@<^и� ��2�aK ���"��%S|�M_�J��I ��ɛj�r⠃� �GQt�T� d�}Bq� U���6��~XT ���$?�{'~�d�vRI���`Lo�Z8𠀷_�,}� "��â(��sX�����h���&!� �B)�*v� �'\z����B�  �����H|$w1	�W�0�E ���
�� M��kn��� �/�4�2�����`����~% �4FSӾ�� u��_1d��s�Q� Hr��l] ��8GZC<?[h�/0��pBd �!���W�I%_�Q/� H�"��ǧ� �r��9 Zg*=15x�:�UA�O� ��`� �Ɂ�0����3��V������g���� ;��QV?�� �@艗� ��%����~ jr\,-a[ 0]���iz{�`���� ��Fa2 ,!���H 	�@Q�� l+��\ ��/W0 �u��.�,� �{��k�� 4�
�.���y�k����~��S�8ȇ  CX��#��T �"�;b� �[��$|��\	ķ'�c��~TA�οp�f�o�d�� E��v��Y� ùON���j �BS=w:Z�~�i-��}��(� \�0�W� �'���f��X�1GRa�h��z �[ͅ�Z�W �}M��O� Ƀ{�K�J��,� iQ�(�� z�v�/ �N�E]��( � V��,^����]+Z	8�O �&1� ���_�I�.h��=  �KR�Q �ø���Zpl�� �Ӂ�t�:N� �V�X������`�edB� �\����H�{)�h�oq�&�� ~���l"�a\�: 0���� C/N)6��;	 �tO��`� ,����V  �ѷ)�?	<�%�@�z3� #�&�<� wɇ�*�Τ ��(�r�|KS����> �Pظ�R 	Q0���8c� s���Yy  Z�h^\%��Ē�=�  �U�^|�	��!w��ส� ������}] ���Q�?0��P�@GU�<��>���;�b�'��P�F���Hq҇ �a�	�!�p ~P�࿋�&��wS �fp� ,%_�g�EO��K�9 ��W��+���@�oY�`�4B6��N��� L����Q e�b��| �I}�LS+�4����k�8L�1 �Y����1�@N��m�f��{� �\�H��oB��"�@5�W�{_`�`�P	�cVU��f�DP�9	  �_���� �����73 ��Pq�$�	@�-ڔ EZH^�?�2*И�����'��~ Cρ�aH{@>�ݐh +�2�� ��E0���� ��$H���d������� ��Q�:�t �_$�h�
� |xBCT��@�:�#�[ �"�� ��w \�J��uT�j�����z���i#�`\�U �bY��@�V��=D��[	�U�1@k��Sv��^T�ч�%1���'���<��ѫ(��- �S`�}�m��bޢ�=���H.� ���	����s��S��YN�����yX��	H�h �OV��(��������}��y�
%���< s�e�h ��2 �*�Q
�(I�)Ȑ�9'j є���3K�����0��B�m��.Ԥ ���� %�y�� � n�fq�� R���������+��VL��K(� �hj�:=���1� Y�g��,�� :eE{��1�}n�2� �|x����> J��_�� a��p��� z�K��w
�X�  �M��/ ��qI�ly�h1a�ƨ!� ��=�:k�SԊ��o��o�P� O4��?�R8B��1G�܎�`[8p��R���h0�mg�����>( �T��)N	�tPƎa������OGІ����!�f��9��D��U��{ ��\>�� �h9pq%.y ��_��nH��`��1 O��v� 麄�C4� WEX%��A,� � �F	� �b{�B2 ۉ�!�ףn��aƠ:��;p;� �����3 XZĿ؛� [��m}�z�t��	;���L_��K��w`t�+�1ص����>(��xwP'����0��R�i�[�� � ��N�� 1��hK"\ *M�b��� ��J��8�؜P��� �0��|�l�v����(�{p���O���	N�B
� 4f�h]:������ ��[��	�S������ �{�*HJ� ��M�!�+����Q��P�M|� �0�Y��,� �D��j��� �Ze����BXY��A �FɴO�(�� $&�W�I�	�`�h�K� �wܺ{^� I�z��1  �]��	�` ��E��W�� ��[��P��&��d������ �
1��ÒyX  ��Y�J�� ���T�� _Ӎ��kt@ �鯫����7�.ܪI�ay����$(�ޥ \sȚ1�0�^��Ű�\���{ .@\(�r� 2Թ�w�p �P��C� �@�8��r�0 ɰ� W1 �ZU
�ŏ�|-��<[�* ;�!��� ����k �Y��-0�+ %W�2f��d���"��堛�� yg����XZz���'Շ O� ���0� �T6�ؼ�$8k	��_Y��j���$��& ��������0���K S��*�� \��1#�V]�� K����- ���P<2I��)��rH�� �N˻'����(�J��R�_t ����̅� ��$����I�]1��;�0< D�
�P�&H K��L�wxЎz����!s 慗E'��X ��gR��t�3��G�p
2�|� lp�K�F���e ��j�[�� ��t�~� �.�	ҋ) ���Hq�;�s�c$��p�k �[��Z�9� p�3K�� �������n�Q��U�����/V x4ʄ��YJ���Ê``���s ���ކ�� �T�|ZJ	+\�� �/_0 =�h���9 +��[�� �Y�i�N !H�]d��A �\���N w��`��� �f�Y2���.�� ��,�!Q p��} sH.���z��{�[ rq ��i���� ���)��`!M3�x�{H� �^�0�� ߔ��nD@�3��&F� }So�h�ͩ�c���Cn�[; Ȝ���2�>J����C�<(�+��` ���i�Q�@[�� 'D؎��` �~X��P ��MJ�_�Zu{����(�04* ��|�D�6�� V�~���/�� Iх���O�� �k#� ^�P��ǐ6�;�8�_��>�-��)r�2���y� �!����U����� �?�B� �5��
���Y+���-1��,> ����/�p �])��d�"� �g�hz5(|p� ��[�� ��h��j>�����T,��&� �̺J��h�b@��$ M��mK� �Q�����jpu+{Bw�ʂ- t	��Dg<� ������x�;P8��!�s�1v��C�U��YP&��+ �E]�@*�|D>a}(h�{2'�YP�1��] ��	˂� ��¯?_�?T։��� ���r�^Ha��`�(�@�2���	�<0hmHO� J�ͅy�r� 0���� �$4���% fpm��@�����xN# ��"KZ��  f��h~�T}� j���2n !I� >�<ZY�����e�r18? ����z2���> R+��[�1k?Q�\���]M �!�_h�r� 	ŨP�0� ������ �8<;E�1j����l �eh� ?�/��[o@ nJ�U^��3M�	�:ڡs����#} ��-����� �7�D���� ƈL��I��ᘜ 	�"����j �=�-� *��Z���� �j�� ���2�O i뗀��ߵkuҬ�b@��U �.�V%K� po�D���x�~�@(�~ J0����= : �Ӹb@O ���� �+��0�2� �����c.��h�8���k 1�y'x��: #ۃ���� �.a]6�i H�$WP�CеV���Ƀ��#��M�� �I	3�� ��� �-f�}/"��輱 :(�*d�w �]-�O��`?rH�6 ���D]�ϼ� ��Qk A�h%{nV �G��'�1] �ǽ��ˀs �AL'�/Z�����`q ��4�D�ѓ �"fk�b ���M���f��m�B�d �3�T�uZkC��q(���\�" ���{4�Z�������&�j/�E� 2�����*(� ��X��- �Q�hHz Zږ*6�$f !������ ��hN�� �m��{�o$�����0�Y�E�� �
�� �� ��2}�	���������W�{0��b�1� _���oAv ��Y�G��Wyp� <���9R�h�J�.�e� ��,��uw� x
�\S#� �邎����W$Ů��n�0LhK���'uHP�	Q ��8xZ�5�t��%���ӝS���*A��)H��`�n�;o� J-�1{`�C� h\����J s�.r'�iB�z��8��8�VQ�}j��l Aֹ���p�`_�Gȵ �8�-�� @Q���� w�J�Y)s� �	!���
 �ܩ�-�K` ��Ps��� 0
�|�� � S<�/�B�}�'�F-�&~��� t��떄ո ��FETR�72����@./ �v� ���*���,U� pa��, �����x�tYr��u���X 	 �!�"A(�}�i����3� �^ ��"��#�����g�� 
	U��*ة�a�=Z����R�0�Љ�%;���1�/�{�<	����F��0�* �Z՟U�� �m��[j�X�(�ŋ� 6mK4Zʢ N��,�CPy �V[����U���p��s�?�� t,�$� ͙�3_c e̪��Y +����� �{���'SUwu �Xq�m H�F���#ݘ[�A�����p��ҋ�E�=(�XD ��e�)��.�OU��؉�-�} !����$��|���)t��@Qhu� ��X�A �z���PR��;�qm> ���u���2@��
^ ��}���B	�~㈊^�)�� �TF�m���k&�=](�!	�y� uF��)\h ��i�"� s�D����� :2�6z�H��c �he��=�' +���� ��a�YI* �_V�>��� N76��(% �}��Z 5V�&�#�/ ����Qw��@�+�h�W� ���%3d� f1��W�� ��,6| �z�f����I�@?�0����o as �BI�^�� S��,���'�9f��j�Wb7��1p� �Z�V)�^q������p,������ � ��� )!�v(j� n�Y<���>߱1�;��ѡ����� ��0	�/GQ vM&�P��� d��K��ybH�:� XZG5�E�A�+�B: '�wN-���;�,���5���4 _��ֱ���y ���)� |� [�@���^ ��U�f���Z�E�R�&����l�@��z��ּ@j +� %�,@��� ��-��S�:d	 �h1�R��+�� AUY [S4��@� ��,�j2	*>Zh�w�޲@%�N��UXP`u��\숗�)>@���^� �Cɉ��M| �Pt�bA��\ �VS	����0ȉކ q�3L9$^���U�m���.�� 䂈������(J��av��hw��c��ѐ��lf���h ��a+�
����� M���cژ�g�<Q �.��^~D� ����p����Y`,
�;�� )��o�|�	�΂փ ��Y�\/;ލ�?H�������c
��X���_��r����Ӿ�·lN� p��P�2O ������ �=��/^QA�w�<�  �j�a��C� ���B� ���-�.�� Z�و�D{R�L +֜�N� .�k�T�5�`���+�� 1�����YD�� ���齣��U*�n�脆�> �p������h��� 3�_J,��(n7O���IM?f�{�ԣ�^ s�Z�g�r �)hF�G�p$ ����� �b�%�) �1�\� :8�^��θ% ��0�>��i:�L��y{��M,��@�����n��Y�@���%��@-�^@rY8��� /#��!B ���\ 
�S0ջH��[��a��f ����@;Z�a`:�F���� J�W�� G��\�_� )���YL�[ �!t
����G:���^� ZR`'QW�}_=�� ��0ӽ� �$�J&�� ��x:ַy_�@��+���p� OȘ���E��:���f� ����R��HN� (������6 @�!�;��^���A>�����}�r���q{���̧�����.ݬ�0�Ņ�XS �>��lcN ������<*��I�`�� �� %Y��M��U��Ăa �B!�Y��� �-~��0�� �&1�G��� B[�ώA8
 �z�D�!>��NG��r>��� ��u3J��� �(0�1y�LXn  $g���}�5����&� H�-�;k��dl���K�B� C$s�� �H7�3�Q<[� ��^��8wi��C��G.�`f�� }7�_�� ���#|4HG(�����P�C��o�Q���S(q t� ��0ƽ�hf! ���P� Ӱ�%��p. ���voB� �]��4��|�1po��0g� )-�H� KX���=�倨i���� 틬��k˚xK z�"�d�p W��-�[ a�)B�^� e'\2��� ���YOf� ��*�/����0x�`"'(u����O
�M\	 VhW9q,KvɄ��A�)U"�;�̟&�����i� �
A�^�G��j��a���h&/S� ���7�y� ����~_} ��j)�R� �8�氂0�9��&ȼ�r��\��j�O�f�ʝ����� b�>0��G �
� ����{pc���Q��1  ���+	� �l^`z�%k �Ȩ�U� �����- ��P�Y)�0���7����c�!��?\
��%�M��{�����6�f.�(� ��<Pv��� 
������ ����n�!?I�=��%[]d ��q�­U�{�@pD
.� XYZ�%�� ���] ɩT;ń���.��#�<���,��h���Lh�@41�O' ��� T��*�v ��Й!3� �/Y����rS �PdK	�� gq���z5 F��0�V�	^u���ȼ@�H��}�Y(��S� ������ À�~��fR (��־XH� ���ĭ�� �%�x-��� �������'�}/��S� ؽob&
@wx���_��� {� ��k���z  �
�㰅� qe����4 ��t�O��� �*�v����� ���j҃��>�@�ޓ1� (�^�
O< ����R�1 ̼� �X� CV�u�0Y� -�5ݚ�w  ^f��k� HJ���L�!8��޸kWƉ�U��� ��X]�1P� ����?w[�@m��J�,��q ��#�Q�"w���������`8D1�"|)�#�~��� ,�L��^J ���2�~>.K`*��$Ip) #؁��+�� \�Ӆ��B��"�E�Q	 ͹8�qJS���B��� �.��P� }EF8*Π�-�>��O1��~ej��y�\z����� �Dcsh�� �Kο�{  ������W#��FJ�� @A0���� �Q�Z ��(���{ gY~�T��� k�
qH��Pn'�	uq�z /d�Q�z�=�����N��� k� �) �_0��e.�(d� ��1�;�MY���!��{ ������>~H�>�2P�� ���v �{��z� =1�
X�b�<dp���^�3D���	�&��� �\��;� �z����`f[�Nbʿ�r|^%�8� Qf�չƆ� K�!�>��t
���h� ���!�]�bXR��; %�`��@ g�(i\��m s�q/���	���a�$�V�2 ��!�� �� ��.ʢ_��� �[� )���/��l.Z�� ���\]� ���^��D ~+���}i �0��
  ڋb���> �4��z��R�'�������H��P�/8�9 ����
���V����a� �'� ��@v ˶ّ�r
�Oai� :�W� @X���+�\�H c0���f���h|@�) ��Tà� 9������b�`[��� ����iK� ��d���?( t�Q���}�,P��	�?��Րa%�ev# o@#�K ���J$�a �cb"#�ܘ6 ���MV� ����|\�� ����u �� �$!���%� ��b�9wBŰ���V�P3��,������� >�@1xzC :!���� ~c����B� �1D��$�� �/��V �w�a y�����5-� �b�������K�Y����E����HL�ҽ?`2N�� ���n�?��P�� FZ��;-��k<l��3P=#�L�~	�V���S`�ZLNC�Z�'tH������L �균�V U!ڗ�9�d �s�ZQ� ���4h�-O �`��i� ���<�D�� j��y2� d�� ��߯�9�@�F̊! �(�^�K�� �a���Z �-D'�~�� �\���� Ͻ >�g �H�9�� ��@���Q�<S :�>��[ Yh O"1%��#!\�@R�f��$ �Zo����� ٳ�p�h� �^���޴鶁m��%p� ��ܱ0
��	 3ƀ�Zh
'zl��e�`���O����,'�z�0J
�7�w� ��j 6^-�����'� 霉¢ R�W�p�;�Y.� *����:� y,`���P ��/�W� >���c�Ϙ�
��u��^`�� ��W���)l]�@�<i۞ ��ït~Y�Lo�(�u��@5��I��z� R�S��)H�X� Ts���{� x3���d ��(Ç'�����Ԓ�0��\S �]�|ýp Ga��E�k�N��!n P��U�0�2 t��1�����J����@؋ ;-A#��� ��Մ@�h� a�����ы�� _��e#�^v� �寅髣�Z��2p�:w/:����ACـ+k�@ ��t��2� W�ѿ� ����(2� *��'��NR ?�^������F�2���Va�-R�t���� �X���� 8ZO2���L*��'�u�90X� ��仟�S�����k��H�#T�0� �� �їZ>.� S	W�Uu�� /;Cf�z�&{� I��W���$  �����( ��n3�t^y�}K/��J`R��?	N��������� _R����.Y�C���V��s�x o�r� qc�Y�P �jѝe�+ �hc.:%פ W�@��[V� �L���� Ր��I�'� ������ {�����T�v�����W: �_��G�Zů�; ��o� =@�0ف��N\������I 'SH��J� r\� ���� a�Ǚ�X �P��hjC�8 1��� -[�� 0���j�* �28��#IP xݶ]��&�% M��Q�K �/[�	���b EU�H���� �\���P�v��&����F� "��9�1z�� ������Ɉ <���*����u4��AR ����nj;� ��_C�����4���`� h�_x��'�
�+@�� w�$�A ��7�O�. ;%���F=� ʸv-ј
(��&@�� �K|�u� *�"�6�� �S�'�Y8��N��|b�pq�f��򌐰-�+ ���'	L2X���N�,��~�L���e\�J����:�<�!d��� �" JZ��I��K���V�W(�O�8 ��\�Q� �����o�� �J�c)�j �-����� !��.��_ �=�ђ�^ �Q(U��}l�8�ʔ��qO����(�@�-���YP�#�� �]e�Q����1'� |�!�� �a����
 [��j�P͈t���°�_~N a��e+�B� �{Kt>C �MW������]���!� �����bC �q��ׁ�� P	�g ��(�OҀ��� �_1/�Y����R��
�Q.��� ��]oE �-���	�HU�`���E��u�� `����1T+�W���[2���� �_ ���b��R��&�NO��;� ,�� _.�{�� �@��2�& �]��RS<� ���	n Lh0 �`H���O�	�YU
� �iҨ!�� 6wTtv��-V^X�+p ��5�'��� ������.l}�<���h�� ����1�� ?��4�O����Q�� ���2�* �|�X��r �AMG��x��c�� PўViXܗW@�`�"��Z<g���� �n�5��
�`Vt���(־6�����&�a�`�e ��< ��9�!�������i������f|K�;�U �Ӊ�Xc�W�8��l� �E!��9 �+V�� ���,	�� ]ivn��� ��[`�|%�10EB�(K� �+�:�� �S/�T! ���� B��Q��;�@��h`^�v�!�@�_�HDE]�)�;�� Aq7/�,a� N��h%�D  �ɼ, aW�'�Sp�l��]� X��h kD�i%tWz[&F.�������v ,���п�T�$z�� �AN�V��?��M`��3D ϟ0�>�� N����; �k���qJh�,�D�0��}�������Y+O��5�@��;�h bI8�FW� =�L����e�;� ��hI� �K��:�0� �T&�P� H;) �c��F;bN��-#�`����>B+�����$��/T� ��w��� ��t��֨����� �"���]� �_�yJ2��;sL�z=�Y�Ev� �À��'Uj�� *KX�0�� �\����~E(�u���jV�bH�
�^�|f 1�3)�Y,?�E�� ��P�4�® �r ��f� =Jaр�qH k�L���t�������w�����$ZWs G�տ<U �-�uDء) /�J��2�[ ����1�� ጽH�J�& �����fV�xe ��
h�=Љ}� x}ˋJ��d���.T�Z!��\?�D+'��z}���0Q* �_M�FK$ )���[Z� ��b�X� ���1p@�s���Z��z�V:�Tھ I�e���ߪ} P�5`�	��9A�
�@0�. j�X�i��N]� �V��� T^�趾`,���x#p��6�w�2nd��������0-< ����\��J�3x-O����� ���]"�:P׌���<��R#غ� �������s }%'�R���� ��"$�w��
}s��� Qt�|�\ 0�D1�∷;���S�ѻ�3� �@�Ȭ ��KS  �\��,t+&3�竤[%���� 4'
ס彻 �$�Oe�S���@��m� ,�
`�� �ҪCN ����'�E��� �kB�Ф #���� ���� H� N�!���t� m�XM	�[�� ��ʫ� 4�3ǻ�� JЮE=����@
���/�6��ඐ� E0��'�� ��8��k� �d�2�+�e��R`��z��	�ڈ��O��������/�d�)�� �����M��[��? �O���^�P�ÌJ�� ,����~�F ���H|�v9h�p��RB 0�L8/�^ z?�ۉ��� ��vr��gl ���K�
;P�%հ��ċ �ܩ��ɺ8�� )ձ��dPM�� ��3�Z ��ڟ�PcS,6. �[^����v&����6pA	�Z�� �M!�~p\�# ��p4&�0 �>�������P�_ ??	b��Xp�V/��k<��T� 	^����@�%�0^��y Ÿ�7 u�)�#�X @�gRN�� � -(�� pi&X��� ��	Pu�5\={� ���Fy 󗄦���9�� ��_PР �W�4"�z����
 �Y�~>x�޹ ���(<� [!��R��D{�G��tH�Q�S$l��K�- F�����.�3�;4���Co�/
Rw�k)J�B* ��P��'���b�2I�#1�f�����>Y{� Ҋ�`�V� ��C-�9�0�� ���^��q ��b?�}=>t1"�!�{��.��j ������=��@洅v �&se��� ����˂�:�" �!�U�͊q���������L�� ���>a	U6 43j`���B ��;��[��$�������	Y�� cJ3�R;���Bݸ>7 H%�G�@�$ x���3� H�/-�NZ���O����:���V@���0�M����K`��� ��'�D6��ټ1��. -�'K���b��Qwާa���x!%|L_? �*H��X�D�@�Sy t�fP��U�! ��o���	9縀���� D��G�!�` �.aY�Vʁ\�Ԡ�	Q�wso ���g�On�����Z5�  �P1�$�����+��H ҽP C��	0�: &�*�+�� �^'�My� 	���~�� #�P�p3�d�Z��� &*�c�>��pO hr'�t T���8����� O���	��9��+b�����f [ �w� `B5����O ��X��	�o���ϣl! �����>"Ov_(��]�eg2���Ъ	w ]�hR�U\P>��y E��"���H }���� '0R����*���;E���� yZ���, �Ҳ:��	A�>�	Y� �V��k�TgN�O`9��o:P#���H4�>��w�U��,ezU�(����Vx>|��2���`c�/� 4��P靗� �	9jH^t@J�ˁ�FA �l�Ӑ�r ]���R�� ��0xѐ��T�	�����^�ꀭd��[ P�AM�Sb� �Ł�j� 8?�P��z�|�@���B ��!�>/�R��^X (�!��*m �V�P��d���\h��yx�Z�#��ǈ Y��	��0�_|2���}B� �vhXf���^��V�:� +�Izw�t ��.�x�� n�+AZ1� ��S_p�I(D�l�(h�2���Ҫ�̕� O�8�ɹR L�(��bSL  }����G !���A� �<�)������\��މ=���M�eH0:�l�/ti�uQ �Pc"p�O ?���ؓx7��/H�""�����*� y|z��) �0B]�+Ƥ���k�"�Mja���]�8 4����I 5�0f�ݴ ��D?ae+] �It2W�K� �'�/��_;��	�R�	�� nfpX& �Z��$;�.����A�[�!@���?Eϐ� ���P��v2>�S �ɻY{%
��s ����y� �I=����/ ����N��NO��%���h(i�)��|\��	_�1��@� �[3�Q��� �ܲ�ZY�A(�1g<pȹ ��BK�� �Wō�d� y)�J'�� ���S	ѩ�� ��3[� �i�]X~? ����<�	 �������u=Ĵ&��5�Ql�3H�1�� �q�h�	 ��X���[�� 1Z�R�8P��* a����p�-bx �)�7o VTNX�� 	�Y�r�bI9��j�c��� ��%0��h 9�`�L/X b����N 	*؋
�=�/��P�` ��5]Un &�����'�F0�Z�� ��7g}�4&��� ���`��YQ��~�y���ȧ��	��0���/8�� Y�3ퟢ 8#�w���� .h_�,!� �H�
�5 �	{�t�P}�� TA�HZ ��+B�� n ��_�� c�~h�x� 4��`ɢ� ���+�� �ʿ!���,,Hx �5��,A� .�j���k� SR��] ��)ſJM�y�����������w�h ~0��\�͟ ĕ� l� ����p��YD��h���
@,�> cr����)���.�P��?��Q�}�J�z �~�R-ZP l"���C ������U- R_0X�M� ���()�- <t�������>���{ {H�* ��s	�k]�2Z��9��H�� ��%�� *n	���"5 6^�ğ����3�@o��M�� ��u�X� H_�$��.=:߰AcL�q?`�� �H
A�8�1��r :� ���` x����%� G߄��?8 �N1�
�)�	SYW���� &k��1�鴿〲�C;/��TR�Q��t�rA`ʮ�5cD ���'�� �X�$�]�}� hu&�a��DP�����O �.'n\�/��4I�a��|�8��Ϙc}Մ .%��� _�1ph��� 	����$�� ��Fi_W0�u� �1��g@ �)�%�z;�$8ƀ�	:��E6���A*�d\ N��.B��	0�$�D`� �?��Ro ��;(à.�'g�J�n`�O^x�`��ch�� ��>3Z�L�����c���� Q��g1�� �n�Yŭ �����h ����m�C^��g���������X�A @�L'/ �C1��}�Q���	Y��[�����m��R�0�O��zk����֍�qSmT{0��_ҰEw�"����>��z����N[�����(��� ��-�!f�%�:�G�tu��@�f ��މI�\ �q`�hCN �ъ2�T�� o=-�Z��� X0͢�y�KT����zc4{� �\]�����q��� BJ!�X@]W �4��"��(ԝ�s�݊��`�^��Y�C�#�h�%yO'�>��� ��io6�4�� �|��dQX� ��P�3�U�w� o��Z�˥��Y�,��X��i *%Q�Л8�;�[�Z
�!��& +��1�� �h;���cU��%��x *��9�0 -�B��V�RUP���s	X�����1�K.�� �IT".� �E����` �cJ5�^� ��!Ƚm� ���9�E
� W��"� �|�- ����&1� h�u[\�zl	&H3 ����O�� X��^�b��>`����)ؖ�xo�@=�I��D>7�1
���v�	�^`C�< �PAU��j� ��K1k�� �ŵ���/ ����+
��� �Ľ >����� &��U���Q ������	��逾�2�� ��s3�!� ���r��Q
 ����ms�������!� �a�K��Xj �։w3W�� �cÑ�ͧuo �%#\r}) _ ���Q^g�*bU �	��.P� ��k� �֧[���z��}X�)�x�`���� �E��< !}/�SՔ9�ҵ�R��K�}�  ��LB(Z� S�AJ$�!�QR��t�� ;����e:�� R�b��S� �Y��x��}� �y����  BA��0/( ��T�� ��B�� �RD�CS�� �WsK��t �l�(���- �G�:*�z ��@h��ٺ�0� ��x�����M��|� uWШV��^���~�5����!Dź��c  H �0(�%�f��[֛� �S��YJT�����Aij ����˾� ���7O�a30�u���C�x��&� �����Yh�\- 	܀���!��Ȅ� S���2Z�|+ r�17uOzr� V��`B��$
ؤ��yk@L�qIɆl?���)�r~��x�B +�N��=���Q�����f ʙO�rрM��\� *3�Ӛ�C������~ ��yR��/5
��U�K9ݧXȢ� ��(�0����	ڀ���[:���+��;��U� ANX���]z�	A
��T�=�>�L�x �;�i$�� VJ���?�;逑��*Z5 ��]n�~� ����B�f� @M1��/� N(+ޢX�G wK��b�#Z �0ö���|��[ �E��`�9� �'W_�\K�-�����vm�����
��	[QS�j�06'�08X� �3�L�Β� P�A����E?�Y`�;� �/���� ��R$��~ �d��a��� �p|)�� .�v���#AW*K�s��~ ��Z�b�� S����:E��Z��ǿ`g�!`F# �Y�F��8&ɀ+�y�m?}rX� @�S���� O�=0��c]`���P@ �����S ��f���U y�x|�l�ܥ�}��@ �K.��	h��{WA7��U�VJ�O� z|{��4�$�s�>��� ��cP�ɰ+/�!@���^]������@�:�N 6W�"�� ���A�.�1��r�>�� F#�"��s�@Հ6� XO��� � z�Y9ł] I��=�\� 1�,����� Nh'7)�� ۄ�p��W "!��F�E 4�14
 N8�O� ٖ/W[�� �a�+��� U�7�0�O�����C��X��%L3���j:w�k��n��� a�`=��>x��	���.�2���Y*9�P�1�f!c� �l������@@-O��Y�<�~0܋��*�v �yഇ�� Ju���޼	 ���L���^�2�8=�ʃ ]/%���� L�-��-�b|$�v� ü���  iGl]�j� ����5D1 �q-�y��%�
'��� "�O^�E�� R�0�{� hN���#� W�*\�%L3��5 4���K �S���c��� M�]	}Y� ��y��-�� b�V�<���kp`��C���)�S�����׀U�4� �Z��_�>��&Nť ?C�ׅ2F�W�<�+���� ��V�%t�� ��F���<\��'_����0 � �ھ:v#��"۱�*�.�U�Y��N�6�е4��d&� ����
 ��t����k����\_� S���� O�&�=�_.4Y� ���ɻ�u�gJ��\0�� Q���� {5��&�0�&�?>�7�p1;���At��Q� �0��(�I Pf��'9��n)� �\>�* ���KX ��}O_�;h/: ���$�0�`����h (�5)�L�Up ���KST�� �H@(��,_��Vٰ�.�D��a
?� ��ڝ��2 �Y(�
y�`�����p�Q��[2Ћ� ���G�! �ʎ�;�J�μ���� #�	�D��uL. �N��B�< �x����/�| n���� �ոi�| P�����" X+�@��b� ��wn*P�f�鹀�0-Q�l�4 Ĭ����@���|k�� �!Z����2Y
��;�D����tKC��O ��ǰ�h� �B����Y[+�Z�z`�!� Q���N���L��A��ه��	 �q������[YQ*�߹� '�h�� ��9&�	�7����[���� @�͘k�n^��Y��2�QA��=�Uģu^�hB_&`��> � ��T��5g��:�1������/pT� {
��� Z�|4�6� ,b�e�sP�v	sW y�x<�6�%�$C Ғ�BUѱ�mv�J0��T����� |�!�R���U8�ܽ+�]�&2���@PS��4 �fQJ���<3-߁��
H� ��~# ��/�E[�� ��R���2!�}e���;�����DW��-`.�N�/Yp���gl {�bT�(O� ө@H5n-՘l $��]3`q ������J 0��6�y�����@�a���	�y�a^U *K\��r�������'��UE�  �[��m�?s�7��������ເ(�B��9�P�X	�@���� �7d��f��,�v� �RM��� 8�X�����e K,C�}� J!�[ƽ|X.U�N )����b#�����㺃�F_�@�#�ɘ� .)�p���Z]�� ��9ʪA W��Zo� )���0	�� P���R��W=F�� *�_�P� ����OS .�w�a��+ ,�i�� ���Q�0�*��x�B����I �$=|e%~� Y9�@��� dU��PI�X��w Q1p��F^ ��D!K��<� �/��$ڢ�U 	��kdY� ���:]�� ��&��Ih�� OY#�}��� Ń\قحv X��/2� -(�W�����p	z����3��P�ه���-�Ð�w�(� ��V�����E�Ⱦ�U� �jp��X� {��2��=P��q#(*��'
ژ0�`Z�� M��`h�d� ��#�}n !�� ��1mrk����AY �N��G�/w�P 1�V�\.�R �x^�ѭ��u�96K�;$;}� Z���(��=~�!ß% �� �6� ���!N� �Y����3X� �^����J����0�Q�j�.�h� ���5�~ Z��#�P��" � �� X1�hZ(�|��5L	 ��� vS@�/^5�4�ޭ���e��O�zZ���`_T <M�������cKq�y ���r� ^.�RL|��b`�@BZsF��Y�@��\S �ꚸ�/Q� �I��V�" ��cA�{L!�y�9#�i0�f�}��� �1v]��(z��B.}�O�'�� ��gK� $f��(�bJW��Iv�B!�@ _�`� �yh�f�� ���2�[���"jn��`TK�) ��3�"W4k *;'�i%
w���sa��#����?���-��`�kg �V��� �1�04��s� ���G��] o����� ͠)�I�X}��e��p���'^�O(�0�<Q���$��A ����]+� ��ℵ� Y�<[�Ch HW]LD ��K��#���E����[ ����r��:���%���aYw�^Z�P���� x�o#+$�@��Z��� '�KJ���
�LV:��X��� 9bh��̲ �����^ �g���1o��Y���;:O t`�|X $�y��? �K��lޙ��`j��� !I.�˒� ��D�rg_K�A�р�/@�1�\�r �m�ʤ�V�� /�R� �-��c�9��	 �p#�����2�>���- 淏F3�+ �Y�x��( �_]��V�f�W���u�`�?�'39�T�/ܿ��\PԸ� �U��{���� 𤻓D2�K��|�����ӄ�� z'�&N��� W!�^��� bM�eX� �9�P�[� B%���؛~ ?�_T� a�T�U�$5W� Lh��>.��_�k�伏&��> �a��\ �B��@�[�'U>de{ ��ŀ�p� ��P0��&���	���է=�3�UT �[v�8ʘ�&
�a���] Q��ҷ���NR	�^M�Y �Z��ֿ��ѝR���x�B D��[Ԥ-� ����� T��)�Xh7 b��͚K% 0�U��)j�#�n��+rtc x���ή���j� -��w� ��EGg�f� 4L\���� <U�x �K��0^��̋3��P�� �(�0�j�� �+�
ū�J xNѮ)%n� Hd���I3 Y�q0���SE����>���j��\O��ծ�
�������>�L�� �3�c�� �[��Y]f ��(	�_�t 2�Yp��] �vW��E 1{����wt���!��O�|��a �݂�V�8oD��	� w{.�J�����!��9[ݷ;�O�z��@鄽�b 3�}�@}�� 8KR�Ѻ�?���)x�v PV>�ʔ�K�	��_�@/ZQ ��"x=1A>�6�`� �#	�pM �Qs��� ��Rl���#=�~J(���	��`eu� 1��3+A0hd������� ���{�M� �`)[��h Z
�j<!��u���c�s�B�U��ֻ�`'�����R~��}� A�@�� ����.�qh!�� ���$��w� /Ԇd(����Y]Dt�8��'�����L����� �F-��au�V?�� ���-狶������� ]\ �b�zD%���x���*��`Q2�-&��b�Ǹ���@�f�<3ަ�4/�.�k ��t���T ��zBM�lZ ;y0L��6@�fi��1(�[��C�����b= �	WF?'z3u n���I> ��1���S N`���� KD}���� �j$ư��4Z �[Q�� -Y�{� ���wٹ%,^q� �S��( ��R캧]:部	מ����C���
�\YQ� �>�G���	��UE�& �?�S�5 � q>W�2�( ��9'���eֶX>N��Ӹ8��V"��T¯ t�	������WH �#Ό�Ք�0T�Qw W���"(� Z��:�� �E���ݡ 	����> $����) v`��K�!��5 ��^ '��͎��	 |ݠGno Th�+�W\~� 0p�
X�� [� �C%:v�����o� W/�M��P��_��� f1�X U)�E�	� O�QN��|* s@Rto^ �,�J��� ځ��]� W$��p�wF�V�r �)� v�����Z}�ܗ���6S,)���&~�%U� ���[��QH �$��	+�tL�G�s��wg��� ��A#�X  C���%:e �t��� �0��\P�6(�[��`�b Y`�Τ�� ��k�i�$�t� b���� �s�.����p4�E �>'� c1~P#� I�=���� !N��͒ +"} �,zr�'ba���T^}By �؜�e_ 燄��=q ��-�ڏ�> c|�d�& ��FX
���E�Ŀ]'P	��q���� ."����X¶$N�> g �ޙ��v[�	R�*����ag���=��� ې� 2�P
� ���@�������!H��/ā�;wR ���S�� ���Ll]P� ş<�X啖�R`���<�=} ]�)�NYG �����LX, �"����h�z����=� ���0�` ��%�2}�>�s�JE��(^ � �+��y� �0�=%�� j裤��A`2(b
٪	��=��" �[0�Z��� ���$!�2 �ӝf��� +�S��{ WR�c,j`]O��1ᗊ�hw�- ���W��Y� X�p��Ea 5y8U���{� <��_T�I� �}��Du� �^�>5JY�r Z��B�XV)^��j�E  ̾��?N�� V�u�e@ǖ�ۆ�� ����}�P� 3�{�T��=��?���v	��� տ�h��p^ ��i��)�#�Y
�w ��`u�$G�����!���e���W ��3�t�� �UV��q\�\ Խ�OAd�!Rݖ��;�3%#�r�� D8^�M�x�:�΀�W�= X�s, ݸq�A�y K0��5ۅ3��繄(����Y	o]:�GJ ��h��� %3�r67{� t�!f� V	��+��$w_�ڟ���hy�[��WX"���]�505��J#��� :F�<�{Y��R�ѣ��D؇! p�/�^�-�HJ�%� �?��	0>^<� ?4�u� �Р:�� `����oT`��!=�  f[�� ^���K� ? �����{� ��yܦ�3|�/9��	�� ]�������0h�
�c��t <�X��*��5M������; ?8� 
2�Z [+��%,{ $.C��Gy� ��l_��  �1�[Z	2 ��m%�)V� ��Ln� ~���нY���hNU̷�>t�0�s���8��:Z �R2㰧| ��^J7�	\@� P��3� �ֱ�Q�.�*
 N� ��/�J ����̪�C��y��"���;� (�� {a�P��m|8 3��oSV�H\?�W� �ͽ��B �_t(��pH �'1\ eQ��zT0�Y��ʇc� �_��g%� 1�>�(�/� \�h]� �tk��� S��	�X*�@�� .o��~�R_��� YQ�;�< Xy�h#/�, ��=8�N��v�zcÐ�~0/>��B�#? r�,�xY8f}��Dr���h9 L��J����
}� ��U�k T��K�L� 81�,�����- �������p��q��zh���k3������R(���#0 �h�b��������L �w���eƚ�۷[w��4� `��Xu8"� \R+ޣ& �P������ _���^"�1������ �s#�2b �_y�:�;�9�'�qk��_�:sKɳ\�l �Q�����`��U� }%�v�/u" 4Y(��� z@5�ʖM� �>L�(Ħ #�6
&��3!� �0�SE��#��Ჺȁ \�"�S��/Ƶ���U�x@�^?�%� �����F}�Va#����)0����]��@��^ g>還'lXz�-����@��k BH��"d�s� �XA@`� o$]RP��|SL��-t�'� �&�d��!�Ȃ0������> ��D���PH:�U̧�gY a/;1� s��r
�(�Y�SUfP�n �Г��̐ �@�	
Z  �[��,�(E=����2`
�)=�1=��#��eB y@�όh�H1v��r
���UjS <`�г���$��5� h� Ϩ�� Kٲ c����bߚ�lPV�F 'X����!� �h�P��� �V�M�� ��YX��T×S�V%����XR��귰 �"���1 ���e�r��	h����P��)��:�^��@ H�G;��R�� �	,��Z/�w ��@uv
h��%q2A�A�Ί��_��!��� ��FV� �t�ӧ\|^ ��z�!v/����_H�Y%W|Kw������[���) �}�]�ޝ��E� ��!`.� �;(��ܛ �eL�Ǝ�Y�4��kV ���mxAT5 ^;�./h>� r��U@�W �ߣl礰�� Ak���`[��=�n" (��*:3� I��q� �C� � N��&�J ��>��_	EӘ �J�YG ���R��X �
C��p b[��l���8	�_���Zσ:��Fl�*� P1���0�y&h/c��ƛ��4��Y) ꠿+�s3� ��W��X� ;���\Oy 0ӳ�Љ��Nߤ��`������K ��e��q��� �\둎lr> ��H�K��z	��_�2̣�{�/PL��, ������&�(	}��X�fh mJ �齖�V��H���) �#�_hz�� ����(a" 8�^��T-� �?�	��y�����@�jt �	�N�; �*�]��&��0��G��j\ ��sa �0F�l���� p���Һ�6}�� �
��+v�	��� �ň�<�1^ ͽ�	���'9�=��Y�8$�n�t �帨� '�\�u,���z �|5e?�\���-��XE ����m( ���<�B�[0 A��] `���Q�5 1�G�� F��"Œ��1=(�+�k �R�`|4� <��D-O� ǬG0_�S �yRb���I�%�P ��G� �'sh�cÐN�HZ܂W����O6�+d ��*0�E��Y���%�A�9�'����
".%� H���q� ��h��Z !2E4o��d @�#�S�w&�C ��zc1
R���"PK�`����� ��Nv�y^�t�}��:�ry�$��_R����u  \5%��d��*i�ȉk��}X����L ��VT��o�Q�J�ȶN	v�t�D��ъ0��SGo�y0	��[X8� �m@-#�t?;h �'N����%~R
�� �ـ��m�,�N��T�%! Ԉ�Wc��ZS��_�(�/!���z���v�� D���<� ��^*�s\"qX� ���-� ��h� ќ��,��� KPL�' �_l�W� d(��Z�2a=/G����aC�H8 V��+�1Mޠ�U �.�RWǕ� fؽg� �-�G�o��~L��#r�rS eF/�p��)D[ n��5���m��`P a�۰���0���3��N��?��d U-�� 7��}@�* �\h�J9 N �M
1 �Pځ��py ���A���E ����2�!� �1'�b*|F�h�NxÔQ����� ����K�? ԯ��֊p�Ay���X�� t���P3� �/]���ؑM���v� Y�P��x� b���관�Z��j��X)�� {��<��� �z½޴( ZXY�N |C[I�d� Ȱ��ċ2�>6��(�>���;�a�Y�A ���X ��f[��� jk�5��� h'BvY�(oM�qQ ��xD �$�E+H�'?%����h9�9�U�Ǉ���� #O����_q/@xW��+�Bh`~ŵ��S� �Q	���5���0�Y*W ��:��., ���魠� ��P���] ���%'@>軀�dА�} �1 �H�� 6hP\qr` �����L�3���S 0��/q:�gy V�}���O����b ��X�T�P -�t!$�i)1���J�F� ���C�� '��R~�M �I}( � ��ׂTK� ��栏
h����*�`�Ep.����e �S*�/ Hqb	�Xr Kv�^] �
���QS  >bZ���	d�j��3�@��� )��Q�?	{ ��^�I��� �(��р<��x@�w��-�1����gpU� �̏�m7 ��~��-8�Yu��%�1�5
X 	��Hu�n ���RQ��> ��[�:�� U��-�3 5͂c��"^�^B`�� A���+�f�����(��^Y �0<W Q�/�+�~��8�`�%jZ��-H
��L�&$k4 .-���+�Z��_D���2@$�}Z��hX@1 �"�[��o �H����� ���<����� ���J>u ��Έ�8��pM:N���O����U W,bG�J���~� ��!�@�'�-� `�Ch�R�u�ZP��H�����<:�v �|����	r> �DY�!��z���o\��I/:˻ې�J ��_�� 
0����I����)K���^� ��k�Σ �һlHQՔ E���װU@�0q�iɟ��\S�
�R2��D� ?��܅,zN �K�p�[$3Xf �(Կ�� ���lpA� iG�_��. ��M��s|������ A���	8 �!��[8I�����v^ +r��-o�7�N �1A�� z��,'�� ���ҋ��� .������� ˒�b`�2�x�����$�)`^� p�yz&UX��I!�
� p�ׁ(K� �Xh6v��w�s:	ܴ� �}��� ����A ��ܠ�*� ��r�,[Sq�<@��%�u�~\�_�� ��[���� ���T���@L��2�0�s��������D�> ����![��T�� J��)�	r�(�V� �þx��^@~�Q� �KL$�\�� -�^��y֦Is����Bht��N T2��=X�� �(Ѳ ���@zB� /�|T�݁ �������r �i��/���A���.��Y�"�R�Ժk ]=Є�Z�Qj��Bp�[X uT�%]b}�Fw�<���h�r8Qs ���M!� yi��zJ�p��w��Z@��� ����G��sP��!1,��1 ��H��7� �-�ӥ� "0���K �HÌ/�: R� N���Chfu�0*E I�te�Za ���!.bA���Bh���w4 @#3�U���|�. 1�]�\�p �-��sM 'V@xDĂd5�7�̆)��(�hJ*�`���#=�w�a�@�U 1���A ���ݞܰ�����[o��F}�\�+��DѺ\������.� R3�!��Ч�2>@�����;&�K��%�`Iu�'���V��1�����Z����&D9�`Z^� 0�QZ� �� %gP�Ŵ� ▦�� ���q:G�s� �@Y��^�d\�� ";�]!�h Z�/���� 1�_�OP$�����PD� �����! Q+��֭�� 1Ū�wk��z9�*���� r��7��t �3���z� ����[��?�%���_8 �R��0n�˘� &3�t� hr6��Y�i��"�! Q�) �v����;0� ���w��sg�X� �]����_���q��n:���C����w& � ���IR�� ��E�O�� �Y���T� :|x�	��Zq���/�_��WЂ ��v�'��y +A־�n���%�ts [�B�3$ Z�����&l�5�K ������ �G�b�Ȑ?^"t��Z`K0�`:}Td�6o��_"�-1 �r���j�� =J��7>��u��S"��0�m 	�v�N�� .�j���� +}�ͦ� >b2�	&o�Ű[ˌ �#���3vY
���; )j+"��B �_~�aJ� �U�%�d� �A��`� �X.-M�Q���P�W��^��%ͱ�{���u=��W ��rK)��>�<�� =���\Sh� �NV zR�LOs `�P	�Z� ���W(���!
$���R���4������ ���Т� mGɹp�k�B :�ʉ�)�P�0�S�����P�� ������]2
0
Fc�  ��	�� ���n��X�@���-�� �Ҧ~,�w~P k?"1F�+ ���ytw�q��P]��/z�Ьgp��p�( 0���Ki_ �R��,�l� у�S��p���|H����W���'0 �"X1�~�����)� �S�fL{�9�ஃ�� �������$�r����[�S ��]�{��0 �%����Ty Q�۹P�� 3���� 	�V��� ��A�:4�� �,�;%`�^�?� ������ ����QC�0 �Y��U�&��- Q�S��i XY�1�ɖ�@�J�o��� e'��� ����~�ηE��(jǹ��� W �F��o(��$ J�5�	Q3 ܑ��2�YWhB�1�+�u� ��S�\��`X�# ��H�� <�w+ρ� a���)�4<�=��C�Ř��۰̀" �h�6�c�,]VU��цua+
@���8�:��{E��Y��'s(�Ni���ڷ	 u_
��4�� }P�R��0� �|!b3�����V��j�� �Y[v��� �?�tﵘ\'l �z�%)�� ��w�Kq�*�.  �h�� � ��2XZRh%�$��. ��&��<E ��z;C��x>�O���|S� �f��LJ �,P��� ��G��� �T�B��{4 rV�A�9 �R�ظ(h@=��1 �:���܄ 	Kҿp���;ؼ��QRW��B��JbX ��I� nM�d�%
 V]D��u�� 8�J��+ ���� ����|-��0ܐĆ�t �� p}E�����!�9�� �j~p�' 稥X��[>Br�iK 
��/ 7�oO�ɋ 2��`�Z�Ū
�q��I�?E�a_@g����$�HNǼX{ �*fP�6 ã����R����>8� i�\cP���M	0��U�'�o�y]r��<���8u�y�鸘ѠLމ�o�	���Zp(�����o�`l�� ��ᓱB� \u��@�Y� R�Q��	� "��2��Z��>�ր�@�)������ �hA!�j.	T� ��'ͤ �M��9�J$ i��[��O �!�)�ț̰f>����%u��k" �8Z Xݴ_�� �
e�3H� ����SQ"���[�`l�	�*�(��������2��6\�s� t���f?Z�@B��� g
Cb]K��%��Y��RpI� ������<!� _h�^�� 2���.	� �,8�/} �p�]J&�E�қ���t<��" ȁ�ؽ��!�O�T:��L� "���}`(
 ߟu9bP���K�325&��� �
	H� t�:��/�9�Gϐ�Ĩv �xԻ1�3g��AOb �W �x�/�K!��� _�ˬY��T �$�^�� ����lS Ҹ�0�� ��\Zְ,҆?�s�h���� _IDxǵ0 �������@$m�l]�_� �8˰M- !�X�IY� ���+�����6� �&��~a ȋ;�f�� �ѿ�����:� F�5C� �-*t�i� ����Wd�\1� }ÿ� �y�航�mh�V�bݠ-X�p �~
[٭��H�$8�I����2`@�Z�W[�
_����B� , ��.V�,��� "%�3�i F1���\ �c��α6P	��q �H�� X ��1h��j�\>����Z� ��q��x ��n���*�!� ������{0G�eYP��� 
��_~�xv �C��o:� A*��z� 	/S ��>D ����[�� |`b�5!A� ^1<�$2˿>'�U$�5� �G� .���HE ��L72
���!���I�x����[h �4�7L�a 1K�tb~%\ R:��hq/{. ��jƗ�>�:�u���7)�Xh�ZԌ; �-���&� ]A�+� )���,�2��KI��� �BHO�)�0�`E��ʐ� 럕.6��-��'�@����{<��!� ��|�H �4�=����� �'����Z$0�� ���E? ��t3*� �vZ�)�����]�^p��`���C���P� �K���G ��Oբ��� �,��Fĺ ��)�_��Qt}| ��	��Vܙ���/���� ���H�,�c �Yr]0�o1 ��U��>ʿ HN�/͐>E;v���P��z rjȡ�5`� ��?�E��9 �f��jB Y\5Rw��%n!��0��r@ ��lb��_�מA	��e��Fw'�Kb����jW �:��&r� 
�)D�� a���/(� ��f;�G�XO;�r&�rr R�W �$𡃒��u� ���t���%��'�SWw�vK_���l[�<��]�����z�AR�qP�����85(��  h����/�� z�k�.ܮ Ę���~ ����}�1�t	 �_^�f@Ͽ�6c� ����rN J����ؿX� T�3(N� ��Ċ� ���"Z�g� `�*��J ��̥W���_������ ���j[��(oV��]"	 �4qZ�P  �7R)<�x �	(�n��{ ���]!� �����*� g��<\0�\�@P� �2u��L���V �i���p�+ ��!Y��Q<�/ Ż%�$5�Z�� 2��r0� f��Gv�:� (���S%�	�u2� i饪 �)��~�D �Z"�+��@����^��s(�1�?��R/� ��N�hM� %�꿡�
S �x�WE60�Ҁ�I8+�� y����^� 0N_ڤZ� 	�#�� �o%���>����� ����
�w� ��ܲ��* ���/��� K'v�PH�* -1��� �Z;�k�& 2�~�A�W  H"�1ޛ� ��̳J��X0� 6+K�D2 �ğ��	>�����o*�B�v�[F�C9��>�� 2���X�ѐ[Q�f�(���J��ďnF� ��	�_� ����`�����w���J��� �t���� �d
��1 ���@�u� 7���f��:�,�`W^ry �v�	 a�񬖚&p� X��(�B�1� �!3�����������
��: 麪+�� F�a��38˕ Q��+��
o��Ժ� �Z_H��� ����(A*� �ٝ��� ���1�� @��ê��|I
*�� ���b E53�`	 [2��P8����S �'~ VUo,�s/ ��Ћyi#=���� \��W���RY	��h@��t [Z���90;%ŀ+	�G,�� �b���AP&� �������� n�v�*�I{z ^�.���M� �Y��}�t���RI��@ ��+�S.�O Po�h�J !	�> ���g�AEZ�-0w���1\�iX����l�����j� )�߉�dhuw ��N&�תT �5�2��<3� ��&:vL��/X�Z2�h�I,C�^��r"P��Pޢ3�;@?,�5d0#A���� ���	@[  +�ZU�h� Ӥ3����:꒖�[ �W���k��΋��]�~ ��x���`�im[�!���_(�{��'�ߒ����_� T%��|�-tI ��
q$��	����}�諊�����' Sm9{� ��u��i��xQ�����
7�����	 Șy�5�@��7 �'�O| �"���V �־�$y�z����ޡ�� k������
-���� ��0v� ��G$�?	�c	���n�P¯� P���'�� W��d�2������P t�Xh�UE;paR (�i�)����- ��L�/� �`�h� Y�n~@o�� �/�XԳ� �[��h������dV*pjN���	�3ܽ�_�S�����yz �d���S;�ҀV����ְL���ta Q�`�r����� �օ�s� j�-l���q� �԰�rP �D�#[��q�_�Q�ѿ@�Ja�(Ą:hӒ��8 ��������b�#Z[̰*�S :陉��m�2�M��&�r0XSfRp��� ���n��b ~a
 ��� {颾'�G��r��O� s��`� ��$[�#�;�{��0
�	1u���sH5�  �����;0&�S) ���8�z���
x)�,�h 3�&#�$߁ ;�t�RV	 �'�<��� w|IA]2�k��d�K��B�pi �I�˾0�
/�$��x�� A�*�� �xf �5��6;������<���d�} ���3t�9](���_
�� �i�  #���H�� g��+V��D ��NlO�v� ^YBK,�T @�	�MU� ��v?���h�`Q��� ��k�uyA��r6 #�Y����������B�rA-C��G���>Q�t ��4��� ����(x� Z׬܄� ����`+ ���S� �̱\C�' @Zp��v"�LV ]13�� $	-�v��8�]��.�@�� U��(��� iZP���	3�
���S*" ��%!����~��A�ե�,� V�Z3ށ	�G��s��)� %�]�k�~: tQY��w2� B_FU� �P���n� xtZ����z耓�	  �[�iW�� �X*�M<z /�Ƥ�B0 �1�j�����h+� @k�x��ѐ� ֤�H/*\;PQ�q�1R� yVZ�41�5_D�.��pb ��x	)���I�WQ�A<pG [��� �����;� .�a��78 N��zxQd �;����,p��@�w	s�f <+ǿ� ��!	��� P�/
�`� S1�邸� �p���OՉH��!M���<��� `��_?���uED@�[�9�u $��^�!�# �{������ �?NE[AK`�	(�T ʱp X���&�Q� h��d�� ⽒�%�  SV��N�� �M$�i���2�"���@N�0�(�fQ����g%�`D ����8sǤ ���� �����}����/i8�C������*�*��r������ Y�>3ȏ�D��� B�j��.�[� SA��F1 �s7*H�Y� `8佡�U �/�I�#X� (*�C���ǀ'T����?�6`5�*� ��(�xXƙ /��,gZ \�ܬ�ϖ ��ԉ���J
�ث� q���'�1��+d�끡7Ѐ����h�0XA�՝ �鑞�f�z���`P��!� i�Z�^��+~� `M�E��)���l��}<�գ��� n1 ��kI$= �P:H["
'1�����sh��6�! ׼�^�a���C��bа�x�� ��bQ���u�$� (����A �Rq}L�1� J��Z��jXvB)>'�� C��� +�ƅ��� b ,X��J

Ԫ������Q�<� ,(�hq*=�bC�#����� ;FYR" �TS��y� �%��[�\�u ������� �}J�֍� �t��.�	X�:Z�L�+~����Ka �Q��|i�@7U��3a ����L�%$� º�^_ ä� ��� ����dX2 ��"�K ���YL/6�H�8x|� �!�
31�\��u�ْ�xE&�ZA m����� ����}Re �O����Y ��Z��9J� �p�鞈[� �$]�	^�/ A��2e�  [�J����@��!��9%��� �"PqUp :�k��v �2
Zh)R>���4����$:%V�/@��I\ �&�H?-d�u� ��c2� �P��hIQ H<g �*YǑ�� 锣�i�����Y���̲*^]�k �͆�2� YʒP��- :rO �D��whT j;���	 }U�����C�P<"� `g�$�@ �%*�(y��{ �ཚ�� ��@wOt� �XT�fHF�_��� �[>��2�8��=I`p� k�q! 3�l��]���Q�}�9�
?����0ϸX�ؾ P�� �([ j�5�"�� �W��J�B�]	X����u ��x�N< |�Y@�(���_&�ށws $1-/�Ɖ���R=��ˀ����� ��Py� Ϩw��1 i+�W�4ŽX� g��{�"� �}x��-	��QG�d�ɣ� ?��9��� ������K\K���V L�D1S 2M��������̮���R� �OH^��P� ��'rv�I�lD� j
�3��P��@�p��%_mqa����[' ��c�.� (ͻ&+EhH�[��;` ����:jm �\ ��J� RB��=�x0{ �Z\Y�gP�=��Vp ;�XZ�� ���j�Q��?�KPz�@�a!�X�齈�-k �E�H� _h���B�	ѽ~w�� f)\���� 	��0���\#Z���� �^��б�H ���_۔� ����B�?��n� �0�u ����T�&*�c���A�� #������ S&%tj8�� +�b��;. ��Yh�u*IAР���T0�M�nհ����� �a�S�+�5�`<T�	��Ur���� ��עB1� �q'>����sd�O�_��b@)�# $� "-�^ |�Y2�	I� 0Vܲ�� � @��6Q(�z ���U��� �{	�
Ar0�� 8�>+�� �h�eɡw i|���/���CX �®<� ��h��� 2!�#H��J�_�m*� �,�`���W )��3��r�pNQ��F�/� �\_�ňñ �. ��S����F
���:`� ��W� (�E. 	Ή��� ^�C>�T��S h�'_8�	"��Y�)�>B �@��'i s:���o�$wl���-���kG �����e[�� �o���R�����5P����` 	1���R ~�
X�*�� ǜ�cb� �_��Wޞa�= �+	�h���ꮂ�k()�Ő� T��	K3� �C�^��	����`(H? �P�+ �����)�����Y* �>":=���vv$V1U;} �d�-��J�w ��W�:�� ^��؍EN �>�S=0	[ 3���k�P +��ɔ= SՅ*���^�γ� (���� ��󆽗�������h r%�n,�� ���	�ݒ\1@��p���� ��#ݠ; Js��� +�ة��V�h��a�
�.H�<� 2׳�W �!wef�} �Hݽ��'��`�r�� ]��P1��r� /�eُUVSq�0Ā� ��	!�47 �b��� �h$-��k��v[)��B�@�� ��M�w* 0E���� a_),2�|�b 	��?>i���Ī���Y\}�K���rd �.�^��� ͍NCK�8� ��oJø)�:�A ���F��>��Y���q  .0��� &�Z�*�����M�[�F���U ��x��+����Go�����a����E� ��i� h����ؘ���50�!� @��"w� �G��:J�� �
'�\l�[�� ��RU����-��ݜȱ�K�7�t =���+��� ZU�X!�'"��Ց2 ����K�} �n_+�0� ��I���H Q�b8\Jf�`��"� �!�h�;I�3b�;M�|ʰS 	�ŋ�D�Lb ���XT@H%cQ��	����_+T� \���P��V��� ټ���m:H�צ ����� r�0f��>��4��� F�a-D�� ݞS]蒄h��0� �Xl(Z���o��}������t�`C/k���j�_7l)�>�&�����Ζc�@��P* ��uk�b�h ��tP�q� �,S*a�Ϊ B;���( �%���#� �d�P�2� �wo�� xJ�[���`.HS�V�3 �f!�{�^rki,��< �O�|:L����'z�@�R�Q~, ����X
S.(�Ǝ���A�� �#�� ��}�� @�LH��� ��ɕ�3qy�(�������J���Q}�R%3�Ӣ� tռ	v|�� D�im]H��S�� _��h QT��NW �=�&�( P���/�a���3�[&"�\ �� {U�*� �����R'�p��[����LZ�����0�Y0$g6 "��~�	�W2K�'z����`����ǜ���K� 6��� ���hv><�n�jJ@�.�� �Q�	� ]�^PI�:�E�3���l*Z���?	��@�����3
Z��'P���  ƻ��Hs �o�S>} �����<� D�����a �!;�Z�� �V#'�� ��f%4�U  H��ZX�k� P1�a�"� 0������ɂ� ���P&	�
�T� A������z�Xo �e����
 ��9�B	 w{�%��x	��C |�W��Hor Sw���f ���X�\W(e�� /�?�� N���F5�� �h�W�[�e���V��MD (���k�I�  �x�pM��6�΀��,�� dºو��ͯ���,s����d� ��N�Ɍ�ꋠ�� �`a(�[0� ������ �n��d� �hN,#87$A�3��1w�i����
�� ��"�Z	� ��l��W���31����^B�ɛu�VP��[K��� ��|X1��z'T���� ���؄�U P
o�=��G�?*��0xh��c ���1P/��! ѩ*���K��X���
ɀ5B�H t�R�TD	#�� ���� ТH��$�e >��� �^1 5M�� �\�HpQ�� ^JVo�
�T�&|����Ue ʁQ3�8/b���<rw 9 ��.^ �%�Ŧ�$��x ��@��� [)��'hc��"��$, ����Z! д6�B��*u�Y�3�^f��W �Ň��$а ��(�[N?��^���H-J K��h{�q� �O��D)� ��xy0m-��� f,
��ԃ �M/��x1:Q����3Ы	 ��'*�^wN ���d
���(����2Aa� .�ջ ��pS$I ����	̈́�.P�8{� ����A�(G� w�'P�4����~}�� פ���9���<A���� ��[��@��#a"����� ZD!�� �~���J��}�˶ǿ�&�p� �-����`?S�+( �Q��k�� ��� �-�5 %Om�g��خ��@V]t�@� ��o1N3� ��Z\S �s��! >�(�]h;� �	��-� ���V/\Q�R����!���������0 �RV�8"�4 �1`*MH� �Z��C��Y�A���ap\h z��W0�� %*�2�b�w ����
\���%�mߥ���#���`|�c��� 2�_0� 1��:���4��6� @�(r����S,1���0 �U��=�yp>���h�>Fg� v,*�X��|c��S��+�Z ��FLu� r̒�P*� �7�z�X-��_�����P �QӪ�B �L�@�A �P(K��	B��S��X���p�_ ~;��E � 闥�W�$[�$ G׀'
� OQ"ѹ& �[��� F�?N���  ����# ����0�Xtu ��~��Ac큱�G肚>Ƈ_��g z�� ���[?����@�J����%*����L	I�'�a��`BѶ �O�`����Ԙ� Ph�Ig	����X(ԝ� U��B�T. �ZicAI�� ������� h�k�7P#� �na>��}4��b�+�U !2
��\%�̽�$ �������@� ]O�A[�� ͆�,�+	�Q�뇵�`�}@��_�jP� ��cV d��Ĺ�� :�_���t� �����p�}J	��Z����
��4� ��[�<Ȝ?{�k� ���&�,�	5 'oU���2u~P��KZ �/��+�^lQV� ��a��2�����3��
�U�J������0�w ޏC��V QT1U�x|���]�L��C��0Ο��YtP ���	��� ���J�2� Ouq3��# �ZU *�(�3� W	�؃� [�� � HA���� �S0�3�� sk���i �_�����S�`����"�Y���@i��e<.�	��UA )(n&R�	Q�"��>��X��9��q?w� ����wH��|�M��o�p�f� �W���,V�P� ��X��E��π=�m@WZ��o� �H�8G<+��z��Q�Ե� �h�M����� ��K�w} (�LҠ��#=&� ��)�A1� `{'q���� �U�]eh	0u����0N���K+ �9_�b��
 ([T��� G��{jNﰺ	1eh m`�����b	Y��ŝ��i$���<% ��q�U�7 ��)
�M�|(t���0u� 	7�P4��> �+KGЭ �����z ��S�^��Ӽ�8ܐ~��K �ձ%��1z�����P�� ��F�j�'}����� �w2�] q�Q����a M��	��]}��!V)a�胅��8�y � �Q(��v�!��G13��.c� X	
�_���(�W ~ҁ;�7 	��u 
rꑐ� 9}��uJP��~�U�׽؝%�	$���ܕ k'[��� AM��|�S�F��^�����f`Y 逘���k 6zK� �"\(}sn���'P�0Q�ܶ�(K��8R� P�˱�| j��fh>1 2v� �� }Dr�4��?:��]&�Ys��TL� ~g�i��:zA� ���{�����>�p����,��� ��3��5 kX��~%Z��-�D`�ï�෕�	
��� � ǉ U��j5z�� ��P+�S �4��(\�x&AK ���R� ���@_ � �
t�cC� ����!��� ����Zw>  ��-�^r2 �����
 ����t� ��] M҂K �
m{�2������1a�} kz�X�,'/ g|��Tn}Z ��;�*�fQ �י#��
Y0�����z ���0ˣ`X"�z ѽG8���	&f�Q3�)�<�0��0�	�>�A�� ��y�v s�(�e\ R����x� ��^;�r�� ��_��� �D5b�Y��n�W�����d�/���� ���WlT'�h~}����O�� ��l���R�_0ԃ�`N��j � �!���;������'p�^ \�0�� G$x��z��
O�t� ������ `pk�	\� q���y2h ���z�Jt� �V�	��>���n^�Pt �8��� �[0o,�f	�� w��Ak�� �aj��h�{} ~��w�) ������x��������'`�[h� ,�s�\V�0JkS���_&�[� �E��߯� 4�����ͦѭ R{�1tx ������w�MK�$ wJ�,��� ߢ+�h�S
?�aR� ~��%O��@�1�q+ �H��K7� �Ue�8;O���)���>��4a���G�������m��/ f��t�� �p6vQ  ��IÝ���#��@�} *޿��dӨLP�w ���R�/� a�!,�� �.�F�h� �c�����.�`�l����K�J �zI�o��yU ���<YM� ���Q�}��%)��ks��� �X�A��P8�!t�;`._�l � %,u	�zS �v{�P�� �D����yR KO��$�U� ,XJ��<{Q*�T ����]��
��ݬ-=���$B(�x1 !��кt��������� _�-o��� 
z���i{~ �0�Ԟh� "�9+�m�<�Հ�J���Q��Z4��@�r͸J�� ���&�WY��3�\@�h/^dy= ��{&�`×X< T���я0*⽰!x� Z�J�u�KL�r 9������dߘFQ�`�� �/N���lK �08�>�- �ߠz!�[f ��g@��� 5�	 �Tckn������ �/�.
�����|G���0À �I��\��: ���V@�� >�7a��\ 6N�%g��	�*�쀕�hIW L�>�[�)	 ��r�Q@���>?_��Z����>C�.u �
��	 ���Ȫ(�'���=�T���7 ����5f(-K��@> ��X��� ���[��� ����o �6�s[8�� +a�.�: ͥ;����f������7 �-�v�����ܑ �&b/�@ 3�Aj?Ykq��^��z n�	%e�	IZ�0}�J!˽O���YP����{���@ZD[h�`1P�E�
�p]N�aK�� �(� �8��	�h@F��O��&�[�	L ��b�Q��PY[A�Sp�, �1/�W@�h ANj���&q e���վ� �6�@��E�?�+˂ O � �C0B�X�~�8:р����V� �_
��%� �)��^�{� C�8Hn�O���[Q섀 �����tX� ����x� zZ�S7;�,��{ ֣��#� W����)0� _m�\�rN �"�a#�: G�h�	�>�@�@�Pz'2 ��b��� fB@ȰIA ���{<E �����	��;.[��8��l%*��H�WB�^�	 ��uY��� �/9�.����1��"� ��,�� ������U �h>�J�|����[�AM�p�� ��]x#��߁�1�!��!� �+Q���� @q�YL[P;�J ��O��� �\��@�);ڷ���eE��؀�k��� �����J�i�8&� /��P��`_�i���<l��g�,��up� h#v�!U� �t��Z�	�D��`���|O 5@���`-��t	���% &hmA�q~с���������"�\Z7(��OL ����r� Ԧ�W�/�^ ����XF9b} !��P���<vQ�-���`A�J?`  U���}�� Ї�*K�F�� �\+�%��~6��'����P��	4���ҿ @�D��� u?���BJ ��2�Ĉ��~�7 F�K ���P���� �ӽ���(���n�1Ё ��C�"��_zvO��w�|b�^��� ߽�)��O�̀z�{=�������0I�p̤=�N �Zy�)� �u���'�<�����,Y)�X(�^�����c��y IfAR�,J � 9U��7� ����k���������^�C)�Ρ/콃ȯ2s��y�1@��/�� �P��Q�k ����ں� �`��5[C�����Eb�=���Ե�U��j ���YSO� pm�?�~'� V�	B��`�e^�m��|dh���x��� 꼅�A|&>J5�rz�ހ�*%�H�� �S�.�@ �o_���Y:����u�&��0�� (W�X�� ��qd�z�:����W���-��;�>5<� B9=	�n �C�b;Q#� ��ǁ�$�"k��4`��F ��o��"�w� k�X�#� �/o)��aۿ	, 0�P����� �+�!��`��M��w�� �Lg:��Pu�� �)#�Y���-O����+�& LPS�$ #�1K��b|9X����� ^/�� ��������Y����b�t� z_��T<å "����{��gQ�v���F �[����O#�_\�b`��(�+�	�R�
-� �)�7� ��Љh]#> ��Z���< �n/��� m���ѝ~I�Z��r�@��W�'� ��h��9�����g���O,Â���� ?�Dhk��p� U �S"��^ ����an
�0��v�;� |�/�5��!���!A�3 =y:�����А^:�W SV-�BH 0�'��X� &�/(�����{Q�ð�h��@]�.'� ���)���<!y �$Z�T��H��� �����S=�| �#�R'�]䑿 �`����� @�!�L0�� �YԻ% �{0��N	 ����]�^ -�X����J9��\���8�O[��z�Dd�)� N�S�� ܐ�37�b) �����Ҝ`��h V4`��A�z TP����x �k2���B (�Y���%�t"@O)�+��� "�膇� [���= ;ؘ�H����	�8�����c��k·�U��\���Ӽ� Y[Za�嶯t
 �,�#	�� T���}��Ű/ h��+��Cyw�{��j�Z	�$�H ��@1~�%��_ �Ө�V�U���`��1� ǯJ�Y�o  �tw	�y�H`�
_��� »I+{ $7 ~�L@�H� z��2KX���X_��$��p"��-�(��C�<� g"��[� �ꭲ�,�T �L�Q�s ��K'��� �C�� ƭ(��5T	r�} ��4V Z'�C\h� !ɀe[���j� `V�	,��Y _�F� ��-��~�I$b�b y���EJ!>Чğ�p�:��$1�ذ
 D�3/�T� _�H	 WّbA�Ȭ��"�k]����°�_���Q� �nҾ�W[A 釗��z{$�c:@��G ��W��]����Q� �� �+-���
����>?X���H� 鹋���� ��\�%rX �(�[�Ad v�*G�b�t p��S)����V ��Q�l��� ��B���� 7Y�_��= �@2�k�T  �1��[�� =�S(,�� �*�A�� }n3��_�� ��6K�P 0ɚD�[ 3����%� EX��]�� mo��q�� s����� �ҳ%�?R L�&r�4�� �	�3
q��a�VX���6R� zŧ�6��x �b�I�B����>3��j�#J ��H��i >8[&+�% p�'�1��� ^閳y��� e��v!�Q%�z�uL��r�� �R��J%�|���-Q ��	LB�u����-�4< J��G�$&'R2 	�+�v� P��B~1� a�Ī�W4 [�E���<w�j�1�\+N��%�K���� �'��\� 퀩�<��L ).��� ��@�Z� 0KxU��[ 1`����2 �X]��F����'�𣂁�@�j�U�<�o���vc �È� �
s� �0Ǆ�� ��N�$ꮥ k�rЍ�R��g b[^�d!�x �\��S� �Zp�V&sY /���حm{ ��c��� w�:;T�1=�o �ͪl���+ �hje�0	 \� ��ұB
���W�z �0��]��M� Z���HG=����Қ�𶹱@��=B�-�(A� �[P�h�E�;	󉤿 O\NP� �ilV��3
r�ZR8e`�� ��i���M%:�����>��~\ �4��f�b_Ł�w��\�DL ��e]�& ^=�����<�2 ��	C���*��M# w� "��^!;�Z ���F_��]����G�(f,KV�"�9`�:� �����Y;	�u)F�b ���_l�J� �BW7�jH�� <�@���d �g�RP2� >�����_� �S�5�}Ht8-)\J �0�w�� ZzO��HB�|� {嬩X� �Ñuן3a ��|o�Ŝ� ��0����fQ "��
& �[�������i@��K�,Q+ŉ ���Ƃ -���c�.��Iq��/���bn� ���E	�V F��4���\�<��C8�X��Z �ҫ��mr�?�5 �7\K��&���qD���	�M}��f4 S�>�ZN��  ��A�+� ��@��|4	 [�uV_�+7 'W1"/�G ��6���`��}?-݂y&�
�n���* �:Q��0�P _zK��. V)�m�&�x>���Q�k� �3X�O  \SV���/�� yC�
�ps���3�A)�pf 1���bJN���;��_ S�F��)g �3Oή�,(��'���5��d��ү���WO������� �7�/�U w�_�h`>D@�"�߃| �ɪ��1�� 7���� F&��Q��%�VWƿв.��EXTu=�߂xw� @F��	S3� P���`�� ��釘�Wvr��`��% �0��� h�@Q�� r�Ts�w'(	 �Ƌ2qZ �,b}ڈ �އ�W���0��`�f� ������ $@�X.� %9���k�?�9ŀ	ݑ�z
�U��� ��� ��	���� �hLƣ�� U�C#q�� ;bH�]ܦI��X�:��; ��\M�S� W])�@� ��293 ���Z� �i�_��sbǕeN������$�J-�^ �= ��� �#�j�W
 I����R�sw��l1�Spp%� �I�5��C9O��Z�1������ ��V<����٩H� �t'�[� � ܱ�0�q�U-"����' �A�/!Äك�.����z�� 9/Hf�Tk ���E��YZ���a,5 BS{W��	� o`�EmJ�� ����Vk�(��xA��u�<�Z�ĺ���[ U(Pڦ	�:���A�~k
Ѝ���������� �E�� 1�Z+ڀd0�[�YXU� �������<�m�����%5 G#���C� ن/��'%�h� ���D� �Q��d,� {�t�`ˢ ��":��P3�@Ð�A�� ��=��L� Z���W!O��h=\�֐HU�M�D��@;-��[ �������؅j��D���A���k�`��� �� Kg�V�?i��h�O�� 4�հ2��%ſ�v��{�u,�� �����r� �دau���2�Р�� 	 !�_�� Ҩ�xY|² �X���D `k	��� 3�i��1��09*� >߾�]q �B�H[�?�Wp�ހT>Y[��N �(��1��c@��ƃ�� s�Zԫ�8 1�(#�}$~8� �[�0��v��zz:gs�� q��u� ��R��i�]��@Z�I ��~��k�1�b��a��� �{q�A�x�{� Y�a	�j�H"J �H��!�w@��(]�z�'<a4��Cː���MXQo �b ��^ ��!*�	@" ϊC�L[ �p��� R������ �? d�0���� F9q"� Q.�N8�ϡ�j �e�l��9�d�U.�`�F� �t-�w�]�^i��S5����Q�g'P�u�YNv�@��� R	��H#{hI�(�"� 醟m�h Xa�Ș</� be��وΙ��-�	�p~����P��#��'�� q�R]!/�g =���*�t�AY�c^y�P.���ʣ8Z�8J��6�)�����<� �;h�:-a ����i��HnM:3�T7��]D�:�����$Q� ��A� �=�V|�[�#� ����o S���O� �Ie��;0ư7:%�`0^ o Q�C�,%$0�� O
�KЕ օZW���;@�rJ!�x�p4� V����� �f��L�uO��@2]Q�@S �3�_���.(π�:�	P� q8W�j� 
��-kQ�� _o_%ͅ !���(J�� m�����-:�hG��p��  �A+������*k���bP���p�v�J.����M�R1/�\:�B�ߔk�h�� `��	2�(��X_�$=k��x�P!غ �'[q˃鎼������ @U�ʹAJ�9(� �h�GM| ��a�{��
�� ��H��'�?�Ѐ�2B�ᮄ�\�OŻ~ ���Z��� .���g ���(N)ƀ�v���~�t �dF���{ ރ�xJɼ �9����c:rU �G���'�`
]�� "CX�O����̈����9-� �t�%�Y�.X C�p�� ��M�� �ӈ��w�����H�/��WS L��" ��@N<���#MEt� .Xh Hk/w��c 2�)� eH����?!� �X S�`�\'S �ː�,0� c	���B$��1&�"ˀ�+[.�� 3�D���\ȃ ��ez�\��=��j,_��)Y]�JK0��.�^ �PT: 	X_ƹ
�髒 �R)}����$�^e@���"�� �K�Fep1�p,��?W�_��w:�"����j �P��Ba �"�^ߋ�� f	�n� 2����Z��0*��+�@�h� �L��0P}�Y|���H�� �D�� c�-�	 hk&1V;�zT��[��@!� 6���I4�����/��� 8/	�r '�����O�2���d�ԉG���J� REk�`{ �H�%Y�� ���F��l ט_�^V���g[O�R��$ ��_|ٔ� �с��k��R���p� �J�O����ⷺ�;K�� ���� �1#!+ɟX �E�šӦ[ J��]B���;Iј���& ]���-�y�������C�_��� �U��� ]�,'z"t� ��M�h�a�!�Q 0��D� [��PW)��r������_t�H6. �uD8�o K�!�)�1� z��Q���/ %F���w���� ��k�6x� �u!��H� Yh273���	�P*�80��$�4�� �U"� �3�/�V�)	�����M ��Z��h&�H{];��Sx�=�DZH!q �Ȃ�:@����|�w�H�8n��!Ӏ��?� oZV���.�B r�lf! �8߹�Б��_����R��j�z���#-�Z���*!���J� �-R�a&�� z����D� �6�E@d�� [:_��-� 	U�!�h�&�@B��l�U8I1 ���M 6	�3߂;�*��u��p� �a�n��0��;v�h�K���(���� 5:�A����� ����X� ������� �(�$e= x����RZk�W6 ��o�� {��>c� |����� K��C
��4��v�v' &���A�r1H��� �@�0�K� ��8� b�e+�	��]��*�'Y�^i� �0ށ�E \H��=�ۉ ��+�T��\�R�ظ(�
�P�'��i�=����U�_��� !B����+�W�@��[�5]Y1<� �����9����� ��� -�%� E+���l �;�aY��Lh���	�� !C�cj.� ���0͘<����>�S��]�N
��0�� �����Ã��o6��[hRA /�2p�����*���N��� �|�qu�f PS����> \�3`��
� W��tT#ڸ���1��u��U �T/P����q
����Ä !L�Y��\S�b��m�� ��V�� )���~��ȸ��0��'�@�$=�x8�\�[��01 �MFH� 7v9�X; ���&��V�!Q	��E	��݄���̭� h�M"���������Qrw���q�k�N�_
���A��� 1��� ��`@���XH$b^
�<u��J��볙� ��R �,V�cE� �����~k ł���7e I��i]L� �,kV���W��/�I��P+O��$`q�Z��Q�X��K) �_F�����r;��؟���� �e��� ���ӌP����Z0�Iđ *�����x �
h]'! ��l �q; �~��<Z ,ѽ0�t=����Pڱdf\@�$n 	�0pU� �|�`���� K�8s$"�\�mt7ˡ��Y��2 pq��},0�'T��&�LI𔋁��_�G/ �"ܺLc��0E�UP��[P�ܶ�.Y+| �Tw	4�n��?�� ��O�D*��z�	�@��%��E��x l �=<-�` [Ϣ�W\Xi !�0��N ��^s�� ��1C�ގ �U�����;�|���p�]�� vL�O, ��%ҡ5��>׀]�ę��p	�S!�L����. ��1��3 ��xNP�/�@}� ��{��bXQ6Ā�U��K��� �b)�]��	ޢ5��½!��X�d HqKZuh�)ї�� ���e�F �=�!ȶ�'#X�W0%R :+a��|2�E� �࡞/� aD"�
�\ ԥ��� �c?�k�� "���y�M�� ����� E���O�'	#�Z�-@�T{P�Q�̰Ap�� Jbv��'(�e�3ܗ���ǰ�|4 *��Խ� i&�Ϩ y J�-M՚8QuT ��/�� �����~B _1��^ S�`��A�>��)��F(�����3@������ �E �d�14���t����_ˢW�� H�$?��1��J��B� l�Z�~m��;A���< �C!�4t� �+��,P�:����.%޷ �-����(�� ����a� D���֩� ��V��� ��Ű��B�� ���k�� �"��3џh  �֝�j��u���@[���\-���?r	�3t��n�`H� 
����y �	!�]�xh��Q��0R
g��R��w�+�TK�Vc�* _$�E�� PD�� o�	�`�_^�x"�����=| �f@���$�	4�) ���J ��
�X�� (�[��� ��S$�!J� �jX
����EW��~�T�^��������L�sX�5x����� �pv��� �������ѹ�|�`��; A�
�*� p �\���9f1��.�"`�Ja�� �$%��  F<��`#� ���X/$ �^܆�{5�9z@`�W! �[I�
� ��;�k�H�b�RU@F�K��Ͱ� ���X���(JUY�0K� ���n.�^ ���[�v2 ޴��Hz� v' �ZD�M͜�Y K}`����=Z ����U��@hտ��;��_ �M�qm/ `�YH�ε�	�[P�p ;0������ q`�*�����U저��B��@�$ f��K��N5��ݺ\`v{�$L%J ���� 1���� ��/��0�����Ϝ��� &6��� �@	�\ ��h s+Q��Z y����8H����2�	�qW��S�ׄ@�e( �R��X�F ��ƽ�Y	K���|��=4� B�!��_� ��T����� ��ƍ�#�\Q���d�ŚBʘ��A� {��� �1t/HG��v����!�[ ]"�%�/LC �)-�Z��� M�7�	��	x��: ���dn ��T�C4N$�R6-�P����	� �m�s��Xh�#�/��o$ Rw9���% �P�Z!��}m �D}s^'y ���e�gX� �@��Z	�� th�3c�&V A��b �^_��v�ʊB� ��.��~�-�E���K�p�{ �P��0�{ (�)�=A�y��� ����ޓ �*-���< �Q���rb� �W��>� ���CI�B �X�1o�#�4l]���TPZ �Qa!��� �t�j@R1'	Չ}���/s� eS"�[�qy���x\>`��s 	�v��X�Nը,ү%��>�`}� �JԂ ��i�:� ���q� �01$j�k� ]>�#���.P^;@{�� x �R����sꠒ���Ho �G��pz���V
> Ǿ�S)�U	/��w .���u���S��P�� N�n~��� �� �-��� sW�����⹬I &����� Yf�B	�� ��$�N�`W ��0k��M�� �I*��;@��Qj�\�`�(�X�O-��� +���bW�$�)Z ꜯI�	,���e3��������JY"�� \���TX� 
+�� �g��[H I�`�҂�>�� �#�<X(� ��?�n�<�,�f*^��k��o���������@(���L�C��w�v 1�^!�e� ��چD��� �	�kIvB� ��� �>�,�zi ��� *���_M�J�� [��:�Q�X:��=� p���"�� 3>���
~ �h�<����)�5�Y!���["��C�؟v�� R*Ʈ��-� q�aˁg �9`̊
[h�� p]/;� �
`�C�p? !˲�Y�2�;�f�ɥ�^����3����d����=�D���� �i���N�!L� �o�� ����� ����0�P1 ��";k	U�8^� 3�Հ�b� 䖅Hl�X[�B��	��� ¾̨P�cA&D�`]���| �2�cZ�O�?�� �Q�)�.�����	V�� Q��D�� a �	�AT�"�p ���鰍 �LfP���Цt$���  ���NSW	�]�B��T��u� �'��#�� vt"�F+߯p�%2���z���� �I��Rn O��2�G� �$V%(ӗq �^H�h�y� 2Jm�&1� �W�"(pݿp�
��u�PVW���!@"�� �G� �I�;_1�/ �@.�8H� -��nV��O�������-�q� xN����M�oR)���5�R���W�)s ���ˀz ҁ�L�9� ��-��l"~����W��S���(��X~� t�I��� ���� ��"h7	� � ��� �d���E�V c�h�7� ��A3ǳ��`zs��C�2u^��0A�1~6��� dP�R�� [�NJ����T �.���2% `�H�А�_ ��A�"�wj�~� �.Vg �H����- �
T	O�U9i��>�q��_ !�.��,C�63� �m�h '�|��� GD�˕�Ux��~�	���9�_� ��<��+��<�� *��$�|X����k����# ���h.���`�/�u@�=-;�݀
����� ��WG�N	 _\�Ӄ+��s
���x)�0e��&V� `X�/p�A�� k.F��� �����P �ƪ�A�
9-�r8�,Y<����!����� ������9�_��0* �2�<!%�
�j��ĵf �WgȌ�'!<�]�jM���k �0Ӻp�N����E�j�0ꕢ�Z�X���G���jy� �_0�9#��~PWŀ$�( �2�\�]�G5��g+0��/&~�Q =U�8�z �^����h �\���� ��n� ��e��&���b��]ź���K" Ꞛ����1�5��v ���Z����& Հ�Y� �+���`�h����� �(� 1����S� ��c/�DoK��X!Ͱ$^��BB�u�|S ֪��,����u:�cI�L�Ԁ��1ڰ�R- �͇q��M ���E|�&�� �r[J��� �;��܈� \P�7���3 Llv��h�� �Ɖ�j� )鑇:� E��	��2t��3�u����&\T~�{ê��Z&�����Ȕ�wŉ �v��B��w��� ��Q��(�Pѻ���y���`D� ��>����g ����E4:+�O�b��A1z�R _����������� h�({��i�݈ N`��	� ���'̳q �i)RuJI� с�6��P ���cw	- �]ʤ��	�0�܍ �K�y) �+�k��f3:!�wuKZ�Ǧ�����`���� ��kPB��.��ѯ�;�d��3���颠��N L�V�CG� a��ȫ���N[�5J�˔� �)x&��0�h�mX� H�Gs����� b��f�^>
Z�(�`� Ry�P��@}�/'�Yf��N8 ��1 i� �������p��fS�2��[�p������v�`��% x�����W� �b�w!� Y�l��, �Ǆ_�A� ���[h�?$�9� �s޺1����t )0�[��h\����ġ�:��=p^���h_�F'� �����fv	]3��~�j��Òp+��_����&�k�b�u��N��4��X =�ZѴ;�+z7 T��`�� )�hc*�%�(r� f�`W<˿ �m�%�)�  �T�/F Y��=��A <e�la^��|hE���g@»@����}� �� /��02��=a1��! E��zS� ���ҽ7�?Cb>�'�_�����+L�;%]�)N`r��b��t:���(����P�̀�>����+�W�Z'� j*�x��I�������<�e 3�O�
� BA��?��0�!�a�<t� ��$	�A`>�� �d���� �n�v23Ҟ [a�EZ,�� _ �U0v�{��ׯ ��9_Q3 o�ˈ�/W *������[�� !�J� ���!�q� �]�0x�* �6V�t�k�}=����X���A�} h�]��p�� �7������L���؃� �����ӊ���\��T�� [�tQ'��hG��Pm0`� g���.` ��	��)� ��X��W��Ewꀽ
��~� L��-g�E�!��0� /�e` �>@*�O� �A����p Օ�:��k i��w��_z��XH�]01��5�iZ��I��@z ƤYS�� ���{��g��� �x�XC�}��f R1��` ��&$�͒Z�C@b�#��HtY /���0�9�>�����N�� �c��#ް�ZHn@�ŋ1 �6��� ���(8���z�� i��^�&GD	I0�ڋ�@	����� {7m�Y ��j�h^Q����P�pF�t��U���*�+j�]=����k�`�� 1[���O NJY��`� ���b��X!D �&H��t ��	)<d�Q,�� 0W��!�b�|�M ,R� x� �h[?�L�$ ��y��� ~%�@��������� �����>�l K@��R�*�B�H�(Ȑ %�-߫�ړ ��� �()����� �n� �w ���Ղ�H�
M�,�< v6P*�R� � �!�� ��j�΀-	0��؀m���� �_�j3t \��f����v�@K4O�څ�� �p!�Y	M� ��������R~8���  �sO�D=����@��ʷ���� _56	p�"� ���wB}� ���|c�VX � #&<�P䤵?a�w�\ 6�+K7���{�?@ �Z\%T��;����_-��H��J&�\�` �CL�9_��d;�i���X� /��p ݐ��:�H4}z��d�������-�e� %���9 �+�m4��� ?=����� 
� �0��� �e٪��K�u}�N�7��=\�0΀��� GL��K�Y��`��� OG ��#�S�,L�������������  ��zN��� ٿ�)�3��ð�0� _�K���U�\����O����B�� �v���� ^�3O� � e���A� P�{ڨ�� [��1�	�. ��O��Q�� ���o�4� ����$��R�=�ꀨS�A� i�_{@�b� X?���)4�JHP@���Hv� ��:�%q��L��^R#aT�X������h8 ���1�^ �Q��T~-q}�$�I[۬t '0�u�	ŷ)��������5w@W0�J\�B_i��� 	}��Uo� x<�l6(�\z�L�� Y�ź���; �m���z����ɠR��� �� )�0�s �h�I�Jf^ 뗈	;]�����趱�K D���wC� g�ӡ�"�.�ZS@U�2m �K֊��n���	c�S8�� yU*�+�H� .dI-�8�b��߻/@ �,Y��5{��A ����	I:������j X��;��W �vz�	_h��[ã��J�!��t��~�^S�� �4�\� 	`3)��z ��ˬ�*"� ���.�( K'�������±4��I[Z W�'l9������0{�6q��.�ěSUX���M�p��� ]��:�~� !�й��*�齇l�+�W�&���!�؏� _� uѯ�|+��nA��8 �S0�@�e��^���,�Zp��y1 �h�V�sb�L,� ����9� ����߼Kv�?���1a!�R0�J;)���B Ȉ� ��-�px� �l��肸��-��/�����P|�L��2V p�WŜ���=C�u ���P[!����	�~� 2��N��' �9��&��o� [V1ؾ�?P� �4^�H�_��=J�� 0�	oh�9 ��.]U��% \�e���X���~|$��I��ϟaF���t� ��-��C��
� �����k�O��@��'�U ��\i/*��yQ���U�j�� ����-Lovz}?��؈/�[� ��bU4�����]!���r�Z�`�������Y��� >E��%B��2�ݵ	 K�#M���}{���R ��ڔ� ��:"+�/�;	Ԁ�#��a�;Y��/�Rf`}Z �잪�L�� �ѻ�ԓ� �H�8cZ�� h0���b��p� 1�Q���2 /"Iw���:u� \��qW�� �"7@w�N<��h���[�Pqc|��`	1u� Ӵ��:�Kx 'e�׶\3 z��g_�<X΀�R��Ϻ;��%jy�� �S�hD����t�[���k��wv 2������1
� h�%�<! ~��"ϋ.� \���g[ a��BM���~	 qS7��0� `�>��@9 
y����� 6��(iI  \1ȼ�% D�$��:�X�����j ��s���* I�a2�� �FY�ҝP� �?0��(˺ /�{HwC�	!0�,���
 �~�Kݘ� �ZCD۞ �Hk#��� ���˯�>�B����,�JΞ�	���ߩ�! VU��~� �gj��P
$��) �1�e�(�f��p�
Q����P �^��t3�j MS����RU ~�	 ��� 5��X�O>� �KQ��!P�.	5? W�y�U�<cO\�;Q���D�,�Mt/ �(��4~%_ |�E���� �\��,�>�-�?A�g��;�m����!°� R��p)-�� _��~� �8g���\�:��#�h'0�!��3���X :���}� Nٺ(��P���J�z���z�w� ��\�VR	�9�"É�j�w@3 ��� �������r�
r��9C�
 �^�H6�0����̝�S�&��@�L��
u�� ǒl�� �����.� ��ƘJ  *8OU�ؽ0 e���<�� �A/�Q��% ]'k"�<�&Q�L ��%�Sp�U��������d�����u���0��"���T]��:+�� ��9�
h�8v ��8�[��l,M<� B�t��\��
� �D� L� m�#��@ �Ը�(�JYH���!�	KD�W2 t��L�������V! G�<����"N�� 5�y�+��4��U@�� �W/� O�� zV�*������N��3!k� uPs���w���`�� b���`>��`�[p �w)�+�ф;B1 U@��3�R���{��_� �o����.�������2��� /�rL�W�= �h<U��F��	]! �D3Ż	|�d���( Pܽ���)� �JD	�M������Oj�[Y+�������Q ���0����t��� f �Y.�� 6:���|� �ʁ����� 1`���*��ҵ�{� ��4��$����bH�� ��-u�_�p�V (�ѥJQ�� [��P+oSX�'Ku�Blk �C���[ R�����h� N* ��u�� ��O��h[ !���xػ o��WZ [A�j�'� �}�F֟� ��.�_hA������� �E)���F< |���^�, �8+�G�� ��>���\� �	���"� 1�y����+nD�㗐��H$�l�� *2�ZR V(�-��A� ��P�	��� �X<��Z�b�֐�GP�T �ܧ��	� Z��O�fb� ���{Y :��C3� 1���.����J N�1������Y�9������J	�� 1������@�ZN�� Ș��l�����[�O��}�?HZ�Ź*�у ��/�� >�Pf��Y&(�� d�Q`��� ����h�� Zĸ
��Kx|) �>��ޥ�( �+��H�� r@b$�P�8ο y���� �JrF`� z%!�׸{� ���Y��:^�s*�:�ؕ�ޑ ������X� �q	�[��� ��'��\?#2��k�e�H 	�X�b\�`s �Gޅ�š:? Mz�ͫ���0<���+ȸ���¿���N� x� i�_�=y�-��5(� ���\� ���}�{u� ���2z��N�� "b���f&	�R���D� �o�U �p�1Y���KG]p���p� O���	 �����
�) ;��(ȅ� &�T8'�� zuZU��r0���1�<������|@��v4 �z!�A�
 �_;�>B?�:\� M���~[ $h/t�� � ѻjZ	 �2"T���-	㰺��V�:�'�+ Œ��tbXӠ�%�&�� &����=� .(��%T� Z�4��A l�����	�R_j������9�h-S������8� ��R�	��� ���0�� ���/�y�{� �h� ��� ߁��0�� �Y[��P �`�#	 ��3��� �� �+���=-)�,���9\!�KwH 
׹ʈ�I� ���z�� ��E�S�� J������ �:�X�g=��kWNQ��Z� ��U�r `�f��b �~�!_�6vH n<:�zܷ ~ON��0��u`�X��̵ �k��օ ^����� �q� �X ]x<یL�Z���Q��n��(ߗW�r��d +8 �H�*hKm� ��U��� �"�pY��d�+�H�'�$h Jj��a� �P]�!̀ 3�SpXB P�/�[�w1�Ĩ)��T|��	2���pH��p0��hxkK qa�f�Z��w�.N�* Vh83�p �Ai��4� XQ�$�b  ���*���C ��=��J^� ��儚�K�s��8 �o Zͭ���"�-^؄��L9�HO�B��*�W ǿ"���}� ���`�� �ƈ��&(�H��1*Cs_%�#��/� ����2�� �a]��\�g��(YZ��s���S��L��c� �)��M ^�Sf#��[H�	�<K\ ��B����S ȡo"� QZpX*K�� ��?����w� _��h��� �d�1D]�X� s=*��6�:-��O0��d'"\�P�� ����2so K�v�G�^ɀ�Z������߀�K��C �i����� �(/�^H�B�l`�R��� ��1X�<��=�*�?�R���m��5.1gА�0� ����Zư� \�~J���?`Ӄ���Z�9)�\�� >�����{T����ޭ��v� :(�Y�aʃ-��l��J� m��R�	 ��MU7`��eoD�$�t ?5���@�:��gҿ1��$n?� ~t�� �j�"��I-�۵ �1��Z����o�.䀉 �]����~��@��RL��i� �f��b� ��Z�,��A �d�1��"��P� �#�] !���8����\�K��aQ
X��#N����� �<�'��W�5R{���H�X$>�ö=���>� �ƀ�^� �z���<�@VKT�0��`ޘ�h)��Ȓ�*'����� %�ի��ɚ ����<�(���O�c�X���5�%���������PL� ���T�� *R�`��Ӹ� �%)p�' K��1�/ �Z�];� �a`�ï�!c��?���� �0V+�hp�|Q�"��L� �9�J[���@�S�V�A�d=,��h�t��_��(��B����&��`� �<�	aR# �z9�_ȉ (H�4JT��l�*\�������� V0�K@�I!Z��U �A��܉٥LS�����Yh&�"� `���w6�݈���O��= ��_�VP!��u����$Ե��� �ߡ���� `3J��5��lZ ���| ��Ѳ�� *�� Ԃ�����x�0i�g ���O�qp)�*���Г� �K��_"^o��� �h�-��[V�Č��Y� ^X"����<<:�}��*� !ك�`U� �����& D�wg$�s �o��/X�u���!���QΊ
b��C� �w(P*
F1G� 0���I �b^��Z Vն%m���$�џ ��W����co 6�G�7 ��T�ykb ���K� ��W��:�� [vQ��;pl���Ќ0Ӊ�U8D��oF��π 2�P��04� .U�N��' �)�]��3�H��p��s�U ?�q�fKg~��-� �P���0 �_�T����� �V!�n�<�^�k�/p�� $I�aNm� T�o����1 �O ��� 2���թ�� U��9�J� O'�T��3 +[��Y#� Wf1�{(~��ʢ�ҫ��_��� % �wކPS�5� �����x �-�XuSpջ��ň�� �"���� H��	Q�2��� �/������;��8%^�;F� 9���Y[�B�u��0� �$J�Rt�}�5������l'X1��97�k� JB���� � 
��K��@ Ff	�]� �1J�*G�)����fZ� ��9W�wT� (���Uˋ3�kN���wY ��R��I �H�z<���.J�` �#�QL iv�YR>&؆� [�
�-� �Ҕsƒ��N�1�[�r�t��P��z"�Ҙ9 �p�h*V� D4���N���[b���`�Q��5�s+j�1��B��h�~U���W� �A�%o��� ԆG���$��@����� 1 eMLf |O�*)� �3l�^&�} �H��&`v��ZI��  }�7���F�d S�	��� tR�O��l�2N!� �b_�������+����~y ���t�	�Y,l`�T�/�n� �(�hMb�E<ऀ�����2]?�Ts�	���c� �ޮo�"K� �t�v��\ ��	Nu��ҘJ *!��l�-h ��IUO�� E�\_��'���h�	£�oC�7��t�� �%zɸ /�\4X�Hy)p� ��1�� � �l�/y p��
�� Z��*�x �[�`�hsr �7b����
:���D� ��C�\�J��z�B �� )�Z	� ��J����# ����a_�� ��И��T���-��� ��H"B�j(�����$�[� ���M� 1龳�"�̮�.V��D�m rPTX���> �l~��W��F'�@�(� �`��)�<�j ���P�L ��/s�_0� 
S��qȗ�v� Q�x�^�_ ����S�x  W�(b�@ ��L^�N ��'�w� ��q�
 ���J���͹���"o�/9pAh %b.�jL� &���a�ҭ �5��ĠR���,o䀸��B��0���� ���] ��_�ܫ� XnÛ��~' �(�|A/j%�-VX�����?	`o$>#�^�a��Ĕ� t���3�1M��o�c��@�֥( _j�0����,�������RD 5���[��0����xG�j�p��^rk}� D0�[�� �����Q �������,	��'�q f{v�[n��r��0��$�.���Ui]� O� ����!�S�z@ ��1 �t�B�W�d��a�&k������?��h��`V���b��S@�ÝL�,��>�R) ��Ƞ�+� ���b%��Y�������_��H ��R���*�gb ��|� ���N���	�`�X���u Wz���'`�(��`]�ڐ J��͋%).�K� AQ/��(� Š�� s1,y�$�3��XY� n�0ʮA�� �h�aV �@��Wc` S�J���!���fp�~� �<0��Lv Q�퇬C	 ]���O`�� R��σ��	��׳�\}?�@	��� ���à�7{ ��2�Z� �a����'�|	�FU�$͒�\�� >��h�E���ϕi����. �و�Q��� �J'[�z���.�������w � �@�O��g��A��	�Q�>B LwrV����v: ǽ�tGQ ����04�?� �K/�;˿��_�_S� �%���6ߢ���A��`�(O��d@�'�Z �� ���R�� �@Й[Z��nH���]2������0)�h�!���� ]@�ed�� 
̀��� X^& �l�>G	� �|���e�~��'�����O��dH��PX��uAZۃ��f �	(V.q�?:Q��R-����p�! �h�8��wv� ��/��[��y	 X�5�y|� �6��0����@V�af@�?��	���U�� !��c��=�&@��\RX�- 4��0�� J��_sT� ��P#شW 	�Vj��/ =��͂���	m~�B 6}bW ^i�uϺm$ lV	���p��|b�_��Wa6)`��"���� ���X��O�̀�]WYu$���	���$�" ���΁ �2���Q�W� >B�4� =��'��?�aF����4X�N� �;�?�fR*v� �ص��U�����w�	 �%-��(���� O\0��ap� ���)�Yߴ��m�U�ZH�h���2R�'=|�I��9A	!�d��{��J�2 ��K+�����\ ��X�h, �Y$ށ�_�*���%�؎� �eR��� �o�/)�� 01���� ���b%�z �>�F�#��݀��rW�� �@ �)�� O^%�:;���� 1��4NB��u� ��J���; �ډ:��� ��xH�h� ���A ͻk ������ &�"Z·�@ �1����08�.K���p1���ld��͈- ���>E�F=����*� ~���e��� >'�^����}| ��4Z�� 2��S��� 
>ԋ3�7|W v��!��; Ĉ�W�ӵ� ��itF&�H� 1/�	2�Q��
�՚`�� P��(��o ��ɟ�p�h-F'1�{� xr�s �E�#	̢P�}@N�"U���W��p"׸� H���ZC��+Yʗw��k���ܦ�x�[W�%
@���隐� ���5�n\��=Ű��p�h�� ��)�6~� �-�g��	A'3�Pa����- �˂�6��/"�f��&`�Q �T!�:����gs� ��F�4����x��pr_��-`�� ��~��ݳ+ �_#��Y� ������@!� h9u)�,� 챵�Y��
 ��{%Zߖ��� ���չ��3�p�uQ^#G���m2��F��I.8 �K�� V[�ŝ"O�b�
�蛘� �Q\�+�,��`e���u��� �Z
��b)� ��_�W�%�u� ���$[i�'��h�Ȟ��}� �ڽ|���PQ�A�i[ ���V��3�� ��١y	�'�\Y; "���*�\&>�� �D��g����tRT���<=��o����)���_h�,2�	S�R@ ��vK0 q�"�:�~! JѬ���9>UL�	[�bA �$� 7����X. � ����� �'V��A���f����̂3_���!Z��n�  ���8J��'S@��%  ��L[�x! 6t�Z~�P �@���$ �5�?�09 �6%C*���! @5d��-�F#@����YtZ��@C1���*���q �!5���
+�b�ӰZԿFނdP ���ܞ2 =��1��r`u�/��F}�h�\�d �����.!�9�f�� �E� %�B�`MJ[��oY���&��*�~f �J�R��3 -.%1ځ�;��logxC��Y@�h8+��ǿ`�ן@M �[%��!]�S0{�b��ޕ �i��	�d `��
Q� �/K&�	� ��'�+����?8��C=���dc4W&[���>��ZǱC���\����d�؁�x��� ��wm)�Y 1�!� �J ^D<�Π�� :F����Y �0��A� o�R�V\�	x��"�;��� �[��<ٗ �G�ۀO��A��\, �e�	���R �y)% �q DI\Q1���&}�-�-��Ľ?
��B� /��w(�X�3v��N�0���h/ipYť֑���vp�{��8��А0� ��G�w�� ���* �i �_{��� p���|��x a����~-i �:�oJ�0f W
�Q�������'�_��� @�:�pL�?�1)�>` :n���O�t-|*V��R���v� �~�ب%:6���
�D��0P�4 ��-�� �6�+�\� �{j�X4�0�� U�:�2i���]� ��+�Q�c�Y������1
����� -�0P�*JZ�pm �Q/� ��z<��%��3�� ��|� L���J�V��P? �hI+_H(E��T 	^��U� Ȓ�-�n Xhvos�˷ �!�*1;�[���(���� ��sjA��������� �1��^Z� b$s�lBy� ��T�Q ?��&�'���I�ë 2�]A��\. �TS���(m��8ղ�@��A =�0���Q� /�.��͵�l��ؐ#��~� `/�5u� Pe'@~Q�$s[�/���� �j�8O�ޚ��� ]`Q_� �T��ciKo �u���f�>�Z��vQ�_xW ���������IC� y��Z� �R�ׇ4#a X@<�n������)	�Q2Ԇq�@����, � ��
�Y���=��-B�< E�-��V
�[@(���0�ӎ�г% U痧YKA�n�?�E����X +�"�_|�<O,��7��R𩉙~s�'��� ��:�YS����u(�BЖ ��=b�[�� )/�X����ַ��	�L'Ky3��>Aq��Z#�$�9�� �d �����C\[�@�< n@� 
��K�������� >��� *����^+��(��0�* _�5>9P ��՟%Xh��^�R�a)��Q� �l(G�� Z����� ��l]�臥 ��f�o � ���yZ�a @	�G���� ��|�/c3�w�B�`>EZ��� %��0�+t�;逖����9� ��h[Z �<��|A l�m�r{���(�q ڒb3׍�"�=���(� hq^��[Q��Xk �C���� <y�+����9�.� ��V �&î LX�Sb����&:	� V� ���XPG �!G�|� 	�p1��^� 
�R> ���PQ� ����X_L� )ӽ��� �ݸ4�1�0-wB8� L�D�% W�\w��<e��()�-�3'ŧX���u�w�@�2;A a��نbH� #���_� z�/�,�	�]X?4z�y.�@�2���
 UK�����C�О�!���:*�9V����b��'� ��H�{�l~2�0[w��4� XnE!�? ��1Y���rO㲩�Ў�7��3� �� 2J�/d~=��p����s ���g&��7��@��o}��8� �TȜ� �K��	S0ݟ)��ص� x�vN7�W< ��*�(p0��Le��,R�U g�LA�(�����t"��^i ��D����X�
8m$��`����o�1 �0�X�� g}�_�[�� �`���R� �8�%�x 	;�b��D\�o��Z�qx%n[�!��Wz���� �{�J;^ ��,��%0 @-?��>�w *�up�����Ր��x t׉(1�X9 �;� _��t�� ���N���O� �@H�T��� �9ނ��,X5�  >!»OBo�e�1�� n��JQ�� ������k�O����&! ؀�5N]����\O���?���u� k��4X�;�݂C������g'���G�K�~� ,&�x*��c��2���/ ����C�BhS[��`��w�P��J0}:�� �{�T����@e���D9�y ��
;��0[�ƨm��`k� ��!4*z$ \�|�@�� ��J�4�9�� 	0�!� Y�@�HJ-��l�Q��.S�� BX!�\�Z 8�>axhy `��oEu� �$�_�Fs}z/
��d�1��������|�[���/� H�q��p���᛽�ڐ 4/��*�9�1�(Y_E��+�;X ���� � P3�?�qOS�k'N�� 0�u�8aq�&�� ��{K�� e(�����
��� 	/�G ;t�V���Z�
�m��PU��`:�F������-l�x� ˽|�d�3� ��^\�D��;�Ȁ��`��[2֜s)���K ��%��o�$$��(Zp�=0D� L��s �\�^%=��P�� ���'vs� h���!� ��_�d�� SC�4���!,D�%p�r�( H������X�^0%�8��b��S�� ;9�E�� ��""}�8_ �Y�Q麅Z*���{��� j������W ��y��~���� ���fZ��  �s1�P� ��H��,��)�OY���*�F 2C��0�	�;@�� l���V��l������� ��R��zV<�%�;�ȋ� �T�	���Lb3U�2�`V�=f�����c�Z�C rQ̰�p�U �\h�qj� �/�����?*� ��N��3�9���2�,�R�"?1�
�=���� ��wP)�	 �W��T;� �K���h��g5��2R��B�� i��6\�� ��_���1r С{+:�9�=&S;��T'y pL/�G�Ybﰠ�R�ͣ	 �T���Q ����5�Z� � 	߀���Y�r� ���P�zL	� ��
|� �g;�ɉ� �1#��O4� �D�hȠez���P��q�XÙз��0N� �9��J@# �����°�9�K���J�ХF�� /���V�� <�J�pK��I� )�C����g~2�a��W  �1���p(��PhN ��Bd�ԛ �b�g��<� ���2�V{ ��	`c��uh�J9I�� i�vRT���Y���ר��P����p5 B��s-��?�ͨ�P^X��	DB߀��x ck~a]� �n�(�%�%8TV� �D��h �B#f�I�4+����� Ћ��Z5	1Ȁ�YW�� ����� }�C�7�x<#� �-�� �����Z��  T�hr�f-r�J�p��T U�򦉥������s���qv`U^�' ��i��9�2?��f��t`0� UM��Z �Y g�]�` �h9,�7��X�����|��t�ķ�}H0�N?��P�9�^eæ�p�`���� ��'AM�8 ��3�_ u���1<Ҝ$:�� �����-7$n� ��M~���c�T��q�� Z)���� ��r��W�� Z��*��[�� �7��,�t�� ZJ��Ł������"d9H7 =S2ͻ�Z$qD oA0��NW^��ߐ s�
����J ��z��q� M�T��di ��,�ˢ ��a�� ���P��Q��V �@\Y/N�J�@���-�*:v�X��ѕ� K!��Z��0  ���Q�" �f`-!�r_4��V�����( Q
���� ����A?� \(ʺ���v�a �n�ije��	Y�g�� �^���9�T��� ��KC�W�$��}S�/�#� � �D�<� I������ 
8n�����<�y P�OsF ���N�% �0|���Q ������;�:���L���[� �gU1Hɲ��B�G�)M�25�
]�s���b�'Sŉ������ V*���Z�z?�������Oui{� (C����Ē ��$�<�b�<u� �߼!��� ����� ��2
����N �ֈ��hŷB@U�YIZ�&���/�3�}@HEJ �t�j� L�^��d@ �+�PXA��( ���8=[� ����ص� � �f)� ����	�:[R*���a�0pV�A}o��s\$ �	�P-y �m��~1����@��ۿ "�l#��U� �0�,Mq�:����/��xZ�v�|�]�J���h {"�\ä�� F�m��	�.���2��@���`|���sV �.Z^} ��wR��?o�%�I���� Q��j�������w�	��I�M<�V�~u%���b ��E��aX� _��̯�M\����jl����(�� ɈJ��V� �P��n�� �S�:\rh�2�'�`	�� �_��~� 	�!AaX/�t^ ��RG$��dHb�s@/��� ��kJ;�� �xn�����z� �7�b�� (���*�p� w�y�����L0�!��0PQ.��J �3�Y���3 ������  �9(�X�mú��J��oż [1��ȋ�D� M��l ����C� �e��D\�.� 2��Pf�1�c0�Oػ}a��A[���� ���U%
ׇZg\��h<ik�L��b�� f�T�\ ��W-1�����Ot� ���W��b�#�2��B� �a��>'�Z �(�f� %�C�;$ ��73B4V X�g�>(�E @G����B Lu�J�Y� ӬbK�XHn�4��.*�>{( ��- ���N�V�iR� ����l� �������:�� 8��&�q x���(0� ����H9����X�5B�@�)�� ��
�! N��P?��/w{�fј^�U,; �#~3uUb�a��w��y�c��3��x �h"Vʋ�E ��Ǣ
 B��4q l�LA��j Ӝ���C��Q�bܥ�
� @5.u����Z�MG����	�'���VS4&0`�U��B</��a���Z?��^���̛	z��a�O��@���I��t '��Ac;� �QL��/R��1z�S*���w&>�
�[ ���1:�_9Ph'�@����	�� Bຐ ɘd�ڹIA 遌;�|Q���S���^�� �Eg���LY�He ���O�Ԡ �-��ț�: ɇ��U�' �u��ׂ-8�lہ�`@,
�v�%v2,���~� U�R�G%� C'�}c�� e�����F� ]1�P��w<��.��_`*�'! ˩	@U?Ł Znx/�&v� �%}��4�,. �X
8�� ��V�!:�(�g�2����F�P�pr�)���� [.��0� ��i/1>�D {��ʷ�3PP�� Z���0YLhb@f.v5˃� �K<�w2X �+�N0J��x�mـ�k����\�� S}"���C(� ��^'=5�a ���?,L
�	��m�(Ɇ%:�-�e�Q�f)j ���]p��~дD 1	��� ���:m��H�� �/��a��c�1��|���X��@�ô3iw��U�;�]�@��o �E�W0��K� )����[� ��{�6�rPt�Ğ� vX��cU�� �r��� �,��.8������ $�'^I�! �Y���oS ��_7����\@兾�J�� �
���h* }{�Z�师������ �h�3� [�0��Nu
� �a��:e��� H�89mv b��z�7 n#cKX�"8���ՋO�Y��c�6r���N �鈴� �3���&�� ҜK�; ��Xù%�/ D�	�QՊ �
�S��1� +�0E�J��Q��OKw@�@W�P��$� ���ۼ�� ���)��	 �Fv>��Z �"�=]�ʿ ��,���p�·�"���� l�)-��+H�:K� ��>�{� ����/��QZ���po1 p�0�n�$�� v��Y L�S��@� ������@*K���vp �����@_ )�S��� R�FȜ� ����0 ��%Y� SW���<.�~ �qӷV� Phe\b��g{���M�0�|L0��\ #�U"�� ��Z� S� M]j�R��,5�$�(�A0ҋ �Y�)�W��{�0���/��# �3`Un�� N��K��`P�X��.S	u����~�� ��ʹsjQ�&>����\2��4�� q駻�y' ���S����Z ���� �R�� f/! ���tz���[�����d�}g �^�K3W�-4AB�t�@��� 6���&�|u���ɺ� !����
T ]ƞС�d(QX3K�E��� "7Wz�� ��fr\	 (�h�U����- "��� �K�wO����m�H�h �+	߰��� �e�'w��� i���/%O��	��T�[� �ǹ�f0�� ������?Z��,`� 0�hw]%����V���([�H h!u ���B�Є +��Ŏq�\(>.� �����`8� @�wZ_�T	 �A����X��p ��S3�m� �D�غ1���@P�%����5!�
�!i��~� �r�1q]X 0 ����\� p���V�� )�^=zK� 6>�/�BY� ��Tɚ�z�?������U
 ٽM���78~��ԣ��Y`%��-� |�\�ӱ ��uV1��@}� Y]����32 �^鸢�� �_���T9=��c��j0ȵ��|w��k�����XR��a@EK~n�*u��m������N ����f2�I�vo*�`�� K���[��� W�#$��%��ęB����t�@�S/�ΐ <ڂ�V���t;�r�Nث�	� ր��c��W t@>��^}�2�B`����� �V��� ��v'�
�h ��D&u%HrRd��!��~>� ]$2ZAW i�G0�,�� 8D��� s/� ����#'� �Ak?,��
&[� 8����D@.�(��� ���O������Ā0g �"q�V��uB��\��Cs��pL�����%Q�̖ �����dy�4�#~��H`� Atn�0J �c3� ��%+��&`. ��$qo� B�3�U! �6�M�*�F���%($��;�k�j�K��3 ���Ѿ ����{<���]& ���X_�L q%�`�WT'�2��wZP`���R�l �Y)�Z ���HP_\ˠ��	�ku x?4F{$�̍|X���(L�s�d��Y ��i!.,�R�]g@��) �q���.� 47҈�Tº D��`�0 u1(&�T �����7PS�V$[^������q��.�5� ���!�J� Ƚ���-� f ���̗ ��Z�6��� �����'� �m[�-���z����aP��"H���Y�z��>�D $X���BI t�	�h, Nuf#%1E "�=	��l n����� �(�sx� $��&�U ����X9f�RB�Z} ش��E���p�<���
�N���� �KVQ�n�x ��D�`I�0���/�W w��jUe?��E .#�ѓ�Q
yt �)�(�h�t3 �_k�-��� l��
0&�������@S� M��Z0� z1
�����_?204Q�@.j� ��.��\ ~��P��0Z ��N��[c k��K,�	L�i�b 1��� �|��M"j0 2YX_E���� �fR�� � �Zt�$�^�Bhz�D�g7�} ����t��^��_Q��0u� U��j�Y�.�z" � �ro� ����hy�� �����ۀ9a� n�@�)�'�P� ����#�P�'���0.��@�G%��U��(�Wl�� �s �̈��Y� ���b�^} ��([�� V0�f<�M}'��=���`�)Ĥ �ًR}Xͳ 
{�ۧ�� �<$/B�� �!�&���� ���N`��X�.L���p��:�93�H��ȗBirY��J+��>��@1�����'<�-�wpf= [������d��AV����[ ��;: ��K ڕ�s@ޖw �ʒ��`�" ��,(���} ��0ɠ�� Q�>�!LF &���e��..��� �i�Z+� ���8��y#�J߳. -(�Z��+�&X�H�^U3ݽ������	� J����Qi R
�,o"�$xU���Ɓ��y�S2���R:(f �Pb\���p� ^#ٝ!��'� ��y�]� ��)/Չ:�[�{� �}F>�PΣ�������a����r�P1 ���G���2°���"u��7�� ����! ���z��&� �'}�Y%a��$x�� ������0b��@ ���LOb
� �ޭ��2�]��> E)�a�HSY h�s���*�[��^H�<mZ)��j r�i�o (۹��ȡ� ��W��K����i[C �/�� �.B���& ��;1u ���� �Y��m3E�q �I��� ��_0��Zzp܀�{ h�d�_b�xq����!������ ��r_1��4{tZ��2!O�`3� %/��� �}��qԶ; 9���k! ��o�=�gv�	%�y�U���@��� g���Z^{W����!�Q�P` s��/�� �0��	c�y�?=bO^p��m  �t�od n�Ȫ 5��KO$�L��$IE�w����{r +!Y�]7n ��b*��� �Z�S���<	�h�r'Ę>��1��[f� ]w$�����+�v��X �0�R� �� �	��JDuٽ!`����Y;M� �A�@t� ~�'��aOE ��&T.��1Aij9m�Ê���� :���J���zPU�[����턐X���$Ლ�<��l&0�3���t~���H�ڐL&@@�ӽ �R��5�����rZ�VYw	 h-
�O0ƠaX ���[��K��� ������=�,*����϶1{0��r��.� ��zk�� ~��0B�x|��s�!�ZV#� SҖ���.-�/�sؾ�d ,���%�?4��	��_����:���pH2�
� ��Z'�9 �{����� S����� �pKӿ�j�a�����&# �]���_�Lq�Cg�����8� �K��!ۿ� 
��Z��� ��f$�� 3��Sh8`�� Ưs:�c&�?w�/ОA�!� ��5e�_�`
t��-ܑJ���X 3��0(�_� �N��/�J�L����O �� u��nӠ�Y]����� ��h�
� ��A��l��Gb���	�L��΋��Z�0��*a_��0a� �v�^�E~U ؟ޛD�2� W�rhj�A}�;��u�N WF�(�� �U+���<�!�P����X ��Y�9. � �E��q� G����^[L�� I;�N����`вQ�~��=��Sj�s �0���bfV�;��\p� N]h_��#;���Mw���t��L��� ���X? [�˺1�"�	5�~� �{��`�0T���W� ��+s�)����h�爐 ���*�\% �nư������� ���qn �!6ȱ[A4 �|��U	� �Ffd(\*� 6�>Y"�?�˞È����������O��:n�s�W�>� ����� .j$ӻı�"����]����R�n��6��j� q�(�.ʗp P�����`� �1�d���2��=����'� �C���{� ��ŮϹ ��QAk: j��O��,�Ơ��Jră ��U��/ ��%��6� ,1�^Y`�	��&R����v�� ���P$b��/!���x�ty��� �(��2�sU \u{�/�� $[RYD1�� @�GH�s�h ��2M�&���� -Y�w }�8��B��,p� "��رq� 4���+|d� ������ ���I���z^ �6	��$1 =���'�M�?P��	�R�( �1ΐz���s. ������� ��׾`�Q (
���,�0ь����u _D���- �����̡:�>
+a���@��N���u ���h=J$�@)�Lˁ �F�?�� uB��$a� �z�!��� �d�֐�%�	\�{� �U�� (j�$r �P��
@��1��	 :�h�Ұ���|���.�� D�m�aQ� ���ч;�] Z���g,(X�x8����@H)�~ �����D� ����}�bA L�n�1�J_ ~K/�8j�� -U���>� ǘͰ���k ��M�C	�H�W J���xK��ʨ�8�5> yZz��� >�h����?��aӔ��������[	��π��<) �����N�4�/;�+�PX����!���� �0�^��`� ��cS�ʐ �3?@�#�� ����aU>�Vº���؁ҸJ�����j��� ��'���	 Ӌ+��� 8N�\`�� _Z���']� �&���:�ǀ4~���_;q� /�-�+� ĠRQ�W�a���F�&� v	 �� ?Z����[��Ü��0� !�+�h* ��j/����
������Y *ݕ��GDs �.���u	Ty&�f%���jAJ �1�@!������  '?�����ˋ�5V֮������� M_����4?�����.��m`�2���:��>,� ���4pv; �n��h&YQ�,����nA;��� �`43+� N[��	h}R|� #�1�?� ���E<�[ ��s�y��0����$�W�%| �ٻF� h�����^1�/�S���7��`�hZ�(� �k�BAم* ��1��j� ��k�e�K z)�L���>��~ /�;�^��?[ �U��1�E *Z���W ��Ƞ��_ �H�ʖ��KH�� YAj��e �#�(,�D ���-��j����X�K ��O|?hC�� �n��Q ҵ ��+��0��7\O� ��c�>��#ֻ�o�� *hPD�"=% �pk;��K�H[� ��s*u^� �
���6[X��f2 �a��P�V+ �\T�y�zt:�{ �D�!���� j#���r ͗_����l ��^��� �[W�>��n��_^w� �P=���h�bI��ȷ0� �Ƶ�J�^� kDzIr�5 ���ԄR M�sH(� 	-���� �D�^l���{� ��?���p��x��� ����g�\Ӹm�P�{`K�> �h�(�HA �z%x�Q|�`)���0 �_��X���9 	���^��] �g�����������	� �2�uLs�� jǠ��xX:	_U �����}��g�h���,��pu�; Q%0�_�@ ���^p��	-!�H �
&	W?F�9ځu�Q��!��;� oB���nY ��U	�:��g ���X]�wQ��k���"���� U��/�2<u�k tے�� ҋaX�_�� <��M#��?u��� '6�Iw�  ���� ,�G�KQ���jӬ���E]"ԡ����S� �A#0ރ����*=�?�� "|� �M
V�T�S�)�!m`?� $t�C�f��I� _�&#��[���vo�` V��@^ ��6�*� ���X�% Ѭ�����2�u�� �Uq�z DI	+ҹ�? ��'�o%5h\-ZA� �/�@�J_�� ���2v`�6p��@���� �g��!��~ �J8F��H�.W@8 �/Y���|< s��N� ���-c$D �����*!� "�?��'Y ��Bg�*��,	���dI� #H��-1 ��Q�3�T ��C������������ ��`�1����	�� �F.��8 R �-L�"�' `�Q#K��� I�*R告� �͓���;� �Q��]�ݰa ��O��|�-�ҍH�>p� �Lq��n�V �2�W�D�UQ`��=�l ��5�� Z��?Ē�x�����5A{+� {Q�p
� ��9�(^���o���_��G @��A� �kUN� (	�������޼������B �	vU�HT]��O_ �XKR� ���Z"	�Yx�yx�� ��K�$%��~ʦ����(� �K��Ջ�{y� �|@I��`�+���`~� �.��qC$ ���m��	���� ���� X,�Q側��� g�P!�1�bXs+�F%&� Ug
1c���6�� ��؊�_&��� ��hRw �'8��] H�3�	�� `q2B�S�p �AU�*�� ���)ѽ � �Z!��Q ̱>�m�_�1� �n��� ��?�J�0����� !�3�_� P*�h���R %f�ܨe}�/|��4j� DJq�dn�R�NE�b0�@��O �����N"���^w�V��
��Xhi ��{[��S���&� `eV� X{��<^�� yp�Mv� �Z���`d��g�ǰ���!� sL_�q�	 hA�U�k4�,ګ������?n� �h�YW�� �+�u�4�@�x�I�!����)� Ͳ��( �q/��vy�c �ߌ� �_��}� ?aR�z*̓�`W�ط@	� R#�81Ӑ	� � 
��Qr`�pƍ| >N���莲 �뷬��\g k�D�f���8 �u�w�������'�˦�^ ۔�U+�Q�w��.	E���C���= KD����\� �h�`:0~u��W� ������ '+�U����_ z���ؒ՗RJ�\� �	��L#��� ��@5[܃� f��ԸP ��,��U EǒO���I�.S_����%��`h�d��A>q����\� ы���� R�<�u�\���_�apK�렙3b�	(�-��2� *��@�%<�?� X�.�8 ��*I�"0�8ω����3��d�/���wp���] i	���@���e�(� 'h�_TR�� 9K�<u�0� ,�o��[W `h�Sg�K������
·�$&~L ��e�I̮ 1���J�A% �x����@�<8# �5���0�]�V y��\
!`3��b�Gh��� �4���a ���Lj�h$`�:�3[Ar�pxv�#�����O͐� �o����HH%��D'/�it�9 (�Q����# ����p;����`��v	��A`�>��k g��)K� vS���� [ �_�i��	8ݱX�g7���w� ��[��-� $zs<��	�t�j3@�!Y XW�o��J���=i+�j�4�� F�$��_� ����8�Y�$ 4�����U��Q]� �C�� ��KY��2k��D ��� �����@}! O�Ḡ
�U ��ث�P% )w�F����J? A�|l P�� uW�� �^L�f(���F.�����xR ��bq&� �9�Z�I
+ y�'�?�����x��T&�C��fP�Y;( �	X ��� W��í�#�� 8}Ѵ��=� �SY�-
^?@% ��P���� [0�W���=]3� �Q���[L}���a �C�4���8���3&	~� Y؆%�>�1 
��w���dQ�@����S "λ3�[�ﯝ�>��o�zK��	� 9�H� XO��$S*B� �^2R�:I5<_�X��=f�Sk�F����Hy�$�a�(�ń�Z���'�=֗s p�H�G�?��N�7]ϐQ�? (ʭX5%O ��`�h1L �ס��;f) �[H�	�~�z�!� @\� ���b鼍
Ir.��>�n�E�ua *h�e"/ �Ѫ@ڹ}� ���P��̀�k���� ��\!��<�	�R:̐�?& ǈN
�7� Z(��8� �� ڜI� x{ԃ��Z� ���en� �[
V���z� ���$Zs� Y7	�۫�t �0\@kh ʑ%�D)�� �|�(͝b�}ԔI�ӏ����C3�0�MPU�%�N'~�X�!�}�� V��Q+p�' eL0��W_�# Rhcv�����ʀ�<	��� \wz%��� �_����m�1ں�I -�82�?�<���q�+��;� ��)��n�t� ��[+��W� 1���	�3H��?G ���[1�XZ�`I�F�R8�h��St�\Q-uk޺M Z��5�
���ύ�	������@����1/ �!��P ǻ��b��Ҷ�����P��	�\��Q3 {�n}H�����!%��p���X|�P�� 
��.� I��Q��L  (�S�	 F���4_£������V/' ��h�s� �K�{�([ ��Z�h F0��˞!csf�.� �ӻ�� ��0���H@	�� � 邒��v� 
��?Z	+� h@�"Դ%�~����N�� a�"˄3��?0H� ��� ��AN�*��$� 6�)�-�? EU]B���  W*�� �ǚ���6 _��7"� �½�����r����p� �f�������  �U�yAYp:%1���Ԡ� ����� fQ���SP2ఓ�Z?��,&�lv�	l���� 9��A�����@�@R/(�1d jn���{|� ���]��� �a�Ц�7 ��w��0�s �>�Ǡ)�  р�bZ� SR�w�;E9 � ��b3�P #����CM �	�^���q.E�� o���p ��
P�:� ;�A,*�����	>�� �! վ;a�#�o� ��@&`[�!\���ݸ%� �Z=��� �Ep��� ����P x+ Q��/�V c%ID�a��U 4X��� Pp�<!��� �'J�2�d ג+`K��ɰ� ���
L2�:��b�y� �j�Kh(-{v ѫ��*�w5���&뱀u0� "��ț��� �pW����9��5 �!��G� �˦V��`o?Q��Yݤ%^c�� �{q� �o��� U�}S!ݻ ����3[��'=zG���V ���`1 ��RÐ��8�)�<�2�X� �H�8w�N� te����* ��k���� [��Y�H �q݀�&�t�Ь<�0�f��ΐ��|$}�� ��%�; ��ec�~� [��?�턦ȓ����Z^M�0ŗ��ә��� �4����:^/�O�
� �ZX�Q� ��0��3����gVPU*���h vͥ�:ʉ �Y*��栽 ^�6�� _����hX� +� ����?C��J4�Bel �N=�P�WY I�	����0
mXP�h�	���Y��L�� ����Z �3�N�~ ��g�� ����0� ��-����� ���`��$�X� ��h�2*�� ���% �C��G� ��/R�� �X6�� N� �����?�b������a� �Z.��!��}&���^�տ�BCZa���<����N�<�,������Zo �O:Å)�  ��]��� G�l6�"(߸ �+�_���b GSu�0�1 BA
� ��`[Z�@YR���8�����b ��3'�}80��l��	 �B-u��2 ŉ�^[�  ��P�Q ~#��ю� 1��F�w�i ��A�}�� =���e�Y ��s��3� J���F�\���׀X�P1Y#�>�kG V �é�̹�4�\ �p��' .!��UT&_������ ��`dʈ�E%�)
Gf��ܬ�2 �b�P�� /�M^�3* ��
#��� �[���rQ  �����A"��؋ 3�<T~'� ��u�xi�v ���GgH /wu#З2�� �v�A� �S,0�=��� �(�a���"vưr'k�ո��� @�9���L0�@����%U�0��Z�gE���	� ��%�hAs ��+��� `���X$�6���0iC �Z[X�����2 =�h�a*�J������@�"^��=�l �FPV�� w�`u��[Y.� ��� �� L9�'�	�_À�O`X Q��w� *� ��:IZ9�y��TL��������?���* �X+Z��	� ����Nt�4 Q*�!�����HJ"Ć���}i൞~���o �
�;-7� %Aݶ� ��������] |p�M@������,�p�+�� w
�GÉ >�W� �6M:�0�1�( �Y�V��� ��	��AP# /�+��\������@�Gr���N�~��� �� ݃+ .�P�p�� 3!4~ "� �I��@ ���	_ p� O[(��'h �kw�5�?���a�;�%�s Y	�]���\ �k<� P�	;�L|a��09���N�;!� .TL~��֣D���9�� �Bv�)�.�*� ?ްO��+[ ���K# ��?_�� 8�PZ1�d
°��&H�`Խ���5+�J�� �P ��:�,�k�(�N�@K�c$I��i����w�{v �h.y4b0 �U�t��j� `&�����3L\#Z���8��t� ��9;! eU�����% a/���?R������`̟:��o{�U��F� ���W$� �,p�/� �+ ޜ��� _\�X�<�3��J��Ԭ Ng���� Xo���"��u ��@��� �i��
�S� tne��^� �k>�~�<�s� J��`Ch�	�a�'-\���=!� �,"��c Vh�Oyx�� �0�ս�|�:�S �߻�: 0ځ��zV ��f	CF'^ �_2�S�� H-��`�B���1��
�_��=m;�>�f�2m� @	��)� ?v������X2� rV�ht� ���5������0��sq#A�h�0�5O ��+����hG&PšDq{O�$x������� _����c� \��h��t�´ٔ|`OG� '
�h�����8Nڠ�� ��[1��'-t�fN�0����I�$7p�X���,�� �4�|� H ��hd Ew�V�ֶ� La݈�%X��� ?��b�u �W��	x�t �ރ�&�f9~��"[��(���a����fh B�=?8�/��x�: ��F�� Ys�NƎ������O r��U��*��T�(�i�H ]e�Iu�� K��oh
�E���=y ����@�S�� E��cz<+`Iw ��KD���	�������V���]���� �#��b�C 5���7��f!�SK�0h �����[�R5r���p�K�c�!����0	�w?�}�� )��XH~�� Pc�q<� ��b���H=LzL��9��
� �u|��� �U"���(���g	��* ؼi5
\p>Y�ھc���j ����(�S �dt$��>^��� E_�ǌ;�kȕ g���rr 4@�1�Z� ��A!� � �{$�*�U +�	�wCH��!=��ؕ:�� �J���#� �	 C�K�P �o�7�� �!�(�O�:�C	�h��cf��yB�S]������ ���W�� �LR\� �0w � �&�O��bx7 ���hVI�� L���]� @<�; �����Y �W	ٿ�� ��郏�� ?
=/�*� �Zd���)P ��$��
  ��j%ג ���ز1(��[���� @���V�G��`� fx����4_��[U�'���N^�w�����ܲ��x�г� =� %(����>)�K⌓�5^�d��
  �P�4]�D��	��eI���  �:�zS1+2r�uǬ%��H�� Z����* ��϶3�ʍ �ըA<�e�;� S���3�Ϟ0�>xC}Q� ܦi|�� �/�W�� +�>�3��: �RG'6�uh�%����}�A�Y`nP ��#z�٣@ 1�N��V��@kI��v�^"����L�a@��@��, � Z0�^h�% R'霠/b �|���S� ��(41 Ћ.2�S��L �@5�O� ��`$͈~ް� ��8ߏIEiV@�tSB'˺)5_��� Z1���k ,� �i��u��� UW�J��� ?;��,ù�.ǰB��2u Nw��,�VR 6$�?)MoX�� .�7��t�%��W��J��n 0N$��M�X�- 3<�ܩt�_��8E��� �x-v� �4�Q��3�] 'pd�� �?�
\� ����،Z _���$'Qg�tY ��K�� �¾U���ݖ�������p�?��y��ׅ�� i��.��?� X$aR�x'�@ 1��V9 �k�#����Z�� ����j b���wpF��= �$��%u����P���cj� ����kE�ߎG�� }y]%8���"9����V���� ��s\! H��O�v�� �mw��5{ b�&2RF(�ī���@��PU � ��#�}J �Z�� \h'bv���`;y> ����Y�X ��˓!�� %A�RQ"+ň�Ǆ�� (	�!��HXn��ZL�����w�X:&} WYVOK�T. ����2pM�^ ���[-(��8N�h ���[������\WU#q�Ł�����\i �M�����r� @��K2�W M�e��| ��/Q.撯 ̕�'�z�4 #֗H��� @0�f^���Q��(�c��Y� +w ��,E �n��;Ҙ�� &)�[� w�����/w��1���3� iYO���9tA;�� u�)#�\ �w�c}��k���<@�:� ӽ9oW٬> SY	(Ѐ^�3p���w���`Y?�	� �tǁ��e, _
�∕f �2՝i` [�����8�2I@�a��� ��ִ�WL� ����j��'�� 2���+�� ��Pp���_�-�?��	 �� J`r�|g lW��3� �2���yI ]���!u���0�X ���y�/��� \x�K	��1��WfQ� #0[�hyYL�? �r��ow� ����j;�z- K�E�\}�:�4�} i�vV�S�~� ���P� �k�C� ��@�� �m����}� S~d6P	�.��D��؀+ӗ ����
3��� �*���g�`h1��`'�f ����UO��X�O ]�[G��K� l���ܻ~_e�S�(֠�5 ����H�����U���@�ո& �-i�wH>!��Pq�/��%	��
���>�� �	~��a�# �4�s�:� cQ�'��j�]�@I��7�@L-�5 �^�&�.� �8`i�?�H %2�h�ov�� ��lՄ�G �:�΃/�L�6�%0(S9�x<ӿ�7/�K�� �3*�� &��n�VZ󬶀t���'[S��h� "DP��V 4�10�m� k�S(�>� ��* �P��_ '���Y�p>V�w B�#�%c6����u�D��������� r+û� T@��%6c�>�b�^������[ !�����0x� ВR��� j v��T�@������� C��h�v�X�g ����KU	��Ω��6.8����;�c �YϹ[<�o)��Pں�� �/R4L"sb܋ \���ޕ ����Vl;�+� 
���1��z��0�Z��U!�>
��ގ��Ay�]��!��u�'� � �Z\��B.ߐ�2輇< k�fJ��,r� �����! �P�3A@B� (���n�Ƞ�1�>*���~7ЅƼ� �����P���5��!F����L� D�����p�3� ��2?p�_p��
e]���p�}H�uy���^���*U �	�S �_q X�vo���X�������7�,�?��8R���N;����)0� �|�%h�O ���E~� Da��Tة`z�L�ᤰ�M�oN�Ŧ�7��� ���.[�S9���^�-��\�� ��!/�0= kH�A(LO��� 	�b#Ve��Z�� �a� �k���מ �����w;V�K���6��w�wr��[�Ɖ�V���X��c��W]�P_mb� �a�ܹ��� G!��b��s��$�N �Z��P �Xɼ��� ��3�k��� ��f�Q�� hL,��-� #��T�<�� dOU�]�h�LTHK_��|\�� �� :#�1 �wҟL�:]|��K���.ZhT _l`���E���d yz
 ��0��`�v'�d^��=�� �L\+O` �d�Y�� l������ ���$�~���`T����@��o����NVH�1d�������3���S�� ź-���P<T选��^i��)е :��O��$�E/����C�)8�� 3�_���L�� ��D��X� E��A�� ��N���� S��r��=@ [������������+����p�[Z�p��!<�, X��<&. P�)�s �-��O�� ���S,Xh Ff��$/�" ��%�;���D����� �� �+�C�  )X@
(׍ ��L�Y�j��fz��ǯ����b���`��W��� �7��)!��|���p�r> �z�	V] �L�Q6i�� �h@x�� ���XI8�	�u 0��2���o h.���ܘ |	c�ɴ��X���o$�G �;�K�J~�ׂ�H��� @&-��5% ����K��W���G�R�� oے)�Z3�W@ 6N�� ����!�/Y[���~�^� Z��1�`�y �����GZEN����H+�=XW �*���bP�"�\���i]0� RJ��Q!�}f,�˵> ����� &ڕ� �i�-Y$�Q� �4�o�9`�����[稚 ���$�K��� �����Ao0 n��*�3�b�͋d
�����s� 'ha	��ۛ(�!ꥸ1�~���S��k���qV���`*K �tvS���hdL�'���@-� ZN�.B� ����ٟ %	��(M ���� q�� !�s�����0ވ�S �#s�L� M��0��G�� �.!R_�[ ���P#θ \7��5 �>��ð� ���$g�)�@�H��� �=!	�*� I4T��A2=�"��gڱ�� z�ā��� !�(�r�9���6lC�
�Y@���.[P�;��u� %.�W�,_��]�  ��y�
�� ��Ya��'��c��Jj� �>-��!� �%��v�'V�I��hP^�? yK�&�d��b-X'�n��� ���.( *��D����Ӻ�E�|�V ��W������ȋ(�玷� P�ʤ %*��Ja��(�u� .>S��w� 襷���\1���-��[O ��c�8^$���_9� (�h�[	0 �"�)ը�� �W2�_|>�B�@�@�z� m���^�Ñ��� ��܀��i�4a��{� �0 �_��%Ͱ��ۂ�ؔ!�QǮϟ�����	� �]�������L ���QUV� �PRM����9b��}	!�"ڏ�� ��W�ҿ	i(m��u��  �?AZ�����e-'�p��ˡZ �������締Y� K������.%n �
G뇱 �4}�<�'�r�& �X�W ��6��:� !0>�@�H Z%h��� ���ƯFg ��|�{�_��i
w�e�z���:  ܬ|"h� 8��*���`���ɚ���p��?aȮ� "�_��H �&��C>fՀ���%k �TH�����C}t�x�p��S Dj� ��\	$�]>yS#�
�>@��P�Q �����1 ��Y�d ���|���L �I�xv��r� K)����h k2@��ߕ ��O����?�d %q� >&�_�� ��O�Tg�p  �h�?���"�����Q� ɧ#+��Z�b~E������ ,���{=!� �:�	sU� ������} �C���	 ��`��9*�@���!� �X��m
�ly ��xU- ����{ �H 5��)�QX�$ Ƒ	��"K�Z��x�b�\�.��sF�w�j�� ��,�O� ���1E����@_�Zr� hBKo��=X%�[�n� Vn�U _%
��	N �� ���ɳR�5@	Q��F �Ȝ,y&�r �sV?���1��\[��`��^	 ��]�>��� �D)�F Su��� (-�W0y�	),�P߀#n�� ��R��X,$��%�y�D����N'`� 0���L)5 ��=+����  n�U�H� ��eŢ�	�)@ ����q �����A X��{���\% B�N��&�Ż��n`����|
��8 �Ւ�t�Z� )�Q��0�q�~[Y�� ({��# �>`/��- '}���0� ^�ʰ[;�Z XL�ƅ�y@��[��lR���S� b�&wY� *�d�)��XK�� S�x���%3��o�p��`@e�=2��V ��Q����� �A(�I�ä4<ap�� 1�Dـg�:����@���(�� dbLE¼_� ���]ޱX+�s��k��#�t \,d�J ѫ�0�t�p ʥ Z��. ��XU!ҽ@ �v
K��� ъ�6rZP��^���S<�J ��_@-��2 ��F� ���&�3 8'��4w�X�`ǅ��� �*�����:�ۀ^��e9�h`0��M� ���1<� 3$q�- ���W�S�v ��8~��4M �
���� �^�d���v` �pB3�� X�]�Aj�� �oH�w�e�͔�����&�4'�� �_ ��&?ْ�������_ OS��W�� [!ŧfЋ 9�`���pS~���	�U ݄uC����� ��dQeW�4 ����t�\�� w�h/z di��\� ��.)T�g �"1�h�H�~�@G�! sn�[Rϥ"t�U^;���� ����%���8�+ �~�� ��SJ��� h�DW��R{�t8���� ����<����)Á�� ���h�����/�`����*Wå��S)ͻ۳z�ѕb�`m�[,3��v ���: ����Wyx�?]f����{!� K�P����A D�z�)�%+�ۇ
s+�lZ��< ���ц$� 8����\��(V�pR�.� Oy��[vk� NA�?��*��ߐ�3ܚ5���V����> �c����;«0ߡs��x� �h^�Jݷ � ��T"v�0�X�I���@�Y� %�O}��$� ��AXw"��Yu��@�hc+�P��\�����f�[���p��~-Ⴠ~b�T[�+�.��jݘ0X`�� "��vO�;�3� ��9j��� áE���8}��y*�`[r�9&_	;�����h��
 �A�_I �Vl,j��o{��A�R�f�*ؘf �N=�g� @��4�xG P�	��7 ���h�J/��p��� ��郗� ,J(�%XQ ~4'8̗ T:g����bRP칾F 25��/G�q `H�Y��ظ� ���#�8gt� �����&0� �V�'|3fX�-����xI�� ���[2�� !���a� �<�Zh� ;����~� $ۘ���P|`�R��S� 3�T0�`V ~�-��H� ���b�J҈�S�� ^g 	���WE( �!?�� )�^ʖ��1:������j? ���,z%Q� �@EZ��yU� �"f	�V ����x/� y�dZ^#�rE����	�� +
��AM� ����@���Iu�*	� ��\o��B��:�ډ�@��W� Z�E�2���(�]*�Q�0s� �0��F�U�X6��Z%�Sx ��f-H�  Ӣ��	�� �;��T2^�!��N�`�D�� �Eu>�9w� *l	�S7�^�3rȤ$ b?�	+��z~����qK� *������]~�^طA�x/��`鲙����ɸ���a�h�e<� ��wԜQ9�W|ՀӾtP ��H�'j ߘiͅ�t�������0�3���� Xh�q˝JW�T�`Af!�f��d�t��0<��(�́�5�� p6�	�%P�LXp���� 
yE�p.�\9|�ֲ��7� �Ƹ08�Z 3�����{����"�Þp}!>h:H;L� -<�VG�Ʌ_�:��mP�� ,R�1�\�$�;��-`���T,�|2Ӂ �:Z3y%��\L.3 ���L� x��t�� ��#Z/� h���!�yy�L�| v���a
 2ۋy��� �c��|/�%h�	�b�^�I���=��( ��_-�. �b��N���Y� �QX[�����? ���Vt],���1`5z�{��txw�@3[ ZY\���* ��0NȽ���:k�y#ﾊ�M��� u
�7�hd S/sɥ���gC$ ��l|� �I 8�Z	 ��5��� �*�@}�f �K�H�� h*� �X�i �����8D���[`�Z�e$ 2����,��1 �w�A��V +���T���^�� ]�Ä$�/	�� ���И� ������ Y���dp�$ Fa��*۾k  }�^�/���g1���O���@ �ha�K" y��C����|� Mds��n�p �!л;^*� ���:�x �+���� V�0�eI�X �qY����9`�m ���D���� \:�;�� �$��^B��	�W(��{��H{aY@�ԃh# x\	�z�r�����Dɸx ���U[]5��Tc䱀�����te�]������#����8�� �X0Q�/*�Ev����� Y�5�{�y� �z�}�a ��
�GH~e ^��,C8A� ��c0W�_�����<�p�������!Q�& 7|�, �� �2���e��PE�*�9+����FW� gTa�G\h��	�RA���� ~.�g�=b ���O��	H�D!�3�(`0�%��V� {�� �\U�%��W��S���yx� #($���å �
����?����LO���1���o��e@ K�rO^�% �D)ߎ��LQ@�	[����]��,�z�u� Wv[�:̓ X�'��e� 	`+�m�.f=S���� ��Ċ��O �n8�Q1a 6�|@��rw:Ұ�e��4� D�(��)@P����z� ���& ���ո� ���'�����O(�S0����d������ U��1 sx )��]�F#���c�<" ��H��@ � ����V�'R�\ty�K� Gk����X!�]�`�S� �o��Ŕ�>�J��`�˒|� y�B��=J Q��U��&<�;&4�TYH�)1mu� B�Z�϶ ��;��<�����] ���3�_!�`;,��F�^�`�� 
�Q���> ���� ���?Ȅ�� ��J��-�B�0� ½��w��	Q� U�h���3NӀ'�[- eK�!|��_���`4.� ��\bC ������!�T+�`�w y�7Q`� �<���� ?#�(�u��p]��صȢ +�&����P��T�l) ��G�� FB-�^%� *�WHM��I K�'�����>��g����� 	���fb�� (Е�p�d Ƶ�Ph렫�B �+�t�b�w����� \;�D�cm� �'��$���N����t+�1Xˍ�u���NKIt�%v A�@�_�J�(a�j���8�� ����d�Xap�06 ��_(��T��t]�m`Y1K�(�w� �N�ae�3 ��KV�۽f �&��^��th�'(�����}��@�Kw���H���N;���u?Y	�[ِU2������J ���q߱� �j��2�<-S�l�Դ p�/���� @�	(%�U\��q��vsA�k��s`�.OY�c �ڗ�MZ[�qnBNw������ ^���H-b �ĥ�ǫ	* +�!N�{�����䡁���)A>�c ����%Jp|� �O�Z9���p 2��z��;�h 4��[��-&� �噘� "Ƚq@�� �P��鿋 I�h\�%e X��q�� X9� ����2�. ��[S�:m��40��1{3 `N���ɇ ���G���/!�� ��{ ���-p��g %	�r� @X ���Q�1o *3(�� %u��[��s��G	Z�L��o �8SN��+���	I�� �?�hb=޴�8�-R�Q����+P�q�� V�/"Ѐ�n��S��Ћ�xԫ �Hk�h' �L���1���� _�A�}�;0�Z�w@k��c/��y��� �>5� 4�ԝ�4<���8��: �h˴2��8l�����PI��C h����[7D��3.�g)`y/� ��`��Q�O+�d.��<�Z�A�� ��4�$8��� �~-|o� )�'6=�N� �SHp^� ��-T��`Qҹ����6k�r��g�@֚S��O��E0,� �̺��$��H~!����@�U%�8���7}00
�?�ڀ{��Tz^� �yW��	�n~%1���a �����ޢ�u׃ſ��b�� {��v�Z� Bкc|K<;�U��ܼ�X� ���K��� _|��a� qD~������� ��
W��� ��M��X<�8� d�R$�s Uf)Ţq��Y�[�'x��TԠ� �Z2������J�)�9�X�x�j_��F6�P� �}�EW	C� 1�h<+ �`��|��� s��c2�F�	�1g��K[��/z�xd�� +�Rں?~ ā�*�1�Z�s �4��� Q/�|U"�� ����j��	�Q��ZK (�&�'VRL ]ʸm�}� `��P�0���,v����Z)JHw/ �zQ����o��[�-0��X�� ���_��y��e�?�	��X]A#+���W@%[Y�P-4�s Ƹ?!�I ��2��`w 8��\��'�$�V?������� �ev԰�T1 ���it4I ����;�3 L	O��w����b���p��� ���x�	�Q�c ��7�yk �2��*L$=)�+b ���zx:����H��ؠ\�� ���7 ����~�DPp�* _������ {���Ph K�d���`	�����J�n.%K�N{<�����@k�Gu� ���+%�0 �O)�HA?�
jp��h1�r �No�d�)��$J��vs �����:�" �	zV�l�� �P��0�u&|ˠ&� ��ر�c �]��x�g��X���0���K?�' ���� �"��<�ּS��U$l �����k��2_�q� �)���� ��C�d n-�>�5�/l��?���E�`��Ǡ ���#.فB� ���0 ƻS��%�i�n��MR"�33꺜@ـ����Mc�]��Q� ű���(���}YC� �[�f2 p�~�xR����0ػj�� c^�h�� ��8�[�C��@|���i �t����z� �V���[0� pX^*�F�]� -�T�|' (�YXh �Z> ���+�x>�3v9�u���%����.Rն�k�����-?����5ظ^ �j��n<�� ���1�R��-���+�����'��P�0��Q��������s ���u��V W0YG��h���-�� ��ӥD%�R	&�肰���������0.��!H�'s<[� o�\�� ��P?�s>�1�Z xW�Z�������LX1 J��*���b ��	�E�� ��r{��0�]����nh��S��2� �6˘!� �8
�ȿQ��Ք��`lN �b��3JV ��%�� ���K����R ���B�ն>�v��W���j� @��Mp4�e!�$�81 �����l�p �@��gX�C; ���A ���W���� �`��_��'vBZ��\������>(� �Bӂ����t��f	[b�T �&�8 /Z�'�u �:�@#� ��b�0 ��,(��Z���V`���& r�>��[���� ���] y�}fh�R �'�9t��� S
�Tph�� Cj�-f� W*���"��ch�b�A�B�q�|�$PEz��	t��@��� ";�Af�װ$ X����δ�*����S?���W��2 �$��] VfI��@u� ���	��^1 �5j#�� 2"ɇ��hF��OKøvA ���� V;R�O{��G�
u@�� }i������� �&+����v� o�M���TUj_i\;���. �z�h��P �ATXl�� ���3��?Py� �X����*�G
�Y�Q�3�鷨� �K��-�̀R���X� ����	��$����� �!�`贿 �6����^� N����_ ŝ���t �̶�bZ~/Y��'|a ���Vi�?$����*t��� ��,_ ^�D��Z��w	���d=�`Ó ��5G-��� :��,h� ^&�y��#�� �P��.4������	�� Y��mQVK��\` �_�+%�| �R�">�����f�-{\2 ��9v�U�SF&��]\�� ���>9N���S ɣB6�rE�'��i�Rw񷌃@nS� �
���? M���]� yd���	�,�1� �>S4�;�.�J �{�'�6��:���8Ep�|� �_����R��y���j �w�+͈�! ���P �Q� ~4K����|�% �8�VD ��R�-���A sQ�Ň�"�Hk0 \x�DiW'1����=s���~� 
�-�+z���PE at��k� dF#�=	��  
���<��R �K1Cݠtd�ܶ��_� �(N���8 oOv�D�P� J����f ��F/�~�Y�zB�9���xe	�p ��cd�L[
���0�	]�_��{�O����� 0��9��J� �>��(�� skM"�,8U J���4 ���7j�������`�R �)���� ��ʉ�N��^�����h ��3��� l-�M���0 @�P�� ������+�3q�Q`Mh Fx�/��� �!�+�.� �i v ì��Ɋ�� $m͑6H8�
j 5���) �\�ׄ�3 ~��>�D����Ÿu�n�h_ ��K�	A�� L�)���(� �a�0��kAC���V� پ����H 	^:�΃] �����z. �D��I��^ ��&4�ft����?߫ q���	,"� �_,����Y[�9 ��4BV�ʾ� ����F �L��I� �7 M�i=�8V� 0�RP��l����� %rOt`�� ��~Dj� Ѥ�/^� � ��m=� �x�Gc���͌�N �P2��� a���w3� ;��k&m0s��h\_E�!Ҁi�"뤥 ���� h2�x71�A &W�$3�X��{ߤ�;�� tU:�s�A� �/bx��{Y �n��4���[�R@�p�� ��#߁��P����Q)�˝ DаF��($O͉ơ��W "�S��� R��`E(�!�Ӯ��Cz�|\ ��e��t� �nO��� ~2G�c}�4�`�	�_T�T�W`d��� k�4�p`�w���� ��m���0� ���#. �k�fS %� �P�s�=� <��'�:eB$�gla�5� ��1��� �>��_$� ���z���`R���M�h�_@�UB�����	���Ŏ ���^�Z� O�pP�!J ٯ0G�݋a��N�~��I��Z B�A���>
	 �1۸ � [;0�����Y�@�S�
HAu5�\`	P���I��.� �,�%��rF }�Q �"�$C��J�_)'o�����ݰ@��c��SW��v�@�c��p���l� ��� 6���� ��^�.�f{; ��'��R�,y� � ��^�A-��/�'��h9��� RT���o ��UY���~ӍK�uq@`T� -��W��J êɺ:�)>Z�LB �Ű]RX�a K��@ �F��9� W_�΄ ���,!H 	F�
 ��3��W� �6��J/)qk ���uE�� �^g��k}��)����j��w�	`�I�^t� 𠉋L���.A9i��w��� ;�ӂ� hro�U��> ��i��B�� ���� 2����L�!r&|�	�b�#� 1C
�� X2�}��R� J�_|� ���!�Yh �-ָRuDw	1� "�6gSK�� ��!�X[ ��W(ﾉI�K�6Z`�~p� [1�V(�5� ;-�E���8�� u�	����O�~��%�� g�]��$����π��	 �h>[,� 2�f:�W��~ �Ђ���2�"���{R �&� � _Z��6�� �ڼ=@��� 4��� ���,�h'� -7�� �����V������^2f`��6�:h �S��WA�	 ��3K"�� P��>�8� ]L� 3(_Y!�K ����h %��ՊE����^�����L ���0�h ��1�3�. ����n���2�d l0��r��^� ş"�� ���銚@ XY�$2Ұ=�ta�@��S/s� ��o[	�� 0�n7��8"^���Y�����w��@������] �lRU$�p�� 2�=�%fr�̀�abX(BJ�v16��*� ����� 	ռLC��z� �)�Ɉ ]W�[�E$ 9-񕬩,�Y�a��� K��A�=E%���5�Ԇ�Q���d�k)" +!�a�7�� �w�9.؀�[��� ����(J^����yK���& �q'��"� �{hC`t� p��M� lK=U���1 ���JO��4���=k�� W�.�Iܧ F���	�] ���Y� ,�P�C�Q� �:1mT�b���9�`r-� �	B��lԺ�Z� �6PUVH��m��j2�H�@$�� �q�; �)�w��� k�W�JX� M���>z �ˁH����� #��'�	  Q_mF���u(� {�Ko��Z���^���'$�� �#���h H��%+��*)�	�j�@���� U(Ž`� �/�]fL�	! �� Ĉ�I�Q 0��;�1�� n��4�� "X�D�C���ܗ�ȸ�K� ����0��&��^��p��� )��~u �P|�i	-� T��`nN �;@��s�΂*ŉ���j�N'�W�0��Lg �+����^���S�܉� ��qfb� ������� ��]��':R��\��h�J 
�a"�� B�P��L���h������Ap u����?߀+��!-z��	��~�F �/�`�c��`*��^��n�2`9�j�
����R�#�@����~-T?�S�ݓ���@#�[��1  $(u��� �
�@4:q<��S �m Q��`6�N ܒ��� ���_�z� ��3`�� ���M(j� �ނP�c�B��, �~�b�x T���.�#;���4�5� ��9_����~� �����5�9DZ�؃�I@�o�� �E$1�>~� ���/M	� n�����\�v �����nyV�� �$	�Կ,4+Y? 邕�j��A@1�	y�@�1�K� :U�t�Vy!뵖�п�M��Ft�rJ� �*�)K�:� 1��(}5# ������` �.���A_ ��I���vw� ����� �U�
YS���)�o�Iv�|=�n���~*��~� S��CU^T���0� ̓��1n� U��.�_�~���ty�`9Q� ��� �^��q�Z������ ;ge�h�V��NG�$b�� ����.|0	9��S��K� �oE���Q��~T~� +Y�S\����!���W��dj JUk��p�H"����� ���s�A���{X b��FWӽ	 #�H�3Β'}j8:���y�0m��[Ȱ�
�Z���7�& S��! L;<K�e��c�px����M7KvW	�u�-��@Q"b ��%
]	�p/,P�_�=���Y 
��]z�\� �'��+�[ S�����XI��V �D���	 �J��_g% pe�|,l(՝���@�7� \#�G�U3��  =MT�q�% �c
[Y���4��fQ�рr�D;?��� �	��� ��Q
Թ$�#oi�?����-6 ��8uY�B}��@��Z��I[�����h� vt�x@W�$ G,	�]�� B�8�<X�������ѐ�ck�X�h� p|�Z �$p�:��I�h���`m0 ��!�-� ^�ZS�̻/ �?� AP	 ��Mwx, �&(~[� �)�}W���g�x �S�ZI�|� a����`�\t���Hr �7��5Z^݅ 
���N�������ٖ��C@Vо��  �SϹ�����X����\P� Ô��G� �+_�Ѧ�B �y�=(� R)��� �ԙ§��� �]i-��b� :�Ef��� 4�UG	� Cg&�(3� X1��/�%� cP#����T���6Lt�� `�
��� � �*Rf�L�7 �ewa��H"} ����4�� �68�&Ao ��l��%t��Ӏ@��4|�$z� TL�3�Uƫ �h�dP �N����Q� :��S���^ ��2�_��� ��P�/To 	<·a� +�����x Z�LG�#{H� �|�P��!��ћ�13����@"@�� �[,޿!� .�~q��1$�o� �?k5 ^�Q>mT�� 2�����t� ,0�OV� 
���� �'�ݷ���H��̝(B·`Fh ���{�J1Y�j@6V�d %�B!��+�n���g_^? `�"��%� A�1=�	h� !T½'<u� s�Eo
X� 1��^��d�M�l ���h1��,*�{A�Q��!���� ���} T�Hi��K��*� j7a\5 �>����V� 	��2�`����������=���S�pg��D����� >����z�s ��w픖��p:��� 3�� ���֐V`�.�� ����0h�ڜ_g���� D=�K�!$�� ��wy� ���l�R1 ݺLϒZ�� �_�u�9� 0
�%ݹ�� ���GI�� ��\�6BZ3Jů����W ��^A��3t ��N6��pO Ȫ2�E��l �5���~K�� ݀���]3O �Q��J�'P
�K<� �ܻg<�}P� !H�jw�ô�� ���K��ً)� Y�{%=�� &�p��xy� M�L5E� �o�����1 8�]0� ؐ� `�e�d��;ܣ��P^Q%N�iD �Gf��,#��l"�a@�LH� �[�^�*o@�x�0�� ��,`$���` �x�� < �ڋ0 �Y(�h��xW& KMD�� �
�0��-��. ��8�O� �P�h:S��E8������+s`�B�� �u�`���r -~�3�OZ( ��@[��'j���3������*k� ��#��dT����	�f��@�~�Y ֍��x ���t]wHq� ��+Lr��[?�	� ��BDZ`.  ���M�^� 0�����6;�ހ;�٤C��\�� �d��� ���
vIڹ G<��pyj W.�%�g ��9Ɛ� o�{�K؇�2������d���<'�w��\?��� �%�7�PՀ ���C�U� �WIp��� �!�>�5H&V�� y����� �����@ �2Z��[ ���S�%��@3�.f�d&�B�t�U��4�L�>�zK�aH� ��!��@l�\�h 4�V�Z7�|W2*�����ܰ�H@|`l�4 ^R��?�>�(��+F����W>�� �~`z0� h��{�(?�r3 »_A�V �'�Y�1 ����J� �B�W��Rm8�(�?�� ������8�,%M,��KR�U��bI�폾O���@�1! �3[��π(�a�Pıwo�Wְۉ�Ȝ��oP��/�^&�2V)O���}n����r2	���  Z9�� v_���\� ���@������ eh-�N�4� �D�O����7�B� v�ZWt��|�,�7�����w�� ��? ʈ�� *m/X�% {ӄ!>$%���@�O� 	�e��^\ �,5ǯ���|������� ;r��N����  ���U�Ȱ$ ���%S>ٗ /����5 ��u�(!���H�,�:� ��Ȭ��w	��$�Ց�� )�o��T��c{`��M@@iVJ 2X��z5�" H%�U�W�8���5Y�D
%���C�H� �\Ro_�r�Z�� /� 6+�� ;���阻�v������D����!h��:�ĸz��>�@;� 5a&�.U� �<~IO+�b����]�H?� ���0�� ����^>�L z�ɐ�$ۖ��n�2 2� ��<�fR ��ͷ )*b�V
��i��ִX`[�0����%�+�:,'U����Ť�y_��ω�� Y^&1�QB�|@ ��gbq�P�ai��[j	 � �"胂w #��q�X��,��ḧ́�0�TfQ�OT� �\��� ٱ܇��Y�~ �V�a��� ;�KNY� H�w/WQ_��V#���}� �D��@�� �`����� r�I�Pױ��z�K2�&}~� '�V��Ip= Z�����J��2��� ��u`�G���ܘ�$�+ �߇O���p) ��"�P�� -z����r�H)y^m���(��S� �R!ź n%�^Z)	� ��tX�:�y0 j;��	<*��� ���<Q���{e��߄�<V �D�-�P 1�H�?_ �	ZӪa���A�2 ��`l ���	_�k��-��~ @"������7�v_~N �vR�m��1��@=�@�( ����Y j�!	Q�� �@+��/3 �2�\0N ���i�D{���~3	�
q|��� r�1ڷ*Q+��$|� �-{%�8��\��*�� ��E�݂T[\7�3@i'��L h�N;�K� ɢ`��M�b\%~0��tޘ3�R�D�*�N�drl�f � �V����h�� �Xſf<�4 [`|�� ����0 �T�<&[��a �'�t��nd���i���#j��l�\騪O� ��4��ʚ ���A���� ,.OT�#�������E) �Mz�H� ]Y%2���L ��	�$�^p�  ��,� o!X*� ����[ z��ё�� xo��D� $�M�|�}U�p������� �S�j��� �n��� Wqp�^F�4w����l�;�� �E(�a� ��~̘`
,��6���- �� 4�$��~�!��	��@Ѐ� BhK��>����;	xpH�3~X �o@���� ���F
ߤ�� Q"�vU �;/[��� ����R����3 [VP θQ<� �I`#��u ��
Q���9~2��jI���Ab`@��L �Һ�}�LCXR ��U�F���]}�0m[ ��p��.�b *����/7 	p_�=Bq��zK AI��F�l ��µ �-�@x ߊ
�������u0�so[ �S���
	�1�߀:���3� �*W��ǿP�� ]���pT�J H�w$k�� ��Y�j @T�%uĆ� &�X2��v ��m ��':�n��ޒ�B�r : �|��Ts 1�\h�e~ ���0���W���Y~(�6H���<�$% �����½�LX`�bVZ�=�� �9
Y!����<@*}��(��`��b��w���R��cK8T�/ {�_�Dt 츀A�� <����:���S�+m ��? V��P@ϰ���^�P3,� �� �'��%�$t����`���!�]s�� �>@ �I��������|`hTe��]��x�9<���~��w�8#�V���! Y�r�^]�q kن�	�i�����3��)��9����B�D�p ��'b3�� ؘ͝�v��$� ֯^		�ay�fe ��C����ޝ^�d�D`�8%���'�F�`� =��hI��5�i����P���鵙N�� ��Hb� u�o�@)� ����OP 56MsV.����@H(� v[ ��&�
��P ��Xh�b^>L�1�D��ނ��� �esƵ-c� Q��~i� ��5����� �pJXOq� )�A+��j� ���K~�� �� ��Z [��%��:�3 $�þ� bN�`I� J���ސ��� ��۽��Qs �E�c�C�t �
�]��w�xFR �9L��� 8Q�H�g2 �!*�x� �
�w�����H�����N0�	���@s����X�U�
� ���w� W Jɩ8��	� )S_�|�! P����Y� ���8�! w�f�e�s� �_�$�v z��ܡ4(�!�@�Xֹ'Eh"��9 ɭ YK���(	s5�� ����, �
��@F+����ܞ<!�J�<TH�U�IR�� ����[��^?�Ћ�� b	��� �Y0�9�� �i�L@c��K�y�v�ͻt#>L�ȣ��{����� 2ڵ�\� ���Ży �Q�T��2���	г����rQ�@}�Ҹ���y~ ��0[ �B�O�w qi	@�_R [h�|P���ʦ��W/������b����<��E*��W���]��}_���s G.�� P(�V����%�i��1�(��a5 Y2*jn{:�Q��]D����� �����" -�{1��Hl2Ý@��%� �ﮬ��rN �����ʆ ��]���� 8c9_�`�!L���OS��{P�'Y8@��#׊� ����a� �M�Π�Y )�-	��$�{�!.���A% s�Y^d ��1�5�[ Z!�/��'� ��-ߩ]��N�g������ 0�YtA� ���l= ��2h_!�{ ��U���^����`<[ ��3)�'� ���+��q������ �����>���(��X���g3 �Y
�VQ ��R��A�� ��b7��� =I1Ł�v�N��xs@��_Y?�c ����t#`[K ;���ex��\�N�O1 ��8[�e!y^ ��Y(S�N�?���=	[�p� AD��k����VW���O� E��\��U _H��'[�~ (����`�����1��Xq�it����� �� �]�0�?�G��O � ���+���.��"�� ̄���h������8>���O�᫢��)�0���/��|�ɀf	?�W��@1�U�H(@��"� �qW�1�afP7��p@����\� ԥZB�Cr�����b�j/>	ȯբ!�2`�|���SA�� �! ����}a�2W �$S	� �_��L`� ,ӿ7�� ���P ���o}:KU A� ��kǷ����f�Ȱ� <0�:XO  ���©1�� �Y�w���~ )@�(��	�5<JtM�pS �D�Oh�m
��-� 1�\k�=(�N����7��	F�zuyU���d��:�����'?�K��1��Q��� v���� G@p2ZHX5J��N�����~ ��%�L- jp�r��� /q����J� ���_�N��� �"U�H+�$�� %�0�a�X^Z���[���� ѝ\���) ߍ_A��#� ���j���p �fh�Zx�G A�.�S����%�q�1� h@I���n���ȴ ���܀�sM����y f�� ��<�޾Lnd�`Gh�@ ��&X� ���ũj K���B�L X�D�{� ���ZY��.Ғ@]HG 2��K(J�/z�X b!�d�� �a�t*�$0c��X�_�>N\�Ӫ��s]�)L�	&�v ǀ5
�� 煇a��P� /;Y�(ʝ�Ac'f/�Wwİ<�+ &_E��ɐ�ͻ��wV| ���N�A�3�ˁ���� u��{�~3x� _����o� ����F�`'C�)M�^��� ��R����ڀ�m` ���(�`|� L���/_� ��w�JR� 7��6(� 窟��˾�v��|^�H����� ��K~g'�k���wԘ�P0��#�k��K f��)�	�� �P�|e�ȶ ]ָ��ʾB���1���J3 �S��� �2aX������́�
U�Ӑ/ߗn:�H~��� �D�τ肢 Q_�t�g�;�с��/��@��)� XS*�G ݑ'��0� �%Fi��+L�� ��$H �b�T<��� 2�X�.*\���Y#�j�J0�^=���bS���Cy �gk�I� Ȣ�Yt`�� /�yބ2� ��WbK} \�����+�P_�IO�`�}Y -��s���N ��a/ ~���d��8IҀ��P�bK�� �0�>O��)�G{���, �Ks��_�%��� T����EbO ���2PR�Y �`���xq� �J{�� ������� t_�N.�f�ev� ���߄ �e��w��� ޶p(��r &=y��� ��H<���t�"�B.��
�ci[ ���WJ��e _��P�&A ��3���j�J���
�\� p;��#���B P���� ?������ %�6�x�F�H�� 2�h�u�za�`��@�@ ��Ao�5 �t���O�S k9�g� *v��YU� <{J�6WR  H�mxY���t�Y �ZV� j�PL:%~:�o��(����" �[Q]`��v>Ko��L_Fǵ`�>Ŷ�;��� �@c�P�� �ͩÄ3~ ���`fS �(���.�Y N1;�
*��	#�"þ��v��� ��U����R�mި	P� ղ�e� ��	�V�fs1?� {��:R��� "ý�Wĵe 9���q@� EY�N�b� �#�� �Z�~a=nĠ���z�����0�0�- l�K��%Ţ�c.c � ����'�3 �k	�V0�; o�s��-�x ����(��* ?W�I@��� ��Z_�Pf� 
�@)�!�^@���9/| .�I�&RP3�� ������gKLK 6��/*&n�8 ��[k�h� �ޓO�R� >����� ������� �:m(�gwY;�[��ẕչ� �$aZ��1\0�Ί��L9.�g ~F )M�!����@6.��˔T/�\`�� 8vdǗxA �7+:��[�\� G��X_�z� -
���	R���*'��e�L�g=������ܮ�Y�@h-�d\�� �']{)=��g�1`�JD ���H�O�Fj����٭i@��3 č�(��� h�J���Mx \�P����o, ��Z�� �梈].�� ��k��� � �[��ZY �,i��G��>K�A�۵bIF|� ~�g!PB_䳞'���@*��, ���ӆXs hR��/�� ݋�O�G}� Yɰ Lŗ�E-���� ��Z�& ˕��
�T� 	+��P�%� �r�hQ� ������� \+��wAt �렍!N� �f��j�\�0 ��'�U� ~��ȌF� pt�b���%?2B�����!�~�� HM��ީo����y@��#��=��JÌ��t� Z�Fd� c��8I�% [��fh� �}����������fx-<�Z��03�:#�z[���Ԁ� ��h2'���u� dt�Q���F�M��\��0#� PVE��a̓���� ���RL�p���0� A�{��N 3�n�)4Q ��	H�J�� $^�\j� �O���R ��dV� ���w]LO f�X�p0���e	 R*�g ������Y �L�H X�:|�� �u4�t��d�0������z'|� �FI��S?$h �$��� OI�^J`� �1���a� ��b	6�����1�X ��S��*��rH��7�K���}�v� ��F
� v��@a���N ��?K�c���ܵ: z�p�h�udX�� Tb����� ,:h�HO�[ �e/+�S^�� U~9A� ��F\)�[ ��hHJA�.�q_@���)��� �M^ -!��:��LS��	��� R�,\��] јa.�VX�,^�S �N����ˁ(�8�Ĉ�Cv�	\�����U�����r� ��v�j'A�@0�Xs!� Ma)���6 �K;�ڴ�! 5lE:�y�_`I*��&���Ox� ��#�
��$?� �h�� V�+�"�3W��#J˾���UPA���P��/[�j��� K�'#��� ��A�W��Z�r:T�ˠ9�[���@ �"�/�m9*� <���� ��1�!�L�Y	� ں:� l\R�6�k 2���߰ո��_��ȶl ���e���i<'�\��h��F���Ⱥ�Z�A�}��� �I�q��� ��N�]/}	����P ���-�f~� �������@� ��)�`/�[ ~��hsNp  ��V#��� ���H�A�8 _�FsBY���tc �Rh�J$)��җ��D��+� ������ى i����z�����#-���"T ��� Y	(�1��_ }'��7�- ��glsOC ���Jx�B Q+:��1G.�|r ;�2>�*��u���o ���a�|�-߆`�)�3 �Q��i����P���?LC,�(�ʝE��0����@��� �,`(yo ����`�~� �[��R>Đ�N?�� (�]�v[���+ѿ2�SU8� ���	pW� dwF�;�u/�' ��U�C܁
�)�8] �Jr��� Zw�HP�% T��bs�� ��>�"��� ���]��� �R��$�^-1�[���஽ #�g7���� z9��.�I� �'��	��q���a�(�/ ��F)�T< �K0��N��8� �B۴���ȩ'�Yu��.hFv� �X_T�a*�	D��� A�/L$�t� 2Z]Y�.P� ��� �Cv� �_��Żr�p� eˋ+[Y��Ė�4�q�$�3�����@���� �!@��� �L� ^�X� 酓�n�; &E�\A�y�f� �ڷF�D��N�2O ������� �<s]��4[ ��Y���! �
�Z�HNaZg�} �#'$8��R��S�'��^~ ���,],��. ���Y (���:lt� �P�ì�ha ���1�%� �/:���v	 ��,`�� 1�
�����4׺�o� �,5�@���-�j�d3 �Al�LF��w� �W�=Q���Հ�P��� w���&D Z�`$�� BGh�������D�J��d %�j&)!"X��Hpݸv6sh�p���"�=�� ��0�q�#��c@���v� ��zÝ�V� ���+�wXK J�������b�EQ����W7r< ��-^J�w��=h|�)�������"i4 3��N�X ���V��� ���z{2�[��O�!cW	� �AP1���p ����H� �h�� �Sk����� ��g	� H�d 
�tuRT�Cn �\2ȣ� �J�U��W�金���@I
�������t��?���߸��Ix�$ ��<χ>\>�� �'h��� i�J���b��(��9�� ���Z���U. [��� P�Ny�n�����{�  $�`.� XĈ��ZL &�a��������J���ϖ�D�� G�ӹ �	X��˸ 1�e)�f� 3�I�� ,�.  �:i�@� =V���G_���. �Ú
'������vpG��k}e&o`	�ՙP or^�� C$/�?��Q ���-Ic�^���~��`,Fxj �$�R�%  �\�.�q�!�e��hNw( ���� ]���S 0A3+�����ǿ�� �� |��o� \��O�8T`���P�J�b�-0'ؾ�a� n �L��Bb 4�u���
����@�(� �W�85A ?�� �#��{�� ���OZ��_��B��`H"E �mW�ГG ��Lq� /����ޒb����[׼ ]�B�����1E;�������m]fWvY�+� ,�\8~Cw
?��� �>`�# �h-N]1�& I�wώb �4��P �%�u�- �o��B�H f�z���/3 ��$~�� N
ꈀ�Q ��c'�ihy� ž�C�X0 �L�Z�� .O��jo��n� ֮�T�hx	B�p2@ gW�'2jR�.!�|��_J(������0��	��t�W �!	�W`� Z���V� ����@W� �x͢p�jl ]������2�J
�؁�� ��������V�[0͝ ��*H��	� ��]��h�� Q �k�x�Z� uG�U<�v� ���@��� ����\h�:E� �^�݁ �[����v���c��`|�< �$S�/'n ���
zx	 �2�}ǜ�:�w���m�~p �4^����	���XRn7�|3 �.�I�<i ���$U/s8���RZ�~�  ɋ4E]��-+���\@�դ �V���1)�]�5.����c�� _Ed/3��N��-�n���d\ :~��m5�:sЀ�G��$�+3%�5���a� 
��	�NH!�| `������-�^˦{���� �B�w�LX ?�N�62�� �
��@�y� (��K�H�
��� Z�9��-|� ��?R�Y�I^�)�Ag�H�����X���l (7�׵�� ��ʀ��&��8K���P#� �})~@�� U�>d0� ���q�xu^ ���$KV���>�v=��	�H��A���/vJ=��'����`�����X��� �� ��P_�h)�� N
���� Lр��h%GD� b}O_[ ���C�$;*� B��%)q ����@! c����  ��aZ�� ,iWx��n AQ!��vhE�P*��� �[ �@�؉�];��vw���<��aK �?���A �u�����K �n髩l�'��|t �5�j=%]�&�!�H�o� �>����Lpȟ��)~�sK:� j��C� 2�0��	X�Ƃ ���( �^���h� ��'g�@� �������( aE!��p U ��/� 9�?���}X�/ rUء��1 ���?Qɛ ƇNl�Y�� �]�6��f{� �h�2Q�N ���w{� 
Y��%S@��QѦ���ft B�@�� ��e���\3�] :#�+�Uu.5}������^ny� Q
��� 2&=	����`q0USH�9���]ā�P@���_Ka�A��j��~�� 2�!@F�\Y )K��(��P��*�U��.:%��1�!N�����o�y �w\{�ӌ�D@0�$��o嵸+���Ҁ�%�A��O���	�Ũ(e�P;pD[&o���h����q�X��	��' d�Ӑ��� �_�؁� ڌ[��0 �;�3��хx� $�<��K� F�H�/�"��1%�����9>j�:� �v�PW�^ �����Je� 1� �*L�U�HW�[�� �,ɀ�X�F�� ��s �Y+�W" ���<�� �*��q˷�;�� �0}9� _P�g:U\H?DI ����� -fwt�\����$`�.
j �h��aU ,(��k�� lZ̶��b PN#��,�� �%�3
�Zhi 齆�2 ��V�����7N����FS �_��	�� �Lv�"��
 ���Z�� �ǧX � sk���/�q�D��1��+.J׈ �K2�; ��/�ňz' ���E� I�ӧP鮵�V"�^@#븐� hՀ4J�͇ i�&2��_K?� �.�sq	>�� %����nӤ��J@h"S�K�@#^� � ��]3s��w���S�,�2Nx>�%[��� b��a X&�zo� �����	�0 ~����g��BY?�b�I�trP��� $�p3�Z ���y`� �/fX j(m��Y��H�_	 ˮRs�ĵ� ��o�`�  ��O��� ��$���;Ǚ� �1l�L��� �~V���D J���vU��o ^bi��mkPH�_ Y� �\Z吸 ��W�k��H ~󟗀�����n ����$j�]gٮA�)+ ��T#��Q-�����)�� ���h�Ud_��bXj��~���ԁ�6`g
 �����8 �U�B�I� ���J���� ��j�1��# ��,_$� ��!�T.�0�OQ`+�א���F�`�0
ʸJ�b�(�1�ȱ4X@� $�2q��-z�:�n ��IS6��%���q�d!���U�H�y �m�� 0��!�A� ;(:�1' ���U��$?<n�G��R� �Zz�F���_Q�� �R��. ���r�� �����, ���驭a*�͝ ���~� ��E]����ݽ���'�� �ǿx�� ��זr����g�z���� ��[)�>�R��l���tHv����ЃT�ӽ� :�Y�l� Z��P�� �xs�� �a��p~- �����
��<�}��)"�@�dh 0ش��� ���*=1X( ��GM�@(��� Ch��� �2?[ ��� �a��U�7i� ���ɜ! +c�f_:����Րj���� Ox5�e��� պ Kٸ��!�Qh�[���_t� �U$��� ��[���F0ƀ"Uqw B ��A��n �=L�Z.����1X�q{ uYh��� :����w 6��dv%�� ��
-Z�* ǃ�{o�5 �EQ`���� ���_ 1j�"�ݰpg ��}�,��@��?�P���z���J��.��2@u]
 �@PT� ��Ǖ!'�oG,F�3 1��\x���W��� )�_� 촞�#��
 ��CԲ2 S���	5|� R�]�����% ��Ƣw&���Oi�x�u ��S;�'�8D`%�[@ �����3�^�����H�� ���M�(�� Ab��TS\ �`	�,����tl��Y��:&�  ���8 ���S	 �N_م!� $,X]�2k$�J �#N �!/�[�	h�ns�xJ�L>�@�Z0�� �[hjN$T ��p��� ���B(� �3ȱ� �-1<��* ������Z��P�z��"y� � �B��@\�������Z���e�(	��o��p !Ӱ3�Z�� �������.0*�k���� X �,S�Rhd|� xD�KJ� E�U����] x`����\ h�[?Q*�}�.�a ł�R" t�	#�LO ����E��<) �3y�-k�0|l �M����V]Ԋ ��=��4~A����; \`��	�c�N�� ZSq�#*x@��	�� Y�lO��Hv!\�#&h@,P��Q� ��}ֈb�`�* �3X[�(ԟE�$�ņL�JR�T%��A �Z~`�F>��?� ��"h�t$�cl d��*(H�S� ��jf�z� �?=�}r�	!j�wv����� ��O�)�� ��5��C]�h���o��_���L��X�`�0� Q�Ǌ�r��?u����!IC��� .TЍ~}�	���u�^��`1����)>�� �<��� ��\^#�� tbq/�L�b � T��� �_��L� ���,��� >�����PE����z���*�h�.@"���( ��젱� O�gn��� &3~9�V� >pE���� �����%� ������ ��1[�(k ULR�Q��E ��2z�� X���rȅ� ��P��ho aH޲�*�L�1�ĳ��D�+��0� ���ê��	�B��_�(� X0��
� ��� �!ˣ�K�� 1����6 \YC�P������ C��/��p;��SfD�O� �Г��~�� �a��� YQP���� ��/#�e� ����"9UQ ʉ��Rc��w�\Ѓ ����p� ��&�/�cQ (�5���eZY����\�v���P�k��bG)��0|�j V��SX� ����]5��� �j̣� X�?��V�.w��H�<�@�l�EA21�!�)� �$����� �S^è���)�� g�� ���8[昄�	 ���k2� :1�b��D ����8�S %��e����mH�^`�� ݺ
�ד� �(�iVt2��[!ۡ�j�Y1 ?��ε��` ~���.���lF�@�GOY �6�9L� 0�hW�{�� ��GKa��1 p��H�$8����h]��  �P�*��	 �aݕ�� T kG\M� 9���͆n �8{���� P����-g ������ Kهջ�k �fZ�ǂR�4 c�_��@�� [����*h> ������ '� �ʁ�� L^�8%��� *ZT�a�̩;�߀����+� l㽄�ꤘ VT^�F~���'*�=C��� Ǝ���� ��
1� �&[VϾ[��sX:'(�l�$ )�!7�y ��2�S��� [�$��)�d N�{~'�P%��k	4����3����9�Y V�B� ^�!�`�����}O��J�C�� � ؀�pU�!���*�� ���hxb-<TXg3N�U&\�j�b�{੻�u��3�ɵ<��	��ߘI��| V ;��y�� ��Zf	�u�a�z 5R{�$����\_4�؝V�R^� ���<� �| �B�_8��P�����q� ?�<� Q���� h?>	}Y� b�Br�ĥ ��#ܝ�� �缭��A���������$�����39�f�x������v��E�5[��@��% k�V;L�a8 Z��wYH� �/��i�� �=^P�5ru d���ݵk� 8-3���@�RY � �z4���A�j( �о�F� 
`��H5Ţ ����}�%|	vr1��'���< ��!�`Z���	0�U���= @�J� �p\��Y��L�
��j$���V (��>�I;��< ;A�O� =�� p4[ �VP��1X� �7Sb#�@ �mΐ�\ ſP�Q# �W�f$��  �)�(������ �o�	��!U� ��S5OiH��`�軐 )���Q-� � ��i1v/�2�Ϸ�g�S��R"!�Ľ� \x���6�_�	lS`���5���µ!���2) ͕�SB�Y��A�j|�`�� ~�t!�5������U� �c�4���z�WN���{�T�.�w} ���# ط��d`� "0�[2,�X  	kho� �g�'�VI_J����͚0q��� ^[���fP p��@��.�����
>� \Y�Q*�*��'��}N hH
(���X��K^��n ��P)%1�� ��h�, I��2�U ���5���) ��c��Y(�ɝ�o ��� ���FGyڟ 1{պ���2˯p�D���=���5�  �zI�� +�s�a�hW.�p� ���	��y� Kx����), ��'�߄ w��0��� H*׉�8|Z�[��Q��L) �ѽ.]��9�������S���� ��*�	c����6鐵�z�+����� \8ŴI��%�"�0w@-���R v&+�Ø� ]�4K_�� &�d��PG�������.Ąـ�0� 1-�Z��j��d; �(À� �	<�Sl)����O��� ,+��4�
 �iu�p]eB-_' ca�
�馑� �����.�S�f�g�(?�$t��>�� ��]�0j W���C\�%�(`T�v�E !��AI�G>�;Ӹ/2p$��/ "����R�U �d@!-�V$���^��H��:G>�� #Ɖ� �L��0[ �fQ��?�M�>��� �̳����Θ� "v	�p؆�N� U�V� �� �d�[� !i�/Ux(�����  ��H�} @43k+8(�L�!V�� R���&�L�1+�!�ԫ}��*� ���W~Q ٹ	=��cw��U��t���e�96 �'�	Su�n�9�b���@"l ��U2V�S�
�����X� ��wF$�\��d�% �������q���E ���\�(�Pu��p�� ��?��> G�����Z#�@L��wXz�	K��J _��W�����`&\ ��6���' #f�Q ��x]��&�A��Z��@^hK8�1�@7�y��x,(b�D�ɇ� �-hb�l.t0 ���'�"��	�d�qF�p:>Xu� *��|%A K�`�_���
� �!�[*	�X�N�m�@�g' �ԅ0�hs X�- �z���/?�P��V8�ub !�]%� -�@c5a1���A���k F"R�`-*� �y,�%���
ٌR���8�,  ʊ��J[�8�����qB� ����S$� .�Q1���P� \��I C��A U��t4|��@&)댉>�l��0�5��A W3�!�~ġ ����.�=騀�"���X�������� h�)�-��� 0��S�x '��l˕߀ �ы�X��pQRc�D��)��P��Z�X���R������K�����W�ĘZ��H;�{ ���\�_ ��C e�� O��E ��/�XF;�R�i��vt�� <V1�O�	.K+���@����ߒ�tC����	��	��`�b��������� k~�.�QW� ��=�|�~� YX"֢��� �9���� B��Z�0+�`}`<`
�X h۾>-w2zuaL� ���u� �lr8��� �o��T�~ _ �p\� ��J���s ZGš�h7f˰ �}8!v�W�G����b# �VI*��Z ��Y��(� �X�}��ŀ���% ����*(�� ��M�PR0�H��&�	S����C0�!ɵ�xӤ�aT^�A��R���`D},�!�N�\C�%�� t8�!r�]R �G�"<1 /�Q��Y�� #���� 	UsP����8 A�)��D�Y Cr�0�� �IX�>��: Zs7��#V/�� ��KE_&> CB D9\�
l�h�T2�uR ���Y�Z *��& �iQm!�� �Һr���(��� ��A�n�� ����I#�P�K|� �"�O�+�� ����s& �D^��hE Hy�ҭG4� K�\Z��,� �Q���' AM�<��H %!(�ZP��V ����'�E�@�Y!����Z��p¾$ X��p��1N ����T��(�]� �HڹyJ6  _����[8�LM�k`G� �H������ �
Pكecq W �J�ȆR Y2�C�� �O"�G�/� v�5���83B�H�Zݚ {�ن�~�� ,�'X%O�� ���Ȥ�� T��	<��,��!���;� K
�^$�E���Ъ~�P!�4���{�|�*��N�&�	8��P$ z9(�����X/�v`�� ���[�HL#��l�e�� ˞ �����JT�F|y� 0\��5�����G`����� X�$�o3�. ��/�͓� �8�T�K<0@���UݐE �}3aP	�:���8i_���K��	� �J�x�]�� ���3H�/�|�$ Y�`��\>� �tV�7' ��B���> (�#�� ��QM� ^ �gP�HO ��	�xJ s��7G���<_���L�����}	 Ѻ,�� ��> �ʿ��I� �����^ ����Wh >�	�~��� �*G�I YX1;�<87.���%|C�	��:) i*P�� ���0~� 5�"ɡUX8������f������/���k4���_��� �~�L^�����
�0Qh{���j� #$[�6k��8 m��)͉ 2�u�{�;���wp����Q������0�V�¹	^�vM����g�� ��.a`I U����hx D_�k��Lw�u� .��%	|N��:�u )�]����� ���,��A ��U*�Sb�z] y3��B@�z�� ~Z
���b0�W� ��v�- �E^�� ��`/��G j*O��}=o�y� �$�� �����>2J �޹N��� +�l��\��.���	��?ʀb�����<;Q�$T1��z?�a �@�3	��u� �|�E��� �)
W~BZ �up���� �����BO P��Z$��` [���:Ki^��@�
\��$��a��D�� d��T� "c�sh#q, ����\�� ��! �XN� �ܫ�y>��;�$��_�I��	3D$�z ���
ڈ �[�2 �X 	��-I�( ���3� �ȕW���x�L{r a�̧zUE�" ��\|d�q� Y �R��������`�ܚ ���40g<� E�ۂ�SP }p��O���1�q3���� �X�� OQ��
r�� 0�B+t�/ �؉$w�1�D� ݀F;6{8y�>_'���j2��� \��b�9��y��؎n� �a�O٬�E�;�M���좋 Q��0�h�� �*�A�'���� V��g����Qs (+��0e�ĺ@󖒻s� �	���Wl����3ːL�'0 �@��6�w�z�����hK�/ ��F���tn����_��Q\�B���@�#�}-b���Y\�D ����% ^ů�/<�� ����  ��1Ҩ6���{�L	��P �cXDoM�^ �ƶ�E�q� �$��b� ��
�#��׀-�V�~t(.�@�\h�I02����&� �����08?�Gt�`��X� ��P�W��(�
��ɓ'�2������1 *�ܨ(N� ��z����8x��>1�9� ��#�f�� 0uhE� � ^-ߘ�T�� 0S��N��L�(a�pb� ��O��$U [ZBV��� aN8�� �$���>	�	W�ҀE���,� MR '��1� ��&s�f� 	��F ��ƜJ� �<K��{ j�Ҭ��aL�� ⟩��o� �ܙDX2���Q��W�>�� � ����D ���W8~�C����	UY]���v��׺2+ ����P O�3�T4Q �-{b�� Y9��� /�����_w� uQ���t!.w� ����* se��^d" 3�{�;� 2Ⱥf@��X�a	�`�����g���:���
��� � ���']�)&ò��@tb��.H\��_���\Ѓ���Ж� *�r�3�� �yKG���2�n��%�������<�V �ǇR(Ĉ ��7c���|ρ�\��A	���^�u����e ���rEbw�9NP��S	���C@C X(Oڮ�W
&*��� 
 �u� �Z鐸�=��x�"J��E~��� �h+4�i%�>� �	�� ���$6»� t�/Ց�fC��@-W�� ���ZS�X� �),ؓ5�R2������ ��sկ��	�K݁��a� �%l���X ����jR�ˆ��>@�v�a���8D��o ^�th ���	;�1��0�y�A�aUh �J�, ��6�H�"� $1�A%9 ��f�| �����/k ��!�L04_�1qG}�P�\ݐ� @)Xʍ�� ��uo���[��P}�j�����O\��� hX�r��^� �1��b-} �@W񊬪 ��^�C�� 5��m����qJ+��Qp3 ���C�n �`[�T@��,1�ط��?2/.Gf �
��� �3�1ʅ�Qo���Y��  ����[���(�Z@��� �Q��2��� �3٣�(���}� ��&N�g	G�]ȓ� �V��s�(�� 2@��U%��� �0!��X#�|��j>`&���' Kރ�^�	�h�8`ؐ�$ ������� 9�閏��� �ǽ$��E1�3�N��o ��
]�	� Y4~,G��V�@� �_X� ��}��~�� �%�Z��� Q��8��� �f�%�_	h$�u '�ӡ�� �L��3�e`<�s�M��f1�7S���c��� \�D1ٸ0AQ��B��08��L&<� �%�� ձ�h���WrP 	Y*�V(� ����R�
 x$��A_( �:�#��WHTFO�p��UP%Ztq ƀ��r:�� J�Gnǂ� ���!}y�h��$0B̽? �
� (�`�\��K�6�>Ջ�r�̑q��w������ �_`S3L ��̵�#\0 :	����V �-��f�%�^@��@��� �RZ��u�� ��h�)#� ,S(�%�����H�A�O`��;�����$� 	Y�Z��\�{��0V�0� ��.>:��� �P���jw��'\H0��5pb/DVr� 2XY�?P)/��� ���O ؤ�Pg>��w����_��S�~��-s\�r2�K��� R0̶,�ր��E�� �P��X��  ��6>���%�^����ˠ� yo	��F� ���d˦R{� ~Z��	5yJLW�	D� ��
� �0��Q� ���W��r� KP��>��*�nA�[ �3 ��<LH���>R� b~�J��(�h8�1�9�	�#��Q�9(K�+ �!Ͳ8$��`@��AZ �d� D���m3s�,��� 5����Ű�,\ � IF��M����i���� ��_��  	�
�b��6Kv]�I�SJ��xM�n�X [��1�#��t� L>Q�i �7S-�E &�x1�	�������2t� BX���]��b	}v��Q�� �k+j�� [0� ��?�]�J	�'�G$��J= ��A��� �5�1ϖ�� �#!��a ��xD��� ԡ3�`��@ J�¾P��� ߉�VZQ�`���h��)��0F" $���N�x X��-�� AH�0����
� �a��]� �st���@�U2\��"q/�t, 3�h�5�1� ˄ָ
��uN�$�s� ;LZ��hL��Gݻa��r>{��6��f[X�(��P��&+� �)t$J\
(��϶�#���	�U�� ������� �x�u�9�}�+��|]�XH{T;��U�6J��8]�'<L\'@� ��)^2� X�,iӶ� 9;��� ������ ��2UP��;�� �o^&��� ( ��Y ����P�� �+�(@;c	ׅ�oޕ� , ������ 5�>�� �B��l�zDX#�W�"<}�[��f����~.	�X�f !���J[q �D��p  ��@ B�V�6�R	 *�Z!���x�%�@�/������ R�qY��p V�UQh�"f ��jN�q  �oz�'�	a����u�Q�<e��A ��vC\ �G P㝴@ p!T����_>u�|Ki��	�� �l	ɜ�����0Z���]�O��� �IW��`�`�ȗ �����F�� B�d�|2��P�/��i[�T�\t ���4�c��X�r ���A�!�^�(CӰ�p:�.For&� Ԫg \_��?��ze�� &�YѤ�kJD#��h�� ���-8f�4L� ��[+��6��_G���� S���X3� Y��{.h/w=W� >�䯴���\(Rbz �Iu�X� @,V�f������@N&����`�
@�/ q\��۝R �$�L���'},x���X]~0��;�3 �)Pݘ� �t2�� 0;��Z��� ��]��
��6�}���d�> ��4L3N2 �ҋ��I�Ew� ��A��� Z��+琌/ ��8�G��gI�t��[�̫� �f1
3�O ��J���/[��A\��|�S� �����
~�x@���Z��u��3�0Ľk��	h Vd=�Ι{���Z� ��^)�xf� �BN���W 	g_cG��E �+�r����_帮 �G]y�,�������o����Xa�uU`�	����C��2�5} KD$X����~.!o]G�ps�[ �"D��￑b*�1�?q ]/���~����V# O��p�`	�n ��^�voP����� \�kW��Z �������{ �K��w�Z�p!�"���
 �&�v�e¹ 5�<���� �zG�T� dW��\�Z� ���2�� ��@j��O�$�-�$f �VP!� {�2wk�6��} �YS��M Z�p�(�� ����[�wOe��\a ��/)� �N�<b�L( �R0�W�� ,��ϊ�� �)�U�d 2�s���h6��zf���M 	��D�L� 1��k�`�����X��%� pER��SQ ��e�H� �#)���O}5 �[p%�0�:����l�2�  Sh���իK�J]���x� ���C�K1�4 e_.��&��$�p�pL� ��H�)�- �יl�t*�P� ��� �	WU!��;& �� �- E0x~�n	� �L����"!�Q\��ЈN ���h�� �XY� dP�=��.��b
-�Y��)�����Q��`/	�@��x�1h e�z�|*� ),/�&Dn�� �jIѪ9'���:�ܸ" ��!���Z N��*'��� ������ �k�"S��x�d:_�]!�Y Q���+ '�ſ�� @C��R�"m��U	�~����Hh*�% �(����� [����	���Ҁ�s��
(�fZ��@��{ d�"6b�>(�(� ��酠)� X+���%' ��|4?*h��J��+�6�0 ����k{�ɹ� )��-�i�mx~/�q�����M;�����t� � ���{� �wq�X��K�Bj@�^Ҡ��4 y3�J	�#�Dr�� -m]�$@��|2�����?�t�� �C+pWZ�y �12���&����\� /P�O:� �,R�h� f����
A) ���1	�J�R;����2�>]^��ʢSW� 0�>"ù� ���u`) џ!ػ�R�} ��x��ʐG�@��b P�O�����?a��=P�e��#�x@��!X0��Jw�H�� /A	#�Xt ����� �1��(�����k�� �<_yI�H��S 3Ҽ�Ğ�� $��h�W���՛� {�4��>���X��f�UD~�����4H�> +�~���X%�B���=w�R" ��{@����|�&�E<��Υ�_"�L �Y�r��=V����@�	�J Q��I��b&��h-�`���ʃcAC��U� �r=�� ��n�#��EMs����	)�Zu٠�I�?e���s܄��8�L�_%���B�� ����X�g �^��ڰ�1w� |���W�Zqc�H�̰�K� �h��f�pF
2�P�� ��Ƥ9 }�^�_�y4��W�qb� ���1����j��ǫ��h� ֟v*��5 q�תgb ��R�� �0)n���g�+ h�=F��8q�ǹ��W� ����/�~v-L	�H����P�����}xv G�uf=�� �Z�]�I?�UQla�1�P 8�R' F�%1�tz; -!�V���X�a �0�ʫI�#������ �i��҄J� �C	�$��j �5\�V�z;Z˂�-�T�%�Ҡ��� �1���!�W�� �<@��_MR�� ���
��	0pZw��K���_g����3����	�X�K|��^�+� !���� ��\�઄Y �2%Q�f ��e����?�]�� rm��H �/�W:���� C�P?˝�9u8 S�*�&�O] ��t�Ƶ|/ e+�V��>�h'���Y���,�Na<*_����J2��@W����I �e���>�H��4������W@����`�n��;� gI�`,� �(��� ��!	ـ�D }�(&6͗ vKB��h�� �[�(����1/��_��� Q�ҹ@��p1��>�� ����j ���_J���M�֢� ��a��gp��� �h��������3��[9+� �&����%3\d����# yq7.���� ��_�$�j�v�Ԩs� �G���\%�@No���4 )�R��� ����NP���# ���z��	������ݙ ���	�k-����#��\��
u��� 2����� �%���\�H�Re���� A���$��/ ��3�?Q�L�ds���j\ �<%S�H	 ���(ʌ� 0�&;�%�8�� ���wC�0��^�G ��!õ ��>��=[X �0�h�E� U�o�j��&[� ���d�$ޙ��`r�X zo�������nwB���/�]r V ����F�0�\PC:�<$���	��Tb߀� @O[��k{����U������ �Y�*���uz!�0���9	�V]���+ ��5������[�x���/��л�Z���'Ƹ��`���a���l� ÕR��!qKH�L ��`'�j �"���fX�*���P(��U���9�x} 6	��i��
]E�� �z�[� b���B/p����LW
0�筤@�������P� 
0X	ӱ� ��x�R1� d�*�<�� a\��	���9�8]�Ȑsh �|%B�?U	 �<��!��� �؄�� J��$K�_
�ヂP��0ۯa]p� �� �[ �l���
�<(j���~�$���w4��De�0�� *�l�^x�� b�]�c����� ��@�N���,�Ba�`!@���x�y�O= �-N%/ � ���U��6� �ӎ�k�G�9�� ���R��s �Aδ<4� �>w	��*?�}Q�P+�D������'0��T�ؖ��p� ��2q�(� �M��-��:�o]�� ����w��B h�6QT�� �\���b��V)�	{/L$�z��?�X��Q�������/�m �_!�k(*��@M�B�l� 1J�%�X����L� � �Rk��h0� �-���I �_��i~5 �W%��������Q�M�� 	�wڟ=�Z ��*ILJ`} ��f��^ �1�	�_� ȻФOd���r� �0���U����?)v��K^�r�I�X &[�h �^�aSQ ���˰� �ݜN����V�=����� I%�����r f)�^pV� T*q��� h�`a^��4<��� ���W�[ �_�Ah` �"�C��D� �;�ܓ������f:�� �ꬅ������؇<$�:㦈0 �?�f:w +$����X �E]���9���@-vNH�� ��͎hQz��� � � ��'�ٸ� �8���Of~Y \�D@_0�
q� Ã͈Q��.u� ,A	� �T�S �W��f�_ t�����@� �r8�A� �K�f�\��=��0
� �ɘA<C���$���]@� ���
�sr1H�k�|Bg�Ӎ Z���
��f���y ��;�����I�mP �h*{�^!� R	�24z� �kC0^�9� ѽ��*Z!~� �в��[a}.
�R`��S�཭�%������ X#�3��l�	���{���m8�X)�ž@ڌ� ��Ș�O ��><�C�����;�B1r� �.���c����SW�XZ� �&_��xC��� �Z�� �L����u��8%�������H�����&N�	�0 /K��rMe���% ���7F �:�zu�5p;
a˻�\�.', ���1�B!����tr� �}K��?J� ��/h)�	�� �\D��U�.�'  ��%�9	Ry�3� �&��V �Vb��W�� 7H���! ����Y�v� y����M(���~nw����1���u>��� <[� : �`�?Y���fX��� Uo���` ����w� ����p�*��$g 5M�!�R+��[�	����G��R#�] �W����>��7�U �!_��X�(�㹀	�| �Ё�CO���_�+�ÀSǈ�E Zh��RT���"�ؠXJͅY �3�%@	��`���B��^ 5X3Ϙ��&��߂!����ёb�O|����� ����� �����a
�%�B��V|?�b0w��_�x� P�#�v����;B���� ����U �`�Y������� 	�X��� ��B0�S@.��D)	e:�I��	�Y� �%��@| �&p�ܴ��O��X}���o��	ȉ�:9�s ��`Q�N<�B���uٯ�LH!�k�� b��w����'�� l8@�T� ���I�� R��X�� �2��q�� ���ɕ7� �e���P�[, �S�\n�p�� �%,�{��R��" ���3��I=xu 5�E�"��� Uj���_ p��s�%1 ��� ]I=���~�H=������N��@����H_~ �/��1� �~�A���� �Y/�lm ���ߘ��0��FG�� ��3�y�- ��sxIe�N ��!*C,;������� ��
!�/�-i��@�_ ��d����G����R�2��%_��k&�mк��y� �
�s�� �_�.S�f	�I�v �0���*� ��,��	�_8T� �X!ݱ� q�`���P B�S�Q� ��u$��� C4閶Nf� bK�t�0� hQ,mJ�L�%�U�� ��C�����[[_ *�ZT6i�L%�Xg �s�al�1� ��>�V*�궎��@���� -���
���w� ���@�Z� -��p� �ٵ���b�X1s ���5̂p�� �1�U� 2�S-^kIb`���R ��	���S^�0J�5 ̢���� ����X^��: ��~�æ2c �	��X ���GY�/]�q ~ao����	.*#�`��U�T����  Áo���C=�����> ���Q�㼷 $�<V���h=ʥ��������� *+нKY ���5��z �Ե��
�h7����ʺ8�\ S�,~�� ]���LzU�V10H� ܁���+�<q� hJ��� �%��5�� �0�
剟3 ܅%�;�?� �0�@�� -�d+��q>i; ����(����\� � z����8 k�}m��[ �)�	 `�!ŀ��|�2�R��<^ �� �J��[N�� �cm�4ҹl?����3�h /X'f�� �����
|�>���r�Аm��B�T� Y��� ��R�8� չn�aD~� ̽j��/��� �#탪c� �u�;O��6 �`qf!�?ً����Z��.	�Y#���4 �)R�&�� %BԚҤ� ���P(�\����M���� ��bf�ٰk �Yz�)� 1����4�J��� W��wXtvL���p�@�Y� ����q� +�S(�\�  �њо �{;�R�� ��e۫����H ^h���/*�W�Q1��L��f�;�À����`����C�#�u�� �]�|� ��ƒ���:L ������n��w,(J�ς+���0H��Q�	n�#�qB2�k��XP��K ��D����P��[�&�^�E����q�0)� �+s��p �h��R�� $��fQ�rP �d}�O��~�T�_�4��id� �*�7���;���0 �������+�K@ٔ�NZ ���uL<�: BQ!���0��8W�C ���� a�&��� )�6��  \�*�t��:��@�p�� +\��P@U�$�2=�`X1�#C hi}�Z� ��!�	*�X{ :H,@�� �	W�)a�<X�O,�Ā&���Hk 2�@��� [
M�������*Ŀ�&� ��7���5 �U���s͑ '`�X���h�c �1��z ���Q�KŶ���.�f1:�ז
 )�	T�2aUl�B��I� K��n"�o :�a��˸�j �{#X��S� �E*�L�� ������ ��rf �����-��'+�U E�&[�M��%$"ԧ ЕH6) ɛ]�m���DP"��N��	 ���IX>�� �l��*.�! ݹ�׺�" ^�%���y|���+��V�`4�  �X�ѨjX��	K`v�A����`�� �)� �ԓS�R.� ^8��/��3�,�T�?s�"��h|�S_3�� ��U�.
� �v�O� t_�$ɪ?҉ |�3<W� -Z@,�����q�PQ�*0yN$��=ؿ�j�ĉr��� ���G�lc.�� A��!U� �^#�]1� ��0�P��b���nk`��`�X�0��Q	 �����H ���̪"� ��8�\Q� <U��j��.��~3P5R�c< Ц1�v�.A�� ��GQΖ�����K�� �[� =%t� ��E�&����LP�Jv_�L�,P�b C�!E�i��]q�GP4u�`ը �%�s��  2H8���Z �!B�����R���6�`: G.�������(� ^�hrx� 2`I_Q/�{�k
�`5�� ��zs� ���΀R����� &]y� �0�r$������ء��*B�5�H�2� ����~6a� �1�?��#�h �D^�}A (ɸ|<r>�=��{��%�:k��_흉�@���� ��7>5S$%�� Ҋ�wb= �n�`E�\;�� �0,#"
� h<`�i�� Gd~ ����1� _��NQ�M>�,�^.V ���C��RNP����t��, 8t ��� ��Wt�)��	�!`� �|k�]� [�>�K�c
 �B�eo�� ���b�j�0�� kq���=� ����^� �N�D-w: ��Y��fs_�N��` ��) ˫��~8� v��7!���Y�a�QP��k �|*K�� �H�As� ���ۘ`n P+ʉ�|]��d��_ 	�KF��H�UX %�PWΕJg�DC}\ ��XSk ���{ 5�� �H��S�-����v�3@M�f�� [�@�~��\�� /ú� �3B�[(���M %\#m�? �FP�峿 0O±z�vo��s@>�π����z< Q ��f;� ��D�m��.4��
��ß�5 (����09 ��:��]�$/�����r'r�g�6�`�X��d*��30�V ޾'&�� ]�!u�_�w���z���>jج�{� r�)���UP�W 	f5P�ʰ?e��O�+)p\;�4 ��4r9{债�$�p�\�� :X#0Y �b��ő`����� �1�P��  ���_v�4Q ���`��X ��ێP�f� =�(�[ �
�2o�S��X^!J�Oد\̅�$��-� �I�wOV�C v�*����2ރ����h�& �a^(V���`e6���1 ��^���� ��PS��$� ��`	ى��]��������a{ـ�hH�D�� 
�/� P��i��� �n�T\�(� ~�Z��1lL�[9Μ:e����� �Z{q�p�.���%�����-��r�����5�@Y(��� ����*� �1!��̷\;mZ��(�.'� 啃V�� X	�ߺ~D� ��_�.T ���hC1 ��+��%�� �`!�-�� ��T��D �/���HL�[ U����� �>~��	P� �A�Q+ ���Y��\�vp�-x��� 	!�~9(h��+WN��܃E� 3�r
�p-�B󸯃 �IQ|�X��Z�v zP��Q� О�G�� �s�JL�d������ ^���XS �v�z��q�$U&{�p�@<!�t>"� �p�,�CJ ��)�( �	6[�� - �!Ё�J��O��Y��� �;��r]ù-K�t� )no��H�R����*� ]����8/K舰�	�o�r��è�@�� �y��_ w�"�E��� F+�˰ i?'|�P��; ��L��� 3!Wܮ�J �E���%p �g�fl: ���)S� ��MI�Xtq 1�:�l2 �"h^���?���O\0�Y� ��5=B��|.�O �J;�6C$~���` 
 �TZ%�m�� \!�in:y�� �����L�) Z�FN�� Y$K�+�E �� ��db ���ؐ���U�t@�5�3p� ��1�Z�4Ր~��z �;������էh���@���  �<���aL�� >���Qc����h�4ֻ'� �"��S�� p��`�C�4�0�v$.�� ,�=�Ў 	�U�S]�)ՠ�t��8��} �y�X���1 T0 �t��6��\��u/� �Kz��� W*����l ߖ,{K<� :u�E���oq>ҘÚ%[�A��`z:R� ��`�A��|ŀ3à.G zː�%�[` �Y�/�RZ� 3e�B��T�*ac��A��Zd[��� 8�wbe� Q�aW��$j`��(yB'd���
�R� w�@�%\s����H���(:�V�{�%���f E'�Z��A�:�� ˶�l����h�{�����x� -y
B��+ ����83&Y G	Uh��_�����2�X�Q �����gw ����|ɮ_��>� ��B��j �b�$&[? ����h�	�j�t�����2�� �?�׵��� =P���S��2� R��5?����K�� �W_%�af�U� ����)Y o�1�^���!���:S_ r�Jm\���],�������9^O����`}j;�g�Xf�@�ö �0p� ���1��.��R�8�`�h�9���W;�ܜ�s�72�ڒ����@U�� ��[ �k)��� ���+��A =Y�x�� 鐔�K�5%���v��
� ]S_ P�� /I�ٳx�� ��A(�^ �h���`+ �B��6��J ��*D�ΐFV(πP���X �����]��QU�q
C? �Dh-�x��� g��� \��MSw K��傏5� �Tj�^Q���O�ᐔ��Y [��KA� /(0	�h��L� ~Փ2�� ��8�� ���C�bHz� �������I eUb�� 8y����%`pK}�(���t�H�K ]�WH�.� 	�)һ� ��
]����p� !��#�h3 r$"�����qMCg��H� t@
�0<E� �bk��	�8�T����c �7�\�� �h�Tk���q��ۀ� �eY���� _t�IC�ݥ4�W�`	S�� ���)pI �0�
��kN�� .bx��;�V sF �փ�X��K��'/���pv�ح���Z���%Y[��B: �PR��A~ c�{��|� �.����D ��LgO�, :�w��G ���
��;P1�� �b��#Ζ �-\�	]lyx��(p������ �Q����h�x
��k� �-�Zz����&@�����%0� ��SY\�jN6��@��	 (�V-��� 1�/�<6�a +Z�R� h�yfn�� �����	��<�ڀ��\���?�W ���"�a/P}|b �E��1��|���ķ/)\�u�
!pP$�eRՀ6���� -��9�%��?���[�0K ݄v�hX� *�#i�p�"�c+�) ~(�<�-$!/�� +���9��(��F@}���
K�E!��,��	� �r?�0��H�$ ��顗n��p6�Y� 3`�y 2�f��D�)�䫨K.F �$��+ ۉ)ӿ`� ��Ah̠B����1��s/� ��V���b��pwf70�c� ]���CE��Ⱥ�� 7�HPV kՅv�����x|C:�P^ � $C� ub`�N�� �J���� 	r����d ���z��� �:E{ǈ�;(  ���� R�]�,MA� ad~��ʣ� \)BP���q+�%ඪI�Q�w���>��`y%	v� g@J2\�p&������Lz �H�5�fXu� Qc:��� ��S��/ ��2�H��_q  ��<���3 �����u 1��`��-q�p� Z�����%4���.��-�8
�6@P5 0� �)Չ�L �Z�g{�� ��0�=�� ��w������R�� �p�����Z*�`�(ˀ��ހ0g \X� I�{˿��U�`���Ŗ�%��
C��-� p'��� �������� �" Z��u!-�� �/�^"�R���¥��h�v�DV1 O�"X~� �s�Q�� dS�BWۼz�0eت��\~����� ���\�Z���U�`� >�c��!�'p[ H��0J� Ο��];B� �"S_�k�lxd �b0�C@2�-	�s���� 3Y���as��? �q�lI���"5�� 	�Fɯ_�'z( ݐ�ؤ��I1���٠`�� -��>��u ;�j��`�(� _i�&��� �����x� ��
@�����x�[��p�0� X�q|�c���) Ջ3�� �#b�[��i���w@�� ���� �Z5��P^`W�aq@�3�~�� S��[̲^ �
�n��j �I��ʮ��_ ɪZ'h]H ��:��C ��lb�*��|�=����_���%`��pG� ����4_9�V��(�w	�-�. Hͦ�P ����Ĵ�
 �3]YS�� �0m5y�1 *�r_��ڗ a������f Q����� ]�k��74 :���$��� 0!ȉ�� �Z�Wl��b�J UT�Q�+��� � &Hs� ��`�&@/ j�_�Da���֧1�Q��? x>�3y � ��h��z
 I�04Jj�� ϪP�iKA���G�Z@�
� �|j�_!k���IJ�
���R�8̀���Xh �&�d f ��_�3L�[�4`�RZ  �)�S��Q�
A٨ě1�bN�G� �9� ��AJ f�����P 	`��
�T� A�%�8�~* �����@�/|��րSѽ�kx>X��^|�ـ����?Y S�2c��[	�������&��c �`R0�[ X�/��� ��Kv���\�/� �X2�Sh� dW耈 �_ ���X O4��* ��Z^S( ��1�����?����@��x�J ��T��ӈ	��<�X J�r ����VQ"� ����0� >`)(�	fR �F�A����~�Z�#�� ��$%�J�� Q1L:��[ �-�c%��} I#R`�@	� ⱝV�x�� Z��z�);$.L�� [(ѫ�� 6� 3���U �1j_`�� /J[ �S���v���L׸��%� �ox.� ���\_K� )�@]V� �b���jn �1:���l��fa{�Hv!'2 �=Z� =�(P~�� �T)�Z`� 0�U����H��*ٸ� r���`�����zh�ء���H�˽)�r�N� �"X Yfh��x0s/��C�3��h�p� z���,�[{; �%P� e� �&9�ȥ �b�΂� �Q�{�p� !_��I��� �~�y�	�U�����A����� ��^�KI C�}�mT/ ��E�R��� 05ZQ�% �$�W� �	�8]��LVP�^z0=�7�� �_��:��	Ms�O ��� &�?<�l�� ���a "�hi��Kȶ2� �׫��ڀ� +���C� 8�Ut�%0 �-�橢�H���Ű� `��[V](�^ �����I� ����>s L��+�V 4�Y�'\�Uf��)�}��1
?&�.r�$�gW\P4 v�<���;�e� b�]`^��IQh�J�0� �<U�Y! �]���cL�N��ra��x�L` ���ف� ��}FN���`B��U< 'l ��cam�v�7+� ��#B2���;�Võ 	[)s�܆  K��ac��4���� }	�hb+JAK>N~�1�*���9P� ��IZ]�M,�������@�
� ���*I�	 ����d�& ]�K�X�B +�G��F- ��u�D�S� �N��~�$[90�<+��� d'��_��������؀�H*l�% ���a��~��
w�`���{j �Z�B|u��I�'�(&@}�% ������N
 *�!�B8L_d�� ��� ���uz	.v�x7� R���5 ����QHI��,~���`o�� �v��G ���X ��� |-�N`:��j �!�T,i�;	�Yt �/P?�}��h��`k� ]�0�_�!� Ba�|ָ1� ki��������(�� �4Q ��n�j�� ���#�$P{%��i����Rsk�޲S-#�|� =�(�X[ ��'�Y�oZ��R �7:� 0���,� ����3S� ��]s�! )��=Y� �6o��U&� �/���Q T�����P�� ݖ��£,� nVǲ)�ѸE;�T`��h (>��?��� ��H�
y�+ k/�l ѬK�0�Y Hŀ�O��I��Ud @)����~���3 �[�EhR1 ��:�o�K��p d_���	�ʀ�B(�3��<��`d��XtS� �?@+ \���蝥t}�
��3]�#�P���0���з �ǛB�2�� �{�I�!<� �$���(�	8M����;Zt �Xrᘭ�v8c�)�� �4��\��^ ��Z��e!$��:��y# �S�31d���@n��}aZ� �L��R�yA|��;���< M>	�� zm ��2��<?�H �3�DG�i�FE`�]ǰ�?�Z�a W��� �*�	U0�9��� ��%��u� F��(w@= ���&�]V zP	��# Ǉ���O�� H��:%�� `��d��P�0 Xt��A� n|��w�����F�<��
�� �M`�Y��{�ݐD �Ε�~��� �I�S�1]*��:��K�#m���
���%�bw�V	�i���;���@=�ـ�0�ݡP �c��Xq-� �@m�"Z�� ��,�I���?u��C��U � �*�(�rt@�9K_�W���/�Zh�0�o�� v�B�� �&��L�?`��q�@��� �V�vѐ�)�(�^ ��<@:0`�3 ��TB�� G��\(���1�����H[ ����5LWZ��pe��3�� �r��iT 1�Z ��h��b=�uN�	��9L����/%h���j�Ɓ���z!u=���U�` |)�B] �؁��?�kP�����A��v�� b��)�Id1��� (͋*��K�D�?Ђ�]�[_!���e�Q(q��� �#�%F��� ۋX�0���(L��/��, ��Ӷ��0� x�\1� <& r�9��˄RV2�	��` :� N����|�B��P����;� ��	�H!��]��#�\�&�X un}= ���-�� %Q�*tC ����3�w�  ط'&�r �W��D1�܂@S��ͮ���v U��
�3+ [������  Z��5y�� ��ױ���ӢtsT ��-Q!
a�k�7����ա��(�A�F�ȓ� 	�5}��ei\w� W{��p+����?��0�1����t��! ���j�:� <��Z�, ��9L�� �ݺ���I>�����w�z ���?��A y�!ѫ� ����Յj p��V�����AL��p��� ��@� 0�mB�?ɒpb�)�@�](�Ę��  �_N� ��,&��bT=��l$R� �'�~ݢ� ��A_p�����%�j����Q�P[�Q ���t!X�� ��u�_D�����;���>>���Q��� �T�R*+�?0�°$J�H iI��nƒ�ް��`J�3��'�Ĉ� ��Do����� �)��b��� �����h-VqF �x²��J  ��qk���� h�g_�^�2�+��� ��} j����9ʩ��A��!`K �j�	�\�	 �p��"]������ho^���`�2 ���K�$��)�Dũ`���Z ����+����A{*��2��W� �M���\� Bouq���a Q������W�e���9pz,�� ���C��g ��	hA iqܬLa� ��ͅP#���� ^�B��V %�-��� S�7�	��� �8j%Wq_ .@Zf)� 	�[�-�O�=��� 
ŝZ~�%X�� ͵\h�;��>��>`���o� �R���~��3�X0�;�� k�U�:�� ��n{�!���a���0h8#� 0�[
ɗ ���h�D��u ��J��������	�� v/��c��� 3޽Y��� �䷸�e 7����~ ����_ LY'�)݈� ��kVH�$ ����2�u ��0P� ��3���u �$-��֎ zb�ڱ�! ��U��b;�k���5j䚘�,��2	��{����	Z��4�O� ? ݗ��RSH� �t|ů��p �K�cU�0_X� �
�Q�A�{&<)�s�`��@�� ��;�� ��s��1 �
�� ��>3_����7�9�]&�2�t,r�F� 偉=l#އA��(�0�i X������.dv� a�(�k
 	�QVW1+ ����l^`I �\HwJ!�{n�Ԉ �g/�±
ZXȀ�9��% �W�ä��� ���{��V =gN���=@�wb�^_��0\�4�u�%Q` ���Z��e��Ez���ذ��LC��1*�~A�H�x� rsR�,.:T� I��$ b��tø��K#.ǌ�,�?(X��| -r�K����,��� ��5ˢY�� (V�^D���>�7 ��h�ݣ�:�B��� �e"#�� ;V }@�Tߏ�\ k���c ��+��v*�/�꘨���S $�W�b�$[<� �C�5 -\v�����3���g 	o��]�O�b ˚Ӹ*; +G�@�� i%`�h��x���@Ǐ�� ��S��fB �]n6Kq�� ; �Nv��	��+ 	Z�>�G�T�NS�D|���d9ǁ[p�V�ܑ�� �	!/� ۾@�e�� DL��Q͌	 �4j�Ѫ@� S2ҷq
�H0� O3�X�Z^S� ����	5 "h��@屼 �0��J�(���n0\6^���:����d�. t� ��#,�2 �>���u՟:B��޸@+�}�M� S�ݻ�tK��	 ��#��� ���0�o	��,�>Z#��.��)ł�h{@�0�S �x�acM�� 7�륛��3{��9� ��wk� �%Z-� Vx,���(��q1:���e�� ��]f|!� �1�S�/ �O�c�ٓL��[��j����z�h��� $��s^#�� ��q��%&!�C m@�]V� ��.�#[� k��D�XG.ʊ�8 n��l� ��$4�6 ���A�����0�	��P��<ݫ+*�ǻ`� �o��('�\|� l�.0Y`��h^i���J;=� ��0���Q ��:R)�w�\�o�^�%�#Z�? V��`~-�����������.��� �� �Z] ������Ip�[^��`ޢ �����$�d�g >e��]���$ʁ� 难�}�sa�Q)�u��PM� J	+Dy��B 5Q�֯c"� K�G	�n&�� x�i�Y�h�>�������� �� �2 ����w�� ��'0	&��2I��~@K�N/�E �`�O��	 �b|��y lT��=�t2��&WQ���ۭ�I��pv��` ����*� Ǵw\"�} 0)��㍐�bT�] ԱrhU8����4Ы��M��	e�B��U����dCF�1M���/��� �?��mA�P���x� �)�4i�� �+b��E�,�� '�^����DX� ��]ɣA%|x�� $���B &�2�"U������}L�� *������ �n$)Vl�J6�ī�Wg2���XR��k>aW��,��ZV=���k�w<A����" Ty/�v�0�}� ��ͅ�� |���P��&/��0�y��׸�( �����! �����[C}� �>Ov,8���>A���:��*��ۉYT��c4��߱	h/�+����8 q_p���B"��`�k�L \�%�D� ���Z���y^�sQ��zM�`;>ӝOp�[���� ����h���N� ʓ���� Ӭ)�R��
�1*� s/��h �e_<�p1 X¡���~ �6����zi ��H�	�Q�Ϧ�3T�t��@ kX_\UP���|� ��WS ӽ{�[�&�4y0 ��̀J"� bM+��� $�!�]�: ��@MӁ���J���ت� 9�:A`�j R�ۯ��_�
CG�o� ����� �hb�_�� �q�V�� � L��P�	���V� 傖� ���3���P��H�� �0X�?���iĊKI��" �'v�ug�� GW��Dh* �o�'!��� ^_�J��� C�y%�8o Q���"�z��	��W| &�\d~,%� ���K��{��H׀��V��LE����N�5S���|S �X0�!U��A�s¸�-`�� h�&/�y ����^K m8��O�[�PH�#@@� V8�
��� =R��^3 ƒ�_���  ��"'-�0 Zh�cL��=�t�U �N����$ �v�B��h<-+!J�CԯG X��À�jypN֮�9���K �b/�R ����~ �Q� �δHK�><1pb) �c���
�~C�k!�"��oA�dI �z��� �h;��� U�/S}+�� ���0���=����� ����!q� b��ؗ�J	�������� ��/~�\^������2�[�Q��x�t ����	�#S!�@����> �oY�d\ �(�*H�iF5s�x�`K ��3钑�� ޿��]<n &�oz,�� ��|�[�� V�W+ݿ �x8gi�L�P<H�Pꣾ N��|'��P͇���a�1b%p3z>� 𻄪d���bP��/�IC�� �Wp7*�F�K��� �"��_�E���t�n�}vH�r ��(���\=b1
���B��F����i��u{ �XA<�>L� �:0@�Ђ ����1y
�\�=�@�fQ��1KĨ� 0�|h ��1���	 �����Y~��KдpC<�[�<(�,-L߿/PI���Q!���tؑ=�s$�آ� �ݻ�+��
�j�w� �$�N�y�����4)} �GX(�R��	� 8����� �u���7R� �Ժ(K�/x' ��I<��h[r����P�����>]�p�Yx�;ߐ| V��*�T�� ��3e��X��`6�� ����z�ݦ&6�d� �����'� �z([��c� �<uԢX� ���P�h~
�����M�|p� �����ׅ �k��R�ør��a�q������h�u��R �� ;�x�J�,id�g}@�Ɂ� ��0��� U�q�� 1�Ä2gt� ?5G
�_����J(��R ��I�E�������? ��D�����)i~��� �H���w\�| ���JSI 2[@.����\y�'XQ�&vA�Ɨ�F[ Q	���:�:�A ��m@ ��w��H�_�^ �(Si�y	{��)��2���W[���qS0	� �F���Z� 6�S���u{ ���=0� 5������;���;�dZ _#D���< ʵ'2CV�S�S{ ��!�h�G5 ��.��Q���2���y�s���  �[�L�R{�����~|/ QL�z�X� M3�J=�� n�����@�{!�0��ʻ �S��W�|� ���7�ߨ�J� �S� ��! �
YDL�E �2�h|W��b�>����E/
�Ms' %��ȊA�  ��GZЏh/^�:@�M�B�_�D����� hL;��ؓP���z���@��V�oĔ�v��S��\�J�1��~���<p� &(��Wa ����Y�Q���t/�^��$�*�R�_�}�� �,V�g�q��3��L� �渷p��J���?0��"Y ��	���?!� &02+Z�x� 3ނ_��L���E '�t�3�hz�Q�XN@�0b�#�@�h�j�����]�J �޺"��� ��կ� �*&����]N�%���%�P j����U �"k���S��G!���� t%gZ�\j� ��^�o� ��$h����P>3�y�YAy�m.�����n6�V��@�\�1�� (�qѢ�W ���� �w^@���dJ��xc���4-���� �#�;��,�+N 0�X�R �N���s���] ��j�G�m����oT��	5C;S����U~� ��Ġu�pV.��m �P��;�x /�O�.�0�:[W �X�̋ ���KG�^[��o$! �h�l�� g�.w�� �n(�� :0�h1,*Q V�����T80��0�^a Z����1� �2@K�/6�� ���j���% �!���	�.[S� >�|/�5 �˄d�� X��P���~Zny0��S��U��w�2��-
��+���n ����冠j��d�D�������b�Iױy��!��Gp�`x��� ���?���P C�#|�'`��� J�y͙�@�@A=_�P X��d�� ��bj� H߰�n pĨ&��,+ w�(���6��f����� 	���>]�u ��ߢ���� ����}�VM �PL� ���
�v2 pY)�Zh b#��O�
 �QN*��9��鬫 �°AR^|G	���@Z�� l�,�y�k� m%��o�w=	���� �`��J �4��
	) �_�G��? ��%F�: /Uq�OPa,)���B�� ��UD%Š h[�I���x-��~O���@�Mh�z{$��d�8�L� `	���h� ���\�J1{ ŭ��`�� P��C; ��:}H���1�f/����I� ��J��� ��
L��� ?���c�� ��:��e� �t��0�\ �%�?�e/ �u!�9�,[�  P�ԏ b2��/a���icI���j� n�q�F%.�� ����v� [.�,��a9��e �* H!��| ���Q�kP+� x��˅���� k��"J��\��@{� ���R�	#�^� �+�\��Udk��;K�E�����:�	��c 670y�� ���!��� Xou���u�,� ʨ�HzX!�� �bΨV��<t����b1�={|�=��Z��A �M����KiN�2�Yw ǵ��ȸU 1r�+�J�:�p ���O� ���YKâ !Ͱ��0� �x�'оU;�� Rڏ.̸��ص��eU��g^�Yoo����l 9��ʦ�	U ���8G��;3(� �a����8&h (^ѳS=X;,[�,�*����N3Z��� �` �F��-h K�u��� 0.��^� 儇	!�\R ��&�,- ǹG�D���B�����%X|� ����cIyzW� 0i�� O�!��ʖ ���	�:�cő�>0�?7��`�W酸�|� P[#�b�������B�X� v��[��U�  �\h�:N �Q��cY� ��&Kl��� ـ�
� �\����� �)�l������{�k�� rx�P({� �_��s�� �`��@u	�f�Y��p��,��]�K�HZ��^ ����P��� �}b���Y2H�`~'0@�w l����; S����H1
0{��^Q I�%�|~{� ��҉���
 8[����!���Ma� ��r$z�' ?����|��>Ћ �Rv0�� �������Z��5�G��[�Dd���!�Y�U�~� �����&��5i��7 �� � ����MHK�S�@=�^ � ��# eڮ��� ���p�b �}gq'�� MA0*�?�����)��� �]����' �"!�^�- h�Ld2�Qj��tK�%����������Ԓ��.q�� �0�3� �,���(MH%b 
����w]PձD	)�� �E��� c��y�� �� h]QZ�� A����
 V��b�H{� ���ځ�u_;���iZ�S	�[�=ք�!��4a�+��@��K ���H~ b�@���W�} �]�2`&�q�d���� �3~�>Z�H)��0�yI� ���qEa�G�߇�h�R
$*�.���m�� ��@�5? ��X"	W� h�H��'�;��_@���]���3s �Љ��1# ߤ��W� ��(���&1�u���	��� %� z0�d�����c���<*_ ��hp!�Y �b�u��	� ���y�품'�����4�~ �h
_��q m��嵇�~�@@���/�t ���W#տ�4XB�`�� �/��΋ ��Xs���C��r��t`rhS@��k��/ f�rs�� �ՋLڱ� �l\P�~����B�| Q[h�6 ;bw�I������00Z .��$? ��2>*A��I��{��	 �\w'�V� �/���&���O��V�Xh���q��a� �	��΀�_/�C�^�� ʼ��l� �j�=��0v@H��<���� B�8�� ��l&6)' L��P� ,��]R`�1�	Z�7S�8�B�����$�	1�v ���>��� �{���,�) �[ �>��W� ä�i�\�? @�X	]zB $�8����}I ����' u�cAW�� ��-���@ Z�1h��d �u�)��#@�^�] P�����U=x^�53��
���c	.���'=�[�^�	Q�� ��?�� b��UYz5a�=@����p ��!��� t�w�7���$EarJ���}4 v~�MY� /��r�{ٞ 9�a��] Y�~��N�2��@�V ������w�.7�� "Gd��mx0�| ��H@�a��:� XM]s������t� �v3ru^�\?R N�V>Ϋ!��` �@$3� ».Vg\�vG}B�߯���*��	� ���G� ��Y�V �/����f�>*��@`�^ 2�P U�gy_ڶ<h�@�TH�"�,�Á �.�wf;�����er�h��$�D����B 	�NS�Y6+�G@��!�)�+\ =�*0& �Zς[�`r8qM�U���6�L4/ R[L@�� }�1(!�Kk3�L��Z�
���f ����dR� |wF�.� 0�X��]�V����S�>�\�� ����<� Ktm����� f�:IO[����uV�i �QP�XC;Nx��f	���k��� .�X��D9 ����%tT ��pe���]OZ�� i�~)HX{0 �O�t���� yE���*� j)��X.��y_�'���ވL���k�w ��ћ���$��v���H� �N�؇�B�~JP�s��>�݅��������2s�AL�
�@�E' �����^X�b%��������z��^��(��P�͕_��Ӆ"��D������Q�O� �3��*�� 1+<��o% ���{�� �d�E]�4� � ��L}����z����������{����+e�"��@��K챖�� JS�����y� �Ӭ(�1i  �x��=X�hcK��b�"��I� V�}��HZ�[
񾦄�c"]пa��'�� Z�έ��=�"�&�剰C� t0�]�_��������K�� fI�J�<9��v ��D 0����Z�0=!H�X�2 ل"�YE �'z��2@v���[���bł�w�@
�>_����*���6� o4� 
`�� ��\Q�SK�>� �U`�@i� ^]�t1�v� J�%���D�  M�؁���� Q�ˋ�>d����~W�o>�Z �Ta@�� �:J�w=1��X��@�HjK`h=���L��� Z�w��d���28� �\X�V��f�ON��c��|L� ���N�6;����`"X�W�J/�]`�$��8�0�E�e >��{S� $������0���*âS� ��[����D3��bi`� 1�?<X��� �|0	Ekuo��@`
<�G� �/��-D,��X5��ʰ� �2XA_�,z? !�\b+���
q����;d�1��0��<������WP��X��}'��`�H�
 �B}�� ��p�h &&*+�(� �f�/J�^��H�� ��!�ha&<�m ��P>Jٌ{��p�X�I}��f����� �$����R�B(P��ЈڸC���:�� ɾK�ц4 ������ �w[���&0��!y�o� 	P�1�ﬡ�����! ��ʮ7�2 �?Ui���0;�(�� ���S�`pg��� Ή (�)r~����u�+� �N ������.�h �1
W��,�s ����v7t�� W<e��>PG 4�Nhjd� ݳ6���� >\YR�a� ���:М%	��)8 �\(&N% ��1'�]HK�`�!� hbcg	�}�z0$��<دu F�?"��]�D ��7�Ah� �C�Z� 9^���-=0PɈ	�zx� V��"�@�~� �Z��� Ĺ�@L"J׌�h'@
��n���	&�-` � ���x�� �V����0 ��!ML�� ߳$�J���K �b鍦N��x������ve �(޳'���Ȓ@��x�A���?@_�T]�!	��a)�մ	�x[:�Q������C� W�V�~�. �Pʧ���n �sY��;I^ ��*��L̨�:�D ��2 ߈�[%�.]��˷!��y�dqK|eD��Y�V -S�\ '���� �߃y�^[�\�� ������:.���? �A��� Xpy�Q+��x 2����� U��$�-�|�^�@	����x �w���N�� �:p2�㯕 ��%#6A�� /gˈ(S���!�d��%� �	)�� p��`�ӧH9d ��!NՃX�� v�G�-F ���� d�����X ��^��"�� ���S�����ء�@q��X ��U
_��܀[3�Z�/��sr�  4+�1y0 ����Y���~� ����� ���Tr�
���$`�[ZR� ��B�L1� ����Dhg fH�2 �X_��Z����ҥ��w�6�U�.�2@�8�*� �#�涽���'�~f�4�q�	�p ��9��N�s���R����� ]0;ځ��Z/%~� ��[� ��`�\�_ A�j��0� �Y3��Id%([���� @��Nk�W��0 K�+� 4�_$:�� F���WǁN� �ZK[�Sf hOGJ�0�H �����x* �����M �X��?W�	��y ����� bg.K�� ֽ%)��� �Q;3�y�"���T��1(���;� Zh�[P>���q�C����4� �~,sTR	
 ���]�)�� L�B~��� ���@= ��D���^� K_��l�:���<�vEL*� @����K d�p�C�W�h]@b�VoXL�� �>���@.P�� ��&�k %ȝ֏Z� Yh�w H$'J:Fe�	.�����xD& 3�g]Z�[�F���2�ȱ��������$]> ��CE��# ��Z^	��A
/xI@� ������R�j �!�� ��/�����# �c��87� �)MX�R #
��'[� �Q�!�(� Z���H�K�[�aF�{��� t�d�ꜲWA�;���p���^�N�,`;�" �XV��� tS�� @G�6 E%V�n�	?����0
@M�&Z?V�����`%⤂$ ��K���0�� ��oa�l� ���� ��_-3�\�SX�m$�
%!Ό�U[�O���� )ݸ$ �\���Lo� x����(�J\^X K�`��! a���g�A� ��%�;��)�X*��'���@��L�&��mT�o����C�$��b���H��WU�̽�^&z� �A�n���t% ����+W�-��� ��!�,�	�U�+��O����[01"�W���v �$ցoJ9^����	\ ��pܙ��
���/C@�	��[h gw��& �) ��-�쏔 �$V��B+�p�����f� 0�U [Yh� �>����� RXDk���4 ��h�>gS8@� �a�� Q0���(�`��"�k�̭��1˺ �nY������5�+���B �ˢ��-D� /fQ�H0�� B��3L�(-9�Ȁ�8�M���~�U�L]� 0'Sl>D!ӽ��䔟�-���*��@� \��}r?.�~��!Z�Čz ���]e ��PVa�s| �~vUTN�� �0�&J�� 1�x���y�@���$C�b��05��TyQ"� ��=O���+�VU@� ��<�K� �~�CM�-w� �,�"�\2� ILR����l�ޢ� -���ɇ�}�$�� ����ΈX�_� �C�����
���`T&� z�/~�ZBCPݮ1`���� q��-�� !Q(J�ul� L��3��H :��!�0��������P �ߨ:�� ��])Oh� ����BlI ����pM Q��	��I ���G"�  �F��k�?R�`p#�S��������� ���&�  ċ3��@[_��0�T1�n���O.;�/ `���F�	G�}䀷>�� ��T���� �3!Ly�km��#��E� �yD����R �P:۶>z!J�4�E1�q(=� ��a����� �e%^&��)�
��}� �K�V	[6�� e�����>��
Z[`k�% 4���:���e~�r`��� ��7f͚��0� ����*�@ �^V��T<' �T� 7�t;��� }#]��3�NZ�r U�/�[�h�}� 4��ˋ(X���;��]o 1%d��+�� /��~�2 ��J��wK��p:����^�| �� FY��� }�Z��� �|�[��G�j� Ĉ��� P@�+K� r����9 �XZ�1:�q=ˮ��?.L���F�%(���[	���/}��$3UL �n5����(�^i��� ���ѿ� �N���~ ?��R�4����C�`Oh��a��U��`Ȕv� W��hDӚ� ��[�ϓ�H' p�.��/� ��G��(%�±�ŐUĳ/�ˁ��L�*�%���Wq��w��u��
�h�~���N� ��$Z;��)ٺuR��ˠ�rY 3�eK6o�s� �dP�߸ 1=a�Us\<@�Pu�}	 X�
�W��U�� ��a:=�e C$"L4 ��[���p �_0�W�P� �簕J��x[���4ɠ�aM�|�D'hs$��-����ʟ BC)m ��U�9� -d*qP�Z �"��Q��� ������B ��oúi1O�Q �����%��J�\� ��!����NT�u_+�/	�t�"�%� 䨠b|�;�� 	�m*rW� ���V����{Q -����A_*�&�@�X`�? �>�������5��xI (������|�@Y�	ʀ���� �j<���r�V~���_u Ȭ�D=������ @��h ���:�1�3׷ ����@寝d~���ҁ< W*��Ƙ�-�I�Y�@rpB��X^�9A<!��������� �h^���"���@�9�|Q� l�:c��j���bY�����񴫈!� �	�����^Y��R�{�- ��W� �����R �$hYP�0� �D���ak ��i�y��� x����� ��� �7� �y��#h AX+����	�H�����-�b�� ��j���;# 	�0i�^� �]����c� R=Sh;,����9b{X>����2���kb�n"��Z�K�IOxq 
�D��� u����k�S�U@|J��
 ����(� D>�2B�3Uy69 +ʈ��ӑ� 	 fn�2h'<j9�w���^pL4D�L�>�`&�q �����.��\1 �Uec% Dw�b�<v �K��2�j�; 	��`D0�(��L�F@�B�= U�Pɐi %�]���"� 5��Y �����K)�� �a�|��	��"���L�e�/��҂:�`P5t� #���ة�S$��'��> @W�*yK����p��$qP���-L�a����e @	��!R)�X��%3p�� ����?���B7E
�@��� ��V*,?H���5��PF�w�� $�MD/� 2�u:;�RW��.�q� �ߡ
� Ǆ��䢽�p �LZ�7�� �"��� ��S.�� �_{��j�sv�������� 0��>	[��~�r�\�� ��D� H��h�6Z��w�s	1v�X$� e�ꋊ/q�1� �+�y�
h/F;-~@d�� Bv@S+�Y�)
d��^� ���S�G r�� �tLC��6���p3�X�@0Muw$ h%[0���z�5(J�)"NpY� ����D � ����� 1	������!~ ��(&��;���O�B�	������ L��#�L�>~V��s�O���[��煑P�;	P��~���:��"$�w ����
X��O����*ZY� �X2�h�Lm��=���#�� �/�-��i��r��ec�`�Xo� �nS�J:`�J��~� R�'�Ӊ�z��� |%w��\h �5ħ�x�QN�������d A�*��-� ��%��� ��J_�Z �u����Q ?�j�a�� x��.Y6� ���A�h�d 1+����C����a��;j�\r� �#e���� ǯ�,mȥy]8���i�FZA(�����n� z�P2|�@�;Z� 6��n*�x s�PB�	Ӂ �!�Z� ����S��
��� `H;��x ��'h�;�_�\�� n���$�k��B�,j���J���� d��Y*E
x� �����t� �iXh�Hkv��=�K���� С����[, ĉ+5����u� ��d�Y��>2F�GPc�K�~ih�>���7���c?Ħ[�����A� ��*�U�,F ]�B�! �LM�ʒ��� ���C�\��:d�1����|�@��T OR�a 0�')|��� }M�{�U�r��]b��s޸H�ΤN �	�������(���O Q�,��N� ��1#k�lS�-I�tаa	 Nɻ��0�z [��c�΃���)+d�����nG������D %���o�~2:�S�̀���� (��.Z��x#�1)�� 
�j(c�i: ۃ<��� L��*~�x� eS��FwA &���0cN��r9����P(j�`\�_�ݭ¿�)��z 'H����,2� *���%( ��!\�I/f vwA�6�*s� �����?�]K2�uU�ڿ" q�	$` ��n�ȫ� �����? �Fy��2)	� \l�S��# �h5ọUH �y8���A%P~�Fk�a+��C��.p	� �[�B)��� X����" ��O�!/	�+te���>���� (߳KX[t���ְ��/���  ��t �U���
����� ��􇀮bx�r	����uQ	Zɺ퀅*I#� -�X��+[~]Yg' !��� ���� �0X�� ���A���!><<&_� �÷�V	�}��^�� ��²�Φ /�z �"����Q�j(�; �	�˳� ��)�R��ZdA4*����o0ZѨ`؈X���Q���ߘ}f �~U	��0ɜl�͚��  |�	�[��<�I� ���.�Rv� �d�v&?�`i1��^��p c��!�3� �0�[2��� �Ƭ�jҞ ���`��� ��Q*C� (�[��Sw�3�K��ER+ؿ�ā�6~�̴�.J� ��X�_� ���� <%U��$ 1!�4���m 	�^�)DR���ـ6�/�>h��9�<����'�!�@%V2 ����e+����c
q� �(�K� �ۊ ��
 ��J?��� ��O�@� ��3`��]A i~���� ��(���* +��u/�� UZh�X����?��.O�Wt ,Hm@�kV R�����b� �����5 MQ�	��Kr��O ����p� �i��� �h�_�֬ ��"�U�[P �$�S�ɸ' "�Xz�ӶN ���J��� G$�����=�5�h�[�����H��P�� �-�Rʷ� oT��  1�X�3�� V�v��[h �tL�(���� �u���ъ3@������^W;# �����'h��wSx_T�Q# ��`�&�����%�0�����i����� ��s�_����@��o�j�E��^� P��:���$����`�1� ��8��tz�z�&���`��#�-���'�!��S ���~�T�[ՒZ�Y�lh\�� ٕ�aQ0 D�e���"\L/`H��"�X'�`����]��������>���XR�H �!F�\~�}���| �U�ͽK� ��`�8+�,�ކ ��p�� �0�k��f�;�v�Ck����`�@5��	�-���X`$Д	�u�4�D���8�m�ah��)�R�y�($�d����&�� q0�[��� �~^g��e =�-��� �X��V��g L}�z�,���*�� ������5�	s���e� >� E�C�����@��.t�� ���I�� �rޖ��\}�K��3�0B� J�ǂ� �m���QC ������o�4�0A���E8� ��: 1TNM� (�	a��e|�nE�
�����X*��� ���@��Ԩ$��{��p��$A؈��<���O\�P�x���͏�;/QA\����6��	�
���a���V	��j�t��%�����btO���D!�} ��R��C��j� ���B �\O<�.� [�si�H�wn f^a��l,/)� �p(�1 »�rm���ы)#:�Y��Z'V(}��n- ôr��ٍ �(�b'Bn\�x�� ��P��?� _�y�`��/\�a{Qn T�� ���5�;� ��X0�JP U��b�]�BLQ �o$��?�h8�-K�`i`^@�@1�
�+�e���`�,�� o���B��{�_Q% ������wS~ 31�XGf����;Ȫ'�>�����RE� Z�Y�H��� P��	�� S�C��bF��GN��"n
 B�1�_�[ h��5�� ����z�DX� 0�)�U��  ꪤo�X ��D�W p���� >�YZ	1}]��!����v��'�^TGl$�#�e�Vʜ O}z����%�\@� �����U	 �!�/]g?�9��� ���`R��A3�Yߐh(y�� Nvq��� �n�K��h�2�DY���pJE� �'t ��� ��<�R0������@��m�34 	<�a� �@ �+��A� �=>0��H,� | ����р ,�9�&�(	q��"O@�bL�u! �#Ǻs�{	`�h6@��H���Ef@��3����!xY��	 ����RA� Q���P�0' �h��U2 �L�&��� .�	ZfR�K�O dH����Οp
 �	V���6�F�f�>h�����p��c�q��S^�݀&_��|ic�V��*T؆�e�� ���& 8 ��!U0�n��	�]Ճw�� \X��/� ��B	�#���1��f���,�E	_�y@��gLp� �.a�?Z"D�-W� C�a@~�?wh�� �V�4���&TW uc~X9�禺 ��;�9� �6���P � +��'��W�۲9���?{ mhS� �>�Xņ( ��@�-�u� d��h*� ��֔�sFL�
b�����y� �l�k��\�� �;�2J� ���&�}� ��� 9��_��pa�j�0�*�0I�	܁�i��������FY
h�>�ix������ ���%���V�� �u���ik q�f:�� �1P#OY� ����:��$�пA� �X(�U��,\�@�A[�Z��� !�K���`���C0_�. �<R "����	y	��tk W�>a��|P��� ������ ���]�/ S�֚��ʧ z�a��?�2�����j�� h$�'���� Y�:�b�P��X R�c�ހ Ʊ�ٲ0*Jاɠ�5}PD���AZ�x ��'�^��.��� �!�@�1���- vN��l}P ,뾪�u�� %N�� ��W���� �7���ݰ��Sڹf�Ƞ�" �\�4F���d��s�]�PS<��݉ ��\�B|� ���<��J ��a4n� ��c/�qR�@�_��Z`����dY�]��w�К �q�'�tP�t�u��� \|�}%+� ��0��c�V ���h^&YԴ�����/ �m�8�x� K��|g����R@�h670��(J����� ׶n�q��~ aQ)YPj_���% ��&ҽ.� zl1˕`� ӿ�j%�� �wxF�˜ D!+И/�&3� X[hH$��;���� [�+� �k,��Kπ|������j I���A�_w\��+į�̭D.�� 󵖾� x� �%�
B D@�΃�2� ф)�Zň����p~�f ����S��i���>}[����b� v.й�`�  �[�/5Q ���&7XJ��������xL-�8 �@�P}X� ����U��E(�<Qˮ����%�{Z?-��j �������^7�} ���	T�杀e�B�C ���"R9 P�z���e� s�?I;x�����(� ����|��vo �7�	FL�[ ������ǐu.
�'d1�R��� �Dl��H �_i��[ I���n aL��\��Y<x��Q�� ǛXiD %.�!�m^9���GO����%�4P��9� ��2�� `�_�� �!�	�Z�I�qK�i�8
�Q� 1g��T��ʀf(���$�/� ��KA �1h�4ӳ ��Q�R�$>�	���Ǩ���A��Ԑ����9�X������ �"0}V[���@�z����(� G*�SL�oz �	�!I� ����G�,� �e)�	~ �ޥ��S<�L������- ��/+~' A඙1?>� �z��K	� ���M��c>XB� Ϳ��[� (\3��& ~�kR�� �B Б�"��F G�D�[- (�R.��E ",��u_�Q� ��B�	É�V��W�װ>���a&�Ɍ ��M�N� 9�=�h��� /w�XoY[)�������p�N
����1�����z V��,��u ~ ���� �ah�s��>ȘQ�����X�� a���V*�) ��d�!F� :r#X,	�/ �`��|�- q�s�#����� ��/I��\�' b��	*�ۀ�� T�1e�4 ���+�� V���`'� |}�4�W�� o).Pց� �܈�]��K\� ���lR&�O<�q����wn�^ �$ =�ـ%�:_ D/�k�����^� ��� ��P)�� �E�"�4� hy�T	�� #[��1w� ���_�u�B��w���g�|��	 ��U}R���.�3� �O���< W�Ҡ�#ە�0����S�	6?�t�,'����  ��S�`���@@��#(��: �
o� �"�z_bE�%���U���=���=�bq��X ���8 �*�W��M��Zi���/ �NѾϤ 4��H� �� [֛���� ��y�� gDY,�B[ ��A1P� �D~%8CS?�U9��ٵ���*{-��ʘAs�0 �LTV'�~ Ј��Z���΂N�R`6
 ��A�.� ��=1��,�p dTϹ0� �h�k�̗ X���] �! �+\Ы(j�r� Ei�/OQ5��Ʉ�� 21 `�(A Y:�Zd*�� ��[��N�x� �>h*. ;k�t��������1�L;� m�N������ :��U6� �b�G�*|k 'mȆ�&�ֹٟ���lv _q �?�1�)\ �����Ӓh� �	8� ���o� �% <�l��:�H �Җp'�.�r N/��ㅿ �o��z8�1 �\�*W�� ٶn� J�O^�:�'�Z�$��| ";_�\a* ���ł �D��1�� #	����
�c������-���	 �U�D��pW��'[��e�  �7�	R��^�� ��e� ��*N�K� >+tp����OݙFP@�$n�J�T ��Z(� /�S	�� �5�VԵ' �*3ӉA�^0�oIm &� Q�GL�M�	"� s�Xc��ꀟ���� ��2 �� 1�+�up�4��.�z� �Z\�U|7���y.�=o�`����,��� �s'W> �zm%D�&�;l^�@�P�$ �׬�2�;r� �0�!�� ��@Ֆ��WM���0��� ���Gu� 1��`�0X �E	ɸZw� h���t_���� ��Pb0 ��K��zZ��� ��o 1F� ���H"��	`D�W��/�!��� �0�X�"e����}�[��=�; �v��T� ��Z��� ���U�F> $�,-h�m�0����z�F���e�4��MO�d���X3�Ԑv��[7�y`�ւ�Y�����a\F�N��i�	!}��ғk�|�`Zʰt  ���P� +�$��>}� Bi��h@.�%��@�*f�qL OKMR�P阰~���V3� ��F$,�s^	�`z�<o*[����Y��� ��W(��� 	��hr��" �D)�2]W ��#���1t ��?2��wu��q����|� ��� �������|
]�I@t#�ؘ���{P?���V9͡�"Tŵ� HjԴ��YH P#���z��~�,�Q� �V����OH8� �X�1<�p(�`�xc �	/Fwd� �Ȝ�`���Pb~hR_����ٹ4�� L� k"���� ͇w�s� �GRTZu�/ e�����	8F� 0�\(�h� Lf���+� N����T|�A�t�(OߵX DɅ��Y��%�-�= �&�oF��+� R��j� ��I},��� �;��ι ��2�Y���	@��D: ��\R�dX��pȏ��@Y����J_ �⁰���� o��r~��f�� "@%X�� +ګ<N�'�M����S��,���+	�h2 6qӤ� ?0~x��1����_	� �Dv*��7�K��� �B>|�<9� �]�~5+ ���f��>V����;� �{$)� �ONK�<� ��-ERئ �"����M/�a �n��| 3t��� ו��)�n���d/ �X��[ �@���#D� V���tJ �	��%��p(<@G���?��ih��)�R+ ���0	�x Z� �(�=[� Ѡ0�� 3�tIa�� ����1�� �g�\�x �z/���� 
R���( Z�򙱪� aJ�k��� �]eۆ�W�9���߀#�G���� ���\^u-� ޚ�؎]. i�n/oR�B ��dpZ���b���ċ�W� ��:��J���x�,@h0.P���]����X'��@�[֮m��>B��vk (�2��j��S,# �B֠�T� �9[���*= L�3 Y��%b��r� 铩�d˷L�@��X%�0�2�N����� ����"] Hwqh8�� ��	{��0/w�X�����.�T� @*�jf9�,\� ���� m���� �3��hK(�\��L<�-�{�}hg2���`� ��,*�z��qT7ш���n��u�����EQ �oTcb��w��e�i;痂W �N � i�U��; �؉p�@B  �s�P���x�}ؙǘ ��K��͕ �Q��Z���v� 1Lk�W �7�!�4� '�[��	c I��+�L�N1��D���� }! ���:��~� �����1�ĸ� ��}XyP� n]�w�( �3�T	�a"��`pݜ��)� ��+�G �dT�� ��(n�N�=4��> ��9����st���}�� Ng1�D��Ʋ� #ȿ� ߽vh��-, 1��B��y N���:��K�^��|Wz��b����!� ��|C�@��;� 
�Փ��� w͋��/Ƶ�_ ��1�^X�] -&�U)�\��� (�O���� ���o�1�0ůrwB�x_��V���{�5� UD���ݲ V�	[W�����  ,N��V��Z����Cт�d� ����$�DS�P�N�0���� d�ŵ�2?p�9=I����7 ���[Y 0�鶢���o�� ��w!���? ��qiǬh 1�@�Q�\wR%�t�?��|(-���9�� ��寏f��RL��^D'�Q��u�[� �Z��[�-v��R��a�)�� ]�/�V}h IZKH�B�wȸ 	�1�Y� �T^��N�s���%��d!/K��� ������f R�ô�
� �Z0d� H_���:�͏!>~ 3X(��|� M�_vO�b% ր��h�Q� ��Ϛ&����� �OG��/]VP�%�Ch�,��>�\�v� ��e�)��U�B��W����v@I�G	� "�����Q�\��-� v&I��O9���A�$���Q���>��	� Y2�H�n� ��%��1�M ��}O��v =�35��� N֧�s��Ɠ&��+q8 鈅�x�� D���CNu� �>�5� �\��^�R( �`�h*�.� 5�ml�S���P�K�g"H(��~���� Iv-͵�� 0�L\MFt ��u{�[P��� ��?:�� U�YfS�� �����>�� �[����D��2 �WH�"�� �R:�~v� kW0��� i����a`+&_2� �����e���G �<�]�
	�_Yި�� �.1� �7\'�)S� ʩ~u��`��i���[4U ���]h�N� I	*�W��Z9����@ ��X\*"ȕs� �d�����1YF+�IT ���"*-H@A(ۀXY���W�T�R	ٰ�{���hj�Z 5l��VBz&���J �	+Ǜ� Xwx_��=Y !��O���
�)�s�%vk �bm�W�q���������K�G �c��W ��1�y-a'>�w;�	��h��� o����29-�X��l�'� ���*���9}���%���ژ� 0|�ǹ� *釨{�@��@�� �hZ��� ��	7�� �����$[SĶ�{��(���t�<N� ����X  �~��%�S$	���US_��d��9�J�������;j� *�"#��C �2���Z�' ,}{P�����x1����?  �L�m0Pԃ*�< ����t�:u �w��rɲ<�_�Ͱ�s� ��E}�Fy+�_����H���@��/�6E[�7�0�R X�.��Y��  �:��u [j��	0{& ��_I�� ������V� �XP�&h�����Q��LU������'v ڤ>*�$�� 1�����u PTY)�M d��/ �VΕ���ذ�0���� '�}H�5� ���rO �Z��;.�C -�U"��w�	��R��ډ��S :	h�`!�� �H�K���� v4|>ʿ� �h���/	~TA��m| ����s��\�7�T: �wIo� >��	���] K��H��xF�����h;M���0/2Y�$4%]����b�
GQ^�����=g���!�#�[�py�N\]��' x@�U���	�$"� oO(�����ي%p�=[ x�p��b�=���N
�Q�� c�AY1�	`��� �����! ϐ'A��Rn��>�a����=҇T�@Ҙ�q 6Yh��2R�>����� 3�[��AFm�4a��~�<� �ʒ	����	w���p��ى �p��Q ��5Г��� ��޽�#����}L�&��P��� ��'���< ����R@�2 �h �Q�� �
��I�G� �S+��ć ����ܭ�� c�K�Z�9 ���(�A �Xp!�ݼR�À��Ym� ��
��� %s�������ט�� ���hܚm �p���W� 땿+i��������f%��-}u@�8�1w���i�@B&�/��A|�� s�rJ��� (�W[_	#� !�/U9�e? ��K�]$� ����^m� ���ˈ ����/D� ���wc���]��p�� �2PO�&�B GAQ �@6�
Ң�O�`��� ���A%�����m�ஔ_�H�� {��0ܲ t �9���7�F�2ɰ`�H�q�! �E���MN 5����2�&�F ָ�A�� />����I% ��xe�!
+x� ��/������2�UE������ү���	��.l*� �(��﷎T��a.�h�K���yj� �>̻	��� n|1!�&Z\7�����3(��}�.�J ~��]�2�bc����*�'��ޢ�酲W�@��� 	C�
�(��|�J� I���0ط ����z��"���������LP�����}B	`Q
�D��� ��Y�*�T p\(/�%�!�,�'���2�q��V��X��d� W�M���+~/��� a1RL ��fQ�-��� ��Z�C>W �:���dث D��ɄҠsZ�| kU�]��>C?P�D ��BW^M��� ����tǝA����D�&�AI��`�� �/\��� ~����	5 �x��B�St�h� 1р��W� ,�Dq��R��ԥ�a�m\K�$p�0`�����?�d���	��R����a ���ؽ��" ��,3=5� �CX�N�6m}�H�� `[h*K�Ԙ�z>�� 2s&� �mN��}���#i~��[ e�)��B ֔O��]�<(��}k|V���� l��,ۅ�ؚ[2�\��y�@� 
��R� �_>�Ü` j��HP Y��J �\A���) �2!�eX ��^�TŨ|�i!� g�[��] - �h�0y����$�&��C �h�Ŭ�����	2_�|�GlX@-B`��  J.���xX�`U�'S �����J>)j ����0� "���h|<9�;�*��˧Y�-�ȫ�l �`��F����삱ʽ�� ���D+� ^�K�[��?�H�V uF�Ǫ�X�� J�8�ے�4�.'��- �H����
,�un� e30��v ʾD���Fz� o��N�� ��.�p� �햁�1*�� ��8�RJ�>~? �*�3��������{��89 %P��[� ����ﹽ $��K-N� z0	*�I�� BL
j��v&Pn���A��f! �B�_AWo 8��.��� 첹��l�� ���31�
� iW	���� ���ͺ���}@ n8�d7�` �x3ɳ1� ���2�������[� AT6�.���`4�j(�5�1��̴� ��$N�_ Q����\ �p)0��`����ʌ�s-��X ��T�|K�� �ܹ�#�M`fj�@�+�V	�% �xhv���n;�����jK�'� � )��װ�L\'�q����g �Y2����;�� ��Ǡ�� ��7�J��´�Y-@D�� )�1�� 8w�Pa��	<��E�����)��c ��$��+zD f)���R�� h�y di uj[���_+佝���0�3����L �[�*�KZH�; �6��L Ak�	�Q1��� �e����_ X�G$��� 6����l���빙 �վ �r�s�Pv ^���2	����� L�p^� )�`�N�2 z�@Oh� �?��D3 ʘ;�i�N�H'� +/G��0�Q� 3���1�� P����� ����R%&�z���[��?���}Q����`�S�s�r 4��!�<A�nb�  ���YS,���� �� ˿x�j.��-��t< )�����s �,Y�ƘU~8R	�
��L����d�)��p�3��� X#�/h-L�D 8E ��U|��w"֠Y��fh�K���j {P�� ^|@��	��{�-_0�p��qA���@�ו�� 1�5�t�� ���@���� 	|���R(x�-�L ���DU��Vc ����	� ��W��_ ��H�|��{�vk 7�b9PhX~ ���3�G ��^��]�� �������Y3Wl����	h7�VU�@�(����� H�"�^�R��a ��s5���"���
���˃&��mU �J�%�P�v:! ���UBp ��KF	%"� ��[ҁ�M 0�hN�, ψe�@6�$_�|����ؽ�� �<��+�K,�p��I��@w�%M �S���h�{ Q��?�� /���e�13 �KY�D�2���k��l ��p��/) z,%[L{�Z �<����!@ �GH8�� T[+�^���S*ҿ�?��P!O<�4 ���H�}��@j�A�9e��Z���w�n��ص� ���uF���Ov@U��j� ��}��ۜ�H��-T�o��� �ܻ�υ���CQ���<h�����s �H�L-�	q TƔ��� � ���8	0(��x�vVk�g)a�����U�ؽ�5�����]��z� �q#��U_� Ȕ�0�[>	� ��C$�A�Hp� �u�9�ӝ�q� ��0���"/ �,GPA�
 �[XS2��Ƅ$ �}>�� 1k��+�� ��	}^� �`q YVT�=N���;�� �:�@�H4B �n�P�����ט ��a� /�)�:�-< �v��"�# 	�_���4�����T "�O^�$�
�2� ˻i�HW� �u��U��B�Ā��� 	T��o-� �� RD�� S�%����& ��Z�� ����et�  |0��w1 '%��e�� A��*�#��h}R� �Ҩ%�\��ˇ^�)y�]X} ��mb� �����(� ���0W)_q �� EQ�� 	�z���^� �eV��3 ���F|� q{�Ċ^�Ӭ W�xF �\(� ��Љ�l��Q��S e����7� �]x4���B ���QV �a�+� ֨)%���x� L�S�	� ���r�8���w@���M ���(���U �������9ҧ��A�7�3  �"}0�`� ��C�� ]��v��Ә�^
��J����z ���q� A]fgJ;�L��>\_!ZfP ֓ �̗Ũc��X��>˞���J��.)|���X9��nC{)ހ7�[
�&4_�,P�l�90�a� 	T�B ��+/��Ǜ�.��w VHOC� �h��޴�>GQ����p��Nh�&���D>��t�����r ������� ��:`z����4����0(���u?�ЈNpC� �w�P��k I��� fS�ڗ� ���ꇀ���UҀܸ��Q H�+.V觐`�ޜ,� jw*C+1 �	��� ή� ֠1�Q T5�:���� >ß����``p'e� �3/�u�k( �J�9�N ��-%غ�m *�L����@ �!��Q%%9�P] �����/���� �캢�� ��I��@2 ��c�ҶJ?P( K3�t���b������E��j����Ӑzt ֌��|= � ���� ��/��%�@k�����-��> %�nH�*&��`L��^�Ɠ�� 5�V���*��4�p�ӭ��̰ �x\9�����������Y!� �7L�P/� �=C'[� �ֈ�����s ��U��%8��� �!��;. �6�,�� �8�%YS<!�� ӿ��
� 	�I��-vb?P#�,�@�؟����Wq��E�`���� ����x_*�1��� -�ƻ� /�V-=�YX (�U��o��� ���L�'�Zn���hQg��Y�;��[��1�]Ʃ�`=�"�;�ɀ?���v �B���t�`�Y����������3�p�� @� Y(�W�yO� ��u�h&{8N��n(��%�� D�O�|]u~�Q`P׸��"-C�~܀*Z��Y ]S���� �ݵ'�h�oԋ��1@��0v�Qٔ4{H s�?��,	 [��$� �C��7� 2���j:t���i�0�'}Ж��P=!K ����ٵx ӥV���� X}e����5D�\���_<x% �V݈߀J���!�_��'P�w: 3��@���mk���ã00	�@�e@�r j�:�l5d ��/�h�q� F�;á	���᠇@)h��������(?�	ʻ-��� ��L}��x3 ��^Fr�LQP կ���� �:�9�.�! ?��X� �o��QZ���M�e )�_!��� U������� 'ڰ�1v
��u�v* [���UhL)�gE��0#����V�۾L�(A��^�R�k�|��1��[����U�<�o �����q2 �IŃ��5 ����� �3���0��ܺ r��� ���n� D�p�R��� �zMEԜ�� *�Q��, �²1�9A���vۗ���LW$�y,�.�G�>��) V4���� _1������D= � ]%#���Q� ��Hs	|� ��4�A'��B���@�z�+`�P�}������� �eHR!Z�J}#th �S�=��B ~e���Ya @�����D g���Д�p:��b��� �R��H�	�  ��o�Dw� aO�1u� ML�|�~p���-�e臷�Q*�`�(��r�H� ��B0eC �Fš�u�  ϵh5�b/��S�P)�:�y�9 �%�(47C�	ʯ� �"v� ;_���b���ha�=�������OZ`� U	�B"$��'h`+@�
�� ��m�}�� ��\U 	��q# ���,ˑ ���J� �2��R$ X����\�"%�t�|��
� �S��� ����E� ���R�n �Tk$֣�H���-��hM 9BA@��_>�(,
`��������@0� �H/<���5X"�'�0�@ -�,�u$�( M��1�'wg`�F���� �A�\��%��)_�6W��2 Z�>fBN����M@��}%,�"Y 1��]�,�� �a�.� �����:Z	 b8�.(�{� TM��� %J�����ۻ@����p� =$�26�A���	���E B&��  ��1��� ��;�,�V�O�lP�c�������%���� �(�ZhTf�4��0���� ݻǓS	_Ѹ@�#��x )!s"+���۸�a? ���d��% �W)4�h t�+fr]� ��3Kۼ�� ��(��x\�� ��B"��yؿ$� Q��t 	�n�����ǌ�(�w�-tg�W4�~Ф2� �_�X-� Y���Z+ �xh���oȰ�q��RL �|%�T��. �a;�V3 꾠F?�m �`w4�O�X�i`~^� �*���3_ I�Y��< �w�]Rj��+���Z�� W�E��.�Xc�$<������U]��!�ýY4��[D +��^�z ��	���{� ��8JQ�� ��p�*���
�>�˶ �1u���P[�h ��_wˍ  ��H��R.Y�Q}3�г��_w� �۰b�)N ��p
�E��B�c�@y�� C�o�:���	 $�/���G� %}�l��	?뼀�!�+�] �ﳽ`�'��\~o*��0��;��H�M�@Sw#Eo ��24^ ȡ��Yu� h���� .2�<߭� r����=>@�(x`0X�҃��`=�� 	ŋP� ���ف�@� ��G'_j��,�?8t�ɧJA�� �0�X1�^�� �h=Zo"�R>裟������#�� t��X��H}x �Y�	�P �yV����/��3�D��Q�j������~�DM��\pVpޗ|�I�(��1� ;�$��S �"������ Q�n�oy�4����Qb��\�g��,z�G �1
Y>F co�@�]'m �(%Q��� [��>�#��L����*����H�� _{fh *�0]��[,T�= !	�3Y %�����k��w�^��� �v� ���'��7�y(z>� �fq0�Z R�rpe�Y� �����: ������LF�����,�Ր� 	��4D� ��ġ�>��� =1��tN�v�f�/L�'�P�,��|IF�`��� �&����(���;״e����	Y����|���&��d���P]�� �������p5H�g��z�$s0 @�"�^�~�����H�� �[	��� � ��52�h�a�D����VK訇2,�Bi��_�ȳ�Z~�M`�d�a� �C���v> ���
�R�P�� 1@q)�>Y( �V
��Z ���Dm���:�� x���Ɏ8����\hC
 Z%YPѬ�$ ����ϫE� �މ��` ��p�}�^��U/� � ��y��r�&��'���� lK
��A.�2>���0 	EX�`�/��rH�� �s�Gʙ�i�@O ����@[�u ~?R�GP!�{Z ���� ���&��P" �~�b3�H��
R��(��5� ڪ��	� �g��N��:J� +A�>U 0����%�`��ܿIwB��;)"��� �,R�@Z�<�ܓ� j��s%�W �b���1�t)�Ǌ����t�(U�J��es���N�������%3����` U�ɿx �5+�1W|3�� ._B��ZȰ$ �S	z!�  �`��,Q K�F��@	q� e�{�^��|�S�j��S��= �������� ]���k�";��S��N &)�7Y@���߀�$� IH-��� a�yS!5  ��/�ZX�� q�t��߸� AR#�&.��# <�}߶H (A%`F�d� *L�^��H� �Q����}��P݋\0 � W��U����� �ߏS�2����"ӂ�x	�V�0 �Z��z ��>ͬ|`� 	0��#�X �і��Z ��+R(� nN<�K¾A?�f��� ���ȑ\�� �{0���, ��X�N��i�}�@�'f�P�[��!È�\ � ��~+ȁ ʲ��{T�� )H����P���3��<��9��6X`�{!WP�?�Y0�>4� �\/���6d��>Q���� �~#��% ���(�AX��./� �3�	29X[���;������ �U�O` ���_��}� �7����� �N��$� �	 �S����y�x�UO�"\�-?s Wӯlb���P�@L�i0"��Y
�xd�h_8���	i �Z��4�Qc�3�|�B^ܐ ������ �
���'],i��F�`� �k|���'�c�B�����.�&�CVO0 �ҾDY� ��)� �Hjg���� Y�k\��� �	�r�p:�O������i8��ݜ+��� 'X�� (�;�K�^[�I�!1�B<B ��@bŮJPk�`��r�� 	'5M@��) _��a�K��OX�t��|mfS��
 �����V ���'�mw "A��2$� �H�`��C�����+Qaam��=,X����[#�� ��Z�Mw� ����Ue!�T�V��`�8�_�� ][��S�ː�&� @/34\~ ���5Jt�9�1������:&������� [��@� w5-,���; ��3O�� D�% t�am�� e��]� 0YH	?� N��-j��P��~���|�F �ل`�-�SX5�`GF�l �nA�8��hF "�~.���u u��B�;q�0�'$��Ш� ���{�~�� Ƴ����zU C������ A���P�-� Y�
 �s�9 ��=5L�K ~�p?��� �%�W-g�~�&����P8� BH��3ˋ�� a�Ģ���ƭ�3� �^�5l�I�B T-1����x� �|X�@J ����� �OH�)�M ���B>\� h��D( ��d@V]� iU)1�pc �-���4�� �mߐ�'� �H��Z�\�o�
E/'���I@� ����.+��1����i��� q�&�"љA��v��U��z� �˶�EW8��� Z����3��a�����D !c,�K�\���ݰ5+ ʞ.Sq�� �B��}v|{�\O������H�x �V�8�ZJ �̃�Xֺ 2	U��zF{5 �)��� QMk �ٹ� :�AvU�5� ��� �P�&��U���� �yq�.�-�85 P1���A�7��B�8Z`d0x�tS� B��䐋 �i�5�r ��L%�(x��� HT�2K���* �aYSL��(0�L\^:�{%��P��[/ �A�K��? ��ZE����	����u��3�Wq o��;iP�Um��w��:���|��LB ��R�q?�[.�U �!�'1���� �[Q�� �0*�\���Iy�z��1k>{ h3��g \����W� ���	؊ X�ON�J� �����Ҹ	|3^�`O���j �����B	ḉ��'@4H,��J�p�@���O���	=�y�|� Qa��N��� �"v<�)��ľ����NQ��_, ���ݖ�)�� ���P�䃒9�/ \�b-"�t $� ڂ�C� Q��0�ȓy� �I/1"��4 ���aV�F��_�D�~�SC�c⽜�J`X� *]�H��)�� �R��`�-q<�	ź^G���� �OY2# i�B�*�>v� �Q�۝_�t ��x`�Z� �%��Y^ ����_t�IZ ��]�Y� ��;&#~p�:�0�1��0�3 ��WN����]~ \����:�����`J
&�R| p�T���?@N�3v��s�# ޫn ��5�J&H�;w�ba @zk�) 
�U�����4 �g�߉.v�2����e왨>P :�����*�Y��H���4�� &�oh �Q�ـ� ��:����O�w��E�����Te	ְ���v��/�^ ��fi��u"����V%��	���~��ֿ�� I�^�"t9Ua���]ā
�3���`뵟�$��& �%�'Bg߶ E4Z[���dp<� jϵ��餀ĂI��_ k����B ����0FJx�!��y�~7��p H	
g�Y U�sG��� f�<���
 !�%C#�� ���A�� �[�,~�H��9�A����`�� �P6F��� ��0/BOvq ��X�Y9�HKq�(��0��8.)�_���0���Ob��w�#�`k�� ���jn��-^��" �تS/ ���A&�"�n���Zp�*m�>TF�/Ⱦ�p�� ċ�i�w�}'_�~���ࡢ�� (Z�E^0� �4��{�U� 5��(��W  �+���"`[���� 3�Z�|��; �nJ��� PM�fR2� ^�<c>�z/� �ͺ ��B�#��"W7� >�y�p9J5���,Lc �>�� ű�B��3�|� Z��a�
� ��#)�0�vX� ;M.��g"x� i��U�������%��@K�� �ǀ0�h�� #1�_�������J|���gZ �'-�`�}#u�_�������	 ��x��� Q�&'}�� 1�Y���cZ(��'$\> �s"��Nt �ͧ!ˠ�ƕ�
,��A (SY�/��v?��2��H � 跚*�(�zh������ nN_0J����-k ��ۨ$ �f�z�k�B�_&~��b�R +[��;Ԗ �v����� �
5:�(�h�v�`�m�/�:��@�����<�p%��U�f� ᕉ�n�;�Tu )ؙ���� X[Y��ͣ� =^+�y���QjI��� �%��������� c �Z
���!W;���&�q ~���}
� ���)�^� �jSAI�q+l�-��{�]9���Ѐ�7RS ��gd��� ����-���h?t�#��� ��	A��8� P��+�� �*K��[� ��k��C��}&l����7@8Ih ���
 ܭ� ���� ֈ#�(�� �'��	���4��Mc����(?��H�� �Q�|��,* ��	��VP� �D��U! \GS�#N)�����	��V� ���4��! ���]�( 	 ���N�#�͜8��& A�[�+��� u�着�8`	��B�0�� U�	�T��]1^��
�������<��HZ�i+����}� �Q���� �~�Eܿ ����UA �����i\�l>� �x���.4�%���A�8?o�-\H��';�,�����< ���3�8u&P�� ��{O�9�A��4�@�`��D�yx|� ��a� ����P�� ���N�1� �3�A��;�Z��Q� ~�����I�>��� FP�N��	��h�����k=[��,G$z����0 �X)��h��PW�� z�\S�p-�t�DI�+J�ap܄ ��/��S��H�b��M P���Q�/�_��� 0�+'�� �p��l��(ۋ�"�Z��@z� ��'ϘT� �.�D�EC����M� ����A+ìw#Խ] ?���g�l �C���� �ĀcW&Z! ��ƺ��z| 7��m@)�.�� ¨W�:�	�px�_`�b�V����N/�]ԯ,�	�|��9��聴`�>�Ӻ�� ��	2Z E�'~9�K Q���� o
��N�Ck+�b�RȽh %t��4 \, �X��� ^n%�~�a�_g1 ���c� ���9�����S�Z������	��WQck�2��.*��� U�ʂ��/b�T���	q���'U �&.�bR�W�9B��!���y pN����� ��Tm[��0 �2��S i��J	�! A�N����� 3�݁�\T��J��h�D��>�f�1��Z_ͫuP`E@~]0f
"�%������� �d��w�y:��Ix&���ci�H�T��!L�_�m@�J�$Ğ:�������� ��3��碎��s���� ��)н�� *��h�n�u�}w��� Sac�#p �����7� H���ZY�2|� ��y�� >�j�t^� �v?ZX�� �{,��r�!�}`.OL(��mx���H�z% ~�X�h'�I8�+��Ń@�f�� ��>������ �����*@ M���Q� ����k� ���yN0���2��+��=P~/ ��'i���y>����}�!G�0���  :�LX�.�� *6���l\� �����ߋ�_b0@�Y+��q[X�:�z��ɫ�_*� �1�� [(�C�7�w ��}��Z]H$kAv ��-5�h,��`�=6CT ���Y0��� �\���8���p�e�D���=ɟ)���b�r�<'[��@�#��Vt��ा� �����K��� �$��/�ƀJ3� ���`��0G��逭�%� �LfK��]B ��Ѱ?��,����ޓ�� N�h�1 %�#v�)Z ��� (�X!�l�^h�f\����@%!Z���:��J�f��� h�L5$ϱ� �]��!m�?l�^-���y��|X[Z�ڟV���9	լ 0� �\h�B$qO�����l;(� �5��K��`4µC�&烹��Y _�����d�� �{h�p P��ZKR�' �o0.�F% �&
�]	��f���I@�}0�  េ�o�� j��O��<���i?��A�1�)�u a?��\�Q� B6���� D�|�T��1�,�@���+?\<�P���� ]�hXp�2 �R\���i�7 Y�&�)fVHG �@�"��w�d5�L�����OB���;␹�!Z�� eP�4>�� ����� d�1(\奈 ��2D�K ��� մ�}J�  ��h��b� �Ջޭ8� ���(�[�� �3gukM
 V~�o��?�� z��+	�t R:"O��|E 1�X�G����-���K������薜��9dG�0RU�� �|��S���q	��2��Y���� �aNn��� �p�,�Z�*�$ ���\��C ��V��� �(髕q� W�H=���?#�_�2���.� G��������r*s\���M��P�� 8�[P�(���l"/�`\��@p 0|���ӎ��18É����&v ^�7��h �Sx��� ��^���R� ���rU'�%5���b�����C$�����m�����[`r��d-��� ��m$ �C��	����F{���`�uP΁�C�w�瀞K�4ą�Ni���p
� �7IJ�81\����&V��R�@_�������B�A�E�6�Q<��>��i���ϐ����h�^��>�09A�!zEPp��'� (����e ����gW �U�7�M��>\� 1�]h2)��,�� �1u��k����r�� �8�.4�(%<�U�ɀ�J��}3*�1���ɺ���Z���4��'
�	�d���Gޟ@��4�^I ��x�_���pa鐰��i\�	z��`��� ��G�$f@9 ٴ�S��5  ��8r����9(���`�d	�H� @�a���W�(0[�;)>���N
���Q]1���/� ��-�"	��:!�ߊ����;1�$#0T� ���.�Ľ ���,x �� A~3��[���y ΍k�� �n����琫�S÷w�f�' Q1չܑ )�4?Y,5�-@���š%��w��X*���7��F�Z �P�N @)� S��0��� G���$Y�W> c����/� U���#����� �X~�(<8۸�w� �_[�� ��	0�^G�>���\�_|`�& ����L�VN ��>S7U[� T!�j;)ی:�K��P<�I,[�S(�`���&�L�T ,z=bŰ� �FN�/�Z ���^ ��L-�[�8w��~�Y�bи� �s�;� �2�$q�N ` RS�+,=�� �[颵	{^��� ���3/ �ۡh�y5b��靋�Oº�_�i �&p��Ț� ����n� 5�)�}Y�	�w^���p~�� iP��-�U��G�`!V�X\�ڨiw�()�� ] ��R �a��_~�8�������r�� ���*[h� <�3+���� PʕǷ��. ���1�Kņ�����yt� {����� ��ҍ�\� �y�;B����� Í�����x� ����#_ �E�.��t�~ �*q��$� �b��V�� D�ǉ�Ԇ� %�cb"X 2�im��G ֙���H	^�?n��]#[�X�9 �P�׸�\o@(`��IXP�� -b�	�Q9y��Ar�1� �U T�w�����d Z���R�r� ᐆP�Q�\Z� ��� �f�P���\HK �h�+W����J��^� ���0r�; Q�s��Z~  U��9�w :]����o ��FXZW�zGϬ� p7%@s�Ȝ�&P�e����2��s(L��C���� �w��h>�� �3S��Qq*�R����r� �P�z5� �M�����%�c-��O�B*���������l��^��x����W<H��R��� �ے�Ə� �%+2��\��� �S.� ����O /�ذ�fA�d��ŀ��X .�k�(�� �z	R�B@�,�u� �^�&�� ���W� � �V�I��+ �B��=ѭq���U S�ԇ\� ����G�>c� �s�}d� Z�)x>�P	�� _t��Z[� +�HA�U�e%��.�)�� >	_��Q�&.�� �5�ۭ�u;+�bG���v���Y�؃� -�'�����t�&9�b�(} ��,=<.� ���1��+ -��^�v )�
�ڐ X �h]Қ�f~��a��*� wb�B\u�- J�:�}��� �~�	L�#�N�'�ƿ G��)t�[�LaX ��T���S�!?3��Ov��>�� 5��C�� �	^��|�P ���_��Lr! �lRq�@�����t���Z�n \A�Ѹ��9~���.��ֱ8�" d+�@=�� ���V
�^ 0�ţ�vXPL?� �k2���|t*���en� ��������,(��$LA��P�:��d3�?$c	N��0�B�P�~�.�s������_�!��^�/�����ܠ������( 	���� xl�ڝU �V��?� �gX��0;9�� '��� P�D�S4���΀���߸G `�<:���\?����5�F�|{ɺ�� dX�����D �2;	�[_ ���'3	�Z�w�-cP�"��k#ω�.�[� �9ʯ�� |a3�1�Y0 �tS�Z�_X<V�ླ���"�x� �#�$�R�P hbpZ�B W�-��_�/ tI%�32�[���
O_	�,��� ���䉤}������Z0�_�[;S���].�	�� �*� �IB�+�%� ���'=vc �KF	 ��R#� ���d'��S,!��A�7�����z�q�~��C�4�	��PZ��$	��T^�a �\��R��F ����"��$�	�#�Z�  �İ�h�j� �&-��/0 �~�*�� �UZR7�e���V+��-�����L~�~$�����Y�e/R����L8���n�
@��,�&`��N!>0\�a� �_��/�d������ Y���� h�S��-( ���p0�$$�^� +%�(�'��b?/ݣ�����g� �6T�p��f�o0a�����3=��� ����2v_��/�)�,�^� ɿ�~���@����JO2��ݤ�}�p��VQ����?�Ԫ����=�(�Sa��\I� + �u~8�X�0Y�ah VI-7%�/� �P>����h�\p9r� �g1�ⵏ;Щ�G��}� )���'��t @��iyɭ�@�������T$RW30�|� �gʧ-i�9 ����"P ��NO��s��'� ��I�� �`�q��%	���l���j���$K ��Q1 -�Y�R(Ɖ �i/��hx\�P�Y�� @04��b��x~ �
+�h�9�π��"�=��}� !�
��� ���:��iB��� h�NA�)�\H= ���`:�ܽ� 8���qFG,Z� �d��]��|�O�8@r ���͖-�d�T�B����� G��L�4>��б�c���g�$S4��.�7) 1
��eQ �:xJ	�^ !��}#�L �8��� ����0� �X���@� �h%�M��) ߮ �W	� T_1��su@ �)�#,�^W���yZ ���1� �}���oa0 E��*��㸿 �xb~p�� e:�y9�����X����b{A 1�_qR��Z �����Ec���>: �_h� Zq^�5�����X�� ��=��
����w0@�k&*`�( �/�2!� ��� �vP�J�@&چ Q��Vy�q �����ޗ �5:�Y�.� 7�J��L
 ��({=1 	���n�� f;���[ $����{�. �8o�J�� "@׋��^4 �|�6�]3�p v/���7Q� ��WD@� �+\��K<X;Y ������� ���dO� )z�W#���A ��@.��_,!��&��S�E �*ؑ� �z ���%���n ��۱6	�s �H�!@%� )LȚ�Y �h�a;��	�kB
`�F% ��o������� �[�$+�+ ��,�U<� ���qY! �(��,��.���� )BSU�}>K�� t�<����_0�!����Y�G����<� �M��uT� Vv�!�m�aw0�`��H\��J���֗,�M5> ����.( ɱ|WS� BV�q.{X%�� �ܑ� �
Q���H�j ��z��8z� 턝"��@���L ;�+K7�#� �ĺ����-�%Pt���N��˶B�|�V�l �UHD�"�|��z�g_����;� ��-�x�:Fy �5�P�'�iX� �6)��1	���1����6j�|���S!��p�T���V�`+�X ]KL������W¾PS��}���`�jhw�� ~v�)oF� Z�w�<����쀸h��z��ALM�I_�V�C� �2�8\]�Tp
�P4A����F"��)�>`������A� ��� �LU�1Bh���E�`TIp2�R[�� h&" �`�S�	��#!w�W`=�^Y� ��P\-�b��3	�[�'�u\�� ��hO4V� �8�1�\�E�]��[} �*��sK�h�U&������l� A��? ,�{�	�X �:2Z�Ώ y�Y �~ 8�5E`�kQK��L�3���0" �/�H� qX �A+( �V����9P=/�J���m�8�2� &���� < h�'����g �nA�� .E!�i ����%������ R�&��:�" �A(+����_3�~�х���� Gh�kׂ� }P�`��� ��!�r� ��9^� # ����3� +�v��WO��(<��-�O`/l����E��¨��� ���b�* �@C�.�
�}� xc���$|- �ƀPͪ
 .�����ĳUZ���)��-� ����׵���>���������H1��yI"��頍���r�>'x+@���7� �	I�*�� X�Gމ�	���d��,w J�;��|�j�V �*��S�� _F-p��L A������0�~��< ��u�%^��[���R)�擐 q����� �Ι��;� 3Nt�9��� ����gi� 醏�J�����`I~�'z` W*׿0�}����HU`�$�� 2JϩG� 0�n�g.
Y ���DV3٨�-�xP����JG�@H�&k�	 /�U��r��(=��\�e Ag�^����3 \k��h�) �7�;� � +����[��?Z`1-�_�.nC���~���8�� 2�X�	�\Hs �i���r b#��!Uх9�@ ���
�����8^�0��[ ��ԘiP� H�X�� 1���Љ��ܶ Y��u� ɺ�7�Z!��N������� "�n/���\ �VC��N�m}Z �	hL"Wշ��X2��y����
 �Q�/�q�%�a[i�Ip�; ���*(�y��� &jX
�<� ���g��� ��l�O@�� 6��X� �Z�����Po�0�
����YH ��'���h�0 �k���O, 1����� ����d��� �ȓ�rV(�� Y+EW���?�����I0 ߐdX:  3V�O��K&1��Q���e'�����/��c:3�w�z�'u�b�\N� �p��E�j�)�0��
��%�fAЈ���q�@��X���Q�a��`�Ζ �8��/ ���Q���>hu�'	G�D ~�Pϰ1�����@ڠ�_ h�@wj��ҹɻ)1�;�A��J ������� ͜P����?�� �Q
�[���Ǟ}��p�;�Z ��x�v 4�w�7i5 ���E����	�P ۂ�v�`ğ� �"ClL�ݓ��� �ׁ�Y��  �)N�B��� %���w ]����� ��VJ)�(	 �OA��_W w��>�zn}�4V9H�����j�࠘?�>�X�����`���D9R��\��� �ʃ����2��z
��%�,|F��<��N�z!� ħ~�K�� 
��\h% Q�[���>��Py!(G	���u��bq�I�}�?%�DG=����S� �U�΃���`è��R�%`�� F,�kV�JQZ�*���aі�� 0W[�PZV �o�챡#�;�,�"_S�L�9P8� ��X�� [�,��?� �p~2WP"������� �@^h�2�� Q`Da}d�� J��f��{ Z݇"w�D��@�1��q>`�� ykH�N�͉ �R��.#��\�= /JC���=�y ���h� B�߁�� Rz1҈�pX���]����0t$ 4�m���מX@T Akz?��`Y���Z�0�U%h��J'%���b|.�@$��=Y��*Z[+�<k�N1P��/# ���	�	[�g �*�i/���PS������r'��e�T� ����)ȫ�\c[7�p�m@�����~F����Y`� �+�֙�� ����n�uP �R'�H�* #���(�q J��Xѕ�9����$�K�p{��ʐZ%�� Y򅹠�B��
�ba�`nZ� �Ђ���J�������[2�EwW������U��a0�. >~�5_@S� �����tg:p��Ԣ! (C����� ʫ�/�r�I�h�HF�$ >�xX=p/0�Q��S���V�{���( y���;���v|_ 9³[T�F r|(Q�� }�Bk�Gss3 ^z۠(
֕�˰�� �b��/�� �� *�L� �A	�3>� �O�B+o �X�)M�� �S���.I�� :��)� Z���D��Lq� 2��*�p�0�j�� �d�|�E� ��;H���1��'#p�����?���xpg�T½.�H,����T������Q��`�.��C?�� ����S� �^��8�M ������� �"򚌞v9 �����3� H{'P��� �cJ�fh l��ѨI�:� 9zFq	�,]"�dH�� �tK�v	� Y�xa������ �����} �D��5��� (�E���j! ���B̈́s��7�
0
� 2�|��8�� 1�ZP�[f	ma���0%L4 ���i��:Ҵ ��):� �J�[��u&z/ �ikIc �b�|�'�� l�Z��B>�Pu�@J������"�@�Z�}���� .����=��A���Y�������:�q�(����9�Z-�	V�@S�k\%:��1��o �؁��7�� �/ͻ�A��T��P��Ԃ�>�� ���E k���$�	 +�hH*T&�� �_�!� ���껇�. ]|
b �}D Q�_"4��~��߀�� O�|@�G�v�x# g$��A�� _�U\���ƺ �|���[� <�ޮ�� �G,�X(�!�`����y�E��[^�(�q ]�#�\��.�� �|���s z��Z��q �^B���fd ��k\銭�S����T[: �(0� ɇ� t�buy��� �|R]_�� ^)��z�oK:�v���k��&	��I�8�J}%����\V'U(|��]!`1�`
�ڦ�� /�bL %���ͤ- z^�Ă�� 7	T�� ��u,��x �3f��� '�IC�ȹ� ���,��1	3�t/x����8;'J?�� C�h_4| ��y*�3�;+���"1)Y#�G�B��@V�� �ܔ��"�?�@�*�
hy. �L�� ����K��}#U�gi�f$�P ����*�X Z�	^3�z�<�/�÷v^� \����4��m���.�C�H� 
'�Fvg{ �32K���	��+��-��� !��I���6�49Z��0� ��R���t@��6� X�H8V��<D5 ��ު- Pmצ"K $�
�؂?�9@���Tܡu�� ��ղj��LAD �,1�*BX]�?�׹r�^"�Q� �.�N�*�e �������\a��R���Y;;���`����/ (�{��~&u� )t-�}C�D x���� ��O� ��Ű���CH�U [3� �F��Q�E�-(ˠ*Y�9 ��L۩1% ��!�/�� �]�?�(�� Ȳ�2�� �v�jy @�uY �x�3
�?O �FP�`Нh �D�dU ������9�J���F�� �	�x�K� ���J:@�`��0��j�2��wp��s�m1 �	�P�Q ϐ������c h��_(�S����0�����M`���Z�:�B~���ˀ� �m�Ĺ��<_� ��H�A Ss���Ԙ������]�S+�~��TYX��B� a���P��|��� ����/Օ���~��7���� ��rP.�*�e��ʴ����Z�^\���>���;!�1�[��	+�HN҆1X�&���`�&�h� ]ď�g�w �Y��c'C ^�X�0�(� 	��7��f ���z#�1h ���r�	 е�Ԫ� ��h2n$��Jd���1�U �v�=�w���*{� @���>B���֓�H���u�3 ���|��` g��
)�� ����@C��$!���"�A=w)�B0_�a*� �O���Q�:q��!���00�p�q����`������.��8 �ҳ�G=ɀ�)h@B!} O�l-��Kn �xX���: �,�Z��� ��	�b}� �Y�Js�I ������ ��A�Nkm��� S9^b����� �DW����!Hx �S:�B�7��@��2 #�Z �W�� ^��\S��w� 䝶i-�W�;1@�� %�^vp�>�� K}S�F�	7��8�sa��9 ��"���WVjx+`!��F �߶mi'��S����K9����z��'�Ր��i�@����X!����^+b2 �w|���S �4��� ��.P�	)�`��X������l2a�Ί
>�_�?���@ �	�X��� ��w��\(�in+!g��@�>�� �<�UB"W ��b*,��
z�����bV)N@���A�WY��h .��	��A 6Qs�j�#3��V��@Q�@ �]\��K �T��%�Ÿ <d�Ì� R����u���K�P��V *`3�P
�9(���A1ʽ�� P �I����P��������5z (+9,���P�"� 4|l	@v�:�P�����;��` �>�O��� ��q���^BPY� ��[! �|�Z2�t S���R�,A ULH�'�Zt �8��+Ţ w��M3{a����R �
�~ ����o �+��\Q�U���h�����H �ݹ �G���A ��P�J� j�@,�XI �~�`�_[��P^��2��܊�	��Ou� ���e�/�4 ���Y�� �E%F�/� C�g�b�RJ !��DLM A���񗩔 ݅������3;pM�hv?e6��P*����@�ؽ��� +����gY K&��� �\�)ʍ ^*�4P�- ����0� e��x=��l(�@FTH��%W! �0����� ���:��T ��
	� Q��iD� �=Ӂ���  �yXx�O ��P'9]	��w<��_^&iUY �6�
�]������� �U��� Y��� �`���8(�� ��TYA�X�;0���`z�)� Q3�L޽o1 �i�W�A(� �@�0N�h& �)�a��d: �*��۶�	 �ER�(qG����PwM�U$�B8L�3�,�잟SZ�@�[\�����) �!��<U��G�悑��{: e�/��|X�Z��7;�� �n�'���) �1˳@�[Z �0�-m��J�;р�#� ���&�� 5P�Lq<��� ��{�ʏV���12	�N+k�i�� ��)�p"h �d�,�	H_ �*ƫ��X y �&}q� a��<���K�܀���f��,1�F����Ѿ�b��X qH��'7@R�ɶ�Z��8вa _��\�X�� y>�! �Z���A� ����'-e L9�lp��L�>>��E��|���@��	mv W�
�� ����k�� 5b|���_V }QH�Y�B�^ LSV� GH��ق7 B)w�`-TX=$��?�V#��cпeh
�� �%�gR�b� U��.���d8�� ��S
�H8Y� z[*�!˸^���p`�� �r��	��h �"�0�ܕg�f-v�˩� 	��G p�TjQh�� '
ǝ\9��uu Z��Jb8�s ��z�"`N �� *� ����0x �|"�c �K��Z��! f��ak.x X����A~�_� 9���[Ya��>����b�2i��  R��{���H._ *��@"� �����A	 �aH��� ��o���2` ڣ�$���� jtL��[� �W�pu��/ ��˒R |'_?� YXo�c� ����F�w #�SPdڸ LI^C�y$Z [��!�Ke�.�`�*�� t� �)����j "�Im2]Fp�?z _�N�Ϋ ȋ	)��G���-������h ���ϘH�[������� ��3��[ ;���4^#�?Q%�����Ds�©`����`0� �y(	ɬ9u �%��� ������3�.�&:\/����8�Hʹ ��:[0�� ����!��%.��@D��� 0��<�� ׀�Z��� �����R���j�K ��*C�L�: ���"W�i ~�h�I�J�\�p�7R��b�i�`.'&�S����¥���U +ʽ����0\�.���k	T�  �Z��?V�`p����(5�� �Yj�X`��Hi��r� T�P���u: 1�R�0.*H;�Q �3��9��,}Bs ���4���:���!و��2WH`�� V|N�qQ~0<s�dY1"��/��F ��.�x��?� �3M�6^ H�-��}`�Z����r�p� �Y3�X�|G K@'��h:���D��� �%S���� �*�`3铃��^%��D(�W����ɦ� ./���69�u�+��,��ͳ|��}� -�] �U�kI�K«���P!�P  ð�(�� �0lὋ<�uA2�5��F � ��V:'W�[,��\}d�p� 10�p��O ��lĺ��� �Ho�� ! Rm�G��wh���j�� �!���|�� H�r�@�h� �f�ސɔo01�>�S]dp�� �e����� Њ�El��WyZ ��v��� �����X�}w � ���P� L�t�7�c �K��� ��τ�A�c� �ŃW	�^�9�5uG��@N��� �{6�c�vu am��; F�D� <^�b���� 2U��5�}�)����E��^Q�1� �~ �+)Z�
�ﴀ(X�����|� �7���l���deE���w`�D� �!P���[C ���u�Ap�� ��~KHJ�,�� ��]Q�	�X� 'ot�y3� �*!��� �_�� �	{w�; (����+��������U� ����4t��>����U��& �r��������	������TY �hxV��c �-b1@�3 �
\��xUXQ�H��M��0���:��q�' 	�hIDH.	�1U����p V؟���S/ ����Q����� ���P� a�1���-q��W#�0���t�� ��B�*VY�n� 	���� PC�W�ʋ�h�@��O��# B�˩Wm��)08�cK ��	����^̐�0�s�.�U"����E��]ܳ	O� ]�I� ��F�x��Ğ ?���p�>=�	�1� s<5�g ��� 0��.� �6�*%� i�1�~�[� ߥ�+�����UN"��ʠv�5 ��G`��	 ���՜�	�{ e A��0����!#�TZ�4�F�XP�> �0��� c=~& (�hb�%^���.�S����_ V��N�{b����&^).�����#��0��&`%VU ����� �J�I�@��:�h�(����Y@X��!�� �V���r�M �L6X%� +�qt����F ��%�A.�� �n(�W8�1���_��A́T� =+
 J��B�yS�s Q�������% ]Y>t@2Z��K�i�  8d-��|eQ�:BY�U�C��;���8	�<@��
��0׉� ��v- �_�U��Ŭ �N���� K���IJO R��0��HY� �n[�� ���_Εx �P\��Iv 1���ړ a�hlZ�gC b��G���qa�?\%� 1�
�T1yB��ń��*p2��c����i�!.%R��1 �����F
 YƉh5�jk��6@������ �ڂ��[^�ŵ@�h� *�V���3 �uYZ
 S�黃NĆ 0�d%�}��#�
���� ���\��\�� e��G��`?6� �oaWt  [��Y @/�'�KD�ùV �A�`�E ���Ѥ>J+�N@ڔ����LOZ� �Q��� ���B`�M� h�yƏ#� mj ��J^ �W��$2LZu������PV~�3˽>�)���?E%�[����� �M�snߝ -f]���ݰ� K���� XSJ�i�-C <T�%:)� ��0ѨϡH#>�`:�\ R�p7�� T��eSZ� 
�t��/0 ��q>���V��kHu(0\� C1݁'�4 *���x �����: 1K(��ϣ�� !�[+� h�r�?C��rU oS��+�!�'��h0W1 y �+��Ҹ�����\jF ��b%	��� ���/� �l�=�2 �F���0�XoE)����������4 ��h�I��q ��z$��� �[�*�	�O����_`�z �'W���qA:"�_��&j� �̏��IQ�[���P�/ �=I|���L�K ���Ƶ� �h)�R뼥 ���a��U/ �"�Pu�f1H�z��|� X�I����� �q��`�1��T �rE��؀HR ��aQ��J.eA,�\K���� �y�Q��?����M��EK����O*��لrQR ��V4�!�"��_[m˼���Y ��,�1���k8��2�'�^ ��$���"��}v ��	��1<۱��K��u��5H[L ,���!,����N$+��;��� �ۺj�=H݁ )R`ο0Qt- �Б�~%�cw��#�` �0-��q ~Ah�m@��0��	�D��\� �!ҋ��,�Yd��O��� �r��J;4���� 
�MC �	���pD�L0| _U��j��.�T{ w��R�v� F���`��# [1�b����DK�<����G��v�R�� ��(>�� ����ܥ�1g��Aֵ��3P �.U^��V] ��')�~� H�����F���2�Xh/#�� ����sS_� ��%i@� &d+�4����������� x��e������ �M�! ʿp˕YXd �a����J�@ˤ�F� )d��bN�: �&��p�� Ǝ��P�� �rh�I�� Z��!x����)/G]PP�}��$�^�*`�N��X�� %h�X�>�r��A9 Q�֨�RS� (G��f��a�)�0ҽ�1߿����@�� ����%)ˍ �4?��L�8 ������ 2t��I_$dk ���ZQ{� s�{-)Y��OX\T�_�?P`�����a ;���n!�l�Z���NU�� �5~8� �9Z��(�� �� �1[Ź�ӿ@!I��� h�5K Df S��HNՄ1 �_�R�� �����O�ؓ \��	#�J� 2��c���'���!eh���* �9{�=H�~V#۾�P*�� a��L�� �^;B��\|
o$�p�=� ��ߢ)�,X=���H�����&� ��U� 0h'�9�� ��B���w�ט 5���� eo
��/WH�)���z��0p!	 p)%&�n�c l��A�{C�t� �H��
X�/ �[Q�0N�aK��&��"��\�	@W��3} Y����s�� hl]��g�8X� ��N�O3'?��wgPm!����[\P�( V1�B�=9�� {Yi��q> 2�����T瞽�h�K��� W��B�2: �Q�Xic��5��`���;V����D�ެ %�]���O���l� �~��A�� O��-����S�	���� 5�a�e�H��{ ��6ځ ����$|�ŷ� ��j�� ����A����#@4��B\ �ň��,% �P��h*_<�$ &!����� �U�w�8- #Y�j�C� ��+��S �`��Y�Kt�(�� ɀ���/ Y�:���D	&���냦?]A�:�'Ӏ��?W����CP�^[�������W��m-vK�ϐx Qɉ��{���3����50� _����� r�	#�Z� �6>�<� a���C��Y��Bhd:I@|pB AO���^�� �ރSV{oѓ����,W \W(ڀt ����u�Y3џh �j��W ~�S���J. ����`͊�x Y�Ǉ��N}R��-��Z��@�x��+ �o�,d�2�/1�4G��܍; ,Zۨ���>�v� �\'
�}!	z���G T2 ^�ĸ!�w� ��1�LU�R �	��i�l<� �'I�tE bYR@a+ʤ �B �e� ](;�)�J�}� v��N�;ʋ=���R��S *z�t�J� �|�9��� ���]� ��1X���� �hS,Z �u�բ���fχ��_p�� \���Q�t 	*�(3F��\��W�I� f�1�8� ����%� U�Ptǉ�� u�Np��RU~�Y�
�Gc�؀�Ήq �]:R��'�"� |#�!{+� ������ X��_�I n�؁�h� )�o~�F� b(O��cz�g 
�P�;���@�<	W���@�8.� �`��X�J�p ������ �Q����	��Pf�!z�q# 1�2w\S�� R�Wṷ��{�������Ճ�Dt�� ,��ƫ �-�z"�d�ꀀG�ȁ �����V[ ��ـ�
A�'%1���p"�� ��醝��P��v� QWY#�;�c J��%���*�y3 ��6Q V����"fz�'���i/0V�����$�9I�t�����ZK ������� �i	T�?� C��[q����L�W���1�"ޅC�Z�8�}��,Hz0 �Ȓ����܉� �^�m ���Q��C>�������-@>�	?�� �%� �R�ۺ9/ݰ��x����)�pXͥ �^�(��|| �5$�b��X-�u D*�����
8h&� P	۲���������_X� -�`�
ǖVb��W���u�a `켋� V�w�e�(�7Sb���> �� !]k@�ZX# �h%�s/�� ��'�ڃ(�O�X^E�@�����GR`��� �����ZY���0׽�	� Xp�J�ؕ�sM� �Ϫt��E� Q�G|)Ѻ!l%���'�o���� ؗ�P�#�` �^"��G<\x ����� ��YE�> ��|5d�4 ��Q��Ћ	 0�/���(K�� �
�P � *&i���_�P���� {X�� ��&�F��T� ^tQHˁ1t�L������ޜy �I��� i��h��*7�(� �K�E�>�����Yk��t �(ӿ\0\X@uH��5� x] ��N�xFP62B��U�u�T�t��b��$�ep�տ tZ�(� +�[�$��v ����"�w O��A����ഽS�� ��c:�I� C 5Xh�� �/\���F@?�U�h��01�u� JAr�5O�$�Y�1�u.�d B��Q�z�²@��R�7�� ��(���J���N�&����^*� �"�?���H (������t�:w�Lp�瀏3�@�	 �_!R���a��`�ܟ���� �p'{�-�{� \���P�� ���#J 'T_%~�j� �X ��- +���8�� 6��D�ƛ� @^|�
P �K�T\a�-~0�����Q;p↎�`o���Lqu{���\�ϥO@���U��X ��+��, k^�Lo�W Ȕ�!��� ��@�'> ������:���.QD� 
h�~#�V���	�^�H��x�
�U�a!�0�A�P�창o�$ ��gKY8�h�� P����q��l~�@�R� a0�P��e OKS����; ��Q�p��3����@��In��fo�&���9�{m�Ȑ]#� |���Z���I� ����*X��  ՝vq3 �0��1;� �����'u�E���� .��V	�Q��:�Z�'��hI �m�vK��z G@�R������{�Y
��)���R �1���9
t�%]2�+�|<qP X��z_��J�-�4�ZhP ̽����O}��'�!��-�`� ��$x<U 8�s�o� ��Q{A��n,+�6 @[p~V ��"��)��`Z^#���_Q T�b�)��� �kBU�pC���Ӹe���! ����f�/��uB#{��"�b*%�=�N�T����_7s>���B Q��V�Ǒ '��/�@��`Qف_)�P��� d��S�=�5>� � TL��O0�<�� �H8^)�2`�_��WmN ����^�} Q	�%���$1� ځ�>`Ĉ��)0c� Jb�k� ���x�*q�7�1��r�Ʒ 6+U�ABl�-���	x����\�o+� �� �`�M��� S#Ս� u)̈́�RQ�
Z~~�<O�f9%��B�H] ����`U����sɈ�.�� 4��f.����ΰKӹ<�N �����H� � ر�:� �%�e�&�?��p��4���:	�R�%�.w j�W�<l! �0��g�`�3��椀��[ ѳo
Ͳ�H� �)[ �� �J���p� ���}hI0��V �� 0����͈K ,�_�x	�u3 %[��V�~JƊ@��'� C�zQ�
y��� �Ui��D�� V�����+�Pɉ��p��X	k z�i�aq�ƽ��Cl��� N#��O 	 u����� ��;�'O� �����~N�r�P�`�eG �t�B�!���EP��P�	��#_� k���%� ��0�Z?q�@:;aU�%����(ҕ�e�p��mݒ"��@���q� _b���Q��� �/s�:�&�SD����� Z���%���	�k/� ���a� ���A����� �K���y� �6�
�;`�(�'��}�PHh �ժ%�
ζ ixa�~X{ T�^R����<�Ԁ����{� ��o���Y ����3>� O�h{,�����-�SP0����Xg� "�\^`Y)� J���Px�� ��4���{p��R I�s[��,����2 ��&v ��Xp��Z�dp-�!J��������W ۿI��HYN�s-@�����ʝ��@�D� n��^��Y� 20o�� �� fQ�wDv	Y����#���Z K��To
%��;�&� �H"{*h8쐁%��b2� S�\��Jp� ^����t�Su�|���X�]˅���p�B�U���/�p��HQ� %�8��^魧R�P �3u� 1���%��D U�x�o�v� VS��_*��Z���Ԝ/X֮��@�F�O��}� �#���E� *���xU��~��ܺ� o |��ŕ�5� $��h�dג����_�6�nHf@�?- gXE�y����[�,���!:  (}\ʿ�P�~�u���k �XG��O�ǘ0��_�7�1�'mv;�.�T G#��	MS3��v� z���)d	{��Ǽ��� �40��v�n|� ���<^5 �Wy`�(�V  
rі+����jy �@1�A� ��.K���$ ��t�G�+b�"W� Nc�%n�H�&� ؇F� Q�.h�Ki� �;!�2�`� ~�����4& ��Б�L i(�-��̧��Z\���t�PD(jX$��|� �4���e�������� SRŶ  ��#�xZO �g��}P�=Q%���"-��W�Å�����%�j Ϳ�҉�`�������� (1�zk��K��{�&}��?p�� �຋��Q V��^�2�"��01����k ~����" �Y�PN� ���-�'���]�`x����} ����K�,�0 m�R?�z	ށ3�OSԵr �˾t�/Ao+0�)o1���	[IU� *H��:V�� P���f��Ku�� �t�1/�V�'_��}cp~�b`��wD,�텻�� �kFt�b ��u"��!�� �X^?��Q�r _���͉�� �P(�ؓ� 
�X#�Y�[8�� ��	7C�_`�t~z �i&.��-�g�)5}I�!]��R�<_�0�,��A��׹� >K��"��Pp���&���գ��΀U��װ�8/��,���"Yy�->���.�\E �8X+�(�|�Pb�-(�0�0�#�[vx6��X 1ѥ�5� �L!���$N &^�u�� �
�h-R.�,Z� t>4"��<�L	 �-��`�x č�3�Nk� q0�wUr* �܈��� h�����+ ~�z��2=X� ��,�Q�uJ[�0 �3Mb*����g :[ͦh@_�?k~̈ )��=��f����C�`i5)��p]9�^��VU���� ЁR��
:� ���F^��z_�wL�Q=��s� �{!�ц#�~�A �ST0m� �*�k�� 3�\h{^;�&�(	 $�_�J��� 9^X���q F��(w04� ����� 	�x
\U���=s) �^RޥC�K-�P\1 UŻ' Hr ��h��.��@>� R �!��1 A��:�L ��tqY�W ����k�F���0#�� P�yL��q �)�`�@0� ��aY��� %�D����R ͑�UV/�h��$�? ��} 
!8�@$�-M <�� ���ՠ����gi[��6@��4��
�b-,>
U��G�	�]	Y��h P�.P��� �U��u��E��m�h�c	&[ŧ ���%s' Ԃ�	��� y�v���A �VaD7��t���X�� $�9�	�� �W;-��Z u%2�]d~ �$#� QRVe�+�O <�,�5�W u�	�!� �k]��r�L�u����Q
 _�K�t�2 eA�x< �X�%ѣʮ 8[B�cy��T�x��A������_�p,*$Yt� �X�	B#�� ��J愑��� �S��>����ً�#@��g��p h_t3�� B��F�7�j��� �d�wR ޺'�G���N�ݾ��|����@�	����Eo0 Ľ���q�H�8�Z"� ��3���	 �2p�~ Vl{�\�0�4v ��(j-	� ��T�n���� �\gO��Ͱ볮��$( Q���]� x��_4��HW� ��g�^$� ���_ ��X�(�׵����S��H���8�0ZH�(kv�<]� ����1���ƥX,+�;�U��P� 3�T7b� �Ug�K� */�$���[ %y�����BE�������8xk�r�A����P{0!��4J ����
�Et1 �K��wF�%�]ЈvN�!�� ��' �d������{�{y�u� T5�I1��2O�!��W�������Jې��S�����P��� -J��/�b 73N���ٿ��W��Y �RZԠ�_� ����0�S� �/��"X��#���S����b
�\~R�p-Y<����E��0� ���3�!�n}��񼰀[���U���h@��u] ���y��� ��"~��_���|!i��� �g)�0
G�:�K�7*<2� |���[/�vx��Q����( �w���1� ��U#3�`�	_;R��N�	V�J���´��^���3���Ra _��	�"Q� �f*7�:� u^\�~�[  �W��e�>q� �5�L��w�&nc{K@b��X)��We| <�VD�(c�M>��
�?�r `4�� /+��W;�2!� �&��(��;`��	��c�XS�;�,��w��9�� �R�Ⱦ3� |[ؼ�^� �-`�E׋C�eqf�{
/�7&g1 ��T`�V9b)���k�
����@�Q/"��vg�# 1�� [���J0�� ��I=.sN��,۠W�a�� �[Y�p���� "�P��(� }4�S� GF��#*�� 0Ҵ���/ c�����%�  �S��5�2�)��٨�,=�H�����1�ǂL.X� QZ�e ���i~�	�%�#��hv�5����; �� ˁ!� X��zH/5�R@�L�Y�@Z�&��~\��$�^�!�� �}R��)�,��h���0��4(�NQ, ��-��I� �lwh�䰯 �.���� #�tN�l; ���0Eˈ&�vR?�1��Xiז  ,�I� �h��M�� ��-T�� �^UQXH�u�� "���{1Q>c�t$і��� ������ke�= $0��] 
)�X��p��q���n���( :�	�P�X� �hÀR��=��&:@��/P �w���}5 n��Vo� ���#�Tu+ '�QW�07�P"�����\��� � |d� "h��:��0 ���rz� .�d�-W) O�0�Џ^;��z�U
���'1� �4|�p0G� ��{D�� �����i���y��zA:u%�s?� ��'��ؐ��������i: �1����� ۰��N�r� Z+�%��
$
�� �@kE��X��-�͎��j�� �����/ �m?�-}�w�:e������ �U�f��� �w�� � Ľ㳨I!��;�>��g�cQ b��WL��� K�0��2�$E�H��/z nC�x�ͽ� ұ����ZY� ����%� "1���g�<���N�$���X��,��N$d �`���~Z���l`�h /a�!�������&�#É �_�z�0I���=h���� �c�Z�� ��剤!������u	�9�m ����ϩ> �/�4��oRm 	����^X�!e8������ �v�Ӹk u�M��\# �v��g�|���)�k����@�� $���5'�`��!-�� ,y ��0�8��*C|G������?�`X�cZ	[�S����̄ �p.�w���X ��N�[ժ! �+��P��� M�'Eb� �_/�3� �VɵKb6 ���Z+I�d Š����<v [� 2H��Z ��J�hb���w� �_$����� �@��k�^wv Xp�R� �(B��~.J ������=�� }�����T�YǴ+	0Z�hO�� FJ�q�*��� Ҁr�c�9 �2i�
���^-�P�0�B&j�����9�x� dM+� � j��h�;��|/������� @�0�:�|�[��� P3��yZ� /4H- �xEC3�8� �0�6&$ l1Z^�z ȅ!�)��M	�}<�� ���E�@ �(cپ2`��vA�+�ɠ'y�Զ ru�Z�� N��i����.�D� �r/�P�RXZ�û���~�9?	��P �[4��rL@�O�֢��  uqٗ����	"3D� Tt֫� ��1��
� �"�E�(��`�f��- R��/��i� <�)1�.� E�K�N�Î ����
�+�I�����$�� *��'Z%� ���P.�) ������9~a�>R� ���;�<�D䣒(� �[h�EKTb�}Չʀ�#�h�zkϥ Q��~� ����"@ )��j���` �v���R��L�J��V�&!X�"`v-N,| �P��!Q� ;Mk>�5�� W:�(�� �ѕ�[Q� �R��-�] �/���	� H����#��"=
_(�U�1^� D]':�41� �[\.΃!O Ck`�5	�Jr@>����0vl������ ihW[e� HSn���}�\��i��`�B�P��:��ý^ �T$�'ʰr@{���3��-5 �pIBZ�s��
ǘA��q��_ LR�n��{� \NY�<��a ���+�����q6�"!)�� �݁���<���c�o����y����\9 ��,ٴE �Dw��) ����	����n�����~��\ل��p���%��<��Ȉ>�/�nAZ��y����g��	�"�5��0���< �w|�R\�Qu�- &!h�>a �Z�R�/wYC@5���=`h.qV ��ԈQ� ����� �`� ��U�( ��vP�u�{ �j���x�����qh�Z2�@��{�Xo( �O���[��qN"�+�>8�2�����| �� ڰ ��J$*�G��hD���i0��.)��%�#���B� ���WG�� �h�4�� ��K�1�%J ?�*����Q��P آ����$1�̺�`Qw� S�g. �}��`'l���"��������%�5�_f�@��Y,|� <��R�+�`�-��y��b�r ��UT \p2
��,J� 0�]@8�8� 3�O��� ����鲙 ���_ha;�� TB2��� �`=�a
 ��KX�C�( ��Q�� ��o\�#'� �qgb���T �S�/�~� e�=1Nq<����[����s�kJ �{�\ �G!_��� �Q3N�p
 7�� +�� ��%�Zfw�s� ��S�^	������r\м%!]���� ����H} 90���;[� �P���I�u kW�o�e�v �D-Q�A %��x��)�sL����\�0�I ��hPеe=�������: %��N�n~>_�/��^�^ hs)F�Ƀ9V��H����i-v�\^�P/��CɌ�R� _��1��vA�	�Y��Рp U�bQW��� ��_f�� )Ue4����ȊBC���VFV r��[������bĬ�� �R+��������PN�!� % �t^iy>{K*�_c0����7 �9r��� �{�0~V�t�!����J�:I��� }[�ɵ�~ �閤��  �-�V�d	 ���Q� �v���h �:%(��5�� s���<�| �/��� JU�o ��%At� ��_[] �a#.��� P��C	R;��������� K�mDOS.	8�`���v�,}}� ���h��Y�B~'ӹ����@����; C���d�x 2%���Y ��Ϥ�" �jB?�Q�K�����z2��\ ��'�퍗���X�sH_QhLq��n?��9y��ZX�� #N��" �|w ����:2 ���T��-�|B����� ���а�? \hbI%ך?�U��~ ����.�O<m��6���uL 	�\]e��58�R��*� ���1+�� �N2M�
�! ��*�k�- 7�_�j/��Ќ nz��p� �KS���� ����� �? ��ɞ{%��n��/�Ԃ�p�W����2  T����0P�u�H	l֤@����bZ۱� ��@�y���Y������<�E\�� ��������u�VCz �p��U�� �K����W��M��� �UE��� ��j��#�64;e@Z�a*�Y K(�&{@�3 ��Z۳V� �J�zW�Q �h:�.��O�+z�d��X 2�h�P��<9� W���I�B �gƝf�� X�PU`�A�2 ��]�˄ H0��K�n "���8RA��8� U
�OT�o ��%����2r�ݱN�+���]���|� R����+ 	���F��P ��C�Xt E�_MK= ����V�)��X�<��'��S�M�0���ܠ� [>�W��P {�MX_����(�0��J� !^��S�� hGD�k���N"�`��@ 0K���J�].���4�;� te�>�c���)_8�3޾�% }�l�q�a� ��i�x� 1�;�<�yV�yk���� �%Iʮ���i}[��hUXy�% F���� ��qTeS� >���
� �f�10�,�2a�>���:P��3 첐��R�-��C ͬ����3���@�k�@� ]�W�y01 ���!��p9*� f,^ؙ��R>-���	��P�L��\��^��?��-���D@T�A�;�� _��B�� R�}�m�e� ��;�]��@ 0��JZ�>|4M3ˣ�X�*� �h&7��� �W���  `-Ko�k� G?Q��|$i8H�V�P��R�~	(KX� s�]0� �Z|�"�� T�	���� ��DZ� �@��:\�-LV� ��'m� 
���J{G ��[(���#�0��HzT�z����/`���� K����q� _{'��a� 8�׹`�|r�!���K�؃ �-��"m��n��K)�h�H��.��?X ��� ��I1ظ�� t�����atq8K���B����@TZ��8� ���~�hN�� ]'P]��e UK���2#j~ ���JL�i� 	�[��P� �rT�D�p� '���nk-���`~gI9 �438�(�����!
 �/,�ų.�� |t�+�Q F�~}�^��?j��!���o��|.���a
�؂��P�g�}Y�@I�V�p(v"#8�ؗ�� w��
��� �;�Q�ض� ��D/_���`��LI8OK^���`/[� ���1SM�! �n�A՘�� _�aJ��� ���
¾O�X��9$��2���� �\�La:��$�Y����� �R�`� Q����@_�I �Rğa�+� 8����e( ��\"�4 ��$�+J�2��Z� I�W���x|�t�V���`s��>�*������QI���\P��� F��̃-D�� �=�+*�4�� �0�C�Z�\� ��I_h�*� 0��{� ��yW˛�u� 1Q��ӄ�px	 ܾ*��A� �Y�0�B(!� K��ټ)e9��`j�α �`'_H\y ��b����� ��_���)�� j]�$	��=�`/K����܀�W͒ �X��i� Mc����T�� �\��L +�.�#�� �n��א���V{�a戠���1J?һ���@����l[s�`	限HX� ����ȼ5y��%[�@\]3�����V����*) ���K����D�2�h�f�<'�߫ p0J��XZYR2̺1`���5 d� wvXu����!��Q��� ���;b�	��������� �Bi�z)��|f /��Q���[h�2�{)��R��``�� C����*z �MJ�O�s�<B�� 
�h���1� �`S�^k� /)]��� ��+��6�`5htN3X�@=�k �^��ǘ��&	_��0���d� R��S��5K��[)� !��0 �� ��J"tI��G��ө �A=��?]灛,#�����-�nY��+��W Q��@ �� �3�}��j� �D��b;�	 
2��1V Tpok@�^�L�! ƃ/���fsi *ڡ�Kj�vl �5 ,1�Y -G�֯SQw� 	�O����M� ${[_�� �~
^�� ��t����}l���[� ��b{�uԬ ��Y�%�+� ��~4� �5�� ��O)L%�Y�-UP�⹆ ��v�f���I������4_ �S=��Ƚ1�U�IǾp	��  ��+���� [Y]�P�� �Z�gxPb:�k ��8Q�?�9�	 L��BIW�^b�À����V��"�p=ې
�_ B�&�� ��Eւ �r�K��� {�wD|��8�u �;p��H� �Y��^�� g&-���uLCV R�b٠�� �R��AD ����[�a�{�{� 4��CS ���\2�� ��� �0���Յn���8 U���;��<��E����z�_� [Z�/� �J>�[�a �#���!i��>�� ���2� ��[ ��r ]�wK�頔��;0�ao.��� Ċ�~c��\Jc$S�;�� �����j��� ��Xhu� Θ���&r'���k���#��z.����<j`�i{[XW� s#5�Y�� -�D������ ��cO&��ƿ�4�`;� <p��竁)��=1����6����O3�k� -T�Z`�� k��}b�� u��0!e. �k 	����@,P�&� ��:��� ��a���H����^ ������^�2������<����~��0� biP�k^ ��o��u\���$���gY ��(��5�� <�
.���)@��w��(� H��u+$���X�!x��h� �����|?�H�`�º ���ՀA�t� sý�'(ڝ #U�X�V�N�¾Ð���6 �&K9 ���:0g۲���'>�ƀΕ�n�Uv)9��	~��%�� ���0V��[12P��� ���nR~�^	 �_&�� @!(ߗ �p�8�C�� quV*���yè��P�:8����[(����?0r�7!��9/nN%�"	 Mf}F�&Ȼ�h�i~�v@��?�%��~�ӄ�%��u:�Y h-("'@KӾf\B�� N����5`lx��0�|YS6 ����e�O���������]&nXz� �8��'U»|@B�Yf��[b�s����z�� ZS8!�_, g��J�qq� ���}Z0�4�󀁗�u! �0֋������$��a�p���*�
B�6v� ��h�J<�� ����I� E�����J
#�-��+��ts�c����,F[$ �@� �
_���3��Z��V5C$��� 1X��H�<(�� P[RbE�!��$��)
�=�T��Q[ �_�ct �ky8̵��*���y �UK���[xz ��S���� �
部�'�ք�5��#`���l� ~0�c!�H�h ��3� �7����x89��%� -����z� ��
k���^����8~ ��E_��� o��OޭZJF{V �!��� �Ch�.�� �T��3�,G 
�!𣉈� }�|7۷�~ ����A�/ s. �����5:ɉ�N~ q^�(�
�  �K%2u5 �X3��Z 7(YM��~� �%�!�h2��� ��P3�W ��UIX#�yk:��w:����	�x*L�v R�&Q� �Z���	���y�a����(���� �t��T1�\� �XÐ�J��d�C�Y���� ��+�[Q�f X��-�~�>�� +0:�_� "���/ ®�R�!�X2΃ 3�h�L��	���,?@�rW%+���b��U� V鱖�z�y �	[��8@ѶG W��C�������[����S�?� �~��*��������� �z���?�b��X��:@���g�� �|��b=���P �ɄMBC&�R ���n���p ��a�ɦ� *#�i���1 BՉ`�kQ��*��8	��-� `bӎ��6Ǔz���8Ɯ B�������VOT��N� ��ܰ'y0�� �Kմ�(V� �R��D� `��8�i|���N�@fB7� �V�a�� �+�0�� 4���Q� 
����0��! ]��a� ��f	�� ɕ����5�a���>Ȟ&��{�P�$��2��!�@�_	bJ� v}6F�Sǁ��u���[�<� ��cO7�� (�\��
�?hR�c +�*�F���р��� %��U"4�X�Y� 'H��� �RU���_�u/ ���wY^�w� 9%���U6 F|E��k,p}  ��0ie��?�;� j�a�~�|��� �E��n<�� [��2L��"�kK�����]�� �S�DR�Ϙ������+Z�{ܼ� ��#�'�
�,�' �1��;� �R�˺O!I���~.pT���,���9�` ������'��^����x��!�� �� N>�0��pQR1Ͷ��^��+E��V �R��p am���#��!: ��V��T J���n N�=���8
i� �gϐ� sA�����0� Q+�O���% @~�Y�i ��"��w�hq����p�j	�G P���� |��8jO������ �w��?�2�/����i��=���� 	V(	�R)� �0�^��3L|cE�1~�=��N��� 2.��Ƙ@ !П̡��?��~�� ��#�-� �Q:b��� Sӻ���8�&�`�鮠 ��%~Ym ��T�`��+ ���.v�)tS`�Ņ���ಀ��"jU ����p�K��+�O�`�L� �?�k��R���0���� �^���p���P��[��Y%`QC��� ����W �g���4���\�>�G� ?� @��W����h%z ۊF[�� #�	�_�p���R �]2�q!i0��T�D�0����������1P%(�{���`�L V�<!� �p4��1� �A�$���ODA|R�@�9 .�`�'1��V����W� �\���1xs�0/����r_ �Nt'T�" �p�L<�1�
�`�P��G��� ������2	����0�&�*�p��V� ���7챩\� �Q�MU�\[����� e���yN �*�#A�k'�s�< 5�]�=l -��)`�D�L�<'��g�� 6�ư�@) È�X�}����=�P�5� %0�·*bo P��q�Z��:K@,$'�!"����<�=
Ү��8 ȋX�(7ݓ䞀�>�9.��- ���t� 15�h=) D򈰼(*Ht� 0��>ͳ� ��� չkS����x��	���� t���z�t8�$\�= ��>{E@x )	�h�`^� c��!Ӂ �LH_9	A0�
�Ġ��7g��������,f KEP�`�� �u-�}���c���8|T�J����	 $RƱ[�� �/ac�Y uT]X�Pd� �Z�萤� !�:\RP� )�[�7��&�4� C�rON������ H�/p� �h@���_��X��C�~��� ���U�jz�0.@����� 2�^@_�� ���
��s pO�`Y�� �N��@ h�y0˵���&/XWCQ���� 6	0�8��\��|�� ���� ��� _� �M��9,KA�5���<��!4�Äl��iv�} ��	���f_ ��y�"�� ��h.���)ȄK1�M�e��V0���N �Dj���	*��v_郟������#v�%��i�_A�	@�M�d���0�U��+Zv�ﵰ2j I�P#�� \(�f�3<����Ob��-�w���"G�N3� Q���/� �.[��^�#�Ny4���g  Zr�$���_C��@��>1 ~G�ڽ�]�� ���W
Ŀ @�����vj��/���Px� U�*+�	 �����$3(A{���Ip� �ѻC1�Z�� �:������� ��o�ԝ堬�^ �(��Ne��;��%��F�4 ���b�X| ����� ��K���}��n �h���,������1��s�w/���Ph 0��� F�E����;@]��M�0 ��%�)� ��	H"�̑<T��?���Ż�>%=~� #8y2S(� �oLwK����A>�)�m0-� e���DQP ����:�!8kH q#�S�,�r���Y���МpR �W������ O�r)�:! K҉��� ��(���� \Z�Q_�$ ������� ���)˲ �����0F �x��A�$� ���]4 ���I�- ���0�,ď� T�FN��U��3�`w�  �'bٰ�1�{S
�0M� =�[��h�� wy!I�DR?��?�b��V}�
 (���)O� ����Xn�x�y_&�2� Кwi�0����+��^ �����j�d���maԆ� }�
�� ��S0� �/gZ�x��}���'��)0��Z� -�V^(��3�+�����~!9�� J����/R �ܚ�h�L4 ��TAaE�� ���Q&	�N )M9�P�r��_\<�2J`� �i;���f ������L� 1�Pta�h��m�5��A��˝��Q��'*S^�\+��rB1��$A��< MU
b3 �1��l�� p���G�	����(1��!�#@�Y���(�Bp��%�r� q*^.�� ��W�F؆�B=�wcRI�$([�'� Q��	��4���{Y���9i��U �<�V��w ��+��	��3"���]�6, +����1 �@U�-�un ��	XaHZ o�f<`�� �\ �4= 1O�^�t޺ Z�Y��UB��b���<���%����)���Ȧ_� �I�t���k:sh'.Ѫ�3� ��-��D{>����&Z	� .Af�S�� -��)��<Zm���e��>��8q��R ׺��m1 ǿ�Z>G������@
�\>���`!�دpV ��>�(�ٌ�,�t =��_�����a  �o� ���[��PQ�%�S�^ ���yW�,&�7 �)��v�  ����h� H��a��� X"b	᯵�Ucj� ~�+�Q ��'%k�� �"U�^ �dG�hK� �![��.�3x���*ND��:h�8\�* �I_Y� ��(�/	nDxb~z`����{h <˩��	W�	�m�l`E Έ�?��˰��e���ր"W��+<%5 P��˸�Y�� Ʃs%�� ��Abl=�� ��S$��R#�ҠJ�� ]����.�
�g�����P0 �Z�tX*� �u��cD' ��9�K����
!+ �H����`�躶�Y���ߎ��+D2|� �{$=M a鄱!�D7 �f�h\Q /(ڤ��b� !��@�� 3���Q~��Z�o&l�X-0g���zp�<�� �/�8�O�T�À�Hzf	 ҋ0��+ �Q�c���4 ���\鵮 �����L�w���� ���)Ӻ�?BQ d$`� �������a]���t`� f� Q��~U.��u� �&4��Ip)Hx� '�tY�� !]铻���	݀s/�-� ���\"�pb�< $*��
�J g]�_!�{e�\-�P�&��J��\	� ��}FSa��鹒n�U|H�w ����� *��$�'YO "��usGi }�b:@����3PS1�
"� �\hqC]L v�7�a�$P��+S�,��[� �}g����x��� �W�1�Q� ������'�����m !fc�Sz H��3K� �,�P<? �â��� ��.���#{$s� "�p��7	 �۱���6> F������ �2����q ��r )t' �ҝYjk& �Rz �NJ��ā��;�\睟 �vV�Mg�:�n �A�� �����'S �\����x���@����� H_u>��B�``�n�p���<�����5��J ����'UP���~[z �)	�E<v L�� >��N�� [es�Y +쐡�w�D �n��ڸ �@�df�:1(R�;h7<���Q�&�A �볚�i �j��XJ� O������� 9� �@'�� \�z�8�W��ir@$���|0Q.z���!2� ���]}� $�o_� � ̞.A}����` �@5r ��
��&�*s��`�Y)� ��Q� "�K��x�؀h0�� �Z� yl��?mȀ�K���%jb�+���c�\)� Z�H�� �� ��, ��z�-h>T �a���|ۋ	��Ċ �\3?޽����K����
Zj����b ����]���e>[X��lA�!����|Ϩ���T�_v���1���Lծ Yc����� �,ޜ%�� ��<�;����� ���D �}(����� ���L� �����Z2�&����{��� ��\V�U?ĺ����@���4ʆ d/��[� ����R" �	V������5�6A˵QW 1�w^�i\�}:,�̶ k�@�U[�ͷ $]"q�?W�K}�� ��vX v�I��p^�P��\VQp�\/ ��`RE~; �1_��� T�nD�,� \����!=�<�: �1Pگ5H����]��\�b ����M�*P �kK:�@�a �!�S�QX}d �	��L:� T]#ˬ! �Y�b р�Kc _� ��J��d� ��V�1��
 �^C�R,]�ˏ��ڜ�/@:nS�v��	 	����PT���f� e���d ���1H�j#%�P���a�O�@���0 �*��,>Yt�-$3� [�Qb�ZY �Ƙ|	P =�O&����_�@�B3� +�N:��� s�#�QS (��`M�^ ��/)��Pv(��:���o� Z�#��C �����"8 =����_��:��� +�)��* ��st��X \�	&���=�� ��?x[/�r��#��9#ـ����] w+�?�� �8ò~�$��� �1�� f��9X%0� �RwWJ[9� �G��3�� ����F� _�h�I[s�Xe� �Z<��J�U�C���7Y�Ǡ�	�) �-y��%�P���l~( 
˝�;�!�� ,�	h�q�>bN#@��(�jr\@Z ���o� �6X�b� <]T��������n��0 �	Z��S� ����� �p&0�~����1��7�0MԦ� �e��\�� 7�š��U rG'���� RY�P�����!G�����kȊ�c ��	�{�� h\�'^R| �%vZc�+0v2)�_JP�Ը ,�+����(�X�q�p�� �c�}�0� �@�X[#�Z�6� 3�UY ����]� ����߿ �C�кgX�	)sŀy�F:zP���e���ų ��#��_�0��	�b��d�� �~�a�D� ?\H/vJ� �f��ZU ����I�X�@�v �01����| ��}�V����=�^�߸ s���H��p	��<`M��pZ� �F��n��4X������ 7V�� <���+��M���=��� ���K���{v^�.N$�s���ʛ &],%�#D�V���ƋjF^S��.0�
I(�� �N�,� Z/}�yi U��a�Y �L��˻ �ى�:��i��&�>^��Q .��;���ߠ��y��z��\%���ġ��t����-�D(��*ЩA ELi
�!� ���%�+� (�Xc ����K�B9 u'�aR�~U������LO*N���x�. j�bHT��<S�� a.��O�\����-;��qZ@h�����w �-���  Y�	�7@�-�����q{������Qm �> �#�B�d }�ȧi��! M�������\�D Ɉ�Ɩ{ ���5h1Fs��y$`<��������0���9��J]�4 	������ �[��S��L(U�����>2��_[!�����	�# ��N�d
�J����� &�O�@�� +�^��]�_ ހ��� ��U�S� ���~ R�hb�0 3�!�J��1�+�*����. �B=��8� ]L���q�����kX� �`Z�ȕQFf)���S1�n �ck��s��:� ��e�Ɍ�/f���F�-���� '�mW��h��	�&�+� ��(C�����K [�sgW �U��HҔa#�(`:C�h� 5����KZ���c!�4Q��ӯ�Y Cd@a*�Ŗ�" �������� ������V�(���0 -�^ ����+1S ���l��/�^@ ���ː� ��,P*LP����H�������ׂ��=��Q� �V~ �^ ����Z;(�>_`�R��@�� �V��T8c U�LS��D b�Ci� ���(���
W	�& ���I�_ �m�TZ� n�0�ІU(-�	t! �~<�sz=Z6�v���Ҳ��h U5�?��� Fӊ�J��� �Z���k��K����֨�0 ����V�q|Q ��C��	�k�� -�e�ӹ �\�}:�1 ə$�;	�yR#`(�q ��kT3�|t� �ڟ"����(�8�}����!Y:� �D�%��� Rq-*�J� x�zN��r~
:���.�@�3[�A cH*�7� û�?��o�J V�$�n;�T rB��h�[��(xJ`, �|��{� ��9��kv�� p���h�� ���]� ^*��v�� ��X�;t�J �����Z ^ܗW��D� �j�V�� �{�b � ?�/!v-� ��\;R���t� �j�F2��f �)���=�� ��2���DH~
�����ѕ��̻��:�B�Ł ���!�H	"�@�8�l���#�^��| <[X(��$� 6}Z��]�>�Q��+�hE�O��«��]2&�p0h�-1c�? ����/U��x.v��"�h@>X��A���u�(����Qo�` ����6hYN 7��@���S ¤"�T�^ U~�%L�y� �ٍ7�0+�� �[ɵ>�	��}�sh[ ��4D���rH-N�pi�1 ]h#�� ���v��� ��2���}��@��X��� ��`j���Ir��&1�_ 	����ݰ �3��u ��e)�vd�C���1�.^/f&T� i����hm|��Q��	LKR��S��֦ �@(H�'l�� ��
%�&�5 q@�(��?��se���C W�Hd���.���	�C�u�� �WG��� ��L�<�0밥 ,���~]n;L	�d��Ȁd�-��[|n��jfT� �]��&�`2� ;.?1� $�I�[T(琢 @��'�o��0"��v���*h�蜭N ���PCQu� ���hU�� ��l�-#Υ�pz�NH�@�8	*?�U,r���P�@�����ͮ%b����2`�� \��@���� ���n� ��M�q$+	��D ЅH� �<�d�� .�	�*�WN �$:��, V
Ӿ|�[ ����� Q�M�-$�JҨ�| =�΍�
�x� 	���<� ���?v[!� ��n��.�� 5K���	=��� ɿ�U�D�'��9���L h����� 4Ip�X�F�	 �! ��� T�`FYh�<��Q ��3��� X�*%݀��@< �V�B�M: S�a��.,>f� d���z��h1@N���� ��ڕ4����@������Q�9���zB�-�s����'��� �Ř�Xb/Qن��}�~� ��i���?<e��;�\�T ��b� ��] �ѹ�^�� )B�ٸ�o �t!�1H�` $c�Y���L�� F�)T&^}EZ��nG �3գ(	��9m��5=��MؑK� ׏�0���3�#�"�&L.�Gp��h�H#�v ���r�S	�yfE��u5" kFa���� �Y%(��';���<�~�)���a6��r@e�� �!����	Ъ+� ���O �-�P[׉�C �ո%�J "�3X��
 K��¨ �����B�� uc���9�2�� ܢ��d�a�n>i� =�.���] �2!��c��i1�h�*I/r!��@N��b��	0��W ���`� (��x�@� ~����<N; ɷ�H�	 �����dUr� �(�,��ˋ��_.�/��-ȹ #�֐��
 �Ŏ6��� }+�D��� t�%W8=� �1�
Q� :����� E�0��J, @�4�f�*ӿ���?໥:. % ���4_s�s�1kf�)ۋ 0��d�����Z3��
I9�8�R���H �`)J��P� !Ђ�_�I ��[�3H�  �X�Z�� \Q�2�40�YdU"� ^]�:�����M �X!�* �]����;�1[����X	� �&�"C*� �մ\�� ��A�&� ��Y1�V�R _I��.0=� ��Skg�� ��B-̱2x~ �	I}u���Y�X�s��5rX�)§��0�́A������^��=1�騕���� �ƀ ����R�< 0��!�$� ��X���m�6\� 8����36 I�g�� �h����� (d��齕 ���c��  ^跬b�� �7~\-0�u�hAi����# ��r���N�<���/�p!J^�mB��)� Y�H�A*?� �ų�OUD��y�������R�	��.K��a
�/�� ��[o�[Pv� ���ޝ�,����X]��� _��x�!0H"W �85�B��SpP���3�Q�2��_� ��s��b� :B�� .j���� QTY���� \}��(��X�SZ�	�p�;]n ��i
+}������(�@���<#�wO��[_����C��[+��9��0 a h	M�` �������c��V��� ��["̘J� 8���X�V\ ������O� ����5t]� ���/zP�9�Q �s.
3<�Z %�uAFV� nb1!Ł�I x�%\U��� �;Hm$rh)�"��I�E�y[�(���`͝� Uf���v8N���c؀,�
� �[��f&�� �ɴŻ� >�nP7� '鱳���S�e:�2�@g����K0����F��� ù�~r�1����LXd��W�+���@�� �4h����5 ����o�Y�F����5���> �/��9 
ع�ş q�(��V]@��� �Ռ=T��B �^��}> ����:�H�� ����DX� m�n�#�Af!��д� ���<2� Dfy�ԟ @F��Y� �&r˳���^[; HYT�*0<>�x� ���v���X�5��ɹ�um ?��J��� �VdP��1�� [`�E��g�;��@��� �v_�*�N $����n� D��H|�.C _
��(�  ,�������Y�E��('?�� ��qpn�� �I�`ϝ�ڮ�Çt P��'����ZQ���{�U�H�� �p�RY� �)	��W 5jn�&�/:*��c���@ ���+X���u�8ޓ QP���<��~�� Zh��N�!-��_��yA ��:׌1W  +%�ZK���\Y
�@��*���� [�~?�J��9�'Z ��M	ѹ�` [S(����F�
 :��'��V;�@�K�3	��c�����.�g T�rj�� ���%D��?*��Y��ia� �:��Z2�V�R���. n�7@s�Z �]�Ȱʀ �F3*�) ��24�lC �݄p����<1N��x�8�`O���� o����$r�/��y��]�cZ0� 'R	��wr�VSfȷ�XO 塩��I��t���ג�'2�^3ֹ �R��t��8�L!��D_�'� ���uT�R� M�-�zfo �̯\� P�Ӹ�v�.��� ^S�0]?��)�� ����,d,!��.� ���^���0G��� ���-O>#�?���l����%�� �YT¢`R(޴����� W�Y��%� ��fS���,�> z��}�K� �!ӹ�k ;�<�CJ �rU��R �f�?����v�i���h�N9 ��V�#(� �ݘ�)����	����U�� '��l#�\<A۹k��1�`a� ���Ji� [��%� T�
�� XH tf��9� �.C�L p@�x:��dM����Jȹ �`�C�ڧP(��0$�F_�꟥J� �R��	� %IA�ѱ��\�_��-����w[����	�Ȃ�:��X�T�c+�{�
�(���v�BH� ��E�n��h����.��>Sn�묀;���� �z�H�����1��ȿ�	��~��hQH� �`�@_�>�-�݀<�ub6(  ��.�	�W0�X�Qh4 bD�zr�V7�HTpW����\��_p��>� GX���;��O˯��0`{W��VC���~��3	p�]�` Ԏ�梖 ��Uf��@� �3�X��A ˿2�� ����,�!�_R{&�� "��wD	�[ �n�*����L�c V(����g��<� U ��[�]��40u� �|5h{���  ����
d�)�����@���G E(�a�\�=,P�� �o �@�G��
} ���%h6t��݇Q +�@H�֘!`X	����$��� �azI����FJ��w`�� ��1��db7:e�����h�*��%��� �t5�Vɼ1���n0����/)~�:� �  3�t���5" Ǚ�Qf	N�(���(2��P���� �Ɠ��$0�щ
��+?@,6�Hs� K�O��	 �o072��ɋt%�%���� 4��.��N=7\�� 2����" )�!W��A�õ�X��a�{�����p/��p����̀�[ �c���61<�`�X���+�P%�A�f�@� �tR��^r� O�`��m �6!�R�B�Z������ �O\6��l �w���DL�w �2�{u&��]�B+�؇� ��Iى�r�V�;L���� @��PՒ$� ��J��� ' �y+��� 0���-��P�� �: ��i��{ S�Z8ċ�� 5��ۈ��  q�H_7K�� �!�^WL� iz��U��NLV�R, 攁��q�Y$����{���փ&ȣ+ �w h^<1��T�RYZ��Q�4��D� �;�0X�_ �K��v�A󉰺�@=ԏ$��������~ ����/�- ����G\ �݋+[Ah� ,�S�D�� �xb����9ڸ�]�D"p (	X_ ����9v�������8 3`fQ"�,� C<.Y�  ��XvitT �ٖ�;�a� Z�e1�� ����K�/��^���e(��- �PwX[:�'�q�`+���O�K�X\��(� � -�m�j�� R%�^�'�=X #L�Tʁ� >!�(_�� l�8�[�R��?�M�I{ �]\������$��@�R�!� �	�sc� q��'��0� ������� ����n���nw|"�2B�� :��W �!@��AK�	�Z�������?��ѽ�cE n%&���V�;�  )K���ʟb��.��f��[&�� ʏ3�d����=j���	ų�*2 �R�t�V� վc$���Pq� 0�
��/��� ���^�`4�2���� ��w�z3�V ����U��� �@N
��	p�Z�S�J�>����aB3���[ ��i����*���/`�\) �;�e��`��/��]�o�{� `�pI0 ׋F!;� ���c� �hd��z�LA	ٮ� ��!� ��Z�/�� >w �j�� J��]�p�S�3u���E��X��
Ѭf ��@��-�p�<(� L�'7p/h�ހ�:�?S ��x,��Ќ<O6�0JB��:���	G�(�2N��I�b�M���;� 0���2%��ׯ�ꬣ܈� *�r����qW��������p�  �f��1˸���m ���@;!�{ ������*�Y����p�O��R˲��
ʌmD���^��	 �"��Q%� v��Y��)} S6��b/k�mٗU � i"QD�r뚦,AuW ���i0/: �(�V �AJ5���F �/��S� ������h�H��Þ�s*�w�`��J��D����?d��e����u@Ӛ�;@k�p��[�,: )��n	3�.H� ��YM�<�Ot\���V�S�s� 0��$y��	��B
�+^��k_ w'*�Jv�:P��0à枘 SOӐ��� K��&3H ������2 �Z���;x� �<%A�����X ���E�� ������@ Ӽ!���`� �K��vSY[ %���� �\��P" �����ꍢw�w� �B�S�Q�_��0�����ҁ�d�>��_!@��*A'	 ��Ip�h�1�\J�a� ���O�� 	-�e ;) �A�����( r]�+�;# gZ�Q� �:W.4�����0 � \�?�B{C �u�qeK ����LI�a4]��/���� ܙ\�G%8���½�����H��P�0n Ab~�����	���LO?P��?^����);V �s��6� �c���� �	����?v���)���h�fzP�K@���6�+]���H�\ �`!ۺ �'�՘=����:#|�!9�2�$d�� �1��Ӷ� ���\� Cf�2sPW� ����i�.��@3ˌ\^�� R"�c����Y������� d��p �J3���!���a cN���� 37�X��� ��b���F�_�^#�t��f�� 箧D�Z)� �����p%~ ܌�y/�^V )+��P�_ �'w��Xh} ��Jz��[	 .\�1<�Z/ ��A��� �,��4 �K�^o��N 	�F��C��X��Y�@���	 ��<(� �LZ
�� ���z� �H;���01X�� [�:���], �Z�v�ԍf���y��� t�\w�a9�� J.�0g  �)b��x��� Q����\�(%� ~2(�u��! ���Zb� �݄LM�� �.���K!��� Ul?Z���	�e&����s���Rn�焥n����%��>�0�t�UV�o9h@k�e� W�n�X_~����A@�V�� X��4K ��'�l�8��� ��:1<�Y�H .;��_ �lQ�*�hX �H�ݣ�v�9}�Z�>Ӱ &� i����z� ��9$�b2 %X��+��� ��R�4 q���zj��)V���9 �˩C��&�� ��@��J�� ;���)�K ^�*a�D.�"Ȯ����n�� ��\'#�p �~��"�� y�.a'XRU ��G-Z� �@n溟�� ���Bc ��퇉sR	@/A��#��� ��n��5���!�郠-1��¤ �DW�� ����V�Zw`�\����X�J������v �y�nX`�0���C��� �Q�ɠ�����Z�����%l� �<
e_�� �d}C1��*�t�D\�E��| �V��Z4_�������?s��|�����x}!Y����F7� ����Jȕ 2_z�IF�� �6hr8C ��9�`F8����B��{ z _۪"� ����Y!�~ �O���n��\UT@x-�[Y +��/pw� "��c!� �W��KZ�m� �������� '�њA7q}	 �QD������
�$8 h��ս `9�קy%�(�&�mo��) 	
űڌ���uL�����1 � �z�) }�U,�r�+ �G3�0 #���|1 �TB	�� �kW#̤Z ܣ�ç��,<� @FN0�7���"J�� ��/&����(�8���8BE �s�/� x m6�����X �_R �ͷ�1
\D ��0�Ah q�LX ��TD �~-Lm
���Oŀ ,���O؂� ���x;��s�F^��*QĀ��?��r��йv 
8h�O"I�0 t��� C��P�N��H,_�`ޭ  ٸ%?��@-�ހVÈ�X�� ����	����0@�.N� � ƴ?� JSP
��u��j�����_�0?"�� Ή6��-��K耧�ģU|���v]E�(	9��.��Hr��p.( �_��!�q ��:�LJ�h�M����Q��/PC�!��8 ]�7��6�t �͈�h�{ ���V��"0/	|��  ��t)��^��\X� �P����H -O�,�Sb� �(�FK��0 �i�Ӌ��[ �P���� ��?�;�#� (͖H�T(�H� �d��9 3~l1��V\��
���/X!�:5�� W�	s�h��ޝy"� ��ˣ���> �T-`?R ,�Zmg� Q"B�f�	� �+���;>�k ŧ�����> ������� ����%! 	 |]Q�=� ���1�a Y�9/�O@m Q+�:fP� �I*�� ~vHov Ջ
�# ڤ&�z�� -S� ��(}�x� Yq�a4��>Er_Y��©LP2���(�'� ������L ��{k��S
n��>�ػ�&� .��* 1)xN�2� #}�&����^?�� Y�L���5 ��^� �n�����<O���[$�} �½��	l�}N ��Kn ����16���Q�W�Ba���[vO ��_��-�q��\I d{'��� 0>~e�4�&��b���v)�t�T���(� X����@� AK/�#�����)�}8��30[ 	�Zh2�f%���] �>'t��/�����1X 씮գ�� ���
y�g�����F�pM�b2�� ��h5i�0n��#�L`(pN��À��һ� �¤���� �5��=��>e��(5��J�H�vz ��)�p_Iʐq���x�%S �-�0� ���'���yu ��R\�85��� ��e�~�릴���[�f>���tZ� � ���\���	{u��]@G-�D_� ��}�p� l!��IPu ��������*  �Z� H]hY^aI-�x����i�rT��MFC���0h_<�] %��~[��� �#eELnK �&���� ��1�amL��
�R�����D%��`X�� ��'�ֶ?� Ϋ.!���������ڒ=�a &*�QU�1_ 2�,��t� ݐ��"[�� R�h]�*N�����!��5��a���{��*�� X���@�% y�-N��5��n;���" ��bY]_	_�f� ��P!3| �HR�*�4�@�8v1Kr �/���P������f]!�Y0=���	�'�S��� GF��� �|a���� 2�}n@�h%������(L�Z�����S:��� �q������z
�P}� k�J1�: 2�S�Ԑ�� �[��#�L�d1 ^Jh�K=�RzE#�`�U��-� 6\R��Dm ��l��h�q �f	ځ�P� �.Z���Qh���D驠��[@\���X�� ���A��o��v����@�# �K_F}2X'��iA�;���E�\o~ �у\2�h �ʵ��u�� ���g���� aɓ�F�h�Ke��������� ��AbO�� /���M, �֖[pr� މ�P�ɸ�����Z��`�,V-Ah3>`JN �ѯ�(n� �0�F��>����Y@4�r�*� �E��5 �!��:U~��)���I�ny'��_P(�s�
�~��XНس ��N���������)�ds���[T�0�� (@J�4���CSW/8 y��ή���@�4M^ «�̱�E ���U/0�t��B ���E
��<b�jG��U[?�� �ݠ�9����ߺ��%|���H��4�0 	R��� �T-s��g �#C��H ��{��[^ ���4  ��o��~ �Z_�d'U� ������  z�F
�R_�?���hn��$� #���� Q�6��� �ǏIs� 
=���������+Kȱ� �k"�敖| �BQWX%���J����� ����(� �|ȼ]����g9�֤4/�Ԗ<��U�`K#�Y��n��w`���_ �I��ª�U��֑�����v�Q�$��Qa0�p��Ք�B���(�E�8 X[*�bc���`qW°�����f)�lʑ:�X0�r GȘ��h ��a���P<x� #�X0�� ���A��o-=�crU�C�3 ���H��R� �:*_@��'��\�� ۳  ف�5pD�js���,;��l"�
d͌j��Rx��(U����� �����z� ��� ��v?KV 
����[�|����`s\V�xA ��1� N�h_�)>���"�}��]���#Y( ��	V�� �xC��T^ ?�+�-"�s 5��͠�i� ��WHhL�
��˲ Eׄ�� ,��� R�̋1�>����Ѯ�K�R�/�Y�s$�����g��q2�*�?� ��̐� �O��b=|vc<7"p�� ��B$#�R>T� ���O�lD�� �b��K����ǧ�8? ��IV ����ϥ@�� f4�&�* ��	�"v}KB0� p�ΰ1�� (�w��IT.�$� ���8���3`�a����^�D��`氕@d:�?z���xF�a ��֢�geWQP�[Z<�x�V��YKeK����n�T�>N �vd{���:���� ����jio��	P������ %�[�� �Wӽm� ���!�
r�`���� �^+%�PM��D��V�|Q�pnu }�v�m0�~��齮��� ]ZkŃ��� ��0�1�. �Dw�\�/� �q�^}��� a�I�� ��w/ FY�,�Ao�����
�,~�.�� .u��� �W�!ڕ�� �[_�@U�M 0�/Er���.���" �^��w� ��Ղ�|q/>���� 9O����#�p�� �9�h&M%�� S`� W���y_=^!�����"� �΁+�p 14m�ƈ���� �U��ł �_h=w�dj ������:��������'�P@|%T� ���f��� ���R�v� ����	{��� G��-�<0$1�/ �`JW�>� ��!{�Uh�ǽ���m�����S���@���,F� G@[!Y)?/ �*���H �6��­U�=q~ -^�	*� �)����3 �_�y̴���N��s ������Y ���h�B5�� �%�܇A�q� ����[�� /��d��� 1�ęh�b��A]���/��1�2��
���� ����%�
����� CK	�� �S�.:�k� �$�'T���(��� ������Z ���X�y x�$YR�	k �KuEL��� 'X��d
?� �N�(��q� �ܶ; 0z1�U�c� �+�/	d��^ޭ`i���A��ʛ+S� �˽{���& ����F�'u+� U�a{�;�r�%�� � ������ >�?HqQ�a�:�>��N�UMh�P>{�b m�4��� �w����)�� ��L�5 1Ү��xa�9T� fp+X"�CyYH�P �_ �
�VK �!%kz�$�@LQrU� s��u�%R ��eKx� $�@� �� 3�Q).�gG�� �ܢ%�緛k��6/S�TU� Q���h8�0��V���cAぃ�1���=�ފ�E���ğ�W� (P�l��DB�Aa~X0�`�_ n�i���<}��.��<S� 8����
(]���J��5���M`��K脡����(��� ,�D|I�	<�� ������� �J������ <e�Љ�D� u���� �Qx�S �ٍC ˗dY� ����q��&� (�}G���՗��P��u� B�J윦ҁ==5 8A�!�;#�X���L]�� Q���3�'ī��TY��.������Ͻ��ոD  Q�0Lb�,�j��J��%��$�ٓ��Q(}�����e�6t� �u���:� 0 �@�h% �e*�La �K^�<7[� g�0��V  ����^h� ��y��m� ���i��^ʦ �Zq~�n�`%\�ǘΧ� hշ��n �B0!Up� _XFi �uY�H(
Ê/2d: )�!��� h����� ͫ�ڛ��Vtj�Q4,�5 Ŀw�Tu�y ��NQDp�$�)\�� A�|Z!� �K]DS/ȯ ���<6q'92a`�� ���ҙk[}pv*+.� ��t�� #��/x���� Y�AႺ� ��HV�d3� � �����2�A�^#�����LQ&7�����q���	�@D���,`�2+��#����H�� Yhl���㱃V�y7��#���5�~3 ��^��H�0� Ç���,� %߶Pv�ΘA	qV��)ܯ
gQ- J����f�H�}`��2D�  ��P#����z� �����x��b�s�k�`�Z�#� v��v����3�ĭ���,+��8 >	͈̃ �Y�8� ��� �L<N�A3& �Y�	�W� v�k�$����u��୤���G�Ӗz �Sx'��fj}����WK��� ?9��ޕ� 1�L��Z~W6&_^�܍��� ��<�x�[{�?�� ��%�|}�(��=��k��g�w��� �'�s�1ަ 9~^(|@�U �C�՘� �Zs)]1� ���N���;X�Q���?�	��t���\ ���*�e]p�a��J��� O��ۀ	�`���ݰ ��a��\��~��X��@�2ܘ��!F 7��P�>` �CW1l� �p��J��V� ʘ?'��� �$R�%��� 0e��Q� ?�\�� �^���( Jݸ\��%z�r8$`�g`�� Xf��=�(��iu��_h-	Q �5��U���q[�"¨&�^A�����W<��w�h� �d{�|L�1��#@��XT >Bk� H�P�A~�U�`�X�N @?(��䳠����� �g�Ŵ ���f	�A �2@�*0W  ��B��ͮ �!:h6@�] s�%�UB5wl b����X* �X
H�J�В�g^zw��3�'� ��ڭ]!��˫$�/_��.1n>�Q���3��!�h����k�q��OX��@
���=����|� ��j�q "���/�P?�R��e@D���q�К��   �S@/P���u��N2�� 	J�B�h��D���k�o��.�?$'� �Y�Z��\N�V���`���  ri�,Q:AWET5�-� �N�U8�S �#�d,� ��tX��M��.I�;���� LU�W"�� i����oN  �Ӂ�r@� ����[� �Z��F��  �Еʨ�����!���'XPU ��������Z YX��H/� =�JS1ջH݁�	ِ�[��FTIx�{ؑ��j���\�#�W�B;�޺? Z*�R�M5�4)B���_@8�I ��J�u� ��4O��	��"��QH�r�KyI���] ��$<�	�9�-�@�羿~� ���fZ az�q0 ��Xẖ��� 4�E�O��>V �YdC\B��������=��<��,�w�)��b��50�9����`���� ��P(L��� �=�t��p�?܀��X�\W�0 �h^��@ ��fS{�� 
>`��a% 	jywȩ� �'�P}��� �v*ͪ�RQ�C��`��(ۈ�x�%�� ����.�O� ����3a�xA��I0�� �rH(�ҋL ���d�ԗ��i�{�;���$�}[�3�� ������/?� ��X�8��R���/j�����4�*`�h cuTޭՔI~�N	��!@���: �Z?�E[� ��c4!��� K�<	��[�h��?4z+ ޥD������v ����8��6�}�_��T�����&Cb��~8�� �'��9� ��1�{ Z�^���Q]��tP��[�&�uT(k��v- �S�^F�h [�f+'
����;�@ŋ�  �P'!�U����}N��	� �9��k�4� �*(�Z �Y�?���<�G�#�q�v�P�o�k���I��.�ľ� �W�8 �6�)�A�j  *��ơ�Ro��v����@?5�����y� $կI�kU�V}��B��p`� ��s-��~j�2r���� �U���{ �>��i�� ���*�̤� �:��]1�,���Z���=��RAh�03�J�z�&�T;�`r��,& ��q��]�J��x/�Q�����]�@��v� �Y���5�A j10�4� hy��/�;��b����G�$5�@��ʷ>y|��mY�0?� �!/n�Uk	p�� �D\$+�X�����;-� ��
 u{a�h�P3 ���S��M
���p��q������z0	� ����ây2 ��{)�0
G �� g�
� ��l!w���o��R�����5
Q� q��JY�&��H Z�� <�EMb1Y ����V�4�� �g��v_y �=�� �B��XU(�!Y@�:a��u���|���w� ��O���+� 6�-�]������@K~� b��嶋) �Ɋ��ø� '�,6�q�� w����`l���)�%�\��^�4�Nl� ��Zc�H}S_��hL6` ��ݦ� �����g:8����X��ǃ����^�:h�<�
�4ƻ���"�A +t̿`;�H P��\!�=(Ǐ%����?�h��������w��o�� �*Lq��3�i;���f��l�� �rV��w��1=���Y#�h`2�ҢT��ù��鈟�Ň�t��e��� î ?8��ږ3 %b
h��s\\� }��lm#����ʧ� a����S !<h�Ŝ� ��^4��R �"�� FDf'�}�t{ ��	Vl�;��$'~%?��e� �P0�Y�B� @W���� hC0}��� �/��-�� '�&�9��_�H��(�� �b�$p~Șv� JD��h� &F8<� �1	R��׋=��$W�8��p�� q��]ӊ� K�@<�<S�����J �:YR�=� �Gc���' W�%ϼa� /	<�VR_,Hz� ɨZ�S ����ح�o<�t #��R���:���ئ@�� pB0�+W ��Z� G��"l�* �`4��+� R߷VU��M ��y%(���~ʗ��Q��/ �ݕ����� Au��%Q�X< ٨Ρ	vz�d� 3�`=P ��' V�� �G��=XD�r���U� (֪�u�� �h��� ݵ�Y}�:<R��O���A��$�\���%�R.q�� >����.��
��� 1�X �=,��}
 ������ i�3ŪaO8wr�~ jn�RXT�a� �^�U ۦᢂ��a	Bg�w���D�=�%ũ� ��5.[�'� PJ�� {�@�aE�� �Z��6�H��ܵ��W� ��U!��H ��Z��d� e+�-?X K"��[u& Y�P�w��d�����T� �!`�R
� ��nB��@ f)���W��_P(φ�nG �h[J�� ���AwS ��:��>! �x���� L�����@�~���Q}Ax��(@_�.1
 �E���h m��ރ��q� ���c�s� ���o�J ��^[ȋ Vy�N�@� ���H�h"�� kt<�������/b$� ���Inӭ< .CN�/ (��չ� +��g��>d���W	�i�"]U �;LIy �-X=����:�}���WVaI��� ������������ X��K�u� M��{aoh�C���O X�B* ��W;��� ,d#!Z��D�� +X�zam �.�� [� �ְ�㠵���+b��㘘� �Y�\)�0� �[�A�h������� %y(X\
�a�v�fpU�"�T]��o �ۄB�H�ځ�t��*��f ���;͍� +Ȅ�9�-��3�}�����h�e����6�Z� ���#in̫�!C��@m� ���%(��>b ���_r, ���y#�z�
����0K�J����1)W�ET��� ��4���+����23 ��0`��!π �Y1� ��rOL�A�)׃�`�k~�����a��[��$�Y�ـ
� �� `�*Q%�	�|?� ��Z,��R 9�<�.�� �1(��|�� ��`0�Y ���ؓ��/��E��{�
�S�.�� P��JȰ �@�-5�
�&������MY, ���ݜQ��f�['X���: �a�ϥ4q���7���r��G8(���f[�ʀ �˵� �âO��N)g��� }��*�A��]��� �Ј�_ �/Π����y6	^@w�p-e:��;X�zN��=΋| _<j4��ڊ
0�ZsG@[����1�� Yp�LhoJ 	?ݥW�� ��G���:� ���	�� Z��w��D.`�� /\��W |�0�Y^)_�� ˺�X��p �%��u�� Ü��F� W�\��.� ���U_���� ��P��IH( �z'���1� /��h�x�G���3�z��X ��b���\ K@W@*��1ÓR����s���Ն�� ��[
�R��j�K��7���D �x �m�>,��v��+W�(N Q��<���2 	ZY�[�� ��u��_� ��Ї�H��#W�b�=Ӌբ�1@�� ���F���@ Cn]�.�q �o��0����[����)�� �	_�RU"���x n/�b iX�Uf�� ���l��H���n|c��t�` ��B\�H�k ]��b)� a�QU0� j���� hOZ �� �*3V�bcA�n���
��_�2wW 9�O��c!i|D ��*ƀʾ, �t]5 �}� :�)3u�����9�bZ� R�-�= �z��Q��?p����$i=�N�s�O��8 ��(B�W ��E�f L���P�=(%�D����<�� 	���&��Ƨ\s �Y� a��0ɍp ���^���>[h����ٵ �3zǈc O�d�m��s� ���0w  Z鞚��Q�K��ܱ��N ː��|�W0�Y"�F��� ��X�Rj ���1!-.���	}��p�� ��ݐ
,�� �DP�	�������������/՚��H�X0L	N�}�PV2�� R_FҘr5�&v: �2y� \�Ad�� ]O�N^G� ݀,�>9U`�8�n�� �KS݂�� F�!�d��=?O�������P ʬ�.�H	( _����p �7
j�� i�������~՛	#��Y�q��� ZRa�P��- qAi���� B�QX:� cJ�e��<*�w o��Q�I ����k ����2� �rsZ��Q	��ׂ[���L ��KX��C ���}�� �*xOٺ�� b����eu!�R ��1�v�a�c8.�]���T ��x�� ���C�h������� ���ˑ>Q�L�V��0����xh ]�3S@ ������� ��ʞe� F�ﲝ¬ ��c��q M����=� @������rH�-��|]�}S	�@��3�� ��6��_Z 1(�aJ�� ��wq���Ȗ�2c������U��gfh�5�� ����3	Ӏ �n�T8��XKj �e�!���� �4�.�:l�T�s��ڈPX��0� +d����b�����[z. �w�	`�ܹk$d [�'4u�M_� �G��� =!��d�A ��w5��<���� ���C� M�ަ��_��� "���u�2k���C3 ��:�	$Q ����)� ��O�Y� %!���^��A�0 ���	 CY�Kh1��u�.��Ǒ:��b ���_Dm L�޶��W�!*�D��I_ ��6�J0�V�~͂����q@J!L���ݠy�O��h} ?!���5.���+��F)� :��^� �c�E�[S �9�y��� r+ʉ�t�\_w ��Ap��� �/T�xi	Q�g��`��� LK�L� 9m���2
 ]��)׋y� ��Lo�W�t���� ������� �ɩQ�� �Ȯ7-�%$?1� ��>N�� +�/�
W� �0��C ��B�Zi�j��{��@�� d6o���X xqD�Շ�F ��{�����@ ���Os ���ba��� h=�
&�ݍ ����W`� ^bu��� ��+�y�!� ��P������0�L� �򻪉  �ST�O��0� ��蛙�wb~����i���T�� ]F��v��UV�����$T ���+��� �������p d�A°��[ ���\h } ;,+�d��� ��w��a K4�?��(�-���Ql�X�%x �ț) �YR�4GoT �V� �h�EB	�y�"�⮐�G\! '��n�c�<�* K��/>�T��� g��y�'(U�Zp�h0,6�f ��}c'�/
 [�J\t� ̲���<r^�R��J�>� �a �iK ���Yq[_�N�����{b�v�+�n 
�֟�c�Z� *�(�� ̭T�5�p�P�R"�@��� �<�-�� ��_F�^� ���hʮ) �馶6^ ũ�
,� �ͤ�Rt ���D�a	!�À�&@�'����C�d�T�Q� �Ж31���^)������n�8�	5� ƞp~�O�L�X�Ͱu� 0�N�~�)� g����� �!�W1տ� _C�q	�����������H~��@*ڿT u���	��Ņ�U�`p�
�� ��B,b@7 �3�h��Hx s e�N������	\�,T� (�d���; ^��� K��b�ɀ8\�| �p��
J+ Sκ�z�!��@��ǞXR�� �ٽ�M�=[,��L>�u�	� ���SXe� ^��N�$c ��P"כu
 s�h�T� ������| ڗ��u��?0r��Ð�Q�?\�����$0�;}��%�xJ!�5���-�9
 Ql�	���� &�)�8�Y�X�0�-$� (ɉƬ+ ���;W� ���yQ ����D��� 	W��Tvm�!�J���VHZ�Cz� �)�j|� 	����� �V9T$��� %�2�APt ��'��UeB{E�����]� �~<B$����q>�� _�ÿ��3�� |������u �	fhg'�
.������Q@���� �mN0.֝ B/C�����$�N>�����r
 !\j�p#L��,HaB���`�� �9��i�� � ڹG�Z 8:���51� ���<]��� ��KH�s�	������n� gy��1C D/	Ѭ!�Z #ʊ�3� �������� �����#&���� ���؃�|)0�X��Ѣ a����7�u��)����[ -�Y�	3�հ��� �����F���C�д$ �mZeV�F� x�o�W: �]`�h�į+��Л'M_� �S����(׼C�xVQ�� ���h${�A ����y��� �����a�ge� ���>ńb"܃/ D��!ہ�]j@�1�)�� �pU� #ׄ����X�P�֪* >�Q���C ��%��uf�X"N9��`� ���dɱ� �/¸S�e�[1�y���`@ł� ���(�W�sQ�N� �9_2�D! N��0� Uݱ>���^ �P)��٧ ��0Jɾ��� �"�@�}�� �>�ОaO1 ����8 3�F4@���@JL��	�_� K�C�'�� ���B�	 i�Eb��8� ��X�2P9pƁ��_����{%����H� !�3(:� ��x�/6�� ���ah�%�_q�0�`W0?���1ѲT� �=�>tה>�� ������L-�� ��� ��r���g i��GA ��pE� ( \��)[ǥ	 �u�d��� �_+��;΄�2�i���tq� 	ĸ�`�� 8��}�ӄ�[�q R���X+�� ߞ3��� '����� .�a�j��@�����Y�5W �h�~����>v
:lF�`��z ��z(ۼ��]*�K�Q���� �����I��/�|�����`���� �֢ 2�h�I���:� `��&�&�{;�����N�� ���:�u� ��ܾ'��؁�1� �Zb 8�Ir���ܒ\�{�N]T� Ŋw��?;܀L@c!pv�~����D� ����@��]�@`>�)�� �^��{	�?�U��/�}������B �	]��bF�62� V�ta>�`�d� �e m`�v������X����_!�L[�7`�
�|往(�Ad�b1�hψpA� I��퐯�ө����Lz� ��N[@	� �K���+�� �c�_'>�� ���� ��!_C���
\N����OV�F��h�[ ���@H+`�\%c|G:� �
m@u� ��-Y07y � ��?��z� �t�1� :߀�"�Z�'g�G��D��	��u� )���Z ת�0RfT�5L�B`_Z�i �'~s�K\�e��`��\� �����[�	R�� �P�_���9y^L����>��	� ({p�y���|Y.U� �J��Ő 'j�W�����Q����qÊ澎p* �1�0�^ ���H�-& 宧���
�P �F�Ӱ���X|o
:�ț �*;�Q ��4]$ ���=y����I���6���	 C��}�4�`�Q(`��0 ��Y��?� ˝N��1b�������5�C� n*�Q�s
 ��$��%� �( �!aN:��i�� ��Ӆ[����t�P��'��p�T�&�C� ���1���P{! H�~� W�O�� H)KE�P�� �`w @G��@,d�� ���'�w\_�9� �\�t%� 5ac
-3d�,��&R�0�� �6���녜��b�� &�H����[�!� �k�d )^��cK��	�e�h�W3���� ��"2\A �*��~  o�1ˉ>�!9Y� ��Q��| _��نo2x $�~�����:�. (м=�Y ��5�n�Xh�e�p	� ��1�w��� �5��/�[� ���K���4 "�Q��aX�� �>٬�X�}%��-��Bo� �\[���hW ��4�0����! '�^��v�> e�W�{7?+���X
 ދ(�OUb Y���P#�}t ���X��1 ����� �(�H��� h�*%Uf�� (�S�q�3�  �"��ʨZ �2a$:���3��������# �A�R�*��8�2 �Z��� ~���SܦF�Im� �!�� ���Uj�� ���k��X hP��#�X��$ �x	Q�� ����0�ԆjW���	�S�H� �(��k��F%_P�e�� df��~���Tغt����1�3) ���8� �	!�^+D�[�����.��� �#�3(�! ��X���P�� _�B<ؔ�� 1ZR�	��괂ǘ�(P&��� VTtRX ?�B�g�EW� 	C��}��S* ǻ��^�o C����MH�*8� V�m��i/pU 5��#�$^K ��sٻ�	qB�ڀ��*����%+ ��U�M @Խ�$�k���0'O;�F��]����/� +���'h@��	#ʹ1�G6��X �����t+� �;�%Y"� R��,b�B� +�����p8��b�b!�(��)���:�@^�" �SA��>���-� �խvn� �Mh0ZW �}� ��z��$�j�� "��=��u�%�^� �9��a� �qW�B�� z$����r:ù�K��I�R�H�Aq�0��;�~���D`�2P��H [/x��� �1��T�h Ou��" �̱1<d� � >��Ŵ&���J�5��(���.,�~�K:��'��P������(	O�`ظ��Y�'��p�PV X^F�� ����b ���I2m-[ h��΀*� �G ��6�[�F�T/+쭯 �_(��0� �N�	�\8 ���h�;� �
	H������ �0��i  ��7P ���f��u&���	)���u� @��Ⱦ�- �f}����� ���1Ջ�W�ㄧ��C,����p�R��g�)��� �N�[@1	 \�l*b�LJ h=%�v���	rY2��/�&�|�}�N�hp�^�q���A��� x�)J��� �3��2� ��[�P�ArX��t�7T����W �/@����� wZ.��P��4 ��H	�ج�@���Y��[�W���]�+�8�9� PZ��Xw hΠ��� ��cu'_� ݄9�� ��߯�R� o]�QM�5$��
 ��"�� �K���X� ����S�-� �s����� �G*���2�w�CT���� ',�"��]SW�6����/��+ �Q�ė� �� ��Z��  3c1G)�,\�� �0��� ���@fht��&������ 	j������ \"gtX�� -�Uţ�� ��/S$�vm�n�X�. � x[�ZV��ľ�a��0�F #�у	�bZ1w�PպB����� r+�� �*ġ.�H��%5p ����ߦ�������l
 ��U2Ә}|���^� �#��[�np������ܕ�6`=R�@������ ��������-X}����JU��$�ē]z OaY��.	!�f��ɍ� bk�Uu�*Y��� ��/��  +��@��Rt fb2�|��` z�'�*��� [�75��\2R K���9����`���F~��D�zАr�F�Z π eR%h�����\E:�jF�𥚟n��%������o=^wmvJ��q1��zE�쏱��4g*M �i_��Z�:vP-V�\� �R�Stz ���Ϸ5�p ǽ٬�Q
 ��\P�>�: -��[!'F �V�y �Y��{P^ k�7��ݑ	+ r� �
�� e��0�`� 	�!ڀ�� [�$��SB�� n"Jk.&�Z�I`��  ،��&�����0�����J�!�[鹎_� �d4Ab�,���ط���� p���SU;���ᴱ܀�"˽�_�I����ys���+^pL�H�AG� ����� ��	0\����Zڨ���b �`�{m'�� �	�Wyx& ��a�:0� �Z��� �rGʑ��A��!pQ.HR�s�&�T"}�� � ��D��c����љ5a ��*��{� ��+��!���ŀ��� �%K���'�PGR#��j, g������v	0'���_�=uP #�"�-�rC?��Χ��}{\��� �|��`">L��C.�ک��~� �>��f� -�^vl��%Za�׀�e�9 �"���` �Z(^��6 �5�sD�� �̥c.¤ �w��� �OR��mÂ ��F��i{YPު��U����h��B��~�� !�Kάk]�p� �X���� �`xT�޽��w|�[^�Ŗ� �`Z�h�(�|# �S���ز-�Z��r*<������h&Y ����'��8{U j�YXx*�%y�\�Ǣ�@3zL�����`�rK� ��ֿ	�)���0� `��ڜ� �$Z�O ���p��- �6�+�! ��
���C���*��rs �<��c���[�e�����X�K�.�3� ���e
� �a����C u����]��gpnh�� ��t� ���W~� ������YS ����I� �81%7�� �P�e�����G f �W H^��a�� 3�1�*�L�4 P뗱��.��[�ɠ�Q?�, m�B�Dʇ� �5^
ƭ� ���%B�@}��N��S	�> ���ͩ�5�)m�� �A��陶+ �xB-o�U $.���� "O���Q�}�~:��*�����C��X�@���$�[V/��<���sz }�{�R��	 Y[h�4��L����u 5��	\�p% �dM�B�c����I�a�XRCZ.��eJ	 �!x��� ��%��r0p��s �E�]ޞ�� 0�_X��wۋ/q �<�M�=V�� >2���1 !�/e���V�0&�"�B��{�".W ������Oc@��zh, 3~a��l|=x� �+O����
��� F��%]��}��5�ٸ� �(�k��	�I Q�DR��]n �p�Z�I� 鍉;Lr���T�._�&-�{��.�N ў'u{�� /�2+(�� 0�j��X�����H��`�R� �E%P� ����-��h����t�y7 k�qdD-f ��SA�W �{@��� �_kbx(}�� ���^\��Q �cH"8U� ���y2bLO��8:(��T� Z�,�� �󾓴���k'Y����h��M���F ��
���$  =tI�̓�&^ AY�!�Z�ź��C���=-����E� �։a�N�Aw� +�]����' _ �$�F% ~�bc�w	 �7ɕ=�� �Tp�f�C� �þ��"�Z �鳐���<8À𠍀�� �m��U�J���� yo&[��2 ���ʭ���/��@��B�� r=q��"�}�內�e�û�3���v �-���*��	�����`{f I�K�0���e�,� �P� �#�!XG �["�<�f��Z �~�ںs�yV ������Q �l^��zv� y�a�����." ��^$�0��'�6 ޿���^��Z 4u�2�ػ  O��*�X#� ���	0K� ��È���} )_"�[Q�����*p�B�K����7�>��=����)��_� L�{ݷ��m��� ~c�W 2���]��� uF�&SE '}����\ �(�@o�w�B�� ���i� ������
�yOs���:�0؏̐�� ȱ��}�[ �Y�d�����
 ��^R����X-�_���1�t(^�p�ٗ@ �� @k���8G;w����Nr���v�L�[|�=R �ܱ�����^�ǃ@��!��S�/�2�����N� D�`����}� W�ݝ^�p� ƀS��Q� h�����>=��ЁY �
ˈ���	�-0��� � X	�)ӈ� ���[qm� 0��Ҩ�F� C/�)� ��A��[� ��c��s� �˟�U�� 89��h�J�̀$3�t� �/)��ZP�qd ������ ���� �Z�DUp� �O�o�%�� 1�N*	��� h-�bG4 �����;D N�Ƥ��$��-����h q4=�8�&N����ο�� KP�<��S�� ����1����Lj�Zh%InP���vb ~T�	�/u �ԗ�$Q�7 ����\� �&}4�m��h��������ۻ@�M��?�u'Q��J
�1�V30L��%/� �A�T�X��.�~�S@"fB=�8 C�}�dJ� ��/\�O�� �k$��A��� �	W\�I=� ��.��yaL���q�� �l�U��� �V��%��F -�Z/q�� �J���rs6I@��8k Vx� ��&��f��� ^�c.�	9 C�_�� �>Z��5 �����O��2� ��� U��
�/!��t=��1�R ��� �{�/�����PP_���(� �\2��Y<����1Q>4�� �5O2�XW������NH�LRx `D&"�d ��ᫀ��U�wC^	��[�d �p4{ٕ #g�'�Z�h���ė��� �,�! ������ ��D9�X�� ��k.���`:,�H� �_X�s�1 ��bO^��TP�� 	�hǾ0=V
�K� A�f!��Jq���<� �Z��p��	W��d ���=�y���6)\�' b�.�Ô �S�&
��P]� ��1W�j�����/�Z�Pht|�^�g�� �VXj��@ ���QA�\���L�O��R! �}0��u 3�B��Ȱ> �!Q�P�  �i�g�� ��	�O��_���5 �H~p\�� J��(�;�� 	�X�ZC��2?���Q� _��u�wXDH� ��7�)��g@��^�ͨ�+f�]��Z��r ��-"ET |�%���s�V��� p7�0�y��l\�� [)ݩ]�+�'������)q��@
��t Нј�{�;� }>]Ĳ�U�E�N$%`�-F������� �X�v�[� �� B}�� lZ5��7���0 �'�H�� n�N�{-D� �0��!ـ &�E��udH �����4� �B$��:�b[�Jछ� �+N��I<A`@�	�S��ewH��:_ ���]�� PһF��JQ�a��Z*�iY0��	+�k� !���EA���*�$A~����E�@��0���r� ��?��K B�@U�����9[_@���R� ��'�3��� _��� �~NX��Z9��=�^`ߒ &]�8Y�s�f�Ai :��oa���*�Ӑ�ɱ,$��>+��G \/�c�(��|��h ����5�&�l��t!3 >DQ#�� ,KE�.�ݙ&/� ~c�X�0�J0� ޻ �V���� U��H�K ])��
�S ~�L�O�} &-��4�hsM �N�K{_�"p���0( �'���	Y� {�t.%2k� H!��&0�� �њ�{�� ��R�� >�D4.ol ]W�����q> �{_鍥� � �p�\<P3 �W�ο���F�KӪ�k��i����1�X=�тtYQ�`���d�K�XO��Gp�V �*�Έ�ްQ[���J�M�Z����`��w ��^��=�x�Y�V��<H���I� s� �f�	��Р�ֱP�@���&�8݉{�Yx �V��%� Xb���� I��a.�'�`�������[W!E�h����RP^ uĐ� �� �1Hyo�e��8��*g�@��4� ���%1(A�t*z���b���L�� �v��1�2� F���cR� .C����P	+�n��)K��Q�}�h�ZI$���"c�&�7f R��w� W>��5�1���Yx���a�� ���_+Q�ȇ%��h�p Z�@�J0o\ z ��C��հ s	<�!��=�/�&@`@�RW� �t�J<�ޝ@ꀾ�M� Q���B���Dh��{�֫��|
 t-�i���!�@�V�	���zp"`_R�� ��i��n w`Xa�z��E<)T dN� nek�o�W�La� 0Ì'��u �F@�H��� ���a�y� ��%��$ 5P�i/
@� �`���� ��KЖ�� ��P#��'o?H� Y �p8�Aw���,���� 
tO�.g'�e�0,}#�2��}�W @����/��  J��&#�`������?���ր�! ň���-3�W �).�S�i ��LU�[_�<@뀢�]	��9��Z���� ���v/�a �	�f7X9R��r(���Q �?]���[ �C�0����2.@�� Q�Bt
 �\�}J��� ���O�֝�+C����)S ��U*з�P g ���\0 x�F�5t�|�@ku��� s͸�Ac�� ��Q��:y �)��u� �_����t ���>�� *�R��� �~@�� � �>"�ڨ �H�(�v� �>�/�;R� �N��`�� �A�� ��D[�7�X�(� �m��Z������(�$h��{��M \�Q�+ ���x��h<��6ec�U+�T� �2���_���h{�@9�>0���!�. ���X~� '^:�"�� $�V�O�@� �Q�!�f -�]+�@E
k���Q!닊a�ܷ=~ �Q��� �b=@�ϓ!`�|��~8X%Z
'� �i��qk		T� ��c� �!�t�;u��.���8,� ��-ݔ �ꝒM�L�4×����Q�� =2�&�R�8݃��*� YZ0H�m@� ����b�U G��.��l �y��_�>r�\&|� ���6� ������j˳#��T ��/�R��(<	ҹKZ� 1Ȩ��v� Ė�q�����XwN��z �ہ(��$� ��"- � �B�d�Z��^k� Vl�L��!<@��O�� N���Y �,F�!K� g�ϐ��^ ������� ����4�( ���^D��=&p�� X#�|� �Q�;�% ���3߉�=Qr�Ig|��� ����P0��� _+��d1���@�� t���9j|� ف�X�	���� VT�$�:~��xC@^p� �bH]ɠ�� �,�G��' �x �3� �L[�R,	
e�{�������p� ��P����{��zԿ`�%?���� P��"�� ����=�p ?x[1K�� W��Z�V ��*"}L='}� O���:�J B	_t�Q��CX*RP�Z/H� 9zq��! �	"���<���Zb��vK��L\�&U�� �RQW� Ai>0�Fn� �����Y��s ��\S� V�5���� Ъ�L%��� �ㅍ�� ���	4 ���E�F+8O<���M�����^��֬�p�P ��[�� ��*������$��`�3�� ����W�0.�� ��d9��\T� ՙ�+x	 ����h1J Q�?���� ������u0 ����!�$�봀B_��,1I��|J@h]� �^ϜY���of�W���� �B��.2 |͉�+�Z �ٯ�E�I( bT��๎ L���I ���d���pl ���7�T &���:��˗CV�/1�����> �ES��Nk�9�	[�C~���"��u� �L��U�ա����w` � ,ث/�g�G ��|��@�� ��U�OH�T ũ�� 5ӗ�)`�N% ��Z�-��qC��H ����T�n�	ķ>�W ӆ�u&� ��ۄ)�	��}ԇ�KpA���6 0����1��� �+�gS����'�y ���k� ��a
CV b݋��T��{) ��erџXo��"�1<�p#DQՅ��$(xη �_IeRq� ����!����'��R�͔� �}re3�1���k�6�� Aʈ�Y?�H� ��/�a�ɘ�F_��G�S �	Ձ�e (-Cͪ�=.��1Ծ�0���2 �
�Z�'�� �Gt(�4҈ ȫ��yV& hR�19;8� Zt#���ao'�Y�߬� ���m�Z�H ��l��� h�A��. ո=9�K����s���j��"B�\~��Q��hC� �<����$�%�R��n���x �'�W�?� ��`[
3 �5�d_O����6��Ě� �N����/ �`�Y
[�9�� 7�Jw5 (����Ҿ ��XvV�7�:�~�µ9~�l� "�؈�<ȝ�р�`v�4���Gg��b H^���s�)W��Z�X�p �^r��$F h#,�6�Wy� ��(�I�J �{�E�� �
�~!� ����4� �E�]ߖ2� ��u�G� �T0B�)R+ ��cl�2U9W�@;���� �*�s�l�p�ϰw:���A��@��ї W������|:��t��� �Z,�^�2��5��?�a�1�c���郋��
*��� �	�&�\�� !�}.5kU 6�	Ώ�� w\�%`< �nye�a1 �q
����B��(w '���o�v�$)��<�=��
��u J���~�- �v2��n��k�x ����	Y����I���� �V�	�vD ��'k\����a�� J�� @�]z�P ���5��"� �����d���o&�~*�_e;� �t
O�N�	���%u�-����� ���(��� ��^/�{`�F�I��(i�V��� ^�����,�V
H����Q��~�;��*�O�P$ʭ� �Q�
�>M���%�����L�f�`6�۹���yJ �����?fȗ �6���^�O��>��� ��_����/ �3J�@X�? %�W�=� [���~���Hp�<{\ xVT-�� #�pj��994w ������%H2>.� ❮��I{.�1 c�}�>]�����K- +ȟ>��0�� �O6�$����3���E���Q lְ01� !Ȼ��T�B  �A��p 'E���� ����,� �0�]
U2� ����@�  ݝg�`�U h-|8!�[� �?�W#xD�,�7� ��Xz�:�����aCU T]&�,� X���Bh1NI��:��2Y \fi��lӧ�we��@[�G ��ZϿ I��|�k�D��*и�2	 \�?����{/ �YA=R��` ��,�)�����$�2���C~}� �k���D�}�H�{�HV� k��%� �_�B� ��/���� Z��	��ܠ Y̊
�LHV-m�' �%!�� ��M��y�Q ��$�Ű���`��>�(�CO�����؀��L�3 <9Xm0o� ���� ��BY�
4 P�����+ �^�,�J���΁��qf��xA�	��$`��8� �.�!ӈ �D1�����/��[Tj�� 3Sf�IN@ �����*8� Y-��4h���(]����t/ �G�=� ��wFvH���S��p�	�z l!�F(���q ����ѝ\� ?�c�/� <��B�#�� "���A�����e`W̾ � ��/��	 s�u��P q2%@�mn  �^OY�; 4
聢��V _vr���: *G����J�$NS��	� _w��qA�>���O�1 "��4kD� �,�`W��lv��^8�� ��|	�{�~*�\ }7�nf��Z�� �N��A2߅��������#0�p���
 ��	�?��y!����0Ȝ ��h���� \���C��= s���Q�L�~>�t �f��ͻ T|�p����L�}ݨ�b� t��$Y� �X1��Zh& b5\P~�B ��R��aAN z�}E�+[�v�J6�ʅ�� t ��lhP�m �~cN-^ @�1�TY��:Ȭ $��|z��z��
��qg�	��u`� �7����S]�! ��Ҙ�%~�c���T����+	 )�VP᩸. �<�M�-�k� �BF�K�V�#�!��_�-� ���'Pk� ��;�,v�^�� �S= ��� E���A�� �pC �Z
�Y�� b�Q�� ;��~�*�x�h,�[D�`���pn#G\���C����e-V���3���	�'�\u�e�z8�� (����� ��0Ń�_���Y!�`�^(i���}_x��p����	S`!ݫ� �w8�g�O�E����I�,~� ^c��%	z� �v�(�y)��E�S�> ��1�%��`0��Z�L�. K½pO��4 �1� ��%���C鞆��w���N���EXi �
_����	1I���������u ����M�=�f8�Q�ꎉ�p _} �A�?%��x� 
�����t�;�����|��1 T
!Ŝ i�K%� O��J�q��:^ۦ� M�� ـ�m��-@ �N^��� �ܲ���	=u� �<�I/�� �f1�>Ph K6���� �
��Ay� �*�ŅE� �Q��]8� �S �|H� ���X�� ��h�L�� �Z�v�A��9�:�J�V� ގ����S a������}�;�\��Q� -[,�\^: 1�Y/�(qV
��H	� �s_y S�ۑ]iB�x��ʁ@,�?

�)Ÿ� ��Ё� M��w�sb|iN�` � � P������c>XĀQ������_� ���\Y4�p�0:� ŉ�f�� ��񎰡(�?)�`�� ��f��@ ��H��$^� �0�\2X�� �N��@d �'��q<��W�����z�R ���%��
 P��I�7�b�0�����#�� R�бL��� |��V�<� �8B���{� �r���p�wѳ:��� �4N��, Ȑ�2� �-�0�PV �8�s^� t 
��_G�fQ-�0|s�ׇ�� ��!�h�� :+L`/��7c�`0�4P! H��>�O s7~5�Ʌ4 ��� ���a�k� 2#�g�U��t 
"�b)�X� 6u/�2pV?�^�j�Cg�I���% �&�N4Zur�����_���C���<@�/���XD��}��L�,���@�� ֭3R�X9�b�| �WS2 ��%j�u�� ���5� ��k�b J��?��(�� E��ς@�� w�`�o .3�1�_;���D �bS� Y	��ۘ� �O�i���_+I� ����	:���5h/ �B� �VK#��=� Z�y쐽���Мɉ�]5� n��LZ� iė��	G�vT��0�� j�¥�ܗ0�} >�ﲹHu@W	c��g�~�����w \j��2��- K'�͗�,�� 馺$�1�\	@	� ^���H; ��5�wt8d�������7�e��K!��):�G} A�/�@9�^s�:	� �X��G��_����`-���} ����L/��⍮�()� �"���'+�  ����T�}��:����U �#Afa#1H c� ���U�젊�8^�i�:�{�����} ˓ۜ	� �U�Zh[\&��} ./��b ��hR��]� �1�����@ ;�Yt~�0���@O��k�� |�:�(� �}$���� ��3I,��LaP C�ۀHW1ѿs]�ɢ@���* ����{�� �v� 9h�_ ɣ~�m$�C�/��'k�_v ���, �齎\%B 4WO�Q�] q��C��Z	nK�^߉l)��H���Q" �T(:�a. �t��&%Z '_�Q�Ԑ ��L�dV�&O!�*��'B���N�5��-�aYW��@���, �q��X �h�<��8��(��}� DJ�C�}L �tAX�I�e��8dN�;���1� ���o���� @��P�dZ ����NcB �=�%�6O� �w�� t�Q���Y���h���^d=�};x�������XW e����{ 7�(�̇� �_��=�M9X)�y⠿U�< �%��>��¶ZV�@t�k|}���+�O� Ş�-T	� ����I 4 �u�C[0�S������ ���o�t9L�L ,�2 r6$� �лN��� �\��"� ��>ѝ;Г0繊�S��P|�,�A� 	��*+� �X�H�A��͉�!���[Vh Y��\w3~k0�N �n�Ƌb B�Z��� `a3�2� ��T�o�f/	������|�2 �O �	� �Ԅ{s���?5΅'�����<�)Ւ|����T \[V=�	�B ���h�{I��ـd�  ���}�t]��w 1ծ�PZݱs��(���O�< ?�M�� C(���$�~4F�g !���]��Hh �Y(���)�Uݟ�� �1���E|���� S������N� 9����Z� ���E ��K������C-���J|�� K�y��� ᷈Q.�� ��kF�?I�$@R렚��\�X� X���\ 3:�G�"|'W�� q&�� c����?/����\�ܗ� P('�[K V��1��� ��L�%Q(F��ci �H|��� �������w ��I����{�J���1�@�ʢ6�fD ��_%��t� {	jz��'e��I���B���y01�*֡�W��i���?;�w �n�a ��!��� �JP��y� ��8O��+�<�w Ʒ���Z_"��&�_�/N��t����4�%z` /���>����-�Vr� �xZ��j�9	
� ,�#��� Ơ r��[�(|J����:\�GÛȭH�0�:�X� )����W� @���k��� 6��$��+�I*R׀VR����8] �
Z�N� ǮF����c&!���$-��j��]��\* 
�v�`�>�0�=^-����`
R��T�L�3[��uu
�� h�����wb ����y�I� ������ _т��?�:s���,��d�� $P! D��y� �u��~�G �y��Q���|��0�$3�P|��	��Jp��>G 1�&����X�L��_��/�, Gg߁xXZ[o�K�R��dy�&z��w�ue|-�l��� Q����X� ��'�R? #:��[� �(@+��l EG�9�y� ֐^J��-; ��o	� �����~b��_vˁ҃oz�W��B��_{h��� �'�ܙP�]ƽ �¦hZ{b e��q��ꘓ�� l
�tچ�|� ���(�_H�ї�`�W��V��[X �h6��==p 2���@�P "Ӹ�RD����p�u�mdZ��Ķ�q�< �A�y���sDfLO���_E� Q�����>H,�N
<��+�A?���[ Yfh-B��Q�m�@͌t� ��>c� ��IW(=۞ ڌt3�� ��y!�
Y;ÀO��u[� 1�'�Jt�_ ���Z6�!. W>K�� #Ё�F� f@"�2��0 �]^!�)��a����������* �h�&���?�˸�}. ��{V����+ ^����� �J2��'k� �E��O(���K:ӑ���9�	� 7���5.n !4@��3�A Ԯ�gX��n �Z%#��Q� ��R!��Y�, �߸�t5@ [�QU�Np ���4��l� �(�qK�J ��`,��l_	��S}8�-�.��U�ȃ�)���L�n��k {%}5P��� ?�N�WR�`l�a���6.^Ј����U#�O�f����˞arp�� �a�M*��� P%�(���& �ZS���9 � ��:� �����h ����THN� �Zr�a��� kId�)1Y ��-u ��P��U�If/V#*Ѿ�'֐�\kv�:Pj��� Y�^�$ .�p��L!w��@6|D�P/  �ؖ*2�� .��l�&�H�4�� ���@ ��N��`K� #h�v��	;W���-ݴg��4�d���� >�,߆�[w����1=�O�"�Q��� �ەX W! �����=�� E8�Ԙ!1�'X��:A:�dj�c�$}�/�� �\h� eN��i�U�< 8��(@X~8��t>�Xf�J��@)]d�H�
N���3^� �`/�Y������|�r>\�� +�t���6 ��nL�4hɸ�[��a� OP.�G����S�� �0�( >%׹�	Ե ��;_�� ���R� ��e�VG<t �Y����xI9S ��F�Xx� [�+��� ����w( W#����Q`��i ��*䂝�x ��2�c� �m=��?9d�	�H �'v���* ˟�x�}ZL�� �!O�bK	�S����� ��I��/��� ɬ� ����w������أ����� �L�91o�� ,*�\5��D �����A��P�� LufX\�z #'��Ol�j U�����,��)^Ѧ�
�� '����	��G 2�(�� i��$ʩ>�# ���"�		���  ��D;� ̺��}�2 �56YQF-�@>CDZ��e|%t��05pL ��ё�� 	�W`��/ !��_�����.�:>x�BJW�t��u ﱠY��� �P�'չ���-O���Z ��>�(�P��z�U:D$�w�-��Z ��1E	� [����AC �ˑ����B ��E]i�s
��@�"�`3v�,�Š��c���s�u����Rڧ ��	����� )��E�F� ��{�/�y7+8`���8���@X�]� �	x���>0�@��� %�r�� vJ�M�Ơ��Q (X��[���� �� A��3E\ۄ &��[' ����5i7X�� h���}6L�� �Z��+� �2�1
�����Y���Up �H��N��"B�@��p�$d��3�X� ��C�F`ޱ
�/��� ������PK�, ����! M���8�m@��t?i^�XH7U<�` ´�&w� �1�L+鿧 �_8�{c��"o
W�p~$e] ȖH�a˻ �\��[ � �J"�3Wa4�$�����T^%H9Xu����Y�).�g��	��h �5�x>P��ZV�_��p:� a�T� ��D�^� ��a�V�� �� ��� �T�RJ
� �A�].�B��<O�#�`n� ������M?���΀�����n��ē �P��v��) ��, '�# �!���M� ��%����R �������e
�߳��Az�_��1�
 2*���!^ �W�L�5� ⁮�9/Jo�?�<�Ĳ6 zrZ�(� !�Ȃ�i��HS�����k'
_˸Q��.rd2�RB �N	+ǋ* �3:������Y��jư��� �b<��,@ �/���l�?迀�V�� Ѿ��̥�# �R�� �ν`� �����%�z`�_�� �	ב��;(��4E���`q��	�:������ Q�2Y&%  pE@_�)P��Z?�9$�K����� r�h�!ڲL 	�[&Z��.�� >��"/ 34
,Q �Y� ��<�� ���ן�'� ̄w���B��R����väf*�%� Xr�+�/[ 1����J�a <2�V&����'~���k
5쩔� �&`2� ��UG.�A �D�z��	��ƭ(����˕s&R�[<`����#�*���H��ڥ���P��ht�/�J�7���0��[9�FǨS{� _�7(ڞa �#�.�i����&g ��F[�� }"���w�T����G�e� *m���kx�\n� �+N�� ��\:�� �^;R�W��N�/�Y� ��B��ݖⴣ� 'Z��!�0��� �TՕ8�� Q�,o	�� �u�О�l�����@*�\"N���qR�2��%�u���nSx+ ���U0� �}���i�
1~� �]��U��t���J-�	B����a��U����#Rx�и!�2���Ⱥ4��L�*�vh�:9���ǁE�V�GJ!1�n��7� PQO�����3���6�@�R��-w�(�P� O��K�� �q� ��f���98�i W�jHyJ ��!ѯ�� ��%T"�� 6�bSLB�� s҂���p�|�I�\tԉ' `�1��.� @��E{�z� �������� !���N_� �C���� �%Y{*a'�9^ �&�NW���^5 k9�S�� Z�����r��Ǌ�� ���� �����(��h �� `UC�	3���"�J���� ���� ����{� �G�a� I2��.� �*#��\䫨Q�`&<��+�<hY 6胴z�~ B����ƣ ��[#�pt -Εc����Ԋ���?��p '�-]rF&9U	 �G�,�x ��ZW
[� ��*�C0 I��dM���A}� �����_, ��Y���T�� ��~��c&�P��}� �:P��7��z�hGt� ���!��8�����ɮb�ܔ15�lB��ײ`�h �J$���ap ��V��'��Hr	�N�G���@ S#Ґ�g i�Ǒ'� u��J�$� ÏP4�� ����<Ԕ �XJ�W��&o���֐��s� ��X����ja�@u�������e�����8^_ б{9�K����f������Ӹ~�V�o .|��[� � �Z�{�	���|�P�2� bܕ��@��Y���H�� yfa�Ԑ��� 2�B#��	 &@ֹQpJ�t%iWр,�� A����oH�70��]@^���B9]��!p`l�s �kR(�$�� >w O -Z7%���b�8|���XQ?�M ����'bf A�ђ�Q�� �!:�ǖ�nM�j��)�^��c ��|P$�%�c�p���/�\ ��&I��E ��a�
�<&��/�_2�6K��H��
�`�W@�<X�P��Q �8���� ��,%��Hx� �G����N����0h����C��K)�G%�t��P�/��w !0�pRN��V����9�^�[X`���i�� 1�L;�  ��A��� DC�,S_[0>�p�	���u� �٧O��B���s���I]1��ï�f�C���x� O��pb*�� �ŗ�g������� *�<Q "�S��E� ٕ��H8� Z�o[Y6 ��hb( �B^��x�]c@��O�<n=f_ �B�Z~�� ���0��@{�$��`���� c��Y8� �x��ɠ�pB
hF逬	È�X(��˷s�u��;�3 GP��(�=Z��zl�W�K _�B�S13�x�pAH��0�� ӆ�WO�� I�8�γ 3 D���'1�� 
BS]V�Itp�� M�� ��H�UY[ \��h�Kg ��!#���9��L:�>I���qu��U�f�V�YS5<��L�{��*9H퉀\�� 1�آ>'� 	F�82
 ��Z��*���~\�)/�܄4�B;� ���#��:�� )����W�O <� o����pn= M�	���� ��R�5(���4s��e���|� )�h�s�_�*�&�� ���� �C��\� [�*��W	�)+� ��#  D�� 	�dR!ͺ�f��`�'��^�عP�Ƅ:��H��$~{�4 XV ���P���� �jK��̘! N���e� 3��O�� Q\�ŋ8L��@SU �!�] ^� r�S�s�	�X
��u�T� �C�;��� ��i��Ng�}� !8�����O �s�' �� �Q����&-� �*@+�T��%�~�� ������ �\��Z!� �.H'���K ��ȑC��:f �� ����j �O��\I �VU��� ��pQql�ϣ���)I��\�
��w�`<$�3�8 @]ʽ�	 �տ��ɹ�_  5J��>����� )մ4��6.��wD�E�O Ġ7>�'�_@��$�]�1�~ �� ���j=�E� �����:�$ Pи�H�` �3�: ���+��� �R��������a��03 V���	�f [���4 � Y�ٷ�� {��ӿ!��ds�`@���S{ �PQ)ڮ�? 	��w.<Y��� [�^ ��h��/.J��2$�����# [Z�	qp0����<����0- @��]�ٝQ�a �j�%� o⼭�$�(OЦခ��B K�g;��[ 	ݤ4X�dH �khP�� 
�1�X�c ����8z B^)!�V�H ������, Ŀ�y2� �x'�T|X <���Rh�F ����@Q�:�Y�O���"�6�ق���Xa� V��c�XU^��H�鿗C���Bp���}�x�|�F�O��Ks %�m��*�H0� ��&ؾ�	h���:�d�0�^]��b��k�!˯(��P�}�q�=O����,R �+�5���?� [}��V&�=������� ������ ����	� ���R�%H^� �6�
$�[ *�������i�п�=��!Ր� ^�P�����'��`Pȫ�]KJ��9���  �T/2�U���ݰ�*�^� ѴGEeg&M�/CZ��8 ����+�����(@�b @��C�ʗ p��0�8�&U9���[�7i��V��� һ���_�� ,�U�$	d ��@+^� ��1"����5 ���J��t ����!�`* �i%|e-&H 1�[�{�.����Q�0r�p x)PF+I�\ �����[� Z
��K�) Y�1�:z� �Z$�BC  �P�9�ׂ] r[�)��=���`�ZY��h@e�[�u0�� ��/G��x!��U}u��{`�� i)��\�G �NS�`� ��%�Ð �f)0�[�( �hJ��+�Hbs P����T��~I�_}"%.`@fR��S �4Y�����3�����q���y� +�[��ͬ m���	��h���[O�V� WB������_�1#퀝|ڗ �!�	Ȩ� �`��q?� �_u�bEW&�A���}�! ��LN� �hn�0�� �P��[��d #()ي ��! ����DÚ�*�$�e�i�a �������} �M�kI�tK�ɲ���ف@�v���KR��H�� �Y+�Z��i�� }h&�U�5���l�� ��X�<��YK~���g ^	����6�D���ȟ������� %wF��'� ��Ю)�:�mC��`�� ��]�"ȧ� ���ZK�� ���T��� ����z�+ �͢�����ގ5����2�B��e{����`Ͻ�\� �3J*�[Q �ذI�`�� ��N6���8 ���>
ڶ�%x�p^��B���.1?�Y��?�D�j buC��V��(�d�>�cd�鯻���h)`�� �K�%�� y-�Z/sR [�{'eJ^ �K��Y���Z�"0c�l�D������H���/+ �慠҃��Ch �^�&�%;���X�:B���� -��I�l� �Z��&BH�� ��4��$�PS���(�	󥂂!�v� ���W\�n �qƗ�u ,_�(�[y1�'~ *�.Օ �	�m��"� S0J��z�L�1��U.�} ~BK��Xd b�H�ŀ�+� ��˰fY� L����^��z0�(� 
�K�?/�j���6�� ^wv���yZzR�������� ��cUb�V� �WX"���!�2�3pZ{� <��K�5��I3��� ��D�(�0:�����2��Ub�w��B  "t6V�%�� �O�5��� ����m;�����V� UA<�W����j�R$��/� ЗJH�, 5g��B�� �6 �(	�}��q'��&ʋ� ��"gQ�� x��M�.��o�?�V��b­ ����w�; �{c�1�� '��Y`2� ��@{H-q �&�B�� ����ܝP ��Z"�d�\���*t���Unt� �d�2�Wx��e�~�@�h�r��[ ���%�� v 5����}g@�@��]�8�W�8ڷdk� �	xL���q ���~�&�����0 ������R`�"_��^���c����a����� S(�w �F|<�[��� ��\�'
�uKi� Z[��SY$�M�bx�@�a� 63�1� �$��EF� �t�IU}w,�*	�F�=�0� �	�XZS�J� h�,p?P� ��"K��� $� յ�0� :ײST[�=]/�1�֜a ���
  (;'�T�&�d������x�S�a�� ��*�$� �t��<?q� ;KzY��йb��W�K�$(7 �q��f���DCe�"���U�� -̶��� ���
�B� ��%����@�O@��� ��_W"Q��/�8p��������U�\�f 'Ȱ���v]Y�2=���ȑ~�AXwh>� h�J����RT|�q��� ��Z��0,� �UP+HΞ��݉�>��u �,-�S� �c���[� X閑��~�$x�<K�.�`��/�z.�eb�j �	,u� ������ ������� ���zV�ys�N�Q�[Z&�& )����;�:YN�����j ��.��Z˭?�7�긋�� ����jtK ��s�ز� ^mrh��5N\��Ҭ�H o1�	�Z 0�/�)ȕ�0��~�� ��1k�(� �D���ut 뢒�?׮��S����W�X ��\|���ؗ̀���=�e�0�hp&�� U@*S��O Y'����4��u� �Ia�wxcd� �P��X �[�QG�yq@  �k]�V #��;H( �W�R@��� ��瘭rM�Dl  ����
<�9R���CKf��) �*��I֐ �S�EZy B���_�@����@㩳�yW�� >��K����� P �&�I=���l�*�U��J�i�q`��X(��s�	1ѷ`]�d����s�*#�YV��  W���?_Z x��62 �ɍ#��L�8�ޯ|��'��WB-�`�c�x/ �A��u f�'�]���l���#!�>`���yn`WM\� �)���� 侲	컨A<�[�sa��i-e(fX�]�%�ZQ&�<h���gI�u���v} r���5!�zj 9�?�_ � �GU���v�� I8���:@�)o �`{���ȏ���ٶ I����Hq� �Y�sX ?�O��h'��� 3��� )} 
�$���U ��`*�Vh� �\}���0� �%	� ����o� ��N'2wH hJ0�L* ]���t� �
x:=�Y� �b����P �Z����`B(\X� �<�� �w�o]�� �ͩz�-7 1[^�V=�yq �b�Ch x_QE����+3�鴭��a���E��ǩ8���t �����2 Z�Q�S&�3.�h��`��1*Zh�jƛ� S']��茕 �O�8T# 5A?��:��� ��4<���� �1����K�X| ��P�/ �q�A�m�;�Hb��؁�5� t/�v�$:'����*`E ��@8�R eV2ɸt��,ED� �$}�! �L�Z�� �,b0���r�]��' �x�E�o) *q��� �[3v� %_�BLZ�	 \hP��� rq��������X��WTZ� I�(R��:{��O\_`�� �|I`��)� ��7��� �~i�4��(�B}�0��JV )����8q *��{N!���0�~�� �Ѱ(�K�� �X	8
A+���'�� ���I�3�מ ��/���o.Q��	ք�X	hMj�{N��E�7��XAo��?��ë� ��l^HU�{ SVP���t ���%v� �&(� �K"��� ]#ש��@ ��-|�U<_ ����)�,:b �>��2#a&�L	�Z�I>�҃��u����L�� �D?��З ��9󴸪3�Փj�������)��@ F�\���镨3������O�����!�	v� ���6[ZLV?~Ā�����rO8�VrM	���A��Gf*�@
� ����v Ye�Ĭ�, I (#��[�p� ���1�_: ҋ�+.�i Q�7�0I�� `Z�J@vW��%3��<�s]=�'� e�E\��� 8�|�pP�DJ%(ǠvH�a �])��_�� �h�t��� u�>gR! ���Q�yW�O��_���/ ъ�!s�?o�'���<��)���q�" ��{u��@ Ӿ�'B�~ ���R�u|��Ƴ�*�X�����Z-0���|��%��SU �:��#�� 5K��f�A.͊ n`����� (���/��U��5�� �(�	 k��� �S#L�m�$ �e-_���C W<�!�� ~2�X�)� п���z� �>A�{�����=@^1�%� �$��9cd� �t\���~�����{�܎�,Q#� �
kx� }ȵSR%�� �nF$
�	 W�z�51��qC ��_�M�,�RT����� !���̈� _�}����k 	ũf��\ 3։x�����[W��U0	�@�+���i ��q�.1�����
4�� ��0)�P%�:[� ^��T/��3�� �s�<:,�����Қ��B�Y� �����j��f�N��1��2- \�|��#�B�L E� �� ԑ17�!�� �Z��[`�B�	���`��ɐ\��N�b �&v�M��� ��[鎶�*�k�-���ľxL'] �d�3`gzF Q����%"� �-���o�˽�'���)�( �&I������ H�^�]N�:��Z� >�?H�9��Y�x4���8�V��_\� �
���C *�!��;�9M�c�`����P� +�ԟ��\ �c��^R����A ��W"8SN �3�~���Q ��nR0��$������v�&68 �JQ� ��v�Y_t{� �1�e�?�M ���olR 'V�^Yci ���`��� �[�Z	�Y +u�=/�RA��^Q��!��?0�@ �|O��
<�������
��K�b<9���E�(� ���!� � �B#�6O� ��C9b������~��8���&x� �3�S} !��^~n��"U��V�i!� �0�A��=> �Pk���L /1�Z���@ \	Їׁ� 3�u��q�t'X��:k��P��@T���$�P��U �G{�Q\�9i���5�� ��N���� #�`�w[�ixVweH	nm��!��h����^�`�X�� ������� �����v8 �#-��[Q ���p�� ���	�� ~ �f�z^r�E">�ժD�ZP����t�c��H~K ��$�U�� _h�3�bW�]-)�@�}e�P�� ��$��Ǟ R��+��� ��	J�v� �b�1��Y �AI���Z����.���8T]�~� H̦J�,��!��F��^*~ 	���<UԐ��YW�� �L��0�� ��K�D����2�����h��D(�]�<
�* ��V���` h�Y�迴��a
��#�R��@�����Z+������ ������K8 ���|�< ���#�� �N���ӂ����� �W�t�՝ ����� ��[��}v� �l���΄ ��ac4s �er<�� ����|� 1#�p�`y ����	P �|�W���ft-��@�(�;!��rP��D�Hn����{� ��1�_� �Xʹ� �/����0�� k�(]3 �vK�,�}X_휋��i: ��ϸc��;o�%e&�� �Z�@�� �K1�����`�;�p���I)�Nt ���7!O�@ "3��޶Ĝ��d���n�-�`t���������~ h_m�M� ����\�,eѪ��NV.�1��`���~�P �2p�t���� ��:<��޹� �ۧp��/�� �!�& �^��[��Ew�`Ö��� ���-GP �d�,��Z�\z~�����gn�l��^� �J)�Q����5 ��Ȼ,�h�O��_�� �6��90�ZA<@-h� %�UD�eW�� �e+�x� 0ݽqV'���@=%��tP	\����{�����~�>�w ������ @��-��� �%V�ƥ+�=��5�����hL� �?�%�\t "(nB;�X �*��H@,�� 1��;�&=�Kd���3� �� #�(a^��%���@�]k�8��MK}.������0�)��]`*��� P��20��X~H �WZ_` �uP!�35 ݋��=U����$�� 6��| ��T�Oꪊ�N	����3S�� n �����8�=���93�#�ITl�.$� i��И��%k�J� (�����z v��˹:��k��G X`�ؿ�� ��աT%S� m�HDQ[� #�X��C� )鋐��uS!�Y�0���
 ��ʼZ;J� >OY�#+� efD'�4�� ���$�ʢ�X�� av�&S>��p1 �s�3(b����������� ��(Ә�)e�@���V�� ��a�q�63 ��I�S#@� �,�_��%� !�� Ҡ9��������@MQ +��.��i ��1˘8� $\%��	� �p۸�l ��3�2�v� �B1n�a0�<.���=���� 1Uw!�yA�]0ذ���Xp2 x�$��_-����2�� D���P�8]Q�j��%�Զ�~?W�i����� P��.��a ��0_�� >9���5� �hVH����Ҷ�i0 ��	Y ��f�}�I ������ [葧� �����:Y9�F�ɰ@�ٸ� ��o��˽ $�*�^ڌ �c>�N����,gu@P<��
eQ��[H0��X W|p�߼ �
!���g�m���Pݔ �Ʀ�(�Y��T��P�P�Ӹ0�������� EZK��H:9��S���B ����WkM �!ȹ;
"�.�3� 4����y|0��c��<|a'�p�] $��v���>����%h3��1��D� �2��t�'��0F3�R)�.����!��Z /�E��Ԉ�L��3U� )�S �1ݬ�
�( �5Q�	��# <zH� �~S���`�P"7B��v� :�6ڼ� �!�\��%� �
���	�W/H�������Z`�lv� �7���,Zf��+�o_�!�Q�i�B@ JZ���H9�-�������� �y�X�x V0�Z^�� ������� �Y��E)� �� ��K���i������� J&�n��^#Z��]b�a��A��&1� E���Xѓ(�� (����:�� �_�r�d� ��(˵¢�2�_H�D�@�% KL�P��>�:������<^ ˥'%�y� �UA�0�! E���[��8�2]	 9
��/H �#���ޑ ��;�!r��#�(��0 �\�_���#��+�ژ�PȮ�;(0����Y p<hH�4���j��8�.Qd ����W�\ -�Ĵǝ�D�c�锃R_�ɀ�Q?�M frSLP	� G@���9[�a��KE��޸	��΢ h�2�N_P\u�)�~ ���J� ��˜��&Rk���Ρ�	��~������%�y`0|� �� ��ď;��R��@����uG �<[��	 �*έPXu�} �'FA	z�.�RU���+@ Z	Ɂ��1 �`�U��  ���
�2PC{� �1Zh��u ��㯅�' �D�L ��K>�b&�@	S�ŋ�<��p(��� ALQ��� ���Vh{x�� �� ~'Cju)ǩ ݘ���� 	Z�mSѬ h*KR�,��� �ɓN'����V�Q{ީ )�p\�M1:ȃ�л/�[���� �h�0�"N ��dE��7����~`B3������F�<���U�	l�C�R �p��J �� r5#� 
�n�1��. �W sJA���[�'z( ��o�\��JUW[�`�8<��L�<����Zy_���� ��?�(ʃ M��ш� ��o�\ �V�- U�7��ͦr ��@���K �!��Z  �ȁ�X�� ����ó�  �ݝp�Yb�%[�H��I*`,B�lU;�����Q� ������ _)g�S?���o����+�\��\Q�q�X[wF�5N>��@�f���$!n ��	�Di|� ѽ�Ñ�n���`j�� 9��2��㌾�  @B	�d�V�?���<�� �XA��^ :�Bq�/� ~��1����	����0 4۸%�>�y� p����q� �h����PU�V�D��%�� Ix 80H$SI ��\�) �[������z ��Y��x^� �!73ȅ� T��E�hpS ��o�C�vA H~DT ��.���� @¾�o��� ���Icu19�/ ����� �tE�*$�����dD^������P
��%�����ps|&�� xU�Y� ,��A����(�_���ps� ��/�D�@Pp��v� ��ʡ�}ӗ��)��&X�
���0%�@`�(�T�4ߢ�B�RW $J�0���;��)��w]	��ZO�71ӉsK�@��ȆX���R�@����� ���1[&! ��ķV�7 ���a�,Y� .���� �ɯ`�I��� .Ehg2 	�fO���ј��S���HRȉ=� ܾ'��^ ��4ޟ:�� �Pb$�5`+ ���>��'Y eJ/�1��?.�~] �hAg�#���(;�� 9�T��� �" YP�w^ ��}�Z�| E��sh�9% /�"�R��S�o��_d�:!��r }��Q ���zOi� ���π =�}�1��t_��;o�-�]Ģ hb[��8 ��G{0�g��#� 	��i�� y����!?/�_��&�  ҝ�R����k[��B����� !�q�P S��B
�yIb��K~��� ,Z5����� L�1X��@��\�,��� ڹ�-
� O�/Z#X �H�P��* ſQ�L�1_��BA�3��rF�R�K��ހj���h��>\���|H ���_�]YJkw���B� #b����{� �,U\�� M�N����eXi- pd'�A~� $,���a.� �}�:̸�8 C<���K��&�
���x~�B����k u6�K���w#�[����PՖ�~] �\Z���{{� ��`�h~Y(�9��X RV�S8�w� �L��l� ���(A_ 
z�9`ʻN:��#��� ���vX VA0W3¿,�����S#�=�c'Ε�q-� �t71�d�t� �aK
�\�L�� lNU�Kb �=��B#� �a�s4�2 �+��ƍ la�8���컅��!�1�` r����I ��/�B$���V��2��~ a��8�.<�Z�i��%) +^ k���ؒ X��r@�.�ڢ5�cI ��(��	�<ɿ���ҕ� �Sb�;��c=( �R�F��1�ZI��JQ H�p��b� �₄P������	?�@�-y���p0���)�3+��;`�� �����V
���G�<f�a#9�[ �p���r X ��YL�� %��'�ѧ1��S��hM� (��>K��޸ ��Q)W� Z*ˁwk��h�0���4 ����R�� �|?�L�� �
S����� ��j��-�9 ؀̈���] J���� $d+��0 �򔗥���:�=��ͨ�P8��Z�b X����.� �(Y��b� �1��fd� 0'�\�a�� X��9�H�F�~����]� 2��A��B  �_�`!h�T }��%�2��s��� ��S��7��g�`ڄ�ٲ�#���	P��(˹A^
��2ǐ5 �1$0��K�r���X Y�W���.Ă���� N������]<�Y����# $;�3�-H ��D�Uo�� �h+R�x c]��W�tu�H �Ϗ	��(= �Z��u�) �L�C!��� z�n���� �Y�W8h0�Q�����K?��!�@�&VD1 9+�n(�� �P���Z^S:�TE�����+�����I�Rr	 �u��2�p� �����x [w^P �1ҋ�
%!њ�r�)�a�a ����� /h^T� ���,a��	��� !^3� �,j){���/}�PQ~� `݉��:�0O����� ����-�U^Vf��C����p��	0��O�7�YUS�.3��8 =�'����s� RIi�)_SL �C�'Wd� �B+T�	0� }E�$�f z���_^ 0���6 K4��W��n�P!�_��A~� Z�D$����0�[�3���-��r R�oA����� ��>wY�H�I�/���� �}����� �n�� �mN\�kW� {2H^�|:���M��\R��Z��`�E��jՀ$. �ʾ���� ��e�D�0��/�q�`z�! �����#� ���ك͸��ݤW���&ҏ� ��A3_ ~�X*L	-�x D��g��.�=+����>T����iY|�9�+��OLψ��?�3 �wju�<� l� �[�-]D� �Q ��+ù� �"����O�� ���C�� f�4R�� �h*y�$� É�Hq�%� /�~`�u �Ax�����_���.�ʌ� S�l�) �[����	T �������� -�u��� X�r�`�{�w� ��%�_+(��"гc��\ �8l��|�_@���� W@���`� p�f� Ӑ�0�Y+��@'�f�n�`J �Aø�2¯3U����� K��yB�w |`UQIՊ�����.�� ������ �����]3�^Q�݀�0�f����L��� *����Et<�`0�W� ������� ����ʙ�� �������&{�7���� ��հ� ����9��� ��Ү+. �m�N�	5Z�� �R՗�UI
ef�� ��}xJq��1�Z02o�v�p�s�:�3� Q��<��W� ����o~|��a�����
"����; ����/T ��G��� hI|ě�K� VQ2��D� ���	:_A �[(�-�>gu���"��V@ L��`�� #ݘi%��BH}�m� �� G����P@]�ȉ.�(�-a�ٶ� ����y��A������� p{���j������иp���Q�"����� �'N��+ �龉%�	W�0�࿳s�Cp����%� ���:�X��Dn����+�P��!���p� �2�|�v�	�1�@YD ��h�<"� f�T����@ S(���#� pX��/����t��}Zh�BKPHP�� )���CW� �5"�r]� ���~N��x}��<��� �2+c) Ϙ��6��nMK�`~ !�0��'�� 9}>oP#����~����Q"��bg	^~� ���/��� BnYҭ!� ��X^��/ i9�}�� ����� ��R��W �7������h�&�I�ҋ �"�b��$��T��Z-���E)ٵ����m ��H�����L��[�@�ů� �2R딾�r
 �:��W�m `��÷�� Ȑ��'X��� �</De#o ���H� ���ŗd���/���_x���϶����2t��@�]����R+ϺLj o�U�� @?껠��DMt� ��Z���ʹ�	c !sѰ�%d� �z����L ��F��1�:����N����-� ��2.�:� XҺ`��g� C�^סYD �)SQ]fq\;�ǀ0���@� #˟�҄����-�'���]�&�!��j�G�x�� |	S{$`� (·7�%)� P��S�D�z�^���pTY+w\�G���� �.A����q��P��\��}vڌ��i�
��|�Pb@�s�^�� �_�@~�/�x뢺s��1 Dջ�z	!� C��0�5��q�C �h*V N��2ղx� :��h-�Q� @���^�c���Z�f	��`8� 9ӵ��P �\xȇ�X �'�3�` %Z�_���q�'�2��� ���JV��հ� �����o,� -�AY�49 \���E��� 617���V`�� ��&j�Lɍ~^<Akyo���Y Z��!��� ����<: �-X�qu�]w1Q�C9�ܵ �e"d� z8����	���_R|%0�Y�0H�x-� Ѫ��o%� �邚;�_)�� �?{��P3�	���c�2���� ��b��W�� ��e�P�� �OQ�	�!� ����ӝ�� ��KD��� /w�(<d �`��\����� WJ��*� s=��hlX�� TR����� ��,�0>۹ L��(��,��� ^�fh�>��"��p%x�( N��e��:�DJ�B�u��U{. 
x��\t�6 �ɶ�|/ ?�h��K����:$�g�%��� ����,K����ج�� 4	�+3՘ �(ڔ?�� ��v�_eH0E 1��sh���02NS	�D���(��n	��* ��e�Wq�x �́���)���0�wӢ�޷C��`~  [��� "�\�h� [sX%F���	�ۀvi@�� ��u�Kb��W��f�Z)��"�L�-�� ��GC[5���t` �
ހ2O� �� �b�B �]���� ؟�V�`�����XH�0Q�8@��(�~k�S�>�Qf PhZ 0�� �#��[� Ł�q]�{� ��E`�F�zN�� ��Q��:��~� ��o�;�8� O�,���pu�w� ���1�
{  ."�Z�N*FH�=v�≋��J� }{at�� ��hO:�Cl ��s IWŶ��լ�%\�J �B!�y��� ^ۿ#���� ]��u~��1�L�; 2�B�C r�8�b) ���гI�h �Q�~�}�/�����u� d�wD���.��ab��*:�/�Q�k�� �aPt�`�N�e �%�e�i�y ]�?�Y�F �# �Ӏ� (�Z��`=� �$�7R� �}◰�]� t�0���m k�#}�$%���lJ�� ����P�X$ZY���� ��B�L�(��_ �Q�j-� �X4/��w�0������&ς� ��V� �ȟ��0H{ j���˷����a�S}�<m�ħ ����A�3�s�0�bڀQ7T� O���L�' 1��lwt��В��d���,�~�>�����7�
 G �QW݁ ���;�$�'9/\ ��CI���K��3��d���1�@|�f:촡6 �=�� ���S���x� r!��] Ԁ 	�
0q����8����P�T�b ��H���AO E~����x>	��]��%^.� ��h�WY����' ��#4���gu� ���Wq� ڿ��1 �A�����Z _����7^�~��@Y�U?�8� S��.��r��@�_�'ԝ�GZɿ���R �w��B��	��0�ES�f�$k�4��9P�� f�h1�9�C �З	�[0��w-��z���(|ؿ�h�� Ё`�c��#L�[ +�_�/� ��O0�T< ��-؝2�W��QV}q�a0�_ �6%��'�� }������;������O����h�z ��	�F� ��v@�,X� �Ң2� S�"+�A� K��'��~��w#0��� ����4-� 3�'t� �����1� ��w`�����(*�WӸ�� ���n�)�/�]��RC�b�J�[d�'�vP`�u� z�3$���1��s� d#�P��������^�� �"?Q�ȋ�;(Ԟ�I@�h�p��| N_R�@� 	٘���LQ� !L���yhTg�*'�:���%�0�� мta�V��,&ǐ�� }3��a1 
����� \���tv���5ơp?�]����[��*@� yxLY��t���V���@��`�.�01А�2  bYT����<>����m�@��&w� �<4�� �Q.���j ����\6�9Ĵ���� ZK��(ibOԉ�s� I��� ��� �<�cJ�Gt -��ގ~�w��Yj�\T��� ���qP������}��0����4� ����#� ���S0x _3o^�� �P��p� )	���� �dV��n�>�z�B�@���pX fS�P��t.�9�&��^����Z�'��Pkȝ"�,�@1 U��� v)��Ȟ�}$:�A i�ٶ�BQ�`��������RK"�����d0Z��x�^����fe�Pǀ��8kt��(N��'��K �^v�4�?L (��:XQ\ �ϵ@�hܚ���-v�����o4�.ZQs R�����0�tX	��D��8� ���h<�2a�H����8 L���5�� jk����}H�r��Z��&�B����_�p%��s�Ј`5� j�� I� )������l��h0P���� ����T-)����cv�X5Ux�@a��@F�4������\�y|��;�/� ��3nO�����A� R� 8�^�d� �����C�Ӱ��*�V� ��k��8�p�G��{� ��eb#ˋ�-�<? h �FP	UR� ��_d��3� �؀�fU�� `ܕB�+ �E.0��� ���a��o� �#�+�� V	q*�R?�ǿ-A�� G!���L� �7���n� x*�P�� s��+µ� X�F����[
�� �-e�� ���J;�g�T �w��b/�5	uh��\�q%�@֟A S�]�� � �T[�u ��<�K� �WZ[*� P��B�]�I^�D��R�����W�-��q.k)�C0 ���
��̴�����j��� -�L��F@#HJ����?�l~41�a3�p�h �Q
۹#� �p�	O� t��U�����`�_� �6���Ⲟ ��\
�h�U���ݥ� �q�(�^��ܱi�� �$��=��kP�׋+�c[�E6�������� ������� [ּN��� ��:^��  ������ 2mw&^x� P��¸ʩ ��I������7`��	l� f�$!�s�� A ֗�� d�>Я�&W �98v�� |m��4���n "���j���Lk��O)4ذ� �'�1ag| &H����i]�Q"/0�W����2JԪж�c
V@�v+�^� 1�X�C}u� 
0�u1�] ��Q+��y� h���$t�� [�KI �T h'R�%� s���U� ����Ik<�9 ����� ��b��Z � �Oh$C�� 5d:�{�,�um'|T��j��`Z'
p;�Q���9�X�&ꪄ ='1��3ή��#��	"�t Ë��<� �;��� sS��Ȩ5 F�y�$a�>ޭৈ��!4�� �<�^B6��]�@p�%�W �t���1*2��b�߸��X�8\�b�oS��
 U8P�H[)%�go�ő�2� �<lK���� ��ES�����ܶO��H �Y:�W�;�`��� S�g���2w A��Ѓ�H ����d�/a "�:�_�� ��Q��hO�Na$����+ �b	�{7�p@�P6��0��V �o����Y1?��%>D�� �H�ƽn͜ X���u� �h/"�$ ����#}8 �SU��Ր 0vX(��MQaJ�`2�xT �k����]� ��}|��- �m
yq  �K��� ����h�0��� ��W|��}� Ґ���r�w�ԟW( f�΂� �"g
���H�6��_����	 ��:�}&c8�B�M �A�x ��7�ɽY� ����m��H��y1�%� !G'��(�PQ�0H �|��O1��/�D�y�� �^�"�\��]H���Z� ���!��b�3(AN����V�%���&�	ˉ�W�?�vQ�$� �8��W�� -a��\:���h�F $�2"�T ����3�\� �1	]�0�,�X�O��y� 1��W� �)x0����Y Z�H$��� _�8 ��! �R��G��/ͽC%��� �T3���4� =O*��җ{9'�� � �N��򁂄0�`X*�a���L� Ҡ���0�s8 ����,hEj �z�$�Y��������_Uvs �?被������2��vR<���|��]�� �y��XٷD A%!�����@0��k�:r� Z�<V��/�~`>Q�@Gb� ���G��� �V(�h3
 F��4�{Y$u�i���/ Z��k�� �O���H��v'>װ;
�� �dP��) �^*����Z �/E5�A �`2�ZNP�V��Ȫ� ď^�_� ?�</�3!� BQj��WS�XC�,T� (H�q��	�!zӀX�� ��[� �kP���-
 ��Ȓ�ќ79~ ٪)�;�� 9"��V=�� ��S��� �����P� ��d�#�� �����AphX�^��z$~ � ��[w��ty�.�I�0�� ����@�W�zR�	��@�[
	���^���w�v4�&o �y$_�<�
���D�v�[�`ي���Y3��Dpƣ��2l ��4�FQ�� S	�ho��-*��u�7��H�n?���P��d�J������p ��0<�(�U��.)��P ��z#�;W���k\�l� ʉ+��]�-[0�`�~��/v�ݻpF��_� %߷,� �1X�8?Z'�ް�_0�@��Q�l��$�Ά� GV[�;h�vF?�)�za\!�4V�hAq���95�� ]fAɜ�u�	w�O  |�-S )��n�� ��WY% �.<�'� ���1�� �]q�bp 9Q*��:u�i�S 1�h)�$��zj�Cv�5�?�� �p�X� �bC�f/�	�]�� ����_ j3�
�r�K ߙ�d�R/��P�s@e�F�^	�� י��Ϙ d�M���	�\��$0 �`���L����Ǒ�`�Pq�kpn�/�̋��ţDx�а�+	 �S"�}{�= '��r�B鰬�mz+��4� ����J�� `��oN�[ �� ����R0���*�����1 ����	�&�6� �f)H���%5`Cy	�Z #������ؼ }�lG��x� ��f'R,Q\� �B��� n%�� �~�!��r	SM�x��N늣X[���~v:�� ��D<� ���O���X̧x ����b�` �Y_r���R�O��=�G ����[�,pu �Q��6T�� ��iK��Bh jz��H�4I,W	l��b�C_�Г���P�X�m�� ��>�y�e!����ɦ����v� �;>6�b�� �����)� #M��Āժ��l��0	�;�z���|�%��p1�����]���!����S͂-�*�,½p��2 ����� Q#�CZ�s ;����¥p� [�W~�8ϱ��Lȴ H�'`(� �� ��<l 8��ğ(->�ڗZ�����Й��ݻ���J Q�D���� 5|n��@M ��L4�TG	}ܰ��0���� k�a@�� �(]%��
��w�ga���_ *��O硭  �[�pH�} :�b-ݤ]Y>� )k�0_��-�(� "���f` U	�T�:�����3�Q��!�B� w�dʞٵ��s0Y� RJ��&U (,����  DP�k "�?�� ��q�1�� )dH�v� �����XEN5� *b�hXPA��&� ���=3����,| ���R�m�'K��V1���z;} �/�˕�F� ��x&�8� '�V�
o  ���K��� 0[�C����u� ).�_RI���u�Š ���D�h���%!��(>/ �=�����{����� FW�K����� ȁ��Y>�; �Q(��� ��8V���4����с�Y1� �cG�q[�u �����S��b`��nC̀D��vW���TP镨V;# �1@��e xj	���%|s�� >`f5��,�8� U�� �#� �[�7���� ���2g!�`Q�JZ�ڙl �����
�� M�b�	~�K#RU 6����]D`C�%ȫ�V�����ئ��pP��� ��G��i2�� T�K��`p7|� �y_�b� ��d���1pe W�6UV�> ad�
@�\K���Ǯ@�.` OA���%� �_�]ĝ�:p� ��w�S? o�7��yv�]t��ȕ uB�EG���V���>���d����;��A�� ��p*Ӣ�������@J0]{^�1�(��I �!Y�&>���=Z�� ~� '�Tc��| �O�:jD�r2 �!��<�y ��Wg�s;��N`���� P1ʳ=<���
 �W���Rig9B@ �ߵXd �����-i��o��b��F	y'�C,k�	� M�/�Q �����PM i'�:��m�X #y�p5�.����� m�a�IU��x&�ȍ)�� ��߰[UK� :�S���H� 0����zK��_@�O�� �\��2���U3 ����0X�Ji��	I| ,<O����Xs� ^�2}ct� �"�~��� �Q��`� J%D�� �@�Z��V��� �1ۡQ ��\(h� !:�g�͡ Z#��+��	?���!��>"8 �ʰn9^�9�� ��B��'� ���0l�����({� \�����
{]�	����^���W� �{dG�g� U[Y��a+����Sa쀰=�4�9���q`@�d��{���XKS���q)��2p� �Z����h +uY:�j� ci��T����л �d%)��C�,?�W������ g�C8���	��ĸ ��\�)&/0���!Y���� pD���"��r{���L�w�)�Qʸ��&Z��W�� x]5z���9E_����Y���� 'S3\ѳIPy��� �� �J��+� t ��f.�K� �A�a�h7!�����`�� ���� ��,&!�� f�C	_�`��5mD�v? ���H�X�\��@G~� �����Q �,��:��H׶��%`� ��e&�W�B �v�E
�� ���}� `!·M�J ��'�/���~�-0��k�z �����.�� N�!L+�"��PTr�Ā�Ⱥ?:��*���b�r� ��v�X�o� �3���*��vG��O�������	�S�� �\XZ) ^�d�_��� J�B3�V���^�� �o�O @�W��JU�(��u�	N��� !_ 0�P�"�h] �+﬽�?�*;_�E��9 Kɪ��@� S*ﻆ4�à{�l�3ɦp ȝ�m ,P�	��E ��`���K���� ��Beu ��)�Z X��������B %�ؿ�qN� ]��J�1. �y�A�Ml$6�� /�3��Fu��H*���k�i`�!��u��1J #,���"� xM����� �(F�@�� D�W05 K���eC�����*đ� L�1�x_� V��P�aN�hi������� 0-�v2$� �:�F�� ��h�"��IpP*��[L��N��"�� 8��Zh}wj �$Q�e�� �*K��wꐯ �(��! �?=�<��#��,萳�'�R�Z�`�O���c  �3.�V� �Ɓ��'Rn�`����h�Bj�����%G�>����Ҁ�uQ�� �X.-}T$ �̋!��S�v�;]�� �^'|	s� w�(��SE�� �J٢o�U`�� &�Z%~���[�����K�\<< U��+��	�X��� �~ev6䝱���_?ʀ�ـh���.h��s��/|�����б [鈫N����%�܊z" �)��Φ�+�/�v�ཨ n��Y^%�� ��jE���ڼ`�*;| lX��E�' V������O�DF��� �Y��GX V��7tR� ��I��L�� !��U�w�FC��P��@e !��]�H$���$�%?, �tc�4���X�2�=�?�-0�> ����Y< �$��. ���-S� �/� ��	�*��w��D ������Q� �0�A�� �4����� E^�w���(�
��% V�c��P:X �^�2���e*��" ��o!ǻK�e� ��H�U0 ^Ϋ���� B����� ���>�H*�& ��� �q�C���t�H�X��!�0�iY���[�D ��-�P�ّ �]�d�; gy2��MoǦ�����>a�y�= ��OSheZ T��@&������W%� PYI��X5��x�_�e�t+ �RS�N� '�!(ږ$>�ǒR3�@Z	�p'# %�2�w�����\�� �@��b5 u���|�����nw�\�%��@1ډ!� ���y`� 0��R��Lu[�ä�� �����x� �ꊳ�f!� Nj~�1ڃ?!�ܜ�� �	���Z��9����3�8� *�u�MW	N �_���1P��� $*�p��j�l��w���ʃ� �Q��6��%ݡ�{�@4.�]��l��3Zu q�W�����*�H �_��y'� :uA��i R�(�N ;>	ֻ�� ���
ڐ�\ �.Kͼ8�Ox�w� H��c1�x�З ��R�O.��= ZI�:P��) ����Ĉ� B�Y1��� �+� �Ӡ �!õ��5w XP��uv/� �S��;���3K��b�	)c� lM �|T��<�6� 
]�eU  ��y���˚�B�VI-X ��ƿ	�hY "T��U�K��m%�J��� �.'�$�R ��L��Z�x:Ow 2���� Y�C�%�dX`� ���T�9?���-!�Xk� ֦��	�Z�A~�/E��Y9����@L�ws�, �1����������Kt�������S��_���~��`�\2���D����	X�+� ���ؗpi ��=���Đ5 �L����p ���Ezi�;��J�a"YpEL Q�X�4�R At��+=�� ��`� C����� ���^�P*���~�h�u �< �^Š���� �mZ����T [�	�-x4/�w��f`��]��`��x ;����? ��*[֨R� o���A�� �H)`�!�@ǯ��%��C�����Q�Y� �,�� X0H�J ��k��,�xŤ`.#9��_^@v0X�Upt��XKtC��@�x��X�7 [ՋLO9Z� =�AJ5�i �l�㣚�H�q ���� v(S�Z�5�቗+��t�, ���zͿqk �|�H�Y ��h����v���@i��X֝�3�"�|���_������!�a]��Y*���	h�V�zvy�r����`n�1��N-$�:ð�[^��>�O���p�I?����^����6���kmz�_�)O �� �����w�� 0��DƁ ��M���n �[Y��E ��ȸgxb�#/ �@ѻӤ �a_fߍ�P �W��p��0�	�9_Yv<��O\/{OP �1����h!)(|�� �0���� J/G��[��I�R�s���>�@��1�/'� L�$�0%���V��-�`"��\p����2�]�I �0l*XLZ �t�)�AI��;ȃ�ۀ���5f��`1a���� /�{�6=f�+G�P�� ��k��|� �`���p���� �W�� ��O�a� �J1�~����������>�@`MM ��0��S|'_m�
�� �r�ZY��S����h�d� �}D@![� ���H�0 �F`���g ����X�Ǻn%(�������c����.pM �]7#�� U��LF@;\�p����h�ˢ�)��,b��H����u��0��ѧ�@��i֢� G�"�_� wb6u+��$�_�<��\��e����l�7�y.N�� ��[�>O ǮAM�ˇ 
�"C��1 ���k�Q�4����y�j��:� ���3/d� ^��+(ݾ%9�}�S�� ���kr�� �t=��PU&��� ��D������ �dz&�� B����	��:��N��^DU�� t��pk.��a8���-��D ��nU��zY _���$�� Ə���2�� ��Gn� ���	��P`�� ��fRQS�-���������o8)� ��LfX�%$ �*�[� �Z�'��� �7-"�1� �KR���� @gC��5 \K���^ �2Pm@1� &\I|8��b�Uec�[�jW�=�zh�+�/ !��*5���gX������ �C�
�cz��\ S�QW��-� �������� @%mP"��'��x�Q��0�5�BҠp$i%X4bL� ��v�� �mٴ!�n���ŋW: [�Oa�Dq �?�\/l@ ����5,�0] �)��X ���`�_(����� 1���3�@Eh�U���#* ��'�ϕ�� (�	BZ�U�^����O �Y-�� �W�T*�\i>�VĖ�k���dH(s�@�[������ĝl Ⱦ�%�F�-}� �ﰞ1� P��57���@����m���P7��c��Z�bT`�S0��#AoRp_�	(����`��?��]pu"� �+K[Ph�� &T%��EQ?��� �Y��L�&I[���� �
-~�x� Q0ڹrL� C/��_�� b��� U�ǘ��Y@o�h `SJ���	[H��@X!�_? F��K�V"ۨ8ף�� W&(Z	/�R �h�j�w�� ��|9Q�z���0`�u�*� ��X_Q/V�<�G�|@��D�H X�0��z�� ):�1���R ��8$јn�� '�0�;� ڳFE �:� Չ���, Z���X� h�N����� ɒ����` JΈ�U��� ��]�_�9� �%\�+�9�H �Z��v�/wܸ ��@�+�L�n �R�	~L���^F��]�-1R|Z@T�����.�+� O�~��n���I��?_��AC �/�Sm�~�������.�ߘ� ?�����	j�H ��S iGy�	A�|? �#�P�g J6�yH�&1 b�����t=��>N�|X�J �;����,���*���Z�� ����4iL� �0z��� �{R�q��M ��\����X6v�Z���&��1����^�Կ� ����|�$;�H ^w+o���D����� :LĐ�Ӣ W��g�s���"���`� W�ò��f� 5���t 1Ȃj"]PݠJɷ B�Y4^ ���/9W�X�� B$���Y)8� �j�a "�%�|��< #�/�	�!;,Ȗ�G;��t����t�Z�j��]�x� �fh�H�"�-��޽��{�2k ��j;�DR���@��U��đ��C��E���k ��/[ �,�o�p�+�� �&A:;r bKWH� hm`!П� ����IA+ ��U4�`w�@��(@Z�'��̀���U�!��� ]�?` �J�ʾ��� Q�h�������@f��gF�J�^@ ��Η� /RG�P��1\��;q $�Q�=E耆�
�L ɂC���`c E�U�@H����%���S#��lz� �ð��� t�e��Dv� ��+
�Q% ��a8��`��� 颺�|3'�.# �{^&"�k)N�@Z�x���׺]@S3L� ���W��B`]��Py� �)�i��3���L��a^� �.�kH>P� �=�0ʝ��8��l6U'�� ��yB� ����ΥL�����	1A����0+���p"���D��Ӵm ʉ�(�W: |�ϣ��) �!Ǩ0�h� L�ڼ�:�z.�J�����︊,�� ���,J +��)�9!� �EO}�`^ zNX��
 �-wȬR�=[>��B�?` �]��H���v@X��$�� Q����R� ���8�'� �@E�[��  �R0bS
�q� U,C�1�a �(�	v�/ �e+�ԡ��0z��� \EI?!�4�@�G:r���[5 E�Ҋ���pP��) �Iq7_~1���� PSh4 ��A]"@_��N��< v�վ�I���wWn�� ǹZ��AyhXmo��@� �ڒ��u~� ����c+��<(�@��|= XW��l  ��w
�,ˠ�_������( }Z;�B  �1���{� �#�p�I�v?/1s |��T�_ ^�o*	2
"����0�V0\h�N.�ǶR(��j� ��-��U	��S���d�BTa �.�<�x��t�^X�`����*�I�G��E1h'4��}f�A�;�c�&��#�= )�g�%`�B	(�	��Y�0�Q.հ�1E�[��P U @�R3ͺ ��p�- Y\�^�U ��l0�j *"���(�
����0��- �P5��W� {���Ah /E6��g ?�TŞ3Z��y� 1�$
�t 5}���F��2���}��L�?lt��� �dS%��� `�ꙉ �{ �01��*}��[���5	E`� 錚��(�� �u������ =��G�;�'r qy(��pStO ��,��Z5��+�����8�u 0���CGo }�X�7^�� j���)�3� ؁?"���o w	�G��i� PTIb��@��� L���1.b��YD�B� }��-U�'�rN����5#*�$� l�-� �)�@��_��P ol�h*�=9f�z����'�� �𲫞�  65&�	ʼ�.YN���� ��+½�z ͒yS�����@5ӂ��� �7`��[<���`cp�V�� ;rT	:l�L� �tA\��> �غZ�Don s��[P��h M��ꢭ�Qd����>�:'�^WbQ�!t ��)z��dn&�
�U��s� �f��R ��/�Ѻ� ��O���e�>Ä �֪K��� �|�'�p�y&�� ���X�[ a�2��g.E ��Ԩ�Z� �ᖗ,(� -#�� �h R^aj�8��G���蔩�<� Xc�'!��� HJ7�b 2³AEPf �K�Hnr<d� ��׶o#�_EL�>H� *S��뼴4�� ��:�-� }��w���!O�n�x�>	 y��D`�wl k��� �h�/9�#0$1] QƯ([�\ ��f�x��	�kN C8�^iv*;�l�gR�kU ��:#Y� h���t( U��xK�軸y ;DI���?��Π����`<2����U��$�!� \��a� ��=��cu��@���U��$��M~o��`^V	"�T^��>`� ��.���Bc,/Y�J�:y �O��K�;{��� �W%)y� �/�H�(� g��R�  f���Q� X��C�7��r
�y ph%Zt�I�`-~��Q�' ��Ċ	Y��O� ��d�� �o�T��Y �Q@n���0� �� �m��� J�-4
!�`~j�i�\���2B�}� U�l�� Y��+���14� �	�h&T O���P�N��/��i@��� $�	� �?��0� �!]��J�  ����R� ��p��A ���'F� �����en� �	`��R2��/�I�a������_+�6T��<&> ^��(%@���� :�i���"\!���G�o��J��$� 6
�m�[#���1�O���o�I8{X)�`��f� w +�,�^�K� �Q�����e�)�p(x�� Z]��`�  v1�[ R���i;� \�G���� ��f�`��� ���0XL��!�t^� ����ػcp �_R���� ���pӀ �x��] ���؋*Z)N�����bs PS�L�� �x�B��x^ ���K	 ������A� S�N���f X
9�[� ��:��_��Z����\� 40�X�^ VUQ�޹� ��p��� 0/+ҫa� �MhDJ��� p@�X [��U�̈  \Q+��ah Sf���B�9t���*��W�p���9�| hJ0Ͽ=v ��5�MW�P� A��/������ ��}8�������@� 2�)��'_X`� ��<C�� �a��1,�z�;�> �Tie)u� ��VP��JL*`Q��W�0[ب���0�H�Jމ� 5��� ���AGh� W.�g-�| oi��A�R/9�� �ٻ�΋S |N��s�g�M0��@ 
	�O��z �YGpP%�J �����XO� �&�ac� _����]d�@)O��"0��P�-r����e��ɐ�U�.�� �_%���eTZ� �گ$V \���3�X^X���� 	���<���W��)� �_����0 �U�]р��1�}����E���b������n� e�0*�� �v�M�_N� ��+h� %Y��(�� ���1�R �_��G�� 0�[ۼ� �����Ez, h�"1'I;�o�k�Y8��4 �@�婾N���@&�Ս  �\(�a� ��?B"��uh��o���R�i� +a��r����
~ ���� ؤ�J������l�$�~ [·4��`�ހ�#��v\w����΀�� XS�T�("��|@����� PX�1(� 3�F6�u�R��L�@��V� �Q�뇀�?��	�ч�F,���Q��>�U0Ъ���H��F����� �!���>���d"��0px� �'.ט�#�}���Q�o r| h���.�Gu ,;��#��T������ +F��@1$�y, %���A閳 ~ؒ)�� y�w�����h�7�_5�"�joq:�� '�%���1 ӹ�dC�f @���3 ǁ������ ���(�N.��&F
Ц)	 B�H۵�D ��oA[+� �$P�� ����O��v, ���;�5k������69�� �bZ֡� Q�
�kED �����ž	 �_"~ZR�� ��8�-� w'����, ~�@
�� �^��Z?GK�Q��["^̹��e]�l�w ��%8�� +�E�$�'~e�@��P�> ������J��z_f��(O� Z'�0x����1P�"�h��B�ۘ� V�j_�b��\�;K��C��l&�(� '�y",��1�H�.�u!�,�W_�$;��b��%�� ׷A��>� ��DF�'#�fP�pT��0 �1�3ٲ��� Ê�m@�X�p> �ka� � �)���]� 2��� @:��-�	 =�ps�+�8z�'�y���� X���P �^���%RJ��V �(ֿ� !�Ή��� _�]��	< ��}�Zbg�u9s�sU &LX"��$
h�D!i.[��V� ���ȗ>p� !$?c�f �5���/S ���.�� �P��Yx������������%�#�?3 �h���2 �1����� �Xl��� 5,�չ Pm>�'����g �:*�� �v�oS ��&���t��:�����+m��P�;�]�B؉� STw�[Q �R�n��1�+�d�ԩ�9kpH�� ����]� ��Bnh���� �KA�S+,�7�� m'��h� �%*�Ч�.��� �,.��9 ʫA4��G�J�K�iY����gX�1�)R"�$<�� �xr�-�`3��k�e� "�.�,� %��1- ���V!e�����`W�$�  s%>������@|2���c����5:p��\
K	?�H�ZB��!��&��� z��k� ��4�ؠ�0;���'���
r� iu���jK� �A^X�
��`d��@�s� ��S��	|�~ �����Q� �:d�����e>u�j��h!?C���4V��`IS ƈ�� �Q ����_� ���T>���B���z��d���� \���O�?)���
�{ ����#� Đ�bGT�� ��&���h���b逵	��QK�2+`��� [�^;�I �/@	Hܥ
5�� ��Y� pڈ�.1��Af���  <����>,2� V�A��\ �IX�'L6��� :�S"ǗX� ��G�Y�'?�? "�츝J~ R�}(r�x�V=���a;��͘� ���vDȯ<�u�G�_�x:ޘ�@U	}w�Ni�� ����Z_� �J8*H� L�6s��b��W�@�� �}��� ������긓 ��/�&-� *�����{'�|Vi�)�_NW/ܪbt�eIP�d�+ Yһ��@�0�R��" oy��Y0� #�Qh�7� �'���d�� e���P
 �<Ul��ƴQ��? {�4��1��	�� ���*SE-��������T^�%)�����`�tF��:!X��iaf &hz)?�; �yN�R�� 壭W��/�l�� �i|�p� պ�3M	��U�?$@���5 �J��K
�\�� �[� 9+�ZK�el93��"@SWF�/0����D�+ kC�T�V�> �˭�P�j �5;O�c\�~�Yݕ��! ���n�(�� �����̓�
���ך�T� a)v�h���ƉQ ����4 ����/�kb�`�_:�� �'�ul���w�.��h��� �7�*��] ����R���Z �&�<��� _���O�*� ]��k���:���Ì�&Ú=;р(��0>�� ���q!r�,�\?�u �R  ��S�xԕ ����4Ѱ �'����-}	H z�����<9�[����d �Z#�w�l������ \�Y� ����R�N� �^t�)& � �b"�v�� �!��������- �'_ǠP�(�� ���A¦xL ^�B����Z �����% �.�ﱳ ��8^��rx� 	݂� I\� ,�<�_K�?����?S�j��[�`�/�0��f�}��h�@�a� ��*B���� ��Ii�te 30*V�`� ��h�N� �w%�	Lp�q�72����v� *�c/P����Zo��m���ߐh��0 ��S����ֶa��R#�*� ;3��+� Z�\]LU�� ��զ���� �(��� Q�����=<n�>��5G�P*��rK �Q�Jڬ$ [��Z!|5 ���bBLw� ��M<&+ �,]�)� ����G�|���ۣv���:_� xPu�m:	* �i#n�` 8���	vq3z ����W� c�%.�� Q:�9C�" �[�	h@�w�f�n����� ��>h�v� ƿ��/��E �np�� #0�$��� ��Q.��K� uT��[]�W �aD*hbE;��'�.ɚd*� �<��wH|�ZŞ�%�a�2�p�-�� ��vu	" �>P�7Ӛ� �^����@�I]���&Fwa�n"��bz]�Ժ���y4:.������N��b3ʐ^�@�%��>;(� #��G� �A���.I 0�$�����i� o��I�� ~�}Y9�� "����R ,��b`*�֘�O�Att�B� hTDmK�� 0տs�� 2��^�aQ� �U1�Ӑ�! �������F#��"��W~ t��IA/, :�	�X��]@�*ĕ�������6ۻ�� �{����C �7��p.W?��XI� �X�2��@�t�� ���0�� \τR۰- �HK�	�� \Ǔf庘 E�h�a�� 2�� �Hч(�� 9������W� <���/諧�& ��`xY*Pմ� ��A�;Jp� ��#(�\k/�}0Ai�u-YT� |�d����#H0kp(� ���n����K�!��7;�\:]h���P�V _�IZ߮B ��+����� �_��A� ���{�ڎҰ� 6��$��y gHc'��uob-~�ahj4 s������@=� ��	� C����Aj;[����C��l�����G���q�8�t �0!�
�X� J9���h��R��;Q�J �Ν��NY ������:���,�]ɬ�n�v����*�� �3,gA� ׍^TeK  &��˶N=\��`�71�"���+��$�@n�6 JX�Z��/�^����]�S�XQ��  �L�Հ5�8��(�!����o��������R�*~A:� �
�zbt� V�x2��ӝ ���n���A.]t�����8۬ 9�����Xc4��@�a�\�� J��-�r� �d��v !�����}� _��O����� 
Z#�X[1� &)�~KR����%������+�� �M�a�QPz�9}��`� K�������� s&��D� m�F��"�+U` 0ԕ��T �������v� d�[�!�) �oaW��� *��I-[� 	R�_O��y�~�0��d \��˗W;	���<�
uS 9��s:�h "��%��{�	�[,���h �21���* �s��� �yb�Lh��y�&�H#o��	� 酼��*��h`�2X` Q�� �W��؂r� �N��Ұ� (�&����h �XZKU�ʍ _�L܌�~� S�T����  ��w�ψ�p�3p[��D ���e�'Z>f� I���w ���L� Qf	ʹ���$p�� x�/��d�xP�J	ʸ �����{�����S@x��y�� Ѧ2��}ٸ �K�v�f 	(���<��)�@n��[-�@ݷR�� \������ɾQ! ��20).�K �_���3 �"�1�!i�@\���5�E=���`�� �uH5q* D
O/�� `)��� �r���3^(�n	�X�J�� 0�{�o�n�����-g  U��=/;� wb�Hl�� }��T{Ru`���?�؁��>� w�qJb~����C��3n yK	���a����� �?���_�& ���s� ��`���8y���I0�p��Z����<ؔ�µ>8�����Z��& ),�
�������철���<RM@�Y%����p�i�E�D3�/�g1�S��7 ^�T�P� hm;e��HY ����S) �������X*JΠ�� �|h^x��/p=f>$�Y����Ω7�� �L!��bC$H�� �8N�)���_��]���\ QI��� /�YW��T�J��-o[�;dQ�~�t9�]�|-�>i�����e������*���%� !��oB��S� R�{n�� �/Ki��΂@XP�JN�Mo�Ә�^�0|~Y9���'ܙu	�ׂ��:�#p�� �[p
�O �E�IAV ���# ��^ �,�!E-�� 	����~�b��H���DY^ ���;��Ͽ L�/(t�>�:[��\E@�� ��J�n��	������ ����7ܩ$ qɽ.8���ͦ E�� �%ؓ�C�q>4B Ut��xW ^Q�C.T (�%���Y���c  9�2+�����̽��>e ��R�E�������ݜ�D�\�� ܼ� ���y�� - �j��cC }a[����
��&b`�Y<�X }�q��v! ٕѷ?��� 7h	Q�) ���"_�
�K�;+��yV^�wg��)Ȥ ���W#T�8*������J��R3� V還���� �)Y��	[Q #�]1
�L	-�@+ ���<T ���(�� A,��qC"���بѴPݎ ������|��;Ջ)5�[J�j*�� ����݆h�Xoa����X�D0��"�R݀ں�` z��J%
�0�+Ճ�1���}L�# عI3�J� Hxi��U� ��]���$Ҿ%�\�p���
 ��H�Ek�� ]�0ևX��� /!�����[ �1O������/*�}0"Z����. (�@2'}U 6~
%��t�}�1�3�o�C� �h-eI�#�
���Α�B� &Y=I���� ^9�_1�0��]q ́��h����RF D/�u�`4?cҀ0�	9S�>����� �!M��	���T��Q)�'4F�R.2�\,����� <Z�U�� ����ЊN�p!<w-؆q �.�j������ �'���H	
(� �1�O�� ��w7�� +��s�6 |� &�X�PN�	��� �J�`��K��'���ŏE��q��
�� -Vʋ\Ow|[a�L��� ��(������8`� ������>�Ѣq�/���=�͡��@�?>_ 8��7L ��0ÿ~ ���O�^� ��ޗh�O ���%��� ���_�}*�(�v�8�{�m��r.� �@C��a��ud L�����1AzJQ����v: �'O�N���������� �=_} �	=�ڮDaK��'zP�i��9g�y�B���&��z��h��"��C��r)�*ȩ2��!�` N$tD)�Lb<��PS�ܗ����@`X �T/A��$���<?��h �#�S �����'�% �[a`0�3�?@����� ��XZ(�5�����A�����2�휀ٸ&\� [#�hܟ�� ����X�7 �5���� ��'2�r�l }y�^@b1H �![9Z
�� �Q�VB� ���,�1M�� �PA�gVL�e KҰp̵x}.��s&f 4s�O <���&]�����	�Q(������N> ��0v ����8�@� S����c �heQ��% <mB�� ���.��ųH@� N��=_ n� �ٙx� �)0�'�_ ����o�a� �KM�V|F�!�+ɸ�� �j���'��2 h7Z������� >E.�|��zӀ��� F`]�?�	B�قC6�Ѿj�׀B@��L�^{� M�;S(K��=C� �LRW
���b�pa�(�H �fZ�&h ����B9݄ ��
��>	I d�'�_#�������0A0ịE��� �_�c3�,Q?P�8� sؑ�lɨ���r�T���z��U�艦��Y1� ���黓�Q L?$�5� � ��P>+)� [���h�N� c���7�i �_VT�� �^f'!�s	��� (.�|���d1!�$���K%p���JkW ��\�? Y �w�� &�[�D'�KQ�^��$�Z��nH����QC�!�; �DXր���`&*M�$�x_=~ �'0�T? ����$� 8D���X���c�� *�:T�<"����ik�}� h�u:3���?P� ��n0D�x� ����X !�*Q^�w  �J,���:
0�� |�ꄺ������ <Sy 1�����!�_j��( �_�B�0�� l*^�k�{� � "���-�� Ƹ���G� 0�hva�� PU�
(� �?J�,���{+L!� �Cyc ���<L���[P/���C�����Ā���H0�[��w�::���EX ��U��½�AHD�]-�Ɛ'ӟkV#����H{��v h�qQn ܺ�<��BU��0���� L&5/I\M��3u���8�Q�*܏؝�2ʋ@_Y�A1� QB��U�κ!@w�.���QfS�1`2�!K�n�H'[�W }�N|� Q��aPk��s%�z���*��Pw�= 0R�dH���@T���� ���>�� ��	���,`ɍ Д�5)�.�
���!ݨ�LҞ�} =� `���<z� h$,6b2 �U����
�������a}z$� \b [;�3�� h>���4�?�'��ʣZ�Q���l� "���	��p��uZ�����E�� V)���	X� ��
:P'�� Dy$������0�j���� +�f�$��� <H���- I���x�e�tl���]_р��z ��W>�� �Y�E|[�� 	����� � �X
��H$��O3�|�+	� [�XZ�	SU# �3W, |o4��R ��'���i �C�ȅ� $?V艾� #��N3�� �b@��d.�o �^���Q�s���[ ��Dt��R�������:\��� v�q[�k A���m��L�Z� 8y�/ �ܭ���6��7~����� H_qK(�X$��/�5�h �.	�=�i;:��O��1�����{`������b�m ��I��+��0� #ց�'�5?�d��(X�˗|�Z�e��]V����S�����y �q)"*� �ݼ�v����6�7�V��/{� �1�^A ��Tѻ��\i@ w4��
��Z��X�:�=� P�#(�3�?v8^�L� ň��\�y x��}�O:�Bl����J^� d���+�?� ��R�s��, ���<)� �=T�1���0r:� ���bV� P��	JYX ��8��)��&�a �q`!.� 2��0:V �%���" {����Z�4w�$H�[ ҟh.�\��t?? 4L���� �R����/�*��3��'򧸔 ���_���7����c �Y��֯� 3��R�_�������y5���D�����Gn�"i@���e �^�V̚� ������ �;ZR0��H4V�������")Հ�0�%����y[�� }�OTPW Ę�x$��r� �>n��R� �e�٘��	 �ZO'�zK�܀��X��ې�%x�����!p �޵X�,�� s� �rY&����\ �џ�P�}�؃� ^:��>�/�9(��R �l���� �^��s� )��	+�z�J=���-���i	 QT�jAqY&��0 ��d�FW��6֮�� O�A�R�� 1Q�)7�Z E�%h#� �>����V	�s� �2�� )e���S�$�-� ��<����������% ���q2����D<� )�`�XJ�9�� ������
Z끕9F��O��?����e ��+�9 ]�}�ؐ�>7� �Q2��.� �*��J��� �p��N-5����b��⒀C9|�3 �hgG�}VU ��xK[Z0 �R�	�
 *ӓ,���;��b���w��q9��Y�U��� m����� 	��w��< _#���D ���X�4�~���9��� K�A�U��Fb�3j#���
�� �2�:G�a�� ,~" F���_N� 0[��j^��&\S�_��� ���GP �U��/�� Ԋ^�B{ 	��@Hh�S!�KK�����BL_J ݽ��aP�.� �������  ��	X� ��U��x9������֒@a�h� [����_ʿ\z;O�A��'0�� 	��1��bfS% [U )��Pt�"ҵ0}^� �F�^�:d� B5�O��{) 	
�_f�@� KHT �� ����J-� �ݶ�/�����.��� $�#��0��)�W��u�5� ���u�OK �zN-ѥt? ����� źg�(z^-~6 P�F��% K��sw� � �V��0 K	���X �ydA� ��a�R䴶\�_ ^ǒ )�V����	e�h�3CW���S 8�yLV �Ѹ�t�H= 9;٫�]f��O@���@<� ����nu ��B���R�!����X�p0Vb 
]� ����e.��Q����d {��h�  �OX�̃�' q������i �t�1oY � ��H����_���Cdk��9f��� S� �� �� [J��&�x X8;_�t>�=/�&�� +[ؿa f�!�h६�N�İ����Ab�h	S����z����ʅu �v�/���:� @��Nļ�!+�4`�%�\r"K΀�q�O� ���0��z�l P�ø�_;� i%3�ce� �.�=L�N ��r~K� Zݩ-�V������/l*�W�r �+�K��N Y(�*�v����������H ٺpAl0<�X�� -x���&��p ��Xh� I	;�n� �����R 0�-��ت���O:���p+T� �� ��\�~���yh�� k�3��]'�����;�@�F' SH6PQ��� M9�T"� ^���+��N� ��6(�1�*�Eg�Ę���2 �K`�� �~s�1�X Bh�S��y a�~�/�?�_ ���}�>��c�)����\���:P# �I9)��X� +Z��� K� ���[��� VQu	��T��Y�h���� 
S�ݹ�ڃ a����R ����!ʁ�z˃���g��a��� ��
� v��f [S醤�@ �x�hU_ d�-K{!p- 2�w�SY�wܠ�٠��� "v<�{- @*������]_�"�"J����>#@�.5a�; ��	�\g�-��zkV��c{ Ƅf;&�� �(J��y�;����h�c�]��	 9�j� W�p @��T+� (Sޮ� ӱ����c`��� ����X>0d4��؇��B]���� 0��A���J���	�`�I ��o�(�`���y �N�A^�2�] H��ž���a��1�З���(�*+� 4��1���^� 0���� %����N��1�p����� �5��_�	/��� h��0.�,$ ��&��s�b*�!�W�q7@��� �]�X�;�s �h.��1\�{P�(��*��� ���Iǿ  �����p� ��:�U1�S ��ڸ����0cKd�� ���H�;�XQz k��k�r$/�6 B\Sw�bW�c�^�~�<�Q +�r[�L
̈́�$  �W� �X2̱?щ=�� ��n�Z����v�'!�ty �-ԁ�.$W9��h�	�	�/��|�YȦ�NX�� ��[�1�� ���@���?�Z���0�Y�7U|D�l��cL�� 9�w(2�0+
�x���n�@�"�Xw� ���)�UYu(s��_@�!���]�@x�C �S4n֚�I ���; ��Z ��h�L������D�����(މ�
�]hP�f)� ����jp��Q# ��P0���.��('U��ِ�;^��<�	T�0
�L=:v���)>��� �ǫC�Tg{���X�~+Pp��8�y�d�/�Apc�ŀ��*=1���!�4d��U�@��?�����+���zط�Z�	�;�T. cT���.�t� IrV��� �	�+�-�!�׋�`�XY�]ӯ0����� ����E���r�qO ��2���'	��t���O�Q]q 2@%���c� �������J@�q��ĝ�o$��m<R"�W��� P j}��� �5���Ww2 ��hMy`d� -���G#�� 
�\sM�	7 `?��e_�u�!��i��>��.�-@�: H
�m�<1������ %� fޥZ{L���.�� ��֘p� �-���@mhOb6�n������3Ϳv�pG�\ˊ Lʤ~/(X�,��`1?"��}� � �@U V-�`(�������P)�q� �Ǜ��!� �O�̭1��-��_�c��xӿ Q����Vv T�"j��X�.qM�됋D�N:��h��[ �
2�z�x���\.cB��h���' (�� D��q��
�Ń [��Qт.n 0�JF�5/���#�8D�,��I�Q�����B~:����"J)a	X� ����c}�r��c#T���  ��%(������������q��� ��H��� X��5�O s�[4�~�0@b
 � �P����, !O�(舟��`�O�� d�|v�	S��@��ߐ� ���C�(�S������� ���:2)QI�\�Y� ]"C�@�1�� :�ȥ %Zhsz��ى.o�0dv ���GZ�0�
�!p��IO �%f~��	� S �D-��Y s`�� �v	�_u�j ��z�4�|,�� ����5.���>`������/�3��  m=�`}� d*�^ØB2�W�C��� ��&(��c|M�
�U3��.��e���	�� y�9� G� xRP�» "Ԡ�K��@ 0繎\��?ɀ 	߁p��$4�"����� (ig��y$B�^U 򧢞cV�: ����	)���ܸ;KVt���3� ����W�� �4F��)j��< )}d�� ���B��\ ɂ��%��� =����1�l	'��)��r�> ���kU�Hc; \'���+� �n3��7��W���p?� �� %�u躞XL$��-v��� &�7Ąٮ%8���(N�1B
�,H� ��!��	z� us?��0� �����p ��鳻��b��E��1� 	�����% ��̼�H=dlc��w�9�X �:�.�21 �^��a�3k )� �S0hdG�4ٺ���VD �<��Z�N �W�XU� щ�-��s ��d���	��
������Kuv�n��LO?� �I�)��� �5w���Y��� �ClT�"�z<Q��A��4���xC}��	���������_�Z̠Y�O��|/ 0�\���o �!�R� (�;������:�ڠ�	��� ]b�QSΎ ��'J
_�l��ķUՒ^�Ѧv<�Z�:����+���h�)�bX���i! �QCO�
	��������� `8O���	 h��/�^�`�}��H��+3�U�MO���� ��� ��QU �w��Z�?� ��k�M�B�:Q��l���%��|i3�DS����N� ���e�l  �Y�r��o��H����Ֆ� ���v� ��c�U�1��8�p��^�C	��S�!<� ��@�3��[Ќ�[=�	rR�fA ���'�,[? �&�� �Yba�+� [:�cf����s&��0p��X��
(	��ڥ_ ���� ,�Ӄ���rA�h�N/��;�(��|�Ɂ  ��;��N� �X_3��7 BM�<�b�] R�4zg��,��?�HɛP�� &[�hM��\�� rHK�c�bg"�%矋��Uq��� ��i��:X �b�j�V�S�1{����*� �[n�)�x� �}jt��.� u��Q1�k�F�K�$���_ ���I� �>��!v�BA1M;��. sp��� �W�4�Յ��&9 �Zl1:L X[p����,�Q 	�ϯwlzP�ـY��I� ��|VA�0� 2�d�ի���Q�Ƚ�/#�`� ���>�	v J��П��bu�`�R�� ��CW4��_Ĕ�d������ ���aB��n ޯ6�d7�1�A;	\��h` 8����Y D�_(���` �0�oOѧ����-�^ f!�mɒ% T�CZj�	�ٕ)�F��� �m���� �Ү����� <L +F�� @(��b�Y�?���Ǔ�����Uԗ(XC�,�����sQ*� ������a^�m �ӈ�J( ��
 � v��,}�z|�^8$�F�P.�[ Z�封p� ��q	Y����[�`��ݼ��2V��*+�EP���r �l-�OÝ �jB���� �k�#1*G�\Q��ӹX@�� ཁ���S�;��j��R(� *s�
� :G��q ��� 4WĿZk� ��1�_p� $��&��Ň�^� _!�1�] �l�y��� 鑏�'Z� 1���YP4 H�*����� ���)�
}�-�u�pI�F�h@i�}�
PB��K/��3�=ZY��~齔����{ =3u�OR pH�5� !o$��� � ]꿚asS����*�<�-&�W���FPV��P �>��-�/u���w0�	�T����P��� s���ݾ7/GM�R���( �F��d�� �IAz.1Z�� &�6B| ! ����Y
���o��Q�P��[ =^��R�
-���C�u�&���+ *|����Ah-��/�C@���$ ߽'5�I! 2��ǹ�� �0E�>ľ�2"V@����+0�(�B� ��|��0a{��>�(��_� �L��8� W��/� ����@;��i� v�OE��� YS�P�z�o��0i��@L��'�e7k�|��36KN��]F@V=�)� �py�
e 錇�X�S�+����Ex� �
��� �_4���� sA�; �@ۉ1Y^R�[���;��T �]0 ۃ�<S\��*:�� �%0�,
 ���9�N  ө�L�� ���D�8�=CP�V(�`	��� �z�A��_^�����$hn6 �/K��G� ���
t��N �čɃ	)��ga��ы�' ��<U�[� ����kfh ��nL�P F����� \��H��Z� Ö���"�� �Y�K��� �!��6 �����)7� \�R1`�#�[�����6����w�7���ŵ ؀ዷD��Ӻ�p����>̈<�hP���� yZ�ͷ8�3˟�)�(���	�\� ���}Nb� ���'+�]����=�m�_"	���/ �����|,�����؀K ��N��Ws� +[��q^d����8�`��� ;HD��� L?}X9� ��h�5b% _r)�9R ��&����( �l��=!�$s_� �M-O�H�5�)���$ &��0��L*9��g���*�� ��B=�/�| GRvp,�	� rf��� �����ڙ���R ����=ỲfcW��>rހ�CHā�/h��S�0K�q ��+�� v5�@Ճ/� ���Q4��p<�J ���n�~�#��)���k� r�b��]�{%�P(�����o����h]=;R��p��������9 ���:� ��?� T�	"�� #��{o�&� ��m�� JE����� �i�ٰj,�@ܗ�`�*�� �ԣ�=Sp�%�PV�K���i<�� �J_F~��(�!��G�X (��7�h2�bQ� ��×]� �4|���r�?/-��́	�5haN����ꝖF ��հ�1� �}6�[K ���L��9h���,��p"��:��h@�� 0ֺ��3U�{�� �� �0 ������u~[�T� ���Ns�&����� �{��Y׻V	k � W��e*t��mO�����b���6BoeG�� ] M3�9^W����`#P�H�?���!w/��AQ�+ʑ�Y{�i�N偶�� F"(�X��	��O�� �hj�� �C��	%�X~VS��:���p���Y� �jљ�q� ˧2�h�r �-�(Ժ ��<��"� �� %�����IDԱS���γG����[�V	� �08� �� տ~ZQR��q` S�'�V���p� _���	s� *�H�Ng��u��d1���X�� �"��P( �^��İ �����#ͰA h�,"��-���٨ �!H �#X)�>		��~��i,�@.�Y�A ��o���h��\�=��@��+�3�ZA�IG�܈�h�`����[� R�ں8�� p��kW�^ �� Z�Yz�$��@ė� ���Zh�P/ �0@�o�{������P`2��� l�����| �LŢ��{�q-I&� ��.��m 1�
��D��k� g��P�0�Q���S3g[,X������ �{i��� �n���0� h��3��uۭ��8 � ŵ!�"k)��� p��+�<3�,�b�B���� R��8��e= ֙��g#(�E ���
� ����sY�ݥS dN���>��,�`k[n	�� ����\#g��CЄ��BV���0ߙ /;.ٿ'%�� �����@��}���J�t ��r�(� ���/���� �6�������Σ$��'�`y"� �UV��� R����N�2�W#$j�@��Z� �n�蓌Q��|[�"XhTm���+� dǃ2��� �!�6"����"���@��3�� 7�9|0òK���PX<�[�� �g�h :�!�~q�;
ԀBЫ�TQ�Oh�!�WR��@8� ��vP�b �T�z�� U�e P�n�c[�Y�@j�6 kn�H� W@��*�]������6C�	��@�_A� �R,�YX  �O���% w�_��1� ��[h�~ (��1�) �d⨉�a[|VB����p�^ �{�/���(�Ōyq1�~�B��6@3���K� Y[\����� �����6 D�(�7~�
r N:�ߔ�<�� ��Z��a �DjW��� �K��2[� 4�~�m�� uL�����,�e ���pF�pY��C����ă=� ��Sk�>�D�� �h_q�Af1�B�lp��?�T��p���p���"<�Y�����b�| ?)��&���\�- ��n����/���c@��'ڰ}(� �!跃' ��H�b�� �[גo�}#~PP��Ws� S�X�*l��-�^���lh� 3(�B߀�&�rZ0� `�-k�t} �Ej�dYu�\SR>"��� ô�� ����7�)IJ����p?OG�߶��� 0�X1�Ӥ?�  ��j��VT^��Z39,1 �*��Y���}� /��sM ��5�x؁) �]�i��>^���\	���pu�� T��ѾxQ� ���L$�O�V��@���^N ���M�K�� ��x)�h���� }��!J)�k�xS|R��o nK=@B��� ��%�4�' ���@5`�#��W��� �����A\�o R"�;I�2 ,Xz���� �W����� �9��\���J��YZI�"�K0�f� � ��g}�RI�qj]�����lb !���B� ��\��*�Q ��ڙI�� ��0�Z��N 9�����@r �[��zΰ���� 50�>[w
��J,�^�Dа��� T���Cŕ� 	�q�[Z�
 o%��i�]:�nԀ�B�(sd ��R�p ���ӌ��  W�V%"ZA 5�`���X  ʷB)Y��h�w+2\��_"ZC@��RJt@�_�[��{ �܆��E�X�:�˰� ��Qh8qu 505��,�P������:��0W@�Z�|���@�L&�=Q;č�]B�۪q���*���k���
�;��xӻGV����	��� ���i�#�^��ر���/?��� �D�ѝ�� h!%�HK�>N\��ȿU� � �&A93�F� Q=Z��8:��a����2���|Y �|�B�� !F�EZ�P� h�z	q�>��d ��4�`H	z? � a�ԅ� ��(3^Ȧq��hm\J��?�=K + �)ض
� ���	�P �%1�b<�c-e R)ź�o���`[ �/� �P��ڤ�θxƫ0�	���r ��]sZ2�l^ ���KL �E��1� P���Q��t���������vH b��A1iU��(t� }p�̾�	 �]I�j� 3y�
�Rt ���)%K���2`Y\. ����|S �;�8}Yp3��� ^�l���+R��<�v�\�F ���0�1�&�[�˧���{� A�#� �:�y
 )P�r>���"�p�H��`�� �
;��D �ї�`Y�S;�t���6K��C_zϗ��TY �	s��� %����vƯ=/�h�� Z ��D�,%_Y 57H����� �̃拡W���:\R�$�q�!�	��0[� ����u
� �����X( ��3T~H[& b��9��N �C���L��%����5�<h_���Z��z!�-��C�ꠙ�� ��12Yx@R����J9 W���!z��nR���r��y%���X=5 �[��4gh ��J�wZ ��n)�x�P���/��R��] ��Ŵ#� �h����aj�_,y�[1����w��/�$ �f�K��(� :��,_�	"?=���BŠs(o�� _���dJ% W�6��2Q ��N���
*o���L�_���g��J���`�\� �N�|ɣMS �����)�H�����0������E� ��Z���8(~G^0s!�\;�,����@Z� ��B
pn�:�� ڑ�[R�v �ԏ/�q!��plA���0 ��[��F��W�G<��S Y�����JB� ����[h�	 ڹ�����|=�H �5�2D��K�_�Mx	��
�"�.�� �V�n�R��h�v~�j�@��Ip�,�j ���������l	^����p�K�� w�zD��. ��Ő�� �꓿-zOr��`"���G)`�pX�/ ~��	��P i9��2� D�����9�_�@�[��. w� �P�G����x� ҩ���&�� ���z�Eh�O�(�@��Q���{���� ��	�L]px1^����l %k�E-��V����T���F����s XȬ��ݮ � O���+0�	[��# �' �PhO<�J �ì/���}�1 �Ш�\V� z����N F��v0�� ���J�:Z��L�$�0	#� V�ef�Bu� ~�����{� ��Y��E 	�!AIZ:�V�����p��Gܰ��`d \�0.�����f�W�@_��J� �B���Q	 Ӿ����q�,��s �H� ����yU�A!R �ݺ�t� ���X��d�uE$0� O�Bï��� g��!���� 	}M���'U ���^�ď �X���� R����Q�]��>2���,0�����=���|��D� ����ј��1	��w >���C� �2�����p7@h�d;� ���KP�z� �6��S�� ��v[C�(0�"B,!��Y'�\���� �{���$�'	������y6:X�� ���<J� ®�Hp��% ��č�b$} n涤7N� ��5��Y����'hт���KU -�S�!L� ����Q*(���I� Z[��P�V����CX0�
 !́MU�I�>�} 0'��T��Vy"C�+�I� �f �_����-JA����}$ !O����/W T�H%[�t� ���ځU�� �{�`W~* �t�Sa����/�,�����QKX�C�  1ź�<� 	�x�\Z�%�tj8��� (�g�'#�I +o���{V�	h]ݔ̵H��Y��Rౌ�G��� "���:}� �[��x�J PQ�\'y��t� z-A���;�r�%��o w��)}s@ 0ٟ𨷤� (�]V�q� 5+m�>�& ױ�C�O��r%�b kW\yQ�-��S: )2�=` ��Z�p�P �jݬ��3��.�: ��� &W��S ���hP#��f��� ����RX�3� pa�� @�5B]�� ��^7� X�_������\]�q���J X�}P��p�� Ή�!�>�[e� ���8����
�M L�`
�+>p��h�@�S#럘 �M.��\��#�� ]�HXyڿ` �������F���0s o�+��� �Р�{�F�O1?���&���C�5�-Zu��
Ƃ�������J�5��٧�` ��[�hY ,-�P\�N �Ψ&3�@����ԭ�	5A�0 ��^�R bw��(� Q0��x� �p/�2\� ��
���� �+�:��_>�C���ś!T  �jB���	��h���8� "���!��� p�=�D, ���
���~:4f�� ��]\���(a,ֲu���� S1;�A�vjv% �]:�b����[`�l_���)� $Ӡ0�U� �l6![����������]� ȑu,Xɸ r [!�) �]�F�PmD��^Q� ���!�� �c?i�� ʙ|R�*�"�%�� �] ��z ��r|Q,��>Tb�e�` �^��1 �ݒ!,(� &�JuYl�p��sh�/� R}�,�oBI ]{Yǒ�'��/ TAh�w�d K���p�18:�<@�0�oE�[��߀��ԅ �܋w�b�� U*��M� ��RO<�| �76�$�z`��*�	8�: �R� FV0mK��
 �Y����*���O�/�1F<� �����(�\��bpo��Uŕ��탉���{�^ p¯�uNV"� ��U�^��q\�"`�� ��c��Z�# ����
�_? �4hs^cgO �E���� ��� N�2�� �)Z���� *�@��pa't��p)�*Qd�|0 ʹX[Z �2z���U @�Yk؎�� �Q�볂��5���:�� �Q1о�>���� WE����Z= �N��O���1 �Y��-��i ��0S��H8J[��0a�(�ˉ� �MJ'� ¾d���� N9B��O��(���,��AX��uw�X����@���H�z ���2K�|��q� �ŭB�&` �G�3�R� uS4�@1 � 	���%� ]����\N�� 	�X��nݍ �Vy�f�* �]�%Y�J�< ͧ��n�� .�]&W� ��ڼ8$�n=	����1hc-�{@�V*@�f�P�� �^�\����V��w�SD����f��p���Z��� P*и��!X�@ ���yX�� ��$��-$v 3[���N �;����k o4�*����F qQ!�
� �(��< m0%��L���3�p��uy ^�a��L6�� ���� P�0`�ͽ' 1zt�aXR� k�?�����"��q�j��=qA��P�����Z� ��,kT@�:�- p�K3\Z ����� 87x-��Z ��JP��~<A^���{�W����� �*�<8� K⟂��� ������Pv�R�{�1j�p�
Y�*�Z�� o�G��� ��/���T ��"���Xg{L@'�������2�S� �R ����,}�\)��iA�z��sN�� �X�O�y�<@���&�%-�	U�|�g��GV�o ���Qka� ����x��� A�/'eBF!���g���~Y 0�ע��)e� ��2�1
\�Q %檣I�!�h�?�; ����� &Ԩ� �U3� �J�ɰ��s�� W��p��� �܂��'�U(� �1�Oc�5�p� �f[Rغ*�0����g�?^:�O ~)P�L��:� �v	$#d �F��"�8�c��S$��X%xȺepU�)��uZ`۝�p��J}@�VRwe����;"� ����7bN��A��P ��ʬ]_� �B)R�8����e-�D��� ��G��S=Nf��/ �	6W`�� *�~�op���x@X`�[� �9�$��~՘f}@�u`S�� �)_����h�d�Ł��* n���Nehry	
�F�0)� #n�~��W���[hGs$��`� ����'��?ORE� 0� z� �N�฻+.�	��إ�[Wp� B0��1� >�x�_�p� C]��U�H/ ;t�!q� ����^2d1���,�΢���@�� c�J��2� �h'��}��C 0��t:P�s,	��������(��C B.Z��HE0��<�����0J&��e`j� i	���� �x�3�� -�j�O��# ���qt�	 �߂��.�0-Y�K^
�1h�fP鴒<�	��� �bd���H4 �M�U)�KZ^!����a��� \`nh��(�O@�Q���?Hw ���UJD� ���v�2�'b�Ï�pO�p�	�� l#+���� ���[ �k �H0'�՚ @h�4��� ^f���X' ���>�ya�W�]�2�` ?_��tU�h �m����� ����P��� (���O\�u����S0Xݠ� J:��i� p�4�����WHK�L! O颷	��
�Tp�� �8�� �<!�Ĕ����.���u�I���[����`Ǳ�m�e{p��n%�o�#�i� Ղ.kj1���|�� <��&wK 6��,��� "�x[�ݽ 1�-�� ˲�,�PK����:��ىp� b���>ֹ 8�`��;�U� P��H ���ī�9�W�`u˫���7 �,{*�Ӝj�� ��h}m�v� 4@*���� ����2a���v�� ���S �����?�)u���%���?c �	ʯw�j��� ����*��� vէ
t��8H�@����5��0�k�>��)�#�pmŀ�ځ	<��l�@Q� %B- ��~���m���� �3�h�"�@oB�U� a���:/� �c���<8 B������%��9
� w��H1�tKN�S�����O��L{�*�-�z����IB 1���R[���D��� K�UY�[�B��(�-`���A7i���zT�(Q"@a�r[ �MIv/�t �
�ϋ!�>�р؇c�	�y 8A���>�� ,3��\(�� ʃ���U�� e���{�gD��ϛ�¯�_�����1�%� �pJ7��K�� ����@�� ��(�	��[���0#
��&�MA �D��_P�]��/0�VF C��{͛4 3ٝlZ/!�%SQ~���q�`C0��$ ���a���X�����`7�pN���K�3 ��������o/`�4 ��61�� X����
ZR ��P����,��V��Ό ��z�15��� _�� ��J��}K ��nr^µ� +���U�N<=zu r?d��\���E� �C �-���s<YU���hI�� $3��(O�� ��>Y����}�QKh��۰%b�1>��lM��"��� v�p��� ��"ʗ� ��أ�o�X��`h�} ���wY1L��Z�����n �JQt������r�p��9� �޸%��R� H��K�j����I/�
�� ��Q��#�� ���1Y %�,x>�{�	+��� ��H��_�@~���CӰ?��8[XY����P �ݫ�VDi�"	�wz�앂��f߀vy�a�8�{����P�������� #��t~���ۓ@L�k� ��	��d <%�P�x���z3Y�Ñ���( ���O�H2 ���X~&��	�؆6�) <�(/]��#�	 Xh�jR*r ��D�� �٭/���,>�)�	ǀ`�� J��0c� X��eu �Y!���4"��@�K��ZS� ����-=	b��eX0� �].ɠ��	 _� ��\�^$q��<���(�p�� ��R �^N�1��;M��U���� D����_|F R��IQk�	¾�� j��H�=�x�-�P/��ϝp: �a����� ȸ�#x)�t� ��i�&޷ �uL�.�=2 )�P�v� ^�$1r�� ������Z�@ �0*{! ��X[��h�QF�?�S� ��� ��) _�8�`� �hVs�QO �0��8BN]��A\h3���( PD��,e��B���/a��~ ��� �v�B�[� $�qQ�'F��5��`�h�� �t���n�E���q���P� T��8Y�$ӰK� ���,�zA��� ��>�� ��af��~ \5�`1��jOƪ �]	�!� AJCz�� �ِ��*X�5y@~��$	���^�bp�P�ʢ���Z( þ1p� ;G>��� �svK����Q^+����:���i ������6 9��P[� ��(��?ٓ�Y�P�p��p� ��\��1� ��%��'q������� �{��x�� ��* ��%�A�ƈ�z����L�/`f�
�럿 <�(��P�Xf ���}q2�.��� *#��!	 Dd�i� [7-\����	��� ]8V�`t �
!�<� U�S�"#2tD�Y/ ���6h ���g�%�P �Y��}>�� G�6{=!�~�� �b�^� -	*��G~%}��I<�N� �1�^��' � �uQ��G :��¸2r t����kf XR[�GPs�\�;&������� �U�� V3 P��hN�� 2�d1Q/��=���I���D��X�5P*������ l����s>�w�Y����������0��&�z]k�N� ���n�H i�,���� !Օt� �>k��N�.��b���Ā��S92ց��%~v���i��Qw�C
 �[}Wqa�D
�A�� S�m'�[ ���X��	 s���A�i�h���+���ʃ���z �!X�X8 �=c~���_�
�@�P7� &����"� �kvU�܀t�&`�� y���� �ާc���� Ϙ��R	��4Њ�����o���- ��
վb$ �[���0� ���x��s� ����z� 2��ˋ/[��`U�8�7W����A(�&��� ����� ��{W��2���zZ�0:� ]���� � ��c�u�$ "�������0&�O��>��( Nՠm�'�[ ��WFٺ@ �Aw��%"�:L��3�򾰛$�����YZ`n};��d �+�h䶀� ��-J̢:�xX;�S��o�$���B 3ވSP(�� ��Q��1�C,drd���� ��D���I��gP�٦A�l� �r���d@Y��ᨓ�� ��!��梈ఉ �J��v�0� \�*�Ah �(�)�`��� 0�6ڀ��r �][�x��4<�܀7aJ� %B����
G& 4T)��c ^܁�%�Z�JE�V���@�H����7%�9X8�����n�`���vk 3S+�2x~?��Z��(�H�z= %|PH�T����^���àW�$ K��@	���vC`��\ � WP���ȇ�?�ʀx�(#�ߝ �m��� �W}Aa1�_ ]0�u���QX ��/؋G�� ���MU�� (Ŧ�u%,]�� ��D2�rh�a�<#������ �]S�Zr �@�"�� �����]yZ� ɹ	P�(uLU�vN�E� ��k��2 X[ð.��} 񤌧���K �J�n�x�	0߼ع�# �関û\� VQ��1��Dy!˹��>S��t����<@�<���P��2[� ,��;�� !ܺ�(�� �`��y� ��˲K� H4o?�� �'u�� ��<�߳|[ ����X2� h�F(����Ni���
X�Gu �";���� dB��� � Z2�[�p�Q �I�X	���t� �B@c�� "� ��O��`_��X�/ չV0�[� j�֏*��� ���P1� ��(	p�!b�y�Z����ĵ }Yɞ�c��\7� ���`����׸],R~ ;$�r}' � w8��N^���%��ppl�Ņ���d� ��?I�	T ����8 �0��S ,��H�] ���D�{��ħ\�3�̸� �O�K��� �N��ܣ�5 �s�O�g ���)1�~���%�+^�B �b����� ��-
�&\Q��� ��>.� �b:HWd�P��a� O��	�Z��Ƅ�� �%g ��\����)@_(U��� �ɐ�k�$	 {��_�>� c����30�n�&X" ,0NC[#P��A $�^�������Q|� �#̰��z��~P"Y��k!���L����A�Y�@pfU'���􍃂��෗�*D<�"��lq��%�ٱu .4Z� ��iO�;� 5��V!� �lp艕�� ��Wԃ,�3� V(�p�z  ��Ȼ�'�Y.� �Q���z@����� �^�`?�5 �_����9 �]�r� �'�b�
 �v�V.G4�w� DڪP /X�y�l� � �@4+�� [2�hI�x �t���+{� ����l5J�Ȑp
�W �ɿ�����Qc���hdao�u �5T���l)!���`�B �]��A� �!�`�f�hX��Y'��� �~Jb"�u� �e��������vS��ͷ:�b[�.	�-��^e��0��I��q���(`�d�d� �T�_&� � �F%/@xq��� �hSz�g �3�/��; �ӁR� �NZ����  En���!z ���4��r� ��X� ��^C�*���@iVU�2�ҕ�Pˀ �~	/j�����b��< ���$��A���p��T�@�'(+� �2��� ��>� Z�A�� ��F���>S��H�#	�7; �)�/a��gn����ƚr� �cUJ`IL+U���֠p��q�ynV�5Q ^;���#b� ����( �֒��P!�Մ�"@깇 �ݶ�>0J ���u�1"ɣ���b� �O؏���
 p4��-�D�M򔿇��1�._!�;*��p�ZLw�x ���'~6	9�4��d�IA�:��p�! ����)�U +O݀X,���� �=�8;�e�����j$�ƕ b�������3�F� ����*�4	-^��Q&� !�XE<���IqO	��+��9-� i�	�[ �V�mNҫ� 0�ht�ZX ����8	�,��^����\�W#v騌���0��!EE�*� ��� ��-w��x���pT� �1���=� 6{��OS s�
�u��/_�'�U5��@���~AG[	�٥ �*�h�y������������  ��^���#�Y;��rQA�{�x�o��c�� 0/���LN� ��.�@�\ Q	���֣
 IP�y��ŝ� ���R_q�� ��И�?� ��
/�e�ic�}'���!��M�j��7��<�l ��.R�U �髄F!�_� �i�� �d�'b�� /�\�}	* ְ����2�V����,=H� �D�q�k _�(8-�O����1�3�Y�i\�.�u��=�� ��(1�nD} 
F���Az�h�(� ���������o�BFNc�� � \��4Q_�~K ��N�/�)	r��*���d�xY ��&�I����5��@��1 �t���:�� 	�3h�J ��Y|.ϣl ��쌺�<� �����f� y������ �b�up�i� ��3?k� Đ��H;U[�WQ>�qS����	;F .(���5�*Q�R��YO� ��
�ת 0����	H ������X(=�@�Q�5 �����z�n8,�[�:�&�� R��p�� ��N0�(_�!w�-@�8�U3�=h��L��� %-0�>O� Xs��5���| +,����h TIc#o��%��l �=B��Q��v ���!��H[� l�W��{|�	 뿢�'�S ���`�5< x!��J/ L�6iAv]�Hk��^B*��N��~� ��+�o�K��;ظp�,�r !`������ �{�}f�� ���.\��V �{	T;$ }�I�褐� ���Q��~�K�%𰩌}� 8��uJ ��<O7�%� ���C�E� �Q��1 �� �mC��Fa���zI���P����^{��� ܁S��,�&����U �G��YQZV������iw�j�ڪ�� -)Td/v�k��1�U��� ��)��2� x*�Z��� ��%��1[� ��0@��Nk<�q�A�?�K]� @��%,��  �~	^�_$����K[�;xʜ�/Xw:��$=�>���%-�����`��v� +���Z XQ�:̥� �����KB"�aw~t��7�lFR$9�cp�� _�B���2V �fʧ	݁���>�pu� �`8��ס��@��,: �2]�Ώ)��꠱sz�8�5T���u�q�� ��_`�~释@nS#O�'�{�� �	��WE ������- hD.����� R~�_��)�I�[=�B<�r�  �n��x�b��	 �ݹ)��~�Q �wydLR9�i_�B��I@�h� �\�kZ��� �i��|/� ��-R�^� 0�Z!�7"�~%�X	����Ξ��� 	�a;����#��N c���+ ѐ:'�)xC �{ �!��|���	p� ���.���S4�#�/Q�_E�m1�0OkfM 9G��� L��	�����ދ�-�g'{��� u��$K�%i�@N��$ �^��� ,\P%��_f �˸�o5h^� �?*H( <�-L~����/�%���6.�0��0(��u ^��1�.������ ��X3J%c�=�������
8� 0�%�ea#9�RO�K	���]� �t��Ԏ�Q /Àh`�
+���U�[�� #����"�>���%��[�����ip���d��� �06���# �%���/� �a���j�2 ��0�Q
�� ���>�(	����X!��zfXy% ��C�ݵZz S��;��"Ѐ)U �12�*�l.� ac�+���rB� ص�R�/%���7��g��Lz`w���@���l��-xw���-��v����	�IV�������Q �փwW��jFT'����"P �BO	��h�*��� ���[�@0�Yk�2�@�F���{�u�P� ���f)����� x"�Q^K��@,����4����͘7uր�1�(�����ڇ� �@*���b[� �]JQU�q�.@���=	u�s�f����z� [Y��$�	 ����(�� %�&�!�
�:^> ��s@� h%|<䨰� �8jy'd�� lhK�>����^�x3@(���" �����b �@țԚ�����ٺb���Pq( �1�x�J��?!��+�M�K���_Da/@�/�` 21�h�<f:J� :�wo�Ƹ4 Nm�,�5�� �_���'�P z� }[��� �*�_v� F���$�k ����&g� y)ڽ��Y�l�K�`t�� �B	�9޶AZhz���ǐ�0��W��_p��iRL �x�~���/Jt ������Xw�} �&dМ]� #��Nb�l \%��VnL !J��d�� eD�½*� ��`����� :}�'�xU ���h�e,�< ��`��  �辤�� ���@2^ ��q��y�d B��Y[h{ u0��f��&ŗ��n��� 
 1�S !�a��� ��KYI��� +��V � 5a�k%~D1���T���j �0;B?Y �3�{� �D5��������>�(��'�t�.�v  ξ�z�ډk �$*��H-�lC�'Ѧ������Y�)@Q���1 �+���� ��`��s
� ���?�a ���4�� �p�[`�d����t� t�N���R� ɫ���(6 �!�X}��k|	;Ջ���vt�A#� ����T�$ �W���/`+�: Ĺy0S( �Z�5O ���'�E a�>:t��N �1)��6� ����� �N�Gn�� �I�c��� �>|�6�J �
�`��� ��Ai1�� ��^��8*� �e�KŷBT )@l��\ %������J8�Q��R����)*����� �S Q��U������~^h�Q�� `��R$��� l��f��Y��)�-݅�9 nS0�:f»�N�h��r2��ke��R\�8�`.��=А��W��1� ��g��S�� �O�z3J��<E+ ����7 U�n����C ��;
�P�	�iz܀����s����y� ��U~	r�J�s����Џ�X?~��� �	L ���GZ�8�=�K �=敢 Չ�w�u��L&�N��Q2 �iB�!'4�<�U�`I�}�bE<��8рl�%��y TGϐ���=�u�X�_�;� �3�j��!n�h6ؼ1j��� 1�5$�YZ� �K+�Ҋ ��7���u- �X��n���T�����0M�l�'j�K��@�V ���X^!� ��&�"� �d�� ݇��+��� znP��� �ڂ��R�^�z}�v%�p)�@ a�,Z��� &h.�{�d*��8 ^U ���j�,����Y +��;#�^���O��wXe�ݫ<����9�0	�h[��`�܈�a @΁����� <��0�n� rN��KDW�:�U��X��� ��l���[(Jظ#��� ���Q�� �@
�J^ �w��~N �>��!��?�� z֠Õ"J X�5��h�E��T]��V�`� �QF�:�9���)�����A�w� � �м(Z�;��5���ԗ�^h�%s@,���) �^9�y�_ �i�r�'`�A��\�2�R�n��}	0��	��^�V�� �"Ɇ�<bÀ��&f!�� �0��#�K:J�s �Ҥ�!�� �,��A�z� �{�#�I �vg�A���.��f���% �E�@�"V �r=��/� x��w>�� �PE�Y�� 0�� �X� �-	��C�1 �I9��AUV(��^�� �퀁�P��?!@�_�� 0���Ł �"T�	`D��h�3� �� �/Q?<��� �h���S��o�n��!��͗]���j�m xIƦ��!Y0
%���3L���C"��� OѢQ�0�"?p��������-�Ya��Hh �&"�	�(��=� ��*خ��1T>@���'�|���}��ǯ��4U@[�] ��ZQ#�k/�x� ~����I� ��$��5\ *�!i�4{K<�ʜ���+��1k �_:�Ӏ�°z�[#�`��!e���T+����P(�<��L�ā;&� ��_� >h	�C����`�؆ָq�* �RM���!35��r�& t4h]� P��ʡ�0� ��_��>P� 8�|%+� ��\'��ܫ xU���iI ��c�1 V�J%��� I���aH��]�0�x( 9	�[���)h#�Lנ�~<  �|�!����K� ��h_�-��L`�, �8O��'3 ��Y�k�1L��D _� B	�R����$�� �J�ѿ�
 a��� Z]�Iίz� �TԧX���"h� �v�Sp� �Q(ܹ}Z�[ b�j���69��)��h��X$�xz U�� Y>�/R�� o��`��S	O��K���9�j��� �4	hpc	F�C ��� �7��
h�ze�����+|0 �)��%4- ��S����y�8�/ & ���ϒ{˳��ѥ.1�#=��8SdT<B������銰 D���Z�� {s�[�~'�)!�	�� V�e� � Ⱦӹ �-{�q��
{� hFς��r@$Y�� ��M�E�:�����[J*�K�a ����Zku��"�%���ŀ�v8���!�hE'0�� �[c���ް) l*-�A�����"�%f ���ND��6|/ !1��~��� R��Ao�b: 5ժ��p �+�c�)���aDw 3��V���u'������,� [��_�/�h��ڸM����c� ^�Г�� _{T.N0;���k�#`���l��� �E8� �=
<0.# �����l_� K���ɿ�
�<���w�z�� �gРY�M3N	��E ���Gaw� �^%���h:_&�[ �~� g	k����ѿJ ��.tQ��/H�0 ��?���� �_0M� X+�h�R�1-x���07U }ߺruvM^?z���������>�02]�Qb�X	h���߁�	��=�����Q���L�6� 1�4aVX"��������p�� �^��?��`�v��-�QՔ��(pP�y�~��VM����]#˽H�" E��ȫ�� :�f��5V 9�2M��HC>� ����i��^���L���[��(��� �N޹�
�$8M��)�u^�O #�YS��-��Kt� p�"  �H�WY� !�d`�;$��x�@�ϸ��� ����|Y J�D�q� 9�.�+�5 ���`-2݆ �$��Q�@u������`I� :3�4 ���1'�P��`&� ¢].��{ ���&��D�@ m0�bz�Ct����8�� ��[�,��%RV��!��u|������� �`��gw^��k�I�a�# �uQ+G>� k��`���_��i��h �!���ɾ+���*��F��a )�Z��kL�z� ��w_�Ț��QN�� ����� 0)ڮ�5�&��'@U��� �%�o\� �X���w�CV ���:�>�"H����^w#��,��O �˝n�3��`O[� a���z�*�)F�2����	�۹.�g9���l/h�8{��z_\��P ���ȁ�X*� ��+�� X��8�K�py�z�qT�Q ~�X�\9w �	���H� s��0��32�\��w�!E ��`R�,�}$d�n �z�ɐ�a�J��$�0Z h1�t���# �'9!R� ��P�����Z���}� �|�@D��� _��V�° �ɓ��
� 9��H2K�Ѥ>*>@�c#�� m ���=�J �df� ��/�!�49�;���C Y����y-��T [��?w�� )Ӆ�Z���\h� ^Y��ϝ���@��-���(́I%��� 5�V�> ��G?u'�0�T1h� ��{��/fB0)d PѸ�5O�2+(@�ྟT��� P�-W�s;0�� ����y]Z� #��4q�� 	���|_�e½� �*�[��c ��1�%ͪ 5�.HU� 4뺄x�2 XRib�/� �3.;7V ��B醭@� _0^�욉[uI�p���φH�#3D"ȸy*� �T,"���7�{���� f84�S��[ +�~�ɕ� �]l�$�� Ȅy�c3� ٰ��� ��&!��W��@���^�$Ц�G�_ "�>��� ��-[�� 僅��0�f����A�P�ܯ* q�iĔ�v0�<����\�8W&!�v r���� ���Q��`��ϝB*��hg/��@���[�Y( �fh�D���� !Ӵ2�K|���;%��A �@h	��¶.�<�p��0�9���$^{������/� �Z�����_E�훀���� $��N�� ����n/t ^�Af����R@Jg�\���&�9E�� ΄  �C� ���AW��Hlf=`� 5�����d�O��`�v�� l `�	�_-ZϺ�%�Kw�� �5F I��^1�� �i��ۉ W s����B x5VY��1�^2�`��lh/��"��pwU ���%)��Z�* �	?�E��?�i�j���+z[%QR���#1��� �`P��x��� R��)�G[� :\�'v��O���Lo���"�P�Y�p(!}� �D��B��-}�Hf� ��W�h 7�r�gB��ۏ����� h��[Na� �Qk�S#I� �W��Y�� u!��n �B<��^]��� $��kC? Z�N���,0$[�@��`7��H
�% .!]L�5� b|��?���|���ϣ8)���A9p�� _�+���|�Pb�-������� ���\h�D� ��ǈ�~!'
�_V�Ӱ��
ι LUޞ�� 0����w��A�� �jÌ� ��b��J�~7P����YH�B� �1�:�5� 3� ��4 y^"׈�`i�u ��H��P� ���0��(3 ��T�V�� I����� Q[?�_�j�+ �KJx���YU�	�S�� �`� �W
 ѿ�K���X��uP�=��@G�J�� ���1\��!�j�AҺ+�� MJ0��S} ��.�Bo� g���\t'>yh��ʜ[�� �?��Sa� J;-N3�� ��ջ�h6	� ��J� ��<�~�9z�	�)DPp'����\�'6���3
�rY�@^U����F��� Z`�H�� P���ްə��$R@�w�
 �&�,̟� /Zn^�� ?s�(Q�[��"8���6Yh �#Z��yg.mȿ	�|�8z�G%�Ev9� I�����1ȷ��ʀ����}�����HX� :�d	�w *�Z[Y��Õ����W� ��!�
�F� �J�����=K�j����
� ��L�q�)怋v�j �ȡ��P�>}�_�� �W�r�������2 Կ�NB-� ����*��(Ƭ �!��� ~��B�U jDr�{���Vԁ�K_`H� /&��4I�~ ���}%!��t�§A��w� ��+Rb�W��0�� u����՘C3�f	��p�\�#�P��%��,wR� ×�"`2�Z�,��ӹ5 ���w�� ��ä��� 3���P� ��8J�?_� ~���U<(z�8M`��0��c� ���+_�- `�n�	i��T�a�_���,��I]	���~�@��&D��b���a�^̃@��S��V G����� �#¯��@ S4׷bT�0�hO!����I�	ո )�"�- �@�uK�� /	.�X� ��{��� �J۽.����^����	T p��ǜ-%=�E�yB��f���k� �n�	R��0N��\S�.����X!�{ 0���`A��� �P*�H�'�u���&h�Z �(ͯ5 ������ �=����`�  ��n�Fz� �*�[� �]�����0 �O���f�@t�+���3 �/z�[� t}~��l� �)k�^@� ��y�D J]�&�C���Z�>�-��З{b pI���ν�\ _�nD%�Q~� Yk��w�� �r8+� ��su! ̏�y� �P}"60X qs�2��k���ʷH�'0�)P ;L��D� h�o��u��J۠C +`뭗�����Q�h0��m���Ր�*�萚_�p�و Q�]Z��@4�2�=��:ч�%�� �f�. �蠤�0 �}�Z�+�݋z`kq��W�< �yd�T�@� H��K�9� �`��p� Nv. �o������% #S��:'[W`1���@� Y�4n�2�>� /��Q!
�B��yG 	HVh�L��4���Ɨ�.�~V���U ��#�� ��)qB�8p[�Ԁ�b�J ��:�>�?�=�!���
�'#��| &���� ��<���@�x������r%Zc����� BX��/S]����uH���[�C(��ї���0 �I��1 *�ѿmwW �g�)Z�`,pX�@�s2 �\YzHqH#� ܃8h�`X��Q� @��) ��} |����Hb8.?�' �i�( *)Y�0/ ��\ReU #�	��
 ��d�`�� �e�͛�- ����9hJ\ �4�t�" ��)�][�Z�*M&�PɦE��� ��Rh7G�b��UE����\ �����
$ �t	�0Uq����zZ�̢�_��	�쀙��1 yٱ�<� �!~L��k�S/��"0���gq%�G0	��)Q�+�'
��.��}r �$�F�ֶ���T�%�R�U�� �|	����< �A��� {�9x&[�O	�b�� B}@�� T�V���2���`�J� �ξ�����v���� ��Y��3����c�%�H?J`�d� ��#�� K<'��>b��:V� d6� S -g��	�������B*��% �{�p�� �^�	�E� �����!�=��FW���0؊X�WQ��E( �H^�	p�LY��. �n� H�h1�fG��4�#s��? SW��_>����u+��`" H�d^�E�[ �:%��� V�AHOw(P� �=�3��� ��_Y@� ��-�`W
=����@j�S���� ��YU%)�TBR�ڭ�\ Ҹ��� *0���J ̗�� ����I�&	{��� %q^kW#2coE�P�J��-O����k�� �7��Ծ�� �E��,	NI �H9������sZ� DY �|NR��ׁ �!��`MSV ê���R� a�,�Ҩ%� mvh��Q1� ��W�� ������u� Ɖ�T��� $��V�A�t>�#��b ػ�ni�8��
@~f\!��aӁ�*.x ���:F�� ��#_�O[ ���PHo��T�� 4�?�	�S*�>ź�W��=wJ<� ���>p��~T��[����&x�e����p�5 *���" %0�P��R�z� �b �}��<ܓ�)�Η`o�g(�:0Ϊ*��S1 ��wx�[X �5��})S1��΂ĕ~ ��^��$�?Er� u��}�,+\x��c��� 17����T�y� 	�݇^�$2Z� )�ַC� �N�?��c�� 1�j�y,'�� ���*\�IOrdK��5`� gˁ�j�2e ��,�x�$�C�%�F ����Eu�� XT7�]�� H�������ZdEh z��X� ��۵����?��Z��w�����	��zq��d ��g���1K �c�[�ؽ�~�.�쳏K;-�u �>c}�tH,K��w�`� ց)�QC�������l�~ F�1�T# @�ij�� �V)q���� �^u�,�� C��a��ǄJ��%��dW ��"�u �� �����w	��1��< )�Eʁ;�v<�&�=���z�c��/��@4]d� �3=��1 f��\uh r��NA���vz���/��q�0w�A�	,1n,W����h� j��� 8�QH>��- ��uL� " ���_�Rɾ��.������ ϋ0����� h/B��H� �d�FT±��f Y$��� i��b�J� �Hxf��� ^F��|q�X�����-߇W0 >1�X!�_xw����h�R �������j0nY�`�s��=��¿��d��j9�h_O;�Şq�Ț����Ј����5�# �	a���s ���!�:� µY��� f�$���� a����P��ŉ���qn���ç��� V,���2x �@n	�����7�`T \W(��*|��A� ~�k8�
� �'��-R9� ��P�%��Q�� ��'s0C��"`�YHj�5�]�9,X0w �������Z'��`(�3�� Y- �۟ MpXh�`E [�*��Fw ِZ-3���Դ�A�� �(�P+��<[�����U#����	�@ su �eY��X@�n1p�t<�O�"���,�v�P~�� <�������h�K0�/.�pk �gL�� Ů�\� �� �ZJ;	�q|4܀�1��[ù��������R(	���?��C! Wڈ<�ۤ ���G�q ���g�	� ���O��[|�J�ǂ���� ��)�~؃ Lq���2 ��c-�SU� �N�%���:fp ��*&eX	P g�3軪 AhBY�q��� �ļ��ܮ '��>Vn_�9`� ����� �[��=�H��l3�Y�t� ���AM ��d������p��� 	�Ts R���<$�� 7 ��d�2 �׵<PCS ���R�* �w�02���' ڢi�P K *��� �H«���|%v�	�^^U�Q i�D��� �Ѱ]�� QY*0�s �[��yczd D0ǩf�i(�� ��w��"�OI�	� � ֈל���zA *��\MȺ$2$�<�)��+ F�0'�xh ����߬� ,B�w~NQ ��[�-x�E���� ��8�t) j���u���LN	��Z�!�#�[ƅ��u� 5�%��I?	Q~O�.`�F�1� �Z�ˀ�K�0Q��%��d��w�釄�a�4ph�������� �_�ݠE�T�K���J����[c`��ޭ^��!�Y��9в�h�}
�W9"� +A�ӵ� �8��WO� <�Gwlp�X铔 ��fm3 �'2�Udn�BN����8��@9k0���"� �}%z��*Hb�͢J� ���¸ř�#P]��������-�� ,R�U�Z��"��Ҩ�zg�٣ e� �	�d�+%� \|NiT��� �
���*� X���.��d\'�{�`	�~mra]�Ҹw�p���+6�ÿ� ��{n��W Kt2(�kZ��!ݔ�b���_���&;�Ĥ�D�����/P����޿`Q�UZ�L� ���ҏ���($�W��9�������_ ���v*�1� Q�f.H�� ђ_�?� �Y"K�����P )�U3�{0^\� ��	�:� &nI�/#�u ��į@�{~; Y_(�f k�ܺ���+ .�S��! �YV�`�f� ����D�� ��L�,ӂ��Z��7A'Y�0�? ����x��3' U��n2$���!�0�б�� ����^V� �p�r�ޕ �B�0[)�	��ὀnh?Ecy>�N�O�@��X Y\L+��{t������ $a�G.� �p�-�� bi
?U���8���j����� &���� ���!��R��)�%�+� ��ڕ�$�K����[�� �:p}�zq ��W���� @l�k�"^��	G4N|@�&�I�X`$��t�	�j�(����h'd�w�%Y ��ݟ���� 2#ƪ3/
� �hUְ}'� %�)ݻMD Jʷa1_�Uu�.p�,� �* Ƌ W^�o���
�a0���d�K�( �Å@	��� F�'Aq� �H�(�V�%&`��14q�u(a� jt��k�� N&�r'B� D��+�~} A��C!����]w�~t	�im� �<յ��R�2 D�/��:�;���8����M2�<�L��c�W@��* 7��(�� .��S�@3+�[ X����� Z����� �됶]+� �	@#���5����9Y�|L �_�C.���x���� �#��u� X�+���Z�2�w V��H�; 'P���Y� A�Z0h���`�黰���|� ٶ�EX�:�.2����|�0vu\	PQ�K`�6W�z�аM���Ȧ���[ 0�Gհ�W��T���`�� ��$����>�)��_��<ĽIH�j ���wY�5 J^���6��<	Ń� (�~���d@��U�
�����Q�C� d�#֑�>:M?��� � 	�V0��Q; ���F�� ����=uVZ*� �h)#>{ 󖟠�2�1���T/�uD 3��#���1��@��<X����V������C2���� 4[���\ �ːꓻ�<LP���S�l���e�>�w02�0J�@� �oZ�I�� Y3��X�ѽ�쀜� ��!�2|� �h����^ 3X�b���	 �R��a�_� �*��%b4} �$�9e��(�O� *:������� ��;kڒ  �"!�_�bv� ���F.�0� ��Hf��(	"�U{@���?_T��%[�Ig ������y� !�
�	� v�Ixܴ:S {&��[w . ����(Ȳ4����N� �_�������Y��G VW �^�RO�Z.���/�� �ɺ�We�� �=`�� �� ����~n���������s ��L���_�t�<i���z-`éE��9 M���@� �v���� ��> �NOP<!x�"� ��<C>�<jՉ� �w>��Ѳ��o���JH�� q5B�\�u ,	%�A#] n$�!� ��ڊ��'S ���|����ȕ��b�;��V������Z 1�s?f��P�'��������(x�� ���g��h �_����V<MU/0���o�b^	�� 0	���{X��ʻ�(8�jb d��B�]�� ��2�_ ݀=ʤ^�{�RCx|K �s"�r &��Z^��L�WT �>�"�&���%��U�  ����@L� �&*�2-��LP8	�Z� ˄:%��=G$ �
�&=���T<c�p�  Q��/g�� ��1��"�k���R��uM���3p��LY h:�m��-��*Fu� �@Gh�X�A�3���f^��I��Y*BK�:����"@髮( ��Hh� ���y�% ��\����� �(�?��7MҼU��ȩ �!�Y09^ �X+؞� ,�^ח̱`c���>�# ��0 h����J ����M	\sP�%@����T��Mw�cA��
�S� �Q�J`y����}	���)�a �Gi$�b�<�͉����l��h����W[[�� ����Mv_ܤ� 
]�� lD�`�	3��t�
Q��� _,���X��Y T�P���x�zX�� #	�h�pu 4�$5��˘��,�`�AU�$p�� ��)���s� �*
���%r= p@�)�U ��
�ڣ�}� B\�m��5X�������:����_3,�] �l*�\+9�W��ZD��	b� ��V��py� <�Ӽ�?֖$�PN�Z�`��X�����\^ 4�G��� �pX �Q_�@��g�( �
�X ��w�� P��1�9�^	񷪐��h BS�2,��=����'}�҂� �d�|_H��yQ ���7ZRUv)� ��hV ��]f��� ��Z���_�� �b'�;MO� �S0� ��f?$N�� ���!:�ӥ;�� i�L�}� �-���(E�>�� AQ�[� �V�� 6�+�@-7 HF?����8*�cS궀�h� ���ଡ�� ����" ���x�6$�;��,�e	 �����c��@�hpj�� WS���V *ɾB�| q'��?$V DWݿv� ���p��� '��~a�?�� ��>����S�Ĉ�P�QJ������/��Wz�1��A�% -X~8��DP?��	%ˀ��Y$P��`�0�� H�ʓ� 黋����0/��9L��	0�2�T�рOU�� w�ׇ�+�F�^W�����5�6 A���Q��N@���D�� BX��� ʺ����h H�@��c pb��r�9� ��\Zj�$R0�$��,6 �I���&x�Jj���`.Ëz� d0�J3��2B�]Y��x7.�KD�*��� ���fh����?��՜�%�PRl�*X�/
�� F�@K!��I_(� }-��s� �/C�>O "�9�K��Q�ȷ��v��Z��e���{%��|� �[����̮�� ��N����'V���%(e��L鍘�Ow�� ��Z���� ����,��� �J8�v[�)]��ԠKŭ,��hC�2�� <�N���� %��C�H+O����ZB��aT� ��� �ڵ�>�,� �uPƚ�� �9����j����B���� s �x�afٷ�VHϸ��$]����) O
J�a� �.��c�����%���~N�� �j ٙ�- �@��z�%�RE
 �C����� <�n�pU�w GC1O�� ���)�]N$ �/ڄ^V�}A��h�*	m��P�0&1 ��\ z�Q!�,�=�ӃN�a���)� �Ʉ�H��6 ��
�� �I)��e 1��	�H�� �|xl\Q TY!'av� `��ַ�_< ŉY���PS
�����X� [��տKH(ѓ��`�o��2+%v�T G���!X`� 7�~�A���N� ���i�z�H���`R�\���� 5�����v�	m�Z�砏�;���[�� �^�)jq	�~K�w���2 ������� �X�h�1�:v\ ,|�a�}V� �-^��P ��Zbװ���ޯ�yC�n�� e��D��YrR )�>ɻ�.x ���EQ��~� �U!��>; K0޵\S ��Cr*�� ��%�H�����3`�! ����X	�¸؀*��&:0ބ�(j�L��
 \��	�Jf �6C��t�,.�W"(y dU�#V ��,v����<YȠ� KX�a%�.��԰�����sy�`�]Bā��H�� 2�ȿ��� ����[%�� ��	���N�x� `��_��'�:I�} ;��� /Y0�w�`������K��] ��>����U��S��M�����f�� bXY~���|�&w (M%0[H��:���p�u�4� ��xc70 #�R�5 �N�2^�ZW@%U�3ҽ 0B +P�� �$t2q��1�ӯ t��VT �LJ�`q���'��v��ȉ j#;�SY
 ф�(��} b��G�@��~��� ��E$"��)�hP�k��]mE�u��� �U^��l�
�h����.p"� u	�wsQ�q _�S,�O�џ X�d@��%3(1�������B0��I^��&
� ,WS��� [���+b� `!j���� u�U��tk��bW�7 m&�U��a 3%�A�h˱>b\ ��]֎� y������hu@6p^��yu��8f�Z�����W��m�%Ґ~�N�q1�j�s���L( �ޱ�	�$�nw ]�,P�~_�$U ��\� ��
����B½D�fi,��o����r0 UƝ����9��s5�W� �����i�ٲ� ����h�LE S��a ��L>	��R �3Ȑ@9��L�Ut;���:��"1?+�sB�t�&�;���Uh�G� ��>�u\J `����|������W$wJ�Oї������}�[�貫%��`�� �.г"� ��K6(_d 1�}��� ��G��c��| �@p�.⣖ �"�Z�� U��;��3�ǌ.�`nR��\�=��� ������.#� �SX�} ���1��Q���;�Kp�`��Xd�O �gߋT�Y����\e7> ���]��[�� ��x-�SR �_�o@�� �C;�^�A� *�e��<+� ���o h���"�U B�`���<�� N5_�]?��ަ��2y�v[t� -)�+�X���X� ��'U���-���k�> w���
[�`B� h`,�2�o�����������0��� ��G�|�P�@5 `)���J�kh ��׉< ��&�1� �C���Z�<pq��� #�G1��EK %>[W�|y;�x���0�R�Z���+ �r�璁�_�)@����1= z��[yi]fp@ Y����$ ��'�,&� ���	_h+P Y�/|�%�O�Q)����>4 j�x}/�dt7%l��`�bN�  g鷬�@� �h�a���B����	�2Ni��P�8%���� ���)�� y;�a�qp� ��V�t\	� �� �H,� ��-��.fX{��즨� G`��0�f �����������;1�Y�Ľ���$T ud����'
N�сp�{ ���t���8们#������ ��j� �I!�Ë �o�hvt�MH�ĺ y1�e�* I<��`.(S=�� nW%	�_�� ���S��m[��@�!���� 3̀p�2 �_-����� � EVU2�K 1�Pt��0 ��`h��� �[�"���n�,�LE. ��S#�3` 2�K�����.�2>����3��\0] �h�ѷ� ��.!�wG ��N�nLf�`u�F0�B�����$� i�k=��\&7t�@d���� �K��0��� �oU<V#�.1�� 5���F� $��58ݰ���w@��� ���^�k�=K�?����h��� j��ƀ&+� ړ��'QG ��z	 h�� �O��6� 3/���Q~� !��ͻ0� NȀ"�W�� �����j@� #����m�QP<�`]CX -�g�1^�����>p �%�q�� �0L�'�a� 5�u�+/���M� ��'��j �`���ŉ mri�b� ΋7XVQ ,!�~�Lt/$�^,� �W���%:^����f����< |1����	y��E ]G*� ���R�ڙ �eT�O6�`y�nZ �鰒�_ ��%8DϽ �Ak�Q ����鞗z�Y�/�2P�K_F ������&�ʹW��`Z�(�	X� b.�، ���?�V��_
�: ^�\���v ��:��2�
C^?�h���0������_:�]�R� cVo���e ǉ	�Ql�! %g��H�9 `T�5��(� 4�F�Ÿ� �/ �R�'� ������(Z�����Yԣ �S
�����ַE �VԶ _�#�:���@�9.f)	������'P �3^��0��Фt �>�	�,�7k� (G*� {4-
F�� )w�����!�[S/�6v�X�v t�_���%�8l���`DU�m�� �yB�gP � �@ax��t�З� G9dL̰�0 �_#�Y-	�ִ\X��%��H�� &�=�Z:���x`�%� W��X[h�� vҚ��ѓ;o���r��K��WH#�E�r 1Z����6O"�����d� �(�q\� ]�~�J�e�������X% p�"�D!b��l��3oP�E	 +��?�0�4 �`�D 92 �ڼs/Xē u�'K|yPD�� �5	ޚ����_}�J�U��������� E���,4 "�3�R���\v� ���
�� ;C�T !�Y{�� v��V������'ă� ��`�^��]R������ ���/C� �	��z�˕>l7Y(2���� p[%��V d�J^RL�ꈽ������y� ��_��(�	 V���N*Ku� ��'�p�,z3 R��D�� ?���I�[.�� ��!�Xf� �+�҆^w�ST��h�_ �txi��ul �TvZȪ� ��� N�X�`�Y�Koz�  5k)�W�0�3�1���w�O�/I\)S���� �ۺd���%���i�_�;\�ZO� �y Ƹ@���&�ϒ-�� a�`�\Z dN_�N��b�p����k!PhCL%��}� �;A{�V� ���D%x�����Lʹ�l!y��Q r���(|��%��2�T�h��W0�:�!� �`�'�"~�P W*�Z��< �w#7�V�[�U��>���9���]h�<yb ����a�1�`��8��^�I��k�R~@�,]!m8y$��"�\����  ���߁��ݡ���;� �ޙ=��- (L��_��	 �t��h�� ��@��JQ0���e-�L�"� �R)��_������~[�ֈ�
K W��%��:���\�_�°�,�h �@LK��(��!Z|���� �涕
0� ��\hw�� ��~c�o����рǫT��"�����:����2� μ0"�PY鍖�����UcD� ��B��L8x�R �	K�%�� m��4
�ِ �^(�څZ8�" ��R��! U/���T�� _+�u�'� �,n��� ��rغ�	&�j�% zb��(�Z� ����� e�^�)};`x}�.H�%$f  j�-�@�LS�,�D땀�t>B +��efj�� '�(�饖 x�Bb�1 L{��ʽ ���,��.�e�	��q��B���X��� �:�.aҝ��I�[�Ą�N����C �U �}F��5��HtŹ'� �w�BI���G V�$�P"h-t3��SWX	 �_c�A��@�qQe �×5��+ >)-Xܒj��������p�Q�o� ��$�#bX�a���÷Q+  ��8p�f�L ��\�wV ��R�2}�@ 8^�H����{)`fh]�-�9`�cRF` &Vh4_�<���`l���z�>E� �T�fN,�9� )ˇL
� �(�TQ� =�u:�G ��-�dX� �ĝ��F� 6
����� ��(svH2� �Tm�5 @��Ծ�V,[Q' &��t���ׂ�z�! +Ͻ,ɉ� ��M����S> ���Z�Eѹ =��*��� P7��?6	-Jz��N`���_���������t1P )�K\�=��� ���� �!����["�� 4��]q� �+-~3�(  ?�J����F� ������ ��v@�3$��[�J�V �"�*��Ž 8���K��1^06���u�)d�n�����Lh� ���9K ��W���v�S�@�áf't	\Vz�`�� �]1�-��qݿF6O�M���3���D 	 �5�c� ؆�l�f�&���8� ɰ�(?���Q$1퐅�� T�B�zg% �@ V���d��w�^�� �XV�� ���Y3zE����(H̓@��8L A1J0V�% ��ph�)�;���[س!���f �"��1 
�ZXx{���#,R	P��`@\�w�ݏ�]��n����Vv�E�,T� ~1�- �[)�h��\3b?�D �'P@� �B�>3�udN��@�f2ͲR���dރ�3���a��J��i)ذ�XY'�]�9��V��> (��*k�>�aj�������NF��%8�T�cLX q-����`
 ��v�V�  ����/ hwb��~� �����D+�w�jčP �^9�)�� B;2௵Pc�ɞ`v�NC�x��
ЋZ9 ���P�N x� �X�.����3�������b��Y �h�Qj�	 �J[S3� ��1�H0#ʐmL�5�����pߗ�����c����� �u�h�!��l?�.�B�"�� ����g�
R ǯ��2�;�r �}�h&0`�x��9pЦ>��&�Ƹ�?���(� ��M~��'�@%hkYO�����:������}J��^7 @�Z�$��� ��9[� �;f�$�u{  �!��]���G$��P=bk\"���:hp�؏����i ۊ]v���É�0��� �Zo�P��e^l�����H 0+�cO�����f�$��- [�	�~/x��u�� ^�9���X 3���N���P ��������^�;���gE����:��I��e����� �6�0�2A �EI��K����)t����Wz�����S̨ ��͛a�8���S1�<�������ڵ�� �aވ��><����]?���u`[� ��A��pf�y-�/=E�4J�m � k(�Q�{�v�>����߃_���;�P���� !� �_��L�k �k�]= V�?��,� 3�����O& �t���਑ ��aŏ� �w�PQ����� ��L�y �X��D=-� ��n�d� %�Xݥ�ɽ �����.�� t�Y�	� E|��(,���_?���2n ����kT� *!�h�AR ̝�\�-݃ �2��!�W �cO��	/��>��Z��w8 c���T �G�$O�� �X�]Q�P1���J���У( Bp���-h  cf���$�& �DK� �	��:�J �j�o!�� �H���z��=B@D$�Om2�̍_��6��PG�} ���Tִ� ��6�\* ��M�F����IQXP�'� ���GZR�= �	��Uс�_N����LpG�P�-,��A߉�}`�]q '�����v ��j����f R�h�)��^ C�B��_ﰁ$�vI�A#����D:eT����`��]d [���K�� �GA���t0 ���(:�K� �A=�[� ^���;��p�c�O� ��i� Z������U ��(�c\!i1�$�XG�� ��~�,3</ ���	ջq� Nr_�P 0�k��`� @�h8�5[���0��ױ��sN Ю���vf 1�e��L���|ܪ\��x%��)�0�^� �Ӻ���}�:	��|�b �*�L)� �Y;��0pX ��ە�A( �Ď"N� �p�@k�x�%δ ? �������j���ɸ P����(� ��0a܌Rw� ��ω�Z�� wD[�
@ m#b��' J3�k^��U�;e嶀��&���7 h�#��:i� !��a�%�Où�#���I-r ���c[� �K��q�� �*��aQ�� �
�A�f6ۉ����-0r��v� ^�u�|;i�>Ӏ���� �-B2���@?���� j�`ڕ ����R��V��[`���h�ȣ��$��� �H%�VR ��"	����K�PGX��*���3�j��� �HwN�u�V� 0kX� �)��3�Q �A~TY	0� %��_8�| c�&���>� �yB��V 0���?;� �ۀ���c�j!� ՙ�*�. �H��RPV�� ��l]��� ���v� 6 �V��o�ՠ�� ��	2χ�4���s� e �f��-� �q�")<�=��Á$� J1[r��(Ui�sDȠ��&�> �(ى=��3 @��}�e\ ���Z2�5������[��� �P����� 	������ќx� hp��ŔB�`�3����� ���!�K� �h�,� @��p����@y�`	Uf ������1N �I ��� J�Hq�b2� �z���uX���{鲬� Ż[���	�ځ][�,ԨG& D��� �d��%	�� ��}\�2 z����o� ���%n0� �T[2��� I|�&�/� ���
�l�Y �|�5 ���ݓ� ����տ����+��*e�O�K ���E& >0ߴ��Z(��ȟƻ/��b�X;�_���n����V
�;�{��l)=*Pw �,�#��t�ڬ21�0�a @��l�I� �����U�� �^Rw��uS �P��\�_ !�������~ �G L) S�'O�"� �q���%4 p=��(롐@� �1�ԕ�� ֑>�uS �X���Y�/8P��� �|�� ���)��0 �N�1h^DTA:�$��܁; ���b'�� Wo��H(w� �����4��_�p��j2
�饌�R��� ضVp�zZ��"+A[k���q ���RI� %uE��3V��^������j��� S#9x��< )�Z �h�i����������:�}�'�b�0���@��$��?=�/`c0�h,L� n��p� ���K˵�>���8��}^h��� 4���&\A\X� 	�>�gāR���`�P�Z� �A��ؠC �3�	���lKu�k�.�S��Xz� ų�/s_� �^;�������@��N\�� %��F�7s M	i^�IO�jJ���EF�� �RV�����e� ��yfu���H��Ba� �9��L �
�͝ZlS���Ua�^`u� D1���E�,��	4Ox ��|i�J�1��8ݡ3��y&Lh'Z��P�H� l҄�\2����`B� ��X�q� �S� �' ���e�*@O ���RY��w  +��/ �q[@�R��H|9�=��zwt ��R�2h+�x�%D��bGg-z�=������� `)Ջ�1�M >Z%���� ����5t�B�`޻����G�،O@]����� T����` ��P���R$aR� ��b0[ L��h�# �_�W/M�:1(�����{�[��J"�-*�@T�ʀţl��~ �~Z������ k�)�=H
����>���8 ������u y�bm��0@U�����(� ���x9»{e{z ������ ����[�*�h�U���	F�.Ǫ�Xh�5�U{Ā���d�&����'T�� #�ѩ0�9l��H~���`X\��� _(���b+��	�uz�� ��yq�h{ &���D�� ��sܝ8[Y]��x2��X6>� ����� �	Ph4±ux/ S@Z��i� dh����a$) ���W\��~ .��b˛U� ����xd)z�P�D�"G_꽠
�@� �'`X�щ\z�˺�C�J� b�3'���?Wı�P �p�� �_�'vr� 	 ͑�� G�䓡�n	r�d�u�%�ȅ� m�*��BJHY�;���QSt���8�N �2�1�]
,�@��J-��h\FM �D�����K�󾁐��<�"pTc?Rv h�]:� ��լ����� �d����,;� ��'_Uxz�sz������w,
Կ Xk�;!� ���$��K&����1�� `�\S�) V��%�nL� Q/7�YA����>�
W��	ɔ0au �h���3�KX��\�T_�z5P��� ��� #� ��� ��Kv��I ������ U�Ն�d# O˼wz4��X�B�h�QDZ'��f �(%/ܹ*E �������Ș� &���8g�'Y�]�P|�F�<s��cj4\_�0pt��=}� ޫ�w��i�
��Y�l��@p%�v� �2	�,�Z |�P���+�,3�� )K���ץQ ��B/��0I�t�G�u ���Z|6iv�@=J��h7;
d��4 kKDwajl �/r��N� v+邕9���R L8-SR|�� Z��I� w�Yh�D ͫ��O. ����?������ ���H-� ���5��TX) L�}�A �>E��;�j�t�VpKT �m�>�ϒ�>l� ^��	��_Dh�=`�>c� ���81)u�Py} v[�(3�'�O� ���r�~ U-/fb��S�� �n���]� %d*�ā����-3Ѳ�@�sj �`��� 'Ki��� !���_  D�0�-[p �F� �\X�`�ri ��y�ʈ� ������ ��.� ��X�^t�0pS� ��[r����b���z'��i<��`8��H� N����?']��?pw����D�U���'�V�;X�x��6�$���"5���� e�n�H�: (���K?�,�*� !� �������s WU�ŵ`� ��0[���<�@  �!M��wP��< ��,1�SQֹt^裔�@ÈPK��	�hl!1��?�p|�������$ `���߽O{8�K��呩����/_�Z, $,j�8 VΉ�!J ���k	� ��ÿ́h�-�c��1� b^yaf)�o �O!Ƚ���M�k��yW�S�em _㡃l��	 ���}�i�� �U�K�u��
��y�� �_�� �L��o��� ��)0J��q��O� �qHa+�R ��]��t��@굤й�� &��C	AS� V��8�"��h�#K�0T���f�A	�0Т�� ykc��h9 ����� �B��`��[ ܟ�Z�0��WMB� /��[� ���y�� �|	�݆h\ �X([��� �0C5� aLU��y �:���$�S�[? �Z_��.�� �/*V:@!�MX�6��^���1��Sh]��_st@�����ڴ&��'R( J���q�՝�7 kZ�hrJs �M��9 
*��e �-��V[ٗ��_��-���z
�Ď� ��o��H2�� ����(�) �
�_�� %�H����~��
&K h% !VZB_� ����v�(΀��3{_y�*��� ��ꦆx�(�!���o��?��	�ԀB����<@5������ �#A3��X 5�1�(� ��K� ����0�� �R	
C���8 ��@N����_S�`������b��`.���pG.��s9 �@�D*-,d����/��Б% Z�v���� m�R�b3�X;"Ѐ:�D����=�.�9����@[�/�)�@�"�N �ɒ��x#����}!ʀ �9Y}'5�� r�Wb� ���G<
α ��)�g�N��t�_�G\���A�o����y(��^Y ]0 XV�u�꧈���:�0��~� ��ƶ�6�K ����.S� �U���	�<�G��3�K C*�;Z�z� @b(_ŬP ���;�N�� �X��!p
� Q�D ��.�	IY�폠���v:Խ$8؅����s+`G� <"ܼ[4A�R���Z�$#���@��h�^B0�:��I ����Ax ?���*� %"&ݠ�� ���\Ԏ�d��0h�N��=� ��g�t���R��q� �#�{��XG ����
whw` s���\&E� �}���A`� ���U9̕��wΘ��� ��
��' y����E ?85���!� r@k�� �	+�X�h�`��2{%YR���'�$k ���+uU� ���}��1�������w5$I���H\
 ��!�)ы�X�` Ig�u&4 Qұ�?� �w���N��ƺ��{�` �����C'���& d]SV��� 8����^ X�K���\��`�Zz� ��3w��� �������2	Y ˹�� h�� Z�kh�i	� O�]L��!���ST@��O �i�C<J	 �!Q��pm ��V�.Ke���O^��*L��x] 8�_q1�
�:���&��m� \��Ӳ�ZW�	����/� �ztr�x� .�Y<���c�;5%�0�����B2���_�%��)|՝��\���˺P��V��p��Z����h�@ �� �K���� J(���{ �����>
 ���0�Xfp* ���Z�� ����q�n��epH4 
�J�����bT��2<.9�1 y�3�-0 _��/�P� 	(�%�)TU ��>�k�� ������} ��z�O��(Ⱥ����x\(� "�	�~hR��&y�2��B��`6������ K���&Pc��4����{�3  U�n�� ��[Zcl�F �	��D������!�u���\}	 ˚���J؁L 3�10� ��_2������� �@�.C"����=���� pcJ���� �y�K��� ��B�u�w� �0�#9���2�߄6^ ��z@L���kAԇ�U��� (쮴�n��e� ȟ��� L�jW`g�^}{ ��IK�N����q��X���� ���"��0�� 9�<�VHA�}c\ fh�B�:�G�t���(� ��a��~1�2����(}.��4 /�8�ec?�H�]N�9�?y�׈�����8M�S| ��`���";�:�#��p�l�� ����W��X L���]0� ��z��4�%W	Ԭ&� ٘�\�I�T[z�6@<�,2� X)�Zf S(0���v���� ��K�<X� �H���q&2����� ���+E�� ��{��WV< 	�&�O�:R^ �0��(̐}������Un����0��Hß�J���`���;�*�>?pX i:o�/ٖ b��c(*Q� ��ȕ��1�)�0"����Q� ?�+ѕ�иTe�ʐ��� 9 �Н��<ׁ�h�K���q�0�ƴ/��@�W(J��2`�h1�?M���%��qY��} Ef/�3�:Lz�9)�_�'�`���������S9v���!�^�� �OB��F��v �_Rhǘ@	յ���c�/�&��� �P�%�_d9"�?'��2�j��tV{��(�J��B�a���o��X�ʇ��E �f[ �h��-<ʲd@�FZ �Ƿ���}X [���q� IF����2 3Z]�W j _����	 �X#�Ғ!� ߆��T��}�0|� 	\��ؘ��|��ԅ 2g�w��p�|%C�@̀�z- k"�w� �:1=�dx�} K�!���H 9��'�?{ ���VD���/ ��SZ��1�o$��B �X�ئ j4'U@�]n �Z��b��9�f�_�뫸P� ��o�G�H�/ _5y��p�2�h%~������L �Z�,�H����Ȃz���[�.̀o����� JV@�'
 K�����h�� ��H1��� $�:����Z�@߀�Q�� /��jҸ� ¯�z�-�. a��oB���=2���!@�{� z\ɰ�� ��[ĸb� qK��/�<� �1)zɧ\wM �Ħ!� �G��S� ��ː�^q}u 3� ���� %����j �x]�8�=��O@���[���Dm���(�P� ���K�N� I)���G�	��0�ٯC 3��o/�" �wE� � 6!_Ii��w�a b%�Qr}r������^���1�_��[����.�*�� :����3 �2�[~FW�a�+��� J���T ~��?�E0�� ��Y�'_ �� ��Ӯ ������]��0��(�de� R\18P| U�Ƈ���6�� #\4�ժF�����+� U��h�4�� ҉�@��~� '%#�ݔ[ -�6k�� {b�� ��\�_s�����~&�UD �T��x�� ܅O���A�X{���#w. u麚Å ��F��_b�z� 	�]��Z� ���Bv�,� 9\�Y�'� ���B�� ��S�֌�I�`Q0[& ��`
�t.��P�.h(ՀpV��X��`��@��{��V�߾|M1��_4 �����k �N>�湢E?h�]��W��{i��'���3�>�`8� 	��P� �R-3�Y���p�� �s�� XhiC?!:�y0Eɟ���t_M��غ�e�|U��A �F�f�Z�?����)�z�� ��y� '�Z�!gʵyd��X�!%y�8�� �ݾ��������P� �-R��>��4q{����� Ѻ����W��kװT� X�� ��f�Q*�Z �N������n:�Ҋ��1��yĞY�2� ����� RX��P� d���m� _�XW�� KDa�U�@�T`Y��� b�l+�J��;-�����k�W90�5���' R�1&� �4�-�Ȅ��� ���	_�(xt��� Q��̌P3� �ܵX�<#ӧ,20��!�f�y� G�� %��JU9�1{S*������ 2��;��� �=Ӻ^3�(��c�����YL :%�Fw��$�b $V6q	�q��Zu���h�L ֕a��i*e>���b`��� l�'9�]�p �h87XN�� �z�y@�>� ^��)��
��E`!-@.]==��L���}�$�<* ��YX� �V�2��Q��  [���"�<� Z�3 %� N����a �HT� F	hQ^��!�@��1�S0� ����� ��"�\P� ����j#�� �]��I�� ����s {��Y�!f� ę��p� �V�"�	(���0 ���
Q�~z �l򞊉�t�FZ��h������q��n�# δo���X� 8)�J��[� ��D�E�� N�1��Fv�&*�|K�L)�|�o>a�i��Ȩ�q� ��Zv N ����������@�0���T����������`�t: �fL�'kv�	%��#C 2���u�J�RWxr�K��  *�p
UZ� �Wys�j���'/�}�=��D� ��lS�e ��bP
R#� %�\�+���I3�{�� �P�pe��X'�|VJ >�J6�K�"� !و�%;[E d�ߚ�� ���B��Ob�[/�a�n�0�� k`��'�Y"-�Q����_`}�0Z!D ����� ��������j��_��`4��� �����3ru �~ˈ깧 4��&�k�I�W��M	@�xP ��5��� �s����� o�¹�m l 	�\�]N��҈ ��r[~����8 �'��� ��U?��� [uL�v�\ �B��S5�8U����1���᭝�`�7�8T\�Pz��0�VS�u��y\2Az������ t�@(	
� �mk�/\j ����4[� � �J�΄����Ԑ �oL��C |E�R韤J�4 ��¯��b�$0���A�� � ^h-H����8� Z��� �.^��)�-�=����� Yr20���D �R�Xoutzg[�0�_��]U Hϳ�ɍ�&��|!p� �'�H��a�t� @~1
�R� �^[)�/�� k\����h �*З�İ�P=�S �to�� �LwN�=�� W��O� �V}�y�d]: ��\�`(����!� ���^����)<�;�T�{I �0#>̥ �^2���!��� /�ZRq53�-F\FٻA��4��K���z`u ��1�� ��-�`Y 0��������4P��� �-wyahnx*̀.%�� ��ɋ�����>�� 㰘R� �?�ՠ�rt��	�NЀ��� ��C��
E �#f��&Ũ	�U�{�x�v �-�C�c��|��1���m0��H_�@Ȼ�n ȦE���� �I�M���	 >�dj��P] V�����2���d��`��Ƌ<�E���b,t�!'���	�>��8��y����*�R|���@��� �~�R߀� S������P���� (x����%�|Vu�������o��Q�;LŇ���X/3w g���x�=R 	��k'2�� Z��A���P���lHN�� ЊX�4���1@�aN�� ^"��@� ���	$�b��F~����uN ����@a�����(� � �؜8�x�<���k/�0���hpl�0��w`A�H�p���6�L� s`� ��5� N����+^���*�kM`"�Y )	����L'µ�D���Ԓ )�!յyY|������m��ʢ�X�=���Q� ��: �-��^N��Hر!�޹����F�, o�����F" ��~ �V�lX�^'��a ���},��-�J���_ԭ ���,[���A��t�%��ڲ�K >-��8P�a �:^��o����#���� 0J����Z��a��`�S���Go�U����Ak� z��� ?;0_��q �C���b{�-;�w��~�xC� !��%�/�{ �X��Dj 8�|&�v/� 9ZF��! ������%)W#�st��Z �Y��-��L	 �X�nq ݹ
 � x�1e� q��+�	P�R� �^)�� ���X�O���h8�d�a�����x����� �%���͉�Q���	Y��P�� �n7÷�� �5_}Dy� ˒w]kV����I�A�Հd�8Z ۀo*�J�� (�1�KL�������Bh�2 ��3��K��Ǧ9<�*G�Z ��8��&�� �䵄BՌ:�:�;�|�_n3�� ��h�a� �,/�l�� ˲s�N� �Ȅ�E�n5���c�x��O?${�h�j�-��� ��T ��5���a��}  �]�� �S����� uتx^O 0Ԏw��%���b �������1I����d����?�� �_RT��:�������p/	� R�$hЄ��Qz� :�k���" M��2��.� �]�8��;+X�[ �����! �3�y/\, ��}Y�%��	} 0&�'����>L�\�� ����Y���
 ��Z��&M��P�0>OR� !%\߲��)^��K��*��~ah r���>��O �x	vpq�`�+�m��tJ��X���TH�P0�S� �7�U(n`1 �3+�I� 0�Q��~m	 �O_y��vC�,j���� 1 H_!��X �[�� 
�7�f�\% 3���4��,�� ��ⲷ) R��C���,P����\h15Р1�Q�}s���>c� �	��[�" |��@{���8�� R�0�Z�L�X ���_��Bv!z� 1�XZ'��A n�6�K�(��@��d� X���V�e	���ߥ;�1�U��z�H/���� �ݒ�B� mk��T-������ �f'�`�j�*� b��%+�_�K� �Y��\�8� �!��e *d]���?��75����� 	�'_"�a� wE�$��F^�u`���w� ��0h�f�O v���в.� ���	ѿ�P �����pm1߸<� �[�A� ��9Ā0������������ ���1�0Vo@+�_�%��v��1�#0�p�|���ۖ�^����}��`�<��� ��,@S�'l ���ˡ�ښ -	�0nً^\. Y�G�� �dA]@o]�ǘ#��8 ���ʗn>�z W�q��	��*Z��!�4/� ��0�K�Lf� Lh�1� Z��ҭ���T�� �;73Ye������.� <�W�5�L� ����>\�.�V)�t�����X����' u��>l� $���ņq ������pM�jJ ��. ����r� �Ӂ�R�j�~�fn (��0 �[2K�� { ��r�&3 �P�	ݖ�r� �K�<H�� A#��=� ��Ș�&�� T[d����2��.Z�0:��F�_�е^��!�����x�T��ur�l@.�~ y]qZC 4�	G ����{� "�P�;j�b �2���W�s� ?��!�1��2��zD��B��� �p?V�E N�j� %�������/�(z]���+@�,�h� A�ob����m�v Y	��� UX�'h,~
#��ږ ȹmH9�����՗�k� Q#����%!e�b�^�`N� y�A��xT( %��/ �� i_�M�D�� J7�X��� �pWĿ�x��Ze�+�	*�w����f:Q���0 ���4�P}C�$�� ��� u9�Ճ*�y� ̰g������ �R{
��D��� ���_� �{�$�� ZY*�0f �ܞ�R�� �{�C�K�=� �_TR�� �|hI�� �e��Ę�������oO? :����tC Å� X�+\�k �=U��� �D\� �#�*ʘ d�-Q�T� c0����=�X��(��?G Q�3�xO� ������ ���̝�� �0G3ڨ�+ ޠ��ΐ���;��J�����Sû`VVuQ4�ۂ����2��}F�3p�]8�̇iIq4�!���6
[��0�Z�>qN ��(3� ^���'8@� h�i;�R�	�W���B��@X�� [���+��!�����$å��`��Q	� �P��K�����B���З0 &�[�(<'� ��xf˗� I�3�,� j֋����=HZ�k�wd�j�u�; c�^PU�B�q �9�% ����?�����J�'�e� �9��g,O��,�f 7��$ ��,�	�^ R�/���(��� �)u����@�3��N [��h$�l�q� �����`����5@K����ɉ� ���Rr^��`�@h�]������Ӌ= B1ه�¼ 6	���r� e� !#��: VS���W��?�31�����K���'I�� YJ`B��� ߬4TǕ� �|�{Ӄ� 9�R�	�Y��i0!� 1�ԣ�  �?۠����S�0,^}�y 烐�5����7�`B)]�����M��#� C���\ �n�SA.�� ���#W�� �@�l�[��u'��C-��\�[4���;X	�(��ᝤ: �Ʉ��95�8Y�ІQ`�R ��!�����@4��:�w^)��������Q9+$ �F��ʸ. L�:
�2b��.Z׳ 4�M\�� }r`1�� o3� ,� ͈�p)�]*Ԡ���\�t؉�Q �U�s Ăe��� ���pP  �+K[��i |����/ _�Xp�([\�	 y"]Y�t  �R��X� ���d�w| �	.�>cP ���R0�� UV;��S*�[d �/�.��T^� ִ������b��B�n8	�h��|��H�V�� �W�3��G� �X$Z-#�� �wyo���� ������E ��9.À�X�� J���OX�<��.��
��@a�@��� �+��W�J ��1�!�2 x�c_b}@�� �!V0�1&B�]�k\�.�>	wy b�h� 0{���< 5>e
%vj P�*�g�� Ll\A�/�����{�bYS� 5آ�?UR� �1�X����	 &�p�%>���Uh<�`��pY��g-�i	�������t�0X�Y ��������fZ��h�W� +�$_�B���:5���<E�
���{����N}�sB ���\�Q�D?� 7�Vx
� Ef!�W΄�t�sX�'��7�Q� �Ba-ùP ��O�$�� )�
�[��K��B��@гX-TO��쨴" 鮅�����%����l��b �����]� �!����<�v. ��	*��s��"��΋�P��iԲ�u��� �S�Z) g��r��� �_���� \V�d1�3��Ā�H�;$V�?̾� � @w�� ���`Po G
�X�Ch�1 =��� O��V� ����_�hB9�"��)��r���ɭȋ��
$J��h~�]QA���C �� �YZ�'�� ��h�0 ���%�qyr���� �h��E� qHrAO��} ���-�� Q�Ǳ3�
 R�O�$�p ^(�W��_V @����=I��Ǭ|�!�� �S_��`I�z) ���1�z�%ԥu�p2X "UӅ7��`�Ѓ����_�$�3T	�[�*���yG ���'8� B ��6�� �$"Sy�T�U� C]�9�� ����Nǿ# Z���
�m+�K���L�h��� fpe� )� �Q곺�>-��X�i�F[�]�������Y j���Em��(M���)���(�0 cd"���� �@�hbm�| )��~u�v z`��1i�> S�f�-*�{� .�4zT��R��2�+y�]��-��g g~�W��2O���bG ���ܴ �\����~N Z(:�[	h� "�p�λz �%T��� L[� K	^Q ��C�� ���$�P1� �D���(��oz��a�5����`� �V���Q����%m�5]��x��P�"!H#����; ��OR���c^��. * ҉�� [���N�
 �h��B^��8�a���z��*�!���� �L���04��1�P�����r�Z�J	��� IC�PÞ
�S��{���`��o ʕV�F[ S0���Y��
�8���?"Z#V)á3����H0 M�����h{ p8�܇���}&��_�`.\ �05���DXS�rQ���L� 1ԛ�A @dƲz��� �Z�?#� T��/ [
}`�h� ��B��^����RW1݅g ���Z�l%`q����?�^&�~Z_f��u��/� ����q ���2��	!wc. K��� �'|u�) ��	\+�0 þo��軭�Hԋ
 ��G�� A���*�8�"ωt�`�>.�0� ���~� �ab�,u# 3�A�ٽ={�)� ��v	� ^R�+� ��4/8tJ%<}� *�vy� �D�������1�za%J�� 
�q\�D<C ��^���zr ��%q� G����� ���<��)ʉ3 �N[aE�� ��Z��"� @����M�buj:F�If ��1N��!L� �Ы�͗ ��Eu?� T�8��Y- |P��y� [1�� W�8�� ��tOK��@���d��e f�w��(�8����|�i�!*�i S���V� �]D��EW��F��n��	��RTE���p�� �}=�	V] ^P��Og+��ϯ|��h�~ ���D�yj��������+� �T�	��i�#:�ƀܔ%whf� �W�Y��� .	��I� �L��0 z�d��3%��<r� q��0� �_���PX&�[x (��/ ,=��%�_9�� �?U
�b  ]P`O���-��	j .X�� �� �@�qB ��!�U�����В�/?��
 �ȿuX��%�n �/�c��+�Y��w��� �	i�
/a= W�*�+��п�l>�O�� �_`!�x �
��Цv ��R&J��g�Cco�^0Őۗ_�p�[�& Xh.f7%������� � ��	�'�N-C�x��^Kc�:�\�9Y!�8)�t��� ��Am+�|��P`�x�� N�C8�.��i� (BMտ��
 K�%ʷb�2t�z� 9��˗�4 ��ݠ�Y��8�]+�Q��\��	`�U []2\��yu� �(���뷘\D$�s ����(��K����21P����y��Ƞ��^ ��c"� 鱲��� �0$��Q�g�V%���ţ��3|��}�� �sv���L� P��0gZ �/ Av��ٝ�� i��5�͖��� VT[�	��9 ֜���09�]�R�B2�x�ںXр��)� �'�+!����1 �LvY&�b):�`��yX]-� �~S�\L �$%� � ��Y�=��I{8 �{F�<V	
*��Jq_2v�� ޻����no�%���$�����D= �v���SH� nJ@����M "Q#�a\�$�0�? ��ԏ+r���x' �$����( �71�� z�2��,[@ `̍��� ���Z�� /Y�a1l+o�S�;��[R)��^M�>�$�f?z� �_̡�d� ��]����� 1}�N2�5; ���&A��U���l�30+�d��h���&5b� ��N1� �-��W[u�Ph�J ��U^�c��  c�h_!�а� ZW`(��F �����B�9 � ��s|*�4������ ��I��4yT e���p��/ �0(ԗ��ů~�At���psK'��La9���i#��� ��`[1� �������m� .�K��V '���(�]3 ���`-h �U����d (R���`o�&�W )[��$R ��Z���� yH�ðm0 k����bY�\p� ��oB�� �L�ı�	f�7��
 Ia� )� [z�=/�V �;I���Y�o�]yő �骙�?����M�aT0�f !+�܋��r/�O���0� ��{9�� �~���Y��X���W+�I(��͸! �e���K�Qy��� .4��BԪ����g� �ޗ� �[���Ջ� w�A;� �Di|�(��|[ Nth\l�ӻ ٌ>am�( �&��1����F��eh����V�=�~���� ������_��[��x��N L�TnfrS ;R����:P�N�*�t��u2� :3��a� U�~(������[݀n4Y�9p1 ?S<-����h�O �( �Y��H]�?6. Ӣ��σ��<1��]�x��!�v�x��%8�����5|��}�p���� 3+��]�i� ����Y( �B���]�X���� :"��t�X{�B��pE� ���UL �[ʘ��A� /(��R� �$�1ˊ�f/� W٧uh<�.��Hq��&�� ��:~�}up (����B	��� �ȰVt��3^���
�\ *W�6�����1�L! �Y �+h�.���b�2�_���� >f��J� I�V�A֥�+(~���
��Y�Fe�)� �����!��Mp��~�^�6B�_�@O̘Ź�������8m� ����Y� �P�V;� ��W�:(�Ɲ\���I�j\)% V��dp�0�Ku������1� i�|5K~%�� ӬȐ�H9��& �	�� ��ɱ�j/�x|3)Y ��`��m^�� �����Xl)���@_�R��,�+G �Zݯ�s T	�_ M�� H,���{�!Y�G��X �`� ����i�v� �@]�a� \���`�3�[ %!Xulj�0� �Z�� ¬W~�ci 2XPs:#Z� ��5����0��G��N[�n�&��� ��%R�p�5 c�j��ҿ���G��p�����`�N ��� L��9 �Z\E��������ƭ��������aC,���ڰRYESlT �u�j��h }(��O;� ݖ��rXD :&�+�0 �{�A�� 4��(���<Z" �+Sq_<:� �,�7� w 湈;G� ��hS��� CF/��;�s��T6D����@� �83�r/%^�x �_�` �@ ����� ���+��T�����-Ulx9k������� %��QN�B ��)� L�]8ohU8J ���t����|�*�!� a��� zpq��&� ��/���E ���)�DC 3���uw/�� ���_\�LAF ����`� �6"ͨ^ ��sB9� �xP�4Ȗn��`L�0̇
���("�_n`���N����W �?Q�ع�� �w���)�[�D�3�\J�X���\P��S�1���������]����g ����O9�"} ���M� U��� .���°;� R�4A���� f�����X*��� ��0\3[
��e�a|�)� ^!�r���(�i`h6V��GHLe�| ����M=�!ϑZ� H>(�����W@�cJ ��
h0 |$�G �M�+ �	U�ʴ-�9�g`7�ڹybPւ ����p�Y^ X�g@�1!~ڴ���U�c>������k�Y�@5
�* )�Z[V�� ����3�8% e&=0�4Rh�ka[Wc�`�� 2����P?���	u���(� ���3JK�� ed�iȉ�:�w,�� �3��_��$/ќ U��-'"�R7��X vu�zh�> l�"pR�8� n�E$�	 ��]�i QPV��-���&��0� @����fE �j0�Vh< *��rө�E4�kK�_���2ZX���r����� �0����v�%����/�g'��@
.�* �0Y(� b~9�J{�=	 ����\)�S��7���x� $h�-6�Q=i�uf�[x�8#��L�c	��͟�Y� ^��A 02@�$ �Q�R��T U5+�@'�	W��*��;%��XF���� ��Y,B����'[W����H1��w�D��y$� ��j����� �e �Z���%��]o��a�� ���:����Z����ݸ ߬��{@� O���� 2����|� �_��}� =�K�G�6 B�
kP V���ƾ�p�A;x���	t='<�#(�	��� ��P) ʕ�8��� �˽IxX| _�H��� q��;����7�� !�~�k}�Z �P���Y� ��̄��� �݅�P!\ 1�.��� @�X�-r V��+��-�^npA�4��̀����(~� ��0Wf�� &�����;��ӕ�0� yN�����A ���Ě-�� ��YT�U"_wOW0�h�[f�8���]Ƚ����w�Y������A vj:�b���  �U��˾� �n?�]s�`0郄���=A���L�P{
�)�3��hs ��J�->�T л'b!��Z�t��z�h �Q W�@���� �c�w��(/�� �Q�㜳�� 	�R{�-߻ <�3���	n!P� �C[ ]�}"���2 ѧ�;�)RV�.�@P��� !���>����Ro�i�+� ��1*Z0 �wJ���,ד ��!݉ @�Y��{�8�@d?#�
��B3͡<龽�t��� J�!���	H�� $��jbZ@8�Y��_`�D�	p������ �K R���:�D �j�Ђ�89v��#��>��r4\;���щQ_��g��cFY��KK� B�������#�\��4�G>��� ɓ��&� }l����.8�^ �I��3���������% �O2�-Yo�U��R���E:� ��C�r� �U�����&���RvI
.*� �B:� �Eň��/b Q�!�{� ����E��S�zb�L�=��?'U� �g�" p�Sh�a��� �;��-[
9F�h�p]A cM;�fQ� ��E��j���H�ւy�� � P�ٖ<h& v
$�ʶ� % �d7-�� ��a׀� �� �	�� ���"�
S��ܗ���G�°�Ke �����RA����i�� �)p�&�]� �(��<r� ���+��b��� ���Y�N����y�	h����C�+@U��JG���bEw� ]���9MT �+`��� �Q��(��� ���󓪀� v����� @Ì� O:����)�Y�1\��%��3 � A����(.ʒ� �U
�~� Q�T���-� ��Uu���������0zXB�/p\C��n�#���M��=�g��\���� �BY@��|� &��dv�z ���`G��9 g��@�� >Ofȁ�%=?Q��	�Y��> T���|�� ��0��ZP Ƹ��u}� �#v�_�]kt� �0p��	S� ��Y���>� �N�d
�� rv�3(X� �h�L�&0��渦 �N`k�a�) ��V^p� Q��Щ�s`��j�ཊ�u� ����/s�D�P�]��.��m!k�`���� �%V�G P�	����0 U_R��B� ��X靵C\ ��E%�/�(�	I���֢���K����� 6L7�wP1S ~(��t��I C���<�� A���׉�� ��9	��u� ����0 �(J�{� ��uS�PW �����#�{ Re�hz��8���@uLg_] ��o��h�
�ʇ���?%}H ;߄�쪦 Y"�ڃ� �3*��0�� �X�ߴ
�� 	����r�¾SиvQ�9���W�����= XhtTg��iJ��rO�.a9b�����/�	pf�^ ��R�u�	������ �aX?�@�c?	��� ���;� B����>: ��(�6�Z��X��� I��
���[�2��%�uW ��e��{� �\΍)���sg�ep��A� �ĕO�	�d� �kB��m� 肠�wںZ �c������p� �!཯�k�;����� �&��D� �9��� V(�����p�y� S"ƉL�z �� ��$ @���]�CR ��[V�-� ��#G����R� n�Q�6*�� �+	�PL�J �a~��*�$yp B�3���� h@]�q��v ��w�N�J� �>hgH
���`�(�\ � �:�0M��������YsX U	ڽyE���V(�1��I�Ӏ+� X��e�V�޾�h:I��� ��ZN�
� 윴�R�����(ۀ��槷Ϛŀ׸[� n	��~�� z�|4�x �"�D?�PW?�N�W͉ǀ�'�� ���3a���Ϣ���=x��zmZ��2��w��xpv )���ep+"�K ��TȮ��ޅN�t�Ϥ!j1H�{������Z]L 2P����HXx� �Y*h�%� �@o(ٟy� ǌ�����\��(�J���� r
�銉CQ��e� nJ�$����(����P �����N ��/(]�db9�Հ&W^�p�J ��Yk�m_�h�����/���r�3� ��(B�wًt�!�C�� _8�%���rAjn������ G[ Ğ�19L$ȿ �����Y ^�釷`y~��%�B�$b$N=� �e��d� j���,� 5�c2�͸%�QT' �h8�� 3�P%0� �	���mo �,�Yx�9ơ5.� ��ѳ�% �~TFu�� �mH[]�r�!^�V�Q+K�'� 0������@��w/�{ i�+�1��9�������)ԅ�����$5���<hu�DO���U T���I�K� +��L�4��>�w�V� ��^�A*�� �4
�&ਦ�p(�ͣ Ҳ�@���p��jIK��P �Y��7H� ��Z4�&n;N��'�G�<�1��08$ۀ�V� ��	�-����`��� Y�(���?t� �qU)�R� 㤒�[��3�w#�T���@�Zu�4� �1E �?�~XuJ[�U��ȯ@ ��+��
� .��X�MG R�FԐ�t���(�d��� ��a�fJ%� y�)_�`���[S�#����� 	W�����?V�����^1�P<�ո� X��$�lb	)�Ry}ܚ.��a �J�/ Q���~�:W`���]� ����?� HZ�~ �_ǠF�7�t@��	�%| ��R0PJ� ��9$cd������ 6�����W0�p@�m"�� ��뛃Lg	M�@ԡb�zX|�X�\ w��R�Ͷ��� �ȗ��/ 阆|�b�԰���W��}e�A���t ��[Q�j� (6��ח� J���Y����
����ƺK)��(���ׅ4F��N� �u���B_L �E�0�b�d ZU�m��k�;*��4����m� Ƹ* � ��b�0�~3 a����\��R���������]�	�Y1v ^Rh`e ����6���j_�|� b V�Y
�|�� ¹�C\>X�� wE_�KR�?��+6 ]��CJ�)����V��@�hU*� ���k����b�(��\^9 Z!���`���M�f� eX�vc� ����� 	�t%Y��� ?�!��\��d} �� S t���*�J��|f��^�� ���~��� K"�(&���lS�L @�P��� ��o��JA���Q&�5��tG �.�HO�h ��B����� 8P�������� 6��k�3���6 ;��*G�	ѯ0+��0 Mv�\w���`8�]���~ ����0D� BV	��ۊT����� _]��1K;� �a�|Z����4 �#�X( �Of���&7Z9��a8���Y�� +kc�a�����`	��T�=,���l��/�$	�.�a� ���t,�>S }�.d��������ƀ�f!�� �팄��W�r����_���D������;� $��\��] %�X�&1�?�����"��#)�$���!��Ա ���e'BC��i����@��� ��G�-�8%���ck��J������Z��=��W����+� ��S�
/ ��<�p#�=> x�� /��dI������ ����%� ��/�����d8��g �`ˀ�3 [����4��"���N���� 7�>�1�Z|�
2�� "�!=#���oF@��Z�,�� n	Ӵ8� ����_� e����d �^�*A)r�H�a���5��V��m�� 3��7�+�& �G�O�8�� ���X�@ѲlhR�22^�� 1�ޫ��x��� +?����`YD��%0q9 �-�߁��� Ղe���B ���@\�&��������	��3�>pCr[� �uZ�0���}%�nSl�d�	� \P���`N {җ��J�	 ��u�I[؎�. �kX��D-9B\�]V�=�?ȸ���(%5�����t� �����C� s��-��ؿ`;��� �� �B�}V>~ �?i���% ������C:�Qy�kST X �WH�E ���v/��}� Aa�`�1��?&�6���ΛKS�Q�X�&�	(°!��'��� ���N��0�s�{��d "�p 	��L�u�  8FH�� ����vQd/��� �U��\ ����6h}��균����S 2��7��D� ����X��$�= ��	0[�q m-b�w�}�|� �Huso �N ��f�$�4���^�n	Ws� ���G\�bfHR- ����N� �P�z^�E ,#��o�a eh%����� �Ү�W��j�o���|��YJ ��8���ְ �Px�X?
0�f��Q���<? �Y^�
�r �Eܫ�F�f$U�%(��v� �-��m~�ͺ9 ?�u��P�Ÿ`kH�w�Q�ˠ��rd�.œ�X(�����R���$�
u�lY [ �K��� 20�.�� ����P�� K�3���2 �0���U �)��#� G���*� ]�+U���� yp�JZ��r X�1�v)�j�(Ǻ��.+�H�'�e����g�q��+�9V?	��� Y�t�JƁ��?Ф�L�� �� a�� �3�m���$����C�B���� S��d+��ň ��0� -!|������[��`��@+ PĞ�"(Q?z�B �0Y��������Z_R颊3���<(���yt�� �Z!�ҿ�A/'��0�� 	�e+�� Y0���=q���� (�3c�}� ���h �RX!T3
 ��{�'�t� ��JI�����U�@��%�'RH�� �}�_P�  ���N�>ɟ���̃� ^!�D�j_ ������J �	�ZBQ). Wь'��:� �(�]��d ���.�O<@�h������PF� ꬎ,��^ ��1�/�q&+� �W�= Ţτ���6�P��Y1��I:�W �a�c�L 2v#����Y ) |�S۶	 �͈UH�+� 3�qN������	����j8�,BY ��5���� *�A���L�V )�o��!�L�r Z�¸��;�8��J��#S 
ϫ�/��� L�42uF^ �gtH'�$!���Pa�-ĺ�?:D����O��uyo	��,��9�l����Z A�/%�":2��?�<�}� �	m�b�W� 滅Ѐ���?�-��u(�X�'N�|�,X${ ��� �u����ܳ�N��W U`�^'J���,�Z@\� �6���V�i ���Z�!=�u��c�'�md�$��| 녡�H_6Z�@0��[J�g� �\����%�oK��`��G ��,�v~_����\�%'a��S�� m����U�	˹e0��JM��� �! �f R�������P "����^j�r�8��.�&�Eu+ ������fDG�� U�2 X�*i" R�A��  ��%^���fa�`j8�cx1,���}!ڷ0Mw|X)���� ��i�V�g� (�C���� o�w�t���B �߈Zh �	 ���&fS�쀷�L�*/������n� �v�XhrN �܊% ��� ����_��]*�`��qo $��h-ZE���_��v�u�r*;Q	���1�� �;W��Dz� yk_�L[9 +hՠ��� �1_]I��T`D�F�;��Y�`LN�} ���P����U��(^
�����:���� A;]�g����Ip,Q�-� 3@р�yZ ����%�^ b�ur�{�* )��'	�p�J���Pm�*� UW��] �[�AZq ��D�&�� �<ux�`>g ��q� �2Q�ڔ�| 1�V�� J	�(Ù �)��1����a	� ��F�,�>@ ���T1h��[V�;��`�t ��1�+a<zL8V Z��iJ�7 ���k��,fb	��0�w���h] [TԹ��� �(j�̡M �h�-������^�\� Ԁ��B(w�<�׀�]O�Ff��=Q���� �� ��A�:���#���Y[���(����Z��xD�����hxpu����[ �a�DW/�,�@����p��j)�� ��A  V�2�[� l���<r� M6�>�ޣ =H�9w��.  �B��[�^ ����Y�:g���0�ݟ��% ��hkJ`�ױ��z��(,Pӻ�G!E�`\� ǫ�����L ��^��:��k[ �Z� ��|�K��� 5��d������]r�� R3ʺ�=k� �V�#���U�R�f���.�v	�i8���bAI) ��r�1	=������@����R�>�� �ٽ�&�Z �`�y�aC�( ��ہ�~� K�Ab|�Q�>����Ӄ����?\G��"���C*��/��� 2�Y=��e;��� U���O �)P 3X��t�(�zw?�G��p��S :�|��� � ��+�LX{�T]������� ��bY��	 3ԸX���`Y2@ -0���D� ��{���p� t�J��� ���5P@� X��IY;� �q��Ǝ�PHf; ���!8* ����({< ���l�H�� �Ř����1�� )( ���\�`��S��L���6�=p�4/ ��	X�#*��>[� �N��_V�)��d������� ��>�C�<Z �\bf�W�e��a�ӐX>�1{��n#$e���[) J;�iS���q�L�� �A�
�! ��C�T؇" ¯�d=BP ��Z	�y ��:�n�9� ���h(|/ ���uٴ� ��`�hZ/ ���4F6"�bkP_��0�E ���K���
Z��عR@t ��q��� ��ƴ]���(0�)���U��߽����n1sk�+E�.�! �	�:�7� '������o 2��`��[�� u��!�Gs}@P �B���(qP��~��UQ�x�.��v ��b(�u ��U��� ��OG@ . ����'<�ͨ��-�� M��U�B]��H�����L� N���~[�+�O�(D n����� ��QV��Mo @�^��1�EE� ৏���؃齸.�Z�E%�;�y�6� }���*���	�J윀s��� {0:�,��~[ l������ ��M  v����� ̐����� 	A:��;a �e3�%��( .���h�G�=x� �A`l����hC����q" _ �{U�&��[	�����h詯(:�ߺ%� �N�$�1/ R���Z���@Ϊ׹��h} �2KW�G �<�,�N���)��*v@��� 6(]R���������p0��@�h^� #�?騪�> Z�p>	 ���h���_)�J��Ԁ ��T�6 %x�+D4 )�h��	��P�~ o�) ��
���	��]P@�u�R� Sp���<���1�b�ŕD� ��I�՗���^٭'���{����� ��"�R��5 �t��Z�<v���y���� �X�e ��+o�	����~*�|��� ѓwn�5}��/���Z�o��z`4�n�d@6�^	 �uX�Kѷ8 ~�1w�O [a� �0 o"{��� �|I���\�0���O����S0����b`�[w� ���) �{� j��_�W�= 2w	Q+}���ď���X�\;C<� �"Y2�z,@/h>�yN�EU`����	���@�	��6� �W��è�/3i�� �p�c<���@�hM`�ӒDW(�߀*>3�;R[?� -��`�ƙu� �sp��� n�?�Tu���� J��)қ�<	I�1 �������a<�!MN��������� ��R輙N��K��#tJz� )�l�v�( ��Z�xr� *\�(
����C�������m���0R��?�z �0Ų�	�r��X�ୂ� ��x�n��.�H �ـ�.  �')�}�	�N�Mn���� �,
Ʉ���p�S���^���* ��TV�2H�8I@.ں X+ђm��Ì�d`Y����|J|� �Z4�T՝ H|���&! ��/ k� �0��� ��
Ly�w :��M�4b!>6� QA�&�@	���S�f1�hb?���Ho~>
6 ��bhVNk Wd�'��_� f*�	�( ��aXX� >E�
�A �I��۹/X���Q`� U5 ����� ���xvU�������� �����:� %��~�� �tkg �
+����N��[+��\��O�% ҪxZD'>����,���A* �J#�;0S�](u�	W� X�z�� �	�*�03�Q�m�����OX\A����p! ̓ȳ��� ������1~ݼ[� �fX$� +/}����uH�%T���޺�qf�^���n\ ���V�f!Oй�ֺܜ[ o8yxK���$^�����< @1*?t��vH�Ѐz�| �5L��9?� /�t���V ��xU�����{��� ���!�1s �9/�,�c 3�:��4V��w� �%��܈� �Y��_�« �Ľ�[����l ��3�S� \1ͤr�Q� �8l�"��'�H �{J�W ��}�P%�� dDX3�.� !���?[u �ۖ�� |��عL��Ƚ���� ��J¨�P�޸~)��� �UOD�^+G�_m�K& c � ��N�H�` 	�����sB ���.��H{� Y!�<��I \PV��� 
���k=� ����}^�q�IR�z۠3�` #�1Nug /����埓(��� �F �@�8�u��N����	�Q���:���� 2��90� ����}Dx- 魋�U� p��9�XS� �ч�0�@���
�_��H��0��\�%���>��f9�-�\ wXzn��LR|k{� 1�+�d3� ���	_� @]ȚʗT �p��x�K��$ �W���H����X� �_j�U�; ކ]"�h ��M}��'�w
,�|ǐ��Y�Xk�} X�ܵ�zE 	�����i}r?y� ����)�R�- w���;�K��XB�v,� �2
�_!���YH��`��RZ�[�à�κ �f�J��c �*Ɛ�S�i0_��)�WX�� l��A� mJ��4�� -t�QZB�� ���JTGO *�@[��`�� �h�C���t ��^{�`ZG ń!��I �,O�x�� ��+�%��PY/��U��?���A�y�c�"Ӕ�ȦQ  `�Li{� ��Y[�� �y��G	�� ���]��F;�4��u��� hS.g:`0]�@�ʁ�#-��B� �빚@Hؘ��vկ\�h��ZA�*��6��20 l@dL�-�	�����0"9��TR��_�V' IU�-�P�%�= �����v'�Ul�X��i��/���>V��  ����}��rD�j��� �!"`V ���F�M��P��I�9�e8⍀/����Z9�_�X�|Hi���� Q)��k� @S�Y�� ��;���]8 �Rg���0�+���s )�}m�����LD�_ �G�"���Q��0� 5)�17O�����{)+ ��_][3�yS �fP�RT ,M�� �.�.eڭ p�j!k, ��]ҭc$ �L�/r@ �X(�P '�h�\R�a%ТV� �_��%��� $5��� r0)�� '� ���e!��:�	~A���ش0���;� ��9�,��+ Չ����`t�:���<�?Jp��4^z��V=�'�Z�AY��r/���U���Q���v��y% �.�V�	,� W�p�A����p$��{&� �+	!���>#�ʜj�c��@�ow.;窀]hBl%���KyH���7u'*D�����wYZ��4q��� ����2�U�S|�����MX�
y I'��>?��� �Y�!�%  )�;tZ�� u�Gۋ�2 ��m|&��� �������	0ɃA8���]$���s�@����1G�I0��S`�$��� ��sh��	�#�P=�M �BH
.�Fi �O^��� Sy�˝h'?��Ԍ���U�@��� �'�p2�Q�8 �Ä_��x� -����!���q��v�{{.��Յۀ#������+�{�y��ؐ� (&t�h�d ��ҫ���+�z'��K��	 �9ƥ����v� I鎝%� K���!ɷZ|F�س��]A�Y*� M!�9)� �PI����� ���~> h-�3_<� 5jn�˵ ����0��t�a����06�.#�+��8ϰ ,O��.�{�1Aj�o��슾  �[��-���N�
�ڋ ��dXY,�s�2�'��1�� �W��P?��8KA?��!�"$�� R*l��� �v	6)�V`ȉ�u�O��(Q ^ ��Z��� s����� ���7�� F��/�BU@ ����| pc��r��JO)aa�2x 8s��X	��?q� P�1
�|� �:�,��IZ �	�-n��� h�R�GK���:o�Q�2ѽwb�a��.&�(� Ë%�u�� *M�	+�\f i�>�� k)��	��� ��`r�Y?�}ߏŀ�]��p�����0�9�ʔ��&�\��^\Йe;�
?��:3��g��� z½1�GF [|Y	��(�� 52{;��'f����	�O�v� ��\��hT���&�� 2Ďy�nm� �~�^���r��{��?�[����, � 1�0�XR� ʵZS�լQ i����� 2
���* �f�&)�" �%��Bt��b���-H�
\� �>�ĉ�HW$=��:�Dś���	��?��R ����� r%P4�� �^LE#�Y�|� ��;��bN� ���� ��X�>'� �t�r��3� yCc�6� �Y���L&<�	S��� ��%6W� �\?�HY� ��eK1X� �U6��?` k��!Z0�r/ �%{��@ hG�8�Q�TNʡ?���؀ɰڒ� �@�A�� ���^�v �K]zN���ݸ�-Q��D��@�`$� Lg"5�ݫ�au� Z�Hf�1� �x�!���:�_ I�"u��`@�p�� 2�c�L0�[ ���K��f� �\�+�$�� ^��Ӂ� 4N�Ԃ��`; �� I�����$Y�� Q���b� �
��N�}S�o>��d\���b[�d���f�*j�<ގ�&��� '"�ك�b; �{�B2�� �C飖�N^{�&#�� �@���?Ca Z��xW h�i�l�� V��k�<��u����\�t �2�R���� !�����S ��7�pTޔ �Pҕ�f� \!�X��R �I�H-�^����w���� ��'��!qR �%�0�O ��w�i�+<�1�������{��)�-���p�o ��ɸ�0 �X+�P�` T�f[��c��sݗؘ"� O���U���!�o��p��h�%*�1���QV P
��N��^��	��In �Ү�G�0 f)�LZ�/��X�9'@p�	
+�ZUŗ��f�*���0�c� n�`�^��� �A���2 q'W�$O7�$Y�� ���X�� ��/�Ip �jr��y �Ҭ�֮� <�*�Y�l� @(���ޢ� �Z������E'�K�)é�����W 0��T��� A�O+��� �"�7�� �S�e���s0 W���Tb��8�K�L�0�� YI�W�hD �/��o� �Q��mH �؍�`_� �013�D�	�m�-�� �UJL}�¦�(~�H��*���9R !�s u/	���P������P���y?�>
�4��R ��d{=2�ۘ �*?ZX NI��� w��=������%���{�L��V�����# ���^ ��Z��� }��z�p�7>K���O��� J��ʄ�/ �a�X�չ 郚H#I���{����X�pX����%���� 
k�q�� � )��� �E�X�ݯ t,�	�T oa��C�\ rQ�;��� �3�
Z?� ����!�Jp¯b�2��Ȓ ��f��D��\� 6�~�'5�!h�`W� ��X��S$ "�󚓰�� ��hQ�* 1��	0� �g6��Hś VĨZO���)Q�èl��@�cDi !�yf�B��
 � XYP *�%#�JO��B2ʋ�x� ��߂����X&� 	[��!� �Εk )�X�(�\ ������n� �M9�=_�s ��;$�1 a� �Ɉ� B�>_��0�[��0&-v=߄��P��fR�Pj� ���s��A Я� ��I ����T� �[7���V�^;�YZ�h�H�`��� _�]�w�-�8勀�P3%�p `��U�X �O:̕h~�,�34Hw����@ ���������P\��_1�:�@�Y���(�5W~TV �|�I�� K�V)��' ���D�=
�>� ,��P�������M�GЄH�v�bB`��� L[�a#�	U��} ���<� @3)�&��9� ?���W >���� ��ըۀk ��g���V$ �T�b���(w�A���e��ظ ��i0�JN���{ ��=�� h�U��k�.�F� �.���Q�� k���Z k�&/��. ���p"`�q 3�hH2���} MT_�O! ��>ɇ0H(�� '|]r�t�� ��{�-1�:X��+d���4�
����ٲ�/�Z@'Ƞ���: �a�QT �� �����.i��P����H��X�؃���� ����	˰v �؄0��� �^Τ�� c��OV�(<�x��pj }UF���P9Ɖ ��p��Z}^ Jj�(�' �d���5�껛 ]1��W� �$�<��� �� �8����V
�q>��v P�s���A{�K���(���$�� i"�q^Hv ε��1B��9�_%S�I�R �?͘j�@ ����w�[>��G�`# �3])B[Z� Oh�J��9�� Sսl���,�� X���3a;��x�KX���L�p����-�� 6ӯ(T#� �g� 	�+� ~�3(�A ��vW�;��;��|a��0Ȇ���R�t��[�2��\�λl?��1���L�� �����.�=YB�d���p�=��Q����H�j�@�kdu���`!HŞ��)V���(�� oCY�Qł �'B�M{>.2���.��yh�#�WA��S&bK�����u��3[ԗ��@�#�H�� �kG´�2 �U�65��{J L1���b>�o fP��U�� ��b� 	ո�+c�7-�Й�� H�|vCz� �T�R.�����P�%��-���1�- (��_)�� ��/��*@� �{bQp_����g��D: ��P� ��<v�(��/3�xp�q ��X�
 �}����hB9 ��)�+'��q�I@v	�j�-���K>�����2	@?�(���	\�0��! ��Yӄ5���⁰ �k>3���a�
h��:W��Y��X���Ā��� ���&�L ΄" �/�:(��� �J��Sp�l  �������ǵ���]`���|"t�_��f Q�ñ�� �Y�2�� �*�v�9�j u/
�RmN�!k	�`�0 � X;�M&ͨW úB(Nq��'"���0z; KY�1�XS�E���/�}% e\m	��Vg �3��8�[�p,�"5M���d%�+��)���_Wf	0 ��+9 ����a[1�����k��;�� �IY�	V+ �W��b�� �uy7vS(�� `%�O�A!�d��H��`v�� [x"�����L�`��݅��:� @\3� ��հ�� [
������V^Oc#�е�& mQ��!�Z S�j~� <�qi��A� �;�������Z�U�h3� ��v��ˡE�av@���Q��H�!��� ���D��b� �&v�ۉt���X@-Y�T� �9^�1�aO߀�#(�	���l ���LFu���'��U��� @#Kӗ��Z01���[z$"$ �����@ ��ؼ���u�a�Iv+��� �i��]� � y��\�6<hs�Wݝ�i�~�<�	ܺ��0.QZ�`��$�K� `��8�p�X� ]S�t �[~2 ��	��� ���u�$�P��� ����� 2^
��<TR{� X�u���0�p/<���^ ���ʦ ��'F}J�� ��lE����{!���='R� w�4���,eP�@K� �	!��(� ��@0[4=����fq�k��RBȻ����'���Q籋�� ���. U�z��Nf��9g'�w{����M�� h�/�<'� q�� �6�A۵��?XU�t ������e�`�>b����k/� [�n�ONz �'��p���q	 �^�!�-����L��K:%��E?9� ��	�?���)�0��Xh6 |3S[��t� ���f%� jOw�ิ �7���K�\�, �-���+��4�;�h1�v �"o#�O�� �*�r�8I� ^�c����|R�i!� � �a��0 �_���wT� �J8}��.�:/X�`�Ĳ��=f���&;���Q�`Z  ����v
�h�m�a�o�%ظd @�3�Y�� j�&Q1����)�`�%��d9�`�3*Ԝk8��#,ǨX 
��麛� �0�`C�w�\�� 6��Z :�$���k����Or�.�(���`q[����� ���� ���W���3��)@\R� �UVa�B��?��LZ	8��}���.�V�s}����A��R^KZ���=���  S�]�! �+����� #/\�\� ��`�h���$�k�\B	 �I��#7�� ��g��� �޼)O��.^L� `���({>�!P��KX �5o��] a0�Q�DPW�v �[��Z@�ژ��Q�,�;2�E �����> �^���K� �`ŽZ��
QF{%#�s_�<v< $�� ��ed�� ��1���ؙ 8l�g��?ހo�+>�( *�P���2� �#��B�y ��@�hKf�,^�(l��R� ˺Y��) J��W��< ɿ�_�s� �CKr���. 볲�(�f�y� �U�������AL�ʁ1 ���I \Zv*��� �Xa)���=[� f`2#D ������J�!bSt���,��&I�ӂ�K)�0�a2� ����#6�`�B�G �X�o�u �wrA[�<\ �{�P�� ��O�H���t+"v0 �P�@�!�� �X_?���s'����
[=%D��d��Z��+l �����| @�Ѩ�`� [hM-aLm0.8)u ɳ��ks� �i�g� \$WxI(�	}E٧�����-� �|�����@�( �ͽ[�	 �DTI�' Z��Aߋ >���M��� �����n3��q1��sJ" �Pܱ�SZ ��/�(C���^J���`�&�X�V=w����]�eC��8�����xKu�l -�(T��� ��F�� �Q V�'0�� ��I5g�
	��X� O�_e�;���'A�/-��P�����S ��\���.�n𯀮�ş �㼃��LN <�
>�Y�L�5$�] ���خ� )0�[��r<�ƻS2����� �h=G���t���N���K�� w��
 K%��� }���� t����8+>�V��I��=��H-jw�ߚ���G� �օ1 E�%v� KHޅ�� ������ I��� ߈^ ����g[ !��W��(ɶ,N��S������ ?�3"�*�ENpy �)� ҇�}A>^]����� 1
��[Xo:� �N#52��H�d���׿m �h7��ͯ _%���VX I@�P�iT ����A�� �72��� �B��W|`xt�g��PY��� $�K�+x �ir.�m�� � E���$�"� ��1��px Y	ֳ'Q ;�J���m�^9���]� ��`G�0� h� �U�� DrS��I��H.W Č!ȃ �Aj�a�k�@ &��M/ O÷�����tia�E�}� .���`��D ���:��@�)�_ _����b�� �D��ٹ uH���s�
 �hX^��?��! �0ۖ� P9����L�� ��!<�%a���.��� �Yv�	�d)�݄-@Р�A�_ ���h�.�FU ɽ��1� ])	���
\ e������ �K��1��� F&��b��ڋ�����?�ʠ�l�x� i�W��ۭ 	h�8~oB�b\�
?� Z�$T��Q�@h�<�F�Z �з�w'}* _D����); OسS-�� �	����H ��Y�!e~�z� �%����a��U���|V��� Iqaj�<�R�(v��_u� A" ���;pSX���O(�x	̏��lJ�4� ��_�e��� ���\�/K 	Ȣb�Ú�)�Q �Ĕ(�4D����C����� �@N��7[� ul�mbW� �����I� ���N����)�22 A$��[��N�_��
�� �'�~�[� �,���� \DO��%#Z ��cЊ��;N� �&���=f�|ѱ���  �%����.�( eO� �� ������ r�V	B�X� �`W"\�E� ��MP�x �w2���/. ���ZY�FE �;I��%�~ }\�:�� �X�y0H~e��:������ I{t�#�� ��q�0j�$a�  ��H��8 �l1��G�p���Y�̀� �QS%(��� =L�FD�$ �b0�J�w �1s��Y D�/�V{ ���s�A ����\v3�	V|4�� ��]��S5 @�QRY���+� A�^UT=]{��
��� ��-X�z� �v�N �� $�RW�n� b�:^�� %��|r�� V#-k��d�e	��@A%Jt�� V����` ~�/Pn���?)'X��Ü А���� �}��CP4 ���1�(� �뾫Ƚ��R��V!~� �=ד�� ����x�^x	p0��?� � ���Z��;W0�}u �J[E2xP����@��� ��L�-tC ��ej�BT� �g ��G;o ��PL��!X @]1yհ%*~�\l \����|> �	���VUi ��+ΐ18��ĴHҞN`�S n����C�5
Ϻ���� �+��V�$ q�r'�:t� � |^����� �Y�-����a���<T[� {�����H1� C?
�Y�� ��c��� F;Q'~�� ��K����BF �Y.O"�Sa;�� ��%ī v�gXG��� ������ 5�Y�z(." �h�g��8�H ��&��., � ʃ��h� ��IO���͸ Y`r��q�Jh�d�� E*�cA� ������� ���hO	�-��p�>
ۀ�=A����0�w�`N1�7	 ��/̜9���ʼ ��.S���iT�Q J���e(K� "����G� �xbl=u3��� J�" a�Y(�*�2t�}�O@�a�Q�!�/@B�� `9�v�$"��ӹp]��� iUa6�H�䆎Q�T�o Kܵ� ��Y[�\ ����!J�y �<ľ/m��;�| ��G
$;���	�`8�\�p� 1�\�&�����V�+�4w�^��!쀁-����1�f)�@�͹�� W��H�� ~n
 �ZL�b%Û���fR! �7��P�� �x��D���>���Hn������t���� ��F&��	�?�GT� ���wʷ �8_��3�#��	����` ��v��X��M�	�T/A�D��Q� ~�Ⱥ,�� k.��P` ��
1�*� ���6������<� 0%��3��@��P���'�\Z� ͽ)ǈ� �-���1Gy�H�h�����I� +���[% ��xL.�� �lzi0��>|Uɜs #ف��z! ��W�d��PX2 ����MF ���^-� 
��'J����.a�<���z" 1���0�������Q�F ��M�P� ����	H��$���A� c 4��(ſfG���WZ\SL ��X�օ6��/�����>���n�	B��_& �
��"��@A�� ��Gv�����'p��R��,S�7 ;��� �ªv_��8B��0��Gh	��� ����*�(�ʀA�� �����������E%��U`���=ޡh���@x	U��G
��P��;�� �=(� ��
�_ ��@�K�Ŏ �t�/��l��H" L'\�D3 �1p
`����*�����T�X ޅ�P	�_ ��ߺy�pJ����\� FNe?��H �75	�l�; �S�����s@s6X:� B��]�)��y�P��� �~�*-�Y`7�����BJ�'�`�"�8�N��G䅸 ��� �'D�Q���w����9� @��Y�,JXh/����* ��P&�_�Z |�RI(@=��u�O�hܾpx�~�P>L ��_붇 �ڻ �)�� ���BYf}|}� u��>w��0�h��I�>J��֒i�7Њ����F�� q����V�ʘ@u�� �R>ā�� *�:�+�&,K��2Z��u ��Q� 	�i��a#>�m'����/� �hk6�c�� ʻ��A9P >����5I�|��@���R���-�:. !��V���	Ǽ&��`�?K$� ٷ�������2��p`� ���V�Q�-F���}�O���j 
�_�R�
��t� ���\P0��&RXZu��2��(�� �X�u�PL-A bj$�Y ,S���]=Ey;0�~4)��`��%�vP$9�7��<ɦ3� �f=��	h�� ���� ���� fV�*��]٠`��Ր���������ڙ����� �G�T'� �I�w7_Z��A^|��� �����0�x ��G��'e��4�!s�.1�� [��W��H˞�hO�)��A��*pŝ=��T��_���<�� �q�K* �5�0Cl�J^� ��AU �~�ϓ���	_]�{���m�U��HK% 1`�(帑0��]���G��|4����@ \��!��<iN��ʄ  �ث�I� f���:B�(�er��#�N}YL���� az��x� R���h�o�Z�d� ;��t�j>����'B��;c`\ �UV(IT^�p�?�a �rWsVqQ k�ߵ��u=� �d�F�� ��ُч����
I��c�$�Z�XVRz�<�m¤�����Q ��I�xk� b��0�e� �.�F�M� �r�xE�� ��Ib8� �3v�0� �T��S1 ݷ���$D� @�<J(�E�� �v�b2�ߔ��٨\?����SR� N(�� �h-؎T�jH ����,Z��xu h��g o|�Z�� ^y	Q[t�Y ���r�H��	Ia^ �����%�� ��� c�d��1���3�?(���;� "��!��|��@Up�_K�0=���7�ib�*��� ��0�x�<�_��D��Կ� � �\�[� ]�P%	��K����V�@�1�] ,�(������	�`h���ݮ!�� ��$��6�}� }��O�� Z������ )�u��� �?�j��Q� ��a��f���zH��_˄%���ָ�L*� �W��7w	$�� X�H'�1N���Qԯ ��m�Z��*|�� ����,�)�1����J�ܑ��� �Q�ݹuy� �G\6�O�Ա]�+���� ������G �3���Q�p'�'� 	O Y�
���%��]P�� ���HR��C �m��0 �!0��Y����9'�s�j��H 1��҃�;�?	P�}���vwD��b�UY��h`W*���u����� ~(���a$* ��z�ӳO�����3�Ȳ.y�t�h�:0�$r ��X�*J ���4z�� e]��R�ǥ�K'�nW`L �h*xXV�e�� ��@��Ŷ��Z��,�� W��U�>g�wM ����?] `�_����9����@��+�
Y~�� f��ʼ@ �[#�Yh �a����X� \�����J 0�R(Ÿ ��S�qPvL?)���Y��hX p����~D��]� �a�E>��� �"� ��I��K��R��L 4H����힤�k��� Z�U��/o}V�T�@_�� �1��?A���_�y��:�����¨��E+���4aJ�Z��nR�t�|A/O���V�#ϵ{! ��=�3%���FGTs���} <��`P�,�$P�+�,@�J 0�B u(�� �ɸ����l���dp]1 5C�H3�KT���%��� � ޯ�y7"8�� ��X�g N�̭��	V �I��A�w X�J��˰ ����l�(0�`��J�����) ��D"���߷�����\�|�x� �bN>������T����~&	�� h0t� `�ן����O����WU0X �<���D�+@�^3�-��*���Ő� d,!i��� Yu"m����U �<��f����ƀ6l�T� �h1���,?~�˜@�<^� 2ZB6J�� 3X�[��'� �� o�\ ��L��� 	G�A����D������ E�>)��Z� �=�_鉦�$!6$��#�Z��p -���õ� t�&���	� ��w�^�� ٗ�G"�ߎ ���E� W݃?�L+	�:İs��Y���2:N� ����_ :�z/�a� ��ވ��� v�OV3Z n����^`� yO��l6+ '������{� ���s��? `P��k�
��W��� 2����^r| �[��Yk�'�"g�7
aUDS0�g������ Ũ )K��'��� ��AqD~�n �`GF"�^! y�	�� �3�첱h; $
�,5&pb��pw���d� �uJ�XUj��3PwT��74%2��� �'t�������c�π��5 ��
�V1�.	�v����X��� �`�1ɰH \#೮QU7�`�����, X�J�C��[��#�Ǐ��� �Q�8��? ����ѝ�i ���
��&n/���Yb�c[� W��X�8�y��%��b_� ��Z�(�� ��4�h�P� ���Ŝ�� ܞ��71o ��S���d�`5��n�" N/��W� ��\S��Y �]�����x?�>�tv�;-�2�� �Wƀ��s������SQ ��^�/�BRzf �]X�� �U ��
���$� �ZS`)Q���z0J�2�W�w�� ���p)�'h �І��|ZB	^W� ��Kn ��`q'c�~r� 8�F$�7� [hSm�Z� �s _+�F�~ q-L�\Q�N	a��Ӳ����d�h' p@�=rv �H!��8�� _��� `�\KH�� ����A0?{� 7�[Z2�RU�����i1� �0�s���� Wo�t\��1 @�~R��E ��揀��a�V k�����\!٢��Zx� -�)�E	Y� �'v�B�Mi @S?
�� �n��;�� �<[&7��g�_6���#�Թ��c� ǧ�1� �H��� ��K%�� ���I;C�� D
���!��5��@���n� �&��I�s��b����� �蚣�&F  #%UK~��,�!8�1|�p�R
�9�ǀ��"�J+ ��_��0( ��i��� �J.��F��} �3=*Z�C����)��t@� \�h&� 0�yH5}� ��+ڝq9P 0�T\��vj�tWb� p���h �M芙 1���B��W��+�������A
��)V��@��3����u�����@������`��L ��� �X�� #_���-��gr���=Ob�����6�}y8d� m�P�B��$(ƺ��*�̀v����r��0�&	����s 尽�X�2>Y �Pt��{[��k �f	�=��mU���j��/y� �X�4���p�� ��	�r�!T���5}=����q� uyL>���* �	@������'
�E� �1ino?� /��,U9^[rpZ��S�RZ�>�ȡ��A�����3 ٺ,��#!����@6J����c��I�a��Vo\w@H���Q	�]�au�P8�; �S�1�� ���	)^�� hVU��� jӵ�:0��S��OF�`vPY�j���z1 ���l�+87�5)�� �j�k�w4;#T2�]���>q�q�l�}XϦ�+ �y�@G� ���c�?( �LO˙ \ǃR�IV�;_� (�/� ��+@5ܨ� ��h��� >���\	� �7K�-]��c���#����+3$	�y��&���ޠC%Lgo�x�1��&P+�@�@�����A 깦��O@����w�Z ���p����(�. ����
�y ���l�(�Y~� ����.� S&��U����H��e&� ����z����I+ \� L�� �Aa=1�w6pB� F��� �J �.-�^_��wtý���5ه�` ����%�W��k ��V����|��񝐿)� �̟Y19�"~����*� �W:�^��"  ؚ��� |�u�Z7�L �*�p�� nU�š�ʺ	�z���\��z,0�e T�p����E)��������4.�3x<�Մ�Z��0 $at����@�
��4��� ��/ �_� �J������j�j��0�S$��1��T�Q UW��� ���� $��{' ���(����q,��I`���}#	g_Z�v� �cM�K9"	ƨ�z� ���~����xN�@�L�5�Z 0^-fn  ~R������� %��Z��.�b~ �P��W! �3uX: � G�d�����ۀ�S
�X� �1��4 ��2�S��_�^ ѢG����̞/@����
R�� c��2��oE�/���}�b
� ����D�K_�-3$`[2���+Z�Gm�W�-��^���A&�M�ha��+��%�QF'��h���?�c ��Y��x �MK�H� G���,��#�&%7�x
�� �e3�� �H�1�? �	��~�=�p�L�6��� g�H^� [����`�v8 h'\���
 K�D�z@-!v[� �j�m�/l�.vh- �
ٹ���� ��[&�:O� 3-_�j�� $ZFR,d ��U��V��;�i N�Ւ)�	.w4�w ��[\�� I�HD%rv �!�)�����u#ڽأ� ��·�$� ��*�� {p�M�`�� ���YV �H���%�z/	-�Ӏ��1�� w�^2�.��_�P[t߷1x	4�Q@`��=˿y��I� g	����G %v��@��&�� �P׷h-< Q��)л�H�� ��:%�l\�P����o�$�� ���=n�p� �Ⱦ��(� f~�Y)a� Ʈ9_���h *�5{|�X "��'`�O
���tj�� E^�O�6:�FV���p�^�� [�*N!� �9�F��dx����Y��� �|	S�o%>؁gT� �*�I]� a ���@����u�L� J��<y{^���&�׷0��T���Â�l�}n ?׾�2��� �6�=Q�� {�mc��aH+�X���k ��L4�6�����q�غG���.�fH O͖&��S r�D���G}� '��@�5�� �Դ%�� ��� �;bG��G�-Xg���L �N`�9 ��
�o�l \[��F,U �ë��#� ���_���aVNz�@�� ������0E$� ��>��� �x'z&K�� �_ �º鬷c� u���!a {e�|���j�<25���y�� @�P�8�� 
����	:�0a�[H����� L�~5n[;��������o`?.��^���7 �[�(�S�� 	U�B �/�HK���a��V��� �DB��N�� WK �&��[�be�ׁ�S	� ~�p��/-j	�����]���CU	 �\�G�  ���'��Q����r� ��|�r'3L���P���K��0 �j����< �5>;�O ��d\���v�kLq ^��	"�����U��� �2�Y +�둡��j ��dD;XhH� �+�E�i, ���m�' RSqb��8��{���1�����7@��Ӳ �(I/h�D:���ͧ@=V�ԽM ���݇��* �\��
c� �����( �b^�)ɳB<���$��`��� ����v� ���(�	Ű�Y��A ����{Q �(�֟PR��^��	�x�Z� A�(�&�}.�� _D�� K%�ly��0 �,�X[!� 	�Գ��7u� �t��خ�� �h|eن�4 "����`.�Y%���L�o�@=,��f�:I��v R�x��� ���:���ݖ�� �%�*0O �7�qh�8- ��զ�I���< � ��v�%�w b������mP���k.�  =y��;�Ӏ�GH���X�� ��Rj�0� &@
��V��`%( ��_+� ����4�� ����c��� �]��� �B��2��_�`��p:l��u�O��� ���џ`_�^���O��:��Q ���B�[W�	��� u�9b� 
<_QO��a*�N�t����	�R3��Ƹ�P�Ol�0��M��W !���<�� ��]v��� ����-�NH)�@�\hA�� ��>KS�`�|�cm��������u�)����
��/GUD-�`/M �}��A�	  �R�>�7� v�dK��A� ��f!l�w^ ��)4]���_��	��*� �5�R(^u#�D���K�n �I�W4� 0iF1��C�)���|+�9�� �z2�^��?@��1�P��[L?��h!zb& �@��6 ��C��Z�����p �X�fP��\�0K( 7��WI�] 1��_�\x ZřrdX�� !k�`gA� ��G���}P�_��p,+
2���`N�L�
䘜M���h]Oc� �u�:����W�B��@2AH��� X) ^τ�� S����<i�Q��c7@���a����C�`��	(��}�?w����-[ZB� �Hv*㰫�� �4T�� ���):�Hu �"�ZQ�<�M��鈰���J���.a�����_�Z�]j;�쀛m��!�2�+�,�-�� �"�!�O R����Z(-�X~Y�%��u �Q¤82�*���W&� E��^S��> �b(Q˪� T�Y�g BL�'���{x� ��>�R����[J�6v ���'�0{�>Q�I�@E䪆g �����,�\)�n��v �X	�^ �TڊVΓ���w )�}˵x% v0��2�S �$�� ��X��qj�T��4�=�3�+� �����)��@O�Ӌ
" 4�Zn�<�}�!\P�85@rZ봃���N�| ���]�`Z=� P��F�'~ B�EMtH�\�� A�W��3� U��pQ}n�$o$B�(kV b�Jh��0 �����_.�i�? � �O�E ����^�� TR��*> ���<��n&��W�O�*���(��ը�@+Q��� 	�C��q�z���h 1#Hc/�0Ћ��VqS�� ���o���['��}��亗 ��5�j��"�:�#l���89 �K���� U����!º�:����9)�\�(b@;�  ݺ���נ� �-zB�� P��`�W�� k\�f �� ��y�g���w� C�����L/'���v �I��B�ɪ �|<���*;H��tS� �A�� 7RU_���/�L��]	 ���`䰵��&x��P@e� ˘�ض%sq�`�l.*� �S�̕�a�F!/P4��s�R Z�u��H]��Ь��+�V�� hGY���Iz�E�ϻ�X#�[ ��u`��<��A��W����Z� �X���	I�A�B3_v �d��\� j�/=�V��̡� ��
�	��[Հ��D3H @�,#˫% !�Q*�<�'�-A�V�徰l�%$[���/��b�P�N���_��`�� ����'?� 4��5	k� SQ��+� 9J�6,Yo ���8�'�1 ��s�Kv��,���� �i<Q��	���p'��^8 >�|�R�\% .�t�u� 1���?)�A�0�i����2п� V�9���Q 1S�(J�@��?�ҒZX D�%�>��V�\��8k@v���10� �0�ꢎ� S�?x\z� h	ڨ� ��P���T ���b�݉��I�
��cؗ X�-QGA�o 9�5!m� v����� ,�'	x�H ��_B�gLb���뀋�/�D ?3���S� �a��Zfx 魻0��w% ���R��� UQ��kΟ9 �*�C�� '~�Ȫ!h �W�V�7<�K�)P�}� ���쿀G��W[N_Έ�/ �?I`w,��� ��\��_�>�)�e d7]�o1�Q���Å��)�G��D`�n}���=@��OJY:����͎̖ ��-��/%�� I]�	��r i��g2Vz�9�' S0.����(���U��g��� )�|h-R �Y޻J��q}:��y�c
�`��>�+��[@�2Ɨ ]%�P����.xy��p� h��[�Q ��i��� (̵�$|/@�%	� P�(���
 ��z���b� ������@,1� ��;��;-:�|u�)G ��X����L�1׏�r ��`�j�� P
�V �YU 	���T^3xt� ��_�=��K 	�Z0�f� ;+QS��� �Yp��[V Lw(�}7��>�$^`��R�@\Vˠ�o�k0�NH �|�@" !��Wtj ��+D� ������' ��:�>�d �K�̀�0�J���o��H�X���Z(׉гE���]Nۮؒ(�p�1P���4�y��
%;��W"�0�z(.)�3 y�_�dU� ��1� 7�A[��J������ M�v	�+�# �6/�[-��1� r����� �a�mC�A H�0tJU�7 9����:�� �}���n! ��k��+(�H������G R�>���a o�.�l�  z�'�1��B �0v~��� 	^_�q@D Al|wT�� ��W���30,�"y��t �>�_��Z U����.	��:�� sо5�F�D �(�V�O����v����ɑ�����U@	��P�� }VǥT?�0���pQ���t�~ �ah�yR���� qN�� �λѓ
�`?��� k��p�2��X4T i�[�� n�|���<���� PoN�!��� Zh@X���)۾�3a蕭 ~�&��� rI������K!�1�k���� U�-ܦ,8گ�"�2��\ ��z�J)����S��A�&��_]�v	�ƀ:#�� b��ɼ}���2�k�?��� .r��٢  ���b��X ����0�J�P� AbǋƄ\	!�@�%Z*� ���O�� �!�]dFP �v�8�hKc����ӷO�����L!�w���#�a�	�I�� ���/�� �,����t'�����8��Y 򭐪���}�� Њ�	m� ��f!���F ���d/rֳ��y���t
 ��ʂ�+�� ݰ�,�TD��L� zJ��5&�%.��!0)ź�"� ��`	
�� �$�宁z(�ۅ �hY�1�� *v�]���6~ur|+@���S "��\w�� <��!��H, �Vl\C� h�{�5�� g���XY$�JF�����P��]eJ���@/~� �Wx4�) ��UɴLi��u ����h�V:ψp�X�# ����� kmݡ���9 o⏠��G� ���]x��� �n�M���.�; ,*/1 �-RɌ.k�K	���s)����vS����Ɓ ��U.�[` P���0\͸ ��@N�!� 
ٟqBhk |_�M.�[��+�`Q�z �*���y#� �F�r��9Ŗ ����� �U)�_� �H%J��E &��/�p6�3�ӬZ�܁ K'���� �i�n,a{�q4��G� \��҆ �]V���R��K+��B\ S%#��	h �@��;� Pv�M��f�QX���|�۠�`@�1[���� a��Q��Z| /hv��g��mKC�ĐH�{V܉�\�h �P�?�"���n����9�K�΀��f2���P���+�>���=3_�T����Iv ��
�\�� ���`^����Q���w v��� ��hqj'\rtג�xpT����當����tx>�G�, �·����W�޿t��L�5 �*�_ ���[��� \v���A h��*�f j��n���� ��QyW%|8x��(�~��}$FzRw4 �g����^����r?��0���f	�Ӌq�7o\P �,��$ 	"�U0�\�j��S� :̷,��0�W^A��@��l^ $1��'b,� �&f[wce��kK��%��j�a�� ��A���q����T |̜�V ��@)���_^W�J������g8�N?����~��|�!	 n�p��{�3 O��v�Ha G#�ä���8yA�^���� ����Lz��4� ����&J����2H�v@���
A?����1��P�ж _o�N���` $��Y�Wh% X�S�j+N,��� .{KvΠ� �� �ѽل�� 2�]߇	ʊR(�@Gޕ� $�<�!ˉ �]_ڒ	 2�h�`l� �%�߬�J� �R>���_� g�K��@��!�XZ=�� ��Y`�(x� �a��k��� ����ǳ��{@ǻ�+�� �h�Sm(ٳ ��Rn���\da�- ����� /��|����H| ���0��� ã[�'� xM
�*)� �\�h�j�8 eJ�	�Y� �X�{� A�`6v���
;ți��N�d��[�\ W�2���uM �鱴4��{ �A�kp�p� �S������ ��8�5�
 ������c ئ�C�<�x�a� ��:����Y	KSC�3�B �a���h�3P:���홐� �{�a[c �3Ӏ�!F&��i�:�Ԧ` 0;GL�@Z t��fQ�gtPW?% /h�7��U�fkĀ�q^b�'��G����Wa NX�8��b )��7օ�$��sv�?y���	 qђ��� p���e[�	?�^� 25A��-@�p� �3�%�s�g�Q	��7P& .�� z�Ļ#��"϶{�`��f S���	�|� �^�-���yq93� �QW`b�[ �g��� u��P����r� ��1�2� *���ʎ �ÃՀ�� [%��aA� 4�8�( �$ !�S��T �I�v�d� �u.�Ao ���ƴ�% ����˧U�#<���6W
z�x�[�9P p���{������ +��]z�~�MZ�����r0���C�d�z���+����_��S V(ʱ'u� ��Y�3�x1�ha�n�@� )�YȜe�'g�X���h¢V��W.��_vA 1,֒�ۖ �B��! �(����iv�a) �YhN�� A#x���kPW|��w��ȋA��D��~D ت���!�<� D�;��9�0 �ҹAr$�ؽ޷e
�.� ���ˢQ�a3�ŉN)��{ ���2� �_b���/� %e���R�Z���S!�)��� ��*e��� ����a�\ ����ь��H���
�h�"�� �-3�F��� ���
�� ,�o���� wE�-�=R���������)<|	��t�Q80M �N̟�pi} �2�\��� ԇ�3��{� ����R��� �0�H��1 ���9E)���@�2���f ;��ԎXv�Mo ��Sb�� ��!�A@� l�	ZS�� uȯ�/���n Ad��`��%8>4$"�i*@� ���
7��0 ��'�� ���
� /�M�4a�c vz��=�K ��}<Qͷ� /�s
��9Z ���E��H ���k��v-�^���� uX.���� Q����*H��|�ֈ�pf�	m���_�����ZD��g��si8�]�#�Y)�	N� �k�+�$�� ��L��ڀ �=[�`�<����o ʶ�I��H.} �h\� @�����:�t!�;*��U �dc%B� !�K�����	l���W��z�XK��豼��&0) ���� h,�%`��R�_��8��k	��vZ@^iQh۔��\�����" ���rx�m? �_�<�#[ ���V� �,�	mN� �J'Bp��z1�� �����8 �>��H/]MQ �p�b\ �;����7 ע�լ(�t/UFV�q+���Z h�D�aH� k��#n`J�P7V_ ;��RU|);^�Ը� ���9M�D��7����k���{@��c� h�_L��+� H�y��w ~��BV���=�? dP-{� vIH�\W�~�	}���@ �D.�B�bt�<�q��Q4� ��`��' ��qSd� _N1�%�:a�� �{�I3 ��n��>�ր����9�w� �}J�� #���8����qx@�o� �1���+� a��^����e 	~�,[�.Z4� �1
� ���9�,�oO5������	 �Z��@�(��[�!���L$ *Pb��.� �-��HU�}� ��"��	� 3����
��F�D~���do��� /*�1ʔ�|B�K�1�W�>]���`��c��iD�{L	 ��إ�XA��������- �|~y^��i P��Vb9�[ ��N�-� ��l*YP Ӿ0����H
y-O����n��  S�6��U*�$��� 1Jz�&���Ƞ�����-�r�� �I\� �pUH5MpY 0����� �ݯ�h ;"�/�y�� '1���v� A�>k�~Wg��0���x ୃ@()_� �P�fX� �Q����(e�[Y̒����.�ft&�%m�� o3� \P��V� �j*��@�h%�B�W0�X�� |/i~�} �R%lcH*�H�� U��D�� $z�2@�R&�!L����. ȉ�Y$C	��^��h?��T�`!Os�w�_��@�5h:S@Zɢ4pa ��fN/��K�ۙ ��:�w��c��4M`��%$@7m5?��I�� +�u��� ��#���� [M4���{ hNl��W� �'���� �[�`^Q��� ��{�vB3 �VCf��* �u��W� ��
t~�O x��欣�z�  9�Wڇ
� oø�&�h$ 1�:�^�z}�R����#������kX���R(̺�"��e� ��M`1� �L#N�uĚ �1�o츐 ;�~ƑP� &���@!	
��?�|��|Cͺh����pZ �O%��4�M~���e�}� �s�Q1#�j��k� �KκX ��C�-;RG����2��ǋ�� �X��� �3�Z+��� _� e���JS����>�8�W12��|�ֆy� �R��/��F `�X	�'|t� �~ xR� ��^eP�ˤy	 G��*�#��>X�wH�a:"_������%4��EWx�5;�����H�Ȁ �K����; �*��͑� i��.� !l�x��K񉣡20�w =�*��Z ���i[(���L@e�U@�%N ��(,��4�R`�2�FJ �����I� _�yZ��z�F2'��V`e�~��X�u �6U��? 7���])	�0���N@�! ��Ϫ� ����b��x \h�)����*� ���� ����	W$� d�%Q� ��@�A /~���G���;���n��lĞ�!�� �Q�{]0� 	FS�P׽x�t���b
����B���hذ� �>}~fa� P"W��b&S ����	1�h �ƽ/�~? a���:�p� ��L2�G�b���U'=� +9	��;�"rf ߢ� ǥ��YO/PP�(�?h����qk�=�r�0Ź��������΃�: _��.?��
�})���J{� ��%����pٸ�+%}�:~N�|_p��d� �r��P�b���%�� �H`��л����y ��^��y�g ��@V���r�d�A��@{���i ��ʀ� ���XݐD�#��m�� ��"� �(�y�N��w�d�����t� .�kf�ۭ8 ,��B���$.p�@Vir U~�]�-XX�� L�a�u|��/���g ��0\�H� �M
����3 ��]A�(��� �����~"�Pa&(�Zc�8^�y����8�)w ����Te�U�s �9o�;Ӱ�	�#0q]P=� �K/(R��� �f:\�A�|:��+�̿��� qY��z�� ���0ΰ��¨/�l���� *�V5r�:�� �
ʁ�w (��"Tj �@����]� �����hC�L(���a�� ��K	���!p�I٘��|e�<�
�ʸB��_�{\ /�m#߼�`x���Ă���HJ��W���\[s �ʬ���;��P��� >�������3}����+� .L���`�� �X*�Zh� i����@D2 ?��s��e	�@�uW �9�}���>�z��X@M��� ?�k��|� S0�Ef^)uҠ�$���	 !�}{��� ��m(@>u���t�ȣ�� T�e�-.�
�����ɰ �h$43�Z 7�OE���X �!������ �)��$_fA��ú������ �3�(�4Z��_�N��t�r@ɬ��ݞ������> �qH+�}�	 Z�U�����&��-�a�H�� .)�N��� ��ty'�X�[ /�����[�f1҅K 죲�b`I��	+��� �a��V@Y�`.�fb0���_� }�@��5����[��A�- X��xc�W �Q| ���u� �S��-�(�I�H��Ze��G^� �3�U�"���sSH� z��>q	�T^A��5��� �}Ž�^ et��BV���pX���0�Z/��S��������J� �/-E� �$Q�y(�<���#���1�}�� �_�WL� (���'�G@ aV*O��<��� 	�CZP($�i �Ї�7� �t�y/P;�� �����Zf �x�,�(�~u���aÀ�! �����&�bS�N0���3���T@��� ������@�������� H�o���x V�y���  I������ �=@&� ;#��2|�*)	����_��� ���0 b(�v�fY 4�B
�"��X�|�H� �0��X f	�Z1�^ ��h"j�=Yb������2ϰ'0��b����W���S  ZRX)�a�,����H��Sw�@���,T ܂�%�H�: 0P��i$ lkJ~�'>q��f��� �����Q ����-Zt]z���{Gu�� ��B�V��� ��;�ĽA��^�)�� 	�!��,w�ċ����$ ��M`�h���@�,��G k"� ��[�@ɼO��$�x��y����	 w�H;��� ��%�물B��.. �\�{Q 3���јdt\83 =H9�]! �Y����� �2�����>[+ ǋ-��D�*�`�?� �����4� z��c�� �0!Ѻ �[R۹�Ç��������04��@q2� �?E���%� t���X-�2 �[��.�f/p��"��  ё8��HB` �Fȁ�	�}u��� R[0� Z��^a���v�� ��*�o�l ��=��+
�^��� �Q���% YfC���$:d� ��6�a  �+>���y� *��(�bX��cw��h�;�߰�� zK�SN��r�o6�+�0"��ר�Z��1��O��o �h3�45 ��i.+�H D��S��` 	؞���* ��C{��� �A@+5`%��8 X[ۄл�r� ǵ>�א �S�+�d���������I�%c�7Gf������ �}?���� �G �K* ԃ�}?�\�Q �W���		�7_^  ��p�Lܶ ��n � ��sZ��:��� (]�3�Lx�K�� �#b�q-$��C XH�%� O5|�A� j��� E����h�w�r}*-RVn�Pa�ʖ��H� �ǳ����s� ����XyA�p�v�P���S�' P��0��� ����v� @�_��Hh5������ͮ0�p� �	����\� Q�:�=?B� ����R f,n@�G#� 2va']<E{�����`�53 ��J�_*�hn�ذ��y����C��(oĳ���̄�;��>���l��ٵ +�χ�	�XW��D���b�0�P� �<g@L��x ٰO���� ��Z�����(.0�dXp�|� ����t��<� $Y�J�;��7��� 0��\��.J� ;ơ�֢< ��#�e�)vKLZ> ��� �b_Y�Xw ����gB�?�c��R^��	�D�� �wS�s $��"Fc/ 	�)�V��3�$@�<�J|b�ߘ�����R8k ٔ��z�� ��[���l A)ٸ1f� 4] �+,(� W�'_�KQy�R` �^[�# �S
���������Y��i1� ���k� � _�e�a�;��� >A0���j9 �~N�1��5{���V�Mp��i Xº�lW�Q ��'U��\�	 �#�w�7�j�"�dR���0�Ju��^�	h "���  ���1��� ]��xKj �T/�@�!�.(ї葟���h^L���%W�0=�2	�Հ�T�/ �C����z4 �^	����� ������\�� �F��1� ��m�J@u�ŽV`d��\9 �z T�b��Wpu:=����2� ;	 ��+1:p�w7}�� $�ML���Ź 0����9I��*@�G ��A��؈J���\9
��3¯��Z�S*��%V�	�A�� ��kN� ����p- '�]|XB!������k�0+ �[���- ��oB�5O�
�1�.���%� -��й6Iuy0 3�[��S 8h�4��� q�c^�� ��B�˩<��5��;���� �
�>�Cu=>S ��3��� ��N��?[��X����PK='0��!���V��" �/,$�Z�� ;�l�TP� �'mw���te���A�:� d���aP��Ec3�"��WX_vOw�s� ?�K�, �4����  /�����0x F�}y��i����w�n�>U:���'�N�q�v�@�f��
 �����0�z� }�Nʴ�l� (-�JI ���k�	��E@�)S &�|A��u /�}L-[�$ cń�������2QQ��,�IP`�89�	�8T� ��1H �*��h~� �?��8� �Eo�]-�&Vi| ¡��6 t�Y��+X��.��`��:U���2�Y�m��`�	�
8�\��  �U[Y6ꊃ fA��Ҧ� �����DZ ��0�NL� ���.�Ah/�~��3���f �+�A�r �;,�: ����s  ���v�� G�	�\�a��>�S�7��L�L /���P�Q խ*�)a2�Vk"H|}�� .��Z�R�� �Ln��~�3`��1��
 ��%���$h EY�?��T= 
�W1�� ��	��q�H 
0ޟY�� ��-#���.UL��\�G�����h���aQ��4���@��UZ� *6�D�0 !��4ߴ�J�5(�R�E@��eZ�qa/�z� #TQ0���9�+�A(�E� �/v#�'R O���� �[ !͒#�\� ��X�^�< ��e0��z V}��hO� S���T� ǎ��\�o� ��a%���� �� �\�n7�3�p;1� �2k���C� TW0K��q ꢔP��" %���/� w���֙xM $"SP��������^1�/.c(l �D�
��0_�Y"��y5�ظ���?��\ �Z{DAQ#Pq���� `V�+���:y)�> ?�C�n��@��������=��� Ҝ�����!��� �])jW�8\�}g��(���<�׀_�,'d\�xZ {��� ���^��?�,�[-���x ���1
�X�6�7H�`"� )�WZU8 �0���u] ~:'a����IG�B��q�E�� 0�X��.�W d�h�(	u{p��$����0 �"˵�� ��GXR�	��|
XSH��	���K������`��X� ����|�Q!?�9���� H���$[Z�G����+�g -N��_T�0��X�H�]4������#� ��e��iĘ� ���(WQ� Ź�1��$ ������$�.� 1(v�a��s��Y ��h�.��:#�&
�W`�� ���$I!� �̊��� �ä	��%�|j"iC]��؃ �Wՠ65� �!Ū�� y���Sf ����Ӊ�* �[�Ε!�\�Hl| �5r�@��� ��,� �u	��� `9<�0�Ȩ��Ð`1�W �o�J��_��f���.�C݁�Vк���Rx`���']��X 23�*�4 �Hѝ[t ��R1��	�=*���D����� Q�V��Ȅb ��*Z�{�p P�JU�� &�bv׺\H�"�݅ ��tk @�2�h�`6. ����_��KV(�~u ��v�ªp��Z �CU!�h�A+4��͝ �7�HУ)�'�@��� �Y��"wB ):W�4� �뼢员 p<�M��[��}�N`]8 �>R�� ��{7� �&�� �\��_�]:J/�JW	����ܨ� ������\�<�<�9 &࣒a� -jt��| ��	�K� ���N�� [���<( ���^�r���bQ�~�?6JH0� ��S��Q� ��`h�B��15���a�=���'�+u%>]� �ɂ[ �j0 ���h�_]� ��&!�K�( ���\�<N: �X'����?��� ���� >����(� ���5��b��Py�\h $��ufQ ����Ő����i~ � �X�L� �����ܝY ��S(� �
����� 	�TF*a����2�؈�N y�=��W� (�&�L�T���� <�|��P ���q^ �-3�v	' GZL�d��cI��@�49�~� ����}Q ��Yh�� L�5*�(cP �Z�W�� �p�?C������}q`[�(V�I���	h�~>\���A�Z��I�u� ���{�����E��r��L�*�! ��z���� K�5���E`�� ).�R��� ���	X�� h�|{�}N.L,	���[� �T��l ��'9�~6cP�ј%f��(� ��ӿb�2�x_ Oڋ��.	҂���2]Kk� �:��3_�x ����R�,��?&��B(O/f�� C�4 ��]tP5_���Z^��3{�e'��A�&{�hr �	ٺF3vl ���R^YKh��$�R�/R�� �y����Ј�Ǻɿ0-D� 2!�B�]�=m#�1��N �*��&�K���� USѾ v�� �Æ�~�����%[�#	� t���Ĉ�q� ���fzU]�`����(��� �s ���[fhy00ս�� ʳ��[	�S��Q�4�� ̡e(�ta[ �k���|� ۴6�1�xN�! \'�i@�+o`�2�4�����h]-:�e�0�(PbݼPO�� �0-v�L5� 	���+����� !�	�U�& �ݾ��z� `wP��@Q}�IZˀ�:�� �|u�^���v*����$� �A����m f���%�� ����0vZ9}T�cv�4�" ��@*�P� ��(ݛ����㖠|'	�1 ���07Kʠ@�|M []�A���� ݓ5���# ҟƻ
щ8)ȅ[��O�q �ˆ�*���+������� ��-�Xv�8�����P0�/0�- ��9�$>� %_B�O^ 	�6����� �Q������"Sj�\:	�`��a�����p0,ډ��� p��K V��sE� \����t ��-��E8:��� ��$W˟���������7 �z��?� Y\�h�<�=�g �	���Qb �A����~8�1��m��#�h�N$�"C�3 �2 �����?S+ �J�ؓ�9�N���P�^�E����� �D	���<kɍ�����Y8�K	��2��R@��!ý4� $.�nZ����z �DY�J�^ �aG�qnw NL��� ]���^��:2u��w8��
<X��\�^ �Z'J�� �z!)����F�5w�f�iz��I[-�)�N�S����C�Ao�]�U�0I|�?;@�{��fq��W�K0d�P�H;-/�Y,e2� ��OL�k��:�T A�q,� ]���� ����L�\ (��[b.���ˡ��`%�Y� <�$������H�Â���w1~ .���VJ�ՙ��Kç���^�� �eª�}� �A1��^{W�����/�,I��"��T��A'Y��,�`貰�K�A��pXԉY ����h�%� aT}�?�Q}� �bf�*�_� �F� k�w~`�3 P�0RX��� S��Y��M,+�� ����m d�!��- ~�_)�q0 ���6��`5 ����_N� �ǹ?���B
�a#P��.* V��'3� ~<D�н0�s�;8���%�p� ˝x��u��,�·�)��� 8��k� �Nfǵ�|X ���b�h~ Y���0�鰸 ��)f��-����@���	�s� ����( AQXY���;����{ ^S�c��v ���<�O�$�F� ����� ]%"��� 1�R	UG�< Q�j�wzN _����k� #�V��!� ��M1ٜ X��'hJ�}����Y������'c܀ω ��L+r) ������V�޲��+��U
p�O�E��5�1� ]��,�����y���'�.9�x �!���� �[�@p����
�)�D� 9\ߔ�$PW s?�R_Q�i됴�����Ead��ZB���%
�v�@��- �s:O]G.�9�q�ݖ��� [Y�`�o ����8�� R���5��m���à(��,��W*��c N��o &f<Y ��q��1���zO|�U������1 I.6�~�.oG ��"�<��G� ��� �U��kAP>s��2�����{�-(�hAt�lb�_z�	��!�B�/�Ծ ��l��% �Vva�81 ��Sn�p	 J����L& 8��.�,3 �J��vb�'��uE��0�&��0����m�`��o ��ϛ-\p<;�~��SU���G .�F�N}' �?U������d;V�f�-�r�0ҾzX���=S��\v���}^jCf�b�@ +�˷��� �#�%f},N ՝���� ��@���^\'����]�j��04�W��a�x��]� �VA�:Z��Lt� {��� ���Hk�,ZdhS*�0
$�U� 8=�|� ;��"�\���pb�י/�L~� �c�?̻�;_: `1	ِ9�� v��A��Q�Z�;�>仠�L���hp��!��z� ������&0�o-2�В�u�1a�����$�
���2�}�� ���K����1��,�	���QPr�0Y  �u���B�Q�������ʁ �	I$�� H cF*s2
 �B�%�K  �<��ʮ�� �S�N��y�� �P�B�� ZY���t0�9u��N��*� ���b!��c ^�4}�����P@`\�8�%�A�+�� �X�\Pp?�'�(��=�c�邢�W�� �J��9�>$v��~���|����@�
� &4��o .�qy���� �\�0�Ŋ �i�x]��>�$���}�J�-#�Z��s�2~�؁q\�/��Fd ���%�f �1���� ��У�p);��ið�{��6�)~����|bv� �1z�[#��]�  �����D�� �V,�S�� �&�ށ� s��,�J �	 ��Ժ�-��Ա!y$.(�� ��ņ�� ��X"V�' pz�P��6� C�
_B�[��D����s I�V);�wm ė�+� O�`�!�, ��X$˟�+� x����Tt8��5s��� �&�z_����]��`�S" �)QR=!�x� ݉3`Ioa ��+�7W� ��R1��,�� �:�a�d.�� �XR�_��W�w�;�-��3+|�pPj��!�z"ܭ� -�t��$\0щz�N�� bD�M�3�<N�@4������ K)\ ��dA���Pc�� ��b�� @��Z
X;�1 R��3�@d �	�}�҆=�PJ^�/й�-U�S,l�z B����� ��s*��eW ��@%�x/ ��p���� >��1�sG*S낀j�	"a<i��/m�� �{����p���[|� y4kdF�� �H�V�b��(�� ���W:m�| ���;Ų0 ��n���|� �G���H O����[���  �1� ��d���C<��im�;(
39H� Vd�rU ������{�(��G����� �	�݃b+� 24S�蘰(	��	�^ i�%�]�9 �O1��ĳ��	���po
 \+ߡ�� �����f��h@�D� ����"i�O� �@�b� ���!��9K� Q�3�/n 7��^�% ,�Ck�u�4g
��Ixi$�qW�Y��# ��GJ��� B��Xh��`�����G�P�%� ��Q3� Dr锨H�^h���*��N �A���i�4B��@H�| �lb:]��p� CW���X�� ,ٌ	���J���&Y���\y~�M>�z��d $���Q���� ^��y1vB8/r ��l�@�H�� �<���(�9��A��T�� ~�	
S�.L�� �L��$ �mk��G)\D	fƊ  ��T&�*��t4��ohL�g~l�� '! 㚙+���Z*��(� `���_���ē�$e�аP ʗ8�+.[vZ 	Ξwk3 j8��&��(��1�2�@?��4�����}�~��^���J�@5h'�y��
ۀf��R 	�o���Lkm �d�_��� ��+�] ��-_�f )�?�R�"� \��bP6����,aO�����ZӺ0��p՗������Q��ϋ2 �Z�t�:� �=҅RI�ZU�# �]y���0 Į�C�h�>J$�( |�ֻ�l ��Ѐ�/���w	� ���*� Z���ٚ0�gh#�1j����V��%��)(���`D� >�AH.vI� J��aG {�-P� �]�!��;V�a�~�o̑�S�� �Mt�(-� J	��XZ��u�����왣���K �<�҃��X��N��`a�>p�Y (�Qj*�q�}~~ ��5��/� ד�\���+�(��@?��1	�^�8/�o$��������k�] /YJ�Cm �ɡ[j,��.�����=�4�� ZS�I��C� ���H���� ��T��ː�.� OY���! ��_�����  �|Wz�� [��A�S��\~�$�@�o�= ����Uz	�$5��Yq��������J= �R@���)_�'����e� �`��[�sw 
\�A˼�W����u���Y=- h�H��n[ õ�2�Ʀ� �V�N*3~ ��`\1XQ ��&�����)�*���. �_\3�����[�Ҁ�-��8 �
���m� ��ݏ��L$1�	j� ��c�Y:��^9B 2phi�� ,�/�F^<�x����	�(>���3��vT_��a ���*�1�`Po�U �p��jx��'��`���R Q���D�F ~�
���U �25�l3�z yth\`½H� �i����P}�"�r�`/ QS��H� �I�f�[�� Vɮ� hMX0O7~� я3�u5?� �'�s�X� +�p(�G0� A���z� 
�a-�|�>������C�p-��I����m�$ ��(_���t��\z  -�J�#�� �p^��������Ī����La� $q�0�8 +H�:��h1 T,$<�u������Vx�zA� 
W+���� #�k-�6�� � y_���XU �!ш'�� [�o�<)�{ �?O�%�
=V����/��E�%w+����1���� ��D���� �'Zk0[� �Q튍 h*�?�m��!�Y���� � ZFh�l"O �B�k��*���4uC �R����h����z�� ��	��W �b�~�dn� @"
J˿���/�� c0�TX ��-��ݒs�  9�鑛��; $`�^i�/� �P��3V� 	���M�7 �^�"Ҫ� 0�W?Ĵa�;#�G	�*�� �V�E� �9�'��= 4��@��h O*�y�k ���3+� [*���� �P�$��� �&����	�b� �i�W����}`���e�����0p��Bs����(�y�;k
 �T�җ0��U�w� 6&]���(}%~�O�*m�5���M�I�0 �h�a˹� �	�\_�4 -��P�#{L $W(Կ��,�/` �"3��>�=��� .����ԝ��àG�ǨZ���XM�� ��H^�#a_)���`�	��� V�!���g� �\�р��� /��i�r4 ��_�lI�� ����W�� �q��1�I �,l6ߘ9V %�Ry�� 0����Җ� ��W�^�� f�FMI	��A��0 &K�ᢹ ��)�PC ��"�xD �� ��k8�#�x��`��z�P@�E"X(į�a�Y�SaM@�rB V�{��Ë���Z˰��� Hg��J�������"!�S)���_����� ���? ���g�B�: ��[�< KA���~� tL�|���nS��?�`�1*�Z(���
����� ���f���� MQ� g.A���;�D���2!�� �}fy� S���(�b� )����9��rc���3���' �d��]���!�P���)��W �1�m�+���FTN��hp&��B"ǀ]k��V �o��aQ�� v��η6�2 �+٬:�  \�0ڮD��1��=g��a(FV�{@�(䡀).�� Z�{�D'�R��������p5�������o
 ����͟*H������؅
s�Ƀ�+�h�R`K�I���w� 	K,�p���9��ö�ɬ����`��.� `�ͱ\'��|Z XS
���;	������e���E����HV����Sc  �A���Yc �/�W��X+ �Ѐ�	���Q ���(��1 䖀��|�:� QZ�V
A9� �O�w0��> !�+�ְ�� ���:��� ����
ZX� �Y�,x��� ���ػ���R�Y��%� p�����2 ��}�r?
x8ހ��S�̗@ p[�^�����v�(��wcp<�X��-+Q~�`�� m��Dېu�_�)� C���$ ?��^�! ��]��h �AE6�^ˁ �n��=��`: fQ �V8�2��"Y���-
 ����)��je`}u�\�1����A�t�$��NY=�} ?�̥1V�؀�'�Ǚ�~Qָ�� ��	����B�$`5�M� / �?����PRS躢1��WC�V�b#� �r�vL X�%p-��\�y �n.�� K�؃�W� xXU���VA�TkVۨ�0��vY�C���a�� ����SZ�1���� /j��� ���9�\ N�SٲJ� ��}�H	# @$��|��0rĠ��@3�R��J�������w�in$����p�a\��t�I rc%"��#� ,K��/� �Xdo	 ȇTe��~���V �� ������@>���� W +���gn?w�[ �S 3ճ���X �{�� �D�Z0��[ h�!��:� z��a��N,��	�e���� ���+� l�_/0� �����y *2�^��A �/$��c(�N���_֨�R�x��Թ]���>� �q
_8�U �~�FMxw�=�n� (��\3* ���*f�� ��}���� �^�! eQƶ�ɩ0J�N\�o�hO� 	��9��B Ď�-��� R��?fcQ3  ��﻿� �n����b� ��h m>�� P��7�2-�T�?���lX| �h�^Q�:�ڋ��R���
�^B�A�m��q���G�j��)�10�Y�b+��/�8�� �� ���B��AhD^m��H� ���\ ��.��K ^?B5Ce ՗�����ҵ�+�u \iK��` *����>l�	�� 
C�K˘� ��l_� �Nʏ{�� �L4/�Vv5L��U0� �Pݸyd �z���t ���Un�_Ӡ��� �;�'hil��u�1���? �7�no |Q�Wz  �-	�v�zI:��
�)�;ֆ:�4 \hRym l_�#���w�pC�[��>�0 ���KP�L ���MC�� Âc���n�[��� !����" ��^�v�{$���b����l������^�8�	��_��%\� �(A��"� �� ��_��R�	*@� B�ǐ����^CP��l�u? W�(�� �{���*���#���ȓv� �T���O��Id_���� �wq�	�� ���jGE��[ �(����v�=�� `Jŀ���y0_ ��Щ�Ns��u�`�#�	���ˀ��DG�	 �Pj��tR���@��Z�� X��!�b �
��Cj� �ʊ"�t�R:����|���:]� �V��S� �$xsj'_��YZ X�~
��ь�x� ��v�K�9�ڀB�� �D����}�v�3�|%b����(߀!�\ � hya@����$>�� �U�^�8��0��W� ,�6aI|��� �9�Ѽ� 1Ŀ5�� ����e���� �������ڃ5�)^!e�E��[X.M���-I �c�a��>	���19`.�'�����W����w��*��2 �&��B��� �)���< ��{�u�!��ì\~��͡ �mH�J/և #�{�|� �X&���	����[J���:��.��{ ��3�uE �`ƀ�%h�Y"��*�D`�� >0rY͆_���j����9��0 '����L��N f�qP� �%��S��� �U2�:�  xȉH�(>�X 
��wV QE�~���à�|O��J��AP{`�.��C�������?�DjV+ݨ������ `�	��M ����#P!� ��ν�ZGV 7�}
��� ���� �B 32�X���ty�v~ $��V�
 �����0����*?�Z&�>�Q)�O΂��� u �8���A���z��-��j� Z#轄&�X �V�`%1��̘` �h�JH��q ����
ˮ K���HJ �����0F =NZ��< �ֻQ	�,7������σf��!�>� _�ok���@l� �K�0*�%��3��c�k �F��ftX(rh ��R�U� ���#��� (ϤH�3Y W|?��ЄU ��X_�1� d��y$,��2�~ a0����; �F`&+�KC$������ϖ * P��Z��.�a�2��� ���Y��
 �ʸ�A� R ��C���� 8����a� {��-�<S� �O�/Й�W ��w�뮬 o5���Z�^[(! ��� w��]��@ ��-L�� ��dB����{ 1��8���P:�*>[�:��WA����!� ����̀h k���*�X��۽[��W= �_:�`� U�(%��9� ���<X� v��2�K�M WV���� ��/��&h �<~���,n>\�������x� ��*ۙ�#� ����W:� �kZ\ջ ��� �*(v��u  ��s���� �I`�Kx�� ��� ��߈�~ $���� j�̴�k�2 ^@�<&I فr��+� �zA��> �@��W�� ?�ǀ��2F�� 
���ڿ~a1�j��e���  >���<+�405��f�$�Q ��;!b��2 A	�=�,;�i �j��aK����B;3��w�N8 D�p@�	�"����ŷJ��電&�� p/b��o��Rn	�Z� ��}�� ~ ���Y�/	ʠP�H�A ��W
���#�Q-(@����_D��=� Y��Jn� �m�C�0���>�%�����|���]���-T�Bg�� ���@�1Z� �S�� ��*�5�bh9f>�j���z ���H_��}U��:*�6.�	��� z�a"�X 0�5�k���>�o��3�����}�=���h���¿"U�] �ʗs�V  �HX6�4�$�`�p_�y����:�//G DEt����b ���.�5 �{\R �Q@;I� MeB0�� �^�]��sO~�����} �i�u1~ h��n��+ ��Q
�� �!�#�h �V�ND<� ۃP
cݵx �K�F�%�� -3�t�`�X����������W ��R���@�^��2t����Y[\��/_���j�h&�ט����;���� ��� �^ ����va>�|������l�6 A����aB �n���@<# T��	X�̵v� ���[a�`�kS�����
�~� 4 G�5̠�KZ���J�� ����PY  �
�?b��*�N~�dG�{ �>��<�� ����xC�!��y��ua�E' �ǂ�t��� �ePfq�� ޼.�;�L2 a�� e�:>[Y�<�u��P�N��/��0�b����!�i�� G��ǰ�,� ȯ��\J ~�K��{������Қǽ�t��,��<�(�I�X� d�G���@�+C o��� 
O��D��r_2�J n� ���b{ވ� �Z��a��� J��!1Io�'�F�� �}� �+�9�"y~*�	��`u� T�Y}m � D����^� ���Oͪ �v��ү�JL!�G�+P()�@
�����8_J��QŹ$ b;xD��� �Y�í�� L���%e_ �ȟ@U�0��
E�=�� ���C�� ́	Ӡ�#��Ȭ�@ш �L����� �t�}lw� �B���V�8"��]������ �����[nܩ�_h�*k�ְ� G��L�,	�)����`���� �d�@_�ſ ��	���=H�=��Ah)'w F#^c��r�֍� �)��~SX0� ��OƼt��(����m*N `���� ZP層�� T]�#�)�U F�-����.J9�0�hO��T�n0 �Z��k1N���f�S�.��E�� ���,��� ���\e�u�9�Sm��K �
 �0Ě�Ԁ�������?D ���]� ���(N e �%?�� �6�~	ҭ�V)0�"|+] lU�����'����s| �4~K����;sy�Vp��@{�� 
���vH8&8��{.C������@g{��Y1X�U,��`��P(����ɗ�}�Q���� X��mV�q( �^�k��U�F$���4ur��� ����� �Q.�9נ�	1�Q]r`= ʴ��\Ȼ�U�y��a��������ڰ�� ����]�AX ��F�7�V �
������\p[ "��3��S U��[/���o-���2�� ��Ay�sv��(� ��	>��SX- q��pQ�� 2�!e:�J� N/W�q��f K�b]�	 �7�jOE �2���J�� )>.<�y��S%X�����.����h��[�	uO��b��� h\K+�|� fI�V���n R��"��z3  Z~OH��[ �A^I� ؽO�tZ�E�5np���
 �oB�vXa ��g4&�J� ����Y� ��Tz�x@u� ��t�JZ*� ���h�3L; 0ϴ��Tȸ( �����B2�q� Z
�@ �0w�	"}�g����X z�<�N�X� ���>B�&� ��/���=C�8���-}?੎��� ��/|I Ԟ<�,6�BEӸ� ��up9�f a��]x�N �k}�Q h�F�_/�I �D�鿴� JƲ	��V �21�5��X�:������*�$S����X� C�<4v  ��PF�a }f@��(���� -�SVe�¸ ��N5Ǔ� ���_!��	 �:��� �?^�G�R�`� ��{9'UwA�= �ݻ_�!.�� ���|h�I��0!	�u��R@��_� ��%����L- ��暵� �5������wz�y�!��� _0�>�
�^%� ���K�*4N �p� �Nf�-x,� ��c��J� _j��u i�`w����U$� X�f:��[� 8�BO��Ǽ�����"� ��*�ܐv<M�� ]Rd�ߒ9[��+�#&��|=���`��$ń�_ ���� ��J��T �%O~�A 	�.��)&� ���<�:����`^�C!� o���<#�d�D����N�$��M. �RT�	���� �#���}��%�A ��	��{'�\QG ���dc� �G�݁���,-@��#/���aP�������� �9���"&$�u�� �]���0� a�/�6tJ3 �B|�~dT� �h�N����P^�i��p�8P���\� )�X���D �A�4.�sYl��_k��&��	�������1#� �4�͐ t$P�c�� �8o"�	( �fZ!���;�ػ� ��$1��ؾ���Q��p�� j�R�E@� �+-�]�\� [�����0Y �tm���B�}��2 X�e�%�� "3۰�-=.h ���k8��1�z3�`� �V���9�� ��
2�	 �!ծ��U� �f��,T)��B�b4�ڒ���໅��pHS 1�F��� J�p�2�|��_����.Dv�	 I�)\�
�i�� l�J�� ��)�	��� ��՞�gxp��RU*���a�]0�ܮ'z�,��� nOcG4e �)�DS�ź ����4T ���";�~  m����H, �^����. �1n��?I�����B��a�&%<> �@O�\�&0>s�� ���2 ����0 kJf	B(zs���;�n`�pǫ ����� gA=]����� ?�v<XۂH����� S$�M�dP �cOIpy�H ��h��Kȹ 3q�8��E ��䤀/t�~�`��+� �	[����� )�B7���m�+ X�<+�,H����>��� 2��!���u [��|�h��V:�c��r� 䴈��5 "I�����R ���N#�	�jp�e6 �����/tXu  �n���Hi4 �?��+��2� wY�/@�)!�l�"�S`k�� >�UQ%�' ^}��$*�  ��FU�� �?	�uZB��.����0� ��c^Z�7� {ÀM[! ��ڡ�>�t �����_ ���?��J5 �!�i	q�Ax98�$��` ����| �I[��S w+����L !ɵ�h�� �5(g��i���4 �n��1�]������� � ��Tݎ�q�`�N;�V�tu�!��]1���8K����}�n���� �ܠa�q �]b ���F� ����-1g��(�;�= ��?�|Q0���~���/����}1�0��8�� � �PA8 �QN�4�� 	�1��U/� Q#�X� (�@��d�S `�-A߈�0 �b(�TZL�����2K �19�� *���{�	�h�b�d��^`ko 8���.��!�A�����/�*	�׀�C�ZN������龚 X-�삌� ��;��4, !'\��| �GX�o����
ky � <\��x �Y�0��`]>��B�q� E�N	�ښ, ���'Yy����f�5p�j�r��.����l�T]�t;>qf GL���	 � ��, �Ԗ��$& �:��2���<�� �UXYR� ��"�q_�v�� d� ��Z�u` �7�����=nt`X��)@ �2ih�p�F �3���Q� ���W��` ��S
ӗ� I���%��X����b��WQ �\��h%m p�xՓ�J� !:?�Ю#������Wd�P��� ����b��	 �r�$X14,^�~�Y3� �ʟі^U PH�]+� � *�� �F@}�V�O ��4PS]�B����@/ ^� ��6�N��e į?�
&F�� z\J�`�2rSW����4� �-�X��� �[��p�Q I,�����0~^ A�e� 	1���K�����s 	�����*� ��oX�2�K��� �fI� [���Q�U \�X�24r -��bTc�.y, ���鱟;�dx�s\�����; �����Y �Qd�?�h�[<� � ����.���hE�C�
J����	�?�ׄ���P�q�U�3o�D�쁱*�� "f`�N蜨�r+�[ЀS��_"�^ L�� G�I��vob�]U��=����O�� ��h&f3� �����6�=�����?7����� yN��! S���K r��H���L C�{.�m7����"�� K�*�¡]�WV���d���7 �Y����^�@��0 ��a��� �q�E�^- �W��D�������v�'�� �hix�� 9������� _O�SY�����Ѱ���0[a~�8>/�Hۨ�t� 2��b8�&�D�+�[��A�k�ֶ^����� 
s�EX��2L�L F����9PӀ�ـ��B� �q'A1�;� �z�Q� ��_�A�Ny� �Bik	�� ���1�Z� �W�D��� UlX��/�H)Z��I���o���`�a� �
��-Z 3nN"�R?�o��  ���� 
���D�WT�7._�%ඍ ���-�� ���\��	 ��X��~��� �պ�����v:G=�}�ro@����� ���]�w�o�����a �҆&�I61-V��3[ʉ� 0�Q��X]� }�y[h��� �N�Y(· s��~3�Q��ULX���Z�� d��� � |x@��c$ �����WA ��M�j��	Y��ʁ�?�����L.-;�*��|+���N=��p!����� ��c\
@` tv����P иY<��\)�
�yE�؀]p$1�_d�����9b� ��%�"(�� �d~Nڪ�� �[���	X 0��u~�cF���x �������8� _��V{ ����[r�����w�u@�6p;��Ӕ S*Ż� �� ؄��=2����`-��%�[W��Cp���3 ,u`)� ��q@�  �t4�mVzP Y�x��h-�s 4�T�2P�x�`I�)�Ğ&��U�0�� ��^2k��h �J �(�� ����¤� &3	��Y ���JZE$� ��r��`x
{� h ����Ѧ%f1��@� � L��w��� ��ETA���|�� k� ���'`&\&�ܪ]� ��i)�z�ȁb1������������ ��ktxPy$T2�[^����������& /��^�~��� ���jF�*���
���iW!`�=�K�y6�p��z�	��wXu����J ����|hy�� �|�!F >�9D/�p}<K5��7{`Oa��P�˳ �_)�1
�n�'& {� �l��b�J ���h�iߛ��P1ke�n+���('�XR���y)�:: ���V]QU��!���'heM E �3�\���7���1�V}�K �\"N�D%ڭP} �T�> ����� ZR饾�#�s>���_�9 Q�� �멘[�� 	�|���� �%!� �5�9�B},u+ ��]ڔ�nP1�� h�d������b��0l%�!��hG䌙@��W[qaQ?�8:���( F�~��m0�?�������l ����[��@ )կέ3 E�RUݽ:8V����~�&z����s��7 �/��tK� b���h��� �1�	N��# "��+b��dv-����;�. ac���~��@`�W�	�;H� ����A��t�FpC0��=fO���ţ���_��2@^����ʢ�ut�R2��� �W4�^�� *�c&z@�� �]���!�_P�[�pM�"5 Z�3O0(� S����_ %���U����/ �0` ����s.�	���| {P�Y%��Aq � ���w�t -�p���\ h�+@��~ J�S�E# ��*ً ���
�>�̐  �����y��Z�tm
r��6�Q ��.Y�����ĺ��B���D.	�H �S��h 3 �����6L����d �bo/Q;ԫ�YBK���� Z���pT�� `�Y�͙� b1�P�	� J��lh�� [����vf-	��@2,ڂ� �@{/���^oT0��ȸB ���¯�� �����-�?簙�^0��|�ʬ�[��n��+�1����̘6�  �����7Q�!d����b��H�X�lr�� �d��J� �Q��[�+s�� �BN�� }��9��#�&�[���00��� 1��V(_�;i� ��7^"&� ����j �T_�����! ��:�%ǂ ��]n"�X!	���Wp��>� D��.HSz ��%Ru V�>��K�h��+���5�~�m���{$(� {�mV�HF� ��J� ����U�N_@��9� �SڬUp�^
� �A��z �'-���u�|j�� ��"kC��! �`�+��| Ȁ6X� j�����VZ��@I-��	hjp�����
ԉ������V���+O �'(�^	a\�U5k�%����fh V��gZ0�2 �l�>���G�M��# ������L5�� ���:= [՘A�ԶW`�U@ը�� ��%gw�� 5�"����Q���,���>����,���/�s�pOh� '*D��ρh `;/I�.R?(���@)�p�JZ�c� _�����&�& �0ф߾ aW>��%� �[��Z!��~@��`Uቕ��O�>(ˀ^�*K>�� �h��� Toj�R �#�_�y �|%��V��=G q_�Ļ� W���B5��g0��Ј��. �#�R��� I��ZT��ː��^ +΁���?� 2�3H[�6�jԷF��!� \0���ŝ� N,RP�d��1��@����EԦK�G%�h� θ��V~� /�1��� �BZ��Yc ��8bS	.�Ai�� ����� +B.'��������4P��3�" ��B�q���AG���[��>�@��E�0b`��%��a��¶.�  �<.��������%f� �H�N<�]����� ���ߟ���Js ����	�h
!�)-�L�� N�[��Dǔph�c��V
�P�r������t!�(/�H�s40)�Q`c��= �sKɒ�@� ZM���Q8�B(@�^I[w �&����) �-��r/�� ӹ��  M'��$5=��:������!Ka^׸Ey� �e��	ց �X�Z
� C���h�	V ��p3�;�� K� CS�����Ӹ<L؈�LA� �)�*�̩�� E��Ҩ=IJ1���]��� �ҏ:X� ��r�R
� ��#U��Z�� A(4�,9ʓ 	�dUD�x{ �
|bk!�(wh�
1�qg� PU��|k �vdA���? ـ2�Q
��"iW��Y��Z1 /�5�N�?�&�X3 2��@t �P��0x�X�a ���bV i�]�٘� w�^���t.K� ĺg��>���`������ 2�BS��Rn\	��y7 (�0w ��t �Qsʷ�o���3B�V~� K��R��+	 �Z�6�}^>��L�:�ˑP�	8�E�Ӭ Ť�HR��GK�_�l��� ����=ܿ �Y���l8[Q ޱ+�0 � ��5��X�C���P��	���{��+�g1� ����� ��Ov��\&R 3H��-�K~���z��P�aL@ 8�����_d�q��
PW �&���_	靅��zP<}CL]|<�7�V� �0��^P�a g)DC�X�������!�_T a�Y5%�� ���MN� ���0�V? I��A�� xQ :%r���(�?� c�X�sZ n')�[�� ���3X�<5,�	��`x� ����˪ Ț(��6^ h�]� �O ��#�GB3 �)�N0(Lwa���[��j@/͒J ���Z"�!���>G 6�ڼL�[
 �p��F�d��C�������/ ��ԉBŐ� �p�
��`0 "�d� Yn� si�w:ʇ�K����?� �	���jq �wr�� ��"_�� �3��7�Y��!� 1�/�l
Z#	 3�\��9� ��,� A�0�X��jBx���y�`p� Pq�I,� 髯K�Fp? �����a	�@�b
 �E ��D�)��� F�r��վ ��H��� R_3 ��&~!&G� 	1�_�s �/�W���� ��#��� T�~G�5 +Vδ.S�	r����ժ �El�V1�^�	���C i� �_�O}1u���� ���ȋ ��\^�� 	O�ܐ����� �Jc�=W%"��|�X�� �4���O� j����0&\�� e�-U�� ����`��{ �T�HZ��Qx����Y�L�qz� �-� ��@H��s��'��u�8]h��`#--0v Hs6F7 u@��~� �P�)�Z�� %�^#�U*�~�����90�P���h9 *X��^�h������z'dJ \L�(�^��?.� ����L�a�� ��w���5>o� >|�� ��X���ֺs���6$1� yc��I �h��oe�~:�#�O��J�� ���Z� �`��0�WA:*�0�@ך� R�x�8�� ���Ź�� @%1!�,Z��fN.��O�
�I��-���� �ȣ��	����w2.�<�}-��)o�EfF�6��uLv �"�_�: �5�;� ��ú�& ����k �jcۀz������)���
�:�@`�C�r 3�H�J�ô�쮐�(r ��|��EȻ  ��^Y�D �����b�nHt��`S�>�� ������� $-�4�9P��hHWO�O H��b�I���DѾ� *uh8>b^����� C��x0J� �;����2�U B	��v�6 �*�f�g�"�!�
`	[}tQ �z�*ؿ	 ��ߋ�T �ZiV+P�0��E3r0H� [�y�]�z��-�@���) �N�
�(���=���^��J�$ ���
�Z)t��d�=QT����r'�wĂ�ta ~�+�&�M �s"�)$#�� 0����(| ����+b Y ����G`:�P-��� R$��c�[ �&�<Q/���eٰ��n)� I��һ���lMV�W/��_`K�� ����MKH� +��2��� ���Ro�'_���A��q%�� ��݂�̇ FE�M�B 1���W��{~ ���@�_� �k��{/x Y:m��������� u�%V)Օ W6�\"xO� �f`RlJ�� D�ST�̞�$�%	� m�� ��@mZ(� ����Q� �Ѕ��	�� ޏ-~`�;m|�d\�#��hKT� �'�}e����V�f~�B�� [�	/E��� �,ZYA�� ��k&�� է�L!� Vj���� �Q�:�F� 9/��X � B1�Z�"~k O�ɲ��y $��򅘼��`Pp�?�,�>�i��u���� K4�Ym, ?0�1���� �kR�	� ���fbhs}���5��� -��$�]� _����A��  �.��9� �X��-�RQ 
���Ɛ� �P%��_p�� '� 0�[�J	������WtKD � ��1���#c>�H= %>��O���]`�\ �z�40h K ʴ5W���\`��q��t  H8T[1o _<��� ��A@�+:�`��Z \��R�
P!ؘ� �� �����氷�r��@�h�����V�Ho:{�yE���� f1�)�Z ρ�yF�S ���z�<�[��5ޠ��%�8k��Љ]�  ���S�� ��%��:�ߴ +�0(����N��  �9b&� MY��� o��	��| ����T��Hh;  �)��� �!ʺ�� 6��Qh� '+&=�[ۯ r��]��ܸ ����d�	��s �5��' W.�N�`x�(#@����d��Vup�|�!�A\��_k	�wc=R��(n�upЕ� Q���B~ 4�Ѵ�&'�,��8 R1�YOZprf ��;�B$����`5�U��>���[���|$�� @
)ص ��5~��Y\a�v{����-���!x��,�N�@V t� ��L�BX�� ���� p(F�C�� �{O��Bt9�=�[3�0g0�5 +X����y`W|�@E9�u�=h3@�&ܷ>k��u�����vr��ːp2��`�w��k�͛�Xl2����E:��!��.�l �/Q��\, c�V_x��O������ɮW��hQx�1�	�c*��t�0� �P��Ⱥ� ����������4 �-�8,0щ 7�;�	 �h�GP�]�\	`'�[�HA�_^���+�!E�Q0���fP�1�2�" j��`K�	_���m05�� �z���	� �VX2�<  �uh�� N}��"׮�X�P� b�h�+��(J�P�]y���-��t��%���H��#�S}� �����*��z���� �\Z F:J�=�j�[ ]h�ӵ T1� ��	��Xbb��@��v~�px `|��,K P���Cc� w�p2G|�) �B
��@�O����Bn�S��[�:�% ��PT ��?�|�#��`V&~B �����l��MU���7���0/Y޳�[W� ]b x������� U҂�F��:@aN1�~� �Ž\��/:�|���h�25 �Io�	<�K ��Be4Q �
@Υb�L�\���� ��+4��#��M�B��Lr �G��� �+ D�ꑇc1�=����ȷ~�A�x �ɦX(�Q�� ��e�Yv� |3�5��U��R�@`Q��;���1Q&!��R��N �����3�5f�����*	�����p�[^��� /��R;� �XVy��N?�� -��@������o�^��(�/ ��5�+�K� ���\��d����U ��8�P �E�\|O�}.�Ң'�\ ⢷]x�(� Ѹ?!���I �<���/�
�Լ S(ј�P ��N�b1 �\��y[&�tv q�{�G���K1_M'<x`CT[��;=��*�\� un����| s#!��g� _eo8a�O�< �%zTPX� �Q+���8$#�� �OH�Ώ��hc>�� :��?	��J�%Ǌ`R�4� j�Wh�ftA 3���1�� �Gq&*�� �8�p�,�
�A �V�o�9�!��N*�m�.:���Р�rū^0�ݭ���l�O�~@y����.N W�l�U�/ ���
�� �@����(�$��m��R���QΏ�A2�W���� ��:�aD� �o7�b��Mz�� )	��� 	\�R {�c� �,�
Y� �Wע@7(X�� t0�P�8�&� �jN%� ].d��f= X�� � 7l���T_ '��}3� �5���f1� ���ֲ�C �%:hdʅ�� S+��oB�X �fX�&��5������]�Q�,*�H�(��[�Ӿptv	 ��E�&�z -�^�b$�|� � �h* Ĳ�QW� ����Y�s!��
LV�к� ��,�X�)z� -[��r���Hd� �+2�"9�� �!��:� �Z&���� hi��I �u�ܮbK|]B"`��yk�,#� �bE	͹ O=���/N������q ���k8i� �5R`c#t��"�I��7E\ 9b�.2� ���,<� YA���Q�u�a|� V�L+� Y�Е}v���x@������C���Ǡ$�� ),�:^�F���_�؀�<�֟/}���VZ@,�(p^�a��� �[X���� �*ܕ�i��LRU �\a�:r� 1!���r����,p�` ����T��W����s����؀ ���T q�n�Ӑ�/xX �tK�W���� Z�ڇ�C� ��_���Dq� �<!�������9n�p xS2�W#� �)*�y�� ,�7q+�1�" e��?<-@w ��'�]f� ��Y��8*�&�F����i�:����`����d��� ��Bmh� +�ꦛ��4� �ǽ1��]K �(t$��-p���A��=�VF
�q�-�	t�gU#�������@a��1XN�q�G9ʤ?� ��3�1�a�5J�[�A�����o0�)��8���P2�6;Ha*m������:S���v#O`dR
�� O4A��H�[�@v�W���.�6�!k�sU���� C�z��	�$�9� E��r{[ ��\�a v� �����_�S� 'X�h�y���H��!���ɠ��{$ �)�#�Z�� g�͖. bN��n	S
�P��3�� �Yu��; �pD؊
 ��rAZY�c Q�Jv�'R��/1�"w_̎� Ƹ��[)�� �d�\�W����X�p_�P U��z��c� �	�C���A Ø{ڼB
 ����^}yX��&���L�H�A(��%���D� )�[1� ƸN ԗ^ӥ���#|Wп�E} �+���H4 Q��!;2�C���/��������^1��=(Z��! ����&��@/V� �.D�� #=��]�^4��|!�u��-�~� �R�g �ǧ�95V i�
hf���Kλ ��1r�t!�ڀ��C��< z�{.�!� D�0U��&[R� �]?�8w� &3�_�J f)���V^9I �A��0� �Z��F }" |��[+��!�9�� nR�.u�� ���P�6�*���� �"��&$5 9R��|� �/�uv, 0�?�8� ��H&!��}���� <P"׸^��Ot'@ }� �m������ �%�l�� �����v!	#q�n�`���_ ��iaO�� ��v�&� �%� �Q� 룳��Xh�x]	�zY��� y/�2�$9��kKЃ
ǻKg�� >���=�� OY��h5H&� ����� f|0�%�]�~�q+ _��#(��$ D��Z�@��̷Bjv�����U5� xg�T	��G��`s �."� ���P�0�^ �U17V��� ;�}E	�ʗ ����@ �)�#��K� �8W���� I�����Ŷ���83�' �����֗�Y���H�Z��	���q� ���Ie	�-ɀZп����r^���B�D��`�'�x ?�O���|��wr� ���䂇{ ���j0ɔM `��F���LK� �YI\Sxy 鲎1��� 	3L@&�6�R�,υ��Pж �yg [m%=� וЁX�T &��ELU ȴ�0]�Q��S:�	��	?��?��ߓ h��Z!�ҵ �ق-��� ,�L '�I^NM� a�P|�� �[�p�h� �o�a!ӻv '���.O�� ������,� 	������*��󍞤)�n� Y���1� ����h������K*�@��gb� iA��u{:	2}��9>�� ��m�Zӏ�v��	h0-�} �$��Ɓ*����j����= ��]b*}�� �� �['!�y��# 5U����0cu~�P�!ͺ )����9 p�J<�, �񀲉�� F��k���H��;���\.�=��_B�0"��i�L��(��~2SG�U�o�)�� ��`&:H�� 	!�+kp��R(�N�8�F�:�/@�Tgx?X,%S���8��"ˁ� ���к4������g�� 0�}��* ��s�����@[�^��j�� �h�MvTb�J������ Ai[?^�Z ��&�0$-ߝ��q�!��� *�F�i)
� (>X�.�_{�L񴀚Q��O I����x ����7�A�t /��Z��'����P��-� Q1ݯ� ,;�% �\m-E� ���Ѥ�7 SW�VB� _����c���R�Kx�� ���]"��sG (��ja z:��^!� A�[1`S�������H���V2�;�J��@	�1x�6 '�j�ZRŞ���� ����3
 􀈸u_�� "J�S��y����v�P��Q0Ӽ��/b������Z�x4�њ ���C� ��	�^�� ��W��([�L-���� /�f'3 �V����<��2�wȠh�ps=|����
���-U���+�� ��?��� �t�m	3 ���%I�Vta 2��@�� )_��Pd ����@Yz�b,�U�X]���-^0W�y��E��[ b���� �~uN7K���c�������� !؀��[^ �X>K�տ 	W�{R� z�Z��:�H�����S� ����dE� QΖA�� y@��2�x �`s�z�l) �Jk�t ��]-�s}� W�45�@������Il��� �?V��%�� �6����� ��dz��� g@�Q� F6��Z�� ��{!��� �$��S�N] 'ֈ�D�3��Lw.5� �-�v@  �����H���B�A(О�%�R}�f|��� ���DXKJ��� ҽ���1 �ȇ���K�;��$l�	A~	� h�9Y ������ ky� ���,C��
#���B���Z�(���� �2O[��Y�.*`� E���ڟ	 c �gɧ� /���,O9�,6] z���� �p�[�-_x���h���K�� ��ވ�P�y ���A�j�@ ���[�c %)J���� H�Z�O-7i�
�5��H���T�� ��(�ڎ����o�>��-0gU���C4u�K����2��[X!������ �� ��ٳ/�F ����K ���:I�n�!��L��� b���J7W ��@�\P�����$�=i�F�H����| 1��p�� 5#?�Q ��>� �Sh �Ыu�|K� ��/�� �vN6�h\g ���A�BY �i�*����M�UDE����G ŝYnB��.[� ��D�# �1�?�+C�|	hk w$��%dD 
�9�˨e V魇�8n��i���� �h�� �o��@:� �R選X+� .�ؙ)�� �<����X 0ڪ�#/W �V>�m���  ���jq�x#�Y���|��� ���[��g ������ u���8�. !�ӫ�r' ]��нh\1 m�J�Hb~� /4��\!L��>��}[���s^��� n���#���@-%"��� ��WH 2� O����J@����F��f�\
Z��q� i*�A!|�����'��?OY*20�  !��H���p�(�* b�_�ʱҿX� ��N9�I]V�P�頽�'�0�  ��&
r� ���^oV�� ��(��~ G�b���1 ��Z��� r �W��� %L�q�_O ��,�Ӗ���� �f[�i���o��c�-�� ��"�n�V�p�%|4��I@́�K8��h���X �^�߸���a���\�x,o ��,Z*�0���eG�`�� �h{�z��� wI�x�@b<0� R��
��� !��kB��u ���4� J ���|@ڻ�y�~�a�1��� (�E�u���癵x�� �� ��%��`����:Hlt�Y(����`�]��܄ ؚ�V� �	��L` �(�fP�? ���UpSJ� ��OAr�?����Pi��f�bH�� XT�)�\8 h��P� ���!m�  �7��@�"A�S��@��l��  6�C+� �(7����?�_>Q� A[0-��Y�c *���:	� F@و�["�Z� <!�% ;�L�YX�=���x�.� ���^��3��X����(��M��2B�c ��]�!f @,��h`m �e	��K��Q ��R������ ��`��, ���I;>!� y��1�'S A&:�V� � �����	�`�� �'X�\�9 ���Eo���|��Z��C��Q�����%�T?X�	vm3�W@�ȥ�� K쨆�	�P�\v� R��d����,ʜs0�� 82� �Z��"�WwdiM���`	>���V���"$�- ]z��O�@�{T ����(� )��U�$�>{�!����� �����4�
'^�� Ugℝ ��!��I��ipp�b �K����Uǐ�t3��b�*� ��'��? �{�NX�� �R�^e��A�н�8*�Y�݊#�H �(e�h�v�� �OèS�э0���`����ݏ� }��9������I�_�4�?k�� �����a �3XxR	 Y!�v��� �o51��� �¢�?>(�؀��=1��I�T )�6p{����`����	�J����U�� '(؁�R& �A^�t J���x�> h&p�^�X� +K��a��O�) *��'Vrf �"�$#�c��V���Q �j�F��=����ih�Vd� 2����C�B �{O+Áu Z��q���f��-���D�΁��@kAs ���K��h�B��=[.�����A����p������T�B	{�2Ƞ��) �ܗ����L�":
����[�� "f�u�`-�1���6X3�� 5��m* q���R���dy<���&�l\@ W��e�K� q��L �J�B�$�-?Z���yi�	ɸ�t:}S�a�*����� �=�ˇ�\� y|��ʣ� ȋ'����}���ʲ���jp<�, ��C8�����A�� 崾�e��E�`N���x��#m�� ��`w.��� ([U��&n�� �����	�*�;��� ���D�K5�`L����':� o��`4�T�[z�rK0�� ���hQ*� ��4��x�:��w �\M^���� V�K"��� �	�̉/]��ǈJ����1Td� #�Ӹ% D*�3��W��-��P{� 1r�&�S$a���W���_3��D����p�(c�
�� ��,^g�����3\0\�Rp"������ G ��z�=RO$�J���Z�� Y�d�[_(� �*s��!�P����h-5:w��b�1�� Zq�u�ٖ�/��c�2��ȼ7 'I��? � �k2�,.{��� �i�J�  �`SV��I �\^F�&��"f�� v˴� ��4��T�� �vY0�S �8h���9 ��־��� L�!��G �i3kT <'�d� �"-7�|lB� }�	Zh� �����N�ۘ�]�	������wo ��ҝh'�.(S��� ���*��p! �J�R��<���X���.�Ћ,�uD ��%X@] Uh.�V�Ā�� k&����(
 	�΂Z�� �)h�� �C�E�"������ň&q_- �g�(��w�l e�v�U��!�"\� q��ɷ���>8� �v5�T�  ��j���! U�a���� g0:ۅ �� �7H{L<�Z�%X���#ɔ���& A��E��sP��� ����N��%� ���J��
������@�?oǽ��HP
 (ܸ�) �o"��� h%1~��E +��P���0u�fRS�|�t�K��� %�B����҇p
� 8�;��' ��A�Yu��Sm1�0�; .D$����X 	̔���)� N��ȧ� �Q	��!j��� qDI���� �r�]#��Hx �SG	�v�NY i����� ,�[��0@s1� �f�;�� Ѱ�jh	
��Jb����҈ �\�j�� �����	J ���?��
 *�@��2�$]�+�V� y�J��i}Ch���  �����EJ����)�u�<`�H_gLks� f���D! �Y�{er� ��.#��8�4����h*JIP˙(�Bn7�d������`){ �#� �_� 0��V��� 5��Yh&���'�0�6� ����\���~��S���'CG��&�)CA�BU���+	J�ΏQ���p�2�|�;�0�$F �fh:�>D��0����" �(�`�.�� ȝ}��{�l�`��± �q����5�` "I�~v��m����a4_ f-���Q`��Z�H֍f@Ο`	�� ��!톘1
X}��~󊠒Y� ���J�.<�� jý��;z� ⃖��O4� ����/Z�R ��\���X� ��� G�- g.B�����\���!2)�pLV��K�bk�f,��L :�����! 9�U��< ��g8-�|%���#0��=rE���Wx4m !��.I Q������zb� ��U���M�G ��-�Np��e&� ��Gu�� R�� >�,3�.`����W ����!�C ;��O5���2���ep\�������a�-��
~� �'!��b)�� m������ ����ZWP ��؈�(� ��D߉��8[!u�A ��I�� Ι]:��� -h�J��s� K��F
oD ^3�-�nt�?rҀx�'�ky� п̃�(� �3�*ZS� �\/ V�}[��y�<d�� �'B�]�G���c΀���_��� �V��B� �Ǹ�-~ ��ȭ a�Q�r�6<A	�ڎ���"���)��/�� v� ��É����V ���
�$ ���t� �}�	��!�B�\ e��? f7�v|�r �����Q~ 	*�����<�?��`��2����7�Qu�̥' eH�Y0��}& �� о'R��Lt�&3�� �T9�U@ �Z�w�q ��G+�k�\� ahK<�s�QB�+��9A�Z�r�W	���C�}�=,�"��?����� �W���ɷt i:3��o�� �]^H2�[ ������ �#�:`���a�L{^o��V'J(@p$#�<�!�@yb
 �/��h` �7��'�4� �Z_Q(��� ��@1�y �i>? 7�HC(ܶ�k��Z��DP�|��1�b���� ��՚�X l%�(�� �1��d� ����K�H� �%2�@��PT�(,٭6��&��8"�@�fY�� {
�r|��H ���.�B&D RN�_	w� ��u��rE�2	6�{\�@���� �7=gb��<[ _װ3�i�翀�lL\ �{������~�vE��d���V���Z  �^���I�>��@UbXH�.��� ��Sq� ʰ�@9� Z���#8�I~=�V
�K�`Appa"�H�%Q��	��D����Z {_�6�%� 9>�« O�k�ʴ
D��W�x����S�_�@J� �X�.�x��������>/� ��e�
$ ֔'Wg@������k����7; � R\S WJ�fj_F� 	����'� ����-�| �:RV0��w�����f;i'��>2&����L� P��� �������R�� Ⱥw�e>�;J��D�"�a- �y@�S���<��o�� ��6>��¸� w�?t�! f���(�PY �󠉎¿�z|��2� p6�%( ��Q�{+�->�%����NB��j UiL��%�~�E������ �� ��� �́�>Ojɼ5 �S�^�x	�wq�@� ��ޜ\T�,��D ��0�^E�yU��I! ý'���;1�X�@��U��[ &��س��% �k0��S(�.V[ ����a:��3�Z�|09ӈ�0�����Ta�ڝ��M W��	��� ��Lנ�I�/���b�`8��jY9*��	��"u�&]�"�����:\Hw( ��2W)ZPD	���݅���yۄ ���q�1 j�z�'^�L{�	� y��J Z��>��.@ ���(e�
��h�0�� :S�,� O3�Q0b �(����E���`�RP�&�1 �W�o��n����������T�����<a�� Q�b"�SZ�,N��Hѣ��������5�ؿ���*���\a��H 7���)Fz�[XO/�9ypb�աL�`PE �|��1� p%�q~�Y� ۼ��m�r: �- K��5�
�@- P]Q��B E �/�x��0 -m�}3Z�qǋ>��#_�������8G��0� &ZR�n
 ,����z%	ɔ��� ��\Z^ Đ��DL& 勥�磧| A�e�/=�}�	� ��8<
	��Y���9�[ ��e��U��H߹MS��5"�0.����v%�>U`�z ��B}���lٿ���:ځ�4�Z��(������/�� �L(�x 1�X3ˁ-�<����)�2� ��eq{/�R��H� �ƾ��� �AҀd;� �SU��W�M ,3"�10� ��QzZÁS ɋ�}�F�4���O������cx)�@v��ź � e�>B�� �@�����W��� 1�� f��w�Y�x\0^�߲;H�_�� (�h�G��M ���aF� Q��[kV �f)�xY &���0�h �Њ��T�  ռ��a k��#�Zr [���}� *�8I@��`��%ӷT ��̃<� �*�	@�� ��0q+�W-���_�ۇ �t���j�� ��3N�/�I	��V|�a�,�:�v�sf��tP'�iF�@���=���I�W^��� ��p2��&1t� =d�A���;؜ ���/v� Ƀ:�d( с��N.�� ��1|��5$4 ��ݽ�� �h��8��`��[G��+��Ah�� 9I?X���� `���Y(��{���~�/�& l�'V_B*�W���z�G��P���k�<��h ���%��� �@�]+b�T 3����;h��� b�&	��: �j��L�� �!�z��1{� �?�_� ���?เ䝁��M �(��)"�wB �̿�N;܁�T���)w������s$�x[V� ��h&�6^FCd�	�H�����qB����9΀�?�Tf� �`���$У� �8s�p� ��t-�����g	 G���f5 �����eM� �V�{��?� 0�GY�<���8� ��h�I]����- -����� _W�`e9� S���QP�]H��(aoDep,=�> x-���� 	�jH?.�zgX-����* �)K��9<_��Y��s, �y��n:��wU4�6@�<wI ��	$?A�j %o�wJ�tV��}6��M��~��*�^@Q�.� 杗E�B��&� 㤃q���,��_�� ���	�� �/�3��z� �|�2��	ǮЁ ,��: Yv!���"atq����l�d�\+2�	���͙��t��9��S#��[N j�s�X )���d�L�쮉�h�-�� ��f	'�P~	�/\U��;Մ� ��뼶}Z8�� i��j�'�"���G�����%&�oQ��ր� �`�_*�3 �;��� ��k�LZd�K��h@�/��� .%]��� ��D�W`5huJ3���/�~ܓB�� �hP�͗1�c鈮��`X �dS%T[F���Kfh����� aZt*�1�
��و��4� 鋵+�� ����Z��'`U�lk!���)��J�b���=� �]��a9T�V��L��c'��@�����1�^: �3+[/�L F�C鐓I� �_����L�} �>�T1�K�����`�d��� o�X��N�%��[# ��c��,�� �B��Yj @8��gR ��į�����W�	�(������X�K%�ٺ�U��� Y0B�ӗ��tOهK��Ä35��b@'�!I �,�U �^E4<�	�Q?�� 1k���.�p� R�P�{� ���d�]�#�@�c
� ֒k3�V ���E�.����� �3D��Ft��� i��uи� �JYf�8� �Q Ϲ��8 
dL���"� PI�@��% 0�U5߹�ïv���}& <ν�U+�pY;� �����  ��-�UZ� E+� �~�� �WvH� T3�EQ(� ��b��0�������H	� r� �V�(��P���� \s��QV �m� �� �s��n���So�L� �Ө䆖� |��_�f ���GQ0�:�(@Z������
���r�S���3�� ��P1
Z�U�? !��u^�q�L��ĄJ��ˀ=�R�n� �H����� ?���x ��N�bĝ q~A�� � *�f[(� G)�Ca�P<�/�\~�$!ز�fڡ��T���J��	M� w�\fZ�u� 4��9�a6��N���!V3�*���Lt��h�SU_���P H�($Ϳ�@ �� )\�_/ !���;��� �%w�� +�q!Lc~ ���RU� ���]�� ���1��,O@I ٚ}(� �[Sk�9�� �:�!/�X�Q��W���S�#�a`J�,J���/�� 綝�1|�0�E�^���2Th� �dM;f@������) � 3����A���h^�%��".�� �!�;� ��Z��%~D�����l� �R��)� �V��%�̖ ��4y,�sp �h��i�lX�; ��5fު"�0	�2�z��ۖ� p���/h� 	���H ��=5,��~M8�8 ����fX  ʡ��2�$O�X� �=�~/n ��!�0a1��S{ �H��_� �7M�U� X��/��ظ7 �hNA�(�� 'IԁM�H�y� ��[��ީ�� ��(�%�}Q���2�^�x�� ��V�S\�`E@"��%��Ԧ���9D1>�C,	���'���:���#�X g{$@.������ � ]`���2�U
#�BV�P]��~�C��1���4'm	�� {Z�}@��h �gj���G #��0Pk�+ ����r� *H�%��/� sb0^��o��8�*��	����+A�Ճ�F`���%]2 |H>���m $��58��x́��@��	>�y ɧ��E� &s���d2LQ��b��1 ȹ�>�[( �V�	�l�� <���_q�� �LI��p��f���p�Y�h�`�L�� ��~�K\�9��(� ��y��1�Z 鲅�.PK D|��vk�= |XY��u��>Nv�  ��~Q ����~� xn*!��<� eQݨ֕�2 �q�EA�0�`����n�^�� ��=����}�R����p �)�[hvpF�V���Đ� 1�XP)�����DЋ����	���n�)0�`�~� �
v�PZ�wS'��N��փ�]\��av���Q�S Yo��ab� Mk��@�н ����5��iL�t $Q#��, �jZqG@ (�\�0���L1�Jp76a�yk#	�p���q�8�f�	���{����[C@ �ܶ0$�r$�� � �����E��d �<�[���h0_�l����ŗ� ���u}N�fe$(��08�=�W8̼B I��� ��_W�2A ��"`hP�5�L��O� �1�0'�Xr�ԣ� �9������8Bt�~����Pи��
���u�< *�� ����&� �J������ Y3[��X� ���9����z�`��Q� ѷ��� ~��L�-�� �a
���� �3�u�=������ ���� �$=���6}���+� U�|f/� �"�I� �'�*r�  l��(�c ަ#�8	�MV���ϯ���!���� ���I�ԠR� ~_2�Lh�x�� �0z�5�P����Oغ ��j�qQ/��|��������t�iw����)��.ό=�9��\��
�� ^�=�Mx� ������ � ���BY� &H����S 9���1�0�n�c`$ޕ 	_p|�i؈-1������ ����[��h���&� ދ�<)[�UV�	���!Çg� ��̀$�8o.�8�7VvZ1�_���g�~} ����ȲRsC�v�%(���"�Z��J��:4?_���U%�����ـ����� �0��P<t� ����K� ���*�/ Z�����ƀHhs�����& _���� !꾂���2�]7��@��Wq�wA'����4��$��L� j�:K��Pl�� m^��!� Z���;W���u ���Ղ,؄{� �DX�Ā&2 �h'P�s�&3ɇF]D�,�p	���E�o ��[��7��ʿ����k &��� �0Ѭ�@ :����2U��c������hw.yU�
H�	䋀�ɯV� q)�`� .��-�� _�B#���H�&��@�>}`Yx��t~/ �b?L�	QS #��YU��s�����y �nY��QR 2�K�ݢ,� �]^6�)�� �_X�A�L��%�t���Ϥz ��h��T� �jL�K�� ����$U6 ��z���!ڡ�pX�ۯ�`�@ ERK���Gf��U��:��i �� ��� J[������ t���ܫʶ H�%A�Q�@�! �h$�?���p �ӹ>b=A3(�P� 1d��$h� �����"���	���-� �[
֟Y�Q 7@��\��H2I���� ��B�����ã� �����k����<`SW �v�D��� �u���,?]u��s�E% �̥b� ��S/Rd����]'{��V����S $��[�	��=I����o�M,}�� ��1Ң Ǯ����f���{�O��� =T��@�X�>��cܓ��_{��^ 1M$C�� �u/�+\7�3?e��`�Ѫ �@�긥' c�u��ٗ���%��b �!�	~"�+�@F�5��20 m�>�� �'E�[� TJ���h.uq
��`� ���[}� �۠�hXB'��8 P���t�� 8u�N�h�� a�I;�`��QU1���.Չ >_y��������q#�'_/\��*�� [��W�� K��c�! ��4�Z�d����u��ti ()ʀ��&� �Lvh/Pw���z�ǻ���� _��#� O�� BF�]� ��閤�+�ׄ ��Dy� �n��PR�� A8k��`:# &�Y��FE �L޲|/h"	D{�U�\��3�-� +K`�VTx1[��v ��̝�R��L�����8@� 3[W�J>���0�,a�`� \���J��?�H��s]�L ĕ�����Ǧ� ^˫]�) �;�h���3}��� �V�1طy�a�kq�� (@*W_pYt� 0�Q
/�P� �"��V3���ѿ�{��DZX$2�|��x���EW0a�j� �r�`�� 5HY7���� _V4����=�:I S�� RPg"�| ���_�D��x�jl ahCR���{7�U� ��y�<0؇�ė{ ��~�6��e_͸�: t����W Z��7��R������M��2� �,��b�*t�S:ʾ�2(��=����#���������h��! :���<F5��� �U����P k�Q��q�>�R [pi�+,�� �^��<��_:�	r� ��1�3�� '��0?#���K5^��9Z`�0�� ���â[^+�0<%@��G�U���9�Qx� h�Rn�^d� �Ȉ�S� ��D��C����YZ�{'/X���+�P��K|8�����L�'� �	���J�� So%Ʋ��i�@��|������(Z�[�a_c���ή�v� {�~3�ni �Zj��*�W�A��U�8��k�~�1�dܠ_���	I�?
 x�K���Y8U+����~M��!%�� ���KV�</�1�00^$��઀�� sp�¢�}Tv�:"ą������B (0%\L� u��+��_�M %��eh��v 'u��\O� ^�6�׽5n�"ٸs�`!�� �#���B) �U!VH[�I�.�Y�ʫh	3� {4w�  �q����|B�\1�I( 0�j�d��8O+ ���P������ ��>��4� f娡��I3+	:�睈� s&6Ao��=�%0�t'C z!��#�]� ��U	�怯���� Eo���h�HFK*(�"�	o��_�,�`���9� ˻ҋ��� _u�|�/�3X�0���s?a���`Z� G�m��.�i& ���ށ��y�L̠ hrZ%U�rv��&Jm  ��
�}� -���=2;� f���8	�p�\�Ki� �<�ý��;���> TXn0�魐� ��N�Gf h�}��p# k(����9_ ����D@&3 ����5��$������[ ����'�|Jv��²��ܪ^~C��Y�tGZ�gfR�@`��	�.Y�ǯ��
ʳ ^(ډu�s�e�4x�����r! `^[�~���ʀ�?���::(�4��3��.�6 ���L G�@T-����0�?��c� ��`�� ;�!�����@��d�� �43j�5 �7K���� -a��}�� 
\��ht��=�E�![�:�".�� Z4�p�� aڕ�H0���^��sć��	��q� �����Q �h�0�� �
C�/�:s�1��)����L��<\�d�^�(�h'�u۪v�@�1�{� ���Ҟ0g� ��u};�: ��
��� 	��o ��C^� �3h?���}~���k� ��iX��� � �U ��D�YL ��[R��\ H0�G A3��� V�6�<�� �>���y����������\g���e��� ��YP��$ywp���u �B@�(-��|�rl,^���ưG 6(���3�>&@a�V ���7�o� U�/1��� T�S2�f ����0� �u�E�I� z����o�� �:�H9`��$|?,@ ސ��c��: ��X	Ћ 2�����A )�1�WjSa4�k����n5Ř h�_� ��� !ʾ[�?{z��%Wg�#V���U�O�[�	p�ڀ%Q��DL�����
 /WX�'���x��G�N���� ��O�:� ���hk*s �J��"�	��� ����C������ ��7M�_�:�4 A�5!��� Ӑ��0� T'��2�]��@)[��  n���rBt�	��� cF��CH�! �BYxV� ���1�&�K� �]�b:�[R�+� ��0 fZX��Qb �`M��n+o ���V��� � �]W~%� pO��ū�1��� �Y�D�[p eB%~��_ z�W�qY!i �侶4 ������� ����	��T l±8[%Dp$��'�JI ��lL��HP;b� "ؕsI ��k���oN��~��������zQ�hG��ZE "gc�~#��uL-U�X\[ ^sV��n>x7{ b'
�.0��(�r �2չ�H u������ f�B���L� ybي��v� �8�E�J ��2!�po5_��1�� ��/9A�N2`�_�
 	�~�/�� ������ Y ؠo�%�i� ��]N&�� ʺ��9�|����Z��MO���$� �F��,� �x�K��	z Ï�wb�� �W�|Y3a?껀��w�>AE�3 Ȉ8鸲:p% ���tV �'�:�\7�  ���1�� ^	ī�3�ߒ@��'K�  �����VS~/�1�~�n`{�� ]��v G61R�7� �>�P�%�J ��� ԃ�� =�	���8�P�� �.!�� ]�X�\>L%?�	�;��:�3��1�\�M9 -���	U� ���]#J&���\�Ę�ն� ��T�Ґ�$ ����1� 3s�	P�Ą@��Z�����D����[@ �؉�/XL�� ��٠� a����W
X<�� �h]	�! ��Ca��:k �
�0\��O{�u1 �es@��H��J��@j_	x �YSQ��~ ��2�[\*
8�/���E���0�$3W�KVe�%{ �6��
P-�3 ���L�5 �V�R���}�H�4 z�C0�p_ �/�I����(��`�U
a��#���������D��x?��N.����N` �����=�;a�N�����X�K��<�� �0�\=�-�v�� O�	����C ��S#û�9cv l��>�֠t 	\���f+ ��W{���P	�%�ŀ  ~�x�i]����؃w� �-�N��h ��]���t+�BP;�����a ��4z
�� �Z$1��� 2H_�Gi:9�΃�������� ���P�"�AB 
����;/� ��_�̲ G�<�액 1�p��I�	?K=����Z �ȹ�~}�X�7�� �����J�� ��
�����$DcJS�ൈ*h'�����( 8C�\3� H)ջsL�������� 	�B]�%�� =�'��� A0�.�	�^3�&����� �!�׋1�� ^`���� "����M(Y/�����	�� �ͤ��� H��_�"  Ցn�}C���M�6������,�uZ O��&q�>���%|r5g?\A�Y�ӰWl� ��sd��ʻ��蠷�VbM Wӡ+	0�()�\̫�) ZX|� 	˺�p{��d
JW�W`�� ��Aݱ$z�(�m���,4�W�F
N���������&�^�|h ��������H֥�N�Pќ�b�%��A�XZ�ID����6z� �.Ш��ʥ�� "(�� �Go���� ]����-^ Wa ��;�l�� 4��&����+�"�n�[��s! ���0Z��X�� ,_��Jy� ��@
��\[ �� �=� ��ha���9�x���a��@�1�@� ��״ H��ߦ�' �ҹ�q��w�5_���Q�O���B� ��8$��� h�щ�:�����+�k�z؈���S<�H�� 2$�C�8�!q( ��-��� �[	,�B��@����n��F X�͚v�x ��Y���8�a.�0$�^$��� ^�/�� ��}� �q@*[� i�_P��b X ��O"�![�@ ʋ(�� 	B�8� +b\j�V�����$�48 ���_IO�������؝�� �:����� �� o��0 9�^�� #Et���+ ���PW.� ꃠ�KT� -Zl�k��&�[@?�1�_ �Q�";�bʷ�u�`�O��� Y0�h�@c K��H��]���'`�� �-���p ���F́ ,�����:��?�����x��� A�9#���� (�Q�[_�Z �X��k���a�@�1�-%�M$X
�` ����.��� ���!�I ukh�d��O:P� L�)�� ��%�2��&{�ɀa�*��� O͠&`��R�� M �(�� 3�%���T�;��Xw P�0�(/ 3����L��V��[��C���艽 f�Ӄ��P� ��V��&J��� 7|�Q���`|m<�P ������$�KJ (�Q"� �X�J��< *�S���M� ��_�b�qAṆT.���� �����sA	�j/_�%'  d���N�� �m���|�4�@Z�~����_�:�V�L�	���ʀQiv�-��� �Y[� h�Ks P� ?-e�yJE�	�Ͷl� �PS� �O%�1@k>�� 	��h
\ Q�����;�[ �'�l�{( ���$�0�X\� nI�-0p��
�\#O���R$��	%/ ���� r�Y_�[�9ʒ���E��-�A��U OY�׫M"$�A �0w�
� aU��.?�,��* ~,�OytS�c��|^�< _p�2�L� Fϱ[UC� ������0���ڸ{�( ��X�b> �#ϽW��[ ��5�0@�i�sF� ��{!t� K�'���&	@,v/�~y�-1| %�L�� M�O�(�� �_8�!� ��-�����a~� �H�
wj<�� �_v��D���g��	R,3�ȽC�W ���{�h� �ή����3s`X� �[lۻ,T𳋦K�y*��������,uEaR�k$]0�� |鎛�;( �@�K��H -5��~��� ���Y+�h ��^�GW�u�!��1LPo��� �GV2�� 	`(����'|40�p@b��\$����  �V +�'�<ߑ �`q����%�@�}����'� �t��W(ˉ �V����1	P+ )½ ��!��h0 ����U��� �1���ߚK�� ɸI�u  W)ݿ0�\ ���c�F� ��pIJ�z�� �U�&��i ���/��E �����HtR�ʁÔ��P 	۷�$��\h=�fR ���� ������L�� �{�'��f }���=q�+ IiD�d�-®X�T7�`<� �"6?1_�[�O� ��at�
 Kޯ�FD��)�����v��3�V�X�6Ȁ�{ ��so��P?0�����Ȟ���j�����-Q� U�HyN��0� ��5�l�&H��| ���@�L,��L ]�YI<� ω�Z�^���@�3 ^$���' ������*΢Z�F�� �q���ñ
�y�k�v���.��X�gsL,��� �)�-& p���o:N��@��c D����(��RnZѝ�Ȝ�r���v����@M�������R(�/��	,�� }QwI} c`Չ�� H	�_湠
 ��?W�%l)'E#�R	�� !��w���k�$�^`ڞP� 	
Z�4�[ �K��cXP �EN�O��H��t 0X�pa �)�[*5�����hbݳϑX�$�/�@ 2�(Zp� f!�KS��	 ��jY�2 u=��f)�d҄����S�
� n�-c'���u `X+��Ed�W���mG'��Lq�Ͱ��9/P�����n3�~X�x�]E� �:�R>� %�A�[2�_�� b�p�{X �5���� (�%��rS _���Q�pF�\ ��� #�{��vj	 R�_"ڰ �Q�%��y��S ����}� ���!�� | J3��0�/��1t��.��Y:4���亜� &��:�?VN;�Ā@* ��X� ������$ �U��^�����(���`�����h� C1;�s��k~�, ����B�3!��סA��0l�# �7��hK[ ��w:}�b<]��	՘�U� �n��b�H\�A�����c��" 2�V�$��1�U���<����#�^��lE/W a�Q�Ԑ�� ��S}\j�� �A�kΨ	 ��nm0�Q1�>�J!�B� ��� �����C(8���p����~� ��XR)غ �� ���9� �QK�V�� `��ˋ�	�@��(c�h�cg� &%4����� ��1)3 I~�F�A� �R�d����o�u�-j:����������Xh� a����%���Hn� �����-rO�'��$�	\p� c���_: =���@�� dB�$\�	 ����?�����Y=�֐�,�� �7��� ���xD	� ��*�Z]�. 0��}7� N_?K����3xB�� ,�_���=�L�� #��Zb�� �L�'�w6 �x�K������	`�;,Z\^���nyT����`�4@�˞(  )��KO	�[ |���lP���0� ɼ����%��\	�- ��� �U��~R d]��^��K��܀꥟s��Ct9��?�-$��?� ����2��]������?���:�f ��;�)�]D����� /h�Z� 250�G`�� '�o�(�3�`
2`Whlm�ȵ4��|� �U?��0 �l���9�� ��\k��u ^:� �_t[�
����ܺ\?À�s	 �uD��� �k
��v�6 ���'z������W��T� �@{C��x{'9Z��罘�J ��2�z�97 \��V�Ǔb@� Y���j
�`�<ڻ0 �I�]�$^�)�P6W� ݀���!_ u��$�� �*�ؿ�� ~�5���I����P��s� ^_F�;�G�й`r��N�����T�X�Ar��q��;�n _\���O��� 	���^}RT /�)���4�� K��� \2�QU���[?�FÆ.��8�@���9͂X�WA�9.�8N� e�Ra�~��
.���"�Y0�L�o!�% ��za�P��$/�&8� �j�� V����^5hv�����NJ� ;��B%� �/�3�#�Q ��'~�>P � ����K��`��^�p�St1'���s(/�5?byW��"�}� ]xo�B�X*Q���0��� �����5� ��&�$���]$> ��N)n� 
����.Ө����y <��wS�⚰�;�� �.�Me�
�&�t� kZ���` �р8��J �^���#� ��/��� s�|���� S%���	с�ۘ�+���Y ^�ɖ�mG% H>�P��� @�)�SU�0 �B���>�K�6�P����%��U �b�������+�sJ �1Y!�[��?��@.D�� ��45���8)��O(� f�"�K.F%noh-0�Y�� ������P J��H��h\q�G�D;U	 1���H�l �.�v�#�`Wt�� 0��X�檧 `����>�	��h`܄��� 9��N�"�� �	
릨4�� y�vq�z�0��рX�| �<���2$� 
������w��Y���If h=OՑ��0 ���ٺFn�A�3��`և _K��l� D�Lhԗ�2�-x�ƒ �	������ i�(þB�  7��NF�� 
�h�8 ,��C4� �1���l-2$��q��p=JX�;� �KYbE+dL' ���,�� �]V1Ϙ��X��
������S?r��j3d����# �sK�	� ��EAW�D&��� {���� ������ S	��%���H^ ��?�� ��g�互�~\ ��d[�)�� :�$�����	�~k)sP�:ꀦ?���N�>��fXY�%@ �v;d���H� 2��t �<X���[?�րA2F�W�$	�_q`\엁'PН:��V����K	`��^X���KZ 2|�V� ����}�ȿ ����-�,��5 �+
yժk�� ZX?�� �O������ �("�zĪ# =�J_�2* g�/N^� �(��kG�mH���b#���y!L�_+a^�tj�/����Ȧ�v���DR�rk�u��)+7 O��5q� �~*�"ˋ �XH�I��.�{��,�&N|��/ZY�2���	�L ���Z�}PCKV���h6 �kg�!�=K� ���ؔ#?Ãc��0� V���j�!��/AX�k��� �4���# 	��łBY c��٠�>$zɹ�:#`m1.� ʻMN��J ���I�3� ��Q��_/�7�B� \��`��}�S���m' ���R(^� ��Z�1 ��J��^ !�Rb��qv<��_���w����.iX`����8J�'`��>��+ =�P�J ���dE�0j S��)��J >�e�`�U1 �C��Z״ WApk��!�5/�L�� ^��Qu�L[� G��%�h ,�x�i�U���jNb��w#�z ��Y�1Ӑ@8�%p �MP/�A�Q�
`���'�h�R3�4��2�]@���:���@��cQ���q&t(n��4�B���)�P��v�܁��? _��� awC(���P��� ����Y0��R�(��w �Hᅘe<�] �_�y� ����$3�� �/hQ��I�A @�nEd�:[fX���K ����y�: �8���ڿB mU\�����'(�upQ	Ph<�� �9���\;�� �1��UM?� z%H�\E ê2�@Dh�bc����\�> ���Oo� ./�U�v �P*ӝ��+��ᾐ 3 .�����t N�(��;T �[S��r�s^ 'pi��+* s��u�1 � ��Q{� ���%:H���yXJٝ����5��"� ]�;X�wnX( ���M�1 3혚Jd쫘� ʽw�
��2�]��� �Kw� 9?��*ǐ� �� 7������]��-��.a��= ݩ�Q�c2��q '?[����!� J�aupI�Sm_��*��C&���J�r��S~�y )�{��W�  ��1�0��RyZ�� �A�0��u��T�U���\Iv�:��@ڇ<� ����Z� ����. B��܋�%�<��p
!��kE����� 	'S�uȎ  ֟�{���b��ܘ0�G�3 ��r	�o�q ��ѻ� ����YkL�`� �)S�b r���;^�s�������U r I)����w[ٮB` �xtv/#��<�����K���3�A� �S (�Z�*���>���������� Z��6ma�,h�`~����B� �_Qƹ /f&=	O˅j
�㔗��Mu5 g�ε�=��_�͝��� �w����Y �q�	Mh �4������ ͂���x=O ���(��)�1�������$���)��& [��QPV��]̻�K�  �[�"< Ł�жhA f��I�0�_ #m���V��n��4����� :Z�sA�� C�(���5- 0���Au� �?��=�� {�����0-D������ *�\/�� %Nx	�s���r����\  ё��wģ?���C�Y[ *���D-�� Z7LM%?� ���&�t�} ����,����J��Ȇ�� _�0	\h> ѵ��S'pR H#�@-�8=.� ��"�� �]����~�I GT��Vy �w�`�� '�^]�7;-d�@\�,��O� !���YX����܀��H@� �Z�1��� `����X ��zD8x�	 Q��l���t �����?� _���x��\�^aDU��V� �3�L)e��^�â��uNr� �r�% ��M
,�Щ ����S��� �6]h�0 O���@��ð9���;���z>����B ��	���EP��] '�z�� �	5�Z
�~��� �ޝ$���ֿ g%_[� ܶ�aS+�` �FI��/T ����D�� 	]� P(�� Bւ9�"m�Z�u�j?ೱ ԁ�ÄQ 2��8E%�� ���f�J:x(�ٖ �AM�/ ��1I� ��*q2}% �xH�����|�-���~8 \�J�!O�{ ���w�k� E���������_t����X[��8N������HW	���\����1 ��a��P��S)�Vf~���Au�<��Z����S�z�ᨊ�h.�`�{>��A��2*�t�\M ��X0٨��Q� �ݘ G-D&�� !B�	�� 7�И=�I@ AO+��*�� �N�%��|S�<?�Y�W0�5��� �&S��~� `�v�bF g5,]z/�3��ߘ��@��n�R?�P[��h�<q�NT V� ���ϔ�J� 	����{~Q�� +a�!�l% �U�B�"W9(4 Y��
�\��R�f�U�7�� xo������Qf�}	 i�4젾Ȓ ,�C��0��� S
��Ԉ'���0��&�Oh{Ѐ�� }w��U�_^S�L�  �	����? 5l��K,���� -���Df� 
�E1W��` Q�I�+��� %�y�  3*��.���� 1���2�[ �l%Z/��S����<3a���$�X&Š�W�� �^GE��) ��	�� |�v@�-��y �P߅�쵸 �ы_)���}� ����Oj����� ���� 1�. Z(	Ҋj������ ﲁ�	�sSf�40�`�q�d�]ȑw !��y��� �6��L��� 1��5���!�^�A��tG*� ���H�Y��.[ >3�` ��*���� 6.V�	B+ �HDߐ(]|}K�7`���0 hn�ӓ <���튞�(З��HK���j��h  i	��^p� ��U�-�q b[_�T�^t'yz�ް��W� Z�) ��`�1Ӄ�ߖ�Dho����κ=
:H0����e,�={���Z�-�b��� @v���Ga �V�ۑ��l |N��f� ;�[� $	܁
u�m �>����A�x��+P����
� �!��F������ ��V
���S� b��1�J� Y�����o^��W �Z4���r�=�j�>�H;g�z �|D�-�A� ��5��1 K��ȋ�� �#��Խ�
��#��U�1���>7_���8zh {���jr� �Pb@( ���K�B�:����N�% di���Y/�o	����Bk{�$�� @��-G ���H�.K;[>��] Ծ3G� m<�h�?K���0z|��X��@��긒��ps��kX��R_ ĳ�	�� F�(�Q�� @�.���� -V�*�N���� �����Uc
�����k ��0j��L_R��\҃x�Z��~ ���Bf �$�L� KQ4Y�^u�r�(�>Sw�� +�a"d����9��	�S!�G��� ��]��  �%�X������:� �8(*��� @鄊<\� �dh�{��e�� !�(�}"��J^�^ @�e�	����~�$@E�" P��A���P� ��3�:] ط��X�ٿ���^0B�P�F ��`� yT�2��D�� ��h��f� �:���>%���p��A ��Qܔ!�� ~�����@���%e����*�1�<���-/��! �ӢH�
��� ��zx�����?�iP-_�|3n�ro�&�4DV �G<$�A�d����w�� Pe:�c�3v� ���p[*�/�Y���� ,�~b�� ��JY��;������N2���p3��8` �+�B��' C �i�� .m���]@?��( ��ɀ�� � �bj�`��@���� tP�#o�� ޛ��h(b�G���!�� �n�o
2�� �㾱�: �Z�H �3���-' [~�XhK�� ��3����#�e�*��r�����n	� S}/KУ ~J�+�Q�XV!kb��@�tK"�̽��D��	� �<�@�l��o��0�a ��'*�u	j  �ŉ�1� =�R�tP	 ����٘$�+'���Q�M E?W�`�?黃x��S��E�`��I�c0[^�Z��$���	��� ZE���=�gHW�$w�X�0�9��Ք�5 h@O*΁� >ٽڠ�( �W��,)_ ��GRD��g!�o��W�T� �-���n J!�؄N��Z�Y��;`u� ~m\ű�c� �s��!"_� �z1�O� ��AY�/��Q	�P�_  �LI�(�z�������Eh`��XZa,d�8����� ���頟x� �ˇ�O���*����!����-����, _)q��F �`ҽ��1 �����
��(
��m?��b��
��!�*�R��(����� ��/ipQZ ��WT_���� ����� �#mQW�0�%8`��M �
�"C���j��N�ZmK3���h=��f ��x���Z ‷�Wd0% ��߭�n�H�~ ba!�8�� ����^�� ���Q����DS#	�>s�`T}b��u����pæ���L�� 	�[�}3���<� ����_ �#P���r�\�kU�8�[���oh2���
��R \��P+� z�1E��j��؝��<� m���Lh�� @l�%+�� X��0Qι ��ʋ � ��HT��u� 	��p�X+ �����ƌ �Y�0p��X  �[B%�D� ��Ō,
ʓ )�Z��!�0�-��ӿ����U X3׸A�k V�j ����i 
_�!�-J ��*�3�	,�G�&�@����۵fP�ֈ� �T���YR8 -��	�vH?� ���*�q u�'.Vh� 7~�b��-R�� �O͸� J���� R�5�ɳ�VFI ⹪氠ڒ	����2��$n8��`��L,ė�?h���F��������
)��>0��.�M����p�K[��CJ�30<v�E��(1����Sn�3`Q"`K� J�}P�w� a���V�?�ѠP@]J���$�<��������x�� ����z2�X������� ���
Z� �'ASy�k� ?����$uo���-���q� 
(�ކ�;���c(�����(��������s�%��e'�� <=��{" �c���^R}·x� ����5��L_�|���t�� p�%#]�[����Q�z�0�!(|�X���2/XAk.� ڄJW�*f$9+ (�Z��� ������ K���T�BV�	>��Ua`�.�� �]_� �"�B�������椔 �iǞ
�8�%r *�R���T.��;�r-���C^��N�
Àx�͐� R�z��S� N	Ȃ�[�HUq "�x�!����]����Ь�-n�`��� ����Y��?:K:���1��\7� �?ȫ	h� ���,��3 �I��j� v�)� �����<�B�г}t� ��0!�.�� Ć'��z�`U����A���I @h�g�D $�=B�7\���q���0�? �d#�N�~i|% �OX��D� vAT� �I�]aH�W�k� e�m'�^1 �bi�:��5 ����#���W%����]�� ��l\�9у�I��N?r� @U���>� �G�g�����ѐ�T ����q6b �閺�3�$���0�Z��h�+�������]���G� "�P��a�Y�5� ��n���� ��*�@E	 3�h(R}5Up���\+�C�R[h�zH�	�3���}|�?4L ��j��	 �K��Y�8r��v����ʀX �i�f!ԝR0��C�8he p-�ɦJ���Q��t>�(� Ȳ��jXRGv }�z/Ovϭ=*�\�������� 	�cH+�� ������?�c �/��-A�X��>�9}�|n�u	��q!U \UL��+ҴO�! ?��  ��u���� ���+&$�(N����S�̟��Ձ� Խo#rt !���݀�x[�����) ��]�}a 3�T'��� S�$5���Q��� <#� �3|�6* L��B�D|�� �䀠���;� %. ͪ8:��!��> �%�p��"�������$9	P���?���� �� #� *���@,\��?�x�A~ 	��Б� 3h1�\��P� /��;u� QV�v�1 7��d��0�8��I����� z*�S��0���.yb# �<1� O\-���<G�@�Ѱh]S ���3	� �"b�Ԛ�闬�' ��V"���MO��e/s� �\A��od��b��pK� B�	��k }8SΈ��` �h��!�Y��o���0�\a�`���`^�۬�J|��0~ �P1tu`p ���;�K ф�Z����� ��"�����0)����� �2�x�IQ`;Z���'X�w�-n�D��a-��U0 �+�°4,� \�bl3�� ����n�� /-7d�� R預��0>�:S�ɻ�4��� �,fto� �-�z0�)�]�sN�`�u�2 ��hE~�l&b�〉�.)�	h
׃F�	��p t��& �K%!�P�{ �^�f�����p� ;���d�sx� aJ[���>���X�{w�b���ֻ�� :���u
����f>^釆 @	����n9�B��W KR!���0 ��Z�'�^ �ʡ��Q�  �T�.h�&C&u �"SG�� ���R��� �Ŗ	��S&���N`\��O `飓y�~ R|�SD�{I ��uOo�� :�3Z@ב ����?1����m���$;v!J�0/�}��G��
2� J�Y9Љr� 8p�'M[�% h�	UH
7 ����;�Z$�:~Y��bB�!'a���u�X�Z���P �n
�i+�|'~��3���z ���$��Q K���.3�+ ���	�=!+�C��;SJ< ��Q���l|>�?��O�J�Y�#�)
@�P� �5�b��� ��F�1u�s���bc�j�����|� Kw��S�BsH�� ��AZ��Hug� LV� �9Bhyt.�� �*J���|�� _��(��P�
�Q��Ip� �+�	ʽ&� �ׅ����8 ���|0 �J�¥� �����z� ה)P��� /��a��+� fh[;�ً�Xʯ`(�]w!�h	�Ec� }޵NB~�&��_ �V)�; �8#���� �.0
*h t�i(V�2�<�}�e��D��z��� �_/X��Z.���| �NV @P��d"<`?��q�Y+ ���(�Pb !��͠ �� ��%� ��&�V8q� �;�1�(�� �ld/������XR_���� ��. z��!D"(#���_���}��� 5���^� Z��l�	�&�q�-� ��{���T ��	���aD?�i=��@	R�z'�KuP�� ����1Ã��Z �ٻ'y�K ������oN.pX�$>	�W�Y�9��C(1��`�[(�����LA���0�T �p�2����΂�@�6�x	y� zĖ_��u�:���h6>��S bxp�i{=+�� �� l�8F�1�֘�@ X	��j�U� �9w���Pl��p� Z0��:�A� ��X/��~N ���,)�`�.[�S �.w�f� ́���v� ���E���Q����(����TJl&X� �܁�� ���*�݀� � �+�f #�h}W�� ���H�ψ	����6�z��Ex�8O��0M���r� ҃�!�$� �/��l ,�̅W� 0�S��)�%�4 [�ݕ�  x�̌&���	"܀�1)�Y�J>W�-@`�� �t�^ᒴp���~�`�# �UT�P]�H v�!���} Z��"X�OW��N� ��(�1'�)�$^��lZ��+��P���VL\[޿ �:� �� �}�P��2 ӽ�|oI ��U�� h�}΀� �Y��R#(��8u�*W3���� ���t���\| � ��$Z%��wD���R	ĭ��P#�
 ����ݻ��$ �W����� �"�)���+�}F�� h�:;1ۣ� e|z�p��	\������/��a ���	��,�f ��Z�]��"�+�I��:��K����|) _���X4
�k��*��[��( �	o������R �/��( ��zܬ�� �*K��˞� a��:��� �پj<�����@���^l���������R* ��c�p{3^ ��,�u<�S ������ �c�V�t� �9=��q���H��PZ|�
�=i��S� h/���1����`B^Y#�V'��Ҥ��fJ o�/�[�2� c�	���u1� Hh7j��L>Fw�����b~���\]j�Z^��H���t��*���� ��r�9,u@� �Y�� N�jL�-0�����: e�	}m���� 0X�J�:�ov ���<L�p���1
�� -	!�Z����ؖȕ"���WU�\\O Wn��Y��� �[�#{�~L����K���T�� ��9Y�^� �c��)؁g�;�� )� �[�o�W:�D�0��!�J �t^�6�N -��0�۫8��P@ƸM*�G � X��� 0��*�����O�����^	��)�W o��\ 
�h�H�-g��G��5�# ��R�>~���Zj7��X	�]�� ��������h� �H�� ���r��D� �Bu�d8� 
�~2҉� `l�/�dp�Zfy���	vg �8ݼ c������ [U4&��)� �A�T���X �͔sNkjS Ch�JY-� �R<T�A/ ��3\�� �(�)��1� �>��+% ! ��/S� $���^ ��ӱ_e�t.��ܼ�������Op��I, x/���%�� HN�!KІ���tZ�r��R�x���%����� P�ZB�:O���v� ���>�,V� �(~і� �����N �9� u�'H ��6�z��x��4�e�Wg��: ;�Gf_ �P��A�)�!�E ��a��ȊN� �D�Wش� ����\��o~6� ����ݐ��{�|�(�[Y���$8k��+��_`��� !�X��	O~ �C���(:�YZ ��x�>� Ƞ�q{��_��Z�x���U��� -cy蔗g���/ ����� ��~@��0f|� Hَq&��2wt�l it� �|���� ����W ��8,ջ�B ��wH �[� @>����95R�2���kDm !�`�È��/h�R��Fb\�� U�ʻ# ���y�.�n ����NO���UF��=Y� 3�fQ�P�-�ֶY ��`g!��=*xB �H�|~X�kep�2�� �/�&�� Ű�$��Q� �4j�º� E��\��&� L���H~� ����� ����`���e� m��.1P��h��KX j�� G�aMv��U^?\� ��K: �J�,��� &[��	 )��`҈Ǘ?�����Z��ʟ ��y��]� �B)�}Y�� ��"�_R����KҺ�q�d~ ua��Z���>�'"{Y�<0�&�H� /�	ZW ȾzN��� ޭ����� ��vJ� ��l�Ҋ�R_(��E��K�� ��A$��� �0��k�@� ��>��-lBGJ����*IQ�$}; .�^F��� H�O�f1�,rBX�]U������ ���bv��xP@��!�Y .b�Q��# �ha$ftO�t~. ��8��!g���򽁀���2  ��HS_�.0��y�L�� ^���v~I��-� ]ҷ�h�{ ���&li 1*����:�?��v����� ���]�/ 2q�b�LU�f�S�>%X�@�+���}	�P3���[� c8�Xh�F ���#� d�5Q,z	9t��M[���# �Z��b�v�]BpW�@�:��K����4�ؿ� 7�� PH�%c��)v ���6��KL����1��O/ ��Xu^Vb' m�t� ���U ِ�,�� cu�ĺ<R U!5�fI��6 �k1'�D�- ��b���H�� �1/��� ��
�[���į�0c�8��s� �,%��� Zy��*]0.�)� ���� 	|p(��.)��� ��5:K��Zw�@ ���57XM��@�!H ������ �e[� d�?ȗ�'��;�D O-�~�Y̥ ��W	� �.鐮&�z� �1_O%0Z<�QÓui������ ��[��� n�N\�f��;!��)�_	�l$ qQa%vbI ��Nm?� ��5S�|��!������9�� �%����� 7h�x�0�^��� gށ�"� r��a �m��b��B����f;�ހ�<x�c� ��N
�l� ����� ���� �'���=� <�K�� �\�8��� �/cI���L���Ë��Z�1��  �Kr�.�W�����6 �y�.����`Z �/$�M��X�@E�Y� �h�V�*+� ��2��j%}6 �(�P�S氢 �R!xKA�x/ ��淬t�&a�f b���� ��c�6
5 �v���Б�~�B���S����.Cp�L��{�$� Н�͡�%����8����p�<H(��1� ȔY)� ^�h8B�K�A63$*p���x& �kT�Eg 1����Z( ��m��W� �c�(�`� �_2��u�HN#���ږS�@X��9: (���l%�#2�C�?��!?ȷk��R �Q��� ���_�?~ �O�<K�X ��*��� ���5� ���Ж nX�0Vt ��21q�T� J��;� ���'�e_BG�[S�6�hr��,?0L��5��) P��:�/��:pl����� �����;�` �h�+�����0�S���ԣ �	^���� ����M� 
 %`G��a Z����",�` ,)�T�� QӹPZ�4 �����Vus�,r@����M �J_��#��8��". ��d�&}9O!�� <%�s �>�1��n a��� ��_�)�d� �(Y��}}� U�-�sJ� ��]��ܨX< [�v�x� K�@�- ��\�B�S ��ɗ~f��et
�p�� ��c��8 4�ǻ2y>	 �G]��{ԒM l��a�^u� h��齖K ܃�g��e���k���y��YyX 	-�v�F� Q���N �_����>[� $���� ؈�di%� �����^ �?����ҳ s_~���. 
��+�,� �K E���b{ �md�I��< !�	���#� �R�qN̮���ZP�5�$�� ?c��3�R��uޯ�^.m�����+ ߾(�R�0 ����P��}gv*N��>���� 	� ��oR� ۺ�T3�W �C�|��� B,������ ܼa�=�F� �P��!K��e'���� ���-��*��P�_[?�E���9��� zD%	0�tk��N, �O�n� ������K���	��\y.� �E��� h0��J]�!}W<�F��;��h��0$�MW T}B� ;�l��@(�'�U ����X�@ ^6LF���,
8v ��xE��T ���V����8���]�pp 
�X�:���ʏ@��I�PU�� 2F
�3Z �<D����u�%�6�)���
��\ ���*�P���r��!8; ��[��k <��!G $��FNH ���(j�> ��ɭ�k1o�7)���3 �䡯HSQ dt+�0� �P(��@� V����� ��f1�h`S ��2���P@<�� ���=�����X`c�uar��J��_B����^�� g���Z �bpWy|(�P]�\���8t� �/[�>�\	:���|��n ~گV	=��Z 9�@�#�� ��R������؝ �]� �.�r �鞺�� �	�pc�/iT� �-]�bx��E�	��u���w{��^����+ �3�䬫 P0�#�2�tx��Sf׉��LX�3 �%���q r5�`�OG�  ���':�y`P��D�Х-�o���,��@5) �Y_RK�V $*�o���k}� �-��_|N����a���� =r�K�lz }����X�B��R�Q�<���ä����C�]�� �@�� ���(O���tם}��� ��qE[�
 �p�.�� "�4���� ���ԜDCHo$� 73P?!��* �
��}t wT^\-k% o���]��O�\�:q�L�  M��S} U�D�];Bq� >���F8'
 ��y)G2a� �4*��� 1����j$�N��c���R;�?' �ڛ��#�Vە�0h��P�����PJR �t����	�S;(���> 2��	���@�!��O��I [�Ι��{ Dh�m�tb�/�T@�`c-N�0�M��`�!�����B ��o�V?bz���� �h���, ���EX� �1�{ˎ �L���j0 �W#���q	�� X�5�hR� C�2����\�T���-=�a�,p�� 
ƋއbF� �CeqL�':^X������� �N��θQ� �������:���$�AػZD��� q�|�5j�.�!� )�Xx��8 ���������X� �k~�a�� �պ�9���"4`Ht��U� �1��� ������N��.�������	P�*@PY.� )�������Z�yv�r|��p� �W2�Z_��p�;�0
�6б�� �%��C� 9�_���i;��Hc� �� �P'�� �}U`��XR�x ��(��@{�p7%�b\���:� 	(ǵd&Zt ��<p���� �����eQE#-�iȄ�w��)���B���b~h\K� �*�0�C `��'��L�.(�ߡ�ip~��-XvK RV͵r�\�2pw#�e YP�
�	�xՠ�?N���7#��/��"o��^��wI�~EUO@��Ϙ� }gQ����� �r{�u��� $	�Y��U� �»gj�|� D
A�_�8�� ���^i�-���n��O,�u$K���@ۅ(�@6�p0�����J��	\�� �g��+� ���1�F ����Ԕ X�f/�����?)�ڀ�1� Y���~Ӡ� �'_D� �%6Jٻ� ,��hK#�� (
����z" �)_ę%�9�E���[� �:]�@*% �p �N� �\��� h�S��P�� DR%/�"M��� ����(:��]ȱ)� �J�м� \�zS�F; �����xXV%�"p��<�pb��ן`�V3O߮���N�uSe� ����q$ �v8ȱ�Y�������N��F���J�� h��o��½�-�{y����	K�jD�!��-��Q��!Z��-�� �����R�N��Z��N|��>�?�0, T�b������� +Ŵ�� P4=
�Q�� #��Y�N ��4��<�}T ������A �M�����} ��^)�!\0�>���� ��|��/�" ��1��3�,��� �g�h�7 
(��_��X��+ E�Y>0>K�8W�����<-
���sx �_��%��q ��
h�MrO����Ȱ%�]� �"\;�. ��,�!�� b%Y�Qy�,������9ȗ >�~jY�� �]W�S �E����h �R��7��2p[��fz��BRso� �X �|�O�0�( ����B�%q�|��b���/�AX� ��"�7�� x����	\+Lեz�P��y- �Z;)�G� �XRb��E �B�a�&!=/y ��;��X� ��1H�� �!I)�( b�f@�� ���X�
 �����m �O�E\X�s7}Hp� 1��-� 4�m���.K�� H���_,fQA o�|!�� }i�$;�� (�&[Qg��?�U��Z̀)>����'u�����F�����:�4`�� �ٽ�����������-hU��^��D�HP� Y5�H<� �MJX����tQ ��a%��b� _�K��!/�� |�V�#,( �@� =���G��u�9	 ���V�:�Ӱ�`��΃�:�C��@� �֙�93����1RfP�_B ,Zu+8Xνܖ��@�S�.P_��(�D��� Z!��H�E>�/ ���%\��+ ��'(��-� ����2Ȝ(���4:���.Z��	�� 
��B� w�>� Yh����P�� ���0l���"P��� ��ϊ�� ������ 1Wh�)����e]"��`��*�lж-��˧q��z30�@��2� �Y�Ho��X� �U<�b k(׃�Կ ���$��C�ՙ���pO (�Ef��Y �L1�u�m���j#�K|�0� L�3b�YP��TX�p�O 5�(ҝ� �'�
Y�$95� 	1�&� �-���(4 t��P2�� r!��Ua�� �.�C�< ����XAU  (K���W} "����ݕyA :nmfILZ ��[��������`W��!d����(w�� �J3�� ������;u^ $߀��������X�� �)���W2 �T�	�nS ri�Q`z0�� �12�.��;���`����� �T��i o��\R{�4� ��
���� �S*ϻ-F $V��HJU �`SضN�(X[�G�h�&1 w��HN:��� �x-��Gf�1�� �5ui, �y�PNj�T7�U��%�� ���#�� �0�[��4 7�A�.�: ѽ�Y�BJ� I�!�A �]~��f� �b��&{^~S:�����Vў@�0�-1�C %�{����n��p��R� v!�Q�ǿ ����H�	.\�!� �br�V��<�?�= ��p �� #�t�*�z�K�@�`DI��(G� {�\S�&� �1���ݤ ֌w�al� ̛�1\^I���n��-�Zژ	<�@�S�!��;�"���V����x�ݳ��71>��| �2�<��[ ��9"��p���� �:%�;'��
�����.�N�����֗��v�UF�t ��(	�,�:��  �@v��\ [�P�uiK2� �qH_��+�5N-ݴ�A��3� \�څE�к=	� �F����� ��Ȇ��R
 ��:*�v�A ��.k�h��<� �K1�*�U �x�\j	0�~ i��U�|� L�}	�Ͳ Iu[���� ^תD@!����|hO��6D� ����(�� ^���.�� Z�WjF� Y���J hXz�`�R� ߺZ�QH�09��	�^���. �=1�g�H\��'�K ��-�Dg� � B���� ��}��[��B	sk� ��8! �`1���;�Z�:sK�����q���]��о���T�1�XR��2���rJ�.���@��R z������ �Vk�Q ���:R ��%��H�H���ß���-8�㥄��++� �
r��T�� [D�36���:|����4�� ��Zh'�#Ƕ���O� ���8YN ��X����<�]���y�'i \��o�&�)� �~"�>����GO#|�Pb�f0�����Y���Z�W���P D9�)�G��u^?O	����Ĳh ��+K�5Z ����e �dh�Ks J{򘁰��˝a��� P��fh,���鹽د%(}�R�Lk���
���F��JΓ�x�`�b"� ���(�X^7 \�Ah�r/3ȭC��%п]5���X�; �t�R�	��{E<K( 4�<2&�y0��P����"� �8�{^�k �`-!�h1� ����mU�X�� �x(_S-� �¶�	���|�����a��9�4FB!�mxU���w�IJ� ?�zx�3�� �S�1-d�� �PY3�X!v �"�h�O0 � ��Km�I 2Y�~)�� "��}��� H���|�'� I-qg�" p������-f[^M �F�e� �Q��� �y�S�� Z��C��] (KȊ
�� u�Ð�A �eT�!�_]�N��'��� ^0�\R�G �>�W�O
>rY u¯�a�� �R��< U��`��\H��w$��#��!�0f�p���&�Tm Ft�&�>͋��Ŭl)� 9�޼C-\ ��pX�R w� /���f,�@��� D	�����BJ�(��0��q��李�@�[@#� fR"Hܟ1 �3�4+M�	�V݀��� �P"ΩĄ2��`����� z�[O��.N�b] ��\WC4� �}n<��2�t� �w���V� ����}� �%�(�;�� k����70��3"��Z� �!Pu�� �ũ�s�,��H��1@��G����0��' ��D�5��	�� L*�[��� x��R�$ ����H�(q ���"a� _��j7� ��&<h�oWO�S"���/� � �@v�OM� ���Z�dD[ !�	 ���K�;Sۀ/�v w�ѕ����G��gc܈�P��)���
�����\�� ��0�y/� �(�]�%��@�������B0����(� P�������~�X��Q��< �2Sd��� 3�[��K��������)�^:BiT��ϟ�v%�+� )#*�z�1 ��o$�v��ɸ{���h;]q��QA-��'�1* �a����W� �������( (b��&�� ���A>�8x 	%�m���9-О;�����Qp,�t|5�X��9~/ �$�^��	Q0� ݈p�� �=.2ʻդ�3����0�Z7�d�ڜ��@3 *�^�r�ԍ Y�`~e�x9�����uJ� ���d[�4 ���c�8�� ����� ���ޮIM^�z��@�e�9 �7% ��}2��1:��Dn*�)� �zxN�D��+0I��O� �n���>� �
'�Y�%Fav� 1����{T �'w�.{ %e�-CZ "�U�� �O��A�R
⺀�>�Y�l� t �1r gS�h^	�2哉�?]� �8���X�=;	��|��8�8 ��A��N�� Q� �IB�d�.hj ��\�`�� r�!��1�?� y��N2�n� a�� ��A�"���2X+�C��m�R0� �ؽ ��s>� %�a�41�����JPS�8 _F��0�����P�>� �®����R3�j��õ;���],��}JPn$ 1a��׃���S@]��4��8�:� 1X����q�3��r� I��� ��@H]�V"}���i�5_ �/
	�& ĠtW��h 73
���A0 ��>�,�q�Zo��~5���VuB l��.�'��D������[m��� S� �d���Z@����3���H ��j�@v�75q�1ZƻL_p,J5 ��a �� xC��"dl@����$�_a�e���~�K�%A��D�y���h���	��"3�ct��V��N����W���,��Q��^*�a6(����r �	�ufs� !�
�Ag[�<�^>� ��U�5� �\�aqT� �K����6n���pm��� 1ði�����2J�>��^f���BZP�p��k� �y��s ò<�@��� 	�P3��E� �M��L� �`�]�Ϙ;����'�,��*0hֽ@g���� �
W�܃�x� �E"��`r f�u��t� �J[�t� ���
���:�82��A@r�� �,� �Cѯ��9č\> MB��wE:P�yX~ W�hUZ�' �Ӿsu�� �+���q��5R���xW +���X�� ��j�;x5����.fP$"k \D!�cI �����Z �
��|�e 	�{��� ��b���]7S�@�5,������ ��jI#����[�� /�8IA�n�?�S����wյ�_�x*����� �PJ���}^ ��G��SM��@QP/�a �YX�pH��h��P� ���"�.1 �t�wL�_j�� ��<Jt� ���N��Mxg !ʮ��/�� ;B��8 ANZk��;���]�Ru�@i�60V� Iݱ%Z=��.���$�  T:H��Wَ �o8C ���5��~ ��a� �.,*�Q��/�ȅXZ� �{��R?�bP%�^��?��� r�߁\ ���k !� S��uA�.}J �^'hH�%��� �+N�����EJ�+�RPU�`����ǵ����L���	��
!臛K���; �B�<��\��N�ǚ����[\�a-Y��u% 9
�\ S���Th�4� ���V��R�_�� ل��S��)� ���h�IZ #UY���� ֫3�%K!V�?-�߾7 D��e��4PT��z��0'X� �ͭC(��?��	������N��J��� �E��)�YӦO�`�N!X@ l#��s9 )�,Z/�5T � ���c�� ������,f-|�UJ���Y8hX 0ĉ��n `y]��@���aܽ �>X��h �G�&�fp� �� ���Y�����q�` �A�
�>��Ve	��Zy� �D}L2!���H� �\eS*_����Ͼ��P@�'W�����@6��� ���S\�����艠� �:g��� �����\*����	0�?�� OgS�(�8���׵8"@�7� �V��!�* ���0�Q
�r;�_ +�R���p8 ��Ê$[X�@�3H�a�R� _�v�
i^$w��@����U(�GL�v R< �.��'�� u�mF�* �	@
�������2��0��|1����� Z�i.@L�
�����fAMX S3���*t�h�V��W�\��yuP�<h��r�X��43 ұ�*�ס䘁 �+��%#�� ��������&7������o�UV�¾�w� �������x��>@� �d �"�$� ��*��{S�@�nF�GKŁ�l��������XX�/]�(�ܐ���vqP��� ~�ƱuTL]������&p,�a���ژu �n@ �H8������k��T�>� ���i�v����YP�y�� /b��_(�o� �7��t ��1S�<́ �I�[���Z�4��Ǿ���ؔ(gȰM
{�P Bm� 1� �#�Z��� 6��T �1-�U���u\Xs����p���'<�����Y���qg��n'� U.�/�S`��
�L���� "k��k(��_	�� %�FwKb��{.�2� �N�l���/��0B )P���X
���&	_���'%v]�\����cb��u� ķ�]��x �g�h�Lz ����:��B %i83��!�/���A�1�;j� Xq_b0�;������
B�����P�ִ�W�`�D ~w_���� "�P�5�� �̴�V_  �������8��� �f��?��&,~��ǵx� {����� >�%�k�F�Z0�)�^`�P���-r���IOAQD����n�� �&�\�h
t#Z� ��K��[���� T+��b�YOQ� ����;�p���5�". �S4��J& L�a��:� G������� Xĕ|�iޢ )�	���_ ��J�I�B���ۼ� �K )|�^Ɓ� 0�{�Z�� ��+K����5}P���@� ��]y�J�1�*�e�%���\�:���}�.���-���!_#�@p��" r�bN(�� ͨǀ�/�W EO�?�Q� y1�l#�Ǐa �),�	h unYC���H� ���Z|\ �-�4�JQ �b�����H.f$G;�AS����͓<;�<}�o��V�ёX'#��� W�]����f� �E��Q��a �z6%���F������&t`
 �Q2�>�'� �@J�u��Y����� ܆� O�� M�t�B��E w�(���#\�P P���W�2 y�i�|�'td�u�`�! �*�;��� ]�[鿰 ��.����|[ ڒ4V�6�zs� EH�mK�� ���,��� ECL�?g�A {�V
(׾ ۦ0H�^�X ��tN߬�U��>�&�� ��)� � �I�J��=c:@�1���l�eRPL'��t�����¸�%0| �	�}��z| ذ��AD 3�@�� _�&�Ք� �cl�υ�����ǎ�b�[A) ��3i�z� �a�Y��g��������� Hɮ���
����ؕ��0 �/ѸX| Z1̀�7� �	0!P�v� �\�Y%������Q W���'L�}�z ��:��+ �!�Ӳ�Pf@���/�8K�$C���'� ����E�� N���x� �[����} �Y�V �]
|Љ׷ ��쿹8_2 Ͷ�Б�{� ��#� �7� JWT���� �����^�c �B��$��� U�F���
��5��
��π�X؁�` 0���X)�6߮F9�Z� =��-��E\��;/'{Щ ��7� J� ��qE�0� }������ �$<���� (� �� ��AƳ�&��@*�Q �D�� Y���9��x ��L��X�J ��3�!� K��'~J8�a����S��|� ���[�K�����	��%" )�U���p��b΀��`��[ V�a���O ���%�N�J�`�� ��D����:�֓ �TR j�w�y�u�\!z �7�tD�1h<C�����A���?Nj�& :�d�R1 ��{����k,����bJ�S
 �-���? \�~׻_`�tr�H�^Z �~[h�D� W����x ������%�!�do��8p �Q?�/��A�� ���7 ���9ZG,�� �	�tyx �@ `�P0 �ځ�!ʋ� �k'g�\pa <���3��?�b�o�Kj%f�� �V�I��� 	2X��k/�E���Zs^��)�_u��RU vTP׍[�� q��.�;�}43�� 2�!Ȉ�Yh������ Q/�0+�Y �K�����2c���-���^�q��4$&�l /f��3��^�������P�H	G)J��R\@�W "�Zч��<�B +Q�C]V�M�k�	:�Ȭ� !m�f���  e��)U� �q��]
 ���P�8{?� ú����� ��QA��{ ߸Jɀ��N@��)���9����C*© Ű���^cR{����) �_���m � h��e�� 	ǌ�7� ������U���͇�Ľ� �v��у� w!9�b� A�v�0m1H ӻ�(���<�_��A�
p�$ &�+�1�9 ��Ղ4�kz �/���� �tW2d�? �n����=� �zTi�G +�o�� N�LSQ�ā�f{�i �c��� �1��4n�� !T�� *�
�� ��1�V�9�������7� ��1�M;*$��� W\��+�R
i/K�c��@1�a����n���;���֝<�� �
�yZ3��: Χ' �ԤD ���G�hNCq� p���e­^�%d����QH��y��ꇩ] ���2�w?0J���L``��#��&s �X����^6�fY�Z� �S�oV�� '��Ue�i} ?7�X�w�� h�Tz�P��`��	Q2ѱ���d�d0����� R��1��l�<�I �]D���� RT~	.)�� ��]�t�pW<T} �3
����ރ���P�okJ r^�	2�~D唲�2�hw���sy �W�
�%#<� u 0�.�3 +W#� c�U�2}r~:���8�[u�_� ������G cX\Y[Ӆ\���}�~��v��{쪑 �Oh�&��8��!N���uT �B�沟p\r���V�́�NS�B:pJ ��8���=��f�� E+#�%r� �Z�(�0�f����e<�3��!��9	�����B؇�P�pq�
L A{��_+�b ��ن���Z ������� [���Y #٫���JDS���hǸ�t� W^�´�� ��)�hR?Y��'�r; �0�u�a� �Lt��%O~w����� ���Ӱ3R% V��Jn�'}��Xj�`p$�� r[�h<;(�7� y���vX *��ս?�� ʵ��," !�`NM/��9󱀔9P� ���]h�_D�	�Ѻ���C�p�Ð>kj 
��Z�� �0`x8WP ��7� � ��@��\ �b9�^�<�f ,�Q�[�� �	I!���_��0�г�Y ^>[�-bRt )�醘� JP��քO�-&`��X��V>#��\�0����� j ���e�#��ER(�c- ����#"��H�� _���l�9� I�X&h;���+/�*�P�UA��(�{� �ቦ�C�@À��_� +�"��% X���{*�H�;�3`a�2�pu�V�����I� ��Ay#(K� v +��[��
e��3���b� �0ԓK%�� ]�麕I h�<��p�� �7Q 5��6 t�ڷ- IuȢ3�� ^����~-t������ |�$���̍Z�3�� �b� �N��s��n�TSR��F�0 '\鮟P ���"�嗎J&�G������ K>��w E1�i �N�(�+^��k ����v�/ ���Va���=�N����ހ�~OKf\��_e���I��ơ�u ��� j�U�q@���lo qߢ�J �׳nZ �WDVO���*�(-.k E�^& 3�Q#+ʖ 
�	��|����Z�Z_" &�*!�e ���k� LN�'V] l�&�ɮ� h|��[����iT���pذ� �4X���y ��Fb�[�� �$�ҭT�z��؀㒪�H��g��UN� \2�Z[YuW ֞����Q�^�� ��l�a ���/�K ���C�&XPR�v\8� �Z	Hԡ� -���k} CbZ:<�� 5|�8�{ �H ;o ��G� �Ԡ�X�
�h!8��P���L2� ���hvN?���� x�.P0	��X (- ��*�� ��V3UHO'hп����@��(� -[Z���� ~C&�)� �1}Y�S ���t	�
�� �Q,��N% �`�S�����O���.�
�9)���},�Š�k^���ڔՀ��h	�횜�bj1��#����W� ��0���s� �$3�P�%|tI)��*�~1�R�J�a��܇+ �Ȓ�������r��Z��@2��� ��V�� ��t��3�N�	e\���/����M �$�50�4� �����^ �U�@pʡ��:{&J0 �߁<>�}� �A7�Q��2[r��B;M�)��u R@���N�� �W_��<�s��~�X -��} �i��?��� *�hd#��� �^�ʕЄo����@�����E� c�ϟ0̛ 5��>��u <�$�U2� ��WpH�,K������hZ=X�� %$��H� ���A?oD �X������ q6{QnJ� �h ���&F{D��ix� �;Z!<�� @���f�	�� �~|n���� "��0�]�X �!_���j�΀�lB� �@!�Z� 8��M��= S&)�so����[	��8|w��^ ��e
�5�~��N0�@��4� �\�w<o�|��~����� 0� i�� 	N�`��Ә�<�����z�{41 �Q(i�߈ ~G	��� �u�=���)��89� lR��˜�_ �Zo�i�U~�@�yH�Z���p�	�9c/�t*��]���f�� ������הO2%�,�u` �?�$F�� P[���@�h7�1�A�`�j۽8%�I�B�[�I�>� ��aTp����6�g1j)� �_��fX6 .��	��wz�ܬ�,%}�^����0�+Z��H� �|�!�"-��� ���е�z ��h����H  ��I���#f�	�!ո��ZԨ=����XN���iL��Pk�� sx���{ ��"�L�] ��h<���~(�� ��ü���[��B�]���X4i���9 ~Q0�^9�����;�1 /�<P�y��g���!'7J ik��wp����~j�g$��$A�xE ����t� {�Pm�]w%�0V�?�����z1� k�K�ۯ����� �X���Y%\��/�`��o�K܀FJP4�	�� ��� ��3�Z�]� 'ԯx�{ ��;m�+q�s5�������� %͊��B#-|��Q�t����VA�� ��1�X�N !�D��J� ȽH��yp_X 9��� òE17v|!�Q� �.�a5 E�R#�ب9�°@úX���L��;�J� ��%��,�� �B�( ���3��� .���]�g0 �t�&|1� 3�ZC��� ?������� �v�%9g 
@��r�� Q�B	�a����@��]ȝ �$Np���[��, +&��( ��������ӗ@b+�`�1 ���g�؞	 �3-��N� �迻*� �^��S��b����z3�_ ^�p¹���Lq� �	fX�Sq�>� m(����!��	�'VRQZ@u�63a�!<�]��� �(U���t� �X�K��><���1�#��%���뾀�P�C���]5@�\QpPN��˘� ,����A`J+�Y����^�0�'�����e��+��� ���A��_| �Z�S��� ��>��:�) ^��X'h�H m��a��\O���Y����i
��9�y���`�% (�tE�_P���3�/����2�]9 ��\�� �-�p�QfP �Έ�t:�����ND�0�w� 3R�2<b8��BZ��������/_�P���5�� �#��}�oz ֦������ )4h���3+t�[#�Y��b J02��"�=��.�ض� #ߤ5�`�� <�H\�bK�=@�A+��0 � [
�ht?�xI #�价�J^V�����v�Xs� ��b�Ul� �`p�J�� �)�2��z̰Cx� ���Q��b����ޠ�O���v3���cB���*�9	��� ~�Zu�0�F���_y�3QlLҚ�N ��.�7�<�	��$Z�� `]�s2^@���r��hv0,�� �(�ᆩ��P~�=ւ��S�0�$��* /����� ~�,����h /��b�6\� @�*Q�ȷT ��W�>}ŀ��Z����X�a	�J(��b�� 	!Ѻ
� \��.�8X$�Vd��r�'�[ ���N��_�`fR�3' #�ѝ�к �*���-P��K�f� �g vZiU� ψ�h�K5 P;��:��� ѷ'�Y��� Z
�MXE� ��X�� ��m|bGi�P0�ݔ��D�P���Q���U�|\	� ����f ���mO��e ��^��Z>��z�J���	�!� #,��SV�]�7��R��`��� ����]� ?�YH�;i�E/� B����� �@w�Ŕ�q �p���#�>�?�. N�����B�Y�.1���0p� <�ɼ[� ����� ���ma���3��� @� ���}��85 B��-<i��/ �4,Z��x J��W���: �N���P#��J�b� �lmnL�:X�K��V��{��+�6 ��h~oP�( F��:�<� �k�4�?� ���F{�= �χb�lv$�9? X�x��^>g�0����3� ~A�)�Y*! �:�m�l� ?LsH�� (�.�r��� %\���:� '��)�U�| ���_"���<
K�9[~ 츒��R���O��7��F ���pk�� ��N�m\�����K�=�` S#�R��+��@�Z("ڍ\@�%�&�DP ���(ߐ� ����	� X�L%�T�� ��`4��S "�U��
� ��d!-(��)��@�0'�YrF1G_�� ?���׽&'ؖ�����
+����A ����G{�\� �eRi�JPh�* N��3�Q���� ?'���W	 )�5�d� 뼟�M]� iB���c�\��Hd,�`�
��τ;�O@��� ���|� ��o]�?�;#�Y�O��w �%"����%:�� �d޿q� ����������� V�ʹ�;{� ��o����$� ��V�� Y��@&Zj ��(�\0�� Μ�z��O� �X�p� �Tr�� �RS���.��5 A*�h0 )�"��Ƶ���&iQ@��� �O�%M �Y��)IX ��vB��L�x'i��j��۹����0@��|��@!�S�� ��"�Q(Z� ��0N��za�C� �я���<> ����0� )��m�f��� !�^��H `}U��� �[!��?E� T]�ەw�Z ��F�n�� rB �Xb�X��! �W��N a���m�3H �T�J��	Z�.�C�DɈ�� m��\i�Q�!��$7���0�u �q�5'��,���\�� ȉ�QĆ�n)C�O�� t���#�rw ����8�@F�㕳ڑ�	�`��8P� �yȄ�H+}�>%f .K�E���� D�	l�&)�^�� �Y� Z�0"O����� �͉�~��\5}K �n��X�{��z(����G�V�]���R1؏ZJ���[ $����+� ,� Ã�} ��3�" ,�.'�n� Xp�]+�� �Hb���\9�����'��[l ��@���,�	 ��<�Ď� �k��}� a�J��Xh�i{ Rw!��p��v�`e�2>1� �t��Z� �h7>�'�� �N	��)v]oX�9�R���we�Ss 3�}�G��ٸH ��[xk% ����h�Q>$���;�`��! �`K
�S�p>�Q��pn�� �h�c+1�8J ��K_F�� �I�sӆ. �*�vXE� �����8>Ze ����5 ��%g��	<���7ZaO���b���� ��d�J�@�� �;��k ��� B���{�Y�����!��,�* 8�
`� ��OQ,�����s
-��`��b���k��9 �VQ��%{ �k���� �2��c�R D$fjI� 1������P��H�:̀�� �V�� �ս���H [���C�� �9@���?� ���[]1o� ����ߍ� �蠝!�u |����� 9�_1e��g N��t�U a�OF����]-� W�� %k8I����_n��<�#��� \ �ah�	�F� $ZSC8覸� �0�Y	(�!&ݚ� �^��.�Q� �TY:(e��,�" �\��0g L���*��� �Ӄ��2X� �h�W� x H��Y)���D�s����Yl{,�lC���	� ��rP����;� �� �Q!�o��.�~�3���[��w����1������	���5a 6y���� K�h`[ ����˽� ,��UZhM �1�K(&x�>w�����I��i� &�����k�T~ �W2�����,�Z �ͦ3� ��	O����� �EHc�K." ���>() �&˨^�WE f�w�BƋ�v� {ia�q�k����#>� ��� g<����^!
H$C� ӹ�g
��ipz�XQh`�2�k�\� /�<}�Yi `0��g�V ]��.� /��c������ ��T����*{�w@)�н� b���z�]O k.��BPUuY�%RM^��hg �����Z �����!�� �p(�K��{�/˄'��5[א���C�v�� Q����� ��(��3�9  �)���6x� ����#�� ��PQ$>�� ��i%h4 (���Ns� �Ļ��"�AϞ���+�f� ��5��㹚=2Y| �����G�� �ht0.�FD��/�_B�q�x`����f[���� I�XS#���ǀ��R�u L�-)�D�Z ��}���"���K��鍆N ��Z(��-! ��˕I�: 	g�Z���R��_+�Cz ����o*=�V�@�������g�MD�w�A���8 � ���\�I� 	h�~'��X�� ��\*%v ��!@W�#' 1�Q��x�y �0��w���{-��Ξ��|J�̌�AHn�p?#�R��/&*�B�2�\[U�4�8�"  �Sv�1h,�D���1[ ��� ���R�' F�A�)�� �� ��X| �ZV0;:�����%.�zpo�|D['#ʠ�J�. T٬�6+�V (�Ύ�P��.��'�X����?��) T^נ�.\] �+���� ��*��8!>���4��tu.�$���a��c)>�;�ې ����
� �g%��fS�H��x	��  C3��e ��%����� i���X�P��`�nqKs8��Y����[�px(D�"�ɀ��oT �,�d���Hac���puI \�:�h�6$�{ �)���# [��9���t��X/dw"���� �}Z ����(�hE�4���́���v��+�_��	�!�Z�� �3@XW*� ䷭�[�:I	���YN ���,�E}�d�
�� ���-� ?��So� K�VW��OBs����_���KX�6hN�+���e�(;����
�'�^ 3������\�p �SR����� )\/W��V� dOY3E��J���!�#�]� Y��B��n����@D�� G��6���19`� �YJ�0����{𱄀+�\ ���_Ķ�&ݩ������ (b�Շ}~^�� �@�ہͥG��� � (�oeh���[>Ex����k��к ���QC82J�GK�dS������.A���Z ����) ��o�`���K�����d�;1 @��o��Mqc=G3�	�-
 �$Q���$��N; Ձ:j��> ��hb�� _���N�Y;^��+�ٯ 	!݄J) �_��ؐ�X�� ����A�`)�������f�� ����J^c��\��;ˈ /(`b�΂� @�Ҵ)����!�t�["B,u-_��C��8c� �{��p�?XU�	���J� �Yw���!}� '��KF��k r-�w�&DR�B3��h}I� d;�K[V� 	F�P�J�� m�/ׂ[	 �Y���b�7O'�g­��*�&0� e�F�qn��Θ� ����u V������ (�^�=
�h }A��� j��U0�[�� ����]� ѐ#"�L ��N��; W���X, ����[� �Ӻ-��> �X�Uǆ94 ���C��� �Z��p�Y�]`����� ��Xe�� [
����� n|6���R~ %�V��鄏  I�Mv~>��� �
(�>%������� ��ګ�-���2��]^0�� 
��Ϋ��	X�ܰ�2��B��aG����  ���`�/ d�񁉒�" �H���{��Q�w���)ʀ8��Y�/��h�@1�}:AUc�����YZ������ i�O���!� �����n�B���&֠ �Kh���,՘��D���Z��=���N��b  ��<��2�T	R_����� �`X�
��:�P��� ��B���#�@�3��� Z�I�Y]H��h��o[ ��8@Z*� R\�"%�� X� �-#� �B�Y�@z����":x}	���e�K 7�u�乽'x� ɵ*�_5�`a!K���C��`�h�i Uy�2��� f��\_�&BYI��x^��, �-}!)< ��ji^�G&~e|�B��fF	_���T������ ѸR�e& 	��Q��;���ZW���= ��^,E[3�Y�
r��1�00V#����U�܇7��t��9.�y�_�ѿ��)�3ھـ�AB�l���
't�r ���W���y�=VO�:��)����h�t��A�>� �$�b�_�J�F �	�L �2mx�Z�� �Ȇ�~�A ��t?�K����|��X��}o��v.+ ���'V )�c�ҥ�-�9���� ����� N0�!Q�K�޿�� ~�b�h �N���'Ԯ ���ˆ,5_�	�`O���r�
`�8ޝ$^
 �mZ1�`[!ͽ|�Y�Ä� &, h4ᒇ�K0fyz[_� �S3����<����@( ����$=� ���g�,		�_؅y!P��b���N����H�0 ��
C鏣��,��f �j[(�R0��z���ղ����� A-�6X�� 	9=��	�h�w����x�� �g��� ���i:X�:	�'1	� 0��� �U���/�.� ����W(�>�V�V� n8�%�b ����I��uT ν0�n��@ F��d~"�D+�#���9�L��G�Z�LX��$2I;�!��</��\*��>� r��Q�	�S ��X��^+��p� J��UC� �@
�v� ��0�	)�. �y��V}c~�����;Æ�ĕ�?,@�c�>��%�@��iً����Z���A��} zV��Y��y #˛$��Wp־J R��NFy�&�I�MY@z��u"�Am�>a��`@ �滨 �r;�.l렠(�2 \-�7u����x爡���(iZ� �|���	�{< źpu� j�H3&ְ� �c �	�<�"��q-�\2 ��%6��O ��o"�h$Q }��+0��� ��u���R��k���,� ���^�?` A������C @p���0 �>!� �C㴆�ENp9 S �P�-ɪ �eکX�" ��!h�2�Gr���-�u� �P+ٸ�JB��땒�_�+�H>� �k��Xh5 ��IH���'?���2�,bd��@��xAZ=XVT��H`�~ 9"�@��� *�nь� �ȭy!b��}� Ua��)+�; Zż��C���� ��3��Uҁnd��-(+����_.��i0�s| �0˻�%��������T�G� D	�x��[ A�E�R�2 �H���� I��R� ��0���#} ��O-_�8 ���!^�� kS���x��{ f)����[ �
�ק�P*ԗ� m��+�J���T��ŵr� ��ӫ4c ����b�n����&hKJ? ��a��P�/����!���� زh'� Kg�ӯ�� ��"�R�Hu�w ^pOb���P�Y�����D( ��U���p� "�ƀ0��+��F�i���$��L��w8�H� <a0^P"~ V	��#����`^��'�&W�, ZNM���aS:ݻB|��1��� Έ'"�� E����7-P��3� �1݋?�= 8��h��[��� ��S�� ~�{	�Y�\ka+ߨ9T ��H�;�� $[Ջ5av!9��@�� %[����H�� 2���`�P
�+Z7� �O�m� ;�t��� !����Q.� g=��	�Pt ���1�2�ru� ���h��0 ŷ9[��P��(}����81�� �'������� :�q	�m� ��6�!�� Wb����Z� ��8���< hzӅ	W"�L�� �@�!�s ;�2hfP �?雗X JV��0�C ���,�^c (%�j2� ���	�h�(w��8L��[�S���A�_ �q*���@�L{�e	�� K7͆6 4�Ȭqۓ ��S��ܗN_�j��f���D�! Kٿ�6��� Q]��S�����^��6�_u�2��W4���� ��[e�B�ZK�Sɬ�h�R �����(ݺ;�/ [`��&�����!R  �- \��)Рq Z��@L�M� P���:+� J�ւ�{� ]FO��^$�.�� ��I�ɘ�ϸU��;���]R�
 ��i	��L��YD�o�렆^� ���C�����h� �b���,EL�� ������l C��^
�RT�PZp�Q� ����jIC� `��O
���W[�� $�)��� 
�� 찘3 Ϳ/�Q'j� ��Z�($ ��ԝ�a�K T��VCAW��N� �E��7 a�<v	�;�x�W?�z�� %_P��6� �t��B��� p�h`eV*��2�@� w��� �^��!�{R �38�.� �ng��փ� ���ɧ� �A_ǹL� �h�Ȼ��3�= V �8��� @Ȏ���#K,�y`�� "��c��N ��[������ ^T���B�W �pt�E`���
���-� ��$2ƿ�_��@6�% ԑ5���� k�n��W G1���+$L�u5����	�[����\�'��@�ɾ_� h�o(���j2� �_�J� ���Ƃ���X046 ��y�D ᯙ�?��K��N�'�\qI|���T̷/��2�%: W�S�[LV��� ���T����:K�a� �P�Y^58)�O����kG�B�<wd� �+��1�|�D�a!/�E ��	R�Fi<v� NH���׏� ��荜 ��iN���D ��[�������drL�� �6��0�1��Y��|�F�` �v:�L%D �	<"�,@#z��!�m+3<p"�}i���ї �z����>�k ]0"�����_T'�P���2t���@bч0��.C�� �ÁP 
��{<�@ 5h�$�}� Z����0ɹA�(�;�w#Ћ 4eY��� ��u���:��	�x�1;�+� {�j�/Xk'3� �}�;!�"���)�躖,����z�-�rF��%���� �as !�>�j�אп{ݭ0�i�FP�� ��0ω��� �;U�!�R 2�0���� �B\}��Q�� {"`�j g�7�i�| 8�{���� 瀞1��^��J ����~}� 	hy��1�$xm� 8�A ,��f<<�×�������$��w 4�/i,;t� ��{���� )�B���0 �9ϋڀEX��Y}�y�s&�+�� ox-�C �	�]`X:/s=�K���x\p�f�'}�pA0� Z��k� ���'���	�P� �L1���s��Y��� \��b���u'Wס�B� ��)�L��>丣]�'^0�&�&X  ���� ~ZI$?���%&��uXzs� n-
}"<u �ע��rx�@�#�/����+�ǔ�(��i%S[�l������	�8҄ ���� ��
+�n_����U�$Q����B� ��w�4$z��'���O��".�ܦ,� G���� >�cL�O(��H�؇X�< U����� ��[��,TK� �"��}��lY�0���B �\��W�('�8�ހK��P  b�X)�	 �2y��fP �d0:��@�:|��7��]/�@�7�� d ���������G%S�L�rU V�%���2 ݉�^�~\�.S���cfЉP�ZU����`v9 ܉�C<M�ƃ�H	��qH�� ��DB��}v� ��]���J�A� .���N\와MH�"&�:��uf��J���Š�4z ��Q�{&��
3�[P� �.0��)}X*#(���������� Ȁ3[���ep B�鍐��T ��(�!^n��z(� \���� ���-d�oP 뷸�(е`���؊{�'�D�U �Fra�A�>`��G�U �n����i./� SQ�5��	� HP��p$ \���K� �����,/s��З� �%|i�|	 H��T �0�K��E� �S��fa9��� .���F�` ���$�ZK@��@���
� �:�?zu � (�S�� ��
���> �=wA�� 9;ջ��~D�T�\$���S ���P>�?[ ���O)N�� �%Sݲ�}q �-�9/dN�x� ��p�%ZSF ͘���j��� ����5 �T��\�J:P� *�B�t 8h$;9�n	�1�)����!�w� =^�uZ�� 4��Yg�� Miҭ-��'u�heK,3 ��C��|�'@�[`����ŏ����ݘ��� �!���t��W#��p�71�:� ����{� ����^��!��p�VC�<�_�x��0�gN�(�� ̹h-9# �_�DN� �W��I�'� ȤbE���������	] J"T)��� �h�v��^�ׁ<�˼��Dd	��Հ\���} �C��>��8���NH� �T� V	��f��� ��Q��!�oB����~X-�7p� �|
�I�� �䖁���npW 2�V���P���<�pqe��G���(6�� 	�"�U��\�! �X�BOZ�'�P�\/bʎ�zXd� ����΀R Ϻ uA.�w ����� �
0�� qp+�w@� ķcM��u�� \�B@�k� �h�NFU�� �͐,�^:�`�'�[0� 5���	 ���ܕ���E�a�YA�f3z $���P� C
�	S��4�p��8(� ��f[��J�$�-vp%� cK�R�!�z� @\�%�� E"�Ճ>HX��
 ݡ���` =�K�0B��[!����N �QW���B� ��K��1�{�������;��RCp�	�=�X�U�;�! ��Qs`	uI��~�M7Uء� .|��y%��;Ȁ����F' 1�?_ �*�<�`��8إ�7��V��s!��X��X� Yl��X�FḧKɎ!�J��\�>z������� �Q��tm�� �Kh�{*� ��ڳ��X1� [	Y�k�T .��`��sZ��6*��	{������_�D b��1�&)���� C�(��[�� :���
+ѹ8��h_ax��� ��~�X�rQR�@�+��P^\����)��}�	�~�0�e����^��m�"��\q�R0� %��� ʳ����T ��JA�#� ��5��D 7�ξ�o�� �xL��'��<� &�O9h���½����P4}�>=�ǅ���	�WQ�� �'�LX�\� %&�����^ h�U��"- ڸ�  $1�mt� �c�S"ԗM��2��鰑���1ǒ�"�,��LV%U O��� ���S�� XIT���	�� ��P���W��^��(�3` Y��F��kVT���@B�s �wP�h�E~���+�L��mS �z�	�y< O�_�J ���AI$yP���ﳁ��z�Z�@��� .��{XPN³� ��Hu� �{��d�w�� Z���jL ���*kY�� ����a� ��$�	�Ġ �'�}~�f�e��t	H޽�6�:�o �K�I�����3u�q��P0�V��;�S��K�^us��R ��-hޫ�ڂ�9���<% �?��o0Z rH�O��� ���楂�dQ�L#�v�О ��3Z[�] t��< �f��'�.�	C �D
�h #��+*8{ ��n�Z	� e}�A`
�GXՂ�*@wƺ� �p'�<2�<;�:	b���R1���5F�I��_�>�Hഋ1 ��~��˔o �؞aN@ĺ ����_
"5� ZB��I��R ��XS{C��@rc� E� ���� �������� L��֟B�&�����l�3�" ������JsO �0����1 ���[�:&@ ��OJ�M�0�� P�� $ek4,�L�o��V�� �bh�&}��Q �U�� []+iˬx� '�����2��h@|��]0�( �9w ��^ �a�~B��������hΎ.��t���>Թs �a!�)k�������4��R .F,	�� �1�R�`.J$��y^�)�����0
� ��~'���q�[g�`�u��& 5��\�F��>g��& Q�aȜ0<�y�Z/ �����7���bm-��[� ��1i���I !(�O��� ���R��l MI�J�+ �p���\&��� ��OP��� �-0ɘ��#|X N�:�xЪ �������-O� 5��� /����1�>�����*�V� �����2!Q ׄ�h�R� �Z�J��� ��9� ��`�]! ���s_�� ��R�@'���� �<��브'y��(0��� S���d��<t� !�-8;�
 X$c,�&P�<Ձ�~����� GS�H�=� .%�A��� ���k� ��殧��  :�`[J9|
o����}����q׺r���'4 s�[؅��Vz��:
_��� �C�2� �Z�% ��j [�a���.�$����@�b��2�����w"�\�h��p�*S8�X����Sl� ���u#����� ׸C
��b
|Ȃ�� ╠�+� ,�����{�����s�3若�\ԿD����~��@q9�� I %B�:u� E��{�!� h�z0(��X��K��ԃ����݇{`'���7XZ�
� �k]�ds� _�Q���� G���x(J \��e�!�j {�s�h��� �8��n"^��F �_�!#�/�;f�1{%6�@��᯷K P�C���� *Aڇ�� ��X�� *>��n)O�$� ��X��
א�i� 6��#} ̴��	�+�����ˀ�B<�� 5�'�) ��+(�� ��-1Z�0 b2��I�J� ��,�e��MV����[�� I�!��e� *����]&u��K+��V��3�5Ы�(�6�M�NS
�L ��d�)���"���h# ��E�Y ��I��� ���tQ'�b�ֿµ�| �C�%�B ��R�fD�� �za��Q</ 8X�h?J� ���4>13�q�Z�����z'B+�P����� J�	���;� �3������9ȒP�҄�q�m�^�%�?@��-4 ������ �_����f z���^��l |b����J W@΁�01B*ZY���%w 9g��/c ����SV12Z_X�d��}�@FG5 � �z�a�� 1N*��� �Ѝ�`�� ��Rs!�n0�`���O^�'2���<�bg������ ��y }�!��cאpHt �m�^	{�p	ݪ<� �`�i� t�9}��v �f��[X���	��T� ���8�!s� �๱Y5�}]J+`� �����z'V�_�4[� $�?����U�����H�� 1��S,] 'P/�qw�8����� �����Q�\�ځ���:� $V�ݾIox`��^���O�@΋(�X �QU�. 81؉���;]� 2܁�%�&�揻���R�P�	�I�^��}�?W��>S��1 �ᔉߋ$(��s=!��<��0�Q
�B�D8� �bB���2
�4$Z-@Y+�Q���gA0���2)��ѳ�����0�3���X`9���h>�R�Q��!�Y����&��j@h��*��5� ����q�l|QA	 �F��[�Xэz>��W&
�v$Q����9�k�
���R���B�Qй?E���y�����	#�>��sI�����K�3��>�> 8�����?FRC�x���~
���]Sl�^��c�[I(�bE���;�t)F�NT�!��@-������v�A��FX�@�Dz�>@�3t<���I��,�nT���7\��R`�t�	Xh�&�d�B8��]N��U��a`�`�E�G3�u�H�>E�X��}�P�|U���E��+�6� @,	�
����4"3Ӊf.�{�>�*�%!a��
�������wT���5�&�+�`�1����d`�d�I�X>���!�1���s`.w801��<�u��t�G7 �p;��R�@��0iaڀ����)4F`	��k�7i�A�D� >O���)f*t�"$[7��b����h�9���	�Y�4��� G,���:�+��t�$6�K�Cwu��q!�J����#�X�X;�y���:�o�7?�Є�����a���� �s�%]9[`*�w�\4$� �¡�o� �^�~����YR N%��{䆽?�w>J��@u邲���R�%�թ8_�L�\��>[=���)�(@)��mi� �����{y�L=	$Y�� �٫���8� ߮�\�}�(T��퀬q��ϡ| Mj������$��Q7 d&8v�kIJC����q��!�Ha����A�z�p� �'��ާx�x�,����蹬}�(Qܘ�a�͞���9'� 航�P r�I�fy�.a�@���{>%��۲���i6 N�e�����1�r�/�W� �]��p� ��$	��� P@=1��\�$Ŷ �9�)�X:�	y  �hA�<����3w �&iy:�e -��ISg�:'� �D5��T;+&�d*�I��] �٪o��"� �j�&� 1�92���� ����r��3��+�L��Z�>��2$ ��pxqޚ'��;�_� ��%~?����qzFш�0TO�s8����c� h�+�V�� *���Av��������k�� 2�%����M ��Y�V�!�� �9n�tM�@�@|� ~"%�^G�Ҳ����{Ƒ� u�3�����  ~MHR�9%��� ���L�'Gp�C�}� g6���?��<l� ��y��tE 2%��>���{*����؃u�ت;�$�#@�a���%w�?��L8Ѫ�A&�����a>�0$���Ǌ�E������/#K���t��k�W� �!a�g�E&.��, ��@����I���O�i� ���%�]��&$S��Q�t+���~����h;�&� �r�s�%@�� *"�����S ��Y$5m�% 3A�	�ڹ�� �U�����!+o�&6���à�@ �����A�Y:��9@t�'K�	5�_ 
���*�!Og� Rz	�X��̪:��qB�8���A������F�Z��0���-�d�L�� �n���?��� C�0�ߋ��VNӀR�� �{����r^>�k�ES�);�'	�8�
����A*�g��Q0��>�ɼl���k�L`\x���� ����٬�0v-�zq� ���"�a�&-�d����Íiw%�0����ۂ:}6��$�< ��@��f��, ;�%���0b �(��Iyظ��M_�	� p�����>�;��C��g�b��I����8��%�`��0u���ơ��8���3���|j��ȏ�) 6�����H+ <e_*�}L65�Xp wʜ��A
��L-����y���V���H����9�����g<���b��˛&֎�������%h!�'� fp���fk�%�@ 0�E^�>����,J&�����rc �E�?%I\�x]����B ��:N��Du����;R'�@l.� Q�o��� �*��O!� �7"�m�%� ��F���Y3��$`\h� ��2��|�a -N��sl6[{� �7���,�N&	�$�8���& ��w~��v2��s����EO���I&�S��Q���p���Uw��^Y��1*�Q�m��{
�J�Z� �D�	�}�X��������������x��� 9j|�0UӒ%K�r
��Xehu���*������%�ة�v� ,j�1> �����݇���=�M����%�����j�@��Lk�>�H�� �u�����t��`�7:M�X��B�/=`��X�� �od[�̔�`:���7�h���eg9΂.@<ZI��B�|�c��/5�Y�J2��h:��� $E��*��t�=�`�M�?���&!�[g�J���@��	}.k�B�)T�`؅N�%��$�n�HI�������␯�F�;A��_C�Ԩ�L&��o�qC����
:���&y�p \$�F)A(���2�����X9���N`}�eHd�|t �J���)��ie=���C �%P�����C;,�HE)��U�i�~���&'�L����A�Ed,�Į_ɀ�0�(��� �&�������.�� ĶUEg�v$�ԁ�!p�� �1�l��uhpF>�6�+,P��yJ�=p e�֪h�� �k��Nv�%����A��pS�?:��H@��%�Z�}� �E�X�(4�L$��Kz@�S�9&k� 1T@��R�.����G����Q���P2�%P{�� ѱ�	�����pӉrS%EH�D��`�����I	J��߀����~.�'�����:��D�8)��1� ��O���15�m�� ��,�V��%/�b\��&]��O� %�ک"+.:D�!����L� �H�&��Pگ�j������g[J�����0�똜vKR��&8O0S���U��P�W%���v�`��,�Ⲻ���f���ل��(i�����ݥ@���?f��ڏ�Ru���)�p6@�� o����K$~�t��`���� �<�\����I�p��)$	З��q�����O'9 �Q0�a�%�n�5�"��u�1@���� 7�i��a��R	�h gO
j��Y� ��z橃|6�	����1p�!�`,����lu��@��;�$�bL���L
 ���nP�@�8���;J���蝩�&� d�O�� o���P�>�v� ]�%�D������f�"0�R +��Gő�P�n�II��L(N`�EfD��<9��q�`b*e��������Q��vڤ@Aj@�y��$�%�? ,�l;�� �&��|��u5A��7A��z� pSި1f6�T����¼�Q$&T L/N�{ ���;��R,Jpt��A �HNE�I2���B�r(�a��\�@�E���H�;0'� &j K��,�P�	o��u^�����$Q��иC !�<�+�r"쥶l�V(�$���x�;�i���Ř3d�8L��$1J)�/p ��s�?'<� �FV�v7�%N�`�6��l�@0� CgF-���� �<�X~(����v	�%�kA�&0���.e�X*e�� �ة>�^���r�ପa��� 0%_:W�XM��ź�����L.�KW��h���ː�8@�6xF�����7�ph�����&�O�
5�N��Q��H� DX��Y�e���`yx:&D�0��9�g��{�����O��C�ͣt�E����*���j�H����pB$���G�>{:� ��ST(ti�P ]��gD$;+ ���r���� k�}�
%���*���9aE �Qc���Y�m������fx�� ��a��~�%$�2<�ۇw�\��Z T#����� o �Ja5������Y�%� �w�S��z J}��<�� ���R�ZK�_��<���� �!	%�~EҳG�]$��e���W,� �Q��>�bX��(π �V)�1�/aZ^c� !���F̓�� `��q		����8�|0��~5 �>Twe�3ǚh}�} h5��xU�s ��V��P���cl�!��d���x0R� ��+�* ����Le��W~�;�$��8�ަ.���D�X��N���d�����|��p��4�X��`<.�7����>��P��)� lUq�z	�i���*��Y$��@����bC �N�9Wd��L���c����%\E�	L���7���������( .Gz���s��L�S����,������A�����+��`��f%����x�� A��x���͘�,���}/ D�<�X ̪�;�$��� �s��\j�&5� ��⻩�V�,%��i�Ϲ���<=p`2L�c���,�� ab!��\��&ج �O2�'P$��@����%t�V���<ߠ�.亸$联��[1�`c;>,�S��kl�ʯ� ����1T�� 
	(�}Z$�ah������e�6A�? �#��>�gy�O��Iʟ�$���Cp�h#�E����o��@;��U����`�-�Q��<�� �T!��� �Ū'+��0 �h�!��	U 8�(��O��q�3�B��� 8����W���|�S3�:��p�&� 9Ez�% ѮT�d�x��Mȵ�ɠ@l 4xE�4a\�=T��9(zy� �%��)B�&�"�Zar��a�j�~ު����'l����Ϩ( H�Y��� ���犖 ��%����.u* ����tt ���kO�oF~�%�I>�P�l6u��}Ut��\͘ %�~n���z��ݢ��4`,��� �B����� *����Y<�݂�����Ԁ���	u��Xx��˶[�)���'�3�O:�i}�b,�qFҹ���?1@����W� �2�%BL�� F��6fd�s���G l��"@�����$��.��v(+��:���3�HXЏ ���͆��pg�����@�~�km'��zZ��:�7���&� ��-Q$�� w������ԯeF0`,Z��њ0����R@��-^1�1�$N�;�� 2���1p�\ו&4`oi� t��T��]�� ���%J��zK��p�@�ԋu�+��{�πt/��w��
&�|�r��� �c�`(�5�ƪ=�8"�xX����� ��(H��ԥ�h��$����7���@��+��.��8��xXK�Ъ ��%�k����1:�D�禈��?NB�������@��V��� 7ub�>;'� <ꂔ8;�k�`D��F�E e.�l�&����TJg�����5�P�
دH� !<�>���W����т .�\_�Bl��
'`��P�v[&���$���p(]	;�'����k���y	p�� Y]��� 	�G,��h �7%��V	+k��3�(�ox�� ��-"�� ��Y�
��<y�^�c� ���8-�����k���~�T�j� ��%	��9��3�]1��p�+��� �E��p���5ܠ!jJ����u��tQ S�#�kL }�-���	=�̺��0L�q��E7�Dp{ �yeN�%�(R#���r���D$�0�������HY�?�bU,Ű��;�1BP���V����k��^+&o�?�ð]5�Ơβ/^��0��]A�;�]��A��	 �x)�Q@@8���04!)�uu�DL� ���Ҹ%�k���}`�53MS3����Գ���']$�ㅁ�a�1������E� K������Q)�W��O[� ��up�h��8I'�����D	L ]�jFW�� ��[��H�� v��@�Sg{,(E� 9Q��Z�2��bc܀�6T �M���:���S�G���&� W�+�Q�� 	�n�\?�O���B��J<|H )s��$=���Ƭ�xv��R�� %[�k\��u��"x��P����#v�iR�w�ݨO�@i�"d�9�F\z�����7���� ^|@0)y� <'J��D�;��������*���0�~�X�ZĤI��]Tn�SL6X���YWw�� a5�SV�] %�^E�[ �t���pÂ ]OȠGE�Y�^�_T��8��è�jT:�s�U �Y�d�]�� �_�S� %��rƿ�u��Nq
9���h≚�٦O8߰D�[]�}����j�@��,� �(6^AvØJ�[�~$�G�Y�y��,�5�! �ш�Ȕ0>f}��Y�"z�q%C�@�$^���@�
Y��qx��\�Xkw�;�`�P�s�L��"y���=``�(�3��
&2w%�jWH�֐&��r7z���/���%>��	�Q1���w��}
��q�R��hza�X.f�}�d袈7J��U~���Ai*�t�oݱ�/Y6��e)@2�y��P�a\C	 Hz�.Y0���㦌E!��3VѨ�|2�&�ԙ-q�D)�3IZQPꠛ���$[�dU����@屨��H�Ȯ��F:��(E�HfV*��,3��X�\@�݄)/y�, Şr}F(E�
�4f�gՈ�U��g�Z
����2��%.s�FF�Y�U������!��W��'X��D�+�رt\�a_P'���6S7��Qz�m���?�yj�j0�IX�פL2�,��5���ky0���q*��xe�Ȉ��(�DZ,%8��^ɪEp�|��M����Q<�x��y�p<���GN��G<Y�1Ṣ޺$� �W�n���`.�'�P� ���X��� �a"n/)eM$��L���A�
 k��6��	�c���{ΜX#>�y V״u$��O�H�fk�iy֋�(g.���t�!R���	�� 4r�P9�M $닫�� �u8�+�NS �>�I�ܭ �U�)���-ǲt`�1��T �k �.՝��P C26W�Z �u����&{0 >��
�i�N �ũ�\g��(PD�B���x< ²/ڛ Є#Ĺ!� ��|m���i������j������e� ����ݺ� i;�%V>2� ֥�fY�'>�w [�}��:���χMvڨX�}7_� 0Ebji:�*�]U����w��=T������-��9~� i�%�Sa �f�`�&� lV���ڔU������<	��k� `�*���\Z���V�躚����I+Bi��f]�����_(������9{ $&�W3�� ,��I�{���R"��͞w�a$ �7h,�� ���ѾŦ`��� E��u�0"VQ�._E ��jh���u�P���K�A���,`�і-���%G_��F�R���d��I� _�VU�f�b! �oy�4hQ "����^��`-��W�`m�=� �x�n���j��5K����k��yg� ��y�k Č�7Owc �s�*al�U0�����< j��FR\�m���P��?�K�A�!���ty up��T6� �rF���N��E^pcU̴�]�$�3�
���O6J#Y�����/��ǧ�R��DxD_	 \p����T��n�{�7PAU�� ��,��� a%��Ƹ�3�g�9U�|s���8R���/[`@�]�̠:+�?F�a�1��Cd����]�8��2���	���� ����o�޶r����� � ]��D�g$�J��|�iRG�I�VrO�H$iT $K�Y�,P�Ի�/�TD�z��|�R��x�Sc=�e���q�Lm��h��l�"^A d�Z9&��e}t /jz�D�J"g����,� �ꂘ��H��#��\�k 䚍���� H���S)ӌ��<� v��a�*i@����� �ӜJN�$|�p? ���7	jwiT"�0�
�������!Q��$fH�4��0(�0#�)_�< �Ս�Wn= �uǛ$��0#[1���r ����q�
F���5�E�R(	\ X��Q( >vR��0��;TU�p �	Jτ_(whv@$� �����J���sS�� !�d�%]�� �߼�r�`P�_	׽��	����H�	rρ���ݘH,���B�	��ѹH�k (��EU�;��!�;c(�0x������]'ԩ�I@ ��O�P����0�j��Tٹߪ���Jf�Dی h�e�ʬ�@,��dK�@HA̢�D<�d�������G\D�c*�W0p*�:��Kݐ c�#2�h0��؆����@t�z���E����]�W��X�e4܂� .������Ҷ���j������{�z�D�t�n���:&�D��R���~@�xmV2�F�Eb�򷌀��{O󏩈��D|�2\���0|r(��M��j(�ZH�t�0|]0pщY�{\2�R/���y]#`X�ng�r���a)��s�@R�	����W�<UB\�dゐX �Ǐ$�Lw�9�b��i�a��B��O� `
:��bc��#W)B^��u��6J@�Q���,��u�9���:{+�iS��l k|-� ��]
Ezx�$A~XM�l\	0���nXX�TDzl���U?���,.=ɀ|�i[��t)	 �0jO$ӂ$|FO�|�_@hwMJ� DS�Z�  ��gÏYq�,�Հ0���~̀���{�P����E��:� R�FK��u������Z������Q�EI��x��t�l�(�>B� �t�W����uI�����E�����x�z�R��٬�����t ��
����X#�`l������ ��ӡ5��1��w7�Tb<R��H ��0 � �a�E���@����!-�{�,ݵ�@�w"#	4�yPܚ|��sh��<�@�٢� w���R��d�E*r�|��cU��m��@`W����Ndj��E�h��	_z��HLw��f@�a��@!�Pe�xb!�-/J�$�h�������PS������LzZ��#�P��)+ ���&�g�رd�H2�H�N(H�d�0�	\��|� r7[	j� �Q�FI��;B䞛|�bx��P�WaT���:b� �B��|\~)�VD���n�C+�qb�Ų4hx�Q�(t���u�h�&R���)ez	�2��v���(0q~�!R!��H���##> ��pz��*�m���zR���P���(ij1��Ԕ��v	C�Dq$rH�p"}D~k�lY$ZHg�X>eBi��������ɻV�R���D]eMJ��?�UZi���>ٵ��.���SjQUHѧ��_��kxw�@�����)�غ~j�e5H����dU����a��f"c��Z�8p�t}�DjKC��H	I�_�w 9�oMW��-��0!"y��8X�)I�7M�]����%�����Dew�ހ��Z��U�(^^��r���A0"�1Ow� ;�T�Vq
B��r����[* �οI��s u/�ٺc�{0�`Kԣ^��,���w� Sn�;��<�Z07<5,��}�:߀����r �������p^ vSis���"vD==�ET��5��(��
���ȅ�;�F��X�9�l
��/�*�yP�R<�ɀf`Q�L ��_TU�#�1��4����h�L�6�0�:c'�jY��(E7�g���� -� 8`_�%�m�u ,ĽJ�����u�2aih��?���� ��q%��}���\��(���`r0�v���} �� �2�e���w�J ji������Y�Z�͐D���{C��:(�Z���@���Y�x�}�1���Y�)��*}� �?�`G��P�!���!A���5�	��� �{\�f�� �ؙ�H����?&UG��+� ��=�Qh�q��)Bm"��\�J(WH�(h��!]�$}Fͥ2!��7�hD�F�1	(�e,�"ۈ���.@�;U�?^�$l��Y2�_����c�1ER�(Q zDZ�	%��� ܡ��
�W?���Q7�c��-�1���y`�i�QR?!ۤ0$�`H"Pd�%��m�¹�0�/K->L\�X@�[Dҗ8�oH0J����1��THLJPX}��ڂAI�*6C(@8\� �X���L Z\�
���`��q�H�jZ#J�؆�:k�g@ ��F��8�[\ڎ(0�!�<|��vxQ���E�rP�w���(�D�B��P�('�B��B�#�S��0����.����c�GP�A�	���z$7O�!q���a��c�b�!q�α�X�(N@g�xǸ��HZ��c��L�
�IH&��c�Ѡ���<2ݰ@� ��^P$]d���I�Sb�`I&$rĶ�(�+��w0������6 �@y:���?��] �,S�) U]~*�(���9t��
���.���DQ@T|8��6'@�;Q����){�0����:S�����x�;��`���[È;�p:��ɁNX8U� T_���?�:�,
�@���_�2��L8/3k��{�,�)@���k.�61*�1x��y�ϓ��G���-t;�	�u6��S̔1Tt`9�4k�k �:�(	��� ��6P�2�`@�1H¨�T	� �l�*U:�@dP7�t�5����h��*@0y��rքI��0@Ք�XX�P~]����B�Е@���1,|@;R0��S�:�`��� ��%�7~Xp����6���DS�:`$@~�9��8���=�@�x�%x�x?�>0���� �6��AR��C�(�x��.7����Q_!�6` ���@��;t���$��=�6S��5��,N��8x��|��x;�,z�`���:�*B��y���g�wM
���9W`܂�!��|(,T�I�	����PT����~. �7R�@i:x�A�� ��,�<�p@T�<4�6��+x�<������)IPP&qx#w�l�2���xOrx|������-�P`u�>R���<�d�A�U�@l��P �7��.�6 �=~�8�_ �;�
�Dx�<I�� �)S,�~�7z�9q��D�.	��(��G,�,P!�9U��~=PJp��W�hڤ4���B�;�4ḏ�xP�/4�{����݆����֋���<U��Pt�!S�+���s�0�f�'���8j_�����|�5D�(�`��U���^0D{ )O�,�>6y�����ĤG�ʌ���0��>�)67؈(�:���Q���G��PL&*|
�w� ,T̤�P
�S��ǅ`?x'��0�(8����DTX�����`�0U`�����5{AD,M�)d���RB p0��q�9�4����[��U�r#�$�u�pb�X�D�p7E��o�����0	�!�w��3�$�i]��"jZ1`�S�dHڝ ����trWM��@_l�`�jh� [�ɻ�.d ����;�7�N�s�Z��tv9:6���lpz��T� �a�s`�}�\ �e���:Pހ�D�T���8O2� "*��Q��42o���tzM��x�������@h��FK*�� �p�s	�� �O�N�:m����q �"k�8V^mE|�xl�r1
$��4璤We� �#'�i�A؎�
�"��HDa@��l'��h }. �����\��~�Ʊ��� #M��D�Y$�[�:��BT��k�l��hTBw�21�q�(��'i�`Fk��Z�#�|��}��䉨 %2^Ċg+��!�	:%ܝ h�|����jƈ�

������w!E�न4��!*�x"�� ;��pj̗� ���M�s���kt 0��1�M>ڕ �m`��SD<H;�u�C�@���/�;���4���!���vJ `�VG�XYdp��O���X=�����C"� ���M��t ~��R�P�� �.Ji#�� ץ�5����7��;<0��w��� �����<1? ����ʸ����`����D��'?T��`�!�<�� W� \�u(Q#`J�A�
���3� �O�aD������!p�ah)� X��<4 ��,/@�����x�|�nQ�yK�Y_ 'pa@�T��� �1���X�P�`-���$s�\��Z�F�����?� g�t�`�<���E�`ܵ30BS�+�4���6s���(�S ,U|�0��֭o�� �D?��s��	8��B) rg��RV� ���D~zp �v.Ꝡ(���:�G(��'�����!�l�	���:0����∤����φ<��0t��S�袤0���� bsL=?AhE�'��X�vus�|��6-q��lS�H��
�1i�����&��aI��3�Eu���^h�{�˭m1!'[p_E$@tF�Pq��0V蔓�)�䔇.['��d ?����ݜ T��Z!l��>8:���2k ��nH#0g�X�Gs(� Q��tqD
�@@��(��
s�[ǌ�A�`}]�	��k�& rh@��ڧ ��*���Y��J�H)�2���`�/�x\� '#XS P��o��>���� S*�%KT��� yW�nǱ_��6gN[�:$v ���E���C9����jܛ ����`�r����k e��&�T� �~�P�-D�G?�+pX�>�#H 7�5���	+|X�����B�(O�tFA���1����0k?:�`d�w&@��f�{�R,�C�� I(~�W����V��Q��i�����aJ��DFv �a)��n��Z���ϟ��!�0pP�&D�T0��
�ML�~Y�����M_c+09� ]�ף@�=��`��G+I�L� F�j�lZ&� ��Ib�x�n��`V!�PLg4PL�Y�`p}��~?�|. �!�8��"LC����Xt�?��6�x�L)pK@�݌�M�s�8-�MS@���k���Luh	´#܆� a�`�sȁ 맦b[>�iJ�1�`��)���$x�����?IK؃�� ģg �dc�І���? J��_�oFs��z�DQ�Y�	.�[��� j�W*�5��n/�p�@�b�@0��@�r�a+ M��)z�:�
w|�,x�9�q�3T\�:�Y�0 I$��(	����J0�B��w'�D�� :���SB�澝�M�G,:tB�a��HtJ�q� a^�X�D�+��8!�u 	'�J�]�%[/ ��!U/�Ȕ\$�G�	DM���3$x�p:�r�w��� ��T�x�>s��FX8qcc���0��wֳG�	 ��_9[�V���\��=�JѼ7tX� ��;PgG ���m�0�� �)�� �?d0�� /�&�X� ^v�S��*ƚSXXJ�|�����4�"`l��u�7`�hQ#�I����x�`�M�#st$*e &{�2�_����deoȌ	ݧw��Ԉ�S`+�8 �R���Y&���$�¹[�\Ȝ����J �l�|��~wJ� �x1����P��sT��~9�8��L��z�q'HD�w��@���:�1�0���Aa<b� �^P�V@ cR���9��E��n��D� �]��#ta�d�� j�~.����
Pe��[�#�8���!�i$<�X� $��p��;�-�?���OU��)�8o� �}.����5�<���)�@��sͧO�	P3h�:N�����G��kQ�T3�Фe�
��XPP0�x��S�`�1������w���U0 Z�\ .LD������v+Y1��ۺg����)�S�G$�P�E\���,�X�8P��� �'0��)���k�p�oeH�Ђ�w2#������И�����=�*0��4��,-��_��
�g��+@x�
.���l�	d��0^�����`j'
5�y6���Rc�@Pū�P0��=�1�"�eN�ؐ^m��p�?�h똈�`XH��-'_�$	�@�5���R$ �-�ɧݫ���u�Ȉ;2�A�K�����`� ~�}�L�x?��Ԁ��&��8��$WP����8�1�`�I�$68`����++ܤ�\!�/��F��X��J/ Z��s�- ��#�F����L��"	+lZ!��$!��3 `X��ϧ�s�2� }��Mq�zL�s�!�� �!�v��j�@������C������X�VW�P���!�N8���V�\U��GC�8"4�����Lc\�P�,� 
���)�;�����:q�񂁥� W��63�:�)���l���_��S���3�6 :�r���.� ��
@g��k?�F�[����j%Є��C� yza���{͎��Ȁ;�����˄�נּ_2<��H�:x# _�]��4^��u��H��ml��0Hs�����$�L"�?�� %���3������`L@B�1���J �ݞ0��Ƚ�B����h� �tF��u�b����4��'[���A�)xѓ� �gƝ�V�Y���y,g����<P��^��5���Xd�`O�|�P�ڔ�b. �p ����)ý,i{H�H��� P�§_:Q�����/���T�4�w�� �pd���kI[K�`0���V?�X]�
,�� �*8�Y�u���`X
[Y�L�>Ǒ,�lh@`���r<�>��'1��p�	<D\
H;���oh�I�
Bw���F��M�s|3�A+�M��L �s"�_�\��D�6;��h�3e'<���d�a�m0��%'O`4�ߐP`l�)����4M����� ���$�R�6��@��o��B l"�ZG8k�� ��*�� #ܦ��`8m��-����y����H�:G>�R�#�%g����c�������;�I�ľ�A	lahh���Ķ ĊAk+/X#������)�Cԏ����)�Xty8w[�v��	Gi`�W��S��Ѫ�rD5���H0)�&ɮ�E�D��y��ۇ��� N̄u�. #�ތT�Vh)
�P>$�@ѧA���L��D�)l���C��'7����;�
8Gv���9%�#�H2�"ÀˤB��C/@y�e�(T���8���\��{��3��P�Tc��� (:w\ �iҜ��.1	�����<C���ѨHX�e�����w&����IhS���]p1���G�oD2�q�� x�)�'�ݴ�C�Hw��3�P�|�	A�6�Yp�4�Ċ |sYQ���+����?h�|`Ϡ�����D��bڲ��<xVAD�H_�A���x��I�@`:��� \�aC%�Ζ o�a=0.Yq �Ԅ-�ST��� KMa'���X���p�����qK}E^�>ܹ�C
	�R4఺[�H�u�(��K�{��+�E��y��~�]�(�$T@��f���>G�,� ����j�;�fL�aI+H������ŗ��ڜu��G7�ɼ.B,�'kp #�?�Ɍ!�e��
u.E��Y�����lG�@�ػ����z�0>A�nw���T�#��aH��#4�t�a�� �YNI�ډ��[P2�(+���`�z���ɧ��(4Cd<� Y��v�`���0�J�L�_���!���\F�r�d7g��k�$�ta'xEdp�4$�3�!�ٙ /�"ر��!�r" ��WK�G���Y��;Dh��+t��K/B��[�YT�a�'����@��C��%��|J�@L���� ��;�G�נ$�B'�� !�@)��D`Tp|G���� �����͐>T���t_����s[�5�N "����U����	h��؞�L?)�O�bP�A��� K�(m�J��ls��� �tKw�bb,q�|y"1�(�t�� W�A�D@�L:l4 tK������At���Y�[��T��'�)�0������)�h�`gep�X�l��,�� ��Z ��� <`���mn��G㬢�0�� G�`�(���!�)���2�����8!3&\W(Fr�[sN�\ ��-N�! �Ӡq���f"�:(�U� ��`�@ -%>�,���PĖD�-��u���s���!q��C�2� ��^Q�{h)�Pȿ�B���_l� ��U;��a� px�ܨ���.Ro +4 C6{jk���` �n>R���A�� ��0� ��Ն�'����"���B���̘���� �C&��+d���%Wv99��7�L�G���v(�TԄ;��D���t�	\f�>�0�m|�bȻG����ʌ@�u�#¹����tӾ|����Q�d } T\!��%v�gȐH�\�d9� ����/��,Q�(`�F��9������X�\"|�ԁi7���`)��X�\�Rl� ��0p� w�Y�z� ����u�Ϲ��>�+�h K��)pR'���J�ox���G`!�*���OiK�����)���%`��,�3�F�_��#�Ȇ�I��'Jg���A�8�]��(Xش���Ӣ����T����+�,>���yǇ��0J4A�qk�ƈ|S X@LҸ����+�2&o�� �O�c �4�~L�� En%R��Ky$D�Da�we;,�#@/!x3B�j"HQ"�&>�`���O�$�U~�8Â��ɏ$�8N8�׈��E�����ʄpA�+ O�����Ƞw�#^2���Ѻ�{*ހ^�4����,��� j����$�t�)�S�+d��Ȉ��m�n/]@�R"��!P���G�D�`f���Yz�3�H8R��y |�F��軄c{����� ��~��p$�w`D�����?��
XP]��=д� �jE�4�,�������s���:w`@��2nJ(�@��R@ cZP-B�Т>V��/	�����"Ps��w ���5P� �f8K����QG$��ౢ�V�@U�� b��ֻ�D� ����z�'e����`ݕ��$_���0 {xc��
�� ��P�G�}e
��ď���R8 >D��y[%�Z�e.��� 0���I�G �|����l��B<�/c�|���.��H@8ꤓ!�I=4 /��:�^-������Tt���.^�BAث�p����� p����^FD7ƭ+LR��u.�)�J����� �����f&���/�����]�w�"u6	Z��ph�<D^��\ T����8mS/����qk���"��3Ǵh��Ys�n�����4���� ���T�|0�H��������u4���T!`|���3�M�sK��d,�M�)>0\d�$dg$�;�OҐp�Q��%C�����cv���,�0p�9�+��e��p@��}�V�!�K� )xB�vJo;�#� l;�I%� ��v=�':�xD���S���T1s�t F� ���*H l~5\%z2-���'x����[��ȹ��=�	�S>�h@;�C4:]�P����%����oJ�]�Ә���@A/,�nD]�H`�%�8���G5o 紽;��yK���7�(T��W�� 쟈�`[����Kq5�	H#p������F`�K(t��`�*"���� ��. T�g�)� A;_��C��Bꢌ\��1�Y���h g�PTԱ���Dr�@<lw��������o��1!.�)`�k����H���� �^PE�Iw���TYG4N5Y�׼�x ݦ�i��� ��ŕ��	 �h��IS'n�`лX%�q"���Al����i�ہ�����~QCj���	�/[���%L~ 4>��	���L��3P��rH [��O�x]�k'	��Д�)�Y?�t!\��1� '<3��HX��G�tR����=V�6h�
�]H<K�U�D�x a�.V��w��P��Ы����	!	x�/3��4�_���+��^�'�]H)�2%�P�W���'����s�ڧ �� �C��x�|$+�&�w���߰[q�=�!�&�jX5�G��m2�����)�1���\�����7ɒ�9��.ʼET�P�_���, ���$T��c/g�4��������QhN`H��6R���J8_s��� \�����'��P��	+d� b�p3�Hg���0k�o>�?�h���s.�0��@SP�t0�/�ē������ZJ���`�~1�����)�2Q�yL= �E�&u�k�w�	���E� k�G�J*���m_`�`�n�|V�o(D�>%�	�D �Q}�|�c �ZNI�,�r���p�*s�� Ѻ�߆� Ý�og�/RA�L戜Tc(��Uyps�`~9D	�38X~$i�8o�s�|q�^>n��,�|��rdIxB/d���5�P��@"����(��� #���B�-hܖk'�Cle*�r�l P�θ<w� ��xw�Y���%�+J�A�$��>!��#0�j�Q��!��I\�<�m�P"[� @=D�&*�G1-EL�`U��vBX��l���륈�����bX}|-���)D�K�@p������U�T#�� ���X>�N�m(��oA~$��l��u�ds/��i��E	��'Get��=�q �N�ă�;\H1���`��m>�{��{B���"Ο�)�: �1~4�m ���gB �6�d�1�sM�_nhs0�?D��x��(������#N�
`�tF�N]�� .ϟ0C^�`tˁ�� -����`�R���p�*���wO���艓�� �����
���옥X|&N���q0�@��V���4�T��Ok��xX\tK��9�HY��`/[)ۗf��R���+�<�%�4�.[���r�,�#���H�dO:��e��ʍh�B��
� �'Dt+F4ݨ��`�;��D�3��Q��rx���,�i!q82��8�h�Y�%�yY�@/�!� ��#�_C��$��(a_bH`sV�P
)�|c�\��3کu@��PF,��l:x#߬�C$�G'����)�J���w�^D�N/�Fp( ���ü�����M�sF�7�!0�Ml�,�n� 4�>i�a��A�1{%<�qk�y.�DD;�'ǂD�H4P�U�x�
h ș��:�-2P�@߻T!�l"+DuźS���k~�S�q���ڐ� o_l[v훿  �+Q���{��p���7T�el�!.�d�%V���M)G0��0���*�.0�B���d�s0�Ѫ�I3�㵗�d�[r�P�T�< �ug#��� �ҼtD��SH�ptL�� �a4��� Lo�K�N�9dx@��`�B���b�`��`��^ #q��T0 �ӏ��ױ�C}��`\��zihxb�vd)�	��J'�!�*�,�(4!w���� pXd��t[���'�t@����h���`��2C�tP��Z��X�:�(� ��V��P\o��þ^�����
Z��R �O���(��Y�`� ���X��Z� �>��V P`^���<��
��]` s��6[;aY�S���a���b�[��
T���L���8l��@��T�� m��] :��R��	4`~8'P��<����?��� 
U���Ny������x:��B�ޤ<N �b���!8P@�T���>#����4t<��G̴$����!Tob :�-�a�Rdj/ 2�dp�Hk!xN���`���$`��E�*�P1�j"���,r��`�aC/@"�����ȼ�[��$��,�@�`��Vt|X�����F�L�E�*��`k	цĴY��

�qb���<�bS�8��H���s@Ȝ!�-Ѭ����G���L g�u�(b��Ĭ[3C,u��X(�r&��k�h���@�u�W� a7��'pT����P$��X� *��;O��m��<)�^�@�M3�D��Tܡ���	{�RQ�PH�DH@l���C!��ȓ�F�$H��Oo,Ԯ$+��@o�H�<��"����.�|).��� �4A�u���_"�&�J���$z l}= �:��RBAI���3��3.[�AU��W.E���vTc�������-5D����k��Ns������ ��p�,"`���ʀ"��h$�G��'W�  �?�!`�4*}g[	�ZX��7�8	麵 !�
�'�idh ��ΕD�8�_�)�gP�²4i�Z�}=�s��qd�w|�JIC�u���[�롨@�K�� ��f�{ �gm��ؽ'��t��0�a�Η�x+# �4� �����;��u��D�&��D �#��b r���6J� GBWy��� �`K�$ Ԉ2C�P�:��	�|�l��K��%�K`�zZt�t�`pJ�Q�j����Nj/�#��8��+��Z)�����PtFC>Mo��d�� 1J�Q���Xl�8^G� ՛x��FK�W~��,`�1_�����nZ��H�+�<���[��`@��������0]v H��y���[z8���U�u����, �T+1�ft�:�!`��쎽^ ��g�Q�U��p^!�/�^v���0cw������N�@1�F�u�M���g�W����p�D��X���	�T蘢:�T�@ w�VJ��qF����C ���e:X#� �`�C+���5�� ���7�v�Uԧu�h��O4�Y el7�;��-��Т3��c��V��?d@ӕ�D�F -D9��l����4W>K�(@?I�H/���4;�u���8�I��d;*��U��퓬��J h����T����`��� .��U^b ���*j�K�y��� ���J�X ����!�1
�b~��`:Q����sH�R ~��
d}��^����t*A�y	����2d�HCs� )���d��K"��`����?��!� v
�ߞ6��h`� �<�g�H��=7����iN�cPn<�k�!���̞��0c����8JA#�c�-0��9���Qp��B�G�p�S+� �?�z�Jϑ0�阼&� 8vxK����!�I��D�z�>e��?�a�����}S c6@��� 5szo�^0_�eC�����#��rL���y��!�42�H��� ��D+�T�s �\ўK�}�0�&H`���� ��7���� g�yn�p!K�Ȯ}�q�wF�A����Ha�@ؚ~�q����Z ��2��T���wI� ���P�~��K(u6e�#j���7��
>��v�f�0w(E��j�|�0�zi,�v�����ղ^��)" ��y��K,'��DhC��/(R�mtt	Q��,2��tC��d7���a̉tL�}��Z���ԫ��E4ۛ��i�"n,B��jk0����|�{@�45�QW 		���Y8������x�`�H�vY��o�� � ��`�1p!��� ߔ �%��Hs� He,י
t����� <�եt�
��D (�1��P����ph���c ax��@��
0�5��M�$���!�;|�H>��5�@�ƹ���()zf� ��?yd�g�];���=)+�.�C�� ���������$F����H%�PG S�pkt'z?IAp ��m:���Q��^>��C$�n	���L����!DX�^����ހ��3s��{8ba�6 <�����8y�����s�`A��t]-��{y�1�\@��[�
c�� ���&R|�e�� iV(�� �T�E�
� 6��@7��3� ;�N�g���`|��oٔ ���Av$c `��·����� �&���9 m���#�"+�֒0�c� ��s ���Y�F �c:q�)��$�uJ�\�` �"С��ߗ�޼�𦚅 �>E|��� hp�/��W9�P�q���0���g�o)5 /�I�b���Z��OP�_!� ��pW�� V���˴��P �_n�ZC>fx �!2�?.�	*bҹ �"� Z�+��D� ()� E��`��`;� ���vU�5w�{��!��i��~�#pv+W���Mn���!�����Ӄz����*�˚�� �׸, j���M��;�� �Kݕ��lp�p
>c���e"ZVS ԕ�;�c�x� Q*���۳�r�������� (q���B�H!�ѝ 15�*�O|�lu� ��}�� ����]{㦘{9hs�v�Y !��pcӀ�ʺ����� �g�cwH!� ��>=�z����`BU�o� ެ��y".�b�C�r����� �Jo�գH(Y�~����e�HX�`� �~ѧ� ��� "�� Y�uˣ]K\��
л� tge��� 
vb���Y߀��J4�N�3� �h�(���7����kp&��9b@0�Ch{�`�pH� /�Nѕ���
	��O��/0h�8n"���	�u�`�����[ Y�cS��o	*�e ��\����`�j@��$s� N�u��H"JA@!Q���:X� p�m"�Zu�n���k*������@�T������| !S&Y"H�֠��c ��y��Õ� G�����ѵ 4 �;FSU��|�@�)�<�#� oƠ-��v�)�{� ޕS�3�|"9�h�e@�:��8�������ΠM�c�0�� s$a!��َ ����ƕ��ti z�����u	�p�� <	ǿ�Jkc����0�� sѐ!�� ,�O��G��1C�}1d���5 ���^W�����t���r�˳� r`8���/�җ(���q����W�TH��=3:� �V$��!� �� S�7����@�2 �Q<����� t��� �g� |��ck�vLC��տ �cn@�!����4r��� �"�/�ˍ�,���Gd��e����:��$*�U�� `d
lhkè ���ᕽ߬�bM��Yù���E� \�!s.�c��xIl9��/�֡�N ��v"���i�������W&�Аs�!��� F B��ٕ�}�b{f e8�<7�^!�B���Pv$�c��Ġ��`)��r���D��h�iZ �X��,�%erL��~�M�x� �� d�,�Ͱ ؀o�c,xP 4�mv�[��s�@`U��͞����`)� s� ����x���c��� A�3PQ�5 k���v�$\}�����!��O� %��9e�uzq��T�p �8�]bt� c���dK
w ^"6�������DЂ�K�s��d@�ba`c�F�~�2"�Z�b��>�@�;�!�� �c�� �+&"7,E��u�|wbP��pw ����� �,�(=�M� �p+�c .ҕ1��"���� ����?��:o ���c�-��}�t��JL�{�gX��ą�� rGw!���,) �� L�:Ѯ�OR�caE��2e�b�`�[��`h	c'V�,���R�۞���g{d�x>�U�� ��|�e�xB\�ޘ��@�a 0"��h�	���� �p|� �\e���`3!�g���x����|b���-Ҿ���<�?��	� ���`S!�tD��t�ps� ޘ���B"P� �I�f�Hc"@�* ߖa��Ǩ��!@?�>�7.K&(�|�A:h��ô'�0�v~ D����t�+�wg`� K,n���������G�� ]R�a�rͱ�=w���3���(t� #�$	>!N�"<�e��&�i�P�v�}*�xy �B�М�\� � ,��`t�c�h�Eė�H�ΐ4=Y7S;w��@V��|e�� ��]�/^$�ń �R"M�\|%g��a�<��^x�[�y��w"
d���� c$s^L��.��3�æ p��!^%D ��}��\L~� 2`<�>�.��D0q�j���C�����>F�)��~�����ڽ����@�JPx�n��[� �(	�f���q�9 iց��&c��}�_K�sw���z��6��o��|R�p��ܕS �Ѐ� <���q@'� p�(c��?T\N��<D���٨hӡ`0������c���Lo��A4Bxz.�[�!��J� ��J��	A�c~  ^�s.T�� ��A���J��ݼ�O�\N0��,��l �>�p�T"e1�F0��&|bǘL��	� ���VG9."�?3��NP�mc�j��"VbX�q#h�p�np�K.E��G��}� y'"a��� �Y� 0A�Q]аT�,d�6q�@�`u�� ��9��0
�c %�n�'z�MU����|� �m��שI�s���Y��=��  "`l�0�b�L����98� 7��_!��t� r�C�>:}S�� ���pq\xt$�!l(� +F	*�P�� B���ؕ9�\(�c�� ��a!���K�����A`�M�0��3DT���i�+!��d ���e����&����E">ۍ��	6mD��hR���֠u^�{�> 5�ȣ|"� �w����m���d��{ P\_#03:��
=�s���8x�>�(/!$`����bk��z�X�d$u�HFz�\�� 9v�����@����V=fA ��=��m} |� ���r ݣ�b��)�����ڸ(f�e���`�#.i��������)
���,�Q����n]� M�`e "��;�m�%,�sx �G�6_����3.� ���!) �W���cŻ����V���ӈ�c�^���Вxb$��l��&��NBA������b�z{��:4P�`����� %���E��c��ⓛ(��� �������lӳ������ѵxg����\΄��:b{�ؓ �����H�� �b"�1�`����d׃8n^|���c<�� �=Ƅ�H�̞͘�u�`o�0�`1�c�t�p�@��������� mªP�E����y "�p������	ގ,� �ʪ���� ��zN����a�N� tK�d"�� �����ʫ�t�`�pt���,�������m�؍QL���p�P 5�+� ���ꢌ�tŇ;	h�,�@�A�/��O
5l�`�?࿭�� +�`��e B�}�����]ٴ�e�RS ��+핬G� T�$!��Q���Ey(�b�[B�R�@l) �3�Y�!_ z� �9ˌ�m�0��, G�(��*����� ������ ���'���C �,c^B:�h�2!ö0�׏�x��p
ʕ.� 3Cp��ZS�O�4�D ���Fḭ d|gQ��"���� $Kn���x c2ҕ�뀯d��L��!R�S�d}	��bL� �u����tZ���!WĀ�~ʏ�>�LLpw/ #$3� n� �:J�YŬ�� ���(�`����^ O�������y�)�O���#n��5D$�О�q���gj�0��A!�����E������ rq�� ��D���}*��	�����~���uۭn���a�� 5������"� �	,�~l�K��@��D�A�<������ _�q��'`�К����?- ��XRg�� s'����� ����znxfk�|ɂ�%�Z��zq }����Ҹ�Wn��`��V�9���T�
]�Y�� r�z�y XQ���?��W��Y8`U�2+�v �G.�z��U���>��9%'p�?�ז �n<�����A��5e�P��;��� *c��\��0 ���2e� �G�1I�� �^t�]�����"@E))q����[��(��_� ���x�� vkR���/su���ֽ�Y��H)z��;��Ŋ�ɀ(�`|e �ݭ�p�8�0�6|.AJ5�E�ԩ�K�չ*�����3�d��;�)��`ȣ�� J��E�>���������zJM �ɨ=t����/���R6�2� ����b�g rHe�/� [�9h6���� �����c| ��2"�\� �����
����v���4��Tp�%D̤`R� Ya8���}<�z� ����? -ŗ�5�O� `��&�h�:cӀ�2��goI�N�B& $� �H���� �~95"SDj��G<�yv� �lI�����?C!4���?/2: %_5�L�o���sؤ�0�5
�9S��� ]�� �a�[�����Nr ��q� ���(���ư�y8��5V�ס�.�g����΃�p�� �!A��5= ��zb�[���6��ajO$��=�PpV��� v�֜����̱� j��W֫u(/���5# ܌�G��
�>��� �.v�l  ��y�5�M �����u6��0���aDF��2���i�V �|�۫�[Yx_� M�N!4&g8��J�nQ5 ���E�F �ۦ6��3 ��4>ӄH �֪xP�6 ����� A�7�pݍ5��8�3ϰ�\��)?y�� W��[�IM/�9��l0�h@�<�1�R8������� ��șd/cV �s9)�� �����vSr���g
P����E&��KV� �x	�����8�p �ʑ
�ly)�2L���u� 1���R���<�m&�x �π�c��U|�5�n���e 12ܩ��8� ���/���P� D���=u�g ��4K!v/�����O�@ ��9Ɉ���x�50
M��F�e�H�?�X��<h������� �&��K��*��߫'��b����8T�y8	� �ɓn�U5 �Ј�_��� )��Xc ���Y_�Ky}f��+�D���L6�\ k�S�K	�� �����d�; +FTm��Mle�����}	������0���
oQ�3� 4�>�/ ƾ�!fsT bA���| 0��6��S U�1��]���c�����!�����5e�V�i��F�6���p�4�ȴ��5�M�f��Ȧ������3��H�k�8H�VlE�����4�U��0��tG ql�d1Ex>��pR	LA��uF!A�����cd��n 
O���(#@�5<S����{0���X� g�ߑ� 3�ۊW�H:l7J�.4c�Sy X����a�� �ɒ9���g�\�����C[�5�9Uyl ��Ȑۇ#	]�>&��; ��H�8-H��$�	n`vy]� -�ǅԟpR�5�yɀL������� i��%�����y �4Y�	f��gҎ�pi�S��-c�D�!���וo����>���a��9�w���e�k��z9�o�b��$ �����.[e�R@@I� B'6��gƞ���<���?���>5��Ș0<���@;���	��M����g� �Ɇ>+�4�\��g� =J"%����5(aɉ��՞p4��Q{�p20Ls O���� ��.�F��)� H�n*�(�����f�N0ڀ�n��8��	=.o�w|�r�� 2����!	 ��� lH��S�5� Lׯp��u>-Z��ɺ���D[�q��Η�dc,��4`�X��.<��"Q@x��Q�J���֡�&��0d7I�
AQ	��C&�qɚ�Jph����2Wg� ��U'�8��8���p|��Ij@��E;� 3����B�u� ��2%i?HH�s������W�Ӏ�׏ lZ�XFR�<8Ѷ��Y���@�A�&qL�\< 9�%~1Lxh ^u�b&��yՐ���<� �[9:��Hp� ������(���~��dPd�g��1�ۘ�/ W��M4�Ț����.�@S����%�3d5`���@�VP{"&���} ��/���P�>6L$��8��T��'��Unpy���\���1�`4� y*B�d��H��Z�b��u��+ah�3ʰ�.k��6O�[��&�PP�����,Ȁa��� F.���H�X� m'̠�� 5)�Ȅ���`���4-0�f���n�� C�5z�Ow� ��h��/Q��w�`�p��3
����@ɪ�7Bp�5��羯 ��x	 *�����a���c=��ܨ��E� P��W��2�D5�IɞEV8�� ]�>����� M����}`;×��א̜ԥ8~�	A<!4m�N��K�}�� �׸/ ��8�����зJ��,#���5����0̎�;=@B�w��(7�� 4�=Tp��b�n�5И��LPdB��@���?&%�� �U�d�l���2V4�Pp� 5��nm�� ���W6��-8�����K")ܪ��8Dؗ�7���n[��t�AV��� ��)6+�ȱ������,?1r (E]N �4�
Ǳ�,�H" tU+�&�F/��?�\� �����@X���}�Q#ؑ Cg�F"�0� B�H�ؕ�-�Ngէ s�A�.x� �J�;�� t��f}�>G� �W!\R�5�� r{�Ȗ�EZGyq)� `�N�F� }��&��8 �Ȉ�	�B�H�&�@�0� �ɳ�5y6�dp�	B����̭ @�s��K�W��+.ɝ�G�V�`��y`�p��kX�K����0`ab�]��=�8� MK̀�T5|��B^���tM�xn�������ÿ�;~,�`�g��Jwf���ŘT��� �eI��}+H�l ~S�B,�O�<&��:��o���f��Ɉ,����s�(B���+�HT`q�8SEX�u�ЇkU��~���FNM� ��&61��0�[�ixl A(�� ���W�Zo ���� ��HP��4��.d����)���� Z�5�Ɋ����V����6*mv���&/+���6�T]�>d���3��O�Gop��״7d���xN�h�hC��D�ա*x� �r�y��h�����! w�v(qEf~�Ȝ��`���&X����� ���5���1���;}paV~�pI�!&� ƽ���g ��Z%����PQ�Y�O��� �l6"�5��e���!3�c���6w�8��\<�"a�7@�D��� �*Wy4��L`HNvƋ�����χ ����W7��ـ�y� �`��0O�?P�t&vd- �ƻ58��߽;��K*h��G�4��	c�&��lU�{(�5@� 2wɋ�������	��	Vht��8�g�W�PɒS�b7 ��.w�@��{Զ��`h/ ɜ4�5�.$�-xg YH�� �����.�` �f%�,��$Icdߊ U����\����(\ ��]Uj\9���� ;M,����` Y~�7��8���u^���0ﰀTZɯ$gs�c�>��+��Hڃb�9��[tY Ȇ��XIV8��u� p��� �i��5 H ɟ�����^	gØ�@�� %ʾ5�j�\� ���|���Х�� �{�=�k'93��h0���E���bp� &�5��M�V�20 t��N����i ����s[�5 7w��Ce��%���@�0����� ��5*1�~F���=�>��� i��Ԕ$5�LV*��(�'�s7�jl[��nA ��E�� R��4��%������W`���È��(ാ�c��%v������_� ��0�n���5<9�j��dWF�� {�\� �L�2��ϐ�\t��b|�hvD��`��� M��3(�5��c��6P�ʈ
�u^(p�Cܪ� -�|� ��dŐX>�,7��-�Ǡ�ΰ ��5�iɩ�����F@����p�ZA�J |��k�� �w+��nc=}�#���(��s��M�/���APE���,���L�0$��g��[�A�p��u��ԁ��e�ń���F��*� ��Wi�M4�{t؀6"��D�J Uq٠7�I+t��p�X 8�Z]���ex�\���`HT��m�E��5|V{�S�C=��<�n�7�1\3e8L�� ����Wٓ�qk �d�C�. ��)Pڂ��m��r���p ��Đ���K�}f6O�܁'��x(p�혔%�i��@��/Dczo���8`�H��| �k��4�,�x.KSF���9?�|���).�ĺ	P-���˅��!��A�2�܁��b,�	������%0 {g�:`fd�cqp�ِ���9�3"�ȉ�������z����P.��	�'�Y��o{`d�g�� 8��HG4�MB@�3%(���_`(�LR�E�5��㇞.6@<(e�8�� �́~ә�P �G�o�xL�LP��9e3���!S14L� �ݱ�o�n(6�����A�',B�D�}���W�� 15�[�6
¸D k�m��?�A��Xs�[�� h �a����i���:���UK�����5 �	���
�� ������� n���ڨ��&娗��СはD� �5��́�T�z������.�� $� �.XU�,�u����w����]H>H�}�Tu��SybH&W��`��¯���0��|^ID=�<��)f��m�n������x�����J�zjP	@�g��,U����H�N�GG;� ���5|:�d ��O�����4H�� J2S���5'�� ���OP$p�|�\��WB�tPR�Pߨ�  `�^�z��9�2f��ɞ�Ȯ�����o�&�� ���p5���,с��~fo��,�G�ϝnGY�@��4� ��X���C���D/N��v��Q t�q�s@�(����>���H �+�)��zEb�n���UV� �;�ĩ��N��P@��>�4g ����^%����KY��,�3
����� q9�G�&��z@8S, $�|69����4��%bz?���Ø�G t�r@�5R�J��]v��ۀ���T"�����`#ρ�W��� 6-S�(5J�P� ���!�P? l����uB�8��p�� I�<C�/=���.l��y��08UZ "�g��2Iͻ�X�h@N,i|��:��L l���	�&4��`?��P�5wa����� ×��23�#6*�pΤ�<������s�]���x0p��xo)Ae�O�$O@'�;ph(Y2���C�>rF<��ʋ�`.X� O`�E�D�������8 dw��,��K��3.�@o�D��9��$�e��f V���U�@��l�p� d���F�q
��ר
ڙk%���2��� �����DqA��&� ���i���5P��N'8Fc����0I�Tc� ��{���� k���c 6�Z��� �����j���R �{ǭ�w��W.dC�P���Klv��ץV�@����Q[��P��؁�nZ Lf7ep ӹ�ך�_��)�!����9��O�EW렼x >B�ug�6��� ����O[5�0�ȓ�@�g8���Z� B�Ϭ���|(�T����Y���Y/�@ܪ��d,�'�,	��,Z���^.��|	厂0@�r uI��jU(��TT��u��!�4 
ɰ0s�*�~�/�}�v\�tl&��Ĵ��Uo���4�>�p�����<M|)x&^2�o�#3�
���$�g���Vp�v���� m���	�M�S�� ��k��n6%D"@�d���K&�� tɨp���JS���h�R�0%��5��� ��z6�[�P�Y}erH��0�� �s Ƶ̢'���2�r� vQ��59�.{�� �+�  �x�l0A�� )�~��gt����X4��`���u�*傟���#ɓ>���=�]�/��x��$��� �=�bZ ��M��BF�4�����t!����5��@�V���0p�tڭP� �z���Iŏ�d@���H85L5 ��1e�9 �2Z�ȹ�7��]>���� ��&)�C�eB?��>Q3vi��},����M8�Kj%�&� 8o��Ձ��L���u��q䰞�6(�� `��5��|�������ov2!��̎;'��w养 �pp�� !U��5��.�� �i�(�B�p����oӈ���n����� ߫ۊ���rH^��~(� ���N��p� ��D�'��}X��G��� 5�����8Y�g"�%M|�� ��os�3`ܟ5�Np`4h}�W灘#�D`HN=�䀖���W �׫����!,N�O�l�K�  ���� �y�8� �pu M���G��$�A$( F��c2�O>S x������	W���l�� �A!��
&��4 Ri��O�����4�z0�g"� ���Oy������`H������� >�R�f� #���II�4}�q0>Y�P�`@�f�/ �i���tP��s�� ���1�>����`� �;E����i����b�p�ě��8J� ���� �� �16̠A�x����e@Pp�@�%��׿V� }8`���R6j͆ �X_v�5?� �4�&ɚ�7���E�c3�-ٖI �mr��!@���H�� �U�/[�s�x$�6\&�<("�X��*P�`,�� % ͓�L{~g �y9l���x��\�Xx�`��l���f�� �!����� ��A�Ȓ(��e���6W��YjC� p����"� ��5���x;	��a[ ����X}�OE��K6��3��`q '�Пa��/f�`�W��A<+�@4�pɰ�����*K��;�`TL�^%��+��?5: �N����u�ge�l Q��{�F� /�E��iᴇ�$���Ǟ����E�D ~p�(�ȓ���� �i<m ���1潰�|6����Z!�`��45��HU|���9�4��� �
��d'��x�<�)���{ Hؐ�{c ۘo�$�DJz��J�1V�H����~ ]����3�R#� 	��&<V	@�z��xv$��" ��'�m ,�
� �u�A����	���%�����`�	h�`�^XX$�l	��A$xSH��8h D��*c�	|���w�s `�"?�紴�.0 ���R��(1������wV+z�L^y,1� 2�����6���a�����H��h
{r&A�>�7|,�Eа�o2�w����+ \%���l�X �{�t��0ݝ��+���n`�_���i�W�p�<��+) 6��2 �70���b �;�|
ɸ� ��G�~$k��� �`n�7�����֝��l�q8v��R�����Hx�j�a����״� j��� ��p�0޲d��(	�����hj6a,ħ밸�G>��x�@�/8��<'>@�h�lץ97X���M� �3k!8�WS�� �fo4��/�����0��� ��'XH�Ȏ�؜ێSN� �?��V�]��5Ȝ���Q/4����0�U�H�8;�A�������K9��Ԡ�X�� ؂OX| $�a��~�k�(���R���k�c�<�� ��'�O|{��[����������Q�l�wBݢ�)�H��7 �.�W��G�_� x��?�Q$X��8$σ�H�b�+��J-���9f����y��k�F��ד~Е3+� ɽ9�Z�� �0$e�N�p�z���� �Ԧ˶�;:6��Ȟ��wN��� ��`�E���;�O���Y+@��4Ș�	�L�W���=?t>	����"(u�V%{1� ���<]HdA���E F��Q��S Weɻ?�{���cg鰐� ��Ε��[ 46S8�Y	� {xZ��\�| �=��b(	x��4c�`�a���%>��WF>���D39��Y!\�%P�n �'B5C ��׽+�8Ʉ���p�{�� ��U�f`�5�+p�2��	�� �a��"|7�N��6���:�<ϖs��X*�8�BG�v 3��5<� ��M�n��p�� L!�����4�58�˪�e%`�#�pf{@p��w��߈$�� �ox����-�����E���/��'t)	Y��Ҏ`0��O�|L��ۅ@�N���mwƴ8�	 ����"�0����� J0π5LH��s�RT��$6Z� �&�ɶp Xa~T5���39�4�.�j|� 6G�Ȯ� ��2�/f�,� ��WR35`ᨉ��{Є��� �Օ����u�-� �}5*`��p�D�H���LN�\� ������ �|�`\	L���$ K����X��4�P����� �p������^3p���~,��H ���f����5�攧`�px�����u� 8��tR����5�j?ipQp$�[p@[�R��Q51��T���W����p��PϠ5�c? 8e�Zo&9{�DJ�����4A�6�~ ި{�������3(��PlT 4^�Ȱ�d�� o�1t�!S�6�%�G�п5A��b� g����6+��T�OL��ѩ� eX�ى!PGT�
�5��3^�k������)D�Q�T�\��*
T��Q��E���6R�m �3_iC��T�בP�E42���F2W�x��`�Qb ���86��� Ӽ�ɯ�l�%��f�X� ����U�T	��H4��f���������h���.��|���" AF`�?���WčX�pF<�zԉg����B�#p`��d�N^u$�ݞa�6q ��w��s<Iw�O �&f�'y�%�z���������=老���@�Դ5����TJ����9�+�Zd�@F_�	�b���ԅ�I����yl��V����Y��[� 7� �q�b�u��J�R�o� ����4cą��z M�o��,&�P�&�l�/����R96���@���;Xf��?<��g�琺Z�f:� ��9�r�!?䀰^� �����5��G �jP��� ����REP~�<}�{� ��Z�Lyh���#�� �$�� �8���� �ɄPv��/�?G�E W�; �8�J��,�@�l���G��ӄOYq��p� ��/
ɉ@0~��]�� jvT.�� 3�IB��f�0Lw �!��s�Q\I@�z1}��! J,��D� ���	@3����l�@���t���(ϦCF| ��#��3{S�n]��0r��!�B�(3��iVW�ȗ>�I�t�M�����%館�	v8��uh�`HC� �ԅ\.9-E�R�2����~$��@�P@Q��-\p�2���<�ߠ��P��5-�N���D �h C��u_8�&��h�w� e?%�H�4>�g�&�ĉ�L�rs� ����8�� I����K�<�Vɥ �?!)��P��� g�屑8[��	�)�tx<���Y/��:JD���)j��0�� =��4���%�)ap��y �3A��]�N�L'R���uh/X�_�AO �`ɓ��2�M�d.x �*�?� �ϳ�dLӀC�
�� �f(��rgH��!�EL�a ��5V��D�t� y;'�t��HX� `C�5��m&{hn ��xUx��D���P��d�Lj��%�h��cGOSP��� �m���S�2��TrD%�$�o��%�$���|�T]|b��n��!#��&�IH�hd��$`���K�f<�\�Т�:�$+�^TB�M+�$.�q�^T>x�;ڙY�I�Ex��B5�S[�E�9�( ��:0�gY�� Ȩ�o ���xd�D��T�2��Ia�� /�L��JT3�\�� �i�V�2!����rݔ�NOF�#b�[��0�}���5?�e�L�L�w����ـ�T�&C� �爾t�8V�'� �� %��5�o�aeu�WQ���� S�9DBט��06z�l���qð�T� ��sM�{�E�����Ȑ��	) ���3-�0O����|#�b���@ ��q�_Q�J� @�%A/
����� �����YH8�ot��> �m�q�ƕH���>Ș a����d\�t:^���a& ������׼ǥ�y��8k��Ç\S������706�p��'^s���`�hp��lǼ����`,���}�>H�st�P�g��C����ȷ���/|���w�s�@�� �f���6(t,}� W�&5���>�"� �Ⱥ�X���H�G�(¨*�D�O;%$1,F���^N�ȵC�:V��b���]�[;�_ ���	��R ��\5hɷl ���7 h&(��� ����u�� ?ե����/ ����5fpL�� ��G%�"0�����T'O�L}\4�p���l��H�(�#2O���� u~D:4�����PȌo'�{�x� x p�'iu"�+��DP��� O�4���>0��pxq�t)PG��|���U��`�oi����n1����VĲD\�F� c��M6����8q� ��U���b��3�`�އ<�� Ι,?pj[�r,:ޜ,� Ȍ�_�'���U��k�bv\��3�
���W�� ��${�f���w �F�˾ue|�x@���:�O�60�� 
,�	����*�ln hv��a Ϧ�\�7p��X������W�y����]���0�n x�%�G���z�Y-��b@�p����շ���H�\k|%�q��[����΁�W����b�e�4�h�R��x�X/24DJ�hx3�D��xk�\�x��%�4$�Dq�!4BB�|�Dܳ�˜xF��3nH�B��T��^a}DgАT���D�­@��.�D�� x�D��xE����1$�CZ�["DySx��#P��Tz�]a��x@�n`ۋ�hߐ�3@V"~��� 1�h��8k0�������5����ՠhQ��� n������.e�����ZG��̏5�j��>� H=V��d>/�0Y�_�% |����)6� �P܋5Sp��킸7�u���ˇ��6�`�5 <=�Y��o��J���^� g9�.�n	oƙ\�Yȭ�m����0�4��0դ@��<���ʘ� K\
��S�g�� ��C?�@6�@�xcϘHiTǀHE9�w� ��+u.�H D����O��7�A�|��@XV'K��H�M���w��`��V�ץ�
E��w�	L6V� �9��3>�\?�k|b � �l~��8؍ �'���G�	�A��d ��"�F����7��_!��UA���2�8��8��B��K$:�:</'�R0��H��� �ڦ y�8���6 ����e5�vdVf����)Ŵ�4���/�4�=P,�L�AEA�Ӏl	{[Q����2��OɊ$	�O� l����P��v���@�F� n�a���)&O��������tv!��E�ڀl��_>����c �>�3�g�A �R\E�Qa��	�h����>@8�0)e�m� pa	6"�#�y�5僠Y����s9�9� �	@�p@�Sq�_z��/�x :��߫��à� �>��������*�e;�-ca���.F��,㾞�3<OS%Z��Ax*��� l�eO�2�p��`H�hG�ϰ� A���G���%`����2���A���N� $��.3�����hɏ5�eݓ�7������v c��4}���ۇ����� �G�+f>&�  ɬT�����N`���M�%�J�5W�� �v�yf	��dЎ�����G[�͸�Ϊ9�e��sP�� ~2;�/	(�i�T4�����`�	M�4�X fĈ���� ���5��
�2H� �e�L:�	���0�W�C����A?U���0�����t��PX�@�7A?]�pTU�@0��5<��Y�w�,�?��_ �@�@����ɐ�5��~�V/G����� R�569^�.��� Gz�_t�~q%(�R�����	�&A �t� J�o\�Qph
!�"� kL9�3,�x`�:6��Y�w;_����F��p�E�ȏjd������_�^�H8�"���<0񷋔�xDͲ������U	Ð�D��S�dk ��Ta�������R�����~`"�����E�$����,��`�mx�����D��خ(
<�� l^��'�R� �P��0B؉� q�0���K�2��a-`���p5���l@�b�% �52�ȒSf���	?�|��C �q���OȐ���PQ��2W��H_����Oڅ	e|$��J�>Ѡ�Y����aĀ<����qؙM�CB��~���5Ve�(X�&6��a �^p�kf�<�I�����9�1��N�_� �L� ��U���� �Ȳ=`oy��S�@�U^��G֐�J � �)u�����6`h_�$�r� ���BL��J-6w��y�u�,K頫�H�.� ���ؑ-�V@��X�:��tq�2}�����=�>Y,��H I&�<�����5as�h��.�����qσ���l�_5и�@���v =z�\��m	��ae�^����q�?�0}j���� �����r��2�``H� ��4�FvL�H)���>ݚC��i�{ ��<7.�Z	iА9w3�y U�o���G�V]
\t�Dc`nޜ�p�� ���r�h ������f��@����n��r���"�H�O�4N� 2٦���Y鋥i����o�j�|��`�g�� �Q�P��5
�Tz��Ȅ�/��9Y	��ڌ s��n ���g�=6�y� ��{���E�5�'�3 nX���,	�q: ����4�j��u��@�@��7d� "H����&��=���;IU���@��6-�(��u2�%�D��耨P��G B�Mp~�5\X�� ��4Re9�J���P����f@��]���]�ЗPw46�	��@�~��$a����H� ��=�Zz�B6��_����F< h�`N�����s��$� `��ז6x$	t� P�|k���3׆�Ht��'s��˔��^L8�e#��v	�K�������z�Y��0f�*��@�ʢ��p�$4�� ���-��4.���:T����{ ɦ1�訠���瞧 ���w��.NE�@�K���P	v ��+f^*`�t��`��kV�?�<8�9��d�X5A���\qu�	/ܖ:�_	���8�i @|e6��c P��2���y��4`&�Ж���"x�k�>�4ӀE�5&^Y\�`��L��w�	e��.4��6��9] (����[0�<�V�J��ȯ_���``�8��ǘ G�����+��2?,��H�"�<����6|��0n��8��༩'������)�`��*(ɚ����X:�����}�}�6x��� XS�q݈>)�`L
��ϳ4@�p2\�D �on��#.F��@m�Vʾ%�J�\��C�X�2�$8����Fu���E�,���࠺۽����P��� �n�5�zO.Ĭ� P)P��/7Q�p��?"�d���y	�ԉ`���?���o�_ �[u(>�e���� pw/ ���\��&E�X�����5 ɭoь2�St�>�dL�Oc��E��p� ��3�n��V�ļX�� l�W�023`R�5� <�$�j��v/JK���) 4��5�|� ~Ϻ���������>���,�>/P� �q��bkWL�u�s\Ԙ����K�շ ;��A���h.�s��B 0�g�%Ă��a!8�E`�-Y�1�gk�N� ��2 �&pT �Tc<kE���v��\8��~%Q��� �Ɏ�X c���H-!py	V�ސ�'Cr ��{ �5 ��(��8
 H�4s�5Y��N�e�� ��FY� �b_�0�p�$ڤ� �mW�p&��܀d	�y��]hV�y ��Y\,Ay�Zsz�S�H�� 8�=We��Ȕ1l����(���h8␤ �dW�n��::��	����+��03���`�5�������l+^f�@��6IS �x�V�5;����N ���26 �fB>��`1�m9��84���e��HNp.����7K�]�h�X S������$5(��u:��q&d�@�7[`�����I�j}�"�G���X��u*/���5T�,@֥��;���Wj3	4���@��<�V�@��Z\`�i�P 7����@*d=ʹ��M�U.�5�|���KЙ�4X��v�Ŀ�w 6�R��6U��\�P����Nގ�������A���O\�bL���ޜr4�K�x�	s��� 4�Ǽۉ �%5z �F�i|�ݗ���Ҟ ��/<e~�5��Ȏ�Pr6\��?�N� i���]N*�(q���y�FXV���b������T#�{?�P�-�,0�r�\0�[�<�@�i�r%�oht��P$�{OE��KP�_3����0 ����/� �L���3)��4u��5p %L�:��`�8�k!��u��	 P):}�Y�,Р�0H�^4����H0pN\�#-�� ��h�����5P��Z����}�.wr��}x<��T-a�ԫ�4�n��P����=�. �����O��D� ���\[�~O���WɃ����z?�P���^U |5Ɂq�ȣ��Rr�>� T�V��l0p�6(9ɛ`p��=��j��2�IU��S\ ��ץ�� �5h��f��8��F�� �蕷$�(¢&7T�	��8_�W�������96.����l��p	���` L�x�Z����hq�wo �]����$��p M����c���@��_ "�F�	������� G��6< ٨�� FZ���< �P �K����3�n��<� �����
x�-&��i��a��_�p�{@� �> 6.�Y�ګLg� ϗ�t�3�	96* �r���5wޡ/KjÀ0�-s�U{1����pL�h�s��2�V�$
���x�ǒ��`�a ���5m��->���N ��|�#��(46�^���]<m	Ɲ�0�&P<#q�3�B�04���yOz;�CL�6 ��4�"$�׻_���
~�q��Br����w�A��L�����8���>���pD��}0;W���� �T��Eۧ� ����38e�p�P`Q��މpV�c���>�C�)?Y�W ��d�5%���ƅ�hɨW���␩�	s�����R@d���r��	�zʀ����o Id��ב�Kuɟk��]�;x�uI����� �����\��1�����:��3f� o.@�����w>(���� �/;�i@U� 5B�Ȉ�۵�ڷ�82�\v(y�����>�����9��A������p�?�1��WeU� �䂳����tQ#r�$�D�*f��p�p�y/���^�pu��%��t�l�~� J;M���JF�8c?9
�5g� q�d�YJ%�L84 �;���i�	�(�3t�`Ϥ������|�L(��C/�x�`��]�����.6�M�m�o��Oڄ �bv7��I��4��N��/fHP��L�ȏ������z��c��Qհ�9F3{��Ƞ�· %������Ly�  x�q	'�n�5��Ppx�<�j�H��PxyG.E���S��8�_��5���0�y(���^��\��U�5��"`�3L�h ?���G���'�(��V�4鼐	�p$WYO94�$�|eXJ��N���������[e����|C��9Ȫ�X�7L���!���\LH%5PvI .��V6��?$匤 B0o(ɰ�p�,3�,��@�$�+NmU|��h�]�������'� � }i>w�p� A!���+��5pp�=*
�����3�I� ���9�v	��Ȅ~�e�Ղ��@�p� s��։��� 5�����I q���BU7�����ɴ�t���[y�D�@<�Ջ�K���;aX�4�6��p�����K�}��( ����*H��Ќ�hÂ�߀ܐW���.ݴȡ�� ����:s�p� ����I5�'&�R���ˤ�/�9���K��(/�U`@`���F�LdM=�?���\�#���T������5P��:F���`���n �(�=�Ѐ���>���E{ �K;��2���Z ݕ5 -�A=ה��� ���/"�&�'��| �M�����|8 �5��9 Б�b�*uxv�������F??�3����*�|�{� �R�]kj[pD Et�q�+0�<6�� ��,5'�?�:���� YX��G�U�b�3X䝀�����Dχ`��T%�ft
P�߰`�F���dd$��v��;"a�0�Y$��� �K6t������� s`E�6:��{��P�W��� �=� ��50���@8����r�����i�,0�� �%�!�ȕ  �Q�w'[&:�,�-D8��4w(D�$d�� �������JX��) G���y�@'a�������ZF ��U�K��%������6w�%��҃T�W�0|2 X-��|��/���!�ژwH �U��5iV�|&�ؼ�bC�l���=ӊ@R��:�	���X�C� t%�.��H�� �ɺ��Q��+���17mӆ:�؇$l ��!�[�V��&��� 3X�8�R@E@��v�����������^5�p�A��3*�$Q.� L�5�a��	�XU)���Y`0�R�u��k�>�4$X-d�i"n0K��a��.	 (�A{��D�z���[g����po9\#�*��D@�B` ��M�o�����A0�0����� �P̖5� �ȿ!vs��\p�8ʘ ���p�3?���5���bvA �&�- �Z�ڼ�N	�,�5z��(��` #�~uJU�్ �*I��nހey����f�������i�*��y7����M��� x�W�_J�(�L�y ����V��/o��`�C�蟇�{�i �Ϧ ������!�L��m�aJ�@0O;p�l��S�f~�1���X����x���<;���|8$��爠��y����� ��X��H��'��.m��,� �s#4�Uc�a�КG(q=H>w�B� �? ��%x��5D�H=��<��u�-S�8��� 9�4���}12��'�8Y ���g�%��.��0��p���EN>��C��s�Zr�H��{�B�} D�K��T9���� "�%� ܾ�B�� iG��K��Th�����Tk��2{���y�Z[ �'8��ҕ���G��0U�9y>�o�+�"H�@4	_&U�GjQ� ��׾� �*���<������˼ �@o{����w�;��v(��|�F��p�3� ��5<�Ț8�����4ՙpb���GW��YHz�@���Vh�:
i7�� ��U����>�� =^岺6!����@"k.9� /�e_܆�)5�偀��+�tKw��0����IF�L��hL^m�7�
�
��,������9��k۟F �H��܌ �a6O�t/�+�wn�,��()��\e{�����հ`�Lɴ,�KӢ�3����EO������H�� G��W�h�3p� ����E?*}NUܧ H֊m�*�����@� �4#�V�8`�oހ��IAf��<�pC��p�ɐV�0���Ⱦ߂��K� #�{�d��x25]��Ң,�bh� x�x�)�����4e��
xN�����K�}���{�T�'� �,W����.��('�`�� N$�s�O�	�� -J�7s���	�#:�������<��� ܻ#e�O���Hz�XD_�a�@U�L �G�d�5H���@�=��~�X�� r�8*� ��|��&�J���������|z;�<d~���	�bF�܀>
P� 5Іm(h�4� ׏�6�~t碨��%=�B<���l���1�I�$ �N�#+��JH�@Ɍ��&��ƀh��f����AF@bc��$�,@��Ȅ��93��/(1��Y	��a��`�c��� �W��E b�w	)��f�:����5�d�� �ȫ0B�	����e�8Q��g.��� ��ȕ`��5���Ze�r(���^r��:��N ���8(�� �/�pl���0pm��� ��Y����2�\n� ��lPڅ����}�f�`��Z��X)9/5"�0`���n�a��.�bLp肨�`�Ȓ~��69�8䇾Ӵj�ĩ�0p�)6��4z�j�����J��Y t&R'�+5�s�5�,�]� ���8q�Uy�|3f�,�.@�1p����������+ T6� Ͻ�1���{` �p60��1$^��v�48ͳ�X �a&]�>�O��� �q��ΐo�.5V`>���l���<�k��Tn�P#4��\P �q�5*�@;I<��Ƭ����g��z,(�KMX`_��˅�<4�p�l��P��>��d�� 4�pV��%@��� �V@ì �$�WP�����v<d����P s��;�|K�j����T����ؽ�%"4w�2��Х p�85�v��*犨L���/�����}p��1@����8�樿��/r i�w |aɣJ���/�Yx3b &�5�$\@>@��A@��,�������`/��B�\�Ȧ1����8���!�ф�= )#��e��g F�]���<C��
���!�8���x���� 2��]&@��q[BJz7`h~�P������ �H�G,�PЂ��Ȏ݀P�u��uK两����}�S��q�p���s��L
���&:�F|�%��r8G��������ś���} @���׈-�P Z�T��_95:�� ����qq+y5�ɏ�?�l�3V�h8�-�H\��Wc�q�x�� ��΃��Xld R&��_�;_��e����=?�L�p� �XyI�o�������Vp�s	(��)�8 �����h�10��������e�(bhU ء'�� ]si��p� ��Cu�.� R�5TnɅ@��y��x�pM ӡ670�(Q�� �3/���VO��p�,l�d�Gj����/ ��hl֥Kz�$��8 8-P�{���� �g�/�+�`�ŝ�|R���\D؀l��� 5Q%8`���@��j�az>�pW ��H5�&�O_���	�V�� ���j�X(EX!�����_Ɋ��q:"����jE^f���1{>p�D�SX�ӝgGB4�@��Oq�3����<�d N�T֝q�6@d��O٦ ���a@�ҽ��r�/J���	<I(�� mTg8Zz��LY��țX[�!�n0ذ\�� ������ז�����g�	� ���U�i�0�*�na�LQ�}�.X���� ���\�5���K�!,�=ԃl�4�D�� ���}�v�[s����QH������ �$��� �7ɢ@n�5Ot��&BpF �41��6�I��+�k�I�X �1;����ϻH�P%�T� �$wm7�ɨt���3��� ��{DZ�;d����Do'֏cj*�z�\�Q�՟Z�|P�b(��0��aQ�8�#b,,�b;�$v�V{�8d� �L��Q� ox��mt� �kEj4�0��-� G�o@tی �I�&	5�8Q�TpJ$�D�	��p��T�����5U�����6�E�Mp� ��ȍ���v`�)B��!�$ ��u9D��S�n���#���Մ	�*��j;v����?KC(<g�w}�PM���(��[~iH�((�2����&�S� }Mz���U/��B�ǺJ��� ����BD���Y<:���hA7��OP�(T�E�l'� ��)\��h9M�]u`:��z3���ik�	�� *��@ P�D���_��莁fz���@Ӟ�b�@�L@;&Y���"J5�NI,�@@�G"@î�a�f'@�����[��� #�n' �E��e�@j�0yţVF�0.��("���gD#C-f��$!~ �]6� .Dt�
G�+�ZC��6��E���L<5��k�8�"�2D, smj�=*�4�$.�X���!��@9@�d<�@�� �)u��$Y�8�/ࣩ����.�p��� 	��xr X��e\�� 
�żI��8�l�)���	�����b ��35jng�z�S�)���3�X�����{� 6�2A�dJ -�Kֲ,rxc �G^�$�LAt aD�T,��]`�0^���  �>��j��<(�t�?H�TP) g��R2nL��fp��&�Ț
��� �\+4Z`{��� Fc�L�)���i��m�DD�L�A�6����T+��c��� !�)�� �? 9����w-Q� F�lyW�k�E@8~5��� (��3��,�W�!�!��츖��9���Rn����u�v���1�!R�I m䧙d��c �3K����8^�e'��`�`&�ns"(9|�@)c�Tﭐz��3�\�s������������D#���f��P��Qj�٪��� ��!�B��&���Q������$�m`�Y5 �n}�0;xԏ��j������Fk�fEAgB�L 1�b��&�u��َ�(���0����� �XfMSe��������r���#�����"��
�!�Ɍ�!P���a�xCB"I ��zMݩ$�ꔀhgÌv4P�P�H3@�}g�eV:O =����Q�4��ScDhٵ)����f7C 8%�j�KSkS@�#����� �� �}Lz��i����fÍv�� ���XdɊA4�S���a� ) �֭5b��4�\!k?	�a�'������Xw�Y��(�0e`��#�3=O��!0�]�f۔�C��P�� �(�e�c2��M��!�C�H�� �����ax���0�b  ����y��
�($� b�`f1q��p��d��;�a�x�0� ��La�e])-��y:X���;�r�Dѳ���R�ĥ��43�� i!���b	����X4 h��9 I&o\�7�)�`��8ȳ<|� ]
�M���� ��kUc�%2h��7��� ����]?�@l�! |{��Y�/:���D�]���qZ�s5��t��JH��V�8��@[@��B h&��_�Z,c�iM~�!/�_i�SgԖ�kj�� (�P8h7ǹ/H�!o8-��*t�L�%�e@�w�.� �Y���=Z�&QL$�}�� ��b�"aL_zy��!�J�T2��cP�#��|b� ~��	��Q�7c���V����8)��� ߬蜟% K�N����[7��2/#�u�P��ʪZ]� �@D9`0,�u�C�_a����u�����L���<K^�Ԏ���f�Q! V�/?�69����0=p�u�ӦHF�O1�z}���T�$8@ ��Q�%^>� $|B6��L׶ߗ����M�S�xfb�D +k�7Mam�����)���GZ :Ճ��8*t�� slB���9�u ߿"�-� �3=���%L�H���[H$|�V	�5
r�`���6��Y��N��R�\�ר���y �7�{������x@�p�_��M��e�"y� �M��.��s�< ��\�7���b i�_��%�S`��01��菄�9�&�g+P��f�q� �|~�<���?�9������`˵E�����=bX,�0���0d*���ZX"X�]�N ��#V�`� ��JGx���Hbt��a�/�#�s��P���V;)i���5���2Ĝq=b,��@m5���)�e\���輭��&8p$�5]�����G���c���v� X�ȋEm�	C�:��To{��}�p�H�B O��)Ң��
�l�Z-"D��y���`d���t�v�z�WYM0���i�@���?���d.X�AL���?h���  ��7�E�[/m�I�@�b`Bh��<Q�x� l@�]��Z&P�p��`���(l�L�I�����4�g0� �:!�:���Ͽ���v� �nt/��pmz���~A��7=�a���=8k0�@V�ht��Qg��xwG��Ubx	�� J�*B50�]90�s� �R�#������ ���� ���t���7 �D��#�U�g�a�iP�P5��')k�L�]|��f�\�9(��S=���^����'�����m��>�s�q��q�.?a�ۣ&�$� �i�\��{�w9�(�s��\���e��%�����(R�g&V��+��t���;�� X��kZ)� � f���V��-T������)R��y`0a�U���� ��'^G�&}h�d�]p��`���	۹H������	:�!h���N��J� q�xUp��)�(����5�g���)L̡ �	:=-�P��DԬ\p��3���ɠ��W���v��!��8v� z�|1D�CS��_��@�T���{$(�%0�ѱ�@2`P(����@F4)�[� ���ޔ܀i�BV�p�0�ryL�i���ɮ\�E���ph1T'Q�u�)��v�C�衯�ڠ�$&�ā! ]Gɶ�5��"�s�# ����q�/�R�1��[�t�0��$�D
`��!���i���6,|�O��L7
y?:�����Ks��<F�! z�=^\� �}�!�K��Px���!�<�� y��e| [�%�2���4��� aF>�[߼	��,@(]'¡��9��6<cx4k`H!�m6j��X�$�D�ǵ�M�y�
 �W�3<) =t����X��#�!�d�� �R�U+<�}-����Mo`0,���̫���P�^�?�A x
!�!�V}) lno�r�� �-�����1 �|;�
X;�� #�]���H$�B�c����� �x��)�s��:! A�^�"��}���s )Â��o��l�%�ഋ��W��J��ɏm�dw�D �;���c1
�׮������B�0Y�6� �����?jf8>vv �-�����$T2� ��Ff�5O �_��.��a��HĲ���s�X�=�b�Bp�$?��f�gOJ�{��1��t��ӊ�#�ϟ��T�1)�[���\���-L�H�v)A' }oB�,�z�	���� D��r�}����
�@�x��(��]E �^��+���0T��:�{9	K���p!l��$�n(H*��| �5M��*	n{. �ɔ�#�C�`�2߈�* �T[�"�K*��8 �g�H�6q o��-���L&T �H�E*�9*���eM'=(��2�]Ty��ʥ@)A��	k!4������@�ǽ$���tF$ !���d:1|�w�H��$R�'�������0DL����g���!�9�a�Ulb'g�aR�0X)�1:������[9(�\l��;�e9G�D>%�0���A�"+����3r�����6���_}@�F9"� BW}��&�X�+,a�.ۀ�i@�����h��e}>�� 4"� D]}�w�%_\x̄� �����u�5�C߀#�L�,@�D��,���X�|ˀ\����$�H��	�M���)<���޾�;��\0�ʰxI8����7��I�<�M�me3!���uu� �oPt�>����mEM��8�dekk7Lȣـ�g pE�=�q�!���0�ਔ�0���� �`�]���������c�#�<�e���|�#À`؂�<e4��ܫ~�����ݕ�i2v� ��5�^(���}9r��&Ŭ�� �$��w�����U�+�����G��E�a�?�d�R�0! �&�r����40�E$� ��R��C!	h��x�ad}��Q�D�A \}[?�jL�<���r�ׂ��5�(�u�!�U�-İ��D��d �r���CsOW� iP��\�H�P��@43��y#��4:txvM�h�ý����W`�ʧ#pn >��&D�p��D�`	[���/��$C���T��9����ñ�� �^��ĩ7rJ�B X�dwFת����B�c�*�T �)��Z�H9$v�`�v�|���3 !_��5�U ���d��(� �FZ�ʢ�g�5��%�K,�&��dT���1���y�&	���`����r���iUI�,����O�� ��3
�c�9�]�K|)����0t`Qܐ/��qȄ�Xȃ���� [l}��L�`<��ჽ���R`��sM��j}����P�4�c=�fL�FV�ʦh1�9�� �L���$�1��!��@8�Y@�$� 0Ox)���	��Ȅ�v�$�-�A��Լ���>�V+G��0��H�[�>�� &UD<��]��B���`��#���}�H��z���0�-��&8�D+`���)��8@����Eg9cв����54�8ŵ7΁�糅 ���)�Q���G�e�d8�����`E��S��)��8p��WPl����]�	�H�#w%�6� �<�:�$pF*|	����et�K�DPd &���`'�I�}n
m,�[���ʣF�"h:�ʡ�� QKo�+�md��2���">8��Oj�I���ʹ#�u^U��0�����">H�y@H���$�;�EZFƀ�̑�͸�=Q�y�K��$�l#o\f$e���O�)��iI|
�B8VܴZ 7�@��럳 ���|Cr
����B׏�0�R���>�#�M@��w	� tCO˪��=N��|��g��m
 w_�������0�x�������E [-��@8w��8��x,��1������i�Z0:�aa�l��P�b};�a�|XCZ }3�g���Y�O$�-"� X$��^8��Z20 $M�X�� h�F��RK)k�(q" ��>�]������X
��@�-�p�.tcLq���;����2� ��|��<� �,/�ƃrHLvtL����ԯ�NE����p7��(�@p0��yLy�uE��w���:��i ��#�-�4�dא��� 19�@|j>�~Q�U��p��;d,�\�$������L2��|�
t��U�����2�,�(O��lcqk C�P[d��'i�#�l�@B]Xo;g��Mi��hh��L�LT�.�����K�,�ﴻ ��e 3w/E�x�`����h����~z�� �5����e>i�Xx-�/��F�N,H���`}A�F1"��X}��O�?�w ��z��S_oG��UҠ 6$/�p��1�X�������;��9z� ���a���8�A���C�a�	�<�Όr� ��v��0��h�]���x�VhHBl�0���Sb��@�|^�=6o$|�{�*��6Z�l�M?�8�����|�!V��aL��� ���Gp눤����&�:�,թ���q��u�!$���|�ϒ�ALX��Ό Pp�7q[�/-9	�<����&�_�
�X�- �"`�p�����P��$��,�T,��w�D	���x�G�a���+)�[�*;PAo�� �d0�դ�L�������%wC���t�� ��
R����cMK̟a��)��q�@�.:9+)7 �G�TTdď <lL�5 �7A�k��x �_�T��4�d	-3/��%h���	�kZ�  �^���%���H�l��E[�W�/#� �k�5��\������W	�l�,	���Z�x��Y���р1p�bl�5 ��f���F+	��@Gz࠭A�3/�#! pb��S���F�ix �jL��:��:�#� /���ݡX����2\�Y�0c}<�Y�̀F[}g��	�OX�	�[�Y�o&��U�D�����b�Y4�⌀�N�i�����Y�/ˑ� ��U��C��&*��;���E_���{<�H��~@!����P���z�	�<�p�,_B�]`�����1 ���U���T8� |�~B'S����Ջ,���n0!l�-���H�T0��V가tF���!���U[�`ҝ5$��&s��`��>����}��sC�`�ٴ}�������$1�dP��P�,��&Ɍ����^ O�羆p�����΁�m�3h� �����Н&��0O��WQ L
ɞ~�G�Ҍ3�,[�Yu��G�
���~��w)��� |��I�.$�4���Xx���f` ��` ۡE��Ǝ�Up����̥�Y}�1[q���s���0,����-Ղ8� ������� �e-[�^���X�0p=��� ����}��޶�Dc���9�1(���,`��9��GM'���O�1��:�h�,Ҽ�\F�X_ lvU\V
�M�p��'�����'#[�8�G����$bX-L)�p��%�2�,i�m/I��&����⿜���[ <��� H.ݥ�x��ߑ�_�R��#1�^) �1��y�Ch�@��.p@:��T �p*V���`r'O��p�X�o�H�UPb<�n�K��BG.v,������y�T�@��	-7z$ Li�E���.?
��Hˁ@N�/#� ��p	����w�� ���M�������,�K���[�T?�h\:Ď��t�~9�dz�g�����DH��R@6���"� N��e�J�Ԕc)Ɛ	�-3�"�� �~H�+���J�t���m���5 �����R~�~�R�� *�?$FD�b`z8ഋv���`m]��r�e�x4�MH1��W��,��A. ����!p�C1�!��z�Q�!�~�m#�H���3�1 ��=�@�°�C��zw��(� ��-Wq���]s�
wG��?�%h���]�� ��C�(D�G�:\#$ ۼ�+;
���l�Ɛ�f����4U���ɯ�H�G�ѮX9I^XL 3��?� ��}�� � ^q)$U?%���"lY�#��X��� �NsV���(�:]� Q�#�`U��~ ����h"��\ ��~B n�&�]���Ю�S #&�> �[}��U]4����Vy��>�u �3~��I`�{ �ԿU�>��HV��H,���'	Āl �u�]�/����+�T��k�G��9:�.x-瘯�׬xf8���\���� p�-���(�W�,c���`
|�� �q��v, ��uwM=Q11j�zN��e<6�˹��Z��ú=���@uA�/z :�L�c% �>"��T;� ]�<�}h�>� U��s>�~8 WJ7F�x�z� ��=l� ���_s��|� t�=�`
��p1��ܠ�z�; '17Ou\8����A+�,#��H�!L�Bw���SF�˄�yv��u�1h���>� b�[t ���C���� ����UA� �W7 �B� �<1�l; �}뚄
�n�C���_ ��<Ot��~c �=g�����1 ��������<�|;��St����Q �7D}��aOv��� �~G�L� 'Y$�<�� ��M� u6+�=m@��v�X 8Ϸ{ˑ�t h�a}+= ;��@�B��` :=?������O`��N�����k����� !��c�v%=i���(�Ƣw<g���k&P�
�G�Q`�> ��~���r=��<	tp:;[\���ʁD��ăv |+��f< x��)����7b�#ѩd� �ve�����<H��u������X� ����Y�$�t�<0�v	�^*AԾ� ���H3�I �=�aW< � 퉿���/M�Y M��}�W|� �=I�X�;��ۀ�nt� �u���}wv l<q�m� ݃jo��|I QX��b ����<V��>sY�������\
��>�ؾ� m<,�PSVY��Ѡ30P_�� ���Ù9 `d<>�:� U3�r���A���<��u͆H�L� $D�X{<�|�Z�����$��1 π]3���	����4�> U|vݸ� JWB=w�����$G �cv�D��<W��\ A5�s	g�6�+�<�&��Yɩ�~���@�1 �&�>ui�Iz�<t�����������M�P,l��;��o���s��Y��Pn��v~1�4���v�%h�t/V�	wC� �\U����$�7?�� H<e-�yt<l� TXob,,��X�� �$Hz D�tv�<C4r��+�Z@����;�@�=���t�L<GZ��A ���n����I�=ul*� ��<o�YUW j�S
a �d�x�Pt,����<���� �s�.�?�����+���4QvL`�	1ZB��A���$p������_v �j�ӎ=̝�x	m�/�,d�.{J� �������S)��^��,�9� �.<E�Ax�-�`*�V�������\��< .���xwHF�D��u��q�F�{ S=��%�G�Bu�`�~�Nv%�pY�<t��쪣��o7H� �-��/w	�ȓ X?_� �r.�]�㝀�x�2��0�N�m$_�h M�����ŀ-�k�1�v� P����0�gT�1�$� eȫ�7ɔ�� �<yw�Ր,I��)〄X��d �yD�v�?=" �?����6�<� g�e0 z�K��<Q��V������ y�$sg��={��f�\(�&}:��3� j�]{��H
�y �K</	P�T\L��� 
�h2�@ ��7̲�<[�sb ���� ���Cc�6�����=d�	>g�]�`�h:��ۧ�`�eT���<#���@׈�:c-�uB�`/�<h� H��U�>��C˄��d!�,wT�v��ǘ� Ob5|�P��B����O]\s�=G_:@p5l ���X��� ��[���v�=
����	�y�T5��,��ro=�χ9z����+�Do~ib�s���N� �V��=y� �z��}������؄.�����$=��1<d=���0w���@Ēor�c ��;���_���[��ȡ���!�n����p�Jy���$,z��K� ��u<��~v��L�x��渇���� >�c�:�ԣ}v
�&$ <'�5�sP��H�4 �{�rva ����=9Pj����ڄ�p�#.3��]� �-<&Tf"t���Y2��8�`�����<�-@�\f P�n�T)1 �=��|/��M����\� ��@f�&���� t�[vp�ԗ�`��1��D\iP���t��Ҡ]��=&k��u&�X� �%��bL���1�pZUH4e_�Ԛߘ�
]U  ��$	T%��� 7���yr�U���aPP:�w&΃�j���3�����M�`L8E8�	+���}�=~ f(�pj��	�G ��S%�=e�� uc<H�� ;t%��� z��^#�"p���p��<Pk$z5���=���4�垀�t$Ψ��;�?�ϡ���i8EO����^{�@w���rŇ~�^�]0��y8=+v� �T�;<��k��˃ ��d箠�t�s�r�<W�Dc5p1-B`UF!�6�"��6<|�}w�Y8�E��7+@��� W�t��:q|�� ��L� �X����V�M3z��}5 �%]
m��A!����4 Gu3B�+8�<�n�
��Ԉ\���	l���\�	N�0KDsR�pD5��y�� �-Tާ2m/�Cz���a�Q�w��.�;Y��54��`,��sv��:oL�4�t`	%~0l=`�2|��Ί�o�ԗL�v���(0�HD/# 4V�vO<�g�d?��L;�Ǩ�,μ0�sE=�^���d�� �Q%t�]G	H �WNE���T�4�7a,�k� �>B�֋Ѓ�<VKuH�����ag�po�0�<�4�rDѹv�`jz>� �e�����v��}4A A ZJ=k�MV�?G��Qc��t
���:f������@I9\:d �PO��T4<�=E���#�x�� :�_`5I4 ���<6���~��hO�x�(�	��f� ?�H,:�	� �so�d1��\�M��ż���*!�  �`���S��� �<U2�{$v� >�aud
=�+Sip�|� DOv�w[�0 2���si�+D�t<������X��V� ��E<����w�U�c�į���X�l�@�����8#�^\Q��l�!Ԓ=�:�A"J���]�<��`d� ��Q�Ӕ�],���M#��LGy 0O����9��$� $�C~�¿p���Z�� ,}9
 <�4���x� ��E�x���V�����,�.�ed ��]<��r9?}	�J�x�@㏢I:�� &���7�T$Q���IE��L�x�v�%�t�6�
�d���+] �X�X* a�Ӑ0�t��h�v��� &7<B_M����"a��@�w�*2� 7��L��]Yք�;�`~�칦�@�}t� /�q��A|RY�H� i{��Pv���s k�7��m*̈́ۃנ`-�tFl�lv"0�~b
8?�����h��p�ف��v�
���m<��w�R)��u��2bp�" `3��s��= ���S9�C|X�$z���5�n��&�0�cW��h_��/��JP�bml!�ణr��@�%J���$`; ��(&��: Z���v�W<�4o 3@��)� Ƅ*���y�5�#P��%iw@��#� �<��5z���{l���VЄ�����2�@�M,l����F)"r
 n����u ���A�\|� �=T�Z���<� L;0(�#� �z��
|<aY 3��섚U�����,@y����~<x�4n1j`�j>���
P �+l�X 8���>y<D�vC!�o��-�Y�d�R� y���<Ig� LW[���&=� �J��{̉��=@W87?A˴���z����vP^�� �=*��Ԏ �MϾ��2��e�l �jL�� v~�="����8�꣙�z 0�4�$m��$n��W�ݵҘ��_�%�`J�� ќ<�϶;tHWP'T���|��D��E�-�@��$ �!=��;<R���{�3W��ɧ�d 5T+�<���/z�`bF`x}�.v�;�'��M�~�{�Rƀ4cr=?�w�����s��4Z� z�"=�+6� V����8H~ �j���l$LG� }z<	�Ǔ	i�L@X�0s8��� V9�{��v[��(��,%d,��gt4q`샡�=�ˑ�U��\�c��F�= ���s�<> TИ J7��ǔ%��<�Z 0��u��k��T"i� ����ӳ����>&u�� Z�AX3��
��w ?�z :7�~@t�_"��P,���z� K����o�<{��G�?V�}Ѹ�,���u(%� �6�w= R��:G�o! 9l��/�`� P~8��V࡮x��_���s�N=�iA�:`d�:ڪ�|L6 �[<s`Pt$zhv� �cy��� ��T�߄:�&^�=m���8} �!�]�WK��p��_s@٘<)	5o��ݒ�{(xNLT����qv�E�`_*S��k�	�
��	�3I� h�w<�;�4� �8s�GW��$~� ҏw~���s (�<"?E��=/a!i�3`h� C%q<��=e��̀J�\9It 0�y$�]��@m�s<:����΀��{	�	�S^��h�wH� ��y���|��� �9��e 'th�v� =3�٭S` dۺ�"��� ��Up״�@y=%�t;H?
&�LX����l�`(�yv O	]�=J� e7U�,0t$��� .�Y; թ�9(�d< -%�l�����[��4 �]ûG���vx��_a��
���=�< iy���<I&��U� =���:!�-#�\+�O����=�g�stw0h� %Tua���Z���r�T5Ii����<��6y|������X	ǀ�g
=w �9�siT��L0� ��
M�E�( R���׿=H�p �.t���:9Xb�����+��_<(�/ ���6 ry
��w�|d��.<lj���JF @�M��u`�@��e�ȼd{	�[���=z��D�y��Z�7;��\�� g�Gu�B_T x���<^%�S]#�[� �E˯�p%�����va;'�	ս��x�`�p��)�{�p� �=bsN�t%=�Ԁ" z�B�P�=.լ�ulI��G,Ż \t�;M VP��%87,�<l���Mݓ��ى�Ӏ�
�N}����=cEЌ�v8|��%�l���e�s��[N���Z�B�p�)��;؜�1���A�N �: C��o/����8��hvwI�
�<!�U���XG�ztP+�\��	Hv  -6��sÙ^0@����m��Y���A��K� `\sT7t �<�3D�;z_�`d�)�����av� �C�f<�)�\���6�$�����~�h� Ju��<*8?�����T�/$��A��+�	��‴Z w(;e� ������0p<���bD7+c���`�p��� ���=��: <hH�;��ظ� �u�D-/ 3i:�4�v T�< %1sV�M*����Ӏ?� ��ʟ<�y ="������m'�S��1 L����pZH�=0�|k��CS�-����H�u���(pD\ _B7'�m늵	8��&$�
�����|�}����(E��U������'Y4L	g�π�d�v�j�Ɔ3X9a���@w:�K
����kn�t�����0@� 3%aL�ɴ�z�]��:Ǭ	�u P"(��m�D50�g �vZ��f
'�4 �DQO.�(��s;��J�g<xt>6W�S��8��a�t ��zv�<�-e|Hp"�,X���ј���9�RQ�lXdHh*��� &+�='xO<R�� ?M�΄$��/�P���� \�r�h<+ a��f�|�e 7ЄW%�+T>#����=ؤ����8��y� ���:������\N��cv����MSül�����p� �k=#�w1Saܴt�7�Z�U ��<�p�L��, Gt�v�ݍ���p��`��ZF�����:L'|@��KE,���`F�v�=��0� R�ޱL�e�&`d+�$?���qlH�d�, ���x�; 7��d�q�p
6�f�&�0 ���dI�<��x�`40���M#���|=��"{8o/�'�(�H{k��z ?_S���EB�Al ��t�� U=a!�/�}�}DK��3sy :;���Iu��HܾU v�a�\#� i�%$+�=&u�� Q�P<X!�_�F�|�)K�g�@������u} � ��v308�&����'G�k۴�5֨�>������H�6أ��r�|x${} 2U<i�K;:�L,������9�6���^@�&��Y� C�8��"D���_B$b���hZ�a�9Y·��H"tI�Z�=��U����d6�DC?�p}�����h`�������xO|B ���h��<��N�ȃ`���h�ԏ �L�Y6p7TD``�i
8����x�c�Hmܛ�� �{�<HL�� u�]�$\>�;��w� ��<|�0�W �-�+Ɋ��6��4���h:��=�v��!����&0,�P;�'�@`�8�����&m�,�:��Eɫf�u�8=h 	&S.lWńn4D~�Z�\=2v; �Y���\� ��� @�:���<|K ��ц�=�I c���#6A�&�x�y�C:�9� Tp` �|� ;G�I��>� =v��i�����C��c�<L],7��� �n��A��ɇ�y��@�R�p�.6��wu@Z�C7���X���d�SN|'Vl�Kt�����:�{X�}�,[��`av>E���^#P�K��A�E��$qRT$�[�(��n` ���
���-,���t�� Ù�0�=In����׈��� �E��tB+J
��<L� ��󦟱��(;� -%۫�@� t��=$$�J7 1>��jX����.x w<0�t2 g���dwP�Ex��
��A���<+�� �d,zܙ�!) ğ�.R�:(bq��� �T �D��O���� �����n�R�8`�.d Q,�=x4Cz�`�- ���M�' Q��#^Ju Tw�=����N��^d�Q���8�7���( �u�|<m	�;�z�\��tWk (�6^�='��*�x0x
Z��1���M���B���S>=�'����t�LW�
���w��Z�� �x��-�/�(�։�<w3]f0�F>v+,k�	=��w�_J�a��m���vT�8)Zl�P@s�#�!��W|����� p��l�<
g �M.��{���N�?DYi��R�D����C�b������=z���R<�{wL��Hy���8tSLn�>	H�i�������0�d�����0��:�� Ykn(t��8K�!Z���}� �xT��v-=��|jՈ�$G���|�>�<�Q��c� "�:� u��ӡ/��磳�0&D� �P<s��}:	�-��KcYJ���'��@�~�<�LWC5��p��8��>E�� �)�K<p_���Z���9�ބ2���e��u��pk �v�Y��>�7���Vu���=�|��54ڌ8�jx�wL �'- �m$�P 1�O/%^P��aH<k � m&
���Pd�h8���DS9/�	�â �=U���v���J��}?@ �8���Č�� 6�~������y�8� ��$��h���6d� ��>IX<���Ľx��u�TnJ` �7���=3|�������#X+�>l1��d�:��F�:<W�-+���LZ8����ߗ�N �=���<'��$���c�B% +k:�� v�	=�/�j����|3W�����rxv��S����c��CI9����ӏ����ɛ7�o�~���g�EbQ�r�8�$�U, 5@���0�<n��,��n(
�� ��d�����]�w<(�	�:�+ �Croy� i#��N��!����t�)<B�&~_`����t �9�� ��Ja&�=8�\o�m�<|�Ԅ; ������_u,�D +:[e|�`�\H8 �? �}�-Lp�<Hw������]3%�u��"o<r��
=q��e+��w�5ݳ N2O�$��.>F��]��s���P�a)6���� &�	aO��*�:�N ŒPτEͯd�)�w`�PP��9�"}$����OP��3�ȡ )%��}��s(�*�P��g�K���y��#�t�%���{K/p	ہ�>̧��������@�$�A�({��� ���� ��D�Y;@??I@����	�h���!,�3��(�8B��1A��  ��*�=����/8�A�1� �5�6���E������c�3 ;�����Y?�C��'�6�� r�=U�9,��X8��Y:� ���f5�]KOT� L<���Q9\Z�2t O �[o
m �^�'ե	�����,89� �q�0�l��f�nY��׬�5�{Pw��2S��]� ������wv���x�x���}	::�0�T �`�ż �Q�Gj+� B�W�� ź��-����Ru�(�gĕp�!�v�{� ={�@�ۗ� W
w~r�H� ��y�E�� ��6[$��#�o|��� U
>��jI�Ҷ`T첾(�V�U(J; S�|�0��/L� ��a+�0l���Ԡ�]eag0$J��a�����p�B|�70��߮ EZeV���� ��1"FK�`d����S0Ջ).N�0����C1���%J��\�|$}pL<�E 3�x�to��U����]�^nR��.˕�EK�ZQа��m >'�h/Mu�8 �rFQA�GN o�/v�#%Տ�Y����?��u 03n��+UP�Q��� !���;-�36	�=!s ��3-�� x��^P)%��Ѡc׀�oh�"�S���x�A,%� �!�(���9ZĽ&Ƞ �
8�0� p�����1�TD�O��aވ�B<��3!��aΌtF�j�� ���� ��5���:U�I��� �H(�j�#x�v$��-\�M�1$��̄]���6�z
Quy$� KR*و���#���>�����dȇ�t�ը*����J�R�\^��jn1�b%� �r��s�_�I�x�)I3����.���t �m'y��y��(���QC�t*ix1�6��F�C�_��!� .�^�f� �tĔ9��2HA�Ƈ�̨��`�4P���QW�.���Vm]^��L�H\�6��P|�`�2~���(J�"��Q0B�20��Zސ����usK-�I�� %��w���Q��!p�@\��H~Є<��K8��į�Ǹ��"��N0�	��0��;�Q^�D�< 3�]Ո޽0Ҋ�J1�X�t�`���`�6p-�D�z���?��x��`����d	M��!���_������W	�ŕ��p�|C\�!ag��� ,��/^�b 
6�U $OvlIX�j�y2 h��O�
R�ڄg�aFd��@�T'6_0�{!����J?�d6nV~?�M�A:�#� .KY�N�qEY�$�>\��X9;�9�e	�,4� �UŚ�����pa��j&%2�/�(��dʫg�����E�@����PM�$�|<`t��Tp�ළ ����( �f��i�y� ���2�#�� �</�=O`���x���~\��qiS���e��!Xw���Ɂ\�j^f"�{`v� _q	�װc�-K�`��2t���1;tl�E�`p��7*l)Hp9�Q.��@>1�ѹ-���� ���%��`(��ʿ-��x&x2��e�Έ!]g�E��Q��:=�D���0����A��vs#&Hl:	�Qf�t 92�v�WP��)!<�5L Q��@@�ʅ�7sX��0� ['t�{�b�I�H ����5^v�1ԫ�&;�H�TĄu�Ll#0��`ޠs����p`D-�Q�X�`�ɇ� �mk��_����y��M��d, �љ��M� /��KD�1n�Xk�b<�,tF�ȸӀ��X �bZ����cG�鿟����
�{�Sp\F3oxn<J�PX��D�Q� 7<�~V�-@���q+&&�
ϟ���`�~A$�B��<Y�	yւ`�A���:0#� �6f���I�@4Z|��4���Y �v���LhQ �����9`	�-��"��trH �DU��P����FK@S` ��R]��6D����3��[�8�9@/��D��%�U:�F`4-����t�$�Zr�=�g�{&H@X�$���tFL �Z���pF`��.	���Dr�x\\%P��0��$\�P�(��<_H �)M�G�@k1��p���_�z�{�bH"4��	�־��,5�@$�8���6c��;0�+.�5w�}tӈhQ��Ht�#.��^�pK�
� ���y�;�d8�ŀ�w�s��\���K�X� 1��甌��
g�w�]_j��bp T�9\	l+M��s����w��I��Z�%�����X�@�W�[� (�E��8�1+M���huΐ��N}L���N��"�QoX�0L`�ԙ���C9H�|��0�E-��m���*�3�L�����U(}�|���M�@gcHP����iFH$���؞9 ,Dv��y�� �`��ISb{��|GD�`�p�'y��|!�c N�=�H�Pm�a@��0���6��y��^��F�b��jNQ�`^)�L.�l����U�x#SߡF��aEUހ�+�}(-'����&\M	��(�
�:- �pv� �wTE܃��Q�u%1����SKD�F��E�c%fQ��Z��xf8'����z2иk-�Ӷ�j�## ��0a���AG0g�s��;wH/�!���#�Ve�S$a߶�����E��̇\P�ğ���$�Y�yj0��U���3�\=����Lx&��Fe�g �Cw��$#���Rg`	��A�e ���#/� �����	S�.@Ed� VF� ���Hk\`���I�@�����ڦ[�,�\FNv<��Su�E���it��l���;��1������D2Wܣ�ԙ��Ӧ���K��~.����@O���Lɐ�.q_�Rg�D:`A�S��2[o{|�xQ��z&��r>�k�\E���<K�	i��Q?́�?��!sx�Ϡ�#-U�0\ľF	�@�8�<� [V�5H��	ܒ����VF�w�d��<�����~�Yә$���R���v�ʨU`^~���%I���F���X�خV�3=��9[]��	"�
�i����58yK�MY��8O0�.=1�(�mdI��rr�'vs5`��٦�Nl���h�Y���VF���0�3��s>	m�IC��Y�(T�7�݉]��~ˀ�԰�9 ��Vv�j.�L�BʹB��; ���3W��v��9T܁�|���˸���%;P�����$C�n�L@�p*�l�?����>�H�����S���^F� {� @3N/C W��U���XIL����'��V[q�0�]�抗3��}2�eE���{�9� ��}$�s�j&�# �oJq�������J>MI��Hݑ��9�^ܰw����`�s��L��Dg����qW��֐��� (�|>�9��1��v�P��������b,��	���K�+y|SP%���A1k-W�0L�� �6��`�~���& aX�Ӎsy��������׉�r<>RML�;"2����������qT5�×o��D���i� #��5�y�\X,_��3��;���fP"���`ygٙĀ�^%��8�0 �J�/�#�Mݴp<2�,ml �N.dO/9� �<�� I�좛���$��<��@H�X���
����m$a���� (&*� �K
xvM´��5e�:���^�U]��	@�C)������2����[d�ܣs{� ������ Nu=�i�5IK��l������~�@���LE��.����,qz���DR`1�yd _���'�`��3�̈́K|���x�Y��Q��3�� �]K�`��֮( ���3#�N mO�Ϟf�("��*��� ����.�JR܄1���:U�0�MT��x3 ���х��B+�,�"�6����� -��ʩ�,F
�<���̀V���;�!�l��J��.��\	|!�#0���9-O�,�y ���Dȸ��U��|=H\��$�h�p	� �&���zC+VR�I��70	�`�@gR�q�༐�&V���Hpf �bI94��
d�|�1�jq����~���	M.�`ܽv"�00
�An.�p��%MBI̥�K�Τȟ�JG� �D�Mj_��>������� �V|$��{:���+W���M!����*N��.b��Gނz�vhk�LAd�O��C��k�E��$�j�q��K� f����\*_M��B�Q8�:�L)H<0�9!�mq:�%���0�4 k��
w+�Y��D�b��,啥��\[��jvE�c"�C�1��`' ������w!�,V��|F�H�<j�2����S�\|	��S���>(J����:$o���`U0��
�9J ���!-� ���D���3O�H�ň�'�y���<�YC 4�jIò�淞#�����UA\������`��/ߌ��|��D�`��eݦ����lR}�[�K/#��i���$��Y ���XpL����8-J,|t ���L�r�M{�	�IW�`'��x�6�Dh[�T�*?�vp�<�j������1ڛKgUaԹ� /W��3(\|̀��Y	9ʁ���
��� ������5_�;phLNHk �+R6������I� ����|R'���i��`:;рe'����P氰])������Q'�2`l`�Z$�X�gj�[{w�ʍ
0��@��ۻ��F�P��j�H0��,W��Ɨ�����S�� MX�.�)*�w����0�� 3-P��IK��U�H`TF�6��\"���_kB�.�P'}��CD�7� ϲ[��=�ņ�v�*X/��,�䀚2S��D~�ϠG,�5W���ە��~*1�5v`
���^e�� ��G ���"-Q9� �����G'_�HQ� f;�w�k'� .�Q����܂9��Ĺ#s�g0�� ?BM>-!�,_b�h�[0X�T �-ω�+���4��hp:RL�!�+m�Al���[� *��`�{K��������J�`�B���'1�������,8P(^F��"χ�SL�D+��@���y�dP��b
�<����:V�HH`�I�L�"����1?Amv����T~`�1��+w9������˨�7�b�����E�f%x�<hl��& @�K�� ����D/5�,6���z8Y@�"�L�;�޸ok���,5UQy�d�<$:�,܄�5vV�����?;p#� �=-ХY��F]}�ZTtރ�e!��z��b\������ `�%�2�ݘuJ��0H��y�, ��/ә� ���Y�ܹ���v%	�KQ�<H�L�'�@� ��M� �_��i`]�Ԉ���U՘�,p�����OFi�D`�)#�&��3 ��z1�6j.ߚ(�S�G�DM`E9�a�j!�,���D�S ���x��)�����^�`��(]������
��I��CA� �X�8���q!���S#��s̀Xi���$-J$ `�X��O�u�DǸ��ՍL����� Ȩ�X� Nc�41.!"/�JXM}��처0�s K����_\�<��(D�a��ZHl/���Ŝ�$���3�s>e�c�~:@��vn�{N�,�L����7Jy8½NPM���,#��]�iP (;N�rtI[(X�� ��[j��儰�J�SݲI ����'��$�oA��_�@@��S
����$�<!T����$�=j@�
V)x�Ѩ���߸�KnD�L�y�~�eo/�#��L�"�`�ˉ��If�����|S�_���$-�oż��c��9�T���E��N`�y�&(�v
�����X�`�5d"x�x��0�r��}������.Z��U�E�=v[� ���=��i�A�6�h S{��y�P1=���k��BO��Ĭ�����1_���� R�e�T&�E����������0\�0�a��,"3̢�0�h ��݆�޽*�	����p�$��@vFM �j0s�&��1&SΤ��K��٤�NQ���e��S�f	i��@ܻ�IZ3ĸ�4+/�#g�_��P��V��\( ��� \ȸ�ĐwNs.�#� ��
���B�\EŐ�=��^��@�3�Tb԰}� ҽL�]��XV����Rt��0p�����7ԴqL������$+q!��0@(��w����,]ME"�H����~뒦	�+x�	��Q�\\��[¨M���8D�`܉� �g���!�_	*�(�� �ŏd+���� ���C�{�$�����3@5�W��{�@@����C<f�Ϧ�h10� )��ܽ�h��;P�����@tT'�IG M�i>S��y���x���� �ܭ�+=�@C�d�g �{΢M� �!��q�� ז�~��b�x-�	� !���J �O��[�@FZ/,#� �Qe��WXlo%�<���h��fM�Qߐ�v��:\9>�ω	3�p`�mt����Aa���Tq1^��lg͟�� 'b�=�� ��u��˦����L��K��I?�`a�3�e=Z�T��k�:�@��r��:ݻ����6�hl�u>\X�):�@�ªZ,q4��������X�����%\��������ܖȽ	]-�u~������h��a��I�Պ�XhO��<:�#� �/߽f�q������C4��L�6�R����4Qm�^ME4�T�$�O\��5�h6 +�I� ���4NgM�%�e ��dØ�Q�4��1�Ȩ��z~ݽ�l�1�_�Ө!�	�Ȍ`�	�$���q7�O�_������2RK��%.#� �V�ý6A�4��x�7,8���^�є�0��nm9~R��(��04�I��̦A �F��H:p#� ����{f~ ��UY �>}�����u�rC�H��9����җ� ��9cxSP�D���~��ɿ��/����\a�@��9g�ң�R0I<ŵ�Q@r�:�3	-��)���D�? Ě|t 0T�q�\u�]4"�|��fd�s�,Ȝ��mѠ�e��������`�Ci �I��ذ-(�ѵ�� >s�,�r/D ���]�SH3U�� !���K<B�t�rt�%[3 ��̸��v��J�!p��S1 �BmP�\6�>�)�X~���,/���H�d.6��(�3�`]!�&6�T��d@_0Dp�x:����<�9�a��l�(�)���и�bF t���=B������Ei�_*�1
X�}w��T��$ 8���#��?�o ��4^G�\�>8�dH+`���#��Hy���z�V�����_4�����/ب����0�v�����h��s`�!����\�*�#.� Q�z���g%��
���X�26��c` �*6���Jڲ�E�ua�2A���/@���Rg�#*��Ѹ�8�u��m딽x���N��H�g�S���0m�(2����z14A��-6�� �YC�%6�MW�4-�� ��ۻT�+԰qz�&[7��b�� P�1x�2���]wS[����:9;b�
<+>z?�O������kK����E�#�j/ڹ�"`�0��ʈ���@��0�L�08�
��O�D�g 6��0�D[� '6��sc1�1m����P��ez �H�2�4%�Ug�.?sRd��]�1��� !-�M\;��j�� J����q<��P���lRO��#��9@Z0I��������a��@��8BA؁�W�2�!� :��`��S�	G� Z�� �e�E;5��m0	���k:r3`Oa���T>��L0E!pY��n#Gq�ˏ� ���%e?3��������:��a�R�\�[�������@�������>�B1�3� T� ?E-à��r1z���*��XC�`3(�i����
0���wؕ`�6sF�!�E'��8�/����L �>'m`�����tav=@.����n�e���'�X8%���z`/tr�(y M����3�^�$!OqM�Z��>�`%�" �3F��/=[��	 �u�,3t� !͂�m����:��� �8�oP����ԋ�@��S	�OX�sha��p�f��|��u^� H`J�i�y�r0�%�jY9�qg��s`c��S
Ơ�߀wM����E"�o��� ����A��!���伾I �}=d�Jx���	:����w�l�{n��݌uM��vb!"Km�i���Eq�>�����Q�� h�r� (���m�T"�J+��Q!I�Ԑ�Q�Kl�n��o��e��tbI/`]�$M7 Q�P2�!4�?� ���h�#�
�H.@{�"8�C2�[���@�?eH�H����ll�b��F\"K qZݑ�� �7�,��8��r�x�J� #ɭ4���T�g싂_0��y����ц�I����}��D{��H"h�0tM��Fn" JlME��7?����5A��3�~�xM��Q� �NpM2�+1���6h��%!�����=A����ja`� �L��DDo	X����5��u�28��_�٩3�"�*H�>� Q����;�#a{�+A�e/�`EHb���"�0��g�Td4@a��<�	!�с�÷���LѢ��s:��-�w�:R�����K0c��!0C?iB��)I�D���4�sM��f IkMX W�]*�������b�!�S�2 \��,�|� �خ�g��)��.�àF�hF���f��13`����4u`0�m�4cEM�����W�h7x�A�.d#��G�()!����5p�����J13�.���"�s���$���� ۭu��&�3
r>���'��� ���T������� d5���������Y%N܈5�錗 =Ì��-! �C��|^ZFz���[��n�`��x�|�! �ڙ�U��(p� EG���a >�m,0�����c�F�"7�� �r���ICs ;98����R�dY0��s|9(���S�6��'��(�iJ���4#X��rt ���\r8!�tF0j�.��X`5��<�x���#%�,F4uu��M9� i�G��ԇ�����^��x#��Ѕ����e|s%�
���x�i������� ��8EP�|7�ƬA�ᎅȟ�1�,���B`$s���-h��90����"�Ʊ�q����i���zڹ
�yr@��>9t𓺸� �#@�0%���|���P��r5向6��Tm`c��%�d� r[ݔ�C��\~�e�ý� ���z������;	{��-1#x�104� Q��޻��F���u0n�{� �+���?H#� V�:<-EI�N �P�i_����?�$�:Ȱ�D����\FF �����IGT	�6~�X��k�JB5����P$q�� /a=�!\h��K`��H�L:���� )@p	R������a1gMJ�AP��舑^�<�HjM��z�� ID�3�s���Fqg�鸄1Gv_� ������C������(:�� 	��2��=ט/p#%�<@�X"h �Qj4,����� ������	���Ⴠr= ��{�k�(�����[G�����* ��.�Wڕ Ơ��#P�\(���� �"��#�T��s���� �׏%����� ����x�kqp�Z��(�3Ğ ^F$�O@�`�2��0!.�)�q�xՏ9�kK���$c{����U/�\������e��Ȥ� ��)<��?$t>	�O�� �9)��t�m����s�0��`�5HZ�		g�d`7l�t�V�
�L�<z�P?���4���Y�si���K`�%���c;�\?�#�a)(&��� ϟGL�xZ��t�Ġ@́��_+�cH��wBO+ts� M��[����zi��6s<?15tL)������)�p�͍-����r`7Q�eB� o� +g��.���H�6 蕔J�n0 �����&���.[0�ڸd>h]`��w%��τ�%s+�&T\FC�O��$�e@ߕ2�j�Uf��G1-5Py � �gn��hv4X�s� ��� �O`@�F�}���Z�ߥ� �s���D0`��<?�
��GY`X����,s�^F ���ڀXlH�po��,�K�:D#I t�Pj^:0���}s��(Ǭ/ʝ�J�8�[� N�pH-E���$��,p<zC)*ki�N�P�����0�U8�؀z��aH��	e��Q������ۘ�Re�#T U8�Z���i����-�[ h��y�&x빀 w�<*6�%3 ?�ې4�h���ZZ�/\~����:c��H��	�e���8 _��oP�=G�,4����	 ��a���gyP���9��U��s�j�|Wi��J�E&�, .��'a8�	on�cQ�yK(�r��}��ܶ K4.�(���ӱĐ��8�)�� q!R��%�E���+�~x:��e�5��_���z&�6���xp�(#�$iɆ���~�oe�9ŷ�@�/:�D�\��觌����)�=W|?����	��$K �/@H��-�������ۧ�Ĺ� 4X��cO�`�=#�x�!�<��)El�` V1�b�ɉ��4��SR��I��%`��nz�GL20$]@!���/��:��Ĥ`�B�	�|���`���9��l"gK��l�Ps��'��(<��C�q� ��L�7�p�(��㤐���.n �����b�_��)I�$��Q[ ���f$�N�İ⴫�8�[qa{s=H hp��t��;ހ���'�<@��aH�,|@>%���`�`y~"Й�xh�Lo�:����\ �i{I�m�`�w�(z���\R�/s/l#! �%�u���K�<C'�)�@Ǣ~��ϭ�r��00��˸�3�z4���68 �~B��9�')� �<�2�|��P) ��R��
���́����!�/k$iY�cL�P4��x���ѥW:� _ A�ۀ�kK�.y��,\�6�Y����4GǨLـ��S���00M�\\% @}��� �v��٣����[4P�9z�������뺽۴|��ԃ� �G��sw�� ��˧#px �R]��/��H
}��0��������En���|:�?����42�nQr�䂎x���?F(@'Y�c�y�MX�X�9�I�L�袌��3EA�) ��YV!���8)9��2���M %���
���v�yH�0�= ~+�xݫ	>�����z0 U 8��(C�HT""�k)A �g� �Q���H05	1�+��scgD�G`5.�K��8��+��S͉B�� TS�/���$`��ٰ�	6�!]D� B���ļ�L����\��c���H@�8h� ���m�W����Ih�s|��67Y5��&��)�� ��D��� ��ܪ�d����~q���Sm@ft��x& TI��r�p�[��0Ka>R��1�p�q@+��)��{���X�Xz\�4� �Do<}�I?z�"s6 z�:��Ԑ��|F���0d��?���j��X�	f�r4��qr ��@Cs����$���4J���D��b3� %5Xj��$�$ؓ�2e4 t�A��,:0�tF D@�䏓�2#YPr�\c�~���z�n���ItU w��X�Ϗ��r�/y7l ZcRণ'�8z�=2��ߠ V�>�Il�A =��&��:�C��-xB|�Pg�ġak��ALM./d#F0���\#G��$o�8�h\FDg����0d�	;N��	DH�������A(�S��(�	��r���V[lu��LF�vaSC7/>�#K�����qS���]?�� �����C�\����%�9y����ذ�ψ��!l�sj ���<DK� pz�qd$��$�MAi�,=�!�ԁ����lL�cp!8Z3��Rp^Bτ�5��a"�.2��� �J�f�IT���)��4q.��, �%���xQ�%�b��.�<Xq@0�x�G1"�܇^HZ��Zp� ���C��(-ÏXyC/4��Q:�#1cTύ��C@��Z�w��x��1Kh�@�m�=�|Z�x��:Fe?O���Y��(�J1 B���&�N�`��?�V���� ��${�X b�+	��z��������'�H�d�+DX��<C	Q�1��n���DCb_ޘ� "���N�Z��\� �K�0	�\���+:-��(z��<ȕ�TϰR� $\����!��o}��A�
|s:��(�ɨ "(�(Y�٧���#�Ne��?���K!ԓ3?;#� ��װ?w�ƻā�����S�٠ �>n����(�$�<����n���r)�\��ȩy�	?1��>@Ԝ�
E��\gy��H�M<@����9!@��X8�XJ� с��ڿ�x^F"v��V�|�%M����i�z��M{>k�#�&|D���||��f���ś%\�f���l.�-g� � ����OIs�Pa�
H3�ψ�������0����1���Ƃ'@W5�D�����/��gx�$g���W�s���=�|�DLA?�$���y���<����.Ƙ�I�L�1� �X����E�p�ԁB��g�d6�p����!�qX���W@�-��HͩJ#��!0��	�J���t����1�P�{�<�)_S�Ȱlӑ�(��E��Y[%�rs�� \F�ZS��CG+���T� �_z��H��=d�� ���Pʊ�l	�by�p�@86"�����
�YU(싙�&����Lh0�(��{xD�H�5`;�X �FA��PV��-�-$����␲10~/�?���AJ>��VP���
m��&)A'<x��!��|�Zj d�F� �(��	+}� ud�|�����&^Q���X�E��L�j�Ѐ�Z)�7�`����4 br��1��H���@xOU�őI���L����H���
	��)D3>�p�m�³��(�IԠmn�h�ę<` Ɛ�,2����I;g��~T	���,��\F<%�ȩ �K���%�9�t��G�D4`R|�ib�^9��*��p�!0pq �*R=��� �d�.���)��|���� _y��L1��ġa���*��r�ɢqy��8��Y-v� G��!��?�����H��� �{q*&��'Y�X��8�x���?HLqiŸn�,c�a��A^R�	���[�pr�� �t��>���GA
�����X"F��91���$�|�{7�/�L����z��p���V�4�:�#� �P������LMRK�h�Q���x��E>�#"?�������W D0�O� ���h��H�Λ��+��j+�##�H1��ؑ����_�`�]֓��x�\�����>Y��f���F��E�z�gm	s��rR� �%��w�|��פ�Z��"�9��e�T �<�m�d�`+��[�1�(?dt�L������.�W���|�S̨(�Wr�~djp��� f�pe�Ӎ�8���Hb �k�	��X�#� ���� � �H��ߴ�Za/�#�
�y���?�AHr\ ��u�D �|��9�J �!���W���I-�y��)=�`!',0Lz����w���s���U��7�4�'0͜r+��W�sn���O�h�� ��x�,
����ۃ?5|�0���'��?�Ię[|X����+H�P^FH =�DY0/� l��!Bt�J��X��U�q-&�����p��:��u�����Jj��"Yw	 a��)��� ��	�J�n�I�w`��.'�����7������xH ����8ͬ�g`l[��Jskx }]�d��&$Q�>����\�i�$O/#D�q�wEs�l@'�e�w%�i4yK YN8w�<=�0a�H2 #�c����dJ��<���qG�blO�̑��'%����� �9V�5(g�oؿ�fJx�0K�8�:�� A��y���	ɕ��<%0O@�� �����'|X�0DC���1D�@x*�R� z��h	�X&�<���G��� ��1�vS����y_���h��W��Dϟ���R��؎�����F ���	�m�l�ϓ�xZd�� ͆Ԛ+�:1&�y�z��mG��$`�bՙ�ШL�p�$q�) ����"�HOx���}��|=�@�$~?��x�A�k��xp��>#l,��V�b�����?e��)*��A&1�ݠq<l�2Y�'Hs�k��J�4;:l#�:HQ���� �$>(���Z9,�CF�ʠ�#��,�c��n	�X�@��_��p�����85�������>���Ų�`	�1�<�S��$� �b5W�$�8���?����� ��M��Ks@`a���m �}u
�P��	�?2`�����'=*Hl����
 Ķ�1]�� �I���c���`��1O�n��i���/����5lD�����_*��*�؀��0h�-�3��*��p���K�����Q]w��@0�篃��҈� ���aP�����8���uh�����Vy�'t��e��`G�'	���y�� `ZU(�?���ĕLl�c4s��H�E���fȘ5�"K�;��Լ� P@z��X��ߺ�b?��@J�t�����O�b�| �ˌmش{� �k��M0�����������~FG :b���$
�|/�4%e��.`Y=?/�+" ��~ �>�R���Г`X�P��gX/D� [�j	3��\ ��k��%�f��B��|�^FH���>�l�%���C���!7��6B0��` �Ӻ<%�`��� �Z�"����>?yӰ�J0� \�'��`�4
�D 6�T�$��Ƴ M���n)�� �Ԙ6�d<�C�Q��! �H`k)A.�Ͽ[g�d�`>� V�Kۑ�-�I�\���q�yE� �P�AZ)u%4o`?�z�a2�|�'��\F� 2w)�L���i��!6� �ۓu�tf���� �Xl��xK��>nd~�z��ᄝ��G��	b�w��c�� �NHI%����&w��W�E�Q��jI	^�Ƹ�\&<��ra���	�Y@�H�Δ��Г��Z��@��1�"K�?̀X,i�("���~vF3s )C�޻��	�h������1	�j�o)�V<pc��ry���|(��gN�� ��[��B�]=$Rk����?HT��b�R(���H5�'[۴�.��ט�"=T��(Q�8�����4|F5 �b��
�n �]%K �d���U1'ks�XžJ\yLI�[�q���p2`BX�ǙW.�v�d|��� �EQn��;6R|��+�0]��s��Lx�u.�## Nf�zt�$����D� ܞ4��[~ (�]#E0���Xq��%�SZ.g��9�Gu����u��j ��;�['� J����1A%LqX,��π�[3�������J�fc 61�:0�OsB����`��n��L� �ȳ-F�n�T��)@@ߛq/a� �p?�4�ݷ�|��|Z�	���\�/�xEG'	*q�&xtF� �[j{����Eb���k�W��T����L,�\�1�	�"*�T�jtF�BR����ŝ�\%�Y����e!��l����1��x��Nq!?P��p�uӖ%4 ���Oazr���c�,�*��<�o�r�����:#7 ��F-��h2�D����.��|}� ���Q-�p�H}�\H�6� ʃ���M`�?5"��oj� KT��Q܅P3�;��M_al9 c	�6| i�$����0���I~�h	V(�T������a�C4����d��>\����-�=��3�)���q��.�3��7 Ĵ���H��g�%���{�	<ͱ��H�%� u1���H9  ��)A+dq\� a`gEM�� x�!�j�6��"4�P#�Iv,��8 -�*�1fj���0� j�H����ڛ����t�H�dpW0�r��`�Z�t����:h#6 �N�����t*�w�$D�I�Q�.� �50a�O��Ip�l�tF2 #�k]27	��?��.�d8�7  �ۑ+��M��\�'e��D`�'т�����a i���g��LBV�X�l�k⍕k�ٻ*Ń��Z���>�.@4)I&o�>x�G}	(X�#�@kL>K�7��m��[�p��y�	|t��p��Q+'�{��?�zpؼ֙V ��{s�*� ?�)��G}�B����j%�ۺ�?�ӈ�><#���X}`O��Õ��a��".����>Slt>(E_�X� �_iD�n��2��g8*�P��D�����N@�������h<k1`����*�����l�)*g4%�/�� ��u�!� ��%�������0����j�~Z���4 �)�K�h/�]�PX�T����EBp���=1ϧ8̍-># ����-�-[�7s� ��+����0����D��	��8p
)Y�(S�x�� ��Rۨߍ�Ny�iz�1 *@0>���~���'+`[� �a��@K =�u��s� fqǑVT��K�����x��m��	��"s@ '9.��`M?�]ё�qF D��KO%4��_�`�F��p�M�4˨t���`��N۬�z���a�XT/��J �-�3�dа2 �f{Kw��)�A&(*�Np��7 ˅ mA* Yn�Z����㺕���3�ęi5 !H.���>-�^�L�5� ����Kv��k�)Xw�l�����h]Y�G��ޜ��m�����BX9�`�1g��H�$Z�t��9� we���E�%��V�I\����yI��!#�{�q;�� �	�8r�N��\v����@���b�u7i�s-�_n� �ʄ�?�+�gdH`��=���� ��A��6)s�����s$�I� �H5'���@�՝��v 0
H��1	�&�{��xN�B1���Q ,>1q��������0�|� ��CW�: �r��) ����0�9�Z�<�/A���������ـ�p�?j���S	h��E)R'����5�
 ��j��H+ [0I��9��c��d��@�ƥ�_�� ���!�rw@ ,�HݳŃ2�i ���^"0V�/�:h'	MB�՚>�� L��Z�k 0���/J����>^ ����� <�7��ֿ	/b"̀��(� ��ڞ��2] ��㆏�,�>�0%��`	�� ���_b ��;?�l\� >0V��2a���(� T��HQ( �8G�0	�/L�8!�t�ǟ�6p���c�1�z�/ 1t� �.2�*0�� �����P�:�8U M(��}�?�и�8U�P������� KzQؠU�e.\��@8ݝ 8��-P �Gy�I.�aH^��ˁ� �� X��: N��n��r*,e xɄY����p����� �7yp=c�0�� �����p6=q2�|�)�TG	�� 3����0����R�L&. �ΰҽi0aB%��X�м5�m -����B��!�^�X�{�����b ;sx�&���Ù̖�Jm�3Ӏ+�p�8�� n���U��<e�ؔ32H��Ȟ�� S�ZA�"��r8�?2åN�@��@#|��3Q�����Ȥ�`@�G0H	a�g 4�h���'�P8#�8f� ��!H�o�d I#�C0+@� )�z������A���=��9���P�
��� �qݐ>(.{� 9�s��3p�8�� }��i6�V(w���O ��kA�%�P��ɐ& 3UE�����8�F�̼@z��R�� 	*��q�`i��<
ј�Ҝ;3^�� T~�{	��U�����$�@���D��ҩ�Kp�
P��,.����8����v���'� ޲� J�r�<`��Ώ 4�;�p��ǁ�4s�8Y�`�@�U�N�3 {gZ�Ev����P�`�ہ��06�0ٖT;g%�·	��{B <����|'L��:s�P���c�3>{���bP�(�G�?o�R`��;*q �D��z�a���?���D��i� E�&��,�4���ٚ�9}*��!�`��4��<��$hrE���_� �Xa{� ]Es���z,�8w���y�λk�	�L�!�]�i;�5�Ч���������R�d��o_@�� �a��dr��IQe��H�q0. HxN��
h��8�W��"�%� �OX�� җ���Jr�������p-�D��"c�4�M:�V���	��t��9 �b5����&��-[�H�(���L�WH8��u�HN� g����i��ec w#<1uԧ�g���.y6����$�7�9 ���mT`�I�	�"��FP�Ai� P6�rYW�U8� `�NᝪX��~��n\���PnC[�ia"O0�ܘ�3b�P4��p� ���Gv�!в�@eL�;�PPݍ�o�����D�˄��1.&�R�f@��0����XR�Y�w�9p4g��f�߻^�8��&�L gc[8e���Z� �0�ξ���Gx}q�pn�ݻO%뀀�t��V0��UT�y�e��� V�P#��Cb���Ą�0�N ӎS3@��@������悬�"br�D���ƀ�0���r^�����	`���/s(�� g 3�EF�D>��2?k0������9�.�"n��(�2��\�Up?`Vz�e$[�� �uJ�8��Th���j�o���m�*$��te��	ŷ�0�&N*!�����G �'Z���>|Y Di��9�"� �K�.�\ex:Hڬ����� ��41��'�)�eX�*�$p=gۦ�� ���c`�3Oj�S��+ [Ð�\$�D�!CS�=ػ�q�&�y�I
,V�^�"�t1FV�>���_���Ca�p�d˘��;��.��f�Ѣ�Y�p׺B��$��#�PX�D�Db @P�� [֑�N����]Fu	"'tPSx�nЎ ��95��A�[X�!��4ǋ��, R�ߵF��#bZE�DQaY�ȉL� AQ�+)Y�j:^����!�)����� &�ہ�,�z�� 1��?�f����{z���uK]��CM� y�娋�[YP�
=�9�S�bs������'/����@� ̐f�]QPR��Obg,�/�էa�d���	_Y�`f�����B�i��a�����T���� 䭡#f|��� �� Zw���-���ax��W�a�%"%"�j '��K;Ae�fxi�FW_È�|�@GWâ����vH�w�)�-! ƅu�vSG��09������ӬGkL	��^��7W��C�f�h �[�H�. �����`�" �(q���H�f^U $��y��R�ZÑ�T#��BR�ض37HdQ��
f�n���`/��i0�:�# 6��P��k 5��}>��MV�� ��'fxH ���x�F �߹&ӡ��<Ѐ��W*L�B�S�	���]@v� 3�3��i,�JB��0,��N��6�������h\�5�}�4$A^Dna6b����f�+�Z��1������ "��_gÎ�Q�h������HQK[WI�'
��B��A+��m2��=�b��� �#��]W��)I�@V��o�/:#���h���W�	B"���`6�}H��.�# ��^�w��I~�w��-%{>)��h���&��PF�m@���7�q���`	7w8Fyn���A�Oʈ��;r�Ңl@�����9�p�ې��P����$���RWZ31Ӵ�8`�"�f������̈́A�Y���(7Bj��+���Ua]�ȉl�DEHU���Q�.Ϧ�tF h�oQ��*U$�V)�-(ڮnV�ۣP�ȸp�k��G��3� 7U��m �ub_��{��Ӛ�Z�ӳ\����E|�@��]�PX����g)OE��d�B�X`\�&���fP���ah�t̔�(������3Y3y�	��<�j�փL��x�  {�i�����&�h�d�*"!#�Bq+���HBB��L��H��~�@��� Οe�+��@S��E��6�#�X���H�������,i�{z��Q[Pf� �B�S���_)j��~tn;��Xv�/!���#��0�7��	��d&� %IYs��wO�	^Szz_'f�V�
6w[�L\F�7�6X���2��Qu6���@�(������O ��W�7[`1�f*�<�Y�a��u#P�� V����!;W9���?Q:�b_��&!���"�v0���ǅ�Q�� ��0&�B� �@%���7gc~ �����7����䗜����`R	f��| �F 3�&�%+DX*��ڈY�0_�G�M/�;
W��A��@�A�8����g�I����%�ǃ���!���@�rakF�xK���q#ZHg(D`�u$
A*, 
�!u\�+�pв2���K)��2/P)��"�G��Y����;4	�By��M��N�z�wH�*���@J8���@:h# ]�Ӵj���}���zy��X�5# ���a��$�P�X��.�����3�h	P��[�?T7� �0��2�B'����d�4)�OI�XyD�	��HD�aJP �X8�t�T+��6���h���C����=.S��{��x�� �	���p�� �,TY���V-Ş�|��[fF }���i�k��!���{����DD�WA��]a��ˁ�C'��1%��� �����#|�0s��Xe�I�ထ�p ��ٰ#��A�P��Q(�2�� ꪃ��63Q�T����[˗�0񹥠JX/�#=�:�u8�D��ug�� ��p���_ ���Z��X���	��g��dc���RД�J	[����T�@*�#� �1�Q+���C�y@���X$��8E�ߐ�v��-٥7a0��1=�j �*�X�Ʀ���%!am9�#�O���,�� �ru	�q�)ń����$, 'ė|�A�%w"���_����e	��$��q�`Ɔ�f�4��
�T,�F���:ۛp�� ���2��|ݠD�X�i"�Z��Mc ��1��*�YTYvF9���<W�># �=���ɒ�b��!�uL1��ب�5"j������NP���h< ܸ�WI¥�C�2kiS�h�0ũ�5h?Pe!�=(�Pj|hJn a���较���ok s&V�� �0[��l��&��+���:4����o�π��l�� &��^?��*	\k�������%��j)L�X��v� ����԰`%�F��Sa!� κ��1����tH�)0Q��_��T��'S�t:�# ��/`$5 ��Te�a�"�3F �+w������[h�zm �N��ʱ ��K>���Af���w��O �UQ��$y�����%��@�tq���|X �(��s"g`�1���-���,�E`H����0�y9'�g�e �ω��zC c%�I��D�9)7�����ҁ�}�F�� ��<:�B��ﯗ+���ƦТ�|�{k��O�`r���>E����B�$��g����"V�:�P�IZ-G�(���J��)�������B���h���\�-�� ��J;|
�B�e�:�ЅPH��`N�� �� �����Ǿ�[ܐ�c՟�K ��b"xg�yc��&�e�+�P^����Ҙ`��F���w9gJ��܃q�����2 DS�g�ڌ���������vG����W��-�bN��i\� (J��#�f�O 0��7�" l��\�	iϢ/��0b���h~�:�Y M=�g\���/�8�{�� �������z���p�G p�q�,V L���%�H �䥒`���P� �Y}�O��X�sҮ�8����s� l�ɷ�� �Z�_�ȑ�<[ ��7���;_������
�<V ���T�	r;�d� �0�!�6��I `|w�Զ����mJ �P��� h�3 ���z���<9� ���Q��^MS�Eǀ[�1� )A���t/ �D����|:�J.@"K��D!P�@��~� �+�㥦�ĸh��s>�o�QL��4 ��ķ�KP>s:
����@�|!0x�c ��ѐꯤ`$Q3Pt؂c�@"� Ġ��5�U&�8;�ˀ�*��D���� ՙa]
�CP 2�/J�K�&�� �a��<�
 ��2��g-����20����ks�P���G���~Vc��������Y��̔qS�T�O :�g�����#H�\ ɻ�>;+�� ���C��^3 ����K����tM �L��ћ�k� ���&�yO �L���� \Uv��8�ς� ��/������D���	y�� �w?� l��p�L�, �t�O�@8��u� {��s�Y�t&�G^���D���0V �
@��2�m�~E��`�L�$Q�\W��A��q ����E �k��l6�L� s\A9����m�� N�S��8j r��?�ܽ�l��p���),X�/'9��� f��	*By�o+��8���r�"������D}�	P��\��� �d)<O��� ��,�y�R�whj�c�tt:��XPԌ�G<LL�2AØh1R �F:i# ̇���:�Ԭ��+���u�fO���D���E ���k�7u���ҿs���$4�g {��~xu܋x�� �FP-��f�����)}Pތ_-�ţ@����L���,��x��B�]G?b�e����w>X��! x�-����?���Vr�XQ� ����CS
G�Ǵ p�Hl�����<A��@�ϽQ�}
�ð`�/ H��Ŀ�L��	�À�UD���2��9���ύ���E��'˧; J���C�U_��Q� h*k���$Ll4$�4i�ฉ��͘�Fz�̃L;��J���Z��O|� ;�%���C�>��F�����XQ�P.
� �C,��G��ɐ)J`�\ ����p���t|7�8]h�$lU0D3�J0�� ��Y�~h�I�P� �S���X� �1��̚P_�/O�hj]���X�侔��P� ����p�@�d Y%�^\����䄠*F� �A�9��,$�9�x���OC��H ���(FB���Y�$u�N�q�~`��F�x �e�`��v�"�8�k �dZKӜ�d(�a�z��D1Z�� ܐ�?�ܝ.�@��k��)9��A��p܎P��{�����`��N ;�.ڤ����@�P$��K� 2�l���.�9w���Dt����\�\�$%L �v��@.�X�m �H��(1Ȑ=��t �X�.rjC� P��F�8�������@�d)��U�x���� ��p� *ܢ��ɵ�����@"X�c^�<R`0x���B� p�%m -s{��&���� .׭X� ��?�ާ� �E��0�(x7�ܽgr� ]W·)M��ˋ��!k�u�S
�w � �K��^������� =��
�C�,|��Nje��p� 3DJ-ndY��	G�l���謰L�O���E�� ��h���:�<���VQ�)GC�P���P���P�1O�0 QV�y֑ ��U'����ok��
���NE �12�r�&���	�!:�̐ c%J�աY@��=����rǼ���xs|݃��H��.��'  �s�L)v%�]��!|@�t�O�*�f��g9��)7[i`O�O8x�
��bXfEk�!!�� ٖ����Ae
��><=� �<]�����?�P��@a\
����~F��8XIai�G��q��t�J��BsS��T
cU��#P7tŤ`� ��B��J��!�Ԥ�/q�=����	�h���V{���b�e�$�;�M ��C�4���.(# ��&��K Jz|��D�N=9�Aȟ�������98�CP�K�;�ؤ�B&�d�@��HC]9y�����$����M�m�FN" 5�Gp!�z�I�D��)��� �d��� _늎`�bU$���m�H�H�p�V�D0��d%��\�A��P�L�t�6�p 4�C \(�cB=s�t�U����n�O)!$��w_M �ԗ�y���\K���tzD�tF� 2��~[�$�v|�� ���hՀ}k��,gi4���0p�I)���q �����V�A�w���7�L�d�Mk8��r�3)L~\�{�»?h��A�S)1���B������1��_�H�k!h|Hav���b�b� %���m1����E 'w硳O3D��0���W@z�Ȕb� ��+��J�ȗ�^	Ě�\�o� ��
��˩�(Ӝ��#�(92)���z״p����	B���`@ìp<�3�s�>�;�oș}Y ������{*h�� ��^��P�l����䠡)�b9�e���7�� p"��m���`-7_�h����!p�e34CI���Y)���I$����� c��H\>�3���������y�3X����&��� O�z���f� IMq�^o �w3�K��#L�<��$��s���.ȸw����@fE� ����vä���ဃEn>3 ��͛/ Ǣ���:`٤�#B��ᤳ�����d�bt�,)n�tXu�H���'�:���^I�H��.�hV�)����I!�� (j�V=��J� ��-I�,��R?I�t��� K�O��+
��g@D�`?��$��`B�����%�0(|춌��w!f��M|��"}a֑'עt�w��>�#���Ǥ��bo@)���{yx���|��(�
B�(\F���h��
	��
x�Z$T2� �i�P�j
���K�����E����d�`��m,	7��ٴb��1��}-O���Hn�!�{�& 7c�h�\�\��}���C���@(��2`y0�5�bX�`*���i��/:�� |��6�MC�&G ,�h�15|��m�]F��;�[�`ٲ� �ԼÞ��|,`$�tF�-�|P�d�ȓ�D@Q��㏲� ����� �'k�h$��$
�oǧ�t�6���I�)�n  
1��Dk��P�AEM`�;�h�5! MV����ٿ��<����-��4l���¹,4 \�1v� �A�iO	� B��|�?×P����$�y���,��Dq�b0nt�C��m@c��`©)8�| �>L��ă�BM��h�� G��-б�J�|��Uoc�O@L���B�+8�?;�ءJ��i�PL �HMX	�<
7J,$���=��Ԁ%�\����_�R�)g�9%�o�W�9M�G�|@*��Q���+�pu���vF� ��+v��	��>�D�h���DR@-?�m���� �?]�=�W����fb�r��į���x�U��r���0��x�<x{T���xIJ�4��R;��� �~j�v��|t�y:�#� ��f}m1�Pp�b�G�D�`����^�e���q�HS\��z��b�P���j���L�豌���1�ĭX̑���9]`pg�HϠ!U̬O��Ĉ��y=�����KS.V�D��F�&�'$g�h�� }���V=G2�W��M��	�<��04���`$�%��d'/+�4�4�0�} ,���$ǯ�� L�]��s T}�+I�c��%[.��8.�a ���|d��$�'CB��� �A=n.���Ѱ��ׇì� �
����� +�5�?2ܴx@Zt����*z'ɑ<-�� U�,6��K��D� �=)!�z|9J�'�Ń���R�@�%kI���D|��P������8�Dû��5�Jei�(Ū�D������"`'� ��xsq��LHqM�E�i���}���t�|�)Y� ���Do�E��P��C�ß��5�1 ���I�� ��+g� q ���Y;�L e�~��<��`�Pc%��H�$7�@v��� K��p�c�������>s$!�KB/�#� �6��	��M]��@�@1wG lAW�0��;��I�7 ́�|���<^��ޜ���d�TC(G�D�`��: �W�ٜ!m����`�Eo��(L]Q�q�}�z�dC��@���z�R��Z�Hd �!��������z V��=�b���a�E��%DW.���`C��`�ژ�@�T�y�GE "�d=&��h�m�P-��XېcS�'?[�A�zĞ���7F�����[���á㨎 8Km�o�b-% �L������hm���NK���C�H��o{�J(��Ƞ�l��i�-?T8�	H���(۫���E�+�JXV���� 2�L@t�O��Ư�RX2Œ�}�D�  �(��X��b��(~@%��`Y�jqZ��#�(�RK�@|�_cT��!f��t�<q@���|U�$'��	h�H�|�� &l�I9�0�Jx�U0?p*�:8�L�y��>@�e�.� �qw��� 6�p���(�H�<"gօ'ώ��� �4�I�<Z�� *�/\m���|D�����}�0^F�r��w1g$`7,� K�hd`�/�D�C4{ &��bU�ͨ��DH� N5�}
g]��J�$���o}U��iI]̓ʱT,��Z�(D��s�XW�	}=�xp�tYZn,>T�zxqh��l��9��c�B�40פ�B�d�@�ߤm�LU�/X>Ȍ���BW�C
�^,^F��`���Tj�[! 4�Q�|{�` J�>�C�-1�BȐsΠ��;)�!-}+uVQ�%��[� ���Ҙ��t��Z-GMn�8hH�,� ��5V��L�lQ�\n�`h�tCDˈȹ������[��g��p��E;���(�҈g��8@��|Y��O�L�Q�PNH� �I:(O?�jw�M���5���BN�4�֤1 Nk+o���z�`��.�
 � ��}���D g�E�=�Y�� �%둢  �O��F2��s�-:4)!2�I� e�O@��ʞ���^F� !��#�w��*���q�YS�f'5l)�z�0@���D�y��W�rt1��=�[�"��D(����\T�8>� �Q�R�Ş���~`N-[% �J���$4va��bH� �'�<�+�����9��ǘl�`D�`~��K�P���y�!`|Mp��[i�+�j�Rp��,��i��	�A+�?�@1�/�>�G��jo�~�*�gyv�&tF� �:;K�.NG	4hk�����MH �Y]coK)ʄ�����'/��w�[l;h#� ���ŤЗ������*�(�i�PG ����/ �^�OU`��X�ѳz��=�!J �b�8D��xu� :jX&	�s����)������� ,�ֈ r׬��;N�'w�T�$�i�ĥ`���z�&=n:bD l�|�8���hVFw���s��;��ɴ�"c��YM�%�zT�����|���;ۄ'�� �z���@�p�y�?����*�K�(�|�8!ͫ��b� q
����U��O4����KR@�v�&�{4	1f=�����~�­  '�U�Dz ��S�(�y\	mR�׈�@^F�1��kĽ��Ґ��� x���:�@�e6uX�����İ ��&��0I�'G%����bO~ ^�� 7��1�M�Wl�xç���[� 	d���.�UC`)�:nX4\*1�G2$h��:�P �H�A�U��N�<���sh�.0ϧ �o��_Ji'P�-�8 ]�8<�	!��( 6�g&�ed|F� `��~�T�@�J�hAFv)�%c��Ot|ie�d`P���@����M��<��3�n-G���,�2B�V�@�a� t�8�C�+ ��[�|Y��g O
C}=��9�� ��,{����ké�(�民����8���0>��s�¨� �%�������1�j|�g��<P>��W�g�d�`�L�}ԕ�X��ml�;��9	��hp��Xa�����$F��СG�/ �̕�p�-�O�|��}fȯ�+ l,�I:'/��7� D�Ă�( d���)�*�b��x~�vF� �,-��ʡ ��H�O��~��!+%)q�5�}���{�;/�#}�\�o�z"bP�'���{��q�b�e�P��q�N*�@0LJ�@-l���>��[;D# *�q���G(����PȀY�b�$�o� þ���&[���m��9�GN�@���\�̬k�t��$P0X������8`�ӤXX�.d�:���s6�Lc�㝋���X��V��vKg) �puS+!��97 k�"����H\9x� ��0g��O� c�t��Ӝ�Хb���(g2� #P�w���Ԟ����E�cIt�8}j ��f@ Q��7~ae��V��L�|b0��kq)CY������/����r��І��� �I��f:��c=x0s ��$�' J��O�/��d����G�8|'%s���z��ZB��;�����k���f�)Q�l���H��g[{VA�`��_���X����F������� ��L]/�#�iׂ%|@��=
;���3�htM՟� �g��΀�;�F� <��S%��d��T ~���A����T� b	�\�
I��*��Kގ�Ō�0P�h ��n��~���`�f��r�}%\�%S@�Rh-��(�X��]=��T��x����!uM,�����w��Am�|�=3�}��g�%2�  �~d"��u}�=�s�T`vFLC2?V��<�����@"ń�j
��r@Ѭ�Nŉ8�{��gM]�lO�x�&� ����UNy�Իa�E�/B����\�ie��a�F̍+��etda�H�3M�;���"f,p(H�%k��IO���P0�8�DЙ�q�/P|,�F�V�ٟ�?���bY� ��=W�7��Io�>n� !uA�I5_gЄ%6 ��T���� 4> �����ES�ȏ%�'G�`b�^ �F��������l[5v�����\༷� M$z���7Tw}�8����:D� p�H�l� �5A�Fk&�e�9��(g�\�Z�d.``�Y 4ԅ�M���š}���D�CJ×'p�0��1�jw%Vd�བྷ�����Ԇ�Z���>�� ����=�ŉP��_o ��G�53=�˖=ㄤ�0�D�&�0��%Kި;�J����C	�pA��� �>���� Ď���:)V%��7'�=��%��L� �D�ܖp�\��g�z酕>+#�{�<YAp��tT|���P)�sߑ�Hɺ�!��K�<o�A�!���:�4��R�
i〇���Ѝ��+t�Y� ��7�)�o�3�Z�1��䊨�� �4u2�7)� ��]�Ú�귄�@��Hg r0�JV@��!����;�'Z�n39� w#V+�1����,��x ���&��D=	��{��8�p� ��#m�J�G�!�N�� S�I�:���-����Ĺ`��RХ\	��a�4#0 �1�R�'/s�@lH�D�gk�K���\U��)��,$A�N� ��Rkٸ�ԛp�����F����b�AL}=?&�
o>0#,�\_e�am�u%-�`y���Z�#�>�#.����Q�V��%�8�"g���A�lK��"4Oh@L�8m �a��'һ���h�Dt+0�QpO5�X�ҭ̸S ���	�<J<a���P�є(�\�1 �?�����L�h:y}O���q"�)�HK���ȷ�@G�?�cV�[n� =̬��B��҄ �*���Q@��}��Zy۬�~��� ��)!�w=ó�@���`������K.>x� s'�M�p[hи��- *��?1��f	���k<��R4��<��_�� +o͒�uGy��sƤ�(@��� ���Ǘ�I��M�2���*���B�	�F=�'hI�uԌ� 2������';�wV��x$�l�0j 	�x�bV�O� |��Q8�(���5m�V���i� �eѬ��4���o��ȓ#�l �Ɉ9�����)�D�H���̧�w��:�y�<r�^�BB����{����淟���wT������H�< ^L&X&Ȱ ��s��oI ��er: �X�B�o)/7��\�b�DT��؄Dȏ��#�&ptF�[�7���$������,�X�9V^F.t���P
_ )�R��g9��W7D})�"�o�x8D3�	st� ��7Mk0 �,(�,{z<���Ĳ�0������h��P]�\�����H��t�<�>�c�).��})�$XY���a�ڕ�=�>�N�������nۘ���z� b��G%�I��<q:�{$H����C.n��E�	�K ��vF��gL�w�%5l}@x)GN���.ۀ�s��}=cC)�����?'��~U����ȳ�b����r�e����]*옓�x!�=>��XHz��R^8J�
�	��0� ���P�Iו4VG|P`�Zq�F��@��9 6P)�_%���L/q`�� P��"ʀ%h�Kp�u���s@��Ԍ��+\Dbü)Z�L�D�����\h�;e}bN�h�%
��H�FG�h2�����0df�C@�����$�� ��gUu��	�zP���㬇Y\�	cUCV�%Q8�.�
�@l�%��H�}� sE	��?�rT}�/�������u��?�`h�@h%X�H��$��O��H�-�54ׂ��� {��4]: �<�me['�K�L�FLi���؀����z ���n�� (�Ł��j� T7��s���"�t�t @�/�1��I�R�w��|���_�� Ǐu�%X<�%k";��[�ސB!fI(�|$�(�� g�� ��Nm=_��P�P�ݻ�G����"a,T)t� L�
���@Y*BP,�#��:�?�STc� �/tP��vm�1��,I�Cp⠥�V�:�J�(P��*�\���sa��B��4$}-;������ � ks�ΉGE�I{� ��J��SC}����-��D�&���˹L�^6�Ԅ� ��n�a�&�D�9�%Ch���J��,E���Xl�� �.ؚ{��DWJ�ʔ�W�\2�$+�:y�%d����ތ� V�\�bC�N/��k���S��������@-��<����M�F冤���o� �3˒�:&ڧ��D��*��t� ��)%��H<|y	��mt�)�BJ����k` ���
���)F�$q�� �F@�,�Z=��ܐPg0��D�	G��y:C�}=#�0s>5��H�\����æ�q�F\HP�Ŵ vF� �_��d	��)��DyܤP�%Lq`,�$���ܘ`k��`p�3 *�h̩!|��!Ą�� ���b�����l����Ĥ����p���y��X�� �/�2���5`�i����1�Q���,�Uy�`rI���������~z� 0-y 1��>�n �t㬦��y�m`ρ��0�q&~*� j�.��F R}�K��)/۴�U���*����hX����� 1��Jo`�|�+�+��'��لhr�)hDì�H����<��^W8����}�a��Ji��#�|U�*qHٵ�	B����J�L-�Z�;�љ��&}.�8����Eĸx�ll��A�$���� Z�r#�vox����(�� � яSR�������8�Z�Tlǹ`� <��J(�	�A\���'t��9�NK�Ub|�ؔK>��.nP �p,z���y"~���܀t�|�+�	@�&��$��ĉK���L5v('w����GNՀ�� (�X�4R�M�Oט��-x����y�:@��舤��	v,S� ���C����d]� Z���x+�}�
q�d�QU�a���بs%�P� �Xr!�=�%0)�'�������Ds�B��,tF�	�GX\�:�T�VF-���y_��;E-!k���Ί/T��@�|�H�`��W�T�^F��^��L�	?w_tP줼���K��uc�h�%6�d��xx�%�|l��$D�`i�:�����W���~���Ԡ%Xt���`�j	=X}%&ܰ��O�+.�<*n��ݲ� ���7j)���~�l�'�q?C'ʒ���;<!#�V�_��/�*�\�K!���=�CVfx(�I`7"}i��)�,H ���<WI�be��*���`@�W���sL�����,7-�	�PpO�������ҹg��'%�
ZD^���D1 �nM&*!e��Q'�鬥 ��9��j{I|��*��Q<$�rŔĽ`��: �U���~ɕd࿄�D@㬣6� (��X� ʖ����01G$"��, �Q��F�5�D0�hc���hHç閰긔��0�"�JY�A��*ɤj�s	/�=��0�>k�_���@XU׺еmx����pZ��TU�,'�����z/��H:g���
@����9I� S"M,e������ j�
���EcU�I|�s��r	SC�0gu���>�p�\.�w��M�����`D���$,����P��y��t �%#+��K�9�����QȏH�Ҹȼ�jvc-K�0B's�x8K\���$�`�	���8� _{��w (-�̰'�_m�O����-��X��)��=�Ƈ�43��� ������8:,*��� ���&L�0 şǈ�S�� ��4+�'���)��r�J�9�Y���x�� q]�7R�����>����^�0S�i)QO���+�u������ �ik�*���|=?-�\ptF��>�H���?�����b���0�� �,	����=?'���@���q��\��("/���B��$F)g�%v=Y�����SdR�<��b�-[0 ����-�O�@y�*����0�<�j����Xޙ���� �L�z��'�w)'d[�f��)PM�g@���e�	�w!h �ׇ��u��	ZxPJw �=�O�\�bH�U��"@� D�F}a(���h� �A� M*H��2�` Ӊj��=�y��씪��\�@rZ��?�Eƪ�@��9�|�W��Zt����@��f<�\}�-���l�@J�>S�D�d��%��c}�e5 (�ϡ7ְ*u)��(���E���I�d�`����v��� |Xg�p�A��.������g^Ҝ���(��%}��!p�|��� y$��Z���;��U���vF���� H���;��NWĈ� ��S;x��N��AQ�K��P��� �THy�@�	G�*�D ݒ�	��?�B��S�p��=� ��	b�����'�� �$�	ig�� �r�������������4�.��z<c��P�Qa�$��ͷ�A�P#�5h�@	.���F��0�����g y��<^F��0�r��z�<�%����(�D�K~@�'���o
_��L�y"x�Ht`�y.e�V G͒����US6Z҈��)�-�&Y�ǘH-�|p
��t�� _� �1���*0�x9Q�O��Ii7��>G�������v���q$*�����$蜘C����6�>݄8�kH���I ��6�~�71��e�����Jms-Ք�D�"Rd� \�bJ���L}�_�ԱI��P*"��Qc�Ǡ���OH"�r�x �ZӴ�:��=j�P�����q`$����f]À�$�6��i�� ��h`�� ������� t�:�<N�(��/��9���^Fy!z��:pp\�A]`hZ�ȸ΀�>��}&���<�vY��vр�[�\nV|�O��.��c�a��2�P�z�A ���8_�Z@�L9T���Ir�֨�%�������q���{�H�@��D}�fXcJ�p���\� ����<� 9D\��BV�y�1�,��~��E�*̴MK|� B%sg� %���X"�b%�g�$�(����b-(/0�z�'�8��~n�z;!��i��kc=�C�pp@Q�^_)ȝ(�����1B
@��f��?'���"��	���Ps�!�q�m>vD +8���� �Nh J�b"���[%z����?v��UwHq�i\D�8Y4U�����{zLi���ի2��l���'�%��Ƭ}=��P*����6@Q��L����5\��L����w�@TLQu�ȼ�� Mf�)׺��&�D�8���T>D�x&�LF ��Y��%� ����9.а�P:�t&��FA��d. ���()!ٮI:���i��`��3ko^�����U�D �t?֐ �� w�����$�mT@�\� �-G�Iȭ>����o(ќ�m�U�tL�H��<��ҿJ�b�*�1��P�襌&�V��xp�)��tmPx�s`�� %勤[�|���q��E�t�osLp(�?P��;څ��>4#�4�0]��u�	1����h��C+������J�AiWX��`��b]$�% ����=�lZ��'����k�z =�f�8{�$'7�-=� �?״X�ս��Ԙ'����R%T��Xv	Ce��\��	�){����J*�4�� '/��܅:��n��{n~�@%Tg �G���3~�%������0I�Z�U�����f��v!:�@�l�Y��ks�S�� �;R��'���9Q����(��� �8�>OϒO���yJa��&�園&���, ��bd�L�GJ����D6I�K���y�|{8./X#-��p`4���t�I'G[�{X���(!c�j$X7�y�c%�~<�?��{\�Q���&^�д��� _'�~�F.7��RO���Llp�0é���I���s�ojn0 C�t��U{NI�X[���(^:
x���b�A� �g�AfA�� ,�@i�P �N��	*�  �D6FV���B����K����QpEe�z\�{(	e��D\�k}U3P�!T��t(�iY ϹQ���G�A�(ٴ�,z �E�"l������X�n�(f��m)�����y�y�3�o������  �<���SrJ��0/��KP��"��K���(z9�<i�@ċ���68�+�#m�L8(�K��l�h�&c�@��#)'G���$��hx "䀄u�=(B3��9��Ǣ�\t�-Ip��L�	Mn~���J��-Z� ����i�S,z�� ��P��; ��eg�:u!�t��h�\F� �W�X�s{K
��M6�`��	����hP���h`�@bc@�%�	U�X`��_�U��� 1�vM,0�4/�
�a��y�,	_�\ �PD����/��O��b�s��%����d�S ��k��J�D|.��p ��_P��y� N�>�6,�ɗ/�2��
U>�G������4�T$�*���;�Fi��J�2�Y��R�:u�����4 `o@��达b�n��u��� ݢ�d`���^fC���Nn�ˍm� ݝ����8xUGէ��nz� ���-֒A(N+�tk�`�!`�"$��&��'���5�����X�Tx@޷	o�n�¹���:��� ��E;q�vs%\��h� dɊ��(�݈!|��B���\c%U�t�Q���X�\���ɺB�Z�ki,�+��c-�>��@�~A�A� ���E �����oa�0�(�-U����Y����uKc��Bs�P$}�t8��D�{"|y%óyL��gm�W�@��yt8'��Y1g��b�*�����Q'�Ī�0���ic=/P L���<��� M^���.;�T0��U7cy2g�J�$Ʈ0	���*^DP�O��`�}=e1��,�)/��w��,�v��&�A�t�P��%�Bv���\#�̏��T��+�` LG_-lÉ^ ��?Q�8V��>��N��t0�@_�^� �Jeo��u+%q����0uG�$�� ���rT�9'Pm��{ ��Q��?u%��IˇJ�+� ������~R%)�!}���Ǥ���Lb���X����|^�J�	c�{��Ddt� ���{v Ӵ������<�}�̐D���t�q� Y��c,O�"��Pr��͵�<�m������Ѱmq^�a�:<�RĦ��r|*�T�a���P�T����~��YXNzY}���q�d�r�}Y8Y� �{�J�(PB"t� ��pEw�3R �c����='W'ȸ5@a��L%�\�kM,@5���;Ȟ�[`\�%D:�(W ,�%H��1l��2���[$p�u%�Y���G�X ._��2��j�m�?�p/0�	7��� �:��8&�y'Ϟ��ɻ���6� �xW�+���C��_Dh}���ϰ�J!p9�9�h�d^ ;�"!��� n��� �oq=@H��|�DKr�4}y�~l���H��� �'*�U�>_�Рp�Ţ���  -)�#r��]Om��:�$B�H�m���<݁����ܫ0�V �C'H)]�F��-�|q�Ĭ;�Rp�PN�,�[��ţC���눈�|��`��eG+�p4(��|'J\{�X�u	gC��X����� ��<p?� ��	c=;�����&����� ��}�O�� q�d�	�{����0���H�] ���Nhy_I�l�:f� ��NV5�F 3=CK��L�\7�N���ݽbW��TD�	�r��&�J9� !������ RKD�Bh��x;����l�?F����3iw���̀՝�"d����Fl�a	Y�K^\X"y��ԃů�)�`_ �4��ɀ2�D�C�}����p�kC�*�x�@]�	H�W�r݀x�Q�k��,�?�dc�����E.����݌H8��}XƔ� ��jg�`�t���� �;���Z|$�I�]+�p!��'^8�=>R���DX���?Q�^�؀A8���'O���� 1�s�K�7N��HJ�l�
�\o��{)?s�(��k�4�h�8~�d$����6.]M���"���4㵄-��l@{���)	�n���w�\)cVP;z��S�ļt�ȯ��%pX�D�l����s~Z����%.�� AHhlJ���耀7#Ĵ��2���IW�L���l'%s`^ C�g�M���m�j�/u�hBs�+a`��3�UI����@"�:��8|�f	(�}�z�E�*Ĵ�{H�D���Ւ�7���R��	/%��y@�W����+��̏&����x�� %k�Nx����oY
Lru}�m�w�T�8�AS����@��0�z�	ۘY-v ��o�ME�,JQ�HX��)*D�$��q���h���$+�� ��il�FW恞j�،��%Iky�/�HpJ#p��|=���g�>�80��� 
ڮ컝}=}�|%\h� �����
R�()gX�I[@'��_��|՝�����ǯ��.��s[D���p�逡�ri\�K���O�?hd Z
,��>��SIv�7:N���`ѕ�'������:Dz��X ���~�Ҝ�Ѿ �E����Aa+���ॕ �a�W��'3G\��^�� �_�"c��9��)���= ��H�?��}%�)� .�8��J9�͗�$\l�趌-kM�4 z�Bn�'o-���O�����7/L�%�B\wMD��V�)!�󼬓�8W�0���g�0!y�q ��tq)7翄l��Pü�|F �����=��%d� T�9�����[���FJ�v�,���{��`H� ��r����p�|*��Ȓm�rJZy�x 2Ǔu�. �
��5h��p�y߸���w�5�x�իZ"dH��'q�\�tF��}MI@hX�%�1��Ȳ�?�S��ǗeB��U"U�䉇�� �7���I^�wY�h`p�5]�	dzivd����[�� �<�M���H34�e��3ډ>�`*��Ӫ�|��#K�tJ��W�HO�ZԻ*�`|�>H�9"`���N*����j(�J�gE����A�0@�%WR��Egz���hေ{����;jZm��� y��r� ~�on_�?��c- �M��(O�<'��\l�� z~�y>D] 0�%��Si�a�9��'�<O��	j_�t�@�ֱ&�.2�Pa�lk�@!���h�\��c%A�� �9	�)/�x�'��@<}�=_���YL3�>m�H�+±w""f��<ë��k�� Զ�L�ᛕ:�	�D%����	�.h�Y��s9D�k��,j���:)�>��d%5K`���
|~C�T	cU�8�� (��FK?�	|�i�5�z���B��i�Ͱ`WKV
?�t8��P�g�q�+���� ��Ў�	�%��I���ؓ�$Q�,%g�D�`�MK�S ���s��sn �����B[Qȏ9iU�ȖVF. �P�F��K\�]8��I�����5˨�x	�B�'}�P��R.�k�\���I��-y\IT�� �GS^�@���,��(^,k�����ҏ�k@V6���b��.��n0 C������d�hKC���0�(7�τ��D��(x+�9)k�zͫ��.�L�����Y �p�Kf(��e��z{��.�)Jսx�l@3R��M �%A�j D�#� a'@dg�Z����ջL�q[�?�0����'k^pL/�[���DHؿ|	z(��w74 �ۨf�'�l^@/m��P�C�B��p��BV9��G���-�	�=YU�4(��R��j	�V�B	+j� �,>�5Y�H�x�`3��S�i�.H`�X�PL�� u��z��"�������/߀�L7H4rM��� %��D6[!�\$�a3�J �1)��<�M^�� �����{���ct�8TRO���U������M&o���ڐ��{������&����p��`P��(M��a��K��耭�y#�}d�����M"ⷳ���Ÿ��i��+؈�������ZN�����m"�F��5~�@�޿&�=�`��5e܄�ՠoWf�/K_~0�?��[Hyf�����%7�-�]v��~q	�դ� N���O$fP���~]ĕ��c`��@sR� �{���&^^�K���CvOZ]�%a��
,W<���/)����������aI��!�e�d`��;H��x�p�h(`QA�s��M=ɀ+!3(.<��� 2��{�� �X��	^�18�b5,�(�A�.SV�0�^?Y*������ !�S�p��wt�	�������Q_;���� �5^y���:0�#�|�o@N)H�d�G`fc�,�/�h�r-}�SP0L9D����0<L� X��u��6�6�Cd��cP4)(!X�W�����G���
�R�� ?�����^�� ��b���R����,_��5��cj;�m���"�8������$��03��(��&�TvF ��6>��X��"�,�~9Rd�0m��L")t®��)y����P�f&U	���g�M�Q���F���Ɋq������ L������I��~��İ�����[j�����7�$�� c{�2�Sn= [�a]���"�����)�� b��S�؃/�~�� %�@����H��&�P )��Gbb�	��.��gW���V�X�UH=ȸi^��x�S�z葿���)�`��#�����I���O�`�H��I �j�*=�/����D������H���q��Wcn[r4$:q# 8-{@�\T�6�������G��� M��QL΄M$k� ���f��@��R`9Q,�&�=`�R)#�a��8^�tP��C!��(3���)�)�����z��()��$j�vF1�PYb��)�U$�������MS�5�B~�# �a)I���&�_��&�� 5��-�)���!�( ��@'��ū�jGt:�D9��_������_��̸� [m%��a�y7�Ϋ(�|D]����WA��P����f���n���?�������;.1�r��]��ӊ����Nu�פ!,���L�hږ�/̞ i�߱��+���s��C��ȩ���1��� �}���V:_PLiQ�%۲jQ?�� Sjz�ػ���i�L��\@����������h����6RI��gDg��4 �Dv���
V�*J��"NB4�E��{	��bf�jt���P��TE��٩�������g�]��I�&��	L>%*S�=~�P`|ka~QX�����}d�5/�"J�%0����,M�|F3pd��E(��P��Y��?���g6zi̿"�Y<]x�O0?.�	ٹHq�ᱭf&Z�
m��Z,w �3��H�1D2AA���d��Q�p=9�q�ȋi��A���!��_<A݃�_�ɶ��� �I�M�)C������\"�(`1�@,a���r����]�%f��Ƚ	�+�\`�Åw���{� �o��H:4��|[��nL��*�f�� ���4	1"@t�~��p� ��IN�0���|����H
��a��;�B��\15���sMLV�� ���E&���B��`�3�`� ��p�!�2�*aă��-�%�!�	�G�(�����_�;&#�7�QH`)���YC�7aKdnM
�3��S��' ��3�!��$���lX�" ���~����
��0I�?Hi*9�� K�@��P��	[�"˂�J����і�АN�+�M}�)�A���F@'�:�mu`k:uAX~f&�`?L^��/e͉�D�]�g�*,�Ƚ�P9������&���į��D���KAЭ�T}����%!YNmES�q�5� }��4��E��{�\kk	�N�S�zU���)��Mo�(	���5Z6,�}���`�f�!��%���p&6BM�>�,&IB���GA��	��y��Zq��6`���S-萟��J��I)��_=a��� �&3
���v?N� a��ѕ�3�}	�Ur� �-_?� �E��y�AT��u[K�4C�8��gA���mt���M#��K#��zq%�FAvHf�4i���# h�W�z�~������X}% M	�r[�4$;T�z��'�������*��+�A��u((���B}��<%��N%U�܀��d{9	�}q s?YV(���%a�<�_��ܵ�!� �- `�ᔛ@4��^xn(@9׀��ht���1yY[a\i`	���)����e���.$5�a�qJ�$N��/ ��$(RuP��Mϸ3�b�%�hE�y�ʀ�';�f 5<�$��\�� ���Tr�޳�J�k��	�b�M�����|Q,Jrݽ2��0.��\�)!a]�8VJ��Xvߟ�l�-ǃ�d�O�[���f�s�%�gb\
)�]���=��Q����@Z�
�垀�Z�p�ض�i_h�w�<��+S�\[� H��0_5sl�b�� �� I^P���a��%�٣�{�J�����0�y�J�@mC(��| �c�/YiINS�ne�_��U��X��W"R��W��5��Ԧ�ER��J�k ����T��J��6A�u7,r�ys|�Nۉ��p�ԻO���%[�=n-ʈ�`��҇%raF�����eB�T��fJP�j+���tϦ���ȩϬ� n@�V���sP�"�-׾�D��Pfs�I8�J�k"	\�H7��s�f�"J e�w%�E�/�]pS�|���`��3��40aLP�_e�-x�� ,ȽC/��z��{j"#'��Hs,�	�	S����?�,ׇ{X����)Q����D;�����N��V*��\�9ċߨ�3��"iA-9 1���-����U�1X�'ۖ�vUX���tI���I��(m ��KP�]/����kļ� CQ���H�J'g��?J[$=� P�;}묁�m��)�0j�&���ݣlX�%��C�]P�c
� 6pUS�X�xMꐹ��	���E���8�+}���ӌ5�Y�*׷��� �v���|�W��sXx�_4���y�t��	����� �y2��Wy 
���������j�7� �6���743p�<�QK�ҋԁiВ�; |hֈs��S�3]go. aIO�jf��I��5�,f��#��-��OJ��9��K����%�7�X�h��0P�Y7d9�	�* �U^��C�u�T�+4��߳��`Vf/���	Jw�n� ���@�+e5��+)5i鸕���|�S֢���BfW{)p�� �����L�&�"�D�P��k`+�M��E�(.�H&��? w���cW�K���T�F��c��뫸_�p'�ڐm~� w��gt�qs���2�7_��,0#�q��f�����@��%�jcO��ڰV<B�E�|T0%B*`�+ȰWJ��Q("`�W�" �U)�!��&nA��KrZ@lq,��16\	�X��~_3�+HT�MA�?,�Q�S3�p �K��'�}�s& �P�>F�["� ��1��3�e�?�:��0h���8����LI�&[OwH�"��@���%���#�  <3��m?
�[��7�sq��$`�g� VM�]�	��lw���a����"���w����-F�h=�r��8Ǜ������@G��;wɴ؛^G���� :��u���0S�ĠY���J݆+��Ar�����nz;k� �a���B%��`���t	�-[�.��$x-7`�6����㳀�=|�t���@��� �8��[+����5'V�z]��Z�xJ�$%�w�������x0��'��T�i��po� 
��)!5`\��Ɉf�%�ae���$"U����b�W)�aX�H[��[�Y%�=հ�������@p������`�}8 ��;{Ӥ��鲕�]=y�����+8���`����pz �`*nb�F\��V� �Ӻ�@����}%�{_�aKA�T���Y��m�����FM��8_�f���Q �[��8_��7� Ƴ+	>��4/J��ͺP����	ݕ h��,q��`KSg7 l��p�$�bW���2�d�#��f�_�t��̨�9�"��, {!��s��� �eSYIi��\I=t ��RQ�Z�W����*� �l|&�f�sK��,A�!�N�J�я��ǭ�p% �fƕ���,+�9-�҂�=
�6j�Fو��� W�b0I~Q/���sp<��[����4]Spy�������8�_'�H�b��U��t�I�iq�hK. !�G&���b�W0P�K�N3�}��|UJ[��XQ�A���%c���"��0�%Pw2��`Wš�v�.wBJ捝0��g4#)?j� �݈�=���Hک��� �F��f��<�ƞ@������ hw� 
�Ԋ�����=`a:�d�f	�,aYtGS	^�����t҇�V���)�>���y�Z���.:b�ByHN�b��{� �̤W�f�)���bV��a��pY&��B&d�F��BLJ���K��+�ف'��� �[��d(�]���ޗt/��M���P��Ad×%�0���[������W���.u��S�^$:�% �����[)�%IŚ�M�A_�1��jو�#�`� .��H�ې����
��p�A8kt9���%_�n ���,䎯�� +���D"q�O	v_p���x�d�Fȇf��K�Bu���d@n�󢎏�ѿ���`���E��IL��$%[SY�  �e���T_�5�����<��k	�� `�)2iT���/��������N!�ˉ.Z�qݬ�`͞x. ���i��I��D9����- Ս��x�|�,
��� ��%[��ц ��L=mǚ4�Y��{��f3��k"�;��@���E��^,���!��J�bAU:Eޓ@�)� 2h,��̭�!i{\�RU+�[qp��-��ռAj5+�ㆮIrs�M�Azd��!/�0��<��u=�[�:n#֠iyi�܄��0�-���J������]��w�� ��
n��#�pu��7����C�i
��g��S:�ZJ_H�s��}��.�j��9�H�����l�^�N�ó��u`�p�M$;̥a� ��@t��� ���H
�Ų�CГ��[�|M���/D�ڜ��е7
�Һ�@���Y��B��#�I�$t&�ѱ	��y"D�A`��Ylw���KI��j�-�2��� P�=�JO��&��[^���(۳����pD&WK�$��L��TS���ʃ���LJ�����%��-����$i�T��,�)(�l��@���� �]����aK�  ���p��Pl�zj��"�H��?��.A��
�/��� ]��I�FK;���e!ٰ6��p�@���qh1	����G��:%%d������%�0Q���= ���')�hX��I�����:�$��sS`<$��t4a[��*�����pP�_��䋍���E-�9�G��' �?/y>���E��_ �}jd��� �Հ�x&�9��? ���BW�/���!�	'�AǷ5�Ag�#W �{��:� q��!����۹�P9yR+�'�m7��~0LT���!@��r���� T��@��S7h�Wm�"+�ͷ��2�j	�+�R@%_�������w���)�� :�t�1p��*��dBmR�J�1����t1�J��:0����A!*+�R�q1��[�J��~"{�d� ��x�,��򕋄�`�h���l�Q��J�ݭ:jd	��� Y]�=�#����O� �)��������}V�8S�
�[+)�	��YsD�!�`T��LJnT �b���H6Պ�����p4Sz��o��<_+Hxk�͆����F­#���ޗL�&��R���N���ȕ���	����!���j�-���@�7{̄ �8���m)�.�j�_o��P����N�"��!ҧ di�&J�(2މ9`��]�����Z��}9a%Xm.������P��=�����NԼ���a�,u:���1�N��� -F�/Y`�Df�:���P��Yj����%ӯH����j`�h0n1��.3�< ���F�	zڀ�T��F<��b)���ן��5~RYv\]8��a�Cflˉ�rqbpw��g��(U9�@?��o&%9���QȈ���4$�%�-n� �h��vR��a�.Q�i��JU�{�1�0`�P/P�E 6_Egnn�2����� kRL�na��%�d�=z�v��?�V�T^Q
.�A�	�J��*n{  �
ԶZ- ��1|~5�y�4�p�_9r�鑉���VTQ*��`�դ�4 k?��qC���-@&q�͔H,���鋨� �ĂL���wN����5'�������gk"�;ȓ8 �Ens��_;�ޛ�P[� �cW�V�/�������}'Vj*`A�cR T�D(��4�O m3��J� [�X���ҰJ���{� �w��S�%��7�K��0�E10#�ׅ*���?���%�B��b��L����J�N���(yO#����QY�V3�M+�F��E�-$ڙk�M�B1����_n��� (�Xc�MPRQ��_L<�Bj`	���!��a?�-�� �Qa6$k�2ˆO�ԢFw{���-���a�����X`�� Q^aP�M/qA��f�x		����V��F `����G�w�@?4��� t�q��f��A��:�_[��� ���2�4�.�Dq�Rv�,��Tne��J�w{Băb��'c��_�L��+(8X���PY�:\�� ݝYo��j�b����{���(7��N���%�;�%��P3){��:LZb�U0[�*�/���G)�6���Q���n�+�����xu�Mċz l5����,BO`؎��P�/L.| h�^B�� ��I8X�[;r��'��xJ�c>ӹ���A��� a]��Yc��$��j��%����ɉN#e�u�W�{;)# ��OC�qf`
��%����`��{��;$�`*'ȯ��j������҉S��1P� s	���cq,������u�/�A�kj �`��^~W �8Q����iE�~q�[gd_ ��1H���O�-��cPy(�//��I�[+k�#�b|T�I{"xYd ��f\�[����C��b�]Z�ɷtY�G��6��+�A��=�+X�),liF^��; N�b[�"	��Y�i���6s,� [���J��Ӡ^�<��M �7��#��	���Ľ���Zj�����a��~0"���TB����} &�.n�z���IgJ�
�0N�~!|�I*1)3�z�I�M�)��$�j�/n�&d��qycyc� ���ݨ7د�@_3��J��"���'�M�q�p��rLE� �KX�P`�OJ� ���'�#��\[$��kV[`Hə��mI��3� ���^���a+Ȑ����*w������8���+"	��X�Xz�_I�D A�c=j����{8
6���N�	�_r�E(+�$'?�JL��Pt`������[}��9+0���?�C" �b!V��f�\���S��!%�́|�%$a���� �A���s�3�Ep���l���%����7�2�H�%�#ĥ)�]�.��|vY:����+���/O`�V��PA�ڗ4��1���"ߖ��m:D�����歏���THK{���4;�|���ϐ{pa�g*sJɞjn] ������T��*�~���k]q�]���Aq�; �ĸ��ac�Jʙl��K��U� �,̀��
xz[+�g9�����V2�"_[�ۈ�ItxE`��I	���Fs���|� /�����Z,LV�_�}%�Z�ih�؁��C��(JJ���0:H��P���_���.�d���ߺ/���@�Y�p���#�[���C�B_ΐo��z�<~��(0�'IK����h�u�R�e x*�LK�N4�2�`tԒJ_�svϷ��)�_y�g����j�-�j��(����3�nHA?O�3ӗV�%7X���ֿ��1�q'U���/D`�}zn����	��j��:�,� R$���8��H�ø�қe�]A��Id��qu r�3���5����q� x�����i[�-@^��]�L~�����PL�Xj�E�;$ӂlX��h�*�)�m�Y�]����C�g8+s������*'P�c����I�c�F#��av��k��@yMiYWHc-x�ɽ�ɴ3�ukB��^�^7wK{eP~�KV��%^`�r� k�T�e��o�[a_���	��(�d� J���:�����g�����K��L$=ެ���p3I��ER�ŀΎ�]���B�a��"�>�f�/���*sB	��^HR�5	0�q����/0��	.Kn��+ �Ym+���TM�hb��_P�*���pq]}���Tr���oe2*�uN�ɣ���� T4�-)���nP��@�IM ��;4C�"�)y`�`�����[ۆؑ�P��ް./�.�T �k���Gu��V��q����چKg�x�΀�h�?-%��戠(i+���/��sݷ��[袤�k?# ̴}���ܕK��6װ�� M6��P��j;�;�n.	ۨYA��f���</u�k�.*= &�g�=���KW`��%�gnc�,��@�& COA�l�(���KR ���$���[_�o�s�Ĝ�N�b�^��T�� W���T9�;�	�h�����cV�x�<��ˈ���E!���j$�}D{���%��:%�b�
�'\���$���4�"��*� ՞����%��m���e�����21��?��]^o�����J_�ʉ���pע< G*oS�PD�����j�݅�_�{�	�"/�l�*����4�	��&��;�f�O�5��"F��%��M��ի���\/�f �+��
�����mw�&uew2*���7g ��ڶF]ʨ�)�1[���FZ���_���� #��(bԮ� GJӅ&WY��9��+��hKvc*���Y ��b�	8j[�p;	����DV��U?�g�1�q}�6����`/���a�O���W�	/j� ��f�������;�Z	�_旲2`#9	�3�)_�,�C_kU0�[��c��7 �J���\��"jΩO�u�t��g�+��כϓ���j1�P�ak!��i��	 ����~�1�ٞ/	�J���p�%�0�BP5�9���q�.K���]��t*)xE�q\����
W0��8�����9`�L	p�a�f�H��J���+��ѳ��kY �&�-���\�V��`�/_��Vq#�����:�[�!�b���!Q	�%��`���
�9��T1*���1n��Ľ���.S���Ӛ؀��H�%��$��v�����	pK!�tG�=���1�	T��X1%+��H�� 5���D+%~��F���
��x�� d!�����%����\��(=�y	�HĮ�i��-_S���J�.F�.+�MǼ��k�0��%��Ņx��"@9y	�U�����`������� �nQ�k���%]/ŊoWV�Q}����Dk8��pK�h���v`��G�G	��?J�#�T���>��h�7�T�J�A��a.M6���ߣ	)�թ"��U8�/�bgU!���WQ�k_Z���Zu$�4���$ h`'}?V�3?�<b�۬�˷�yJ�����`��3�	�qa��+����&X
ӑ��W�9�_yY�'Ml�I>��@�}�_
�i�0x ��rm��K�h* ���U���5�����P���%I"{�y� ^N�f��3���aId� �,�ɽ���<�B�͸N]�4^�@ch� j��޳�FZU�#�����[��)1 ��C����r �r�e-�=���_hI�~���X(,������o������ `�|f�->Ka����?�\����-������ ��:a$��|�U��)��	��QEG9	S��)~ 1���{����'�d��0ң����A�<��Qo���衅N���� �d=��FP	^��?u)���gYT�� 	
�7���h'���P�S��`�)�EVi���C�/��}�����	�+R�0��}� �X�Ӧ��{	�p��Y�!�@V�i��x��'��#!_!���C�^A�a:n���B����$��ɑ��4~�+k�#V�<�
�?���	�B�,���+u��jT \�C��*�)X`܀|�� ��u� V���鸪I,p��1a��P(e�#�%��"�� מ)�����D`s��}UD#��t�{/0��`W�ŤP ��܁���\�/��_e�S�P��FS�3	�+�b�%��D�,�gV�`���ϱK$��(��w�O�L�0�' ���2�`#$�����aP�d�����-E	>w����?Vdl��K+쉴�_���L�tEō@����R	x���[Y�E��{�?*��D�0�[9't$bL��& ��(�;����b�'��]m�|�Kbl�3�� 7�NB�z�_�.�/n� �����y���u�`���%�T`�6т B8k�I �gA��m7ғCq 27Q�)P� �K�a+��*�N��ߤ�dvV�Qn)R�d9Xx',�I��K/�9��N���>��[`�K��A���j�J|'.&�ު=�*j��I`�Eǋ�HB��\E3�Q�������j��_������Jۢ���D����	��l=� 81�_5k��z��j�>��
�=��4 t0�2W�������0��-�_��j�>��O?���Nw�b!f�/ǿ�U��J�����[��b>��?}T }�3:��<K���C�f{��q�nPL�~ ���$�tZ��缈��5
#� ����^0%"%s(��r@+\���ۦ1SV�@|� ?�"Z����n)[\W'v/� LI�����ћ%x�������DH��	���&�y[�U�߮*I?��dKH�{��B����.8z�A���wl!���*��V���	�Y�`��ӫ0{�!a����b���`�j�)j�s�[�ץ.Pj�#�t��f����B��,sa�5]?�Cވ����=�+V�j_$���N0�iM� mq��1�\ITH�.a[/�ư��� �e�p��{� E-<�Wq�	>D��u�*	U�(����\�a�qP]wkH c��fպmN�����"��v��U�}+%w�o3��)_�XV{2��\n,R�Y U��Ǜ�v`&�~/�݁|a閬sqDL+_P�J�%`�$ ���4�"%�s���	��_`8�a�@u���"#1�X��t> �N�2��Q�]A�U��[�@����V�D%@���LKP��(l�	�U��"��\�?	V�-�j�7��I�i���Ӛ(�`:�Hz��+$J�-[�%�7O�[�Ǐ�M5Q���4[�ò�P�*�a�� �+k���;�j�GN����@�mA.<;�}A�q+�M;�Ѩ�g� Y�Pm�9 �!�@-S��{��q+�^#��8�.JʱJ��KnJ�{��T8��PQї΋�'���t��͂�1
�:%'Tuq��[��	��t�A1�i�_�#�oP�� ;_	��-�9x>������$�� ��#``-�%�����]\���@�j�� Pdp�)��-��H :l?׋K���C�7�.V}�F���e%�)���)���	�P`W8%�aN��,�{�ǽ�S>h�������Xz}@'#SM�ľ��<��{\�סe� �0�� M"�g�c_���}�8e!y��SYR��A�Y�b�@���S_N�K�(����yg>�+^%j��f�����, ����vq�L���@��/�^�s���؍/-:ڬ��(��K���|��w)�5����N�L��Sy�1��� ۹����ZXn蝀I٭��罘��@C����	�q��� �8vm���x%�����M���[��$����_!�t*%�g���~� �����M���`�ah%��.�&�)����R���_ '��o@��}ɚ�2�� S�|_�&N�S~�8#/]K�Y�U �Q�wِ�:�P��tQ�F �Y�\{��� a+��s>3�+V��F0S�� b��EXs�1ُ�^9Q2�	�� J򞷚�ZX�|v��5G��::�$؂�t
Qv����򦅪�c\h�]D�0�;JO���]���Z\\��\@�a@Ű%A'[��ƭ/uʩ���l\S��TF�Q�'I��1� �+Oa ����}3�8ޔ��z��l����	e�B��):\"K�y����"����^����PЪ)���B=#�;��A /�y���? �����?]���z':�2�A(�{�P�U?�{iN(���/�Njn0>��Ox���J]`��}��v�$�%�1!$�ǋ��	�3|C�I �zz�s�c����@�_�eO[�����O�5��i� E��E�O���E�%z�I�[y)������E4 �v�A�+�T`� Z۸\?�c:H�5$N �Wo���މt7U:axЗ�u�_�@#	0��K X����g�����O�.2��\�Q+��U�`~�i���Vw���"���?�~ f�CQ����/a	�qH��R��@�`@a[���3���k��:ni�� :�����O��"��F�HȩZ� ��4�Qz� �HϿ�s�x��� ������[��nfM;��d���t�i��}7�	��82�j�M��|Z��ğۏ�a̟U��/�BӶ���@`woZ�ȗW%�s��\3'���	�%<F �'���K��_���t��	Y	j�}®fJ�Q) �I�|��|Nr��� ɘ~?�/	[$W���VJ%�Z��	sO����n4%�TZpRπ���mA���.t��� ��?m�`3��Z_�x_�a���N%ym�����Kv�j?̽��rn�.�X��}�+i[0yI�L�<U��qg�����jz�����J&�V�[ k��������1O�$��@��Ӓ�0�����p���&�:�b��8A�s�?Z ��[�q	��J0���ڥ�(� d���_W�	�����*QI%dI����M�	��qJ��+�uK^����ѳ�I3�I�,�ˬ�:PLUG�`�3��<	�d���1�%QY��9K!�u��8 @�EF�:&^d���д0�[)�I�^�� �¯�`� ��Z�e�dK�?A�as."=)[7+�A\1�~$	��%Q�B�PͶ�w�e\w�E�j���BİM ��T�r���Pe�����t���Q(���@ xp�g���&p�&����N�	��x2��%[T�9�L�@%��p�q��`c���6F���|=�`���wn��_��p~r�eWJ$��Z����/�&�'��}1��){ޒ�� J݅6��{���q������!�ϵm�%mo�����_��E�"{�n;kqK�&�����+�ĉ�a pֈ�6�z� ~9�5�t�0��a��f���\�P��t�K���:ZK��{�e�/" `���a�vI�n9'���\���W/i�y�`��K_�ԁ�wK�� �HT�� �g_o~?�JV�1>j ��-[tZK��`P)��*Z_@l�%�a��OW퓏��% [���j��^��]�Ʉz�x;������`���ӵ�@?�$���5,h��.��T��WJP��J~�X.���6Nj0r�l���
�欗{0�� u�N!����*�h����	?����jr *��gW~�ۀ0�^�{������n	��p��c�b,�0Q����Uܕ�μ4k�/.-�?�7�<���?;g�F�|@���e��)I�[�*�C1�YUnm�������?�����P����-��@H��&'[8Tog�@/��d��Ҋ�W1n����'��ֻ�0��N���^na\�0���HJ_����J�r���@��̩CٯJ����+(�܈��?D1X��ϸ@�G�rt��JAV`Q�畾O(a�̟�9RT!w3a)�_G4����A��:$z����T�^�N��:l�] �+AT��cL#��J��_�J`�*���$��8r�_[k��9������	ؖ��P����	�p ,#�`��M�D��V�b��Ul�%�ɐX^�	��W�^��"J�c��M��n`�Xug���=	P������{���Yz%��o�������;�p(�t2���h�*-^�dj�n�"̯���Z%+fެ �!�x��/ ���y�()��V�<�D��P�?c�/��W��~BN``�.a uƁ�UAR[t��!��**���EZ���>�� ˜+Vҷ>_Z��9S�ഡ Ļf ӟ!�C���m3d`wl%�Nlΰe��P��˂��c?��t[	��Y�DGP�=�Z�'_�$�N������n�� E��m@ѫ{V�	�-P�%[_b�wFv)-A%QS�{�p�C B:Ƙ����^+�D��R��l�������aX/ �#�ѱX%���F9�� 6���9~P�1�:s� #v6{3��N[��̽IAk�z-%�j]M��d�YyGx��+�|U� m�	�%t<��b��P��ݿ�m���m^a;�%�������/ڻu�A<j*���7� ϛ7@;M�O�@��";�4rj;ۏ�_�������s�MD���������. �r���p��\Q!3�*D�j��ib����余�h /%�:g���&��,�5G��9%e1Yis�Rk�V)%,�� ��P��@2E؝_��.��r2�z��X#r����d�� �dWw��� ����V���+��o�H�pfI���տ6�=��Q+%���v.~p�51	��]9~.m�NŹ�(�����*-�fS y%�A��Hf�&�p�q�V���%����Ȋ�K���uu��Y$�- �a�ic� �^g�% �$׳�y�	�*��d+�P'� 3FpŎ��� ͌����o3���\f2�LIN�D��V�(º,���+2��V����e	�Z��ET}�Q�$�ؐ�XV��]�IR���Y�)XJ�ؕA`+ u�6� ���E���GFj��� ՏȒ��@��@-�U��@j3�OK�p���`��aY7���
냕	h�Y��p;�+�}���y#>�@��_|B�`���y�a�b��=��KNE�+ti�����%�������4���zp��[`�ـ��߄t� WVf	#�,K� �ޟ1�*�'�'���O�5m1Vq��
�p����{'f�p�J*�6�I$S�2_[Yc ��fmB4 ���Q��
�����,����s��@]&�>�FC.��N[��5��@��,�G��*OzV�����j��J|�!���>?#���`B���K�����,}��:�Մ�޳�f/Է� .�:��r{?�S#��+i�)��,�zZ|�/�Y��j��).���@W��_-PVd��|���i�[���O���+�q��)�R������q+ț���]@�Gk�'̓�j9���������	CeX�< �끽}	,`�[;Y� �L��CRt��5�2�_�Щ'�i2VO	�)Z�}���Kӹ]ܒ�QL�s�Oz�԰݊Hh���0`bX��m��NM������k����^�-��2f�i�Z_�! �[�V�����x���I�
��h����0v�	o{�p��N��P�E��`��t��?�Հ��J?�!�쏀�.@H��w�yZ�1�ݷ�����`�W�V�da��BҶ�(�� �0a���"�8 �9G�T�	�YA�,Af���?��[۲��u����½�$߽�� �2'WS�!%��1[0�g�"�ؖ�kx{Ex��$ʮ�)h���T���X�M�[��-V���Q�=[���	P���1���\�K��P����,V�}~��?������*�J0CR=|��s�5��ւ,;֓FdTu�E!��1�9'qj6O\ M	�^v�~��Y�o��������ѝQ�	�.��Y_��+����
T`Zm�`'r/^Q�6� ��%GT#+��pa'~ȥD��7�5C画�J�i��7�� ��Dv���j�-J"���f� ��}�K%�R�� �a[P21��1I#*��	�/�YA����l�@�A������ x	]��Ň� ˓ ���+>P��Z����*��+Y?�Z8�S�y�X�|Sȑ ����B;�߀1{��]0+�o�+��+5L�5���-�OA�HX���&��D����~ %�a7�o�����`��)�%��]�ʤ� B���i��Sm��1n �an�кZ�<� ���j����mDkg��N�,�Z��쿜��	�)�!���O��>���H��;aIg��P	��K�������;����£�,T�8cj��Ꮹ�	/�)�Q߉�ٮ?[���"���:�ї���)�Ȣ���X�����тMjnnP�iP��.�D| �*/���@ ͑e��(.P�cT �MփVZ��=ݤ��D�χ�«)��i��3�ߑ�+`U�����(��~�b�N��^�Xm ��Bq��[?ϻÂ!X�:ANU#S�𧏚�bi�q'[�aސ�Cӻ�"�1�0YoA�Y�����]f�BJ�7�A�;j���ܽP!_9�0��3 �G2\9D�"�~ ��MO+`)X���f���aJ_�F��Y���-Y�P� ���>3�ї#������V��c[+��2��)�Q1VWH������3+q�j���
�ٖӛ�dB���+Y��Ѣ�%O� V���t�6v�@U��/�A��bP�)�:��x�O,�ńc(8WW��uq�I<Z ���T9杈��A����~?��^�p?�(Z��%ˏ�{�������Cv���V]�sr�:����(�8�O �[�3��b�U������y�8t[�߼�_>�e �r��^�y'a���	f1��������:hdֲ9�nj �ٷ�W�dx8�N���$\��+�`�a&q�S������  0��a/�H׳%���֞���Zm}0���&�qF���RS%P��2��>��++qH�E�|�N
��1��	] Y��>R�9b���}��/��P�����(��D������%'!e�	��&��󉝥���+�Ԁ5���J	Ue<`Me����_�I��*���������6uOw@m��_�0��}_�;��S����M*[=�ܤ�p�w&PS2��#�zr�[��L��-���Q�C	&�;���@"h�0�p^�G�#.=3�˛����`Z���G��%��f��O	��n�T6p���q8�@O��lH�	Aе5J"�Z`��m@�E�#�YA�%anb'���֟��~�z����&�Vfk �Z:�J���k�3 �X��Fs�O��X�20����N��e1�z����V@�_>� �W�!�:]ha����*�\ĭ�ȑ�u�. ��_���x�٦!U����i�NGb�'���_��?��s֙��A�@@	�G�7�h��0u�	9i=!#�&܏�`S�?;�/i^D{ @]�s�%n��o�XnZ����� 6| ��P,�v��FO*'_/�,މ_�]�r�t��>xN�l7-�T�PB� ��g�	�$sa(³�Ws��N� {]?Ѩ<�G)Z�� uf��V��_��$Jj\v�^��q��	6}��fbib��:{���Oa/+��EþF$�q����.(&N����NجY%#��S��q���s�v���� �����\<��-v�%B�}=��B\� A�������!#�}�=��x)� A1>��:PJo�'���:$����f���6]��S{���V���Y'M_�Z�Bu[0}��i{� �{w����}`��MV�X�).��^����H�"(�-���$P��*T ����c{�-�6�S���U[��1k|E(O��P\ 4�B�܌���~	�[qv����AN�� �ykzL�� {j�/��@r�2u�
_�����[_m
d`����rjQ	������Q@>��p�������?J�#�}�-�_V�� W�A}�[�M�@��Ge�+��R�$|��c�.(�:����������h%��	Є_	�8�ӝ�+���!�y&�K�-`w��/�t		��0����5H#�%�S��*.8�B���	M�n|��@�����bX���q����ƈ��-������ ��W��=�'O�zbe����| fq���1��%�Sڧ[7P�� 8C�pNd�%���᰼�'�G��T~��!��n;#�����[��cq.O g�	��e%���_��t!b�6�+�J+�O��K&5�[9�	q��2�aKE;	(jUm��&��5H�t�ڎbB�\�¿�\�I���	�K�����јg���,ƕB��v{� �.3�0xyij��� b��K$�\
"G��	��ՎCv�R�5^�6�[�sp�>z��9�����`w���J`z�`����_
�����+|�� ��utL}��$��� .6Vp	��d��=���IP`ؿf(GaW����@�%@a�0�)�!i+i��O���3� (_�����t[Q����,�NɰM 5}j�*��[�t�a5�%�������/�b�V\�&R ��,3�U�,�СB�\p|��M"�p�r@�%q��T�;�� 
��� L/9%�(�Ḱe��.#aR2�[��U^<IߖB��G7L�%����T�@�wE�l+ȁ��7p�$�	61����M�݀�嘪�ݦ�s�y�C��[?���	�Iv*��#�9�p��	��or}E<χ��!Y�t�<@p���NĪ���R��	[n(�$1�H]��$�\�����?`�#�;�����gZ^ �_L��O P�/8N�'Qv$�Go4a�]��ӓ�A Sn<AG ���d�=.ղ	�h[q��[Fw��7�][1p�/%�V��<��I�%�ã��}J��Ԡ=�{H�kɕ >�вe'+����s�\gz�A{Y(�,_���QW���qV{��܎�I�<8$@�{ ��5�	VY#]�� ��}V.l�(�.� ��S���-[���gZ+��J�I"MH���o�n���		%:�AE/w��y�<U�O@�)��G�T�\_�W�&���1]m�T��P�J�_Q��Ҳ⍌(�`���0rW>�$b��P��I����sw`�:�tYME�9ݶ�%H����<�K����u$�T"E�HAf�za�T�� pl-����%I,��ގ� �oA���Z��p\���؀��a�jU�gW�� �����@S'
V��_��5R�ꛁ�qEC��9-h���ܿv.*�3r�����K:	J!}ο]���B���MP�a�^mI��^�m��)��"ku���[��{Q��7.�'���O"A���4.���m�V��W�-v�K��o�\��{�L��	( r��\���m-
<]�>>����W���@��7 �׋��Z;H�N�JS�d�+�3I*���?n�%���}�PtZ�Bj���3xxi(z����e���I�e! �th�l��PR���TL]�1P-@3 \N�e��~� ��0�Α���_X���S*�䪧�J������<���PSRՒ}7ĀF��Ŗc"� ������7��帀�*_?�F���,��Մp
�`R���uT:�Λ ��go�0`���>rt�4�@p��ֵ����a����N�����K��O�	��t̺ˊ	0LG��>S�]iY� ��W�Ύ�$d`�V��/����X u!��}���xc�����c%1sdн��כ��W�(���8b�m��h�ب.];�`��'{�C�_8"Cɥ|��[��K�G����T��^�5a�1��:����*Q�pD��,P�M��&��(������O�`<���)�]E���d���(-�,�
����5�(u�ܫ�]Di_�7��vW)���ZE�*���Ng H_����J����k��"�mkk�p����C|�Q��ݒ��<�\��ipn�o�(Si[��%����_�������^����Y� �-,��7�[�d #�����\�0��� Z�F��eo%d��5�'�|�����1`�]��vEa���	�R)DzwPԴ�1_a�	�Q� �z8�K��&�x��q��!8�O��r	�b�g��15��9�P��jMa�}��)����f.j� r��q����Q#'	7�	���+T�Q���z4�m���� ��)9��� ���h��@	�J����l�c^zW�� �;�6�i ��Ǌ����&��p���8���
�s�H'�H�YRm���h^��Ѓ# H�����w��{�"���p��q��杜�KwR"��^�"� �x�����K,���Σ�^d7U���� uI�4R���y s������8:, ��Iū�����	E�!iͫ�n2�H�b�7� )�?a�u'�;K ,�9�PO.1I0t��lg�� �Z;]7�{j���)B�\�F0�
s(z��|t� �_'O��i��]H���K�h��@� o�s}���rb���)��� �ބ^Cw���m�!�|^���6�Y�qKڻ@T�k�`��]�
 Ռ�3,��+<�v���i=���C�o J?lpڥ<[tؙ���L ��������-x] ���$�a��ћ���w��!y�%��/��x������0'!P��p�[��Q6�` �T�* n�:��Ӕ�e�x� �����Ӵ(�s��=������O������T@Y�$ ]��Q�,�h�  ���W��(^�� `dIR�D|� !Z��8�h�~������<k m��Y���~��L&ߎ���@Iܠ�E�\M=�ր!���� ?<H���]��P�Znmڠ8��I7;0X��=�۹�O!~ K2����n=8#� J i��(�<p��_! ��F����j5^�������z�X�9 �P�d��`�#�Q{ 2��b�/v�ZHX���|4,��z^5 ���x���H�� Z˙l�[�o��@%��A� +�;*Q�,��S9`�b��^���� �Lj�$��H��Q Q�LҀn��>�Fv �b{� P��{�Ty tF*�^b��rn���׶�SPU<��^���V�N ��o�]�hB6�p�`s�Z�����0\��T���n �?�D�� ;����J �1[���>��� ���( �VZ���YlS�]cL D}M�� s�d�� �;�l�} a��mPsH<3].NU��I�(�}� a�hB#� ���~�d��� Ǜj�Mlc1|H(���S �k��Nt�xA#��6���%0,��}*2H���m�0�j�g	@�!\������q� ��E#�K� ���L=���*����#&�1\v���_��©�OCQ#i�1u��m�� �[*�n"���xD#_�I���!ރ���&�az� �T�f�F#?g��E|;`h��0�Yy�ԇ�$�!:g$k�%C?�~ �N�o�R~9z��P�����ԡP`�e�@�a���s��_�V$P�P�4�ױ c_��X�% `˩؛�K+ e�����0�ay� 0�
�3�WP�`��,��H�ACؼ�����U }�!��� ��u@7�8��R�4��s ��w����� ��饉����!X�@���i ��"�CQg�h��9M�9��`?�DE ��9�d���H�o(��� >�*�c����<�����1��l��}	��Ó�� 8`�EW������/� �� �.�0������pXO���W3  ~��ٔ �vPgf<�L'�������7 ����[�� av0�{C������@���W��*�Vqp	��#�<�@Ӥ�����X���`�;?��#�'1��o�j< /��<�kq��[�1s@ x���G� �MP`fs?�;f�! �wL���Xÿ(\^�	r� �5��$ؠ ��ɨ���1o��Ӑ;��:0!�j���.�� k@��5`QJ���E`-�ʺDt���^�ר���f��` ñ�jb� ?������dPf0بO(�.��H��� %��h8) ��s�JI �Xh`*��=08;O�+B6&U@t�(�T���xv=-Sw5��V����'d�A���# ,� ;s��V�7�0�@���C(]Z��8&j��G<A�螱U,��h������㼨�Ĺ@M������-p�n��م� ����� ���_�!cŚ�4�a�#���]n���\ ����J�	��Ҙ~� ǰ���[`8����D�^��]Di T;�5����m��F�MHcv��	�-M ׽�_(���b�`�|A��`٪�� S�;'<T���F�*b�H��0b�{1~G��ۨ�ዔ J�g0 ��K�_HY$X��꾸�Ѹ��I0��<�����X1q�$cs��5�R��?�+\S��#� M�cp�D�M��� ^����
o�d�~F,D���3`�%#&ݑ `��� ߱����iIX �K?�N�#ܢ����݉<��d�FH���c��P�O�	��(^�y@ͮ��Hw��? h��<L�`�s��DQ]:�~� X�	�q&0<i1��� lI���X�L쿌M�cNs�@�Md�쎱��IG%��1@��g#i����*�J-�>"���F��ѣ�4���u���j��� L�;P�������5��Ԋ
@� $���F-:O�<R.���{�� Օg[z��O-%��q@<�d06XJh[�p�<��ċ�����x U�c�$j\:O�?�9��"�^��* �?�k�I�p���H氣��	 e�ʉ�:`���@:�h��K;��mtd�\i�=�� QP��[�T`>P� 5�������a9� ���� s��Z�
� E�'��: �r�l�=X�@��[ �
����>��X�#SԚY��� b��+E|��%�20E���`�'�$I�@�;ei K4~ߧ��9��a�ײTRH E��h��[=c6�`�4�f��ԂA��@C��r��p��;��Hݠ�쟀���� �M'�)pU��^FPR1,��쀫3)��"[��.��(d�+,�H2�|"�EY ��@�h�Foؚ��7���N� ���R] z�V�"��0��	����fp�C9��1�t�Ad�Q`ښ����S�`��qC�� X��*]	d��w+a!��%$�/��0o���%e�H�� (���]O�g�bV���i0�)� ��"��;�c&#(]��"l#�M�c#̀&+M��,�g!ope(�%1��ٸB	EF;��Њ=�$`0M������@�m�jn��*���q8q� �k�m�p&ں2�X��ը'�-@�K�.~�^$,���@=��\@L_��i� �I��Т$P�#����� �sc�(Jްa�@�� d0|A����0Eq��]�U�x�����=&ځ$$�mr�A�!�`u������f9����'t?�tۿ ���x�'�����?��P �8�P�2��g��FQW�<j�?ckq���9PCh�f�"L� o�t�I��dهf���πWAL$>�֒�n	�j�a��S�G������y�IJ����X�W�N>�����`	��d��$�{x= }���;�P�D`��|� 8��yw� �ҫ�{���<��u) ��%��P�d,���٨�b� L��!mw��uz.+��$dL`��#��6�l���T,܀�<��jL�+Z l�^Fp {���$�81��#��JA��)��T� Q�z��"���'c" E2��b��#�J��ӌb �f�3`#ޢ��`g��0GM_� y蠻h ��;մ/{ J^�8 ���V��� b/��:^� k�~��<3? e|��n��� ��,u�ʀ�Ĕ�[P1�O.�c �h˸� ����V����9 oq�L�܂ ����t��$}�~O� 2�1��(���e��<) �z�RX������:S��?\���+�@���E� d��2��|�)�
H��aCXR��@�y����۞��#� ����\��� 2)orF�4p"O}S���P��g�Zt?� m�4���2�FT{��	lh��u�7�*��BF ?#t�zV���	?�C�P�{Xnө�E�3���*y�6��~��J�&�0�* �9�#f�uX{s��k���؅� ��18\?Vly�e3_g����5^� ��{p<���斊���([p����s!������ ����Ӱ� F��Jm5� ��E���@ ������T<�Ѐ��F�gp���R�ܟ��4�6{kݡ|����1΢3g ��n�a�H� ��k����0�w�,�i�k��s��ڦ������D3nS����q~k�U#'f �����,�} ���!�#�� ��T�髇u 3ۉlQ��0H�� �]6k"����ڧ�߈P��^t��z!)g�� �E\#�Qa U�Vs�`�e�-|���]C�� ^�}
(,� �^Uq-�5<� P+�L�Go)Q�� N��
0��YW-�'ԋ5IQ�z أ��
��,�� ����� ����|{'=�o��Y��6��>� q�/2��7Q�O����#���}x�P�(x� �ދ�ɡ� m,lKׇ��~w(����@Tq�� R?��D�*T���A���n�� ڇ� ���0�[Z��T 6R����~��2w@�89 |D�3]�� �;���{U���� I�]�,�/ הg5Ys�����xDPԳAXeo��P߲���f��j��p��
��݈�W �Qm�-�}(�� x��6 ��ER����:N=�TT�6j�/��<W���)��z����� P6d-�jӱ�D\RN�Q� ���{G� ֗!�:Rj ����)ղ% r�4���R �J�_x�Q�:M����� 5��~L���@*�,l�sX ��?R���-�A4����%`�i6T	���a rPt�x�� $d}U8� ����� O�*P( �.���u~��h�C�H�A\ `sP��p�@'�W��&�\� ��d�r���	�U�$�py���!AO�F0�x �)C��w~	 �SQ'�W� �i�~*�{�?��y�T�jU����Rr0��	W��}'P@(e�m �"M�ۧHC9�R Y�ϲ b��o��r�w�n"Eց$����VY�)Uτ��r� x?(;RmY<'��=�7L�|� �������.	{_o/���xR�� $��� L��5NϜ
�z�%PШ}R ���Qt��0�'�E�����.|�� 6z��CQ��i�����0#�pw�( �OGHQ���3�]\8�+����H)9w ��<qV� �QxH��I] �k�ag��0,�6��9Q͠�R\����Sj�U����XBH˪����*�@Q�&��)FK���֝= }�1��p��Li� _b�P�tN��ك���q�~�?�cU6�����.`!�*Z^�v��9Ò )fN���:'P	��L�����,,�%DE}�Mf@�N ���2@h����XI��w@T ^�YE�P�0`��� ��G��O6 �Q@H�I� �Rs����y :��|�� �Tq�-s/�EQ\�A ą_�� 'M�+@J� �73)�2[�	�P�O	4�d��=�v?yT�����*$= ���B ݔ������ �t	��M�3fU։  �l������|��Ђb �[�4<FA`)�sh��x/w�;�|`��o �ݯQJ�Y��%�7����.`U8��o��H��xz� Dp~�f�<�]�R6�qѫ�"nK-��¸`�A ��t����+ }WD�X�F �Uh@��H�HB4>3A �����d�����|[4!�0l�Rx�5�`�-�',>v� Լ��;�E��TQF�h�$���(� �Wm��퐢������@ڮQz� 9k계F�6P|��1`�0!Q����o� ��`ɲ| ,���=���{Qg�wP��(�W��?Kђ,� �.M����= �ԫ��PbZ ����,G��X�ܺpq)��:�Rr&�
h /Gȷ� ���(>m^� �w��|ԯ����CgU?�_9��+�<&�ϴ�͡,O0�� �RÆ��H*.� 2��|!�4�W \�R��@c��b%uDB|�@�� �㹱n{§&�"� JY�T�b�Că��������HM��@��P�]^��|�2�/�z۶<�|>�RФ�f�Y}��=
�[�����H�0�K��4=�V,� �s���|���HkWy�P�	��4& ���f}�S� �*v����Q�(Dd���e}' ٿ����p4����F@T�R n�b:~�(|J�r(���=� Q[��R���H���������@�^xt P�jN��L� �ܒ�� �ĴH�Y#� ��Qm�q<�n '�)ɫѲ�~|�Pe�??	�'2�8� �P�ْ�J06�
`�`�  �}y����Y�v|�<�� 	�)�L������m@�KE��PP�Y&v:8ta����2� `�<�Sh� ����Uq���C#��Q@�r�=�����:_�Q '`0�{�2`����ܧ �+*���3K��4��z=0 ���#��ܸY�<XT�,nHԋ{� o�6� j��x۞��s�;>���2� R��; �yr�P}Y �۾��+��q� �Q���R� ���>���;�u����*��D�Q���r� �Ɯ��*�&�t@?��R@>��À,WT c¬���MŘ� .-��~b�@0�(����'d}���`��vy)`5�U��L���� 	�C��&}PH~9@��|S�1 ��RH-�� ���NO �ܼ	+�[�xB{���'ƫHt�T�ř�X��>(3:k,]P�i P����h	a<�2q|�$i zk.L�!��� {�|�����z�e�`k�< )�}�8 yRa��P!���F����),R�Q���nE�� ���q�X� �eܠ�k����=��t�3��&�wt�īBe�lV$�� l%rP�� �W6�����ޅ1��ł�a��W� eUk�g�6���C��[ ��Z �� Hy�R)m}� 3?��0�D8Eݧ�=R��yo>o� g˅X΀ �}��ܲ��A(:Lz&��h�� ��=��c��p�<� X�5���� �.�Z~�ǘ|FI�,�".(K4�H�i�d�3��lr�Ο��0pD�Q]����^Lh�H� �1$�|U� %s�:CQ3 ����-�� D��Jݷi o�«�h����zQ �M��P�01}j OF� ��i�S��� RGg+T�4ܓ���lj��ia V}Ne����*���WH&�� i�{�G�:
�B݌= ��WJ�;l
�&��� �m��IT�Z)���h^S��{ͮ���9� �ӿ�0*�ME!�� ��KANl����@�ݤ�>� Ud[��z�� ���N&���0��pp ��BqR.\� ȫ"Pa[�`��3Fʿ$u)�ƣ�@�C�n
W��8��S��+��;�T��Ц�sU?Bb	+�F����� �[��{߸O��|���ʍP�� ���_�)$>� 	�q(����G�m� ���(WAb�|���v���݃8,�k� ��}�V�;��P5������ӎ���!$ ��vL�� T���B���t��� <I'M�� Qf���C�|��-����D���S� 4�U=�0���6�C��8��Y���.�: ��֔9=T^H���1v ���H�t��Ȁı)�� VX�t�|� ��y�o@CF
�����$ �!��:�	��yt�@Xz+.'G�3��`\��&|j�RC0�\m� 7�r�5��(���Q	��-�D\p:� �2���� ��?޶Q+(��@5��~.�� {�ȵ\ X���YPF]:�Ҏ|�b��P橾& ��/�jQ�Rm�6��X��.��B�?-#� �[A${?R��K���xg �����fx%p]&���:���+* k��V���0�� <�+��� ДܖP}����<q�|�2 ��A6RV�����peQpH9���d���9ʤ�	�G�:��[! dg'�,��c���k/\Q`F��mZ@�K}��< ~��z����oӀ���L�n��8Rwe�Fs.�:@	���h7�N ��{+������i�KX�*,.UQH���(V����R�� P��G��K �a���� %��
'�DmK��ܨ� �a�Z�t��|�� ��#��]c �r��X)Q�,.���`h&:G�0�@|=m*���� ۋ���W�%q�hq�t� D+˝�	 �F#"Q': ��O�|�
/ ^�]���# J?�2� FQ>-��L��:'��|*�@���R9w�Q$���:�p��|��~�(21+�ZPm�`zW K�(��[.�1����>�O}�R�~�xf� �T�3�W��ܞ�@�.9���H%>(A 럋��a� }]<��Eu� �?l�Q�N8P'( 8̌���v ���T�z�iya���I �X`�Ǣ �ܳV<�|� ���	
b�R �ܵ!C��q�LΧ8� �{���~$V�&, ƩT/:}d,F�$0(�q)�b?�����Rk�7Q�td� -��ڶ�[��꫷��0��a�T8Ƒ��� l�n�К#!�f {��J�iQ�*��x�l� �K��{s� z��to�x^Ra����`8Κ �1wr�8� mٵR�֣�^~HЮ
p9��d	r;��mʉ ���IrV�M ����ks�,y�:��$�� R$��[��{)�:� ��PK=��?�	6	}RSX��� r޳*�b ���pl��Q�"+k��A��P���� ��#�>�^�d|� P��'�e������Lz=�@� �0HmQ� 
ӫ.7���%RW�����ˮ�h��T�\� r��w�$��\L�K �7m�8���w��|}�i�*����M)�, �Cč�@6�U=�ޙٓ��p�9�$��0��N����ܨ@�U��R	��ր�J�<�-���`@�d Ev:�|
���Z�0w* �����#� Qy��i������ ѓ�#*��Q��XPҦF �����(|<���G��t �_z���Q �A��-ښk�|T��������3�G�����.Apo�.8{ �;yl ��3&�*�
��� ���8o�{�m�x+|�`�����>y��۴K�l%������ h���4�&?�Tb������e�O,}� �R��KT���)//<�l�[��PE؈t��Jk�R�Å���~-�g�%��S/��U��FH`�R��A���Qc���px�{�@��� GIQ1�" ��}�;ym(Eݥ 5HQ �����pe�dt�������0j._Q<0n;JL����.��@�#�� W���$�G彦�$k>�}�1� �,����MP8 T�0�{���Rt �Q�y��`0���� �;�P���!�R�ܠ> ��x=��U �/�Ģ�P�HCIQl�m�T�$|� +���{�v��� ��E�- �ca��,ܴ�� C�F	 jݖP����_�b'�}P>�/E:�+p�l� Hwv��d�m�u}��l-�4 �.��Hj�R�,|�_�b:������ �+�c�q hu{R9�< H ��r�`��0	ТN� ��Ǫ� �w�Q��*T	FG�<�{��vʩ�ԁ�Tݫ �/P:<��~�.�n �� ��� �+0�b\��l�!w[
�* �����8�s��^Xr�L�h�>�S��UA�m ����p CvP�ܺ��r� �/yދ���%�J�0_[ vր�#��`�@��| �M����>Rق�J��@�$����	��A��6�,R=� Ι�����@�|U�pDR �XE��r�~?�� �0�^X	]�'��qL������ڌ�Dv��
� .�d��� �1��yR�x����"[�I�ܠ���X�|�9�D�R).�ƨ6�`�&p��� P�/1�D�R)�π�n�W�>��L0Z&���`��iJ:�3B�V�����+�����X,-�S��Rj�k�) ։?�ʚ���#B��@��S �%wP�5��y��\�U�W�P�B�<��zR�*�x;"���V�����ẽ����n�@�ڰ��,	
�� l#��]�H�lw8T�UF��������#���@ظ;�*�Pq���� hC�=�� w`��R�A�Ugx��`��Pt}�Sn��sp�Ǭ�]����� 1��yT^�AC@[�+pG-�PU���h�T� �&��� W���ּ�ܞ�`(?��
�ɜ��9 �Z����+}6O��R'�@To8 ��J�[���`c�/�t �3��Q�:,��lێ�<�C�$܀�i�H����Q}u9}��tl�\<�e�6�ï��{�#)��,��[�>�`�U��|.�*��_wj'|�P�� �L�(��B�}N�ۿ؟@z�.� �U�6Qo�$A��|㠆���P8Q��7��&�� ]�|}�%𢣘�.���а;�HX�5IH�(K� ��%Y"��d wۜ���@	H�(� v�QK�K���̵�l�� �zAK@���|���!t����� �3�|.���2�/]@h�9������'���zϷo�`dDFt� ��1�����;�oC��􈺅 �nYU��q,��<0Ht�	�l���p� �Qa����H }2��|T�	P��ப�w�X�,me�^�}3�*���4,Q ���m��R u�TM�; ˈ"Q��Xm b�1�@�PsH �Rpʦ�ͱ����Ę��U�x@����(�HJӼ� JCQ�6�P��t �L)�߈\P
�D
���D��@鰸/�{�AQ@�0��5 Ӻ"�bR���O|-G�t�H��I]�ҫ�xk%�`��� y}�ڭ�G� ��.O� Q�۱��B<���|������������,m��gۀ����oP�� �dU\	X.� �wv����o��z �����Q���G�Υ�R
(���ڋ8 ��+z��9k%?v)]0��6\�d��߀q�{�~���\�^PJ;f�j ���0�x����O	k�̚�(��`L1���K#~?��P Px �+H��G��J8%QT*����A�������?g� �S�(��k� �F��N�| �ܧ��V�zG8{����\h/4 ��2��i}~X	�&�� �QJ���y�VI$��������b*�ޱ`(�:�;���_ճ�+�R`�b)���P ��;n� �8};�e]P,�K "���C$RP�gUk�<]s����F�Dj@8΋5NQ��Ly�� bE��I��s� �W� (�E��� R����4=�}�9�; �k�.�X#��\��� ZQXb��l;d �q�/ E��'��$��8�:,���TP� �`�IX�x�U�ۼP_�`Ѐ�\HY��,�@��|����5��� (O%��d� v�R�9q�I ��w�:���P�-y�
f��> 9v���FC��ܳ��pD� �Tj�E�F�L\��a	��O19I'&��d��<�T����\k�`���*P�R�# _x��X٘�� T�'A]=���vf{�@Q(̤���� �%?zqU3L'��h`� ��>\$N�����v�H�<��j�FN��@�g��9 �,6�����#��CTE)�?��_�U>}���� ��SQ{�%�D'f��(y�H!��G�ЀQ)tB&�A� �v� ����ߥ��/�Ra���ʹ��Jk��`� aN��(�H_��'��U��������5:ܲs���z����0? Rh�|�5��
Z<��� �#���?x�A+��)� �(���L���Y1���	�ZH P$������ۨR��a���ś ����{Rצ.����t;x.X/�c6��0��|� �=*���|�� �l?���*�Q"$��s�Ɔ`#p��p}@�B���ک�Sj�wP���ٻpհH� *���=�Z��́[P���n�t���b`ۘ&��G�;���ڈ�;+R�{p�p��<p^��X����� �PQ̅]@������j 4�>��7��������p`� �L�'*u۾� H����- ��9Rӯ �Hҏ��k�'QG�\�y|�� �Ru�hL: �/��j�� q���|�� A��~R$lx6�c�D�)��"pH0�| &������U�����M��~
���3��&�� X���H*$�=���`'�v�H�KXH�� \�!@��X<E�}���ؐ+�Q�;�p�� RÕɢf}�#� ��ROu�o�4�dE� ���� ��&���:  ��*�<�H@�k�Q �a��r|b�o}����d��S�RHp$�sC�,���� ���>�� ��0nQ�1H�( ��������R���"�0Sd/��i#��� 
{Ia������R,t��� >ݲ��
� 4���8�%�Pk�t�uR�� �䃄H�Ā'WP�o���D}���{���� �+P�L�«� U/3���E`	����T�ZG)��O{#����Ik>X�#;"!�0��Y�� \Dm���x�RVW~���Ϭ�^p�6|��-'8p.��v ze�U�6�hZ�%@�tǏ �n"VqP�� �R+`�� ���1}�E� ��*�'�J���P{yFW(=� t�	+��O�d�i�h���``�|�t���� ����� ��OjdU��� ��x�/���\Y(~Ï�6*��T&�ӄ=<,	�Sp\J!tе> ���MQm��� �̈�.}'	#��� i�/����88�Rs�!��`0�ˀ��.��t �\��b����� >�ߜ�D�j �(�ur�3����#xR �7��W���H��(���?w�l <���(�Q��!�)�]O�>3���0� }@m���o�Q�6Y � sݧT��5j {�#��
.Т� MTj� \å����.q��d�Q�б���l��k������U�u �j��[0�(J��2'8�`���gǇ���mP
��_��)�\�(	/0�@� �P���R�q���H�4�ہlǡ& �˸��+t�	b���D�2�=�$Lh !�p�"����h�P��یKX#*��\ 0��0�c�;�$0d s��lC1KS!���~A�T�GHP�R,]ش ��\���J?4 $�$�˾������^!��עO�ldP��*Q l	,��P���W9ܔu��2��q0�%Me|R� ,b��E�0��0_��p����'��@��N8Qo�R��������>q*.O��@nlQsV��� �g*��
� ޴{��q��XR��N��� ��3G�������uKJ`i���� aUFΙ��{y���4f��� ��g�����$�&�	�M�9� ���J�}~ �E��n�ͪPܨ\������x�vPb�Y��ӳ����|� �.�&�� ߴD����w`_)H���!+J��_��(��*�(ZIs��	�"T�BaG{��@(��*֖�Lh���`d�@�����%B����-*J_L s��B'��1�dS���@(�u����+�I�1H#]��`(/+'b��� Ad�� YKo-��� Dj
�Ux�\.� T�N���j��~ ��>H��sp*pk�hƢi �3 C�19W-�4 ����f/��y�+��M�*��? ���snJ��[}&�'��D�:/ �5��?�*�� W$k;[^|um ���{�D�.a�ϵ�
uL�+�a�6��u4H"��}f�!m��%�/�H%�HpGR�ܻ�� ���$� ߬��XP�	̨D݀���s@�@?�^�@EX��x6�w��ډ�x�=�����Q ��Z	�21\�� �E�H��� ��=��})�� /���[�N�4@Q������2�?���>ԘƉO �Tz�\�'?t�0w�<`U 5�bj'�R�\�S @¾�D-�r@pKO�k��0�o?^��� ����I����lvs�\�)2�,Չ� w��1���_�H/��8�?��Q��`�(��^-�� 
�����
�ꫤ� �NwP��>r *U��t������_H�^d |ʉ�F�@ݏ �ۼ�ĸ< �2�r�4]P�\�4�%UJ��)� �4��]9��%��x����0;̄���}�ޓ����l��P��Rm �,T�:V3��N���яB8#l<�`R�5�� JY:��et�	zoQ0H�*pG�P�l^��� ���;�5��A�R:+� ���qX=���*}T������|��� Q
�@�� �\^�i.� ��*�!;, �O��>R����Өw�l'5ʀ�,v� �[�"Q��c�ٌ��)�u,}d/��O$�Jm`'�� �R���Z� �|�)ܤ ��A�U�<�P�� P���N�5�7p��iŁ�� � ���� �R��] ,��~�2v/<uz���|0���=�P���3g}���Ef���R%n�_m��8=�U*\
(@�� �m��� �z�ho+���:�8�.Qf�/@��>�� �\�����:,9�|RG-7��	}!��V����]�z��;	�~�
e�� ���qչ���@H� F4�5L	�R oe�k�V-u�.Z� *'ǕR�hDQ]&�����1��,�-p�+ ����Q*� ������Ԫ���� �mK��B��JS�� �2�P|��Ӑ��� ��)O�[/@P�ħ�P n�hdj��>-}R*�O �Q4��{ :�bUD�E�?�Ӂ#��y��/$w	W���.ho�p�f���W�< <ܿ�> (��V1�K J�R�%�-s�x*�a��"�0�`�wy�J�����H��*Lh��� %!�	�S���5�O���� �09RU�Wg_�vJ��p�J����/ �6<�z%x e܇�=aR�.`��8JH�(b��R_��ʣ�j�'ګ���8�҈Xh��D��$�'�d���������b5i�0��!��eI��ʌT~=��)̆�CJ E#�ͬ�a]������E��  X�\��k@�-?
w�T'�P!��@p�H�����m��w=�N'������ ��䔰f>�d ��P�fR~F-��ʸ���U�z@D�P&��� �.�� �5�OxSܵ14�.h`R۾`� ����}���
t�� ��S�$H�CQK��`�q�g��5$0�p�ߺ ���Ƅ8Q��WF�M\ۜ�I|�!~Y�"4�  {�-L�%���� �PKf���D~|���{�S4��HT�n��r�`E��{�8ܒ��4@$�[(p�����OT/H�2�|��G�*��p���>�i�`��_�4�N 6�1�?H�H8��
7�R o�P6�<�Z�ަA����j�$�����a�?�H��<�T'Q�`��
|�:�������q���`C��� ��new��ģD^�'R��9#�8I �X>��4�p!XTx����B��tT��|��=N09^���q,|���/�"�����NT-}���WET��(<�4�= JV6�_&��0���� �^\+f�4�R��-�{�ce���ߐ�d}S��-��Z�P� g)k
����v�,8���EIN� B�$�|&��$B�yx�3h�y��Q*�hk��IhX�� ��X@�]}D�ҙhReH*$9��qp���'$��4��hl+i8Q ?l���ӡ� �� m�;S�6�"���ۉU���27�|�;�l�ܸ,�1k�PH�G�*dJ���a(`,�$D�� �0HA�M �	P-�<!� ��%�.� ��U�(�	�R�Q�ƌ�OK'qhcD(��֠2Qj�S XJ�*�y�頌2 T��,-X��L��Q��A�Ȭ� ��&�R*��s
�;�����@l �z�b�>HMQ9� �C}cL�h�
 �I�Po6M���E���x���� ��%�y�-��`�?�S �\���_�i���>NW��;���������0X� �~������ Q��Kl�=�� b�P*�� [�4"���-�Bhu (�lQ ��k�sfq�(����T�-,1;�H
�� 	�AcU�yp4��%Xm@�t�4�U	�1���9��ҲC�}� �z�S�$wPm�� VisgO���x9�&������N@�f6�ڱ,l�?HxPb�"J@l3N%D�P��LG��8&`��R�\�Ӏ�s�s+K�Lp,y]P蝨U�%@l�+9�}��fcI����&aӠ�Yh�P�|G�.}�q�)x ���䷡���kԔB�;0�f|!�{q�W���J ��[p�D(�a���� "�|\~������F]J" $�|@�fd��D�l|�:����|��т�\��+�dܶXhq�#��9D]6N#A����c�(R�t���2"TTb
�|40�>�2�\����)V�$� 4��K`��J�i���T��9p�d'�,t�W�+��������"�XR�1�Ժ<�`GM�ʻ aUJO0�	 ���L�9{	�eW��o`��Z� �nQ�.G��Z�������O������B��+ DQ-�w� ��*�l�!��`PR_n�P�ǈL��������m.�=Zn.���R �"i^
���Cݡ0�ې5�O᪽�(�� �ki�?�#��NL�h%	+��K2�w�U�N��:p�ܺ��X���Ǐ6�g{ jQ�� *G4�A�v�� �#݉M<�H [�JQ���,8��I .�����x� H���ʱ� �}<�~���@Ni]*�N�FQ�nPM.�6���@��K�� !�����t" h?R\��SM�	���t$H����У�h� PQ�b�>DqO�AE�,��0
]����+  QùMN����x�ӑ> �|�Hh���J�5�H
� �IĄ�"�@�G��@�	�J�dI��iCZU�,�U�	tP��$� ��Q'�� �7���%.� �r���X8 �I{�R���N��t��,�,�X�WD���z�Q��,�� F@T�
1[�6�(+��dU@��P$%F K��|�3��{� �y'�:R��8Tm� {�x��D������В )�|�JM����Q^���( WaJ�}�����yЗL�Z���/ �����	�<����K!��8�mBl�s)�tp^ ������8� �ٽ�rP�	�3 �ˤ0}`?p�Wlk4�b��\@���	��<�O\�'x� r�q)ӱ\�&�/�P�QJ�GU��:����� �Hn�Dȫ0�Q-w�� �6Z 5ܳ�g
M|�Q��i@�	�@H�Pׄ��l��(��+M��A�:��d/��]�v������fDܷ ,1��wF�:��l��X��@
���0p\�$��ӂ����� ܶ�b2���0�
4��U�	�@l@ �+�V��Wdv O�z���(JQ������	��I] ֟)yR lTvM��B (�+#���os�H������0��<A44�ؐ&�r�E�"ВFh$Q�`�Nk��}� ���&v���:� Rf`O̩���H�� ��
��"nM#L�p/�����<|2� (*N}0G�.�;8�Q����5J��Ȯ7�oHX��-z ��Y�x@� 
L� �Q{%; k��)+Z�W&�|�� �h����`Àf>��	�،#�|u й& W�[8�7� �բR��h�����?E|���vu*O羉���`�b�|�HY� A��|�����lx�Sk��u��ā������!4@Q�p�0,�+�<����h
 R��ʹ Lϯ��+Q �e���RT}�`��%��-z3p?��,��J�������LC���;<�ʀ�b̸*u@yn�F�}=���ţq4�a�3��tVK}�� ���� �([���~.��`��R��ؓ� γo���Z� Й�7�b� zRi9�ª�o||E� ��hUݑH����{R>j�5�V�~�|�*��aN�ȣ�0�Rp�@�)}B��<b�1C� �Kv�3HpoQ����Ԭ ��������0u@�.5��@������W���k ��"��|[�2�v�0����͜#w�+��*�� ��E�Pm,>V��� �ōRO�HB�Gj�����C0�F~�X��}� Lp�'<��81-{z�%�;I���e����h�(� �`�}t;s��KDg���I�ș�0 .�*�٣�E��^pnq,A�YFtHJ.` �}U�$����hi�<&�(S�Ħ� �p�x����[�(�P_ �5�*W�� }�+��� |Ymt�@������1
�TLY~������o����P��*	pH�T�(?��)��~� l
��RH��=���6@8ыh	�����r9RV<�!�x|J��3?x�p)Y��,f���  �J�}���|����$��� �����-�Q?�q�RV:��ʲ�< �O�껬Ë.�P,(<�,4"�6�Bg�ˮ��|����k�(�n�V`|B���އ`�^T��>���d ��E��$,e����k�f@4���HLԼ�=h��Tqp��̾���d�W8�S�lQ�����0� -x� D#4J���.�� �ް 
f�h�ό�<ڞ��I� ٫�v0 +�WZ=�o�8���tz]��_��H��Dcr 70}�6N}l ܣS����\(�0�'Pو@r�"I �ɐ��d	���Kxhu�(�]� ��!�{���Mv�H �b���?%��4H���7 ���2������0?�|�!�E�F��('�Kŵ�����,2h��[+� ��z�Q]� ��9%y R�ǆh�Hb[$��g�*�M���Rs �c�f���ZD�8+�*} W/mK�J|�pP �0����?��^�ݐ�  ���K�Q�6� ��:��Txmt
 0ybR�����XPl��ꈆH�JN��Ԥ�����r� 'M�)]� ��&y(���Q���R������9 �����T:,N7�l�� A��*i� ࡾC݀3wO��J.����UuƤb��|j� .�(��¨�[�$H�� �UV�-�|cy� 7r�Xj_۰�  5��H��R��|��N�vz���+ ���+w�4
�P���0�� T(�u�ۮ��!����n ��VQ �����\ �ۄoG�s� N�|?�k�U�j 
PI 631�L$��|�ݶ>��p`� ��{R�	 �'W�2�|,d���j�$D	}�>�
  	���P �`��|��p�� �n}�D��� :x_P�d��w�#b/�B� ����V�+��n��Rak�K���x �����5 � �ٓ�n)8��&�4}�@�	�q*��L;'��n~R���%��	>�T� �c���Ls�@�i��`��tΤ���.(�h*� �J�Pt�������@%�$f)<;0��}Q� ��%i�NV�l� LΊ���9z��&�l< h���,��]��%�`�&�[6�� ����3\p2[�F8�m��1�nE����Q�Z����+�ABcB�_0��� +L�ۍ� 2 }l��:�- �G�������QJ��0�B\�� ��z9�U��w�+��P ��p= �"{� �Z�����P@V�5H�Q�qF� "�< �܋Y��8�ߏژD��� �^Px�� T�96�Lݺ a��g�|�*�`9�/Qr�JҪ�,iѡ�`�qN} ^�;k��P�%@T_ �Y*�n	��<�t��KИh����pD��dR t����s��pH/��*Qj`Ɔ��
PF�w �7ًK� 1�)oQh�MH�= �����D����+��p�gCm���� {�$�c�U *��,��x��4Y��X�|U_�py�m��g���(��/ G��"LQI'�<���E����$;�a� ��"��P� %V���~���4ec��{l����۫�R��K\`����|PT��?� H���V%8 D�Rk�2� 1~rJ}�� ���5�����RS���Ҥ� h
1���H��(V��\�#�Q���K��@��5��� 0O�R,Wgd9~7�t��� ���K���*]�s�ن0�6 �pcEz:��>݂��Xn�p�3�QI b`y�ݟ� J��������v��WjO0����" �J�u}L��PL?�yG#6	��`I��{F�~�.T��|8�)�5�>��ڢ� R��A@P�|p^������l��
`l6Ðl ��,Rf�� ���۲� Z@�emN��jnQk��Ϸ��@�}*Z*ˀ!�P�����ŕ�� YS����� ��b�o%>,%��XDź�(�Ɉ���+܁���`xƦS0'(��P�����Z�[c-�)_���*�i(T����=�J�" �'�Mm쨮 5�A��֩D,��I� �_�!�e�^���aQ���Q�L��� 1���"k/���!�x��,� K�[,�W�{�4�˅0V��D,�i�������0���s�����K,`Ց@��9�V�Lp{j�&T���yT�0�`���(�!�, M����t�wN���w���� � 2(O���� �e�ؖ�>�� F�k��� �zEW�`P� �h�_vi{�� \�`�s�o p�6��k��@���A��{U�aw��W>p��o��" @�Q�νF,��vW%b��wa�n� e��m�O�W�]8��+i���U��`�� ^)�0RJ�_�������? �������Z\1B� E'��XL2�N��,0�̀e)?W
�y@'�����U>!���c -Q�A�|�h9��=���Ǫ����D#ط�y� V0�'��t�S�ǃ�rjd@I���[� ��#��~�* E�7��4:�Y� �&�9�� ɕ�Ӝk��">�����R�Ƚ'� P���T��$�̓;�� �']2�Ďy���Ox:���&rQ�;�T}.? C�s�F;��m+e&�1��w1�� �@`�_(˼ WN5����0a78r�] ���9}�FX�0:;^��DȏrC ��U�7�s�� ��j`�11�K� �x���� ;J�:2� ��[*x��� qD��7yPTH>�〩�8r^J�8�6:�����;܆3�t���`%Q ���
�Z3� ^��6�`#)SȐ �b@��>"?Ilu��J)H�a#��YС���_u�p� �� �sDy���Z �<���˕	�WmS�G��0$�(&�dx�Qg���5��� ��ԩ	-0�.�H�)�]��2���E��! F\L�w�)3}A�!cDt��`�=_��%
 ��6�w}�7ꅡ��j���@��H,���OiY�<&�K]0�� ��`ys�o+J  U�Xw��_L�%#P�)@�U9�H]�c0N@G� !� ���K��f ͵v��G��AD�� ����!��qL 0I�'��P�4&Z�#/�I��L�΂��� 	C<�󷼎����H�7s�.Ni�ؗ1�Jt$,�����5��� ��g^�)[��M �8~��4�}E)- ª0:�*\�8�X�< �۔��Z/�� �6�<��w�vM����ʚ\	t����{ �0���e� 
pyZg�i4��@h&+�h;M�K��-��tIk����\��|���0;�F]�Ad�@���9?u&�$}� ������Y�Z�����;�]�� g��#шP��S��'V�s4���\+�&s1��*1�;���� ѿ�f�S�
��t%�����F��h>L�1~�!Dk9�hH����H��GTr&z�pY*�*�L� �������SA�LׅB������T�F�C� �⾢��!�h@�0���l ?kt'�7������w������� `���SG2zb(̋�|�2%Q`[���`��!i���>�V��7����3�����H�Z����?���&�wt�)�TB�K >��k���?�ف�%��H���`o��i��X�I�k�����E �S�7gs�X�k���P ���C� �ݰ�w�踑�&"'e`x��Z�ǑQ=[8Iʴ*_��<y��Bqy�������@�-�0�*��*�� �}�.�y ���u��DR�49���>�p 8C�:����\� �
5��q�r� ���6�@�p�AX��r�"_�Mx>v}
�m4Έ�H�M�I��`O!�j, ��rpC Ls�y�%��|�HW�X�`��E"�ab0�p��\�.؄� �-1�5 �Z����8���B �P�m,#A�>�E]!�N������� ���WC����<t�.�/��uJ����gâ]} ��"��fcW0{ A�b�P���M�_��#v��������N֛I�غ��s�	� pZ+� ��e):���\��L�A� �Gl>#�xj(�`\o���=&F C!�L<�� ��1w0��x���ܩe=�c� �(�;,L W��`�:ے z����U��w� d�Z�� S��R�2� ��Ot�_� �:�M"�� ������R w�:�{2��tD�^�P�-�0 ��TZq"3n���`��컄e>�#��i ��1��A�� �
a���K�|�_p�Њ�M�A(�oĆap�|7 ���0\C�9| w-@�$�x� T)b�ĀXA9*�:P�o���\<�"�A[8;Nr`��@�$�}@AÖ�\�>X��ʐ(P0�h��D+��ƊB��/��t?�qw@��2�#)y~^�+�GU (�@��o�#z�{9e.q$0zL�߻�#1�+��֎�@��� �Q4q�߂Z�'0 h�ET�X���w(:��D��*��(!\d�$��� `L�����X`K�'N���I wG#�Y� Az��]�H��tj���X&|��#*[yx#X���R��̖x@��ĐG"44N�$TH��n�ME�>>������T�V't��OɆm����� }����|`�ߒ�gg2� o!e
Z�輁���Ձ�������Mw���:�Z���!bG�w/i�������(���HHw6ھh
VЖ���(ÆE1�
���Y�X�@&��� �?h�k�$H7vLI:@�DW�Ƙ��k���>2[d�9!h�Tb����^Ip�D�Ax*��Z2�@�P�#t�����!Z�v�B���� $�%���Z1ݗF%��� �#_���mf1�y]��A�l��w5|JUO���1�0q@��N�k��h��iD� �w�^��\ y��.�lZV�s��$�Ċ)�H�=��( ��s\���<xXCj��kۛ�R8� ��9�@y�����>z� ,B%C��[~IM=\ ��3�x��{ ��ɵv� �3c��h60E�`�Hk`'I^r	4�/��n�Qi��0�� f4WY�3V�[q5����p)1k�ELZ���5U��S��f T��k�"�,�;7U ` ޏw� B�E�5=J�q�m��o�`L�fh!?4��i�� �!ް �E�31�Q 4���c �����U"�։#*� ��1��� �jxr��l`"�)\@��m,S4� �=-%�_v�� H���O�,�<��� �� ���T
i'r`�:�mp��F�&�u�� <egSl|.�����MJH� ��4���)�}��_>������!�y)�'`���,J �L���-����� � M%K`:X�=7)�y�ˀ&��o���^�C�pBdF�?��p0���o�M0s����0	�!ϷL<�K +��j :v$����z녙˺�O��H�e�� ��'��4��1>�@�Qn��ev��!��=G�
�`�* ; �Dvp��=�: P!�bП����8�|��)�:��Tz���6I���\{t��`4cÔ��̃� �(Ey�^/�g�@�@1����� ͙�T����c����܈ &
�`�RO�=�Ш�0`��@�Qޛ�݀_�@�Q >�φP	��
����ΡM-s��@޴ �L	���� 3���7!�PW '�R�wUy(z\C2�a�=��H7q����j1�S���샨�☂z���+��T�AÙ�9�t 5�s�U�Q�*�rD��Gɜ�U�/#�V���Ps$�	������[z��IgH9�U�F��iq%O�ʀ�����71F9�a�*�' R��30� E<j�'@*�7H�D�~�����3$R� ��woS W2��p|�k�Ӓ (��`IJ��#�ű@ ��<߹��Py��8�! ^aߥ�1#t�c� �!aD)����|�;��&�X�� �g�U�����Ѩ�`k��cs9 b����5�, �	�k Iap1�ܥ��|?�Dx��0�L ��d>�& ����2j/C�����D�~:�E��h�Y�{���y}�r�����8�Rx��"DQ���lNr�#��y�y�-
�!5���[7 �A�H�dG`���� c�\��l̐v`� 1�j,,�Cs�D�!�C�E��  �nc��)��P���օ>���� \f�:�� �(R� �r�xI������8�����r ��h)X�6����`�X"^�7�H9
#���"ل@$Sa� �� ��WYTDx%˦�S����
Q�L+at���B���V|��@��1 �;����ۮw�)p��g��������P�����	����!$
	�������`�!O��2J:%.H� j ˿�Ih���P���3��P�,�:[. ގ���PN ?�K�Ba����@�8��[ ⟒�3s�� F��Ya�&��P�I�p�鴐h�{Ij0	)��@���s[8����ێ�.��s˔$P^u� 7*��oqS�>	�p[����"��:0U k�z��t"�=v �,�jЅ⌂�����a��R� �9,���"�r�e�Xv�z��+'p������و�/��O$� e���g� 
��uo9 �af�n�/<}�r�x{�@�0kd�s�����@PγYVC�"(�M�[WG0O� J�h�� m���������a�2R�<�H�#CE`s@�$y3\�d |�ȔBF��
O�?�*���=�q��sY�ա B<�g&3m�F!��={�/� ���[xr �
v|��/{$+LS� �v���'?���,�=��� �. ǟ� ��ѐU�� =�1�5�� ��<��gA��K�3ҳ ��̡ R�]�w�HN��� 4�Q���,zV`.���=�ӅpC�q� R�Zf�S�����(J��6�� P�j��^H ɛ��ֳպ(,��Y��1|V�=AxQ�Ap� ���4���.N��6Md�| �`��һ� �Un�z� 
S���E�p� �^R�ա� �xB��{�C �����$�;�QM�5��2���I>� w�����	�iՃ��C�)� s����k?�� 샢��S�f�� �D��w ʁa>�7�h� dx�f�4��`�Ze&� yV�r�?G� ���ϕ��� �FY�C� �U!��^5h ħ/L��� {����r� �O�q7�� �,�j
�Yf<����9�0`@��(�;\���˳t +�^r�ao		7���2P ��;��݀ ��L7nߩ� T>-�R�� ����?� �װw�n�� �Dv�d� 7����&���@��f ) �6!�ya`Q��KJ��� m��T��� @�z�� �u`�^�� LT�����K ���g�wv� ����M� 6����@ ��`�=�W����o��� 7T6�x��?g����Oi� �6z$�����%E �Ǿj}	8� ��^� ��ۀ��J�$�{ ��V� C��P�E69�c����>����A�O�u��%8<�(z���<N} �����C�8 �6��>���JYe��*��䅮�@+l�;�� �a?E�@"��5��@B��'
��k�.�%W�V t��9� ��D���KrU C�:h��� �}��x�9D ��{l$�7����� ��+�I�����h�B u�!PnR�� C���dHZ.��䡀Хe.�7� hN`��:�Ov�Gc�n� ^�"���i�mN%�݁T��~�#g���2ڝp� [&�n;�B ����Y��p
��� hF�Qe�-�� ������S�G{ �yL��z צ��aY#" h�9�U:�� ���=�t I�/[Y��  h�Hl�&�;$���������m��h0�yn�[Dl����� �)&�cZ;�=�� RϹ�
4n�h򐻣0L��<��:*�#r� ������ A�Pߐ�U;c���4F���n�0� ������Y� ������� u��͕;�	q �1�7֡� ����M�t�;/>�;ĳUIb������ ��э�L�
��+�����to�����:��5��  \��$P�������҄��:��� g���� &t��Wh�; y{�謡 ȿB����%P��� 6-_�� �����?�� �g(5�A����=����僞�0� ��7�|
�RP0�5 ]o�U�����ۇҝ�h�/ �J{��} �OҩX�U9f���-؝���� �zT�SB� ("�K3?� �1���^�� ���k`i 9��������|� P^gA�'~� ~w&��+�;�`�i*<��	�4��� ��,�@L'm,��� �.��� W�jK�	�g �k�s�-� �a|��ܕ��fA%;�� �젖��� H� ��?��*�UP	� �(.���h �]�ܻ� � �ɍ��;��u��˹���p�:)�ܼ Qʭ.���|y� ���������ZB�h�}��T���8�e���H�R�^* �S�b�\C� 
T���;�������;���� ǂ8�L� U����Օ� �ז��t �q��� ��0�L��=|�q. ���DpfՋ�q �۝� ����g� �ׁ=�@W�qC ;1�͆�߇�� \��g�*�\m+�2<�������ټ����ے� 2���S �G��viL�,\_�V{ozD �	gO���mP��/ ���.���c>,� �_�RQ<@�q �j`g�)  ùv����H�}Pc. %n>�떃 ���P�N�<����É+ĀD>�!���ހV�b� �^�3q�<E ~��f�����۽�ѕ�
i�E;q62,p�H ��݇�>k����V%���[�`���`}P��i&�]� ��96y�,v�,��p�N�A������)Xe��ݑ�O;0�S%g�����s2$�_.�/`/m���SX`5�9�W/y��% 4u�� ��9�/�J�(��Q�B$�K��{��,���(�� �tߖ���VP"����o��P�?��=��;�p���$������.pjU�e�I`G��� V��'��^
�����%�u�wm�" �����ڍ��$s�*w_����k�� ��U� ��R໖�",lȔ 9T3�r5xm������<�܀�g20����6�����ވC�kH0@ ���1� ������^�8c@������� �Ɛ�uj ��r�迸�`� pNV��!�F �Ր��������S�t�E1b� 
�N��&p������7�үE֧�ˁd�صq@��z=���h4�S��)� ��}-p��] ��8O*��c:b�r$I�% `7ֿ?�p��<pO��������^��<�� O��=� �2�����0U�p/� �7�\OHo L���臸�H/Tb�\��Qղp�qz�� O51غ��#(�M�`� �x���0�5[�µY�,�� "?�\��0� ��YI)�nOӯ؂5��p��
�´�� �[Lb��2(p����Qc�?���!\�@˜�[�u� �lO��)�#?/��XL���t��v2��ه���� �b� o�}�Y� ��p�	� 7D����- b2q[A ����� {�|���H�+ �C[�#E�4 �Y�	f�}S�F&���z���yZ�%��@�f[ �����-@iūƱoe��l� \�ш�Z��,ˤK UY���g<%��۠��TbԮZ �3��� LS'i��= �W��N�� J+b�Z�YS�jڇ\��� �_&����K5BPZ$���i�����@���N�{�]�q�vZ.?s� X�,�\Po/~��t��Z��lb΋�^" �E�Zx��H1� �
R�_,�J���B�lϗD~/8�ʝ +����w�}� ��b�ZI� 'ԅ�ѩ=
|��i/]8j�� 3[*ʤ��}� Y����[ 5D����}�z^ ?H�R�b�;)Ȁ.Q�pP�qmc]���Zr�w�=|��{�YW,����E��� }�<�BI���Zl���ʐj�UX7��� x[a� �	z�}r��i��@Rm��Zz���e{E ��L�6��i �������H|3 �Nl��}���&�1pO��[!#�v��|Z�Ԧe�h 5�.za[��� o%���t3��ː|j<�T��`�)�R@�C��!� �����lZ�gI?�w�}h ,&c;��l/$@t� ]|��YO =�_o��: �ka�d�R%bzZ��������,��#}i��
{�o b�/ZA�&� 6�D�_L���� �-�%8A}�?oU��Y*�8��kĐGu� qi��ӼrZ �m%�}N[@ #1`���_� ixE��� Û��.MLdL �>_ �i�b�� zou��J�±@[*���̘C{ls���m�GY^�ۥX�a�[�R k��m�}L���XR�:C@9��[�]0���w�Lj� H��vE��-�b�gŀd�Y�:'���k�:@�����X� ��}�6C\� 4�$
�do��aD P�Z�2Icd� [V���{	� ,dvsc�/ ��S�Z����|L��C���;�&!bŞ����h�
^����ŀ/PBl`��\3�(��s�5�k�}�	�W�Y��3`' ���y{�]�7 �W��u1jn�E8(� ��}D�W~�<���>7K�#���08jf ��$��|-��lp� E� Īb��Z������l�S ���� '�}�ơf��Y|�r���m�9F�UV -q�Y��^���[}�sv(,�!�|0���1 �J��~��^e[f
�P��5j�T0�2�Z<o�$e��H7*��h�)��BL`ޓ� ��<wb��h	��� �D���l��� &�|��`[��Z���bjop�*��q�&�J� c[|�tDe�p���ӫl���`|�J �|I:�rt FD�N��Z�.�( �㙆����}0i[!�{�b��}�����VE̤��(�ZJ<�` &�䕃Ԛ��D�� L+Z�v}��<�� Ob�|j8ד�4�Aq-r�p���}���(��^��2�� ��F �EQ;&�: �oa���$4�`���|� 
�z/Q��pWTsC���U� N�}��1K�� �ku�_�cv���A��9o ����I82 C��X�h�0��@�V��S5�׸DB
 �"����� ��va��ic,=W���r� ��
d>qD ��Z'���=����@�F�0�p���߮��Hp&mfo��;��P��������;W A2c��*w�,�% ��&ax��m�Y�+iC���N	�넇c`1qV��R�n��6�� t�E�{�� Y:��D�| %}�?
���( �b�A�P��p �W� �1��p=����6m��C�q�� ���|+I��a�@Fz
V Q��p.�  �L��e�n4��/�E�v�;�AM�DH{ p~���a1� �E��;>gA:#@@Ċ�rZ� KC����>H �`
��,p^ Jh��LC�j�w��;> �� B+��R�xH�`a�	�?� ��pC(��yV v���;����F�@���r8�(�p>
��Qq{B� N���Hw� �֓PD
# ����[q �Ō�ZK3&�C��VTq_��	H(�,#������-3���DJ�A"�q C�	�co� >.F&�U!� �8� ����� AyC���� P;	�G$�@	+DV
�ZC@q?Ǳ�H��$g�J�RX �c��)�
�8"	5`؅pD ��e[��>ߍ��d�� �a�nK=�bk��l�0~��⤽D��@����b� ߹�C`e �F>����h�I��L�����b9�R]��> �3�A�p� n��
\�� �u�����`�p?5)�y�r�t���'} ɳǻ�� �z~�$C��8���H޼A��p��\����� ��h`D �.~�w�J
1� 4Q���ބ���+�n�t;��o!Œ
�ܦ>���e�s��04I��}�����Ϭl��
��t������4��b�M�.�t�q�S*9���Խ#D��+$ϲ���3���Xb,�M;iX��� ��a6�Y
��� ������Bs zH.|��( ڞO
�ś" ���L�f	�y	��L��2 kT����n��� �C����S	�B@`�4^
��V�v;�M8���^K��f�"l�����m��jp�X0R;��� ��`؁o #Ӊ�
/=>m��C0k�NB�HM���z(�Q`��`t�\\ �&P_X&Cp�$ q� s��.�������`��(s���A�8� ����T^.p�| ҷvqY�� �C���=� �Ė_0�"��L%��$��
I��\'�`8�(���N�p��� �P����A@�w�/S����Dn�Y
:JA-��ʁ���g���F���c��[ `p���ƭ�$�`��v3� �q���w
 [�i�B���C*N�G���}�� 
�!$�K� Yq존s��=��4��/� �!�ީ��ώW	�0���9S�(L� ���`}0�	Ū2������:�l+ ��rB��	�*p�>E�~ ����,�8��l��
%�(iZ
���&S, X�MF��J�Q�CC$�	����Z��@�t�L ;횤�H�� TC���~ ԇ
��"�X��.%��o���Vq̀�	NE
"]��@z�d��(��J�`x�c{�5s��\����z�X',�����K[�s.p�D  Q��lvj�2�m
���>�+�#I"�����@��3p �ga��I��.�	��$��$���G�;:_�b��e��*F �
T��H�D=D�P����c�p�}rn ����R.�&~d ����9�x� ��L	��x� �o0(qT��/��)��0KVe\�GPH#?q����3/��&k Ce��6�p��DpV���C
 ��waq�tPKg�A Hh� Dᅋ8���P.�7-J]§�a�@����r0("��k!���� ���L/Գ5�~�K&�\�E��l��ayM�`����zX-d F�0�B� D��+�� �)��d7�75�p��'�"?�ǂ�
CnB��LV�>c\d�]�N�,��o��L��>� �[a�/�d���$MC�cD��N��rÍ&w� ��5���Ƙ0��v��pk� ]��RUj�gC�ꂊ'b����0h�@q�t�}
�Bˮ�Y D1w���l[q��S� �o�x�t� ���{�IZC ����0�/� ]��%�9�eC����b�x4{��Z�#����Ktk/�,� ���z��r��v
ƣM��$Zt z�<������.� XU�
��&]� X�Pոxr�T �EM/�u��} �I	�� ���Ց
�� ��.�-!	�>qĀh"��%��k�����������&!Q� ����y b���Ct&[(��{F �幻��S-qg�8pl] ��C���� �*OpB\w ��6
Z�' �����kN\�h ��\C�x� a�{
2��Xb�D�`�0��P~T���l-�����NY2�D<�'zJ� �GC��Κ���
-;�A���w|��!C�9Ҹ IL�K9�����V���L�  �Cs��X��1_p�6�e� �ԛ�D# �x
'�C^� 	*{ �TH���c�|'bm;8���`,8u�� #�d�f�H�` �D��kA�^ �=�� Th�J�����b� ��3Ð�q 
�f���Qs,7�6�0��`T lp�� �T��,c ׭�M��8`���S ��U�qW$�tX	��R�v@t >�p�@h`�Nr� Ժ�A �L�ՌD� ꃀ	!�Hpc�Lł�2���r�؈&m	C`� @��.�Y������$ߺ��w����	(���.�q�jR���f�s ��Q��<�� ��dn�ED '|NC��J �w��4�К�DT�}8 ����޺�����'j�9� d_s�5��� f��p\ F �ߜ'���C ���s���v���WHiC�|� ��9�(?g��ЄL�B3�eձ[�������if�#�M�O�	$r��p���Q�I ���E5������J����� )x����g ��a�,�ָ'���8S��|T�:�/����D�>��� 6b�F�w|ə#����Zn	��=C@�6@�s�; *���Ջ�����%{�벓�#w� ��;�B����`��݁ �Z(!�>�f8�Y�e�?vJ@�y�c"��Mk���FwG050�� ?R�f7׏�D٬�2UTۀ@��b_`�]P��[�Z"_^�)9��a���W���uc����s�$^���Մ b1ү"� �ꪛZ[P�}�z� ��+fШ�)EhX�}���� Ǥ����ݖ X3UB�	� R"�T��ڎ�A��L���0 1���?V ����m���S '.G��R�D ���#v)�| ��ua��_���B͔J@hbЧp�`���<��q�8�(�f��� ip g2(Y�ޫk�x�P9H ���,�\�7yb ����p
� �����������b�H�?����I��T (��hm�3� �a���ɯ0
YA��֍�6��a�(·���[��@�X�A���RJ�=���_� �[�C�t��T�����i�`f#	�! ��ѹ�k�yn5a@�	i��Ň��0�w`��a�H4� �iݿH���&!� ����G��I��=S.{�P(��:�c3x��rL�7���!Ro U�HC�%7�5&|���!�(/g�e��h �_� ���䋕�U���ө��B|�0��j�ǈ+����@���
�W<^� f�[�� "����,���	w�d.�"�r>��t����X��亁J�fݧ�8� #�I�KA� dBiXى �q]���j}� -7��p#e 5�]��nl �=>�S7Lc ����?���/���,� ��i���+ �Q���H;�s �>J�j� nY"�6bt�����Cz  Nam�_}QGy�z�k�[�T�ˈ���"R �(����z ����y�Q��^�[9� |�m�0�u� Ug����ƴ?N|8 �F:�nD�� �f�e���]K�o� $��t��n� �ƿ�V��l����A�KC ��P����o�Zi�nNL�t�e��E��[�� 1F���D�� i6���� �<z�$c�V��n��[����{���Ĵ`A��(�L�l1�i{x��_>h$�D�Ga�!��� �?b���AQ��Hg�rb���C�*͌ =Ja	Ӗ�����`�΀�^���Gjn�� �84/T@�\l�x`� �mLR*T���0!\�p@O�G�A �c��(��?J��f]�g���1�H;J�X�!�Y�]�,�	A��U����s�M��w\!�d�Q �|⨘���P/#� ���/l:�^��?� ɠ����҉@��ؾ;�X�`�HC�Z[es1�(a:�D) ���0�T��a�X<-OAK��Jol?�Q��,�v]�8N�Jt�>�aa��L�� �� ��&����䫎���L>E�P�	@HQ�e< ���
����1��"X��H#�T�Ow� R���Dx�(&�W@%�[�tlLJb� ���>������Jނ�A0lb��f�XKD�# �����ϭ0}Z�I�qY��f�#� pK��?9 �J��e�W�A��=�&��AW`Q�N8���M-ilHd9b��P�� LQau� J;�ѡ�X5Sr U3Sg�\��F���/�5�=�T�C�4���j���θ7��2 W`���  ��ŋ��g:#� ����q]��.�F��H���!T#�����=��f8��%~ (q�� cA�O�V֏;	i�R0��I���Qw �!�{�-�b&fZ��8� �}.&��� ���>mZ��jN��i2a�YK|2��D,	��/ �J��ꨴ0�,Oj0^F.��U�pfm�� ��4�OZ��T�����Xi����:'(�r��(�mb��N���0�Ea ��D{|T��0*�g�hN<R�" f���|�d ��c��3a1 ��Z�*N	�9�� ؏'��(��}�j��"? =w)h�>%�O�l25ȷ  ��}�)� ��D���(��P�7 m�&�b�~v���}pS���:bzQM�I� $�����B�{9 t&����G �`�. y�s����׮J�@��XCg �!a���\`����~���nw�'���.���_�8 >q�׈�jD`R���;?�� �'$&�t �m��4�� �]ґIĝd���� Rr�Q���>�� Q
����l:J�@a��2� �B*gux{�/N��=��G��Z�XϊR�`C��-���
ͽ�N��SR���n��`������F�&�ȣ~���� Ω���
�<�✁X 倲VQ�v��
��O�j���wRC�� ��n_l��������=����Q)���`AS�9�s# Fj-�'�I�����{� Ag-$E�U��#H��Ftn^](��Ȝ5
�Dl� H�@��]>wL@��
�� ��U���&�i"�������V�T�HW]ˀ���6�I�]��~���0f���(",�e���������K�� �@E��҇'��7���1Bj:5! K��<�ŭj "}Q�v�`�O��.�5�20C���ʇ ��8-�0ȏH^:�I(oa[J�#��S K�W(�XJ�o26�,	PbiK�Lei�x"Тւ�����YP�4�`�M!>e��H�D@dJ�	(�o���BE�_CL�)V@�RP��,*j4�"��� �Z�����������E$HNR�� ��ۚ;/T]B� �E��lxbX��2=:8�����o *�b`�HC�c/ �`�>Qj��`+a�զ,�8ڰ J��0�Q�<�iKcgy�HsA�H�\hV"]���2A�ы���,P��#�	Ī��H	��I��\vJ [#~ǭ�^�0ᕫ��$�h	�Ou(��@�|0����*��s�<�/�;=�rA���	
q��!l1�]PA���q��8�O�n��o���Jp�������@��3��̓ �R:b3y!����2QۡS����W�	H�1��p
 ���PZ�W�@�8g���!�I`�b����l��(��C"�|�@�} V�WJ�������K��ۈΐ E���"��p �����
�@���I��6`��	V�^9H�]���A�ߵ$����R$p�b�P��"�N@�[�i�\������[�� ��	"� �����b!��h�x$$0P�$�),�Q��܀Lb(S`d:�|@�A
K�"��\iT@��C��K弈��bS( K�~ज𛫌^ XR��)ߐHE�3
���}���K4��Ϸ �7�T���� ~F��>E�0y��]��a�qL�8 �BoQu�W*4)�>Y@	V��RK�������g�@8ip��F�xT��$���币_H��SXh�
����x<�b/�H��C�;���`ԨU},��J�ݘ�:�^n ������ϡ��7AOEh	�w���E`# �@�����J�@d����~ 
 �xU�O ]ܛ�0� 8��W�[���x� P���ȊO�o]�B�a��w@�Q	�G-��� ����sn9���e6X'���`\��H:Oԗ����T�� Ka�1	S� ���]��n� �0o���=/ ���Q�� ƫaߢz^ +�qG֗ 1��~�� ��.L��:f�So/G嗐6a���8%��P!:w1 ��S�
'곃��6��� %�C����X���w {o�I���,������4�f�� �a`q��r �p^�v��b�4``��H�� CwU�jK��ǽ�O�@��^ ��ɼ	x$>|%���Wk��EdU|�|B �����S���h:� VoX�� lR����="��>kw����W�x�aȁ�#�@�� ���
�v� ��� ���t��2�^o۔A QYP��&�	��1o���4qp���p�,X�L^Б�?�ևNEf�X�O� �s̺h-x�"���B�4X�@ǽ���2��nQ�7 ̎���0�T�p���r �H�!.ûz ���~@ �3+�p�9��t �WF4.�Q �\�0D'����o<�t [#�pZ� ���B��`�!~��]��P��3 xSmF�4� �Yv�h��֡ݚn'v*�1� n��/����vU;��@��
���^:jo��ފHx� �&��#NU �T��� �p�ް�9� O��7� a�� ����h O�5��� (�k�<�� �q���`@�U���<4� �j�I��>��AZd�ae $��Y���q^���xp��D/o�&�fl� ��}�R� ��zw�� ��%��M!�o�e��#�E��\UO7߀��k8�x?��>M+-b�p�� �d�2C�m�wXW���L	С#g���.����>�U���F� :�R8���~# a��^�Y�!���ȓP�A��G��	�� ��� �1�2���w����6�B�\�`^U"�C��$���.D� z�����!�� -������z�?n��{; �l" A&|� eNWU�!�?�\�%A0�/�
ű�y���Y +��M��!�֙��/C3���~h�;jW�XUD����K{��<�q.�\ @������� �vg��$�:���&:�O�!逬���]����&p#�kO�6��`е{�� ��P�r���Z��h�`�W��&��p/� ��!�^�S����@و��.m�  ��2�:1��zWE}��$�y	��& Ȯ˂�	�_BHར�b�[��m-��Q��n�,��ܷ�l� !_��6� ��Ćދ��$�֤ ��G��yxB�����`�� ��p�m�Fyv\�D c�i?H]�w� ��<�3� P���lOs7@��`A�Ć�<���\- "�8��?X�� �G�pL��	A�j� 4���#L>�|]ŀ�Fի{� ���*?�|o�����fW��4/��y:o�@��\u(��p��7" �0�u���p�m ��!"V�6q�@ �J0wX�$����W#<GP�N�� vfjw �� �Y��x U��>ܯq�̲�|�=:`�ܐ�>^F�ػ)�(��O� ?�3�� ��a����SЦ�!��2�s/�|z�x� X�>���pYnr�,`�?c �p�!�O+�P�{��� ~V���Ɯ ��`%4Zi�� �G[EL���v �� ��!�����> Ej��1 ��(����x	`�za���!�L�[@��*�	<Vq ι<w!|9 �p�?�c�Ղ�j0L@
�{���o���p�� 8�A]�qu ��)���� 95�c$!� �3|����0�n?�Hs	�e[�,`@ŵ @e`��A�,��Z�e���2O� pa��k*��د!퉋���T<[�O�pѴ Ho	����{� ~'1�TT�(��C!8q �ᾬ�t�?��K㺠 ���6� � e���� ̒޾b�� >��_("��� ���l\9�� �kt�*P����e �9��y���lՠ�8 �� 4#I:(�� l�a�i
-�}���!lwPǱѵ���X:0��)f� �A��E� ��+�!p(�7 ��YY �\N��0 �	<��qQ��� D���"g�����ɺ=�S������=+E� ���bpf��[�q9�O�V�s� :6٧��� ~2��}!��*m{�Mܣ_r����c�,}|^K�ׯ줋 �<khm�� �5繝� �ؔ�r%~ ��=�md6� ն��{��\t@�7��Q 6I^]�rԬ��Z�ùd�`D; �N��b�w6 l�Ls�M0�X  ����fY/�Q�7>X�l�P�Գ uE����V @�}�[��;����ٻ^����m �Za<���� �#ĵ�L '@�s=�I taSKzdX���/� �~�s" ��g�ă8� m�ڭot� *�n� ܏[���h�L��j m����=��H&Mq%��0���t� 丧Z}�$s��r����� ~l
���*�Zm �>P�eh=�̀�`���� jÂ
�ti*:k8�S���ܺ�>qn ��H�� ߋl�!mO���z�:Ίd�ه�"b����Y) ?�Pf�w4y�v�֠8�	�T< �	��� �j���/� �h���� �$�\�J�C 	e䌗ք ӊ'�g���X?���E(@�tb�c��k�mQ[�x��Ws� �o ��-J�f�L���[mn��lq5�J�� �z�# �`;x�r{� ����gA�� zI���> ��~�Կ
 ��ܪ�] Ã=�xrQ>�,}o����u����b��� @�~��� ǯ�L�܀T��r{�3=��<sW]Ug���� i��Z�ۈ� �����c�	 �(�2�� �^Yn���}�+b��@��~q�4 DsB&p�����)`�W�y�`��_�B�s`}Z� �i=S�� �C׊��,W _t|z�lҏam<J����wr����7�ɹ�>H_��M��]`�ǲ����(�Ɛ�~��� ʛ�m?�� lHjD��z� �'u��Yt@ G眺�r]7 |s�n=�^�C�
j�	�u l��Z�FsE��@8DCc {�Ō75rA��@)8��iʽ��X�$+ ��o�k�pB>m� �l�`�{��At�������&��}�ЋÇ����=��w@�s� �Y�<5���Պ�^%�� BLÏ�m1P+s�0:��LGT lV��Sʊ�rigct7����R�X���ъ�3P��tʮ&�
m� ?�s�:c��~w�d��q ʍ̣XƿS �lZyd:	��Y� P�}��H^t<��-x�m2:O�� ݄��X1� ��Dl<Qs13����� �q�~�im	ɡ]��E��H����l �ys۰���W���6`��} �B�s������'m8y,�8l a��D��x% w�1䞔�	��W $�Cs ��p�}G�Ԋ�;�ݕ��	mZ�]8[ pܠxL� @�9�n�	�k:, P��me�V��a=�� �g#}�| \xL$m�Bt������H�}�x@��T^ VG|�r��0 9<I}!M���;��܇K𮸆 n���r*r� �fdL}�t� ɉ��H�xEs ��l,��� m�PnY�&��c��-Ȗ�
���l"��Ŕ�7�×���v�|�F���l�Æ��ˡ�<�0р��� 氺�$#�'l�|D��LeÀ��� ����jC� )�m���� @*�Zڈ󣘜Ӑ.<`�0h��mtW	��0���q<����~�8� �lʌ�sx �D��a�k�Y3 L�l�& m�w�fW�O�� ��l�A3NnH�H� b80=�G1 o��I�l��� �EOc����&�҄��&_��� �f�+!mg���	̼L�r бt�:�-�� �,mf����\&��h ��}�C�|�,��|z�:s7���� � �̋ɛ~e���M��d�u�k��TC���tp��N���m�jk� �ۥf \�~A��Ż��y�xb��o���0 ����[R�$�N�+���n`��M}� ��l/��j�{�6��~;����: xIt�8�a, SWm�r��t�잜��� ����u�NO�# m�`�%����� !�}Ҫl �$m���X�, 3�����ʮ�I����#;!�}{s��dq�����}KH�� ��Aц>;-�|��t!x�7�}�"@�.��<;��� �m�R�� �a��E�\�� ��Zޓ���l�]�;�s_&p�]̀XmU�8%� ��(������sIn�@}�&@���+L� �b:���g����sf��[ Ca�,c�b!}�CY=��'N|��w �q��HH�� ���*�0 m/N<�}�n�]�~�@[�}�&X�I��`ԩ @_�~]���F�^����(/������"m�p,< �����@�8H�� ��O�M&�� p��l�k]rz��,Z6� �~�Th�	��z ��D�l� �Nu����j=�JШ�t ����Rئ vs�V�X��K)� ��. r��$5{�zs��E�!��wf�Y� 4�n�% ��_���� le��)��?ʨ �~�CeKu �����" .m��s��&�4G�'p�b����ɐl���r�N�6yf�P}�$!Ṗ)U�h���4�)��k�H����)�����<I��Eg�@P�C��L��1�}Dazq������c
�.@8�X "��@�}�~�����x�F�,o,�5������Ks�~��ב@����	I��c�`�F�0�x0�a 쎾���ܖ�\kl0`7 9�E� }w����.����X����luJ �!z� � �͋|��`sO�9�� @t�:Q�� �csu�h�~���P�$�X� ����Q"��~K�0P�S4v��z�D|@���� &N�~}Z�1�;��ݷ{�&�M�I�,OT�2x(�����[�L�>\t:���@݊��1q }������¦����Ԩ=�p���`��0L�����̇�m��,�& �}�0���<�) Yկ߼�X��~ l�����u���D��z��Dq�������p`V�t���}ow�a��_�H�Qs���@�O� D�o���$�Pl�vF�1�
@�P�ml��$��=��B_�XL����&n�N�����6 ��ݸ�q�~���}�`|A�(o�#u���tn=�[ �}�z=� �EYH
�Z �b�^t��	�*=J�Ї\ ( w9[��L�ctՂ�l��	��7ÀXGj�� �x%*��b< n��lg �0H���.Y�"��m�, ���>\t~8���� hѤ����T��( ��q}�V�~��0�u4�ʮ�|&J0ۃp�R� �:��}\��_L� [�-� �Q���rxx> Gn��f�}�E`�z+���aD�pЊ dR|�oB��'3Y��u�X��R2�8@Ss �	6Eü,.�=` �}�['JH)��
��Enm W���~@*��^� ��X0��e_:I\9�&�H�FS�R� 4��4?`�:z� �]m�dUu� �}
yw����k�@�[;:ʸ sZ]���x��ي� �&��4�Sxn1�@�mL}�o|���	�k� F��s�����v3L�OB a��`��o #&�l��9��� �Y�� �~��؇X��0�y�l.�m�{�g�� iI�}�� Ats�&J�ٰ� ;�o1Vf�XH� n�}��B��`��k�ഞ�.�p� A�Ż� ��x����| ��)s�5����w��G��h���?# M�ٌg�l: �5=��DŇ`P�} ��~0������;�l�)� ��c"�L�:=�G ��b,����}�qi�H��� њrO����oW ��M�f1�~w }�\�5D��gs�K�	l�[F \�`�u ����}��9��:�c�� ��:* b�f�Z���|�| Hd�7>ʑ:	tE� ���� �W��~�r� }���y5tS��:�^����k�0 �w�-� ���h$, r�f��l� ��mD��\�~&��<ŝ ��i1	� ��l5+y�� FC[� �� }�dK����M��ۉ x�	QS�7���YH��>�ML��9t��Xm ,��|V<��	w�� lO���� ڪ��[m �x�w/g�,�~C&	�I�N� ?��"	�s�o�煄c����Kp�t�L��O��� `�lu�b��.��V�jv�����l(���0�� P:�Y�x}HC�\���8�� �50m�9� ���AM�6H_� ����*�L�0~�s@c��}���F�"�uz��7Z&`���,h�ď�a��h�ހgP��I	�`4x�P��M�~\`���kT�ͩ�%/��4����\� [�M< ��m'LkJ��-"�Ht�(�D�0����x�:y[��ʑ�,@�靨�0M�[ma�8� Է{�:�z<�r8� p��
�Ȇ/� ��1N0�YP	�8���2 �D��/�l�9�j}������<m�۩�,�� �_bq�l�� �a9I���"��o�a>t|�;�&��0��)�X����(���V��
oE� [t��U�څX�d"�Pi���Ó�(� �c�S}�� �ؼu���8��?5�*]���li�oc'�*^��S��
qm=��H�u>Z�݀��E�<Jq @�f$�� E�~ �ԯ"��'}:���8��`�yLs��9�w�`h�
�:�����t��vԉ��x Z���>4czÂ�"�E@(p~���r' l���s�rm}î���M d��N��� c��H.I��y@�zǋ�7 ,�Js���ח�p���� qQ��}K&�10p����.� ���6� ]��?�b��H(� 1Ӊ��9_m��r��D��PE'9d����v �r��Pl�ws08�:�6��X (Ŀ���2W��P�
t���֌��j���e���=����p5(�6�Lƣ �g}�
� �l��Mۜx�,�,�>�?3�L}�g�,�>���$�� x2mx#�����M��۲��� ��̩am�^]t~���u�W$� �>��h�c�_鑴0qr	.$���68�}��,�Y�" mͨ�s�=Q�܄y�)`,_I<�4:m *���Կ,�a��U�o�l���xN|s�K�d�@	�}�F����+"/msE&I�b�a�zR�@R�!1�h��P�*��9
m�f ���O� HVj��97� ����ع�� ?tL��lv�	�M_`!�� �~!Zh�c`Y|8Qb���LN� �G�����}���4`�E��cm̻4U�A�w �F~��%���s���( ��l.O�y|;�W���@���I �k5pGq��X���#���>� , Qx!�c k�NZ�� 0~�z��׿:hр]��En8��}uv!@�ޕ,��\0X�х `�	&l�;� ��BID �E���o�>��"h������İ���(�ֽ����� ?fg��`!.1 o��YW��k ���~��qv� J���z���py,���< �sg��^����8�w�N ����� ��=:��� �a��w���$�x� 	��]RJ�@-�˻��H�
t��TA�zĸ�psqf�@��Z�������l1]�h�}_��% ���n�W!6�z����p���9 ��'�{/ F	5U���:� ���j�P��<�+\���<����@� ؐs��O�����\�ԫ�TD�Y�� L���̜AU ���( ��kn��9����z���Iu :�;�� S>a8�����[����L�� x�6m���� ���{�g�<�K���XԌ'�h Jjhb�W#*�O)�����5T?�4!���� �_*��}�4׾0���!�<���M��ß{��ì�@�piWJ!�8�.C: ��=��v�O��ʷ���
/�������Cw��a�R-� ���ؽ�?m(Tp�)���|�طvnY>ל���uD��} ���j���,]#��v��?��(Ӝ�c �R��V��(����1.����_�t�z!Ө��8�%�xޅ}�Y ��' TK՘ �?����F�����\�@��� ���Ν���_�z �,׃X��� (@ h-����@>�D��a�]���&�t	�_/�������� t�תJ8q�M_�	���N F�wJ�bu����5�Y ϔw�� X�36't�
��fF� ��y�����cʒ`-� Y�N��m$z� I'W�E�, �d�v� *g�Z�
����z8�9� ]q�IY�S 3/M�Q�d���7հq��fX ���n%ܷ� @�\�<�� I��ɀ� �eSr�� q뽋nJ��9�����C�Ь�̼ hu��)B��R��@�.��| i/ٮv�w� ��UT�~Vtƃѹ����Q 3�B顀�P�H���ܣD&�}�R���=�p dp3�K'#�Z�+bϐH��� l;��?/<�2�zA`5���HD���O���k���X3$7��pw���d��(���:� ye|8������ώ +�n���Z�!�[�� �6>�� =/r�A�u�m��v��}yz �W�x�G��1v.�n@�s��� �:�M��� ��`lW���*�����pU� ��2��P�[5�Yy� �Q��3���(�?�O*� N8�A> ���߹p�$�����bHY��مP��K����@�(T X����< �`!� �^m��$�0��0�ּ>�� �dEI�y �T��U$��:=���ἷ�t�͵x� zL/N�%6�P�9*If�Ӱ��) �_�n�H 7���2?��W����%��t����	2 ��* � ڲ����i ��b�2�U
�e�W��������}���0��H��=�M3��] ����9����������8Yc �K�.�H�Pߨ��d��܀�9����� �4�U�J� Säa���}��ߩ���S�P��0"��i8��� ����0�<G�� ��u�����I�U P�a�� ��퍹@ɽ�(� �A?�0��u� ���m�.�˅�bp�>ɳ��?��@�E� �p�Ն�e� o��
�ǯZ8J�xP3�� �ډ��v�C �1������ ���/9�L���1���=�  *7�w�����Հ0& S���.mo ��~�?�� S��R��vb�u(�2j>��=z��w~kn��q���y1�:�e� |�S�%{}�� ��Y�F��� �V��L��"wS	��,x����~+ کyP��� �TR��W���	�ܮ�����i�#�Õ�M^?� ���2�bŌ�Ā_}D�tS �`#[�k� ��R���Y �\)<�} _��~��1b w�xU]�M� �����4iG 3d�{��j}=�q����A�N- ~�מ��M�q�iU}���ح �[ƽM����C 2��4�
�ؘ�  Ă~�P(� ��mw�R$t�����!��L3��8}�r��K$`R�t��L_{G�.�C���}���<,Q�o0���F)�Sم!1ۀ�s }0�x�aL<��t	�����g=S�8 ��|q7r}� �jI��)$	QW &�T�M ��g&a�O }����NR]�Mc��Gx� UZi q�7� �@}�#�� �l�G��-�Hq�� �/5�� �~�R�r� ��M�����8V3���� =��%~p� �� ��6�,:�� �$v���}{\��Qa�~�=1��c�-ʒ(�� C�M@�2	�8��88�O
6�/�L9CK����}h� ��s�� Sz����� �V��*֝x�d����B	��K���L�� �x�i�$� M�2G}6 C_b���L=� 4��S��p/`�����y�� $B��@����L�� 4Vs+~$��D� ��� ��(�
M�v�iNf]N}�K��o� ��S���"��@��T}�� �~��{��� �	]�^�?� �Qˠ�Z(V}ۢA�t����v-K�@]dAnB���6)P }��&eދ>���0� 98�5�$� �}�p�~2&����s���M[x� ��!o:UH~��3@i�	� ��\�Xε�=.� ���MFP���t��>�8� �;Z	��>� M��5q����~��0��_���5	L� x�\#�9e �~�P�}�8$�7L�0 �ܰ!�$UA(Q�cB�T`Ś� 2⪟�0��3��/��}��P.���  �"le���� �j�߾����{IL��40Kr) <�
�.+ �Log-�Dĕ~�R��@ܓ� ��P��i�c�M�R}� ��ny��C� �Lӏ�5w\$9d\���~��`�;�pA�� �ɢŤ�?}���P�0# {�5�QX��P���4�i�	x�}2��~��p�� �
��m���	F��ɀ��@���~� �H�����	��� |���$,Fd��쀔C�{�<~�=�&�PEQ�� �<6��}S��} ���閟�X34 �T�e}�t� ��H/�k�	��M( ����� �	QݭW�k �~����v$�2h �x�,�	֮� P�;��b}���
��� .�r��I���S笩 ��� ��(z��p�9*� %Y��}��P$������;D3�0�à���;&�>��@���\\��d-)���%�� �~���t�<y2 ���n�ES�@�ق� �}�"h� �*~��zKg�ǒ��c��,��@�'yT�}���h�ŭL^� ԗfS������ �M��
K�$�u8�6���� 5\;�".48S �ɓ�`,9�L,^R� q��Mv�� W��z��t�� ���~�$�/8Q@Ay�f��d��/�`��* ^��8�o�ؠ1_����C�@��}���'℔�{$BzT �q
k�{�� l� �~��}uLq�#)ɗ �,Ξ��� O}ѽ�~�ɕ6fK �C��`8�ˤ=k �S�P��a\.}׃ܞ�KS`�8,����X� ����}�t=�~ F�AU�5� ��@�� ���}��g�p �!=���J-:���A�5m}��� K��~d�Y y�����zL} �mP�/��	J���ث��|��vU�� �C��N�D\'x�藀��SAY �R�G��U񝍗�]}��`���a1����ʋp<�:� ��tr09�t �e+	��N^�Ix9AG���m�&�5�-�wA����I,�Q�	"���8>��$[�@���~Œ��$Ǭ�H�� ߠFi��R����X�M 8�`���C�W�L��8�s � D�`�e� �%~��r�� Rl��]� �.%=�6-�uL�а���8ᐝ?� �E�	/mƀ�{�' ��N}�?ڀ�|�����@�"�B~C���|EcL��� �6R˦0�Ԁ�Y�$
O4���Q}�; � �Aj�.{h�B��q��}	#� ��ͅP S^��ں����tG�xg~/ 6~���\�L=�9S;`�Z ў���5�� ��~�<@ �R���MްH�xq"��XX PF}�~�e�D.>�L��d��S-�lbW/� ,��Tz �f��'�0ܠ���XRPL������� d�$M[4���4�8V���@~�/F16`�����b09p J~� ׽Q��	$:S(p�~0���t���3�|��/�����x` �t�	'��Á�T�}�9��H�?b#�Βp��
N�+�T�ή> 41	7#�� Po�"�)����]��@>�~���O��\�H``���`���,�,���#���ߧ>��.�dS�I�����h�@#���&�	��C �r��6Y��tL �A[{������:�����k}~��������P����`��Ȩ�@����T���A��z���
�D���� G}��Q� ]R��I��� ��NogS� ��|z�X}�m<�Ţ��E�0��	�4�?������y���3� �;�1q�넃Ӊk�؅�/$�ē��A�%p�����G����M0X�:}� ����\r���Ø�6�B�!�Յp(:�q �xd�$k�>��L#�wC�8  ֑��� }��!{��|�*���� 9�n� �R�FT�m�=~���$kf��QDp� ����e.��E~��NZWA#�K ���*����V ������^��"m�y� �%ٸ��t K��}�_(�����6 �Q�/Mi� D�Wr�},�� ���?��/ O��~���u T�!�ID�P� �C9JHFm��M��,�Y_�a����}��+~ʩc��p'�Nl �����S� O9�p/�"~z� �{=�n<$tEH0~�Sz�P��V9���# ��{8�"�� Ҡ�.qilS��~��`X�j ����_�M�m�:Q��$�۹��~�Hx��'8R4 ���M�6����!ay"#}?��=��s>�9n���ۘ}�� �$S2 ���JL�Nc ��ʏ��~2XW��M��D ����t{,��@�zyk ��a2s����ϸG$����	p��3 ���5Ϻ�&����"��[�Sq��h�N�� ą��蠶�|y ��I���$e*O04ˠ��K�B����3 ���ʕk+�a���rh�ӯ .b4*�� K&�u�c$��(e��=� �X��#�*<�� �ל�� SG��)���/"ԒԞP ���B�
 �4O���(��PH�g�@q�t< �1�N�R, �arA�h�� �s�}��m���� �S�� 
�����^ ����W�3�p�`����n]�^B:�	�9 m��7�>t�W�������|X�����ಝ�4@ a����& *m�c+8� ��6]��ɘ�W{�ӊp��@3�� ������O�I�@rm� ר���0�� T���=�4��Nb�����	 ����4�K\�z �˔�7aI��`lc@���n ���V�0�� ����m-�`�� ���W��� 2�%9�Fr�d�7�ft�:��|^������ �&紲 4�%LO�� ���p��c� K�����n�Cde�������VU�5�:�|��Ǐ"8q�N� �����o��ޏR���<���  OS�_UL�#��(� 3V�2�q+�9W�t ����^��x�@�2M�� ���tP��آ@]1f��d���Ap��8|�k'B� ��iA� (!��	��&� ���H�h$�f� �+5�"q #��I��c @��8�VJ��ᕚ ~�����=:]��s����a l��b����-���@z�` �H��?��z����f$m=��U��4�&��"$������V˖�P��r�⦙��.��� [g�*c �x�z2e�U6��� ���<F5䀤4R�LZ`.��
]#���5_?��ُ2&q�7����~��5=y����L�<`���X�E��ә�IB耿q�٢�vؠ�� t��݋s��X@@��x�	O��(4��� �;�+��Y���R��8P�� ���6<P���d=�*���ת���C��L��M0�r��E �Ժ���[��:��π�D�d���]��>3�"S05��u%��j��@�.��蕞��D��@�e/��X�4� �����4�	�-�����m�	��� ����� )zF��y`��+ŗ�~�)��'� *��<�C�\`��� ���Xm�?|� ��B�Ǣ}Y�i�=�/�k�2#`J�� �3��~�j�Gs�A� `P*:/�]µ�#�&b��e;���1� �M����� 0;�q�Gm;"���d�#�Y��/�k	X�7� D�^�D	[j� ��qX_��H��O%^.��~� ����� �O��^4��Ϗ`"i�]_�є��1#p�fU%�i���_Ӫ4�t.����<�5�q�	L��0l@eD8%c\�,�� �q~�PZ�!|@��F$zP DY��� �O�J/��F�L� �����VP;[�Mtߔ��* �ѠC�ho�t�F�`�_[�S���f,}��k
�4�\�N_��6Ҵ ����iV�|@HS󠗵���p�����qc�Ё[� 﫣��F� ���Ţ3� �Bh������ۀ�w�m׊4�|Y`$���85a�6��G��T����r������и��"�Z�%W:�H�6,��|������! r������ ��1��{!�.e�@�A��N lw���;B#HÜY�}A.!�( �ꗫ�&< ��rJ���U �!k����Hi� w�����h���!�0 A_)#]��������+m�ݟpʧ<��$�`SV� ̹d�L�E �X���Rs��H�O&0h| j�#R9�c৐��. ���>�45�!� ق�� 4_��๢�� ��k��+�(�7��H����f��������;?�Y���|XԌ��X`,5w z�ˤ����pMB���8ऀ�g�[ �8Sh�+�Q�{�%كA� ��b����t]�58X�&U��`L����;���S�	�B� hds��;��UpD�:������L~� >�� 4���QI=xW���T������,&�2&0ey� �b�6������N`	k����@�8e���E����0�� �FS��#�X=��N�w���[	��ނ��$�;��3E4�f��`!WM��-A%6�?� ��c�yO ��;��w Ⱦ&V�Y�9� ��60�Q�{r1�`�Қ>��U��f Ԣ�j���15�����Uɝ Z҄!�L�� ����[�3%� e��o#F ���@�28�p�
����{�$�r����e�@�MtI ��7l4!0s�.��� O�M/���U� u��,�V h�3�	�PO�8`�U�QSLc0 �碋��p����\IY��:V�H����ԟ�x� �ݤ��S��;V��w��@%��ԯ?� c��괥�|�肒Y�8
W�����8���~�`�L/���@����]� ��?��ǎ"XQ�C������&��0
������oH�A���`�� �cdO�C� [���a�06����οG��xq�� W%�*��G/��~���� ����1��G ���M������@�*������x~�6����ȯZv[�@n���x��.�s�I���O��)8@�h�X�r �K~�`�.')�|��f �� X�bi���� 	&y���!�X{qr��]	����:����"��dp��� ����'��- .��h����3iY����z����PJ��x�@�L;tЕm1�W�.&ӱ�����C ����#�r �\1��`x����y�����֜�Xڀ�q�N�����q�	��V� ]��������_ 3�P�v�} ���ӱ�ZBV۶W��:Ѕ; ��fiLc]�08b��O� �d������� 	�������.gp����~�4 �wnz��� �'��^��kgX��Z�} iӔ����L�*� �o�0��
�sӘ�d���
���(�-�!�Gt�B�P��ޅ��D?��Q�D��;����Am�˪��DEa^�(��S��7�<D�8񑑃�c��|	@�=9!�b����&��3+d�o7ڤ݀�H�ˆ���W"�wD�t��w�M
}v����,��%s���o����L�,P�v�-�W�m�����o�� ��sc�����ޚ�	 �1��p���� ��?�@ G<��J�{�5�	t]����#bD�V q`R�z ��k��7S�� 1�Z�m)�Y3UD�5�qBt�� /^<���W JNL�
�&��S���(��� ��� =>P������{/���F�#�,��aʺCF��ZY �A��ߠ����` ��l��F��ГcgV��yRrE�$��[ �W��Ć� ]��h�B&��x�����i ̌]� ���� c�2�N�g�w[H���1w�!����� 0�
D��}�ts��[ v*W��s�t2� ��ǧ~Z��^����
�4qM��3ž*�0�;�p���{��侭����XlQ�^R��{t�x� n�:]kߦx�L�ۋq��h� H�1V��>� ��_�I�.W�| Y�:����z� o���,���� E6�P� ��9O��y� 8����Ȅ�%PK��뜗����:�� ��b��m� �P*|�?����~���/���|a y	�?�X� [�
�|6`��! �o��᤾.��󉶰5�'�
�M����r� �����p|� �����FMt�s�� ȾN� ��\�0r�z[ ��H���� ����N�B���t���KS� ���Z)x�:~����dɧ��
���bp����ڀ�	۽��%y��d���XA� ���Sw������hQ �(�����@���~ ��0���B �\���=z� ˝�	w(���m��]�^0Ͱ�M�����(�+΀�6���8 pV 12�ƍ|\��.G� ��f�(~���Z��b�{���%磀zW n]f�[� ����9E�� ���Ź$�9F� 58�
Wi~[|�����=�p B��g�#X���\OI����J�0�p��
�;�Ā�?b����j��@��6�W�.�ٰc��\�������([V� �
���܎9�������	G���:� ^���Z�r�$�~$p ��SnVgD�{�[�b�Yp�dD�p@� ���\�r�4 e�ѻmL���@�4~��������t�"��4�@�X̾�s�9��:�<ǉ� ��MY����"�=0~�5�2���H�r���Nh�-⬯V�J��E���WT{�~��`j�7��l���]ЯO:�� C¾xduI�]�0 8���^��� ����ү����)@��n�H� ���>@��xy���ׁ�N��؆B!�`�����О&�p@�`� ��t[����o��T�^p*`������<���Iv�p�2�����l�oEJ���k+]� ��&}�1�:��*@ù��tX 2�/��o` &Ѐ� �?uN \^�Y��) (�,���f>'5:� ��`���2>yR�ֶ��m��#�@`���^+��:=>�zz@�_:� �4\x5i� �ȸaq�9$`L�@�M�(ņ�G�P�W>�a�j�-m �}��`.��:���H �uA�S*j �	�iǃ�� ��UC(!E����/ט�j�&�\O 
��D �V]8��,6$� dK�D� شi�j��� �@�?��� ��kj& � �՝�i�7�h�s̠�+�����=���
ԫ� e\pj����� ��8Z��c������]�o�	�~j���өܠ0�����݂�W��u�`?i�X�cp���j��,��h����bR� �o�i�e�Xgy.��泠�O/&�f��bД��i� g~�ިʠ �̏��H�馉�c��Bj���i_�F�Rl ��H�(�� �nU3�i��f�^��!�����(�G�,�X�i����[Հ��D�z��eo ��ad��� fn�Fj�e�8�)�a���n�8�K�3��Hj�A�����0T���Q�����|��e:����!lj�%E�`����I}��,;V��(�$���j� ��꤬4Sq$�xq3�a� � j]��iU�N ����,��ͪ�j��d�DԢ�����\
K�i3�������Qj�B�m�"?z>nM�\���c��������j��M10�%���)S�@�sZ����T/���Ȓ�� �`M���BӪ�tb� ���*�#� ҇�.�Y0q%p̪�	�CT����� ��i��E� ktL������(8��[J���
�c�!� ?<��� ���-~@?�ؠj�@5^�Y� �mF�R_0od�)���r j����l�p( PO{��� ���9lz�/&Բ��?x�Ǡ>��N)=���2��i��[,��;�0�f��>��<�}�b�����,@�߼�c�
zEv� �����T C�i��Gj��'"�(D@ļf��>�ek�<9@�l�d��u�f0�/p�E����$������i�
�`HڑC����p���?=fG�&5ԭ8��� ip7}ˈ�v5k��+Ɂ���0g��:j�մW`(�By �����uG:�4Է���� �|Jc ������d�R��Oxj�� =��a��&ڦTz�T7Cl���<�I �5M� ��g�0ʪ���e�n�#�9 ���uY�ڝH@lѪ �`�8�Ӿ4���H��Y�\⸑�|��I	x�g �%�>��T �n�r�mE�L+>xt �߽�c32X]$���@g�ؒ
:�}&�L�)b��|��mx;$�����	�L��D�`0�HIUi��ѨjˢP`��8���J��Lb��� /�C|��� ��cd�Uq���� �ɭ{?	�oLj4��8z�@�N~��D2dC C�%�~ե���$�< �{�J��� 
�4� ���H�rg�u��� ��N�b j�����i�)�����GC�X��s ��vYj�T��� P��p�� Rժ� P�b��e�\�Y ��'��� �O�7�W���5jN@9�Ճ�i�X�����j*��} ��6��?i��Y�\�����`�	b�!� �� 5�vj����K� ׇ�E�X�j|� �$�p��b�`	��g�.O�V����@h��`Ÿ<te��i�Uup�|l� �J� ӎ�g����uj���p��? &ԗ�q��*�� ����ȃm$J&H�h�'��ʩAĐ��g|�9������s&�� ��H	�4�Rz`��� 2���Xխ|7\H_� ���� ���~&6h�@`��i ���d�`c�C	���"��P��k	 �_�0�2�cr�%�Q������`���,�? VL�i䩍A���.��h��`O��U� pc��~x j�2\�[�8l�
aި�T�Y�CI�� ��i��t�ܦ��`�����CjvJ4���i ©�7���m��lt�h��� ��j�w�g�X��E@|���� ���O
!`�Hv���V�D�~�A����Ǩ�=��)Ì0��y}^Y�HP`$0��Q���<U�K�_l� էS/]��
�r�*�}�.�!� ���d |��˅��cnp�r��'���P��iҀ�d��../X<L���}��p(Iqӳ��~�5�,%R�̘�$�#l��W�`�i� ��l�4>"�Xe�����q ��B�Q�'�Ni�: fP�E.�v
 �N�Md������lք�10��H��ɴ�>�d����i��ć���nBv0���/^J\�����֢ �i�wO߈�u�A�_��0	P,���p�'tY @�;�F7g d����ا{�	�S�6 ���4�L{L>X��x�����H`HaqL^�i�<�Ԓx@� ��_����c�d�f��ɠ��x��&b���(,��,�]��l9/���p<��$!��Kt� �<02`8�ps�&,j �4]Rxn�^�.(��*�B�aѧ��V}��0��%�i��3�R����@���� )U��/q�(@H: �f��W�$�� Ȇ2o�f�[��aa��OqmU��x@�o �ڬ� Dj��K ���L�A���B�D�� /�͵�k.|T��\,
��=�r�ʪI����E� Se�*j�� ||l;��<���~��0a����tܠ��gӇm��V��v	�({�pJ $��ŉ) h���/� �M	z�Z���� ��W�Ԭɔ ��'Ð��� ��)!���	��j�l +�0�
ת����5�8��� �M��,Cs$���� f��7;X� �j���W��t�2HT�I |��hj�4���I`��	�e۳�����f�s`�G��i �e�|�2	0����ƨ�M�� h�P����cl�CWJ��k�p|���?4��!C԰�~��l�"؆!@��x)�Dpv�\�h��+�����.����&��ڊ#P�E�N�ʖ ޙ��j$�����R�����a�!j���d�m�i����L�ô�)~v���F�<5�Aj@��I��T3�%u ��Ԉ���I��`H.�d��ȀHs�8�u�!��9�jv� �����&�@��
�@�Y� �J��ӸXz, .�c���H��y����}a1 �-�G|[&j�,|e��Ѭ���8:���q��Pj�zp�� 	X,�ĄO��6���z�Y~-H�' 1��i�?� �p��l� _s��47+ @\�.d2|� i���-��P��xX �� LtRj��ӶL8�����>!&e�� �W�0z?d���� kӨT�/�H����U��Q�j��Â�a�`�%b��������xP�8	qZj��3�����8����U��v|��Ʉ���
�?�Ek�ÏC`h��!.�N�?��΃�
���d�C��{���� 9� ֬N���i��,@<�� �4��/�@� �i�z3� ��e��O����]*�DY�.R| ���@?йX0zP��6v��d��Z��ذ0L�5>8�6����@���b ��#�%j!��0`ӐW�	U���\l��b V��}��쀨���d� @._��s�� ���vȣ�P�r�i�]�����Ut�-�w@��#=*DY�,H	�Α���Bs���� ������̄�d|��i�u�A8dB��@�c�T������f���P�M���ƋB ���. n�&�a��G��W���*�@�\И �Iz��xp i�rj��g��SJM�� �����?�w��i������~%ԵP0p`h�e��j�Ɓ�H?`��\1:�� ��@��_� \�����T'j�z �!���l�ܤ� ���!��@�\��9be��Z�+T�����t`�:�� 䵃�~|֌L6؏�l �^n$ء� @%�t�2�]���f����Xt 7��i��U��d1,	�L��v���Z�u����Th�;<B�7(� ���	P_�lX�[�c���~`@�� �3�V!Dd\�$&�� �M'{��LlHp <�����5��ή:ZpA`0h�f!I����Y����ũba�TW´)`�� U�!�o�,�% ��f}��k���L��Qdh����8�� ��Ϻ&M�eU8\A�� ��0���D㪞�#2p�� Zɀ�i� ���ӛ��/�#��I��k�����) <��-Z����n�Lڼ ���uv �.�P�i��] "3����z��[�CT�jJp�T ��Ҫ�	�# E���i�|�D맑.���L�ت���d"�L �2��E�e#3X�0�Q*��`^#�t�3�f�y�����_��q�(pd� i�����}�wmb����1�8���h�=���?X�.l���gr�@T�q �Z-D3Hj�\���Y�T���U�����rCH3L.��������=�����d&; ~�A�����Fpl�	�H�sl �XM� �@!���,������d���pEi��s �q�c`�ԃE��9`L��4� �(R�<��%�����B3`|��r�7V��Sֆ���� �ZTݩ2'5�P1j�`v؂���>�}$�2�>�`�B�s���?�f��W:��aҸ�\ 2}j\q�i�.�	ue���Y�<��i�;R�r|G�8	ʺDo �L>�9s���},�IЬ ܏X�,��2�ഢ6 j�`�z�W��2�Ƙ�H�Gx���� ����t�>`�t	7��V�3u��1:n� F
?���VAvԂে@R��al��Ȩ �i��:���e�A?j�� nt��`![&,{�'A|;�C1�j�K�i�P�f\�R��6���Qu���@�T �i�	U���o� &�,�T2���� ,h���+�Вu �t��ͪ��Y�o3hj�P��y� �f�-�=X�&Ɣ�?�1�t*�p�����5 zv���S� ��̪�����%�
|�;Џ�tdCv�IpD���zT�� *���o�i���x�q�-`���� ���v����a�ٳ@짗.#���)4�p�\�  ?� ��Uj�'7~o�5�K4��(���Lr�@d�)�t�x
ΰdH��H-A�0=ԜZ ̚{��s>���C �<jfN �� n�i�Jk7�}��t���@�b���a�' ��ɩ�i�%�X��u�_0XE��6z����)J	�T�l g�"j.�:a����(4�aJ��� ��$g��'d����h9S ����C���i ��se����|�l���U�䭟 ��i��? ��I�_�L���S��v���o�i�
�u4� VC�x�R�A<hd`r��|�[�we�y���QD����	�Q�-�n ,=�t��q����P��uY�/Z����G��H��3 �u�X�� �9��<J�Pp� d6x����PH�� ^��|�W�Aq��i����B �sd��� xt����1�8�.�	�P/��K�L��׿Ќ
J�X�@ �iW��G�t,,;:� �pJ��\e Mk�E�Q�@; ��3
�(\�����Q�-��]�@K���!Q� 
/�\���ՠHQ�@�u"]��HEaˠ�����W&Ќ���eJ!xR�#�.���V��w��fU"��r���C{t��ι�!�����Á�N]dT�"V1:��{��*�<�B 3���e 姃,��\� �;���i �����7D��w� r���~.����� �������EC<��O�W�Hi(��]`yL}�h�|�x�V@�-�d|�zZ�H~My�:�P,�TUaiP�"(yԛ��)k��	�>7 ��y�� ��:Z�d�-b��Me"]�'+����5R�8��:Lp�A�������5���� N���3��QЛ�bG��j�L�x ��ѩ������od�
5"���PM�8`P�`:���`g9��o�����0s!��o�UM ��&1z!)�y(yr�;˗�"��>P�̛P%-�rB�4���R���0}��7��j��°��d���pdPH�`��#}����`������WS�a3�r������o�����} '�\~���� �W��B� ��h.���� �\�[b(֌p�iY ����� mh�-��|7��/�&�(�� �����D��� _r"�LK��B��2𻸳a�� rD=n�� �+�/F�?lP}<�� ��u!�3� ��^y'�{MP��q��i��X�}��� �u�T��! ������� E���҃ ���\)c�j0���5;v�.��o���p�[��a�`�%�QVXT�i=�J�,�.1F��I�*������'�S��#�]��\��`�!=� ��e
P�:�%��Mi% }�����YŢ	`!c��K �ªr����h�[ >�l}��N� �������:1��� m�f q�C��z�#��8 }�JZVLX9yD`8��! SZ<]�'
�̗(�ڀ�@4��@PL�N� ���)���>U�;� �Q��#t? |� 0x�������L;l� c@���������0��B<.oݨl@wD�V̸@�$�3^�; :e��]��M��Ǥ��E� �yI v���w�5!�������/� Qid}jt6���`<�� `�a��)�|������3~(y�ǐ3���o��ɀոc2Z}e���t�\�*� �%���� �#O��CG�^o�ҥ? #�r��� �������^���n���&� 6,��X�F�C�������� s��h:�[ ����?�� nu�-Y�W mf6���� "���\�FN���������  ��P�� q�ն@C��L0�#n��w� ��TFq^������J�� L��M��� q����#;� ã��"�uw3P���R޹ )��a�k^? ��|��� ��>i������NSa�^��@ 
'���2��#�73 ��j�� ��4^d�C ���y!��f@��<i�0�� G���5E8�zs[����`�0f �?��*�)���I^�h������� ���{Ͽd� ���Ȅl, ^Ts��y ᮷��*��Fd�����6[���PX^oG�@ί� fx�]�_ Z�塥��Kx +fcl�^�� �����%ut��'`��� �b��&^�> �Ez�, t|������a��jU����]����H_A���@�U9��D0�JhX�] �C�2����� �@�> �W2�ʱ ��]�SY'����X`�q��� ����@^���]��U���4-AŠ���� ��d	%^�:�2��~1��v� ��`\p��8��ő=^S�`�������O�i��� �ק/!�*� -�
h^�������ޤX�  %me�^������� +�Y������}�"5 rp )�F�]ٖ�a��!Ы� �����{�_�u�^#�f"5� ����%;� ߺ�b���]v:�[���/�x�{� KG��)RF�|~A^�2��Y1� �� i���Ч�$����H`��V1`��g�K��8����$�� �|B@N� �^ުC�'r_�X	���=v� �o^��H�� �J&�t��(X�B�SI���  Ԙ��]�i�<�LI� �����9�� F</�E ^��v�`��Px��z��	��/_���C�)�y�E-�H�@4��$�� ��S��P�� 	��'��<u,�� �V,s�X�dX��1^���_�;f���F���^��׿D7��Y�؆� 0�h)j%��#��x���>5Z?��&0 �*�\�Y�^��&���b�x�BA��{�l�����1u�e�6 ���T��]��	��P� 3&<�'�?����P�Βx_���H�VC}^��PJ��9q�z�ۀHT��<�8t�?`���ĸ��EJ�C0о���$p(>���m^t `�c��v� ��i �d�n(�.� �v��M�� ?4�����^ �h]��2� �w���g�_����� \�p X����^ϻ(�!���`V�@4�
-d��	0 ?A�5^�v(,~� ������p�h���^�X�� �9��b�X� ���ϝ6P-���BV)���b� �8��U�(�g�ĥ��]Y��+���-U��U�� r�ǃ�J5��I)X���]k Y�}��gD	�w,� �70�>\K]����'��F(@S�H�{ ������h%jz10؅ ^ՙd椗?"��R ��T����7�����pľ� �'"�qσ�+���#$$�C J�]�W� ��uF��w:`��r� DU�~^������[d��ߪ�F��Ѻz(ą!��D���� ��eؑE 1D�A�N .ހd�}��� @_��Z�w�GD�r��p��u� ��iE��t��Jz��ů��@#1� ���e�rE���_��Ϡ�/�����x� 6$Q�M^�c�2��@�oxE�ˏGM�@:�$u ���������6��0��X��1.#8��r�C'�\�D���T� ~�h�
��!:�) B�kr�Z:��oE�!�=�x�t7�� ��X�����E���3��>] �.�Nz��)m;�O �����C�� �B|��E?���Rgp�X8 �/�����P;�% �o��ޯ>8. ����}������o�4K
ޮ �~T�ũ�0�b�WM�@E1��	 k�y9��>�`�B����=5yR��t�������v���6x� ,J��ߜ�{dF�5�R�������b٩(8� �/0��S�'�Z2��_��.�-�stF������0�$<��?x ƙ"!hMH� ��鳥A �E�7��&v���C���D�h$�@nM� ��U�߮�� ��ZC��N� ܾ�ýE����#M��⪒�[  |J.�^� �M�I��(]ߕt� )x�"� �?.���@n ��5���0~�pJ��ş���-�&����̀�V{�CP�- ��e�[�H>�  Ů|��	�� C.Ά�-�` $�P�S!���.�  2Xx�0�q� ����\��<��������o����1��,���r0���զ��+w� �E�/qϣ �L�����^,��Qr��Ц� �����5a� *�:t�������&�"���%��E� 0>�N���_/��4w�4P�� ������}EQS�񹀨.��$�ry 8kl���nE��s� ��V�z�ŝ>���u7��Cc�-�60� �*�/�k3.3a4�~���2 C�`yE3l� S���4�T��	��@%~�� �/�_^�Dy3�+@�#��.����Hx�z<���o�V�u�b0 �N'���"Y L~�;մ�T�Gr6��.������@��ys% �Eʘ�^�X�� ���.�ն��B��=	�5�S����M%b�E�-u���� Ų�U��G =#VlF0�9 ����P�E�:�h�)���ղ��� �g�J�tΓ���� P����3u�` b�2��  nyjP0�r	�.�d��4�*� �F(��ʵ��\2|�)EO;�
^�<-uq�	�%���C�^&W޼�p��b d��5قE�\,|�Ljn��m���u�� <�k&C�¨-������?����<8z���uǛ�p)�OY ���9���e8�0 ��.�uQ� �g��w�t�:&���y܂����Q.���A��#��D<RC(��� `�.ǘ�Mptrxߐ��EF`8 ī���Or,.q^����\eߴ��kCp1�[Ϫ w��2�\:��0��� ���E ��(�~zژhR�u-n�,�{:=��矌/CԂ�5���+�-�<<1 ���*.��	z ���t߃�� �r��k����� Ϋ��Z;���E#���
��	=j� �.>V� a�%5�?�t; ���V�u ��%x�4(��� ����a�� KzQ�ˏ $A.�?�� 5����{+E�� H�D��c 26F.����zZ�#���0�6t� P�E�-4&��0̀���.��<��C@P!�xz�^&�A��#0�?,oָ �v	�cH'� ��޲K�_MɕVq,�r�3��Ƃ�`@��� �n�i��;.�o��C^4� ������x�����e~�E�<ҏ�N΂m����G.M��GH}N�������]as�hS��o����α��/����`��o����`�b �=J��.����zH)�͋�ؕ&E���>s.���y����`L� ��q��s+!E����T��o(��\�( @�u{ݸ?U�mE-#��j��.����L��_$9�t�z!;�2��� �\]}��f�	��T�{� �`��!�D��* 	�9I�^A��~�r�v�Ⱦ[!�w���q WnK�	� >�Z�I2��� !�u? 'G}PO	�l��
 U]֬�)� j8!�\��z�Q�_؁	
 ��^]v-�%�7�!��~ k�M�	E�̠[�<�� ���d�8���
	��IE_���i���!�7�Q����� ~�A��f	i�(�� E��˃�GQ !����
�] �A	| ��H1.ܟ
!�P��2�K��'IO_<� &�P�>��!n��V`>��t�_ ]�	F r�#p�̣>!�:� �:`x��t)�]�� >\�6�!�,O'�F,���P>���Y�(\8� Ma��]��� ��L!�w�� 	�jY�_����\ (�cb��! �Z��	^%ڐ0��6���][yw�?a�k!��xFMQN�]�@ln R����yC|�:�!��Q ]��^0f� C$�?(�G�$'����r�9?_o�A�P7 ��'�!f�*���������,���>&v����B} !�3�H8��Y �\�	'N>�!�)~���M�<�J��P�`EH�P;0���b�IJ�v� !�af�V��]�&	R�� !�b���C��� �8�t��n>N� [	)F� �aL�O3� !�Y:y�&�{W�{d�����T�#���!�m�"�VI�^�x
BFi6���3��������tV@n=��{	Y�N�I*jT�� ��	��_��%� �Յk��-"|1�D8�i�<������R�	u���8�<lIn�!ȉ�] �ƛX�`��	:�G\R��@L��t/	��nI���X��l �#��A�7 ]צ�_!�( �M�����EL��	ΐ�����j�y���Z �(�-[a �+	L�e w;�K J3L�L@' ��=P	X7L Ip.��H����0T�S�1?  zt��P��$ฒ^ 9{�.0 7�`�0El�'�!��༽Lܼ O��2�#	�'�@D:�.OU������( �J�����]�	@��@oNL��\ ��Mf	��y�^���p &����!��O h�3)�X��_��N� �Z!�%��!뉘9��!�����<6���N d�-X_L�	�S�+G��'|��9 d����d�f�F��� ߖ?�AN� ]ۧ�Y!�> ��3	,<�� 1D0QZ����^e��!�% �M�7�ĕt� ������������9L%�X(�D���h.�a����h$������ 7��	`\������������W!�,@��_� fu瀀-Չ�����H(S� �m��YΌ�as�8�P��N��!Z������8���0Q1]9�s ����T�!� ����e`H�
]R�2��6wài����\�� n����
�Ô]JLp�.��d+I�@���`>�&Xw�	�D|M����7r�~h��HN`���^_��W 	/Ѭ&]�<���h�!����S�a�[ �L���\�'�!�:�� ���V�	�v	ϩ �l�4����&E������d�@^]�x;��6�����,��"| '��;8��	D�V\ ����Lw�&!� �[4�M�|ZŁ� !`�]V:l%�04z8��v��H�� fI�6�!-S��\�D��r�o��E�@43H\$�>fXnz�W���0=�@�vFY2^:���6~ }/ �i��!��T��t�8����	gAc8 ]��t� ��HL� ōP	�jzI�lc��}ߏD�p�$a@�ݾ� @sW�(]uS��:�� ��E�!/:[� �PT8")���	QJ#�-��p��r	�!���4�� >�2q�|A L��ȨT.�1�&0 ��^�|  NA]��	Kg	P�j���!&�t���vu�nľ�}��L A���"�F%>��8!�����i���B�tA[��`���T�,�<���:  zqJ���D���! mup"x>>�P��p?nb|�>O	�,`JR��ـ��v�� =	�pI�]1�� r0"�Dl��%�����}ȐH])��4��.������9<�������]��0	�\��  �$]�q�qO��!���0vfY�]߀ ��<@���<�C�� ��QS�>} �	_'Ӹ�Ƹ]�� p/x��!z� ��R	�nY��而7�.>r ��)43��>�~о.u��	n�m�q!���ž�`�Xu�;���Sx�,� \��� �H1T �F��]����	8(.���� �H�� �6}^?��z��a<p�;��߸/@����<��p)]G���ѕ�!AĈ��^�)b ��i̒a�¨V��Cp�.>�K�� 8�y�� �]_�QnM�	l1(#��DP._� !�E�|<̀0O\���H &���>]zb��>l�}��E6nˀ�`� "B�R��� �!ł' ���?��t�;�!��۝|���5�)=?|�`:(� yi�A>+J�Y�_�,`� vI�1�dG��	E ��^�@G�!��� �$? �k}"a	�@8R� �
�!9���^d ��\�t��� `�/+	p(�����	�*�7 ��z�X�xI��´X�6���aN��x���?����Yq� (X�	 0(�KLF��$�5l R!�vr��6��iC)� ���T`��0���<�` �"����]|�(61�X� �y�	Ѵ���~9��WM3`�q��B��ET�L-|�0 ��d��T���]up���E�!mK�o����&Pk�%ʈ���x�� �o�,�Vp T!��9�cM�����K� �]��?���pSɑ$`0�w&^;h,� d)�ξnp��p� ^%�g�{��|��N�<������p��), �VN/�$wڌ ����:��� ��~R_���x� �p�	4�� ��n��!�:|%�h ��]3P4	.À*�NT��@�s��>|��|�ّ][!P�;���� ���-2!� �P���&��^� Ԟ��;���ӧ��L��` �}�^���).l��s��9��<e��8�(��; [�>Q�	p F6Py�Ҿ��!��"��_�a�J�`z�s��|N&D{a��٭8���nL��m�ʜ�|�x^�P��h�γ�H�-�}	,�1Q �JcZ Gِ� �!��,P�S��G	Y�x0�q�\�n����,!�XE ��2� �<�	��� &�g��印d ��+K�i40�T��8�4?�hL�L>�8ݤv�
n���� /��Z���sS� ؃ɱ�H��|:fH������x���0ؠ _k|����s�x: ��H�>��!�[��새� �\A*]�ݐ�f�<����C۾Xh ��kJ��P��+a\pU��0o<j����P`Dx'<�͓wt�s"B^�P}7���x�X�|'a�U2Q��!� h�U.� 8ޑ�R2 ���	�/Ѫ�q���U!�����>��j�]��t�I&�,܈��|��=�	��Y@�?��!n�z ���v������6 ϙY��~�\A(&�u�\�sŭH��c�F�|'�8���$`�Xyt^_�@�p��� -ǣB����L@�tLU�����C��P�1-�H	�JI�`��SH{�:�.r�!+,`� ���&�ؼ		�%.��z�iL ���Qƙ`H�b$~� �rz�ޮQ!d��Ф���6�]7��fIX�,^@��x�%&�H �^)��-�FPAd"ဌ?j�&Z�0;��#-� V��*	 ���r�5��V�4�D�i �1��A	�[�+0�xpE�!:� L�_ "�t����K	i��-���0أ,��Q $n	<�ˣ��A�@�5���P ��!��1^�Atf`}i	XD ]�E���l�H �����mx_('��b�8f���Ϲ):�$���жL�]Y�?�L� s�D�6�!�� ���<�/-�:��.3 �8dǬ���4�p��ST �N|Nt��
�$Q��{�!�^d� H��c�]���ٌ�V������ �%+�-[�x��d	��
����9��<0�#8�UM-D�@�h,H�* ��~9'�M�N%	�\>0Rz�d��,.�l�Q�1sB�W�I~p9�Z�����6��.�Re&�^5i�Ӹ�fy O6���E�������}�XL�h��"�
@L�tL�G��0r�,��'� ��l.�_���:o��@�]�ܨ��bzĂxRИ�tZ�� ��	�}9?$\]8u����m�| �!�w��,M"`�%@��\ ��`�rؘ�p .��p�sF��pX�`��ipԾ�P����B��V�4$Ah�<�� 4��6B\7�	� �	Z��X�\-z��s0h� ̳ ���]�ᡀq���{`e��t�̄�.��Q��^�c 	7u�]�b��J�)� Ե� G]�`	L��p C��$������`58�9�7������k�
$����8��o4�@"�|�2I��[�� h5�+ 8��"֩ G��,�A
5δU(8�@L8��B�9f8��:�����Y8��-2��h .8��~wx��D|�  CB�	y�P��`A}G��3���Wb|�Z�%^�'�9U���s��S���0�a�P���{,�L[@ǱQ�IM =z�~ �FDG.�fWBy����嗐�LX�x ���&q9b�<4[$� S�\�� W�m�̣q P��<Y��D zZ��0(�� I���%�<�� �O{2R���SG��4 î� ?B5�y�J�{C,9��X��� +���mio�Us֓����?.O((	�X]���+�ŀeI�1;�Jo`( �M`("<� h|
R>������S�V�z� �G�j��� 3ӧZ�?I�Jw@[s]�Y��'z��^�m	1gR��� �2����A�P��0�G�h!)�W��: ��w#�P��?;�8C��LʏHz'L�s ��ı�e� ��J�Ԑ>:�!�2�5g7� �K0��s>)EF@��IN���[ w]��0������| w:BSU�uJ�D� �=vRHO� 0�8�)L����"��u )_m��t��,Ѩq�hYԀ�'od���T��n],r) ��
9�4d��"G\�` *ɻhxYF<}�L�H�f@_ ��E���\����ϮqL��Zg�7xa�8n�m�@do\S�}u� 9� ���J� ,�s�� x[1]��*� Ӥؿ�Ȭ6 #-c�����)
��r\B�R,�G*��)f�l�-��(� �����)�/�x���ʯ��R\��@��+% E�I�jm�B �o)V"�;�̝f,-�w�r{�c���آ)H d>*O���'El^�	�3_y �"ը|�} (�2d)F� �L[�J2�]�6�m D�bC�����_�f#,d4�q�3�)�I{AZc0 �L��\ �r��'@y`��u|"��ܥ����Z��x� ��͌!,��LX� 0L>5]� �}\���D�G9<��-l�s�՛�Y`q(Z�;]@���\& �v��Q,�c�m|��@�G�x �� <KC�f �,j9�!�'���$G�� d�(�t��Mn8) [z]h���B\�NA��)�D��Yrĵ�x�� �ȡ~'�[Ҳ)���и
r��!�`�olm�%&����K?(� @'wEb�",Z�z��|}��˶W�@@��2$B�c~��%�5�]��\Щ� -���)�,���!?M���߆���"	��	U�~ȷ�P\Q���� �,'yՒmF% e7!��S�ckZ� _9��Q��,��"����I(�W)�^&�V@�N��c|� 6in!t�l��)ǌ@���`���f3,n��� ���'��.5 \�()N/gw�j���# l~,�8Dj N�(;\� b)�42�k,��gZrA�A�n�����\mOd"h�p�`��,l� ��ӀpZ\��'
 i�g]P-)�,��\��[�(0L��&���m���f�䱰� 񹠈mU� ,�΍��' �x\J)A��&8�m�2v��p����d ��\(M"�)��F� ���,��c ��<PA(T������m�yR��@�,h� �"��l�@(?��t��!��m���& Z,1�5=D L�N(�!�) �2�V�$�|�l���#�b�Q(�~�)@M@Z�Y�KI�P\<�πҔ I>RB�)�l �\w��! Ñ,7��x �)2�K�\ x1�.0�l}8�̸,�'���ļ�+�=�!��t��,݉���xe�t +�@�)��&���(�� E� 
T��hj�wn ���BLԟ \��W,��(�x� Jɪr[��) ��@%՝�P�8t�	�i׽���
�q��g�An�;ם�, 0���)]��R�Ǟ���;�,Yg0�ư�$)�� >�&=-��P�� �q� a��wmeO,��tx�p|�~�>Zs� ��]#Ty�|�� 	κ�' \\�� 0)��a	\n�]r6C`��pL��|Q_�D^zѦ���!��q"�a`��P8�;c�_�WV@4� �'ݢ\�$`sl�	�!��A�0,xt��I�n�� (5�m�x� ?��ta��7�����,�Um�����P	P� -\��� +pc)_�%0 �;ۗȨ�'�pf�\��y>�R���M�%,_���l���	��{�[��-��0�L3\�>0���x`�� �Nr>�'m/&��9ĭPb��jn�!�@p��$��T�g= �Ɍ�,|�6rO�����y��=���@��� Mǐ`:y�m$��	���L�9t�(�B����|\5 n�.�lLC,�����t_�?\�[oTL��w��b�|� "�3�)E:�� �k�6,�>�g�l����iR(]�/�������`�(휺,�`o���@�J�\���Q*0�e
�*H74X,~\�.���@ Wc\��l�v�9A�������;�/���������Hip !r,m�;�# ���Y(D[�)�|�� ?T�إ�, cn�#i����(L^y Pr��1���b,eħ�� ��m�C �'�@!)�Q��4@�o�m ;�,�r�
4 �r��Q�؂lq00� ���\�6 ��d)GI�n<!����`�,�}p��C+���s�(Ȁ�v��{�������)������C'
7���^���bj��F �'vl)�� ��J���y,i;���pb����KjA�f�����;dd����O�n��[�5 7�)F�L�� #�ylB�?S�� ���G\K A��i)���|m�ovI�C�`,ad '�[<��\�>�y��~�����]�pr��Qg �l�F\�V(��"*/@��HU�(�����\���}�0�3aY�����s���oHt�>��/����L�� ��wRl���: V�S(����\�4�3_<�a�� �t ,0�}�[�˃\��4��/'p��H�L�x��n�����.\X8� Vh̞f� �!��, �+]@��\�:)�6u�#�`l, �F�S�O7�X�� =e)���u<���l�&7L�%.B@~��n���k) R�o�,���8,��D >PH�i��?���w`)�g��sl	���H,.�C�)�z|]{��7P_y��ho� ��^�5�Il�Ոl��a\���(���{(��]�<���C&!���dN���X�����J��+f�� W�0�����,��,�|ʑ0L��;���#��� �n�,�0t1 %3�#��BZ5�"P")��zL�D
wUr�� �)iv(�j�[�5���Q����0�m���| 1���:�@��R0LB W\��T,l�ś �6t��&��0 ;��\"�c,�!n�-H��  e�R^(kP )���*?,o�g�mL����-P(
aJ]�����k���o 2�Sm,�;�y ��#�7��H�� zA%eU�G,T6���nb�r�\W  k\'X(��;GВ�>���+���P�m䟨��2���Y��Ϳ$^E`R��)� ��xi�jI�\��`85� �)z>[=��Z�A(�Սi��� ��4���\��7� Xc��Eni}�~\��Z옦p\��]�� ��'��m*_'�zD��� ��
L(Wpϒ� ��\�m�V�$M��܄����U̹��z	b)�J �;I�:�&������TF	2L�n��a���(�&�G:,�c�hث�X�dH�0%�'P��m�M�@�U,��#�l��)�0�K��, ��yH�9�&z�:]��{�8 ."4)�W��/��o�'����~pWE�0�*�� ��x,��g%l� =c�#�Z|��(ו���7����mq��HPJ�^�l.� �AEol�50,L�c�0�� t;�a)�{<s9�T�m[,��FK> `�oe� <)���?�8$vTo�a���&�p��)n?@��� ��7l���\�� �<B�)�vJ^]��0��� '�墡$,�(-]��2QnZ'��\ 0�)��Y~�<���7����J�P����m.��o��q���"�i3Pr�@��#���F(��"��] � ����,��Ԙ��Z�s#q�?�	3�°�mOD �� U�	|�=s(Z_���F&��/1G!�C��#�w�	�\��(�;0)K� �XAGm	M�� 6,0Vz�g~�h�[R3���,�At�\xr6�o�`��g�C��b�y(���)D8B�����K¬(�\sca�Lt0x=��A�o�
*!��,8 �Rh~��[ꨞ<,�x �Z���Ðd�l�B(��zaZX����no,mv��CH��ƥB��h\c��;�P)M��n#��������Pw� +<��[��� )#�������R ��X�#Į(y��)Q.�D�g�B�mS���0}+�%>� ���w(G���0!���ٿ� ��uL?�`�������4����0L����mn���Z��I>B0e,���N,�$Q���R��r]- �)���x�SwF P�,��! ���x�)��L��|�9�m�+,��,'~�� _IB��|k� /9F�L�J#Us},�VTr �A��'�-�r,�(�d�		��m>��a1���H��	�]BXT��@2+�!E���P��Sr� ,\�G����| '�T�� |d\B�)��"�M��0 9� ����E�3](��}����	q,_@x���! �#��l�~(Ǭ�)W��� �yh��Q�* PU�`����pu�M(�r,<��g���� ���m&�� w�@<)�I �n,�~em�� ���W��<2�
�\#���� �	�ᚸ|yo$�i{ R�z�[��H:��_p��6~V���8�&���rX�d�1@!'	b�.Řh �}�P���8>���\�B� ��l�)2_{�[� ���s�\�dhC�a��;P�ԁPO
���p�G }�2<Mg�o�!`��Er�� ����yYX=\���~�C���!$v�� �i�'؁��,��eG���!�a��Hl�Ж� _v\Y�%*�j`�
���?�� al)ߍ9S��@m\�|���(� 4��;�@"�[_+	ц�U �>��Bߘ�*�LQl`� s��\�<'�p�l����!4�r�[������H6X ?����M,� n���vK� ��x�,]����D	�O�r��
�~> ����'���F�`\�(a9M�m��8��U(���� �p:%��
�:@-! ��)���(�_�D�d�h-'�/���Q� W�)�=��$%��K� �*�v ~���Zj�)@s�	J�\�&?L6I��c0���.��`	�ix�͡t	[_��`�'�zl;�\ �)P�5�GrZ,H�8�j[��W;�zv�T1@ ��	�\��/�� �`?�S�� .�f�)O9BW\g!�n`�8&H��\zmE#��d��o��i� ���$P��\�at�$��X ������g��F����$� ���{m�����+v&�pXIJ,|��	���
B�I�m�H���	ۂ�SoÜDp���e}u�2	ݙ��_hXx8cK �B�):�zE�_���kw ,�Ng�m� ض/ n��e#}XH ��F/!�$���,��ݻ�#� �"J(��l�P,4h�s|�rp�W�)���v���Em<h� �Ξ�U%��\ �)����Q�&���"�|� l�o)���'� $�LŸ@�=�I�����;�1Xڹp��_� �/�2�b��
L\� z|[f�� �uV��T��&Q( ?3�!�zIAڳ'����5 R�tC��L1(�F��_&;�\H�&�LH���+@��g�o�- $?�A( _��8���)���&�Q2�,�/�� ���!��-�)Ȯ�; q������?�,!� P���QD)]5Zh`h�$$�6�-�X�<( w���)|�t:��BA l�R*L��,��Q: ,�0\�ޣ���~�gl��@4�nL�by���\;`\�O��Y�%�|l�X��� �eL-B(�ܛ�|��`!�,bD� I,���xP����L�l�����Fb$�IoBr'�Hd�t� �)�{F]�x<8���Q.i�
�m$/� e&�p�)y84��-	�x7��r�`���n'��l�G({��!���ù \�m��,l�����Z�$�O��U+ ��r�M�m| ,�Y�ev���$Ѐ� A��dJ���}m V��Gn��I2�0��%o����S ԏ� \H��)�!�pQw���J�֓l��aP$h S|��)T���M�=]�,r@P��<�6 �L �^\�5)E"à�� �a,Pw�oLh�p`0-�]<}�s\b����D�g�l�C�^ZL�����>�'�C� ��҂Y{>���H,����_�����Ĉ� 1 &�h��+ ����)��C/'��A4?�I�pZ.�4��&���*��(��ڮ� nlm[��9 ��)�!�>C ��2,�Ƙ� ݸܹ�\���+W ���`64c�	��qPg�d�,N@�5����'����<\|��;�j��"2��=m�n,͎v��R}*IZ��1�� �Y?d�(���g�m� �|�!�	<�y�Ԑ�]/��6G!��ya�D͇��Sc����I#yr�,΢؃ݣ��~�pD%)�����]0�ɗR�9'�~�� �+�s�g\*5����N�Z��l��Ln� ��(LC�Z�U��p;5v��z�� �)�2b�L`
 ����w��2W��4���0ŭ�,m���D��G����~\9�`�mx�%Q`İ�,̙�� !h~�=p(���`:��}�8m0,"�"� J�3M(��u�E}� [B��,��3�{�Z�� �SK^�W�)� +��m�}tk!�, ��Kd��
�͋'�)��@�����,;�� '��Q%� ��A�L7)� �@l`�Y om��3����<� ����)��X_��&l����p�����]����"?�z���~	`�`g�x�)��t�J���@',>m���Κ�1h�w��\k ܶ�@x�Um�G�<g{ ܙX���VK��t�

n��0x4 ~�]|�`\�f)�I�0���7� �6̬ژ�
�J\[�0�i�� ��:9(hm%<�,�s�7P'	{x]}�L�+���b���C&�(�D�Q�)\�|��4�R(��%�'\@bO��~�n�ʙ�#+)_� �&N;�IlK�UZ<�P	DȄ�� ����,`�3�%{�!�ƨtί���Ę(w�<�&#q��s(
5k�\cwذ��Urv��|�In~ 4�qu> �R�)�7A�o��m�, 2R�\Ow�Cg)B���`J��A�& �
�/}�)� H�B(�<@ �wS�"�E�,3��!���i V(H^�)�$���;d:�'@� ��h�a∐ I(�����6g�}�R���\�@3r�BH��U{�&���Ұ,:W] nŴ�$~�K|1��
�"��­n��� ?B}6pA]�R0�����:�,��n#$���B
y�X?o�P��	�Md���� �~�/��p��Lr(HV�?� o%g��e,��D�=��Yg�n�� .N�iw\'��u]�)D�}: �_PWUrН`L�N��	�2�������k1j�F�D�)���� �/\�l��.0`;��m &vh��d�h��&�h ��@(��}�z,����5Ø�%�Dh��� }(N��'8x[��L�a0k0�q n>�&��|� ���L$	xmo���
���pp�1%ԦGScN�Ld�	#Kp��T�� �(��)V�t� ���&�-*�h�{��F#�"��D�DtZ��*N�GO\
|� h,�$1�D�i@&�� ��5Y�����lJ�����>�B>�X��&@�� b��l��9���%t0�� 4S7�95�=UN��+�\- t
�J�Zs���jE�7M�V8 ��d�� ���>M�3y�H�uL�Hn�9`0P,~� ����w�>�\}��|ı��0,e `$��qm (R7z���T�訌D0��n,r� ���޿��.����T��Z �njm ����'��  )�MF"QRes,L.�ވ>�|Z��i��)�/k='��!�l��܄ �*\3?�&��h �c�5��Z�,H�1�\� �)���] ��q�%�{x[1b�� `�Vt� %or_(�"�)�<s}�Hj8#*%�����գZl���Ե��o<A�IO��L� b��CMd�1��� � !it�	X�]�h=�B#c���O��)�(����{��>v\�Q��,4�/�n�0H�J* )Jѿ�ȊJ:Ҽ!��kKD}g\s��+� i)��,(�Qx��������h�( 6t��@2)��<R�Y� ���%�Ę/�w (-j�]�58)��y,o	x( /PVXa@	�[(�R)��R�
k�D�,*:~^?�t�7&�wȨ�M�dU�'��@�@
l�L���r]f�T����܏?g%���	�-�VU\�Kf��@4�Ci3X���l1%�P� Ǳ�d��G���c ���@��YU8��s����_���#�)� �"[�Mݺ��f@�lnx��հ1`T& X(Pi8t�	j�ކD��~Ԥ\l�@b#)���&ĦMP雚�%OxQ0� JqZ��)�������H6,*ct�'e�"����y�1v[p��n�E�>��4* �9��m ��'�&j�4	Q��y�$pL����1)a�<� ��Rm,�.r`H� �� ���	)���� ����mi���78 ,��!��Js]���@a�����7o� ��B̈4@0�+�` ؼ��Q��PL�������"���3��x���� .஠� �3X`�< �J(�&�)�4"n g��lH~� ���m��KQ�8� �1n0"gY�m;/]��j@�b9� E(Seik|�=�~H' ��E<$9#|y%�1xT �%�>���<_- (nQ���(�F{��Ƅj�:�������@�� ;�����H͆(.}�tc��`�p��B�MҀ�'`�]Z�D�F'I�8��]c���m:���C���~>1\�@���RFH�\�0���$��V<XUv�H� h�y��BXs>t�t� �%� R�Dn�X�S�`�N�">�1s)@��u�ch& M�O�k |�@0�4[mL�h�SH: �'@�5sgZY�p _�c�ׁV9��n���qy~Ө�� �{�m�I�Ja�@��ݚ �����3��B��� �_PZ�#����O� {�c�C� ˞���?5Z�"9� U�uΉ|���i��<���a� ��7sDW����v; ��[ ���|T۝lZ�"��̀���ߵ���a =�ͮ��-(5��b��0��n� #1���N� 5�:%��o� |�.�_#�W� D�֋䎻]�kq���l+¤(��v���G �K�) ��S��iU %��#�k h��r��� �iE��� ��K�NL ;���wݫ�� �e�ψ�:.
gr`v�O�6�: �o�2~>�����8�r��B�z�HZ؈Yp�0�/`����ɓ��6��O3g@� K�f�D���Ά.��>�� �/�Ȫ1秐� ��*��:� ��ϩ7�bz ��(u8�P.=�'���ԃ��q!�6�b��r�aġ�lTsf���`�(d����M�S����;�>��Vg�cө��' ������ ?�G�>�N; �@�M�5 8�iv����}s�\�Ro�r"���n�OC�� �͞q�o�����<p�Ǒ� �sV��{#�@��N���wI�H"�`�p�7Ȩ�g��_v���[o#�Dr��VA +M�'،�v �R�9Κ����&�6���P�� �Qh�y� _6��r	�.;b+��
 =��pػ ��g�� ��j\�f v���&�u���l*��!�� �p�H�n8b� r�2�Cs!���� _�Q��v7pg 2 ���r�o�����JN� rX��l�hptX�� �Z�vx�c �oFr�%��3���!�ܨ��9o���V�d��� �2A>�ֽ���k�:r 1�2K5#���(�._&�.��0L"� � �g> �qB��� ��.]Ajg �	�v �r �°!-��R ���?�Vf �	�rP �&�aP �њ�ݖoe���T���rv�&̀�h�z�w �!'�n�� ��:��T�J�j��n�r*�x�uO��~��"��B ���w��p� �ڨq��r� 3�sn��� �l������Q����D�rӐ��=���`!��䐤 3�I˓� 1���rǘ�k���f@�v=� �"s��x� mr�[5iB��k~3�`  �؎��g�|'�rx�H�u5��`X�lP�~�>��[�̐� ��T������W� Mt	�R(��if�9w�p��©�>/��X{`<mY��q�)�rNb'�z�[2����l �T�mqR7(~��`�e&&�d i�cp��P��:`��?r�H:��0��G�,�9��~�A �����>rx}����p� c�*�����:�J �����r��	@�A� ����O�l�
 i#��,�?L���rfQ\q暏� ���6�u�cA��c՘8� ё������� D�_پ�C�����@�� �6��Jty� �)uO+S�bo�rI��q\M&���ѣ�,����	rS�N H����>�>l�n���/a�A4��0�'�iA(@ӳRlk����qH�P!�i 	|�/9�,��� 8�p�D M?2�qr4:�]&GZ *�۹L�����,�������.Й� �{����T%�
��72��@�� ���Cr���� Yl�������Æ�������<����)�G�v��y�dW=��+�;��Z��>`w.*!�^���Y=&"o` �y��	X�?A�`;�����������l'G��Mr��!�o9F�{�$a� vz0,W,��)=.�~JO�0����W.[����e@�r o�v���� wp�~:�b�\6|2+�0Vpl�L����T�~�'��=˂Į0�L��?�sK ����v�u��:��@�B,l���l���'�Ͻ��t! �\ ����D,"�� z�q�[ތ�*���U�$�r����
0D[Z��q�@"%7 ���9!n� ~g'U���r�l�z��ؐ�F�/i�����^�H�2�d]��9OQE� �Xr�X	�qu
�h�w��� @�s�\��r.���y�`�� pL�~ ����A�:�X�d�	���`�r	(7�*�s է�� �Q�?R0�>r�L,Ǌ�μ� �n:��e�.G1�W¸Qrh AZpj�Ȩ�(LR� <]��N��$o4�!,���`�@� (�n����� �b��F�G -�r���C�=�$��~�+�I��^xW&u������ag�u( $e�q�Y�r�� �¶�-G�"��$�.�n���rЃ������8��|:?μA ��w���.�r� 1���~ү�X!TQ���C �	P����H�` ������7��VY��}�0�j�or�%E@�<��$��<DhER�I�\ڱr��n�A�����ʍ���3]jt
UW�㤾���Kԗ�:�d��:�7Ǽ@Q�p�=sz���m<B�����r0`�8.�
E�?BB����,� �O�����Ю�1o�����,=)� 3�{1��?K @p��."Ɛk�b;���� ��U�a�@��;��%A�gͅ���~�`� ��Ι�_����d@ď�gJ��@�p�� ��oVq�".��	�h�<�I���
"��7�d`bs��4ro%�v� �S��L��.��� ��%*�jz�H�J tbBk� s�ͦ1�21r��p�0�c��vK�6 ����0����0Lf	��s��@~��	��2�!A��I ����qD0�H��h���� �H��UB|�r�. �k�=�, ���`a�Nd��[������r�HY8 `�D�5�atxn7[�(��aE^�ȶ�H�<Ӛu��̀HƁ&"���B�@�� �|���rA(M]���<�����1&n Ǣ �r��帘 m�q�X	�2Ӈ�:QM�r��ӱ�6@�qֲ?)�B���'��Q�/�cè���bpȩ� HKMGN3��.*�Ѐ��I� x�|? qF]~&��,>ƨ� K/[��r'�mJ� J���~���h� 9·����g��d{ ���ϙ���[�~�@�r" M���׬����0.��m�8�r	�q����������$�P(�+�<��KVx����� 9�ɾ�ao� �{�pˉ���	�b��c�Jt� �}�����@&Brs���$��n��R���`x����F8� �k�����ۿ$P����;A��!21H�4�� |n�$W���Ub�h�(���o,$ ��w�?��n`�ߓ��>]��H>���A�� s�^Q�x-.8��g�w���r�>{,�(�c&��L�3���mp}s|a�t�\���Ϥ�� ,���{l�>X�wW}���r �\s�ڎ9��~S��A��{�>��k݁(r�(�mn�� p!�^�T��@6�Bx�{�rN���-C����� �a9.o�~���#, ?L $Q�����ί���Z$H�p 0O���"
��β�{e��|�8�*�ǰ�aC�#�Bl��e`H�� �zg�t�f`�r��;��A�7� d��]�5	_y��h/ITq� L���?u� l����@���PѨu�%�F71�(���$�[��q����LoL ��h�	��]R,�6?�b) �IL�^x�K}�CԚ\��x�,��L �"�e��H��	r����9t � Y�Θ��-��H�Ԡ( uw\pf��$ȸP(��&I$w�����8��2�����/#x;��=���r����P�5�U3���N�`d�0z*8~� �� ���������T� �H���Šr*n �J�5�9N��|m�H�;l�g��r�-K�Լ����:���`������<�e�{���0�B ����^���f`�Jr#�pU�α8�h�� ,H��|� r&�#ue�K[� ���w�t	�i㳀DxZ��&�.� �f�F@_#�B�Z�W<��3	�����-��[ 5��R�~3`��Q��2@�l�A��0� �	��Ό�� T�q�,n՗ ����0�� �r3.��(����s� �����d�^r�6�=��B(���Z�<��� Hs��E�	ˏ�P���-�r���|T��$a� ��~�_c���<���J�zcR�
�j+`d�t� Z�WN0k��.��|p�j~����-&ˀ$m������~o�慠&�PQR�0W���	 <i�{��,� �q�<�r �81?�!��&�k| ���ם�aSB!�r�h� ������ �͎�Rq�<���rS�<�(J���ܻh��+Ҁ�ex
�P��� 8wl�±���>���� ��>�x>�� �r2��P�d��:��p�?Mד�IzpD��0��_$���<��HK����������g��"{tVf(��!�6k�0�� ���pZ�m ���rd�����> ���s ��orn�J�$�(���.���	����`�6?����r 7tZ$��A:O_�8���b9����0��q"j�X�}��0�p|�;��������L��5(��"h���1/�dO� ³rs��B�3 ���S ��2�:�L���/r��+,l� ��7�Kr���M�� ����g���P����K�Q@�����H�(>���,Z��������`�٧=�� �ƛQZ{w.�k�˾�Ov�~
��4��
���G���P`v�?� �b���mdy Ԧ���r>p�����]�dc� nAP�1.�Gu������a���� ���es�|��J����%�`'��g�
�h��� ?*V]d�	t��`�'��ݹ����Qg��y��E�� #w �r�
Tq�	[NP��뀘���,��A0������������ l0 !�gqFp�D(�9�>{Zx^�O� �:�w�Z*�j;��L?h ��������D<a^W��d�~� �p�0�����g+	\Ё�r)ao��^vZ���W� 5O��̗�p�� �"����|Y\N Rк�;ˆ�	������n�y֨��r �Vz�hs�����}� ����IF�9z�r4 ��p��$=΢����"� �r@��P��x� l[������H��1�c74��K?H�ȲT&2�@T���ͻ�� |lÊr
1������/���`�� }OŃ�T|�H2s���B���Db)B�� L��M|ېljcQ��&݃�2w� �OUt_��[;oΓ� ����B��p�ϋ|h��w����T_��r<4�0��~�* � �����q�i�� ��Fr�1z�8G���� b�]�T��jDy�Ƥ� �g �|�l�(胔���n���7���} &�xh �!��p��^��V�`��{��&�������X� �p����R��4S�q�>]��`N�~	<�OH`��Q�d�d��9|�gr0�D��oS�`���T!�.�/�� �ݾo6�)&q0 �J���$+���k�Dq�.bLX�: �B���� ��t��T�`���9�5@� YZ�E1O� rQ�"u�w�`�0�_� !�.�m�
 �/��r��t�|� *pꖿ��0J�p�s� �m�3�ЏP���&��a ��d�,�����ANb`��x/X�\ ��P*� >F�����'iS��Z���%�0.Q�w��q�è$����x�{.J�0@� ����kIy$���Pe��+T��OA�v�^<��-`ר��4�u���e.ШRJg}� �q���Wـ�Z.�3|a�́G�R0�Dt��[7� Z~'(��!�M��$� ������nJ��u�]-��*��.�����5�/:�" �r`N���$,� �o���g�H�q�इ���G^����x��sƃ�&�mvK� 8qL+s՗�.© �zP_4���R�0�Z���J�?�!Dr&�� )�=A� �B���&���\��1�]�,�,�����D��̼ �%@��� �w��� r���`�� ��E�39�2��\G����+�������h��u�&X�"���tr�j�7,��P���C`hc�ʺ�ৰh&�ph�A��b���VΘ��8bK�|r�P�;�����L"N�i�@��%?ϝ�>�	�� �1f�F ���vp�r�);	$�P�$�P?�H�:0B�r4*�hTq��oȤ�$ �sS��|����X� ��#dGu� ���so�L_ �PB�w�H�X`�mu㐂�Pĭβr�Ѫ~�G�@�#��.��T u�=j,��r�H�O'Q*�����J� �?��/�&|�T=	rO+�4�3 ��s���x6,�,@V/�@8D���=�k�ʓ`�M) A��R��Κj� �(VpF"� *��^�H1-�h�r o?���[��q�4Еl>��o'�I�8H�y���nx�ң rd���V��	�����Yq�s�I� 8쬏or��$���[<��F���2���&���ߘ��轉t��P4�|���������`�M8��dR���h��7]4�Ѯ���������n��f`H� �͎�;�rP�@�F����u��a�#����]��L��C�p��a�' ��,��9�������`,��^��H�����@�-�`HPqtt ����r9{���� 
�!�L�3�-�� 8`G���i�r.	�|L?�_B�=*��0-���` p��@ ��z���>\]| C�	.��Ø�\� ؕ9��@&�>�Aq�6A�msn�֒��?g�E�z�Y��p�� ��4��G��\��;c�� 0H���L����\Y�♖�x��`��&{��_u�.À���C���ԇ�}k�ɰ(�K�&͞L� BJ�1ɽ���b �Pr%���>��Z9�O�S�@�6��	Dx�@�� J.jy��Z�����N��hIb�
P��<o��Հp���Ρ�9d��	C�:y�E������@ 'W���N�� �Z����s@!�R��r����5 ����F��`�2Se���`�4h☠L�L	�����+ ����1�����j�>�� ��Or��x6� h#8f˟!��l=�k ��{�_�`���0h@qrva ��~�_�����R�z�&�~@�K��B^�P j\�'.� �U]�&u�\��`��@YFp��n{�;>���t��)*�@8�Nv���g���b$+�4�� J��q¶7��m� ��{[9
��r�-�p�{i ,���`q&:�$�_<7o���g`�>L8	3�=��qze�5�|� U���_\� *%n�y���M+�XP ����t
N�^3�8XY�~���f�'��A� �8 ���� oL�d !���rF
¡;���\ ���ѣ�T�@����@V�M��^�7$T�x��9��D�R�j��,�&�{-�� r���4����O�*K�� j�H+� ���s�2z�0 8���pĲ���Ho��!6�$�p�,��H �_c���/��T|@�� ��v�6b�g09��G*��dWF����0.:�� ���یT� r������[����!�+	�� �eS&�p|�_��tl�n�-��U�����Sr i2v�o΢:w�~k�!n�L �B�=���O�wb m��3�%�\��$ l �Au��h(s�� Kf-��*�\^$N��+`�v�2	�3�4�?Ā��L��$qP ���[��{��b� 0tӤq��U�R� ȜsO�	��p N�! 8��9f��m��/�V8P�j� �hZs��?(lz2�������6 ���\;�~�!��q��M�G�<���I�~p���Ęl�QG��Y@�sP���M�wmh�=b%���tH٤�1��'8� z�^;�lK #yj39=�N �6��
�d ��c��!]$�S���3(�/`���� �H�UQt�  Oå��-as�) VN�PH �Ϝ���0�Pw�g�~�1��x%��N\ TIE|M:�4R��Z{��O�Q �) �N�������lQ�� ���pS�-�}O��N��~��x�u���M#�僐�J��C�F|�[�lg���Z�K��L ?�	�O��P���x� Պ��2���tB�M@h&� � )�LN��l�(���-�|Ā$c\�e�Y@�O �N G�s�x�k�n�l��#��d �?*�N[��=K�O��zw3�a�m�Q~2|d� I�oN�, &`�<��c�(�T� �з�4�	���lt� �A��)ʫT:� j��n=� h%�>U�$�]N�-�J��L̎�;�@t W���l�}��X�O�a؀)���71�[0C���	��Yi�He�n�Q� XLT��xI�(�+ PO6*�F�)@�NP�'���b�A���,� y�2��ᩄ)�vP�S�MߌO0�xV: ΈHl1���B �DN>�}|	��m��3���L�^��9��PVc  @O|����t�P �N�=�1&*�0 a�W����^��A��\��l����Ha��@���� �c.^�l� �����a�X�"FY9�0�)��J�O y�/���wc ��xáܜTC�� �/�t2�H5�s �YD������e@ 4����I�� #)k�]_\	 ��y�O&}`�*�I���N،�~��~R� ��`)mbN �'-5�	�Ȟʀ�����* ��O��PN� 1l|;�r�bxC*����� .:�m�QWHd�	%\� ��>$l�P��˜�d� æH6O?NT �>�'ύo)�k��{�!��ZL�LQ� 4�钮�LH9T#G�dc��@���dZ��h��/ �a�܏)o��$�H�����G)��HlI��@��� �/J��O��to�bP9`���mX�� g ���yn�OY!��q>o���]@v��y�"��t)�N�1}� �:u��,�(, ����3��N"���Bx�	jh@;`` i~N)�P��X�,N� �Lb�a�xp(�;�x��,~N�� ��bz�J�+�r� �� �E;����v) -N�T_�e�:�:Ld.�(	QF���5���D#&�L����iOF�<�yNA�Ֆ)�p`�&a  �8QY�
`�i% ��拣vj)`3�X� |���r�%Vt�1е��i�`謰d���B)��Pa�/i�d,p~d�rf�U�$? qs �)��V6��r0 �*�A�x��u̛�`p�	|�F��L�\�M}'sAƁ�)����\z T\_��2qbg��K�H��d� ���� �W�l���>X� m鯽'INǿt�ӁD25l���`%X1Jh)���n�pH��L|� dF�s[pM@�pθ/CFW~��v�b���l���'�9p�-�`L���j<�yߛ��)lS!��-�<��(�а�Qe��$lx�܏ޞ �c���|ǲH��lP�"Y�p�\|| %f��0*� ���yN� ��m���dU� �~X�lH ?�k�߽�OPﴘ )ryK��l�:� ���O(�vF���N$��</�>Sl�  ��~�Og`_'�H���T E�ܱo�t� 4��a� =5iEK�Nu����!ލ)S~ΐH c�9alQ���Fu�r P��n�_8[Å�,���(���.��� ONF%,&��:c��/q�逹�l26�{ �shj��F B��'ݔ�� 9�<�� [Areٗp �u���x; E�(���� ���K�r� �t��B"?��s�h~����C'�D�@�����A������ 	pC�Z'|� &sWݛ,x b\����-J!j(X�_nKxN�t�C!J Dͻx:�?~;yJ���2x!]f�J�k-��gx�/�{JB�9��+x� ý:2JB��nex��@+�xk���̱��/�*"c;��.@{�]%@#���$%b���'/ �_q�3��9p�L���C�;儎��M@rg$��@�W��m�p�a,���k�q���Lʁu%s@��XZA,t�`�1y�{��v�c,�з�o5
��t�W� J{�^8n?;4R��YZz(�t� -)d%�/��$D��  =�}є���'�& �!��O���kCr �~�D�y�Ƙ� �,���w� &MB��d=+�4�!)EBv�3 �����{h��>�v�'��˖���F �$
k�	�>!Ҁ
y(�`� Lh�XM����?�����`�}L�!F�!/���3��K+���!�� �xd
Y`�C�F/��q 2�r�jF`���y��a��8���J �fV&�����f�Z!��U�Vi��h} 3���a����j~������� R�?�����$�9 &��Ӌ@%q������&G�E���~ �X�-�]m��s �Z���z���x�%����^u�-хK��^��g�L��Z<� !�Q��ez7߇ @�J�����xi��eo �Y�0�� Rt�G-&�ex%�g*�R5 Fr}�������y�J{?����i�U����ph_g3���<� ��0�J� 	m[�y��}�x�������;(i���2�����E�@���2�s��J��H�� ϵkI�w$
�����@8��o�	. ���o� ���dVc1� �C�����@��� �|y<����gh��C	��m�Ekh$^����!�P1Xv�}�2��kq��:�)(�p��a���=o�"����� x�,�qv�R>7��&tʃ�)y"���bg$, t��7h'�����%c���,믨8�Lg �����\� ��.���[���:�����<���J0��>�� �,{�c��m��s[��iΥʥ@�s�<
��3�<52@`�y�c H�?���V�( �.`0�U ���8�' ��r�Ƃl`/y������&�F�"��� �clB@��44���P�&���X�������e�x>;� �<�^0 1fav
�������X!( ��%�V��� �ih�����X.0����x� ,HjQ_�i���� ���}Y�� ��5�v^�`?H_���G���gIM�0Ӹz �\=�#�v�η���i`�h ��U�et� g<���[ LM�@��� �֬�bj ��(x�P� �6!W-� �"$U������|�;�� n{���0vt PH+��$� |U|O7?�/ �XFS� ���'��� �^��,p �԰�l�� 0�v�EX@ �|�!�炧�KD���8��׍����U v)�m�*b1�i��XqrRq����O�E! �/'�:6xw*��5�,� æ̙��s	��2 _G3��$ƛ�u҇F@Ӟ� ������ ��®�w|�'&�m%| �D��+'�@u�H��cd 9����F ����jO~��N� �R�8 ��<���=x�N���E��� �H� ��n�Q�� 0��lO�?GN��u4�aW0��@�M�1����I����h��S �}l�� ���o-�� �
Ov�J� ��{�y�: m�3�P�����"�����t$ J��~L� [��yRv� ��1�xtT� ��%P�Fl ﰆֈ�mA J�x?H�( ��-�:�;�� j�=�t82 ���+�Q���_�����/�V.JW��� E����{�\�� HtC���3���{�W0� i��1��x�8�<<׸�w����K� y��k>�M |�u֟������S�D* �s����a O�W~�E �G����� �șg�$�` h�Pr��O���U�/�`� _�K���# 7?�X�P	�1J�{ L��;dv� ����`����_�0GOfy $���^#�V)�� ��xԪ	ϳO�@� sݮ5ek n�VM���(�K��E/ kw�y��_U�Tԯ��Z#V�ؗe�O�a'lI���;�n�T=�n L�]0.����H �A O%xΤ�� zv��$����r�^���p��� �&W��K� ������$���:�ٯJ��b ���0K� `�|
��y ߻�v���~ ��?
|�uw q>�Jڱr�TֆO�\{L��-�x�3 ��mB[,Q+5 �֎����>O2�# �+̭Id ���,W��H�Te�I���=�1}Հ6`��f������'�. �K�5��e� m���ѝl9�N_��Gv���v2 �P�yN V|U�q9��
>�&�̆��%w-4��YP,�y���(�V�n �ɱ�7%�����=�W⦥� �����'� ����ߴ ���OC�'� з�-����8����W �U���!.� Ry3ҖO��|_XE?����� �EB�_O���0�{���� ��VH�� t���3�Ԉ;z ��g;֞���DШ����k�_�U�� ��TX���^�0�� p(�lԓ ��cO��կ�+��dB����Z�.�����۝ O���ER� �N�}��$�z�����ߩh�L�< �:w�_K Pe���^���*�x��N�7ϪM5�bm��@�H.��Ahn֐q`,y &����HOX� ��w���1��e�?�,fD3@�9�ϯl�֤��-� ҏ����:��O��\�=�L�Y Pҍ�5�9h_�e�X�Q�O�z��� |��#v��u?�!�� @��Y(���0��@�& �-�h2��!0�yv���2�HPYB�����Z]<֡8΀����7�/�F*��@у�� .�����>�NZ/���x�a`oՍf%�.�\J� ��'�E���Uo]Q�"�� ��i_�V�x�*Jv�h�� ��]��\����.8�H�&��@M��?!<�G�����~A�� _����y��]�C�Y���aw��&� 4n�9���mIO�P�F���j�/(Ԝ���?o $B�ߝ�xIll&Ҹ "�B�*� �L����4 �����O��y��UX&��� ��������aF�\��O��a� x�)m���h�����bX ~"�%�J&�w���`�P��,��_�8B��C>�GJ[r��� �~���3���z�{�4�x�N�'�J�����ԅ� ����� ��E��9���� ������W�<�?�p!��x��� ��DK_���� P��Ԑ|bHh���t����t�\�tx�q��  *7Ŭvd` �X����D����5� ��9�f�y; �b�jO�K��� A	��9�ow���N��x֝B�OM0�j&�����Ԁ�@���3��ӗPғf�Sb� O���P/���͜)������# =w��_]}�|5\{@b9Շ#����Gi�N���$_M$ ����HeG��$�;0U�J�2�p���<���l�2i�E��*H���,���u;�i|� ����=�dX���n����d1z�	߾y �bX��Y�Wh�&��4�(���hԙq ����x�PV�UL�� ����!0<��B|�P �L0L ���`e�m�֋��A��`�F)|��`��İ� ���
D_�X�|.[0­�� Ҋ�̩����Ϝ����}�-(����Hޖ�������������Sn�OHFl =$H/�9t���lGm��:\����
n@�5��Ρ��0+����їM��f2�GO�@���y �ve�ݔ���&���u�W��Ǭ�
� |y��������rt��o��^�_�	�.-�<��pQ����� ��XN�5�O֯��}���l6���S�"X��u2�8.��S$`��H�?�m �u;��`�i�-��\M$
+�@4�ـ��d� O�ʌ���� �ճ^�f�Dp�����]A������ )[��� ��R��917���-�Pq��&��Tx�"���h�����Un0�����D�,��:���@ �&	4���8���s֧r��H�~ׄ(_� 
���u�M*$�� �ق�-�%����t�;�ίq/$v� K���:���H�mB���oLp�7���`��z�� Z�pJ��:%�u����U��I� 8�N���V���t�����4 5��J� ��O���_t �<�Պ�L���v�>ρ�?���O�u͔xxF�	!Ђu�0	�`H%��,Jq �?]�1�ɀ�(x#�> �Q�C�� �E��dպD9� ���W���ޜ@�E	O��.,y8�x��$�FU�� ښ�^�d�u��@�O:�=�y�`�) �U� �V��zܿ!҉��1р�y�K��t J�E�Ǆ	C����Ϡ�W�_�H ��ϯ�@�,�0OK�݀#~D��
�������.X�� ��3�`��P�}b�]����رy
�U���	��������̚�\ԇ�@���� (-�Qҳ�t� ^� ̼�4_O�pvX5�҃�Lש\*`,� 7Z�0WO�����E�H/=�,�j���� !�;��}�	Mq�ՀL��r� N��E��K���(#�~���`�������q�=�L-���`�L�W�� Dԫ��^����M� �7 <� ���l0k�q^ 5�r(��� ������O����J��>��1���Z[��p���y���"ϧ�D|*.���ԯv~��r�����UX&�qd?�|z�P�&-$v�b�H�(��y���Ne�cJ�Ր�O�H�����U�L�׮D����p f�$!�P� O�����x*?_�?��2A3�/[`$y�z�r����B�(��NA�����DPа���h�q�@���4@�TZ��=� s�	a����Wb��Oy��/�lb�k�u	�� �ˊ�EpB�PL��O���3�4<� $�[��u!V�Zd��] �=�jA��� �p_���by� r�g֬ ����3�� ����r
����Op����h�D=�i� V���S'EH�` *�x���
?��� ����B��	��$�]��S�e�J��-����Qͪ�x, �hTR��O���םT�Ǡ0|q�� ��.ቕ�! O{ge�-��*�A��x� �D]�� Ӽ�����9�Eވ�#�����GҒyYӀ� ���2�]�L� ׌�v6�:�҅B���|�
-���5>/Կ��\? !l�b��O ������:ږ�0T^Ƹ�X�dp� ��3��;Oc
�=U�(������� ���u=�N�:��Ԧ�p|U��Y<��0�9�a� ������ %z���F'�ʠ�o�@�b%�K5_����( �w3��;X��҃��`�.�@�ϸU��;��Q?��O(3Ű)�`��RhE�eOL�8D������>������|���>j�RQ��Oρ�|߄DJ&x|	�io[�p��4Jqx�`�N�^w�$}�l ���,�@N<���� �]p�����S,�� �%�BǪ ���<�x$%Q ����g �Eȑ�˅ �@֭B_0�s��@\�;�a !�N�<�OH���ѝ�Ԃ�,%��D�O���N������9����򴂴�a0��`{\�vM �x���_��g� ��'�� �`��iO�h�R4��� ��t{ ���L��,hrHHq�W���O� r)QDB6�: c_�G֘��y�w�S�����_��ծ�y��Di�|`��U���'�P��&����:���NF ��`��ܐ� �kz�N��t>�� _O�J%��ձ5/���� >�~���Yq��y�ӭ_��P�� \GO�b�xB��վ����\�@ ��N����R8f ��Pyt��0 ��?j�7� �a����{��sl��఩�t�{��E�XO��hD9 ��gzZ��|%�.�ld��	{w4dV8�Ȃ:�Y��ς�zc����@ .��Ԯ�&(<~W�$�����<������H1t`�:� ��*q�����4 -�ëpF;yG�¬P0x7sO&�L ,ƙ�{@����h�|2���a�o�q���iD��}`V����sAk���N+� 6����� %<QÒE�: g5�rj�]�.�\�: '���N| b�dO��R�8��愫n��:�o �>PO��'D.8�`6m��j�$���
�>_A�x��) F3�iz�\��r�9��������e��N�?�`��qOp� �˖�� �/��Ո���y� �w����(��ՂlU��d7 �쓪���L>]	��p@��.�\(� DP��u����k��&� �s�R�idx�%�� ��mW� �Ȱ�cX�oJ� ���Eߒ�7��?�,ϣ;���=S�G6�����$��B�#O�0�Z@ Ll0����J�x`-��&�H��T|�BA�p�0�N��G/?<�����n���|X�P� ��f�8��E\j�# ���TԔ�FҪ���O�L�?J3�D_E���2�O���p�� 3Z��ΘV�%�~!x���!l��?[� �S�5J�d��'t��Em�� ��� �k��z����`����������9 �N���زH� �������4��0���� C&4����N ����ѹ�� ��+��V�xH�P'�h���.i�� Ԫ{�H�d�����A���p��JA�� ���S���Y��:����'y���>C`�pM�[f��D���10�*:�v ň�ِq�Ϩ�	O��_#��J��G��x��@�9��${�>Xҟ`�R�1Z�p�0��~[?ϲ�S�IY��b�-������A���� �H�y��P$����V6� şr��T�ؘ �$q}ղ�|��] P"^GA/Ͼ  ���: _9f��8�����Z�O,��!�;@�4��Ƹ(��y")��x��K�E������E� ��&����ғi��>��<� �3�Y۔M ���!��L�Վ 4�fu q-O<��Vi抳�?��h�0����<�Qy>�c 
�7�/�&*!��i�� G`��Rn�y� b|�vĨ �����B�� ?R��A�f�y�V��- Q�;NՀm �֤��� Y�)BČD�� �G'n@�
��N��pe����=4�� ��A:h;JCET�D�td���pwX�	�PN儌���qH�P'@����D_ ��h���)���� 5�+��"���|�$ӊ�w�D �������W�m��J�
�P@T�MOS� t��Y�^�?���� �3���N�a�Y�0s�3�o�eR����5{WyZ�UO�Ty�H�-�n%S	T�N�7�N�H Ma+ߦBk ���t�%�v�"�|M�L�j���J˲
���0LՆ��Sɨ��TyB 5�����"�� ���3l)p&� /��N2zO|� ���q������:����7x���؈���4�ZO���{8�^2�j�+�H�q(	�%r0��9�ҝ�0��k�v��� {͍�_%��H <� ����ܝ�����D�<ä6�,���
��� D��K8�d�u������+Sr�0E4�Լ�:@��� l���=����0o �\ҧ� N�T���) ���h�ߟ ��t������+� �a���� �e�x_v	P��W�L���
�,�l�x� ��r�b������� �-��E֐�J,�yp���� Nr �������d�� ��H��F��Vw-��R`�P 3Z���z�$+b� ��>�֗������.h�$>H2�>O�k ����0��ƌ������*|BrN(��� �f�Ɔ;(ʭ��,}��2j_=mfOXԜ��Q�r���N��d����%�P���Ovl֝W��qP����D��]�y�;�@�r� ��Tp�ҹ$ԍ����]�e�� ��F-j�0�4Hr]�\D����uԅ	��I�h�Ϫ��^9��3'��xw&�U�@�CQY��cO�A�`�r[�7��@0�w��,C�5O� T�EuՉwİ8�1qp��l��NTyBp(�T@��#����Iz���,�� AoD	�t�9��JTy|��1�s��dH�޿P8 ��B��^��tt`��m
���s �5m�4�t�T [��� k�ڇ�s�l|�4�tY;��ছ��-ՎcL��?&�ԭ e��:�0r��S�\H�4�0��;���֗�:8o�pD��|���D ��	PC�v �v��&�� �xu-��XF� Y<��y���|���[�9h�$�<p ,
�g�6�=e���y� �H= �Df���m��ta灓��>@l ���6���Ybxa�@l�d>���)���0�Y�<!���-�e���8g� �� ��W�
�7��΀,��D���@��y�����@piՓ���:gy�x�>��~tM�! #�C���AHaP=r�%���	 ��Mۘ��B��  վ{D���^ �,����� �`2O%��F �^��� ��_�<��$Rl5�&O���� �c�^�%���ɿ�øF�l�������n3G-6�`�� ��D�|px� � �O�L��4k������0N��m.�� F�/1��b[�)Aȣp������m�O�M%��h���X�H��$ĝ�yQ���]Fx�`�>��ŀ��dIt�S��hMŀ�A�F��TБ��G�l <E�����D���GW�6f��mN�h�I2Ih�N���0����`��*f�S���� ��_���D1k�=��<��xfî'�?M���z�,J�{ x����[j� ���?:O��Ĉ�^�$qk}�區˄Ӳ�O������8=�ԝ������� thN���6J�c��Qkt�_��b�$ ��4kJ�R���<�G �b� �Z&PL���8� ��N��Գsd��Ux��O� piϖ����DJ��8�FV$���m�ҿ�T\�(�F���(M+q�����>� lim�B��{�� u.-�p�����!0��/d��~� ���xq��	P�`Z�0!��$Ք0? {l��	��x ���7�qO|� }�o�C��/��<�&�8��E���]��X��H��%1hA!{|�p1N�xb�;ԙ ��L_X�Oa+(����z� �{yC����l� ��O���>�:w�| ;}?���H)r� |�w�Ab�~Oq��U;�N����_���ǝ��J����D�8�]�����"��j�O�'�<����#�}� ƤH����5hD�G�ِ�Ԙ �8�P[�?-ў����/�I�����ax:�����$T� L�*�8Q$4e�
V�����:ОN��o빻"����\O���XF� L��1�T��Q�!�I� ����<�$O�� r�Dӡ�/vo$���K[T���3 ���N�0���_������3�������zN����t�l&�[.V�y�������^�֘��u� ��,�:�� ���"�<���_Ow�+( : �W �/�[�ָ�H�4&�0 �]�7J�|
�薤� �EN?��&<���g�>!@lu���玤v�0'�d �I։?ߔ�ܫЃT%ːbM���2�­4�� ����� ��|x���2�T���h0�i�5�Q�0�C���J������N���u�\~(D����0Hz�� )y��/F`ֲ�ޠ{�+��M~���&���T ��y�<K��ܞXs�{�|���%@:�=f�,��p2�(��.�M�'�{W.��� �Q������td�(,�	PT�Ƽ
V0�<�'hJ������g�MTLd���V
ࠫ�`ܡj �ظr��z�,�)NJ���F��R_b��h��٤D q��P���?^�8Z �n�����!K�؟����DNA|J��� �vUͲ#Ճ\�( Ԕ��Z�O�x�W*���4�M}��0��D*@z[�� )8��"� �Nm���܎�����@�'|�+p���k 5�]�~���T��0��}�GM�)��� j�f����� �W���_���͐� ����u��h�3l��,��=,>%���	��Ed���b0��ԁsM�Orq#h�V����I�>L7�pd��t�[� �����"µ�0���nK}~�(��q��4D��䋂�&ϦR? ��n���� �+ʚE�,��� ��A� ,bu���8|���;�Կÿ�&��� F���7@�A+�@���?�?�Epz=	��@T��j�#``�:osu&�Ĵ��R'���=����g��:� ��+hO�Z �d���� ]r|o�kU��`��h& ��3�1|\ɴU�%�j�gv<��c�O�Ô�܉��j4� z���L-���M[�����:�^�NF�� �BEO�Z�,�Ҏ ���!ՠ���/|����t�L@PF�q3.A�nO��,R�s�	����EӺ�T�9��JU֧���\��n"�@$�I�	�_p�%�'pd@b �ۮ�3��i�ҹ4�bP~�\��_�x��,8��Y���d!�l"�U ������� x�z ��72�D���:���� k�J8���H��L�*@��MO��8����mͺZ����(�G����y�N� �~�'��`��x�d �.אOl�Hʀ��Ĩ.΀� �қ���<ѯH��۝�<6���2�X`:���*^+�\h !��ϼ��cnO �[G��￘� �%���~� �@��uP���WH��d�r��ڊ��Y�NXh�,���5����@�ރ O.Ea�є����9�I�NV	�5�����[ 2�R���w G/��F� ��U�,����L���H|��?@(��sA�r5 9�4n�$��� @��� ����c�Ϝ�G�@ئ[AL:a���oH��U�c,"Z`�8��D� �Y�h�����w��b�tPX���N 4C%$J� �.ycf��ظ@`�P�/,�9��	�Z}B��<\b��xO� �U�{�% �ǐ������՜��@OW�	�7�pkW� �ԙ�'H���I�����b QT,�J\\X��=� �����U ��ǼZSf�Lm� O�nj§�LB,>�(� o7��ST�hu`/8_|.� �Ӻ%ҋ��u� ����#�x� �9πU�\O�(�
��L%� ��yK-��ф�g�z"�`��4���H�@�Pr�-O�����s���P� ��3�^�� c�ֆ%Ϙ0HE�q�v�ɻ:�hw�ԧ��0�;���	8�<H|NAy�w��.]@o*��� ��l1 7�Q֊�
��璺 ������ud�����|��&`�l �׀�J6,c�dʩ  ���7�ϰ���С�W�D����{��-��ľyH�l �_/d
&=`�լ�i���0 eM�K�O���,�"�$�o�ĵb�O��0������ Bӎ=� P����Հ���
we�����a`��JX��9�� ����g%jBO� �L5ϢJ��`�:- �*4%� O ��TD���7$�0D S$�K�P����� �q=O/�
�>H�@VE� �p���/v� ��O��n� ��ԟ��ցR(� ��W�ݣ�.G�(���ȃ|�R}u�*z��A�� ��ğ��g@ ��
�L��Nu' ������ �>n��K͘�<$,@8:R0�d cZtO��m ����v���`L��L�&(-�ٱ�`�<D��ƀ�Y�R=����1◴pQ��@��� D�x��4|<�c ZB�AO��}���t�k:Vc���@L�B. �����9�*(�e�&�����V�jbt] ���;����@��>(��z�
�ǻ9s&%E,O���Y/} N�҂f�n�<0�.���/����@��&g �>�;�w-AH���%�����G��� Lv'6�p\�u0�kp% ����A����� �FI$ny ]�-�:̾�&�M/¼�]�T$ـ�I�6sy � ݔ-� ����H	��Kg ��B/����ǅ�(� ��Ld�% u&Ox �'Э�8�B0����Cr�9u� <Oׁ�2#�P X��X�ߛ|x�(e��Zp�_���F��d�W� �δ�����Zw��]i��h��ҕ���N��O��MU�ht��D����I�%w�X�� �s'��j�rS�@���z�����y'`L]6F��_�TT����B�Rw��� �	��1�'m���5���0j ��<�E�OL�hAw:�^������	(Q� "��&5��]��U���1o(A�!��jY�����N#��`@�r���e���� ���� t0��8�n� ^Ԏs��E���.����R� ��E�� ��Ü�(�$�=b��Êe�[7O <ϽF1ߋ5�? ��v|�>��0��D��`HR3��Q��1q$��1L�K �Ņ�G=����EMB'��z�`�+�x�b�F�yx�\�p(Z�O� �
�J� �xC�����69�V��J���'krp�[��	-�N`�� �i)=���(r�� 7`�S��� o�N����tp ^b�����+H�lȏh��O�z� �C*��>� I���l�՘� P�\H"��N‴��ڴ {���r`T�$����d��P}�8��q�K�T ��ʣ��Y��Cg�4���;ru9b�N�ј�	�2�$ �j�������Z^��ɨ0�U-����%�XL M���.H+�J�s��pi� ������XD�g��jvZ (2��[���� XK���5�%0�Xq�tBU�;�^'ҰJЀ��&�Ӑ�4� ��uIS-w���A� P�	�����@BN+)fT|��Xt�9���xB5�`����r����(�Ы���_�;um���Sy`�3�X�\	�utxa��S��l� N�>�/�;h��V�� t�� 5���^��i>�NL�	�T�jp���`��CX7*$M @��Jr��y%����o4
���~P��"DB��@�ꗀe
 mP��j�i��y�� ��Ԝg	�&��48>2>��t%�6��o�֒)�������A*��L�0%���p?�v�l��p>��	n&]@�͋��=� ��̢�1O`ʨ�:���� ����y<=�Uؘ�bQl)8J�$�e�:�'�"��W���Ϩq;�d�����P�(��J��PZ8��.D��,�A�@tp� �Ȋ��8�� ��>�� T��꓄~\��9 ,�l�?ޥ�&�l��	�ҀW�Jx�% ��> ����@,�pY;��֍	+���D��j��vk�����{ ��@ ��h'!�Ȑy�lt4����P_TW��{~ ��$�wc>õ@Q�3Ϣ	�NI�n��M�14m�u� �$$.R"��x����^��(ɟ,���� ��UO�`lI���k-���g@ ��= ��yb��CH��/� �����p� �{d��z <��Ծ� �܇���
q��� �#(P�y>^:+�ՠ�|MN9���0����� /�$%��,B����W{��IP[�_	R�.lK�F�P0 �ѭ���]9[- ��|��rq���T���4�H��AΘ؍�`c,P�ے4��k�8 Έ�q��ԝ��#A��*GX���<9��	�.$��,���]�{�'���<��LAL.T�� [�EQ�Ω�^�fV]~��*18�k+���H�ND |[�I�"���Z�@`��0d��H.�@y�� ��pO�n~N�Ę ��&��yZ갴l���G�4� $����st� ��~������N�TB����C �<�����m�g7T����ԸT�9b;�j͸�t<R�Dѿ����Y�2 �z�͛ ���Ǿ�a/kI�c��� � 5O��B��l� ��ç�-������_�������} �v !�i�O��n,|+'��O�(y�\M|	ܠo���N |����&/q�'D� ��t�%.�����H6ȍ�]�� c԰��H�� ��L�1C�+�,������=^�(p|� �y����ҝH�� jO���z�v W�®��x�����k5!OM �-��&� =�w����c ���">�[L	�2�Z���-�-��� J��\G�[yȀ_���-��H M�6�XD���~B2�GJ?t�`T5�9E�@N�����P��<�U�$�o!�Rpo*�h�R�#�҂�V0�����lGֈR�Ox�y��紀d�L)�
	��HtNI:��cV| s�R��U��Q���&Ix`/C��RsmNֲԗ��B��:(�L!O����r��m��j�d&�oh #���00��� ���4e)֞�����LՏ���c�� �E��:� �s��,�$L^�~�T� ��'OXtH ��dN_��9$ �2ؕ��}bV���
T�W ڰ�>=C��/ZF����7@�T����V���L3�H�	kׇX*���;�8/� M�����v�� p쓆���|�7��@)"�^�ZJ؀P�c�%��[r."~�ԨW��o ��uX�2L Ԟ���n�L��%Q���m�T�ʐ� [Kw�U��C�� �z �=�D���)�A���.������� ��"�O%Bx�w<v��@P�6�H@^��4 *3�ۨ�N_D� ;��N>�y� ��Le|9�\��ȗ�4J�E�C�8"�H;8J���"#�0�d=����-���>��c]��Np�U���2U�L� ��e!�2:J���Gήy��H2h!KO��$H�+'�F������o�x&-��$�lE�V˱�pI�/�p�~G��KHy��w�T�Ϝ �XM��,0"x��y ���E�/ r8��-L|�8`��������B�!p��|7��ȞU����LY5�L{�=��#.�<�!χ���E�0t���9�Y�0��±�v�=(wֻ84X�P�x��@9h��0:��=M� ��,���/�9Ң)�ĭPb��,6�	���x��������~�b4���@�Ӳ:$r��-�yh���f]P�	 ��������;Q���� }F��	kjz�l�C9;	D��<�# �u�DO}� �G	�� %�MeN��O�V�
b��&� �)u�-U �Ŵ���C��h��
�Z��,� �w�ܥ�i�%r Myvx{R��E$�#�����'z�A�}PT"�[��	�f�l �L�X��BE?�	���  �%m�.�]V���Ʊq��=w	��0:�z��<ؗ�Q�] \���C }�s��I�f,J�@���%�p0�!��I�D� Jf��R8�	�[�T� �6��S	�3o� 0����s0 DxX�� ��6��H�8&��h�nl ��Y���Pä���|T�x� �O�󆰝 �Z�t+�T�X*0��C���do�~� �V�	�X^J��Լ�0����
xh�(�n�?��5�SO�J���9�����y:�| ,���b�;O��n��j��87� a$�J m����Z�~� 7��P��j|wF!��%o�`0\� :��F�Ы��O8��N��ƹ���w����Ƌ�Ù��AĒ�` �[ɲPӸ@H�0⯿���M��6�Ԩ^��X>�ȃ��2?�Nk´� 8f�n�$�H/��	�%�u[E�H3����l��x�X�x"w~� ,�d�
tyLx�|� �	N�PtY �
�`�[.D�F��UZg��  4�Q��PxSjC���g�{��=�� T�n��@Q����p�T�[��� 1�qVZڨ� ״;�RL��a8횜�KY�p1� �_��6�y´A3ܵX��,c[
���� T$��6p ���e/ �[^��6�� AZ�T�� -�R�]�}^ ��	[�i�2�\Z^� ���� FK?[�ъzW�;�e�Է�%C�E��\��d��R����_�z����g�@�"Ar '
��Rr�� ��D��6�� MZG̀Tm� ��.��;!�����q�[p� Y�%�T� ˫5�K��� X��]LE\ �[�ʘ�+�x�w	 �����v�H2/�w��==U ���z�R�[�� 8�J��2E� �\U��[6_��� lu���R�k �O���ń /KV�o�� ��[�32Qi �K��RO��$
N��Z�w ;G�[LK��ulc�<Xy ��@+��������[��K��"�Pq��Ie���d��	(��� 4�Ɏ� k���T��O|���� ��[� �)Zm���8qЀ�[��8
u�Ĩ F1߱YZȑ�p(�G�*H�41�:�5еH� ���'Z�u���;�RV@�U�� 
K9��*~��(Za]{?04}Vdpx��@�y+�-$�Ȅ4�0��(9��R���Y`*_�tԵ`�Z� IW�1k@��R � ��;� l��Qf^�LZHy���%�#�!�5�9?� �I���[�$+yt k1S��U&�T}�`9"��QZrb��x�������܀P�k:x3p| _��[O������>P� 4a ��+K6Aw� ��0TZOռ fp����HMl��EF'e"�[=�0Q�U��B���������RY@d +oT�Յ���" >��&���5��\nT��z/�z�����r_$���]� 0��Wv���{索 p��#M(��,;Q(=� FjR0�� ��OKZc^,�@X �f�0-��dx� �nv��[|:i h`�����R�̾����Q|��H�p8������m� X�7A� ���`�h�[�o �{:�s�:�� F�=��Y�x�ȴ��Ti� +f�3� 6��8_p�5��, D��1T� ��+j�օ�OL� 6�M�zv��j���: ?��`<�Ơ�����DΟ,{��
��;k�`�x��$K�l$� ��F��M�_TmP�ӬR��	 �<����t���"Ā�$uZ �����*אd1ꂨ����[VI�����OH��g-G����P)�3����sh�m�0���e$����1Rq@�DdP��檙�P�@�H����F�) 1��\i�9wN��ɀ\ZAy ^*-������ 3�m�~ �y�
�%� ��9��mP�{pF��!��;s"��;p㈽��@wr�`!mI {
S�����Hm�G�X�Մ��Y�(m�s3	���@�4&^m=�N��A;��mB94��q����bume <��M� �� ����=����PL 0��\F����VX�qpځ����]�"���>8��@����@���]����y��� �8�x Z�D���T����xl�@XpT�@�P���j\f�&-��a>�����@O�~Z@�H���89V6�AD�j�T~� ��&�MY�� @��Q��/_����+�͔��`-����A����$���HI�6��2o `!����9�bl� !UQ,$G:V4��! tX�D���:8p��XA�'�?6���h���� g}��
b� |X��)Hй ኀ&"�d(=-�.���E ���� �R�������D� 5�ڱ;�� 9:�RK.ь��Vt�= ��]�6�۱�GwŔ� ��rX��|j aJ�Ӽ��6Z��ܤ@�})`Y���Bt|U��a plg��00ո�� �,^�V$�F�A�+����O� �,��M(ر\=�N�nf~�h� @�X����t %K^QFPAUVR���������8L�| A˚HwZ��bO�\�0� *������!�ڎP@�Y�����T@�uz��X@k���ZP�| ����z֦���V��A��,�;��G�0�8 �>o�L��`��RAg�`�ł�����a��!t�t<}�1�6	#L�`�?�P(
�
��.V���� ٚ���H&h� �}�Ǒ�" ߝ�G�]���# ���'V�g[�h0�3P�Ȳ�V ��T�� a;��_S��|mP�Q�(�Cxf��W�7��L�]�'�`��޻l����E|��F@��x}��N�� ��܊\��H6d�f�����X�ٲS��>��3� 17��g ?�]R�` �ؠ���9j߀vwMx��.a� �c�; g��iP� H5Q��9� r\3슘�siU ��q,B8� 3��� ��gs(>��xb N<�cp�� x�gM�sW u�a&#�ȕ�? _]��Zp� 3�	�@��{ �C��=��ݐ:<p Ocu�����. ��w: v߹	���8����S��*"t��nA{`�u(��� 0��<�w�� ��)��� ��!_�5�M C0�� ��.疜��x� �z�iI��x����p���_k�U8�D]�&��@�$�%�ɂ �|���0 -����� ���/�� �u7�@�Ε�n8 �c��^��57�8\ʆA��܅i 3�ha���wo��\V��	}� ��r�@K�<��D4� :��ى�~���l�֚z��� Fu3d �(D�������,�N��[�(�<�z-f���X@��� (�pm�>A���V�w�`��2�qQvA��� `��� �:)�|�~ �7��%� ����g^�x���~\瘒��$�� GBp-�`l�4���7��2���? R�^ f�������6�LJ ��Y�%�N ����8ϴe���sA�<8	 \�F�Y^�Mzĸ�����d���@�h�F�4(���Lc _��ɲq �o<>�r�� @|���^��  X�4�x� 7t���'��{��	S�� lMf�X��{ (��g�0I m�̅��� O�D��vT����*�^`B�m��cM��g �W�aF�rA8�@��p8� �7>��/I|,��| 5��\!��+^@G�۱��}'r (��vb�n� ��U�ΨމM�� �5ц�A�  �x=��Ou�О<K�8� n j�|G�N���O��S�� ��k15��6�:^�`��E�
 !�W��Fu~ /���ω�1r� _%4���Iu� �5]H6�S� 3q�omC� )�_P��<�Ρ�UI!�ð�E&s� ek�Q�d,7$H+�`��kt� 6ɕ�@��*}���� W)�B��\�|���� l���[ �5^�A�։V�LDԨ�<�*i��:k� �ھP�&�� ��
BaX�	 4k����ۀP��J I���5	�>�q�V .w�l����� 'ȉp�^���������0Ո��]	��,�\�7z tM��U`O�<F�A �!�m��D\�a p@�\}�y M=x�;�(9����@L�Dc�� C���#� ӕ�l^��;��&�R(�8�S�Ђ������~,��� ��H�Q�?:�a �%Fb_�Xs� .���i逰��w05' ���>( �:c���h� ��QP�$��� R�\��<�#���8���`^+3'��Їq��C�R`�]X3� ��^F�!=zZ���jc.��� �u�)ˀ,�� ���]}�� @=�RK�F�>e����t0�2�d�  p��r=��	#���,�j@���b]�`*��[������ �ؑ�?]J6���d�� ���* �A�1�듐,@P6.W�2�\�
 3;ώ#�^.��v����Iq?,�Й�x;E �-��x @)���C�$�l � ������oƉ�Op@��?^�Q:ކ���8��� ���7���=� FAN�Y�c�14 �Ϭ���k�^� �8�{��+���n��e��� QOF	� �X@���iq_���{W�7�Q��Lp|P� �A��dU��0(�v��,��@J��Y�u�c�Е�KLk�=;�	v�D��በ�9~0�Lt�<� `3��}L�RqA�� �+���� J�]�L� 蜺�ĆX_v �V�F>=���Da�4�y�8��4�0w8��}9��_:�l��Tp	 �����E� P�9<u��|�N?�82��P�_�a8^
���S�|�y'7� R���>��oa�^����5/�89�
�eY%��+�@�~t�˘��#�y��?\���;�N��K� `[�]� ��y���&� g�?��e��	 ���>9�ϻ�� y��u�^{�O)�*l ��%Qd����hA�0�2s U����웘��g�� �� +���S�w��蕇����������h��4(�r�;.��_}q�
�@�v�� p`5,}-	I���j�&B ���#F�^��� EK���0]�P�s�YA�Gd�,�g��:� �NeU�Y{6�R��}A�`^Z+q#������d)��`d|{����'�lve�� o�,a�����.�<�c����㱹��:�� \�S�D�� ���h㓔ٕ��_!l�f L�74φp��N F�S���>��\��H�ʐ	$	^�Bh<<Z%�S��U�hИ��XK���Վ :��\Ġ��X�$�v �f�F�� �G�_��	:�v�da�.�wu� ���fi?
��Y�� 9�\ = �y84c���`nP�M]@�N;�Xż �(o���h���7��= ����݉:#�9�ܿ���[h��㖡�! K>�x�Vc���ug ��,�	�M���Tڰ�:$mqP����ZQ �nFXE��K �ƕsp��H�`����C��cM�H���;����`dV|� �o_RFW�� �=m����<v���u`�R�G��>�Q���H	��? 8��Ն�@ȧ�\dӉ=��@�2 ZKg`3����X�ՀEya+���XO }$v�
!����%r��\� �����L�V������+���0�G>-���q����>�8�р�<H�I9G �6��wٗ?y���o�W �#���Y��z\���(� k�V^
N�d�s t�$0�8?_� ��1!+SM�,�H L#_���W�Rc���m����SA^���.� +`��U�=�.��s�H�	� 6�<�̳���:~����_�I`�0�Љ ��~z��� ���<ڕ� �ʉ���^O� L=�q~� ��)��~; �,�i����G���#�(���ޕyr�@P�S[z�(pt�\i�T�G0Y���x�8 떛~��=�\��!`�`U��'K��}pX�XPT u��W�5B�i�\|l` �#(�Ǒ��qf^�U02n ɉ���u���B\ �
�o�J�A`��� �R�0���'��	�b�������A���<p!��wG`6T�Ҁ@�=F%������qA<'� "n�� �#,T�` ���q�SR<҉Q��$/:Vj
��Z���7E�[.6����`��q�����+g`2ѐ�V�78H�%L�a 
?�\���ӕ`K�@�CІL}�A� TK���� -�D�ust����V & ��<l�B�9� L��������N��
����1�w
�����	A��lΧI��$����^)��/��ie� lf����5� �Co=�j]�xW p�;d&��$^:]��É��ex�(�� �6`�ZX8�9Ɇ��@ ^ �U���L�E��H5��Y���b>2����!~�|tH�,@�.-^�C��)��:�;s 5�����\�0:̖	� O�[<�lF��� �X�K�!_�ea=��@���w ��(�<C4R˕�'���ծL�,�F&?� �@�
(�P ϕ�Ba����&��� ��;�IJ�1T���&}� ��F�a/ �f�@6�7w��!���h{.P�Y_Hw� &�>�.��A�Pz��N�W/5_ �S��.� ��oH���B}��C�V~`ApNL�3�Y���UI(;!Y�"�<^��,H�>T/!^�J#���f���Z��� }��<�E&s�����0��w��_��U>@W��V�+ ��y���A�p� 7N���K�X��B�D�AԀ@ xT)�#5���[�;YA;�&B:p��)J�`��� �����ھ�~!	)P��9}o �z�>pS�`](�:':�~�B? (�չ^T���� |+a���}�a������Faԗ���w�б)=V����r#Ԍ�����,��#`�aA_�`�7�:�� �d��| ?�FG�f�L��w1 a�c�� A!N	Ez2㉾��}x�\��0�6�� (>�i�*���6.�x�B��@�$10��8J� Sl�P�D$~�0 �(�
�=4E`������y� ��?����V{k_�	}� tz���	����� Æ�H�� j(�7�q���|* �<�k|a�t���_������ *��ũ� @uv��Z�� �Oyѕhm �ڣ[Y��鰲<��.On)���@R�ۄ����8� _�t7F�i� E��] �CK�k��t�� W�G#��Bu|L ���h$׳�o���?`kԸ���DRe��.�� �A�_���@yiLۻx�@(ύ����¶��1� �d+�'����LQ	 ����Tk(;���E�D���f{[J ��kpّ�<���@�Ldv�c��_��[գ|����L �g�e5u@k�� �<��Կ 3�(�Z8��� �N�s2����,���< �g����"�������	�_����@4��� -B�|y]с ��n�9<�� 7��׷+I �x�/K]t2p�>F΀���� ��INP�6l�%W�B�y� u\k���V��䷴U� ����` 4��M�fs 㚓\�r� u���^��� �R��,4i���#��� A�_����8��tk��@���r�0����#�8� e�"�rb M����� ��w��un�Y �7��ۧ�E�Ǵ>�����}f %9kV�}3��_շ`l��� ���=� �����'t �ۀ]c� �&:
D�� H�!Kk�<������������;Hf8���� �e�w��-�|���@ ��Ҹ] k����1��c>�q0`V��� ы��6k�	3Mn����5@�Df�l�iy�ҋ���������` $؃&(M��< r����:C�K��$�����V`p���̍��B�b�*"�y�D1'���A�Ok�R1$4w�W�8������5ɩ~� f�O�<P�=��V=$�����퀨����Y� ȇ��(��� ��}���4[���V�L����7+ i��s0��9 �Men�,�S���‑�0����%�LT��!�b���i� ��涠�9Jt�$'�\��0f`�	 �k���T]� �0o� �����e�~~;RlH� 8Y�4��{v2�����; &���k�^����0	����*��㮀�� <X�� ~T����R��Ԛ ������ ���u���0�����{�r\� ����V�z��h���d�9��iH��t% t�S�����$����4�!��6�>&t)��� �l����S��� �~)A���W�?���y�Y,��\
C��X`TH( ˬ7o< l���ۊ�@���ӯ?j� }�Ԇ��LZ,�� ���J�}� ����B�j/��
�� b�ud�v����R5�X�s �r2�\W��-t�!�����4�/����}�F�R��1�+aLB�6��w鐈��U?XA��. ���B Y��Lw;�9cW.�Xr��|< ��kY{��pZ fr)c��] �[/WX@�� S��3p7a��[�Q�����k�\�`��ܠ� ij!�c�.Z��'|���Ѝ�ra�YT �W��Z?U� ��m^���`������)O �Z؝>9`0nV(R�Y����&��S����})�f��LӢȀ��6pPKA)P4a�a~�y�%B=Ǽ G���ȿ# ��N��T�,)�r��Maқ= �ׁƎ��(�*,fp�]�g ����� v����:��0tUO����fb��\װ���{#�|2 ��ކ��d 3������ �*������P�G!�v}�(�Ej������ �}s~�T#�b�{J8��ƥaRAW4��6�o! �{��9����AԬl��aiM`�z�;�`��J��� ��sl��{�ޤ6R� z=W�;�*8@ u�"��Khtc��g������� 4So�� K5��C����'�ni����?H���5;��@0�k0�� ���J^��� 7��5�E�q���j����N�{dm��O�S����$��[&��FЀ5�N����ڕ ��f8�T���/_
{�$��8B�?��W�����\�� ��a�S����f�֭�9m ��G��4NF����O��$��90���=׮|�BX�<mP�Y��q����$G�]3�l��ğ��C�H�o�B �[���{��Dr8	��� X�dLl��{�ŕ \S)n^�4t�"@Q��(x�lZq� ��0�~i�5h�P��eD���{�ń��6C��4!���o�B�F2�5(�@�?2	|�a:�� X!���� �'�)������T��Hl���b�Y `�_��'Qh�=� ��,Cʯo�5V\P/�m@�qq2>t!���n?��������9[���O'(�a��4�ST�P�l �`$�$��@��u�k�lԨH�������(v�$���(���P��iHI����S�dh<<��������� � �`�-Q@�  �d� ]�F���=~�I������	��@�%���_�g�q��c��$x6���`���I ��S'� %�C\�#�d;
+6�D���$y|�Ao�%$�2���C�ko	¤��  �h4|t�܀=���
Y��l�a2�� ��D��\o ��0H��*��<2(�$̉��B�j�ǅ�I��/��X44�A`p<�O��i#�������| �a ���o��[㜚P�cBU����D2,x����H�|2A0� 48x �Z��)5�� ĭ��lkq�X���Q� �c���,� Q<b���:z5�%*Ɛ��_�� 3-�f�@qML0�:If��w ���(�TA�W\�1}0�44Bүbd8Z���R�$hI�R �}i�4�@�f�A٘ zm���7u�(�c�\Qb���Z�g�����A�0@��@���I�}(�	���2a��$Б�IQ08�{��Jv${x�@uM
�4�I� (r�u]�����`t���K�p(o
�H4�5cʻ)D�D��"�3h �(	k���\Ru
H���O� ���]�$�!���ۀ���9�&dh��t��3lU�R�HPg�OH�Qd"d���s4��9�od�;R\ ��V*����|m�w����q�H��SJ�A�`������Dz�}P�l��g����܋_\��)]�S��g��Bm1G�iJ�� Y%Rg�T���������@��}���X 05g\$S��{hO���t��cE0�6Tu@,/\@�W�x͹�BI�+������P�j4S�z�f���dא,��$��b��`��S8�IXj� T�yx$H���S ��<�J��T���*�1b�A`-�ƍ%8���d9����tq�����WL��c[��I��X���+@��3h�_ρ��foP S[���g�=1(�P�5-����#c�ؤK?�L��a̘�Fd!(b=@0 Z-(�!���`Q��������F�� �P��s��z*A�BNq�ܽ��? {�b_��l�᥋��j�	�R�� L��Q��8f�k8�����2[�$q��� �?�%��բ��_�R�ss�S4D��=��,��b��ϸ��� Wj$�|Nb08�� _�h�X�Ā]�$͔T���%Yh����p�!��R��+N�o �<��(��
�� Ke-�{��
���d�`�JH�|T�g��t�%@�k���=�xWd����@�4\%c��� ݰsrYU�#�F�Z/1ħ��%�6�Jb �֙+��4Ff$: ��}�3��r`0��h��\�l46T��`J�m~�s�f�,�	��"DQ�k� �$�1: �[:ʩ�P n�X���>א�� ��{�˱� �b��J	� .����Zsr B�t��Iy� )���j� ���/7saq����nXI��{`�� ��|nF���@T�))b�0D�@�3�O�a�� �Y�G D���A��#a��b�M��u ��Fn��rgxt���C�shp�q� -���*sKzt�Y��W�PM�� ;0
��n�лV��0q���*�(���G�c��,�����A
6���X�}�[y3���~��=�B>4�6P� �� xT� #S �qB-�g=Z*����x9�( ���ʓV��*�v�<�� �[b5X� �"�֧��I���0}1�P�� g��:L�� �ɯn�(<� RQ)�2��`�I����*�q�,Y�X�� ;+��o�H)Ihr����I���Π��V� 6ԲѝN} 5T���B~�Z|�Vr���%7 \�P@�+��t�T���Zd�t� X0M�x��(ݠ�q|oр=5���0�ݹ�.W !����b�4|�zM7�Ҟ@� �R����9 ��7_�,� ��Y�c��vy����B�:�� )���e��}9`	!6���ئ���&/ E|BKϥ�6jwp89��GC$	� �ۢ�����|�g ����nT�q�vQa$ �c� m�?`�e��asx8�;քt�`=�E#d�:������|����)��~� +�k4����es!5� n�+���(�����x6�� ��VU_�w z!5���y����������?ֽۀp|�9.��i��X 7#5*�^�_� ��t�S��U�b�&�0�Y��Ȝ� �� �G4:�m��X�Ho�� �،D�� � 4���So �p�Jd&2 �)��޴�-�Y=jDz�b�05�}&|���U���8����:�I_0	�!a%���|�^�xk�j]Ʀ ��~�Bi� ��S��tG���/��h�X����3���/��M<�W-�T��D Ÿ�6��lq:,f����&Ʈu� ՘����6 ;d��а��gP���`��| m1���}�acHkA ^��q�@70q���;����� �a���n�0@��`� yw��塇0��8@�) �/�\l�n�����&��a ��J��,�Ŝe��:��`��o!��p��� '�3���z�WI�0/A ��FT�d �	�^9�Q��� 8~L�6�4�8,D ��Kh�8���rT]�g"���@gsy��ٕH�b\���h�J�iz@�kT�*��?�c�� �����[A�< �|�*Ѥ QYz�H � �!Ջ��� S��=�s� �����u�П" �D�'r�21�[:� f�3���NH2�ԫ�	�\O���|�;Ò���uڐ��7�L���&� ,�"I�w6r����Y��a���%S;��� 5#��̄&n<|� �r�>�0 4�}�	U
,8���'�cx���|��`\�<�u ��34�0�$���d��r���"Tw�+���J�R�	�]���8�ߤ�x �v�R���� �m���`9��&z$��|S(�r��pH#ls���� ��O?���| ��5�[��7�2\�?t�� I�Lo��+r�0�ڤ�8>�@��?D�>s$ �R��W� �;Hry0N eS��U��3 �^�Fw߼�|7 O�	�1E~c�;��r��u��� |�w�+��K r��y�t?hZ �7�6�T �4���|{ ���2�m� �Ul˘7P�\�Hb�Y�5!R� *kI�\�H<܀���Č�k �4�|n��zI�d�E�U�O� ��|� l��G#� �,�;�� E�rN���s��2T�[V��X���8��p :v���w�9 �r!�*��x. ��@R�{�� HZ��ł���_�� +5�r�]�J%�T��;�� �����Av��T��@�*$�l< Q���|��( T�rO�}oZ�|�IAs�Np�f���vD��|z�Ư�Ì,��E <>@��U��0�;� r)������ w����.�8f �d4L�U����e��|�3��~�`����0ز	�4�.��� �|�IC	��r�L�>t	]R�m��ʍ*��r�Wp}�e�p��;�SK	��B�XM��rJg
��sո����	@�V��S+�@�|r��$�W�4� �aP_Ĥ@Z?�q��˩��}L�2:�8��Vfh�`�`�S��mHK� ��4�pd�eR)N� �52 v������ ��%�>´�Ӝ�4ø���s�˸� ����UW�����s��z *3-%HbM������\hL$4	&u�׀��r�ȏR �����~����`v����Ŏ	hy��R�HG��d��:q� ��7��vϘ� v+��ߏ�~L8�:���(���Zr��|>7� 2��!�H,�^H c?��r	���<I`��pB8����4��Rs�������|~ɠ��d �P���[��,	$ tJ'\�" M3�a�r�z�M�̳�w�G���R}���ߍ����"l������À��@�\p� ���U��cl�t��� ��Ks�0$iVu�:�l5�
����"��4q�L���iň `r��b��E��S���@�Q��U)^���|�= ��#����9�h�)U dr�6t<�
5s{���F�F`'�	�s��	� �[��qB>�M(� ����I� �)�ګu�|.U�dȀ8i*Ә�I"�tO` D����r*S8�̤����� =6����0�}p��3 f�/UqH�F"�a(�=$� �_Er��]�fϢ��@ȢP �n�>Xrtz��{G�xa���2	]E�� @���Q������S8��g¥85��� ]���:���Ez\�B#r�� P�������`�i-�����V��m�� �:�n��R� ����5�%��4��h�}���|/�q�v�U��64@`d�t�� u��yAљ ���+i~E�Mw ƃ̘_ ���s/ܤC��q� *� �,S�L .�T�V�?���r;+��B� <-��� ��9*�7kn�Ô�8r��� c�m�q�D>w���S���|rX-�9� t�L�DY�� ��?T�&Z�Wo1�����%$��ܵ|@�G�t}&T�b1�� �<�Bݧjã�k�70�X?P���,��0��Tsg�� XC����m`��v$���� >r@�5�ك��/D����x� &���}�:Rm4�Z`�Q/���9,@���Kc�x�|M�F�z2�o��f�#P��X7*1J�Q����S�p �o���=���~�4� �ci�.	E�B �!�! ɊGt�h� �W��	�g����$���| ��)a�st+އƄ  �)�2"{�c���P�T'�q�@1 �䏧G�nd�i�'�v���`D�1\������
������� ����ˊrTz����$v2 k��1��P>�5�!�z:#
`_]��:`!����ٮ� r�7��_���zp�0@��-�����k�_ ��Wi' �=��/����̲Z˵�e9����(RH ^�`
�7"�~4 �񛼺#���Yx	~�gW�?�-`�`�`˰F�����]ıy�!�jV�n���C�B��������Ŀ5� �4�9��8�|��\_ ����,X�����[��0{�@ćF�u/�����\A.�&���`?�g��/s�Jf)<ɘ �*���p� ��:]��=����r0�e�K�� /Eu֗�ȭL�������V� 6�/ӳ��5q� �G��4��{ �����] �'�dV�/m�.@斧� *���b�/ ڒ;ļ� �B�lJ�V�_ C�U�Ȧ�'�(���w�x�t�X PV�(���u����;X���d/0�C�|��� �֟�R��s* i�L/o�9���@2�VC� ���ʯ���0��n�:x7zi�1��"������ k9�/�'D��<8*<�x���=��{u@6� G:�-���Sw�k/���T���� <M��\�J  �%/�N��l�H�������^�� �ƻ_/�$�ųt {x069������"��+�"�)�`�o�p/�z� 0��$ A��ۙ� ���.�� /��y ������D ��Hb���5 ~��=��/"kV�������� ���ɭ���/05N������T$R� �h>�� O�)���+/q���X�D��*����{12Cc Df!k �/m��P %.�3a ��錴ă@��ip��/0�n��* Ό�N��0���- �`:t6���:�[�����p$߁��< h��9Q"�VU.ڠ� ��AS�v�x�Hh�$#l	Ƈ�0��� Q���l�- Zɚ�߫�! ƌ��5�/ �AMlx�V? _3�W�Ȯb$�%H��&a�-��A�8��Z܀\�5� D��k-�90��� d�Ve
�����˖�����3�/n���������� �(�� ��a�<r�;G�V@� ,2�\�^� ��.���
 ��{��߈�/�	�> �����`�RΦ6(D/ٓ�УH���,��@ ��iɮ�p����I"1!�Q0��>Ϟ��*��us��d#j�9� �C0��/6�9 = Z����  i�vn��}X	��S5 �o���������	� �NT9�Q_�T� �qȯ� g���2���<y� $u}ަ�p�ܐt��.n��Ƞ>=� ��D�Vu/J�^�Y@d<�˃�{����2�\Tb�/]��m �|���1����� <��d5/�aT ˆ��j�X��Ly���3p��/,�ޤ	w ����= �y�]�J7 Ű��`���,��/���Q�X�	��{��Ζ ���\���� o/����[��}`�J�g����/x���eu"�	_����� ������	�KŤ�h_1�� �>��+˼�`��!%;�9h#���l1wĪ�i�G�{՘0 �E�WT`� ǌ/;t4G�,��^@��ܴ `�����&ư� d_��^�5G �\�I
g�x.D��e����%H����h �r���� �.X�Н��u 'ȍ�_"��`)i�4�J� �2��j����"Lp���	�ݒxǔ��`p`MU��� ,n ��\DG :�a�,;l��� .�Q{ Z>Y|��P?mS�1�(k ]e:�I�3,x
 ?�ۤ2� ��E�J$O�����ɍI�� �J�| ��W���(K�A��`F���=`�I��'w ܠ�Je�n3 ߮�N��=c#1C���z F�ݚg/E�'�+�4�t�nJÄ�ڳB����=�YS������X�z㒀��>���.)i� �G�q�#$w��U����Y�A�����bu� �ߪG!:�@�F,ۮ ��CX$�`f� � �15�� �w�gC�_�uc�������>��͞@٘�Xef�HB� xW�� ӬN��"Q�E�~`��nxu�`�hv\���p(0A�!���TC� �iyF��L>0����{�fh��iR�l��q�H�1}~���`���P��zh��E�w0�4YC�c���w�h	������iq|��(��w#�'�rkD~���4"\���u Y�AP�{(z�d���Қ]f�� 
I����	�Ѩw����9 ��n@�YI�*2.1ހ!b~u�r�xp�Q%=���������W�����r���9� [�W�g�~  b�.}��0)�0S~��0����CU �X�Q).
�8 }��m��O��VԠ��% 5
H�4����/ �:{;*vt, � �-�^��	�WD����J, t�4K2��� 9 ��r��J Gj32
*� i����N�^7���- �f��]��M��u������s�Le�l��=�Ԁ�h"�é�|7z�g�vQ��kl>�Zɇإ�� ~%$�gw�� ��&�,�3@��� Wh��2"pB��H��:� ��- �óZgxS
�@�w�˸�v ��NKx0� E7��|M ���x&��N%6��Z�-�|�O���#����y| ���\�! �_}��B�L� ����� #!����s� 2)�3��I��� lg�"��u0���@j@�.�� �ҳ��� �K�'�lZ *�Ȗ�mo r�~$_y ?�L�����G�p8��� st�FN+O �V2~3��! w<�*�;n ʞ��{QxF ���@4�'���/ �t��2���@Z���s �xU]<�[ %nM`P� H�÷�!Z6��<� -v�L8� �\9 ~���� ��C'/�+ ���<��B� V�sOi@+� wM��>J~� ���[<�' �G�о#43`lx@�.wW�!�Tn�'/l@�q�#>9~�ĕ�zM	�\��`p�^̬ )��(4S" ����x��L 1 ���<���$3���DB�)%�6�	��_o� y�|@w� (�;�&�R?�� 9�.fi�����b��������L��-��o�E<� ������ L�p9.`L��_^��-j�	 lLU���]�g��8 ��_M�p `c
W��A K�1��p�fH����0 <+��?' V!@K�Z� u�$R��_ �]�Y�p禃�B�,  1�퉮@C0w9d ry�Ol�$����L�A�M�(f�� ��$���suI x�	�[yM r�"CqS60 �i!�'ܥ �\uvs(w��UqM���.�� ��E'j� |��rD�� 5��Lt�w� ~��(�fs�AX ���>M���. ���z|���5; u"8,�� �\h�x�tM	�0���
��Aw���fL v�7���j�i��ܒЂ� 
؈��l�#^��B�U���� �	"�}��-q�&c�' Ck�x`�FE��_�p=N'� i�XmcH�� :�"	�� y�' H˷ }���� l"Fp�N(q���w�[B�`;�,"Ϭ@̤L z�>T��	��g��j @&~�l; �L�Wa.M��O�'׹n�0�y8w�R�M�2GKZ!� q"n��\�\�o���4~'��M#{`0)(��cW�x;E����lT��ށYi�����P���p��o* ������� .�'mas��L�����`�`N@�I��&�@�!�.0 ���-~$lp ��@ki�Q �S�O�L�� ��.|[��� �G�i
`6�, �- Rz��� B��'o� hc��l��% i�#F|_��<?w��h� ��D�/���y! i�$V^�(Ww7 �ր��k� �oB�Wl ���!��� �J`�-� �Ul(Z~@� .�����A��'p��-B;���8Ϋ"��s#� ^%	�,���?z�!l�o��$� L���_��� g'��A� �yܙ!WS ���.k� D��8�Z�H�� ň~�M}�X��=�� ޅ/�w .3
Ҭ� ��hym�l�E~ hG���� ��o��D �q�'��� �6�Gz�LR|B_Y����� F{� �wX"��� lZBL`�#R8®�0��<%���ݭ,"p ��.@EĠ7:����'� �Z?y�/g ���l~i� U>�^w5��0h�F��'`�`"h�V�L���\���>`���1`��U�0 hV��]���6$�s��J���e;�c ӗ)˧�L ��%�p�X�H �V�^2'�"�kDKC\�g ���&;�pSp�8�e.9ve���x�02���˰"'>� ܒn׿y��4�`��`� ����&@6��S cֿ�	� !��B��� `�◾�-%���CH�i# ���qp�\< F�R"�saųB�L��$�[7l6�) �' �<�p:� �Y���L�J�? ;��!tP������v�.TA���ǟ�[�uw�L.��ʃc�])�"A�
qa�S9�G-�k0� �ql���\�8ޯ�N�^ |,q�p� w��մ��&LT�X�5�9ܘpz#��l���\���"�h �1��>�%� �8U :��� �5r�_��K	$&�!�@��緀8��,�n� B7_t�p�� c��'s�*?� �\��&�L�� ��c2�T�.���-� �#� ��wΨ wl	X�+z�9�sp� O���0 ���.<��f�Aȋ� ��'� ���&�c~�� ����Z�%� �M��y &G��Ek '��.`l C�
t�L�����il�`��~4����*�`8;�\YdPdi�Fw&����!V��� z�MY牍�'�$�D�l�+�(	�bqqMS 4g x�㱎� �����x���pM���|ݣ �K�x'���7�0� luvMn���	i!���8��������x�J�g�p������ �,�s=��A؉Eo���ugH�48��9�V�i$�.� ��P	m �qR�u�L?˷����C�|�='��[@�� FA��l��1�s��h�;HƈP� S0Uɨ ���L���NWM���¨��оq�=^�@\~K��?�� �oA����(�����U"C�a!4�?iz\��XR��� /=A'L� z�_�k{߸� R��H~��3� ]<�'vpI� �lˣJ�x��Li���d�b3�Cl�������_ LY�ܿ :Ȣ!�^�� JH�`o/��� \ZW~�$ .cE4���ǧ����t�R.��<hL Lr�Oԙt1����܀��;�p�����tMy�iO�p	-�=w�nK~`,̰����.Ruvm	2��*�k��,;x�[�W�<c1�ߪ�sY��i݀8N'�;�M�rvms�� O��j��:tN	���"������fͦL h�](�� &~P�� N�)�R6c 1�l�&\!F�����m�� (�l�c�S���Lv�����! ������;Ck�0(X�$�L%��z��-(ၬ���@=;�7| ��So`�u�%����`1��Vhx�ٱ5� *b����:�� 6�j�� �y\)�ڳ�CK0�Ȩ���!�O�i?�pp��� �9�4;$_���A�G��`�:l�d6~!y����,H���5� M�o��l �\[�x1y8�'�(�O@m�.w#,W�����aE��8 ��~��ufںd ����S���M��(���dy0��L��8>%fi�ESȣ4 lw-��#�!pn@�M� ���.#ulP�@� �<~& ����Nٖ �tS@Ϩsl�Pc�L�$PH��z� ��j��� �"Mc�a �wD~�Z���0�̳�wr��K9l�\�>�x,ޓ(��'# %�qs >�̕3�L[9of r\ts&c ���}@!L��b;uO�HH��@uCW{���X81���.�e�l^Zm� �������s&]}� O+�HI4�'m"��LG��L|s�ӕb.���H�oD)�s~ഄ9*���!�� � 9�L���$��+)݀�怹 욱�'�NS꺰L �D�c&����R�\A �MK|x̣'�.�t� �?�o�	 9�'Z& �Lq�R��y��Z�8&�v��֓�1�.y@��U2d��r��8�"-�΄ ~loiM�!�"���W@�xEܺ@���� �`Ym�� yS#�
ī����� f��	L��� ���� ����j+q�,Z}�.�%&�ˆk��$� H��!��8ٔ�j4��$\D������<౴�� �kݼ���!Z�,��|p]׎�B���l�X ~�sM�iNT��<�%w^�$�� '�٨�m�,H�$��`�w>�J��$���|1��Lw�~��p H��n
u��3��h 2΢kAf��h >@V�~����� �.�'䜨 ��$���a��.S�  ׷�'��K�j����o����L0v���_�x��>8p�E�!��8��n@8�� �ܜm����$���? ��'S V�.��dt��(h����b(�� �p���u� LM[�bE���H��B�@��jM)S����Lt�R��'ˀ��)v�%�����[<X0� -.$�F�/a���*����'o0 I~���Q��`�`|�kV{�0z� �%uAO��� M�N�L�z+ l�GJ��W�'���(��>Pl��*.{��j;�d�-j���}&(_p �L~>&. *��	��4Y������Lp{�)O������:$�r h���}�'� ��6H�̗p4l�W��x ��$u,��H 3�@މW1p&�g�G�11�U��#%G<�h���wH`��0�a��o��i��;���ne�L��`�)E�� Wn,lY��� n!��'I¸]� >�z�E���x� H7�wM ���2a�4��ِ� B���f}�"��,�< p��j ��.V��
�����J�b�*n%w}G��Q� �s���Wݹ L}F!� ٣%Vm;�U "��	u��,j�⅀ #(C��I�y�;�Vo� �s��5��s���q��,E+���&�|F���_�� \".Wm�䙶�����K�&,S�(؀Ӷ��� J�?�H0�Px��&at���'g�pgiH��
��JIpy�`2��Ep�$X� @�P9�쑸� ��LQ'@��9�h��p��+�?�&�L@M�J�|������j	T@*���ol C�"f����vka�D��z	� W!i}6���S�h`!�+y�o��0��((L��<���aC��X�	oE~�����p@�ŗ&3�!��9�Ā�v�{�MP6%���gx�7��!�*���0k�SE�!�"&1"�	�_�����$>� +k�LR-���CؓǸ�n2t��O���� �@kC��z&�I��K
 d��� y3����s! �Lp@)lcb�K��A�z 8�t�H�� �2�L5�*Wb�}T���Km�tqP Nl�)]��<y1 ����'�\�A�L���D0%o�`���9�T�%��-����`@��` ���~��LjϢ���p��= ����&�l� k�~T�L ����7�3.���������q�鲐�������|�%w� ��l�+��.����]��.�,7�J��@��d}&ㅳ����Lh8�i������ ΃'����w=X���F��;�� 5r��v�A�H�lz�d�� �s�.�uɰ�H�$v @���tF Ծ)����� 0ia���o p�,���JZ����2�ɠ��,x Ao�s,&#h�<�t��� �)Z�ʀ�'��	��g ���s���8�h�M/����t��8�����ď��X��3ȼ�bۿ-��I~ 6�%Zm�b�p��</F ~'�z��AH R�f��£ 
�x-.���b'3�,��y��@K��Lݷ?\� iD#I�����nø��t:߀1^p�ZK h5��NA��;�yВ�	���ԛ�mŸ��L�n�,�wl���S9��h�"c����$� O��[�9}�L�p?z` �s���vdi ��Qgo	�'Z#��Cܡ���k�iw�.p� l{�C�Y=�(�d Q|M����XdY�q��☏�����x+xM@!ɿ
�E�|KH���j&9�o '.�Ylm �(P`�}��q�R��M�����Q\�� "�!Ä|AI�PG�w�� �� sO�+�M m/疉'1� ���bu&n�����Ny� L!�w�9~ ҈Z|{� r!FNOϨ V�[mx:M?�ă����z8lV�v [�4�2�@�{-'\�z�`�nN��gC� 
h\��s�4z���U8?��y��B�}�x�� H3o�,n "ZdT$ 1VP���.�^�
��4>��l3Y� L׼����䨡p �'Oam�$s�5��!�Ie �hw3��7�T���F��,@� ��Lb,>vs���V*C &c���T m#z{Mt� [�s��E����1�Oh(CR"	��oϋ $�[W�� f��H5�� �yƫ~� l�Z"�U�P�� ������,�G�¢��L�<_H-7�L h���S���X������ �ᱫ�G�lg ��~i� d��b�� "M|�1� ��!�'��o��Y�{���PB�k`+8�v<	 p#�4v !ܓ������" *4nW.# a�ͭ N�"�����.�� ^�z��_����c�$�r��p�0�וg�L0)d Y~H.� x�&Xn����HKm��a�Z���\  �gX@l� �?P���L� ��!ޟoi~G�Az-�<�0�2���d �~Au��Tw} $n���t��  OK������8�> .�'�O���*H�Ή�!؜��x�c_c�π=�JeiK �W�s�� \�k@�ǁ��LCd'��T̨Q �.b���U��[���� ��>&�Kx3$O+L&( 6��E�;�~�0�`P�xu}�����xA-��w��b� ����<��K�v��t���>ǸvE '��*hJ`K	\urs�Ԭe�! ���c4�� ވ^[!Ξ Umf@��G���x����<�{r}&��..M�`O &�?X����>_P�W�� �z|S� ��LgQGN&0�u��p���
��~��<H�� ��`���� y-��tk� x?A2�ˈ�5�a<0�x>�oX� ˍB~��M�D�'�L�p/ "��7�0��Ph�$ϵs�B@�~��R?��x���9�٨�r��m?(A�iĚ@D#.h)?��!��;�x FJ�?������a��>;�� �#���iL��c��� @�׾�I���`��^CHT!�? ��0���^�A!)�G�$�y�UFR7D'�$j��1�����_�%Ws	J�	� sy�D��1��+��֊��T�˂!�� �5��g ��ޕz#'���s+]��K�x�L�FmP��\]�� �ǜw���Z� ���s婔�!�M�`�L(ә����K7
1̇#9_��!�3��YxL�\`Y�o ��|h�l� ��Q�oz7�`��'`R��"^Q+ T
d栞�5 ��z%�.?1" L��X���P @:r�� �%�S!3�9�h�p��ofg1z� H��|B�� �ɝ�s�� �h[��^X�u� ��s��������!� ��P��\��>� ^�z}׍�雂��2��s�a���xހ"�8���p<" ������h��Gp���IX<�X�Ʀ3���L >���:[:h;�� .� ����4�� +z��i�oI�QT����'�\?� V�I���t{ �Y�v326����F���;�5E�]�:jO�d��A������� FG\Q������j���� �N�b� �ȍ�����o� E�Yl� 3:z�$y�� �i_c��vr� w��a�N !E�b_B{� �SZ@�sg^ ����8�5{k����FOS�]� c�R1��!5�c��f�m� \@� ��
�� �<P?9�s qU�>Z'z ��IX}� cK?�~�28�E�3=@U��Tu��/I�n�)a�ܼ��Wp��H�٠���qZ ����Ar�� &���g��� ;��>k�. r�)���za���݀x"^ߞ�y P̛����@���0�H6�տ-���a3H�����]�{� �m͵gR��q����8U:�������L ƳoA8&-� �Z����?�Dx<hR��H��mv	)�
���=G'X�Z0�8A�^M�&�l�� �3�
 ��nO#��"�F!�@��y\C ��%e+g>f0~�3V��N� �5�> �-dAs�!�}����n�f�p��:L�G ����3�� ��I�� ��&�y�gW��0�,�nx �H��#��9�-�1Wz�6�����0VL
�>G�X� ���H�.�% ���y�a�����U����ES ��T��(�a�  f����� S��zB`� ���yx���0`��>��Wm 9:XL�z\�K��}�� E��`�8�@3�	�!e��
n:~� ��s�uWL�e܍��Y 9%���mM���dɘ��hYi�� �	̉�w �0���q�T��Ԍ�����n��� Ł�������x}���jΩ^ŀ�%	-sY��W����b �Rj�&5�� �.LP`� ���ߡk �᣸��� ���OeS���k	�٭�$��|�|at�7 � D�FE�m��pѶ�!�F'�甜	�� �Ó/�s���*ؠ�":);>D>	,o$2����c�`���o�Z�Qi��4���P�� �.o���vl�a/�	��)PT�[:��y��!��z��e[�1c�`� �uy� �Xh�7�D��a�A�lM��8W6��  �X���� ^�t����$�PYh�k@Еr) �����N<X��l������7gS�M����˰��: ����������G��>� �A%��RE\��ڀ᷸_ �sc��9���U^��"��q�sA,�:C�H !��V��r ��7' � �s�|���~� 4Ydp㸛 b�tؽ ��j�n@]i\�$0LP��=�w �e@!����ߐ`�S���
�R����ׄ"�C*  =�c璍�Z�92� ��h8���v�:U��Gfp(A��']?��y����M{�H�¥f�t:�o��^-�!Ў7&<? ښ�o����Ǫ��K:� D2���AL Ӟ"d��O 0���D�V�1s#. ¬�)&*����'j� �_ Q���& =���#U�$��7�I��s@�>�C_�� �$��%� �'�x�[�� ���*A.w���}���Q�'�B�p�b�� d��܆�/ ��v19���o�@����8�q;�z�H�� B�؞Sߖ� @�l*g k��v�#?�98 ���V�� ��?����0�(l����1 ѝO�	a3tJ oǠd�D ��l���(�'��P\H� 2c�3�&$GD�g��1eyԧ��r Z��:w��� N���_�0'P;+({w}� ��>��\�ϯ`� ������R I�6����Q���; o�R�iȰt��Ն���f4~=�c���H} �-�+��0q�J��Hdc��� ��	���]�ن�c��� �h�O��� �!p�,��.-9� ���gx�tP����t� -�%�a.�h q�ہ�;Q�g���=	��vX���h-a�Q�ܱ�w+,�> b8r�"�I����'� ��/@G���s [��qɶ�r�	�S�[��. �.ç��pX$�ɰ��?�룠�N���=��H��,�	k�ԓ�v3@��f� �U_��۰� 	��j� <KOU�L ��Y��љV Ϳ=��Ȱ� :��̨Qc.a݀ �z'�� A̂U�V� �����C?:vd�M�A��� l�HU��2� �}�Y�L� @da�H�Σ�qf��c�Ť��N�dD0ɀ`��Ǎ ӴeFB_Z
������ݐz� p:I�Ѡ��h[r�~�v�⛋�?�%p�`�80�(i����J,A�`v�`���3��k ����^�R�(�P_� g6���� k&����>c $��
��_��m d�)Fn�����@\��a�z� ^��F��)�u9���p\Φ�v���ρ�t ���u�e ��w>p��4A�3P�� f=M���� /�dSbK37��
��]��s@FD��!ŀ0��A��r$)	W �?t���g��`Pޞs� �R�%Ü�, �S]��� ���C��OIַ 1�R+����'����cFfр0V�[���� �Że�� E��aޑ��RQ- �gC�� z���~��r��@��L��]�\[؍�a  s��mX�<����4Oȳ�!���/@q�����G�D��4L��`g�wV���L������G�8BT�02?x��8FX ҙ"���U !�ZkN� ��>���
�+� h�x��*�[$ �� ��%�ۥ�:y2��#$ �Z\i	��t&2�������u� ?�`:��x �C�U����HF_�`0���@���y�R#!��Ɛt����N;��H k�n�a�:���� � ��vP�j�J>� f�ȣz1] ���v�*��ҼcA�߹:�� �tb���8
���lo ��FW���������z� ���2ʶ͘ ��n�t�cx~,��s0����^�6�I��mG�E�ؠ}Խ ������XXBF �KR��0= Wt8�d��:��c��!M � ����Nzܨ�2�P!t��n��d���D7� ����L�Y� ���>WEg�TpA?�|sN 6�v����y .��!���QT<)c�xh;�������B��b�!$��qr�����Un@�V� {}DWZYp2]�"�Cp�K��t0�P �� �H��E�k�=wA�y� �sU�����H�<��j6 ��$Ӡ�i�� 'HǫFr � �D&8�����2���O�M�#�� �kb�^� ��A_�;�f`�p��w9z�tޠ�Ȼ�� �[<�������G`�g-3(p�`�8�Y�C�},��0 �Q�	|�#)���܂D��<�.ߩ� ����y��z�%�}�&��� wd�2"��H��P��H�A�Lr1��$�� ��&�>�( uA�X{G� ��1s0��F �4�ʊ�� 85�R� ����|� P/\.v��p6w_b �~�� n�k�c7� O־Nv���<�Z��)���\��q֟������?� �rSP�vX `1u�[�4��o7�8�V�L1 ��wN�Q��˘�K���CU�1�p�v� �Ȯe����&v���cᴀ��C��\� ����:� xI�1�nL�`dub@i�� ��>�$��� ���	<J{; ���O7?P�f%�πC��m�=Uu�ؘ�t� !�&�� /U��r_� �"]+�Ѷ ��j������me�_���� ������hd ��'�j7�H}����L��w��>��h�CD��mu �=�ϔ+� ��\�8��P�	 ��Pr�Zv�}.n,<���X��g zu�.J�G �/�k�{�� �VդM�n�<62�88Qfr ��%���t� ��=eÂ�� Ld���)� �I�����:D H�:NwX R`�}�f� /�+�w�>���
}4�`��� S�8��:�| �X�Eذ����:�����$�A#M ,!�q���b ���O�K�u�<1tk��A� ��L[���� w)un:� &F'h�C�d�]
Ӆ�M�Lv� ݟY%2C�B�����lT�F 9H|Y��H�� f����g;Ġ 
�ǯ^Pҁ Ou��7�	��  Q�G�ݩǅ��D45|s�4���r���0T�5|���"��H�8�
�q� ـA{�j Tuy�r� 9k�Ҩ�ĩ݅������$���&��z 5��� P�e�� rZ�d�L?��倾��#c hq�*"9/�(N��,Rd��`���d��� !5�G��$�48OH u䯰yTK��ϘL��� �F���4 MR|ly��\| ʗ��U ��ku����>�}P�x �p�@�f;�,�`=��`
 ���	x�Og��o�H���$��,�88�����L�����0��2���S�" '�4��Q �r�I�塐� �ª�D�� �4@�ǿ� 3�u�*��7V,��H�$t��[�rl ٜ�n_�ϢW����������6(�v����t�wn`��$iꞭ��IDXF� ��?,���f����\������K��Sߒ43�Μ }v 
ǆ�������Ao�q)�e�P�&d*ۮ��ځ���7� ������L ��o����W$TL�W4ݠ����ަ�y3v�e�9�Aۑ#��z@��������u��>�8Tj��T88TLe �ݷ�	+�<����0h5?�� U�°,av�hȗx�;���> �t? �ٞڰ���Z�������5�����
��H �g�V�(:� ,-����u�"�M��|����ip H�* � ǋ���1 ��}$2��H�^�U�VF�| ��nݪ5�I0�{zҶ :���hэR IT�%v�Xd��w��=��ސ�L�R:쀑7r��x/���|o@g��n�$_�h 	q�TϚ�"������&/�X=zu��q�3L�4v�E�I�:l3�H��ɓ܄�)�H��Z5�H�: f����"#v��20c��)�h���)t?����\*ܐ �u_�ҩ�/k��Tr��H����$�M�:!�g� P�0v H�'TÕ �]�t���� �j�/���~1�`B���Ύ�� �x<�NfPL�P� �\/�gb ����*�P�� !&��3 �@��;�Qu�\��।���@�F�ODd�u��8\��/�)��\M�ݏP����)\���!.��ޔ\y �n"�	��\�)��,TU�����,�\�8\P�!@��.��>��lΦuA8� G�@/��� &��1�}�I �ǦE����F��~��p#m�8 ��ƪ����z�6��$�p< J��4���?r�&8�9$��@��E����`I��`�;g�2G�8��`y��P�TM!>vd��R=�%� ���}?'�xH&`8��r	��]*`\$������ �aR����|]s�`�� �~lpe#/q�ǲrO _T�3��`����� �f���4�1��;��?����ޠ7X�q� ����1��4 T�s�8,� �������V v�/�x�����)Àբ�� S�a��H��� ��Q(�:{4�x����H�$�D���D�d�@ .5��P��� �4���p�FM�C�Z�:>�l��A!����@6���&W ��]�i
8�3ҡ�U@��b_��I �6T;5�� ��v��8�' �4xA�S;Ӕ������ (����D� ��&A��T��Y��Τ;�z�؟��g(�F W+m4�q� �d�H"[8�v$�a���
�4� �G��^;�{���a@w�ς�!>���|"��!6�(�2<y���\x5`.�v�������K [�a��g�C s�ͦ^��=(1I�� ��� �h���đ��6��w�[Ű�ˠ qQ�%� 	
6��.�� Ŏ:�?kQt9[�xG��)7N�`�q�E�}b���M���� 8����2P��: v��RX��F �"�V�|� ����'۰| �%��M< �jb�&vtY\�L�~�����m��1�2��䜠`�V@�8Z=jh
��b��� ������4�e!�� ��L:9u��T͡1�C�H�׈A��8e��m)��o��Ѱ�1��']�Hw���C��|����Vs��\)�͔@���ly]��A$k��!e^ug ��b.,��L������Шw���� c�p�x;��8Ñ H��wv�C��/�{��� b��9x��B�O� �?�RM�PϷ� hvL�p�o`�#�b��8����S�o0 �X� 7`^�3��� +N��B�� �ch�dA��v���Lc�[9K	 ��m�u� �O}�d� Q��KFC�  �����G$p�>����[ĥ�@�H
���}Cp�����!�`�nfe� �pƹ?�����A5 �.�Nb~E���o��d��{�i? �HFg&��$�81��X�����` M����]�`��;Y�XNFS%H�� ^0m	������ �M���0�'0=� ���>���1�Q�c� �`���of�T�p0�1�jHr��ng��}�!y S���U O���#��,PR� O���;�\��6D��_�Yx#�X�N��\��&��p }��WKL�}�lw�C z�\ 6��!��S $)��\9�����G>@���"���>��,<�������a��� R���{24�- �`[)`}�(0�:�^� �rGq7��z/ ��άe�W_;n懢[�f�\��ь�m%g2� W >	��ۊy�ʘ O�Y,�/����؀��!�Q<X�x+�`���!6Ԙ7!�= �*i\�ȏeZ������������ jOt�Sh�isK ����� �Ϊ�P���bx�J���	)�� ��r�x/I��:S�@`o��2�L?�MV( -�����ty �7EY�t_�8�K��N�]���6���sH� a�����2�,]��L=�� ���0s:N��O�$�_m�� Z��p\]B���⇦��"���?����J�c7��>i����n: ˚�6�Xr 
����R: ��1Ԡ�P I�/�x?��� ���G7� ۼ������.a�H\Z%���i ��N��9 �c-ќ~����퇡!j ��@ϣ�kf 	�<��5# ��H��/�T�@�_�
P�`Ѱ���!͠��+ܲ�������jݭ>/�
��M`�.��~{����&0� G�m�!� )Btl�0׋���	�i`k���#3�2��jẅ���X�0��@e�����
�� �5���s�X ^�x��L RH�^�{��ꄾ ���`�QG�&�ذ��% �u^���?���VN��Q��L�>�l���_! �p:`�7{�1 �� �M� `&��(�?ꏖpI�v�+�PF��C�� 5\s�e�� X�i�O3 �!F�N�������:Y ��ُ�};  �4�,`��D� ���9KO_.�L�"Ay� ׬��9�k� m�{�s���j��]z1��D�ؐ�U�ﴞݼHv"Z���x��{O�X�w������0F-/c���1���f0Vĸ�_�<�m�L�pÿ�/ܠ��j ���s�~8
��� SU�.�2skw�@�d
x}*Ą�y��� �'���V/ ,�Q%иS(�"p��=	��{��ː�g ��E��Be/�˴x�0�Ȁ��|Ph�E2�1�俋�B�� ���H~�=JI� `�k�� ^���i?�`�g� T�<���!�A �^�� P+�FW�� �����˝���{�M� (*��F ��1�Q�ao ÷2�7#� :��~���(�xU? ���j�zt�7 X������ M"�6�{�������	�7��x�Q*������\�����Y"�^�� ҍ��]��KtbFE����gY�*8���:�D� EUO�`��"���3:��B�)���oIŠ����@,��|��h��P1��x� 5�����t����C������x9@������Zw�: v������ňQ��A7����fPo�K��U�`����3P�#���aW(:��� ԅJ+U�Ɔ�	���[]��S�}`%
J���L�0��p�:� v���(a���P�2�(�A��!8����� _�y�lD*
w�NkX��r����J@����<�� ��]��
}��7�<�����A0&RL�&���bӧ!\v'D�H�\B�@7k�S���D���R"�T��.� G��>�`i�Rp�F��h@t�1$����������m�p���{Ѐ�RŘ� �)�FA�� #��mޝ�V�W��f�� Iib��cT�����k���e�}ه`pXw�z{Z�p �6 ��?��� A�e�:�c �!ǹ}i8��?�
㆟�⁐}Z�3��>�B�,	�Th~Ŀ�Q�= ��]w��N��й#cq��zJ�D��Gt^H������4� K�j|V�e��Pp� ?��O�=!$bM�.����Ȍm�8�Y�M���s �`:1I��!}��/@��P%R�i�'��0g{(\V� QC:9u/dp��yY� nT!�i0GN e���� � �r��s0M�
\2���:�@� L[�Z�U	k.$NA�M�}^�Ҙ�������ֹ ��1{z�* 
~F�5	  Uh��Zu z�E����}Q�P���3f c%ƉGL+����@�j��� n;A����~W�!�Pu`2Qw G/
:v�>�e� �Ȋ� V"�hm3i � �'�Q�+ ̃��XZ�H��0�I�@��� ��T���tD�zu���6��T�<h� �`
�/"���J��� |!��jhv� �1%X\Lq� k�]#�'� U�J)�h� �y�\�D5 U����+P� ������ �����Y��&@v=����ttU���ҙ�@�G� ��u��d�3��zb~��� ��*	Lu�|>��U�ey �3�i�w�$Th+#���E�~j�ӕ[�Y�� 4,֬�:a�:��Fm h������;��]��=j <եA�
d �˄����~�	�᠝�U��� 0d����AA�)� _�?���/�=�i{P �R! ]d� D���׽Fn{��C��%��:霄b��z�v���-��/x�q8' ���_�.��ҹ��~��� @�1��m; �X�9�Z8d�@�W" n�@6% ���-xzPr|������n��_U!�Wq0�� �"h���( _���!�)�k� ��ο�i�c�.� J���p �j0�) _.<�F�{"Y@2�m>���b��J5ji C����: GWV������X���R`�v�5 �=Oؖ�Ҭ���|��k� ��@u9NוN� ����½ '��R�-��\B���u|����  !��/>?� -�@}8��נ7Df �� N�)������;h<z ޓ#j�^�g !o��d�� �����[rh{�ݠ�0�.ydx M"Iu;��|����S�O k].�z-��>����~`��F�� O[��-$^������4� p+�O�����A ��)���	�(z����ޕ� ��[�fO>�zs�D m^7*3���!��{ MZ�\dm�q �z��� ���t� |0~�PQ=( �S�+t�t =6<��e- !E��3�� �/ϴ��s {4���pJ�)�od������TC��4i�.�u� :��֣~���U$ ��Xv��.� a6����X&L��
7�Y��<�����6t@��8" �i ��J�k��	K�&aS� >����Hp+1o�2墘@�
�
;ѫ�� P�>Z�� ���4F"U7��ߌ,vhYD��$]�8=w��F *���� p��D�tR8� 5����� )�χ߷	�o0�P�i�l�64�@�U� 2��}	�x!� քp� |��h�,W&�c� Q���JV��+c/݉��XL9����׻b@� ����$6t��zR�M7&�!ni �:I`v�d
�����%U6A pǴ,��
�׊Jl�Iyz��/j���}�-���z�e�%˓���x} ���k���i_[����`�@�h��נ ���WG 7���Y6q� 8:�ן&g��ܖ �#�� �$�75el ㆴ�[�B����n41�������G ���� �tP�e��$��� `,��a �x���/h`�)��60 }�i'�w�0	��3�8b���(v�u��(�0�`;M p�,'v�]F:@(�j��� �frBa�Ӗm@��¡�9F��� ��3�\o~�������/����L"p �W�p٩�`k�EM%�3
�w1������ ~�:X�a�������A0�mi	�p-�<\:��Z��@�%�ݟҰ� ���XL� �
�� }K�05�B�����pU׼�8� F��kߵ$�� S����2�=��b� �|��E� ~O�غ��0 ��"���M _t��7T�1 �%s�﹊�W�� ����6o.g�7~��*�O���RB4	v��� �[7�,�	�.��@�KQ\G, �ls�/�� ����`�GB6k���Ώ�s qԈ�֚��F^н9��M��D�{ A�x6����r��^t�0�� =���\� ��VL@t0 �|�u�W�c��e�[nj@��1 �D�{����� ʴ�C�>�� @��U\X%� �W�C���SQp &��� �]8g�{� %�@�pW* �OE��|� �GIN���������Z� �}O]#�A6\�0 ��U!�(�^� 0��sb��$/�X��A�`���('���c�7 CE�^��W �v��&p-�� g��ԙqނ 3P�έa>lW��	����^ tTU��� ��d�3_t� [>�r��X5 Pq�H�G�?p�� ��x� ��$�9g�c�6������� ݊�Vp%.t� R�ܺ��� ����̈́ }X]P�	�w$ Fp��Δ;��\��%�������C 7��r?�L��6� ��(/r��#�����g6� ��^�ޔ���x���k�����)ŕ��.��F6׺d�̦T� �8�>� ���u��k[#��x�,s) �u@��z� n�Q��P��ˆF�������Ԅ��<5� Uƃn~�p�vN�����I���5�S��-i ���@OR c�;|Z�~697�ي���4Ӻ��_�2n� �&~x ��BӨu� ��\/g>q:�^�|X������Mo�H �<�"�� �Vҩq�^�DF���xdB�j�\� �w� ��t���8 u�I!kd�� ߅>F�� �ޯ����x�t� �i�4���zJ���˅�E�d�� 5	��O��~:^� ���pz!3�AE뎩��r� ����k��� iڥf|j� п�"�Q�p�l�F �:�A�i=� �����K`���Iا �Z���b�yg |/���z�z��= ו�����������@X�������(G�W
Y���¸���eQ#S�z@�� �DH���I� Ͽ������:�y0~ � �f�t����͊8X��  ��� �r�F71	��$D�s�{!WID�q����(�=UvG;!)����f�\�,�ΰw�>q} ݀�����	Z� �����~T ��Y�z6� ��[c���,�#�9 �~l�}!�1[�0��� -��c�OV� 8T4�D�� �Ʃ=��k>�⁴�|��� 8�򃜉�Z �3�H����LB���ѱ����M@�Hxs8�4���t[��� �����E�L4|=@i�5���z��w�t@0�� �v۠4��f?�w������9,g j8�6��� |¼S7�&�y� ݁#4;�x	rã �����Qq�1@�s���! ��ۅa��6 ��E,�p> ��x��J
�9� G��[�.LP� �S��~_� I������h:Đ �*����֘ܐ� Pr�m� �hc�(ګ� ���/�������֐h�����рTq>��R��)��bv��<�;�߇�F; ���� �i�ɋ��@������U���/�}�K���D7��Ȅ��G�_E���v� [=�q�}� <|g���RA˟�C�e���v��V����=T�5����D�1{HC(?���6�j	�	���� B+ה;G3�Y�}�p}� O����,g�,j2C�ɨ�Ԑ ���|�A� Ь<9;~/>�D�y�zF�t��S�70p���9���y�}�|0��7�0��?:�B����O�Rs�+�  ��.� q��a�}|{L�L v�U����L�� j0ߪq8O �9#����=�,�l��Y�<��x�6�0)q���|� �4J��0�X	*Ex� 7U�� 4�Y!I�d8���|�AQ ��xIs�{ pӷ���j4��i:�S[���z~`I��ڪ������>8�xHE�g ���p� ��jXp� �v����C �b�҇	�8~�BV��y}�)q<M ���?�tO`�!�=�f�q.���	91V����C}B� �����,f�yLLX�|D?IC �F\�[M>*��5@�Q�8��D��w}�`�k�:R�V��{�З8$� \_'%��G�ZTR@��i� �ab��@�[ c����7;n�����pp��S9+��H�*H 8s��O R�+���
�rSt� �ǂ�2-���&��I�:��(�&��8 R�f,C�����w��o) �`#���:G5z�ȃ4���8G�9�������j$�h�����~��5"����XW �%��\E Y�r�NU�P� β]�TQpZ�-<�3�Ԥ��C +����|�x�  `����Y�3� (��R��p�0GS�	��(1� �;��0S٤�i GN��F*`j��1�70���oA��Wp@T �FB��0(�O�+�F��;�!g7��>|!G�𷍅�x'�~�w! $���Y�;����Y-��[��YmC<�C~aCF�S�@~�Fu���(����$V��	]� |o��8�:���JV�t �@��=sk ��R(�[/(�\��&�'7��p��� [@՚�À��{�-��,� ���1� a!�oXv. ��;f��ͶĐ"246 ���h��� ���_���4�����għ0�?�IF�qq��Xt +�G�HLO� ��!����e �a�/���	�#F& ��aH�� b���ډ �R|��F/% �9W'��U �D�(g�����|�m � ��C�u ��FO�ci�����0�k ���<�	� �wV-"� ��
��1 㠗��#E ����J]�񍮅X����F� 3�mΕX��� .*�@�0�~H�� 8�[��&��G������Y���� �'�G<, k)D�v�S� ��/@|�
^�����XP��`t�G�������y� �{��s�� S��wa�P�{� � �OT�3��x ./��\ �bEnZRX1 N�Ϡ�<�$G� �2Bq����G	��}Q)P4 b�0�� ݽ����k ��Gw��{ ���.�F ���X�A" W�z��4\��^��*��
 ���o?Ża:+� �#;0��F$�D  ����0��(K��PJ�6/@�1�c5\�` Ug���$�� �4�	��u�`��{��}�<H�p�]��t#F����s6�W*�;���Ğl�� Kұ��]<m����wتpr��M� �N���� ��iC�[1��~^�x� h�� ��Q��^L>?P����@���� �3�~S��w�� n1�ބ�c�^��?��e�H�\���q��5�u`��Ҁ� �����*�����gJ��{9 ��?�Y@� �1	��3���9��N&]�56 a2/���.]A�ڝM�C>;*(�� �Y���+g �J�q�V�h`m�{�A�?�I�@ ���S����t�* ��j�{��� ���Hx� ����L��5��R"�8�P̑,�?�>��\�3@���H$δށ/2�䯺	Y��T� E�}��y:�x�d�a�T�:��Bx�}T�_ �(Ы�����@=�P�m�
>�zQ�7� .d�q���~��<����5	�º� Ԍ�u=Y� �×��� E���k�� �lZ�-ƀ�V�k� �ۢ0�i�T�! �����z��i�����<矞� ��Q�/�9�\�@׫w:���4$�纣�� U��S�3y| �4�}~�e�,f�N ���Յr��^������x[ f��7՝���W�����G�	�1��{#��ȃ	S�?� <ĳD� ��ˇѶ��a�a
�"���8�*�h �i�o �=I6p�!�+� �U
���F&�z�Y �pP��+L�� I���� ȫ]�ڬ�d�3�� �+� cmP6�QY����( ���5� �b�o���@�6qF��E�*�4 -�ݤ`ԧ��>@�J��u��o��G��Be�.�D�(�k���l"���ɠ$������V��Oe�*B$(��(�^T!��
z6.��`Fa��@\ q�ܟC�|�(Ѩ��� <V���H� �6w|���ed@�?1:�t�HG�M Nú/"�x�Qd�����u��],`�8 ��P9j�\�t��"Z�`��/�L ���r��y�O ���,| ;���Ɠ0^C���xFP�6��$����"a��.�z៕��g�j�0 �p#^��� �o$0��}lTQ�<�N K,켉#d�郷i����7L\�;N�	=��
f� ��~o�� ��
!3�u q�ݔbCz��5��Z3�<<���o�!�G(ǂ EW��/@��$d����XzB��}L�U�V�� �3��D� �7q��pR��� lX���@zm�]H��60�u&���@��%'�)�Lt��Y�� �W�ƍ3�O��a�_��+�f����/o�G� d��F�50�i L���R�����^�@c#�x�$��PAN�'��C��D�i��R��P��@$��4� �_ 1d�[bB��`p25��G�J��¹rӛ����apٲ���7��h�&����� ���>8�w�
�UA�� �p���[*�(� ���{J�,"bVS�$�fПA��%��WHd�	R�0�8y� �]^��JH�Z�nf#��EPp'���L$�6����c�L>��)�������&���<��� P�'�+�q ���%<�:l ��k�Jq:�`��(��Cg�>����8zz���ɥlD1�x"���� ���`1q��&6���=�"
����U$<� ���9�j� +욈��1��U���!p�T2�t� ��7B�[�����=� �䆜ۇ����0�V%o ��7��&�� ��?�fAR=����
Z@����Q�i�����1�H��ʆ)�x�\;��`��[W��c� ��`�&�f0,%��']1�4��&��^����<�t9�J��f\�C��= %��� +�n�RQU|w{sȠ��T�@d WRo]%�
6V ��"����f�a�:�0��!4�h�D�u�e *
���CH�C��pJgF�:(���
kB8P\�#���pr�3wUOjv�V)I�p�����W�8��U���U���p��P�epBG�_^�L�p|SH���p���(;��T�A���k��)#�=��W8�qd�0���8��J]�T�}p��HO���"��H��8�!�LHH��2��(+Hq���S_>�����"��b�0h��l>�}�dJU!ȡ'L�hrˮ�����q��w�� O_F
�i�A��al	����iH�d�#��bh"f��9(	|HN��^�����D�	��!4h�_�kߖ�Y
hȩ"���X8��"��Nܟ[�+�4�7�d8@3�RƜ�ܚѓ�9Hi�8����!(�X��F3
��mp𧵎!hptӤx�Gk�p��F��7��E�$�8k� �	7iH�J���h��/�+HX��p�#��(a%xl�)�0�>��p�Z42jhOp0p[2;�&ȿ��p��pǨ2�T.;��Ua}h�pZ�%}(x"�p={hpHk�*�
-*=8B(����p���ޯ��pu�5�h0kp�K�;��� ^8ՕŨ�+�83�8���|�plr����G��+�H1�p��8�(2��>َ�����ƽo< ş^~�vpD0��]�8!m��{��bF�=ˀ�-�a�8������Odp�(}ꁅA>��+$p@�b�af]!0��ec���2#H�Ş��)W��� 1�����	 �m��Zq�a ُ񚂸a"��@ U+��h�p���L��> � 6^�I�p �,X��k�� Uo"Q!�";��(RJ$���`e�S!P��$�����w
<���Ĳ6!8u��T@ǰ��t$��S�h��`EG�T|$�RT�*`�G��L����H$��H'�S�R>�#�>��� ���0�#�7�$4� ��-9"��U��u�'��h1�������1@$��(�R�D-��`�h_��� ����.��,B}� �ɉ�! �x�����'��.@8[�!�0ɻ:��ߺ�j$P��[��i�?Ls���:�a��g�X�׋�2�����Ax*~	����L?�P*G_�)����aR(վ4h#ށ���:���&��buF�@�C� A]�!a�I9�ҏ*����˵�> Ff#�n���
@���� *�TƔ{�&�WDh����ns�Mp� ����"���� ߝ�1������T�ճG�3R�����ؠ����z&0`�%1�:A�v����PIp����L��o�oȧ 7����}|�D=o.+넀7|����$<s�K:��Tr �}�Ѩ;6ҼLF|	k$�= ��7�.��g [L����b6���a������V? !��7ѻ�rNB) ���ct,�&�: �<e��1 �����ĲȰ8 ?�s��ו�v�F$�,�I�]Y����!�%� N ��p1�5�
$��t�z��ɔ�$�7L��~ʌ�0
ҰYk;+$]0��%�SH�|0��&����H��<�s� �뉴ڻ��ID �X!�+`�G�{�� Pk1��ɍ�(��TӔ�&���@���������ʮfu` r�2������{��C�- �|r��+
����,�"0�)�k!X$:QPX5��m�&�|�H�a�.f8�� ����� ��OXp�0X����t����H&�1� $�Gnq�T���7�/0B�Xz  	�d�f����hg���@�ud�@��a�NJ �'+pz��� �h4���bo�0dH��
�  �E�TP4!� �Y�KAh�\�� ��|���ai�ғ��=`"P�[4���D0�0�v������)���������*�"� ��׬?�J�v�<�]T�W@PC �;�ŕf�LVh㜛p�A�����|�O�H|r��(j�� ������� Bf��	��'1��&@�ѹT�GB?*@�R��0������ΞBĬP3 ݳ?���|)4�Vb�ǯA��Q0��R�ơHST��R�am��,��$�tP�G�A �z�=�~`� ����B�Z�t�Cj@0�ȧ�h(K��m3{C��4Ă8���;���; �L㰖 ��?IP����K�dy1�5b-� pD}�>��	T���:@@�#� �ʶVum��x��v=�,�����" M��Kkv�J@���m+	�Bp���wL��`.��LN�=��4���'����D?�T͝`�P�ccYgJ�CA~�H��t8���Wr+�X�1a/l�Հ}Z���M#*G�@o���1 ۳�뺙�W Q+���C�: D*i����o�,�kАf * ���"d�X̧ 9Jo�,� ���Ơ��v�%��� 3��f=1q  k�MQ>� p�mFly��`fT��0c*6Dw ���o4e��� ��f��� �A:R�(X�W ���p�q�v2���6�Xm�B��c���4j��0~ ���S(������+�DC� ���[=lA xn9Ph� ���M�( ���H4�8��[�동�0�ָC��h���#� £�)��P?W�
�%~������,��0D) ���rV�O@ɼN� G�%m4!ҿ��D� aZLx0`�ՂH��P, �v4��P,u� 8>G�����!��;�"���p��ɹ���
g/���a<]i|`' ���b��`��$2�j:^,��ՄlQ;ސ�*``�TB�^������@��@	�5�/�����%Z���m�<wc`���h6� 쫃���
;P���Bn����"t���*@��0�,zP�0Z�� Y�ԗ܎v
��;���2UKb�E����)����쌑���C �o���KF>H %�^!����iC��E!`�h�ua7�F�1��J����{�`�2��v:O@ �<)=a;БysP V�(�Uo�\�1&��E�� ������\;޴�0S�>�G�P� @��r��f�Y�>�N%�l�1B��t=�`"! ���^�J8+
f������oA�<�P���`+X�̀@QA� ��KS����#Bx!ʥ���`$�;n�� Џ��(�'H/|�*�����${�!B���@fK�7�/p$�U� �<�,�>�h�$d OW���H�T��!G� �'��h�g2�[�NP��	��tW�8,&�O ���N<��0���s5�,� ����� �{d���MAT�^��`�\ �Jr<��8�y R/6�ۨ>$ ����{�e �8#r�0���x� A_��c{U���X};Нk|��Z��C�F���� �A��4��T�h]�� H8�Β��Y�n�vfذ Љc� ˤy�;��a����!��WM7�@���p �J'<�"��;3�	���&j.o98 �v���)�G�o�S������B�㌸�Id��t8��AƃP�� ��t4/��1"q�)�90���� �xi�h@� �W��)B2�I�X�Lt "�{��a%�u��H�g�a�:]���B n"��%� ��*����&4&��uÇg��о� ��Jm�;CT�<��a��2�!���% {(9)�=���A��]���Pf��@���"� �<:P��� N֔�\ƺ�x� �Ł�h`晫q�16/j؍�ހ`-���[ �0o�\�b��P�Cj��� ��<��RN~*P� nA�K Y�2u��O�ح$9�� Uz�	H�sA�T ��7F���� m���1� �h}�虫΁����c��ɀQ}k |�u�>�� ���C,;�_ G���
�	� �a���v��x� ��Չ;�+<�� 7 Z�IG�n ��j�� �#	�c|. aH��bQP� ���%+B@dU�R�Chs_�j= l��<���������Ժ�bpD/eQ�ۓ�by^ >@� Q����i� .B�{�,����
���0F�zk!��Z!)�Q� J0�@�p�r��?��) ��/T�]�� �Px����� ��)��g	��� =��X,���zSI!p��2��1����@��*��.0�{?t�\�$Ҁ�K��� +�����& �>�kY��� ��j9��Ӭ �~��81 �0���/� k�ɐ�\r�|s�*� �}.��y'
�P�	_�T4��(���p� �<��A٫1	�P0� `�4 ���hN��v�{��;�lrS|<=�À��"���pMr���`�1��� �|:���d�M�S�ʟ�tÐrF���jG�͠�vF��n &ҍC�� ����a ����m�b�qXΐ,Be*� ��֟�Y��� \8I���ƾ(���Y>]k �I��;m�9��sp�* ���2������d��Ae?>+���TG� Ѧ-��(j{�D�>�)7��� Gs
p�m	��)\�q��t�@F1&�Eo}�A��V���@m�� �n��p<���0E@P˲� I8�y��	 ���F�:���?-/D��y xT��Қ�tbՃ�����,Y{^ oQ�N9�1 ��kE�� ��0Pl	���.�� ���M� !ĕC�%ʔ �[1�R�q� 	G���,�$ �k`�I�E���=	� �o]��/J�����-H�<󨾸��`�3?��Gl- 2ћ�5q�
RynDpb�m �U��e'T��E��2P�����r ��V� 㛿�� �h۱�B:"	�8���p� зUR��#� Fd��=�E�[���Vxq%��X R曩��8�
�=)W{T�gqO�ap\��! �8�E��2 >�$(�(�W�q��#d�Ӎ٘�3l	�)V� �%,� 4KRm�EJ �)"F�{��+�;*U��@+�PYp���z��8"�#�EA�UY8�9I{0�����l!J�� ���]$y�Pr�l�4=��,�=0g�8�Sp�w���A_@�u����7��"�R)E4
j`�á"� ��iAҶ�SW��Q���%L�Y)�4L a�,�pX� K��OT�li
�lZ!�zGR�4qX!����& JI(���A� �`�Ww<�����k����#P� j� �7T`-��?Ug�|_�I�>��J$��R [n�
�� c���đu� _�x3��� �=jn)`e�������C fܭ0D-rG L��a��h�@�9}y ���$Q��)wjT�*�sB�#͏0Ȕ� �gj�ec�B������_t5Uq�ʡ�n�Y	QD��ҽ@X� � �Q���o>Z�j�8*9��8�Ā8��ړB�D�R�8D�`����TH�� ��G��<����@I
��g�)���A�� ejO�ע�G�	�9�Ӯ����8F^O��]�� ���Ow`��U�y/���$�Q4_����� ,J�83��E ^�G{�D�s�		�4�8���iO�A���p�Z=E�P+i�
Q�H�9HP�
��'I�lI`�x�hE"4�^��A�`R��@v3��e=,>�i�p-�Ҁ��4�8�r���T6ĳm<_D��~ ��*hrX��>��{Jù� eYc�M�� ����m�� �cW�� �V �;�Ap��?dT�,��h]����c zq7�Wž� Ko�ם�f<?��h`��\�JA��n�à�
H����*�W�|��p"e8-������L�w���1~�@vWB� ��K�| �$.^��?������Z��vO|����i{q2�C89�� hv�_f��[j]�n���`|��3b-�8�6 n}�Y�m��@��4�ˊ��b� �ǝ��?����R��rq�8�3������s������ xS���bN�9�C��s��8������Pvl������jÓu���$��� '-u��;�� 	N���k�� W�H�GP���ͨ��5�� ѸЬu�[_ ������ ���:�Om=�v ��Q*8�[pD.ƭHiMH8���5ڸ�H~�-�������7��X� a��˺�� �뗰� �i.�[��& Ý��y ��߲�U� ��x�F� (�&�0�Ǝ�G �y�h�nKt� ���5�j� ��B��$ q�bt�Q[���_ �j&.
� ��݁�p:4<��L��z/��g�<m���#Ĉ���`mq"
�UL@g����#Z�V\�ly��
���^�� �_j�bF~�q	���!�g�p�G^����j>C� �zTi?g ��0�F� �)�*�a% �ޅ{@�^9BC�p[;&�x' ��?���
�UA�C�3R ��4�~� >�kyܔ� �t���Yo�Q��,��X��6�}v; ��{�YH�,�� �p�J����1 7�����؅ �S��x���W�J ��B�&<Dl� 8�1�9G�M[�Sd- ���4rD,�b�}�L�<��z� ��X�a� fR�P8q���L �i��Q�P/*� 2���+8w����p��T ��rz��� �vt_��_��8��8��Y�@ps� ���,;�8"�@Wr`�ꔃ�$9����������+� ��(�0@�x d��e��ơ�#�k-��2�L� ae�\�����H���&�ؐV�l��8p� A+�����xr�/7�脀��͒Ĥ���+����� zF ����;|Ȋ7�� ��d��} ���UI� �p���Ñ.��4M�" �Y�#��� _����º� i�hb� ��L�B� 2k����[S���.��67�)�YR��{D��b \��<�$:P!�B`� |oL 8�a<�Bf$:Ј����uD�p)#�8�I�7��	:��������఩$��܀[㹶�c�)��G%Z��$��� 8�0 E%�qm� ���O�!�,���:��FC+S�����Ĥ���� gܥ�֝`�u�Q���p@9��&8\ �!;��f�&�@P�6�"�UH�� �#A�b�i��^ ��:���?=)+��ۼ ����X� �Ƕ�X��1�8�D�S�<�T��&�LR"����w�AĴ�Q��7������q&���p~�)�^vꚄ�&P <�u38 �+2 T�W�s�	������6��X5Hь��phjj�l!pJ0�Ī��jނ!� ��C=S������i#��F�� Ӻ�� #W<P�MKIX���l����ظ�4��@��1���eA��c�
3)��T���\�L,#��Z�`
g�S�ь+�8��d8�3���q�ع��	M��8�)T5d �<�c�� I�.��� ���Z�сNA����E� ]R[���� Wk�Dl�g�<��������h� nj�;0�ؽ�N�`qӑ��=������j7 wBs�  ёl8��p,*��C8Ҩ �+��~�VvY -(����#t"Цz���pC)D~ �W^�m�%09���*)\ �Ψ��I�t�x,�>��.�;F�@_@�j���NXP[� ~4������� fEźυ��8�D��,�W�mG�7Z�q2a�j�L�u�x�<@aT���H�R �â�@m?x�����!��.YDđ}� �\3 d�ʹ	��61�$�u4Y��b�����TrP\�D#+\�#u���L&9�n����?�Y �����qG� M!���Pw?V�Ĕ�W���r �����/�X)Z���pH�kv�;-�$?�Ty\���6��J�
�w���\�T�����3�������	�������j8 ��+�<g��&���ޗ̚ l�B�
����d�����0��`%� ΐo�9���蒯a���q���r�c�\����b"�����ؼJ�Q!�ɡ�⛨O�p*�!��dŅl �p����G�Q!l �&ܜ(�{[g�0�8�*ҙ�|�Di?�P���};�4GI0�3�K��"��?�����*���W@�NU+&�P��.�es��$�Pԉ�6hШL�Dl:�,� ���P�� X�,=<�8�����4�0�pճ��4��>H4��f��$�PSQq�"h���Uܠ�� ���d��X�7U�&S��[�
�C��]@I�D��	�:�|��D#��Ow�@>7QY�M8�z6�8�7+�#����� C��*c߄E@g(������qp��(����X� �|�8�;R�$�l�Ģ� ����Y������#�� E������kY��DČ0�!K@!8�(�ޑ�%t
�W���!9�Lz 8�	�LPLipL%r@n��İ����lAL�P����N�6�% $���BD �(�S {��i'4 ���Ќ�S�ພ-8�9pp����\!r��`��U�u?ܬ�(�����3@�M\;�u����ay� oI�� ����6�!L0%M�d��L�� A��v�b
T��#��a��'@��}�0���e�8dupi�4E~���z ૒�H�:��@�k�W] �����g#H��^���xU ��M�.Q Vfq������?�B҂^��}� �]��3x���� `��^
X,xs��zqA
��
��z@�W�5O�sվ�Ѣv�8����C�Ӫ M&RH}WV�R8q �Q��
b�>��z9��V +2���O�6Ũؒq��MR��Ľ<� "��ȴ� �����$ �	�N�W� {�q��`�C P��H�"�OTA��F86��� �r�=f	-��P�8 �N��~��6�H��F ��9 `���u�V���� @,6ނ�zM��J� ц�����v[Q֕ �pf>g�z+(�J�ۘi�Z ?{��x����NWu�� 6���B�@Q�FA����N ���X	P��
��i�Z"��WG�e�q���`��� ��4�gWv�8B��q�V4�� ��~���M��04
i|�~T�l&��D��L(:p�
�<L FQ��IL�טhN��t�S�zdPH�� (M��J�8	Y.
"�z&�P��@Lyd���G����ʓT �N&q(�A��ۘ��8nެ��|H��,=�B �~�#Օ�f���0z}�uL�܆�Ǡ�J5klA��Ul!�ZlH�Vl��Vl�I�h�h�l�l����jG��B౒��V2+X�>�d�#s���ɠ0Hk(�B���n)�+�}���L�� ��#IG�=�	��1�#@��K�8?� ��&"�����2���Μd���pI�P����d��7}y� ��X6Y�� N&J��9�� �W���� 7�PG�v<a�@�qt" M��1$��y3���7�e� �	���K��a
N�j�8B.�� �R/mg�DLKөgCj;9���r7��I����wM@|�1�b�X�F͐�p���31H
J|jB��/�vw�:���Ƌ8����#���ߝ$�7�f����p@�i� ���ٕ(	5�-B��Z��9M%�L�]"p��)Kbρ�n3.@�AtS�6\aK��Ԁ��ⳣ^ǩYw��h��k,C �J�}�b�)�.؂J�G!ҙ@��#�������B#�`��Q! .�����=+a�yD�p��29�8�	$�E4�$��>@�a@� Hd�qC�&d�8c �]$��!��:Sp�B�٩."4�T������}T1)c�/��LA�
��j�i���1���T���K�qUPܢ1!��Nr��
IJ܏�1��B��@BPNL&���LY-	�ѥ`���Bp>ɑm�gK��)���RD��K1*���8��_5r!�I�$�(��Iy��^ܡA������L��"�  �ԡm#��/  ����� ��3A'��@ G�g��1 �"�BV�0 ��:~�M o�O� '�]�dv p$��2��� Y+H�/X�|=��b��=P@TB�� �zg���@����H�=0G�@N擶 ��[_����P�g ��]�D�/>) ��U���꒗�i!r�!��8 }(�&�p��*?�Ѩ �@�� ix|�9��%��F�|����*��wWI�Е��R�&� ���ƒUs8I� �P�J 
�4�(�A [U����� �����]� ���bD/�� �3����)	 aՁ��`K�4 >OU��"#C����X r���[��w;>\��U��ӡw� C�pT�lB=��n��;�U�+ڐ  �ۂR �'a�"������T
؊pQ?d��Sa�=�1^��!��\8ɨ��Dn������p�
 ��� vs"p ���{���� �}I�_ۙ�#�<rU�o" �^������ ��t��6K �-Q�W���%#M*a��T XO�
�"� ������? �k�Gs)h[�$¸� ��LƋ ��@��~�s<�iTp|�;������]��08A�@��[L��T !+Uhk����������D �J��r��p	F�[�f�9�v��[� �qS�u). �^�f2ߋ����=���[�K�vJ*)�Ӳ��~��T�����(�NA(< G�]����P� 6=w|\�m�! LH� ��ĸF���p�AÆ#��!'a7���f ��N�x�}"e���X�{�)Z~�����"]%Q���M�Ҕ��* ��B�� _�m�<;�'��6�1��Z���Ü�n�y^z��8q��� ��Z��m��H3}^� )�?���� �P�ȵt��p�@�^�) �?;5GF��d�/qu����
)�@x ��GmM�=�����9�(xE_��U��qئ�;�x�����
�T�v $�=�S �)�P��1� ��r�Ơ5��b�^߮��pY�¼ �t�Ci��'��$>�X�XG;(��u�Ŧ�,0�5���&�q. 8s�1\�)�T �*_���<D�Q����)�(�ą���6>��@,���1�i�=�PT?�� ._>��K<x"��O�@��e�).�TBf ��. ۆM��7�s�)#`�S�[|�0�78���w�
i.������A
T*�DK8��8/�|�V�(2�@|k!-�C���A��ATк�9ڦ�Ҁ4D�P�\Q��*�		�4�@���G�Be�/��#��8P��IL�f����Lp$�����M��8��8�_a-54h��/X���s�֝𠄬�*���	p����.���e&�v� u�W�ؗM^� K�T��d� v��"z	;��G���!1X)o� 	����р�eJ<W:5C���1fKt0 ����و����	�M<��sX�(�Y�"H�G���������m���ybLݠ���*&20Ľ =H��t�3hë�6�'��פ�GuV�1D��ߠB� e���1���ǅĈ�DJ0��������Q�Z�A�3Բ�Sp����� �2׆TA��ԨoԬDy�`��W@�d�p83���]� ����th� �N�����[`?����H)P(��� Q!�֓=B�� uf���A�t~�T���,�֊i�� |�hI���+~8�9� �x0� �Oe�ի ~9�d�Jy9� ߖ�XnD A�)��c H
~�L��P �Ԗ�Y� �n�ꨀ���~�{	�T �ʊ[���Of�� ����kB>������ �6���_�X�d���p�T�]�8n����lI
 � ��(��2ؖ
�I�Z� ]��}�bB�݀�e�(Z�2�����ZEB�ʘIP� ��Y�l�B p���$_2b��n�18@��~� ��N��y�� ���ד�AK�Z�tq��ˬ��[���URU��E4��Ȍ��QR�D4 T�T0�q+ 2�t\��ygH�W4&�0Bҁ���Y�pC��^�PT4�	�� ��`>
�T AO�i��`�~�!��	 �&��"SeY�[)T��l�����$��Z�J�r�lq��?9�R24�eD�A�'L�4���&	LT���$L��lĻ�������Pr"�N��(�)�d�t�0AjRf�U��L4>�l��(0�����9�$�t ($9�� �Z���S��x�̕�ŧ�@�5��1TНd��p;����}� ���2����zm ��鑛U�a �-~�x7�� (���%��� �F9b�OdXqg �C�&���E}l?�_��¾ 8R�7�
X j��3����u�>����p�Ǐe�c�8P?�k^ ���.�� `N�d�/� ���I'� 8�_�p�b` �^7sd�~ &���[)� ƚ��.� g��?�s�Z���;^��������w�I�r���p�k�5� �w �_�h��G! ��;�� Q_���mf2 ݉�R�U	>�[	#� Yh��2����>�����ŤH Ԙ��߆�w7�?Ĕ�$�@���:��n>�U������o2�@����;���d3 Ƅ�r0�Gh�B R�c���V ��Sj�d~� ���t��x���pp�;�+����$.�f����A9qd�]6�� p�[�œH�����iBP`Şd Pc2'Љ4� �BrY7� ���%����9���v�� ��Qӿ� �D�+��F7�d���<C%hW�ՠ:��_8|�����þ`�@�C_`Xy���Q4��g`�-eɭ>먀3�����<<� �D�=>��w  dى��м�U�1��t ���@�F�oYga�C��)0W��u� k~���5� ����ֳ����(� �'�j�=-& z�e��>aX�x �?-�L[#��r(��+H� >K�XYuǩ%��.�~t=Nl��@�k�3e�H	W��; @k�W󋝽 �+�A��M�0z� T��a��~�+�c b�6�쉿� p4��
#>L� �gn�U T�Z�+�]A��;>�$u0�|#a4�y �������@"��B��c:��.� ��,U( �Q�>�� �'�z�tE/ ?Z�xկ��<d�}��%�jBv� �AFߊ��V \ƀ��E��[����-tN� � a�#� ����m|h ƞH�߾̡ +Ԩ�(kc ;�`g�~� D����p��ʼ t�qSG �$x���I ��A���� 54#
eH`���^ 	�ل��~>ơ�Aէ^ �#Uq��4��k�*̰�:� ��W� �-ƙw2�} m�&;��g� �k��x �8����� !�9�JL �|G���� �� �7yu� '��=� �x�M`*-�� ǻnE+ƍ;L���tFJ�`�\ �k��:�` 2M�7a 0?��1E�t<{� DL�Pl�64 � �HC�@�3��E ��>d	bvY ��T�Đ��^E8� Z�������P�0�G��B/� �c�E����{ ��`9�y̲@UE*����s��:� �X!���Ï �I��.�J� �-�zǨ)�?/
��1��_��@;ա .��Wb�< ��n`����k���Z\���o�J �<�(�3%��[Qʹ��u@�qV��@��[|�\��!�	+&�pM�j5����2@��y{��ϮD�@~�� l��m�M�3�����˞�%���R.8�o�t`�ڪ�3Q���{� 6]*e���� 𱻎C�i7v� ��8�� 2nM'�<7ԗ\0( �bu$#��E�Ӟ��= J)�2��i ���MƮbX�h �G�y�0�)|�-�$'CL �J�l �b�* ��a��1�#t,ɏf���Y���b���}�H�9�������so �)bD(d+ 	Vw�HLgᒣ� �8���=i��E�?G6dVIp�S���p�<� @*P�] ��E�bF�G��R-��hv� �K��Sb�� �nc'dJ� �"���kb4�� m��o���h��bK����ft#"������q� ������i. ��b�wg� #}�aEP9�� �l��!c*�Ks���k��$d� b:�?y��)�� � W��0���FX*�?��|g�L7�h�� R
�*}������ ���sӆ"Z���*BP@�PeP��f�r{љv�  :�.�,b�� 9d2�B���ɝĠj�z(���2Vfԏ& �i%Mյ������`�35y�\*q!���bc}�@
���Ġ+�ۇ.�5��	d{� �j3�T�%O���)��h�*" 4!Vtc���=��O���(���e�=���!� �&b��� ��k*.'T��	�"�5 6��8 
d^-F;K���(g���7����_���^b�|e͎# ܏u� D�	7*=� �j��/��� i�&��ȕ� �����b� �{ۍp>?�u d����O�Y #�z�V*�|�?�Ύ,Fc��bw X���!l�
#zdi��@��b���tG �7d'�����h@���R���R4� *��M��b n<��QN����@A�^���ܾ�k���.a��W2�����9ר>��� :	`;di �c�5�Q���Y���@~�>��c�`�i�Y��* �y�p�rA) +?�7�,	���;�0v�����7&�F"��l��~9�a�� �� � L�Y��*�<7�
,$P� �Nb�1;�� k?c�(:�� �0/4��8.���:�a ᵷC/� �n5��)�\"� �h>��kf l�.��2<<�=	��Ŋ�[f>ۀ��d~%_�\UI�.���i�B	 )�T���_uU��0X�9݆�}Y��ٜ%p( ����m��:wk �a�Ӡ<[ڤ����: ��sqlSt/�dV ��{Ac (���ba�.�$*�^���KP�)�����I&�v� ��;?��H9�Q� Gl�U#�x�=�р�ߪ����� �_�G��a ��s����٪2�@��� tn�����c Yd�QG2`y'p���r�[�q� ��`�9c �"-�j�Q�� ���9��� �<G?�n� �a
Ki�_A||å�;@��6� H���[`3>�c dh��V����V�j 4�T��&~��n0����H Ҫ��q�= C�2�:ؒ_ �L�n��� ��zc�`�� �w!�����IT �n��8
B�@0ƪ���� ����Gmz nJH�`IC �tO�cʟ`a�鱥v� (DY`�n 9��>��[�f��̰r7� 0���.&'a ^�Ucy(�:8�
 �4��?l� �����c #�z�^תv��@���$`�ʾ��,c,�z� ��G1n`{� T��x�aP��@�:3� rX���v�4 �]���ض����`���5
 3X��c���= ţ`)�Q��aO���P!z��p<:����@7G�nR,:�`������q�;Q� �u���5#��I�@6��� fg���& �ʴ�#+(� �;��nfyH;a����D(�l�`�9W a���Go* c�߁��!q� �n�	��<��Skr����gQvI�"�D9�t�)�Ƴ �
���aWШ#�� `bEl��0$,)P ���u˶�aN�`�+t���D��� >5(��Hx% `���n���v���;$cE��󄃞ܰ�ͣ������� ����Gj� F+���Z������OΪ�@P8j�k�� ߨ|-�~a	'��`���w�J��⥾���������� �IeaQܘs���c�3b�O�̠8�L���r�)��ŧ����aٽۥ?�{� k�`T���%r�p�����B�`H���� �&a{xw*
Iz�q� ��>� Ϝ�K6H`���aA	8%j ���go�� �#�]�b�(D��&�n�oϒ~@׌�L�X�m�y�^��X�� f�JA�6� �hd�k]��~"tC `�z{��ް� �������͐ n����]�<�Ÿ��@�Z��c�`�$}�:�� �aq�c�<3 ���ڡ k2�<�\�e�Z-��~�`�� `N�_��V�L��g���(��&��=4}����� �8�:� �cř���t�n��=:0��")�E�R G�JƟr�p� dv'�����~����]�ފ�G��%��̺�,�-�	��L���p���r^0���!P( ��e�U���)��� �h<~� =cR��`�� �-���!� ������ �nV��aY� ��k�@Рj �M��esU 7_P��> �`Dٖ�U�QM.�z�e������+�Xs� ���i�x��%5������xzX������`0�O@�v?~.'� jq0�\6 T
C1�n��4 cN�o� ��� �$Qݤ��WH�h h��`V��m��>���@ ���|��<ˀI��aj ��bXT�� .+���N����`�j �r �q�&XE3NLp8a �����13BpF���^ J�}5����q��< Th6�.��n����Ȫ��=Q>�@�_��"@J�ǠS �S<�!p��x�d�u �bKGU�l�pycs�a�r��m.�� c�)k��,�H(R�U�,�<�3V�� ��)�� ��H-c��fd�J�1����� Мp��:����N_���1I�H����}gS f����} 1�׷Bwǉ=W��9�$$�� O��t�\u6 �y��"�� %E��'i\.kg�j@C�� ��F�f��>�: ����ѡX� �l�8�v���W�l�T���O�hg��,i�)�� ��޴����������_��wм	 ��O��� ��Y���1[ �Hr�g�p�8D��t ��dC�F8� ����T�h��� im�Zg�z(<E�yR �DQF�c+ ��i��'���g��@x� <5�U%O���{�w�<��g9��l��0�36����F G~t�g�Y���� �EW� ���,�rG� !�sD�5�� (�W��U ˜�V>�;a�MdoE5 gk�@��W��vzF��Q��<yI{U
�/Ӏ�W�:��|�A��T���H���ϯ��#�Y�� iX��~��e �8A�t`߶�w�N�� }��W~�xY ,�<� H��]K)3 \�5��Wb�<"�L� �0��w it��6{�ց �W�"����� ���kqFv �?is��V L,�Wq<JXĿ� ׽b	9*���&��W��=Xg�� ��:x�� 卵�4���6p @�+?\� �h7^�� ϵ%���D X��9��V� G5�ޅA���x��W4M���hv7���pA�� ܼ -Wd:���'XY2�0E5 A�����	4 9�W�����=Z�|x| .�!-r, 3yH���?���8�;X�P� y�����@� I�EˬW� k�9Xr}��*���!�s �L�'#��8 ���W��!�Ϟ�f����� pJ�ۥ��Wr;3XH2vЯ�{� �b�?�T I��'J�j$RM���gNͿ p�(V�8�[#���pHz���,@rՌ8�N�s^���4������JX� zU/�F@K���Z� �W�s}P���^�2	�7�A��� ��-fw"��֫O��1I��x]���A��UD G��/3�� �����ƈ:�ߏ��X�@�xZ�l��=i���} �F�lVt�jU*^���}X�z� �����`��@*ј(�a�/�v�l�����ߨ��J�ۆ��qK� z)yLB�+k����;�P���Z ���lGB�� ��g$6�Z4��'��� #k ���z7�C�t�E ɓi�؁��<%�*H�a,|���1�?���.�� ��D&>���Q��`�o�'� ���C䲐{�(mj�2R�}��� �N+ۑt���0׶�x� j� NƮ�Z� 2Nk�a�>B��������z�@(����(B�	��y ,!0�cG�R&ZI�� m����	d��� @*0��!C�P���QՒ �u�)�I
k3!�?	ˈ� ��h4�D<I��4yJֈ� N��"�̈������S�Eз��Bޔ�N��>�\ ����C�x@�R �ıt�*���8��I��	?��T���H  x��=m��AAX�lS���35T �Eф��?<;�|��;q�Q����=+*�`�#,G�xg(�*)+ `���4�B���TC��~���>R`���6
�{�����D�,{��1�Wx ���@��y�BO�@�U� �@����f+�"w�<��b�5�� �N|��㏗�Q ���"��>CF�X�9P提��R�W�@��x��!TSQ�xҡ������WΛ� BB�1��[{�^ .��N�����bC�W
�v���J�_������,��}
�(D7���9[ w��w?/�!㖜���p�L���
�G��@�	K`j�_C>W P7�eT<
��8������,R7L�(�>C���i{
��[���:Q����By�U� u7�V�|��  X7�.�C�F� �Ub�x`� ���+�!A`@7/�E�DE�@k�x@C���U�r^ )�``5��D�E�, O��@� ��G���6��Ξ`:�8	s�(/�!G�0��Ϙ\�.����9��8�J��A(�� �/� !Ε�ǽ ��πB7kFY�׼���@�Y ���|� ��C�ߏ O�[��m*��H"�8	0�A ��! :�d�Z� ��7Q>E�[Be^�-�Hȝ�?Z��V��p�C�X��r�8��3��5&ZU0�A��c� j�D-,�;��y1/Jh���! >h�z��� 6f*��m��0␀�3'P���-��ޘa����˔p������H��t��@�_�0��kj`�`�=�U�6y!����ڴ���X������1�1B���K���d^�5�`�@����H:L��30����T���2�4y� m�� ���Š8��?�2)Шt,�'g��0���N�a5�CHOP��{�yI������m���ɚ�����4 ����<.�7f���c�A$g�1��9����= 
�@�υ(*`P'��t��V���G�`�B��;D|b�"=a�ܿ"�L�`N�����8 ��(���(>27�{� ��aQ8��8��:ع���i��*�� 8ʶXȢ�CA�� �6�hb"Ѐ�$�p�$!v|�x&z�P�B�R�J��@�co�X��ĉ��	m�*�Rl��i6�Ձ�<J�pd���B
��h�kn�������XL,Z&��7"X"�����4��1�1������p���o�A0��*������~�S�;�Ԡ�p�lR��t܋�� 
k!�\�8�3��6]��[��I�\��k�+t^ic($`4[٪|nZH(]�HJ�#0U���i+'�@�P�����1�l�� �H�ñ�_2�^���PR�J��\ jF���$ :��ɹ6�9\� |m
yD助<�����{� �Hs�����*�r8-�P' ;��O���e2%[xb8�G����X��dMwt�3�ap�FEs� ���p��$o
1C��;B�9ZB7����P�M��F���E%10�$��r`��q�G5w�ʚ<b#��L<3�ĎT>�H 8t�Sf%$�:�#����n֦�G�;[!f��2�8�ۑ��<ݐ�ȭ�3���2L<�⸔�)�#h
���d�q�VRx��Ј�B�#I��x�<�2�Hx��c'�<R�0h�xY[C++���b�d�q��B�<!�x�3��1�!��!Vّ��?Jx~��Sb��8�܆S�<w�َ!+R��ň�A��ӽ0�)�C�184�����)��9�g�P�Sc0�w��ӦQ 2eNص`$�C����U݄��H�"��`X�B3�$�7�#	�9|"�� .$ ���Uj#�/�w
�����
�YQ�:D��(��? ���Ʌ���X� �d,�˲1�0*��<�{ML,�@\��Y�6��8�@#�� ����5�"KÈo�ͼ�`ӧ*��xdS��0�Ѵ�AP��,��,H���윀� ��C�!	R֘T �;3�ӨT����hP�Tf�����
��M0��yŲa(:ּb���0�؄�7#���v!�-�@�C��W��<"�3@��:�9��
a,��0�.�烖�:O�����)Ə���-��H����T*:H���N�hD� lR�Q���̠� �@*RKx
���������O�}�/�7t�'2��)$����v���<R*�H�$�(
�91�^�`X�0w(0����Ѵ!@i�
CB��W� ��e�"�iK��^|�3S�(Cv�`6@�
����4�� ]�i����`��XDL�t
�
0����#��Ot(����'[��*�q�X�`SX	����P����`߱/�|M�x)�,	7�1��@�p�!�e�+F��A�x�:�$-+L�⌷TH��i��@��N��p#�0B�EC*���-&�����Y�x,�p:�1�Q��5��#L�D�xi�&6V�`/�i���f����[ԧ,�i�n �0��Y�O��D	�!
�*\�e^ )4��zD�	�Y�O8�	7��-�2�H0��Y�)�`$$XQs��@AP%�gtێƘ;��Q�9��Lz�	�B���OC �6N�����#�lVOԦ�:���=`-D�	{7��D�xyP�O�evr��:P��������6�(�!s�8'%�|�<�Cd �"&MT�2Rpr��0B� �UB��݀�V$"�ɨ��u,��|�<(`D�r�M��af� ������x�< -���{�"�Iy�H�&�P�
�!�����9(|J�[]� 	At`��o@�3�9H�p|��X�.@�˸�D�~
�L�ͨ�1������=�%`�(��XD��I�PH�R4TUR�P �f頻1~-��V'��J` $��%d?PW���������R�M�7<, \�z�wT���j�|	��DN�XLև��2(H�h�d<.��I��rb� �±���T�q�ːe�"Ո��>p��;���.l&FզA�� �7���'�T�ش�8詠�V���&R�8��$�l�KQ�$�s��2�������a -3�(iT\���
�P��\��ڌp�w�@��D���Dl��Bi� SD����5{6���܄"a�Q`O�נt���%o�1���꨼}᠔�q���؇M�Hww�����OF$��8-�.P��(�l�%f6t���D2>/���5�1�'�	4@P� �͘�oW�0`#��XG΂Rl����!?�E���U���6�1���C�DHT�h� �I�}����J�p�(jh��`��O��f��n�/����X�pp$��b���� a�Ǻ ]a;��f@8-M� ������P���8���O��̺(`�0@%�K�@�M8t��Re��"�/$2TR �N'Ӊ�ht`�U�(��@��<����"F�w��� t�╖�y��EN��y��!�ԩ;�d����w���C��ʲ���ܠЖ��O4���~�\"#0&�x��!H	���r�  ���T�ˊf��qB�c@0���!�I�
���G(�.M~IH�D�Ź ��^��?�'!��D�`&#x)�! ;��HwL�#q-D"�2P �|&x{H�a�ɝ���)<h̆i��"%z��͊��R�ز�4t9X�LB�N3d]�������)�TY�L�a�Y�!qt"i
�"D܄�'�ۋÇ"����n� �E��3?W�̅R�c����T�ai�x8Pŀ�EǪ�*�0C8�����TNG����S�QtK���p���2�H���[�4��ؗ�DXx�)��Cq�3�������*������)3���z<M����d��Q�s U�;��8p'��%�<AD�B��!t��Y���&eT@1a���XLRZ����H�������P��Q�C� ��U�p}� ��$>����:m|��Hr��i� �����5L���U�'���� ������� ��:�s7���4b��h`�!r��xr�!T��V���~�®�`��)�6�(��һ ��eC�B�lH�(�?``+�� m����r'�`� ���n)D �L�0j�r� ���k����8� 2L�3��lI>�L`�:�a�Hr��p�g�!��a1��+��| יL���D� �[iJ�e=8^,�x�d��`ia�#H�� �qa攃}�� �s{�A��)︤�'n=������3�	* !��82x Vu�%�\��}��р��l�6`�@>ş2iK�B$G��!�62��=0A�����G(���2�K/�i�|��_7 u�fS�s���R���B�N<~�	|@��R8z�5����X� ��&�oaEW �t1c�S 
�R�է ��5,&-0}t��;��  (�]4,r���񊉤�N����� YRg��Mi2���� `�:(�� ���uM�y�i�e�2R@JЦ- �[�t��� �M�+�;7 ������ Bت����%E~nN)���H?���kV�I�З�=K.b�e��� ��{tǐ	�����Yf��I� �Ì`��rǯv��@ђ�5 &�c��Q�}  �w�4������5��0�����B �wk� Ⱁ%x��7�A� �Q"ޥr�\�{,�X�t�ʑ�y�Ȟ��&��f��X��'�xdG�]*���R��q�K;�s��l�E���:�� ��&�;��:sG��� �� t�{�� <W�
>1q�t�����9>�Wn�w���5�`>�	Y�{} �b�~� �F[/���}�:���wWsJ��3 �d������-��̇���.���騧��ݪ@�$#������^���R �5�=M��:�y�� $]�(�|�@��| �0}��(>�� �p�閭 �B]�x�������W�-�0\��p������=�0#X4�M ,�]�լ�(H�4m���sl��n��Ń0i��9��@7� ���p���lѓ}0�� �!���8��:޴PS1��ϟ)m9�R�x7����C�;}�Н| ��J��G��(A��@�����Ա�r�a\�0�KW��p�}� �t=�H�H�� ���BOs��� �Α5�d�r/�[֧��P�&��
�P�H%45; �q���@���ݼw�-9���`@#}̑�ŗ4�G�6 �ɶ�� 9s��[%�A���ʃ����;+E�n�j瀓3�! ��9����f ݨ��#z�P� r��Q��ˁ�Y�聠��ڪ �ݸ\��W[j\�A4��.��a����πztf�j:ד Ӵ��=�7$�D�(���/ ��=��C�ѫ�@$�����s���]�= -��>�� �h���'&�K0�[�Q����}%����rU�nx�,����xI7 %V��&8� �����;ӱ����]���H�ߐ�.I3j�8���׭�=�� �T�I�2 �q��L�� ݟ��ug�x|;��(��`�,Nb�R��T$	��,x� S-���|V=��$�� (垷8�&��(j�%P��,�d�VElf�������ܕ Hv�Xe��:o��p�s���,�60����$�O���0���
�S���¡����� �@&�a>��:X� �^'�����E0���ۂ�����^�� �� oS�Y�T�RH��P� x����'�X.�L$h�b�q�7��i��5�Ƈ�`j���,��	5��Ci��ݦưd �,�P�����dT�-������(&ᅋ��@݄��q����1T_����G� �M�eIU� x2���v�LN' �<�5mK���X@��Q�+�����L�� ě�la�epp $�Cd�(U��@���� ���|����$�������@���$ ~�� ��j�g� �1���)Y����L���ZӋ���5����TmQ��'-p�`&��ϊ��� o���S': A[.TR���f�v;��/���iT� 5-�� �t�I_0�� e�O9}���:��2�8 G���7R��P���� ��ۧ��/�� �J�<�d�t�C�ډ8��Xg�ۗ(��G9'	��$�`��P�HY�`᳘�uxI&��(��x�L��� ��N�hIL �e��~hF�0�Ƞg�Ȁ��^P�k X�9�~g���R$����N�,����'?�JKXĐ�w ґ����,p`Q��O�b�膁6!�w�|*�	�� 4UL(�h���P)�������}/@ ��� �Z���o���]R�Y� �`ܙIy S��C`˺4`~`g@P�����S���N�����G���a�}B�'� >�X��N��D�7 $�Eا� �\���P� �.��� �#
��� �;�E���B�~^�����g�Dд��=�H��(=��z��� |
h�,�%�q��4���p��O ����Вx`+%�H�q�ħ�&��\~��=69��g�(8ظ:��=�BF��ج=�l�ݾo6p�&�����| "�/jW�P����qu`he DL�k� ���9�[:��W̞h ��!�LCM1Fp�4:>��[j q�� �	Q��,��i EoJ/��uXb���D�� ��LpY�֢s� ��� �S�I$� �YM��How�>�IV�C�1��g�J$���|@ 	�0Y<�$�� ��Lo���p�O�v���p����@=�qtP�7��e;���	��@�"P��0�����i�̧m��� P���*����q� ���p��|��,C�P�]'I�پ����A����Z$�ky��Mt�[��Ғ�T1����Qz� ��N��ǁ1�d���m]( U�,LW�t��k��n4�\�0*� �����7��d ������� O�f��G	�ި�qzĀ�P�D�1� ��n>Z '�W��j����7 p������?��]7�@h�Qy�	��6"��} �� ���<W� 1���z���0�hp��(5��P�dWԇA�)�o��,�8 %�ku�xCZ b�6�������0,_a���xhX 2Y�t\�	��.��V� }j�?́�NZ�p�Q �,$���ըP������R��cd��i_ �8���� �+tW�H� �*��� ��8)����=A�����,,�@ܻ�Mv ��	��J�'��E#����$:Is �k��"i���Ѱ L�n�\�H�� �f1B:��	����(�#�� 8��<>��oh�3�� !(׏ %)=О���|� ��@��$�k�<�J^=s:�� �`o�� �r��h�$0-Eh�: Q�Z=��#�l�>e`��	���2�Z�H�c*U=�������|(��� @�>��B� �%�_=��=?R��I���5�)�� ��bkE=��\�pD_� g��0�A�>d����j�
�8w&K�Px�(y-�ƭ ��3�J=�� t�d=|� �@
�]wI<���>nqU �=9��M��u�rs ��*Ȟ"�O\��W��=��:���(����It��m<h�@�"�/ 5=�Z�N2� �tw�*��nB^<�� �@�� #=�fw�V ��&q)�/� �3li2�P���=	O�Bq x̦e���� �Sr5(�o��9�X�����I� ��E�>�~���Gm�p�;N�H�,=����X-8r�X�(�.��� ��"uG�x�]���
I��� M��j�� �A��F=fs\����j��>#�+m��)9�r�ty�x�<�9�'�)[. �aiP# �S��'= -��$ w�)����"��r|p��Y���8�����m�bx��#|�X�`8Q�6ŨS� �r��c� ���q�c50��W�� �N�<��)?�����*(��c-A��@�l��U�@�w�'0|F V医��
Pr�� �ړ�(%+$*�P I�a�r@A�F�>^캡r� 6IYH)߰� ��5��gN	�yr ���x!c��'q=�� T&�,���	G��<OQ��߯����d�Ќk��6ie�� ?Bw��(pgW�ACþ0k0:>Me�{��/��	 1�طQ�% ֚�n���d~��A
����4��0�@G��i������"�@��B���1�ᾀ8}eׁf�.8��:��@1�u$2^�ߎ�/'C	h�gy�k��{|^��2 A�Ϲ>����@i
�ъ�gɝ0�������n��!�h�~x� �w	c�� �+�YFS8� �[����ھʞQ��C_ �G4��� ��a�@c[ �ّ
e����s ��4�r�h� A��
��� K�^u/�� �p\F�9���g��� *��,�´ 0:T�3&�}��I �h�� Q������j�v�6W� Я�.�>=��>d`�v ���"��Бw��2� e���
1 ���Ȯ; �����c�: �y3��AC q����T �-�0'G��(�N��m�R�Z�;Sw3����.� ���?� ���SC�� )ѿ.�]- �P����m���u ſ�]� 
_!� ��ܩ�s7���z�x*I[��-hD�ھ�ce�������/��U�����\�?�<=*�v`�1�@���ϲLP�z� :D��ƈ��\�t ��.�?��0] +���3����k���Q	��׈!� �?���t�^��%p��b�E �<ik�$&>��ߐ�(��4�]B�Z����ז��pR��Ơ1���ЛY �D��*54� qo���? ܑ��0�Ol鏨֍����V'��dHl,���
Z�����E%t���ת$��: �ܒ��@V��r�Q@����
i��"���<N@�E1�O ���� ����&�;� yGS�%�M@P�6�����0>k� ��w�˾o�v �uJl��N��(�?�z��a��\3�4�x�B0&��� ��F������0@�i���R�����@��W�z� ���:#� {���2M�>H�� �(��4� #��%�2vީw���@�ģt��%�l��O+�, an�Yq��:��@p���l;Q�Q�1ƀ�'x_ ��i��	�Q\���� $�d�c{;���h�Ԑ��� �	���i�� �|o�z���X�� &l�CVڒ��v��dS���8�� ���6-\aYD)�2༡�0��.�a XAq���H>% 	Q�gHb� ��OX�$'>�H������s.��P ȃ5��(%$���ꔟ����Qޠ���qI ���>�l�H�׊am@�� .�^�2��&�jLPKိ���tM���+h������x�<	��� �~�$av�H'�����xA9 ���ݿa����^d8�Y$ dT�윱 �q���� �m��9.0,��<>�P���^� QGX�u���$�����9�T��� ��W��z�ƣ��9JMTI�.�R�֗�kD���{b��V:����_,, ��m�����M��l��(��ȝ�������)l�
� ���Y�P(���:���&ΥT�^8�}_a�!ù��M &�N��4������$bk� (Y���6�����FU�~���ύ	�n� P1/��� �֒�	��]l� d��4E��O0Z@�����dX���h��� #i}�kF QE�$�u���7.���(�C������r��j5����T��Cs�N���;�tA t�)��z�� s����q��X���������� Я���m� $�C�ab��'���E�q ������L�X.�~�}�X�=�ڼ� �P�q�3��������a���ܿ�_�`(��"A�:�^ �|�t0 �a!��Y� �[d�c��H�o(��L�<h�"1i�jC�y��p���0�X��Q �G��/�g�"���(���A����0F��1�%��8�s� ��!V�(
 �)dJ}���- H{�G5פ� ܕ*#(�8H� ��<L�9 �u�7�d@ڰ� l�ͤ�*�tw �R��-0��im J܍Q< �Sh�{=�� >N���k���!@�H@�G�r�S�N��p��� �<�ABޏy!���-ŷ��?�Z�\���Ay%]�T ����� ��b��٤�0�Zm+�S� �H���,7��;p`�a{Ak�Nf@�����2?d)*�?إΤ N����G`=Y�r�� '��xo����awf�F4�1��K�~��c�2��� �Gj�E�-?�70�D&e��č�H`�žh L�>CN��a c6����Y�$��`��uO[�����kK�� ���	ML�t� �wh�G-i��*�bM  �O�k���A� �����Y{2�0��<Ϡ5h����!t�o� ��\%� �kZC	P�L��.8�� Ekg�pAPfI�! ]koSd��$P:\�Ԗ��D��O�@�������C-:0����`	� A�x#Y'
��F^+ϣ5ϭ9/���[s*�u�j�`K� ��V�|0��lO��0�э�	!��� Yr{�u�'=�P��2�	x���R��͹@����>�P�'������ �Wߨ�Hk0�G)#Z�� ���A���, U��z�W�J��)H��p������ �;1I��8J��ȍ�g��'1�@���� m���ix.�<�� 
W�K����?�� �e�Gw� J�D줩�c�6�ߛg9��FG�T �_e��V�b&I�.�R�o�^��� @�n���)����3�����F ����B� dq��u��T�� Ul^�#:0�nւ�-�@�} `�Dq���Ir� T���O�j �G�����S <|�DBߦ?O���k�G��}).Y�W ���]V nHů��?������dy� �"H��T9c �=�!v�r k���)��� uF��.G4��e=��9@��*3�.7
ڷ �)P� +(?�_ߕ�IԮق�s� О���i�+!���/\(�k�F��>��}��)�꾀���G���R��`a�{ N+��Q|.:b! ��Y&`��HG�nsU�dJ$ +r.��)�� ?����v# ���pt/&9?�M� ^I+�0� �E�7�����b�n�ݷЇ
#�Y���.p�A� ��n0��Ϙ߽�Qe��=ZwM� 9�);G��]��0/ߌ��4 ?�g�<.+~�񏾬G�����0d� Ml��E��_�HӒ)J���8�� ���V��~�&|H�%�G� P.,V<K}�=lǿUp)�T �^�o&H� i+��F�/ ��X����ֈ.Y�y�G�x; 9�q*�1&��W<��[@�@7�.��F�@�������>^f�9��]�	��I8[7@��o�L��A���A���(�s@.-h�V ��Z�������a�'����H��) �gMk~��	q|Ď �V�u� <���G��0�kcH!���z�� A��;�n� ��-?��|+�l�����G���T ;0�� x�Q�.�	��ôs��d�`��� j^�n��V* �d+�����Z|߾?�@.��4&�L �!�i�)�oL X�2�$��4Jp���(CT�� ������ ��)}�O7� 2x��8�(��$�� -�c�"� W��S� ��xe�)4	��Fp 4�PU])>C��� ����S�G� )֕5+�� aV��	�H� �$Nk�� _�yHѓ)�LD� �./��g:�� l�ڈ�x(�G6p4_�.L M��]u�HZ��#�b/� r�G�H���olh�%<���������e�M�y���.�`�WL6)9
��ܛ�}�5�+n��".�Y	�)�^��E���h� =-�>�x�( .��)Z������8p@�9ߺXӸ&��1���'@To�s H���R���P�� �;��7x�).��L Çw��H V�"�>[�|t;�q��E��@Gǰ� &ӿ��	�������GX���	Ģ l7��?	e��l��>3�yT�����(H��)$[.U�C�8�� �hL�9��?+;�O�gC�防J��T
�?�ӏ��A,�0hYP��A|q�<u �.���)�U&��z�<���W�p� m�-H<PČ� ���%�yf��)��(��w�P��00�| ���' O�X�1�0/ߨ|�,� �ܑ)[�t������S����c(���d��)K���-T$XH0(�D�M��)��92�X�@��� �A�{� �2
Ζ� /�I�y+��Cc�8@�Lh �i�A�> �v�=�)Y t.u��� fl�5�g 7)��.�Y��8Hǀ��?���!ܜȉ�Z��o\0L���pm< ^����7��e�C���}�'Fr���/�s��� G �xP�f� �,��Ӯ%p3�)��-+�}�Xj� l���&�	Wܱ)��@?�<� ��zb�� s��u���0��J�)2��� �H�]�~Y�X:
���	����@�?.^����&��$l䓉=U�X�k����� ����"[���%�E�����u��J�+*?�{`mL�}� ���_�x� �)��+�D�<L�O�uH~@�=9�k������AX{���D�`DIt: ��o��G� 9v�R.�  p�F�~]Q�&�5L N�y��A7��)���H�E=w�5�!��ߪ8���%�H����@��� s+��8#�C� ��~�T_�G��.���`����)����� �nf.rIy.m+u���o��*`�f�?hw� �J+Ÿ* ��S��?�l 2�)��
��Gь����{�*A�'� 7��9��0[b�	���AG,"�f&� 7���WL��K��૆( w��Y�]��~�;�����) �GB.V�	Tߌ���!�@�k�� �iZձ��z����8=��4��	�LW�����!<#( ���qscZtߝ�ˣ����ʐ{e�:�� F�k+8��� Q������\�DF� H�+�`k R�M��ƨ-߸�t�/��c� I�!pQ�i�Y�/@$�w�K��=$r� ;.�`{R��X�� ��mM �n�7��09.g�+G�@kM�ְ��H�lL\ 6��w�+.$���=�Q����p\�s<+�J���b�F�xzG�4�2:<�i&_E{�B}.��j+H�@�Et� �/R߭�p�n��L��� Kc�W6����)*��l�	��Ǆ�hvJ2������)�Р��:>y \p��4�����w@a��� t8.#���� �h+�����Ց ������ �
+<���>X�� h�G��
I����� (�t��M ®�̕�z �0Ґ�?�z�	BG�KP]���İ>�<U,�Hp��@|��� �*����G�����)��LF^ .?pbB;�H+� PJ�y��x�VGo���S�.�H�?9f��Բdx���1s.�nQ�R6�0�� ��G��@e$��� 3˲]�� �VJ<��)����GQ��D ��xBN+?��)"���\��~p�}@�K����<�e���ǡ���ߨ8�n�<p̦1D ?��G9��X� 0Ԡ��A� �ajߥ�?� ��b���G� @.4ʭI���D���`0�`?ݩ�.����)s� �HP3<s�,^�d {:�ڰBw1�)�ˀ�R��] ���L�ߗݠ������.�(�E����>%N|��T&�� ߦ��P� )z/��GM��_��@���}U�46y`)�ט�7G^p���kJ��?�7���&x�\�D�)Q�@ܡ� 9���_T�\ �g���B��� ��G��.� �+[}/�e;ߧ�|@:@m���FP��� t~uS�&�������H��)U ��c�|+Ḙ sG\߄y�!H W���T��������o� �	�ɨ<Ϝ�i���(���� ���q^tc�W�����}�0�h��uwc ���U�Tj#=iB�x��L�� �c�F�{H��)��A��^�&�y.X�� F�C�c�H�/eqH�S�ɛ��<@ܯ����)[�`�ø�����<���@4v/`����Qz a+��u5z_W����9��1~o>���)q �xK�_�� (G<C��<�T ��������Ԭ��`�<�&�7��aL�0� `|��m���}�$	�N��$����#t����oH��/� a Ȭ�X Gp�%&�Z. �b�R��z��%�����)��	�	#�l���Gs �
3�M�7��0Ht� W��-���l���i��>�?je��  8W.��x�
����|[��Y�FpC���+� {l���ָį��t^]G@Me-�(�aX`��G=�yR� �1�)uz	�?H� ��_{���LɄ.��<p	�e�( ��q4�P%��0��/y�9f@?ߢkN ��K�z�F��)���#T��	Wu�.� ������a`ɜHٴ6�OƔ��0�k� 澡�b��ME�' dF?��j��&H�@T*�\H����{u��G�� �ºh@� 0+*Q�(L^ ��r���c���pL�I�z�)�Rp`|f_pU0l F�о^g1�)K���X�ےG ��-]oܶ �d���Ғ�	��)q�D͔�������$* ����)F��6}�0��O�����R�|`��� }��\��GL
� djz9���wH페pq�H�@-��I��.�0Y��0�Az�XUF���'*��r���Z)��Ye"��� �,��)r��X̸��V�����7�X����GrV�6���,��p*$��J����q�%OLj9
GS���; �!�㸪�~�gD^T���9 ��Z� ��嶝[OHj���� ��� ���*�� ��[��� i��B�� nŘ���8�$d�O�Q ���6�9� (3���q �X��EĘ�اfG�N`p)
�ΰ��H&.,����H�9�~�w[�0 8t�矓���G�S� `�|/.�-'��!�7CF<y/=3���K����(4��c��3>���>~ܢ|��� �Eo�QU�5��T(ꁺP�a��LM�| �)�s�I� !�S�|� H5�s��� �E�V���� �
w�a��j���S�� 濉@��>� Uʙ�x�P��`��H�v���O@��R��� )P"�3���;�_�\|H�F�j�<�	 U�����>Nێ� MLBh ��W��.lq�"D���ۇ\è�ުy9��CAX<���;�� ���ώ�GV:��\�G LH�� �L��j�l ���DGr���N���3��,{��u'��}�/L��T� G j]X�ι(|�����i��)J��-��� H;o���N<�_.��ɝ^��T�H� �� G᪩����ݔ�?,� �W�)<�
��Z��GJ�En\8u��5 �v�Zk�j�G�4	��n��4)g���; �luDq/H�$��T�] �v��������nlo����H���G@)Aɨ���<tz��@
�e�p h��ۭ�H)	���� �0��[P��B��r(��>U2 ��G]��X[ H��`�c� �i6F�2����8w݃�G!��ZؾP�|���8�\H�>,I��� lǵ`3�&��T �ү��F�eb�XݭRI5T�x*�cv�<�3�kp8�� O��@G������?^=Y1K �7 �9�6�oyXzI$�.� ?Fr�� ����xA�h$a�6 /��G���H�@S�YNc��=��f��y� :� "�Gl>XD �tb���E
������S SjV��~G ���%��{9��H� ��+�����]��8���F�X��]��:!���,Û~;���G �"��f���|�-B:��?k~��o(�H�� E.�ٚN��:�	(�S���� `�_9 IW��V(o v�a�kЯ�Hb� )_�H�q� G�9�ͯ�Pf�+L�� �Z��w�߫,t@(y���;D�<�@��G>K܇0?��:���I��W(�ӭ�|��@�C�����. ��?H�&xG�����w���j>m%��	I� P2{��<���hǐ�>Q�	]����Kx�|�ՋE��]�<�\/H:q�@!D3��K@��)T����=.nP (��A 0�@��O$!�܉d9��eJ lyf|4 �Щx?׶�(	Έf!P��ڀ�GL�a�� �)�3l4�p�7S�8��@ w�G��*	f�>�`�� ��Z����V. 7#�l� �� Q�p�����d�o����_*y�~�H.(���G�x|L��8f�r�লx���� �0Oo~Ӯ;�Ҁ�C�K�Uiv	)ג�h堡'ڎ�c y���ߨ(���<M� �Dm�H ���&J)8	��.��e,	�GX� ��yjI :^���K�8�?�����RX�+H� ��/�AF��3倴 �����)Á��sVL ��׺��&��,?�L�jz���k�3���H b�{�Tz �d�x�S����3�$b���G(:�Z�YO���pJ�(\'����^�� G	V�߽z��O��Av�3�$@4�G{F0�$?p&`E�9.m�`X�pkI 1wuC�2TH �X�����WS;��p=�EAr�>�> �s�~� �g�#�� `�>H1��<����H�OR�@��� ߞ?��&Hy�!IO\��liH��X�7���x�O��0I3�rE��~B����-��7<<HH�E2�	�sØ ���L�(¹ �秷�H.�uFJ��@�쯏W��8�tc �MG%��w�H� ����֯� >ѭj0�Z�x�G �*8�]�R �T�2 @�)�ߊ�F:��H��X�C�����`�T �a��6�G�S|Iר�/�WM�T� ����u��Ԛp���K��q����� �1v$���l�*AWx N��`�B�p�1܁1��n@�@���" ��K�Mj��0[n�%��8�� K��Q�B~* ��1�[ �d-��6 
�\��rn� ����l��-�=m�0��%�(�0�c��:��W���ɗ���q�N�@��w� 7U�:ݴ�'�`*�B��}J�Fx?j3ډ��	K���-G &f�A�[�����	X���������#�g��sZ��t� JҖ��X�)Iz�.��06���|�U�p���^�Ԙ�E�F}Ze��uU�T��E�ۄ���n����%���� �bR^��A�	df�ŀ�'"�) �0+Y��� TF�h��)�߿������\RJ^��2�j�#6íY�	�k@��UZ��(J�. $�������ҝa(�!.U�:�r�� 8���6��nO���ߤ��t:}&�HiB.��WpQs�,|�� `���b5F��X�\D��7�~ڱ`<J�B
-��b�� ԥS.W{o��ߕ\�e�<> 
��)�&ə��.���YR�  ��l�Sߪy�� L1s;)�&�R�< ֢��?x>�, ��3JR�}��~ P�+U��=n���H]������7�j[y�+.���)�� r��%�÷�Z�����H}��G ����Y�m�?��$y| t� W�m���v�|�<y� T_7e�)Fi�B�^. �+G�_�߻�GnP�z�- 7�WI�)ƘB������� U�We%.]`	��T P�R8�߭w�d�$��q�� fU�jEG� �)�=[�����q:Ѓ! �'2��;i� j���C��� ��S�ՙ�d� Up!�iSʁ��$�� �	�O�Z�� ���i ����]w�I:k��O��C׀(����=�� �dg�ݐ�E˃����ز��i��H ������� �|�vJ���f ��7x*i p�9�.�Z���j� j�94�`7���i�߸�� �@������ �ע�iU:�^�@6�[a�>�3���AE����:�2 �о���7 נ_[�ea�(!�6t8 i���>���?,���8��j���q#��B�-|���s��'@P��� ���F���i�9�����N�Aj~�s
R��ɐ�V8tj����h�����"�� i��B�����{�>�$ 3�u�9�	�zj^���[�pǽ "*����b� �RjrN� i/��&�1����>���sML���"�l�!��9�]�<�� �|m�f�u�H!ν�� �º��{�iHJrhY^��T: [���� ���?i�:�+R� ��>S�� G�d���3p]u/� 8�����>�Y�ؠ�k~F�XWC���0��@�f��נ�:r� x�8��Y���0�@�� ����<����T|  �����
Sj ���,Q�� $���;D� ��u�J�ɐZ�P�� ���`c~��5 T����+0�k�i�?o������UHA���qpk��w�m /i I�O�2�4�0 �%	�x  ����EH�P8!L������$��� ��w#�P�@ �d�����x�t���q�p9�0x�pXЇ(���vB�Lt�A)H�_Ŝ����� zg��S1$��4� s�����?�P��-��@�z3��sXq@#���(���� {��С�����k9P�X����u��?� �M$���ys/V������W�$p�P S��l��z�z�F��(aL� �Gaj��4����= �LsL n_��x�����c0���ɓ������l�6���u����iES�f������X�{�r()� M|xFI@j�> b���W��L ur,�iC��� V� ϼ���gjzP���
����ѡ�R!�0��\ʾ�pza���#dC[U\L��TX�Giw"P.E�I��� d4��,����8TNZ�����d��58
���j���t��еװQ�:`��j8:��������J��{ ����~�� ���\_��� pRnW0Oq�]G@Z�M�� �ln�t4� u�8����l���
��X� �+\vB�t� ��#� ��A�]���TǤB��i��
�H�	Iˠ��5!|��t:2�H�Yh}�q;��8� ����ǬI�$i1tQ�� �L���y| ���D���hNI�8 �O�f5��,d��y2_p� �D;ʎk���r ��(�,6� ��g�.�� �̠A�E� ��4�w~� ���Q0�S��,� ��@�$���p΃�; �BIm�|�� �i,+?@��(�����Zӗ�P �2M�i `���8a�? q��������7���r��i���w h!u��r ��
��<9����L��2.z(���Ӄ �-�a�nV�)�� �@t� 4oj���UD��ɀ	��� 'Y8Ǡ���Ğ@��h��(� N<���. ��Y�~�qt: <���d�+H� ���' 2n���9@�&��d���ӂ3(, ��\�zw� �btÉK�=���X�70Џ� �f����i:o%&�c���0h� �|��H�7�����0���'� 0�t<8� *���vy��zdƋ"���(�-�_a+�� 5�eb��Y�:��;�.@p�~���~�C�	�n�h:�7�R��w����D�t��c�����ˠ`� �Y�ug+=�@)� ���@z�X%�$�>�`� 탬���� ��M�yC��p��\@����: ��!N5�V� �^v`��.w�x �'����ʩiZ"u��C(p����i��oaY�:�JM%�䯄p�Zٶ�L�#1��1�>�|� �J�����twR�yᭀ��@���I?B�d���LaFt$>�P�������*���E�\�^�V���E����Gg�U"H�S�ʯ���)� *1{��G�j�+���]C�+�
�o@4r#�<��"\�iݏ���� �����Zpd� O�b�t	h���͠m�0'�*��@��P��&�9��x�`˪�C�L�@
���:��=�6p�.���/ ܣ�e�I�r�a;G���W0�8J�	�>�cp:,>u&��P��E�����|l
F�� TPi��t�ĴZ@l��
g�ʀ� ם�$�)uv���҃\�� ��,���y�H� lTipX�Ad�I����Q�����9�냤*a���B9֓��R��b�'���@`q�� +�Q�~o�8����$�� ���� �����X��°:�a���	І�x�=6��n��:�E��J;
�'�p�����p �Y�頛.G�(<�/i��<�y1�89��Y�&�݀ d� �w�U����q\L�P��O*��3�� H�pڛ�d��/��� �X��q��}h���C�@iwݻ��	�=� 2)"��s��LQ� ��G��`�it!���s��)�	C�	���*�H���Zݠ���,J��`�i�G,�RH ��D�t� =n�����	I�h�8!<�����[����M�&�CHX� �Œ�9/ ��D���;�(�jm| ��s�3�;?�@����������B:� ,�5�<����2�6C����
4����X�1�dz '��+�H�{�`(. �Jz�� ����F���.%�(;��A+ ������ .T���N�� ��z*�Z�� ���@/P︧xB +!h�w�� �"��Q�P*:k���H�A�|��P̘�H'itS�|���R8�h�c��]�v#D�C��L���L7�~�������ZP��� MӃ�@��Ct� ��̔g,8�� 	�U��F�����e 3Vނ!�r$�s���:ih"g��� �'9�Š���	�t�+�2�@L���l����g��s�ar�¬ �6��(L0RLH �����O�	�'v��|�;�W�|"�y�`�qëi��6�"�W&���q���|�{�n�X:7 @�Z������A�d�)  g�X!�e��?@;L$�y�ɼ�,�H���r]���L�H� ��[50fR��i�/�t�l��&l ��?���F� ���:�� �mܢ�b�� �Y���L aA!ޚ��(f:�X�B�B��,���ft��u���R5��Y`�-:����$Ĝ� @�U��
]0��_w��S�� i��������ve����df��I �Y\���j�������)�Ka�B4x8�� ��^p/<�����,�� Oa ��OD��� l%���^[c�hط�� t_�ɏ�0�R��\\��Ց��P�D��5�ꉥ�=d mLHzt"��[�p�R`je����9��!oA';V�9N4 D�gY1t�@FQu��\O���"vl����4�� �?j��i2�۬@F7|�-ef�<�� �i����1.ٿ$ �t�U�� -����� �yX��������P��� �x���� i��� ����� �l�y�P����<D�ܥi\zk 0B��X�/J���:<�*��!0�`��ø�� ������ʡ ���i���$hR�H� ���@�.�x -i]f@��JBĐ�`�sz�������M~_j�pC�8ԃ�av �3���
�������f��N`�o� ��{��u �'��iJW����`>��ߠTڥ��bL(��0j{���&*��S�`� �싣�
� �����iA���AU��B����v2]����r�� ��z��	�{�X�� ��",6i����7��[^ }����rP|� c!�q#̉ ¹�a�t�i�+
  � �Ç��9���#i/�Ē�<ؽ��j��=3�NZ��� -bI|���:�1J�dA��p����i��B�8�z.4͐ǹ¼��SF��B�@�����ZuѰz 8��	� 2�Cc�9 i��j�� ፠o�;� Py��<� @I���iX�y�`��C��}�B�L ���5��x�@��y������@�`�r �� �J(m�����A����d��ha `�i ���`��J�����zC d�;7�}�:�>��������@k�է�t�(����x�L�' lLah��C�i������j��@:.�X 7J(;�� �gz�sQ�� �iV@jP� $���R�&�f0 8���,Y�	��1� 4��/� �-�~��޴Z�`
�@��K7c� �Bbd� 35o�7�^�+� }(gp��>i8`E�FJ����*�b�xD��iLǀSu`��Ѓ�|V	��z�$gw��� G�h����/��00x�� �B�ݛy� �;i�J��� ȥ~x��HX5B*�Tt��A�_���x?;6!�N���	AL���ːЂϧ�Yp�����s��H���Ш� �5-�oj��c��y�q@��L��EM8S`�ioߠ�.� ��0��4�� в��u�+f�:��6*��L��n�D�E�r�D� 0Zsj�٩V�Lד��8a�O�J ��U��H&p�M���@�3�I�����ph����!��0 ������x�=�� Υ>Jw� �ecjp ��𘉐����(@�0~���ň�M���17n��-��u.�7��B�� �bj� �D��0	T̠_����ୈ�\��	�U �yg�s������ �@#r�$����g�k�x��չ$@��zxvf2挨$��. `��mF]sUK��켐��p�\t�����]V���t�0w�p2@Hp�o�m�=�p`- �$*{3.��� A�]}�����P�i@����;������p`a��Ԧ�Oe �i����.\�:	�L'ܫ�C��(��9��t ��YÉ�?�3�r�<��N�Á!� @iIUXk�;�V�(\���tO��e��@�'���� |��c���)�.1|�� K�VYZ��� �B�z��� �T����P oS���a~] �v������ Eg�-��ϐj`i��x>� �m�B��H��u �G�^j +?�3�a�Q	j���Gb0�)5�!	��!gZ0�� r��F^>j A���0�b�`i�_�[L����d�!SW���?�$��1t�� ������ 'y𳿣Ё "��A�� &s9�p%E�L������� � �f��K�d�G-��f$�8 ��ߠ�������|�`q�V�7 ����>(�l�yb���`n��$Cx��R�8޺�& �5��pi$ �d[��=O �M 2����p `�e����` �y%}�p�<<�h �,�u���;@ ��j/֯o �%ㆠ$}L���v K�0*� 9U:�pN\�H%�����
�� .�x��; �ȧ���#Cp��@�s��൯P��: �O�V_0>�?�
�6y� (�Y/D�x�s�>�~�4���V�&��f%ܴ��Ƨ� ��Zq���x8/��"X���p\)Rt���HؗwE4��aQ�ժ�R� *F�p�_o|� dQ���� �c+��i�� �k��pl� ��ծ[a� ���3}�9� p$~���]�p,l&� {�v�S���!H��tV��%5 � q� w�G��� �7`�'�A� ��.&bSp� ���i��% Y�L.���((��M�I�/���q���W�p<�~E,���Zj�`L6p������7 ^���$��3Q�2b��^~�x�I��$R� ��� ��ضFp� -���ġ�xB��� �����X		
��pu��-l�:�* �N�����95"�p��?�l ��{g���L kx������֠v8�[p���%����� P�߄հ�9pƓ�	� ��W�����b��z���J �����t� ��p���đ��k̀ʫQ�i �9����/]�%$������,���}���� ��
���`^�(����l#�b�YP���|�H�{[��'nY%�	p! �Bd/2O�>�Ip�;Η ��Y���p 2dh��^H4(���K��TY-. �%��p��?�Ї8���F��q ����6���$�� �c� ����Ť 懥�9������z�I0�p �=��ؐ�1>PB�č�8�d����Z� �^�6 (��| �ւ%�Ht��f&�`��.)�3�!���\=@ı��b rP��a^qL��f&S@ϝ���ș��x�8����Z�r}�\`�f t���e���!R@�H_&fl���ݯ���߃X�tW|'�p�o���y���b+� $���P<m��p���ӎ� �dZ�����$�b���=�f1(� G�sͧ�{ 0F���_���:��`� ��i&�(ު�� �J.���N�[<jp˸���C�E����W����+���^R�f��%ePU`��)Gpn~9$ΰ����D', ��?%N��� ���o�}S(]x�<')&/��ޫ�L��>�=��A~K�ql�p� �Q%|��(� [��spj�<�M	:��� �������@�q���*/� ��p��q�.x[��>w�6�� ���}�p]�U��L�.:%6�R#����}�p�A��$4�1���{f��'�:�! ��T�$���ǫ�A��	��x(�� )
S��qw��+���̃��,>��|�P� ?A���D�F|�#;\�.��3������0ع �'Oo�%Xv�X��V�p�~L�� 5�NoD2���%\�
�Z�܀"���L� ܊�����u� D��%����@�ޯ� �p���+�Z� �>�ϲMK% �<����q�ͺ�7�(��k�A�ǌz�0���E ܼ��HA,dk�/r��bE8���*�g��� ��apҷ���� ��@���3x��!> �f��������hy؋Ua�ȏ��&P�Ő��3܄��F! ∺+(�I�n�7 @%d}o��q�f�v|�@��ـ�BT��-AH縘�[�ڰ�put��������3�q�jײ��72� �ԫ�b�, �;��Ggq,��<����,h m}��D6��:��`�q 7G�JAo ����:NM�E�8 �R�_�0��-��T0`P��I/�d��i�<��y� LH��O?:F@4����0O���.L>q� o���]ɝ @�^|���\o�_D�s��`�xG�� [�\���2R ~$�Zj�= և�%Æ�� �s��_N}:ׁ(\2�������?�u� e�X�n��f��t�ч{ԯV ��KP�>�= 0S�E�Ǐ ���6�ռ�87��S�p���4L��鳖����=E��`w��C���X��DGaͿ ̮���<{����!Ú=����3���<�?�� S���l�LQd�]� `'E�Џ �G�o� _/.�0����nHp ���� OFTt�Dc �oS���2 �NH�u۴�`�p9��D<^�.T�� ��j��<�����@���sw� �.FRk�fDP$�y����)�l��� G���� ?����a	WO���F�\��n��%�� =ڮ��v�/:�;o�D���b����<�� �d�^Bږ�=��w�ՠ���,-(��L��0�(@��a;	^= F[��v��>���.��_Ԙ�#�зu��W�Bhr@�������x�D�G�S�L�3� �� �o<a�
U��� ?��k�$��	u�� ��j9���.��(�>x�u �O�~�UȨ�@�`0��/(1x�6E���s� �9����l���'�H�1���R��;�&�0� �l_��Wq�>d&�V�jy��� ����<:�X��D>�,T���-#�9���<�������'�J:��8��O�s�j|�`���]��%�x��� ܏�M�\t<����>" d�� oݳ*��p�	I�  ��/&�*��p:�f @ �$����$M����tx���jɘ[��g���d���Ŏؕ'����� ����*��2��6�T����-1@e=����T�����&[p��X��Wo}� ��
Sƞ�� �@8�b�4�|� /��7F�g���\�E�ߧ� �WT�z=�� _��X��DH,�����K�p�%�| �a������5< �=O�ìL��.��� ��SP����Xa$
�&L�/ P]�S1��(9[0�p�Z�6�V"�i��0F�Y Ȏ�T��dL�0Q� r��tO�&<e ��3����z�Ic]�@48s��/⒁�+�w(�������D��76�c��t��� ��͏ ��B�E�l ���?��g� }�42ڏx�;Î�� �h�Y�H�H�,�qˉ��d�߁ܛ�о��)� ,7�9� N�Q���,�2���
�G�Lx��t{��ppv�������(��mr�{|5��p!l@40X�* bV�HE�m ���o�(9 �I��n�� ���x�.��<�P$�� EaN?
��c� d���OuP�\ ʓ���|����U���$a�E�D�����\$�g� �@����l�F ���4\W�
:� �8�D+�� l"5��Q`A��H��N
�ob���ꑀ8d���;�����8�����%�N��I�J��Ս.iBޮ`����H�n� �X�-���s [;I$D� ��Wd�H�� �7�����xmS��[�DXj�c�~��Q�	�}� lM�4� ���)�DHLf�	Ү�
���3�J�`/\ j`�P�<
�L�� �c���_EK�L�.�Z<%;"D]ڋ��p>M�`��	���Q	��������,� ��H�`E��~t5�\A����z&�<d� ���P� K�o��MW��ܴ��h/	�D� P�C�X��*�S�j�	[�
� F��U��x� HJ��ߘ��k���%��Q�A 0ot?��\ˠ��E�����C�T�ܘj�������������~ ]���:����;��3��:9 ���=X$F�b��{� �R����>���Tw�� L0��~=5�B�����$����d��8 ?xU$l	�3� rA�߷ͬ���`L SO���[�D8�P�t ��8�V�ЭPG�:֑(
��+VoD�0=?O�Ja$�e ^a]���; LYU����� E� �h�-^���_�@�����" ��(��i��B꨺��?��`q��@�Z���o�V�����l�$D�b��=ƴ���,#���@���� \���F����`��͓?>:��gRt�H�p��lH�,����!��>��& #�[�\ b�7���v>L��@8��EϬ�D��'I���~��� ج��Y=W|d� ]M�U����<���9Ƣ ��G���-m�DO�%b�Ŏ� f�a4��� �ND�H ���dz���Gx�4S���������Ux�:3揃WE��*R�$�\L�n�� ��ӏ'���Ax��E�# CHhepU߬=��F\�΀ D4GE�:x&���N� 0��\�D�W_����JEH��!��aVk�[��uF &y�l�e���E=@��orڬ�9���;���D\Վ<���If�J�T�� F��4��h\@H� wvl�D��{���X���p4)A��h�z (��D���З� �WK�=%L� �f�;�7\2^��D����cO|� ��?0$�8�t��% S:��i�"t ��)En��/�����e�b"�u?N��gXP.E/2��z�_�� �$4ᱏ0��m��^��*<J�t.E� [�L`f�	("@��D8�IE�/H�4��A�_P�<\�e�� ��=ȟD�=GI�� {Ls7� �ʅ��<���o�������GLPX� �$K{��� ��x��}a�E�P�/��f@���A����S�
�E��?X0���i� �Y'���1�p�.�x�^E��8 ����U% =��R�l��	�O� ��5��DT.��!�E���x�&/��|�� ���&���@��@h��%�x��DF�aE^��?���$� ��p��V�h�Dm�H�(cp� .P���ԤՆ��<2f� j���D�t�.0L�'�@���E�e*q"ĝp@�&H� {Ŕ%�����`��Jt�\΀a����~ D�.�J6��`t�;HQ���VB�<����!  PV���	�y����n�� �%?;E�D t�ʏ���&��x\[�@�I� �,z1@/Ƭ��5�ux+ �Ej���ȹD,�n@���l ��x�9^IH*� w'��. ��0�@E��P���x_L�9�� +/��BF�K00*��DR>�ck�//փ�f���+�%D�������]g�~�&�d�x�1\@ U&6����~+��D~���Lf&�L#�@�xX���P=F{��=�ĕ�u�e��a�0�D�/X�!( �u,Y9�gw�����@�	� d�����'��|a�A�Q@J��1L��/;�.�����9EZ�a �,t��PS����׏� U��l��5����=oBW��'�d	l� ��8�D^�H}����c�.%�M b�|�T���XQ��z@���ac��$
搋�@ć*f������(�RE���]#W.*g���m��a��P�DvL;U/ ���@�<���i��F�T�;
,�S;��`>�s&!���1�����%� D3�Eo߭(�{�a�J����_�nG��Pt�ĩ,D�� pi�<"���0m�p^��= �UE֩�Dw��&�8�z ,9���X�����; �DM��\��FQ�� C��֏Gu�Ϩmp D�� ���8$?�� ��BEǤ���F�7�xg2P�C�\�0t� k�ݚॏ�
�|f���@H��?���x/�8��f%��h� D
z�[h t(�N��rF`d;8��D�Ci�f�)��Y_3 '�h�E�	I��pD�:K�����|�����4�DB����X��`���  �ܬ�Fp�`<�<ӀC.��HYX؍� ����Z�E;b��U\�>~_�+�(@�E��6
���> 񬳉o���� L`
�6��b}	t[`�#J�pنr=�eP��Ԡ��� /J�`�}q?s쥯��:�@(���� ��k �7���p �By�2��K���D�X�$���`���%�D\�9�`�I��� �y�� *'O�{�o�0���I�� ���`䜀�� 4�{�l�5�����\̀:Ո�(,�, ��H�Av\?�`�(pF� �����<�X�6ݘo�?�u�ԏR9��Z_��0H�a< j�:e������$;ܪ�Ⓦj9�1 F|Ѯہ	 ���OCea�� �p0��㔌 �#�&�u �!��qXV0�Nw`�~d׵Q����=:)@X�� �'5aՏI�l�N^��2!��0GtFMԊYo������>�G�_�p�2 ��akH��H�e�W��	T������:l���$�_'��3�i��`��+��?oC��U@��t2 I�ڝ��h�"D<����Y�lQ�0��В�;'X��Ga��� �B �ܨ������h	^���  d�J���L�Z�7F��jT��� �������X�L��������`k�~K���J��0B؇a� ������
���ʎ���S���k����=�L�/���?
��0vH�
	Є������uH_K*�#�m��p�_Z0��R�#FIC����͘	=����%ծ�ӫ��)p�\��Ƃ�T� G��j- J���g x,��	���x.��&dg\ː� �L&?vP �~q��(�a����� �,Euc��'���l�����Z 5E��p� �����K�/E�[����=��9����f��ٌ�Ga����� %��@�t;�H`\E���`rJ/���8���3����:�:�U���W�$��� Z��H,8I� ֝���P�دe?Cp���u�a�<�:>����Y1Mt�'k���@�� G�VxwD����Ŝ	�@i�p$ 'ߘR*�(8E�4�7����߀v�Z�r`l/N
�Kň��t2@�#���\��@����NT��� U�+�ZD���&��L�ͳ|v��РP���0 �6`W�5��i� �U�E�&��J� ؖ�rs ���U���F�;���S�.�@\� ���7�& 8��3���[z2��������cą�v�ά��8_l��[����q��D��T��B5�~K����� 
m�x�����ԡ�>/ ���IB ���uO�/�&J��g���� ��a�D�2�� IHO;���w��	� �t��5�ܑ8$0  ײ�z1p�� J�e(�۪���i��s��_� '�v����<
M<3��À�᪹B ����sRX ������T��ժ�w�:`� ��H�W������u�����@��4�e 9x�p�ެ�!d���v�s�V���G �&Ø%� v�ʬ�fw���81'���{=�H9B��݌�����t��\������ӈO��G>�l��mL3��g����s�c�е� YXL\,)y ���N�l ��KX�|�9�3��/ ���� �����J����o�4��IU����%�s���뙢 �#�<���t,�&������-��<~�@7��[rS�F p����>��Q7� 9�X�b�H�8@��[�Q1��%��O����� ��^�"b��� A�!@��2p�Hb�Y S����W�
8�lr�#4=��������sm�����=���8,�Y/  O����G9Q��pA<r� ����5��:iG=�w�NȆgC-�(���P�nTs�	+��c ta���=��
N ɖÄD��"�s
��o۫���� �[���� t�֬�),\s�x���EvBA��h�&��o-u6��`Sݬ iѿ��=��2��fh�˘h ��^؇��`]0I�����薓�Z�H\r���z4v`�0	U(�R ����n@*ؒ��<�����0H�H.�x{ W����� ͐�J�eL<=�W�h����0l $��P��]��X�A;�s�ɠ�h���ig�(��X&9P�(P ����(��sǠ��ǥp����b���N�S��7�g��rj0;���tVCS�.��ϰQ�� �#����2 }��*|��Q�`����p�X����(*wC� ۨ�^� ����ku�� D�>�J� /�q�o ���SG�Ei��A���֏����L+T�<���m���;�P�|�$LT�"I���/��=&�P)w�L�`
��T9���yx��$py��巶�)8�9��`zt�c� �4$~&� ������ L�6s^��> ]�ͩi�	`��c�a'�`�pҘ �"X��}69U�Cʬ�=���v0s��� 	V�;IO�z p4�-{�� ����sV ��9��SM �\hf%�� $�K9�L����s�y^���F %�Eg�eq����;�s`v�<P� �Zrq4�l-;̓2��گg��s,p� [�\�L�g\�&!��½�@\��� &�sO�Kȉ�EP��?�w���� tم�s�@7�U a�B�Fg��3����s� �N��qr������8��1IiE �v)L�W �
VU;s��|O	�D<� 8���'�p���X���� ��r��Cѣ���E�=/�Y��s�r� �m|W􄬵 #�3�j&y�%��<����� ZD� �`r��NW@)�1s@:Z� �����N SV#��W"(�z/��@Xm����v|d>.[Δ�\U�^ =�%rn;s�bq����wG:n?�8I�� W/�t=0��� >�m�\W�0�& �蓀o�k�s�4�ᨈ�X  �)\N tI	�W<��1�sR�|@��������5�Y� Kі�Wv= s�L�h�bN� ���Z�P���aA�р�~�z�/���Wt��#�0����(_s����@u�	3^���	�Ec�n��p�����q00�_6@L0�$�tEPs,\�>��]�����A�q/�W�ZL+h >������X Άӽ�<�j	�O'�L �([�WLu:�lAs�\@p��-�g:K� ".���3y�� �Bh�sLM�p�\� �S���g �s=%:V)H?� �f��͜��p�I��8�Y( L�����X hO�yP�"	���l�Q���r
� �RJ�� ~��?Ζv� G|⚰7<�p �Qs�&�L@\�[T e��#�I��{ĐP �Glr*�4F���M� �����s	tw�����#�S�5��p�Yfڰ����T�
�
��n�i^p�t�d)<%��x�w�(G� ��6q�v������w�z����>;j�� Zr�9�������p�sPC�L�S�^�!� }����:��s�@@J�dv4e\>"π�{�U ����Lgd�s��XW��@�D�dhhj\�` E|,	�&r��GtTȃ�i��`D[t���f���n� ��4��A� ����'9���8#rx�>�
	�"��p�}����༥�'���s�~@	�X�P�����a�`Sx�v��!8ހ�����L�-r���`��� 	L|wV��Sx���-�� DiNa f�C{e �_]��|-�����/1ª���G�H��W��2�d. 3JsMUQ5-q�c���"}Ɯ���Bk s�| =���~(q ���� �#	����~Mp�\K�}���Fhq.r8`�����s��|>�\�pH�H8  Z	#�oL������1�v�>
���&ep q:��=č`7�mt�d�}���"�a��X�Z�	+L"���/c��V�>I��j	]�����p�(Ә0��Ψ����#�> ��@��Z]����Ï���UV��s��C�oG��H@�� �`Va�{��3s�-�/@�1�I��i� ��g
sF��#��8L�Z<5�2�`t�i0t%%���2X� |��]{R�
H�I� �=uʩ����v|p���$S�F ;x�J�X���L�|�6��D���d 8�9�.>0���>���������Aj#.F!�-8 �y ��$7${j�`�u�(���F���8� $բN�v�� ����6�p ȟ�P$h�n bw�R �q�W�� �@�~ �nC%;H^'��}EƲ0��� 1K�M��^ �p�C�� `�u�D�n 0�	+Q�� �ɻ��LvZ�"�� �={�� ˗���)O$f������dȫh�%��Iv�g��qa�� ���X�����H�hG0�tN��x��#z�a"���Ɍ ���Ϸ�); ��(2��$��Ǻ�bЮ�� ���ȯ� ���'��[�`��0ӌ��pZ����UX���ټ
;�B� �c��4$D�9g��m���)Fp�$$�(�b��� :7��ۯ_ +mٖ�1�t�8X�-w#]脁0*�,�� (�$W�@x�s"'Q��ʄ�����Ν��#7�՗ZK6 9�[v�V�_#lo��p�! ۟\�p=�x��cV�EY�`�ŃI�$�a`4!{�5�U� C��&Q1�!���:g�����{H� ܁�K�I� ��!ل|�q���2�;��������� ��\�f�d�<�s��Q$|l}eZ�-�!�a��@�R��`hT +�&;��gH8��K��2�k�P�]O\�P��N����6��c�A����)�>����`n'!�9��}6 �wK%Ϙ"�c$)������ �Vv��Ѽ.�D�5���P�L#V{|y*K� ����}lj 4��?h���Q�.0�[�yw�)"U����{��2�b� A�]���ݚ ����YQd9�H)���@�W� �xga��ɸ�$��T��[�P��%?P����ӝ���w(�| 3Q�� !ʙI�(@iO�髳<�p��Px�O�4�%�H 80���)�Cc1h`. ɿ�����
��A
�����|8����7تި�1�$��̤���y 0\�uܝ1W�(h���c:� ��n<�\�6 B�#
y�X'*� з����tIxH���) %���+� �ЦwW � ���^7�v�� �FI�Ã17q�(�u����l�@�+I����N�G�0 � ��䡪3�)��'���� Qv��ȣa��!H�3Йu(F�"� ș
��U'*V:�
7�"ߠ ���\�nH����b	С����"t5 V��jf�3H�l��u�ǃCy�}�F��F���H(� əckK�%|���*υ�+�,�����2� �$�Zy2��@��#�� �0`+9�}
��Ę	�!j}� �u募�+y�R��;q@: ��������^z/�t ����9�R_� �˔��%OP���R� (F>���` �,�0��l��\J�?�ـ��h'��orƁH4X � � Oh*j>��� ���K�N���$�`8 +P���p��7s9�u�M� ���������1+�����`�ё'�s��S�D�2��(�mt�8˘@��v(���@ϙe� y�	���M(����NE���H(f^Pȱ��%�A@!��p0l6A�N@����O]��!'(2��	/���xY� 'ʗ����eT"���% ��0�$I�R�H349g�a�(؛�`�6@��E+~�A[? r���ʿ �`��K$�J��34ߐ�����,�g�`}����"&�{�-x�[��o �h�5�E�*>K<�`��@�����&�&��lān �(�����2ԧ�Y�RW9hx ���0��1	�� �?F,t3. ��0b�I
�� �Z&8�� FL7���DX�n;�����8�0 o�Y�h:>t�&�� q,�9�#�G������s� ,a��| �-�l�
U� �����Cm8��.Z���' �D#�j�e 4�,�Wӂ8#�`,2��� O�?���-����� ���tJ~Q*�^�U?�H�b�+ 0,�s� ��5tN8 ��mXk�9 �����,���@�=}e8k�R ;.qY tB���U,�L �X �f�P�x:���-CO��� �W,��� 9^<
�X��8lvx�[�0����,���S:�Ě T����>ȵ��� ,��  (��.�b18�\���i����M�o, 6�&ҟ��8ph�`I���?>�p(��:~� ���*�89�4�Ϧ���+=dR��,�Y9.?��@Ƙ $�P׽�/�<GV�6P �p�r8��n�[X$���� �-�/�ж�x��q,=dh�8�:�"6l�3�iv��� -��m��q?��&^2� ��Q	�� `Xtی\,p���nl��z+��蛀l,ӐŠ~������-����o�[áU��� m/�~S,H Qn՝?Z��^e��9,�D@=�T �4;S��\HaP �8�|�-k�]���p��� >��p�� 08�O�|�-��m	� ��8�� ��A��kX�|�S� �Ď�zt,�(�J@��$��8�� ,\Xۅ<#�%)��q� +&�T8;:�WP���������,^�����}�-P29�� KCH���Hj���:mnDay��X��@\�CG,l[�.A���	���:�`�~28:OS| -ёD��B���};ݓ���X*�p(	�3�`��-�qK��:R�}��A����J=pЁ����&0�� �~Z�=ye �hd�8�� 0"۰U�-�.f�� 3ȗ78yun�Y�%�Ў&���IX�D^,� �҈�M:JrH��( �F�Ł\C>�L 8e�~
nq]X@,��}������`ER>�8���!uUp�(y������D���,�>g� �xm��?�$���Q���,�Y?(�8�o�[�9�
A<ψ ��C�:�8 P���Π(]�l�U$`u@��S<��`�� ���j�Jwc8} i?_#� �-�l�,����@Hq(���2��7��,� ��^]}��� ��TCގ����P�<� w�+���'8ˬ`���i��[�:6��,RmӇD��B��3����[���AVy��1E��>��֘-�8[���2P>�3�D��+���J� �[��X��� {�^7�� N,�-� .,�ɘC��Yb�f<��Ԛ �
�zG�� _,O�}٢ X���Q?�8 �������h.��,�Q���.wB5�@ (o��x г���{S}`X^�a�83��	���AP�;ip( �a_8!r~�$X�l$�ջ��v��4��,u���ʜ�?��  � �g>]��� �=�,��`-n��E���B2 B����dk���� ڞh<0s�|���Ĳ�:`/��QM�Rb74~6�`�
��	�%ɐٻ? 20XK�`�Hѓ<� �3и����@�G����x'���
@�����`S�"�� �*]��X�F��� ���-+�ò.f�`��c�:1n�8�_ `
X��T���ڸX&��hd8	��[��&ޗ�`�XغD ��!��=� �~X2�85S ���=�&�0� @^8A�o�[U��r�x>��!<*��"L�4;��v�9�o ���Y>
p��0Ҡ�-�,�M X��8�rt =�b�h���� �d%Wse�}X 8����;��D �[,��,w�pP	�����.<;W�`X�!�"9�`�D_)B�p�5ga0����=��p���GA�9yQ�-����{PS"�� �����]p�|��� �D���� ������� ���9R�ݪ 
];��B� ��"��� ��C��ͳ��}´�2�l�Z,�m�} �E��*��n�+��� ؏��'�≀�L ����^'�UM�$��G|L�<8-��r�ƃq�L z��Q@�)��I�C�]���L�`�-ٗ�wr� �}K=/)��n���ܿh�0!���L"0;Q�����S��l���85���c%1��-dz��A� b��X�P�M�� ���l�n N��X�rx #K�>���,�v0NM:٘Z ~��b�T�pH�a B��/�Dt�'�e�5G�f	�! E�)]�A}��XA��`<� ��m�5n��������`{���N��PH�JfaG\��d��`n�
#?h X�:�e�:#����NGV�`ָ�|�q��*�F.�
8D�]��aC����p)��'W�( � �gC�O��9�~V���|3( o��.*��A �5�Ӛ���H�<s �� r(�� ��!@��6u߲M0̸)�tF�n��I� ��VŇ�i�R�� ��]�t�n�8( @�R 6f�X��`�A�~>����$-my�8�*��W-�A����yt�'> ީ>���  l���ŏgG儶L���%no!> 3zM ��Δ��r�:˖�B ?��.�e�W$�Wx@�u� ������� ��Mj�� �a@k5�S�����!�D���&� ��Q�����^IE@��ހ" kw�!˹^�|� Rɉ6`|�s>.�7;�s^����:��u CF>]#�'<�yJ�q�� n��ޚ��O�~���=�H/{ KV$�7;ە �l���q��D�W>��1�)m JFTd�#c�X�t��*��?~8�q�E ��,$�����;�!��� ~���t�,>+Ā [��1ޮuOf˧����x$ �(n�>%�}"�B����1˥ m >��;u��	kR%{�[������8 �A�F�-PԪ> ?�8����|�U`� �9�C6>'1:�� t�yF N����a���������:3�7�%��>��uܘk�� $I՝.˚�<�� ��\>a���?C�.��A�f��)r�Qd�h��+� _��' �a̭U�� �`)�h*
 ���L1�>T ���p̹N�	g�ʊܥ��<>�6��$����� 8Ǆ���Q:{:�vԖ9���/$w�>A:��Zr�(΀�˙� 
�_$�%K�`��]P}9;D���&�����y�Vr�w X)$�l>� ��=�'�������<,� ���)(w-8>2�Q��� �ktb ��2ʁ{��>AZ �̫]'l �^Ù\N�� �Q
ԅ>c�
U�$s� R��V{
���D��� ��M>"��0⽐� �]�k.g�4 �X˯W_��
�t�C���p���3�В���5 ��Q��v=a>�&��#e�qH�P;�t �����i��� �>BJ�Z���.����U�n$� '���>9@ pȥ�o%�&��( uQ��ʎB������`H:��1���}��?�P>�3v��I0�:l� �Y�0�PP�&�'�HC�Ėz�[$U���s����Y@��4��h�C��.0������`0ݎx��y�R���1�,��p�G����̣�� ��t�(����%9�� &@�G ��=8�����4�<D! /*W�@,�r� �G�.B�&��J��X����z�@B:�| �<�I"�!% �G	|� ��㟕���% @�P�D� _�!�QG-LF^5ȯ�Ep� "K@l�����d@v�	DG� >�݀�%�)��y 8Xk�H̰��6�GS ���x@���'D� E��c: ?���%6�G� O_�CX:pƌ�V@/j�P���G>��:��w������ϗ��U��2Q�*�X�����%9:~�ɢY�@n�K;l`��Gj::�m�4�%f�"/�� U�@��'��crG#-�B�(�|9^L%����tR:4v�`�Q����dcMG��SI&=��0�t�?��zGFdp	��"�NV*� -Ϛ;�f������M��G|Š�ds .R�J��|4�`�@���ZD�v�� G�SL.�$)�n� P�"��j@gP��F��0��(�A��C�>�_���]�9��	{Bn=����zz��c?0��Ј;���w�� P�L�m�t� =��Z�s� \��
al�� jb�����;i��M�S�=\- ���1Y� �VZ����@�c�g>�w�dꀗC�y pY]����2�<A�Sn-��J�� �v{@�%��H�G�g�u�IC3�Y5 !o{����	���q ݚ�<V��z�6�D8hF�n{l�Q1+ ��\z�R« 5���m$�=o��2TxH%t��; h �b�[����!k ��6̷��~�wF��=�`�g���a'�E��ޚ� �o�^���0d��`n�l#�k�v�Wj����!H��8y@Ȭ �Y{pc��� �>��4�ż ��H�B`�YG��<P��v� ,;8�`3��Հn� �e�?�Ӏ����ѽ �V=�6Bpt �faL>����j���f���!C����[
�a�� ��w��S���(5@tbJ<r�q�7C�
f@�����js�����R,�!c� �j%2� O� ;,dR��-m����a"p0�b�U�|EC��ԀHjR
��Pߜ����� ��}�Оue FB9"��8 �����
�� Q�%K(� ��P!jC��
Y��g�*(S �or�곅 0��Y����*(0�k933pf'����-5`�<k^W=�1�m ϰVJ�`�D���Š��z0XQVO5
cw+$�܍Co����/�`]u;i�8@OI 3�$��X?�@�*kc��_D&�	�!k��X�n��s������auZ��+� ��D%����;A��c)� ��o���V� �L��u��I,�� hU�Q6�$�Y/{����b�qd �@N��2E1�Zc�!�P�4�d�O�	-�![X�ƽ, �����O��l�Qx� �$���cF�JG�DvB n�t���Z�BX<� )�F�W~������ߐ��D�<�1��܅G�WB�8��ɸw2 �DLH�d���p���6?x�8aP��';�$�aHR�c��o�	!hW ��m�e��y� ) _�I�]���{N�.�%��<e@p�Ă<�~AN6�"H4J���o� %�t�� +=��D�� N��s�5X�$c4�Kn�&��
*ډ���$��!m2�k��6(�#d+DO���H!\�]0��+�l�,�^Q�ci���8-a v\��������>�+2N�0h`8ڃ!���c@��1]b4=�L�a�FS".Q��|��$ ǜ��R�#_l�LWbt'P幟�ݼ;����!�y5��M->��d4?�� H�S�7�� |�q"�B*�'�%1��L,�ϫ!�Pa����t�D"]J�mxG��W��,���-0让8�j��A���P�@��`����[P���(�l�� �W§�J *� �r4#�Ff�<ER�+�Xs��| ����H,�H�@#t4�W�G�g< ړ�:�{����D%?`���J���2��;��<`O�l#�[/T�h�X���#�Ñ�j�6�M��\	a>� 
[�ޖ�" ��ۢ���XhD6��.et+�>� �2�]���dY����R�T�3�{��bI�v@���}�2������ tW���~5F\"/�_�o�,�1D�UZ`7=�)����� �������M�`��=��2'��~UL'���Q]1E��ȶ� ?� y�Dz|�<./�8^Fs S�)U�P�d��8y�H����N�d��л�C9 ��6��D�,�� 1�[
�=�+�ߥ�5��b?<4	�{�8�,.O�7��f.�'��?0C \��I�+
_q.��^�a�Io� i� W�,=��Ł<d mO�1���.�n��F��pU�,b�g8���j�k�`�ֲI$�8����ZhbO�������H(P�x� �`~z�#�I�K6�$J�3��<�A�=.����i�9�`$��;�D-Lc�#>I�b���$ eV��8���P��	��	�O0,��'@��QVĐ`���`�Y1!� �^z���Q;�Ԅ �ѡ��x�uL�@�4mS5,6nlB?z���y�r. �b�e�I�Qz���|��0�!�]3 ;�0-=�����<OoE�MGݗ��p�Z�PR�a����`�_��g�\�/ đ��& vj0����� �׿��� 6>�?�!���l��d$q<x@>���9Ȩ�� �o�-��F ��z����T��N�b��������aA�%�3O��A�z��0d��1����h�˂���^tw�8�e��u��d`=������vY�92 �'��8� 7u� C6�EmN�@�C�M�%��ڀ��o��#5���@R��]�IU���i�u�?X�N $� &}鏒��z�1 �b;N<D��\�ĥS �$�	���� �Ԟ ��֛ޘ5aE<�����R�PR�	�IW���� �m���p��� R�� ����TAh���D�VLH,��QM�u� '�����������e�,�7����k�"�}|K���'�a�~`}p� o��`1�n�X6� dT���|�U��{�e&Q ݍ,�y)z��8KGԯ3��k�WwcIPrXm� �/�ጁ��;���J<{@�~��D� qZL�9�	�,�⼽�\W�{���7�ڧ��@d�� ��n�g9~�O+�$��5I�������y�^' t�U�L�<�.�P�]cH�"� ys��E�/F&h?> Y�Ɨ���J46od��S�:� ��{���m��D�خ���k��? )L�W�=�d5��:��A��D8 ��߿@�� �+�Cfd�9� A��s�L��>�R+f�?�a�x͙#�İ\!�' LCGN~�Ч0L4,Ҩ���	�逘�i�zT���b�`�NM �e�>�B�` <j����9=�+�D�	��A��ӧ ��z��;o��|������@Zrt+�;8��PP���N����c��;�ʀ�8X����7��@W��	Kd@�H�1�8�w��}<.>3�'�m �yҌQ�H ��u�4\�d��_�����T����>��� h���wP+e�� `􂔅f� 8�7�U�?�� �	�JAkQ.I4`̂<M D0CV���[ 9whP�2�l o�(��!���)�.���
G%Y�l��U���\6��X%@8�7u�"<~� ���U��a u3٩�%��՚��D6��|L/+��$��V� 	��������}��mJ9� T��0,eS ��hp��'jl��b&�����e�+� ��8�s��z��MrW��� .-:�#�=�_u�`�(���� ]MP�1� ���!h���T��� ļ���_�azꄍ�Ԋ�q& �$"�<�A��ʛ���p)0�$^� ޅ�m�u��RGL� ?�,Lm��$�J���Rr���8�8�p��>�L/���4� B�����ao;ໟ�zﭩJ�DL���HVM@�����vcY��ǹ0KB�`� 0�E�f�������+F`9�᣻ yuA��� �X��g���`p� �Y��1��U+��?���
 :��x�LG����jd��  Й�w-��=ـi�%B�C��I�����gAz(8�� U�2N i Ġ�
���V$�z0�����IJ	�-�#��\=����$�3�l� k�F�� ��c�	�D&� �ކ��8�����,zb�<��t\Sa��{J�X7 �Xޣ�?�� ;����%�P-��o:�j� A*5�ɖ)0vn�� ��M�{�ٸ�?t9��b���+:��XpH���D,� ��f��h���$\� 1���T���O<�X�i6�2��z�I��~�L7Az .��5�F(E�Ӑ  �CM2{��<D�@�P�h� �7g[y��<�ǒO��@0T�ʱ\�Xe�Z?��L����u'%(����]9;�8�D�/{�Y���,����|�2��cҘ8�I���0�Ԥ�	�������������WE��IN��ִz� ���E�\���%J���&St܂�NU1`8�W��8]0ɚ�� S�����2��� ��I]��;4��с �8a�@l��Q�E�hHC0��LS6�������U��!�����łD�\� x1�~'�d�	�� 큞]=��M���e��{[L@"δ��9Ll��x2�Ԃ���8��I�JB�����\��A��l �;+`EZ�! ��Rb�-Dz ��o�qW��� ѷxQ��G��>���Xk���s �=d��{����4a�1X; 8� E�͙�!Ǖ	��Kts̈�%�����a\[����?�#>�k,�DPc!Ԓ���W �BsC��<	��c�����AM����.UȨO X�����L�@��<|$��01`��h��Nq@���X~��'�^�m&t<	����lqUzN�@���;6��,��{�_��&b�����)e)��>�&�Mp�	X����! ��΀e�X ��7������:��@�"�h����h����/e1��͛��44QH��ދ��~: Di�<�l��mǅuB�9H7���p$ R���m��W�%H�p� @�`���>��@��J{���%�2s�?<�V5bM�����1z���B� /P_� yV|�$bDӘ Mf���P�&�: �3����R���l�n����ǜ<}@�f �B= ��Z��. �:��Ez�� L����>_�B�$��� �Q�ݾ7�6��z�Kr (X��� /ǂ�n�vB�
�=��G/38�X�{� Ԉ�]�L�c��L�T���{"�%�3��'_�L$8�� �\�b�1�$������a�v��cY�@L���� Ӈ`���d�t��7_�T�Q��ʘxX�4Ӻ��^>'8`Q�� H����c�B��ܭ5=��t/i�,/��@�� L�I򙳪�:zU '������?�%0�/��f�=�`��[4 t�!S ��&�V), k|����>C�",�t�i�q��欖�r�� {��~�� ���?�X[,���G��-����}��2��̟�� U���=���(JA�����t1��"��T R��a�0!�\d��1첻Z#?<���QKaW+����&UiD`�������O�H�7F��Dm+��@=Y�й����;0�r�L@L� �o�yvz�W H�SM�0�P�Qy��*v�A�@��L�-]8L�u�����H(���#�C�^I����3� �o�	;E���� ��XDo����d�<� �x~�/ͻŇ,Vت �ݕ<�׼S$�M�	�߀�;�Ɛ���h�ZU b�D�@_�JKl ��� ��Qً�E8�L2!<���
=����&02�� ��+�H%`�b\W���?0E�H��Dr<��� V�RmU���r,�4C�d�����PD�� Ք(���q;�+F�/-ԝ1:26\���7���Jd��t���S��=dH�~ 5]
�̻M��x�O��az�o9Eǉ%� ���+D��x l�`NJ��Č Pr�e�Lz��pf��?D~� o3
����u ��}UaR���Oz��*`{�����݂4U�$�o0ߛ�}<6�9�%I���r<�>ϗ ןP���bm͖��?9� ����pյ�:�Z�  �;�0aD�TG���ĭzi@�ARCDB�P �F ��S1��� ��RL+�	Px�N�8!��&��@�� ����W�K?��8��R�D�w:��� �����'�%AW�D�� i1-ϧ�"�5��`^�!�L�]�`�̯@;\�Z�e�mz�} ����'��l�`BfX��<�����X'��]���ڵ�+��m�/�Ȑ� �ޑ���8� �Sٍ�"�6H�(�Hc� ]mR_vZ yDޫ?���@tݚ߼��3�1��D�U%DO�p �����@d����<� ��"�M�)� ���= ��vD�L��p��#6�^�Pͦ [d)F<ܴD�y҅�ڐI��rA�",H� `�o��-X`p�֜a��s���ly4�� �G�Q�#'t��>�h�n�}v�H�.��� �b`��z�ѯ����OVc��X9��� Q3EO��5��@���"��t6`����go�J�:1d&����<�) 7]�9N�\���������؝2{%�����p��8�z��L���8��� ���oY��t(;WN1��uȺ�&V��J��b� }d��	[B ;��+|�Q6;�RΈh �A��/xn�='F� �m��3���"��OI�(4?��>�2a��6�"8	�Ȋ�� ���b�>��ٛ''1w��L<�ے���U�Lp�����ax�Z�N?J�� �CB� &w�=/ ��4��9ï ̲STU+�\��ն��ԁ̴; ��ɤ�Dؑ]��V�H\ٷ i�S:.�f q��X�3a �+6�7{���D�0�+#CE�4�x�5ǁ�S0@10�Q��>6�����h�U`�2cXP�"-'6n��B�8����9 � M��<E"�`� ���Wv6f�(ژ	�V?ڐ�i��p%�S� ���s6�>e��|`�]! P�l���݁�hªv챈�>�)�u�W����,;|��R�pHN 9��i�� "'�e�� /T����Z2 9���8�+��1�0h� L�b���%��/��f x<� @�dCU��t �VA�:O1��!kU��lP/(<üR��n��K�����@ɍ-�Jc�W;a�N���$ �͆b2og	�&v��$$Ì��8����N ��b�6-zRD� ���'�B-�L��	 ���,����>�6��,������0\R����3 ��Z;�� ��oܝ4c��O��DX<��ַ gݭ>���b} ʪ<{&V9=����JX �`���|��P�7;3p�����0o�/6�� ���;��7�f��J4�Ȅ�����'2ۥ W,�#z��$T���-�7,����Y�+�x�oO�O�z��ą���xb��*A\�GY�oOC�Z��������9�.���%��� �uT�����6�Q� ��{�e�9��m� GSֳ���:n� Ƒu1�ߧ.��8xR���tgw� y ��ց��_ @�H�����<�y@V�� G�Ҧ?�1�8:	 ��d�)�[N����P-�B'���!1�LS�����tB"!X���|+X�ǔ�@��، ����Ʌ��)4��pg ͎����{��6�,@3�V\W<��dX =�|�a��ִ�c�;� ��.���,M�pߒ�k��̤a�W�^į� +��	�f��<^� ~�t���C/����� ��k����az`D�<� v�N �ԏYT�Z,ߨ��� �H��x��(;BP ��ZD� ޜ�z��J�ٝ�6���b Շ��t�Q| i��6m){'��8��`�"����&��g x�m�$Nt`_�� R�`��Bn p�����ou( �~�a��H<���$��Y�o��1g�;��)��%���(>]�`0�?� W�T���V�L���r�� a�Ymx��l��Q<�cyGs|���jP���\�9 �����G	 �m'/�� a_<����O�h�aV�$+���. �G�p�� 냛� 0q�.�z�9�]`I����x;D��9�� ��gЕu�rjl��_\����cA�y�x�.�n0�]��yc��g� %��<�̰0i{����gR�� O��v�f��b`1c�/р�'y��F�0���Ġ�|��Q���63Lճ@��2 M��k��AB b�V�����QE*�1�!˴p����i�j�i��P����� ��)�1�� �W�-a�H����Ϥ� �����Q=��j�#��"� �{z�H���ƹ��4�Do��8�k�z���`�iN�F���� M%�U���N�?�Xa�x��Ţ �B�3�i�xM��0 ��u.�op�j&"��� �aG}��>��8�@<���Ui�� :ʒ�d��`P�a��Lm�(`KX(���%���4���$�z���F��yjL��� �GN@V �27Hhqp����o��= ���!� ��:z���T߰7�!��e���qY�5v �"C'4F&
��8��@�Z���Lw������Y���0�BR�� ���g��M�4�k&��Ga	�H�B�$PU���&<����0\dX ��	c�9Fؚ�8��=9�� �� ��|�3�X�,�z���1�� [/�|qwH�8 �����`X��:��/ Ff��<8 ��;��#�Osd� ϻ����A�Ԙ(�hD> �m�?[�`�9diF��<���c0|9I帀�j.A��4L�A��V����/`v�� G���Ǿ�� ����_U����@��T�]`�I�ǄH �R�q�Gj�ѷg6ڪ�.B�fվK0����Hr1�'Bت����"�V�qD2�w������!���Q�Ht�Y�x��u ��Ǡۍ�Y ?E�!�)B?s�������cN���5jԬ����� k�_��U�, &y��T��](H[M�sc���0������ +VǍ� s��
q)rOGn�* ��:-1VK��
8 �)��X��"�?��  �Ud�_�$��_H$7�� �5(`��q ���3���.�Kx>dN�|��͍�%���5n"��i�u,Ð��\�2a��VD� !;����I\`��OE J��}�7- ˉr�H�a��&��`���@ �e�C��Z<FN�7PP0LlK�$,�oLc��� �%1�B��(�ȳ�o"�B8d�����G`viҭ^	(��3�dj��p�B�l����8�ė��1.Ϛ�@*m� c���vU�Z%�|ͯb�jy�p�IhGo�� U��Ѷ��:��l��D�s/`�þ����&�;��p�oT���j�V �2���a�*���N��]�)	�Ew��l�>ı�8Bo%��f�i�|o'��`t$V�4��4 Jm+�MSN C�F�䀘�bæ&����Frd�-9+!�Z�!j]y�� E���U�X@����"fT�H�@�P�@>/`x����3��0�  ��ד��[�@�찪� &)Ց��u9����a�R��0����ްD�	K\��෯{�12&ߏ�� ������� �b�� ��<;>^�M\ҏ �j����y�P3�cDS�`�i+��,�i�"٦�@�&�6N } ]�&*(�8d������1.�b ��2���Ρ #�q������ؿ��1# 頯L�(P5���^	� dgF�V��5	�J�� ���;��tR��А�1L�6`ҁ�	M@�
�H�Z ���������@�1�Yݗ ��78��,��> @������`���[��:�8��4zN �B�){ Γ���^�a�
t�X�#���a�$w�5�@7
�">��j��c��d��2��ʆڳY0�I�� ������8s�k�@$w)�.�1�Q~�����}��71�!y�?�u3}B\����"M��>���%+?0 � 6g^a�/0`�Y$A�� z�ޮͷ'�	k�\�@�1Ӏ16�r��W���N(u &@�#3��b�F�H���EA�o d9�Q�_ �5���#����ma��0
{���Xxޞ��S �����ܯP�| �G��}ݝF+'��� )	#wR�b!H��*�O�VD��X�"$�m�F� ��� �@�)p���[������0��a����P?�+ ���҈GP "���(����0�A� �|׬��-� N*ƚ)!a�Ov1�1C z�
"��5_� H�Gh���� �^~C�V�a(�r� ���*��T[�P�� 
�@�r�H�H��~���� �����\F�I��L�D� :��L�k4~����Dӑc� �R��+y ��Y�E���1`Jj�ϴLx������	�<� (�w��3��!+�����4�nX�$6e��8�.2 ��9�	�؞0�He��� +A�>���
`�0�(�&�x<�ԦA��������] hB��@M�)}A�����ڸ�P�� R����5�3خQ��8[��"��\�|�|��9�	ŋ�/�BD���r�L�-[(h�	��@(\oYi�* �҇��F�$�� '��
Hzӆ�DA �G�p��)�[ T*��k�U�
q�թ���IN�0[VI�?4 9)���3+!`��ѐ�x����t�b��RY<Q� �����T2�鹜�m�nB��PX�\���%��Ҙ&>�A�b��5� I�P@8�?Ø��Q^��:s��`��9;�Y�@|�D�f 2�$}�I�K �h��ZFR�^`C@x�x�,��Gx 
����n� ˽>�p�_\��0�s��)�,cY����	CSIpB��h>� ~F9���@���X ��`4��G��T�f&`0��ң>{`�H�Ƭ/^)���2�0`�A#fC��w�4��Ig ���w���� p�����1D�����~��Bϻ�I�L /ғcW�>^C<��ޜf�@����(9�3T`�r����"�Qh �UlR� B��f�>�(��J�� <��'���_�?��@� ��,^�n�W �Q��fV� ���{F��� +�w�V� 1I,H��~���<�{�̓���$�mU���K�a�&(�� ���8l� 9��t���0<��p"@&q9��� B��&s�DP�d.;y�:_ ���
\u���>�� ��l%1�qL=�e������]�$2�\i~r�� ���K���X׈���`p�~�8�	�%$���U!�0)����7B_�E�Jն	rF�\��ԑ�̓�8����,Q| M^��P��B���>���1L1��?��V� Tֈm�����`�.��(?��������:��$kD,�8 ���L�")b�%T�]"�����������| <�x��LP` ߱A�,��*@�	��-&X@�	�0�E5 ^��`��d��9��|R �\$�7��0�I+V���B�W� �������bbH�@0�tR>� ��v:���ta�C�9�� ��7�߬�� � 3��xҍ�0�옏��XF��H���'���� C��2� \����P���pXY��<�p����!�r���c�� ��~9�f
$��`l�$|=��Ŕ���H�.+30� ��pv(8X��� .�}����&W�D+� R����,�-3s �L��� 
}����r3 oeR?zJ�E-��`죪� �8^��ɥ ڔ�
έr��0)�1Vx�%������c o�� 1*O��s�E㒚��� �+�:�G?���) ����u1���q�#@ͤ�H��������FC�08-� ¶��L�
r��a*;!�\��0>i�6�< %�~:������ �y��f�&��h�rG� ��	l:V�	P>��������(v0��?ȉ2:�Y#��w��(���nǶ�b����"S�f`����2�8�9��3@DP�x�}��u�\���*	�B �]�z�2��\���@A�Њɞ��M:�D�lv'�|�`� ��9[� �|������$��শ�p��t�K1 lr/&za�n�+�] �� gRO����E��[�D�@�������U n��%�1t� 5枟�{,�2��ܔ@�ҏV f�[�$�`�� ��MɢN��{��ֺ��~����'Y�E�k)���� �ͽ���N1@l��G� f�䳻�=�9$�'��j��L+� ���QӍ��Q$ ��[����X@;H�)���hK Ș�\��L(&��a����k�5�90m0�A�Y��у�ށ�#����MȐ� ���`���� 2��a����HA���D�j�� Uw��e� '�ȀE(�`�q��c�8
�I��٫*L�ȀjP^H��'��B��@t�< ��E�|����g���y��9������*���:|l���u� �`$��-KF�l�ə$! 	�v�4W�ա�Y��Zy� B��A���20�	�aK q����b �W�){[C�Q0��g ������.�PY�(R|��f��P�@�_C���&�=	�f� _%L���Q� 5���1ۈ�r����#��@Jz-P�	�?���cT'
פv���{I���)\����
�����烀ǎ7�F��H�Vи1;Q)	3+�@��b9�r ���\���f��,,�{Ь� �YV���<� �9P�Ժ���@R���"� Hi��v�j1ζq@��`�� ����Bm���(T��
Ka���������~AN�y�eu s��=�B[�X|����d��o���Y$�@��w����Z<0� ��Q�Y��u���-rl�U$�� �j��hL�rL|/�G�V\@��T��r��� 6�����a�,��7A�0[��lR���^O%2��]\ԯ��� }��[N�˃ :��ic)<�&��@0F�q�L�\x�FQ��|1�T���<o� hfڍ���v b��Q(qI'�ܢ���y'����@�5�+ x�{А�,DW+�
�)�ޤ0� �2�ӂ������ �ؓ���� we����p:��,2τ ������t	�����%��z�Xa���ϧ��X����PٯмӘK	��(��.�4`���e mB	jn(�/��l�&b��)���@^+"Yg�>K���`$��˝\L�0���%� ��ǖm�?�Cr�.2+�`!��	6ſ
`Tx���(;�@�{;n
�z,��!	,l�J限�� 􋾑Y�[���ǰ@�*@�o�ܲ� I��<�j��xߜ�+.���ǻ!4���/C�� �|B�����`z�n����Z�kS�i��#`S� ,ǥZ��'�ɐ�� r���F.f1�@Owyh�d;ӆR�`7��N}'��֪�a Q��!j� ���k����?.F��@�DR ̀߆��b�$B0�{Tn�ο�����(�1D�� ,Rv?.�a �ܡT�\��%��@ 3*�Ws�w ��<��9��0� ��zL]�?�bk�Q���̧\���N��Z@ a��@j,Z����X�8�%0�1n�����튵c���RI1�$�Z�*�m�T I�ҮP ��l(��b�N������ؑ���JJ�8� �t,kdwS8mC'
����n�JȤp �vPŷ��N�JgV���ӌ`FG%z�ǲ��@��u1�v1.p��
�3y��;���g]��0�a :2�=BG��d _�a��݃�� �@��=&�H� R\3�ڐ�L�	�|%����-4Q	Ĵ�a�c�T����O�C��P�ŗ9�h֮�D�[\��"���~�$���_��D2�	�x ��Z���~R�K0��"�t$����1	��\<�2� O����^�"|����B��T�\Q@���-��v�>�/?���@� ���6gB�`�0)���㘣�����2 ^�y��� J=���rP� ��E���c��� A��i� \ҿ��U�ۄ��T#Hl����2C ��D�s� ��3 GxJ
%1���hI�F ��\�p���(�DE�� �Z�م,�R}�~�Hp	5xܠ İ*���L��P��� Ab���"����O�d 1�#�߇ �^A��N��Q �b-8�H���N�@�pj���-���G a�0���������/ �C�7�� 'eQ�noh�\;�08��b�G�R��fW}%����@0*Dܓ��4_.	\F�*>�� �8���r̐�ob咻��y� L?N��y �*��k��Q	�5����G��Xjk�d]\���� fAI�� ��Jh�� ՗C�]�wnR�� �v�zY����2�{����\��A�v�	~G�Xa�� 8�&VD ���N�0���'$�� ������ �sI[�{,��*'��  ���R��J~��ǭ����b�5~�su����tM��	+�8\�?�����OTπ��[�ޘh0�z衬�|�N�˴	��9� T-y^� 6i��2��A� ƿa�B��
�CtP����0�5�� W�e
����X�`�u����^@�z/� �Sw!@ɐK0��8�-ۘ8�*�Ђ���L7��Y�}��֕����3�&|�����4�ʸ �VB�*M��u =��]��.�`K�� �<9y���� ����劘�\����䒐 ��J��G"�J�(,�>ܵ�b"���+�=@.���v ��V���
��T��7��Lu��z�/�w(T�@�3�20�&�cDF�!��3 h�(z���1��I�R(�k��e:�����|w`�~'PD�z�R��~ج� �{�ݛ=2���q�l�.nX� ��B�]��+ �����	�H@�尧re��6�X���	5�Ĩ�O���� �@�*�ՑP����<L������A' ި̚L+� c�/����	��%�)$�E@nb�� *�Q.�v�����@̨� .&>�9�{~QJ)�tF���W�,x��,[=|`Ko��q �Ǩ*H/֛$�'��x��Vf�u]	(��P���� ���G����,C��7' *�-HB\�l�� 
���|���������T�iȨ.ˈ�^��u�d~�O��D�̴� �'��;?����\�ĵ� [�"Rw��@��~??v����GB���҆�Nxc�ԙh���tw����[��G!��\-?���`��x ��1��͹2�ߞ�u
P�R���AFMP#�
� �↠��YV�jӗ��=� xo
CڠD�|�}(�����[��^]�("��`Q�I�d��%�G|��+��:٪��
 ���0m� ܍��}1 ��hd������� �N3?��<<����%^�p�Ԅ��.ѐ�0�� �(V�� ^�Q'���	���Ś �(b O�:U�a �TC�6��	L3$:�8ۀJ�N��2}	,x��	�鋄�I�(�O����1 f����2 ���|i�~+#�D����0�� %�e�� �r�	�5��Ĩј����x� �Z�hK;� �dpBX���1����l�(�tc�b|��Eo#���� r)���������m?%P���&&,�����TH6. ��$�c �s��ʹ�	�����tI*�2�Щ��"ld���88�������،�p����+�Q�������y�� �|J,we�-YL�	������^ ���-�Z+?�}k�D[���_�d
�}'ƅh �u �����-x��:Ö��Eq��Q��2�ʯ�g*2 �8�� �c��>*i}` ��Z.]5��24{֥��FA~a(60��"�� ����g�r`� ��;�@N+" ���	��YX �ɂ�e )�A�Mk�� #1����������4��_,�.h`�C���r�̠�\����!^��W������&/���@%IsY	�V���݀�����@�:�]�6$���Zה܂0�`d;�H��X�'0����2c��{ٱ�Pv	~�1�t�� �,ki��� ��O��e�	L���hDb�	��(8,t`q��
_����@�U��-���� ;�L?��\�C�>��b���*" ^M{��9)�W�-p ����k	�x�~,���sG�(�+L�������3�!@�&9Lw��Mӽ� �]�����[�̗���                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                      (       @                                ��� ��������������������������<����?���������������������������������������������=������<?������?�������������������������������������������������������� �� �  �  �  � �� �� �� �� �� �� �� �� �� �� �� ?�����?������������������������������(       @         �                        �  �   �� �   � � ��  ��� ���   �  �   �� �   � � ��  ���                                                                                                          ��p          ����wp      ������wwp    ��������wp     ��������p      ��������        ��������        ��������        ��������        ��������        ��������        ��������        ��������        ������          ����  ��        ��  ��            ��            ��                                                                                                                                           �������������������������� �� �  �  �  � �� �� �� �� �� �� �� �� �� �� �� ?�����?������������������������������(                �                         �  �   �� �   � � ��  ��� ���   �  �   �� �   � � ��  ���                             �w   ���wp ����p  ����   ����   ���    � �    ��    �                                     ��  ��  ��  �  �  �  �  �  �  �  �  �  ��  ��  ��  ��           0  1u     �  2u   (  3u�4   V S _ V E R S I O N _ I N F O     ���                                       D     V a r F i l e I n f o     $    T r a n s l a t i o n     �T   S t r i n g F i l e I n f o   0   0 4 0 7 0 4 B 0   @   P r o d u c t N a m e     W i n d o w s   U p d a t e     4   F i l e V e r s i o n     2 . 0 3 . 0 0 0 2   8   P r o d u c t V e r s i o n   2 . 0 3 . 0 0 0 2   , 
  I n t e r n a l N a m e   s t u b     @   O r i g i n a l F i l e n a m e   s t u b . s h a r k                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                            O�00g��ۭ�-ݗd����H����ih�Yȣl�q��c#\��,�����}	f.���*���/N��\�	�J��4�n�~a.C���P!�OAD,hXn��K]x��g�m$�"A�6c��Z���$��M&��A��Oh��3$\m������@��Wr<�7K���Yc#�c%���1��Ò���L�*�I\�?�g�E�Dʢ�7F����7��&�"��G���ߒ�e-qP��`�S���>z�9v1�9a`��
���Rcݱ�%gK�GԱ�m�@���%#y�'�� �>��_��<L�q��0\%h���zo2kG�Zk�=�z%$�6rV:'j^ ������s<�.eK-��%����">�"1��?�˰��zV3*4����D4SӼ�f�.? (
 