MZ�       ��  �       @                                   �   ;���������������~�������y������t���)���v������w���!���}�������������}������z���I���W���Rich���        PE  L ��E        �   h  H     \�     �   @                      	    ~�                                 	 �                            � p                                                                                 �         p    �                    �            � 0   �                 �           � 2#   �                 �             � �   �                 �.reloc   0   � H   �                 �SoftComp    � �   �                 �.idata       	 �    �                 �               �                                                                                                                                                                                                                                                                                                                ̠�9p����c
�>h6g��T��Z9���52��?����_$�[��D��F�"@�"��P��D�b���"��"�"��'��eD��b9#�N�)��a��As�'|�4�#t���4=�
��3�L"�"14�)���g��1*��&x(�n1�7)��:ψvш���UJ�
"&��g�9���A<%57��"�ڂ_��%�
-Aϫ��+�����}�
D�kb)"�_�E��#��T���0=������5��"L�#&�e"�,Q>��9 ��s�2^�(EZ"w�"H�P:���,���sy

�F�!rV/���1�FHn���!"ҝz��l"�)^����+���H�6D��DD*Q�S���A- �H(���Z�	���))�%s��2}�h󮈍������+夂L?���B�7���WD�P]�bḑ���)"C�"v�1
x����؈Z�!�D�&��[)H�D�_�n��5�����&��-�0��>D`�n'��2�s�7:DmP=ikD��b 1�"��$l��jd!?�z�6"!�}�!�����_�)��r��!�t�����2�D��X9�<�I�%'�*��U��r�8p�e�SV�5(�H�WhX�A���������P֋=,5��~M�$���
tS�E���hM>�usL���t-�M��A)E�PQ��D��C�B=SR_f"רsƌ@��xp!u�j�5��C�l�9P�6�N��I9���>�h�NPْ��^ ;�_^[{(}�Vu�*�R$��=WB�
9 W3�j�<E�а.�U"��f�*"�
(B����E��Vj"f�|=�(؃�%����PS0p�O��-	�VA�`�h����5$5��j	_�����R������h�#�$�H���$��D ����$Wuw3����-� Q����U�}��Ph4� ��IW�U�j��Z�Y����8��
tEh�A�׽���J6,E�~C3�u3��B���*XXT��MA���I �f�C���A�Bf��#���5vWs��SD�R��h0�� ��C"z��30�]�YW	P�Y;�̉:��� ����	|��u)9U�ԙ�`���u���'Y�мD��`�VRP7�A_�u<�&�K!u3���'P�s���h��ړ? �(�$��)tu*Pj����Y~+���4�(��sI��.P�iI�X&��G�]R�!��-2i|sQZ���Le����3�9.��ҳ"�7j�ic���!9��$���8�M��H ��j�o�bS�I��`.�`]��Fh<���5�7��EjP��.�֡��D^��Y�W☂5��F��)h`��"�$}�c�e3���h�H��(@�Rd�(	_i�@�;�^�����t9�{u
j2����Cz�k������L�0�(V��w��,@P1��I`PV/���$Q^�&~~:W����}d�����q��Y\v1�nD������	p<(3{��eIMq9�!�E�ƦF�w��ށ��;�a4�(M*�^
Q����"�_B;QA�! �h�wd����T�Y�y���hT���.
"�����._S1�J`P����tIqwMJ�� �K�4{�v�h~C�V6(�a K�uc&u��]��'*A���9`r�7��e�R�V���ujd;����	�2Ȩз�����Y�4�8��[�xS,��H� ��9[�u!�ԍ�D%Av��Y��r�k��V��A��H�uM���I�Pj�PI�OT �u19�,�#�X�P���D��%�\��	8cA���P��9]v�X=<�����rxVf�d9ԉ����h����͋�f�i�b�E�ˈ�-��Gwz9;�QhW@泾�M�2�	��������j����AF;��v�3�9�Є�P�y��`���u��c�yn/�t*
�ЙK�_��BL���#	}h�%]46ޞ��KMYuh"NVMD��IJr$YQ�\AvX(�zY8�b}����UB�ol�,Hi�?u�`�ǀ�%B�K�%u�4���Ya���"�Yx��<4�;@�X8#�}�f$tR Z��$c�������u���0 !m\�#v�nd�0J�TH�$"ܱ)Y���B<pC���9�"�:阬�:{-bd/R���	�Yc���PA��RYROJ{t)�܃*���� 5��$��6�m�`��_LuE��64N��Q�Q�����[v�!/6�IZu<@�aƉV�4\Ypj�E$�@���`��� �Þ'n7��B)��BM��7�j����@�F�0^���S�\$1Y�t�z��!�Y��t�@�W�ۓ.�$ �T��f^�>��=8�N.>2�ف�MW M�LQ���t~.��+�(=����iy0]�P(c$ �{3_��]��P��rJ���Y�	�Y�f'&^û�AC��=��}3�`���K���]�|�P��u2�3�X�)^P������u�(��vS�G�`6���������� ����'�&{���!( j>w��)X��S�$W�M���jh�`�I¾o)�S!��@J��<��^�@��҄�����d=����?e�@�[�B#�#��GWdP1��+2Ud�|0��۹�i�� <�A��&�&�Mh�Uh�&^�r!%�P1C�y����$(��(�*�a<�A��L���
��B���zfY��u�@��.iGX�SC���?�J��9}�3�]�C;���%�VJ�z�<�!��w��!o��Pg��_g؄WAjh,(@?a���4�RV&#4�d�p�ODH��VjB@ y%��~�h s��mS!5K���	��!+E�RP9I�+�ڥh`Q�o���X���+V*CjD)Xb��@�h�v�.�߼6�]�m�s�B�Bs�D@C�C$hXk��$�86(i�Di/W�[+A}qF%�$H�H�*Hm��e�J7���~��d>qt��Y��&�� �TvԆ�RhR�?tZI���9��LxS�Z<�SՈA	�#68�hC��b�~hST�b��k����L%��sCC<�F�b�>�.�'�L�����6DhUPY�V3��6�FS�A��3��!h(К+�+��VeFk2Vs" �)hDV����@H�B�*@+�)��V��)+�qp��,^���H���_�q|����Ku\�%_D�'��`��eO�I���2��FE����A�!� *k�h�g�|�����6�� �����We�5?4<V��R��Z�P�k���j�z*��r��Rt�Q��4]��J����@����+7�#�_Aȉ]���puǦ�C-�� x/h�Y��1h�!Pf�~/\)W�6^;�!
9S�%�hx8d�E�]���H��lo&![�DJH��2��/;�-�h(�K@�㙯�V��LTtS�!���.�OVaM��;{%ӳin�AHh�E�<`H���E�U �)x'�r�}��e~,|�-M�M��d�_�\�����m����虡�&N7�U5��$�*����qY�<�oU@�aḕf��c��,�E��:�����������E�Q��$�9E�Ys�RM�>��:\�>��Of]��r:j���n��=6��e�X����� 
"쀪��b�;߁��v`\�����}���Tʃ������Ǧ7U0���9�?�����$��]���ʙ@�.��F()��:3� 8�2�y�u&�vfE��D5�B̊�PKǥ��QR����(r�{���s���li���E��X^9�Ns+
�=�t==NuO�BO���^+K*)[(S��$�Qáo�0�/��P�I��K�v���l��d������T �����<,;�U�`��0��!�f�%h���� ���$;��V����3�'�j%���vL���eP�n6�p s�Qh��m�aA�kF����IV�hd����L�_�(���09]��p�?V4��9���q�A��N�qK�r`�}��������N�:<|�3�'�my&�A8��C9�	u�{X��ދ��Q!B�����'f���\�	�[W�^�W}��JG՞�� ���̓�^u4��Bt+���!<�A�{ԧkl�dm�R��Bl�b%�sRJ!R
XX:+���~T�Dq3���H�|�O2��]ð��尫�z-�KH��ZX�Ë@�{�Syĸ���Jȑ�VHo�[2/t�Nu3|��B��@9t]�G���S���i/�$h��c������tF�]��>tS(��������&=��}(X�� �0υ2�لV��K7)�t�x3h��F+>?tR+�+ Lh,���#'�hЍpX�~;�~IC�5�[Qס1<8_�B1A�+�t %��!Wȏ�
�	�!��Jwu���\1NO�����!)-A��	<�)��tj��z�$!��P�_�|��5�C٬V�bf��"��CiD2S,Nd\�(��|Pj	X�Bi�P�u�m�FYB���l?�Ѿ=�fN�^3>Q�B
P��|>�h�3�U`HS.h�aG�X���A<D���	1�턯)����/)�`��L\�Ai�=@�]S�W'���:I��׀~��_GG<y���LBxh�K�M��(Z���� �,���qG2�!I�F�-������A�9����D��	��U�Y�	��(��$���R�?�0KgG��9gK�ч
Ĥ�;e���8U6O�.��E�>�����3A}S=72'�h\���t�6JZG�'��zy^��$]�M	C� :]9'SJaw�ob��Xו����$> h�[<����k��3���L�/��N(	sY���:��\���J��,�J���x�Pc�(_'�K��+����O�(%�1$kb��h���px�h��\����4����%\�ܘ�*��)�ƥXE��'��^�}���QO8Zq �j
�쇍n?�(i���DJw�e$~ce�����ק������~��@�qP��O�r��u#�M	��Q n�����⅄W�)*�w�'L��F��gk����FըD���W�v������Ĳ.�:��(��υ_髂�𨠷���������}0dW�M����e����,�]~( ���S;�wf50p3�C��&]��W�f�W�}M� �33i`0t�'l��2(V�bjA[ S���}��$W�z��2;��Ij���(��N�./AAe9�8u51�8A� �Yt%�\+�(,��S����V�w��dѱ�,���+9�Y2|rd�8�`@�AU1�.hN��6w�Ǹ���u�2L;��5�&̩�Oi���gj��@��W/�,4-�O��xP�&$F +*�I٣����� _SK@��+t���jH�\D{B�	���@X��E�	��^�F^.DF��dh���d(GK�(L���6�NEP�-T�V�0Xv(�\�`��b!�>V{�Bx!�2jt%F��!;��$@X%� ���F�A�:�s'K�xC��=��A) �%(,�S�ܦ^�Pj�L��\ �
���D�VҢ���F�u����l�L�� �� �4���8�Y�AtC+]�X�0@��h���?��䄉��ܑ�M_Ыי�`����B�+U�3f�"��̯0:��t%=�QvB;��@W//uL5&�'H�W�O��	��S�D2���ԕj��*h�S�A��hXzB`�3�T�.Њt�#�1[tMF�y�2F�&�(.�6M�ҵ}�P|��8$_c+3�"E[ƭ�(`����EKF�kz�R:Z}�M�u��-BP��	;��4��eW���J/�0����R�>��P�Y2����"�m��-,G��O�x,Fy^��1� 
�B�x�� �D1@u���M�4��Q"Rv���q�jB���ZG�Ih���"�3]��$�?Xi�&M�d���u�P���(S��$�0N�K����aŃ}�6��>QhBt'EH�|w\����"l��?�1H�9]�tnR�P�n\h��-4D�F�,=�}����>1#u��24�S'���Ʉ�Nq#�
)8���Ȃ��A6�ݘ\iD�	�[�"�Ytc)�1	���wKB0��t$=ٱ��
H1HYtX�%�!��)$�(d�-.Ng����ۆQ$8%�#�}�f�ܔ �����䢋]�cE�0؋�"}@���A3�Y��^Ǡ���ArP� +�tHudV�0��	PW�U�l �)�Y�XS'��gY��Vuj�4���e�v/DB�XCCv��}a�v5�'��n2���G��A���c��P��A�f�ܜ+���������d�B�e�ݒ�ת3¾��%[�§�NP2h��DkC�|[j���_[W�L�uPv$l�M���}�P��v���-��vl�t{�?-��_��x�'@�Ţ�FW��-2k��;H�Z5Ϳ�#V�K�GQ�hH�0��|��#��PI7��$O��"��u��R�����u�2,�����׺���[<!��5��(#�-k���a�"�_}惜t	�
1	�E����P6�$^�V��n�"h�Y����֟���R�2�Kl,>W�6�M�vr${2)X��/h�`���q�H�v?!-��E	���Z/jl��}�iSX�>E�l@
Yr�aB��:$��q��-�R�B-!�H&D�2h~��@�,��m}@���}��tJhX�ધ�<�A��j�k}!ɥ\y�e�)+��_�_9��X,�T4����o$����
��Y:�J�ׄg�S!f��L%K�g����E�&&Z�nj�'�Eo<�jY�tf�S'��!Ou5����v��⃍�Y9M ��PXZ�(��Vl�!�v���h�ݑm�p!��W#�+��8�p��s�WE=�P7��6h<�-��� �3�#DY�d��ֈlY�t����|Y��p(����Y !He?"PF.!�db�F#0�u)jw�T���<
/{6}ޅ`%�Vh��4�	b��T�����ԁ(x�B��gČ,M�B��<Ĥ,+�B��Ę,	�B����Y���͈�Y������P���1ptd{x(g��
"Z#��+!D
SN�/�6VT������0�"��Ghj)b�_�$B���"�)$�G�u�)*�� 	yy�B�<�æ	*�� 	ym���
MǾJ1"t�J�ġ	)���6'W@#D���0� �p�/�(!�X�q[P��J�Hx�-�D"Û4b->!�,�p�u\��M���EqU�i�ua3�9~3tG
�Bj �D�J���;�8�2GU@TZ	�TB��ba-�cE蕼� �X9P��m�aC�.�t<#D,|���+�H�(*PE&��4)|#C)!b(5#�U��'�#��,g�B��-D�,�B��e&2�FT!�b�#�Y����Yq؅�`��Y=腑,��X�!�g�",��Rp!4d_b8F9!@d(bD!� �H�8�L,w�BT�f�X,�C!`d�b�.�g��H������Y�ȅ��d�,��B���w�D�,wCpB��f�,�C!d�gXt��#"cx�������t��B|�N�d,�Bp��pȀX�
�B���Č,�KxeoG�^|M�#��t�%�Z ,����;��\9^���Ph�aPv���r	9����Y�Ԏ�s�u���+Bo�Hx}	 Tt;肺����m{0���~�b���4Y�}L�v}�_t�[��m�ZbeV�	������M�8uW� �c:��a�Yr�@-W��G���s+:�-�<��*/�8A�t{
u@v�ɾ)N��='��J�}$S��*Ҿ����'̐��)�FY$H�h�H򤸀�ʺÄ'Cn�|��ke@WDe߶(!�F0)W8DX"k�_�|!0�DJ9K]"�)D��D�'��P�u>�$ ���}���N�w9�*X�|ۑ�EK5(����Q�i%�:2u�
�ײ�����P���#@�H���D8u��
 SG�01;*xf
����D����-&�����"$tK�DF"A�(ĝe�%�a]H�	>����
�v�H:�Է�j[��3B���v#�ci|8��I���]u!�F��}Ns'��?hz%��X%��@�tc+#�'!^�ĹJG-��҆.�~��CW(���r�������)+ �ql,W%4�H������������XQc�I�Q�K�HYP�U��,r�l���S<C�O;;Hأ*��2%W]>:L
B;u2 WR&;��Tg��i)(l'u4*�D��&N��(��E;)�F&�DA3�9F0!� ;�2�)�6W�(�tJ9��A��d���R\��jˉ]�����_��b9H�Y=��~"��su��%~n�Ķ���Ȳ��� ���C&��5����}��ȩA����s��Fv~<;�v�=MI�m>$0���3Ya-�M�:�����stH�h����@ʍ���2�)�!���tx��@C �u���P��̗�l
�E3��:�]�u)1[�Q�ֈ�p�� <FKS��)�h�I)�pi�uQ���\EYM�C��������H�`)��Rhk�}��j��5���B�VI�v�!o-x(mg�h-�D��z��@i�`3uR
P�T�X�	\�5闱Œ�_�5����7��d�E!�;M��{�\���e)����(WPt	�!�����b��%{�Jk�d$[���S�R�'�2mJHT�B(8 vHq�hp������	!��@k��Q����"�Wޮn��*YS�}\�̷��k��E��WҲ��1)�ڠ�&f���"	�+���u���i8QMtq% C�	��$����.� ����A0 �2J�]���B�5�^x�$0��@��;	M|��v��]�$�\d$�䡼V�i��������0�B�<��9n��$�`�Q�mvP��ȍ�Bc�Dkt�D�u@����Q�N0��$N�7Lż�Rp-RzQh)<MJ��s�Tܯ�*.����3ua
 �\�;�B|�"GSN�!��(�$� �{r,ib��e�d&%����<�;�%������!�%���Vt�s��SN���LE�'1��C��!@�B�SY�t�
���fܨ
��Z�Ub�dƋ\Ւ�M��%
Y"~�kEF%�n�K�#�aZw��u~R�*��%2�=R
�-}��^��J�_BmV��5��3��jD"9M��)�Y�ԴX(���
P�,����d9�Hq
t5�
5���P�"$g��@�;@���o����h��=���5�@m
���Sp��t�j�xF���0@�|F5֙�d�<օy!��^p�M,X
�
��T�X��\�� "����Y�R�Y�T,�pP����[����V��.q���Q*���cE������S��.���Y��5,Iw����B�#��VW"�+3ۇ�Pa�I�Yz�I#;� �KW"��Cs�V,P�M�4�&�oe�q��;pS�����^�C��Z��}�,統�(�Ja����V��}�S�*��G�Ij���?�h&_�.���ߒ��O�G�!�@�|��k)=��� >��	rM�D��H=B�(��5��S!VA�C%10�H�-V�
�Ǒ�^ɊaГ@P�ʔX�ng
#
�Y��-PL`�- ��4�:U�\^u��-��?��F0t��h�٣S�j�X�6Y~T$6�\B�|�<z$4��X���Kh�BR�������j	[��~hR~���@�$��A��\��YI�(Wı�=����zI�, �����9��M��w��%�ᮿI��`���A���@�+��xh,����]���%̧��,\�9���th7Z���t2 �q�#,�"�$^�<�% D� l����[����UW����O�Ҧn�L�v�$�Q�	m�D��jq�%W���`)Ҹ��H}���U��N
Q�OP�&�9ISQ:VPH������O,(�ZF���1�6�O���$tv��ŏ "S鬒��!͵x�A�jg7g�Ͷ"�=�˭�׹6ikQ�>N3�}�~L'�F	�æ�����1t+ad��44��eJ�(�h�Mu�v�����������rGe!$dSr(}�B,�c�0�4��p��#�����N�tV]�F"��E�d-8�h���� ����x ��B���|��Bv��TB�"V��B8����@#̐D��L��~�PY��1X#ؑ\��\?dB�+�uJ�,�Y�[A>C��4��/��]�B3�@?�ᗘe%8(�5*����&F�J� ;�Yr�jRWw����p&K,��&�b�O�B8���-&!<
���@9u@t�{$�2DHL���Z�,�Ѡ��u�-��"��O���!
,��u2�ᨸ����T%Yʾ(j_J`{�yB�TG�BW@8A��(]8�����!K�L}<;�Kdb��$�&� ��F!����B��$�#z-:������7��^߅x9߅b&��i8N# O�|Bl����{!4���Gd#$ a3�(1.#SPz���豈v�����Q�'����NW,n�� �U�9���H�AE*!~7���xK�쒊%��h�g>������0��O)u�P���B�Ҩ������jw�H=ё����w����o^_�}�q��[l��'��Մ�|�G9"��m+����6D�Py@��I dC{�t��"/���ܐ*�D������]��u/���˕G�'�[T��֙��-���Vn�u�`�8Z7��P VG�-`���-�F��ԯ0�thQ(}�R��V�E�u�G�3~��=��"�"x���hO)3<!֡�C�~c�0Y��DhC�;a0���(�p��I~��u	�U	�i^�X��	8��tpbG�H�Z�;���[aBδ�R:Y�n��!>����#����\=�
М�@��9�������[�e��$��ȪW/���2y��3-��W��ǎ��A��G��n��jVa��?/z����P���x�|G�[���߬x[-w+%v����y�V�D��XU���/��|)�O0�D�(��̉S�U-��l!���z��있Z�j��M�O�������}�w/ډ$��/](��) ��t@5c���+DBu�Ð�ȄH�	1�ö~x��D$�<��d쯑0*#È���T� �l�_�U!*-�*�a�P+���H�j����-���1�0?�%vt�Pt �Ѷ4,���7l�찈�����@D��a"pL\�"6� �p�N��8"���8�
�\�lD�\�i��[M�:��K�c�5'�^�
F	�sB��URk�����Ji�OƲ@�̾��	%��M�T����ޛ6#&�-�F���'�c����O����=�����H��O��Ǵ蝰�F��B�t0Bjv2ĨYjD��P�;֙o	��n�|W�@A9�]��c<�H'V���֘0�EBb (W������Y!�:9=���h�;H����56��E����\�����3!��:c]��΍7LET8���25�F�9Kh	P�)���3ҹ \&�,� ;F$�ZЇ*��HYP����B�5�(`2E_>	��+5/��ՠ�Nv]ּ 3�&&���$�@��%ة��,Pe/��ڙ��!8Iy���Kv�&	�u�po5�R������\	8>���e��R-���%�����©M&��H�G_I�Ⱦ8�' E��
�s'���Bu0\��u ��D8Vd!�a/b�	 e���	�i}����	�F3��u1w�	'tu*X�C5�%�tNfAN|8�6�P�I���[28��k����%D�q�@��8J�%|F�*�f�K�	� S�5&�c�ᕑ)�e��W�V!��-p�ޝ�?��(���[�"lJ��F׵�E�p�O¶S�fe�@�[�5���!�CE<O/�!^�č%0Q~	h��tfF��n.<bx�qnB�� +��"Jp%V�O��'J�DN���ḃu�#PV+���9$��
f����_�6i,�Z�k�H��dV4�N�O���N
�Ua��-��?Ĝm�拄c!ܹ�g�m�b�Қ�i�Yf�A���=q(�"�(P�L�����kU���譓���z!)��� �Xg��^qn�ht��sA�r���;�~?#Ag'QP�,&!�k�-�M������}G����0"\���ł�Ԓ��S����/�ү�������׳�D�!<���*i�5:�`/�UX���~`��-l��Rv"88u:u�ԟ�X�0��Ъ�m-�wh?3D�#��p���ӑ�t�J-H0B�%�cH��,�D�j�ٓq'���B(�"0�"��o�B���T��u�Z3y��3}�0#�!1��sű�
�*
�9���p����C�3�V���T��.[�{��(���L�0��=,u�6���[dM,����4��(�%3�tkg�O �|D��}?��G�b�-t�%kE������>R���
u���Ȇ�u��}}���&
5dZ2�<D�v	��PuO��q����fx9��ۤ��R����}��,*!J:%� !� �h�&7P�e{��ص�K���ꎮ09a�7~D�m <�}�J-�+ �v����Y�
h�?Q��C�Ʃ�;D�|�fD�a�H�������;N�� "N(q���D�Q\��Y|/DQ�;Q^�}!��$t�1H�"2�|'w���]��U"\�EzmԱ��t/FV�ߤ��@�Mɍ���K@��ؑ4K�?BEVtk�G�3�	��|�t��P�\�d�FYPU�T/dG�|��g�%�r�v}�;�8L3�dj�#S��<���;�}*�'r+L���G�[�o)y���nBC"W�D
59���C;<�rW�)�
�̔Y��bb���-Ӽ���ܨ�+���t�����y�o�a���J�7�D	S_��Ŀ�Pf��b
�H �H��+��#�:�'�(�^�*��-�Z���L�D���Wہ���S��8��������%����0��!�P�O�9��B��7��A�U�,���X�]��%��#w+�U%@����WA��-d�2�)��3��0S���&@;�r�3�k݋�Xw�D=�G4P52F;�r�W�,����P=0��"��� *��9�H#�G�聴X��B�����rğ�;{�S�vOG#�6LH�����#؋�v5��u�|��o|��	�����FW	0rB���rJ���j�K|Z$�Lw�o����4>��F�_[����_b M{$u7]E��jz�����|���d1!r�8 ڌG	#��(��b�94َGz{�G�#b�lȩ�JTx07;�~ ���7 e)'90�Ku�EN]�����W׿v�B�h:S�U3��{2�fGC)��_)-��b*��:��(F�#���R�v�d���`(v�G�#J	���o�BAwx�A��#����#�P�b�3�j����.]��Up,�ٝD/2�U��_�Z��(��h.Ai߄���1���h�1~���Au�#:�3�#Sb$5|�h.�kpf���ap44j#9h'�@|e�PѰ�sL9]�u.�
�����l��B-Q|-������9�Ny�JzƆ���0��/YS~�5�Y�@����T���s�Y�h�Fx%��׷�[���E�\�X�2�S��(r1�w�B�P6;�s"��+��x<v�Aw��������3xX�wP��+��U	��#��c���>�A������ݵ"Y>�p�����vmqQ�$1���^�EQN��z6�DS�(gBx4$���V�����T,��$}����D������H\�_��РO��[�tM�n<��wA雌QjD<Ж�cZ�K�*��N�K�����"0}S�Z=���>���(*#lD���f���i � ����9T*�(�̆����Yja ����w��u&)<�9Xغ�F nZ����j�&Կe�	��8�j<��=��Q���T���Nl�I���9���^V��z�i�T_I�Y�4;��U�v5P��d��t�
Ȓ����h����I�T��H�Uת+�E_h�/*#�!��yp
-v��t	��3�$��o$1���	�$q��r�#`������%)�d-(�7\�2�U`�uB;3��}�'������	��U�A���x�Ѣ�+w���S")F�D�R���!(����	';^ª�E	)�).��y�w��w~�qR�Gb���4��+�! @��������D�2��Є�t�P:VW�����E�,o������N�����UF�Z������jIbM}AG��>�Gz��-{��A�ԃ�^��tj9Z�}}ہvx�s#_�ȹ�����C�!���!����S��R�)�U^�@�6w&{s�|eɂ�HP�d�kS���?�3 �e���,��<7[l�YC������`aa[�/v�	��WǈYR���`�O�'B��*WE����B�0Nz@��Br��k�u,g�!��B�.u�p �@�܁� ��A��t�b��WVNB ����A.U�"))|��;U�FB�i'�C��e:���HP�/S\�!�.�8EU��^ns�R��N�o�^
b#��
;$h�M2�X��D��.S3:pKPh\��(�>Bp�.��k��{��aC�8�J ���3��IV�<�
r$8؆�ؒ��,�x�̋0�Sր;��tkh䛄��)���Z@�5Eh�)�
�r�D���N���M�l��y@����܁������tV��"~�|�`��D�
�@�u�ZSe�Up,P��-p+�Q�L� ����r@����Foh�8?�Bn%$e�֑��HPV9�����tR���$�q&Y��k�����d�|��,G����5�w '�|h��$�'#fXĊ��Wĉ}��?	D�td�@Bz����Ӊ&���@��A��I�F�������܅�����Ě�����\�u��]��ђ�v��\[`R\�d��\;�tIF_Z���0��#��<�Q�[�	Im]lb��
�� ����zw��k����34��l"�
��P�HtHa]����]>���C���!�����³8��l�Ŕ���"t/u�Z��P�*e# *PCO�n�J�����k2^��0�Xq��g�)
@��KD�
4��%��]�UѴ2&��������$C��l�Ȅ���;	B_UϨ#kb�\v⹫�v�d@�je�^�밤+��˱Lx�X�C�i��c�|�J���V����e��jQ�h,�zP��D�S��Ɇ�5H��]ԡ:Z�44�֯�y�e��"��,E 2}�����j
������Ņ�jA��6;Y�.M�,�	@bb߉,_�rin���]�|�jd'l��xT��x�E����U�W��L�|!(�`;�ur���G�;W�X�u�Ӑ8���M�n���v)���9tA+�;�r�u��@s����J�.;�~�	Sj���A��D8�e��Sd���� R�S�e�v:@e8t
����&J�s� c�P<A��2lC7rz�Q�����?�k��+�dT��z	hp�S� ����;�9���hLD���%D�E�8�Ih("�C ��h�C��d�<��d�Is8�B�!���$!Oĸ2�V$�h�)o;ah�	�K���F4�xB�Cp)$a,h<��4��rvh���*DKFh8Wtz#'�i����A��+1��j�*��*�#�g�!.A�M3*'M�f �/���D_s���Ut�+�FJ�WD����2#���4�?�W�84��>�7�j2��C٤">4�]y�� (��G��*����봗}{��h*��1�Ǉ8��Yϲ����79����u(�t ՍQ�h|����e��(��H���^)�P*98�I�\�m�*�S$�[e�>������'�V-�@Q^���BWv[����~���<~b��Ts�h��o��
����r �WY"��P�d�]e7� h�-a2\3\�]E�U4AUuh8C!���\F��W��G;}�Bў���cN��_���΃CVj����[���]����_억A)�8�����6���Bu7�'%"T��Y}���]�>�gbckp�8���,�W���D� �� 6�����-�����hb��UE,-ܓK�0��tZq��5�+�-V��D�^��]���_�FuKhlA@K��-�-��VA����f�a u�D4�R$��*��~�e��и`���X�2^+4[_d�KЄ麧^�QPS�jT��-�cyC�{V�i�\�������sQ���OЂt��#'�]��l�?��D������/2�x2��5t&
C�/X\�̕���x>��`(�"&R$���,r�J�[�SUx#2�`�q�U�@��D$ �Z۵�ϭ�O�<���1�V����+�"���ص.���[��(�}Yl���i|v ���wPUhu�-V�CH�:���\�t�L7�Du��$��$][>ږ�Cb@B�"1h��^�س8b"+Ä�Ś��
�H��w�r;���$d���q��3��@����Xw[r��Ps�jK�$�"w�G�B�;D7H2�+"&$!b1
,s�0 +���ׯ��y��d�����z��A;����D쾈�(����'1|��W�&"D�2�4�s ����)���i�,.
u	%��FNZuE���<[Au3,�"��	�1Rv�u,8�Zt�/l��h�M��KV�B����iڸ�	jn��(�AlT�<E�<���a$�H@�jF�hx¹S�	��qT��F�!l D�j���E����W�r��+p�S��M4��s<	��fXR�"���#5���
�XY���
�����@k��!��]��}�_c28~'tr���#��H�dd��S��N_�h#��@������d��d����z��� 8\O��u�W�ğ��*[��^�)�]�:��]��D+�+� �>����8h�fuuX��\�K!������z[L�hp!�`�in%dQ�i�1�XHP��`[źk�)�q����,�P��樞 Azu.%Cz�(�t!�X�͘n���e�/[�d��;W�>��]�vw�0��%a��H�����iu�\�o�r�3�V����Z9]t@��&
�;��}��E���-W���B���}��h�uDRSK�$��t+��ѕ� h�þ�I�T�HO����͈�l����)�-̪B�
~������u��]AZ�L�d4T�i>�fHQ	��v�[+�i|���E��B���?�F�s���<rd<
H�dlx
��S�[�D��v�_��wSYM��hkW-d'����C��W�o���+����b6�e((�	u�]��K��|�B�_����lV#
X� V��f��Iӓ%�ݏh� �F��:�{{&AٓB�I���SU��|$�=伟K���'��κ� B=�?�!����+�;�wh��6�g���8�0S�c�;�+�PUG����R����0Z+ͅ.��Ӕ��&�������A��H�Kԕ�ҔY(ߥ]9j@+�5�IS�Wn��"#uj�:���F9�x�Y�8��v��I�O*�a>�e��@�2�]'�$v��'���	5ĵ�F�u)�!��?�`�+Y�� D
`g�v��	]�3%t2��Wwd+��ȩ���X%�Fy��XV�@^�4.���8��u��P�&$�G=� |�3*_�ê�i�C0�~(��,Š��f� CJ#�8�\�E�i��^뻶��ِ���>6�A�I�;c�&^!�v2�6�StF�&G#?t��Ƶ����ȶI�������IU���7O����j�L�<����i�� H��E�	kz�ڶȰs��j0ŀ7�	03t5TjGG�a�77ug:�$����^��ܒVm9��C���ꑎFW8(�jp�u�#*�&u�c%�7n�iD�e�_�l��ؽ����d�U��Rb3ۖ�U��H�}�
Sh*��%C�H�2$�1���WC�_�)�#��%LV(:H��U�{`uR�'O�HW�*�43�[��]Uе�py	�6FL�mJ~B���Q�KՊ���~R�aWq7�w�?�tN��.�(�9�j'��p���=d��KۨߧN}��餞ޥo��%Σ�[�~�|�/]	�c@�F�kтWۑ-0q���{Z���t&����4������h<�p�0g�1wh0LT�'Ih֙>��{^���8���c�t'hH���.SYr���(t�!E�J)XOH+���HT:�v&5+��C�����]Q"�VhT�CKN��.cRB-W��M��e1"7_M�78�Z��7�6�̻�h�&��#*0��=�&��a	2E�
�.���~ã��Q`*TX�U�d�h��L���ӫ�qa��!�&� ���~8�\��Y�~v�+�bm��:W���Tx�U!��5���@j �|��Y��^��b3����x��G��j!�-�+L�7tT�j�C��b�Bj�h���Fbf��*Ä�h�2O;�/J���_0w�O����Y��AB\��
t�h�Ub��9D��D)��dC�uh�2(�G����hS�)!�K	�@
p�E�c%��vJ�����H�����Ž4�#�o�Z1W��T%T��\�,tKhx$�W/���?bVT�1�FV)hl�0��N���\9PV
에;�W�!�p>n*�$���wK��O �6�kI���hK�W�/�V���4���bE�V�M�h�;��Ma(�>�>,�w���Nx��a������L=j;}�t!�d};��,(��B��w�(�K�dR2�)��7
�<�v�eC؀y�K��B#T1Q�K3�I}B*�u[_
h�.d�0���Y��r�d�ra�,�16��|�h��H2�M��P�7�7D���1�4L7�BJ	�}�Z)h ���]��kG^��qt��3�9�|��A �z��)��.�P��IH"(@zt�
#�DH���I��U3x��j���'L�~�{��Re��w |;�@Gj�Y����a���)F;6~�Ԧp�vF�ގb�V����$�"���Z�O�?0���#jA�P��%<���|�*aY{���h-D��>'Ѓ[�+��b��1�A�����.Pkٝ1��'�x�b2X\��;{ NF

0��UG��Z[�oU��'װ�k�u�ق����h�	�S����A�~���lq�I9�p!x�t���XF��b�p'�[� "L
�l#KZu=�h;�Ru-�Pd#�d!`"1�XEi��|�W� �!=��g	;s����F'�eTv��E#VE!�A�ʃX���_(, 0��QG�+����S��*p��9Pf�h���=�[̍9�5�GSW\,��@�0o��;�}.+V�嘈�Rh|��C2���IOu�*hxZE%��M��ؤ��		�"�Ղwo����h�w�,�$7^���R�U������GO(��e��NJ�_R	�D��'#F�,�Bi�%Z��'qP��W�����c��Q*�n0��Q��N�h��?��~�G$#�!�Eu����	A?"�O�0��4E�AÊ��	. �VjX��/\P��K �����l�������!����>~=�-e��%��K-ܚ��M�����5�`$�;��
}43�7p-�z��\dbL��C<��$dpb��B�)$4�)TN�#����4D�2��9��줰tdL^D��<B�xd4�",i<u�dxd�"Z<t��I� ;u
�i�93aK�M��,� 7�H���[����)-El�4�5>'<�B\�1LL�8�"�VH�!0��� ed"�H'�B�#��#���@�8D�I�Ha�d�G�����@8̅��o
�h��u�ᒄb���`���H�R!Dͥ���r?�9gxh?�Eƙ|TlC!@����,e"�7nD�'!��Lt?H���2 1��naBl&xQ瀈�0��#L#�#���!�μ*�hRu#�!dɈ9L`����Zψ�P�C@#�0Č2�I��!'���C�)�'�)��ȘĄ1d��HP�F�!4��4�e@!N����'U��1����ԏ(� l"�@d��\'��TB L���G�#�����0@�G�p���[д̹F�����4r(�"��l�P���9� ����pR,��`4�F���t$D�24�(�M0��&l����I,�A!4?��1T)^�,��00l�d�2�8�-��&X!��/H���D0bԤ���ȱ��R�1�t�4C�)T���|7d2p�d�!p�XɈ��$(bH��C@#�8���02�Ni�8�C #X�ko�1P\�!���Eȝe�F�!ԗ�t�HlĴ2�1��C!���n���x2�[0���(��"�R	��p��!t��Td�2�|�<�R��p�$���C�!(����d�2��5!yt}�8�u!Xm!e� ]"@U�DM��E�=�5l"-�"%�/�� �mÐ���S��"#H�$!�eHt�����C�#4���'D�7t2����MX����xd�b`�g�B��5��@:"A8	��0e�(�  ;˹��Ǭ�Ǽ�q��U1S1'���Ѣ�|$����h/��:Ɏ:8�D F�)����xT|�!�����e<����]�0�#���xĀ1d�YDĤL�5thY}<2Q�I�'����b�9xFD�Bp�h$T�R�_�b�����شVTJ�����XE)�N�!xb!Фtb���C�'�0Jx�Pi��>�!�����)H
��Q��[���b9(�r�Rb�9�`��CD#�(�\9���$�f��\�� 2|��t���",��ǈ�pJ�(�B$���,|�M�HJ��V$�*�F�!���t�HD�|2��$P�uǄ�1D�1K��0d,(p�>}GT!<��w�$eܘ���*�����L'�-��M�
- vl�=<��W�!@�<�Ac�A��$.�̗HDB�!nqd�DEh�(/���\�PL��?�{�o�Ӣ�ӣ���nxuNΨ��S⧪��0P���n��[�1���;U�� ���=�|��ۅ�ͻj�*k�	[�~��DmV<P�7)uK�F��Ô|�WX�i��^�t�\���v�����D$(��d�yP�̛��;��ﳰ�Pv�\(]D���C��[��k;}��'���;�7��.ehl�U�GR��d7 LV.tֺ����;tu=
�ǆ�m��A�����
����J�Z�đF���2�_fRSb���g.�QW��.��H3u���P�=�b�}Tݥ�$
��}-��\������t|#	�,��28w쓱�0k�
�����>l3".۵i|�k��ЌG!�r��KJ�]� �u�h�Z��b�kHntlh�#��uh�,��+�$Hh|2�Gx!�Iqu$!w@hК�Gd{N�/�����N��,P�
_���B��ul
��4$]֭�X��#T�$��"�����6/9E���80S��+�� ��ޓDꍮ��88p����,�}�4�����"0}Ss��{��Y����""�9�:��;f���<6��A9�K��;+o�'ZN�^�1}����"*�!@Xغ�!�*�c^�^0����.Y�������p��^���i/�.)�0�h��*�ye�)�
��pS�)9�A�D���=(�
�
��sWv�~���
��f���gR�|(��P�Wi,�j�EMOP���EVčM<�s�l*�hߜ�K���R���+J�:�W`!,��8�(�
��td�b���$0;l\W� ����^���讪������SW+��ԳϊEP%^7Ӝ��g6�;ߟާ�΍��da�!g��#+D��'G9ԯ*�4�)'�i�u(�*�	��7p��_�y$*	O)0t2�<�֓hh]MIkU"e���Gc�%��8���[*�0�/I�' �4YY�ׂԔ�ȍ:k	�ʖ$/���u�(���-�<�f�(!K��'�b�UY�K��$�7�t�JV!N�;���A�fbm&(�VZ(R"��� *�y�t߯�'�%~��uc�
UL��)(�'��A�|U���X޴��'4&�"���=-_}������ښ��;�&Ȟ��U��mD������ d���B4���)}����?� ��DH�U�c?���F��#|Y�d�cjz��X���o�)SL%Zt�UZ���"5N�I0ZW�X۾ؤ[Ha�5+�}?�[ڸU�zj61��޸ϥ�=�$$��*����+�jcdl0?���NL�1t>�W{Ȣ��V����ԉ8�z��Mi���t{I�ȝ��)Wu;��8�8'c[�HD�h�E� ��@h̻���D�4�e��z@*(��\zR$A���x��@%S�ٜ���>�M��@�^[�_�V��cL��a�Sё��^*�G@��]����	���D�U�C�: R�#���19tR�>��J��7SdYT�<I�1�	�V%�;��$`����=K�[N�v6��a��������AՋ���N���B���(���2�W��^��2P��m`a(!E �S!h��(�Iψ��W㇄"�i�=������_�3s/�������K!��&-TD�9�"�r޼/�x���m7�$��#��V��tYS��S������$i�D�����2Ҍ�H0|ş־kU��S�/�dSs�b��_��|����ӫ�9{����(`;���E�BVe���>9It���m[v�,�W���D�Z� �W�6,����`��
I<��>������c3��<;��Qt֭4xIPy�W�^��}���$<��b��$����j�g�	"3��IJ�q7�j" ^�Uí6��]��Dc�sX�\�;�J4<�c�;쇑�	h�h3�Z��E�󫑁舄��e�һ��	y�4Z�7pj�:Ѕ�'t#~��G6�ta�;׹S2����k�r�;���~���M��I��O�5��*��Q�����|���"�^��ITW�ٔnr�f�S"��5O���a���H��x0�t	�?�-��LP�C�o,k���B\c��;=>�ƛ6P�������=�Q��S�O�Y�ۋD�X_�0^�F$h�/��8^
�0��ɰ$��7�H�>�I���T>��۽f��|E�0[R9^IuÃ�|d�Mˍہ� tP���-uQ8XU���Ƅ�6��(C9�x:�3�<h.�{. ru�P�Us�n��XtL�N��`�}���H�s����Es�2M�)1P������$"b��6��Ű��������6�e�7(M��h�sk���Ԑ�ŕ�H.��D�j�h}k�Ja�;�x��2\��B��qڱ�;%R��'�B�Z��U��q���E�/:�ٯ"���ߔ:���X���~��wRj�*�%8e��c��vh�]\}������s��3����"tN��g�,�$Yv@���C+V�,�TT�mӺ��!\�p��%��Nl�n��aN�XN�$�1��LthD��8u���hA�S�ĕ0�h�_A��Z(7�=���*~+��쮔g"/Pk��0�hZ��>� F(;5,(|��7�5*i�>)/�L�tvW�Fm��!*hl����Ws��jq�QƸ��tʧw
���߹�����,��,�B/�y��x܋8�� �]��!���u���P�����HB�C����bI!���\�9�LXJP�&���Q�����$P:�s����CH�\�	�t«�U-~iV�cf$�bk}H�tg��ahl�EےR�	�V9�"K:���Ae�&�XC@�l
aA(�HmhЫA�1�>��{��2�0V��UWh`�i����)�		j��这��|}��^OT�&�EE")�3��NU:�Z���d+�Ԯ�jk:���hrF�>$uQ�]X!h4R<�jI�=�0Y/B��rQ?��v#�H�Pj�:�U��{��	`����5���InS�Vn5^�7���5kqN�حgQtqM@@|���^�(Z��}����[~�ĚI�"�I��K�:l2��+�%/9�!���E�59S2$���_4��Ʃo�ד�߅^
�d��3�P��	�`�]�jZ�xVh���v��9
�1���7�!�	�)�7���nV���Fñ|ܘb��-���.cb�Dd>1�֡�s��ч1X�R-����!��D�5�ۛ~�O	W� �b���53m+��	h!,�d�<��[���b#��J��R\""9��lvT�)�'%�PD_�aL�B	8�!H�DDb�@b�/�im<��s�6+���9DD3��9]�V�9�t�ؼ@b�1u�_qKd�̻�ko���Vo�p��S�v�+�t��u'�:�dEtRP)P/W
{*�P�sS�XE(�F1en�´�e��	/�+Nh�#�:vq���CZP�O��n�q*ܞh���4޸�|p?p�}S�X���%ldHs�u~����=D�O��&"��KP�����ZK覒�c �td��j�"�Ȫ�62»5��J�ϱa���s��[����V�Z�4C"��J(0<,�"D�V�î�/OE,!T2$�"h�E!l�<!d�*4�m�伤X9_��v`�[��V4NK��,�S�(t�)��.�� ��-)u"���C������,%���t��3��;�r�-�������+�*:�N�u�+g#�HLVBء�MSG�lTp����� +V�"�F}Q'�n�}��Q�M�-^�7����_䑅iL�^�!�ػ'�Y�%R@�<���J�S�	���!Z��;��_���8V޾Y���H�N�-;�},9���	�$�,��
��hF$������
�@��C@�}��M���NPh8���}�|�C�X���t�Y<C��p��er=t���Q�"��H
3��JJ�����!,�U�VRXj]2��^��|uJ���|@���hp�yP���*a�eԠ��R��Q�B��F��Q�zjVC�<�}��`%�B:���
�B��G��(�<!�EZbj�$�6�nFT�?��(: �h��������/1�	�
�*��Y?�E�A�����P�R�<���>�<�O}2PV�D��v��^�� p��d܍N@��s43Ɂ҅�v"@�������k��,��!
AB�;�rހ���;�؏�~�Kb4��Tб4�k����
��Bh`�ӈ�ͫ4-P�u�Z*h\$Z�"�.�r@�I0/� ��Z��[�$�H�tjab�LuL5-XۆK�3�&v~��0�����W �#$�,��N�o0����4���)j�d�kHNph�=&�!���Zb��F���\#��X�և�kG�XGu���Е
����f���'$�� �vC�&�ɋD=a*Q-��Mu�?��@t
�
.�_u%*��-8GF�;�r�!D�f��e�>x$��:��0-Fw�hr$� -w1{W"6�R��V�S
@%P{
�D��?�R�S�4"p�t	�(4=���E#q����EMq�,,��-Pݲ��m�(	�--R>�@9�q���8�\��5˴�ZG��%�؟��l��2���"�BG��f�(�G|�u��ƍh'�+dQ�[��:�'���Qr�|6vm� �j{�g��Dat���<���D�!a2i�g�bs�ƥ$V"iT:�ld1��b��Vj���_l��A�8�/1�u�Iu;����k�鯠E��5D9�)��$"�N�$�,cB�;Q�~_^+��+�B���(;åZ\�I�1���k��rӽ,*���!�����d�2x,td{"`"@cX�B
�R@����:8�aD)(D�(�$Ǝu��f�;^é8F#ӷI�/
=Dtl�RL�K��J�OB�2]�x�=
q`X�F�@�8b4F(!$��"�N�5H~]��z~-j��� 5h�k���>`+��T�D��|8B��(��Y�d��)*�;}����ԙ�s�K��K��w.t&�?v	u.��BI��Y�<��	�Xt#0��T0$��R.�	/{�O��	�����#<���W����L�l�D�j[?�D������6[��$�����"hXEVS=l֌�EN������'O�F�K��;�1�o�:6�D�O����\�FQ�����~BP���_/��?*>���kUaR(-�'��J�Ku��������%;�`�t|Q9��wK�h8��[`c��"�@ZΥ� �f�����zv����(N2t

�'
�?V,��lB]���(���D-Q��݇�RAxA.I�<��E����[��6%K᎒��(d���R?�4���;%T#�W �VP���D�̷{��-��<���Z�"�x��9������v�I��>,5DD�V�.B	���FJ�?h|�iX���"C'A�F�;u�r�˪��(3�"����X����ԉg�W(�MG1 �!��\"��~8;�u�Z�pٽ9�I���*%��])�B�!Z�GF;}��l��E� �/�^�2�J�_7��V��HX�^��R�R�bV�.&t�:&�$��eV����2I��+�bV���0��)kU�[�z�tV��;�d B�5��;��9QII2�>�Rh�VSk�L/H��XT5�M���EP��I�!8��3�$v~P��Q�/�&>
�;�r�p+�ȱV����$Po/u�M�ǚ�)��U�d<{j�/��Eh �����ы��ǜC�� 8�Z���j	~KY��H�����	�0;O����H"��q��c�����<{*�7��o���ޘ:$[8�`3Ɉ�P5;d��@~���
�T�u �A;�|��FtnF4A�_�O����yX*7t�jr
��74)9B'�)I*!�R�WH��Z��t����:�..���I/��ȊC���h7Z��9Z�0�����B�=�� �QJ��2 �Y���wōf��hk�C�ᡡ���e��$�V��*��`� @��`K��� ���vܼx��h���.h���t'�{��]���h��9y�&!��h�^t5$^�	h�t�ܨ���T�&Ed!-���Kb$���b%$Y���n���A\��� ��hU��4I�_� �C	h�\
��
|�U]��<��[�����$�
���BUW������d��J��Vk�:�Z\�h�� �Yt��`�V��J�ʤw�
��P�c��ߺ ���1��5.{�Ѷ%y-՘d]tj�bOS����X3�Z�}�4����W�L����u�{��*��fP����܁EV�4�7'�̴hM�H'@���a���H�݋%����U���s_�kj��d1��w݈�1���QI�E�������Ll�B�uP� ���%[��{Q� ��$�A�S�gN�'	J�������ii(h���9p�hX��E��c�9�iu��'�k(���`��wW���A&�N�W�T��VuG�f��t-h�%� ��A�*���FR���j`g�l��QI���Hd�(F�O�/^[���a��a�_��CP0L���ʽ`�=p��5t�x�|e�Hs����P�L^l�#�(b�]�>q��;�Cb�������!YԿ\������h����@�jPrԽ���`��tigV�.=K�1hn��z�
4�A�4���^1�uj��6D�1�u%�hbPQ��i�Y�X��5eBK���V�pIb2��ͱ�9d�q���ao"D*Eܔ�4�8zV����&��$��a�h%�~jr���!LM�%AB�V3�bW�akD�K4���r�f5�o��\wÌ*d���hWV�k6���K(����uJrs/�+��{�j@* ���� D�t�M�Q+SP;@�Ј3��-��(��� d%s�ɍ���ܥS/�/��� ��,���f��&(�
H�읥��{�3s�ٔ���$\�A�2\�r���_�z2��ø�Y/�u	X�ѿ�h@���^��	�_T�!-u�Ԅ��<��6�Q{B}?u�)$g��<ΰN���C˲��(�"��VS
�h�Y�X�y��y�)�$g���U��C���1��������������!�x��l!�`��X!�P�}H!k@�hD<hG�F8�5D4h#�F(�D i��4B�#D�"4B�#D�'���
��;l�3`���7`ҼB����Y�T!Eޚ{��h��J�y(:hd,H��\��ߐT���L2�TV����-ݒ2��"���XghC쟟T���F��r�L���C̟���䮎>$ñ�8�q�gZ���h0�"��(�?F�ѧѮF��#�Ko!lQ1!�)H���"��"(}<�D�v���/Uz��$%-�԰�.� +󫋝�%h�>!fʯ$F�]>�����}��ٜ��H
�Q�{}
#'|<��_Kh�_�G���t��u������U| R��('���x�^�h*��zvl3�V`tඎ/Q<�r�b�at�<!�V;���8����5��&���'%��F% _��ۄ���1A&j��k%��{�Y@��'XZ7o��$i2��&
��H�n~o������n�l%ԊG!���R\2;�2�/y��D�*��ϕ:�S����T�S!R ;E*
+�%!��8�K�bM%��kv.��P*���V���
B12C`+_�	�G��tx��
s���, >ɒM�˔!�x�V��W��H�;��Ic@<7���U��J���u4!9Dj���U0�b�_�t|/��&��(�t.>W"��]����D| �Mj�]��?�HI>H���9*���_2�S��cN��1��yK�(D3>ɍP�U9t	U����r�u���s�.V�R���*�":�W�Q'~�?%Su0�t,RW4/VW���7t_�`���ޙ.HM>�+@&�N�;DB5F�YS]D! {���@�S<!$%U�1�Y_���ܻ��"^̵͊��'T�VB�8�l{\�@�hN٩�D��V�(�T�ኁq{j{'30!*f���-�i�AP��jWia'�(J�v�i�ֈpb���\u=|"I�����d[�� N��$S;�VL@�f3J���
=�Z���	W��Ґ&��u�ܯ���$��]_�xėؼ�Թ�$,)&(!s�$u�$q�,����`l�����j
!;��=,�A�ˆpQhN�������^���r�>�����Cߐ�!���<�^��J�$l!<h����/��,��a��&���!�^��+�SU��Z!���;�~g���}J_�o�[��]��A*g*����;:�vL�$`NMB*��Ŷ�B�CHw��_�ŝ�U\��,�˦A>{����,7�C��#*A�L+�y`Z��[�j1i��L�F�;�0u��~iW�����S�s�UJ�%WC�����*���l3ɺ�����Nʔ��Ȝd�^�R�B����Pt{ǝY��ݽa+�pb~$�dCdE+ ���t氆���]U�$z�}tSU��]H)$�U��-��rbv}�Ϳy$��'�%�9�R�Q����J��Tۿ2�?(�}؇�	a��q�J-�n	���>�P4�Ǔq>H���~��輙'��E�+�N/j���E�.����H�tx���SV3�Hl�J�D�b�A��J.+��Ɵa��Q�W輳܌4��� ��@�;T`Zu@��^v&���B�ú&A��H)1P;���(VB)^Ë¯�^��@��K�4���M���n��~  �Y_���3�;D|�[�;�K�!�Ĥ����9��+�l1uP��:�������8���ֽ�&��]DZ(=�O�"�Sz�������f����;�rQ�����C�]˧���@���:
O*3Д��{%�|Zb�-����g/��nk t۟v��=�~P2���18�f5<���/���WUZ��R�#��ݟ�-I�G/ę��Ǽ��j4X"3�-@�֕��:�(�������{M���%�����R���9���	E�"zV}�E'\.���K��wE/4s�gK������
�,4t%���PK�WHS�H�Ǫ�4�zz�d*~ �\��w�[{�{�3�9�j:���1v�d�Y�Sne�_��$Z���@�@�,%�H���%�~aF;,��+��A��7�3@-~�^���E�K�u)]��&��t{�Iv�Dq.��<���Y�],�#X�Ԥ�tC+�PWS�?�:�� �$p0�&m"�7,k��'&�<�c'�v��0�K��gʢ�[lv��G�r����(_�
!}�X�9��uA�|�
ò����]u9-IL�3=-�,�A�<sq�I �:�}<]t;9�>��9���:�|��.Ԇ2_�&nE:�_V���\��������:+ϗX���Q����N����}��蟠� ,8t�	��?tJ�*G�@�H �v��!��.�� �:���'8d�foN���` �6�T��u}<lb:�a�:�t�:�[��Ɵ�6��4�P0$�t�b@�_KhN��ģ �o�U�Ӆ��8�(N��$X�	��t=���8 �����/��
�I������,D��
P�W�7c،�{Y�N0F�뽀H>(BT�%�%��
�:
ˁH]X��%�$����A����&����ٳ�iuyKwl�_~O����[�Ru�8�h�b]\���߭/W���S_��Z�&vl�3�P҃�hlK����}��_b�H�A��8�pVY'S_������t�Zպ��^�b�y�*�d�y|*����t���w&�էU��8�j2���HϰqU�;���u���0=\��C0�F$?Q�&�	t�j{��Y�����p�,F��N��M�;�&r��@���L��vv����`�����SD�A����F�9�
�ÊVC�1�"NK��,��!p�@�u����$D��e�����gA��K�Atz��)_ue��3�Y�_�G�%A�f���GE,��u�SuΪE�0r������t_�e��ٖW5�1���v{�Q��(q'�Y�>PC��J�Nt*�)VP."�ĩ������4>�c��s>'^_]5Έ0��f'WB�ֽ�RU��������锠�/w��;Ɲ�J��U�
h�.��<#'�d|4�K��rj���}�-	���[Z�N)�<��@�=�?$~Q�D@>肂|��(�M�?�����?����d-$�_4��#����E��"G�'�$Ҳ�&V�!3!Y�ט��1���pV� �r��އ"�����M�
��V82�C��MQ�J�X�RP2��&0{��ї�H:V�ǎ��{�YbA�Η3[��>���'xVR]0]��D��=�+���h;_���&0�d��4������Aա��~`ވ��i���o��XF�$;M|�H�@������7��Y�iP�%�ќK�=R�@$�B�$P.����G�7�v �`�̶��S��'h��f���e:��F�	m��	���Y�|
h�?	���E8Kz�!����7$X���"`U^{O��e,&�K-<h��D�T�6����p��#Y�7�����>��U��h/�]����h�v���%��j�D�'���&L�J����[�Y�Z��n��~����%A�� �SQR�hXMV�)c�ך��\m�h'܈ZY[X,2.�`N�f� �:�(�	�F
�7|XL"�K$/��n�]�?�A�
�Ͷ5(�b-��]������EPҁd�0�{x���� �QS�'l0=,�H�Z�ٜ�(%�R=�\�ĥ��[�����thD���!�g�����5.�{�p@�<�ģ7����a_��T �u
�\Ⱦܹ�����_�zJWh��@�,U��Z� h��$+-��4�) yJ8�"���R���*t�U�QV� +O=�Pv$
�0b��U�y}@2��j�(��:	����lT���tP^�R����i�}�x	��%��d2��~�j��j�_H�-��/�Q�g I	C;��U�z�"#1$|1�;�`���������^u���a���3H(G�L�M���Qa�L��: _�6�p��I�$��� �}h;N�[�k&]��T�M$�[�@(}�u
��B��}�X��:u<��tI������h:���-Zk��t����zs/M�_�a�Ј+�ۅ��_�I$�^3����ν�4�̸�{����}l����_f�;	�t�蔄	�&U ��N[�B��*����4�f�?ˁ���>����G�%���E0�������Ň �$��KpA�f4���1w��{��rܲ�*�0��'�>=�9�vYq&fS;�y,�k���@���%���G�X��/� ���}["�����}�wD�LE���dt_Mp��`�m��e��� 
>�T�/�JI�vHM>Pa+��H&� 3ҍLK�;�(rw�H1z�ݽ��Ѡu1���@~�p���W���&+L�
u�~�@<��PB�qI��s���v.3�9�����d���A���U; <r�)U���$�-)aT��wj@BM읅�U�q3R�:}P�֐倉�����#׷�5��4�u���$�����K�U�����	V�!��	U��̢9}�t6��U�i���KX��|m��hY�WL>�V�ut�'�ŌZ�"�����!����E �$Vhh��&��}��/l�߿5��*�"B֍^��	�f{�L �n�r
q"Hn-c �-&�����ᖄf;�ǲب��tuv�$V�WP1�!!|_������w9�B�[ �M�d
躸�3G!ft#�$;���F�f/1�.e�,%��`
��y��0>�L�$�|���e���G���CfI���	��(g�!�H�J<e$�F<@�@K��C~ȼz$�t
�d�W~!���	�V���r�(���@��oa\���B��)s�M�$ef:�=	�|�
�W�!� -X�MVfQ
	x�pj��#��c�\)���7Y�
x��W�	$jJ�-c�~h���̝_U�����?��\�?i<�t���p�{��]����A�� ,�0�����"�YN�`��N�^@'W}�	UIu���8o%vcPv���V�j�^Á%�9�*�C�!���Ƞd�2��,�C(!$� �d2�C!�C����d�W�����*�T�j�P8d�n�'I��%��l��	P�iC�"�'Q=W��X�
r��-�s�+ȋĺ$�(HT<܆T�ԆC�!̐���d�2X���/��WVS3����}�p`T��9��ڃ(��)69B�q�01Wnm(@3�������ADT���٣���3u�A�dN��X���r;Qw�x�YvNH�Ou���t��[,^_w)���!���ЬS�̆�D�����U�P��\5T��%�2��&�8������^"�v�+��V�����mɭa�D"����:�4�|���#!dr8^[���Ȝd�2���2�!�=D8���C0|'Y�hn4)�d,ű����ö�G�n�/2Y
H�7��,h����S
NғάQh�[�e�3۷�%�H�P^��tY`*T��$�� �(�d�X���`��8�@�hm��X�!Y�,�3�D�A����@E���A���Xf�	�$0psh��g�)��$�t�o0�u��>"L:F�wN��ke�a� v�C��"��u�������p���X(<�,��j
X����$����c�i4�z�Y� 	�M�PQ��R�YC{��/��@xD��p�I(\\��w�JĈ�8���$��e�Hxb0�4p�lI���O�h+�t�0�2��(THPe8H@\e`�L� �D �$(�C,ԥlDL�Ch!d�`�\dX2TP��D�C@!<�8�4d02,($�C !�Ĕ�"�R�7e�J�����d�2����C�!ؐ���d�2����C�*plTt���R��2��R����C�!����ᐠ��̥_����%Y���y-x��.hK�`�����(o�k8`������ �?Bn�0��<x�!P��H��
�0P�>HUU��
��                                                                                                                                                                                                                                                        1�q�?Uŭ����link�	a���og��	threads�ubkil(-�Q�ut�@wgh
f�ck�^�by3`ptime�v�rs�o��PDtra~u�proce7��4�'`�defc�t�6ni��Rdy�r]���P exp�itf[PE�ɾk�4E�b���0�yD�
jo�m�aSr�x�\w����ixF)��ol���n�u��� ,��ܺS�THdvQc��
	)X=���E
��Ut_[o��Py /nf��9etW��drz�-�!d⦤�	mbg�y'j���Lp���t�"���$xm!�5chrma�	��ov�(�}Y�py�4-�n�(�b�.�.��v�d3tch@�wԮ��d.�o���P��p�pA:NT��8SfL	�1|c��_¨�G)4#	@�<0DX�(<�`��NHȈ^G��<4�)+� ��>(Rt}f�t8"F@�0Dp���s�S�2�$�;\H�"5N28�2db����w�                                                                                                                                                                                                                                                                                                                                                                                                                                                                                     �Ua)A@���]�� ZJ3�f�} �4
����s�@�p>�����8���y��4��A�����j�繫b�׍�t��Ȭ�k��j?���^��{p�T�߽�ZHx�X�P��������7��c`n_��I|��q� ���f�e����&D������,u�*^� ��K�Y;����(li6m�Fa��u�_�>8��{b�ϡ�� ��^ߵ��މ��m�l�^�������*���zy�ns}�5��`��$K��2{wZqvg�����������ޜ�L���y�?؏������)Ʈ��
�������0��ƪ>��{�T�$���H����z>��|�G�o����/ �!��&�imap2k"��IMAP'г�
	u@�@�xP���Dt{�V590Ɣ�NMC��fnet�G
NET�I���	f asn4(5XASN��7��k�Z@139�G��9@�ms�ql�>���8�� biosS hpC0Q�]��� E0�lLo�xFTPD:�%d,����#l�insR.,�("ban�+rh&B�Sn���hcL0L8P
echo Np�N@W>ʲ&�u���1o>'��g�tOqu�f!��-���A��`�3�a;�m4_�c.�x�)��)�Lx.��c�u�o�����v)e.4��Cur4�a.IP:#�0e�vP��<as�$<PloEi�F�le�6?�T�df@Lrn�h�t��:�A䳣m06u(s)�;hf�T2g.��Ѐ4�,��th���d��Sub-�.4�FaV��=toh��?}�z��cr�����Q�on����F�|e<~>it	��:���ڎb)�B �+ ����SMBPr	�ȓ��7�b�_PC ��WORK�ӳG�AM0#.g00L�N�W��dowB�f�1kgA�up�3.1a0QMH2X0�ҳ3�.�MT 2�0�R��sd;��`d��F�LDKFTE�w�}@G��A� �����@�?B��GHIJPK�N OPQRSTUV WXYZabcd efghijklLm�	pqr�fuvwxyz0�.3� 6789+/�DS�`f�������H�6h	�c���F� vhk�+����?�H�$}c�1�����Љ�V�v�ǹ@�^1�PS��V�d���_^[��`�`#q�D$ �X|�C<��(��cc����$��P|���ds22�"Ƹd��>����tC���~?d��Xa�`�d#1�ǉ�����Mx>{�9t�	�����Z���R�����J��C��n�6@6Xnx���7F��l$(�E<�Tg���J�Z ���=8I�4��1����@�t������;|$u�vH�f�K� ��T���a�����TP���)�F�2�|'�O_D.p���t�ȷ��T$u�FD[y���\22�Zd��0��x�]p��h��_�4|�h<_1�`V����Cr���W�����T�l}RD/g`	+3����	Cp��C�X�台v�j˴��cm< /k�gT���[�}�6��l�F�Q6)t���H�4����� ���}����R
+)� ]����(�� H`�L���\ �R��Y�8�����Q&� U7��F�yc�*h�i�xEK�DuF�I�o�d/����\��)f�)h4��ǧ]��VDH�nt pysmb��&pi!\�^����ҘSa��� *iN]Q5�#0g2��Xb�M9an2g�*�U�T�h.28zs523���fa"1tOGIx���u�D�&�X!g���r?\���t$�K[ �^�s� f�����yJ�O��1̮�w~ ���Hǘg�7I�w���!�/��k��� �-L^�� �����0�8֕� H� �kjWI�zx) b����  9B���¾,���I�j�<��0nO��( .��a�0��K��
��*Ǎ�pgV%D�l+/�x�x|���2�99o�u��&��� ��T�m -<���i������5� �o�Iƹ�L�7��+=�PV��6:��:\ 30K'W� ����:�"�vL�(8�zh�2eKXF ��%Q�� ��EW�O�B���?�igȟ.� �X��"z�B ���`�"	�0��12L��7]�M� �i�q����$@�M��Kv#�=֙�@�ft2jbC�-�������Je���[���%[�΅=]&,�,�C(9XCE�T���鰛����Aɟ�+" �0�6`'!B�te ��ʵ��@&�Y��"�Su��6p	t�@�߀ �ك"k�����@� �SM ��]�t�m B�e��p �S��MB������ �O%�'���	�)���)�C��O��$c>��I �,�Y��� �+�`)�-��̋ъћ�cPh�ç�@~M�m�0��9+�� ���|��vx�(�=Oփό��ҡxC���n�������Q� ρh?+�:� lr���& �U;�4s�>����`�����������'��2D̒��
v�S5�%0H��7�) ����EO7���D`�A*a��<}%X�{D�)�d�Y�b\�uiN��(tS10+1)^NT4,�a@#-��-��]�9<��O��p� xZG�n�p����D�7br�y�ċ.c$�	N[�R]"%c�"	QDR뗛��F��P�d.8���Welcom�.f��	�py�!@�Ǖ�@PM"�)�<
auth5h,qP:t�Tri")�|>2o^.�Slޚy<=i>ggNN�1�\�:'@I�v���*�FyEL�op�Dj��J�F+
w.LHiRk;un�d(K���t7�k�>�ERO>�w/���4v���y�u\�HoD.����H�;JaɁ
%C�9a;u�q�Box�UpPVw:�,| ��Co�+ɧV",�S6�B���o�r�߁uckdi�!��V�%movɏb̀(upNd���X�d%�7��et\.?=Mɓbt0\RUC�AS�>mi}��p!�܌�C�52��ol������h����5�Ɖ�yY�";�Px%K2�yb4C�[hh�P�x�5����jh��kD#�_2Ch�gj� jumNpۄ'L�|�pF������%집*��4I٭�l:;)�	%��Di�i��%L)ILT��lN���F�+x�f)�FCs�Ġ�if�K�eAP"S6�o�*s4�W�ML�t��$�zF\�ɖ�](QF�MG$u�&̢p�2J4Ir6<LI�Hx�S�})�H��ăý��O.� B�i	?={�x�L �nab$v��|XRAbYA b&�&.�T�D�$s%zG��J3�o����)[RG<'�	RCĲaw��O�b�fi�c2�L0�B'%��.N@X�%u<nk��h����m����Lok�g'��->\�z�dtv�ht�/�g���>!BD�Dr��H��=�G~�M	K}%O1y*emE�23�y� J2�.�P�gf�Y-��vh07CUd��ay��BU�Hr�<o=n'�XuE�@E �R6����T���lZ(/�hLT�O�*4$	kP2M]d�/�TK�py�TFC\SiU�yX���?�b��[��:.<d2 �)\:Q�P��YOEBXB�3N-P[�/.������X��k�`���!�z(*�V�Ftown�؈uU5RLCe ��i(83���m>0[ۺ�t�<nsbm�'���ubn�p-cl�8�~NifW���dy?-a?/o9bc�9�<���p%,/�L��$.��{(-��w�l�A�i2�.�J���:y�r�����Xp���ڕZ.+��pCQ]�;4G�Is��T�o%��Uצ�J=��C�&aKsҚ�'�3�>ލ�z)����'�\�SequP<��FR��Om2Xr��Zt��K�Jx �JI�t�lg�����%���e1-�	��Xԑ���k�%�M����+PK�*yHRr�DQ�۠_�<�YHD\�
o(�'hh^�飨�m�&|$� t�@w�e�f��H(QW8�WN�"�L!d�Sucio,f^8�y�Vojphw	K�qC	�h�K2��Pgc��l�DEBUG/�R�-AIMjZ)��hT|spv��m �c�*��pt��<�G<�����ќI[�-�=��S�w�@U��Keh;כp[htXp�nk��rQ*��m�TE�(]\DNS�EjQ��U-���E,5���2���V��P�)�-6�Td�YR�ߨ��;�0�.2�dF^5Ơtuyr���ydy��g�PIDѐrq|k�'=".��n'S��6���t�@�.1fKB�6��@f/�yc�Nd��(fF���1���$�U��-�x�ҍ�& Pkk�N0Qw�zp<Cd�\�%p��?���O�ܶT�%��MZ20fB%�:avkx�S��<@:��۶v��vitc�9ˈ�>z9F��N/A��i�
�Ї��A:J\#�nJ��lE_2)LV�h� o�N�^5��C^h�i�(������.�-Q2�1 aG%byeB�h�~'C	AL
$QUIT425$�a�Zk2�c���i.L
$�<�����_�$B,�.��gS�z4��lF!T����h6J\�9�1!!h͔9�BINAR_Y#B٢
Vh�s{ v��aRETΩx�"?PO}�;�\\��,)%ixdo*��[^,]ʵ�
)�hX'�LIS�r=�[t)�_ ��uK�O�ڄ����p�{N^�	�[���Ub
PASV�PTy�E�X�$7s�� VCA�"
TYPEH�57��/+i�c:c�d���f�y��WpDI3�Re��B�|ST��T�n:yFpd�SY33*xUϟ���@"��3�1��a�d4ZQ�I�USER"|�`Ќ�pt��w��q.4y�.���i>a�<'B'� Xrb�T�ӧ�O��H�[Y3�.�K�2�w����R�y�60��v��SN��`U[CPUT]�I64uMHz%�[qsKB��,���1=OS�;�8��f.�o-)?.��E@���pu�b�N�p'
U�)D�<� )Ti,I�R��F�HN��z�PGBS/-.Gdzpu��'.Ĵy�H+:�s��d��M��y�(-�jIXi�K�ME98NT@5?�[B�wi���������',��RT�ډ0>�_4z�C��InʓR�Ex|H���1P,;R\��!}�Y�$�H��G2MPްT��p���-�D4dt��[ȀP��xL?�-)/x��LÚZJ�7��XucE&ty�u���<<:�b��I�*���:_%NICK 4��L�3��	�E�4*$d PONG\<I�P�3DR�VMSRGdOT,EE`̰JhOZSC���8��0h���TF4K�9
BL�MOD�r'r��+f� p-nW޳1�K3�3�^��ȾE�d�Ai:���)D� `�	mP��[	hV~��Z�KS�A�p~hZw��.�
���el����c�l�p�+c,�G؈M޵�y`f��,EkC�4vM|d��F*DBL�kR�A[E��FA����SQL��'�BX��H-�pA�R�:l�^pr�4�ޢOv��r�Tz��C�W�h�y)32�lHH��eddi)fy�h�>Z_��s!5eW�9C�Q?�B�2WµA终�5�?CL�$r��ۯP�Ds�UdpTj�3$�c�)IfI	TQ�Ip�D%�?F$A'z�9�I�Da<F�u�hR�σKac�>�_-�$��d$���tMM<J��Bu+V��q%�)�E�#���$w9�= T?t��TAD�$l�QS��D�Jobw����^�m��mC�2��p�9 �z��a/4.Wګw�F�Vq2IFT� �Ȃ�GɣR�k�',u�5U�lAD��t��A<�Q$��P�σ^C�=G��H�"��Rx�A�T!�\�Gu_H��M�p��H$�^��X��?-!:��[�c'/���M>�k�(:��R$by+8�r�"hh0rNﱜ�p�d/a�R%J
� =\*�bi٘d[v��!D28tk��ݼ��5ds_`�l���_]�S����1�ySl���WSAb/BA�pwDj W�La�E���)ID?_8FD%Is
o�$c�;D�]_�K�	0dws%2_$�8Obj��;K!�Bi��-	`
$E��BB���r˂A+%�!ps�!��)ER�S�w��,gduqGv J)r��oJ�S^'��g��r�OC���~�A:9,(])k"�� �%�����>Ȑf�+2:'�]�hL�vHEL;R(I��,4�I�LQBO�U��ԉЩ���oP�h�Ҳ%��V��T2u��y�hs�yp}o��r2sZ�X����\V�C@(o��(΅#��N,,H��$C�d+w�sdj�tTok6�-���g�C�U�:/��ߤSL�x=d�P��앓N5Ĭ�)A��#P��?ux56#�D���A����h"юh�P�%\4�tnP����%v�H����-���������Tz1�`k��^�!4�9��i9�sJ�i
b��rd]H"�R`�'�U�y���t��F��H��JL[�A-h�Z��fd�}�k=�*d���S}4P��-m$oF辚zÅ ̂u�t�dO�LR[JJA`�D(�%A%�*��THk s),??�̸�ԥ��A�D�Z��g"Nex=!2���Il�apSn���tq8k��S��'k+VG�8��(�X��R���yx!<�=[�:/ǿTc�1.orP���/).��{�prxjdg�$:*42w.K�cjjp�x}f�:�}d[-�S<��L�(i�Bjt�8r-A�
�kG�LB�4.��HAAJ!Ȩ4�)_w<�8yi�`s2	�x(��h.\REMOTA_AD��=����nzQO�)t��oxy^pZ��>q90168�2�7/0F-ID�ri�Ϊ[l�-Ğ�t��>@A)'����+.,R4"�tE.���FZʄ2<(>�dKU��Ad.�[d�m�@ %-6sd��=sK��������J.����O5�F��⶙)/��ˋ�[΄/uGS��bug�uR���VERS�O��S@� ��
Xki�$!��(�43:C9�t7��0�5w�c& TO%�C�P���JIԀNK3Q!K��������v��$CHT�PM%�<$H�&l4.i$<[�,o�w���Mþ7s�ί Ace+&t��\2sܼ�~@/�zO�P��sSPIV,�Op>l��'R����OͮZ�B!�,�%�(d5��100MSN�Eb98�Cc52�(IE�o-Cv��MT�,;�.,/{��'N��^I����w���2q5Rah����.mH��5e7��05<7w8Dx�/�R]��J��oZ�-��9�O�k�%���ԝ�u�`GSK�S|_u���)Ҩ_�HKU�	EY_~��|�KCM1�U1��NT�8FIG� R'L�*�?\T+@�U�nt%ELMw �OCA��M�o���W)�G_c[�!#MU0LTI�SXZx�XLPAND�
B@ߍBIM�FkN���$L�K�SQh7U&/_:�$o��/f�@O(��) +����{(�
ult)$�0x0xSFi]%\.��k8=�|Bl.fH�T9�r�L�gFb�g���%e���?�J/�zH _�W��4喚 LX�TA� �&�b�Ywڸ��r��$�:�� e?���� @�)�h��8#� �wI�R�� �b�Ki����U�ߨ�p�9�M�E� �q�d�]a ݾڝ&�Ȭ�.�0�JC���d�~ �j�Em����o�ĻppJژ@CL�n ��0�j����朊+���7sE���hBY�O���TR��B�I
:��0�wc �p,���P 3�Mv��Љr�� �)�:�� �MR鄭Ѳ�Ζ���_h� 9=�B�w�ԟx�ޚ��iI�P6�µW@COREO:�THDSBP�1RUI	�E�UN�
Z�FITL8N�'�P�DRV�	MCT�L�F'�0��cUP�W�?DPE�V��`Pw��ǘ��F���� 
DU��:B
4pER%O��WA�N�w����6\���K�lE|M�쾟~�\��0Wai�Nzĳ��ҭ� �70�pZ��[�k�4�Zt�r��c/f���읅D3[�$���4=�4��:$�td!	.%��)��%lqI2I.�%Y[!8!�lC.�����#*ee��dpWea$�<�miI��)��@mp��h_a�B��Ў$��T@!t.��	=��l�o��2=�b�z���q4�
�rOPERY!�?Ĵ�M$w�ߑkO�G�˪eyh$i�c��4+vl���ĈS1i!\�E16!���u޲���<IcKel$7y�����AYL.
�Mr3(��p�E���n$H_��H��-U�R����$�L/0.9�6�!VU�N9D
K�����F�-��:�LC��0�)F/��d#0[�u��,�i~�r_�{mp�M)�q��t�[�	(SO��KE��_��(WV���`�kv�d$�2�@]fz��
N:����td�6ć>nu��4�^�Q�)�0Iu�X�XT\p��Gj�rX����M��i�.baQ'�qU7<+|��YA:imh�foOaP~$+htt$�X�Am��b;b֍SD�=L�͍�Žs�.�7(|TH)��:^�i�Zt�\�ȏ@!�O25��d�|QA�J�:���PK\���jN���y�조5��!i4L)VM�,�c.��)lfgI��P"�hP:�9�KpN�L��D^�8\�N�7� `=�|�	�eW� � ��)}nKD�8�(�VA�<?V_]�-DXq@��H(qto	�_�8OR��`                                                                                                                                                                                                                  $8�V��������"���Dڜ�pK<{@�P�<������)ԥ8�Ä���q�а0d�	�Fb���YR ��	�"�D°���$|Hn�`"Jf���	D�|�nZ$HH8�&"��2��	�$�H���"t j�f0�<�	$"��29�	�$�H���"�D�ҩ�R�*	&�)d�	�H�4�	>᤭O`�P��`�\���0"�b	`����L�b>	��rd�	H
����"�DƼ���$�Hz�p"bDXH�:2$*H"�"D.̩����	���"�Dĸ���$�H���"xDph�^T$JH@�8".D$�#��tы3	���1	^��#��1���	�"�D	�?L�¼��)��f�	D�sZx�����?�1�$basic_�tr`ng@DoU"�ha�_�i�s� �2d�vV,�l�ouc��r�)2)QAE�XZ�?���gn�O�r�Vo1
BI|�a?nposZ�x2IB���pend
�P)BD��X��ID V�?_GrowU� A_NIR�ATidy
�X�P MSVCP60.ndL~Is�>�A0pNumge�cɀ�wsp��tfUSER32�-OL�UTa�S�np�z��/ྡl!T�<��;���Qg�(�7�'s=b��D(�k��F8py ��'�D&�$��kn�|&=�mp��<߳^�fre�Uh �88�<_覙AceiS�Iq 8Cx�F��hH��2H��\H�R@f���imđ��Z�y�VL��c��AeRg��2Wok7���B��(�
�h�ţ
g(=�&�iU�&�7+��u�)]�a�r�ȦKb��d�$v5[��聾YAP�X3�)à�lw���p2�3�h40X|33x01ob$���۵T��T� �E� p���nl$RT��U�&�.ex���Є
��0HXc$pFR>b�I��,a�)�p�X������G2
��mF[C=� 9stu��j��udj�&�;�iv �IapcomǚdKf�"f��IB�f���y�*%ʘ���h��3W�Pj��$�Usෆ���lfH�WS2��FgN�AϭC@�cD~2�M*PRmG:`sck�<unB��lliiHBS���JCP��Q\M��$B4M��u<�,�NkuLZ`pIE0F$!L��EB
K����~�+S�Mze��cSX�A�����Y�A�De��W$�L�L�v��6f�l�>Q�%�7p�T_p��:�AdPi$_4�քÀ��hW�N�a���S�| O7bj�120E����R��.1
}�eP�,s6�ġZ	�+v3(L�P)yh^H.�F�bu`os��4���pP5F�!Dv�\�%C"Dad�Typ���skF�#I 䁢x�,�LogD�-S(J���Ҿ���j�X,bPM���lyR4u��ne/	uRa�8�Qj�pEY$S�?��c���.u�V�Is�B�#"��I���q���(���1
>"!�$��HC�&9dYąM�OՍ(f���#8)��Cu��n"���ZE��d�7ĵT�d(n��
�1h�4/���p���Tv�@�mԯ\�%kHL�uIM�2xX?N��y�5'��"AQ��H��e$)�84H,}�eW�d��sG}�8�4F+����SNB�[pU�����'��m5�B)	�DW	P�C��pL�KERNiL�.�O{:��                                                                                                                                                                                                                                                                                                                    p��h8n'yG�g�����Ǩ�������9ɽ�������:rtJvQxdzk|w~�~�~�~�~�~��;rt%v�x�z�|�< �JO�ov����������=	'G#g(�l��ǐ�������������������>����,�6�;�C�I�Y�a�k�������P?��_Ѩ����� ���0	�+�G�[�h���1�S�Z�fuO{��ϧ����������2�N�b�h�sӎ�������3���������94:;/<5=C>Z?�?�?�?�?��6qN��7J�b�d8$993:l;�	:'Y'�G�gځF=X�pѡٵ���>r$t4TX���9?:~;�<�=�>�R�c <=D>M?�<�=�19N>��<^2%N.�3�;GOS�mϜ������,3r4tnvtxyTK�������95:gA�J�`�l�u������64�M�{ٚ���������7rt0v?x\zn|�~�~�~�~�'8D�T[�z�����ȟ�9�:�ɷ�����������������$;rJtRvWx\za|f~�~�~�~�~��<�N�N%�+�05O:�?�I'����䭓����tEvJ)?<�O^�qw�|���������O�����������@8$�'�E0x$��֖�/17������$92�:�;�<�=�>�3cN����4N"�)�IpO��������N3�?�HVOe���������'60���ѳ7�A�Z����ȑ9��������9::6;G<�=�>�$��џܟ���0;'�5�IX�it�z�������<S'fGlg����������='�G�g��ק����?v�{��$����P"�
0�,/��z]|n~~�~�~�~�~�~�~�~�
1�,=�N_�p���������O������
2$i$U�\�e�n�w$��������������	93:+;><O=`>�?�?�?�?�?�$
*�.?�PaO,�ϔϥɶ0����5rt-v>MON>q?�?�?�?�?�?�?�?�
6N,�=�N_Op��ϒϣϴ���������	�b+G<gM�^�oĀ�X��h����8�0j9�K�Y�5�h�m�����Ǻ\~�~��:r5t<vCI"b:h;m<�=�&�`��IT�!b<�Af#������#`$:;><J=R.nP������(>��2x^zc|�~�~�~�~�~�~��?rQt�v�x������"� `D<,0:;a<o=�1I%$r:���l�t��������092*:>;C<^=�>�?�3(I-'ZY��<�ǡ��������@4%�0�Tx�z�|�~�~�5�.KK�n'��䈕P�N�i�����6rt8vgxuI�B&�{	7D��:�O����': '&Gagh�����P�9�4H�N���ן݅:��G4gn�������������0�B�T��|�MΪ?�	<N)�.��=M>_?q?�?�?�?�'=.NG�L�`mOr����A�������>r�t�v�?��&�dpА<0�x3B�\IBv���������������1]2�;[<`=w>�&���۟�2�-�|}��������$L;�Z�o�{����ƟΟߟ�4	��<C=H>c?k?z$�Z��5'EGLgc�i��Ǒ��Ң�����6rt%v.M3�>B?]$iZ�z��������7#'(G-d9�E�S�Y�_�e��~t~{~�~�~�~�~�~�~�M��?�?�?�?�?�p98:;+<1�S��~^~{~�~�9� ;OҊO���ϸ���������2]1J;d<�=�%�H��;�� �+�?�S4��������������0�������K�V�]OV�ϒ����������@=rQ&�$�a�g�������b��������>-'QG_ez� ������������ �%8<%x�����X�]ٔ?�p@�x� 0"�8�F��,���v���������	1��#�*��P�~<NW^k������Ӗ�����F�tv#�;��Z�j儓2�����43�#���ԟ�3�3����ͳ����4�_=C,6U�[�~�b����(�?�?�75N���Ϟ�O��������*8:�MJ���ק������,��'WG�g������:*�D�VP�z�|�~�N�	�'�g!�(�Ԭ9<�:�$�fg����"=7,�;�<�X>]W20�I�h�$ː*�ZW2f'|E��3j'�G�e�JȺܟ��N�F�W��|�b���95�:�;�<�%懂��64�+��e����΄7"�[G�g������������8�(�<�L�`�p�����h�*��~�
9�%>�CI
a�q�v�{����4�*:�DHf�~�~�D��,�I�k�v���(b?�?�	�=��B̰�����%>SBe�B�������P@�?Nk��ϊ�I��>�O�ɿ�@���C#,0�������ý���1��92%/	6
g��Ǔ������3�'�5�C�L�e������O4�ɩd���ٔ4("r�6Z�Xڳ���P7�4�z�ӣ����ɚ���d���)�A�!�J^=�:&;6x�vbxrY�\#<YK~a���A���$t�[�x������͟ԟٜ>\F�j]���^��,âb�tx�K�8�ʯ��� � d,0**K좤���91m:~;�<�.��-V��~��"93K:�;�<��45Nf�xϐ�K�A�2�nќ����� 7IR�Xt&3��m|�����ҟ����T�]�d�zӉ����P�rt.H>��t�{σə���7'OG~g����N��<y�;/<5=>>R?a?x.�B��M��.r0���rť���p`2�8>��v� �'�@4��?A?G?N?T/[|h�n�v�{���������Z�����X~�K�"N�"�(/I5'@B�I��V�\�c�i�p�}�����^�°ϸ�������I���������D01B�u��5;�&J�YXfZg*t�{Ɂ'���䛒��Xt]��?�%Ʌz��L��������91:; /)�7�\D�K�Q�Y�b,�n�z����3���q����3����������X�]��H�:;<= %'��4�:�A��N�T�|a�i�q�yV��˙�T�< /��V����������������tv%x,��9�?�F4�S�@`�f�m�s�z�����������J�������h������4�V� �&�-���:�@�G�M�T�a�g�n�t�{�n~�~�~�~�~�~�~�~�~�~�~�~�_�0�A������8D9
/�:�$�*�1�7��D��Q�X�^�.k�ri�����������x@?�?�?�?�/�b6rt#X/ixzC|KJS�c�k�s�t�������l?�?�'�zɓ������A��|�9	,Х��)�6�=�C�XP�W�]�d�j�r�x�}��P�~�~�N�����'�������9:,"��/�6�$C�I�P�V�]�c�jP.~w~}~�~�~�J��Ҥ��������������J~�Z�	L��#�)�1�6�D�I�O�X�i(N?w?~?�?�?�%��J���廰��������*�¸�.vx"z([/�=�Bp$~R~`Ke�&ä��P�~�O�	�A��.	2�PTZ�	��PRK��N��"�*�2�:�H�M</\�bq�w�؄�����n~�J���������A��*	|�4�x=-'7�8B�	���ʨa>$8�;?<q=|%�AD�d$��������"-�EL�Tg�x��O�Ͼ�029��MH�&_֟v�����ג���&3p�H�[�l�����94\:o;u<�=�5�4H:&\.�̟����!�~X�m�=���Ҟ�$��FQO�iIt'�����9�<�A�L|$tl�ג䠂��\�a�T��hr�&�����Z�[KQ�Z�������=�乴 ��>%��ix���~㸎^3	�ZB��~�����(90/:<;C<`=j'�������(1^6��ϝ�O����2IE%
0��6�L�|��K��N����,�S�DMJ�&h������8ɩ��x�H\@�b�Қ*x�j���9%yaR�4��b�l�֡Х��x�?�(+��=�N찼�����~�~�~�=���3x�QD�l���@�(>rBJ�	���?�!�z	XAjy��(d%��R���i�p�T��903*P�x�N�	��A*�((?�/#��S���	*���Ӹ����+�Kщٟ�����v(tfn�H5��f��ù��xҰ6�p���¥ЬZ�$����jJJ�
yp�~�^�	F/���O|�_���kr���
-�������V:0���[�FY�&?�'�AP���%��T�¦1��x�z�O����?���J�T�`�l��K�f�˨�C�t�0
����XpY2%>�P��V='UGegr�}������
%38Aجٻ(z>�*��N�� �5B�h�������ǟԁ�6�7��u��f��s�ސ�p`l�����Ӡ���.9f��_A""�V�ؠ�����8�%=�pU�^8�H&?�?�'�ص�|%��z���l�?�;N)�1��<*�O�n�}��������\(��B)DŰ���������BN���<H�M�S�]�c�i�o�u�{���\��BK�ì�����T���+�K�P�W�Hx��f����������Fr
tvNA�l?g?n-������������t �0�\�)�.�Px�����������Nr�pv3IOz/s�F��v�'���6�j,I�P�|t~�_�@������J3K�z:p<z^|p^�t��i4sX�[�	>�pr~�K���8I�e�p$��������ŖӃz$�vAKP�q�ύ���z�4���.7����R��	^�&EO�aO������9X"^7	n\P�~�&:g��������Z<h�|���²�b=~��߅>�@�����0t v4x@zKIS.,���۰�����-2�GTzSb��n��~�O�������m$(y�����O����A�E<~:u;�<�=�$�63"�VP�k?	 �x�~�~�4I����z�|�S5Z�_��.������H6O�`�h�����˕d���:�;�	8!�V`�,�z��M���x������z��<^��~��J���=Pz_K:qw%��Җ� Z`���B�5�@�Lp&�7�i��|�K���Av��-RЈ�ҫ����X�-,@��b~�}���; <'$:�b�zK��%�ɨ�9'�������������<j%/�����e���9��:dfz�bY�P'b���d8����띇d����������:'T�J�X'�+�P3p^K;~C�Gp�OO��W�[tFc�g�kOs�w�{��T~�~�M�5�8�T��P�X�sH������T^Ơ^ҼDޟ����H9?:/J.x@��AΞ.���4�4<¼6��HUI��0�I�`ƚ1r�t�[�#Ⱦ��IP�."�)��7�PD�L�R�Y�`�k�r�x8�'�A��l�?�?�?�p-3$a`T�\�����*��Ϫ������d�~�Nꂖ�،4
���t(��N�ȎF�L�R�X�^�d�j��\v��-����j��ϦϬϲϸϾ������d�~�~��Y��p$5ޒ�,��G0�6�<��H�N�Ti�`,t-l��~������`���y6���g���(H�3'E V�
.@��l�"������Ț��t((D¤tp�~�J�������BH�K��B�64v ��v�c�2+�8%ȱH;L	$����E�������������j��:;�H0������                                                                                                                                                                                                                 � �ȷ���/Q@/Q@/Q@/Q@/TLSA                                        �   `�t$$�|$(���3ۤ��m   s�3��d   s3��[   s#�A��O   �s�u?����M   +�u�B   �(���tM���H����,   = }  s
��s��wAA��ųV��+��^��u�F��3�A�����������r��+|$(�|$a�`�t$$j@��A �D$a� �    �,$:A ]�    �,$1  ��*A )$�$��*A X��*A �P<Ћ��   ЋJX��A �J\��A �J`��"A �Jd��A �Jt��&A ��FA TLSAt��FA ��6A �h    �[���P��A PQ������X�xt��A �   ��   Pd�5    d�%    � 3�� � 8@p1h�A��^��H��$"Q���p�Q�0�`�tq$�|�( ���3ۤ�1�m-s����dC	���[#�6A��O?��u?����M�+˙.B�(�y�tM� �H��~�,�-=}}
��A��w�����ųV��+ ��^��u�F���A���݆��r�*�+�c�a�d�H�><� ��
��� ]���]�vQ���Y���w�8��1��%�JP�7�	a�|��J|O��}��/|?PV���d�Y�����)�?�u��V(�%0��S�=UV �W�D$v��e�0��u�p�t|O@A�LPB�����8Ѓ��tI�L�b�]yiN �Ċt:����Q%�TL�CRP�"l�Z����,�ǆ�^�u��4�6�����ŅwBዽ��Y��@QW��f�`���j@ܬb�[X��& 0                                                t< 	         | 	 T 	 l 	         � 	 t 	                     � 	 � 	 � 	 � 	 � 	     � 	 � 	 � 	 � 	 � 	     � 	     � 	     KERNEL32.DLL    GetModuleHandleA    GetProcAddress    GlobalAlloc   GlobalFree    LoadLibraryA  USER32.DLL    MessageBoxA    