MZ�       ��  �       @                                   �   � �	�!�L�!This program cannot be run in DOS mode.
$       C��S�� �� �� �� �� ��� �� ��� �� ��� �� Rich��                         PE  L             �                  �    @                    [<    �p                               \p  P                                                                                                                   .text  G                          `code ] ;M       F                    `.rdata  c   p      X              @  @.data  [�   �   �   ^              @  �                                                                                                                                                                                                                                                                                                                                                                                                                        h����R��#ɉBZ#�$�����$����X3�W+|$�|$�_ ��!   h����V��|$��!N	N^3�Y��    �� f��2���
��   �Uj�R���    #�!rZWSR�+T$�Z3�R�������ҁ��r�����Z���r�d�@0�@��|����|���p�� ;���ph�w�P�ą�!H	HX+�I����΅Ǆ�$����+�YPh�����$����D$Ɂ�����S�#�$������#C�� ;׋��    8l$���   �3D$�+Ɓ�����S3�$������#C#������ ��   h  @ 3l$ف�����Q�+L$���#i8L$�	�� �����Q�̇�	��h�ׁ�����S#�$������#S#���$��������    ��3�Z3��� �^   Vhr^3����q��4E�*R#�$����ҋ�#r��r�#���j�W��;��!w_hr^3�R#T$��ԋr��    ����l$��P�ć� ��h����Y+���	+�3�V4$���3Nہ�    �6�    #���������[<h�c�W����!G	G_�$����X�Cj P��#�1HXh.���Y�YQh.���Y+�Y�V+�$����^��j W���� �W#T$�ՋW_h����Z�ZQ�̇1�	��h����^+���������Q+�$����#L$���qp �	�|$�1N��   ��(�   ��m�[h�u?�P�ā�    !H	HXhiz�
#�$����3�$����L$�+́�����AV��3N8�$������    �6�π� ��   �   8vw�MPINo|Z�hh   $$3�#L$�+�$����������V�$������#N�� �6���   ��iz�
h�jzih
���P��;މpXj V��8�$�����D$�	^^3\$�[�  S3�[j@h 0  Sj Q���    �A��?��F�$�����AY#D$�Xj �Ћ�h[E�QW���� ��G_V�݁�	���Wh	���_�_[<��}E��h}E����+4$#�#ۃ��C��   �"�p�n��h   $$�    ��V�$������]F�1^��(j Q���    1QYT$�#T$�Z�sV+�$����3�$����^�R�$����#�$����Z�K��$����+�Q#�$����+�$������3q�d$�ҋ	;�����S+ہ� @���    �   qV�ĭ�s0�.��3ہ�    Q�$����ϋ�3Y�� �	y Ƀ�h @�;�+$�ހ� ��   [<Wh�3�_3�_R3ҁʷ3��   f�T��C��>��J��13�V��m�ы�V�� �6���CS\$�[�j Q���   ��R# ٞ�Qց�L[���QY�$����+T$�Z��j�S��z ;�!C[j ��IX<d�$����XH����_�    ��    3�Xh ��W���;ǉO_h��_L$���������P3D$�+�$������3HۅƋ ;��Ӂ�   3�Y��(��(�   �k�a�Gt����^?Uj��(j P��;�	xX#|$�_�[h�p�R���   �K(Ah   $$��    �JZ+�Yh�jziV#���  jhl�ؿQ��;��YYhys�P[3�3\$�+�R+T$�3Ջ�#Z�L$�Z��� ��W������GO��ys�P�3�_h 0  j R�Ԁ� #��Z+܋ZZ�   *�h   $$j h���#��   ����������=2h   $$+$��    ��������Ћ�h,�"~Q�́�    ;��AYj P�Ā� #�1pX��RT$�#$Z[<j P�Ā� 8t$�1pX3�$����^�Ch`3i ����    +<$;��   ��`3i �V+�^����(WhE��_+�_��E�︃�(�   �C��>��h   $$��(�sj P���    ��    1pXt$��^�S#\$�[�KVhxm�^3�#�$�����$����S3ߋ�#s�� s���8vw�MPI�� ��Shxm�[3�W�$����#�$�������_#���$����_�?���3�t$�W���m(���)+Ћ�#w#�w�?;����    �� h�<  3��$����+�Q#�$������y#���	��    ۃ�j Q�̀� �   67���	/<�K(A�'�	AYD$�X�D$h@{���    ��    +$#���   Wh@{��_�3�$����+�$����������PD$���#x��    � ��$����z-3��   ��U��SVWh����W����    ���__��2��+�[�]��h�mΑR��ɉrZ�$����^[<j P���	xX�$����#�$����_�[x�S������C����+;��	   � 9~�,���h   $$�#�$����+�$����+�P3Ë�3Xɋ ������+�{ j V���    	N^L$�Y�W��c���_3����S!�Sh�S!�3�+\$ԁ�    Vt$�t$���^;��� �6�� ���\$�+�P���X� ��#Xv #�X� ��$������^�����h>h�Q��t �މQYT$��1���Z�3�hm�9R��#�ۉZZ��$����[��Q�$����Y2�   Ƈ��RBj W����	__������CK���t���� ;�+�#\$���1j��������Q+L$���Pd���3Y#���	�� ��W������G���t��#���$������������Q3L$؋�y��    �� �	����: �U���S+�+�[;E�S   j R��ۄ�$�����r+�$����#t$rZ4$^F;s�����j�Q��;��	   Uj[��67�!AY�$����#D$�X�S$j�W���� !W_h��3T$��$����3�W|$�#�$������3W;ы?#���+�+T$�PD$ʋ�#P�� P� #ۃ�����х��r�Cj S�܁�    �s#�$�����s[h�V^+�^j S���    �S#�$�����S[�3Һ�V#��Z�Q�$����#L$�Y��j�P��;�#�!xX+�_�S3\$�܋{���� ���^R�$�����ԋZ��    �   �qV�ĭ�s0�.�h   $$���Vh:?sP+ċċp��;�� ��   �^��:?s��                                                                                                                                                                                          j�P�Ā� !xXh�C����+$�#���   S޻�C��;��    �[`h   �$+�Xj Q����Q#T$�+ЋQY+�$����T$�Z��Þb�h��b�h=P[f�   �� pz �   j S��;�1K[L$�Yø   S�$����[�hZr�+S���    �S[h|���Z3�+�Q#�$������#Q�#�Q�	�� �� ��   j V��;ǇV��~/�3�$�����V^��    ��|�����D$�%�>3�Z=P[fj�R��#��|$��}I�!BZ��nX#D$�+�S�$����+\$���3C} ���$�����r�A��   j R�Ԁ� 1rZ3���	�\w �W���'b��w�   �@y�?��j S���   ��"�p�n��z+��{�$����#�$�����{[h	�\_+��$����3|$�������S3݋�#{�D$�=:���΃���   Wh���_�_Sh���+�\$�R3T$Ƌ�#Z�Z���   ���qh   $$��   +ˁ��c�\$�������Q+ʋ�#Y�l$��	�   �\eh   $$��    ��   �� pz �r   ��j   R3�+T$�Z��Z   h�fQ�� !y	yY��Ն}j_3�j�Q�̀� �� !qYhx��v��S���3�$����S\$��܋s;������� �^��x��vj h��ZV�   ��>��J��1��m�3�i�h   $$��,  h��G���$����Ɓ�    +$��    �   ٞ��   Sh��G�3�3�$����������Q�$������#Y�ߋ	�|$�|��   ��$����+�R+Ћ�3Z�    �#ҁ�   �Ћ�h�.�P�ąǅ�!x	xX+�_��j S��-f-^�$����[hbg��VS\$�[�B,  ��ha�|vP��9T$�!p	pX+�$����^���   j P��;ف�    �X3�$����3�$�����XXh�;B\$�j �+�$����j �����+�[P3D$�+�$������3X�L$��� � �� ��   W���_;� �?�|$�.�L;ǃ�+�[���;B@<f;xH�5   ���e���e��   j Q�̀� �A�$�����$�����AYD$�X�h���Kj S��w { 1s[W���֮��$����_�-+  �؁�d��j�Q���   �����h   $$v !yYj |$��$����+|$��$����Q��~�Pk��#y;�y�	��$������� ��   ��d��;���ǁ���7$|$ށ�����R+�$����+�$������#z��������c`޿���ۅσ��8���   �   ��$�BS�����E�˨�f�T�@���C��j P�ą��    �X+�$����؋XXhC��#\$�+�+ځ�    P��������q��3X;�| � ;Ӂ�   �	   ٞL���83��$����������Q3�$������#Y��	��$����|���3   Xj R����� 1ZZ��$����[���[��;ǋP���.|D$�XCV�$�����$����^��h2�G�Sh�SF[+�+��$����j \$��$����\$�3�P#�$�����$������Xۋ �} ��W+|$ߋ�_�#ҋ?�K(A��   ���SFhp� +Vh�8o"P��x �߉pX�^��(  �Ёǖ��h��罅�+<$��    ��   ���   W#|$�3�_h,��hF��R�ԅ��!r	rZW+�$����_�(  Vt$�^��h����R��| #��JZ3�$����Y���T   h�4�W����    �   �=2� 9~�,���h   $$�__��q^�[3�Q3�Y�   R3ҁ��ٿ;�3�Z���ٿ3�aQ+�Yh��S+�$����[h���W+�$�����$����_hL��h��*h�	<�P�Ā� ɉXX������+�[hp  ���/��j P�ą�#�1PXҺ�/��u 3��$����+T$�V+�$������#Vr #�V�6����Ƈ��R# ٞL�	�8vw�M��|$WR+�$����3T$�Z�0  h�I�+D$�W|$�����G��    �?��   P�	   �u
{���WD3�Vt$�^�=PR3�+T$�Zh~mj W����    �D$��4�G+D$֋G_3D$�X+�j�S�܀� ��!K[3ρ��ƀYGE�Ph<[�4W���� �   �'�}r�@!W	W_h��8#T$�j 3�$����W+�$����+����W��?��P3Ƌ�P�ǋ ��    �n��z+�!F4]ң�Y��   +�3�3T$���    W+���3W�   ��d͂�����������|$�=�?�� ��j P��#ہ�    1XXh��83�$����3�P3D$�+ċ�X�р� � ��   e��   �[h�  R�$����Z�D$PWhc���Sދ܋{��� ���   ρ��P��+�S$+\$���{�    �#���   P3���c�����$����Ty +�X��.  h�jziVVh��m������]+�R׋�3r#ҁ�    �t ���R#T$��ԋr8|$��    ���   h��m��� +$#��   ���8vw�MPINo��   ��$  jShZ�"�[3�[j Q�́�    �   u
{�y3��yYhZ�"�_3�+�$�����R3T$���#z�|$����z����D$�ȃ�h 0  �   a�Gt��h   j j Q��p 	AY�X�Ћ�W#�$����_h�jzij Q���D$�	�KW���q�$����+�qYV����[�^�@$  jV3t$�^h 0  �þ��h�X��W����    ;�!G	G_�������ЁȾ���+�Xh ( hJ!iV��9t$�!^	^^�$����\$�[j ;��Ћ�Q�$����Y�D$W+�_�$T$h��dV��;�!~	~^h*ϵ����4#�$����j 3�$����3|$�3�V+����#~z �    ~�6;�;���   Q3L$��$������3y��,���qV�ĭ�s0�.�\e#��	�   ���c`޿����xQ��$8�$�������_h*ϵ�+4$#Ɂ�    ��   `Wh�GʹR���D$��y��� !B	BZSj R��;�	ZZ��iV��[���#�a����Ƈ��R# ٞL���8vh_p5:Vh	��P���    ;�!H	HXL$�3L$�Y�"  V���6��#T$�+�$����Zh �  Q3L$�Yj Wj R���	   �)�O��kh   $$1ZZh���G[3�3�$����������W���P$f��#_�q �?�� ۃ����G��h_p5:V���	/<�K(A���$����}��!  �|$S�܇���L$��$����Yh �  j h5C9QP�ą�#�!x	xXR����sZ��Sj P��;χx+|$��xXhnNX�+�+�R+T$ڋ�z�   ��Y��*����h   $$�׋x �����_j W���#�1G_j +�$����X��nNX��� +��$����j �$����D$�#�$����3�3�Q�$������s��$��3A;�#ҋ	�    ���Q#�$������A�� �	�� ���$P�   c`޿����xQj��$c쁁�$c�h   U�ï��j P���    u �P�$�����PX3ҁ���;�+�+�3ҁ�����P3�ŋ�#P;� �Ѐ� ��   hZoީV��3Լ�j P�ą�1XXh3Լ�܁�����R���f+�$������#Z;�#ҋ��#Ƀ��[�&   ��S�܇���3�$�����$����Y��V���+Ɂ�   P�ć� ��3�3�Y�^j V��;�1^^;��$R�ԇ����	   �����_�ujV���6��3�#D$�Xh   Uj V��;с�    �F��G��$�����F^�������Ё��k����    ��$����tZ��Xj Q�̀� ��    	YY3ہ��k��#��   �h   $$+��	��7Q3�$����#�$������#Y�   K(A�'�}r�@y�Y�	�D$�5j���   hZoީVS3\$�[��  �� �� ��h�[V��8T$��    !^	^^+�#�$����[��S��j�W���\$��|$�'D�!W_3�#�$����Z[<�����Wh���3�������GQ����8+�$������y��8t$�	��$������   �_�[P�Á�����A��   j�S��;��!C[h2r�x�$����X�� #�3�X��2r�xI��   �.�\e:�H����c��Q#�$����Y#���WhQE�`_�3|$�|$���������S#�$������3{�˨�f�T��C��>��J��;�#ہ�   ShQE�`\$�+�[��    +�[��   SR3�$����Z�$P�ª��P������@H����#��   PINoh   $$+��$����D$Ɓ�����V#t$�+t$���#F�׋6��    ��jS�Ł��L Sh�L [3�[   PW|$�+�_hZoީj�W����    �   �!w_j S��#�;�1C[h�ؖ�X+�3�$����������@QL$���3A;�;ʋ	�   (A�'�h   $$��    ��   j W��#�#�	G_h�ؖ��$����������R+�$������#B�ً#����X�i  ��z+�!F��j�W��;�!W_����ͻZ���ˋ�h���pP�Ā� !H	HXh�6T(Y�P3�$����#�$�����ċHp 9�$����� ��   j V��;˃�$����~	~^h�6T(_+�3�j 3�|$�������P+�$����+D$���#x�;ʋ #Ɂ�   V�$����#�$������3~��$������$�����6�� ��   ��   ��#�3����t'V+����t'�   $�BS�����E�˨�f�T��h   $$��    3�^�QL$̋̋Y��    ��$�����	����Vj +��^N����r 3�R#T$�3׋ԋr#���$����#n�ы��   ����R<Q#L$�L�5��w�MPINo|��    �YQhL�5��P3�$����D$��#H�� ��    H� ��    ��   +�V+t$�3���N#��6��   �Jj S�܁�    ��Gt����^?Uj1S[3�Z�BW#|$�3�_�Q3�$����Y��V���mPh�mR#T$�+T$݋ԋBۋ��   3�S�$�����܋C��    ��    ����_  QR3�Z�Jj P��#�1xXhnOcW+�$����|$�������V+�$������#~} �6���3�3|$�Vt$����#~��~�6;Ѕ���h���%Q����������=2� 9~��   ��qV�ĭ�s0�.h   $$�yYhnOcW_3�+|$�V3�$������#~�   ���c`޿���ۀ� ~�6�߁�   �rhS�4W��;��    !W	W_3�$����Z���˨�f�T��C��>�z��K�Sh�K��+ށ�    V�$��������jӋ�3^�� �ʋ6��Ɂ�   3�[��YS#\$�\$�[��(Q+L$�YI������^S+\$���IkP[h_p5:Vj V���#�1^^��g�oh��ڌ[�a  ���!�j P��;�1xXh�!�_3�#�$������������S��-��{��3{���    ��	   ��k�a�Gth   $$������   h �  j SS����ܘ3�[��P�ć0� ��U��R�ԇ2���#�$����#�$����^@<���   V+�^�  +�#D$ɸ   j�V��#�!V^�Z��o   P���_L/W3����_L/�� �3�Q�$�����$�����̋y�   �z+�!F4]ң��	��h  @ j�W����    �!o_Q�̇�	��#T$�3T$�Z�X
  �݁��Hj W���� �    1G_+D$Ը�H�� +�3�$����������S�$����ދ�#C��    #ۋ�D$���[<Q3�I�᭡�9�� +�+$+�R3֋�J��    ;Ћ�	   �c`޿�Ձ�    ��Q+�$��������9��    �Y�KS3\$�#\$�[�CQ�$����Y؃�Q�̇1�	���   C��>��  QV34$^3����m�3�i�%����{$��    ��   j R�ԄD$��1JZ+�$����+�$�������o���+�Yj P��t �HL$�3�$�����HXh��o�Y�+�+L$ف�����ART$�+֋�J~ ���    �   _�u
{���WD-b�)�O��h   $$����ha�W�P��y !p	pX3t$�^��   @�6   ��Sh�e�[�W#|$�3����_�l$��?��   h�e��+$Ɂ�   ��   ��0   Wh(�-�_�_��(�-�����i�h�i��y +$;��    �����*   h   �$����_V+t$�^�  j�R��#�!zZ#|$�3�_���E   ��    ��    j V���D$��    1~^�|$�_��  h��5R��ɀ� !J	JZ3L$�Y����   �@   Pj D$�#D$��$����+�R3�T$��3B��;��9t$��    ��   H����ٰ�� �    3؁�sWa8#D$Ɂ�����Q#L$���#A;ы	�   :�H����c`޿�h   $$��Wh��ٰ����MS+ߋ�#{�� {����	E�˨�f�T���   3�3�$����+�3�P���3x�� ��    � �    ��   �   ����   3���   S�$�����$����[�   h.��R����!Z	ZZh��n�3\$�������V�3t$���#^���    �6��    #҃�3��$����\$с�    V#t$���3^#ɀ� �6�INo|Z�h�&g�����_������nԃ��   3���   SV3�$�����^�$j�W���� !G_WV�#t$�^�s�Cj P��#��   Uj[��67h   $$�H+L$�HXh��L$�V�$������#Nv ��    N�6�ǁ�   �R�$�����ԋJ�� #����   j W���#�	G_h��+D$�+D$�RӋ�#B�   nh   $$w B���    �   !F4]ң�Y��*����d�h   $$��+�X�hΝ�mW���� !G	G_����hZoީh��?^R���   2� 9~�,���qV�    !r	rZR+ҁ�s6�<҅��Z��s6�<�k  j�Q�̀� ����!yY+�|$�_�Ё�$��h��9PP���t !X	XX+ہ�$���   f�T��C��>��Jh   $$+�PD$��ċX��    � ��   ����3.Ih3.I��+$�    ���   ��(3L$������AV�$����+t$���N;�;ً6�� ;с�   �� I�   8vw�MPINh   $$��B���3��R+ԋ�#r�&g�����_�r��#���   S\$�[d�0   h)U���+<$�    ��   W����?��h)U��3T$��$����j �#T$�PD$���#P����    P� ��    ��   S3\$��$������Sy ���#Ɂ�   �Z�@�xj P����ʇx�$�����xXS#\$�\$�[;o��   j P�Ą�$����;ƇX�$�����XX�[���	   �n��z+�!h�  h҄��S��;�!s	s[��    ��4iހ� �W+�$������*�_z���w#��?��   ��4i�,$j R���    	JZ+L$��$����Y�Gj P��t ��$����1HX�+�Y�G��   P�X�?S�܇��Á���8�X9<$����h�"��Q�̀� y !A	AY3�H��qDIр� �3��$����������Q�3̋�#A��;��	} ��   S������CK��qDIс�    ��$����x+�+�#�$����j �$�����$����W3�$����3|$̋��_��    �?��   Q3�L$���Y�    �	�T��C��>��J��1��   h_p5:j R��s 1rZj R���    �Z#�$�����ZZ#\$�[��  �Ё�]Sh���][�\$�݁�������Q#L$��3Y�ȋ	��    ���L$��;��D$�I��[�$����S���09��#{��    {��|$�g����   ^]j�W���   ���WD-b�)�!G_D$�Xh �  �ú�c�Ph��c�S+�$����+\$�܋C�؅����   +�ā��U+D������S\$�+ۋ�#C�Ƌ��#҃�j Q�K(A�'�  PQL$�Y��hl�Q��q #�!i	iY��SVPD$�3�X`h+/��Q�̅։AYh����3�$����+ā�    Q3͋�3A;��	p ��   +��$������    W+���G��    ҋ?Ɂ�   j W���� 	G_h����X�X�U�Ej V��;ˇV3�T$��V^T$�T$�Z+��N  ��    +ہ��R�Q��    I���R�;ʁ�    +�3�$����������R��$������#J�� ���    ��   ������c`޿�ՋuW����?��3�[uh��g}#�;�+$�� ��j Q���T��1AY�$����3Ƹ��g}�   ��X�> ��  j�P��9D$�!pX���[��^�N��    ��h��T�P�Ā� t �XX�+�[��ȋ>��#(v��#(v}W+�$����_��S#\$�[f�j P�ą�	HXh��Y�3�$����3�$����3�R+�+T$���J�    �ϋy ��$����u�����������D-b�)�O��k�a�Gt����  j�P���!XXh?�o[3�#�$����������P���� L3�$������#X��    �� � ���j�R�Ԁ� !rZh?�o^3�3�$�����$����+�S+\$���3s����    ��    �����6  Q�̇�	��D$�D$�X����  ��  h���p~ +<$�ց�   Vh���p�������^;�#���$������������Q�$������3q �	��    q ��   f�Ph�Y�p+�$����������V+�$������#F��� �6;؁�   �D$�j �#�$����XQL$�΋�3A�� �	#Ɂ�   Ph�Y�p���\ej 3�#D$�XR��$������B#�8�$�������$�����w���    ��   +�X���  ��    f;W3��_��   f�Q+�$����Y���  f;V+�^��   Vh�xR3T$��ԋr�ڋ��+�t$��������S�$����#�$������#s;��   �Ƈ��h   $$���$���� �];ρ�   R+ҁ�x�   vw��+�j 3�S\$�+ދ܋St ���   P+�$������3P#�� ҃�f�#������  ;P#�$����X��Ҁ� I������o������O��k�a�Gt�a^[P#�$����X�� j W�����o�$����l$ǋo_��P�D$�X���Vh/m��R���   K(A�'�}r�@y�lh   $$�   ;h   $$�zZSR#�$����3T$�Z�u�   �U�V3t$�^�FhF+�R��;�#�!z	zZ3�_���1  �PW����	+�_hbg��W����?��D$�3�X�uW+�O���I�0��3��S3\$�+ڋ�#{;�#�{�;Ӄ�h�2��S�܀� �� !K	K[h�I�0#�$����������W3����#O;�ҋ?�:�H����c`޿����x�� ��   3��$����+�S\$��3K�ߋ�d$����H  j P��҇x��f�̄�xXhE��+�$����|$�+�V3�������3~�   �J��1��m�3�h   $$�� �6�� ���_hE���	   ��R# ٞL�� +$�� ��    ��   ��Q+�+�Y����   Sj Q��| 8�$�����Q3�+ҋQY3�$������<K��   _�uh   $$+�Z�Ë<K�h&����uh��ΒW��#�;�!w	w_3�^�R  ��j�P���t����^?Uj[��6!pX+�#�$����^�E��E�    j R��u �J#�$����L$��JZ�Y�Uj V��;���F#D$�+D$�F^�������Ё��L�)���	;X���"�3�X���L�)����   h!R��V��#�!N	N^L$�Y�Fã5�'h�5�'�� +$#���    ��   E��hd��RQ�̀� �QYT$Ɂ�Ё �Z�~W+�$����3�$����_�}�V���6���#\$�[���-  ���Avj�P�ąl$�!XX+�3ݻ�Av�|$���f���3��$����3\$�R+T$�#�$������#Z8�$����Z�������   ��-   ����Ph��P�+<$�   Յ��   �CW�$�����_CSP#�$����X�����SWj 3�$����_��T��>��;�+�_j R�Ԁ� 1rZhT��>^�^�u��%��h����u��ƻ��ƻ�E  R3�Z��[��$����L#Ʌ��  hwPA8S���    #��C[h�u+D$�+$3�S3\$���3C�    ��    ��ʅρ�   3�X���u��   ��h   �
{�3�+�3�$����RT$�T$؋�#Z�Ӆ�Z��� ~ ��   _^P+D$�X��	   j[��67��h   $$� j�Q��#�!QYT$�T$�Z�����Q�̇�	��+�$����Z��&  �y9E���   j�S�܁�    !{[��P�ć� ��3�$����[J���   �"�]�j W���    �OL$֋O_+�Y�{<�|x��!�jGh]�'#R��;׉rZh!�jG^3�^\���    ;�E�_W+�������	   �������h   $$3�_S��    K������    3�+�$�����$������    V3�$������3^#ɋ6�� ;Ѓ��0   3�[Q̋̋y��	��^W3�$����_�� Q�$�����$����Y��E��������   �xQ��h   $$����B,�\S������CK��B,�\;��[�U����h   �3D$�S�$����+\$��܋C;��+�$����܁�������P�$������X�� �   ��m�3�i�%���Ƌ �� #ҁ�   #|$ف�������P3D$ɋ�3x;ʋ �����$����t$�j 3t$�t$�^P3�$������Iȫ6��3p��    #�� �   ���   Q�̇�	��h"�&Z3�Z��"�&�� U��S�3�[���SVWj P�ą�1pX+t$�^�]��j P���    �   j[��67���	1XXh��J���Y�_��������W|$���_��    �?#ҁ�   �3߁���{iR�$����#T$ҋ�#Z�� Z�����   j�P�ą�$����!xX��������O����Jp 9�$����+�_[<�s|h��8�W��#�8l$�!w	w_hz�,^�^hz�,��    +$��    ;��   �[x�;��	   ͂�������$�{ V���6��h�`6[3�$����+�W+�$������_��;؋?�ك�3�+�$������    V3���3^#��6�    �����`6[�3��©��h�������+$ҁ�   ����O�g��O�g�h��H9W����!O	O_3�3�Y�W#�$����_�U�j S��| 1{[#�$����_3�j R���   T��C��>��J��h   $$	BZ3D$�X��j R��ۇZ3�$����#�$�����ZZ\$�[2#�B�   �Ƈ��R# ٞu �: �����������Wh����_+�_;E��   R3�+�ZF;s�!���j�P��#�!xXj ���AI��{[�}������GP3�3D$݋�xۋ ��)�O��k�a�t�����   O����� �|$�U3�_P�������Ё����    3��$����R3T$�Ћ�#B�(A�'�}rB��ށ�    ���S$�Q3L$�3�$����Y�r�CRh��T$ȁ�����V��n��m#t$���#V��6�    9t$����Zh�8�$����r +$�� ��   ���j Q��q �q�$��������θ�qY������F��3L3�    +�^j S����1K[h3L3+�Y;��� �Y�Yh���V���!N	N^#�$����Y;���   hs.�IR��#�!J	JZ+�+L$�Y;��k   h��§W���|$��i}��    !G	G_�$����X�u��u�	   �c`޿���h���h��rQ�̅Ӂ�    �qYt$�^�u����S+܁�,�[��#|$с�����Q��f����#y�    �	�� ��   ^�$��������/������Q+�$������#Y�ދ	;�Vh���^�^h���;��Ƈ��R# ٞL���8vw�+$�    ���� U��j S��#���$�����8(�	{[j Q��#�#�1qYh.�DW���   _�u
{���WD-b�h   $$�__Qh�R��S����    !S	S[#T$�3T$�Z�E�P�ć� ���$����+\$�[�uj S�܀� | 	K[�񤮹Z+�Yι 7��h    +�3�ZR��VhK�^^3�t$܁�������R�$����#T$���3r8\$֋�5�;X���"�p�n��z+��   j R�Ԁ� �r3�rZhK�^W�3����w�|$��?��3�3t$߁�����R+T$���#r���8�$������$��������QL$�+�Y�]h���W��#��w_+�$����3t$�^���S#\$�#�$����[���UP������@H��q�T��+�XRhq�TZ�3��$������    P+D$��$������P�|$�c9�� 9L$��߁�   �j W����    ��    �w+�$�����w_3��$����^3��P+Ÿ��ܡ���3ā�    S��$������C��    ���J��1��m�3�i�%���z �ȃ�h��ܡ��    +$#Ƀ�3��   �8vw�MPIh   $$+����� �D$�Z��RT$�+�Z�]P�ć� ��+L$�Y����   _h   $$���U��
�D~��
�D~�3���D��,P+���D��,�|$�O�X����B^�h�B^�;Å�+4$���   3�+�W+�O��[1Wƀ� �3�_Qh[1W��$����#�$����W�$������#O#�O�?��    ��   3��3�P3�#�$������#Hr ��    H� ����   ��G��aZ����Wh��3�+|$��$����������V3t$ˋ�#~8�$�����6�    ����    �#|$�|$�������V+�3��#~�} �6�� ��   J��������#�$������    V�$������3N�    ;�6p #���[^_hq�4�P�ā|$��b���XX+�$����[�#�� U��Q�̇9�	��h\F�1Q�̅�!q	qYSj�R���!zZ��������O��ǖA��|$���
g+�<$��    S+ً�{�    �� ���   W#|$�+�$�����ǖA��� ��C��>��J��1���3�R���C�b#�$������#z�� z��ʁ�   �]��j�P�ą�!pX�������ց��S�;��^V#�$������S�8�$����+�3�$�����$����3�S+݁�I����3s��D$�Z�Ҁ� �����   Q3Ɂ�]��   �u
{���WD-b�)�O��h   $$;�3�#�$������    R�$������J�    ��    � ~ ��j P����$�����Ub?�pt$�pXh�]���/�9Ձ�������R+�$������3r;���#҃�3�#t$�#�$����+�R#T$�T$���r�� �#�;߃���P#�$����D$�X;��N   hn��.W����    �+�!F4]ң�Y��*�O_3L$�+L$�Y����h͓K�W���    ���G_D$�3�X�u��S#\$�[�u�uV���6��h�Ǳ�#T$�3ԁ�����BQ�+ʋ�Q��    ;ދ	�   �ĭ�s0�.�\e:�H��    ���Z���Ǳ��u�u�   ��t1��t1��������D9�V�$����^�T9���$�BS�����E�˨����_���[^_j Q���	QY������BJ������#��Zhm�{IR�ԅ�#�!r	rZ3������΅ʀ� +�^�R�ԇ���3�X� ��t�6�q�0 f9{1o��s�2/�#L�>�<jkT֙���:`�����@��*`��O�$�^���s�w��Xv?y�.޵���@E�v,vk�AI�� �bp����S�*��*�pNn�{_�2�4��'kdp`K,ns5����E5$|d/��$�J���7�Fk�*��bh篹�1�'q�Q��,�w�~��Jo�-��Bҡ��a,z�1bƠ,}4��5�">nir��(F�8�T�ӓ�Y���Úo��R��C�#���? {����e9<�(�|�#��)����'L������Kg����x��M+��4cW���	teʐI�8ta6R�)G&BHq�)C��<U�ox{�$�p"E�����-��8���c/ϭ�-�~XPu*ha�5���E��Tj���z F��tJ?��Z��n�J�N�(��V(��.4�~;\IW6>3����A�_���96��kП�B�Z�������o�B*���;9 �rF(=�D��㧨pz]r;o��s�I�9?}s�d���l����0�@���vr�h����&��.�!%wv52�>d�L����&���5��B�g�t";T5t�RLu;��y�s/
�Rؒ!��k���u�������s'�����_���C����%�7G �X�b��x�:�YfH�d�m�O!4�NZ�%7�]�rXo^0�P�����<�'96���8�ޤ�p�!�,�e��}:���>�K����Z�J�Jn�
I�7���Goa h瑉D���]��r��m�=_�'�ك�WS�֜^��H?����
U�v,��P���QQ41h+�����ֻ�h����#:�z�d ���_�&��sC�)*!�N#��b���K�g�қ�zlE��6�Jsy�k���tB	�KYzO��vr�h����&��.�!%wv52�>d�L����&���B؀��Ҋ�t";T5tΉ �ӎ�Me8�C�͐.�����x_�5h]g�U�O�2�Ɇ�\,���lT�����)�)n�KP)�MntĢE`����hR?<Z�,�D�*��	"����#E�8ta6R�)G�
���"��=�ѐ�XHr<=2�%D�`�6!�bĽf���9���\��+����&��٦J1q�a��wU��F#�3�7k��צ�o@�Ȗ��o�4�O �����;Y� &�/�Gl���뙀�?��tNZ�r��G��٦J1q�a��wU��F#�3�7k�_( _�W������m�ђ��7���B��8��ϊ�D���k�i�%i��̣������;E�4:AFAi��E�ah��2FdR���c,a�kBZ��;e���f^��}���qC��|Z�눒" �a$�#X0�縭��`��b/"�Q�ob�FpL��n�Co�c|��~1Vbv�m�]�+ơ�Y�¬�tq�3�2��y��\Ģ;
&�1�U��¡L��_ @��ۿ!�T�z��ǿ�\6�����D���w��b����m�O!4�NZbӞA��<���x:j�����<�'9��q���/�y�H�����Z��n�Jl�� ������ӹ�B�b�߼g���4_l����d�'��p�L�#ֹ��������-|_g�Y9]߱bT��uZ3d�9����	˚M�L]�Q�	�1?c �qC6����l����}Yr�n�d��k���M>�ϘA�K$r̘��:������l"4�A���67{���U����`T]��^���s�w�G�۠L��£k�X)��vO��y`�`v0��/��2̈DC!�$��u��_{���B8קB��6�_>�v=��я���I�CKJb_�`?�7V�blCH'�t���pſX�]���u�2?q<�߷�έնS�6:�                                                                                                                                                                                                                                                                                                                                                                                                                                                                  �q  r  �q  �q  �q  Hq  `q  zq  �q  �q  �q  �q      8r  Pr  `r  "r      0q  "q  q  q      �p          <q  Hp  �p          r   p  �p          pr  4p                      �q  r  �q  �q  �q  Hq  `q  zq  �q  �q  �q  �q      8r  Pr  `r  "r      0q  "q  q  q      � DrawTextA GetMessageA �LoadImageA  �SetCursor user32.dll  c EnterCriticalSection  n EnumResourceLanguagesA  p EnumResourceNamesA  	GetModuleHandleA  2GetStartupInfoA �LoadLibraryA  -SetEndOfFile  `Sleep oTlsSetValue �VirtualAlloc  �WriteFile �lstrcmpA  kernel32.dll  # CoGetCurrentProcess 3 CoInitializeSecurity  � OleCreateLink WriteClassStg ole32.dll                                                                                                                                                                                                                                                                                                                                                                                                        3� �u�f��                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    �1��橲��*�Iq��lE�i�����"�@�)�{iȃ�bMp�>��
������m�,�ʯ��:�V��A���8c�9Ql|�u{��@+���^"*N	�����k��tȧ�/)^TܤCt-kqO�`�����C׽O]�G\�#AK)�T�I�{��}�)$�++ZF����7ֶW�A5�r,)޴�8@e)�6 J�}�y�dQ���HTTgD��h��!�~�����VɬeP��˾�M�PG�NK��Q�,D����͗M3�z���j�	��o��GN;����{�L�8k��H��6Y �0��[�S�F�q-EKRNcu����h�OjP���m�$�~�0����)߮bq��_��2${��C7!����P!�qϘ))Ï���8HΠs�^�lC�4� b�� �i�2E�(K6K��M��od�f�|�W�;{�M���Y.9hߖ( ��ajWN���L�WN�;�	���Q���2
8� ������H�jblLO�� Olss�ωC����|��0�Co�2�HDd�Y�K~mz�ɸ�z������4����K��'�����c��v����tJ ���y���t�
��2Ro4B�#	ݼ⯺�t<�Kc0�{����A]��T^p��W��N��hG�9�M6��ۨ/s>#���$M�Ѝ��J��LQ�Pߓ����S�����i��D�vzGT�-+���b�)<�AM1zUp�^R�M¢lO!t?��-*�2�KY�_+䂕H��C��&�3_��W@P��R}Hf!��@��5�B����d�-2�g�1.��J)+|�N��� �/�E���zZ�\���?�0����2,3���]��L4��`���D�5���%7g�u�픖&�+cw}�Z���q'�:����R�衘��YWM�˖�-'Ba�,�'�଀��V�l�Լ�<�{1�`\��`_�םG��AR�p��y�~�����b[n����'�o<���KI���4<���	�YU-��]y��<}{I��.I��}уn++��ti��e;��=e��2'�,Tov�t����e�u-_q%��h����(��=���vE+�5;�-:���Q�䱌�}t� Dٷn�u/��� oKbԧ5s(O������JiV9XТݍw��J�p�>��[�6g���	l�tv��5W[|-IV< �����k��Fx���k���Qk�gI00\����>_u~�,>+槗�}��%]yb�a0����v}�DY��߼��Z��YG*=?j���}J���"X���Q������٪Ӻ�Vg�}����ߘ��E�vZoғ���d�-�BX�`�����>�<adA8�8H}'���I'g��|ʟ懛��G�7�J%�l��I�É� ��+\{*�h0f��B�O��-���'+Wi�
���J����M"����d��G�<Q,'�N�x{���T3�8YK���a��� x@֏)�<�z�p1�9xv��-���Ò�<��;y�W���&��yC90^d2& Ĵ�ߨ,�q?6�[|"��/�qNXdp&���ؑ�W��ϓ�s�@[�������b���o���TG�3< �Ӛ�i��)�D�������7"[���q����p�~���*�y�N���3���*��[Y�Ea���X��/�+�A�����iL��5r��yd�pA>�;��<��=PY9�����gۤ�B�m�x�<JK2��z_����������;�Gͳ���tr����`jDy2;k܉���V`W
��=��i��ib����F�����`M���E������AX�5�~
�<�h��U�p)������DK��1gw����"��OrW��4dC⺿@������},82|E'��#�R1>
\ �.o�0f5��*|v�2��+~�m�N(��f6��B�3⊅�����]�Ef���RQx�f�Mm��4$�~s*�O���x LUR��,PO�F�K|�W��ce������3��GI�v���bnݩe�I��%y�ǫ����Z��P��L�ն�l?�=�x݇�đ���T��?�梞ԕ��{����2 K>a�U53��a�X���s6�qX%�p&`�۟�pS��
'c�5�n}� j���� $An@���x�-EOB2�=a1pY�N|���*���Cr�k�� 7lk���OLSF���Fx���%�PKzw��tp4��%^�S�#G�QkJ�5���p'�'���د���K#��� J�9��^�� ��-��p�B�g�Uȕ�OZ�������PN� Y�������T���Фo<"�N;�f��l�@&j�4a�q�h�C͛�ϊ�*�'��N�"i������Š�@�S��"`���q^���ؾ|~H�zi[~��E5y�(��h�/�O��[n�B�9ȉ�5"�,����ީe�;(ȴ����̯������(q����d����:tn_�`<@�&b��b\���! �i@I�VJȃE�xD�|6��>O߹�@�����8b��E}8]L�+d��39�;h��dx�N��:E��:�� ��e\X��"���Sa�t0���yF�! �KM���˔A�x�RV�y��� ��h�딬y�Z��Tga��KM����gj�A�6+�ɨo���L�Cg�֮m�U�)>��jlT�g�Z�tN�ݙ��f�����8�h�ސ�l�X��c��b��5g÷b�SY�5ӭU�]�V��e4�c�dO2�	�;��*R%O�ai#�r���Ve�j�1.�t�0� �y��ӿ�/�:�
{D�w�A��]�ىa�\�X��~{�����*��-�k(��XJ���3�y�QpZX,���r胔kk�Nԗ�H�;�3�A?����I��{�4� �}v��<֓5���J�l�2'$pǁUy��Q�#ѹ�Y�����!.��+d�	��C����9�*1ɶ�Q��8��5|��9�P*��K� ��cm`�[L3��;��>�W�������Z��Q��*_����K�ܥu<���i
�-��G��̀�1�B5�{Z�8oYR���'[l\�����9��=�֌o�eI���<4�'F�cMPV.��>���1�x �_���$A�Te��j�<��Aҧ{���y~�H���=�7q��0�E �R)rU^n����i��Q!]Il�Qz }
p�, ;yϪ(���Т�M�m�N$�T6
C�U�3�R=@O@������}h�2?v��6�&��}�g����C����_.%"q	��E?m��CN�ۑ�)w_U���$�!DB���ACIq�d�+�[O/�z�Gl�Qemc����؀�N�Ȕs5�O�L��#�5���m(�7II�����;M!�6�\�IƋ�BVx+�
+�������z�Iڳ�w��r�(�"`^c�5�qY���$(� �?����ھ�� �:񍺢M>@d�J���E�����H���2˸�kN���/ΰ���i���>�uE}ݚ���g:7l� �� =���Y4���{?�ͧn�� 	1k!).��?����D_�V�E�R�vM�c�J�O�*� �=jD��w��N�f��oB��A�3Lae�`I�=O2��۸� 0~<-{����g�"VHR$�'2�֚Gc�|�;yBɰUѦ��rzh���	��^ǥ���&�-ſԭ�3�1/��[���M�^��o�-���z���-j�ٖ�s@]������4�g��r���;^â�n͇+Z�Ox����F�#�2���M}k�}��VnuZ�a��O����ZT�CC��.@L�i��g��\������'��
ݧ�؄�uO����灩�%����7g��L��E�|̕��PdA���� -$�\���HK4��]��"f)�緽щ��@`�D����VX�jt��^P�o��<�����%���ML,x
^�&l��\���B3��ťZ=F�l�r-[��f���f1w�K�>���M] +�q�*J*L��X�<~�W���w���DƼ��g=�$D-���_�gE����]95�St�՛�!ѢT
����x��na��2�����q9�Hm]D/&WJI��i����T�0�,.��Ҩby��ંVø�f�@�N�&��:��G*Dň���+�L�Ң�C����G���bR���b9D4�:��]�@�&��zb���j|�?v�OȬ���t�s�;��Dv�c�%-�`��l]⫥)B���O_0��@$;N۫\^��Y�]�b�p�������}�,���g�=�Enc�fGQ��۔T��Q̙���5���ǝ���&�E�E��ym'���Ӊ��oҳĿ��Y�R��SW_���U�y{eC�2
O�G+-f�!���$	�&[Ȁ	Ws�{��q/���8/Dږ��r�D�L]x�t�VS_���)w��{Ԩ�ab�}�����������������?���j��$>8�8���O�^��?�`�޶G���8�O�5SSas��X�
�Ø1�Ȳ?�L�f�t�y��IiiʌƋn�ե��[��/�{��1��~�^�Ȑ�a/�0�v�X7�n�N�{��۹@_)"#���E m��=�f�rvb��?��U�\6�fI��r�vp>3��FI�&-6�)>��Q�͉�u͡���oE�V$�������o�v���4f����8�j�/4���2���0���������Y&ș)?J���7o��Iִ2����D||oe���i�X"$3+G>��j��^󓢼L6�`Һ�goq��2m���=4[�S�vvk8.�u��;?��:o<�����iG�s{��w��vxkc컍��8m�^f�x�O��g ������l�^BA75�f}Χ#���c������/H	)M;��(%ҺuV��Z�O�9`��e�Rv��ǻN�0=�U��@�Ec�a�����T��gk6'�>��'�K/�� ��l!�絁��yn���7����^��6pg��d���M'c�I���U�W���kS�q������K�{}-4S�V���,$��^�D��`Te�!��jЇ.ia�;�V�t�-���>�1��T{������9~c����;�6H(�wx�o��.�?����J��� �J����+%�.�>�]z]���nd�4���Ѐ>X�5�
Jb�K)����:�=�UAS�φ�b�(({�z����@��O�^?7!����Uㅾ)�� g{��Z�Y�RO+�3�HM��tE��"�0�HC"�IzF���q�@e����6��٤�*;������.����Ѳ��n��4�݄Z{/�.��V_����dE�`ρ�0jČ� +qx`y�ܩU�����H]��� .��Q��i���"JB��ؾ��)��������ne�]��a9�#B��3�8�l��xDP�)��$M�%��1�{�;[@�ࠪ��O����%��j��څ>r���t�:4�a��t|��ʼ�:�o�R�_�c`���%ZL�6[�h���F�Hl��t٨�`�!e@��wL`+�i�����b��	���������d�b`��m��Vau�]A�R�?<��W�N�,ĕ0�aY�0?���H�7����%]͙�
i=6���G(^�j�S��IP�f��/� `��]� ����Z�a��N�f����[7�{�Y����=��0�sZ~�'P�[y\Y��m�)�����k�3��)����GWxn�o�?>p6̹z��}g&]ji&Ѕ�bTN����K%9!^��Ӧ�J?��&�_���%�DL�]iIɄs�'n��L�#9�J�:���\�4����F��*�9�i�q���۩G����7F��c���'�nF�d�B��Xp��mI��ݸ\�(ˀ��I8y�(H�Y zK�^	��	���XqP"Hz)6�,t���^���^c��]t��x��0���2�
C�]!Da�O�'��H��pl�+��zh��7R2�3���Nf��t ��z~��`8���<��SBۮIRD�~׋:>sg��0f^v�Cu���IY^�ts�L�'���n�醌��Ķ���+�<X�����p6�@�>����"��
�D<)|)R�[�{���`�?��� l\q#��T���T]�ρ��X�ڿ����Ļ���L�r�Q�/�r�lF��q��;�.��Ԗ/BQ�N�ڰ"�*��"^�ӑ���<)�Жc%$""g�)��{� �2n�J\��w4�=������k5�w���o)��yJH��X).&D�R��#o��b�l�S!T�(*�#�j�8��JD�!����*�dA��@�} �\5J�80���w��J�$��3S���CC�pg�=m��u�=�s.c�Q��r�Z>YT�$D&=�l�Ua*��_O��O��&xm�x�=�K���� v��������e(�,c��Sĵz�dh���o �?����G�~\�O"�p�W7�V�VT@`3A����_d�a{=ԋ�<˰���(����ֶ��m^�ɓ��x��E�AF�����i�� �*od�uٹ��@7�B��U��l%���<Մ�p�/ =6���#"�%�[V��lF��g���W�o���RW�֙��d�֭�ud���~k�f�\4k�Hh��*�܍���@��B�)ȸ�����0b)7-�Y1d'sZ����\��#3����Tl#�#�1!��(=��7����y�w��O;�7
��E�A�!brv�8㜾��(�4�un-��MX,�6�t��!b+�3[q㭨��S��ܫVU�{tX`O�
��� (�$�K�lV�aa����B�	�b��{�Q�ٮ�@yvp�W�I)>��Rs	�ud��S�K��J����rQ��N��i��`�� ����
��$�#Q2ޑ��J��k��A�Sa�`5��s䞧o�V��8h�]M�|�"�9���$ W��6x
v7Q�7v2�3]4TɚoI-�+��q/jCI�v?ko���iz�%<�� �qW����|�t߷ܺ�,�QK�F�P<֥ 6�#���5f���x8����~� ���Uއ������X��Bx���w ����W��1� �˃K����@5B"	8���4��7+~0'i��c�"��/~��][�ɡZ���+�V��;9ވ�/�F�6)�CO�}a�o��� VeЂ�[zQ�(���w�NN(̇�AQ���C�����Oc�[&�bҺ\^ت�2���
��c����{d�%>T^ѡ[��w����ʩX���+i�i�L?�*�x]	�e �Y����K4&!�N�p-H��M���������S�P<�w\��#�a� 1�/��{~�+p��j���1䬢8V�V�D�� ��.28��#S�v}�r)ze����p��묂��D1B��*��&HO�
�Յ�f�!�D�N���A���v�j=؃m�@�}y��y��μ��74�'v���3ISG�%�&N?Y3�'L���Q�!Rb̡zA���Z���i
����6�~�6�u]���Z���)��3�kq@�?tk*���:�kKn� �QXxsjQI]$坙�=��}��5
&�X:C|����O�9��8����������v:#��I�(�Ү��F��8��FK�@�xA`G6l�vA�z��Jn�ت�����FQ����i�u��v�]y#�%A�3��Ŧ��:7\Q���}��s:����&D����z�����g�ϧݥ�l KmXbF��+�/����EgX��36��.y�K���2"^�l�V�l@�1P�U�������qB�f43;�Ω�3dЌ�����R�9X����'��LH�/�c�,���|I��q��	RW&\)\ ���7Czw	����{D}#�G��AA@ [��TD��9U7�ɮQ�b��u�R]a����P{�sS�]���Z�8��$o!��hKHjE��zS�N�=�ۦ=_ޠ^	Dg�Q�^ �,�T�|�)t���������]�iry��#�p�E틖u�A�J�g�1�P��O�o�Aܭ���[&�`Y	\��Hd	�nۗW�zy��A7��&�r+��:oL�m���XWCo������Gښ���ps��*,��K��-�A���?�Oѻ�n��*09�[pJbJg5�:J�D6����9��Y�������IFQ�� ^��o�].�Ȍ9}T�sBfr�ڐ�0��"�O�E�"�����mx;��]knB痦90Q��x�����m�e3�K�@e�ԝR�S	�Ε�US����k%�^�r�	 V8�M�͏��K�f{�F��(@�o�R��}R3�o9�5���o�����}��'a�i��	R��bO"���q��%����%�%~��N�k��1�� 	޵�]��w=אlu=��֒�AYEU-3dBtS\��_p�n[��}�CсJJ�o���x��(��{^>_GF^�g[)88�M���:�r�U��a
��};c��7�F�J�t���4���<L�m�@��N��2I�b#H���^B�W|�w,L� V紳����[���ᆾ?� yd�Y R[j�>;�Z���O�$�E����[fwor�6������[$����+�T��)�>IڊUí�u��r�G(וNۧԟ���K���l_?	��
��x8IG��{+Y�����{����3k��oj|��l��#iv�?��X&)�����*q4_��f�3��U\}y�V�{��4����4K�gj��@](��D�!~���C=]e��P�g�@	ו'ȑ_�J�Ԑ��"�i���C4��c�<��.2F��(:<\���<5�m��'N�v��Q�Z+b�gG�v�1p�o�����a���7@���E��D���-4��ĸ�ͱs�#�'�?��Dx�2��IE������������Mq��*!����:�O�^��S�1���(�G���?��<���!�M}ז�7�J�Ͷ���R��!��O+�&U�њ��	0
��Z5u5!.���5����y���I��Bfi�g'm�!e7'	+�,#�B���?� �	/�[�IH@��O��ʘ����?G�^7�}�����!�/�N~
x�nD� ���ֵ}�b40dK�X
+���e?�s��;m�������d=��C��W#����4�TE�f��6��6��F��ؕ:���C`��n��������{!�)JZ�r��*�2*O&�3sB�"w�C��� �ٱ[Ced�\l�2�u��� t�t����`ck������m�ƈ��0]Z�R��)�MN4��(�z�B&�%�x�W0_^��W�.�~��_����L���u��G>��	�0�<(Ww�B�ț#\6f��l��_�@b"~�KS7����'4L�o������RT(<�Hz?*����z3T�ĵ;��:�"Cj'b�~0�%�X��2^TuO���,�f�P�W�d����U�W��ض���&n>Q(��B@�(v1�i��%�7��r`ca��μu�-�JW����%�7*#�[�T^a�Ј�C����6���k���zu����´P��l�\!s�j��Ƌ�)0(_���t�_�;^�Kš>���������r|4rp�RN�8,����w$u+�`n���/�I�ȮIk� z[��]~2���޼ٿx��J-�@�l��w��n���Q��1 ;2�IAp�_U*�~xE2u��J�닆��R/��_��.���]�O>��c�8� ���Ak�R�T�7��Q5.0c�M~7:���O�C��"���ItՏ:Px�\ �����&��xOd ��W��C)�F��Y���AؖH�B��*Z���gp߮�����i���k(ůi8@��\o�cR�6*Z��y�p�R �J�l.��GH^�<	y^M�*'�TG�֣,�B�
Hm���!�iV��O�U{+�c��9����⍆�I	�7�ܧ��a�j�����4�խ�t�v�^x�(h!�y+#!5�r���o}�mqm
��aέX$�U�+� +���#�d���LpٔbZ�{��p���J0�0∹��k��_m�=�$�EF�(������3Y����J;���~�4�4;���X�$Hz��/M?���5�!�2C��S��uZʓy<1&V�.�W��I�<��e�W(���owᾆ�\]��Z�.�T]�*f�ۨP�R���SMV�C#?r�6�_I�G�2�<gkR>�!|.	�Ԭp�������~>s���"j&pC�;�7��BNTP�oO��":u�Ҟ�4���J)! �4[u�����v�o|an#���_5劾��-��������Q����C�r��g��[��;�j���X�H�����g�)V��W)	%֔Ж�f
��i?JO� :m\��U[ �׸J~;�L7{��Ϫ8Q�Sh&�*��g�V��A�{���ɞ�r�fC��1�������+(o4�Ï*�@l�W����{7�h�\��r0]����7���Q�:{,�$�{l�m�Xk��d	d=zm�$�֫	�Ft^�X%E~��'ག�uwg�����ҍ�}�qjȼ���?֎gy�)�����{���_ �w`��s���V}��~�[5�	8ݸ&W��ն�'4��(�	x�Z8#W75�������MJY�7?95-V�����$Go	/�����0 >��Lɼc��V� ���U��P߅^��aN�0R������8ʑ���R��b��9�����n����M:�pP=�����}�~����i߹M%�m�ڊ j�W?�w"F�"׽h�-���}���}
��n��������Rm,���f �&�"�%%�!_c��H�#�3�9[��sQċqI"+�h޳4+=1d�$!o��4�^��]CAv@^׾�(O*	���0TR<;�am� �"��L>dt+6��"&Vn�d�ۤ����&-{��xc��w:Pm�^�ew�	UB}�y �ס3��<(4b���#�!&A�LV��=9pB�{d����wO��>�TK�TC܆؉dl�.�H��p�
''��Z��3h'���'�O�ÌۚFv�D�}��K,Շ�4�ۗ������W�Λ�6��ŗ�5x#�u\cb��-]���\�4���L���1��,������'W=�x������1���N��j�/)�<�(1
�=wY����ݦYAg�4+��|���ƌ�j��S�o�j��>�#1q!�}�*��n���:T����V�k�e�������R�i������"� Ov\�$�_����z�W��Ͷ�}�fP-��O���H�"�w�ߧ��}�;�j 2���>�|Ōҩ��(	��9��$�bY�\�|2L*��R�}��V�~ qI+r��6l�� :���ndl�����Hڻ"X�
�� ��Mу��c��4/��V�t��C+����?ӥ<y�T�ż�'5��Ǣ�N�[��ڢ�7΢�+�A�8�ް�E�亟Dn�w�}��w��O	�F)+,f���鴛�%�M�bk���,�\Gc<i[��b�N{��F�n,����������}
Lƺ����캧����Gk?A��E���5���{���vR��z�.㸰�u�p�Ϝ����k#�!� �O��9f�J}*�SWir+~B�/U�B�{��1p|�^�(iJ�q[ԇˁ���U�4�)����R���[�خ�T�2�󛌗��n2��dhiY��dm�b���p��d� +�a��E��t6&�u����^Z)�j#��b�e��e�?�N�P�+����Nr�-�h�v�%��m~�lg��+�����'�ťbU_��M�Iڨ|��0o�L��8a����Oڐ]z���AyY��){\��:H�$:��0o
[�zF�i#�b�Vd��T^!�E���j>9I)��������1�3�$�J%�Q�z���If�&��0�����7�֏|�H,�������K%U��Ŭ5'��\���j]�r���}��~P�WY��hd|�NÃ̆=0�@�xz!1a�!ɧ�����r�4�~T!4h����'�yH-7e��|b˃�ca�_B��8"�Y;y?<�_����t��d���s~�����6���F<s�e'�%������	`m�t,�ϓ�%�ܣv���MW��-���|�B�j�l)�I�66$��!m�^o��tK�9A|wƋ��}{�͇.�_$G��d�]�~�~/�����x;���z���*�����rZ���wc��l��#�fO��n	�̔�H�%)v�)q�*�N٫i]@��d�۩?,�Z�~�57ce@,���s��v�ue��u��G��"4�*
��j��9�nhu�{ZѼn���Xf(7u)�Sc�
��Cn����.
K�+�~9	 �cn`�q�w+;��Kr�O�},��ك���h��4�cb������[*�ĉ9�+-F���Nc���K��e���s�c(�u
�f�Y�Eq<*5:�v�j�k��\"��X�:���vv�)��aNAr�g%�ӻin�|� ���8�*�%��Oٷ]�p C�WR5S����ļ�EҚ�_�X��!�k�b��i& ���B���g��:!����`('��zG�Q�%�xR��W^R��bz����V?v�N^z�����r�FC�����1s�oy�J�V��v�}O�¶�K����6H�z@-
/��kJ��'����~M���U*E��l�z32�m4��B�̱w�T"�
b�H�ɝD
+�v}6˕\n��d��,ۏ�F�����<�>m<!
��_�E�Z���	,ޠ6�݇w_?%����Zv����Z�r��s��{��!@��Z��˧y��Y(��Ѐ�]%�^-�
׼2�*<ja����b�k�j��ZU60탛k��~W������ZM)!�с�,��/�:D��N2����nLJ>:۠���wU��$�a�%��D�Ӡ4[1���x�[��޾*(���D��P₸Y�UA
���n�IO�"� �^6�K^�Sg!B��`V.���CkKUSP��RTU���aV8ji�f�Z��!@D���	�L���t;�唓S�z��X �rE��Nx�A£�������U�ʧi{�	��������TG�`�O�,\h�����$�4~GK���S�Y�TWh��#	~Nt��ɜ�L����s&D		�
ɜ�����0��c_�����V4��<[֖�7��9˛ݰ�/A�1'GE�ݖ~� f�7L�^6B&�4*o�&��\<��-Ǿ���T���Ф��9�j�P7��t�T�����\W�H2�M��f����t>���G������T8��s.�6N ��7�X�Ez��%��8)	�6V+�q6��9��g!˔�-�ǧQ��]��|"g��<n]E2B���#-����ZSf�Z�o��\/�K��+�O���&V�����c*؈����q��'����o�>���k�}m�R�$:?pI��=ҥ�ᷗ��	
�(�·���k�3H�e�_�ȅ	3M�[�,���/-�-T��G�����c/+*1�I}Zi�`P����z[� �g���i��&R�V|M��7ĬŹ ��`6
T^Q�S�B�{Z<QI��?���E�����1�����b��@F.>[�'K=�9k����ga����񗢺���>�������Ԗ~[q�d�_�*3'�J�����tm�<�̇]ñhw6����h\�C0�����{zٻ�IP�U��e�m�vh]��	3��4@�MNN�6˳��_������-���$_6�!��G�@bcs 1<���������Jwus����U�(�_~�.?~9@Z,�Q�']u��j�b�3�	\��&ȵ���w��#ԕ6tBǤϙ�A)�/e�E��Z!�!�D0�Ny����~�_Nt+S�f�`e�AIw�Y�oFk���~W1�����w�ps/���B��(�K(��G0�_�.X��ј� �]A�-�e$=�l*n-B��,T�:db�ٰB��<jVq���X~����kɍ�g�I���gB4���*���f�*ɋ��h](o�m;a��qSn�b}�p
m�:���7��=8ʷ�8Re��֌!�M��ZNQ�7��?�w
[4&�:��]��,������d[s�B
�m��`�4s�$�����Vȩ�J���UB�IXyzK$��7T	�, E��O���Z*�
��"l14 �7�7��Q�Y�����I�g1�3-M,�*����HLͭ5����z[���P��}��x�����G3d�̶-X�_�Cr3o�\�F��iwMסt7?B�9���A����a�����y�Rg\�5�U��vI��x]{=S(�ڴ�zF6lusЬ�a�lMy�´��c�6���^��HL�
=��cjLu��g�x^�����2�����z�u��ڭ(�7�j�ضL(l�
$4�n������$���]�⅍��T#��3)l������چ��W'��U|����(n��
���i��F:?|kĸy�5�!�/���S�t��G";��&1�<�tk�ԧ}��(��2ރ�d(�~�#�'�0��(�G�� ��O�.�Z�x����R���f�5�8�U#�.�u�T"�e�/�~�JԜJ�� ��[�'��������ɽ�SXhV�M����)рj�����At�D؃�o��[	�6���L�u��Ϡ`)�R��уu+.�뵀���s� dq���B9�����#����c�M�����@��*[�;�D�K=N=1�J��7�xM���-ػ��%�aTtY�"۩O�`���Я��,i���ˍM.:yX����n~C����v�L3]X4s�֨kل�|�G�L�xp� K�[͜n���,��L�1���ƨ�C�#��Մ��G���F������"�p���h�E�J�I|�kyN��<vN�1�h�F��S���#�C����jyz����N�b:�c�R�l�y*[�o�_�ۘ���c�e�O4�3UL)-��u^�_Dw��`S:�nοQ3�Ҕ����v�P�тCQEp�z��\���11.^��l����b�`G�9 �p�Ǳ9��'��F�!o�� ��$ˣ��k>Ԉo�%n��SX�"H0�b�l�r�F��xNO�qW'����GC���|VY�2ч�!b )��s��g�ಞ#�,�0��i�]`;�ݫ���~xd%ӮK�4?K$E5q`�>5�X�u����]u�3��B��{l�`�7����j=pwse�V�4u3n�
RT{'���w��3�3$(	��P��R�P�_w
������֛��
���}����z�������(r�NR9���!P>߯Dz���v�깶x7&�φ�N�N�n�s�:j�u���fɓ���M��Ձ��mr�Z��g�N��)/�4�6FS�� �پ���(:��db�k��Ｑ��вi���TT|[h���w1��T `�
qevJ��qI�QP�L���~l��Rcy�%�W��7����4f� ͟�c|�֥��jS^.������0���˽�fqD��I>��#&�$ޜ�I ������j}s�3П�(`�@u��)�"+�*�8Y1��
�w�ywO��E�	uVN ��z�?��\V�	�1�������T�X�+�^��E�>�岆,�^.�(���ӣ;r��k��\#�����[}(;���-��3G��W��<[K.?���s�EE�<�(HF�+��)m$�5��qo�A������W��|O��{Xq�������]<�o�Ab�y��1O��	��{�}�ʬ�ǃ��iO&���a�Í�i.��o7" Ν��Z.,�C\�>���7����$��ԇ�#��k;Ƞ�6��JՈ�_�e���.+21*�i]�"#=d��iec��k(Sᷙ�{�Y��?1Q���G��~$1M����rEupsN�ƅa�����r��+	���svK{���ܥ��>a��7�]�k�f=L�'�X-5�v6�u.��B�W	:uLn�%�>���R�3?3ʫCD��4��ձ'� ����E�!��$�8�z��E^���B�eǣ�(֟1T�D��������ٞW�]�b�W���μ��P��|l�>h�����6����T���`�VU�v�<:/z�&�GO��-P��R���g��_�Z�WH�p���b7�1D3W�)��;@���c�D5���V� ��|/'�m[�ȍ�ђ�)�b�h'�~sa�5�:�!T퐢�<*��E�3�Bc���E|Ӈb�)>䜨g��{���dx�����3�ڞ�ۤ��{�6h�6���P	@KMO���C �4���%�,��f�;4���;��ʾ�TSr�<�[-�f 3�'ڸ�~�\:<��r�i�g�;��������	DK�����-{:$V�N�4�Ѹ�<���=s��Q�_��J���0�u���=�Z���-�Y"g���hY`��ϒ��jcX�I���tx\"��������B��ŤzvJ���PK�}~ę��LV�fҕ/MQ���>˷7�Q��"�e�I����n��*h<������ӽmI��]�V��y�~>"+�sr3//V����㚶z�(L���<e��{��[>JA[n61�K��MזR�u}p�.G�vZ�g�Q��ZM���,�[� /xE�MYeJ��� ��99b�'z��l�8���$s��<be�ư�`�ݭt���G��tC\a)o)���P`�x��F$�#'����y����3D{J�7�%�E�S}�#��zq��2Fy2L�S돒O(�Ø'u5�.��#fD&��K�h̴�A4��q�;�0�.d�x���vg������ԩEۦM?k�_�����\נ�WbG��MD<����,��uP�t���e�}^K��Wp�`�d�bM��0\}������	�7z��}������n���M�2� ���v�a��a�K:�ৎ�������w�K{�k�ʨC�B�V�9�d-Kv�`/�1&��U��C�O�J	��u���<��-�(8��V�@���U��.��*g �F<���Oar��#�zqh�Q/?¬��|H	n��,�|�#ꏐӿR	_FU�]��Z9���/o0*&,�T�.[�=c9/���Gk�u�G��#�z��s�Wt���}�����\��~-��$��w�]�� ���ur�g+W��۽��܀�[O-�㍳��}�3�L�9ʎբT�ـ��7�Hf��,��#����ч4�en�'n�]�n��0�����(kh/y��Ʈͬ��4���rŏ�c�1�m��%��fݞ��i�vֶ�5tP^�9��J/�8�	&m�u�s�d/���Pd�0�1&��}�)V����W[<�,( e�=��B�Ŵ��T8G�:�$An�����om�nR�#]��iV��$�vc�GA������Ʋ�|'@M�P+=��n
��b���s���.�oT2R �}��nnDf�HR��h����U>NHs��T�0��z-�GLa��#�؂����s)�Y�� <�q.u��Z���r�n��y�����m9v:"� �4uθ���X�\h���M'(�����*�g���li����x���~\��f`k��u����-�M�0���"�u�ѧ�&L�(��^`pj�^u���s�KK�sz�k#��G�B�����J�o��\&B;���w�WU�0u,6>�u����H�P����9�ңS�@��m�\Ã�!m9�����".Hgy�|s��0!QG-��j�7ܰm5��� ����{�h��vU"�#G������9�x�qi�me=�����鐊��?��	�����x�[��w�m��_���H��.,��D�";��N��Ϧg]Q��c��h�D�?�FÛ$�eaEY�2;*��n$�U*�w�de*vn�%����fխ屬��"`�h{׫ef��FE-�Ԯl���(r�0�&Ó��Ó�B/��-�(;̴��۽�cjBUU��oP�
nǟc����29thm���&�u��㮘I��.f���Ɉ�ǿ�?C+�v#�o�W�����?B�|J�qm+`�bL��cNy��2,����!(Y��v`X��H�h;��2��P�S°�(,5Mx[�۫	ս�k��^�����Y��;�Ė��؊u��Ц�fk^8�<KA�����a�'���p�>��<y圱��WU78�-t�U��IkOHv� �'�
v=d-x5N*;�+�tzb�V�����N��L`_�y�fHm����Ӕ�8[�M�!nK����OF���� 0��~��W����?Y/
œ�4d��g/�O��;0�5kB R�������|؜4ʉ�;;�ԯ�ɨ����s�S����1`�*�U-ǋi��g�~�7 TW���9��f	R�1�� �Z�"J�6����1ׄ�7�F�;q�i�0_7������"��c�lt�������*��U���ב�}N��W2�"��/'�S^�-�h�wHǡKS��7I1��g*�ܳF�4��(��JQZ�r�*�H��,�t�=��/���j�/���d�ʙ!U�F��t`�������V��Rxu��jRc�sM��HnbLXOz1W��/���O��f����v��D�h��,�X[�1-��Y%ص�c����
��hg�A��i2�V^�'�>����|Jۓ�%�,o�(gBUި�b�:@����������XKǩ-�QN�_���8�16����"�^��� �"�AxxdȘ,lt����t�����>4�_U=6�I�@�)#6\jd.g��5�17��d����N-�'�>>MK���`)�;�s���O��܃���݆+Oy>|��h�"ѫ+kX�����攋`6����!�ad�M.�9�n�:TA�k�ր]#,�q$�UYR��
��h���œ�*���eh���4X�1�.��a>h�����:U�"`m��fm�m��=뤥?E_΀R�� �Lw?=?�Q��w���4�����0q�&����3�t��k� �͖���;�<��bY�s{��{��k�!������%��WB�w�ֽ+�6=[s$r�F��b�<����1���(=�>��4�6��&��CwQc�Q�̹a�&�I.�Τ�C����T�{�2�T"�=�2������K֎���������!A��K.��n���ڐ��q��5�)bCuEL#SO35-����*��ed���v׵��-;��I�8�+U_C�	FO��H����&���9-͌E�v���e>N���Y#�InM�-/yF���e���/�W�U�'|�5�DQB@�̤Ș,���-�㚈�/'��#�۝���adh꿚Sm"jz�.�M"gt<U�_��%���� �L}���F�>�M�J��oΦ�0/h\�M�J-�sck(����=����"{���Ƞ.K�����9�#�"��'�f���Ͳj�:� ��k7o3�w�<�C����*跘;fΚ=����6�wT����b�������'[�ut\a��)�_�omr�����M=���g�bh5^�Rj)%�1)ծ�Ϩ��[���猽��쨸��F�{>�5�,�$�*��o��Z�B+����gS��$�Mܿ^(����C�F���`�5Pe�8�W��|ԛ����;�7��&M��l�'�G5�N�Tt�#/�A@�6ĦN�/���NukF
-�	s�N���(��	����-_�J��r͡�:��j�Ϥ@�-�u�)�h��
e�F��HS+E�K����1X⧀��K�hC�q@[��ޖS���~6m �mڂ"	i�c`�|��^nWys�˜��*��v��/�s���� ?�ܖ��C~bt�U����������Ne��fo�A y0��iL����3�ѵ��V@�����Ȣ�����!�@Mw;z����&kZ���|��:V�j�d�j\;8rxfqBC��_=9Wc�_,�!��9+����o��j����˔�_[e=��_���t�uٺ�2��L�޼��:��%������noluA@���[!a�a�N�"#V�����Ra��Z�س�T�s�D��ȻvuU=�,9A�'���]�4�8T�I�Um xs�,��S!w��q:��7��'X��m��Ku��Ņ�i��B־N�Y�[脴�e���s���k���a�1*j82�UݕB�A���BWP7_v�u��"� �wp��;�t��`�VY�2*���6��s��3�t���+�C�����R߱��=f�E�!�D���X����dM���i��<��
�o��@H��_��8���NdP?�(�*?�)��FJ��qd�h)䖱(ǀ$���/w�=�5
=�B�}�+k"��)���zVʁ���8{0���[��0�e1�:p:��k��wv�m��#�0'	t��ƚ�M9l��s��������٢�=DI�d��c$bV����vs���,��ч��;W�ph������/�uH#ew`�S�����tar�G����7��Z�k�#�O��GXo�A��[���C^���)	yak��z��Y_��0@�˽ז$ �ʍ:O7�Y/8��6��	`=�Ӯ���gP-����)1$.�����%b*��#\���=o���B�m�������]꛺�-<��-��90�/�&���cP�ZOO����3�2k�{S��K��C�8QJD�?p��t,}`�*��\^��9������LC��O�"8�PLm�b�L��*��싸�����͖��7�)�a���Z�$ĸ�M�(l����^"8�Q1�%)���7_,r����)�t����=�q���+��"#�I��{�a�d6j�g�%��w�T�#��f0�>��)^��S�1�EI���3���sA�
ڄ�I=^. ns�~:w�*"�0��I:+i ,�]��:ܜ%�`���^�8���l
��K�[o���bH���	���/pp�X�`6y!�"r��z�\d����Q�ԉ�����z'�P?e<����ص�XB���hE+�u&����K�a,�K5�b����<=9�*0u����yeM���z�tԴ��&��XY�F]d(�7�ӈ�2������5�]��P�0�#DX�Ε�`�w��t]�tRs'���L�X���)�`&�0���#�Uc��	 u��3ة���4u�0i`�#'�(N�C#ئw�$���|�5����L�\a�Ǐ�'��U��TsspJ��'&��nu����%s�G�:u�'�Mp���.��kWi,�W�����qUH6��k���~xte5�ھ���(�^
����(%�l��6S�/q������$]�(ګSa�+�Iݩ{6��rr�����_$��k�֟d ����|�E���|{����т�Avz�!�� �C�� /)��	���џI|y�k�,Ď��:�eM�sU��12,�B3/�¡;��$��0�*+We����|/j����_yf�$iV>��$��������p�9�z�w�s�ht���4˔�/C;�&����O����(�����x�k�U�ύK�C�k���hBj����c����sO׎"ѹf�L�Z����]$���Z���7�Ǧ-�����+@��&���h|Sf㞄���f�gp�[������F�ڱ%hF��q���U��{K<��/L?N��Cr=e����,�>�O�VPS���ڠ�r` $�Բ��T�:�r��ͤ��NیoX�<�a��̪��<;����F{��G���0~�S�/[���^�מ��ާ|k�-��z��ӝ�.�����{�-�v��+�����e��!��j��,��ծ�x�1�~���k�-D�+�dv��(bp��tz���ReWKf�@��[FEa<��s��R�~��_�H�u��_k'�`���Uk^�f��t����
�;d�%t��?����lel��D��Ϲ�B�����θ�w�M�*zXf�?߈䙄���dQQ�� 3ܬw�Y\�sE5e�gX�i$ ��A��x��,)F�zC���ʴ+Go�p�3�!�i�@-� ˨�H4�s�/�����m�'-��G.���^�	�#İ�9�YI}?Pv��VJ��D.e�^ ��ҮX�L�ء��� Z���@���Л��u�����3L�|H�;!��^���s~^+
��5�^b�Ajܲ�!y����7>G�]5�;įN�d�@O���oH���j��	��'�i/���x�`����éO`��S;7�)�2����x���v�gԼj�0��y�-�̯K�E�c�UyI+���ۿ��K�cԤN����섏E�Ni1�H�%��a��|��<�"b&���C�������f�>��	��Cv�0ʑ,;����h��((�>$!�?
����u�:�>��4��z,�U@Q�	��*����3�ŮZ)��m>ߠ��<���w�y�A�ks��)n�y G���N���a��)/��|���y-�"?���꩎^n3��w��7k��7tW�y"�y�0��''�3���T� W�>���M����B�B����>+s�ը���O��H��ЈW���jE�>�u�Ҟ��%`�+|d������l6wWl�;��	�
��� U��F� .Q"��(9�w�jC�S���p��*�G@������^혊m�#7��CjH��_p�gs%ɤ�mFN�&��'�l�?���t)�bf_j�+���9�\03;z;8v�8Hhp�)D����'��)�U�q.���+=�$nS�$��&Q�A�j�T����W��ӎ��3D��R�X8�폥�"�j�k�תHSo?6Eb�(P�I���GЫ���jp`�Q�_���m{�wB1�IX\�n}�W�F��r#�*�+�ϖ�'ݎ����b!�b]7$	C�\�v�p��&4jR��kʭ������+<���B��/�/f�`�ʡ�텅�c�O�#Z�P[m��hK'���+��D-;n
�M��������n{>�9p8м\U��H��Y�f 0	ID�ӈ�XfBn�^��\p�Ǒ�a	<U�4���}��$����	��J �X�5�y��w��iA���f���{R=�Y����^�d�I�6Ս
�,��"EJ���;*L]�r��=��K����B8g�o�g���j��I�q[W��.���֑*;���Q.0c,�� �E2�(��76$��� ��o?��ނ�i5��!���?���<ܦ�O��8��*l���!	n��\坓6k�p4P����&k������
��Y�.�� s�CW�/�1����*�6(�na���B.�]�"���N/��8��b[C^��֞���y�c&���jf�D�8NeӜ���<*��	�����Ş��4x�͇�ļ��v��z� �*B��y6y�������ʥjrV��k27^�� �ɵ�h���9�O��s�rQ�h'��欨����U�C��2�zd��,#X��}�a� z��=,/є,�dח��uP����B�ڟ��I�&������Δٲf;�.�j�Ҁ��t�����[d�{���L��K�
Գ�,���Y�R��`�=��ߐ`��p=!�?8�,���[�?7N]稾��C���]�P�2�\E֘w�@"�m�]d7П��Q��Pk�RL��v07��.�.��|�Ü�Ɗ��b�v2a'h!5�T!���Vk���e�/I��~��y��S�����a���50��������9�Wi7�^���i��4Ⱦ�1Ch���Ђ�P�jB?ĕ1O(`s�W��)~��s`����g�k����mb���z�$�c�o%��Uj 7�����ئ�U*b }`�/�Ӂ4�8M.2�4�����	�J��X�*gD� �m�u��W��xI��lS�fP��P�� 1�-�ׇP6�)�u
;P��ߢ-w�{Z��Y	I�ux��U�k|r-tw�'G�[���[_^e1r�ߟF�c����$��[_$IU0~�Y���z��;#g_ÑZ�l���5%,�8�(F�_0v���q��PLpfxbkQ��>g��0��"4e2���W$���M�c\�
p�֧j:�c`@TEKpP�aɹ\s�]����ݮ�>.�_�|@1G�B����/�����"�<� �У�D���c�-��E�`�p'm�/�dC�h���hZ� ����m�v���wMZ��d3�⮆(iH�p�AQ����s�+��!6A`Xh*%X��RI[�&d�����cƂ�r���l�؂�[�����0��׬��������{t�> �s�p��<�����0����Ў*�>�3�j��P�9��YCߵT�k��T�b[S��4��I��گ�\�w���*������3�89���@q��T}i�	�[g��,�V�����v�:�H��<ԇ��`��ߖ;I����@%�9� lyNg�4]&t�=k�V?�I�tb-�ψ�򝒼�%tg"42�\X�ɜR1z���<R�j �n����[��b�����(Ix&���BϦ��>h���4sʝ�|����$ܩ	Ex�]�Z���~��R2x��"�Jn�8E�o��x
�%Ζ�c�gG�2�bW�{�$ p1�{��[TS)�����yO�Q\�ֆ��)��^t �_��I��XUwR�E|k&y�ܴ��WAS��C���xJ��Rn��u���!|+=�2���+��o�͊�-���.3��^Z6�!"!G����J���Ԓ*��w.���ꍪ�BtK.�M��OU�uH.����Q�o��O�����>R|��T�Zv�쌽��Z�e��7s_l_�)����U�����H֤�����^/(�[D�>*���4�/~5:
jӰk'������Lm�v�� 93�3�r�$"g,���(���PJ_��/)�<�m(e�Z~�0�p�WC��L� mΫ~8TT�+��|%��3���i٠����K�S�~|N����|��_��3E:c(�z������RL��5�vA=�.H쏢N�*K�s,d�T�����.�׫�\�Ar�/l�,i
x���{w٨\�[A��'�wɍ�,Q�K���2�Ҙ���jg��C%��4l���0�l�JwT�1��Nܯ�c���|���Q���f�M�q����E%�A�L���v�m��O�p�go���tX�\$�i�Vx4)Y�R��b.�Aٗ�)���.��z�wЎ�@V4G7fދ'��g'*^��c.Q�X���>���=�Ŗ$~���B<�ߵ�E�q�R��������pZ\:RY)�S�4��&��<(�-1]d��Q�-,�[Eg�/�ܥ�BwY�޶f���C��w蓶�"�I8���ށ�q��Wƍư�t�\��oY��_��O	݇4o&h�	��4f��{㱖�b��\0�������b*q����@2[sj$+�l��9���d] �=S��js�J�p��j�Q�y}O^���MR4zƓ�j�&~�ݑ��z�ʹ�rJ�@���r���X'���?���>A[��݃[������H��o�o�p���1�} �T$�{��<)7YE��I�[�����2N��C�cʡ�x]`��h���=�$���2	k+��A�HPAQ�>caA.�#��i�kh"�˥?�K��_m�iAqeo^�Ŝ\��(I�b,�����b5�\5�aۭW�@����-��}k{	.����+�s�i2�I
��|1X#�E����	cT#s"���9A��M�[5�p\ԁi Xj��Ӿf�>h:�0jT	�$��b���
��z�4
Z/8�H�)X��aF��~w��F�@���o�$��NMHk)�vQ����N��� �����:�%�#y�G�*��V�Lx�h{�f�tf�Wi�|,_9C�g���Li{5z�|��yC�ae �ar�M�-e_� �� ��ɱ��,*��Փ�-b�->�ُ��d�C��Tb��DF�߀�E�I������?i��ko����DvkVˁi6U��A��yy�����#���J���.�*�tA҈��^������e��)�(��x�8���q�r($��`��y�?@'Z�R�j����֢F'�6�r.G]o��ݾL���g���Iۭ��n�ŀ�/�j�/�)��U*��VJ��	4A��Q�w*�^6�@�_�ɍ<Ì$�y�+e��(#�|���M�
T�"[�_������	 EQ��DW���5�������J0�i�f~Ic�k�:�,�-ᬉծ�4I��1�\z��BD�0�k�^�������O7�Y�l��٨Fcv��оy�T����ʪ�W7���z��%o��ȣ^ă�f�j��Q�����H��։ӵ�� b�e�#G:���R���ɲ�7(���j�;ែ�"�4�sTQ�?��T�*��W����o���D��1�w\�T�*씁��󃺼%@2��;~%����n�`Jc�?9[����wM�f+�K^��**p���-��rQ��Z���������I��؃,p��2��w�Ʀ(�P8�J|^�+��L`�7�炱�[q�'oN�ȋ{�GȒ��-�&h���o�2x�β�F]c�!p�8 Qoh�����$����?�n}֚cUq�x��~�sO���	#�E���%�O)>�)D�KD�[y�$=����؊d�H8�>�𽪺��>�ʡ%ĳ���J�M0���Ta>y�f�b�f�����'�PLE��ê@��JI�4Cb�x�#�7��'* �V}��)���wUF���So���r�#�?W��@%N��� �*n5�J\Xs���)�>�,!�$��e��UD��Š�A��/J����A+�����߭`�������v���)�v�� ��f)�#�xû�DYs r�x�k�v�_����/!��Y��5z��#:��@M�y��-�}�;�e���*Ys���^./(�3�2�Dm[܊^ꖅ�@*K(�\��0B������L�VX�姚�ڛ�"7�.�U����"�M�c���QӠ��7O�`�Ŏ�YA{�npz�l�	��#i���q2\��M�S�5tmD�?���G=*H��Fs�h-�MA�:c.��E>��A`l����Ve#4�j B
�|F,�
�I�kt�Ս�S�t2R�O7Z�bF�9�1���q�Y�c�3Z;�ÇG���7M��>��iRk��tȴ!�={5�l�h�k���LI��Hq���|�� �������=�J,e�pX�O\��xc��s>ts�aT�J)����@	��ۇ�Q��3P�G��@����g�F����7�����/�<�`��d��ݐ!������U��(��s��bn~�ٗ����t�2�$��PuVƅ��Xsl�/t��^�X�L^��ށ Y;m�GH��ai��0 �a@q�T��� ���O�����Qq�H�ͷHW
�� ��?(uY4U\2&�Bl3C3?�wr��-8`�<�dKuQ��\��.�	ǀ/��G<��!0E�t���eCJ��_������#;����t[��΢�JT�ve�M%*�X��%��&��`��� ��UP, e�5 _mf1=>7�5���Z4�ߟrS^o�Q�ڔl�jM���tn�B��w�V�a��߁��X��+lLM�m�+��ͽ[t�w���������%�U�(R�v����Ӆ��ɹ�����u�$�ȗ�:Ø� v7�RkW3ɓʗ�Mqh��xuU4V?'�b��w�c���|�V�5�u�8�U���	��4�&��8��NW�}����Y���3�>M��;C��vJ�s��J��7K�"]����V����|�����7��$�&Ks�i>�E�����lF�7G}�5e��4�ĝ*b�Z�J��N#J������23K�έ3F�P�IHJ��G�"�rڼ��q�v/�V��#�w2����A�R���L+6er���(O۞;Q�m[��>�]2�5@;٨��G�x����d�q�'��_��w�V�W��"	�ؔ\|c���nP� ���ȀA�����[��;޶��F��M�r=!�7l�NilQ��Rg�����������Q���K@9f��{�XR��&.B3i\I�*��z?LE�L�]E�?wñc*O��&w}�t҉\�X�Cr�؂8Ti�<1�KN��a_�
)s����h?Z����F >~|��j��6h�m�����^e�&.�Qs��X>�}$˹��5kq�7<�GD)�W�Q����ۄTo(x讕At5
��N����bk�����i�6Ǡ;D(��QWDj%=��x�m�bvnw�c�na��	��j[�n {r'��h�^p~��?��?�4�E���X���Z��F���򵴐��v��7A������������������].�9���0D�!��;����NFs,��{-�0ٸ���R��(1���܍%6u��b��9έ��"��;��ԑ[��cG���N��y��ݯ�{dݏ.1��v~�'2�Y:�#��a�k�DM	d1��._C���&�3�����1�����x� TfJ��L��;`p Je*ЇŚ�|?��%�W���y3α��j6��\
��|�xg�&� J���bs�?�e�y��-���ٻ�GݪT�¯̠~��%�O��:�`��5u�s�P�t��EH�����ò$���H��n��Gx�S"Nb$z;�X+Sx6��H�!B:��8�w)�1n��5�ѕs�O?���<}�!�T��.�@RVMYMy8j����A��1�u�>�!�V3�QU��u_P+�e�x�DVk�1�)U�wdj�v�;�f��I ��X���ȝF�b��+F������r��R�O��|0�|G����#��&�rD�U9�$؜4��Q8M�
�q�/m���]�C��t"�]�'D?��l���j�?��+�L	5�~W^���ҲT����/N\EaL�nE�[�������v�T�pC+�2�3���a��//�Ulx�`�֙d�C �G��JѮ�eU�R�OڲY�\p��]q�?f�*`t���"<T�gOd�A;Y5?����2àK��JZ/p�Xsl+b��u�	q�4�
A��6�>P�'�R8�ޓz))�1d!>`V���gZC��{���-��o������́
83�u����?LuajS	��bxw�E>��9�SG�Y+�2�(Y�47H�~���iwCܚm�Ҕ�I�!�Ȣ{{�#*,Jx��[�ݑb-���X	:��9�����ySha��n�bI�h�W��tg#*�� 5tơ��He�a7ӹ쟠]) Q9L^'�a�c%��%� ��D~��Tų9�?�"'�2�G��ω�#�Y7��3�)Ɋ�pY)7�7��+E�yI1���7�;�����N���dj��%נѝ�Q�[ K=8�
�Dz����q��|���\�J| �Ί�Ҿ|=K���}B��y�^N[��y�;V��Z���O���+=��z{�~���o`�W������1��uS�՝ٕ�J~��k�Q�t�с�I�UK��� �%�ԩ8�V�u�x�K�����hSh>ͮЙn`Ih
Tx����hNiA"MC��}�c�P!7t����Yp��؛qGPCz��� J�.~Q��OLE|5��y����-��vj(��]H�I(�煸��h�#M�j̘�S �x�(��P��Լ6�k�Lc����:u栊��ؽJs�]�W�{���<Mܑ�qH(�R�ZO�`��^LQ� �`��'��m�	�fV�ҽ����?U|�Vj��������␊��](��L6���{7�ߜ�*�p�pMH��a�{ը.F���~�N�B������^D�h���fZ��ܼ?Q [��f� [�^E�dh��Pini%ǝ2pgh�L���H�^u,V!ɡ�GZn�Νwc�_�i�y�ꐬ��c��|9w��eC+ԥU��$-rrU�]g���#6(R�@,J"ĵ4��][����]_��
���XM*㪟�ΠȲ��	�c�<�;����'S�=5�����w�M�!�=�}�8�S7V����	��t����,�4�K���x�)�$/H��)K��!:�h���2Q�Sp��Y� ^ ���e}�63g���6�j����f��Y���\#V��V�-F}�X�.�P�v�P ��ɑ�� ,=:��%�y�h^��q��#��lg�\�4��r�_����F˓/��5�r=��bK��g��6�z���5����%	T�k���i����Ɣ|m;��r�$����ԟ]^5�m�Nɛ( q���p�r���`!�>���˙:�]��D��V���s���5�&1���"�/���G�A�=|�8o2��� uE�a���*���i��4�f��&������쇶ޏ�Y_c���!������s�1Ȑs��\��z��R��LjR�9ί��~����c� �~J��X�K(������O��x���/�R]�+��so�}��C~�҄�iqbh��cr����+q�՗��,�G��h�>��8k��������^]���N~>&"�
��0�mS<")GJ!�9��N����9cJK�h��(*@��
3��#���"��zʗ�c�a~�oQV���H��/E�`��T'�o!�1��5y��l���-(���x�Tԛb�V�thI�����C)d_�!.,���L���p�)���"��/T{N�7�ql�b�/�*w�
;����b�i0�Y֟$ௗ�i��?$!��o����,�?Yz���c�X��o$i��Q��(%��W	2o����Ci�W�����2(�Z�o��1����n..�� 7
�:�
�����Q��j��P?o㎷-�8�R]00���$��f�lͥ��=�umƌ2'6Ja���X��[N��0�0GG�r|!ڄ Nԅ�Up��k�Y6����7�7���'�+4��P�u���-6�����A�>�a&V�C[�i����	��p��R�ۻ3K^2 �!_�:�h|.Ω�t��.����K��"B��X�\q���E��y������A�7K�@��s�4�e+����1i���t�^!�D���49-8�T���H����%c6K�����,ZWu� ����f�C䧉�q�mV�v^�(��w)\5i���~�t7��H8Y~����GR�k�L���A������A�Y�q&�k�o�{Z���±�O�?t���ҿ�j�ߩ�f��z��)Р�z��8�G��u_����l������Ô{SE�d�>F�{���gy�"�s��rA��{�
Q=B2��FY���=ŝ�*����|L}��� ����G$��ܮm����"��p�1{M�&	��~��!��[�� g�ݭJc/��w�|�Ii���4)�SQ���ԲӮw�K��sH��*����.��ۓI �����Ɵ�Q�vom2>�5�p�|�)
��@����B~�ȳ7�q����A-mD����]I�J��%G���A�נ):��t��\�y��ve��ȀDP��:�^T��C쮷y<+Z�I�n����d��ۻ��c��csJsdx�$�Ԝ��y������2���;��C��t��W˖��BF������*����0�Z�4t��D2ꑂ�(5�TC@���}���+:��XWetZ���`��n6 ���W�Q�K�s+1i5��pY�]ۯ�W`�=� d
�1�ԇ���Z=5Z���\�yU�fSv�U<7��|<~����ݹNV��0���u73�V�$�=.hM5T�V򽃧8�����q�O�b�n�3,��h	�ao��^�m�#8��f���OO,�����t�Ŷ�;#��X;?�<�r�@ה�B�R�_�8x멜A	Ȧ<WN��V�:�y��d�A�2q�X!&HY$>D�#h���S?��Y(�3��>b�<�� VG��A��:8��z�@��~	p�Z�Z|�I^R�m�t�����Kί����F/i�c���`F��7X����������]�M��X�$����Dfw��?�-9��;N�f^�ZJ��_��_� F��=W�JO�S�J4���z�Ѵ�N���_x��]�5���z�#]I��Zw���0�en���)������Ar��_'!�j��r�NR�A�n��C�o��\�i��4v�$\$� �Q�:�1!���ܴ1��ɰ��H��qG���֙��ȸ/�W�����7}th���^�߼;��:=�_�s�"L���?r���~��#)2b��a��"�.���F]o,��I�J<�u:�(��e���So��|$iܡ�t�uH�B�I.�7�;8�g&�?����K&�P2@���U�"c�=����sGٓ�=1�oZ$����r���%����}Jɟ�b�vN�Zin.���4�^�]��PAMO޾ 1�Ԣ=)(R��S�����Qt��[��ig	d�x�Ǳ\�a���Ď��~Wjˈ_���SK�Ώ���!��T,+��.� R"�v3��4�(�O���C�q"ٺr�O��`�¾n�2��|N�{�B�``�+�yݝ1�g�Gz*B�k���L�q'�1��>�۹�s��x�nM�Ӈ�k��Ͼ,�w�-�|��ՐO!���A�Ъ���B��y��!k6�����
���`2����W@ێ?�\��堂�A�RtF>=c����T�u��F�\mx&��.�5���܇��=i�N�t��4Y&�8Qݐ8��yA�=����C�IQ��<[�.U��}�;F���b�&k&�מ��i2'/H���Ǵ;����H���v�&M��
�Cx�r����Nd���O��-�^\�;�oV������ĔZ�V�D<�Z�����j��7T�f[Y\��C���lA�͇������a � ���cF�9�U��βtMe��
˒G)�Ο?�=�p�?�}y]�A�B��
�^���Գ������*�r"����Ѹ��0Q��Z�a܏�@ �x��2���HIҌ��U]�E06����u�d�����4�Q�ל��e��f��Îb˂�b���ZWu��ŘwB��Ȥa�v&9m-	i��c�p���4��!,y�lw�j ��NB��i[�[�K�jo�������K{U"�z�Ŧ�N�>9[�.&u�&��Bˑ���+�-����B���o1ǦA�n���&����òh5�O�x����7��4`�p|���)���gu*�H�5�XsS��d��D��ް#�D�Q�m�����-o��CA
�#K���3���������(�MWl�����f�����Ϩ�����{F�':�$G�f�ػ'�����d�G0��0�� �.R����wL�)��Q��j���G���l��}�6����=�Y��n�dD�NY���ZP�1�m��{�#���j�T;{e͋s>!G�{o��?���EX��4�-�
�Q���k�����Y{�R�Ia�a޴����J�ʹ�w*�k�W��(�2
q�P��wyW�#A�K��b��LWܒ�|���T����<�FE�fy��P	�x4�����$�i}
��R.�F�b��r��F�U�LH�Gǁ��&����V�;���&m���� �o�Y&a�5[�����gt��P�d�E`�%
ק`"'!�{Q�@�,��`O����n��a�Z�֊��
Y|}�c�� Տ2�p?#�[`(����`��T��gQ��"wQ*Qe����;~�8��@0�{]8Y@V$��3�E�(v�d�3�?w�r��+��h��O�i�gtI^e���J��4�dT�"����5�FN��o��$ WT�>��đ4���KT�t�r5f�at�:��Ԏ>�L��V��H���N1uF���a�W�^�?ڶNgv�XD	a�L�8�υ�����??o�����sھ�6�����N��+�|�D�C0��R)�u3�40����a�y|�`�Xf��p`���0'˦P���n��XZ���xFIk�M���� M�x�����Fgn͓�$�@~O=��R� hb(^��4GM��P��IJ�RW!`%gsfS�z/xj��������@�ѩ0ྑ"/�<�⋿Z��+��ЧI(q�Ik����mVwM-��!�������^1#���X �E�^��xq4ܕ��FDů�')���ӂ�f0t��x�� 8W��z�|a��ي?�W����ݨ�n������0��BuZْ,cܿN-�qR&r^b^��8����;'�6�tx�=x1�E�_�)�v�K���?���W>��"�i��|���c��u�/9�^=k�C[�4��+BHcz�s0�q0�~@���^-����.K��~���W�kR���#��_���|8�g�g�ΐT>�K�l7\*�=�(}��̅��.'�x���Ե�����S�-�q;��@]S�!����֙p
F�z��I�i��v�vu�l�`�%5[���DsVv!_��P�b��N�nS*=.u��X?n#���Y�G�c�6�$
����z}���=,�}{xUZm�i������`�lCx:]��7T�����{U���n{@
�c��G���X"����t홼��O-h�ނ���y�>x0'`�'�o�C���Z�P�y��w̬�B���3��K���no����t�e�5�⚃0A�r,�;{D'���`����+�8U���?V�3�P�R�Q�TRD�fjy��g5m���B�L��׏H�Y��c�nW�{�B����+#��!ta�J�_Q���ӟ�a�	
B�<�j͠S��6&��}i�̀v�I�c�����;��9E�'��.*� c�V.�U:�Q ��ۇe�5��\���f
���a��_y��������
r^ ��$�m�"�Ey1�l/�P�uD����[j�PK����/�e�1��L �A���k���� �}g�Py�8���5��+�^�Jq�_��)�\�  �f!,�!O�V#�w���?|eJ�*��%?�?+����f	(��~V�i�=�!L�=�鋷F�k�bЬam��4��j�R��9��!���z�nj��!��
z��A7�r#ܨ�wX�:�]��\��q����{(�uܶeG+�u��|hD����a����I>{��V��I�_R�DXKdk yŠ
'�.��0���0QU��ͪ�D3�"�hT <�~E�K_h�_Ԋg�ld���`�p1mD/��A�谌�`eF�#?{]�^"��#�6����LR�yo�C�o��=Q:�E�� ��K�L�)�>�*53���um��%\Ꚋ��x��@�@<(��}��@HW���v Q�)S��8�Wţ��I�*N}���I�4��5�܂[l��RR�\P���f��$���[ _�`p�vd��9��Ǡ'!��HkT�L�ՙ=��[��Ъ��_�(!�'�~�h�cUgt��]!~��I�Q�`�Ӑ��.G;z��&#^ȹ�Vi6���Q�n���/[�-�?�[3����~����%n��\y�G��H-΂�x�XA�h���U�7��{��y.g+ī��%�C�y�%"�H���{��@I;0�>�ŜV��:��s��N�Q��㮹�'��)�\�                                                                                                                                                                                                                                                                                