MZ�       ��  �       @                                   �   � �	�!�L�!This program cannot be run in DOS mode.
$       }��9�l�9�l�9�l�9�l�8�l�9�m��l�`��:�l�ű~�8�l�юg�*�l�Rich9�l�                        PE  L ABdH        �     �8      8  �                              Q  �  �                                �F  (                           @J  8                                                  �  �                           .text   �  �  �  �                 h.data   �1     �1                 @  �INIT    `  �F  `  �F                 �.reloc  �  @J  �  @J              @  B                �G  �G  �G  �G  �G  H  H  &H  >H  HH  fH  tH  ~H  �H  �H  �H  �H  �H  �H  I  I  I  (I  :I  HI  dI  tI  �I  �I  �I  �I  �I  �I  �I  J  J          ����� �             U���<SVW3�vw
�IZ�4(H���u�5� �E�P��QRZY�E��E�   �}��E�@  �Ẻ}ԉ}�v
wt���Z�7��E�P�E�jP�� ����   fP��%fX�E�h� P���
   7E�X��c�$��u�E�P�� �E�jP�E�P�� ��|3SU][�E�P�E��u�jWP�u��� ��|j_fS��f[�E�P�� fP�QfX�u��� �   ��$Ë�_^[�� U��� SVWfS���f[�   �   4RCr���E�E�}�s�   v
wt���Z�7��E��u�   fP��%fX�E�P�u��� ��t�tfQfY�=�F  w�ePS[X�E��F �E�j�u��E�P�� ���e� fS��f[�E�P�`  ��u�*j h j j j j �E�P�� ��u	�u��� QRZY_^[�� �% w s \ % w s % w s   U���8SVW~bF8���A(b�E�h� P�� fUf�ڠf]3ۍE��E�   �]��E�@  �EЉ]؉]�fPf� fX�E�P�E�h?  P�� ���   ��$�;���  �5� �Ddk Wh   j�]�]���;ÉE��\  fPf� fX�   WSj��WSj�E��֋��}�~bF8���A(b�}� ��   ����   �5� fS��f[�}�]蹀   3��E�Ph   Sj �u��u��� ����   fP��%fX�}���h2 Sh� h h   �   �u�3���� ���u���  fQfY�}�h� �u��   3���� h �u���S�u���h� �u��փ� W���  _�u�u��O���~bF8���A(b�E��(����u�5� ���u��%P�   X�}� �5� t�u���fUf� f]��tW���u����u��� SU][jX_^[�� �U���  SVW�} u2��  ~
Rv�~:��j ������Pj j j �u�� ��t2��t  PV^Xfǅ������������E��E�f�  �E�f������f�H������ PS[X������P������P�u��������  �������������� ������ |������9�����u2���   �E�f������f�HrsB����5�X:e�������  v2��   ~
Rv�~:��f������ ��   3��������f��������E��p�����������ȃ��P�   Xh� ������P�  ��u2��ZfUf�ڠf]��  �E�~
Rv�~:��h: �u���   ��t2��)�   �   S���hT �u��   ��t2���_^[�� ̋D$���t���@��� ̋D$f�f��t
��f�@@��� �SVWfS���f[fP��%fXfS��f[�\ �6���������� |�~bF8���A(bW���  _�� �6�|�������� |�P�   X_^[�U��QSVW�
   �   ��2�} t�} t
�E� ��u3��`fUf�ڠf]�u�� Y�E��
   �   ��I�E� ��t(�u��u�u�� ����u�E��u�	  �E��W���  _3�_^[�� ��������������\   %   %   U���XSVW�e� v
wt���Z�7�hDdk h   j�� �E�}� u3���  vw
�IZ�4(H���   3��}���u�u��� YYhP
 �u��� YYh� �u��� YY~bF8���A(b�u�E�P�� �E�   �e� �E�@  �EĉE؃e� �e� PV^X�E�Pj�E�Pj �E�Ph?  �E�P�� �E��}� }�u��� 3��  �   �   4RCr���}���   �e� �e� v
wt���Z�7�h� �E�P�� hDdk h   j�� �E��}� u�u��� �u��� 3��  PV^X�E�Ph   �u�j�E�P�u��� �E��}� |Kh �E���P�� YY��t3�
   �   ��I�u��� �u��� �u��� jX�$  fP��%fX�u��� �e� �e� �
   7E�X��c�$�hDdk h   j�� �Ẽ}� ��   PV^X�   3��}��hT
 �u��� YYh� �u��� YYhX
 �u��� YYh� �u��� YY�u̍E�P�� h� �E�P�� �   ��$��E�P�u�jj �E�P�u��� �E��}� |fP��%fX�E�   �u��� fQfY�u��� �
   �   ��2��u��� �E�_^[�� U��QSVfS��f[j h�F h�F h�F �~  ��E�P��  �� �� �Q�0����F �I� ��� �u��   ��   ��$�^�[���U��SVW�   �   S���P�E"�XP�   X_^[]� U��fPf� fX�M2҃a �a �� 3�]� U��QQ�u�E�P�� �E�P�� �� I o C r e a t e D e v i c e     I o C r e a t e S y m b o l i c L i n k     P s S e t C r e a t e P r o c e s s N o t i f y R o u t i n e   S�   ��$�hH �>�����F P�   Xhh �(���h� ��F �����=�F  ��F t�=�F  t��t
fS��f[�[�2�[�U���SVWvw
�IZ�4(H��������{�������u
�  ���   W���  _hl �E�P�� PS[X�E�Pjj h �  �E�Pj�u��F �E�}� }
�  ��   �   ��$�h� �E�P�� rsB����5�X:e�E�P�E�P��F �E�}� }�  ��gfQfY�E�@8 �E�@@ �E�@p W���  _�A   ��F fUf� f]�/���fUf� f]j h: ��F �
   �   ��2�3�_^[�� �U��j�h h d�    Pd�%    ��SVW�e�fQfY�� �E�fUf�ڠf]�e� �e� �$ �U��� 0  }8V^�����3����IQ�E��RS�� ����u	�M���E���E���jXËe�M��fS��f[3��M�d�    _^[��U��fPf� fX�   fUf� f]h, ����~bF8���A(b]� �U��SSU][h �u�  Y��YujX�
fUf� f]3�[]� U��QQRZYP ��E�%����"�XQ�u   Y�E�M��~bF8���A(b�� 

 U���<SVWV^h� �E�P�� �
   �   ��I�E�   �e� �E�@  �E��E��e� �e� SU][�e� j j j`jjh�   j �E�P�E�Ph  �E�P�� �E��
   �   ��2�}� |�}� }3��k  fUf�ڠf]hDdk h �  j �� �Ẽ}� ��   v
wt���Z�7�� 0  3��}���   �   S����e� ��E�@�Eā}�5  s`fUf�ڠf]�Eċ<��A �Ũ��3����+����ً����3��O�����˃���
   �   ��2� �}̃��3��O���fP��%fXj j h �  �u̍E�Pj j j �u�� �E��u��� �u��� P�   X�e� �e� j j j@jjh�   j �E�P�E�Ph   ��E�P�� �E�3��������~bF8���A(b�}� t	�u��� QRZYjX_^[���U��WW���  _�Ef�8 t@@_]� �U��QQS�
   7E�X��c�$�� ��tXv
wt���Z�7��E�h� P�� ~
Rv�~:��E�jP�u� ��ufS��f[�u�������t3��,fUf� f]~
Rv�~:���u�u�u�u�u�u��F [�� �U��SWW���  _�� ��fUf�ڠf]��tU���tPfP��%fX�=�F r@�=�F w7QY�=�F u�=�F s�°  ��   SU][�
P�   X�A�@D�3�_[]���%� �%� �%�           SSYS32     www.6700.cn/?b                  �           � � � � � : T l � �   2 � � � �  $  + P u � � � �  3 Q p � � � �  ) L n � � � �   %  C  _  z  �  �  �  �  "! D! _! ! �! �! �! �! " H" l" �" �" �" �" # '# O# n# �# �# �# �# $ 3$ Q$ s$ �$ �$ �$ �$ % 1% V% u% �% �% �% �% & /& Q& r& �& �& �& �& ' ;' X' u' �' �' �' �' �' %( E( e( �( �( �( �( ) D) _) }) �) �) �) * !* @* e* �* �* �* �* + '+ E+ f+ �+ �+ �+ �+ �+ , 2, L, g, �, �, �, �, �, - 2- L- j- �- �- �- �- �- . 6. P. j. �. �. �. �. �. / 2/ N/ f/ �/ �/ �/ �/ �/ 0 50 R0 m0 �0 �0 �0 �0 �0 1 51 T1 o1 �1 �1 �1 �1 �1 2 62 O2 l2 �2 �2 �2 �2 �2 3 53 T3 t3 �3 �3 �3 �3 4 %4 @4 [4 z4 �4 �4 �4 �4 
5 $5 B5 \5 }5 �5 �5 �5 �5 6 /6 I6 g6 �6 �6 �6 �6 �6 7 77 Q7 j7 �7 �7 �7 �7 �7 8 ;8 V8 s8 �8 �8 �8 �8 �8 9 09 O9 r9 �9 �9 �9 �9 �9 : : 6: O: i: �: �: �: �: �: ; -; M; m; �; �; �; < '< M< s< �< �< �< = 2= X= ~= �= �= �= > <> b> �> �> �> �> �> ? 7? U? o? �? �? �? �? �? @ 2@ P@ j@ �@ �@ �@ �@ A A *A @A XA sA �A �A �A 2 W a O P Z S   A b O ` b  > O U S   J ` S U W a b ` g J c a S `   J ` S U W a b ` g J c a S ` J   J A ] T b e O ` S J ; W Q ` ] a ] T b J 7 \ b S ` \ S b  3 f ^ Z ] ` S ` J ; O W \   7 3 F > : = @ 3  3 F 3   7 < 3 B 1 > :  1 > :   J 2 S d W Q S J : ] Q O Z A g a b S [ F   J 2 ] a 2 S d W Q S a J : ] Q O Z A g a b S [ F   J A g a b S [ @ ] ] b J a g a b S [ !   J R ` W d S ` a J S b Q J V ] a b a   J   J A g a b S [ @ ] ] b   J A ] T b e O ` S J ; W Q ` ] a ] T b J E W \ R ] e a J 1 c ` ` S \ b D S ` a W ] \ J > ] Z W Q W S a J 3 f ^ Z ] ` S `   @ c \   A g a b S [ 1 V S Q Y   J a g a b S [ !   J a g a Q V Y  S f S   A g a b S [ @ ] ] b   agaQVYSfS caS`W\WbSfS AgabS[   !&#ac`dSg&&OZZgSaQ][   !&#ORbO]PO]OZZgSaQ][   !&#Q]RS_WV]]Q][   !&#c\W]\[]^Q][   !&#XaYYc\W]\Q][   !&#dYYc\W]\Q][   !&#d Q\Q][   !&#W^Zca[aOZZgSaQ][   !&#[[ab b Q][   !&#Wd`R]PWU\Sb   !&#eeec&cQ][   !&#cc&cQ][   !&#W[UhVO\UfWcQ][   !&#bZZW\Yb]\SQ][   !&#QVO\\SZS%&Q][   !&#c%b]e\Q][   !&#c\W]\'#]ZQ][Q\   !&#[[a'#]ZQ][Q\   !&#[Ta'#]ZQ][Q\   !&#bZO&Q][   !&#ORO&Q][   !&#c QOWYcQ][   !&#[[aQOWYcQ][   !&#Q]RSQOWYcQ][   !&#^cPZSZSQ][   !&#cZSZSQ][   !&#%b]e\Q][   !&#bdaS\R%b]e\Q][   !&#Wd`aS\R%b]e\Q][   !&#bZb%b]e\Q][   !&#UaS\R%b]e\Q][   !&#a[aaS\R%b]e\Q][   !&#[[aaS\R[]gcQ][   !&#'Wd`Q][   !&#[gOR'Wd`Q][   !&#c'Wd`Q][   !&#c\W]\'Wd`Q][   !&#Q[^"^Q\gOV]]Q][   !&#c\ $#Q][   !&#c\W]\__Q][   !&#dWSeOZWc\W]\Q\gOV]]Q][   !&#c\W]\\O``]eORQ][   !&#Z\VSW[O&Q][   !&#eeeTP]ObQ\   !&#Q^`]POWRcQ][   !&#c\abObPOWRcQ][   !&#gQ\fORQ][   !&#eeeSe]e]Q][   !&#bS[^ZObSc\W]\$!Q][   !&#\SeWa$&$Q][   !&#Q`SObWdSc\W]\agaP]ZOOQ][   !&#eee_gcZSQ][   !&#''SQQ   !&#eee'Wd`Q][   !&#[UcYOYOQ][   !&#Y]]f]] OR"OZZ\Sb   !&#eee&TTTQ][   !&#c\W]\^][]V]Q][   !&#  % !!    !&#eeeS\R !Q][   !&#e%QZW\YQ][   !&#e %QZW\YQ][   !&#c\W]\Q][   !&#QZWQY&ZS&ZSQ][   !&#abPO\\S`OZZgSaQ][   !&#[[a[]gcQ][   !&#c[]gcQ][   !&#[[ac[]gcQ][   !&#aV]e[]gcQ][   !&#Wd`aS\R[]gcQ][   !&#Wd`c[]gcQ][   !&#Wd`[]gcQ][   !&#Q]`S^R[QOabQ][   !&#[&R[QOabQ][   !&#RQeeR[QOabQ][   !&#`S\`S\R[QOabQ][   !&#TWZSaVS\PO\U\Sb   !&#PO\\S`P]fQ\   !&#eeePO\\S`P]fQ\   !&#OQbW]\Q]]^S\Q\   !&#c"aYg''Q\   !&#caYg''Q\   !&#c aYg''Q\   !&#c!aYg''Q\   !&#aYg''Q\   !&#caYg''Q\   !&#cSbSQ\   !&#W^OZSfOO\geVS`SQ][   !&#eee!$#bO\Q][   !&#eeeeW\]^S\Q\   !&#eeebO\W^Q][   !&#OZSfOO\geVS`SQ][   !&#XaaPOZSfOO\geVS`SQ][   !&#\a #OZSfOO\geVS`SQ][   !&#aPOZSfOO\geVS`SQ][   !&#W^OZSfOO\geVS`SQ][   !&#^]^'dQ\   !&#fc\W[gORQ\   !&#WSPO`b b Q][   !&#S``]`\SeQSZZQ\   !&#Ocb]aSO`QV[a\Q][   !&#Q\a!% Q][   !&#aSSY!% Q][   !&#\O[SQ\\WQQ\   !&#b]]ZaPO`YcOWa]Q][   !&#eeeYcOWa]Q][   !&#YcOWa]Q][   !&#eeeQ]^ga]Q][   !&#c\W]\Q]^ga]Q][   !&#Ocb]aSO`QV[a\Q][   !&#]Y[]^VhQ][   !&#eee\QOabQ\   !&#eeeORa!% Q][   !&#!$ORa!% Q][   !&#eee[O]VSVSQ][   !&#eee##$$\Sb   !&###$$\Sb   !&#eeeUXXQQ   !&#UXXQQ   !&#eee'"'#Q][   !&#'"'#Q][   !&#[g !Q][   !&#eee[g !Q][   !&#%PQ][Q\   !&#eee%PQ][Q\   !&#eee!#$%Q][   !&#!#$%Q][   !&#eee!% Q][   !&#!% Q][   !&#Y!$'Q][   !&#eeeY!$'Q][   !&#eeeVO]c`ZQ][   !&#VO]c`ZQ][   !&#eee!% \Sb   !&#!% \Sb   !&#eee"''Q][   !&#"''Q][   !&#eee'##Q][   !&#'##Q][   !&#%'!'Q][   !&#eee%'!'Q][   !&#eee!""&Q][   !&#!""&Q][   !&#&' #Q][   !&#eee&' #Q][   !&#eeebb[^!Q][   !&#bb[^!Q][   !&#eee!bUQ\   !&#!bUQ\   !&#eeebbXXQ][   !&#bbXXQ][   !&#eee#'%&Q][   !&##'%&Q][   !&#eee'&%$#"Q][   !&#'&%$#"Q][   !&#eeehVO] !Q][   !&#hVO] !Q][   !&# !eOQ][   !&#eee !eOQ][   !&#eee#'Q][   !&#a]Tb#'Q][   !&#eeedQ][   !&#dQ][   !&#eee&##Q][   !&#&##Q][   !&#eeeec !Q][   !&#ec !Q][   !&#eeeVO]RfQ][   !&#VO]RfQ][   !&#'YcQ][   !&#eee'YcQ][   !&#eeeb b Q][   !&#b b Q][   !&#eeeYc&Q][   !&#Yc&Q][   !&#eeed !Q][   !&#d !Q][   !&#eee##Q][   !&#eee# Q][   !&## Q][   !&#eee_c !Q][   !&#_c !Q][   !&#eeeVO]YO\ !Q][   !&#VO]YO\ !Q][   !&#eeeYO\ !Q][   !&#YO\ !Q][   !&#VO\U !Q][   !&#eeeVO\U !Q][   !&#!b][Q][   !&#eee!b][Q][   !&#eeeO\ga]Q][   !&#O\ga]Q][   !&##'%&Q][   !&#eee#'%&Q][   !&#b!X"Q][   !&#eeeb!X"Q][   !&#eeehV!Q][   !&#hV!Q][   !&#eee&%#%Q][   !&#&%#%Q][   !&#eee%$$%Q][   !&#%$$%Q][   !&#WSc\W]\ !Q][   !&#eeeRO]VO\UbcQ][   !&#RO]VO\UbcQ][   !&#eeeZR !Q][   !&#ZR !Q][   !&#eee!$'Q][   !&#!$'Q][   !&#'\WQ][   !&#eee'\WQ][   !&#eee%''#Q][   !&#%''#Q][   !&#eeeaVO !Q][   !&#aVO !Q][   !&#eeeZSbV]bQ][   !&#ZSbV]bQ][   !&#eee&%#%Q][   !&#&%#%Q][   !&#"#!!Q\   !&#$VQ][Q\   !&#eee$VQ][Q\   !&#eeeXX]ZQ\   !&#XX]ZQ\   !&#eO\UhVWYcQ][   !&#eeeeO\UhVWYcQ][   !&#eeehVO\Q][   !&#hVO\Q][   !&#eee $ Q][   !&# $ Q][   !&#eee!$#Q][   !&#!$#Q][   !&#eee"#!!Q\   !&#"#!!Q\   !&#!bUQ][   !&#eee!bUQ][   !&#b][Ob]ZSWQ][   !&#eeeb][Ob]ZSWQ][   !&#'''QVOQ][   !&#eee'''QVOQ][  %[[aYQ\  %WYOYOQ][  %aOTS__Q][  %!$aOTSQ][  %PPa!$aOTSQ][  %eee[[aYQ\  %eeeWYOYOQ][  %b]]ZWYOYOQ][  %eee!$aOTSQ][  %haYW\Ua]TbQ][  %T]`c[WYOYOQ][  %c^`WaW\UQ][Q\  %aQO\YW\Ua]TbQ][  %Ydc^XWO\U[W\Q][  %`SU`WaW\UQ][Q\  %c^RObS`WaW\UQ][Q\  %c^RObS%XWO\U[W\Q][  %R]e\Z]OR`WaW\UQ][Q\  %R\ZcaYOa^S`aYgZOPaQ][  %R\Zca YOa^S`aYgZOPaQ][  %R\Zca!YOa^S`aYgZOPaQ][  %R\Zca"YOa^S`aYgZOPaQ][  %R\Zca#YOa^S`aYgZOPaQ][  %R\Zca$YOa^S`aYgZOPaQ][  %R\Zca%YOa^S`aYgZOPaQ][  %R\Zca&YOa^S`aYgZOPaQ][  %R\Zca'YOa^S`aYgZOPaQ][  %R\ZcaYOa^S`aYgZOPaQ][  %R\ZScYOa^S`aYgZOPaQ][  %R\ZSc YOa^S`aYgZOPaQ][  %R\ZSc!YOa^S`aYgZOPaQ][  %R\ZSc"YOa^S`aYgZOPaQ][  %R\ZSc#YOa^S`aYgZOPaQ][  %R\ZSc$YOa^S`aYgZOPaQ][  %R\ZSc%YOa^S`aYgZOPaQ][  %R\ZSc&YOa^S`aYgZOPaQ][  %R\ZSc'YOa^S`aYgZOPaQ][  %R\ZScYOa^S`aYgZOPaQ][   !&#eeeOP!$#Q][   !&#OP!$#Q][   !&#eee# !#\Sb   !&## !#\Sb   !&#eeeVO]Z !\Sb   !&#VO]Z !\Sb   !&#eee&'Q][   !&#&'Q][   !&#eee!% Q][   !&#!% Q][   !&#eee'#!!Q][   !&#'#!!Q][   !&#eeePOfc\Q][   !&#POfc\Q\   !&#&%"'Q][   !&#eee&%"'Q][   !&#f`ehQ][   !&#eeef`ehQ][   !&#a[O`bbO]PO]OZZgSaQ][   !&#%YSg\Sb   !&#eee%YSg\Sb  %Zc]a]TbQ][  %h\[_Q][  %O`ae^Q][  %^QbcbcQ][  %b][[a]TbQ][  %eeeZc]a]TbQ][  %eeeh\[_Q][  %eeeO`ae^Q][  %eee^QbcbcQ][  %eeeb][[a]TbQ][   + P u � � � �  3 Q p � � � �  ) L n � � � �   %  C  _  z  �  �  �  �  "! D! _! ! �! �! �! �! " H" l" �" �" �" �" # '# O# n# �# �# �# �# $ 3$ Q$ s$ �$ �$ �$ �$ % 1% V% u% �% �% �% �% & /& Q& r& �& �& �& �& ' ;' X' u' �' �' �' �' �' %( E( e( �( �( �( �( ) D) _) }) �) �) �) * !* @* e* �* �* �* �* + '+ E+ f+ �+ �+ �+ �+ �+ , 2, L, g, �, �, �, �, �, - 2- L- j- �- �- �- �- �- . 6. P. j. �. �. �. �. �. / 2/ N/ f/ �/ �/ �/ �/ �/ 0 50 R0 m0 �0 �0 �0 �0 �0 1 51 T1 o1 �1 �1 �1 �1 �1 2 62 O2 l2 �2 �2 �2 �2 �2 3 53 T3 t3 �3 �3 �3 �3 4 %4 @4 [4 z4 �4 �4 �4 �4 
5 $5 B5 \5 }5 �5 �5 �5 �5 6 /6 I6 g6 �6 �6 �6 �6 �6 7 77 Q7 j7 �7 �7 �7 �7 �7 8 ;8 V8 s8 �8 �8 �8 �8 �8 9 09 O9 r9 �9 �9 �9 �9 �9 : : 6: O: i: �: �: �: �: �: ; -; M; m; �; �; �; < '< M< s< �< �< �< = 2= X= ~= �= �= �= > <> b> �> �> �> �> �> ? 7? U? o? �? �? �? �? �? @ 2@ P@ j@ �@ �@ �@ �@ A A *A @A XA sA �A �A �A                                                 G          2J  �                      �G  �G  �G  �G  �G  H  H  &H  >H  HH  fH  tH  ~H  �H  �H  �H  �H  �H  �H  I  I  I  (I  :I  HI  dI  tI  �I  �I  �I  �I  �I  �I  �I  J  J      ZwClose PRtlFreeUnicodeString  fZwSetValueKey �RtlAnsiStringToUnicodeString  aRtlInitAnsiString 9ZwOpenKey dRtlInitUnicodeString  �PsCreateSystemThread  �strncpy �PsLookupProcessByProcessId  G ExFreePool  �wcscpy  �_snwprintf  )ZwEnumerateKey  �wcscat  : ExAllocatePoolWithTag �ObfDereferenceObject  �ObQueryNameString �ObReferenceObjectByHandle �_wcsnicmp �wcslen  �strstr  RZwQueryValueKey ZwCreateKey �KeServiceDescriptorTable  �PsGetVersion  ZwCreateFile  �IofCompleteRequest  AMmGetSystemRoutineAddress �strncmp :IoGetCurrentProcess z_except_handler3  �_stricmp  nZwWriteFile RtlCompareUnicodeString K ExGetPreviousMode ntoskrnl.exe      �   3 3N3�3�3�3�3�34"4�4�4�4�4�455P5W5�5�56I6c6i6n6�6�6�6�6�6�6797�7�7�8�8�8\9l9�9�9�9:�:�:�:�:�:�:�::;L;�;�;�;�;�;�;�;<!<*<3<K<y<�<�<�<�<�<�<�<�<�<�<�<=6=C=\=y=~=�=�=�=�=�=>6>@>�>�>�>?????r?|?�?�?�?�?   �  000*0F0L0p0u0�0�0�0)1O1X1�1�1+2k2�2	3>3J3S3�3�3�34484~4�4�4�4�4�4555\5`5d5h5l5p5t5x5|5�5�5�5�5�5�5�5�5�5�5�5�5�5�5�5�5�5�5�5�5�5�5�5�5�5�5�5�5�5�5�5�5 66666666 6$6(6,6064686<6@6D6H6L6P6T6X6\6`6d6h6l6p6t6x6|6�6�6�6�6�6�6�6�6�6�6�6�6�6�6�6�6�6�6�6�6�6�6�6�6�6�6�6�6�6�6�6�6 77777777 7$7(7,7074787<7@7D7H7L7P7T7X7\7`7d7h7l7p7t7x7|7�7�7�7�7�7�7�7�7�7�7�7�7�7�7�7�7�7�7�7�7�7�7�7�7�7�7�7�7�7�7�7�7 88888888 8$8(8,8084888<8@8D8H8L8P8T8X8\8`8d8h8l8p8t8x8|8�8�8�8�8�8�8�8�8�8�8�8�8�8�8�8�8�8�8�8�8�8�8�8�8�8�8�8�8�8�8�8�8 99999999 9$9(9,9094989<9@9D9H9L9P9T9X9\9`9d9h9l9p9t9x9|9�9�9�9�9�9�9�9�9�9�9�9�9�9�9�9�9�9�9�9�9�9�9�9�9�9�9�9�9�9�9�9�9 :::::::: :$:(:,:0:4:8:<:@:D:H:L:P:T:X:\:`:d:h:l:p:t:x:|:   @  t  �1�1�1�1�1�1�1�1�1 22222222 2$2(2,2024282<2@2D2H2L2P2T2X2\2`2d2h2l2p2t2x2|2�2�2�2�2�2�2�2�2�2�2�2�2�2�2�2�2�2�2�2�2�2�2�2�2�2�2�2�2�2�2�2�2 33333333 3$3(3,3034383<3@3D3H3L3P3T3X3\3`3d3h3l3p3t3x3|3�3�3�3�3�3�3�3�3�3�3�3�3�3�3�3�3�3�3�3�3�3�3�3�3�3�3�3�3�3�3�3�3 44444444 4$4(4,4044484<4@4D4H4L4P4T4X4\4`4d4h4l4p4t4x4|4�4�4�4�4�4�4�4�4�4�4�4�4�4�4�4�4�4�4�4�4�4�4�4�4�4�4�4�4�4�4�4�4 55555555 5$5(5,5054585<5@5D5H5L5P5T5X5\5`5d5h5l5p5t5x5|5�5�5�5�5�5�5�5�5�5�5�5�5�5�5�5�5�5�5�5�5�5�5�5�5�5�5�5�5�5�5�5�5 66666666 6$6(6,6064686<6@6D6H6L6P6T6X6\6`6d6h6l6p6t6x6|6�6�6�6�6�6�6�6�6�6�6�6�6                                                                                                                                          