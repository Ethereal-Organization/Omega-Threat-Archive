MZ�       ��  �       @                                   �   � �	�!�L�!This program cannot be run in DOS mode.
$       A�u��&��&��&���&��&\��&��&��&��&���&��& ��&��&���&��&���&��&Rich��&        PE  L j7        �            d      p    @                   �     �:   �    @                        X  �    �  `                                                                  H  |      �                           .text   P      P                    `.data   �   p      T              @  �.rsrc  �   �      \              @  @�,�<8   �,�<E   �,�<P   �,�<Z   �,�<d   �,�<q           ADVAPI32.dll USER32.dll GDI32.dll ole32.dll KERNEL32.dll msvcrt.dll                                                                                                                                                                                                                                                                                                                             �Y  �Y  �Y  �Y  �Y  Z   Z  <Z  JZ      lZ  �Z  �Z  �Z  �Z  �Z  �Z   [      [  .[  H[  b[  n[      �[  �[  �[  �[  �[  \      "\  B\  L\  \\  p\  �\  �\  �\  �\  �\  �\  �\  ]  "]  6]      T]  ^]  l]  t]  ~]  �]  �]  �]  �]  �]                  �oe[�E:%�㮸�:�T������Ʊ�洴$�t6bR���@ �ݍ}����*  ���ƍ=/@ �+   ��G  ��4�ǁ��  �@ �s�ȉ;�HfZ�U���pV��@ ���<"uF���t<"u��>"u�< ~F�> ��< F���u�V�w���Y��                                                                                            �9�fT ���p�sq�����$����u?� �q�p��%HP���3���u%%��  �u@��������H��u-�����u2;��u>uغi  �r������,��t(��t�4��Ju����uhv@ �tI�t��                                                                                                                                                      �AVa�GаЧ2��P$s�W������@�;&6C�g���;�)�p�+6&S�w����+�8�`vKFX<g]�(�@h��#?5�e��&�4�s�[#�R��Ŧ��g�ET��Ġ�k�y� �����P4P(�M�\������@$@8�]�L�,����3�pp�m�|�<����#�``�}�l�L��֣S�th���\��ƳC� d x���l����s�0T0H�-�<�|���c� D X�=�,��^/�BЭ��1�	�P����A�����@�&6C�g�HЈ;�9�p�6&S�w��+�;�`�[FV#����[�I�t�VF3����K�Y� �{vv�'�԰�{�y�0�kvf�7�Ġ�k�y� 놖��P4P(�M�\������@$@8�]�L�,;��k2�pp�m�|�<����#�``�}�l�L��֣S�th���\��ƳC� d x���l����s�0T0H�-�<�|���c� jC7�X�>�tc�Gд¨��P�s�W������ �_GB"�u�؈;��p�6&S�w����+�9�`�[FVc�P��/�I�)KVF3����K�� �{fv�'�԰�{�i���g�7����k�	� ����S�P4P(�M�\�����׀
2]�2�L�����ó�pr�m�|�<����#�``�=�l�b����S�th�Y�\��Ƴ� d x���l����s�`T0H�-�<�|���÷ D X�=�,��c�GдШ�	� �s�W������@�;&6C�g���;�)�p�+6&S�w����+�9�`�[FV#�����[�I��KVF3����K�Y� �{fv�'�԰�{�i�0�kvf�7�Ġ�k�y� �����P4P(�M�\������@$@8�]�L�,����3�pp�m�|�<����#�``�}�l�L��֣S�th���\��ƳC� d x���[����s�0T0H�-�<�|ڮ��c� D X�=�,�O�F6��t��2�	�4c;r�S|R����8C�Ȳ6^s�g�WZ������Ўw����>��`3~v&#֌P��+�L�#n~63Ɯ@���b�s��3vv~"�İ͸��P<>��2�;��❆�$l���#I�	P�8�ՙ\��b�y�<�y��K޴H�,��u���@p0-���(=���|�`��}�lk�M���P|��\�v���9�w� aZ�[K��F�,o>���# �/�C�b7er`D�~�fI��-�"�ך�?�I#��=S�����dX��ȵL@�Q&f)L�刐�>.��p�}as(��Di�C9�`�1B>#�����1r��t�KS��F������s�fs��OаȻ�d7�̉��h�+(�B}� ��8f��(tÜ�J�Y�ti�'�{cH��}0V�.��pp�:�V�{� M#W�6�#$���@�L�C�Iӛ7T8$�|�YN����$du}@v���8���$TE�p�O�}#�>�~��+n�{#H��PSΔ�ԛ�&���7�S�.ċ�l#��"�/�c�Ԍ́���2��.3ĀY�+�9�2���%{���љr��OrDw��s����?Bt���_z�7�k��t'Rd!��ƴ���]�gB�N�7����,�M����ti�'�~fО����@�����^i����fs'�`[��zQ��$M��'Dm���x�6)98����H����a�b�vX%PH��1p����XGUIH��=�ӵ�{�KtĘ�2,%�c�s������V�G�8��d3��8��l���rw�����K����C	�ܯ)��fc8I��4쨹�����s�U����"'���V���M���-9�hs��#{�&�{ϛ���w�1D9�M�\�k���j�r$@8�(�)����Q�Ս��+>��*�[5`֚�``�{�z��$9]`�W����������O��� d &��TL����43�3���8|�n�|����	H�Q@8�8��0�MQC2K�?#�F�����3�W�/P�"�3*�S&C����Q�C��OV&V(�i�kN�?<g�$<���X�6�`YKJuWUd�f3�'hv�b����bR��}���P�8�%0Dc
4���n���!�@�ws�U1�4�M�Օ� �~xC�Ca��α�H�,���Hv�T X0(E���=��su` ����m	+�]�P @����ը�]��h8`xΖ��h�	�,u�?��+��p��o֋���e���ŷ+��F�׹ķ�PKFM"\�N�V��C�[��k�I��&�s����v3�����(s�(2���K�9�#3�#�XB|��XȽU$�Z����q�Y���#��1+;�HAy ,L`�o�#糼�8�S.�)S5P���iV� ����@��Ύ�xF��(���@�����<&�uW�6"�����6�uLd4`m�l�	L��Ԋ+��'�6��<���aɂT }sxp	�@	|��PT5{)���ve�h;�H��|8�8��*���دEH/W��i�U�ٜ��Ĝ�(:�"�o�;#�9qH��gF �C�ZFS�D2� ��X>�������g��:ћ�@]��<�#���N��TS�V�L+Ok7�i�.�eމ�C�,�$�B��@��Di ���s]u�/�����0�7����=�=�DY�S�u'�����[pMC\],�Ttd`��3X�Y�K�|`��/B��n�?1���4��l�i�4|��47�ڠJ����㠱=3�Kd6�[s䥒�B�fZ��ܸ3�t���� נ�ŋ�W
t�1���;H�7��;�.���Ұ�[��g��Y�e���E��\=wx��r�?��KSu�I�Ԁ�����@���P?�Ե��'|� �n�-_��H�['��� 	�T��������v�s�떃��]U,p8�� ��#S\L<�DDtp��#oHJ�"�;����0�}�_2��~������$��|�Y�L��p�Β�
�&�#L���-&��P/7�J�U��c���KS�e\od���0[��՛�Gd*
���y�?���G�����73[���q�/�w��}���D2o��9�`AGU��̣/0hF����ZP�
bb��;��]� �{f�'�����R|�P�n��@`�T|��k����d���
�U\R(��vI�|��3R�$@83̀L��0YI<�U�돃c��X�<���^g�dT3��Y�<�L�VϣVTP8$�|�YN����$` ߖ�(������׾0Qc��E�<��C�斋�߻�0C$�)�sBvc���Uhn�atI�E�f�7��K{���3��hL7)�`������ C>BFS��H������t�_V&;�noP�I�� �����'��K��[�=3"c�Dʧߒ3�>�p�:%z�i��@�i�4�����`b�Z�\�J����a�.a!F�)�0�z�����pun���M�˦���x`���X#��Z��V�t|�Y����� ax����l��j�s�ZTZH�-�<�|����cH5@X��tl��MQC�W�[D8V�	ٰ��w��1���-�@%2p^�͌��>n���CYEa`x�����'���:H"�r�t��Y�<���UUFۗ����>�ԈU~fvx3�<�1�R,<�*H��)������g�xy����%-�T�I�)��?��@�����?�������*I/V�$<�l������ d`C�G��V���<Dm����6ϾƙC��Tx��<�l��	|f�PT5��5�<��(�c����Z�����Kn�/�!��L����|�K|Ec~�qDS�;�#?�g�+��](�I�ɥn+����6�S��_FV��'����3rI���CbS�k����Y��4/5�G��	��l\�ks�G�7�,# �B���l�����6�U��M�\�ێ^���@$@��y�9̔��������I�9�*��&�`n`r���&ۮҿS�zt�,�%��̫��6�����8h���k�Zϫ�L�-�ԍ�	�� �5$�=�v�O�%�֨��	�P�z�%������@�;C6C�g�R�[�,���76#�T�{����9u�;FS����x��r����KV26+}~@#�Y�� �����'���$�-�i�,vfFh���0�y�������P�$�������������=�q]�L�0���+���@��i O{L�=�ZP��Dh����hiP��(KcpK6�P
�P	@:�������4�)���}[�4T0�-)0��mU��ۻ���*�f��Ðl�h\ͨ%'�cD��s�oI�<3N!��C�N�O����S4�u��#N3�r�������`ɝ@V������r<W�dKVF��@���]NEd%��/�ԵC��i7u ;!��W��g��y� f��C��!\H�Hޣ�떃��@$Ǟ��L�DO���ee|�Aa�9�I��C�encN���T�Lޕ)�{�q�����ͦ4)�K^� ���L�l����*��5Z.�S�P�����c� s�i�a��)G#'�p��Ш%	�P�S3s|��X��s�(�+&6�P�k��+�)�C�#F3�r�g�}y �^D#&;�mo+��ɡ��KSE<GD��˙L�0�~ސ��lX�D7��0�X�������R�D=�dy5cs�U���E�\դ�z-�Ѵۿ��=�I(�BYIH�pp����I�SC�el��x����� ����do\|�Y��9V�0d���Yh�	 ;�0Q�q8��yS�n��_��ߧH}�,��Ɍg�G���n{�R�c��z�R?���غ< �>���g����S=6�u�V&V�����.~���/)>�����;�L$��KS�k8��7�K�-�輍���β�Ե������?��H�['�VM,�����g�1�H�H�4H|����i�(<^8�7�&�Ӯ���6���PhA�T6�FC�e��U��}��`S�Zt���/����0� ;S!�I�A�-͠��6�oT0H�{�i;�`�S�/@D%��(#qtX�F�����E�R�G8A�yKc�p��7��f	jA�+ޕ��t<�)��a�Y��5��N�iRx�b��u��a��m �@��K�� 섙s/�'��O7k��(�kvX��a$�Ћ|���ט��"y���A�\/�HF��;s�P8}�I�Ӌ�?� '*M)l2}���<�uO����Eh~�l����ӗC�p hޑ��0��óC� � x�HR��^J�s��߷Ŏ�O��	l�<�D X�=�,��c�GдШ�	�P�s�W������@�;&6C�g���;�)�p�+6&S�w����+�9�`�[FV#�����[�I��KVF3����K�Y� �{fv�'�԰�{�i�0�kvf�7�Ġ�k�y� �����P4P(�M�\������@$@8�]�L�,����3�pp�m�|�<����#�``�}�l�L��֣S�th���\��ƳC� d x���l����s�0T0H�-�<�|���c� D X�=�,�s���bж]�΄�P��Vv����Eİ*��W��|{�򳦐���T�PR|�������Y<�U��ڤ��Y<���1pc�L�l��A>&�Z������Y�{,0�r�:łl/�Y蘕�T�R��wWc�N����RH �N��̪��5��uj���Rqѯf�����=����E��=�yև˿a��޺�')嗉�����.N�i��������Dѭ.�?7iy�r�1�'�7�Y�[�;x��l-�>@�j���;�)�c݇��I�tS3�3�[�fʕ��K�tS3��+�#ہ��_�4'��_8�ɁjFMܰ�'��/H���:���Jg?��=h���:V���8U?��Hu;3���~0E��� =��u;3���~0E�����H���:V���8U?��=h���:V���8U?��H���zΰ�$%��M(��zzcΰ�$%��-H٧�:y���Jt":uY,�'����i�o",'U��	�ztD-��������~���7H�쇑�b0䱐B5݈�r6G��^��)?���3�yeۜ�W8؝�R��yۼ�W88���?�n������8�+Q�N�9�����8�+Q�n���|78�z�뿑�z�E�|78�z�뿑n������8�+Q�N�9�����8�+Q�n��[����x�]k?��y�[����x�]k?�n������8�+Q�N�9�����8�+Q�n���|78�z�뿑�z�E�|78�z�뿑n������8�+Q�N�9�����8�+Q�n��[����x�]k?��y�[����x�]k?�n������8�+Q�N�9�����8�+Q�n���|78�z�뿑�z�E�|78�z�뿑n������8�+Q�N�9�����8�+Q�n��[����x�]k?��y�[����x�]k?�n������8�+Q�N�9�����8�+Q�n���|78�z�뿑�z�E�|78�z�뿑;D~���i�Jۆ��DL��'i�߹3>\��s!�������NЃ��a���W������
�_�ۙ�6~K�iŒ������rmm����{75^A�����Ί¯���-���R��vT�϶C�F�R��03�!�5��CJ��wa*�h��Xԝ�7�;"C���~@DL]Ə�x�+i^BX��� Ĺ��y:�d�l�Q�����[S��L�4�+d&O�Я��Vj�վ�:+��p�����W]Q x(l�̮H �� �k)q�XŻw�}����P��^��}r�b}QWI����߆�k ���r�G���/ŷ9�3�G �]�}��݉Ý$�ʹ��,Y�\�y�@��3��x�T�Us��7K��Bl:L�U.���Y:J�X��#ʂ���Z�1F �*>������ç׏�-�/Vg��&2,4�1"O��U���:=�y�;�Iӡ` f��|t�����q���Mc*%x��*�#���-��p.���3}�j���GY�vG�䴻g�qQ�0�pqrmz�:-¸�����q�P)*��.il��ו+�40X�NYCH�ĕ���K�i���T�_Z��`q��>�LGh}#�M}�`U�j����2O{�r1�'d�[��*�jf�[�7O��ʦF�A���(#�j�0�0��-ц^���P��Us=���,�$b'���x�u��?Z�w�痝��^��(�OD2�@��m�Ҭ4��|5��@H� G糭>@0���M'�~5��x)^軬���S�����Q�f!6:!���T�-��Y R-Uf��v�dB��i�Af9 ԗ����*���w��$���&i������e?��x�h�C��vf?}��*ðZ^���f�A�1Rr(G�U[3�[U�>��sn0�V�>H�j�¦�Z+`8�B�V������N�@s3��އ<u���;jI��H�k��L�D�/�L.�o!SɍPK�'��l.������8Z� (R0�T�3:�0\0���L{)rK��.�O�(tҜ�������,��lA�}Ů�lm�܇D�v�*��+c� !����(�U��^Y��t�-�Ś�Ҩ*0�$�`Rv���}�WX/I������`�R���j���`I5�}�,}�L\��`&E�U��p�`�}w.� ?P۹�U�3Z���/=��C��˚rC��}�t[������L�>Q�F��9������0^�Q�O���YX˸�����6�Q	��g���m����h�s�,����>;h�� Z'l��eϳi��\t���R.h)�-�%C����H/1��r��`c�EM���3i$�Ks��+tЖ������_l�%B��X4����^ӆ�?O��]��zmT�M�2���&� 4��Z&-=��m��Ԝ�1��_����WrQ,%獪�z�2�+�o��"��n�/�Ƈ��hS�V@r<ٺ��Z#�$4�����N��L���8*����U�U��ȋk��!�?�63���rF�9��Gj3p�Lx�/��}\e+
�xI�8n���i�C��V\���2�5���XX�u��(�5U��Nk$���q�g������U�j��U����6��_c�U��̎�O��)�O�i@�4[gp�f�F���f@�sp<�T��A�u[E�n��A!·O��T#h��d�=�b�f�1c�{I�|]�^��ZE���UÓ�\>>:kc�r���16;0����4��>O���S^�Ѯq�+���4�
�y-3��BW��or��ٞ]%�ۉbT��ػ����S~�*����Ɍ���F���_8e���]���4�c"(w��n�}V��Y�AR�֪;��.�H٩:��Dt��Ǿ�g`�<�Qgʭ��Y%dhyDJ�+ߏ�w^���(�5��˾�*8��~�²v�*Μ[[�2�Z|=,r�-��	�dʊ���\��(�X�F����[��5Y��~��:����� �2�[N��=��ӑ�����No?Lt&,���Js�liP��_��ǿ��<���̄v.Mdh^��*k$ i�#H�������W!��}Hl��!ْ�2�O�_T��(�0EǸ%�|3�2����[Lm���'0�����TDFQ2;���SJ�cQ��6-��lGtׯ�-Bv�`�.�5���r"�֖_/��͋�i1
	����)�u�5�|d17J�9t��R�����+]\�ڮ��H��$E����#��Y�q��OR_:���?��W4�i��?��t�i2~����p�]I*�����}����ZI/��c��S�G<�w�Bw����C%#դf~DױP��S	�t�_U��H����2�r$������)���t�a�B�)u7gd�mf3���ǂ��pV��oYP��|��q� �w��,	z�K�O"s6�EO-�ޥ{��(�U��ڽ�0�1a���=�`Az�I@��j>7����d�X��+ԢEa��Ld;7ޛg!,�0l��� ��y�o��ФH��[6�;~���VR���XhO�;�"4d<2�ף�>M3���9FH�qM�v��ˢ4!��C5�����r:��v\�(�<��8{��r&�	�;�/��O���'�ζ���)i���܀M�U?Tjj0Ro�w4h�|r�Q�3��kѦ�~�*��Q��cKՅ���qG$���d�\�љ�5ʽYl�ʊ��{b���ǐyd�����0�� B���^i7�����-	�ɢ3[�CB�9
:��X˚ -es��������Xw5�ΨM<���܈�4�H0^bȇ��p]�ˤ�y�)�P�"�!%#_H܎���e#-�r��l!n��A�5�����	!�#�ʰBF�ҟ;_K�=7��ʿ�&p���/�u��d��<_�8���Sad0�,��zG6Y���%�)-i�1�ʟ�L�+���\]�\w��$i�5��=9,$�t�w��X\����rt���π<R	,�;�J	H�6�KBIX��(���gZ�]�0[^�g�C��%���
_�w���/��7h��������|*���g�{P��N�/�
e�K�o.p�������n5��ᨐ�9U��� \�5�-�~W�}���ޯ"�/	z!o0��f9ς4u�0�z�11�l�g�`��/�Ҹr���&�ޣE�r��7����Z���z����{�7�G��' ��-�)�݅��H�@�����š�r��ώΟA� 옶&~��#������T�f-�ܱI���^����S��{x�,	��������9��T�)���z�g�����k}�Sp���v�'T	ʷVk/Z!|�V5�~���y����B���W�U��]R9n�$�x��S��HғԢ��9�D��1NνΡ�{4r��I���a���x3i��F�ɷ�=�/��]�Z�^v����y�K�<����$X���e
��z]��/�;��f��)j9CA�hd�K���,��2T=�&'ge��ObKxq:���m��֐.ve�X�(�qT"���V�B�V3X*��ݚh�`,n����r`#ꩂ���E�-9�8�u���v3B#�|M�E��40�
p�d�/cp��[
k��q�6�kx1$��&)SD��[(��/�e�`�� 5(Y�+�@)�C �G���)�@k.u��z���%R�=���e+~�l�)�v{�;��b�҅��H	����|�n��"e��إC� 0r���;ٚi�������k$��P�f�!_능�f艷N�/�,���蒂�+9��=̭kV�h���(���}x��3A1�G�~N��Qe�;#������!;Z8�):@��AO^giH�,�P��$y�D��6$�;�žs����M��΃��I �P� ����L ,f����|p^x�M� ��6F��{W�7������[����X�EWЯ� ����=�5gWO{�3�y��&�aԶl��3�����+�I�h�8�i�������ڞ�?mih�(�HΙ$��4���3V��q�F�<:7<%rFb��Ο�$JGO{����S�cA���Zc�����:d���랾�(�x����M��ѝa���bLQxCu��fX[9OSxS�ɋS��� z|)l5���=��	z��)���I�Yǃ���PҚJȒ�ځ����$�,��j�K���lc@p�u���g����f���{VZ
��P8��Z�ߪ���g��"R��8O8+��j�u
S���?��v�
�O<x#fڷ4���c�Y�mF�3zJS�*�Ԑ��8�ET�>�TuVo���5=]s��3~�P�xU6h?~���MΞFn��ې��*q��T� �`�Dk���L���B]�i�RT�)�R�;�@jS�'�}h�g0y=��zW�<ۄq��=&zm<��8����iލ(��*9�\P�i���s��]�q�[����R'2�2�<�V���~z��99Z0$qmh�H4��?A�eX%ׅp�!I��7��7�tV�v��5w+����a�%�؃�nu���d��Tq��D,�'��ͅ�v8���*^�nF�"����1�!>��a�j~f�躧����V�frf�L�V[��n��u��	0
"�W�K$���K�MB���Oѱt!3�t��9���!3���4�|f��,*�O��%J^����������[�>fɇ�f\���M�*�n�j][x�Oj/�lG�/����A��+F4�oE��o%�LP�S���Xt��d~|-#3���ί&A�Wǅ�@���'%��7V8!>�	��%G) n{�������K�)�s������L)�L�3�d��5�����~KP����|���7���-�N�=O����i�o�y�s4����q���֠��ܛ��
�a�S�ỳǒ[��4F7!�++a�04����a_g�DT�Q�ݷD-�y�o"ӏm����Xc��ɜ-�g0,�4<���Y�����<�3�����2���ԯbyo"&kcB�>M��5IN<�3
3�Žn�"��ܟS�L���S�;��ͱ�5���q��	cW�練�c[�0t�FX���렵2�|�i*��c�8��o��*��X|���5�-��.�$�Z�/$������1j�a�cvr@�b#���k~�VF`o��@��Ń|���z����#���"79P��D�B��f`(�j�Zl�����+<b��D�mhB:6l����=-��bu��H�?X,��� �/?��y�~0tOO{�����P��2�0�,C�˞�h�,�#�J�U��l-��X ��fT����af�M��.u,'m;��f�0�纝Oq,�TW��1�Ոh��jB�y��k�p3l��uI5]�/����"��r��%�X!�D0�pu��o�m�6��_v8>ď+��QYa�A2���sV�e��т�o�1N�O]5^�q,V�Yօ��w�t�0����i���t|U�Ur���H�xZ��d��ip����������Gt��Q����u��<XøU��:�`�+A��Z;s���]$�hW�����S�H�\}���5�j�W�
#֬��{��N�����M�'z���:�d@7x��N"ػk�#VT!	��L��@���_���%KvnD���f���Bc�%PӕH��UA��Ҩ���m�=K��_�ϽH-K����}U�n��~��o��ηO�We��h�f�I�h�TN�)�!f�͖ښ��Ϝ�}��q�����v �B9�?^��6;�y��0g��b�H��&&��ł��q��W���S �GL�����M�j�\�����,^ف6f�ǐ&� <^�1l�(W����6}~�(�X�[T<�����t��Q����++��FnDSK�ﾯֿ]WܽE�ڞDw�.s i���N8�J;�k�!�s����1�.�.J�b��#��K��ȏ&�%������J�ʝ�eA���P����I��!����P����I݆eA��C����RÀ	��Ea��C����RÀ	��eA�3�oX�"�@�]f��
3�oX�"�@�]�rr��W��8��R��	��LRʥ��:��Ry:	��pr�=���d��y:I��(�[��ؼ_�}>I�Z�u�����S�R=~	�>�U����z��R9z	�|�A�e�[X�e��l}δ*�`o�uI�^7�a�8��(��=���m��z��xٮ��kϷ��VQ��!��;��7��M��2&��"��F��!��B��@]��z��������p�� ��h��ȺՃN'�a��=E�w�`��CC�~�98�d~��AK��%��͢��k��n��d��Vյ2��X��j����%����Ȍ0k��^������ݟ\�`ܟJ�R��}��M��@��s���׻K��'�\L�^�5~��6�OI�r�}�+�-a��ר`��b����:������~��.��/��S��\����;ĕ{\��z������r��[3�}݀b��V��T��Z��H��S�� ��.ϤQq��X�'^�62�RO���P�Z�C�O�-?����J����pӍ<"��/��H��6��^�,��l����^��4��w����z��a����{:��U��J����w˛#��4Ӛ+޵W��^��G�X�+U�)l�0�HLΔkh�(Q�Me����T:�4�O�ڑ2��[��x��0#��6�.��[G{�f��S��Ѱ(�co��g�S��є?�w{�N�4�s���a�[uyO�l�éV��}�[��O�R�4�)�)Q.�W��Tj��-�)Q�@P�	�T�^3���hĐ[��O�,����
��[uM{�0�3���T�����t�.�%����_�n��1����)������EǼ,;����A��;��fа"� � �|$��ȁ��t�5*������1��5��3���,��~����.��M�� ��^��<��]����"K��(��Q��+��E��e@�^��f��}͊� �j�j�Y+%P�pｴ�"�Z�U�(��0����aε	������+��i�r��,�Lo�)�{A�r:��A*�+3�on�2�:�V�J�����!\Sr�"��l�����N|�xZ��J&�WM��j[�r��-[�gs�0,�Q6�RC�%�z��Qɨ3��F��d��]��y���<�E��C9�#�Mz��'(��_~� � ]�n"�#<۾]v�%�8-�O���It��u�C%�Zʏ;C�aI�h,�s/�L�C�aI�h,�s/�L6ʏ;�,��`��C����*oۃ,��`��C���6ʏ;C�aI�h,�s/�L�C�aI�h,�s/�L6ʏ;�!	�(l�3o�V��[�!	�(l�3o�6ʏ;C�aI�h,�s/�L�C�aI�h,�s/�L6ʏ;�,��`��C����*oۃ,��`��C���6ʏ;C�aI�h,�s/�L�C�aI�h,�s/�L6ʏ;�!	�(l�3o�V��[�!	�(l�3o�6ʏ;C�aI�h,�s/�L�C�aI�h,�s/�L6ʏ;�,��`��C����*oۃ,��`��C���3ˀ(W�`C�x<�}�GĊ[�^[�RQ�~�L6��"Q�F
�c�	1�i��K-�G �f����3�.O	���ZJ��s�ĽO
��xm�A(P]j��s�y2>�u��ϰ����s�y2>�u��/P]jZv�����j�p}JZv�����j�/P]j6�X����*�U]O0=
6�X����*�U]/P]jZv�����j�p}JZv�����j�/P]j��s�y2>�u��ϰ����s�y2>�u��/P]jZv�����j�p}JZv�����j�/P]j6�X����*�U]O0=
6�X����*�U]/P]jZv�����j�p}JZv�����j�/P]j��s�y2>�u��ϰ����s�y2>�u��/P]jZv�����j�p}JZv�����j�/P]j6�X����*�U]O0=
6�X����*�U]/P]jZv�����j�p}JZv�����j�/P]j��s�y2>�u��ϰ����s�y2>��5j��@�;&6C�g���;�)�p�+6&S�w����+�9�`�[FV#�����[�I��KVF3����K�Y� �{fv�'�԰�{�i�0�kvf�7�Ġ�k�y� �����P4P(�M�\������@$@8�]�L�,����3�pp�m�|�<����#�``�}�l�L��֣S�th���\��ƳC� d x���l����s�0T0H�-�<�|���c� D X�=�,��c�GдШ�	�P�s�W������@�;&6C�g���;�)�p�+6&S�w����+�9�`�[FV#�����[�I��KVF3����K�Y� �{fv�'�԰�{�i�0�kvf�7�Ġ�k�y� �����P4P(�M�\������@$@8�]�L�,����3�pp�m�|�<����#�``�}�l�L��֣S�th���\��ƳC� d x���l����s�0T0H�-�<�|���c� D X�=�,��c�GдШ�	�P�s�W������@�;&6C�g���;�)�p�+6&S�w����+�9�`�[FV#�����[�I��KVF3����K�Y� �{fv�'�԰�{�i�0�kvf�7�Ġ�k�y� �����P4P(�M�\������@$@8�]�L�,����3�pp�m�|�<����#�``�}�l�L��֣S�th���\��ƳC� d x���l����s�0T0H�-�<�|���c� D X�=�,��c�GдШ�	�P�s�W������@�;&6C�g���;�)�p�+6&S�w����+�9�`�[FV#�����[�I��KVF3����K�Y� �{fv�'�԰�{�i�0�kvf�7�Ġ�k�y� �����P4P(�M�\������@$@8�]�L�,����3�pp�m�|�<����#�``�}�l�L��֣S�th���\��ƳC� d x���l����s�0T0H�-�<�|���c� D X�=�,��c�GдШ�	�P�s�W������@�;&6C�g���;�)�p�+6&S�w����+�9�`�[FV#�����[�I��KVF3����K�Y� �{fv�'�԰�{�i�0�kvf�7�Ġ�k�y� �����P4P(�M�\������@$@8�]�L�,����3�pp�m�|�<����#�``�}�l�L��֣S�th���\��ƳC� d x���l����s�0T0H�-�<�|���c� D X�=�,��c�GдШ�	�P�s�W������@�;&6C�g���;�)�p�+6&S�w����+�9�`�[FV#�����[�I��KVF3����K�Y� �{fv�'�԰�{�i�0�kvf�7�Ġ�k�y� �����P4P(�M�\������@$@8�]�L�,����3�pp�m�|�<����#�``�}�l�L��֣S�th���\��ƳC� d x���l����s�0T0H�-�<�|���c� D X�=�,��c�GдШ�y�P�{s�W������@�;&6C�g�Ҁ�;�Y�p�[6&S�w���E�U�R�?*:#�����/�(�@�$"#P��䀫.��n�
W�Sܱ��{�i�H�&|�Rӷ��k�y� �����P4P(�M�\������@$@8�]�L�,����3�pp�m�|�<����#�``�}�l�L��֣S�th���\��ƳC� d x���l����s�0T0H�-�<�|���c� D X�=�,��c�GдШ�	�P�s�W������@�;&6C�g���;�)�p�+6&S�w����+�9�`�[FV#�����[�I��KVF3����K�Y� �{fv�'�԰�{�i�0�kvf�7�Ġ�k�y� �����P4P(�M�\������@$@8�]�L�,����3�pp�m�|�<����#�``�}�l�L��֣S�th���\��ƳC� d x���l����s�0T0H�-�<�|���c� D X�=�,���Gп�+�9�`�;\6!�6����;�)@p2�k�(���6
 IB{�����u�b�
�S�h^e��6���lo}$$Ls���B�O~!lC5;N�C��+�ˆ�M�_��]P�Փ�s�]`O\����$�g{g�+�2�a��k4pw�w������*�����H�H�����S�?X�X�s�y�k���j�)?)����ɩ��5�Kz�:�:����꺀�̍H�a�~�g�М��X�;�Я�! �-����n�H '2&k�7&:3����W7�$�}�%���q]M����A�R)2]�euh�H����e�w.Pu�x����$�5uKgi>E�H�4�͏�D�V��TNYY�x���XT4F#��$�W,1o4p(�m�\Н��]3p�p𻑩���E��3�pp�m�|�<����#�``�}�l�L��֣S�th���\��ƳC� d x���l����s�0T0H�-�<�|���c� D X�=�,�                                                                                                                                                                                                                               �X          ^Z     �X          [  (  �X          �[  L  Y          \  d  ,Y          F]  �  lY          �]  �                      �Y  �Y  �Y  �Y  �Y  Z   Z  <Z  JZ      lZ  �Z  �Z  �Z  �Z  �Z  �Z   [      [  .[  H[  b[  n[      �[  �[  �[  �[  �[  \      "\  B\  L\  \\  p\  �\  �\  �\  �\  �\  �\  �\  ]  "]  6]      T]  ^]  l]  t]  ~]  �]  �]  �]  �]  �]      YLsaSetTrustedDomainInformation   AdjustTokenPrivileges � GetSecurityDescriptorSacl �RegOpenKeyExW g CryptDecrypt  � EqualDomainSid  LLsaQueryTrustedDomainInfo  AccessCheck y CryptGetProvParam ADVAPI32.dll  �PrivateExtractIconExW �IsCharAlphaNumericA 	RemoveMenu  7 CheckRadioButton  � EnumDisplaySettingsExW  � DestroyAcceleratorTable � ExitWindowsEx  GetCursorPos  USER32.dll  � GdiPlayJournal  \GetOutlineTextMetricsW   BRUSHOBJ_pvAllocRbrush  � FillPath  [GetOutlineTextMetricsA  GDI32.dll ' CoGetCallContext  � OleCreateEmbeddingHelper  k CreateClassMoniker  [ CoSetProxyBlanket � MkParseDisplayName  � OleCreateFromDataEx ole32.dll ^GetProcessShutdownParameters  � ExitVDM �HeapQueryTagW gGetModuleHandleA  eSetCommBreak  �GetStartupInfoA �ValidateLCType  ZGetProcessHeap  � GetCommandLineA �VirtualAllocEx  GetDiskFreeSpaceExA [ DefineDosDeviceA  WritePrivateProfileStructW  .GetFullPathNameA  � FatalAppExitW KERNEL32.dll  � _c_exit � _fputwchar  \ctime 
wctomb  C_wtol � _fpieee_flt �putwchar  ufreopen _wgetcwd  1_ismbckata  msvcrt.dll                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                 ��.;+++�k'�{Ơk�돠.;+++�k'�{Ơk#��]\��ܢ�2�|D��)sA�΢�
(��TU�:��w2���)s��΢�
(��(��(���TU�X]\����8�oO/8� !N�+++*oO/m�/8��~�oO/��O/��O/��O/�oO/�ߦoO/�/+++r���e��w0m8��0��9/O)oO(�/O��9oO*)oO)�oO*��9gO))�gO)9_O()O�_O(le~�_O/��/+++B����oO/RQTUP�k+X]\^������/O8�oO/��*~,����Ө�)~,�����Ӡh7(�ks(蠃K( �[(آ_O#�[O(آ_O'�sd��wEl8��o�+(�����0/O~�oO'$�/{�_O#�/�(�oO/ /md~ޠoO/��VTUP�k+X�S�kK�h#�*+++���m�\����(�*+++�E�~�m����h/�)+++��`�"?����h'�*+++��,�I����h�*+++��W&����h�*+++���������h�*+++���{�����h�*+++�G)'������hK�*+++��5Р�����hOP�k+X]\^����Ӡ�\���]'�+�++�+\���]�k�+;++^\���]#VTUP��X]\^�����\�]K�Ӯ�~-\�]��^X�]VTUP�[$�k(۠��ꏠ.;+++�c#�k+X]\^���gO/�/O8�oO#���+++�?O(��m'(/O�oO'8��5+~.�m�-�-(/O(���^��+++�x'�/O(���) #���++� �gO/�ޠoO'X����oO�wO+?�m(/O(�ۦoO�/+++������/��~����u'+$�p����oO#*+++�oO#��VTUP�]\^��A��8��e��ym8١g.+;'��9�;'k��~)8�ie~VTU�k+^����X]\�Ң^�n��f'�^�n������~��m7(n��(�(�[[�(�k?�f#�����^�)�n�3+��(�c_�^�������(�������($�k-c��ynk�n�8Р^��7�(_�'�g��o�(n�����n�[�k�o�#[�n�+(o�'[���n#�[h�f�~�TUP�V�'+]X�폠.;+++�k'��'�+0{~�[�cPU�k+^����X]\�~�u#�U�m'�n��/�+;++\�+���X#�n��^��m/�������n'[���X'\�n�[X�f��^�n������v�+_�n��[?�f��n'z����n��k?������^��n�������*~M�n��kC�^�(i?�n��n�[�+�+�n�[�+�+����X/�+�XOTUP�V�'+^�ZX]\���5�+++�e��8�����n��v�+j�^���������V�@�X++++S��k+BӢn�P��k+(^�(آ۪++��]\X�ۦ.�k+�+�m�[OTUPRV�^�ZX�*+++��y`3����Ӂ/�+;++�+/++�+���آn��n��SK�n��++{k+�n��k/jk+�n��k#+o+++++�-��lۿ���"�[�v���'U�+++�ρ/�+;++�+/++�+���ؠ^��i�n�PRV�X�����Ӡ�6��������P�+���
�ز'�ݵa���é݅F�Z�҇ �5�ȗ��̫�wD��:S]�                                                                                                                                                                                                                                                                                                                                           �                  0  �               	  H   `�  �                  �4   V S _ V E R S I O N _ I N F O   4 ���       y    y?                        \    S t r i n g F i l e I n f o   8    0 4 0 9 0 4 B 0   H &  C o m p a n y N a m e     M B E Q E U   C o r p o r a t i o n     L "  F i l e D e s c r i p t i o n     S s y d u o r i   U t i l i t y     8   F i l e V e r s i o n     5 . 0 0 . 2 1 6 9 . 1   8   I n t e r n a l N a m e   g u g u h 3 2 . e x e   \ 6  L e g a l C o p y r i g h t   C o p y r i g h t   ( C )   M B E Q E U   C o r p .     @   O r i g i n a l F i l e n a m e   g u g u h 3 2 . e x e   D "  P r o d u c t N a m e     S s y d u o r i   U t i l i t y     <   P r o d u c t V e r s i o n   5 . 0 0 . 2 1 6 9 . 1   D     V a r F i l e I n f o     $    T r a n s l a t i o n     	�                                                                                                                                                                    