MZ�       ��  �       @                                   �   � �	�!�L�!This program cannot be run in DOS mode.
$       PE  L �s�@        �  �   �            �    @                     �    `                                �  (      Dg                   p 	                                          @      ��  �                          .text   ��      �                    `.data   P   �      �              @  �.idata  H	   �   
   �              @  @.rsrc   Dg      h   �              @  @.reloc  �
   p     :             @  BI�C8           MSVBVM50.DLL                                                                                                                                                                                                                                                                                                                                                                                                                                      ?�@ ��@ F�@   �@ �@ �@   s�@ ��@ z�@               �?  [�@ ��@ c�@   ��@ ��@ ��@ '  ƣ@ �@ ͣ@     x@    E�@ [�@ j�@ ӟ@ 9�@ ��@ �@ &�@ 3�@ 3�@ ��@ �@  �@ -�@ -�@ ��@ ��@         '  ]�@ ��@ d�@     �@ !   ��@ ˤ@ ڤ@ C�@ ��@ �@ x�@ ̦@ ��@ 1�@ ��@ O�@ ީ@ 6�@ G�@ :�@ ��@ ��@ ��@ խ@ �@ �@ <�@ M�@ @�@ ��@ ��@ ��@ ۱@ �@ �@ J�@ V�@         /  ��@ E�@ �@     �@    j�@ z�@ ��@ �@ �@ ٵ@ ��@ ȶ@ ȶ@ �@ ��@ ��@     .      ��@ z�@     �@    ޷@ �@ r�@ ��@ z�@ ��@ �@ U�@ m�@ ��@ ��@ κ@ �@ �@ �@ �@ .�@ B�@ V�@ V�@ [�@ s�@               ��@       ��@ t�@ 
      ��@ ��@               �?      q�@ N�@   Q�@     X�@         �%`�@ �%��@ �%��@ �%@�@ �%�@ �%��@ �%��@ �%�@ �%D�@ �%�@ �%��@ �%��@ �%��@ �%��@ �%��@ �%��@ �%@�@ �%��@ �%X�@ �%��@ �%X�@ �%��@ �%L�@ �%H�@ �%��@ �%P�@ �%��@ �%(�@ �%��@ �%��@ �%<�@ �%��@ �%�@ �%t�@ �%��@ �%�@ �%��@ �%d�@ �% �@ �%��@ �%��@ �%8�@ �%��@ �%��@ �%$�@ �%��@ �%`�@ �%��@ �%��@ �%�@ �%(�@ �%4�@ �%��@ �%T�@ �%0�@ �%��@ �%\�@ �%4�@ �%<�@ �%��@ �%��@ �%��@ �%��@ �% �@ �%l�@ �%��@ �%0�@ �%p�@ �%T�@ �%��@ �%H�@ �% �@ �%��@ �%�@ �%��@ �%P�@ �%x�@ �%\�@ �%�@ �%8�@ �%��@ �%D�@ �%��@ �%��@ �%L�@ �%$�@ �%�@ �%��@ �%�@ �%�@ �%�@ �%,�@ �% �@ �%��@ �%,�@ �%�@ �%��@ �%|�@ �%��@ �%��@ �%h�@ �%��@ �%�@   h�z@ �����      0   @   8   jh�L16E��7��PX�               mscomm  MsComm 0    ��1 ���d�J�F����R���s�Է��B�����!�:O�3�f�� � `ӓ                                    �c  �b    frmKillAntiSpy  Form1  B #�b  lt  ~b     	 00   h  �        �  �     (  �	  00    �          �  �      h  ^"  00     �%  �'         �  nM       h  ^  (   0   `                                      �   �� �   � � ��  ��� ���   �  �   �� �   � � ��  ���                    �wwwwwwwwwwwwwwwwwp������������������p������������������p������������������p������������������p������������������p������������������p������������������p������������������p�����������������p����������0������p�������� �30�����p�������;;��0���p�������;0?� 30���p�������;3;�3;����p���������� � ���p�������0������3��p�������3�  ?�3��p���� ����������p����p�� ���� ���p����p���;����p����p���������p��� � ��0�������p���pp� ����p������ ��������p���p��p������p���� �� ��������p���������������p�������� ���������p�������p�������p����� � ���������p������������������p������������������p������������������p������������������p������������������p���������������    ������������������������������������x����������������������������������x��������������������������������x��������������������������������������������������������������      �      �      �      �      �      �      �      �      �      �      �      �      �      �      �      �      �      �      �      �      �      �      �      �      �      �      �      �      �      �      �      �      �      �      �      �      �      �      �      �    ?  �      �    �  �   �  �   �  �   �  �   �  �   �  (       @                                      �   �� �   � � ��  ��� ���   �  �   �� �   � � ��  ���             wwwwwwwwwwww������������������������������������������������������������������� ��������� �0�������� �0�������3�;�������0���0�������;� �0�����  � �����8������x� ���������������� ��������� ���������p��������p� �������������������������������������������������������������  ����������������������x������������������������������������������  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  ?�  �  �� �(                                             �   �� �   � � ��  ��� ���   �  �   �� �   � � ��  ���       wwwwwp�����p�����p����p��p�p����p���p��p�0��p�3��p�����p����  ���������x���������� ��������0�������;������0��0�(   0   `                                     7 6% U   D) W, U9 N0! `?,  y (y "|% UG+ bB0 Ot8 'G_ Io :W} III WVV sUS kqR bYe Ja} fee wid ujs vwx �   �f �s  �z  �NN �SS �_^ �hY �he �rk �ut �nj �tm �ys �|q � � � � � /� � � � (�& �% �) �1 -�$ 0�"  �/ 2�6 $�6 >�: I� s�6 K�7 |�< '�; �S =�F 6�F &�x u�F W�O u�G o�s ,�C 1�K 6�Q :�W K�c C�e {�n G�k L�s R�{ ��  ه5 �9 ��1 ��Q ��M ��q ��h ��v ��t ��{ ��} ӒR �F �G ��C ��D �\ ��V ʕf Мl ��y ƕz ӥf �i �l ��b �w �x �v ��| ��t <�  F� L� T� W� (M� *k� f� k� q� x�  n� x� z� (v� @|� iq�     �� /�� v�� _�� [� X� _�� l� �� �� �� �� 
�� �� /�� �� �� '�� *�� 8�� .�� 5�� O�� J�� t�� G�� C�� Q�� I�� Z�� |�� _�� M�� T�� c�� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ͛� ۗ� Ě� М� ⚎ ᛐ ��� ͨ� ٦� δ� ݵ� ʢ� ԥ� ٳ� ୊ 㲌 � ��� 嶑 � ̴� ֺ� ɹ� ־� ��� 弢 ��� ��� �ژ �ՙ �Ч �ɮ �� �� �̑ �Ê ��� �Ȗ �ؖ �± �ħ �ȩ �Ш �Ө �˶ �ʹ �Ӹ �׷ �� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ���     r
 ##""""""""""""""""""""""""""""""!!!%���������������������������������!%���������������������������������"%���������������������������������"%���������������������������������"%���������������������������������"%���������������������������������"%�������������������onn�����������"%�������������������ig�����������"&��������������sno�vvvc���ns������"&�������������{{ggy}wccb{{n������")������������{wwv���vww's�����#*������������|��wvy���vvy�s�����#*�����������ٟ���}����}}����ns����#+��������������������������n����%+����������{vv������������vv�����%+����������wy~�������������yy{����%_�����������������뵫}����������%_�������������������������������%_��������������������|�����������%_����������


�������|����s������%_�����5nom/-/�������|���|�������%l����I,,
@?OML�������|�����������&l����5SQ,
,OM=DGG4�\$�蟵�������&l���双UQ7OOML4477�^������������&����H@SUSQQOMLL=749H&������������)���I

LUSQQOML=774-

@������������)���<LOUTSQҳK,3334--@������������)������UTS�
,--22-J������������*���֎�UTS�,,--42-t������������*������TS�=7744J��������������*������/TS�=7741s�������������*������QTS�=7749��������������*�������TQ��[R7R���������������*������������������������������^�����������\������������������μ^���������������������������������*%��������������������������)hVVV��������������������������*�hYYYW��������������������������*�hhYc��������������������������+�hhg��������������������������+�um��������������������������+����������������������������_���������������������������_�������  ������  �      �      �      �      �      �      �      �      �      �      �      �      �      �      �      �      �      �      �      �      �      �      �      �      �      �      �      �      �      �      �      �      �      �      �      �      �      �      �    ?  �      �    �  �   �  �   �  �   �  �   �  �   �  (       @                                     7 6% U   D) W, U9 N0! `?,  y (y "|% UG+ bB0 Ot8 'G_ Io :W} III WVV sUS kqR bYe Ja} fee wid ujs vwx �   �f �s  �z  �NN �SS �_^ �hY �he �rk �ut �nj �tm �ys �|q � � � � � /� � � � (�& �% �) �1 -�$ 0�"  �/ 2�6 $�6 >�: I� s�6 K�7 |�< '�; �S =�F 6�F &�x u�F W�O u�G o�s ,�C 1�K 6�Q :�W K�c C�e {�n G�k L�s R�{ ��  ه5 �9 ��1 ��Q ��M ��q ��h ��v ��t ��{ ��} ӒR �F �G ��C ��D �\ ��V ʕf Мl ��y ƕz ӥf �i �l ��b �w �x �v ��| ��t <�  F� L� T� W� (M� *k� f� k� q� x�  n� x� z� (v� @|� iq�     �� /�� v�� _�� [� X� _�� l� �� �� �� �� 
�� �� /�� �� �� '�� *�� 8�� .�� 5�� O�� J�� t�� G�� C�� Q�� I�� Z�� |�� _�� M�� T�� c�� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ͛� ۗ� Ě� М� ⚎ ᛐ ��� ͨ� ٦� δ� ݵ� ʢ� ԥ� ٳ� ୊ 㲌 � ��� 嶑 � ̴� ֺ� ɹ� ־� ��� 弢 ��� ��� �ژ �ՙ �Ч �ɮ �� �� �̑ �Ê ��� �Ȗ �ؖ �± �ħ �ȩ �Ш �Ө �˶ �ʹ �Ӹ �׷ �� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ���         �������¹�����������������������������������ۻ��������������������������������������������������������������������������������g�����������������jnxxZs^m�������������ww��w{���������������x��}y��s���������������������r���������|}��������}x������������������������������������|������������s�,,����|�����������,@OM����|�����������U6,OM/8F^^����������ITSQOMC74H����������,/TSQPF764,,������������US׵,,-3-�����������UQ�7644R������������QQ�=74m�������������UQ�>=4�������������������������������������������������μ�������������������dXWW]������������������pYYb�������������������hj�������������������l�����������������������������������ϰ�����  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  ?�  �  �� �(                                            7 6% U   D) W, U9 N0! `?,  y (y "|% UG+ bB0 Ot8 'G_ Io :W} III WVV sUS kqR bYe Ja} fee wid ujs vwx �   �f �s  �z  �NN �SS �_^ �hY �he �rk �ut �nj �tm �ys �|q � � � � � /� � � � (�& �% �) �1 -�$ 0�"  �/ 2�6 $�6 >�: I� s�6 K�7 |�< '�; �S =�F 6�F &�x u�F W�O u�G o�s ,�C 1�K 6�Q :�W K�c C�e {�n G�k L�s R�{ ��  ه5 �9 ��1 ��Q ��M ��q ��h ��v ��t ��{ ��} ӒR �F �G ��C ��D �\ ��V ʕf Мl ��y ƕz ӥf �i �l ��b �w �x �v ��| ��t <�  F� L� T� W� (M� *k� f� k� q� x�  n� x� z� (v� @|� iq�     �� /�� v�� _�� [� X� _�� l� �� �� �� �� 
�� �� /�� �� �� '�� *�� 8�� .�� 5�� O�� J�� t�� G�� C�� Q�� I�� Z�� |�� _�� M�� T�� c�� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ͛� ۗ� Ě� М� ⚎ ᛐ ��� ͨ� ٦� δ� ݵ� ʢ� ԥ� ٳ� ୊ 㲌 � ��� 嶑 � ̴� ֺ� ɹ� ־� ��� 弢 ��� ��� �ژ �ՙ �Ч �ɮ �� �� �̑ �Ê ��� �Ȗ �ؖ �± �ħ �ȩ �Ш �Ө �˶ �ʹ �Ӹ �׷ �� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ���         )�����������_�����������_�����������k�����rzbl��l�����~���������疢���������驪��������1AD��������aTOL7�������T�--�������T�E4����������������_��������eec���������r������������������j�xZ�m������������ww���{����(   0   `                                                          ++ 79333333333333333333331333333333397++                                            3
374I4O3P3P3P3P3P3P3P3P3P3P3P3P3P3P3P3P3P3P3P2Q3P3P3P3P3P3P3P3P3P4O4I373
++                                        373x2�3�3�3�3�3�3�3�3�3�3�3�3�3�3�3�3�3�3�3�4�3�3�3�3�3�3�3�3�3�3�3�2�3x377                                       �__��]]��\\��[[��ZZ��YY��XX��VV��TT��TT��SS��QQ��PP��PP��PP��PP��PP��PP��PP��PP��PP��PP��PP��PP��PP��PP��PP��PP��PP��PP��PP��OO��MM�LL��MM�3�4J9                                       �aa����������������������������������������������������������������������������������������������������������������������������������̙��OO�3�4O3                                       �aa��������������������������������������������������߿��޽��ܸ��ݺ��ܸ��۶��ڵ��ٲ��ر��ׯ��֭��լ��Ԫ��Ө��Ӧ��Ҥ��ѣ��С��ϟ��ʹ������PP�3�3P3                                       �bb������������������������������������������������������߿��޽��ݻ��ݺ��ܸ��۶��ڵ��ٲ��ر��ׯ��֭��լ��Ԫ��Ө��Ӧ��Ҥ��ѣ��С��Ͷ������SR�3�3P3                                       �dd����������������������������������������������������������߿��޽��ݻ��ݺ��ܸ��۶��ڵ��ٲ��ر��ׯ��֭��լ��Ԫ��Ө��Ӧ��Ҥ��ѣ��ζ������TS�3�3P3                                       �ee��������������������������������������������������������������߿��޽��ݻ��ݺ��ܸ��۶��ڵ��ٲ��ر��ׯ��֭��լ��Ԫ��Ө��Ӧ��Ҥ��η������UT�3�3P3                                       �ff������������������������������������������������������������������߿��޽��ݻ��ݺ��ܸ��۶��ڵ��ٲ��ر��ׯ��֭��լ��Ԫ��Ө��Ӧ��ϸ������WV�3�3P3                                       �ig����������������������������������������������������������������������߿��޽��q��k��k��լ��ڵ��ٲ��ر��ׯ��֭��լ��Ԫ��Ө��Ϲ������YW�3�3P3                                       �kh����������������������������������������������������������Ҩ��˝���������Ŷ��vhr�ʓb��\��ҩ��۶��ڵ��͟��ɗ��׮��֭��լ��Ԫ��к������YX�3�3P3                                       �nj������������������������������������������������������޿���w��k��o�̼�� 9�� >��;���L������ܸ��~��h��t��Ď��ׯ��֭��լ��л������[Z�3�3P3                                       �pk�����������������������������������������������������#J��!C���a��V�slm�R��c�� N���=��B�ҎO� A��!A���k�����ر��ׯ��֭��Ѽ������][�3�3P3                                       �rl�������������������������������������������������8]�� F�� G��7��scj�:W}�;���5���%���bUa�o]_�;�� H�� F���ut��y��ٲ��ر��ׯ��Ѽ������_\�3�3P3                                       �un�������������������������������������������������*e��:���)��� L�� >��
V��9���4���'��� ?�� A��U�����q��uww��y��ڵ��ٲ��ر��Ҿ������`^�3�3P3                                       �xo�������������������������������������������������]���W���Q���0���e��(���9���4���.���	g��h�����������{����e��t����ٲ��Ҿ������a_�3�3P3                                       �{p������������������������������������������̴�|v��?���V���P���J���E���?���9���4���.���(���#������������@|��vjt��s������ڵ��ҿ������ca�3�3P3                                       �}q�����������������������������������������8`�� >�� B��G���P���I���D���>���8���3���-���'���"���������s�� ?�� >��ln�������۶����������db�3�3P3                                       �s����������������������������������������� J�� U��n��R���O���I���D���B���c���_���+������������������ W�� U��(Y���Ì��ܸ����������fd�3�3P3                                       ��t�����������������������������������������F���`���Z���U���O���H���C���������������YYY�Hq� f�� s�� ��� ���������)����ɗ��ݺ����������he�3�3P3                                       ��u�����������������������������������������c���^���Y���T���N���H���B���������������YYY�Jn� l�� z�� ������
������*����ݻ��ݻ����������ig�3�3P3                                       ��w�����������������������������������������~���N���Q���S���M���H���B���������������YYY�(i��������������	�����������߿��޽����������jh�3�3P3                                       ��x��������������������������ө������ۻ����� t � z �q�G���L���G���A���������������YYY�+o�� ���������+�����w��������������߿����������lj�3�3P3                                       ��y���������������������#� �"y��r��m�Ȫb�
������(v��L���F���A���������������YYY�+o�����������*n���˜��������������������������mk�3�3P3                                       Ð{�����������������c�]� � � � �s�v�1�I��;�Y�5�P�-�J�A���L���F���A���������������YYY�+o�����������6��������������������������������ol�3�3P3                                       Œ}�����������������-�,�I�m�?�_��� z �
��:�W�4�N�'�:��J�%�y�'�w���������t�YXW�NNN��wY��͠�����B������������������������������������qm�3�3P3                                       ȕ~��������������۸�y��W���Q�z�@�b�#�4�7�S�9�W�4�N�.�F������,��$�ζ����q�c]V�LLL������������������������������������������ο������ro�3�3P3                                       ʗ�������������~�H�i�:�J�o�P�y�J�p�E�h�?�_�9�V�4�N�.�F�(�=�#�5��+��"�+�%�~�S�kqR��~a��Î��������������������������������������ο������tp�3�3P3                                       ͚����������U�T� } �  �/�F�P�x�J�p�E�h�?�_�8�U�3�L�-�C�'�;�!�2��*��!��� } � { �{�@��č��������������������������������������Ϳ������ur�3�3P3                                       Н����������2�6�*�@�<�Z�U��O�w�I�n�D�f��ږ�����o�s�$|(������������� ��{�@��ʙ��������������������������������������Ϳ������ws�3�3P3                                       Ӡ����������m��_���Z��U��O�w�I�n�c��������������UXU� ~ � � � � � � ���	����{�@��س��������������������������������������̿������yt�3�3P3                                       բ�������������^���Y��S�}�M�u�H�l����������������WWW��	���������	������|������������������������������������������̾������zv�3�3P3                                       إ����������������������X��M�u�H�l����������������WWW�%�9� �/��&�����|�<��ՙ����������������������������������������������˾������{w�3�3P3                                       ڧ������������������������L�s�G�k����������������WWW�$�8��/��&���)���r��������������������������������������������������˿������}x�3�3P3                                       ݪ����������������������?�_�L�r�F�j����������������WWW�$�7��-��$���0�"������������������������������������������������������ʾ������y�3�3P3                                       ୊������������������������K�q�D�f�������������jjj�UUU���M�}�b��)�x�w����������������������������������������������������������ʾ�������{�3�3P3                                       㰋���������������������������������������{�~oa�LLL�LLL��������������������������������������������������������������������������ɾ�������}�3�4O3                                       岌�������������������������������������ݵ����n�[WR�ddd�����������������������������������������������������������������������������������~�6�7J9                                       紎����������������������������������������������������������������������������������������������������������������������������������pp��ji�:"�?$9;'                                       귏������������������������������������������������������������������������������������������������������rl���R��� ��� �� ��z ��p ��f�}QN�?$UB)I$$                                       �������������������������������������������������������������������������������������������������������un��̙���R���D���6���-�ٌ9��SP�B%YC(&F.�                                          �������������������������������������������������������������������������������������������������������xo��֣���[���R���D�ۓI��VQ�B%YC(&F.�                                              ���������������������������������������������������������������������������������������������������������{p������g���[�ݛ[��ZT�B%YC(&F.�                                                  �������������������������������������������������������������������������������������������������������}q������t�ޡj��]U�E%YC(&F.�                                                      �ĕ������������������������������������������������������������������������������������������������������s������{��aW�D(ZJ(&F.�                                                          �Ǘ�������������������������������������������������������������������������������������������������������t��߶��bU�D(lG/+U+�                                                              �˙��ֱ��԰��Ѯ��ϭ��ͫ��˪��ȩ��Ũ��æ�����忤�㽢�ມ�޷��۵��ڳ��ױ��ծ��Ҭ��Ъ��Χ��˥��ɣ��Ơ��Ğ����u���t�                                                    �      �      �      �      �      �      �      �      �      �      �      �      �      �      �      �      �      �      �      �      �      �      �      �      �      �      �      �      �      �      �      �      �      �      �      �      �      �      �      �      �      �      �      �      �    ?  �      �    �  �   �  (       @                                              3
874I4O3P3P3P3P3P3P3P3P3P3P3P3P3P3P3P3P3P4O4I373
++                        875x4�3�3�3�3�3�3�3�3�3�3�3�3�3�3�3�3�3�3�3�2�3x377                       Ϟ��ۧ��٦��ؤ��֣��֣��ԡ��Ӡ��ў��ѝ��ѝ��ѝ��ѝ��ѝ��Н��М��М��М��М��М��М��М��ޘ��3�4J9                       ͱ�����������������������������������������������������������������������������������̙�ᜐ�3�4O3                       ɲ�������������������������������������������޽��ݺ��۷��ڴ��ر��ׯ��֬��ԩ��ӧ��Ѥ��ҿ�ᜑ�3�3P3                       ̵�����������������������������������������������޽��ݺ��۷��ڴ��ر��ׯ��֬��ԩ��ӧ��ҿ�ᜑ�3�3P3                       η���������������������������������������������������޽��Ǖ��ȗ��ڴ��ر��ׯ��֬��ԩ��ҿ�ᜑ�3�3P3                       и�������������������������������������������˝�����ͼ��vku��^��۷��ٲ��Ɠ��֭��֬��ҿ�ᜑ�3�3P3                       Һ������������������������������������������Λn��h�H�� K����Q��y���u�ܣm��Ɠ��ׯ��ҿ�ᜑ�3�3P3                       Ӽ�������������������������������������� G��A��sej�8���4���Ja}�c\g� G��4U���Ï��ر��ҿ�ᜑ�3�3P3                       ־��������������������������������������V���2���P��;���2���n��[�����1����y��ɗ��ҿ�ᜑ�3�3P3                       ������������������������������������`t��T���M���D���;���2���*���!���������wnv��{��ҿ�ᜑ�3�3P3                       �³�����������������������������*h��`��Q���K���B���R���<���$���������k�� N��ͦ���ҿ�ᜑ�3�3P3                       �Ĵ�����������������������������l���]���T���K���G�������www�'G_� n�� ��������������ҿ�ᜑ�3�3P3                       �ƶ�����������������������������|���N���R���I���a�������www�(d���������������׾��ҿ�ᜑ�3�3P3                       �Ƿ������������������Х���}��Ш�  ���8���I���`�������www�0t��������n����ݻ������ҿ�ᜑ�3�3P3                       �ʹ��������������ϧ�  �.|�u�/�;�Y�1�J�B���H���_�������www�0t���������������������ҿ�ᜑ�3�3P3                       �̹��������������ݛ�T�~��)���9�V�0�I�
���1�=�E���p�TRP���t����������������������ҿ�✑�3�3P3                       �ͻ����������ͧ�U�E�L�s�K�q�B�c�9�V�0�I�'�;��.�� �c�@�Kn7�㹏����������������������ҿ�✑�3�3P3                       �н�������������O�w�I�m�D�d�K�c�6�K� �0��&��� � � � ��ɗ����������������������ҿ�✑�3�3P3                       �Ѿ���������X���[��R�{�I�m��������jjj� ~ � � ���
�����Ԭ����������������������ҿ�✑�3�3P3                       ����������������f��P�x�G�k���������jjj��.��#������r��������������������������ҿ�⛐�3�3P3                       ��������������������D�f�F�j���������jjj�#�5��'���˭c������������������������������ҿ�⛏�3�3P3                       ��������������������S�y�G�h���������fff�>�:�-�8������������������������������������ҿ�⚏�5�4O3                       �����������������������������ʳ�zm`�QQQ����������������������������������������������ҿ�▊�8�:K6                       ����������������������������������������������������������������������������������������ە��>$�?&=D"                       ��������������������������������������������������������������������嶑��G��8�ދ6�Ղ5���c�H+`G+$@                         ��������������������������������������������������������������������������`���1���"�ɇG�`?,tQ1!/U3"U                          ���������������������������������������������������������������������Ǩ��΅���T�ϖ^�dC0sP0 0Z-@@@                           ���������������������������������������������������������������������Я��ؖ�ʕk�bA1uP5 0`@0@@@                               ���������������������������������������������������������������������Ѱ�ͬ��`B0�T9(:UG+@@@                                   �Ԫ��ڹ��׶��ִ��Գ��Ѳ��ϰ��̯��˭��ɬ��ƪ��é���������ᾥ�޻��۹��ಓ�㻢                                    �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  � �(                                             373x2�3�3�3�3�3�3�3�3�2�3x37        �{n�٭��֨��Ӧ��Ҥ��̡��ɞ��Ɯ��ę��������������3�4J        ��r����������������������ݻ��ڵ��װ��Ԫ��ҥ��3�4O        ��u��������������������������Ӫ��ԫ��װ��Ԫ�￨�3�3P        y������������������ҽ��~�W��ۚZ�ɞx��Ө�����3�3P        ȕ|�����������������O���h��6���z��u�����ï�3�3P        Ϝ������������������;���E���E������
���{����ű�3�3P        բ������������������U���e�������{����������ȵ�3�3P        ܩ����������7��K�7��_�Z�������7���1��������ɷ�3�3P        ܩ��������}�M�t�;�Y�+�A��'�Uz;��ض����������̺�3�3P        ܩ������V��N�v��Ч�"~%��
����������������ͽ�5�5M        ܩ����������L�r�����=�F����̑��������������ɺ�: �="C        ܩ������������������������������������������xl�B(tH'.        ܩ��������������������������������C���C��@�G+�N. HY7!        ܩ������������������������������ܩ���v�iH3�O3$dS7"%U9	        ܩ��ܩ��ܩ��ܩ��ܩ��ܩ��ޫ��֣��ܩ��٩�-                �   �   �   �   � ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ���n�$ Form1 . 5<   Y     �  D F�*    Command1  Command1 8�w �2    List0 - - '  '   �� Small Fonts�2    List1 �- '  '   �� Small Fonts�2    List2 �-   '   �� Small Fonts�2    List3 7- �   '   �� Small Fonts�    Timer1 �	  #  N  �   l�@     ��������     �@ �@    �             �y@   l�@     ��������    ��@ ,�@    X�             z@   l�@     ��������    P�@ P�@     �             Lz@ P   ���d�J�F����R��                                          Gd      \@ '�    ��@    ��@    ��@    t�@    ̈@    ��@    P�@    �@    ć@    ��@    ��@ VB5!�*             ~              	          P|@ �0  ���         �   Lz@ �y@ @ h   o   v   w   Mscomm MsConn  mscomm     l�@     �@ ����    ��@ <�@    �~             �{@     �@     �{@    �{@     �{@    �{@      |@ ��@     < �@ d�@ @  4    �@ ����         |@ ,	 0�@ ����H|@     �{@ t{@ �@ �@ �@         �l$��  �SR     �  l�@     �@ ��@ H  �@ �@  �@ * \ A C : \ D o c u m e n t s   a n d   S e t t i n g s \ B e n \ D e s k t o p \ v 5 8 \ W i n - S p y \ W i n S p y 7 6 \ A n t i   S p y \ M s C o n n . v b p                                                                                                                                                                                                                                                                                                                                                                               �z@       l�@     Ȓ@ ����    ��@ �@    �-             @    D�@     @    @     @    @ 	 �h l $�@ (�@     4% T�@ d�@ @  @   t�@           H�@ � ��@   @  D   ��@           d�@ �  �@   @  H   �@           ̀@ � �@   @  L   ��@           (�@ � $�@   @  P   ��@           ��@ � ,�@   @  T   ��@           ��@ � 4�@   @  X   <�@ ����        `�@ � L�@ ������@ 	�@ �@ #�@ W�@ 0�@ =�@ J�@ d�@     @ �~@ �@ �@ �@ B�@     4@ �~@ �@ �@ �@                                                                                     \@ �~@ �@ �@ �@ (�@                                                                     �@ �~@ �@ �@ �@                                                                                     �@ �~@ �@ �@ �@                                                                                     �@ �~@ �@ �@ �@                                                                                     �@ �~@ �@ �@ �@                         5�@                                                                                                 �l$��  �  �l$��  ��  �l$��  �5  �l$��  ��  �l$G   �  �l$W   �  �l$?   �!  �l$��  ��0  �l$��  �74         p�@ H�@ ����    `�@ �O�磶I���:)
    ��@             �@ 	  	         �~@ ����(�@             �@ 
   ��@ ��  ��     �y@ �����@     4�@     ��@        ��  �     �y@ ������@     $�@     �@        ��  �     z@ ������@     X�@     �@        ��  �     t{@ ����܋@             �@    ؄@ ��  �         ��@ ̆@ ܆@ �@ ��@  �@ �@ �@         ԋ@     mscomm  frmKillAntiSpy  modKillProcess  modMisc vb6To5  System  Class1         �s�Է��B�����!ԇ��&�"vN�����̾��d�J�F����R���X�z�OE�H4BE�s�*O�3�f�� � `ӓTimer1  .=����h�8 +3q�C:\program files\DevStudio\VB\VB5.OLB   VB  ��@        	   ��@ ą@ d�@         p� O�3�f�� � `ӓList1   �N�3�f�� � `ӓCommand1    List0   List2   List3   :O�3�f�� � `ӓForm       Kernel32.dll       RegisterServiceProcess  X�@ l�@    h�@ �p�@ �t��h��@ �0@ ����   CheckRunningProcess_SystExe StripFileName   Split   ReadUntil   Command1_Click  Form_Load   Timer1_Timer    GoStealth    d        4  <   ,   (4$ 
   $   	   kernel32       GetWindowsDirectoryA    X�@ h�@    t�@ �|�@ �t��h��@ �0@ ����      GetSystemDirectoryA X�@ ��@    ��@ ���@ �t��hć@ �0@ ����      CreateToolhelp32Snapshot    X�@ �@    ��@ ���@ �t��h�@ �0@ ����      Process32First  X�@ @�@    ��@ ���@ �t��hP�@ �0@ ����      Process32Next   X�@ ��@    ��@ ���@ �t��h��@ �0@ ����      CloseHandle X�@ ��@    ��@ ���@ �t��ḧ@ �0@ ����             T e x t        s y s t 3 2 . e x e        \              c a l c . e x e        OpenProcess +Z��J�Wj��~X�@ X�@    ��@ ���@ �t��ht�@ �0@ ����      TerminateProcess    X�@ ��@    ��@ ���@ �t��h��@ �0@ ����   ,          !cu��I s <�@ Settings   1   #=����h�8 +3q�"=����h�8 +3q�   �@  �@     yO�3�f�� � `ӓ   \ z i p l o g . t x t   O�3�f�� � `ӓ
       -       <   F o u n d   a n d   C l e a n e d   A n t i - S p y   :            \ s l o g . d l l       � +=����h�8 +3q����;�N�N)�q��*=����h�8 +3q�!=����h�8 +3q�Class   P�gv���3 +3oVBInternal  8�@        	       H�@ ��@         p�     � 4 
 �? �      GetVersionExA   X�@ ��@    ��@ ���@ �t��h��@ �0@ ����   WinVer   @         .   O p e r a t i n g   S y s t e m           =        * W i n d o w s   N T *        * W i n d o w s   9 *      ,   VBA5.DLL    __vbaAryUnlock  __vbaStrVarVal  __vbaVarIndexLoadRefLock    __vbaLineInputVar   __vbaStrLike    __vbaStrCat __vbaI2Var  __vbaStrToAnsi  __vbaWriteFile  __vbaFileOpen   __vbaFileClose  __vbaVarCat __vbaFreeObjList    __vbaObjSet __vbaVarAdd __vbaEnd    __vbaFreeObj    __vbaNew2   �@ ��@ __vbaStrToUnicode   __vbaLsetFixstr __vbaOnError    __vbaFixstrConstruct    __vbaVarForNext __vbaVarForInit __vbaLenBstr    __vbaFpI4   __vbaR8Str  __vbaInStr  __vbaStrI4  __vbaErrorOverflow  __vbaAryDestruct    __vbaGenerateBoundsError    __vbaRedimPreserve  __vbaVarCopy    __vbaStrCmp __vbaRefVarAry  __vbaUbound __vbaVarIndexLoad   __vbaStrCopy    __vbaVarMove    __vbaFreeStrList    __vbaFreeVarList    __vbaVarTstEq   __vbaFreeStr    __vbaHresultCheckObj    __vbaLateMemCallLd  __vbaStrVarMove __vbaStrMove    __vbaFreeVar    __vbaObjVar __vbaStrFixstr  __vbaLateMemSt  __vbaRecAnsiToUni   __vbaRecUniToAnsi   __vbaSetSystemError __vbaI4Var  __vbaRedim  �fĤ�I�x � 8<�__vbaExitProc   __vbaLbound __vbaI2I4      W i n d o w s          .      W i n d o w s   9 5        W i n d o w s   N T     __vbaStrI2          |�@     ,�@ ��@     ��@ �@ ��@    �@        ��@ ��@ ȓ@                     ��@ ��@ ��@ ȓ@     Ȓ@ �������������@    D�@    ����                 `��@                ���       `А@             00           `��@                  $        `��@                ���        `��@             /  	��       `��@             /    ��        `ؐ@             &&0��  <�@  `�@             ���/  ��  �@  `��@             00�0       �@ x�@ P�@ x�@ ��@ ��@ T�@ �@         �~@ ����           ��@     �@ ��@ ��@             d          t{@ ����           Ȑ@     ��@ ��@ Đ@             @         l�@ ����    (�@     p�@     ����    MsComm  ȅ@ t�@ ��@ ȅ@ ��@ ��@ ȅ@ �@ ��@ ȅ@ <�@ ��@ FilePath    sIn sDelim  nLimit  bCompare    T�@  �@ ��@ intMajor    intMinor    strPlatform ����������������������������U���h�@ d�    Pd�%    ��  �ESVW��e�3��E� @ P�u��������Q��   3�������V�J   ������J   �������Ej�u܉uԉ�������������������|�����l�����\�����L����0�Z�����@ ���Ӄ���u��c  �����������QRh<�@ ǅ����(  ���@ PV�Z������Ӎ����������PQh<�@ ��@ �$�@ �5��@ ����  ������Rh  �L�@ ���   �ԉ�|���������h�@ �
�������J������Q�B�������B��P�Ӌ=��@ ��|�����j ������h�@ R��P��|���P�8�@ ��P���@ �Ѝ������D�@ �E������������Q������RP���  ��}�Uh�  hd�@ RP��@ �������M�ǅ����    �D�@ �������\�@ ��|����׃��EԋԹ   ��L�����T����
��P���h�@ �J������Q�B��X����B��P��j ������h�@ R��P��|���P�8�@ ����l���PQ�P�@ ��l�����L���RPǅT����@ ǅL����  �x�@ ��l�����|���QRj�����@ ��f��uX������������PQh<�@ ���@ �U�PR��������@ ������������PQh<�@ ��@ ������U�R������@ h��@ �I�E�t	�M����@ ������������PQj��@ ����\�����l�����|���RPQj���@ ��ÍM��\�@ �������%��@ ËEP��R�E�M܋U�_��M�^[�P�U�H�M�P�E�d�    ��]� ��U���h�@ d�    Pd�%    ��LSVW�}�e�3���E�@ W�u��S�E�u��u��0�@ �Mԉu܉u؉uԉuĉ0�u��E������ �@ �MčU�QR�U�E�P�MԋQPW��   ;�}h   hd�@ WP��@ �UčM����@ �M��\�@ �M�Q�T�@ �Rj���@ ���   ��j�
�M��J�M�Q�B�E��B�U�R�H�@ ��P���@ �ЍM��D�@ �M����@ h�@ �"�E�t	�M��\�@ �M��\�@ �M����@ ÍM��%��@ ËEP��Q�U�E؋M�_��E�^d�    [��]� ����������U���h�@ d�    Pd�%    ��PS�]VW�3�e�3��E� @ S�}��V�U3��M��}�}�}��}ЉEȉE��E�� �@ �E�M�8�Rh8�@ �p�@ ��u�E��U��MЉE��E�   �0�@ �U�E��  �M�QR�M�PQS�u��օ�}h  hd�@ SP��@ �UȍM��E�    �D�@ ��j Vj�U�j Rjh   ���@ �M����t$f�9u�Q�A+�;�r	�l�@ �M��    �	�l�@ �M�I�U��� �@ �EfG�\  � 3���;���3Ƀ�����tU�M�UȍE�RP�U�Q3�RS�u��U�;�}h  hd�@ SP��@ �UȍM�u��D�@ �E�Ph8�@ �p�@ ���(�����j Vj�M�j Qjh   ���@ �M����t$f�9u�Q�A+�;�r	�l�@ �M��    �	�l�@ �M�I�U��� �@ �U�MЉU��U��E�   �0�@ h��@ ��E�t	�M����@ �M��\�@ Ë5\�@ �M��֍E�Pj � �@ �M���ËEP��Q�U�EЋM�_��E�^[�J�M܉B�E��J�M�d�    ��]� ���@ �U���h�@ d�    Pd�%    ��d�ESVW��e�3��E�@@ P�u��Q�U�M�u�u�uԉuĉu��2�u�j�P�ER�Q���@ P���@ �=D�@ �ЍM��׋U�R���@ �0@ ����A��   �E�u�P�E�@  ���@ �%8@ �4�@ ���	  �ӍM�P�U�QR�<�@ �E�P���@ �ЍM��׍M����@ �U�M�QR�E� ��E�
   �u��E�@  ���@ �E�]��Q���@ �E��E��]��E��E�����   ��P�U��E�RP�\�@ �M�Q���@ �Ћ��׍UčE�RPj���@ ���h��@ �#�E�t	�M��\�@ �MčU�QRj���@ ��ÍM��%\�@ ËEP��Q�U�E�M�_��E�^d�    [��]� ��t������U���h�@ d�    Pd�%    ��p�ES��V$�W�   �e�#��E�P@ P�M��E�R3��M��E܉E؉EȉE��E��E��E��   �EȉE��E��E�P�U�Q�E�R�M�P�U�QR�u��E��  �u��0�@ �5 �@ �=\�@ �T�@ ��t(�@�@ �M��֍E�P�%  �M��׍M��U�Q�E�RP�����E�    hƞ@ �
�M��\�@ ÍM��U�QRj���@ ���M��%��@ ËEP��Q�M�E�_^d�    [��]� �����������U���h�@ d�    Pd�%    ��   �s��SVW�e��E�`@ �E���E��M����M�E�    �U��MQ�P�E�   �U�Rh�   ���@ �E�   j��4�@ �E�   �E�P���@ P�M�Q�U�R�(�@ P� �����L�����@ �E�P�M�Q���@ P�U�Rj ��@ ��L����E��M�Q�U�Rj��@ ���E�   �U��M�� �@ �E���\���ǅT���@  �M�Q��T���R��t���P�<�@ �M�Q�U�Rj ��@ ��t����M����@ �M��\�@ �E�   �E�P���@ P�M�Q�U�R�(�@ P�u�����L�����@ �E�P�M�Q���@ P�U�Rj ��@ ��L����E��M�Q�U�Rj��@ ���E�   �U��M�� �@ �E���\���ǅT���@  �M�Q��T���R��t���P�<�@ �M�Q�U�Rj ��@ ��t����M����@ �M��\�@ �E�   �=��@  uh��@ h0�@ ���@ ǅ �����@ �
ǅ �����@ �� ������H����U�R��H������H���R�Q��D�����D��� }#jh �@ ��H���P��D���Q��@ ������
ǅ���    �U���@�����P���P��@������@���P�Rh��<�����<��� }#jhh@�@ ��@���Q��<���R��@ ������
ǅ���    3�f��P��������f��8����M��`�@ ��8�����t�E�   ���@ �E�
   �U�R��t���P�P�@ ǅ\���T�@ ǅT���   ��t���Q��T���R��d���P�$�@ P���@ �ЍM��D�@ ��d���Q��t���Rj���@ ���E�   �Ẻ�\���ǅT���@  j��T���Q���@ ��|���ǅt���   ��t����M����@ �E�   ǅ\���8�@ ǅT����  �U�R��T���P�x�@ �ȅ�t�E�   ���@ �E�   ��t���R�E��UR��  ��H�����H��� }#h  hd�@ �EP��H���Q��@ ������
ǅ���    ��t������@ �E�   ��t���R�E�P�M��EP��  ��t������@ �E�    h:�@ �6�M�Q�U�Rj��@ ���M��`�@ ��d���P��t���Qj���@ ��ÍM����@ �M��\�@ �M����@ �M����@ �M����@ �M��\�@ ËU��MQ�P�E��M�d�    _^[��]� ����U���h�@ d�    Pd�%    �\  �n��SVW�e��E��@ �E���E��M����M�E�    �U��MQ�P�E�   �U�Rh�   ���@ �E�   j��4�@ �E�   �E�P���@ P�M�Q�U�R�(�@ P������ �����@ �E�P�M�Q���@ P�U�Rj ��@ �� ����E��M�Q�U�Rj��@ ���E�   �U��M�� �@ �E��� ���ǅ���@  �M�Q�����R��h���P�<�@ �M�Q�U�Rj ��@ ��h����M����@ �M��\�@ �E�   �E�P���@ P�M�Q�U�R�(�@ P������ �����@ �E�P�M�Q���@ P�U�Rj ��@ �� ����E��M�Q�U�Rj��@ ���E�   �U��M�� �@ �E��� ���ǅ���@  �M�Q�����R��h���P�<�@ �M�Q�U�Rj ��@ ��h����M����@ �M��\�@ �E�   ǅp��� �ǅh���
   ��h���P���@ f�����ǅ���   ������M����@ ��h������@ �E�   �M��EP��  P��|���Q�8�@ �����������R�������������R���   ������������ }&h�   hl�@ ������P������Q��@ �������
ǅ����    f�����f������fǅ���� f�E�  ��|����`�@ �f�E�f�������  f�E�f�M�f;�������  �E�	   �U��MQ��   P��|���R�8�@ ������f�E�P�������������P���   ������������ }&h�   hl�@ ������Q������R��@ �������
ǅ����    ��|����`�@ �E�
   �E��UR��  P��|���P�8�@ ������f�M�Q�������������Q���   ������������ }&h�   hl�@ ������R������P��@ �������
ǅ����    ��|����`�@ �E�   �M��EP��  P��|���Q�8�@ ������f�U�R�������������R���   ������������ }&h�   hl�@ ������P������Q��@ �������
ǅ����    ��|����`�@ �E�   �U��MQ��  P��|���R�8�@ ������f�E�P�������������P���   ������������ }&h�   hl�@ ������Q������R��@ �������
ǅ����    ��|����`�@ �E�   �E��UR��  P��x���P�8�@ �������M��EP��  P��|���Q�8�@ �����������R�������������R���   ������������ }&h�   hl�@ ������P������Q��@ �������
ǅ����    �U�Rf�����P�������������P���   ������������ }&h�   hl�@ ������Q������R��@ �������
ǅ����    �E��������E�    �������M��D�@ �M�Q�  �ЉU��M��\�@ ��x���P��|���Qj���@ ���E�   �}����  �E�   ��h���R� �@ ǅ �����@ ǅ���   ǅ�����@ ǅ���   �E��UR��   P��x���P�8�@ �������M��EP��   P��|���Q�8�@ �����������R�������������R���   ������������ }&h�   hl�@ ������P������Q��@ �������
ǅ����    �U�Rf�����P�������������P���   ������������ }&h�   hl�@ ������Q������R��@ �������
ǅ����    �E��������E�    ��������@���ǅ8���   ��h���R�����P��X���Q���@ P�����R��H���P���@ P��8���Q��(���R���@ �ЍM����@ ��x���P��|���Qj���@ ����8���R��H���P��X���Q��h���Rj���@ ���E�   ǅ ���Ԋ@ ǅ���   �E�P�����Q��h���R�$�@ P���@ �ЍM��D�@ ��h������@ �E�   j�d�@ �E�   �E�Pjj�j���@ �E�   �M�Q�U�R���@ Ph�@ ��@ ���E�   j�d�@ �E�   �E��UR��  P��x���P�8�@ �������M��EP��  P��|���Q�8�@ �����������R�������������R���   ������������ }&h�   hl�@ ������P������Q��@ �������
ǅ����    �U�Rf�����P�������������P���   ������������ }&h�   hl�@ ������Q������R��@ �������
ǅ����    �E��������E�    �������M��D�@ �M�Q�  �ЉU��M��\�@ ��x���P��|���Qj���@ ���E�   �}����  �E�   ��h���R� �@ ǅ �����@ ǅ���   ǅ�����@ ǅ���   �E��UR��   P��x���P�8�@ �������M��EP��   P��|���Q�8�@ �����������R�������������R���   ������������ }&h�   hl�@ ������P������Q��@ �������
ǅ����    �U�Rf�����P�������������P���   ������������ }&h�   hl�@ ������Q������R��@ �������
ǅ����    �E��������E�    ��������@���ǅ8���   ��h���R�����P��X���Q���@ P�����R��H���P���@ P��8���Q��(���R���@ �ЍM����@ ��x���P��|���Qj���@ ����8���R��H���P��X���Q��h���Rj���@ ���E�   ǅ ���Ԋ@ ǅ���   �E�P�����Q��h���R�$�@ P���@ �ЍM��D�@ ��h������@ �E�   j�d�@ �E�   �E�Pjj�j���@ �E�   �M�Q�U�R���@ Ph�@ ��@ ���E�   j�d�@ �E�   �E��UR��  P��x���P�8�@ �������M��EP��  P��|���Q�8�@ �����������R�������������R���   ������������ }&h�   hl�@ ������P������Q��@ �������
ǅ����    �U�Rf�����P�������������P���   ������������ }&h�   hl�@ ������Q������R��@ �������
ǅ����    �E��������E�    ��������p���ǅh���   ��h���R�t�@ ��x���P��|���Qj���@ ����h������@ �E�    �&����E�    h��@ �[�U�R�E�Pj��@ ����x���Q��|���Rj���@ ����(���P��8���Q��H���R��X���P��h���Qj���@ ��ÍM��\�@ �M����@ �M����@ �M����@ �M����@ �M��\�@ ËU��MQ�P�E��M�d�    _^[��]� ���@ ��U���h�@ d�    Pd�%    ��   �]^��SVW�e��E�p@ �E�    �E�    �E��UR�Q�E�   �E�     �E�   j��4�@ �E�   j���@ �ЍM��D�@ Pj
���@ �ЍM��D�@ P��@ �E��E�   �U��M����@ �M�Q�U�Rj��@ ���E�   �E�x4 u �M��4Qht{@ ���@ �U��4��h�����E��4��h�����h�����U��E��<P�M��:Q�U��8R�E���U�R�Q�E��}� }jhd�@ �E�P�M�Q��@ ��d����
ǅd���    �E�   h�@ �U�B<P��@ �E��E�   �M�Q�U�R�E�P�$�@ P���@ �ЍM��D�@ �M�Q�U�Rj���@ ���E�   �E�Ph �@ �<�@ �ȅ���   �E�   �=��@  uh��@ h0�@ ���@ ǅ`�����@ �
ǅ`�����@ ��`�����E��M�Q�U���M�Q�P�E��}� }jh �@ �U�R�E�P��@ ��\����
ǅ\���    �M��M�j �U���M�Q�P|�E��}� }j|h@�@ �U�R�E�P��@ ��X����
ǅX���    �M��`�@ �E�	   �M�Qh@�@ �<�@ �Ѕ�t�E�
   jj ������@ hX�@ �C�E�����t	�M����@ �M�Q�U�Rj��@ ���M��`�@ �E�P�M�Qj���@ ��ÍM��\�@ �M����@ ËU��MQ�P�U�E���M��J�EĉB�MȉJ�E��M�d�    _^[��]� ������������U���h�@ d�    Pd�%    ��   ��Z��SVW�e��E��@ �E�    �E�    �E�   �E�     �E�   �M��EP��   P�M�Q�8�@ ��@�����@������@���Q���  ��<�����<��� }&h�  hl�@ ��@���R��<���P��@ �� ����
ǅ ���    �M��`�@ �E�   �M��EP��  P�M�Q�8�@ ��@�����@������@���Q���  ��<�����<��� }&h�  hl�@ ��@���R��<���P��@ ������
ǅ���    �M��`�@ �E�   �M��EP��  P�M�Q�8�@ ��@�����@������@���Q���  ��<�����<��� }&h�  hl�@ ��@���R��<���P��@ ������
ǅ���    �M��`�@ �E�   �M��EP��  P�M�Q�8�@ ��@�����@������@���Q���  ��<�����<��� }&h�  hl�@ ��@���R��<���P��@ ������
ǅ���    �M��`�@ �E�   j��4�@ �E�   �E� ��E�
   �M�Q���@ f��T���ǅL���   ��L����M����@ �M����@ �E�   �U�R���@ P�d�@ �E�	   �E�Q�U�R���@ Pj�j���@ �E�
   �E�P���@ P���@ �ȅ���  �E�   �U�R���@ P�E�P���@ �E�   ǅd���8�@ ǅ\����  �M�Q��\���R�x�@ ����t�P  �E�   ǅd���    ǅ\���   ǅD���   ǅH��������\�@ �M�� �@ �M�Q��D���R��H���P�M�Q�U�R�E�P���@ P�M��EP��   ��@�����@��� }#h   hd�@ �MQ��@���R��@ ������
ǅ���    �   ��V���ċ�\������`����P��d����H��h����Pj�E�P�M�Q��|���R�(�@ �� P��l���P�P�@ �M�Q�P�@ �U��MQ��   P�U�R�8�@ ��<���ǅT��� �ǅL���
   �   �NV���ċ�L������P����P��T����H��X����P��l���P�M�Q���@ P��<������<���Q���  ��8�����8��� }&h�  hl�@ ��<���R��8���P��@ ������
ǅ���    �M�Q�U�R�E�Pj��@ ���M��`�@ ��l���Q��|���R�E�Pj���@ ���E�   ǅd���   ǅ\���   ǅD���   ǅH��������\�@ �M�� �@ �M�Q��D���R��H���P�M�Q�U�R�E�P���@ P�M��EP��   ��@�����@��� }#h   hd�@ �MQ��@���R��@ ������
ǅ���    �   ��T���ċ�\������`����P��d����H��h����Pj�E�P�M�Q��|���R�(�@ �� P��l���P�P�@ �M�Q�P�@ �U��MQ��  P�U�R�8�@ ��<���ǅT��� �ǅL���
   �   �:T���ċ�L������P����P��T����H��X����P��l���P�M�Q���@ P��<������<���Q���  ��8�����8��� }&h�  hl�@ ��<���R��8���P��@ ������
ǅ���    �M�Q�U�R�E�Pj��@ ���M��`�@ ��l���Q��|���R�E�Pj���@ ���E�   ǅd���   ǅ\���   ǅD���   ǅH��������\�@ �M�� �@ �M�Q��D���R��H���P�M�Q�U�R�E�P���@ P�M��EP��   ��@�����@��� }#h   hd�@ �MQ��@���R��@ �� ����
ǅ ���    �   �R���ċ�\������`����P��d����H��h����Pj�E�P�M�Q��|���R�(�@ �� P��l���P�P�@ �M�Q�P�@ �U��MQ��  P�U�R�8�@ ��<���ǅT��� �ǅL���
   �   �&R���ċ�L������P����P��T����H��X����P��l���P�M�Q���@ P��<������<���Q���  ��8�����8��� }&h�  hl�@ ��<���R��8���P��@ �������
ǅ����    �M�Q�U�R�E�Pj��@ ���M��`�@ ��l���Q��|���R�E�Pj���@ ���E�   ǅd���   ǅ\���   ǅD���   ǅH��������\�@ �M�� �@ �M�Q��D���R��H���P�M�Q�U�R�E�P���@ P�M��EP��   ��@�����@��� }#h   hd�@ �MQ��@���R��@ �������
ǅ����    �   �P���ċ�\������`����P��d����H��h����Pj�E�P�M�Q��|���R�(�@ �� P��l���P�P�@ �M�Q�P�@ �U��MQ��  P�U�R�8�@ ��<���ǅT��� �ǅL���
   �   �P���ċ�L������P����P��T����H��X����P��l���P�M�Q���@ P��<������<���Q���  ��8�����8��� }&h�  hl�@ ��<���R��8���P��@ �������
ǅ����    �M�Q�U�R�E�Pj��@ ���M��`�@ ��l���Q��|���R�E�Pj���@ ���4����E�   �M�Q���@ P�d�@ h��@ �[�U�����t	�M����@ �E�P�P�@ �M�Q�U�R�E�Pj��@ ���M��`�@ ��l���Q��|���R�E�Pj���@ ��ÍM����@ �M����@ ËM�UЉ�EԉA�U؉Q�E܉A3��M�d�    _^[��]� ���������U���h�@ d�    Pd�%    ��t  SVW��   3��������J   �������3��e��J   ������Vj��E�8@ �u���������������������������������������������������������t�����d�����T�����D�����4�����$���������������8�����@ ���Ӎ�����������PQh<�@ �}�ǅ����(  ���@ PW�A����������Ӎ�����������RPh<�@ ��@ VVjVh4�@ h,  V���@ ��@ �5D�@ �=L�@ �����������]  ������Qh  �׋Ѝ������֍�����R��  �Ѝ������֋�����������PQh  �Ӌ�����������RPh  �Ӎ�����������QRj��@ ��j ���@ �Ѝ�������j ���@ �Ѝ������֋�����������j3�Rh  ��|���ǅt���   �������������׋Ѝ������֋�����P��������Pj ���@ H�������  ������������jQh  ǅ����   ������ǅ����    �׋Ѝ������֋�����P��������Pj ���@ 3ҍ����������ڍ�t���f�����P�����Q��d���RPǅ���   ��@ ��d���Q��@ ������PRh  �׋Ѝ�������P�,�@ �Ѝ������֋�����������PQh  �Ӌ�������T�����\�����D���RPǅ����    ǅT���   � �@ �M��������4���RP������ǅ����@  � �@ ��D�����4���QR�x�@ ������������������P������Q������R������P������Q������RPj��@ �� ��4�����D���Q��T���R��d���P��t���Q������R�����PQj���@ �� f������ uM������������RPh<�@ ���@ �M�PQ�;�����������@ ������������RPh<�@ ��@ �����������Qj�h� ������=�@ ����j V��������V������3�hp�@ �����ډU��   �E�P�������@ hp�@ �   ������������Q������R������P������Q������R������P������QRj��@ ��$��$�����4�����D���PQ��T���R��d���P��t���Q������RPj���@ �� �ËM�f�E�_^d�    [��]� ���@ ���U���h�@ d�    Pd�%    ��HSVW3��0�@ �Mԉe��E�H@ �E܉E؉EԉEĉE��E������ �@ �E��M�P�E�U�Q�R�U�QR��   �UčM����@ �M��\�@ �E�P�T�@ �Qj���@ ���   ��j�
�M��J�M�Q�B�E��B�U�R�H�@ ��P���@ �ЍM��D�@ �M����@ h��@ �"�E�t	�M��\�@ �M��\�@ �M����@ ÍM��%��@ ËM�E�_^d�    [��]� ����������U���h�@ d�    Pd�%    ��<�USVW3��M�e��E�X@ �}�}�}�}ԉ}��}�� �@ �u�Ph8�@ �p�@ ��u�M�U��MȍM��E�   �0�@ �U�E�RVP�  �ЍM��D�@ ���@ ��j Vj�M�j Qjh   �ӋM����t$f�9u�Q�A+�;�r	�l�@ �M��    �	�l�@ �M�I�U��� �@ �UfG�$  �3���;���3Ƀ�����t:�E�U�R�M�PQ�E�    �  �ЍM��D�@ �U�Rh8�@ �p�@ ���G�����j Vj�E�j Pjh   �ӋM����t$f�9u�Q�A+�;�r	�l�@ �M��    �	�l�@ �M�I�U��� �@ �M�U��MȍM��E�   �0�@ h��@ �
�M����@ Ë5\�@ �M��֍U�Rj � �@ �M���ËE�Uԋ�_^[��U؉Q�U܉Q�U��Q�M�d�    ��]� ���@ ���������U���h�@ d�    Pd�%    ��d�MSV�u3��W�E�E�EԉEĉE���e�jP�ER�E�x@ �Q���@ P���@ �=D�@ �ЍM��׋U�R���@ �h@ ����A��   �E�u�P�E�@  ���@ �%p@ �4�@ ����   �ӍM�P�U�QR�<�@ �E�P���@ �ЍM��׍M����@ �U�M�QR�E� ��E�
   �u��E�@  ���@ �E�]��Q���@ �E��E��]��E��E���u��P�U��E�RP�\�@ �M�Q���@ �Ћ��׍UčE�RPj���@ ���h{�@ �#�E�t	�M��\�@ �MčU�QRj���@ ��ÍM��%\�@ ËM�E�_^d�    [��]� �D������������U���h�@ d�    Pd�%    ���  �ESVW��e�3��E��@ P�]��Q�E   3��������������%   ��0���󫍅0���RPh|�@ ������������������������ǅ�����   ���@ P聼������@ ��0���������QRh|�@ ��@ ;���   �������5|�@ �֋}������f��֋Mf�������+�tHtH��   ���@ �   �|�@ �   f����@ h\�@ R�Ӌ5D�@ �Ѝ������֋=�@ P�׋Ѝ�������Pht�@ �׋Ѝ�������P�Ef�Q�ӋЍ�������P�׋M���֍�����������R������P������QRj��@ ����E�M�8�@ f�f��M� �@ h��@ �(������������R������P������QRj��@ ���ËEP��Q�M�E�_^d�    [��]� ����                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                            (�  ��������h�  ��                      v�  ��  ��  ��  ��  ��  ��  ��  ��   �  �  �  0�  D�   �R�  f�  t�  ��  ��  ��  ��  ��  ��  ��  �  (�  :�  J�  X�  h�  z�  ��  ��   ���  ��  x ���  ��  ��  �  �   �,�  <�  H�  V�  h�  v�  ��  ��  ��  ��  ��  ��  ��  �  &�  :�  H�  Z�  n�  |�  ��  ��   �� ���  ��  ��  ��  ��  ��  � �; ��  �  &�  � �6�  J�  \�  � �d  �j�  b �x�  ��  h ���  ��  ��  i ���  ��  ��  ��  ��  
�  �  &�  6�      �)/v��1v�<v#>vϾ/v��=v�b0v��.v+>v>�1vUx<v�O0v�;v�~<vy�1v�5;v� .vȥ1v�e;v��3v�0v	x<v��/v.2>v�9;v�0v�3>vR�/v��/v�<v�x<v�y<v��/v<v<�;vJ�/v��1vn02v�/v��/v�)0v�9;v��/v*'/v��>vݿ/v61v��2v�/vV*2v�<v>�1v�/v�5;v�1v�B1vJc1vY+0v�:v$|<vUy<v��>vr�/v%�3v$K.vڹ/v�/v�2v�B1v;v�(.v��.vԌ;v��/v�6.v9~;v�x<v�y<v��/v>�/v��/v	y<vDs<v�.v��.v��/v.�/v�>vC�:vx#/v�>v�/>v�$>vĸ.v�B1v��/ve�<v[�<v��3v�4>v��/vx�/v�/v    MSVBVM50.DLL    __vbaStrI2    _CIcos    _adj_fptan    __vbaVarMove    __vbaStrI4    __vbaFreeVar    __vbaStrVarMove   __vbaLenBstr    __vbaFreeVarList    __vbaEnd    _adj_fdiv_m64   __vbaFreeObjList    __vbaLineInputVar   _adj_fprem1   __vbaRecAnsiToUni   __vbaStrCat   __vbaLsetFixstr   __vbaWriteFile    __vbaSetSystemError   __vbaHresultCheckObj    _adj_fdiv_m32   __vbaAryDestruct    __vbaLateMemSt    __vbaVarIndexLoadRefLock    __vbaExitProc   __vbaVarForInit   __vbaOnError    __vbaObjSet   __vbaStrLike    _adj_fdiv_m16i    _adj_fdivr_m16i   __vbaVarIndexLoad   __vbaStrFixstr    __vbaRefVarAry    _CIsin    __vbaChkstk   __vbaFileClose    EVENT_SINK_AddRef   __vbaGenerateBoundsError    __vbaStrCmp   __vbaVarTstEq   __vbaI2I4   __vbaObjVar   DllFunctionCall   __vbaLbound   __vbaRedimPreserve    _adj_fpatan   __vbaFixstrConstruct    __vbaRedim    __vbaRecUniToAnsi   EVENT_SINK_Release    _CIsqrt   EVENT_SINK_QueryInterface   __vbaExceptHandler    __vbaStrToUnicode   _adj_fprem    _adj_fdivr_m64    __vbaFPException    __vbaUbound   __vbaStrVarVal    __vbaVarCat   __vbaI2Var    _CIlog    __vbaErrorOverflow    __vbaFileOpen   __vbaInStr    __vbaR8Str    __vbaNew2   _adj_fdiv_m32i    _adj_fdivr_m32i   __vbaStrCopy    __vbaFreeStrList    _adj_fdivr_m32    _adj_fdiv_r   __vbaI4Var    __vbaVarAdd   __vbaStrToAnsi    __vbaVarCopy    __vbaFpI4   __vbaLateMemCallLd    _CIatan   __vbaStrMove    _allmul   _CItan    __vbaAryUnlock    __vbaVarForNext   _CIexp    __vbaFreeStr    __vbaFreeObj                                                                                                                                                                                                �s�@��        X  �   @  �   (  �    �s�@��        �  �    �s�@��        �  �    �s�@��    	 1u  � �2u  � �3u  p �4u  X �5u  @ �6u  ( �7u   �8u  �  �9u  �  �    �s�@��     	  �      �s�@��         �      �s�@��         �      �s�@��         �      �s�@��         �      �s�@��               �s�@��               �s�@��         (      �s�@��         8      �s�@��         H      �s�@��         X  p h  �      � �   �      \ h  �      �	 �  �      l �%  �      @ h  �      |E �  �      $N �  �      �\ (  �      �] �  �      �` h  �              h4   V S _ V E R S I O N _ I N F O     ���                                           D     V a r F i l e I n f o     $    T r a n s l a t i o n     	��   S t r i n g F i l e I n f o   �   0 4 0 9 0 4 B 0   (   C o m m e n t s   m s c o m m     0   C o m p a n y N a m e     m s c o m m     8   F i l e D e s c r i p t i o n     m s c o m m     0   P r o d u c t N a m e     M s C o n n     , 
  F i l e V e r s i o n     1 . 0 0     0 
  P r o d u c t V e r s i o n   1 . 0 0     0   I n t e r n a l N a m e   M s c o m m     @   O r i g i n a l F i l e n a m e   M s c o m m . e x e        	 00   h  1u     �  2u   (  3u00    �  4u      �  5u    h  6u00     �%  7u       �  8u     h  9u(                                             373x2�3�3�3�3�3�3�3�3�2�3x37        �{n�٭��֨��Ӧ��Ҥ��̡��ɞ��Ɯ��ę��������������3�4J        ��r����������������������ݻ��ڵ��װ��Ԫ��ҥ��3�4O        ��u��������������������������Ӫ��ԫ��װ��Ԫ�￨�3�3P        y������������������ҽ��~�W��ۚZ�ɞx��Ө�����3�3P        ȕ|�����������������O���h��6���z��u�����ï�3�3P        Ϝ������������������;���E���E������
���{����ű�3�3P        բ������������������U���e�������{����������ȵ�3�3P        ܩ����������7��K�7��_�Z�������7���1��������ɷ�3�3P        ܩ��������}�M�t�;�Y�+�A��'�Uz;��ض����������̺�3�3P        ܩ������V��N�v��Ч�"~%��
����������������ͽ�5�5M        ܩ����������L�r�����=�F����̑��������������ɺ�: �="C        ܩ������������������������������������������xl�B(tH'.        ܩ��������������������������������C���C��@�G+�N. HY7!        ܩ������������������������������ܩ���v�iH3�O3$dS7"%U9	        ܩ��ܩ��ܩ��ܩ��ܩ��ܩ��ޫ��֣��ܩ��٩�-                �   �   �   �   � ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ���n�(       @                                              3
874I4O3P3P3P3P3P3P3P3P3P3P3P3P3P3P3P3P3P4O4I373
++                        875x4�3�3�3�3�3�3�3�3�3�3�3�3�3�3�3�3�3�3�3�2�3x377                       Ϟ��ۧ��٦��ؤ��֣��֣��ԡ��Ӡ��ў��ѝ��ѝ��ѝ��ѝ��ѝ��Н��М��М��М��М��М��М��М��ޘ��3�4J9                       ͱ�����������������������������������������������������������������������������������̙�ᜐ�3�4O3                       ɲ�������������������������������������������޽��ݺ��۷��ڴ��ر��ׯ��֬��ԩ��ӧ��Ѥ��ҿ�ᜑ�3�3P3                       ̵�����������������������������������������������޽��ݺ��۷��ڴ��ر��ׯ��֬��ԩ��ӧ��ҿ�ᜑ�3�3P3                       η���������������������������������������������������޽��Ǖ��ȗ��ڴ��ر��ׯ��֬��ԩ��ҿ�ᜑ�3�3P3                       и�������������������������������������������˝�����ͼ��vku��^��۷��ٲ��Ɠ��֭��֬��ҿ�ᜑ�3�3P3                       Һ������������������������������������������Λn��h�H�� K����Q��y���u�ܣm��Ɠ��ׯ��ҿ�ᜑ�3�3P3                       Ӽ�������������������������������������� G��A��sej�8���4���Ja}�c\g� G��4U���Ï��ر��ҿ�ᜑ�3�3P3                       ־��������������������������������������V���2���P��;���2���n��[�����1����y��ɗ��ҿ�ᜑ�3�3P3                       ������������������������������������`t��T���M���D���;���2���*���!���������wnv��{��ҿ�ᜑ�3�3P3                       �³�����������������������������*h��`��Q���K���B���R���<���$���������k�� N��ͦ���ҿ�ᜑ�3�3P3                       �Ĵ�����������������������������l���]���T���K���G�������www�'G_� n�� ��������������ҿ�ᜑ�3�3P3                       �ƶ�����������������������������|���N���R���I���a�������www�(d���������������׾��ҿ�ᜑ�3�3P3                       �Ƿ������������������Х���}��Ш�  ���8���I���`�������www�0t��������n����ݻ������ҿ�ᜑ�3�3P3                       �ʹ��������������ϧ�  �.|�u�/�;�Y�1�J�B���H���_�������www�0t���������������������ҿ�ᜑ�3�3P3                       �̹��������������ݛ�T�~��)���9�V�0�I�
���1�=�E���p�TRP���t����������������������ҿ�✑�3�3P3                       �ͻ����������ͧ�U�E�L�s�K�q�B�c�9�V�0�I�'�;��.�� �c�@�Kn7�㹏����������������������ҿ�✑�3�3P3                       �н�������������O�w�I�m�D�d�K�c�6�K� �0��&��� � � � ��ɗ����������������������ҿ�✑�3�3P3                       �Ѿ���������X���[��R�{�I�m��������jjj� ~ � � ���
�����Ԭ����������������������ҿ�✑�3�3P3                       ����������������f��P�x�G�k���������jjj��.��#������r��������������������������ҿ�⛐�3�3P3                       ��������������������D�f�F�j���������jjj�#�5��'���˭c������������������������������ҿ�⛏�3�3P3                       ��������������������S�y�G�h���������fff�>�:�-�8������������������������������������ҿ�⚏�5�4O3                       �����������������������������ʳ�zm`�QQQ����������������������������������������������ҿ�▊�8�:K6                       ����������������������������������������������������������������������������������������ە��>$�?&=D"                       ��������������������������������������������������������������������嶑��G��8�ދ6�Ղ5���c�H+`G+$@                         ��������������������������������������������������������������������������`���1���"�ɇG�`?,tQ1!/U3"U                          ���������������������������������������������������������������������Ǩ��΅���T�ϖ^�dC0sP0 0Z-@@@                           ���������������������������������������������������������������������Я��ؖ�ʕk�bA1uP5 0`@0@@@                               ���������������������������������������������������������������������Ѱ�ͬ��`B0�T9(:UG+@@@                                   �Ԫ��ڹ��׶��ִ��Գ��Ѳ��ϰ��̯��˭��ɬ��ƪ��é���������ᾥ�޻��۹��ಓ�㻢                                    �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  � �(   0   `                                                          ++ 79333333333333333333331333333333397++                                            3
374I4O3P3P3P3P3P3P3P3P3P3P3P3P3P3P3P3P3P3P3P2Q3P3P3P3P3P3P3P3P3P4O4I373
++                                        373x2�3�3�3�3�3�3�3�3�3�3�3�3�3�3�3�3�3�3�3�4�3�3�3�3�3�3�3�3�3�3�3�2�3x377                                       �__��]]��\\��[[��ZZ��YY��XX��VV��TT��TT��SS��QQ��PP��PP��PP��PP��PP��PP��PP��PP��PP��PP��PP��PP��PP��PP��PP��PP��PP��PP��PP��OO��MM�LL��MM�3�4J9                                       �aa����������������������������������������������������������������������������������������������������������������������������������̙��OO�3�4O3                                       �aa��������������������������������������������������߿��޽��ܸ��ݺ��ܸ��۶��ڵ��ٲ��ر��ׯ��֭��լ��Ԫ��Ө��Ӧ��Ҥ��ѣ��С��ϟ��ʹ������PP�3�3P3                                       �bb������������������������������������������������������߿��޽��ݻ��ݺ��ܸ��۶��ڵ��ٲ��ر��ׯ��֭��լ��Ԫ��Ө��Ӧ��Ҥ��ѣ��С��Ͷ������SR�3�3P3                                       �dd����������������������������������������������������������߿��޽��ݻ��ݺ��ܸ��۶��ڵ��ٲ��ر��ׯ��֭��լ��Ԫ��Ө��Ӧ��Ҥ��ѣ��ζ������TS�3�3P3                                       �ee��������������������������������������������������������������߿��޽��ݻ��ݺ��ܸ��۶��ڵ��ٲ��ر��ׯ��֭��լ��Ԫ��Ө��Ӧ��Ҥ��η������UT�3�3P3                                       �ff������������������������������������������������������������������߿��޽��ݻ��ݺ��ܸ��۶��ڵ��ٲ��ر��ׯ��֭��լ��Ԫ��Ө��Ӧ��ϸ������WV�3�3P3                                       �ig����������������������������������������������������������������������߿��޽��q��k��k��լ��ڵ��ٲ��ر��ׯ��֭��լ��Ԫ��Ө��Ϲ������YW�3�3P3                                       �kh����������������������������������������������������������Ҩ��˝���������Ŷ��vhr�ʓb��\��ҩ��۶��ڵ��͟��ɗ��׮��֭��լ��Ԫ��к������YX�3�3P3                                       �nj������������������������������������������������������޿���w��k��o�̼�� 9�� >��;���L������ܸ��~��h��t��Ď��ׯ��֭��լ��л������[Z�3�3P3                                       �pk�����������������������������������������������������#J��!C���a��V�slm�R��c�� N���=��B�ҎO� A��!A���k�����ر��ׯ��֭��Ѽ������][�3�3P3                                       �rl�������������������������������������������������8]�� F�� G��7��scj�:W}�;���5���%���bUa�o]_�;�� H�� F���ut��y��ٲ��ر��ׯ��Ѽ������_\�3�3P3                                       �un�������������������������������������������������*e��:���)��� L�� >��
V��9���4���'��� ?�� A��U�����q��uww��y��ڵ��ٲ��ر��Ҿ������`^�3�3P3                                       �xo�������������������������������������������������]���W���Q���0���e��(���9���4���.���	g��h�����������{����e��t����ٲ��Ҿ������a_�3�3P3                                       �{p������������������������������������������̴�|v��?���V���P���J���E���?���9���4���.���(���#������������@|��vjt��s������ڵ��ҿ������ca�3�3P3                                       �}q�����������������������������������������8`�� >�� B��G���P���I���D���>���8���3���-���'���"���������s�� ?�� >��ln�������۶����������db�3�3P3                                       �s����������������������������������������� J�� U��n��R���O���I���D���B���c���_���+������������������ W�� U��(Y���Ì��ܸ����������fd�3�3P3                                       ��t�����������������������������������������F���`���Z���U���O���H���C���������������YYY�Hq� f�� s�� ��� ���������)����ɗ��ݺ����������he�3�3P3                                       ��u�����������������������������������������c���^���Y���T���N���H���B���������������YYY�Jn� l�� z�� ������
������*����ݻ��ݻ����������ig�3�3P3                                       ��w�����������������������������������������~���N���Q���S���M���H���B���������������YYY�(i��������������	�����������߿��޽����������jh�3�3P3                                       ��x��������������������������ө������ۻ����� t � z �q�G���L���G���A���������������YYY�+o�� ���������+�����w��������������߿����������lj�3�3P3                                       ��y���������������������#� �"y��r��m�Ȫb�
������(v��L���F���A���������������YYY�+o�����������*n���˜��������������������������mk�3�3P3                                       Ð{�����������������c�]� � � � �s�v�1�I��;�Y�5�P�-�J�A���L���F���A���������������YYY�+o�����������6��������������������������������ol�3�3P3                                       Œ}�����������������-�,�I�m�?�_��� z �
��:�W�4�N�'�:��J�%�y�'�w���������t�YXW�NNN��wY��͠�����B������������������������������������qm�3�3P3                                       ȕ~��������������۸�y��W���Q�z�@�b�#�4�7�S�9�W�4�N�.�F������,��$�ζ����q�c]V�LLL������������������������������������������ο������ro�3�3P3                                       ʗ�������������~�H�i�:�J�o�P�y�J�p�E�h�?�_�9�V�4�N�.�F�(�=�#�5��+��"�+�%�~�S�kqR��~a��Î��������������������������������������ο������tp�3�3P3                                       ͚����������U�T� } �  �/�F�P�x�J�p�E�h�?�_�8�U�3�L�-�C�'�;�!�2��*��!��� } � { �{�@��č��������������������������������������Ϳ������ur�3�3P3                                       Н����������2�6�*�@�<�Z�U��O�w�I�n�D�f��ږ�����o�s�$|(������������� ��{�@��ʙ��������������������������������������Ϳ������ws�3�3P3                                       Ӡ����������m��_���Z��U��O�w�I�n�c��������������UXU� ~ � � � � � � ���	����{�@��س��������������������������������������̿������yt�3�3P3                                       բ�������������^���Y��S�}�M�u�H�l����������������WWW��	���������	������|������������������������������������������̾������zv�3�3P3                                       إ����������������������X��M�u�H�l����������������WWW�%�9� �/��&�����|�<��ՙ����������������������������������������������˾������{w�3�3P3                                       ڧ������������������������L�s�G�k����������������WWW�$�8��/��&���)���r��������������������������������������������������˿������}x�3�3P3                                       ݪ����������������������?�_�L�r�F�j����������������WWW�$�7��-��$���0�"������������������������������������������������������ʾ������y�3�3P3                                       ୊������������������������K�q�D�f�������������jjj�UUU���M�}�b��)�x�w����������������������������������������������������������ʾ�������{�3�3P3                                       㰋���������������������������������������{�~oa�LLL�LLL��������������������������������������������������������������������������ɾ�������}�3�4O3                                       岌�������������������������������������ݵ����n�[WR�ddd�����������������������������������������������������������������������������������~�6�7J9                                       紎����������������������������������������������������������������������������������������������������������������������������������pp��ji�:"�?$9;'                                       귏������������������������������������������������������������������������������������������������������rl���R��� ��� �� ��z ��p ��f�}QN�?$UB)I$$                                       �������������������������������������������������������������������������������������������������������un��̙���R���D���6���-�ٌ9��SP�B%YC(&F.�                                          �������������������������������������������������������������������������������������������������������xo��֣���[���R���D�ۓI��VQ�B%YC(&F.�                                              ���������������������������������������������������������������������������������������������������������{p������g���[�ݛ[��ZT�B%YC(&F.�                                                  �������������������������������������������������������������������������������������������������������}q������t�ޡj��]U�E%YC(&F.�                                                      �ĕ������������������������������������������������������������������������������������������������������s������{��aW�D(ZJ(&F.�                                                          �Ǘ�������������������������������������������������������������������������������������������������������t��߶��bU�D(lG/+U+�                                                              �˙��ֱ��԰��Ѯ��ϭ��ͫ��˪��ȩ��Ũ��æ�����忤�㽢�ມ�޷��۵��ڳ��ױ��ծ��Ҭ��Ъ��Χ��˥��ɣ��Ơ��Ğ����u���t�                                                    �      �      �      �      �      �      �      �      �      �      �      �      �      �      �      �      �      �      �      �      �      �      �      �      �      �      �      �      �      �      �      �      �      �      �      �      �      �      �      �      �      �      �      �      �    ?  �      �    �  �   �  (                                            7 6% U   D) W, U9 N0! `?,  y (y "|% UG+ bB0 Ot8 'G_ Io :W} III WVV sUS kqR bYe Ja} fee wid ujs vwx �   �f �s  �z  �NN �SS �_^ �hY �he �rk �ut �nj �tm �ys �|q � � � � � /� � � � (�& �% �) �1 -�$ 0�"  �/ 2�6 $�6 >�: I� s�6 K�7 |�< '�; �S =�F 6�F &�x u�F W�O u�G o�s ,�C 1�K 6�Q :�W K�c C�e {�n G�k L�s R�{ ��  ه5 �9 ��1 ��Q ��M ��q ��h ��v ��t ��{ ��} ӒR �F �G ��C ��D �\ ��V ʕf Мl ��y ƕz ӥf �i �l ��b �w �x �v ��| ��t <�  F� L� T� W� (M� *k� f� k� q� x�  n� x� z� (v� @|� iq�     �� /�� v�� _�� [� X� _�� l� �� �� �� �� 
�� �� /�� �� �� '�� *�� 8�� .�� 5�� O�� J�� t�� G�� C�� Q�� I�� Z�� |�� _�� M�� T�� c�� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ͛� ۗ� Ě� М� ⚎ ᛐ ��� ͨ� ٦� δ� ݵ� ʢ� ԥ� ٳ� ୊ 㲌 � ��� 嶑 � ̴� ֺ� ɹ� ־� ��� 弢 ��� ��� �ژ �ՙ �Ч �ɮ �� �� �̑ �Ê ��� �Ȗ �ؖ �± �ħ �ȩ �Ш �Ө �˶ �ʹ �Ӹ �׷ �� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ���         )�����������_�����������_�����������k�����rzbl��l�����~���������疢���������驪��������1AD��������aTOL7�������T�--�������T�E4����������������_��������eec���������r������������������j�xZ�m������������ww���{����(       @                                     7 6% U   D) W, U9 N0! `?,  y (y "|% UG+ bB0 Ot8 'G_ Io :W} III WVV sUS kqR bYe Ja} fee wid ujs vwx �   �f �s  �z  �NN �SS �_^ �hY �he �rk �ut �nj �tm �ys �|q � � � � � /� � � � (�& �% �) �1 -�$ 0�"  �/ 2�6 $�6 >�: I� s�6 K�7 |�< '�; �S =�F 6�F &�x u�F W�O u�G o�s ,�C 1�K 6�Q :�W K�c C�e {�n G�k L�s R�{ ��  ه5 �9 ��1 ��Q ��M ��q ��h ��v ��t ��{ ��} ӒR �F �G ��C ��D �\ ��V ʕf Мl ��y ƕz ӥf �i �l ��b �w �x �v ��| ��t <�  F� L� T� W� (M� *k� f� k� q� x�  n� x� z� (v� @|� iq�     �� /�� v�� _�� [� X� _�� l� �� �� �� �� 
�� �� /�� �� �� '�� *�� 8�� .�� 5�� O�� J�� t�� G�� C�� Q�� I�� Z�� |�� _�� M�� T�� c�� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ͛� ۗ� Ě� М� ⚎ ᛐ ��� ͨ� ٦� δ� ݵ� ʢ� ԥ� ٳ� ୊ 㲌 � ��� 嶑 � ̴� ֺ� ɹ� ־� ��� 弢 ��� ��� �ژ �ՙ �Ч �ɮ �� �� �̑ �Ê ��� �Ȗ �ؖ �± �ħ �ȩ �Ш �Ө �˶ �ʹ �Ӹ �׷ �� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ���         �������¹�����������������������������������ۻ��������������������������������������������������������������������������������g�����������������jnxxZs^m�������������ww��w{���������������x��}y��s���������������������r���������|}��������}x������������������������������������|������������s�,,����|�����������,@OM����|�����������U6,OM/8F^^����������ITSQOMC74H����������,/TSQPF764,,������������US׵,,-3-�����������UQ�7644R������������QQ�=74m�������������UQ�>=4�������������������������������������������������μ�������������������dXWW]������������������pYYb�������������������hj�������������������l�����������������������������������ϰ�����  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  ?�  �  �� �(   0   `                                     7 6% U   D) W, U9 N0! `?,  y (y "|% UG+ bB0 Ot8 'G_ Io :W} III WVV sUS kqR bYe Ja} fee wid ujs vwx �   �f �s  �z  �NN �SS �_^ �hY �he �rk �ut �nj �tm �ys �|q � � � � � /� � � � (�& �% �) �1 -�$ 0�"  �/ 2�6 $�6 >�: I� s�6 K�7 |�< '�; �S =�F 6�F &�x u�F W�O u�G o�s ,�C 1�K 6�Q :�W K�c C�e {�n G�k L�s R�{ ��  ه5 �9 ��1 ��Q ��M ��q ��h ��v ��t ��{ ��} ӒR �F �G ��C ��D �\ ��V ʕf Мl ��y ƕz ӥf �i �l ��b �w �x �v ��| ��t <�  F� L� T� W� (M� *k� f� k� q� x�  n� x� z� (v� @|� iq�     �� /�� v�� _�� [� X� _�� l� �� �� �� �� 
�� �� /�� �� �� '�� *�� 8�� .�� 5�� O�� J�� t�� G�� C�� Q�� I�� Z�� |�� _�� M�� T�� c�� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ͛� ۗ� Ě� М� ⚎ ᛐ ��� ͨ� ٦� δ� ݵ� ʢ� ԥ� ٳ� ୊ 㲌 � ��� 嶑 � ̴� ֺ� ɹ� ־� ��� 弢 ��� ��� �ژ �ՙ �Ч �ɮ �� �� �̑ �Ê ��� �Ȗ �ؖ �± �ħ �ȩ �Ш �Ө �˶ �ʹ �Ӹ �׷ �� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ���     r
 ##""""""""""""""""""""""""""""""!!!%���������������������������������!%���������������������������������"%���������������������������������"%���������������������������������"%���������������������������������"%���������������������������������"%�������������������onn�����������"%�������������������ig�����������"&��������������sno�vvvc���ns������"&�������������{{ggy}wccb{{n������")������������{wwv���vww's�����#*������������|��wvy���vvy�s�����#*�����������ٟ���}����}}����ns����#+��������������������������n����%+����������{vv������������vv�����%+����������wy~�������������yy{����%_�����������������뵫}����������%_�������������������������������%_��������������������|�����������%_����������


�������|����s������%_�����5nom/-/�������|���|�������%l����I,,
@?OML�������|�����������&l����5SQ,
,OM=DGG4�\$�蟵�������&l���双UQ7OOML4477�^������������&����H@SUSQQOMLL=749H&������������)���I

LUSQQOML=774-

@������������)���<LOUTSQҳK,3334--@������������)������UTS�
,--22-J������������*���֎�UTS�,,--42-t������������*������TS�=7744J��������������*������/TS�=7741s�������������*������QTS�=7749��������������*�������TQ��[R7R���������������*������������������������������^�����������\������������������μ^���������������������������������*%��������������������������)hVVV��������������������������*�hYYYW��������������������������*�hhYc��������������������������+�hhg��������������������������+�um��������������������������+����������������������������_���������������������������_�������  ������  �      �      �      �      �      �      �      �      �      �      �      �      �      �      �      �      �      �      �      �      �      �      �      �      �      �      �      �      �      �      �      �      �      �      �      �      �      �      �    ?  �      �    �  �   �  �   �  �   �  �   �  �   �  (                                             �   �� �   � � ��  ��� ���   �  �   �� �   � � ��  ���       wwwwwp�����p�����p����p��p�p����p���p��p�0��p�3��p�����p����  ���������x���������� ��������0�������;������0��0�(       @                                      �   �� �   � � ��  ��� ���   �  �   �� �   � � ��  ���             wwwwwwwwwwww������������������������������������������������������������������� ��������� �0�������� �0�������3�;�������0���0�������;� �0�����  � �����8������x� ���������������� ��������� ���������p��������p� �������������������������������������������������������������  ����������������������x������������������������������������������  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  ?�  �  �� �(   0   `                                      �   �� �   � � ��  ��� ���   �  �   �� �   � � ��  ���                    �wwwwwwwwwwwwwwwwwp������������������p������������������p������������������p������������������p������������������p������������������p������������������p������������������p�����������������p����������0������p�������� �30�����p�������;;��0���p�������;0?� 30���p�������;3;�3;����p���������� � ���p�������0������3��p�������3�  ?�3��p���� ����������p����p�� ���� ���p����p���;����p����p���������p��� � ��0�������p���pp� ����p������ ��������p���p��p������p���� �� ��������p���������������p�������� ���������p�������p�������p����� � ���������p������������������p������������������p������������������p������������������p������������������p���������������    ������������������������������������x����������������������������������x��������������������������������x��������������������������������������������������������������      �      �      �      �      �      �      �      �      �      �      �      �      �      �      �      �      �      �      �      �      �      �      �      �      �      �      �      �      �      �      �      �      �      �      �      �      �      �      �      �    ?  �      �    �  �   �  �   �  �   �  �   �  �   �                                                                                                                                                                                                 �  000000$0(0,0D0H0L0T0X0\0d0h0l0t0|0�0�0�0�0�0�0�0�0�0�0�0�0�0�0�0�0�0�0�0�0�0�0�0�0�0�0�0 11111111 1$1(1,1014181<1@1D1H1L1P1T1X1\1`1d1t1x1|1�1�1�1�1�1�1�1�1�1�1�1�1�1�1�1�1�1�1�1�1�1�1�1�1�1 22222222 2$2(2,202D2P2T2`2d2�2�2�2�2�2�2�2�2�2�2�2�2�2�2�2�2�2�2�2�233333 3&3,32383>3D3J3P3V3\3b3h3n3t3z3�3�3�3�3�3�3�3�3�3�3�3�3�3�3�3�3�3�3�3�3�3�34
4444"4(4.444:4@4F4L4R4X4^4d4j4p4v4|4�4�4�4�4�4�4�4�4�4�4�4�4�4�4�4�4�4�4�4�4�4 555   p  �   �9�9�9�9�9�9�9::,:0:H:�:�:�:�:�:�:�:�:�:�:�:�:$;@;D;H;x;�;�;�;�;�;�;�;�;�;�;�;�;�;�;<<<$<(<,<0<4<T<\<`<h<l<p<�>�>�>�>�>�>�>�>�>�>�>�>�>???$?,?<?L?T?d?t?|?�?�?�?�?�?�?�?�?�? �  @  000$0(0,0004080<0@0D0L0P0T0X0\0`0h0l0p0t0x0�0�0�0�0�0�0,1014181<1�1�1�1�1�1�1 2222d2h2l2p2t2�2p3t3�3�3�3�3�3�3�3�3�3 44 4(40484P4X4`4h4�4�4�4�4�4�4�4�4�4�4�4�4�4�5�5�5�5�6�6�6�6�6�6�7�7�7�7�7�7�7�7�7�7�7�7888!8,818P8T8\8a8l8q8�8�8�8�8�8�8�8�8�8�8�8�8t9x9�9�9�9�9�9�9�9�9�9�9�94:8:T;h;l;�;�;�;�;�;�;�=�= �  �  �0�0�0�0�0�0�0�0�0�0111 1(181@1d1�1�1�1�12<2X2`2�2�2�2�2�2�2�2�2�2�2�2�2�2�2�23 3(3,303L3X3`3x3|3�3�3�3�3�3�3�3�3�3�3�3�3�3'4O4�4�4�455%5+5E5`5�5�5�5�5�5�5�56#6Q6y6�6�6�6�6�6�6�67!7'7;7@7Q7g7�7�7�7�78!8B8m8u8�8�8�8�8�8�8�8�8�8�8999W9|9�9�9�9�9:::9:[:m:~:�:�:�:�:�:;3;E;V;o;t;�;�;�;�;�;�;<Q<X<^<o<u<�<�<�<�<�<�<�<
=4=>=T=]=n=~=�=�=�=O>U>[>a>j>�>�>�>�>�>?W?f?w?�?�?�?�?�?�?   �  4  00,050F0U0g0u0�0�0�0�0�0�01111$1.1:1t1�1�1�12/2G2Q2v2}2�2�2�2�2�23)3_3p3�3�3�3�3�3�3444#4,454g4�4�4�4�4�455#5<5R5}5�5�5�5�5�5�5�5�56!6L6\6k6t6�6�6�6�6'7;7v7�7�78-8Q8�8�8�8�89-9K9o9�9�9�9�9!:\:p:�:�:;;/;W;a;u;�;�;�;<Z<n<�<�<�<�<=3=G=i=p={=�=�=�=�=�=�=�=>'>b>v>�>�>??5?]?g?{?�?�? �  8   00`0t0�0�0�0�0191M1o1v1�1�1�1�1�1�1�1�1
2-2h2|2�2�2!373F3^3p3�3�3�3�3�3�3�3�34'4L4�4�4�4�4�4�4�4�4�45[5i5�5�5�5�5�5�5�5�56666 6,6W6e6�6�6�6�6�6�6�67!7-7=7J7S7�7�78?8S8n8�8�8�8�89G9[9v9�9�9�9�9	:(:H:Q:b:i:�:�:�:�:�:�:�:�:6;?;c;�;�;�;<<*<�<�<�<�<�<=J=S=w=�=�=	>>$>>>�>�>�>??'?^?g?�?�?�?   �  4  0.080R0�0�0�01!1;1r1{1�1�1�112B2L2f2�2�23)353O3h3o3t3�3�3�3�3�3�3�3'4v4�45565<5F5R5X5^5d5�5�5 6`6�6�67(7{7�7�7�718Q8W8m8�8�8�8�8�8�8+9g9�9�9�9�9�9::: :K:U:`:i:n::�:�:�:�:�:;;;3;L;R;�;�;�;�;�;<D<V<g<�<�<�<�<�<�<�<7=@=G=M=^=d=�=�=�=�=�=�=�=�=>)>?>H>Y>i>v>�>�>?-?;?N?T?h?�?�?�?�?�?�?�?   �     .0>0M0R0x0                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                  