MZ�       ��  �       @                                   �   � �	�!�L�!This program cannot be run in DOS mode.
$       �m*��D��D��D��E��D��W��D��/O��D�
B��D�Rich�D�                        PE  L p;vH        �       �  � a�     �   @                      �                                       � �    0  p�                                                                                                         wjk      �                       �  �wi2      �  �  �                `  �wv      X   � p   �             @  �                                                                                                                                                                                                                                                                                                                                                                                                                                                                jO��:��K��z��z��z��z��z��~�N��}��z��z��z��z�����z��{��z��z��z��z����U���z�                                                                                                           p�  0          5�)D4PF 3  3  3  3  3  3  3  3 �   @�� �	�T/����   ���萎  ���E�,���Tx�I5� �n�Q3��e3�}z3��3�_#3��73���2�*��]�5��i��P�R�����Gw��DȎG��UʏK�G���38 �G�1��w�G�(�z)�Gy���G;���K��Ge�|�6��GGn��Yi� ���w7 .��cS-." P�a� �+��M�3����zp���� �6� S.Z��P\E\P�4X�Ѕ��P�[J�:3��5-��\d� �쉵}����#����%N0� C��,t�a�u��IJ��T��� ���g����������K&�6R�TU?3Fh�} ���1� 3E�F� Q`����o ���^�k���P��WPi�Qɍ_�X� ���
v�W��a� �����ƢM^V)6	 й�"_[_�?_W�S���c��:�^�� �#VX���a������k^j8j�	j2	 �O^�ڂ	 ��WY�5�t�jы]u�MX\j�M�6ig���H
 U�q~'y�.�
Wm: !�Ra�P�\��1a������* {d��SW[�p�Rx~ҋ��ŘtɹV5�XW��\W�� ��_�yU^���a+[�� g�O�=����:Ӄ'�y
$�6� .�Tد��zt,W��ivH._SQ& =��ּ ��'��"�T_��t�����f 5LjD���-����� ���~L�ÃV�W8��r� �:�6�<�Y��n�u�#��Tu�P�T��j�U�׉� '����9��I ������j�� ;c��3���������� �8;q��j�U��>����6\n탘De
d�yz�X拚����b�"�0�V��1<7����6�e7t�����g�b��Œ�3�	��!� ��=�T� �3q����t�1�fVK(��΁� �ڊ�� V�P�{���\V��AV�3�s�W�D��( �OYw��Z��~E�aKM�?�F��A3������ *������<
u_�k�(�zu�o� ���^��S����,+��œ��A�q stL[��t�ݓ�ޖ����[�N_u_���`�(�F�1c؆�(� �ɢEKP+�����*��E�NZ�Z �ƅ[tX� ����B������F���a� >��%��p�� Ĩ�t^6ȁ .��oM���+�J�S�yV.]� �%W@x�2�y�@g��9��$�F���څ��_��FqF���%��$�ke��vW�0���?�� �J�'� �y�Y� �E�^���^	r�	���M胬'*'��N�}qIf�9�m�M�%Y�+8�u�Uf��@�C^�Jߋw�����KE�t���:W����@��h�?�%��܋�.�z4MV��+틘)L_U�_ڔD�Fj�`�~h�w�r���"3 ��-Ʌ8 �3KmE �m!��R8���uF��P t\����D�>�����(��=����W�����Q6 {�" w�s��(S4�_wDtaV^���~�}p�u�6FN�3i����:�w1���R�_
}g�\��v��*!��g! ���DzwSNb�޻'��U2;�[_'% �rͻ"w/�" <7���K"�.e� ꄝ�F�" �f"ttԣ;k�W�>����8�AVДY4 ��@�A��_[ �QhE�V�=�'E�uu6�����`�# ����Ht�O{zd:�P�� Rb$dhS$ p��F�$ �_)��$ �|$ ;� ��  Y%Xac�tV�,��C]�Ԯv���3��d��z�oj5:9�-���&�M��;�S�^�eg)��xۥ��㫨�僅Z*�P�6S)�>�z��� �ZLM�\�5U	]�|>~�;qr���-�Ϯl�U(Ce��kኘ%�d?��z\+t�]-w����Y/]�Lj�dW�7��#s9�[��K�ѣ�oa�b�5~�D��0,.ja $�4�%���\��E��YjVP�8. ��q	����@iU{��{x-%zW�Li}S@|���i�#t]���d�^���XL'���{V���
4x��]�L��0F��x8x���#!�K�	P73�b���,:��F�)����p`k ��h;N&!Q��.H�R|���K�j���(��߫�,�f�owX"xR����e�mAXC"�#q"*  .8�[�ɗ�5P�̯��������--�i#:Oc�j_%7&�&�86E$S����A_�u��)M�?P.�q*@\�	�޹��\�7z�2o
�r����+
��L��:Õ/���z�&��(�bQ?ش��'3l�8l��(Rd4���W�O�)��p?�*�%2J�T����6d�G:���U;�0{�Qua֛(�u�#n����9�K3�!yQ(#GFX��Ki�+�f�&��z�un0�&!�o�5��?��@�� +�F=�]v�8�*>�^�#����SР�>L`#&�H���G'觻�L�� �/KCE���l����PuQ���\>���BW83�✌�D~��f��$��@���Q$\zd୷U
T]ڿ{���9R�@)��<�`MTP���h?���>Q�`��_��qqi1Q`�ѭ���+�p��(	(�)$SѶ�j��hZ�h����t�Hl�D�1����ӫ��W?,�i�#+�h7F�^C9ʮ�w��Y��EֲT*ҫ1���״��?��$�/XT��I�_y�2'���A��Ӝ�2@��D����1"�"o�֊n�J�9��o��}�=|���Um
�:V�g4���=��>qjyu'�����.�3N�p�f��I13��gINw�2*y��pb�O��|č�����@8�r�c̙S� �Ό�u��3���)��p�!�R�^������������{���Fx��
.�6�����|��w8��3h6N�y�:��5?М�r��1��e���b7��ӸK���W �J�O}����Ѹ�Q�q�@8��w�v�Q��B4��P��D��r���ѿu��E�?���;+ɒ��[=��(�-��*��mD��w���+u<����0��t��Q=bMP�)�#���G�jba��a��uVO����+JE;&��|f\&��|�z�����O��hvh7�d�W�^�wl!��+Ȑeo	����he�	�r�R��_#x��f�Z���ڀr��ä��C������)g�N/�❴ ���R����j r�R��Y���:ɔ�V��u�juh�	y{D�[��^�O0>E�����\��#UI�Si`x'�aj@�2=�:5SH��&E��ϔ;42V0������N"O-�V��*�C2�f�:V	��=���e�"Q�j�o��I���\�fi[��N��E`t/1�niJU,W}�&�V��$�[��4ˇأ�����@�����|��(�s�����4����I���-�u�R��m�e�I'i���'���n�m��]�X����S�g��_�*Z�3X�c1s�#|F]ˣ3���dP.��=�';B}2��꒓DSڈ~�8��	��;���X>����)>ȍ�6_[��n<��_�<�^�Z'u���n��W'�_KT�E��K��0c�R��X!y�*P�2)G�O_ʬ9OM�0C�;�4��`j�9��e�ǈZ��磷`�QL����9�y�p�Ih� c�sc�d����:��t�hH�h=�_�	�8e��\�D�#j�L���cF2!o�o���6BC�J��വ�zw؉�a�{���0*'d�h�F{[�_�	P�k¤.�x��N��O ���k�
���Kn�IPq�N��DFE��ߐk_M��qG��$ߞ�j���]��o_�`�o/��Ct�����M��`��_��jJ=�,w�˷�(�i�e�>���3�x5�u+ �q_'�7���2#q������D ��P�"�j��Vw��DR?A��A���c�y�a8��S�W�փz�($�Ez;�C����0����v�O��|<�|q���4��!�i�W��ku74�]};�c��"�y�X�S�)_�ܻU3��W���t�N���{�b^��/zZ�8N :�&E�T����3	X`���[��T:P��5��%��:���ܵ✵q��U�E�M���e�m�U,��7�b��0�fT,�N�suF�4}��1ǵ�w��K�V����TK�e	덡}?���kB���g1X/dE�XXF��@Q�u�'s�oԌ���Q	 \����SP�X�Wxl�Q���_t����Ա!X��ah2������i����)9�Qz�^�"l�(�tcf�
�3�� l-����c�ӟ&���#���6�a�Ka��^�3�je=b�V	b��
V^M���o�W�lo�+g0�� u��XP!��n�liM�����kNr[��J%A)��g�
�a [�X��ô�aO�\4h���U�a6�_*f�'d���S�i�p�D�%���b��A�"P����,���_�����M��_�y���!�a�fd�k�Q �{C�4F ����`rg�؞^���yN�e���H�e_F���L0�z�=rW�CգF�H���M ����x.^����E � �T���8_�72[mLb�ɑr�c��:d>��~��A�g	Z�g�� "�{:V�4�9@^1�;Sua#��TTy���d�b!h������e���ľ?��-���v>��1��ӋY�0�Zc%R�����h����|�5O� �7Yq|� �m���r�����@>nA���hdi�by#-:W��n��d�"U*c�r$ꡂT �O`�.v�o�~��6�mB����gwj��-`�L��	���!2�~υo=��gTph f�3�D���qӵuU�6�zK�5�Рr��#a:��QjV)�B����`�;$ G��s�3xW��DlKM�p�O���<�3Y#�](K���:��cJ*��b��IT.*&� �p���sue��k��O .uz
��A�g��v�p#��ځ�s���W�����q��*	j�+���������)��V����_k[�i&_D�� 5\@����18���K����g(��?k�P"�i�f������u,���.Ԛ����ut�+f�|�f�R
�s2���vF��t��!v�CT��L�ra�9�����46n:�M57������A��G�S�[lV6��e%Ic+��2���q�qw)�h����\;-���������b_D�{�3C�-Y�%bjѳ��eeD����l��0�0�$�Uh��&��(w�]�Y��E�P�^��ܣ��dA�t�_y ����L�T'E����cq� ��Ou $�#��KY�FV�{x�#�� .���p�ijw���x�K�.�tZأ:�%� ߳r@��ohhG�%"� e*��fv4ԇ9�D���YLLH��x�pD� � 'g�w���pl"ϲp�4칅"`���KU��P��q!O��R��o��Q��vq7�EwIP>�\M���ȧ5��̚�/������F� �%�$���L#64\�"�����ʐ�~��F��36tp�r^炗�� �e�u�'EF�==�X:��g�:Vo1�ns����i� �P/�ϕ��~Y!������)Ե,wL�nY���l@��F;EH/_6�s���5�������\{�jI� 9���$6�(z�t��;p�uWB��.;������K5�Y����v�6����_��GLEڮ �	�'͎�'�@0m��א#�\ՙ�vi�8{�
�'�czxR;sh�%wp�/|Ffg�ʀ� 9wG���L���W�XwY{5 a�%xh�V�ba �;](�����땙���� ߣo��B9�nU���_����	�*���WZ)ra���xX�}�HҨ�%y�/�S�iO �Ԧ>�h����Z�/w7�/& �1s]�D~�A����9��sa����z�)�9n�!�mB-�`Ac{�#d�Ѭ3Pg&-�=��P�/87j�,��𹜌B�}�4c���6�o�Q�bES�?|��L,� 朢4��a��C�\�|9��Y�I-�~ W�`q7���	1	����P% �C�ED Sؤ���s 3]t�c�ձ�=2��
�& �OƐ�nV���$��s� S�0�T��R0q����#���K�6vP�}L�W�C�S:��p �P9�e�� S����k>�e�mk�N9�Qm��H�� *�eKlxgjx��վ�y�� �x��,��"ҝ�R����^��AV{��ʢqhK��M- "H�w�Ѣh�M�hVg���u��/�ll�:3U�ƨq�7w1d Vo�EK?���������_8����MPؗPv�N �:�\jꊯ�:�gO#�K �E�K���cw�t�Ϣ�j���G��N�����*fa&�� (GEb�f\���'��螼�T�
�o����UᄄKJӕK�V ��jpR1c*����9T�e,f6\?yGǘ{�������ͱ�a�n�(-		#O�U�z2��ttu!�
�(ES�F�|X��&+��Q&v�z���0h�3� ��e! �[�����`�yq��g���|8���>d�	#��ύ���@L�&�������g�� �K�f�g��]P/1ͺw�l�cG��� �Q	�C瘻�M�BBU�3�׉�~J���z�$�@/�yw��z�F$���
����ݟ�5�� ���)�ܶ��(�My*��]2ht�T�:��id�`it�%�d�g��i��z�婋�y��$m��y�)����8��j������dM !������F�@��_y>8�窷�?���+��+ � &x�C�y"�~�$�T�����֙R��+��j��E �gC��֢X��\��#_ڪ�� �j���AEP�C��Ί#a>�5�19�	oA�nn�2R�$��I���Ɏ��4�UiՆ �A�V�o����k�Y"���E`Q�j��'�aL��x���Nα7f�N����1�?Z��P2�E���!�������t�^t���@r�d����;�Dyu�I3�������Ģ� �}RY.�sp�h�%����p�FFL���.R;�� X;~��B3�$��։����|yeq����5\������_e���������$�~w ��� f��Rḍ�q�ѓ�Y!��Cя���w�#!Ͳ��5�r��$L^㺾<~A?dh;;I���:s�[g' �3������D�⭏7g+�w������1t1`dQ͝�M/�)����kI��e<�XYq*�u>&�sRh �!�.�n����\1N��N�C�[�hg�O2��v�dd�9�����l/C��Q]_�=��5T�9ܰ�i rn̗R�Ze_�~x �}ZX�_�^���<��.;�v��j��g��/B]�H+(���`Cd���E��c��SY�z�� Q.6�:d�幌 T�y��U^��\�UħE���ř�uF� �e�I2	�`t��b��@��12�5�њH�)�EU �ė4�E��{�#�,^��Q�O:K$V����lX�2�?Lt��	*��m&�e��� �Ío�h���e�\\����E���t��Un���,����ʤl���Z������>���] E��� �zstj}�~��KJcIu)��`uy^ �K!���2FIc#��l�ΌTn^���)�]ݼ�X�4k��� �L__�)���$��
���C�|�T�����Pxf=اu'i��}�t�pwD�#~X�8	�	0٠� ܫ� 8�����/����篅�[�Q#J�/ٔ6�PB�a��i[d��8�!g~��_w�E?!H
��uYe����Fn�S����@�0x�z�K2���!#�8ʿ������W�z �ÕM�������Ȉ��m����Be�ز�	�`{n-�N �p���~2�t 28��s�?�}���k�f��o;s���J*��d D5�?�I$t=���h�q&��	���'����qo��LM!x?꼶�d�·- I�օN�x�����F��B#�/�jj�S"4��&�o���z�%�- kb�Q}�O	���	0����,�Q��{���k���2�ֆ-?m��`�o�� �:���HP�o ���5�X��F�"L�8[�.�s&�u�9��t���"9A |_n}�B���8 J�9 �� $�EN�S=	( �t�jS_�����{��95��0�_��Da�j�x��i1�pl�V=����s�x��o�P ��w�Q�0:/
�|�<��8��Ⱈ@`�8�3��ʰu���S<��ث��Y�Mt!�l�Njɱ�p�xZ�̺���y}G���q���i��$�)��f�6� Pp�_�c$����@�a\�:�v�,�_��w�w�1ݚpJ��٢b� kr.�h��Z��MD�(&01���m�W����� �A΃��_�/�u���Z@Ԓg������Yzs�ت��t37�� �����R��]{_����Xŷ-k��ޤ��e�
�RR� �y|v̵芘H0��G�.��=an�q[�G����@q�1�_3�p6�R�?��5 �W��ιq��߫?�δ�e]�.�TF:��)E�������R/d �4�t�#Q=jZ�䔗p&Iz:���ݱ[Y�Ŗq;�#Z��SP�8�r�j��B���P 1���3��������Gv[C&��^ s����=��O}�H�#��j�[��=��44\x�L�]K���oyD���6�>ѓ�L���N��4w\,da�d��b�g���MK ��~yvg;��s��D�1m ��O���g���s�2{��\� �����F�H�d��M���bnk(Q�v��B�����Gb��ؓf�#*�ׄ�"����@?��I���]k�������� �� ����������A����x�l&j�"Ũ��@R�ȝ�l;>~�������2���F��O{X]�׋H��uA�C��X�E)әX\vI��� ;��Q�}*[q�泔)NvFxB���|,o��������ؒ��\����0
hE0-+ =��1ڨ��>!z�V���3�ؐՄ��D��33�ᕍ� �1q�6�|S ���N���>Fר�_ʑ�s!4�`�����0 ��Ҕ�܆����d��^ k}��tq�����2jL7���KDP�%>���ӊ�M8�}�2�� '4�� Z�U(�e���}�^dp�]��JUj��m�O�����  Q�[��l��K���HE�z�5��<ZBL��V�`�	��=�F�CWt�O Y�޹V_�l�qq��cT{���H� �6	���Ex:�Tq�k ��Ӄ�1�v��t������/�=��>�S缛��F�I}bTV�z��6�a�^�=������ĩwݦc�!A�bq+�U���w���~YG�s�ZK����o��b���4�m���I'����N��� A��%����VI�<\�ɻ��Q�T�'0��Z�sl�$yŸ �A�5L�;����q8��[�ۘߥ���Ĥ������� �Y�s܂�g-��B4�0��4���A�fP�"9�ΪwC:�؈�/��M���mz��f��b�~����H#i������� �c�A�e�|f ��u���y��������7�}��e0��aD gWPt��&"I��@�:
�C����x �5��̮.���>�i#��Ns��0\��W��W=n������hAaD*�v��ex?j����2� o��Śʩ�*��^-j������	��?MUe3�$��<�}Ј7"��5�0����#�t�����5�����۱88�ӧ �������E�QB���D���9ࠤA �未
�-���z�����?ү�$3�.�f�ޟt��Q�\� �B�{�&u\��]�߱���=�;�����'/V�:d	���z��y��7�(G� �>��SEGp�J�5�>���[�|��y>��0n��H��w�:����N�B�߄�gsZ ԯ)�ۧ�7m>`n;c����q��SpL�3j�`���<��7��]�ΩI���3��W`���@�?�%*���,��L��Ɉ�5�+F���0���_�N�������A��N	��A�z�I�����T9���8
�a�-Dö�!$��� 3Tj�Ň�+|%r�1�Q%���3���@y��U�'Z,Y�
���kt=���a�S �9¸�hl_a�v%+��sP��' �uu8��;�"zӍ{����fVݮSo�R��X�cٟ*�ↆ ����ۿ�Q�Z��W��ÆW0�_�}~�W�qn�u�A����x��K�_]ߍ�� ��ښ�3�$�.W_7��ƙ_v�=�б#���bL�����LcK]�ې�Kj��q�K��h���ZO�ǀ�G ��_��]"��;Ϧ�S�u�W�5��*��hU�hv�^��s�~����@9,p�[K
%����F�d�^iOZ� �C9��+ ��Ǎ>�^��eP �׸���4��
��1���&@b81�h�J��X]�C���GL�<���Y�~��D��Ռ�9���Ò�u�� H�MM�j�a��|T�c����r �w��c��^Vs�؁Nl׋jZR>L�t�<����#
���ہ�@L�(���uEiK�G�݅3����~Ne($_l�V�x�6r'��Φ��B)��}t�,�ǡ�c�SK��L�i��eKD�|���X5KA݂27�W�i$�mp*-u��&αYlvZ�b�����;�A�+� ��S5��jw��f	�  t\�S������t�����c�'#�h|C^����0��8:QӜ3r ����rНҥ���$���:n�G`p\��#���Q�=VEbN�n��l8�`X��@�lvOu�鷟���� k T�N�"ޓ/=����
��kT���)�H^�X%���M��C��^HS�����U~�=L7X�6?^ڒEn�:�cdTL\/��4��}A�c-KH~�u�3	{� ù~]�mI<k4��H���suZ�H�]��V�V�5#�h}�;o��ȷ/fG~��oz㊹�Tu�W;�$@���\�zRi�oz�B�7¢䐚�|�[6���U#�������U�f1�x��p�w����-��q�LL '5��WE���{��Q�!0��i� {���&����v����BvQ�A`o�_jX	!0z�-%�M�y
7�0M�-���TF�8�n��c� 9u��8 P��G'/S l��~�_3 y��WD
=Z$(�5焦�� ���?~����u���wü���U��� �Kxg�(V�চ𷗞p9Kquy�>\?�2)%��/{u��y��m6��F��M��ru��x�%$�T��� �`�#.�Oj��z!�ܲ���P����^����4�Ա�7�2x�8�m}�^�! יZ�k���585�ۀk����0�h{�~����%@[��b����C��E��;l@��tЄ>�ͫ�����e���@����]�?��u���]��
x��e��>�]�b�5�H�m�OL�5&��VY�7�@=��D���:�Zq
8�-��l�Ȃn����~I+�Z`:1[o���%[a�g��Wo��/�I9��N����Y���8��il�0և���� <�+𨜼E��Z�N��x�Cx7�2g9|)]h5��K�տhӸ����)����lF��;띍-�(:܋���q���5O&g7-$۩`�n�g�yx}mx�� ����|���I�����?+����R��N��j�j�*%��.��Ź@W
;�1��� 4�І�0���� ��>0�
��C�B���L@y��� �>
	��NqG��#+���ǜ�?Ⱦ'����}��#��w�Ytϼ�B�>s?���L6�$�ߗ����̤�Ȱt�.����Ih/ �6|+���]%��J5��<��v=Ǆ���ί"[?�;{P�@��!�A�����T���=��b,���N�����<}&�@t'�mvX��Z2�'������Nзғ(o�9h�4�	�4���1)��`p�Q���V�\�tsq,�":�������3�LTX"(��*pq4>����(�o4z�2�a !�P�]K�a�]z�do�t����,Z0{R�aݗ7.�
���sذ�DZ�H�Q"h�
un��ƕ�zk����܁I2�'tPd��z�!E�4����R+�i�O�kX~�>ƿ	�z��t2�g�ڏJU��y����@5���#n4�T��@�r���`�����P*�j#���#�p�H�v"��-�h�#�X�Z��l��.��D!)B�$Ten�zc+D�L��ڃ�_R����S�鴤t<���hH�w%"-���+M~e��۪5�n�\qrc�$S>d�� K{�%V��jBE��d����t*�\�>�I��;ȃ+�M$q����OVD����>b�a%����`��!6 t1F�tr�I�t�#�T�uG�fG�I����f;7��z�(%�(�5��c������<��X[����z��0��+#9��g�j=mz��;��8>�]�����G�_�[&(E���f1��I�3(��7��?�,��^=�p����Xg<��S[�����Mьz��6z�C����Z�����3��Q!R�9 |��J�N���
1��W�8ƴv�  ���˃(�
%�b���]}��T�'�=�o���^�1��p�Q��D0!��]q	��t��� y^�q��}o΋w`���o��$�t�y��N��HeKW���d��C�_��� {x��O��o&+���^:�}�d_m�u��lj�`pb	I��)S��$����|�����'��_5�D��)qq��|*�fW	*�U�M>(��z8}���uj`)�ީ�Jog߀Z�t)��@�A��ŁҴ��ʯ��+
�4�'�U�
�T+��G��������p���AyVo�L�~�響�l�<�l�����10�tlٴd��c��OS��ߤ����(�v�/�=�d@+�2�¾0�f�p |Yy2!+#/�@�T���O����{3�e�v��f���� >0�N�!6
J�	����Ē�&�Ru�T�Cz��K2뾦��xx���џU���g�;q���_򹇾:0�������?II�h���5�{�k����L��� Y
;uJ�_������b���h��Ȱxm��9NP�e%������;>2��7R�d+H}O���J�xJ�G��16Lt�Z�tk�,9���=L�����noEڍ�5�J�E.�@z_Q�u���s��Qﵥ@����)0�re�`ob7䁹����%s�Z�L��ÙT|5Jc��v2�ov7�=�kN	�\�P��O��-��� ; ��/rQf��X����}������W1�Ir���l�,k�/�Ɓ���U��
�Ri��b����6?���jlW�=g#��+�1߷��N��N�9�h��,�T��Wlh�&��5�w�����~"��'�z�˫�"�gԎ��%�����.���:1Ϣ��kM�Iy�i��)��{1a�c�QTS �2ҫD2�Ǵ���r؁d;�����f�X�,���,Jq�9V���(���'��mo�=;?�v@��R�o^��y��{n��S��)��zي�{���9�&a�/Bd��S��U/y�p�%����=�k"8��ؼ8zٸ��E2�eH��) :�G�;`R�(�~k5dK�>?��ۗ&A�%
�Go�F�항2�|�'(�W��.�n��V4�V�^&5F�\���(�()r7V����� ��]�ۉ��]ok��[��	�­�jЍQ�B&��f,ɖm��f���l����~�wM��I����8BW���V�� �a�'�L�x��,�|폥�������K�h�*b��=Pe�5A�W�@�g����z���	�}�V�8�����؄魶�Dw�+�߿0I|G�Y����5��Ī���p��U r90�w��1��K����/�5}3�`e�e���7��T�f��4O w2=j/#baG��'�1�SGɘ������~1}L��t��0��c-pa�#����A��ᗇ)q��\��]:Y���J��M����?g���sG�(�e�?���Y$\7�y��w�>�~����A#�@0)���	,�̀���(��$-'���dl�n����d�AL�Z`Xf�A-�������VYe,�aH��P��Yy�����o�=�2���;O�(WvsXckS�fy��}��b������O}��o+��ylҽ|c��P9@Ɋ��Ck�a�2d�+�GܟA\΍7�#�vHP�o���Mr�K���Lz6��oⷂ�ad�q���W,��xUu��,�
�������=g-��P��A�])1nK�#�Τ�+8b
���=Ǟ���Ҥ�2�
(�j�V��s6G�~u
&��lj�L�jX��x*3L��t��H��Co~�J
Lh�֖�?�L{�'ژF�$3Ќ4e�"����|bA�-��U ��b�����%���ٌA1(���H,�s��7�K�hl��Kv���7�	4��{������8��6-���#�z���e�}�-�n���*�n'����f&'�fK��&�P;�+��H�j�x.b�j����-#�)J�^�rE$TFi��q ���<}�j�2�H�/�V�"ϕ�{�
�"��z���� �+��;9���?�L�d��Rܔ�jD`	?�[MYt�;c����I�3��X-}�U[�a\+�¬9J[�O���D��l�Yn�rIo^��d@�g[��-얓4��W�r��!�2�cs�[g��X����$���٪Y������Ҫ��>j$;^3��>�����i�8���y�"�7�<a��a��Iq6�o%LT��9��]��Sd;zސ�R {�t*t*dԹ41X�+��
%}��*���~5��5#7E��u�/�_�����)Ig�S6��Ġ#�>mí2���U���WJ��H|�qS���n��6"]�� �O �# +Q�6׸�'�'q��D)7��a�6�X��cJ
w�\�r��=��蛑b ���vC�vΗ%m�/��w��sz��͕z���=n�;�ĺ�$ꆔ6�of��sK��A��&7�#�, �q���X���)[լr�x��1E�������L9N�@yF��8.b�2�}���oGm+th�MB9�_s'�(qR�|-}3�9�:��Ӑ�0�r~[�0B���Zk(��J&;>�;��GWr^�1hf��n{O	��g��2�J`�v�-�U�_T\F�^�'�a�F~�
X���#�ʫ��J�� �'U�iQ�e��9b��g��<�iƑj��f9��=ԕ�s��L ����CƮ����T��ڜ��1��y{��M1�٘-l%�sD?���O!��*���H��VzK5�H����U-�@�?�e3���n  䧉!Y��z��_�:��"��;��1���3��t��2���S���?.�4EYZ���(FE�E���:�/?O�&��q�ܛ@��7�xmY&��AE+ܴ�y���BFh��
�t�g�<�>�U�X�	b1&�]�v�P��<!�\T�o�7pa�)XN����L�t�������sZJ�\�%v��x��@4���o�r7.��GR9��5t���23�\0��\��էD�A�(�����o�vJH�N��k�������(������Ξ�̓�E�]��"�����A�P���<l��I�~� =*�ȫ��uEAQ�f8|0J��A눇�U�\�9jM� t���d�`�?ǂJ<v.|��-�-5� x����;ˢG��3n7���*�ToB?��i�
f��98�Gpq6�"��L������x��f�����]`(�Rk�=�;F�Dq��}�uaC�:ЩWcH�먪���GQii��}�J�����
�|. �����X���F)� �9$X��N!�?@�ˀCk 4恊U�"]C4�����*�e�;!lMf��ʔaγ0I.�g�y��jB�U�>�7v�'+���{6K���w��4�����OE�*�l��<'�=h�A��~�8}��ɥ<�e����x>+���>�}Z���?O&�WS�\��I6�I�L�~����dq��b%��:�p17;o��Maq�s�K���~�)�wt$oNb��߾�7�T��c6QI�N�0�|Y\���-y�$O��:B׍G��}h�q�%�SrA�6ո��Ʀ:�/��&�FR[̒��?�u} lcZP=�����v@�r�eh�b�;��S�G�S�SM���c��kO0��`!'J�Qh��x�}_�@o����L1�YQ���`��+�V�Vg�!B��9���y1�9�oB�T���&��RA_���I~ᆂ�y���zW����O>bV��S)#���z���u�����h>��������S��>�р�֏Z�PHD�F.�f�h�����=��u�T��wc�{N�|�O��D�\*�71�l�́� fX��m&� k���k��P���t��7֛"��zUٰ����C�����w�BZ:��X�ZF�@f��u�q��]�<Vx��7o�P�>�O����\�\9(��u�+D�sLU���H퇉��rp \�q7�Ǎ-���*�?T
%2��E[&W�Ø��H�-ľ��D�Y�=��<X�t4�-��u�-�$�I�.��P�?F�r���P���Y�E|��1{@i!_���Qg�X�^iH=kBk|mb<-��e�v/Z'e7�q�M��}������)��7,�^t@�x���I �_+��^�:6U;�����m(�}"�M[[�/i�d�B��?���[��!?o3�M���0l����7��O�-r%F+��՝������/�D0�%��	�Xr�]���*�����I)|���p��]<�1a�eE�y�<�V��}��� 65"a9�J�]���^��C��@�sw�%�%��������*�US��'�\��S�M�-�n�� �H�*�����PٟXZ+9��ڂo�� Τ�̜�#��i[s�OVDU�F>`�IR)����ǥ܋���G���x�?Yv��eB|TH�o��OM�N��,(�(Șn
��3d=a�E7.�@jq�Q妣�DϠ�n�SgQC^�ܧ�e�C���ql�hZ*܇l��_c��
>ڵ�� g�f�6���(�0Al'����J�p��A�v_�y����G/'��x�c�d�)�WT3�aE��(�oZ����M���[�:�sad��4�~H_���ɏ��
Sx�� �_Z�2�]l�Q2i�V'k�~NA���)�mX����Ff���F츭���e� ȫ��V�r��^y%�W��̖�j"�˺��	�b��E��2)JRp:��{UQ�?��g������oK8#f��a��T����X��|(�
h��m���TQd���|�� v]>�D��I�=hN{B��a�u,��Q��a����D�����uS��� |mI�=��t����	ic�Ď���%�?ʽ�}n�w���ϮGe��n'G=�VT�.x��K��H���@��2P���ն�O�8�x-5�r�Z���At�j��b@��.�������4ҳkGݦͣz� ��(������/�F��8�,?���{8*��I��C���P~�7�r��Lr7ܿ���8��h���Z��XտO}�@m�V��sl�S(�F [wV��\�2��J��U:��#�&�8莰� �?�NTj�|�n���lp��P�Ʒ������/q�Z�h�q�1{�<c����}�e�=@��>_@���%�ۏ�]�id<�YA�&
H�ު�%X��7�|�+��SƢY9NL|pI��/�D��Y�����n�%��s�J�p��E-BQ�r�W�<\hDv"��������GrX�ق�Һ��,�ff#"�g����a	n������1%|�\ɐA}�pjC"�P1>e�N��X��K��&Q�������ps�8C���Rc{�LR߸"g͆��_]��LGm��*����s�'�o$��93tfg�D�;l��Te6�["tv�n�#EDUF���ё=~���ϕ$�/���S <e�����D���Ǚ&K��ىd��r��� ���yqq�>hv��9��o�{��K�v4�H�D��{T�c���Y��D���>�QwL�uҚ(�y��n���A(�%�g����%�#JSR�K����g��<���;xk��'��+ ���&�W%����ם�G�Z4��<�4�z��&�ܻ��t�J'�02A�,�<���X�AD�������B0���(&�M Ԣ������y/OB��Z؊:�f��F�u����O�
�;K!�Ԭ��
/���Q�8^q�ћ]��3��K�
���sJ?�"eF��>�|�޶{��ŭj����j���cl�=��b���)�%�\Q�W���8}��z�г���	���<��F�5�Q�"�3��4���j�17z���(���˻EY�Ӛd��i�^k��u�+�:|pp��~g(���I�B��XVs�kr�:��?yU�oA(5�����>y�D���/�J��jO������SY_y5o�PG�)Q�a,L�v@+WƩ�|�K؃ ]���M�}`�^��P�j6Dh�O�K�A�o��l� �!;4� �nǕ�t0�zX݉ )�`K���ͨ\o��T����]��L1r������M��ŅF�":�1l��S=3����=�\��ʾ{��A��r��/�TE0��0�X	�[R�^��<�
���Z:t�a����4��s�bK0�����T�SEm.���OQ#�[~WY�}��8�˝op]ai�H�=���L�o�� ��0K Ӗ���kA�mՐz��Fo1���,'�u�O�	t߉����R.�n� v?�\�˱%��]^�8���!��;�o�n�W��L�`��0��)@�ێ���3D)�ʣP���C� ��x0��-��3yZΈ�_�p�C����`��)��z�]��mr�����%5�Ae��'���1��Տ����T�}:f�[77�-�s�L�3���e([�1F�Q�E�͗'0����Cq@�i�lΡI�����#g�<J>��=qF�c�['���+*`��&�? �WK˖����%���#�?�}�	��3<��Y���¦񧍈��&�2~�À�AȬ��%L�ī����������3#�|4��`�yǗݱ�P��4����?�IV��=�%�B7��Y��5Xqm�[��l�WL�^�fXT��������z�/e%�;�R���(��;����0����n�DS��A\a��RS�/�n�!I����ۥ*�Λ����P�`��C�i�V_�g�!m+6,PJe5�v��œ��B[W>�1h�܊�U�t�]��;/��K�F�ɱ�pf?w{G�*�d��"^��ꖯ��;�9�����=��y��%H�td��?jly�#�֥qڛg�������9�E�6�Y'�e�`v/��n�(/#�V�S�|3�=����ė�s�H��n�Wh��n�p^�-��E0���ٲ��nSU��t���`��+�<�O���&邸����A�]����;�����
�a�~������S�o-H"�+%�&�Wg1?X���d=� {+���COD�R�J�Hac�������m�h���p��2ߢ���F�ԗȠx��2��T��/t9�34�7\�BQ�D���3�09�������Ƨ<A;s�ї��M�ȩ���[��BG�ԯ��=��,�4^-l�р>����6�Xޯ��+���-m� �X����E�|NO[0��dݙq����I�B�ZNR٥a���v��N8�^�T<�-X��=fnś��cÛ<,�L�]��s�NW�>[�,g�a��o����v�f�]+�D��[:M)�gO-��������;]u�Q�H>��t'�4?�4\�ݵ/����0J�~�� F��k�t.�P5��֠_��ǖ���b��)�A�r��˝���$�#� a4"E������O?�2�3cc��5g"�`5������ an�����˾F^��zY��2�b48I!��󿚢1)��SZJu�l��+1Y����B��/օZ홮[i#�<P?��2��f�1h��������9р�6����O��!c�	�WXC���#1���^�7E�Hbs膦V��3�q�׹~�@���bi$��)�_������4��բ���A]�D\F�/�9d�ծ���I���x�%�Vn��8���J�a)�\��[ѡ�=^o��x2�-�q�``z䚦"]����, C+J4�/X3q�>����W�C�D��	�`+�"O-�ᰵ���[8��%!���
al����N�st_A���3�e����^�����(���JK�B<Y����*J��^��A6+����EN�_E4A�?'��E�t/������I�]�tƳ��.�����E&��7ݵ�i{�7���I��{gAk������$�E��!��ي�C�I���6�m�擢	P:�#:�ش/�#��U�+���	���a £D�����V���E�!3)���At�/A�����{I��i��F��ѡl��U��z��T��;���.����.��{R4t�d|_]Ze��f�q�4����Aߛ?M��Q��5�JI��-�,:_�98��6����M��¬]2��<��w��0A����Z�%2k��+f���1�	����o�[qſ�AK����ѵ�=ZA)^l�6���M#�]�$��#�� ��1����T�D�]9_�i�H1��*lV�'Q<ESP%�#��;c�`�A?� �꿮R1��%�_7��r��bR8�f�㍭ް^�:m.7j��I<-2#�M�戝��>m����ƪF���D�sd`t��51�}���m�Y9ߪ׃�1�o$p!��B*��p1L~���Cr\r�Ny�H)�R,�-AaN�5[���{8}wm�݃WS�p_��:�W`Z��Ɲ9.��d$��3��U2��pQ���1{W?�s$���4*9�4q�UT��r'5z���*m��n.�1�,�&�E����@����S`��=���.�M�lz�i��Z��[��b�YZ,�+��D2�/�~��*@�;D���;�_T�4]��fI��<�+A���H8����~`T�p�����}Ox���y4�s��(�9��f��铚�D�77-����-�|�om�pa��L��YȝF�ڷ�)���Jya�f��8��njL�y[i�в��Ψ�?�OX�F8J�蝤e��Ě˚	ټ��6fdÄ@xϷ�a�HX�u��87��u�̭Y8�![�6�n{�7�&L���ƒ��Ӧ�&��ua�߻�Y.!����0�D8�N'��^���ToR�$̉�]�k�1�c�S�5�??����U?�?.�|�
1��g�>EO?x<66�Б��CY��������m��A�x�]/�٥ �t�-����pw��}�ˀ"�O3Il�����-q�3"�4΁�~��rfɲ3�=��:���'�#^����~=�������|������"4~�Af�\�5���D���X�n�a���(h�����k`�47�**c ��}^q�0�vJ���;�2�h�Յ�%6̣sHl��9?x^���D���t�Z�\�G�s����D[G��8�`�d�R,HΟ�o�XW��$j��JOr��-�ҳ�����1�ap�Z=�}���y�)�QDܕ��H
��G�곁`�q�hv��<��b��v�H����ھD���B5�:�{����K�ޒ�W(AéfGB��#iܥ~ �D+R��@	CT��:I���r�:l��?T������'m�^J�@����������b	뎧5�ɸ�y�^~�weB���M�o��4_����1�_�GW^�	ʊ:���>��B%D�ͬ�!%L���ea��S� ��Q�!�e��% :�G쯚�| �C'�����ad�;Σ-|�1�L\��3=�P��Vh�o�Lk\�*��'�����w=�mM�-��x�]��?�k�(ܗ���$����������%�ow�:��}�I���+o�۸�^�S��j�;�PgH�1�@n���]�h��Y4���I����FK:?M�]��z���0Ҷ$��:S8�f�߈=C��ԙ�)T�g]���2=)��Z����C���X�4?
7�䣣�2oS@ު=��-���v�BO� 8u����Ό��C�:��"�� �!���/�
}��lL-�������r]��!� >���V��1�8 �I��Xݩ��"���l$�l2�KP����G�O:!<t�^->���F�1aQc"����7ƅ�2�#�L�`�eB�E���q�	�/�7����������nΒ�oګ-�ZU�4�-��>p�%o�{�����&^,�-w�#_�K�@�S��F��$�W�MJsZ<1߀��?IA��ňlj�x)��\�Nn�0#�##��O�dno+��#�h~Q>ئ,aA�aVJQvPx����mh�[ɖ�Xu�,��EO]:\a�����F!��vHK�7��Q�����x2h�h�{�t`�x�z>,���C�M�Ex���1;=��*�A=��5�A��{�"���8�q�7?����'BAz�$Ȑ�0��Ϋ�Q����s����T���0��4�ze{A�!կ�aJx9���Օ�5���^)�S<��x�$�&G���uL`�}� �w�r4�GN�#Us�+���	Z�Wa��TS��)�-�T}�{"��,��Q���e��,�P�}����B}d����ܥ�	�I�
�}�Y��V #-�����;H�"4�`j"���tk�n<�����XQ�M2D�����?$�M���y�� �{�o�\����cP�}��?� �tu�[&E�YB�.z�C,|j,��M�]���4A��2EK�2�4�O#9��³�+;�%?G� 1�����ͅ*� ��"د��1��).;��CJ53:"�S��f��N@�Ǔ�x���7��}#`'��N�`$��݂9*��>���aG�	�JȃK3N%!���1 ���[f�'>(�1! �w�m���j$�
���t$�-���>%˵	݁��'H#g����~��B<�ێ���6i��NI��>�/�P��	�t��e�����S�%�<�x��" Gi�����W�$����*� �{�cc�%@6�
�z�j�_%=27�� I�M8ڀ}K��?n�np{�q�h~3�G���@G��'�<�*�ɘsfhW�ס6��=n�����2��20�Xh��L&�s4��������B��[ku\�|y0Aa*�������,�Q?�s��x[�9 e��a/&^�8]b�t^O�,j�c����!��5��=ج�����}���.�
�-��� �݊Yx�e��l�f+S=�.t�u��_���������d�����j��s�g;ehii���_�Ey��)�IS��)f�-�?�*��u�p�MTf��3��Xj[��h-@������u�`�ƾc��)����&9�15T6ie:~��V�۲�wB���,�����,��Պ۩%D������J��aj� ]M�J���n�%��S���F�"L�[s�-�	n��^/���
�zJ$0��?�<��E�;�iw�o�~���"�����P���8~��WS,�F����N�,>u{y�G�� pDS�I�4>��Z4�ƥP[ʫ���
�\�5�m�:�\�V(NĎ��s�b)�P�ţ�-Ǣ���8��Ӡ�
s]�ۚz1������H�j��·TT$���:���\,�w�Xw��I�^j��9�i�T�tJ;����\�>݃K\u���J|���-�W^t%�Ye�7|B�L��lsn��rb�Ǌ>s��LW���#��n��R_���T��2��8��˸��֗�F&��y�ga�n�j��|�+�����,v���t%CA�J_�^*��[��a�	ލ,he�A��Ǧ�vY-�@�p.�����������4������ w��j�/.{�O3��$�&�k��`ڂ!����6=��Qk�� ��ES����m�,�&$�-C�B�jV$�
��;n������*e�� ����hХ��0�
c#؟�]�oY[����Ч�M@$�Zs�$[|�iܕ*GV�/*QB;h�-�5�"k��A���}��/��+��GΡZ���I��nZ"U�soH"��D�	�c�?7޿��Us�Qߥ�� h5��{^'���� 3���}J����$����_C���/hf��Z�����;V��k�|5r��a�*�U�����Fɤ�4\s�1��2׭�*՘�@�ǝb>d'�M ��
�pv�0��߃�wH[��1G�?��?������db�4�88�!3�9dƣ\��8�9a�H�*��lZ���M�W���D��q�$��\t6(�0ʊ�V�H�B��m��Wʿ8C�����j�iq�Sf�������@�Lr,F�-�0�M�6�s��(�j¹����7���#�������Cȓ��W�$O6�/���$��Qb�+��אָ�^�+�_�=U��vЦ�Uބqj|��Ʌ[���-c"L��N���F`��P^d�G̷"d |mܵ�<K�w�A}Ӥp{&%E���%+[D��cѤw`�)���r���
��.�h����hH��������\rl�=C�W�˥r2'�qN�>�ҹv�n�'E�N�<�*?� ��^�~�B�ǻt�KZĉ���~(���2����@�q�_�e��)��;��V��a��XE�#�����>�ʡ�/��oj�|�;�35i,A��0zn��(K=�0�k����ƥ���v��X��C:�$dn23�[�Y;��U%+޴�zsm;E?�D@��5�l�{>����ܥ�##-��R�oJ[�� �S�s�6:;W3�K�"D�+����a����T�~6���ZlE�4o�<"����ժ�����z42,�y�f9�¸���ׯ!���bէ��=�2|���e6�v�8��1�<@	׆ԅ?�)��8��Ȩ"P����͚J�%����V���U$U�/��[�ˀ+�ф�h�����.�"��ˆ)\R��L����(%@<�7����7��'�N��7�<��/��J#4�%u4�z��5�哊5y#�ܖ��9�¦���J�mrY-}3�گ�~�y�O|�#�W굢j�--T@��(�:��B~��n�]��`���V�4R��~m���zZ��_�!�h��ځ<	�����Wy��;ϧܖOiT�w�Ӣ��#����`��E�5F/	��M\��/@$� �'��lK⽥s�3 ���-w�z�v��c>;C�S��^-�t14���v�DaY��/2)���E��5ͽ	��t �	��Ȕ�+
m/&��tH<��L?�j:n���u�� �a����v��?��(}����9h.�Њ�D��w����ҙ�^�]Z����K(�ota�� by���lTF��i��^�~�SHP�ef�98e��+�^'�#s� �<!�i�]�p�e*mRm��S1E6�0-.pG��i)C(�;Ҡf1t����o���-��1��AkRʹ�(Gu;j�#' �n�ҚlN k��%t�r��[ � �:����f|�?�H$9�	=�M��px2#q��2�����0<}��d���+��[�07k�"N]2�PKW���xeax�F=���Yfa�D��$p�{m/Us�B�Ҷ۪H�(��v����'#���0������r�&,�8}dV�=E�?���](���� �s(:����Z�(���������+kH!7���D���[C�ei~M(A�$@�L��S���.C�Ob
�Z������b�p��"���k/˰����Ih!�|�+��!���At[C��($yA*�.<�]}�L�͑AG�RѪ��Z�B$�N�Њ+܃>7���բP��?�+���RH����]�^�mA�sN�B�������\ho�LID���L�����"��S�Aq�D9a��Zw��O����J�j� 4PV �E��=hV��K�����ױ���η�D��DO�G?"a����E�)$�8��ؗ���C�G ��;���lw��M4­�$:����E*�e>��"�}<ʈ���o�^Lb��:��'P��1])�';z^�QV�ԩ�2��}#;'�N��"�r����c��y�޺@���Q��j���E_Uvq�<{|��]�)fw���#�)�	�Ӎ;��)�>��"�������ZBHg}��],v��*C�g���y�\(����s��,v�AQg��"c����hyk����,P���͖�̞eu�U��|s-��0������K���/���ԛ���#Q|J�5��y�N�+l�#4��%D�z��".�AF�#�e�$%a��Ȍ���<9��T�M�2R@�Lx��R���1w���L:��sy���Ģ�;7T���l`@
k~���6(U�����&eZG���kk�|�~{��Toq%�=ud2"�g|�}��MT9i��}!���a&PZ�q�����fX��1�����a=4���W.ع�a���:XY��ϼC��q`���ުblhQ%ԗ̊�-��_�6,�'� �����\��3>n���C���ql�1��Ul���ێ��V�Z1/��=2Ϋo[���f�E�; �c
q<��ړ"�e���Pf�$�?��r�^O1�G�?�|�+�=L�n���X��XO6��J���r��4?�@��EnW% ���=�§�\?�Q+6��������$�	��9Ģ �,{%���ݡI�Ή%����E��i\��4�*���'C'M�2v�`,�dG�J@/XK��"��ߢ� �3M���\@k�M#\4u�>��.wzv�b]D3?K�Y�.-Z����H��^=E�ի�k�6vãI&�:b�@����m�5#��r�*�B��q�	,޼" ʢ��Ӭ3B��!{$m�7�/�F�j�R��c�߁˨�m���8-�:��B�?f�C�S�7V2x�>z1>�խ:%�:�[�Q=�>�I��Q��i��t���r�N%�ꝶ�3ق39Iw�Ȥ0`3nq6�_��=�q2����'~ ���U��A]]����R�@�=@>��^��%]C�~n2��S٘�����3��;E���"P*��6l* �n^�Y ���\�1Y�56�bu.�Y�o�g~���/z%
�鷺=W�l]�u��]#f����������41��k%�5�<(K`��w���?(I�1*��f�ZP:�^N��{;�IN�H/{���!�w�p���P��]9<��`.�&�����Qy���f7����a����0��>M>$Z~W"�n�Oh�w�El��N"J�D��OV7`�2��n�����m{ ,3�����bX�"N�;�jTq$�t�I���!ɓ\\i؉5�\?��_D��2AZ�����=��Q{�9�K;�>�[��� >w�:{:��y��#�e���WX�#�z���"4���s�(3#i"��^E� �W&t"���OR��ч�QpK�`�ղ��x�h�X1w�K^&r@�����>�!�<�_p����$ J3���4~�P͚Θ���!+�T���F��|�E	FZ���o�ԝbj����^d�+��������D�!#���:�7�L_^�
����'�>)/sV�#ӄ���.�dR�B�Q��hƨ��]핞�ѳ���%�Y 	:;n�y�RfM���S8�M�H#M;H�c�5��s�?(#�Iz�PB/�şW�h$z(mx����@T��4;p��]��-?���g���'�J�]��x����b�&S� J8m)�������*���\%q@�?gO��#���{��A�!��a��R]�*����"�[����N�xc��s�������LC����OϹ�=��*w�@�C����������s2W���B�ˮ c[�sz���m�VR0gCM!\��[G�)Ac����Օ���x�E��=��c���VFU���î�5`qD��)�����E\T�i()w�#�+�>��"2���׾^�ɝ̲�*�	;Sr@n��7F��j��nU8�?F��]���F��)ϙ�a�ks��S�o���av���Z*(�"��(Gà���g&~6�s��N�g�AZjq!t��1e�qN+*�����ˁ;p�HȎ?�|�)RZ�t�sB�r�,�ɑ���m��t ���@���q��l���o������ �������jV�ҍd��4y��'�&�!���.e����V�竽��r�'f;�j�x݀V�����Et�?��Xo�s9� "�w���5���>��M�>��⠛��)��G�&������L�XVs���nq�����LQN�`�O���)�M���g�1�N�h�g�Dt��i�|�y��$�h;�;�G���|���'�� uL��@��5���e��L��;�����N�Ā�î�	n9�q$���G�O"%�2.w�y=w�u�8mNы��!�޳*�L����-'?�┎P��\7�I���@��G��r��XR��j�@���-e1`�U2��s��*>���x��9�+���R{C�o�!�-�1g�����vZ��:yu۷��Qig3�����Iwk`��rB ���
�_VgqǪ��R$9�M5�:�����WEÍ#�S)zP~�ʪtU'��kgL�Y��&�+�/��|홢#�T\��MS�=��b��ʨ���NTG�: QEN�֘2�;�PM�I�w:cU��v�"ce��J�E)���i�E������in��K��pU�[o�I����G2ñ�U/���x�AV�l��+�JB�R��nc��z��]-㷱N��5d��"R��Vn]���?G���7���Fe��.�,7 E���﬌!0�UXwU�<P�:l�����o���5�����~`z\Q�
F�F|�O@.pש�n� �m����H��
��d���0'N������n��
�*���e�B�(�a��Pi[�;�L�n�;�]z��\Nq_���R��J�
o��X���"IZ"8v�4�p����H:�[����G8���iQ�=��c���.���u���?��%ovR,i��/���$�@��IX�������\��W�`=�$�h� �����ؽcR� 	Kj1i���]��A�6�B�}����֏]	K2�^�}p`ג���튕a�n��,��Q��/d��ntשތO��V�#�>�K`�m��=&P��^͂#>��&	�f|<��C�7�}��!��=X"f
⛙�Qe��`8�?�Q�ms��Bi�Եj�����k>ob�H�=`x�������j%]�;���B���6�N{�����~���af6!7�P�+C� ȯEe��8�OTq��ۘ� kE�!����R b��ց�Q#a�dmD0誵��4��ȶ�a�o�/$]k����}�RfP�>м��9�x�v�jW��RT�!� fKUs���6��u�zd-�JM���E���9s�jc����۝�1�%�Vƶ,Hv.�fcΘ���ԋ!��JՍ��х�E�`����3�|�ֶ�Af�����C��#�2i_���n]	�ED�("��aMHv��~�4���M'(�t�&>N\K-7ZnC��R���
!�X1W���]ڎ�s���Jٓ|+�@�
4-Ym=�'�E#�|����c/0���_M���Zh�5e%���L͉��r8E�X�q0�-T|	�|�j5"m�Dui=&��Q�*�w8Ĵ�~���m��Ň%��I��q�]m�j	����L�eB�|`W
�%���U���}9�<�Of�x���='�R)5dXO1+�tc�cܒ�F�-�ޫH4;k�p��.&�.]ד���G�K�\o���b;�������r���7n�h�k����mЭz+?��K7���	�Y%� �g�S��v��� 9�b]�x�`�z�y�?�t����oT�F]�>�S����ov�(&�>b�=Uԥ���J�. N`ˑ����6< ���h尓�����Ini�����:���Q����^M��ԫ���2j��o�7���S�\��s֖��dYM�`z����� ���)Mpcwo�q�CQ6&��1 �s���s�|�������O�~���YO�9�&��@j��`_�d�w�	�{i��T����A�Ah�Ќ7�;GR�x:|�%%�����!����+Ir�.�Xf�:�G֌����[^������ `Q�ɿ�BB!J��	�,l?@�b����{~>\��Q�i�؅B�x�Q���G]Ir�l��j C{�վn��f*�߱�2��Yɏ��!�|��>��%tG�h |��©w��k^��l"�I5d��sO�0�՘�����@ye)��[�	Zx@���-bgG�&�Nx�k��K!6���<n�Y���AV�@����x�/Y7�c��IwC��Zuk���k���0�@2s���W�}�J�+�iE�"��N#�F�R�m�%6��ɞU&xʌ^��+��U���K&P)>�ҁ����6}��u�]�9�jwj�mlҩf�<�QM�/Wn�>	�E1uy<�<%� �q�ӺZȍB�' I�+Pp�@J�@�5%��A�Z{NY��,�R�ΎMN󇪽��|G�b�s���c��|����l�H��Sw:��fѼ�ф%���`�m�
�N��|�Ӄ��/�TB����[�uV���ۂL2�4��N�}_�3!u�ENpZ}���$A<�~k�s�<{Y*��C���S�Yr�Ո���ǂz��?~Sv̈�j
���1+<�/g��E�R:�}k�͢�=J@�C^r'9t�b0Zb��Rj��$o�v �"�8�S�d��/��~��Oi��0���"���A��@0��ffj��K�����c�U)�Mo�Z5%iuԡY�^��t���t9d��`T�f�w9���<�'�	H�8Y�>���&�bPp�we�7t��ʥ�h_7qQ����pR��(� ����J�D���'j0۴�,饒�ov'y�^�9q
�+AZǞ��qJ���{.(���#�E��o~��9�L~v�_�dQ.k�r:P$�Z�����#ԥ�3���N^r�kstS��N2NA��O���5��<����F��	��������F�>����+e��e�	ŗ/r۹���3Ia�}�Ys�ֹU�o�6	�펣�S�0[�z���.?��mG����?�<Ϻ��������зȵ	����#[dK@�$�v^�)�����_�):����O���������]f��u�gv�Y�>��cȡ��CJM����o��,�����S�k�߻�Wc_�*���P�6#����$Hu@����o�⎂o'i���$b�m�6�۟��u��te���R`ף�8���F[s&��t�8���I��B�`ݚ�KFy6���&b�Y˞x�����26L[w�����t�{G
�Lt�|�����%�{�c6$�����U�SR6�'��� ��1П��&4�;����Ch���2���/�>R�M$~����m27]a�|&�eg9}�9Ub�y�|<�_.� ג1M����ȉ��Rh"-7�������x���!��f�nYW�q��5�!A�1��dj��n��ƪ\P}<U�=�8���fc���}�M���+�fXAR隻�1@��~�V�HM�P���O+���䑑%�,y;�u)G�¸R�>�����3�2�cF����D`����`��$/��%�w�)s!C�5�����1���&����9�y�L�S����bG�|�
��D_���C-��-*�H<���Cw(ad�E�N�n�����O�q�˪�������C�-��ʊz�?�vo����V�����L)'4O<qhyq�a��5��{�S�5��NIk�����.������4��'�â�v�]�o�	�̯�rF����a8�Ӗ�3`�;D��w�o�0?�[C�/I�a�d	f�[�9��z�0�;0�f*95������G¢�E���L������0r�7��Q��VcՆ�6��ᵙ#S�_��XuFq0��}Q��e��5(��ow
|}��V�����������9�����6�"��hR陎����}A �.���N��	����עmkݯ��PU�r����4";h����s~�����TcFS��S�{����:��g�����7V�y��8�����0�B����pɷʄ�#��EX] ��,�`���V�e�,,)��9�2��Qt4b.:㐿C������d�^����g�۞}p���g���h���'X�S��n! *�)Sš�g�W^k�ܚ�q��q����dǎ	oL��D������x��꺍5w�{�L-�Ϭ�A��p������hI�ar=ŏ�~}{��3'rV���Mrv�޲8��������H����o��ja�%{�cjW'�����/�A�yǼ���S�����ֻl��B��.�;�l� "�P{�7/��jI�p�� �Ŵ9�$���ݏ���؋"<��յ��ba8���cc�S�	&�������{�K)`<��'��z�9��VE�ڔ(حQЂ�-j��j�K�����/���x��	��q_g���?���&����'J:w2%ox�s C����Zӽ�rg�c�^�@�XF{i
 �&6�re!2k�;��������at��5s����A#�B�E���(�,�y9p�[@��TU+7_|N܉j��5�a:����z,��^t���bo��a�(�7�Gr0N�o�,z�h���c(}�q���F-�Y�O��n�Jp�`�w�e�z�����m 5.R�ψ��`|����ρ};�wޝo�"�����?l�e�oŝ3t�zt>C����OGz���.֚��rʃf��ro�����-�mh������5@�;��I�0r��Y�g��0H�(��nA7��w���g �l�A�g�Gڀ�p�|��sW�ɤ�+�ʔ�,N�i��n���ϵt��t�2(�^}|\���e"u�J@!]r�%��,ѽ��3��s��ۄE������-��.~�x���)_\f=~�Ŷb�wc"�F�U��N�7ZF�J˭��Jc:���S-�+z,�˛��v�z�{J��k�+v���qe���{)�>�=~?i<7��xȡ������V2�䄮:��K�.��{؅M�	��~�"�X'Y�ښ��}��pcW��S�*����,ףB��98���O���.�`2�%􅿃�o��nV]gS-zBOAU�F�H��Q�q��<~����H.�d;jf�SOPǯ�z≏����Jô�
Ƕ
����Hێ[9�%���T�t���ph�:��*q�)���4C�h�/�H�x����>o%��K(�\�Ɲ0�l�t�E4�+����ǰ�W�
�T�"��/3�uс	)��n�Nކ%�V��(V�y���#��y[H`�ѤWw6�2��Vo���$2�>�������~�����A��O�PK�	wL䑰j[���2�"���#�g�tQM�;f�P%�#Mw�� ��R_�iڡ�mj����?Y��e"z֌˒�1��b����2Kk��	5���>	� ��p;�O5[
��)��b�	P+�cM�0��� 4��j�
�O�:-[�Q����1�,���"��R}����n�	�(3nPL�J�m��������6�숨�ͬ��7�T'��������<L?s��ɚ��t��v�xW͌��H���L�����)Q)�}���嘹5Qt���u�Sg�)�欶��F�ω�S��.�ŝ��}J<g�\0ǥ:
�R�6�3^�u1y e�_��h�}3��3"��=� �tY� �vP�~�I�x�\����V�Ө:��j�S��~��W������R�W���>��߉�JL]�1���û��I�k���16�3'wD,�ҽM�tpM���~��"��UV�����	GI^*���f2���s��3��V�"ȇ�8�_��\�̍E�?���X^���d�,�"��tVΖސ�����K�X���զ�4e�����h�J����G��4���K�^�C������u1��Ds���S���uD�1ֶ/�҇�.�),b�(�z@��C�=���BVP�<�(t�Lf���B�~.����bٞ�\���&ىN��]���m3��1���C���ԍ�m���/�Þ@U	��"�k���Н0�On�a�~��+���4�	¸��!�D�8,ܫ�ħ�f�Z?�J�W�%�UN����O��TP��d\G�v6I9�
dEh�TѬ����n��0J@�������Aݙ�JA��G'i�:� =KꎧJ?�7�C�i��뻘+�LUKr�~�k*�_�x�$��KQ5GM���-��[~���.9����Z�e`]Fd�Q<�H��l���^ˬؗs����;����h�(����ڑ
�4�_�0v!ײq�c;�V�N�{���V�����9��N7����w8Ri��Q� BX�N�����$5�����2a�.��+F����1��1�?�c�/v��@�%^��؏���B	���|������W ��.�UU���X�h,��������6�ЬE��rK'��Ń��
��m�	��W��{�߱����Ë�l�)����86l`����|��^=��DGz�:�o��Ug/��&Ȇ��
�>��xt�� �=�b^�DL��������� �2��rܭ�ä���eI��R�~�$ފ�
���9#�h����&$ 0�EV�L����i�6��E(|z%�D�@��x�t�$S'K����g ��k{��@heΛ��Z��aX%��(ߠI��g�ǜD� �ܠv�a�_�,���,O
�Z\nĨ���r@�5�	.�Sp(Fo���ׅ�2�HP� b�L�k7�Y��6<��EZ9��,wx85�N<݃`�(���e<�
�N���6U%0n� �ti�ҥw�BrV�^`��De�ׅSo{�/��ǂ	��*���*
�ɟ�'w2��\�3mX�5y����
������f������3a �$���b�?
&�9�� Q��a�5zo���p��1��)8�@&����� ���?"h6!�r�=r|�,�m��������������!U��1���V��1:��=�.`�;�����c�����M��8�Zj���73���R���T+��p��`N����
�:i���3M����^g��"�4�U�����.�I�ctHPu���Jб����n3Ř`����@+��[�    ��4$X��&�$P5Fz  hEp$P_���n  ��    ���  �å
  �Ź�  �   �
   �����Ã�$55M  `���kV�ƭ%a1GGGG1	  KǸ�  �=4'  Q���Y�����Ya���`����X���aaW�+��    P �X_z{��L�  VN^h�  V��^f�Sh+��L[[f_����_R �Z���Q0���Q0�D$�PRW_�ԃ��R�8 ��8 $Z��hg_{X�    W� V__VW���.t���
uL_^�   ɵ��]��X�Y�j`�4N�-�^�WW�T$��Rh!   Z)$ZW�$   X�� �$���ċ ��SPXW�4$����6Vh   ^4$^��^B h�9�[�    z{�tu �   ԹE p-~m�����t�>A�7.�4$��P�B8$������+�X�� "h   [�R��^�$��R�<$P�4$����6V�$   ^��C "hU"e_�    rs�>`���M�ta�   �J��0q�T^^V� 8� ���7� )4$^R�V%��O%��Z�>SS�t$��� �<$��#��`���T@�p(  T��}p�K�4ݣ�n�y�N!��_�g�4g��gF��g�z����k����P�����K$Tm�se��6��ώ���5�j�U!l<k��W�@�P�������F�?�.P����;��z���5H&=j�/�`iL ���w(	�ot�,c�{�CG�uh��}p��w0�)8�|�ӷ��Zq˞��\���4:�N�nm��d��d������Y�b]��]���lV�}X����u�bW�T�����B84��us/�o�
���k�����^=������4®���S-kY���~���L���6�;��_���d�n�\J��4C��]���4?ƪ~-?q3�Ͳ�!�0� ��� �<G�- �8�GuC���ܾ���9V���=�v;�����fE�����A�y�u`�;�4�@$(g���z�7��EB����:���l����u��#�"9�q����1Kr	���5F�3���yq�֩���Δ�EQ({_��6a֩|G�N��}X#竿"���CBuh��u��uϾ?���9�>�����7�<����,�a��?��uu�>�=J���?��O=���~}ո3,Gy�οD��=v��Ku����[��Wv6<u~rwַ�����(1��g�&�݄s�ؠwpǘu�m<>@J2��Z�=��0���ͪ߶2���2�8rp���ϹzuC*�s �7���E��1?�?>@6��/����7��w3|�?�>>A20���8> ��ڨ���P?Ҙ޿4���9@�7��N����ڨ�}�x���1Zɻ�}Es��l@*5ү�����?^e:,@�5�Q��4�|ug���$��7���A�4�����(�us��4�5`� �����ڠ��g���KCK8kꝥ7�< ��uX���4I@=�`���x���%�����{�4A��˭� \�?��C���*0�#=}=A�+<I�<uwZ+DIw<��CpK2+P�<�5*��ܑ9K"gtm�)tS�@,lI;ut|-tI�:���FK�N�8f�KO�-ܧ8Kt��qJ���9�9;KpC��]9�99��»�:��a8K��ˎL=\�:�="�%8��:K@ �ɿ7=�1 �4��uЃ�G4���_��>P���=B��U�����>Pɦ��
�nN��� ��4#�KE�F4h����ʾ4�������4������47���Y��4|������4��>����+��� !ߌJ�3�9��G����վ�Y���ڙ��x���I��]1����[��й���4������l�?���l��l��xl[l��7l�l���m��m���m�.am��Dm�]����m�4���3ЮqVв�{��������4�����5#���G��$j���Ѯ���t����������$9���[��4~������4�����������*��4M���o��4�������4�������4��>��4a������Ԧ�����4������40���R��4u�����Ժ�����4����!��4D���f��4�������4�������4���5��4X���z��4�������4������4'���I��4l����ثd��������������4;���]��4�������4��~��9�dR���,��O��tq��*�������4�������4۾�@;�d;������$���T���6������42���T��4wܾ���4�������4���#��4F���h��4�������4�������4���7��4Z���|��4�������4������4)���K��4n������4�������4������4=���_��4�������4�������4���.��4Q���s��4�������4�������4 ���B��4e������4�������4������44���V��4y������4�������4���%��4H���j��4�������4�������4���9��4\���~��4�������4������4+���M��4p������4�������4������4?���a��4�������4�������4���0��4S���u��4�������4�������4"���D��4g������4�������4������46���X��4{������4�������4�Є�d��n��/>�����뺯���T�ش;�%ˡ�?l�����9��\����`�4-�Z�F�� ~K���02-����������>�~������y8�W�P_�Ŵ�'=����5�~�:���Y���7u�T ��u��(�K�O����+�9$�Ļ���r��=���lgK���v�	t�1�;����ث�0�v�h�BK�y��w?r��x�p��zn�v9��_;��M�u��~��O�✌��L�Z4~OP���#
��~����zu�����nK��*2�4Cl^��2˵d�oa��H��(��d%��+�u�+��q��1^�E�� � �g��	��+���L�ΎPs9����Nj(�$Ԩ\ef��P��_��c�@7}π���'g����?-�ς7�U�����g�˄��6�@��d��P����p����7���!�u��e�o�b_�����[v����wA���ҥ�������gs|!�Qt34&"|�M�j���TB����z�h��d�g�X���!,�?��O��;�������+�'l{�2��Ƴ�e�<����v��rה���qgiϳ{���^T���x�U��C���0H8g������j�$�����!X�.t��L���1�t᩸^�hl�k8���dfm�H���s+?�Ő�;C�j
Y�?�����y��V��B7���[d e�=8vD����34r�]lW�O�'�f�DξR{˛jJ�����P�&�A����s�rI�p6������������7�ݶq�G}?��;�wmy|�;<�]�������e��G���s���KP������w�|�h4=7xV5]s?��#8jԆ�졝.5�A��|�_ ��˥#>w�<�y;H(fh��>���$;��>����O�	�i�-����~�]�4û��>�
Ȫ ���<��~�#�u�}��$!���$~i��;>H�,�j ^x ��#�Z�z˾t�FUK 8��/ʪr����)��#ԏ��g7@�����-䧻��z.0�z�&���l�$T�>WY��)��Ѹ�=[�<4�z^�R?0�	����a�5�#�(�gXe��I�,5x�Rj��t�('�}�"���e�{��$��b܋#2�i�FS�/�):�4_���4�X_�$��0���K�� �.�J��m4��/������_ �<)K@�]14��s�U�4���z�@�v���a �nZ�SQ��Xx�P�;�1xI�p>�{ ���mȴ��3`�ݺ�p禑)��C-�ȭ�u�#iR K���+b�>������_�T�6�5c�"
,	�4JH��ax 2b����BT�ж����Y$ ˌ�椌��t�*��1�gτ:*��:��?c� ˮ���s�7�v��U�jӪ��.T?4]�agND�t���U����9N͞6��"�s"�"
0�oe�ڀ�����n�����K.͚-q�4;"�q c�i贆o���� \v�GZ�K��n�	���D��r� �*�*�ЅY]��#x��S]��8��&��K��t*�2t�95�&+t)�>, T���g�K���JP�@�a��1g�39D���` �~޽�T�d�0DIZA�Q5Q��O>x��� KP�<f�f�ÜN�Uqw��Ej�@x�[�W��`� ��i|�W��s	�OKӇ7D�{A��Od�L� 7*��C��F�ݼ�{|b�U'�w14���� �3�6�Ҭ@mR7�GR�#���̎T �������]�������t��N,4�� K��@�+0���"�Q�R�c0}����X�ӆ� ���.@ڳQ��nm�}}')AFK��M �r�������)@��y�Bo�KjC�O��>�P~FD� K<%�\�5	�)|5}���,G�T�	c�<��JԸJ��m��݉ٛ�Bg��@�{�Z�� �6�׀���P��h��{��"�+��H�� �6��q@C���^�g���� ��~:5ճ{�kѻV/�D��	0�,FKb�s�
��G�XY_O��=ah)_�ـφى@��0)K�v<�����L� K�*�b��I�9:�����
�$�MǇ��-����1ta~��Z�iu>�S���Hp�̀���T;��`�>Լ�KV�;�u���X�CH&�o�L߭��������?�C�@ϫ��;�(A�M�6�j�w�%z��&�����xq̟Լ %�Z ��'��� ˤ! !ֽ	o�tɯ�5`�0){|pzh /nȪg�8�ni�	wn:S�4z�uw}� K�0�>�.�ot�+�<&�>��736�te�^պʰ@qf�>.@I����Zhq3w�<��t������; I�ce�m2 o��#�қ�+6^[>Z�P[}��$�.��	�:����ה���b�;L�?�E �
����r�5v�wm6A�*�Z������ K�M�����)��Vʤj�ŏ��B� �T�;g*cK:F�c��4#ǔ=j4K{��=G�t�C�><=K��0Br����i� Og�yx�9���?c��MUFNi�r8FI&�@KSJ7�	��4��i���H�7
C��,��g� k:��k�C�|V��0�����e\�能K�M� x06�˂^_z~I�	Q�]�C?���媤��� �!\*�6�=�8|�f�0��Ȭk��[$� �ݎN�=,���B3',�|Fi��*�x[��8������ܜ���B����N��UM΃!� ˪�	�x3��u�;<I���VѰA�D��zW�� ���$TR`�֭#�=������1������ �҉TA��L>J�tD����LhGT��z� �ט*�� �AL w�GQy*L'�D3����B���/G�� ��f�>�F; ����g�B7�����5�� I�I��-`�22���O�~`���u�yC:�ᅱK4��$6J�TAC������FЩF��j.@�˱� }uˑ�e!q2
1R��]�� ԲA�u�l �]��=�w�,�Ov��j���^���5�T!���Z��In���U��Z#�ϼ��o��ymG�DH���A+�n�Ϭ@/M#9q�5꣊�T}�8#{�!� ؅;J���y��zw:�z�>��1�&�8�ܢ��� K�2/���U�x��?�
�ڹG�F��q�u�MK��n�Ѹ��;�\B`��H�<�K9 ��]|s)B谘�\��q⬫#�In����K��#���RgA����Ûx*`�N% N�~���>�=��/�u�ӯ����#DR�/§ ���dk�9.,�
ʀ�B�1 �d����Y<�k� ��D	e|wJ�&���s���Uv�����{��N��+y���_N�ρ�@{Xm�9ⳓȋ�d���*��?p}1[c�>ǹX'ԛ��71H=��K�-yC/�e��c%��;	|
)�"�I`M?>��K��$d@:u\oc�瑿b�qã��qxP
�K�}8̺`v@�R
A��jNYtC: �I_C�7� K#N$K=�7y�مN�!];���	Sڟ��� �	�tm[cL<?Ũ��6�S�AC�c�~� �e��{�%Bg*�"꒫�37�L;N���B˱� Ii��)񓺏=俒`09�`���aKz�8f�K� ����x��kk|�U
��'ߙ@�hK��^�Iԃ�����B{��O���N�m�,�(��R)�������R��?%R˥� ��`������Nm����^��=�l�<�� ���v���7���Ѧ��E����~��e���� 4�D�b�� i��++ռܪQxt�u3b׃�H��؆8�Ix��k�CKB{��Y)B�_	���'������yLЅ�ݺ�)�h�G�)�O�] �E�I�*�$�0���0v�' S4D�| K(�̖h}3�ED2���}(2,�ϻ2��	���&�[��R�"u~�}� �w�"��Q�I�ș��Ϳr�D�(�00�KY��ĩN�|h��dj g&l�E,�,?��Ju[j@dE�+@�j�|=E܇7O�`p�6�
��y �S��Z�K����a�g�����l��#
��Zƈ2˙�X����Cz>V=���ۑB0ǈ�6���)yG�Q 5v��K�)�Cs~�#ney�y�Y���7�+���҈ �B!�-�*�=��<
X��$�.`��@�>���k#/N�KT��#�p�9��n�{��3̅���	+�����Çڙ� K�r8*��\R���u��L�S��Q�4[�����V0��<]ͻVC�d��K`lrD6Es1�G�Ѐ�2(�8�$��>��n'��Hmyi78�H�d�M55 K���,�軦-��)] �2���4�O�@�K����	��l���S�R�!B8��N��;K��N� K��8+?�m��^ �]���!���`~ɾ�\K��09���<��d���w7�K�F�&�Km���9we��W�Y	!�*T�ˌR<����Gg^_ ˂��̕�S��Ϭ�k�oR��� ?���8OJ4O����G�+�[{����l%���^�X� ���:��H���(�s�K8x�1y /���D.����cyy ��5�3�}qW�b�1�0�}��r��d�9.˥�Y1�����?�n�)��a����`��9��}KHw ��Eg���K`Oq����t�����'t��x����1��W�}|ŵH2Wu�Dr�$�b��G_L�8��Io&����	���MF���WDyt!�s"��G*�Fۥ�F��~]�92��˺s�
����}@���+������MR�5�S�)���s��D���s ��G�T�O���9a�D�������8<J���d��M�fo����U�yL� �7��5�y�t|s��;��n<��R�Z+|8�r�2�C�v����g�ߡH�nv�ٛb#��O4��}�x�0�mr��?��Ó�Ѣf%�[1�p~�^zK�b `B{;���A�Q��g���U��c�k K�v���'<��_UY�BG�[�������M	G�H��^�ױ�,tu����K�j ��Y��N�\>������V�-im�#N���Ԑ�8dY���&��(M�gtUPŖjq�k �`�����z����08�8��k�Q�Il?ͺ��Q�ȍ��'���T�����:��ہm!C��㮬�sf ���g�3l�^ȳ����'S0ehn�7����g̹�E��}�!d��o	K������]����ܠc %�ѶP�U=ri�K�E �k��PJ�௯��ʌ�y�������� ˚F�����H�=�,��IM�J�b䘦��䑘a ���ԚMK쥛Ii�*������OĂ�O��ڄ��[m*��ҁ����˲��j�t_�D�x �$^�]��'y	���">���Q�5��Va_�_��[�������Z k=����̄;g���4��p��I|\ [$u��س�)�$�
��8��[��;8�Ң�[ ������y���J2����u;�e~�v�5Cvu�
μ@&��,�m�J��YK��l#����h��;��Q�i��
K��9m���]Y���$�x,��o ˱u����*������w���vH��_�W�5�i��H�O6a�ޤ�V [�������	�+��_�g�S���{d�:^ f���X�C��'W��j�E��[T>)*◦|	υ��|�ꦮK|N�Gw����Țwu��GG5WQ�P�M��t��j)(� J�U \N`�d|�����QZV�E��³���Vvq��6�P�:e�A������������(~��n�O�A�8�r��,Ȇ��� :�vσ�G~�;�K�m�R�(�~Y�CѰ0]���Q�ݷ蛡�]s%���4.� �Z�F���0-�u[�y�J�I�C��e�̉1�kmiи=���Ho�ÿ��X�V� ˨D�Gi�in'�i�h!c<�hvM��������bF���Ķ�F���tDKd�M�?�`����ɖ Y�%>j�Bj�/�G�G]7�@W\L����� 2������ؘ��8eH Ku�����Oڗ�����(�-Q�*������K1�1���_t�xz�����}�KbaBӕ�ʡ��$�{�Ԕ���s/��K��4��y���w��C�o���D �;��u޾��n���a��)}D ���P!\��1 �=��Ay�mV+H~@�C"n��!�?���<�sb�M���q��aB�˒��P���e�'�G$B"�+q|]!�R
K���� �$S����'�O�xQ@@a5��せ�]��]o�V�Ԯ�4�V�= ��!\֩�m���	��<�=�د��~@�X��܎@YXG
�Rm�= ��Ьc%ڠ�g�cP��".$�];����=�ղ�� �	�lo{�R�ꕕ���.9�G /b�;>&�!uψq�+�a���B&����?27 A�-�{�d�����U����z��V��>L�Qě�̐���wG8�X����g��Ff���9#♌��6��.����w���'���x±$���u�>������״�H�Ǫ��$�T�>\�7<I����wլ'of�;�ŭ�j��4� �2��q��ƕ��F�ʝkV��Xo��_�,��M���ܞ����ڑಒ� �w=���R�}�ڀ��2��@�z����P���џ��V��4-��<HظI��$�Ƙ����0H���z���I�돈��ҍ��©����a�[wdl~����Bf�D�5��$G��
 ����⭐Um��u`2�6�]���1�r��{���ϓ� K���?=�����K�ջ�۹9������"&��D-4���m������qY�.�E�r�E %���K��}w����t���;a� �
�kfC�l�OpO?��ƈ�/������@U�o�Yfj�m���y�J�=��׿�qFq��[M=��`���\o�ׁg��������(h�NA%���C��4&(�����4������H�����a�45�A�����دKc�|�@3�$qHu2BQ��'�3��|Z��$Fca�������t�v7%��?��ATQ�7�&���>�}G2�F���ݹ��$������t�5%m�6�����XH��5��������_H�����[��t*�3�����~Iv. ��9��|�"��>�w3d��C�� ˗Nt�	���]8�L7�C�0]X  �iVI��4�ظ�v��C6_���-t3���������ypD�x�=�c81]8mz^���t�5!�Ծ�9�����G�b8<w�d�j�)��t$>v�$��i`h�������a<����!��$����t#�=�݈��5�o�2�%?$� �D��ֿ�>T��t3c#�_�nQl���9��˕^����`���.0r�+����ƀ�Y΀���g)*��k�C���!���g� 4M���o��4�������4�������4���>��4a������4�������4������40���R��4u������4�������4����!��4D���f��4�������4�������4���5��4X���z��4�������4������4'���I��4l������4�������4������4;���]��4�������4�������4
���,��4O���q��4�������4�������4���@��4c�T��Ԩ������4�������2�TT��4w������4��uT������#��4F���h��4������k���]T��M����7�=�Z���|�/ԟ�����q����5��pe�����d'�͚���4栺����P����V��Pq���>��u����Ф�[���Л��G���\��U=�����@����߶�[���ф��4v���;��U������������������44���V��4y������4�������4���%��4H���j��4�������4�������4���9��4\���~��4�������4������4+���M��4p������4�������4������4?���a��4�������4�������4���0��4S���u��4�������4�������4"���D��4g������4�������4������46���X��4{������4�������4���'��4J���l��4�������4�������4  �;  3�3ă�@��(��8  ��	  ���	�H�+Ɂ��g  ��m  �0L  �    �˴;  #�����^��Z8xz��Z8xz��l(  V�^1��-   ���8(  ���А��"  H+�P���X��V��4^�����3���O  ~�W2�-l_"��(�FN>S��.r���y���w˴@i8��;Ґ��*4�2p�t�q۹�3�]x}��ZiUH��z��S�n��HCGŋ2�4�nRK"�^�9�y#S��!Rי,-C)R��"|cخ�eS{���s��\�%i���o�-JPƣ��9����Ap,�,4��x�C"	k�ٸ�>""����>���/ڋN��j%p�R�����#H��˟K7��f䁷����18������6R8o!_�K���?�Y?($��*��������2�L��|.	q�P�l�z)�@����D��T�:�I��pm>v[�-~�i�΁�@xT��@x�4$V�<$��Vh   ^4$^�>P���k(  ��X�>���?��T^^�+�E�~nw��E3�wA��`���H^�ƵKمU*�,)����T�0gL�E[�c����aI(�����<�MT���<�M�$RW_�ԃ��SR[��   ��[WW�4E�<$Y_�    `+�a)
P�   ���X������P��X�   ��-�]����ԗ*���)a5q���T$�����E���8���(   V�$   Y�
W�T$���̋	��V^SS��W_PP���ă�� ����UӁ�Vx�,��   ��LB "h�`[�    rs�)|��t��   �ⒾHv�Ӱ�~��TG�܃��D$�Ph   X)$X��C  h   [�Q�D$��T[[��H1�	��H1�	�T$�RQV3�^�̃��	Qh   Y$YS�5"������[�    |}�)~��=   ��������j��1S�� � B�t)������J?I	�W�m.�oO���
��Nj�ѥ�ff�$��V�1��   ��^W���   Z�TYY�$��� ���a�2T���a�2�$� VW_V�\$��T[[`��!j�T��!j��$��R:%)��R:%)��T[[�d   ���8h�q��%�Jh�{ͳk����W鵒�2U��,��:U��r�Q�qS/�5%Z����[���V����,�8�Qd<?���o�i'ά����*R�|$��VW_��h�F	�4$��S���J�����[����+�S��^WW_Y���n!���n!�\$�S��h@fq2�$��Sh$$r2[)$[S+�$[�$����� .T��� .�$V^SS����h#+�|[Sh#+�|[1$[CK+ˋ܋��W��_VBJ���tu +�xy����^Sh�F[[�   xy��7   BJWhwy�J_<$_P�V0���!iH+�XW�T� ��XMa<$_������tu �$��T^R��N)�T�4$^Vh("^4$^SV�ƿ�#��� ���"�^[WV3�^��I��I�#   ��S�)	h�с���+��W0n
vd����ZS�|}�R��_W�,$�   _�����?��aRR���$RR���$S�$V^SS��S[VV�����HPT���HP�<$S�TH",���1�+�[VhNS+^4$^��R�,$
���Z����ׁ�`(��
�����8liL��8liL�t$�V��SS�t$���ȍ`@���  ��I|Q6�����I����g�z�߲���\;C��ä�TL�Ӗy ���<��+�%��M~@�	���Aο�����r^����^����!�����1�/�'�{�"�4�d�H �yh�<��"��!T�Fvh�w~��G-%����Qut,�!|�qvjy�9�F��"~�*E�Gہ�'�h�fdh�����6�s~��)�cڤ4-ۈ*�8�,|��t��).tמݹY�5��(%B���,�XK��W�L�5-��~-�T��gS.�Y.�J��P떕37�}/���/�L�xH؋J�0ԁ]�H3ٗG|1��2��P2�D�k�C�b�2�B�۳@{3L4�ۻ>4�!^��<�4|����:15��"��8�5��*6�6���݀6�4�̻�!y7���7�0 �(T8���4�m��t�g� ���>�GS��y��� ������ �Ѳ�%�� �?�+������Z���0��ɔ����\�����Z5��?��Psw�P���J�2�7�H���m�d���������p�I�u6��=�0�l��	�I��O���H��n����%mq����ݱONM����#����wu����ӳ��q����ۿ��{�C>^ �6�KA�/rL:����I�=ou��\�[���F�������9(��..V�.6��56��9��.E��	3.��iq`�'q�.1�/�����/d�m/��X��.�/	����/e�q,�����7�.y;���.��/b*w/r9���.m�j9��.|�./	*�9���.d�l9��.��φ�(/`��+�^�u��n]��2�K	z
�.j�B/ka���?Z/i�7�*^�ڜ�e̊9���.����z>d/`����L{/~��~͌Zk��,}�&m/�.{��,xX�n�.vݔ,w�(90�q�h!�	pdt�.p��s˰�Y��.OԧN$�9	�.>ސ9�.<�}K��9x�.9$%���MGW���	�,CɆ�W��.A���K9#�.֧��_�9�Ķ.in�O�.Y#-�F���V�T��Rn4��P��.�v-�G��.Q�,�R9�.����Zi�'���轰���.�����ż�_rCѲ��.�)V,��9PR�.���9F��.q�9�w�.�:�.���Ӽ�kU!mc��֣.��]9�v�.��.���ե��.�^���Nh{�_��K�.�*�-���Ӛ�.�j�՜��.��Y��&�.���u��i�26�OaM�q�E���9�s�.�ƱY��R�V�Q��9ܨ.݄j����A�9�.�W����R�'�����o����9���Q�.��-�9Sެ.�E�.��S9"5�.�,�.�}-�8Q%Q9;��.q����7���-�����R.�̦-���� �/9�0P.��W.�D%�S9��R.�V.�>��(V.��z9ѣU.�iU9��T.����^\b*�2C��W�3@m�oWZ��*ˁ"��<_.�$ *����8Y�9�hY.������\.��X3�A\.�9��!MLU�m[9\�Z.ThM��FZ��+.'�iY.ٴ�*�jJ���\��=X.�P�*�(�T[.�H��k_Z.��*/�I�(E^9�^.=>E.+��9\rA�*�vR!d4
�9K���4<��n�5@�����X-�9՜B.�<Ґ�*<��*�@.:�j�9(�D.�WR+6�9+�G.#�B.5d�)%B.3�h+0AQ4F�a�&A�L.r+,���M.I+	���N.�+b?LN.�,+_6�$+ �Z]�M9ffM.�=3+�[�\L9���ѽ�F9��O.]�2ҹ_F9��N.jIvP�:'ft.JE9�dq.e!f�k�pZf�g�ipZdcd�o�sZb~�%�v.i7�T�dӛ��9��u.�b�gu�t�p.`�B9�]t.��+�k�q.}��`%}�v9h_v.���a�.w�O9T{y.�.n	t�xZE"N9@x.��M(N�XG}.LQ��Z�|.J#LZ}	4(H�	��jy@{}Zq�K9$�|.� J9*|.��IZv�(Ax
W[9#�~.(qi�[~�`�E9׈a.,]
N�g.V'DZs&DZp�!�!�t�T�cZw�JZt6�(Q�
%�\]�(��
�Ic.��@Z�)�(���Z�G�(�
��p�g:� J9J9g.����`.�܆Z�ԓ(��L�.�<~)��hZ��f)��9��k.¦�ol.�*I)���i�@)���j.�tOZ�@9�=m.��k.�5�> &)����x}�po9�<o.�C�9�n.�9yI��ҡ�)�qe�Y��Zd�Q�Z��>9�.��.��)9�.���z�|.��8Z�X�)�6�9 �.���9S�.J��)�Lc��.����P׬�ӥ'�;�,P����J'�>�-P���o&�=�.P�?��4%� .P�@���$�'N/P�e���#�*k(PɎ���"�)�)P���ƨ!�,�*P����M!��+P��� ��4P�"��7?�4P�G���>�M5P�h���=�f6P����<��7P����;��0P����p;��1P���:��2P�!��:9�/2P�J���8�H3Pl��7��b<P���6���=P���5���>P�����
�7���B[A�����eV7����� �/AW����
�#��O��-��"�f��<,	+wM�>JX �T���.�a/?M/�\.z�u둳x�W� P+F�G{��7�'nz&"�52�$o̔�p3�C=8q���6�>��4��G�3y��Έ�8���>����uc΀���\J�d�I'v��O��GZW�L��7�	'YR5w�/v�/�3Km&2=m1�n0nn4L�����-P� Q,$iu?��T;qP)H�3m�����q$?q&#�r&"i٪���kw��s4^�}�sL�K6����A�G)M����b�={&uM�Y�l0s�\w&�q
���(Op�?�[�2~� t')uB��2zmz?z/�{t�v&0no+f�Ǵ�J���� ���}�}&��~�t~&$I.��/���$�%%_��� ��=h  +���3�	   ��	   ���Ã�_#Ƙ�r����L@h	|@Y��4<  #��3���Z[  ��˧����   ��   �`  Ã��    ��r6  +����   ���	   H��#������YS[���  WS3�3�[_1N+�-�H  ���   @3����	   ��   @3��3���ƐR�Z������������C   ��B�ky�����I���xF|_hg(4��ɶ"1�U�/-1V.3R����r���6����d:{� �%����Ƽ��t$�VW�$��Q�V �����u��Y�R�h" ������+�Z��$��SS�t$���(�1�
rt��F$�k5����dT]�jڶ\��B^��;]�W�R`$��-O��<$_W�,$%2A_�
   ��6[,]6�Ձ�n�E��n�E�|$�WS[VV����V�7��   ��^�7WV_��s  ��_�7T^^T__�>��ܚ˱b��P<%��s��'����Kë�DlZ Z�>�#�<��h�Aj�rC�N��5��ݧn��=��&Z��']��I:0��d�{䩅��+t���x�<��9�x�������mp��䞅�QP@�V��;�[)3�c���'_��j/1O�
 �(�+�W�����lϡ�t�'��p��+²7����b�g~�4�E���⚸������0-z���B2�5Y  `5�  �    �+����D@@��i  +���2]@��r  ��+Ɂ�~  �������h�  Z�����R�V�   +�#�Z�� ���3ž����� b�;�wTL  � ^�ZR��g�    `%y'  ��   ��H-�]  �   3Ë�^+�+�Xt�� ��  ���s� ��@   �D���
   ��@�-�w  0FYJ�����_l�N��g[>��O�.�zd���R������5�]�6��lR�Z����N��\�X��Q�	���G�?2��G�V��w=J�U��9����ި���;N��*y������:���pJ�ni���E^J���)�(�c�%�$�c�n��)�8�H�zI�����e�n��1j<����mi�^�����u�x��~0F#eFƧ/t�סI=���GSK��	t:dg$�L󱰤�B��;\�(՟���&.��3 K��F�1\�#֚B��E���Ksڿ���W��W�=�N-������V��c�s�f]¯-�x�o��Yڛ��Q����S|�X��+v7��@ '�F�����xu!�a�l�$�]���	Ş �|E�d�g���o_������䋝K����l�,nA1��|ܓ����s����[�+�v��\�4�(�8n��l��L���H�3?�4X_A,`m�J�M��-K��/
�C�J(�q�Dl0|:��� $����$z���/Q5����/�� �4zP	ô7�[�T�'w�,bA��g �A�:(��ZY�#��Oy���@��:%�!)��n�kO�k�a��3F���5'aБh�����1SME*"��'gᭁaF�Zr~F;.�5x�Wy�
jVUʜ0tE֝��P�\%!y1��g�\K|�{¯�|��(��&YD]Iq(�k��:� ?��nx0=�[վ��Ň7�~�Z�����KVt5��~�ޟ�&E�2�~�ՐbMPL���D6�o��:�o	�ђ=�)[�������w�o�[D�i�d���rJo��.�E�壂��B�܃��X�i%�M=3ޒ�?���R1i�ֱ�jk�U;���.L=�?�*yW�غE��ނ��k�b\�������+�4h�t��Tӡ��ߓ�l��Xo�]V� �_�y�����0t�˰�|�<�F���G%��vл��v�����m��k=qR`���a%@:� V�A{����G��c�j��nAwq��h�v�F*9�r�)��@�=��0�S�<u����>5�������<~�M���\����em�x�}� k	�:� \�W�pT���Wc=��z�\=KV�kR�mo�J�P�ǫ1D�hm����������������K�N�`J��� I�mce���l��!��/Q�}�/�c�����g¹��B�T��T�/r����1���羽i�T�&p��q�Z���Z�9�Ұ�����[Չ�2Aދ������x��~�+&'��[��nv�%��xm��ӐL-FĻi���U=����c=�q��%4<8ͩSe�][m`�� X�v������c�53mp��y�ɢ&�c7���<QJ�?�A=%$�2�#��=�kC)����t�����1���v�T̬h'���~w�(L�
�uCjv$
;R=�����]�������	���;/��l����i�����Û�8r���wǰ�h�P��d"��P��9�b�E2.>��(|'���
���VEb��~��Ŕ?�?���	�&Q��OEJ�e��Wr�s��~� ���R�H���}
�l�U�?[h�`�Ar
��$.�g�j4�f`Aԧ<;8���^u���v�G��sXK<�X_�c*	�gl�_�T�������M��$>1����,�c~��gc����% |���+n��:E���?+8�F�΁�b�����_�e}�t-���lh7�ᐒNV	GE��?��5�b��xi@�Bf�刘������t��4���*_��8a:3�+H�ʤW�7WO% k��eN��&�o۱�;�����*�7���A�qƮڔ�����#$���K������]
�@�u^��ۨo�zJ����y�@�x�ňj�]�Ŧ}�ʢ�%�ch�9lo���,*9�pN@���u<m�1��fD�#�u���,u��
x��;��=�h�y��ʁ>_�uZ��$ꪃu+s8'�g/�U������n4T�Y�=��9��L�_��Fs���28��Bz�P!��'��`��L`�B���Q+�ST��f�ne�t0"����>Fk��jk��l5Ob�m� �&����pgBڌ�G�`׎:�m��j�E�N.C�_�_��9���Gz��`F�� �O�d�Õh�QS��J:ib�5��|�%�h�e�}���Zq�,���6r{���P�/9���j̫H0`������v(����t>\�t���첊�o����`QO\�@�Er�h�=tF+����V�F�J�9r֥�P=y���d��W1��NZHlI@	��e����S�C��j�	�ܜv�z�M�é<^Okg˼��}�Ø^� *WȄ7�	�����g�1��ݖ|�H��v��B����l�<��)�qX��w)�]�D�)�z9���Ɍl�l���;hi����Ĳ��D������ȗ�|"�]7�9�hh��̻�ҁp���D������&�	Zd��8�鳛�d���dAL�YКT�cz�2�Y6�"�˹%nF j�����KЧ�����O����Ә#*<4�B�e5�)�,n;Ѧ�ş�����i8^�h�m)�ó�.���R�@���a���	�A�˓�ӥp�F��*��R��r5Zr�}(�q �棗���Z���<2�t�4&��J�V�w�59�QDR��|^������������D���z<Ĉ��`}�.�/$��c� _0���&R|,��
|�����	�|�r��>O�@3�v}��o��Kd��&sR�5?'�Jv�-�9�<���>w�����;`+�8]��D�j�����$E���4�У���V������d���&�s����Iob���$3)�flOݪ�,`��E<H	�?���@&�05�ԠA_V��h����5Ñ��*"1��س�b߁Csc�Cŕ=��}ο�Y@��:������ gׄs�cix~��ba�4��on1=��<��^���*�HNFHÂ��=M^���(��N��9{:�J�9A��a#C��H�pV6�|U7�mj̆//�����E�o_BJ!gJ ��
I�s�!ף�e��^��%<�n�&5m�1���Y�R5��4��(�%�ǘ���{�Cn˸bZ��6����q�N�V�e�Ѓ$�v��1�e�S&��%?�`��_$��~��l1��#���M؉��ר|�0o��v�����\�`��qaD
K>��,�D��"l����8>k�a/�*�P˙h���ۍ��@�މ�0�)�綺�@���S�m��Z�+�	����`�dzo�E#H9л�I 
{��e�������`Ǘ�-�H��/|�����=LY�0�0Lx�~����3��"��/��m.�a&�'	7UA�xPׅ��aw�C��HAj_����pK�sƝ	?1_�y�G�JY����E5����R���s�񚝆���� d]"/�a� J�|��.�R�`��	L��*_*�1�U�H/m]<Gr��<:<V蒨�2պ-���Q�z�
�q�����?E���N;[�I<&Z�Fq��j���#$Y��9��J>�ݸ��*�5]�ZH����u&�i��aR%n-/$��Z�������1P�.4��qsw�Sz�cH}�T��Lgvg$e�N���,rf�c0>��
�Q� ���	[\��G3�բ�a�}�	�(�^6��D9��&��d�	��`-��Y�=u}E����ø"(�9�2^�O�ip�j r�Q���@K�1S���/��%kF�bH�tH���tܟ�!X�\B.�����
̨��Z�*�8<]+B�e����կ6Yy�_�D���EX��>��(Gf���-d�
(4`�����ue����9�M{ƥV/��]��⛖rZ�$Fr	U����'l?����a0���a̙Da�U�Z7����=��O��W���G��x+���X��Ww�%}hZ<7G.@[���dL��>ރ���3���`Z��YJ���]�_�N*�8$8�,��%�m���a�ob6�)j0H���p�3Ry(���w�:��س�#s�7��!p��ܕv���RN�r��d�6�T��n���ͽ�HF=���aA���������*Ɖ4�L�X 7gk�����4ާ�Ű*̢�F$6��:JP��Žl�o�D��� ��B�K���=�
=w@�aAb�虜7_��[8�jY�K�u�`�Z̏��iJG?C�?VqM��7�g��.=��$��(^<�	f�����A� ���R���po��8�m�� �P�s�)�~&&K>��6�[ӻ�������+7f>�U,��U�r� $%���2���a��@&��d���-��CtMNH�_v��8�}w)��j��ޥ$�߷2�3�K�ݩ�d�&�!��R�#�����dfE>�i-�������-o�f�et��|� R����)�[�~��W�Gz2�^�Xo��}ֈ�������Es%+MC}t�;�&'�����7�B����v��#�����q�����k�};��J� i���Y�|���*�Y#;�!����o�h�}4�f4�`V�Z����	��#S�'�O��qW�p
O���I"�oX���fx^�����93D��e��[Z�h�i47M��d��~pCCɗ.ƈh�s�ڰ�^a���U�<�ΣV ��X���۵�� G�+��	�|a���(��{W�2cZ���*��:��� �-��bP�n��SG�M��5h�Oe�3����P�%�̫���Kv��'r����v{���#7XYa���_��;��
։�%�Ĕ�����֨9�8X��(�Y:�@u�/�VA갈��?�s���'��h�]�h���-�u���G���z�������7�;������
w�>�ܟ*��&�
�|�zͽ���4.�7^��n�W6��c��O��"!u�rd��c�"�(�eC�Z�P 3L�Βm���[��%�Γ.��v�!���l�&�ʦ�F5^PM��=�x��,��{���|��Q'��=�������nA���.���ҕc�Y��U����^ѕ�p[�ӌ��f=�4@�7Tt���̤�}�6sf�H;+�y�������M�Y��(�׬\����u�w֞efn��|�T1���E�]�9������eO}I��X�c�}�\�o=N��`WFƹi�\JecS(-Zg���zs��c���E}�2��F
��p�\1�B%�����Hr�1�W\�	sW�!��O��*�n$�xّ-�|����E2�5FB�!��x]��N he�dr����8+:b�&nb���	{����>m�����FF"ۢ�&���Zۊn���w�0�c�V�7!<�+F���u��MH��h�N�U}F� z��+�ğ1�i�5�������i����3C�Nv�Vհŕd�VM uD5VA�q^��xFmd�<>���F�(\��/Mǰ�R����*:!��B��MB�OGw���dt`Q�'uTn
����'�������KI�,�$[�_b�46i���;$o@4ۡ'el�D�U��t|��X� �E+�i ���On�Q�"6�]� `C�'���:r+�p�Ec%��Kw�e�뇮H��e��XT��Q�]���{��6��]U��>���v�p��:p-���z=|�x��&���m6��!.�����g�J+�֒��B�x0*��o�Pa��0������3�����,
�VO2��7-*���r40��$���f����,_�����-��Ѿ��g"�����4gUY�?�_+x���{Kity:��L(���`�c����6TU)D�qO .���Ww.'�n,Z�[k�d�|�3�j����}�@�o%k�?���ߘʈG��(	s�H��a�8��G!̧¥@�i���[5��(]�1+`;�+�"��k[����,�����z�v @�n(�^�8���3/lQ�cPt�[bR�?
sf˕��n���%d�!�y���P�VV��ρ}^?���rj �H�����luV�ԝP(���K����^Z�8����Z�{��J�`�\Y�'&dN<i���À�������Y*$����)�j9%ܚj�;2��CP��O�Vl��n���H@��q�4��aab='"v�D���9cUz���'�����j(������ŉ�wfVЃZe~T��B8+j���Ү\b��Q���c�4�4}ϸ�P�Ҷ�R��i*WၨuK��5�s�tҺ}M|I�F�7��F��r��s�Mvx��LŐ��H�n��tPF������f^w]��a\�-T<DQ{����$�Dr��%���I��Az��dt	c��c��X-J{/)�ڿ��^y����G�Z���L��4e�e
�a��ꍚߙsqbp7R���+y��n_�C�>�!y���i�4�s�yϼ�Oǩ���l�uT�0n����0K}�Tecw�P꘬�D�8��b�!�YI�k��������m.�[����'�
/�����YZV����|�o������ y����� ��vA]����Ĥ���8�c��++u��v�qV���/��J�\���t������y�ҟ�&��ï�+)�I#�.��vP���?�;í�F-r��$�ٖ#�dP�/p /\iD�"��Zc�O37p<��*��xTu�ơ Yq����	�8[��%��H���+��F��C&��}3p8��@r���P��.X`d9P����yGt�g�%F@�g&T�ɐg,���$o3*.����m�P@M�"N�r�@�_�d��y�V�H��$�?%��Q�����YT�e:P�o	{��f.��6�0CU���PuSȗ���5��0�6$r&�xX��K�R-=��rV��^d�Z+��f��N&��a3�ɸ��N�b.K�!�BQN*�9ȫJ݇@��1Rg�>P!ſ�j�CJ�T%�N`��'��F�V�vg����rK��I+z�*k�o�bяZ�H��!�q�f�7��BZM�8h�<?���C��dye�y�03%,�[�oHT���j\�������$��H������dl�����[S�sW��D-�S	�kdևLr�Y�jZ��l�K��V6�N��z��4%�z�Z��ȺҀN�&��m�;ePɿ~��z���a�Y�ӣ��XS���al4$��B�Aks��>� ZTo˱��F�t	4���K�A7'X�X ��U�1i��� �1�:6������B~T:�lP��06���m�d�>'�@=��5�f��0�o庭�����gA�/Ra�?��o]ħ�J����h�Oν�"*��CS�'�e���Iײ�5���y(Sڬ���sW���6�f�J���fc+�3����H���w�e/����Qlq�:��Q�v��<�"��+V�����ǈ��ۥO���`w�ANm�i����!"�zd��'��!��7q�J���H�	���i=ا�FW �g�x��n�s����?�W�cK�A9���߷�E���-��R����f�X���(�a�e �Ǫz�U�Tx�~/m���Ì�W�ƭx~����J_�e�b-��{����q���� �B��,ϴH2n@pV��
?���(E�O�0{q���%*��y(�{vy�,������f9~�#�`�g�{�I�z&[���?�����`�)�gTI6E`z9��[z'-�Ō�:�px���������g�{����57�:�^�1�4�Tz�`_��t�޻����%K0�?>M?�~b��q�X���ɜ�!7��O���q���~�X����\ ��D��M��}��G�Ϛ/��\aB ���{;��j�/8x[�NU��&vɏ'���o�(�� ɍ�=���Heb�$���^"m�/�-�%�-�ή�<��Q� v�/<m��@G�y�yl�����+��}�G!a+����7wYk[��m�`�;P�c�'�ϕf�g�I��/m�ّE#��oؠ�"�éS�w�ĸ8u�J�U��G�J�^� Rw<}�P!`G� 	{�b��Q��{`��������)TLb����X��Z��p�@">�b��1ҷ)��3���o�g<�^[�y+\Ⱥ����f��ك8�$C�̻����k�/� m�ؗ�dJr�U	�xy��IS�YN���:�vT��S��Q���k��6]�Q�����5XX������}]���#��&V,3~.RW9�z��B�<�M�s�(i�RZ�-����4i��M	���K��C�K1�A���_Z-K��)̍�~�#g��Ө�S�P��{����К�-�)�׊s�*t��&���7��3�I�-�k��z�AN�h���l�Z�8Ʋ{س�k6X�s�)H��)=�U�U��g��!>�6�N��F�V�[;��~���V�:�������gl~~��2�/�x�t3a��0E���j׸�U2T���ϓ������h���oҊ���Ԅ��<�I�0A���]�����Mg�,�����=������.t.K�G�&�ƚ�ŉb@J��=J�z8M���� ��Σ�	�%��^�)�:S�$��{��8��<n-���
��*3O�4\BSeTa}6�I��d����PA^���� v�����?(��e]:�~�����,����M��S����G�|7�O��EMߗ Sbs-�R㏧�1a:�AS�AU�E$φ��v0-A ��<�J�wv��?����8��g�Fj(�z�s��B�������P��T�7��4O�����5�'H+�E`�ɪU�&��y��̉Y �x��<�P��0N/߾�!ՉՉ����1L�h�$����k>w:q�`�b�Q���Nk�7����(Y�M�s���$Qk�50�	�c�L�%�$��#�!� W�����Fs�[��|�㾲��:�h�F��C�$�1�sS��*N�E�n��� 8�o�
�hVo.�^i��ۃ��W��}pv�-?�o��6"f[�v�{���W�+��ʪYofXw�����;E����pz�@�Hh��Y���;%��ġ�i���,t���l��B��Ч8[����*�o�4/�s�p���2�\٨�Ab�(�BX0��)ښsؼ�}.��K�6���3%�nM�{�<��!�c,����1����kN�8���.��bG�l��>����27 [G�8N[ 	�l;a>�3�_]��¬C�i�1����:�������p�@i$��O?����6.Zo�{�@k��¶0 �yv%�����&��r�2��� D7�Cwt�M9y��#�4�d{�o��V�5�W��U�<:�6.�~��AZU��鏗c�>,�S��cE�~�&��n��m��d}?$��(��,��\*��%G�>�ra	�O�n��"�5gN#82x�39e�_6���R��w5��w��tѴ���ϪB�;�&@Q,%����<�g���t� -|�����f��i��y�k�Z�
����L��zS�Xk�|�s��KK�yF���gt�GekH�Ed���v�N%D^��9Ɔ�i8��8)R���sG'M��-ؤ��������T�#�iQ1�@��U�g�
��J�5�����0�
�5%3�O���w��G�)2����_���Y�� 	�n����d�����N��
Һ��w2��߈���3�2`��7X�R�2���z���ߊ���_��6�ۯr!�����FI�h�Q��{
�6�4V�Z���D+a4�\}����}�:%AK�x��e�v
����[$ZGG�4 ߫�<1���eʑд3A�h�/���R����V�s�?�E^���C �T�M�{���h�C=@#�ZSU)W���cf��B��C���_b��g�w�c�x��2d�e.�;���ì�;�Ey��x>����خ>����	3�gЀ7�Y��.,.����]�U+gT�C�6��J��L�|�N�o.�vb��\�hxjLk�����ol��8�va��:�J�8��!��.q��-�C�
B�ǥ�ټ+�o�v����esM���h���j?��d�I"y���o�l��V2� �~nȝR�&��T0@���c2B9	� �7ſ�M��̪~��i�W������'c�0�TM�h����<!�?�eѠ"�/�e_m��W`Z�M"�$Z�+`��*:P1���'#�f pMF�y��S�3��%�/�Ŋ��o�ʬ�ƒW��	��3�j���o)~sRT�A>1-/� �͈���Ѻ�`��$B���z�cțH�>R���_��l����T��h��;}RG3��vC��O��y�4���VBO�^'�bs제,�����]�>��<�m��Ѯ�P��;`��S��@s�D�)Q�~��ʫ3}/�Bl'�^T\��n��Q�Ú6-�����ώ�پ�_-~�79vPl�b�/zQ3cO&1;��r%�Y���}�C`H�ӆ�R�W�;)qi�W�(0Hj�oa=̵��<V���o� ҃��B��(kG�m��5���x훴j
�
YD�J@�%��g��G=�����X���1
���+
�I����eq�qe���`i{+�=w�M��k&�>��Q$��d!�D����,���x+�m�{�k�����������d�V��ρ5!β�d�����7��O��-�՗X�E�wx�ót�$7)d_���c�-�N]_��.�:ݢ���q�V�'L�̝��؎��6�q��0ʋӶ��.�!� ��@�tn�%d"��A���k��� ��L��Y������l���e���"%��G���˄�Wű��>��QD�ań�(�g}���D����ՙC�S6�������X
 �P�p��<SO^�_���&��?q���d3QD� ��$քN���]��'C�x�h�E�-�B+��p��N��\T=ǈ�7i��k�5T%��v��tH;����S����)��M��Æz����nuc"Q�5�4~��|�J��ȂE�-A���)��Z��fPژ@�U�4�+ө�z=�+>y�Jx�	�9�ם?�<n�$�b��6����Sd��$�"�f��W�k8k�9^�J!�ƕ�KC�����1��]N��,�bYYu	,[�D�T�ʧ)���(x���=Y����:u,�{��l���O��u0rd��C��N�ӑ���#�>b�P�qB�q��E�c\�@X�PϭpR��h��"��������<%m�B90����@�{�ޢaW�����9ċ�:+\ݳ�ı���*c���]�Z�#�2���
w�v��"��1�J1uV@I��]�H�����Q�1�
P2;� ��:��,�'�"��"bF�e��CE�w2�kYI�K_~�Ac�ը)��Fa�,��Y�'�<�goܩ�&��i��8E�����Ӛ^]bw����������k}a&T�Aغ�y�i�>9x4�J���>5��,�]��B��(��[�zo�kM'��Z��P#��S*P�ʆq<n uԨ�ꔄ�@��Ȼz�Pg�����4����h�Rgt'p��77��O%s�*��Nm�>��Y���;ZXEh�8�'�o�~��/�ӭ�X]Qў���i ����
|x�7��T���4>QFi��?@H��Y�@H*�?��!N�ę�F�R_����GA�&umm�5��{9W���9J@+J�Ww�מ�����g��)���R>v͒䏃\ۓJ%ڗxN����_��ͰcZ�<��~�W����xPP��o%EW��N�44X��Xo�a�4��x��d��9�`02���ݢ�C��y܈���>�ڷcS�W�+aF�n�b�.r�YN� ϣي�Vd-̏��txz�U).�.����1N2��jl��卌aPI����h�H���b�$� �Ōy�&��5 ٝ'�X9)��c?
!f�a��ӳ��2C�����쵺ʘ0%&�p�f"X�*���5��!�q��R�16�i�E����iK�Z���;����aG=E B�m�nu�(��Z(H�i+R��F�g�~
	ȿ����X��c���/p�+���&���k-!�o�x���X���yϺ#D�u��oq�-��IO��̩���M0v�c�y�� |�'�m�G�K'cM�SH���>n[�q(��<�+i@
�|�D��8dT��G�.��(�G��"E�4ك����!�����Dy��g䚹���i^vݽMnm��O�@��;�Um��
דK�M�.ň�X2�Dg<w����}��qc|<,��ި�n���̞��B�
�G�d,4H�Uae ���h�,����ov>t��~�hK���{J��S��,Z*S�X="���]c�j����)^�Ɯ�B��52���r�[(���b�g3p����c�:��%bF�zHE��8ا��i�yQ�����=)sD�n�fP�Ȥ�<�z^��LuDk9�%m�ШC���H?�t���b�J�M{����u_�306!�+�=�tG�?���u�yo�ڋ��=��,�V���1�y����;\�;^�u�pA�{Y)HS��
 ���3��\a�m��8{��(PBG�`�+�D ��E.��dR���z)�ȃ�a�x�g�~{EQZH��yF�.�E���WBV�
$s�J)�ϑ���k�L�s�CR��3tNerG��_>nw���2RR��UH�iEt�v�_0�'�"b�]�E�V�=�`46��m��it�.���C�B>*90,NH<��n�J���	�قU�S��USR��a�x���e���C���3�U+�t���/�������w��6c	
Do� 5n�r�=Yv1�,�ם_h���;�<Yκ�(��s��#�BD�ۡ����������W���/���jH��>Ă�������i��VH-g�{mmCSs�Soh��$��=(�!y�ެ����Fګ*=����6&b���Y1��~�ߝ�L�0����@�B;M>�u�]��w>&�CG���Кi����4mN�%oY�:а���&i%9�?op�W�4��]jv$�����X��H�p�����}y��K���	m/"���
"�9���ޡ�V+P�Cj��5���=�j���28x ����6��(f���0�80�ر�����K-!ΰ C�Q�]��
�N�=���P!�0^�M��0���Y��.k.Ik���Z����n�:����n��Rӷߥ��c#��G
�i�6ٌ�ue�Ƭ�6}����)��Q�s}��qP��ДN�'q �u����:.
j b����&�P<����n�"6
a����2o9D,��+?+�{���`�/�E�k0��0�N��S��>����Ђj��	:��L{c'�^���>�{!xi���Ԣ+�%[�]Q�Tb��0/P���}��g�n���eE�N~D��p�h�k;'M��H�?� �O�v��Y��!Rl�7"��of��:��5�pU���H�W��+RX��NU1���gy 9��Pl�ʷ��+VLVsl��
���ۚo�zܼ>�t87S�����WR
i������s� k��p�׿�}�9�2c"�j�����p������&U�rLۤ���P[��Ln�-�N����)����n��������Y�٢�\U�}�QEN�2%b�N���-�>�"��8�l�\�uSm���R���V����2E�W�����-�2��S�d���?U��s�ղ���� ��~H��v#��$xd)����3�/-���j�	���ĺ��p��s����Tٝ*1m�Z�0��e	�J�Xy�f,�s&Xd�]�}9���Y�m�n����$�]C|H�ǈ:k�kIs�Du�,'K�������:pΪ�g~�4W�y��N���Q�1	s��-1;R�Q��+�ZG�����呶l:~�>Jq�ZcK���asNo��y�2�u�
\�&�C��=�I��'���X��je���'%����G�.�-f5��J�k��9������oV���]�,�����3�m����=�|���G���	�f��J�n_3����`�3k��A�x�3H��[��H�dC��38$�
z��i#.�ʞ��D�9J f��Bs�R���[�����w�1$ј�!Sn �,B�`���.DRE�+�fYD�1Ҹs,Ƅ�b�~�4E
�*T���+L�Ǻt����O�[�.�rM�j�Y�*b�ve!��f���,���?PQ��Y����?��u��"��69��(e.=0�;�e���a~ 5��NhV;ځBP���[����b�M�M-���t}K *�[/%E���N"x�nv<�1�x7#�5aJ��5=8���P��pjTLGK|JQ���C�ȍ�����s�@^ع�D�Lҗ��}$+�3��c�0%{��dM1��޻]��h��՘~�JI��j��?�pX�K�0�F�ӂ^��<�����~p'��3�����
C�� ��L8�$���������)�[V�,�En���P�����4ﰴr���c~t�%)�s��� �(�Tb����0���G6> ��9�+�Ԥ���+`1�1$��� =�
� Ig�B�V�ɞ��ss�X���CQ�i��K<��-x����W�z�~)��P���[�y���O��*�j5�|��e"���O2vv��S�~��*}��d;)3 �clh�$�zΨ"a#྽����{T�V���-�[Uʖ�|��#���6��tV�q��
����-��F�ŕu�����`���� �w�ש������A� �9gC��OZ��鑠H'<��Q�׫%r��Ż/�a��P���*0�u<iv��;K��Ї�(4����C �`�5���8F`�[�y��N���]� ��"�T�i�$E�#��A�a���N�~�9g�鋗�d���z~�qӔO>��8��!7v�h�d(�Ly$��^ur��fp��M�se�<g@q��E����j*ߒ?�/�g�2�y�S��/ߤ�\Ʀ(�W��A4`��P���%8�:��P�~�>j��"�j��!��?������&���2�I.�_J\*7-�_��Q�+��(�ԚOo���n�_=����Gj���h�*�l��G���;�T
'�qʓ\��5X!��Ul�����i31�a���BƣW�	l@ō�7G��|͇+�=��u� =P��m�bi��@�+BP��[c}%<�'0��^�)/��ȡ�c=(Ēj��ڢ�c�S���"7{H޲��H��ӡ�~0�������R�����Bd�|pc�Zi�[�o��w�����h��}�f��B�ָ���!�~J�=�F��B��_��'ٻ��>Ph~)rAhR��ýC�Z�O�܄�
a��C�W�`K��.A�8�`_\P�9%�xn�)��ׅ����ؤ)A������&B#��Hw�Q�٠#��RVs��$���+�_�F��v��(%!�ao������JG'Xs�p�7���๦,YY߮�7�#����D��.�i��X�)l5�.�d[Ή<�,�g��4�ֽ�R�j���{gG,A�� D>�^Q� s����)���h�
o$�Q.).�PS�*Vu�B��ܞ�X��K�LH����iwksE�V���2�B�v�e��ڸA���q����O/��b�~V	�0�W�����+�4���8^���)��>��1�����Fm0t�{���o�B��u��(����{Έi� B��o���%�a���9�/�C��]H(����5�2YGu�o��F��N��s�����G�g�AN���A�G^��-�n���E��РE��,��!A9q��QO�W7 ���̫B 0�M<j���Oh]����}��Iz��H�@NW�i�I��&�z!7)f""b��w"22���3��$�L��31�85w�]u�h���˺��^���X����
1�y�;���!fۢ��wr��b����ZTOE�
��ek�m_G�L�pT�4��R'k�B�fJ�ܶa��%��VXy,s�=�We/�>M=��NW�x����ZI�̡ў�It5���z�*��C`���hj;�&�,�lU��`*b�n���HT�6���}k�I6��4Ɍu�1�.Q	%?�;(���սk�d�[�'we���R��j2�y41�K��wn,���j�>Q�}�>$�[�Y��>eo����yO���/Iug+�;���v~�b�G��w"���9����AW�;[F���\��,��\���$ZOMiN�<T�Ģ��6F5'��X_��!���w���yg�+���E�`DD!�����suѐ��O���#n����u��Ͳ�$�[�]~��Z���&�
��� �O�2n�.@�4���q�*�i�^����b�O븟ZJF��ݚŘa�gil��u�ʱc���]��~�zu����:m���k6kq.� ��}z`��.����Z�g5s"���Bω1����]2/ٳ¶���=H5-x���W`�z̰D2�?B���n-��,8�Y��������E���̓��� ό}�6@"����{�B\�GD�����83(��A����C��K�W�����^xw�'b�#���2��Cٞ��w�2�i��A)��G��8�~x�4�<�N��cT�>Z즟nӉ������w1������h��?-�����G�m ��!ٚ��Mk6��S��������I���VM,�0$dH���<<��\�>�E�t��X� O*f^*.�X���hǖg� �!�ߪ���I�2��ly��
��@x>�F]�k�����:�-aY��m�j�\��xh�I�]��u�'�	-ѯb�M*ys��FQ7�a��u�(gP̪V��,b�z���^�t�ӺG��|��!��k��'�"�D��}'�ڀ��͎�4(ccD��,��C#0�3�o�7&l)2�_FZ�5!\?2�eiƎ�RwO����\2�^�ل����]F�p�]h��)�h�9�H@�Jp�e$өZ2����#��)k�i.�$>��]ݖ�L�r� � a�2t�IFd��v�*�tm�?N�e�b3#���U�/��R���en~[l��K�"
xB���3��U�Ȥ���G�
�<�P+|Yk��a��>k�����hNL��_�NhGg�b ,��]��ŵUW;�����F�t��j�a7|<��c<�8�7Q�����eqm��":��$HccY��S�Tըጠ&;�I.tӥ��L(1_���#J9�Vk�ͺ��X���;�#;�uX9JkKg�$8.���;�e�/�g��{6�@*#�r�c���/�=�j���\�&��E+��ym���{�����~�#���*@1��lY`���,�.m�73��7.�poC hP�.���s�v\�X5��V�}��փ�ߪ�ҥ`mW�:[�R�? 	�i��l��l@+e�:��:ӽ��v���V*R�%LC���
;)l�Ԅ6��9>&%G`4�� ������0<ó��H�$�Eϝ>�U�N����������#&c#�� r����V{��zޅ&�� �Ƿ�b�ت5X��_�w(�I�E�)G��Ql��,$�%�l)��X�3�"����iM@V�̄Iw�.d ʎZ� w���9�B{{r�*�gA*u���%+o0�iJ���n���!_�W�A`�\��_{ǚ�U���&���Z<qp�Ļ,]1�>������� �����b���-�K���a��j �X�Dz�[�0�ip����|w��tE���Mo�Rg<�b�
�F��LHИ���9���]���0�[�T��_�h��n��E���*����<H�����c�,��BB�J���b������]^,WɆ�@c�~ltO@qIe3~s4�T��y'�v�.$B}3��m(��Q.�rb�B�<�ֵAx�zC��p���m�* �_T���2�(�p ��x0a[<�4���Ğ�~�-�4��y�hC�b8��M��D���|	������.�(Ta��l�fۍ�x�:��@��Η���B�j�]:�L�/��7K&Xh��]o�R�2,"�"e ���4��ޠxCB����(ʯ��;��>�~��GV9}��<�� a��_��ޏ�qFl��� UL����o��q��Z���s1a�������.�|�w��:�oc[��s��r�ĤR�4�O��$���D�O�)�4�z���@o�*2pM?���'G�d_�4d��[�÷E�혠��b.�eZ-H��DVF�5�i4b�����&ǹ�Bn+�F�s+�Q�eU�_�r�a�宸���3~��]����Lx
����������J��5)^4�-��wg�M�(�:�_����9�	4$�I`��[���kF#�LJ���1��X�6yd�{�$֫ec�Ϙ���
t���3�wL4h��UO����p4�1�Æ���8LS�08jrPB�������[v�a��	B����~B������'�ƍ+EC�5�dc��O=ܰ�����6K2�� ݇�;�D������B��V��F��5(�e�8:Q����Y}�������x�ai����p^��Lg)���b�a��"�Ek*V�n5=�f�0~����`�U!����ad���D�Ҷ�=W��ֻGy �ي?���~�3z���/M��u��հ�����j�>&Y�y��S 4m Q	���~�Ҹ}>;�hۘ�B��&�f9/-�P��4JگE����>8ȟE�'��FK��o0#���J�}UW�Q�}?�E�&��Sh)�ֱ�~��2,$z���_�ro��l�������TR��c���<�}�-ߙ�����z]��,@� �	�e3?�,l�U��6��t<�9���aW�z�	dɑ�`�r�=].�C��)�aA����+|�7d��)H�W��Bē�+ ������;����|kS�*99Z�����c�3�L���/��ҙ0h&q�Ȓ}��##�BY0�7|���c��D�a̓!	�,�Q�28Ѣ�$iӔj1�҄������Tl��SCY:��pm�wH����E�JƳ�ĆTBL$�(�F��}����4x�L�-���ԃG��c\���zэN�S���[W��wx�f������U�B/�2""ԯ��>���Y��-w���zx�VAMł� (�%@�5]�8Q�p�@W!$��!G���9�wc}���s�M�'b�\i�r}y ��sr�i
sy���D*`����g I�����,I�%�ׂ`jZ���ETq�k;9ktj�VϢ��8���Ӛ��,hm�CXz�.�nX��i����ԉZ?x��qpm댅���V���n�X�MLEʿ��@�R��u��"��$�r�G 3e����
��^���+[2 �y(1�.h`�!B3��rX����tUk�Z��nL=*�$<<Z�5�����Õ�}���c���/���|�gH�rX��ۭ�h�����*�L8���ѝ w�x4/�̄u��ܱ�]�{"REt���$�tL��'�!O��ɏR��5�~�f�[(��2�S��v�P��Z����@����!�XIٞ  �*#D���4i��x�Jv#���Ȑ�'�ʆ$_D����,�=v*c��pXm���%�m�����Τ��Y��]�X����S�{�"��*kr:���(��nß8�B{���E�w�KSl�A�:횿޲-��F�0A�Ě`-r\� �ɥ�Ow�8� �
�~��H�akvU΂i������Y���g�2'�	 4�t� n\,�[�F��M�{R$Q�:����)6@[�O3��(pO�ɆQh�a.�[�P�QR�B�^ҽo�yNוy��%��	Z�5'�W�s\�ҕ;.�ϵsJ���}&{;�44'�[c��(� �d�s�n_E���a���Uݨ��(Ǜ��e����v���%�V�y�#�R7fl���6
�Z�������7Ɉ>>�r,���S�HH79���Թh��r�QDX� >"'0N�1J����eg�>��S������}��A�7kx�}�#)�jj�a
��j	�d�[��fPY��W4S���.-sZoYb��؃�Fj^x�ݙ1.�ʸ>��1���� �z0��f�ۆ�x��8� D��	[�{���R�4C�{��9!ŻsB�a�2���E���VUY���]$�-}��s��	������GzUm����f�;񁈿��GҴ���q�j��u���ج��䲳λē�$쑪�I$z�Bb�x�FhIlΊ���&X�H��Q��J�n�d��']L���r~W=�]x�����o�s�]�T�%�υ<�2�dt�D�Gn���� �#L�%n���ps��̶�V���޳��i��wܬ��š��9l�k�Y]�p�F��ڳC_���~*�z�Wfڪ� ����s�o�fi��Ю��Xx��5��lZi��?��/9)ka-��� q�zc�������X�~���: O}���F_�h�A�hs��?T�Ă2&��'
�!9i�ѷ�IH�b���_hGđ��]S���3~�+sF��SQYc�^i��Jq��}�o`a�s�p2�!Å�h2{��^N��tj��uMC����bB�b�2�e�ܲT~#���c�D�K�Ů)��~��~�+$�)ٝĮ��Ւ�J-�y�3���k���^����FM{f|Vqp��ڻ����5o���U��ØHb���L�����+�JƏ,и�����i{e��*_Dؓ4̮�L�$!8n-�Bs�h��o��?s~�똂�k�=��}b���'�$5�(B�1~�:�|p�O�=���Z��.������r���q���ݟ�la��R����V��*�@����Z�3�m���Y�t�Z����f�����Ze���KUv���oH��~��<͖O��h���l��0�mN�4ж2���ZAb�EH��`��C_��=��jVj�}	"��M�b�_�F#u�&�Iݠ�o9�O��&���k�䂬���f�|2R��Dje���Y��<�r�=p�p�& �^"`�P��v���cZ�c�"Tq�f�J�(�~����NtlsxtƛP�ji���OIߚUv�����,��3���:8��Obi��}��_�5:a�����V�z�)Ѐѵ��\1{�FgZ�~9�´�6���B>�	ޱz��ܯ��Q�lo�\���E �I����Oy��b���vГ���.�����n4k���F���f�w�P���{]��i�^�����6�/�~�F`�2�9��n�"�Spjk��;�2�\���R?���^�c�s-�u'��rv�=�M�1R��N"4�۪7(g+��լ�q:���^q����y%&��� D4t�o�#��!{�Η߰0hᗔ��I;p!_ٻՎ�V�j�<Z��2�8;7Ð�&H�y-����z��+�;�=�s�J�E(Z�
��VL]�T�k4�q?���%�fqh��7V�aPEm���{��Y�K���F���,��,�"�bx�1�I�����)��`|.4yp!eC#b�k�<��B��h�jUɖus:�lH3�z8o��(�d���}^�c����?�-T��(�|<�[�k���"�;P��Lp�=d�����^v���yVQ��I�)&��Z��0�
�U�o�%��ܿ���7$@�N��śSE?����L�0B�@+�3#�������b@�HE�;E��:9ں�z"�9|���V�;3pSO��(8:�8f�уw��z��S'V!�),Rنt?�/��f��z=�p��Rvw������Ca���i�������'"K.���iCE�/�׫�F�	�Y��U�[Y� �ap�� /�Ў�ЇmU>*/�r����K�A��W��	U]����?y�����aU�����&^]�XU%��7����i+0���u̳�a��j�إ�n�J�ȕD��T�-: �X��7�D��^�(}���S�+X����RQh���oϽU�3�Í��f*<z)���3t��h)4͇2��]J}�y�����z�H,��dH��1tރ���L*�3&+C���b�[��^���O� ��k6\�d��S$ih
tBu�|d�PV�/�&HC�^
԰�|C$0"��x�ƞ�7�Xrl��Y��_��5_l�pXV�Vű�w�&N\���r��J2�)�R�����?З�/K�eeX@ž��&%�+yj�\�����k$�'���� �ǂ��y�H�a�+��k_�Y�uk�z2����;$��j_.ȣ�*t�
e8K��l�_��n��֡���F�Fw�"�76T��*J�t:-�n�5ڻ�����w���fS��u�>��#�[+l��x�9qXĊc��/��,��A��w�eW���	l8c�!2}��^�2ɳ_�N(��Ц3�4x���k3�����X��&�YÁ6M�5��4[��d�E�m{�j��8�4�>�t��˙<��������8%_���t̽sy��l�h�}���	���<Ǳm���6s{[���m#`S�2� 5`<)m��tx��x	F{M��7�`��	��w!e��]ma(�5�hw̛��)�[���&�ҍ�&a�h��+rg�+���'szl�P�x�P�T��������Ƽ.�V�K�.gs�--[��x��`�@�g��\>�}ʤ��im_����@�h��O��H�Ӡ�����u]�Y�P�cA���0ڦ���<w�u�����օ�A���^�+|��"�T����G�^�TU����u?��ʴ[tö�-U~�d�޽�� 끶Z�O�)�@f���"�焃<�p�q�&/�/���<����A
w�H	�]�t?��|83�ge�1'�����qʇ
.|wWJB��ʫ0F���k�t�I����.��s��y@BS�TÕcm�S$��=ˡU��.��� �(}��[�>�ǞN�Z�
�|A�/�{��_`5/�C��(I�"(���>7/��_~[�2�@+?���%���J�2!�r���+@ڣ�2Q�[���L�2v�[B�}�a�<�6E��a�mG����[�2�~��2����y�_�ݹ����p�n1�۪���Ƶ��Q��8�Y��&�g��~�*G5C�}h�Wx����)�M�.���Ь���aU�H��Y��U�0���W���d��g�@d��[��Gp?J��s��"]*le�VP?s�7L2u���%6Ot "�v��[j[3O*~e�;G�sKmҊ%�VU�ry�sR�<(v�S\�uC*���~�1�:Iq�,Z������ѻ���;���kW�}����}�T��թ���_Zĉ�${I��~�!7[��Xx�ыD�V����*^_��n����Ʉ�^b�Q7�U����8~M}=+���bL���m�^�㱘 ��c^�UnR30/��@zu�х�6��mU�(�+L�XD�������� � KⲼ��"W��Ib�;���)�U�f��������UT�6Vi׻�b$F���v���l�f�U̾+Z�����0�{�ư9F]W���0�Ԇ�"�JM
�{{��n�%$����$�T4�D�bP��!7�>�>��8=t��ܲ�~�d샔*���ehƳV�d|LH�K�-�xI���m��D�~����i��-���}o���=B6p���,��Q�������9��+�>1����J�7$��M_��k�������!�1c��Hɫ
�����E尘�W��ۈ.�j��J�����ke,�:�c>m�A�c$IT�H�oQ�ag�3�9/�
E$���W�-)�я#�͐C�%�`�7v�b��� �о���=�y�s�o�	���A�HjI�ب@] p��ޠ�F=w@�O��묫����B�2�P��46��=<�l�$F�����&�� ����a4vp�#�9�_/�H#/O݆��`{	�)��e-�=p'��\ב�5�W��*0�9`��=(/�~U�Z�Ǜ�����X�hdsh_�,�W:��}��
�@�{�����`�5�c}�tWo�;=�8��%Aǉ9���búI�� f8�/S{��5��ȸ�����]_��t���U�Ҳʮ)����ހ�� �}����	�P��n���6��xo����p3:@����1�c��_��;
Vބ5�k��Y"mk�ۑW���:�c�q $���*#\��MVs��z���� �������|v��"I�t7���N ��q��AH2(��|�Ve���iZ�|6�s�;ru/jP�C=��|����V��#��P�*,x��5R�#�7UQP�J���ҽ,S+�5�U��L��9�J��hq�]@�X��ӚaiZ�8v�B��c^�׀�b�xBcv��b���үO��is7���o3=�x��/51_�ஷ�����.����o��F  :/�o>�/wI@�p�ic�xZ+�j�4���2���gp�I�cY^ԧ�%�u0aĒ^��M��vӏ/��ufI=��qMʧtKpLf����B��� F���	� ����e�R���!˛m��q�Oq��-�Ey�����3��87�@���Ln|��P�c�(m�r�n1�R84��|*�+q�) ���y
�����&�� 
���EoWUg���!31�rj&�8%$�O�^��p u���C���c�1�Q	;�ԮYPB���9����<gV��&l����PL���Ǫ �!��a�,]	��7�cw������0����!�I�^����\��n I1K;���|V���{�Db��E��$[bV����D�HoC=bʬ��v�=���`5��*>
,|��:H7Pb�h����o�[|�A���\��:DiHxb�z�L1+:��~P�Ӛc����)���5��X�n{k̠���f8��f���h���X�>�i���o#��~+^�㚡�clP��8P���>6*��9? �@o���dO8�攜G��MY�y%��d4I���Ew�yh��Bk8��S[n�St9F� �y�RT�<u�4�w�R�/��u[��+La��d	�hD�mw��¢�D"(�q�r�W����ȕ��/�ػ�s��SF?��\�k;��1qI��3(k�H�齼����u��}B��_W�8�	w1r����ĉBa���/t�@{-54�%�;r���B�^a&��&L�'bA��H���2���NŮ��fp��V;q���&�{G���4�h`(:�/�E[)���A�������ӿ���uP�ݬEEj���nqs�X�)l@c���A�M;dt��cN��[����$ u��p d������5�9J�Q孮�ع1� 6���)�fI�"�:�Qn"}a�����%  �bFfC<ˇ7*����ϔ��{���u;��/ Lg�R���If&�J��3�7�>�U
�Tq���J��k��Ȗ4�-�k-��~SLe�)2
��1Ƣ ��ճQLpG�`M�Mm�=	��v�V uz���x�^Ľg���	h�����V
�Ͼ��1"�P��.@��e}W�.aO֧aC]����#�	������Mjx`n� ����N[0M/%UĎ|,M ���f�us|��܈���m����"��S5���/��{�|%1�&��?����n:2YM���mzX���A�N�I�枊/��*�iv/k��ߏs�)5x�({@K߶K�E������ܭ�%u�r���Q.�Y0%��r�Z��釷��UH'jUVbl�اc�(�ŧ�R�� ��(�H��)I�����Z��(sy�HM�FR%u�Fbb� �sIX:*D��c��b_�765�z��3��a��OL�4;5�]gZ��H��x6�=���&�d��}H"�����D�d�rᓒ��x;O`
��(�I��齽G-�i<V��H�A�G_ۮ����k��r5��)�c�ޮW\��֗���'s��f��S7z����N��ϒ�u0�oj齳[�R0o����)Q��	�B��)�HM.���s�Qg��fu�olL&��0�̃�)CA6���.͊�̫��p_���R����^1�ﯦN�v�#��G*w�V���eG��A$գ:��8��Fb���7yQ�D�O=.P�k%����s3
P�G�p��&n��;�??�R���.�Tb��#�֭����6���u^���[}徰ɥ�&b����d2�Dv�!O�_C�gcgl�JheH��)0��%lH��0#��+���B�.�H_e�[±�f}��@M��w3��£�����O����m���9�}E�'(���C��Ԗm�ǹ'w�KU}��lx{7{f�'ى<p����9Y5�g�V2�XE���az��c�,V-h!�����`}���ʍ�x��7%�;.�C'c｡H<��@2��+l�*����ɂb��д��7���D���gd����^$�d�K��n��]��ǈ���+P��M�o��>��ݜ�,*���T��6:r��79njOZ�mR��(T���r�e?��Jk?D�mL4.�n����4�� ���ҩ��^pݒ�Û��0+�Pʵ��EB�/��֙��\��	�]MQ"Q� ���+�;��P���(Dц2��FI�u�?�/���͑֬O��8��r� ��/>�ZKh
+���i�Qx�~��nH���3�����5֚n̗����aP��f�\���]�J�:����ky��H�k������x`��d��×�b��G��f�X���9�H���T
�������E�P��) �|<s9��I��Թ4�UG�M" �$IC� �g\Y���n�nL����:�5M�Y��B>��E�GM������w�O��LIа"��K��4�����M>��G�X+xd���+\����&X��C��?���bO�z2؈�A�u�.dl����sS���`W2��4���^��iP@�����y�e��Ѡ��p�8��s�H�C�h!�����Rs=(R@::�M�)����BΟ���6�K�;68�6�ߵ�@�\v�L8p�_)����՛S�W�5���`x}
|��Ý�xa�-iҜ���'�K��7]>@*����;d�!^`*k>��ф�b�Q)����W�+�R�'��F��GA_Ds��:q��AyV‸/�#�_��RH�����I�\W��?�L�	w �w�s8�
ٶh�f�����|��^�P35��3��𪂠�ȯ�����Ԫ*�7-��C&c an'�s1�C����,1�A)͎�2y�WQ�{�㟨o^tu��^F��Yd�d�#�X��!�"V���"\�K���~g�̥�����Q ���x�S��gF�9(yXg6\fRjƮ����D>tf��,��3�ʴ>�I�9r�EΛR�3Dk��ʘ	p���h�ݨp��3���}�x _P��L��ڞd��߷'��'��5ޠ�⅍��7|u�g�zG��M��r?#�Lݾ�y�}��AI�ҹ�ILD�x^;aސ����n$O�Ŧe^s`Rdb���?R�r2��6/�I_4���	|Ͱ��B5��*/��c�;e���jP�?Q���]�U��?��f@F�(�
ei����wA⻂
| �V i��ޢ����	�����\�_Qw	�9 ��*1g�ce������4��DfN
ף��{l��.]��[ΔNն[�B���lqi�������@����
��B�����\a=�q�ص��X�۳i��q�K΂n���0VI
iu�G����G:K��&+92� ��9�_����|��=љ�CS�N'�D�F-�Te�;�qÿ�	P��_�縅sL:����!s�w��_ټ/��� �NY*5��qK g�V�;�-��'D�߽"�o`�2�Z��ý�:�I��a���@���������TO?Z>�]�0Y�(����صo�B�K�A��ўW`�'o�ʾ�4��huc]R��hCŗR�p��OmP�4<�r�?��C��I�i�Щ7��(i*v�  v�Ҡ0݀���ǿ����Ud���Z���m+
C�B�[ul�|�F@��_�qx��R�=�IYي;O���W�{��4�n;ϦY٪2�����ʁ�0�?7�B�a�].r-�z��ћ%��O ca5v�\���ܭ������P��Ơ�>�_�)�H"
#Ž�/2��[{��ar��7~&I��s�<�0�51Z3R+n��yp�E*`@�[r G�r}|�Yҹ9ҵ��%�ꮆ��I��*��L�]���xI>Sl�Y�D��A�Di4s���o��:s�]�N�E���Э���Π�Aj�������f)�B�i!��v ����V�L�)����x��O�\7��y6�ST��ǔ�����e+�$�QK|b���/<����ׇ��4ġ�K���g��-�Qp�\.��.��e&�v�1z��*˺��tyA4���J�\H��/�!Q�L��[���!y��23'��L���@���[a�(q��UN�^ 4��;D �p�|�f�*#�j�#��	�����Gb�PZ�1)�K�����peO�,�O0J�(V�Z�Q�#��i	v�FJpl�3�9���?����ǭ�iu�:x��hH�X��v�\����6����(D_"Ry�jmy)"q	�h�4����l� c>�Z=fEiT}���j� AD}���suV�)�/���:�Oa����x�e ���:�a��v|L�z��P,fzcQ�'��_�X_�ep���=��	�l]�ΐr�i��/!c���,��A^��!z��L�<�*��[���-��q�L�4� �=������c���C�d][����1����&�½5���Q�)V���F����c�eW�e��$��0;?Ԃ;����D�N���~�f�O�6������Q��#�F��}7�o}�̮�7��׳o���_�qK�ԓ����X��rcW�nV�;�b1J!I�~W��i&[uz�t�&,��yl�~�dkO�k*W.�KW:]>%9��;��T�ۑ��4�@eY<��l{yP�َ���Oc�|X��?f�U��f�|w���ݽ�_m�M��|�mr�� iI1E��qtV�V�/�ޠ1T�8���k�vk�\�K�n���\m�8�m��`�wE&�����p�K�|��U�2[�|�)���b!6|A|�or�/���g�B�Hr�9e�8�hD�Z����pPm�̷�~Ոn&��,��9d w�B�ȋU��(P8nvK,�f�oi��
�Z]A�Ɋ������.a;%ĈLE,~lD3����Y�M�2�wF��$��B�T�0�K�]�Ss�}�p@Ҧ�����P�z�W��
m&bR�ݤBa�5�D���f���jO�A*P�zї'*�!�ÙV6XYg.�.1c��*��s8c�NP��x��6&BD�̝KQ]	ګ�,�fƝ��L ���b��ę�� w�
�����_�:��h���+����3�'��s�OGV���A_�7�b���6s��w����L�2\OKimz��;I}s��ɀ}�`�� �ߖC?Z��$�..سv�($�[��*���b�V��*�u�S֏V�}���Ɓ��or�_3!��\��� rL��*����F�$'9{�B��u{Y:��u�׊����c��s㫝F麭�
��m�(~�y`�nޏL��$t�չ`SJr�9 �PCމ�D8u
�h��-��L]Id;Xٷ�pr�tH���ʜ+Y������3-`]�Jt�i��w�����4W ��LyΛ1�����_>Pfx�LW���;2�� �"��+���Ǵ�W2��:�Lg<�?��8��ELS���!� ��P�i�	�N7��;�nd���c�$��{RN
�C�ہ�NXd
6��~.Q(��)�B����|7��7!Ӛ��Bq:��ң�)
G����n�F�`��W�AAH�²�����7?�PQ��a��V�8Wׂ��7E<|��w�!�fUtv��s�M�P�e��k�+\�2r�����.��j��Ų����ʟ�����g� �\��Q�#��k�	RUk�i�:����>��|���f� ����ǆb���e�!�c\��u`tR �����|1��ȦQUy	�%[a	�:|�~�V����qp�*+c֕���{�3�N/�d�)ZR&{��ػ�5��]*B�]�I@[|��H�VT������R����L�yMO��8a�0��*��I������ò�U\�� '�t�^8�{Q��݋��b�����@+V�%�M�/ۖO��q��=�uF�R�ËC@.7�Ǿ��^�:~��T���`�P5#�iY���O(tڝ�l^W�^��%Ԩ��a���vw+QG�T�������*,�m�~Vg�mM� ��X +��ݏ*22����~C,nE�w�m����B��u�xv�ه�G��^;r׳2O`�H�#5؄��"�Ь��l��;|�;��-Աg�[W4i�.���弋� s��%�Tm�"g�*%��Bf~�k��>�K}�n�a�:,�<�k�wy�t�uY�U�3����8��Ƅ����-�	�tB@�:ݤSs��6� m<��h����R�4���ĝ=m6v3��!��z��
+� u�`��m�y���2�2�3�w�-��E����Do�3r<#�4b ���+
Ό:�L�]�v�U	�+�`��V�
���I��]����d�2l
�:�!�Ϋ��˹�9���p������,� c�Dpi����⹾�Pձ.fR��CQF=泌V�'_���6�LW�[�{&pl�;~'5�v�#D�T�L5Z4ԅ麒'�L��LԤ������$f�p��}s�7V�F֚�	��]�>C��(^����C�-�j A�l�G�#�hV��"�2��e�`�xk�����fs��_�к29�g���2�	�K�����&��u)!h̖������V{C���n T@D���I�{ʉ�1����%��ݭ$.j �Ӑ����xU%n�եa���8�%j#�����.���"<���*5����!�B"؄�B���a1 @14n�-����gBy����]Dg6�2F";�@����tHҚ�Ѝ!��B��:�f}���FYY�c1���}�u>���#D��I�'�g��u�f�9cԕdn�f�Hخ~�Dß=l��#������/�����-��5�Al�d��ݟ�ti�&��l��OO/�ӗO���aܾ�`T�!b�t󂬋BG��ؠҎ�/�׸����^rҐbQ�#\�����R_��|ؤ�ϋ�V�����O}�p�)�/�a���� 2��g���) ���t5Sx�ݺq'�(J�JB�=V���'�L�y�НĒ�Nm��0%��v$Ḃ�[�4o\vB}��By��7$�F�_2�@��9��]�1�(��e�ҷ�����R`�qz���*�;jPCI�͇b�+��-Sլ$V��b��s�f�-hy��:I�"rl"�Z�h0�K۱"O���Ӝb>B,;�MS�dI��z�[oZJ�c/0+�w�l.�+� �0>-8P�U6V��l
[����6�[HV�Ub�	���2A��}����Q��S�̦N!�p�(_܎3���O~��}��3}�c�?��B�F�Pq��G<�#���q,��+�}��T��_G����(�\w������D�C������U_ �ͫ�l�n�~��L(,w�b$�}���*���L�h�����B'�LEE���E̶п��Sʌ��^�!C��IO1�i��ȼGI�2�C|E[�ɒ����78'"#�����Cd$ �2x���@�jl�#��w�{
�舾Bl_<�iI萐�S<Oo�Lb�������%���E�_��Z��@t�:�4 N����$ ��e�$B��wc����/~��xe�`.�x-sQ�&���1� �յVWZ�-��N�MR��;[?]�Czxl>!��������YX��h	^��"	ޡ�`Xk���7̓���p�8����J��=(�q�:m	g|�S y�h��K���T���c��br��p���uƴ/l�R���vo����0�!��֬-���qb�L����I�� 
�M7%*�?}��ktl�F�1�B��Q��k�D���1x�	7�
����~��s>Ӏ�w�d&�I�ɭ�d�G�}�&c{���ҩ1Qs�?5�uFZ�G�*�jk^�;�=j���ђɵey���1å DPYc�4�r�ySAAa�i���������Xl�]���dNpL��2����$�9b��xSŠ�_�<��N�� YF\M�=�Q�A�h��&	��Q�H[�#k����iU#��֊�K�πOO�,�)��ޭ�!�6&��'&�?�P���9��mUm�B
�rZ�i3���FU�!����9u��Y,^w�[},�(�o��K�O�[ڃ&2�0��4v]8����5� ��)��u}�J{v�l��a*�����~��V��
}3�7L�4P�y�a���@��ׇ[$�b���Z;0�~�������4'�̯�Z�"����K�MH�� ���/3�Y����"�u�龨��ќV��o]�Qؿ���U�e��[�'.�i�=�ʣ��o)�]��;����q4A�BR\���e#b�=6�8�b����|*wB��e�]p��Dg���n��C��;�.�Q�)e�#`��I��������Ѕ�ٮ�T�C��'�T���6�@݁��359O+��1DР�x��y�� �L��UjF�В�>�n������%�-�X�5O�dZ�\�P"T����/�1¶�r�Ń��no���a����ǂf�;�_,8�������v��6�خ  L�"�$BHӏ&�W�/-�d�X`���y+cH����NT�W�S*e��=��&H����G�F��)�����W��ٚ/�R�խ������^L���p��9��@<r�1`�Sr�w&�P#� �<��zr��h@� _�l�o�/�����=y���5��"���)j�#��o�ι�ͭ�I�XZJtHrZ��\�6e���?`�J[���ҳ�>Vi�[�E�/�e��%�̼S����6��^��,���KY����ۺ�B99�Y�	mL�B=�-�����R%7�R��[�g����0$���;ETZ���6�\X�
~���[������Lk��1qD��@����{E�~̂�/���J�r�`��fU���9GmD�W
<���2�K��b��A[��A�E^��z����l� �Cq=�<�Y��gPR�Ҹ�:QRx0W����ؾ��E�kgû�n2�c��D斯��.ƀ-*�]I����)鎶�
c��3`��2�����8rv �D�Đ��"ۡ)rJ%�ى�s_4D6.��^��AډT�/�K�#V��Ȇ�ـ=�Y|��$�m.�Q"tp�IixH��k'tL;n�m]_���m�E�&��ؔ�|���֟��75���C��Ђqgd����_z����e� ���XT0����ay��ǟ)@��QI�	oQ�iG͟���?8�q#����<��3B�ۦI`�{ޅ3,�[���T�W}=}��^d��|�p�΋��'ۊ���6�	�,�;v���@�;�b^������_����f'nY�Em��C>��3���Bcϼ�������w���C7�o(�/����T`m�r�[�E��q|��bT�����_����o�:��M����8&�v1Sv�]S����yO"ɶ1�-�Tv�ށ��O'd����ܓ�1ZC7D��#�ժm��C3����y�l�����6�y�W<�GƐx&��Ɣ&����e�렐&�S�����]�K(}*?�#3�]O������e�HT8��x[��&%�g���d�Ьα����/D�;�g9�"��B�������k�7�N���,"�y������e�Kd�q�ͅS)���KR�GM5��ʯ�24 %�ր}��	o@Zl��0&�Ia���<���rw������R���MU�1�����m[c�U���e۩Md��]��?��8��0�{3�ցP�D}S�ˠ\�52XU��%^�^�U�7³�X��_ֳ��x&k�e
�(����!�;Zշ,ٜ�C�e��h��c�n���0(�.OM������?�׃ؿM��>K��<]�r�㮊!1�Ta?�*51}'骑�wA\�7ZT���|��-�h֜�E��e�!D��_�����n�&�gX�Lz���1O�1V<.3������ˬAA�],d��BLY�8=폠X���q��^��!�-	 �V�p���1�}m���� ��lrb:(�נS7Ҟ�w�w�0Q�{�GL�`�~���d�5'��v�#�����@ۜ�����e�H3�l�a ����:�D�����2m����#�|:��8��)�<���{(�R�ٓ[(���bʹc��C���z	nwE��Zӷ���}�����*x�æy�����z��gW���T0d�~�Ha�D��LJ��s}�7�k��}yO����F�mU��[/��?��h=,GEʊ��3	}Oe�)��aJ�e�c`�y�2%��M��xzV)�@�ޚ�'��"W �P�&s�f������:eEux�Šv�#M"�p)w�
�ߎ�!�Bx�S���Z,7C ���9��������|Q�X��B99Tw��{�����}�U�ς�;�� �ZBNR���
Q�G���U��\�<D+n�R}�n��	�Z�*����㞱�\0��m�"l׾�{�]������Kt�G�#|k
�b��Y�ல� ��i��_�\�\�{�Kp�N�V��-o�������8�|Ŗ�
(�]
HV�(���鰈HȐB�D�J՛�)cs�}�P�h��NX0�vY�8�bG�C
���a3�.��7s��ࢵ0l��Ձ$A l(T�]K�:��:���.gz�׃lg�Y�g��o5�Y��х��S$*��k���oA��Y��������v��p��/�n��f�Ű�`�>`2O���@$�t{�y22D��k�nbY��VU�N�	`��M��яߟ:h�0
�31%��?n&w�1�WݩW���|U$���(��}�9�"�T�<�'�u�5Ǳ��zQW����ֿד!R2�6�3��d��8x�~>�ฐ�p��	mΚ�hܧu�V��NJ�X~��b`[<��;��3»���Ё��)��SҤJs/�5 �,DmEcjIdS��%�ژ����0�H����	c�F����[M�n�6�/��Q�^��b�q&%������ʜ��7�YZ��K�Dé�<g�E���cߚ<!Tha>�QH�e�[C�~�NP�AT#����Յ8U���������tE}��D�bA/5�
��Z��K�
�v���R�df.�2��>��w.�`ܘ~	�W�$��gO�_6k�C������}w��������*�Aq�p�ʙ�2�ls��Y�zI�S�����c�-S��z���u���Y�� ����ؑ����治�q��\�K������=y?��}����3ј������ɖ�8�A�E�&Z���2?�Ӿ�����/�4m]�[e��\[.�1���Z��#��4��U#_��BEL����~].�!�G�:5�(��H���B�hڬHfxc�W��\M� ����z�	��U9X[\��A�h?נJ����v���tg6Y���8��� J��-���7��{�y���G������C%\3ά-y>;���0�P���~�|�8hʏ�?�.Su���m�bۆ%��L�v�M2���x�Wq�I�-(ew�q�~<�'#�1D�W�H�������)f��,�w�:.��S�)�g��9�2Uͷ������`3���ȅ��a��R��>�6�i�0�f�Ee���Z�3OT*������{�k:�(n+�RTAԘ�����\-��3���^�z!�rט#a��fg�I�aD����0A�_[D^���C2b3R��ad��jd����F�z��q�c��z�Gy�#y�d�U#7nj�l�w��UM[�L�ԅl���c�� �Uۆ�)�rE9C�7�`3�|2L���?�l�ڐ���״(���C�րn����!���,TӒְ���� Oe*4]:����lg��]��,Ea�I21�8���up9F���a:,Y�8���}<y�R����3��U�ӆ�W�L�˛��^g�����6���bb����Hv��\���C�0�Ғ�A�`�J������mo?��v+Fu�fD3�i��8�f�NV��o�>�����kP�������`x=���$�I��~:-Q����Z���'�.�)E�?���5{��;��eo��λ�(_�0�����rJ��0�;~�r'^��EM�C���9��6�պ��#$7��+x�̞b�t��`��f���ܻ>%��r&�t1-���L���4�� �:Z�[�6��r��ue�|�n���b�ؓ�x��Tڷ�z���b�k��3�)��>j�< #�^hoj�9����:5��}�Di| ��v�^D�$8A0OW��h)e\����u�W���Q�NؙrG���g��ȆE�=A{� �	�*���KPUz����D80���8���<�C25�sy�ˋ^����c�T�ð��ݤ��B�`�p�D�i�2�4�)�����az��[T�@��Т�j!�#J2c�𗉒12��|�����l��u�6�1��D��b���-�2ݟB[�U���Yj	:J�c��)��`IB�z�֋��4��AM��jM���i�!vkR!�|���8G�*&~mT5��� ��}g[�.�Ї�!�8���q�E�F��nm������l��?���>�q�-<��]�x�6B&��j_ i��N�c޴�0�H�4+%"�����Ct[�2I�-z�#���U�ۊ�yA��=sR��L�6H2���2���w�Ӏ��//ls׾Ӓ�cj{<DC:��������Lj?Nuz��o�h9��<5e��(8�g���������N`�6���&�2�C*�ݑ���n8�uZ�[�Q���nJ�$����n�Y�V��ݴn��:l	���w�VW\ͮ�]�"��p�e���!l������+A	���2����q	#Y��/��gT�6.�󣢟��7(�:�����|S��4_lBSH�ّ��sv�ي��}Y��:5� H���/7���e��	EF����E d��P��.�N�E4G�a�2f��v;��/��Ό����#��;4;���b�އ8U���ڨ�6�!��!_�_���ĺ�������hgχ�_TA7��/_����R7�9K�@�
��Ⱦ���M�uo�0�b���i���<��q1�S����O��k�Ŧ4�,�^z*V��@���x�,n�� Ίݮ����;qf��u�G]������#V�k��(�t��a��Bg�[�d19���۹����3���vb��t�g��=�Nt���k>�ț��&�'C^��&R�C2L93�#�_TS��dMϺ9�"��\�@Õ�'��L\��-�E/�r}��,�q���.*�~����!��o׈ȿ� ��r\+c��|��DE�#d<-Dk�7R'\��9Ip6���j4����ݴ������!%��m��7�ea��9!�$j��H��^���)Z��Zz��>lP ���屷R{��6f�a�]�U*��/l�m+A��>��Ѹd��Ã0'|�^՘"�Z7U�����$�����
ئK�Pe��r��Yn��飉!o!%C�5�ݷ"o�CN�x��X���-=Qm��	MrRR��M�g�,���t9U�/���4�|�h{��T@����5�0�i���]�)�L1D9�[�����Q�A�Y=�:qԮ�rYJc{M!;�ᤸ�Vl<. I�1�u�U�e٭�`�S/����3<�m�hۓ�Ra����N'A��C7k�R?z[K:'�
s�����(N(SQ�����#ms.��^�q^�r~�T��0p�^3����*rL�f;	�����J����kk]�A���w&�.B�Y3S�CC%��H��dkr{���ǣwDq�����1d�_�ѾB6W�/#�e�a`ٱV�?賥��F���B�z{��{ۋPB�
���#i`+-w���I��{:�v4"�N�6��)�~����(�_�$��%�j�����MK����!>�z̖L#:����|v�����\�#e���>��e�/0�e.�%'H�fs�ڡ�ka7�F�n�2�ۭѱ�n�#QN��r��5z=@j*��c�{�C�q�\;�؋��m���V�* ;�8Iq�uz'2%��д��+�NB�C���@�O�0Lr
5�I�ӽ�"P��9����������?BE�Ч����vC,c��y�#v�[�N�����V�!�Ä�֋�SeȂhv��ˍ��I�H"C ו�~� ~�d��H���.ү�G�<=S os� +{�x��aO�6z�j.8�I��j�q�oxc��ˈ]�6�yc;)7C�4<��mD�dn��K �;#�H�^*�	N��p˔|� �ER�3��Ș��B���a�����hFY�Hz����Uͯ*��>��.˂rT�*�T4����#���i �y -�QA6� q�VZoX�M9�%J�#��pQt�q�[�IՇ��|�ٻJ�W�6"M6�,�01�rHܰA��o�E��Vl��Lᆴ�S�����P�)BW_�!�������x��~t�+"�=g2�<���r�N��e.{�&nZ�B����g�S�R��`rRj�A��(2b� ^�~Sp�vk��**"�aku|K����YW�Kw�5����Ht�q�b{�і�����(����d��8�B�%��l}�����4�Bs�G's
Z��m<?�|�$���; �r��_�M�OG����Ja�?d���JC�x=�Q��]0`6�Zj.+Dt��r׷ l@nDB�����LH�ID��n]v�#��2QR:��J�Zoc:.2���Q6Z�9�Ct�Y���Ԝ�Y�����"���aPW)^��U����Z���OQ����:gv���Dmh�O�S��%��H�A(2-Iތ�*��Kq����{צ��:d"��i#�>+�-�$������ӑ����B19I�F��]tC��L�:��T��O�����NWU�ç��_��Bw�Z5t;.�ؿ�|��ɲ5G��t5N���?�
�#{�u��k���&�c��41�Ğŗ+3&*|��̻��a���Doˮ���PE|�J�1���8?y�÷_e���}y�_�.ِq7���t�L���j�bQ_O^,VMrم�����9���ΰ�	{�����ݻx�F~"^z'�v�=�#��TO��^?��Hi	j�iu�Jd�weK��%�2��@��/�Z�ͼСk>�S��9Ww�W��	Z�W�:�9�2�R`�B6�������D�SX��:�? �K-E2�"z�Q�?��
��T�
0���8��m�u�t�x2��ߙ���D�k�rs)��& B%<�ǽ���.[�B�.<M�g�SxS|[����k��,]���%���t%L�$4�e®jy�Pp�q��T���\=5����f6�{��*�W���$&�S2YGy~8�3_'):'��P��mn̼hMg�s�������]�W��|�8|�0��/L0.й/)�6���W6���2�����?�@�(���2�n��;�E��v�>Q/�����U6Z���ْ���ƪpV�{3�2�4����u��!o����
m*_�h��-�� S����,�M<��H�t�{�3l��f�Ox����'�k�U_j�uރ�ك�v�9.�[��I;b\��q�`�5&Y}�oL�����9�I�4�r� ���Vc��"y�w$.����������f�Id���"�6��>��wB�bP6x��L��+��q�鯖 ��InXvpWt��;ItL�m�,4�jЋ�+�bX!9�v,՗ ��Z�D��箔¾*殑���+��g�a]�-�+Y��Ole<�+G��&bH��ʊ
�]~Ar}�˰�נ��Hz�n��ye�H�f(�qq��{���k��4��Qj_ 鉡RW}�h�?���"�g���;���J����*BB�,mňԥ_�q��<	���/����+T����T8"?�(b�QEɻM��*yh]���o�����xwȚ5b�)8ȉ�0iW+��-�E�z��������愈X�\��	�E�lψaT�ze��B�<�Ƣ���Ь���@�{��D,��nj�S�\C�<���Xu
�O��,�Dyg~���5�]�4u�������~N���_u�a/$���3��|p�Q���4�.��LL�+EɠS��˩C�i���
XV�|�j�KX�`��`9U���g|.Ŀ	��D�`�}7��&�J5��r d�����1�g��2�сr>u6:���E��Tr�>Y#��9�s�P8+�4s�{�mT�Uݐy��Ӭly�?���`o���𳹅�w��iw9$S��If�̃��$1y?��D��<����t+�t�j�H\\��YT����h+�YF���=�{0�^�*�>3�J�"#�j*�3�A�q�
��R(w�hdV�y

��+�	��
uk�+�[0��%�V�",9il�������5�\_�������'Yl#�~Iܞ���T��Iy����`�F�m,�, �8�Mb�^��lX?�U_�@!��� �Ꜻٶ��fIRڴ�жg��wbR3�P58���0��i7��)Ѽ<��l�G*WUCS�}��% ��k��M]ѱ�>��������\�5@
;H| �[����6U(t����'	�wV݃�eT�	��5�|e����`�Ww)rJ���"+���~�[��%On���c��R�oC��]'fF�Q��1xG��me^k�i��;S
~���-��I ��6_ z�x�xFӶ�v=��������������fܥ�ptq�/�����܈^������\V�6���Ȓ���T[`<�]�/`���}6��� #�\�{�� K�s��Z��keJ%F:��ɳ���vTؐ^�>�D^���ԇ�r���H��$���j+x8�@�r1��	z��8Mox�)#)��-�zrsA��jL������dw��ry�DWI��' L�r?6p�v5�b?T���r�<�W��n
��Pb����	)�ȑU}AC�C�/�����ĵ��~n�>#�PTe���^�ƨ�SP��s�Fn�:I3���9�� ��2��x�v��Ju��#k�TM��"{��&;t$�(���	�S�uqMY$�<^Bݜ#���5D�ⶺ<��>�[�"�����ඏ�t�;������.���-arg���oo�E�&���+�( ��c�̻��@�0?m��&���"�Y>�
����_2�6�W��S/wj⮵I��õ���F�f�7٥�#��:�y���˲(�2jI��D��ȦR��fƨEX�f�=�����{ה����� No~~���!�Ry0�ӶΥ)������LـW���\��Ǹ�A��̌I%6�W���	����%�{ �U=����jr�s#���gO;*O%�JQ�{�7q�#� r$�݈�x(5��t�t� ��j������U�*��z�h��i�)?�P�1����6Z�{��b0�]�����$��a4�q�Q���G�_�U��z�dB�9��B�_�ljw���5È� � v\C��P{n�Jr���� �z��k�[����U��9���Sx������9}���°W~�A]��M{vr�!���C���[�Ò���&��T{|�������h���qlC�f`��t�\��u��tlt���O���=3+`�T�?j+���j�����5Bl����=N��������x�ԧ!��v+0Z����}�j71��ө�VU�8�␈��/&^�_]����J�º>��7�bǅo'MҕlE*�I�p�7�q65պQ0��˸O�)�E1��k_Gmʲ��Mc���
����L�$�x0�]w_���7�GC񀷆�Ky�L� O��}��[Oh
���!$�sa�y�I�ˢ/x���u�$lޠ�m-AL�SS'�æ��!r*R+�����y���TIA��zw�Z&N ��U�19���fm>��@���OZ�gb�5u��&3��a{=K�+��jf��S
�:���y��>Z�A�w���*P�	=Ưu��O@(����;��+�وo��S�dO	��!# �r��۫Kb:�!O����Ӟ�B؍�	���5��	f�:$�r:Y����1�f[�9���j�z�J�� ��th�x����?s��Ds����G����?��(�D�̰�Z��٦��������'�\r���?_W���|���E��$���Ǡ�5F��f�±�+�^7�� :�dz��{���Ja�8,�ۚi�k�4ifׅ.s�?"�Ľyl5+�Zη�G+�FM����*kF��ۼ&��(s���qM�U-*�2�>O�<��`73z�� h\�Y�aZ��)$��k\�<��6�6�8�����5P��`�SѦ�S����dI|C�_�J�hu�&�@ˎ��g���Spg��AF���z����`�S
���$���9Df�������`x�I@nhk���C�7}�D��9mR-q»��'�� �ƽ���+��Wh,�,���)Xm
S�H�j�3�lg��A"?�~S[�*
��fqk8�-=�:S��OٍS�� _�?/Y�"��_��o{�`��!k�%�u}_�X|�`�؂GU�ɻkn�C�o����r�^������vI��YqG"�\/?+`M�Ӫp�p�x;ɖ����
�cI��+��zߑ��\6�m^�HG��t�����钰�ꛖ{�s[�}I��B1��e�keau{+�*pb�M��Pw�*=�?����������)�3p�m��uH)�30^�U!��_Ww�f�>�d�4��1J�EY�3T_�����6)��y������8�Z����_�����+��2l��(`��Ix.rxrpE����j*����[�ñ�E漻�/ǭ�4@G�P�N�s���d1E	v�'/-��Iv�a��e�EԠv��ix�X�n���;%�/,�_H#��N*�M��W`ݥ���$�퍰Fԁw�s*6t�uχ�TTp��Oy�feK@%e��u��FRP��Z=�#]mb�8�2(48��j�u=6/i�D��	�����0�-$�W�ß
5��ٓD�Ͻ�T�v���3��~t���x�cV�][t�ba"j������^�I���G�W<�M���� AH��P����}eB�bz��s 3��ü�|_<.�$��Oz)aD7��Cζ���(f(����g�����,x�D�V}N|��Q�G�?��h�H�>x�+Ή�v��(fi�ʮ[�qr�*h��p`,V��1p��˂��p(HT���<�1��s��nݙд@�m��R��{@��%FM���/��G}m�jG�´�?���ۮ>TG�Q��Ԁ*I#�H�F�NB-5;Au��nӄ��"��|�!����]T�(���F:s�o�,��<��GY3��*��M�D*�V�{ ���A���Ny/�$P;�pP_W�����mŹ��Ĕ��6l�V|o���ŚE�j	N�X&�z��������.�fy�2f�c���<�j�׺U рC��_�+�k�_ޏ�@�ya�E�r��F*T�G�b�V�rZ_}��R�?�%��1V״���3�w0�x�b-�Wֽ�W���nU�4i\Ɋ�~{ރE�PH״�P����Қ��un��ZY��=+	z���4��@�w��wQ�t�����g�^�=�^�k�{nC��gW# ��mEW|���w�`�mZ|��0�B�e��
7 �eD�>����(����t�{;��,�~�h�6m�M�/^� %�^G�=ƶ��y7��.�C��`Ab���ϔ[��}�y�'1�bu�7�{\xܹx���
O�h�/�|�q�6Y]�h��ʖ��y�Z�y4����.*��Sf���!fE�ܫУ���-�����U���`y���Hy6=۰�k_�z��L�Úޒb�߰~9n_�� ��@�T�d���x�lr�k|EἤA6��h=�*gSC��pD2i�UM�a�f��5!�*����ұt+�S��� l�h|q�|8-n�0YͶ�oNSE��I��3LUʹԆ�
K|�0~`���񉉦�0�뗜��/�p���=#��<��Ӏ|�HtP�����,�R�?ч�GB�-�{���n�y$@���J�x�L���ݻ=�Y%DTn��D-3��[�v~�끒\J���U�2�&����<���̒+Ր��C�c>�C}/�v�-M����z��O%+���M4�B�^MB�rQ�V>������ ���D���72n�=�G���ĖO����.b0�1�^�;�t����	���T�S��a��B�tc���������՞ܥE,$�K���hh��������EE���lm1|�I�P����s"�v�w��{وc���i,Cy� }n��T��P���0h����zagsW��Rǿ"�������!~������'���PȔ]���{B�l���,δbg��:Q7�E��XN�Q�v�/o^��G�4�]v�Sc#��.�������E�2f�92�[7����
]��Am��@��"vG3i�i[�b�}+$<�ף�`[�Ep���-j��w��X�Y�5��������[�H�l����|a��t�����X��0xy����g����|��W0��.�?|X&6�l�N<'/�/��Dh-����=�����$�a����U���)o��]��o��M�9�kӬiQ�^�^+�*3� >1`�k��elz�T�h��ͥ�\w&0��p`NЊ�$���A��^���:�p68r	��2l�yѵ^þj7���aF�~?��_%�A�,9��� a_gZ�������J���2J	Bf>�:��F���ь�����]g�_����V�wߐG��t�
9�o���T���@.#����vU� f5&q>p�d%�Z߉�L&΋��A܈�Ζ<�Ȟ���+Fx0s�(���nO�3Y���cz�^�ӌ����{�W���"���nA�@���7{:}��]����6�g�д���{�&�	�Ə9xu��ْG��Ν��*ۀ(�dv�~�y�uuV�C���=NB>����;�1Zy�q[ܬ@�Z��k|\��`�oL�.�w� ��{�Q�r�Y�B��5�u���M�׬�S����*�P��9�����q8�	�����	���6w�\⼝g������uj��R�����]ǀ�K���J5.�(�����D� |E/4d�]g�r�C�,�O�>�I"�XW�����>��<�~�]wvw��uzՠ���́H�`f\��o�7ђj�ZeX6�F[��f3�~w��ΩzO{��ʞ}������I���3:xe r﷗���Mn�q޿����E��J�C��Y��\ȹ�s��/h��[w_9�Y����Q��燃��oOy�����4�s�� ��GJb���^�ȹ-b�:���6�4�SJ���=g��2�a~��^��%�֭\�e$��V���OX��n��٘�>r�c˭����v��J�$C��}]_<�!��f,s�L�f�g3I�����p���:�jz���3�ܼ�L�����)�U�;J.T���e�s'K�@d��;�D��(�N(�hj0�I�<�?���#rmUuuEA����=砹D����	*&�#�Q��Uci�f2�(��*�6�a��R'��%��sl��2���3^��ؠ�OCY��R]�_�֪��:Tn�- P� 6�b����ź���
��7�Ȯ��2F �L�'D+�6��.���D��V��t44�������3���U`�x�J.GYەֲ�vA�ՅD��=��È!���ڄ���m���������LB�7�g	���Pk��I��+:��-�i\v�f=�����c�ύv Q�*���Py"�2�_h9�mo�Uܚ�~��5g�0*�A6V�w���u���䉘qB�]�Y3��j *�Wy�L@4I�uG^+����&�	hWΙ��-�P�G��}�^���ߥ�������'�� ��}<�m�
�)�s�i�-\��i��I繛R����q���U������_�d����]�|6��L�Vfʓ3�5[2@�4�OO���"=ܸ7W(xB�A�M�L:�M",�M�%�Iy��@D�s~(_>-�P@��<�P�%&��H�h�i�y�x�ɮ����+m��V�JxU�]��,���▗�]G�4��~�5X[�Ik)|�����k�h��f
^��y���(�ŉ���ͿxENߝ�}�pf��^8t�G���<�AA0������-
x9��.s���&Z�b�H�f�f�W������í;�b�[���3K��4]XXt�!��mD�L#�1"��Q~�>���xP\�5֝��5םψAL�4�+�k����H4��3'G�"n����~5w�SۛZ;�[��x�}�����$�s���!�I�|RO��M- ��V�x.�m^�W2���A���l���B�na�ޏ�:��Ҿ�+����o��6+�(�qW�${]tw�����2���'�obFhv<���M*#E��s��8������XOjQ
]�D�[��"�:כ�h�brӻC��0d-��v��RS�\���d~��p��p��#���_(�"`�7�-D�����ĩ��a����_䫒�O�`Iٮ�-���- 뻏_@U�|�gr�����-�	*OP��L�b �s*�-m���^�.���8&�JaZ0�Ꭼ��\%VM�-�ڇH�=��[��G")�rJ�6f���x+�*`�Ң�	��L�����i0�`����ק��:6�@̩�4�4~�U�q5�Y19�m�1�k��i�Wc��>Z/>)�t3 ��l����D�$Bv�ΔR�s@��w���:tY)�r���χ	�P���-�	�eF!@�ղߋF;���fW|�F�	c��.1�w��Ʉ�~:	V��Q��Q�������[�*������%^�����Ȯu�b6ݗJ���V�L�lS���d7��0t�<tc�am���:R�kA(ϒ�hUD)�B���8�KTR������f�h����m�^W:�#��h�:y7�wΝ>[(P�����)8����|��%�[�z�|
�!��`Y�������4��[���C~$Y��c����z���-�o8�Ĳ�21����v.+s�?�����I*m���z�p�(�)�\�6:�tr��6gH��ŏ���w�.����][S2��R����3,C�T��J�(�Jio(P8U=T]�n�TX��XH�%��&wu�qYxFV0�psĩ.#�yG�l�8 �	FN����x*?D�����D�*���Im��@PS.���GjN�F,��t�#�8�z�*����X��9�3^�X�)u� x������f�򀭾WdR�J,{����4���!�:|ZU�^�������V�v}�J�9��UeA��L��5��������6�\B��d�Um���,
P��'�5g��T�=�O���N�g��O(QF�3"�"���-p�,Q�9�~�,�dx�"��� o{�l�Wn���Ȉ��
�?~]�P�U~g�G�J�u�r�^	�J}w&MK|=ȷ!����h�g���[� ���30����g�u��:��_�i�d�`�y��7�~N�ft6u82��N��B@�kO�Q�<msg���Ze�Y���	c�,��$��
���7)q�1��E�Ѿ~���k��a\��3�~|��Ș��Py+�+�*��&�=��C�L��Cg�5�2g֔���e��̑�h5/�:������1_��iWbiҳY}c��E$v���Sͫ��QIwI�ɟI��`�֑���ƽ�<����嗔T��ρl�.'V>�l��ߤ q�-5�G�bo�cpkw[3���d'���\�he��t�BS�>�0�Q��Ϥ4wܙ@�}gfs����)j��MDq1���`Z�3�f�dM�ԛ����Ӊ  ��r�o�+�1���ro������ʮ�}��w$��.�< }��Qw��:#�T���dΪ��dvl�5b3A�^��Zi�r�UM�\����)�8e��'���z�X��P�pP2��#Ж#���U�;E1�Aכ��-�{d����0V���.� �D�po])�V����Q �wȌ���5�>�[,Y�}g}�$��Q@O$V	6K�� W7+��W�7m��aY��t ���eN��F�oM�9����,eH���J����9U��b2�󍬒Qw�=��qM��ɀt��	�)�f��i,?~�3��X7��@��3�w��ŭ���k��e�y��WGH���	��x�T-PpK{k���G{H�ʅ�+ص#�X�AfjM�\X^�n_�P�$G�㡨��K n������g�y
(��x/V��%����E�B�I�ɟt�s�ׂ�9����BVX+�[�4/LE�%�����5��Ƞ��X�>������Vt)��G��~��~T�>��	�<�*�;fe����Wq��0�q���1��&�҃����P,u��XL�³���x�lZB�8J�/�+��wkC��\m��a�f������Uh}QY��7��(6�P�6�1
��7 ;��0�!��NM�&�w-X�-�s(����U�<K�&tQ��ڑ%QN2޺�ə߅�A��SP"�#��t_b�&�`�_���*�>��S�.��A�k?���7�#p+A���4�$�}�߄Y�I'W8Xq��,�*�9o'A�Cg�	y��Ѡ���C���
�h¡#��`X����]h {�:yb����4�	�����z��w�E#�>�4��D���T��>[�$��.  �Lp����z�4�&b�?��\h�qe��Q�2�����Kq�����C�Լ.����f��|��h��ym��7j�#��:�z)"5]���/��jҸ�$��n�:h^!ۇ��]7|�d7qhLM�ݔv�Ї/�#��i ��W�E����C���yW��i$ox��%Cnjw��Z�5�XÕĪ�莳rbk�(�#b�����^~�߿BD�H	��,z���)d�H�vZ�#k��q]A4�g�R�$�����>�Һz �`H��ZL;�b��S�g�Z�J��Ã3x\�u����C4����52wu��j*%�1��c�'���ӏ+kr�Ww�4�*Ă��e���%&�T�t+{�\�C�����VL�t�SV��*����{$g�=�ù7���$�0N�b���I���O�����x)��=_3����GN~:\i7�$�8"�%;���d��.�@�D�T	u�BL'�0����(��#r��2�˄�3�i�i�6�9'�a��ָ��E�vG�MX�A���Io�h�1o���!��P��~�]��j�T�ۖ��O�)ܶ8f�c#��>�� ㌭�6k΄~�k$��Hr��(�}�`���?�:�w�{R�\<����Z^b߫�������B<�>?�ru��S��VȜ�?�.�S�v���l�a����Չ�k���(�*+�X��g��r [osC\�T�}>X��N��Ĩ�Ҿށ]xx��.�������`\�2��R����f��}\�܊d�!a��n:x�4˭��i����^�0J�]�'�J��n� �'X?w49�{ W�u�Q�.�)7��D��D�M��)�E�/�x?S��X+����s�D?�X�C2.��A���@j�h2�y: !UE}�&:����<��,���f1����^!�2� �ƣRև�l���+B�cGs'��b�*g���"�:��:�d=d�*�mvN��׶R/Uf�������P�8א�#����^�G;Q�= �@W��� >�߈`�d�nz�S�@7)#�:����Z�����yu4٢n�ppq��$A1e��o��{�d�"(%��)ˡ}*���ST�W��9�b��9��3FG��|�����AC�F0׺�c�ݷ	5�NM�Zg��q}P���
�u�1�2�!��1젉����{��>���3P�K�{����0��i��x�=��@��c�l(�87��|Y��S�$1�<�G2�m���'o��d��ۇ��,S�9|�b��j��`=��-3L�S�<�AC�@�b��|�$�vr����`#Cs���~c�	B1WY��z��_M�M�K�hX_ɓ���}>w��3K�q�
Zj��ҡ��^����bi5��F�I)����1lJ١�Fԥ&В̣_��@#�;�z�Y@�!߾	�9�A�j꤀X��>���F�<�O<������9ƺ�OW�<Cϭ�p�U�J�>'�.�ynj��o��ű�4 x��U<F��}1X��lh>�N���z�A���a���/6=t�}7��S����⧃���$��'�:�p��+�0��!9���,�k���_`�)z��	���3HOI��!$�~PYJ�ݬD]�,D���T�F�h�v��nF]_O��%����ݣǏurp#�x����{�Z�l��P���VҞ��x_�If����օw��kDS�AB�s?|s4�͒�b�l@���j7��Wf��an���"��CQ�SA:D�a���k�d�
w�VF4R3^�d�<Z~1�`��&�)A����yӹ�a.�!{q�qj��?��~�b+��;j����ޫ��v8�������6����.H��N�*G8��,�muu?2B��Mnm$�;���I����� -�x1�s��L���X�T?�e��J���ZC�fW���Wp�m����h��M���ݪ�UbiQ��]y���������+c�qx�Oտ�����(a�=�&kS=DnP�p�k��/|�v�|�q�û)pe-|B� Z�+��z�1�kݚ�8l���c�.^�� ٱK�5�������a�?��_�&&29�zs#�S�Ϻ����g4�5	=w���12�gU��5K�v]F\'@�@���$̀|OG�0�T�"?�H���bV����,~�d`���b,����2 �k`�$-��g�<K�HHb�	�Pi���r4��o�x�﫡�8qy�7���Ky&b��e���- b�5)�H�|Q7Rt%\E��ߴE��\�~�|^��n��V9��X+P�D@L�������J_M�O̓T���y  �k�� �#.{Xev�� �)���ٙ�;lB�2EQ����{�yEq���2���Mh�>���!��iՈfť�f��'�r8�wR?��=�m����;TA7y���h�����<#j�5�q5��2P�)��|td��X���#(љ���S7��.U��&6�Q��@�ψL�-:$Vɻ	�B�RzLf�r#�is �9��-�Vr8O^��"�9x>�V8tA_��2�\��<]��b���=n塉�儕`Ɍ]bML�m8m��YC�:8�2|<�+J��y������D!{��S���G��I��|0�%���S�ysz�[`y�D������6����o%����6�7nWWj�sͼ����qd×G�9~-�'��ᢦ�U�`&��;�\ 'hX����s�@6�.�^@	�Î��~Y��
�U��}�HSO��\sb��d> 嶮-ݴ4p����	��d4�E!/�9#��5��f��p�QF���rdە����8�)��yqҡ"��1L�kYt������*o�-�b0� 7��� z~��C�oG$TK��}gQ_���}�V.��32��e�������l� �JJ��}��OR��Nix�Vg��m�y�y���G���m�Q� �g焆
ңlUn�q�`���|j�p5�w��e�P�k��Iq��52���0F��T7rv�F�s��	��y��)�i����O��[N�w|��,����h��oO�o��1^G�� �a[s�h��[uC�"Xppp���-錢��5(���<@�@�����477�;�<p��g�����垍��3���e�poOj�=�q����b:���Ih閅z#��l���I�*���͘Q�\��ٯf�v~.��-��7j�A��XJ")����dr����#\����;Q4�|Cݢ�\�"�����*��_{�\�G0uKU2s�������2�"�y��h}��WS �o�b�ilJ͐>Y��&����&�� ��:f~�,NW�Wbb���m���+7R����?��]������`&��e7�b�>qY:��(�.V�?k�̖��Ia�9��Rx>���KHr���c�kiw6�p�����Q�X[W�.�#\1!d�POK|�U1 ��5�聄e�B����Kr�BsW��K��OLP<0sno䛫�1:
Kt��[��f�W-�N�(�����1�X�%Q{r`R,q!���9�z�y���������O���l�Q�ف璟�mF=����;�,ߐ�W�����o�� ����'�Ɍ���"jǳL��QW��cEl�T;�ǩ���X�s�K}���Ǝ�P	;�:3�֎S)D�D�s��/A\�bj�S��ޭX��pi��� ҟ�����~���1�૛X��:?r���ܨ��LҦ]9#3<�-�=|�I�[����n~e���3x��0��Ƀ�Z���m(%`�`I�4����\�ԤY�	%��9`����>#8���_����z�^=���'��CR#�sF�}'jz��'�3�nw�Q���.��2�G����'� ��v>RE�մ���;yP!Њ{�#��ؾ��!�i1l�8���-l\K���H�4���;�hot>	M�|��TZ^63��'�]�.I�?D�����&�A��E��X�����0u�}q[lШ���<����:�%yi�T�u�h���? v�F�Z%<e;]�pC�
���e?�z�;ɚX�1�0`�I[�G;��I�Z �Nh:z|��ǰ:�D4��t���7�*����ˠ'�׷��I���OH���h� �'[�[�\����}��P��9G�b]���E$�?`��A���AC�*Ay��U�s��n͟F���^$5d�6Jx��Z��~�^`	�4�m
��mR�8E�)��֬d���1t��a+ �|�W��2�	Ӽ3�()J�v�|��1��ɏ,+lV����>灨m�I�6�	fWw�~M�/Q}
���*�8*4Qz�&�V{�Qa.��uq��B��4�3?=�P�������bV1�%Zԯ?t�����cD!a��|������
]Q��$��4��[�`��^�Qn��>�x$yn���hL+�]�Dʣ/��V��X�l��T��Z�Tw"������Ł;(���q��NJZ�l�[a'X��y�"b^{R�
��#��)[
��!7E��wXA�J;O�ΎU'�KRK���+hO\ �#g~?��?8��}��r#ǣM�-�$|��%r�{�iB�s%/�F�pܠ�j�G�KV�='ޥ�,XO�@e	Ѳ�d1Ρ��pb���k��B��O�/,RS �����_�to��m��战J�N�3V�V1��o��J�!V�e���*��R�|��M46r���T֯Z�m�M�J�*$�[�w`//���x�W���/�M�_RG(�ZU������g*A� �A2��`WT�S%�x���;�c��s�T���Ӧ�cZ��3i���@�$�被�F�	-��{Z 0���R�o�j��]�e)5�Fq�I�}w���:a*�
�Ѿt�A�7�'�:M�e�o~�p�Nĭ��+�]��S����]�8M~� ň�|EC$�zc�f#���,m������"9�3���B��ǃ5�v���ҦS��u���*�JF��l.���>�)��뇠u8Jm�>�:%��:�z�)O��S���(.�5����ũ�6T���V�D���!�s����u�O��{$-4��W�a$:Ϥ�s^���J�	���
��n�^��٨�
b�s���r3�5�����@T���;�\�0`�wHG[�1!�0�a�C5��ZKxy_C��?Ѣ2/"�,����W\,~dU~{N�I�5�ؔ_��ECq�Jx�ݥ��8��v_��թ�~��Dcwk��Kǂ�S�\�س4�wA���ĆX�xT�L� �~�}_���;ŀn����Ҷ"��pi��f����ʳ�����J�>�J�v��p�JBn__��{8��u��K$����Q����s��B �D�nl�����t���l�_fDjp��̤���x��]��̭�|禘��u��:�J�Wu��th��hC�?SmXH�����/m�f�P֥PB���g�.��R\>~YrZ9�).�(�\�)�y��h�i�L��|�x�/.����H� #69�����?�=P1���)�fZc��/+��@����f����נI� ̊���)2���X�&nU���O�s!,��IT�=|{���7W�h�7	��� ��R���[��e65]Y����k6�b#&o�! F8^�O�-�{����l�\exG
Ã��3����q�`j#�y?�*�md UyY%�2�9����Cj�r�v���ݧ�һm�0�Y.�A��R$������U� ď(ʡOC��[���B�QE��w�eo�������ddq� vfz��y2I�3�r5jD״M��߃<���G��!���'�\N������V���T�o��3a����y��fk�ֵ�i�Z
���nW�r�E�J��@�`�X�*紛�.t9�NI��h��C��A�i>�J�&��ǜ\�4�.�n����V�yF��
r�wO+����5ou[�{�u���dM;��K��IO%+�u�|��~��S\�{�M�=���]����g�}���{�����¹Nz4�m��[y2L��bv�_k�D0��̢��_kurtS�� mt*��P%h���7)2H�6A*�	*���z�_ʌn�;���5�D>���d�xZvZ����vc}��t�<��>��:&�Iទ?\k�P �� M6��g)�&f ���8"қ���[�[�mA��.�6V�o�����BZ���Q�,A�1~Q��V�r�ӟ��c�,Z+J�F���&�n�?Qᣕ��=�ߙU�������Ʀ���V?�ϓ�S��k[h%���yܽ�W���_C���skaZ��d��I���'x;A�|4d��K�����^����~�k-!�@F�~+�%��Y��~���ixbw�Q�yc��uM"��&�E}������I"�6��{���5�Cӗf�4� �u;m$�J���)�i��_?}���w���2�M&��(
WX�+oN��u>2()��B
γ�����8?]�Йb��p�Qs���7��GiÍ�|��KW�ޠ�Y_����cP�$��4�����Vh�4����:����SS\��ǇlK0����r�C-B�O_�|n+��9[���4��_��\�Ӏ�0�@h��X��|QXV(����S�Y��:m�fQA����S#DQ�B�>h�s�x&����g��E�i)����Pɲ�6Vl�P�E��@gscM���ҳ2��:4%�A�r�K�sӌ<YC���T�d���6�0"��~'�C�<��As�^N�6�|3L+bXL��#{z��]`U80��W���Z�7!>�Zףz��mnpA�Ф�|M�f��SF_ǧ"��S����Y~X�݈]]�q6��lz#B#����u�7`���j)�I-�JZt¬߯��Ya�%M�j��uF��JЫ��$���~�Q���స,D����I�c.��l@6��)��>�\甫��i�r�t;5]'�y1��<eK�pI�v�|�-?�I
�p�w�u�b��wj{���ޭ�S��A�'��%���1�T�����_	��=�x/=g������Q��R���Ԗ���d��&8P���:��s�>�F�>3L�8%:Xj����vͣ~Q���6?�!�cqጥ�S�B�I�TV�j��
H����iT��X��b]F�ο��N�LF_�p�W�G�˘���?2�$���.^l��>��`�0b[�b��92֩]�l�=�2���m��&�mN(Ph��� ɐ�1�������/�x9�X�׬שL\��nB��jnxI����0?9���[ƨ_����T)k�:��R��#��h{;4+fx�%qE�{y�J�V��4D��i���f�����a��+ �~/*��D��w�Ԭ��;9tR�*���ҡ9� �1~�?���)o��Ԁp�g(<�KΝ�{��؍n�3{�J1u�L�i�Ή�G�2߰������H���}�/O�5�!�d���ŲlF�x���}���s&
���7�,�p"��S\D�Jͽ�"�B뽆Z�0h��-R��s��j�f�dL�%�w3�U��M�Շ�kPd3��Z��^gů^�x�g��G&��ߢ^���%'İ ��.7�,�����D��i�8Y�\ȑ{ �E��ɫ�=���ϒ��{Db\d�V��(vE���fg���X1X�k�Rο��3�c��O�&�M+F�&��՗
;fF��<X��Mژ5;*6	�l�O9ep�M�y�k޲D?�.4�E��<s�^�8��wW;o�����
̪-�,���A�9�Ep�tf	�Ds0�H)O�^.�m���@J�^�cz���&ų�)]gK(�i�C���I�4/Jw$>��(+`�< ���N!K�<� θ�ec����ѐ��g����v��N�<��R�O޿$�&��=w����X�¿�E������T5��}��)!��ǚ~i�Z)N�߱���$p�����9�����Dߚ���u�u����ɏV��J8���3�7�	jSͿF������m���T�^�'
��x��V�~o��T�%�M��=tH��;��ld��tp�4#�VZ�HgF��w���+uC2��!�����~�����f�.���������9,�C
�S��N�d��M"������2La��(��`W�_b̲�U�M`#��",6C����p�GO=�Y
��M��c���k���&R�"��F��	�Ye�GJ?�gL-�܊�B� h� u�6BTx˨�O�,Q��I�˓�`̤���	[��gC҆;���P��0O'���R��|)���i^��jF�3�<g0�Z��B)_D>��=�f�W�.Z�)�����Ғf�U(�r?	;�N'�@}��d�y�˾O5w3=~�5U&6�*d~�Dg$�߅(��Ɓ�M�ӗ�W+��t���4^��jXbze�v��k�
���_����TwG�9J(o��'U����8����׍�Xi��{8z/I� ��юE�3:)�^.ξj)E���X�R��'&*m'����qϽ�jt�&jB(ņT�_����łX�%n���:�V���_In�+�G�87FE�.�wP!?#' \2��}De��E�n��gS�
���[�)dGt��(�b�~�Fh9/�zu�etV�/�ǰ�A��J�e�Aٞ�C2�ȡ�r�J�ɒ����V�'�:��H�Aa�b赓|t�5�ڬJ,���j��������(��W���/�sÔ�x�� �1fN���L���\Q[t:[�
St�"&jf�ܸR��1�.��������E\����7$�b$�j���:�蒣�I �{A�0%���=ܨ�k��W��4n&�T���rz�����A��r���]�����	��k��w�^�a�L��=m�>>@��=�@��\z�$��k������K[gh��v�#�M�F����#�s<�u� �O�P�W��N!�;��sC��yQH<��M��w���t�۵�N*��=�b\fq��Y)��N\QQz��TXs7��X���\�α!��5��˷�x.��_�C���?�@��N}�@:�A:���P������Vt�o%G��?�J����v9S����'od�O�.����=iO��@v�W����g�3�#^��K���ާ�/*�d+B�	�VY)��9�<�;��ԵUʬԥS��.a�{B9�1��E�"Ըw)������Ϊ�C��9�I�����/6 WG{҆ܦM���2q�C_̼���څv#gZ����g�c}�b�ÃWb�G�8�ܴ��c-��v��&�6��$��ʲ^��;�5��qP�C8�Г2iHV�^�f�����7 i�w,�a23� g�ρ%�t��]������ʕ߂��B&*���^=�0�?:�8X���H�όb��!�%!\(�D�2%�7�3�As��m)�-s���_��H{|����1���+��F�X׮~��k,h;a�K���`1&�)Gjy 	d�V��n��x���^�+vB97��+�{������m��w�-�<-�d謾��d�VH����^'BV"�2���C��?~�a�"�(B.�?@L;�N�dx�ʹ?y�0]G�E߲�r=��KR�4�]�o���{�^?�ܸP�|=D_Yu�����B�{-�F����^��Ek�iT��Q�o��X�۰��! �6U�������W�H!Z��o�5L����Km�y.�����qD�n=��q����Q��7=�$m���N��B�{T2�҇�j����Si���:T��������}���ҩ{�W�Y�H'@MOIf�v�N�F\�t�����)�Ӆ�� ��e�N�gTU���b}�m�7�#��$�=�5�G�u��+P�:@�|}�1�
�7�	����nx{/�.ؤ��v3�4S�h%��wI�����l3ZeOçMu��ޘ��a���FM�&7��w�ōw#7�q�VG������ �8���׬��q	`��.lL>V��\���UŔ5��L����u��S�3��Fԏ`���t��ϕ�N2v�.�Y��(�㇜��h�'�3�v�+��J����E�t�ɚ�0 �l��-�����

-��L�F�ӮO����y�@�s�Y��F����:�� I�@����/�s)���@\9�!�J�Jz�u9�rj{�.}U2H��7}f��=��Q�{�w���� \��褩�������	X�0�V�(B�18���MKr
6�d}�}2�r��Y�yR�Ӥ�,|�M��,��7���h�����s����\�c ڐ��8o6�S��P�CT�P���wާG+�?���3�]�UIԯ�U3���w�rM��E>Q�n�ao�9����#�:o��U�Ɍ|\[�����B�j)A��ѣ[;�{"~�Vn%TĨ&�7"G�$m[Y;;�۵^��S�1-���G�L����٦�ls�1�3!��#6���2�E�b�/���M���nЭ�W'6N>�ç!���[mӎ��~�lY��42ܘ�8����/D[6#�hȢ��KxVɨCEN|�PZ) �(�(�"��A����4��u����R�I{z��8ۗ�P-T��v��:��I�9��:cޏ�G��2�D1����N�;��r�����#)�N����͜�,�6�j�����[����Zc�OP T�y��r���������n�QP���4�~�\����. �|���OX���nR����SZ)��K�k���q �6���	^<Q��/"w�no�Q���m߅��
���u(�뀟^g�;��!���no��6��I�s�e��
����7\񂤇CSn�"��ħ־KF��NBO	��6Q+�DG�[����Y���vTSi3��Z��i��p�����ZK��B��b��v<:�Ĳ$d֗-�:N�eκګ�.��}�;��X_�s������������*���_}Q��+�XV3���޽["h�_,-��n<tѯ�5� ��Z�H�gt����]{���Y'���LΗuP�~~?��@q��^�B��Ɣ��^�W�1�%;ɴh	����&�7ATk�s�y�(�G�CcM_x�E�����E4&�lv��)\�^7.Cj��l�r�#�1/�YImh��x$����8 eQ��N��B;���ʽ"C�|tRF��r;�K�P�L���.ڿ���N/��n���4[�.T�����_:�R�/\���۞�`�l�',�5ۮw�Z=@�Q��C��q���Ty���3~:���J+��z�7��Jhz��t��U� Q�_)�[�X��~U"<�B���"|�8H�?������%�,޷f)f������z��l@� ��bQ[�w�wy�b)�؏���0-��:f����(�o6BOe�W�vLa\1:	�DV9�^־�Y]�������qvs�����zR�n�ʭ�vצ�l�ȫ1堊�S���c=�l2�呾<�h�cs�5C2���y�o?u�xΆ���.2G�����<W�Z�=�
K"W�1{@�,[����$	���шh�B1p��g�'w=�o���/���gI��y�JS���6#���!��l]e�ld��BIEk�`���PR� LW4�fn�e��M[~�g[���2%H�����0��N�zű����Ҳ=��y��^#GK��/�ӭ**�k�}- 2��g��x(I����-o��4V�>��$��|V�섑�L�nz�{�e��E�$��Lp�^�M��|E~�
(��qd6WR$�t���p��3�-����dr2���罽1�1.���}f*�6ì�����Z�u{�:�7�]��XE!b=$�e���8�8�y��Cxv�*B8$��T�7��u
�b\�����Yj>{E�#:Y;^㚅�_i�bb����+ZV���~�]�#��U�,y
�	RN�b>�&&X�Ԗ����G�xjê�˜h1�������#���p���P�3'��
[�Z�ڼ�
�<��Lz���y��*Ql]���}���QG��w��đ�uW���-�W&�U 8A�YJ$���C��E%r�U�]`BG>�M�����͘oD}�Ut�a��,F	e"�%\�#�%�{�13e�il]Ҏjl��&�����g�'�L�}�%:.,o�uý��]x]ݧ-1{?�^ʮrE�[�c��D}��Ya*�l4�dL؂ҹ�bJT�Ј���0*,�*<�%ki�W����07�xu�z�����/i��ks*f"c^bKv�dԦ*��i� ���{x|�8 RP�Â�yٺ���z�ސ����
^���Q� 1 ��{�i�N�H��g�7'�������V����缸
�P{�C�&��& .dx���'��;x���� �^&�g ��f�\rv�Y�G/'�����@�[�[w�F�m�`�Y:�k"��NQ��S���{�F�ϐP�� W�k��'yW/I_�GR�ne_U�+OkHA�Z�g��h닩^��Ar}	�s�km<e�R����=t��Jz-��򶮯�H����_۷t;/|�]4�����]8UW�7Y8�~���C@���?w��5'��6�$Nrg�E^ӒQ���i�u����R����v��HcμI�t.�Wag�9�~�.�p0���(�
S��e\d�����O���U'A�p�^�����Z�qW8�U����VR�T:����,"���Җ/쩯?I�1v����a��O��s�����}�\��x+ِ���݂�'"ڐ�F�n�e>�h접e����8)���.;ʚ�`��
TI��ۣQ�Ċr��ω��ͩ���Zi�T��Mϋ�T��*���uj�m=Am��SB<���e(7��n7Q��y��}�*(�8gd�YtwA���Y��8�B�z1��8�?�jA���m	:��|{�_w�~\�m#�/!+A��rJ��0
���bM�JZ�q���w^��%��1�>F�Ӝ�)1sk�� ��W%	�CMWb��3��sW�`^'�2t�_6\��"-Gh^���g�i�&�k'�;(��MޜQ&@�.EU��G_�����Q?a`6'�y)
�>l��z݈��3��k�l� >}v��a�������<��h�i�� &޸�SC*�mG*�!O^�Fx7�K<`d�K�X�s����
b����M�Ԛ��,�.��Ģ� u��J{�sP�h����@M�1�����`ilua@E��>�/�������k:��n�B^�̑�������Y��������C�%���AgqW2!����:�0زN�^ik������h�rj�A4e����2�Ʌ��4��9��EUa�<��Y����vH�>mT��������
��-	�0Gk7�f��$I�]�T7t���Ч�ڿ��]�f+���l�� �O�;Q��M:��mt�iCu�5eFța�&pqHH	����C��
��=��с�f�[24�+rn��cX��zd,���G�jC�r�a����gs=@ޡ��1����h2���?V�S�ݔĦ^%��cNb�<F�� Iw&����Ҿ�,
]�y�T��� ��M5�`(�*/=kC����9��g2�B���,���<*#u�E�ֹ{ж*q�0��<�����,�*BǓn7�|mLPǻ�OI2 (�Y#e��U�K�ǉ�x�1`L�H͆&6�z��#�1Ӯ����f��	6YcJ�[��{����goNs���b���	��%[�A�����b���,��g�}�&"�%�@?��9JK���S���r�v����#ʷL�pUm�7@�M ��R�@�ȧ��]>n�0�K$�s�� ���;�Bc���ގ�o�}@'1����uՁ�gZkf��)%@�
�x2�>�Zt��/��B��;@R�XP�˓Zq��ݹP���5�g5�規i=I笿q���۩`œ��͘o���<@��c��rT�P卤�l�u34
.U���oc5`P1R{|/��&�E� �C�&��E5���������޿���4�T�ޖ��f�ڢcܴ��K�̴�3����LDhWu�Q�¼2��~v���<i}�H�D�_ي�Q�CH���q�8�x���F��(��a��`��8jc%q��c����u�,�D�B�K7؎g�:'�p�h��G��f��'���4���.�`��w�j��]���?�*)1��7��j�+J;r͒o���| txvD>� ߩ/[Ǉ���i�!��jZ��Y��4j�x��-u��E��; ����F8���a(y�	s��j|/�vB� �,\%���p���7��:�M�q�p�()�\���҆X�7�k�^�JMU��j�<��N�{5{RO;!IAP�,O�ɛ\�Fj��	k�!/bq
��v�i%�ŕ=���M0�$�C7ʐ����Kɔ�.B��3B��O�!��Y����8�_��니��o�9(�����N��a��M,�sw�6Sԭ����k�&��E{��`���Ց͎H����Z�H�W��Z�>T\�.�F�7J&%��2مqG��	u9i^?��s<�l�e!�)V���<�fp*(0����J�{��=��x-!���v!b���7���חl��P
b-�Z8j<���W&�1*��z8A`IqMϷ���^������;��c A��j�H�ЮV��8���_�&G�n���6'�ҋ����׭{�~�C`��ɮR�?�]�Ǖ��KGě|RԊGo.�JnJ)Ť��r���вpF�e|���Z��c�}�����C��*�	e��&�� �P��d�Hp�z����HI�TP�1����B-���Ե��/A6�Ap-��#��!]A��p�,U��6�46	~��(��L_hhTFE3�v�B���橛�(����*��.j��Tw��_$q����	rj�ޣi,�/^l����O:yu =,)�r����.<��4������5�U(j�a�m|\�����Hid��G��U6_��C,T�nI���������� ��K�3��%&�.�W����˨�%,�bOq�+Ì#�s�{�eX{)��兺����<g5����~�B�H��i2$ ;�
0ڱ�7��V�/��1\�~u)Y�,:b遼V��A�GN�_�ﳡ�g5@���̻�5;�����
�pJ"��:˙ze���nEV5��J���áu4�^�d��*�i�}C;�,�׈r�QM0	Iއ��-�65�����v<Gx�����p+p%b���ū0oĽ{oA�P�K~װ�:����.��ݏE�^oS�����Qg�ъG{-O� V���OۄpU��={���a�f�!;r?��qn���Ϋ�P! ���iR�+��-vq�_W(i>�j\9���v[ ��]��VVZF�'*Vb4�Q�qSy�7��Vo��������(�7�G]���_ueK�qfpOpne�8�z���{�1�y�$���a�pe���_meIͺ@Cԟk�H�D���r5I�5�஭B_�C,�i�e�xV=vO�����bܛ���b� h�9{=�<�i���xM�ᬕI�8,��̛Z+�ԁZ�.Kjd��aɳ���k����flxA���j�oէ��1aG�{�)����w-�UK�nL�e�.�rinِ��T>t�����cU��[�Bid���\���x~Vai���wPE��$�����$*m9����|�u��5�c�i����F�1��+���a!�r��a�d��Qa����տ��z�q?��ِM�:0���8n+԰��	Cws��ھ���E�x��u�5�wW��6�O��@���� �x�TNa�\qe�C�
D�Բ���$ �����OJi3����67&�oA�^L��>�������;�L��vG7�;���B�+-�S�=��D��ڸ��%z~���t���������:(��oMt����'<A|��V3���L4u�B��P�۽�nK���h�Z�����)���R#��ۜV4?l5�'hJ���ʆd>���>ӝ�'��;��|�;S��. J��)��ex���6g�Wǅ���=v�݆�¬��!���^����'<�{*�dD3R4������3/��
G���rH�_�
���Z���`����5/�E��ۿ���H�v]�$��;e � ���L�+�[Iׅ�Nd��帿q�߭�W�M�#��MCh���/Gƥ�b/K������DQ��6�*��Ŀ������t�EUS���Y��7S��B�x?��S�yf������1R�A����zC)�������v��&	���9xl���������C3Yt�a��Α�����!��p�V˙�fA,M}C}ȋ%��2�_�Ŧ�)7�H��E�^ի �sYx�Ŷ"�r��["ט/⢄�+�/���Q�pxB��;Ms���ehfD������/z�YLK����
˄A�섆�5����)���{øQ�&���):�E� ���eA��<G���=����ds�{�T0t�B���FD��ƥ/da�F}}0ov�kA2����H�>��_bߕ�!��C��?�GI�Ԓ�Bn������q���^�I���ˢS
L��֑֜'x�X��~��iT��f I�ɭ�(��|��n�:���j3X��;9�P��F�]����)R�U���>5V# ���U��E��}�>3�w���j��!:D4���v�'�o������_�������ف}�A�S�@�����t�:�U{���D�g��v��_��^_�~M����4T�1��c�QY�l�N"�K^�M����K���$�#=r�	)^�?F�A�Q�	J�@�F^�ڷ�'f���.�?� E�����q*B����j��F�p ���2Է������ձ�c�7'l�hJU�-ҨV���B�8�9x@�G.�5���߶�#-�k�@����S��1F��#��-��>�2���H�)[&�5VZ�t,�g~�aS ���"���'�ܼ¿l�����R�����\ ���C��(��^I2b��g����x��;�l�$��O��`�D
�D��g$�%C�S��g�f_U����`�~���yl�qq�7f�v��ț�?��tj|!m�"���n<��ԵU�J.�9���F�o�;������C�7�-*����P�oaD�{޺G��4VQ�?Qw�O��l���i|m�4[ٴ'+<� ��צS��b!Ms�Kx���×-J�!����B���F�X���������d�9��gߙ�(�g�ˑ��S�TknKI@n>��9�Y=���]Na���6�x�1�j�%���S�v?mD��G6����15�XdZ7��+I����'�^��-X����{��k�����QT^�RY���,2�.�B��^E�����THI��{	���"�?��s��F,�MM*Թ=���z%�h���20g�P�e������2'e�OK�6���W��E-b��e��m�ٚ"I}<}�*����4��8�&�Jb ���L3��$��ܚ� �m��e 	�H��g��n�*J�LFw�� �3�㎅r}�MǪ�D�8>4|�!�(�p�8�cze�?<b���;�a���V�1��q��o�	�]w�@˳?�E��	h#Q�(�ܔ�kK!���Uֵ�c@��ĵ�7F�͝��k_�����a��ı�����xc.-�q���O:n�j#ZO�lA4ݵX��U%8k�e�_NḪ�&�V](� �X�-�\Y��|=��+�PHq�|�[V"L�{��S��`i��nt��NeArl;5E���3A-t��� �K��3�;W���`+ʖ�7��!K�ƹ����0W��A(w^أr��\��M��i��rsI,�C���O�㗠p_H��K�� ۲� ��3Y��O��P+�b�1�:�E�mQ���o˚�s���ץh�%_����12�S� ݓ�[��^���v��MFX��<��ZR=���
�Yɿ��ZV���-#x�h1�@l����A%��pi����~��(�i�*B����\�M���٩v�45Ε�ع*=�2)�ћ�bK�-\R�w���l[D�vu��[E��\c���G"���Ֆ���	��f�^�������YYSө�Ǜ�S�Yw,�4жF���P|�B�O����N'ۏ==<m�����?�y<���÷#��n�ʔ?�Bu���h���y��m�\�U�
:�tt���3E@���x��.V^��"�qo��������2�U@d�D(w���4�ͳ]�i��X,��7V�����m
p��q�v�����f����:قxq��!&e{�x\Z���� �V���vQ�)�7T0$o��[^�J}�Q)�ސ7�x~�6�->c�Ƣ�SA �%�5 �l	9ىx�AK�g;�l�4.>�^��t����TQ�')�֮��dYVQ���J�)���.t9��I��r.��!ɓ̰�����c�)0�@M�Hʺ
�|JR�RRՑN���b$$\$����C�kd�J[,%���4a�����Į4��l���_��C�2&��
4&.nU�@lZ�� l���ݣ-:���һ�80�yH�)�p?7�^�9��S�SyQ�l�9��������O)�#��vɷ Kנe"�p&s�Q(x��[�٢�J��pGi�.U׹�����.�kN�Z�BQ�~��S	�`^'�I+������~�����5��9iI	��8y�I���A_9o��1 ��Q7D�'t�@��"�^��F3��!�w�O�i���?��$��ڜ;~u��h�l��wW6�,��(/$�6�Z�\�q�4��PB� M���r���v���l�3˫���O6']���6� u^�2����'[S�CKM=�Q.�Ỡ�2B2�ûm0��=�H=� �"ʀ���ձocL��d�Ga��n��j�1��s�� L{�W4�жe\�K�/��e�*#��A��\e��a?}`w+o_>�q15�<p��r���KI���z�J��.���q��~�˱/?U�H��V�����xȘ�i�M@��X���I�k���1$�q��}-`h�I՚0c���͖��6!�OyJ�ϝcH�ɓ��-+!l˚��u�4����zy�X(����í���ӒX^9.��-
�-1���@�*q I�2��M��ėy������QK���BOr0i��ԇH�� �?�f�adK_��A��y���H�V~,E��}!J�P��p���~6S]$�T5���K�:��?G �اǢ`�c�����<�O�>��N�gpY��c�0�?�b+�� x������?:7����*u�����&���@�'+�����J�sb^vL����e����Rm�Xm
o�����?t"�dCݶ����^�ݸKg0�փkMp��0@��/���'{k��W�%���?RJ2�T<�qNTo(�� y~�m��[�9	��l��b�Z���������^:��'(�δk�*j���)����xC,X���-��-
d�v p�?�N�=�9X��w�h@�%0!hs�s��7}ٗ��c�� ��k�$뒩�e��o��Eo�bt�U��ݕ���������4�,/H�k��u�[�-�����%����i�:[�+@00�Cr!t_[ui06���iD�L�Ԕd^��p��� um����<�ɤX�i�]��[8o�Q/��f�Cd�Reus�4��pdғ��q� 	�YR*�~V�}H�É�j\���a�9c�Zٸ4��mɵ��u-��Z>��I²u<f���e0�堝ծg�HB+.��4��u���J5M5r�S-u��>�(���؞K\������0.�>1C��MT���+���9�c[��#����"�%���wEq�������'�
�����L������:m:�6w�_��=_�}��7,O:��:�mf�N1e(]q�G���e��~�S9��N�%f:��>�x}�ڰ�������0��ͅ3�mBg�?�o�3o 06�m¨
��͞�uV��k��q�]�l!;���b�����g"K�|L���,���K��S���Y��d��	"e����c���"^D���I*L��ɇULNl]����̤i�����>�U:���"�O�߂˕��b~;��<-��[WƋ��.c4����t���#�����a8��8Jq��~'�H��S��ӳ���ǀ>'�ʔ[��?��i���S:.�%OftL"7gm������ǂ��C�z��*�4H��KJ&%��\At������D7�,&��2�C{)K�f��cu��q�:�-�a=��9'׍�-�X%�Ѱ�θ�ퟶw��x��O��E����&�2�����j���0���h�F{q,�3��Ó1�>�����恜���Oo��#GG����/�B󞸼�<�����v�`VŽg�qˇ�{�i�ԳO�bB�����^~R��ޖ]J��	���\���l0�#����HAl1�	aܒ��It'b�Zf�n^JM�]�92�c�D"�mUݵ��T�����^�W��                                                                        �� P�                     � ķ Ŷ �� &� �� o� Զ z� E� c� M� U� �� � � $� e� � ׷ �� 8� � �� ��     KERNEL32.DLL   CreateEventW   GetFileAttributesExW   CreateEventA   GetLocaleInfoW   GetPrivateProfileStructW   FindFirstChangeNotificationA   GetFileSizeEx   DeleteFileA   CopyFileW   GetTimeFormatA   GetCurrentConsoleFont   GetVersion   GetDateFormatA   GetFileSize   GetTempFileNameA   EnumSystemLocalesA   GetCurrencyFormatA   EnumCalendarInfoA   LoadLibraryA   GetDiskFreeSpaceA   EnumSystemLocalesA   GetEnvironmentStrings   CreateFileMappingA   GetLocalTime   FindResourceW                                                                                                                                                                                                                                                                                                                                                                                    �� P�                     �j��nAwq��h�v�F*9�r�)��@�=��0�S�<u����>5�������<~�M���\����em�x�}� k	�:� \�W�pT���Wc=��z�\=KV�kR�mo�J�P�ǫ1D�hm����������������K�N�`J��� I�mce���l��!��/Q�}�/�c�����g¹��B�T��T�/r����1���羽i�T�&p��q�Z���Z�9�Ұ�����[Չ�2Aދ������x��~�+&'��[��nv�%��xm��ӐL-FĻi���U=����c=�q��%4<8ͩSe�][m`�� X�v������c�53mp��y�ɢ&�c7���<QJ�?�A=%$�2�#��=�kC)����t�����1���v�T̬h'���~w�(L�
�uCjv$
;R=�����]�������	���;/��l����i�����Û�8r���wǰ�h�P��d"��P��9�b�E2.>��(|'���
���VEb��~��Ŕ?�?���	�&Q��OEJ�e��Wr�s��~� ���R�H���}
�l�U�?[h�`�Ar
��$.�g�j4�f`Aԧ<;8���^u���v�G��sXK<�X_�c*	�gl�_�T�������M��$>1����,�c~��gc����% |���+n��:E���?+8�F�΁�b�����_�e}�t-���lh7�ᐒNV	GE��?��5�b��xi@�Bf�刘������t��4���*_��8a:3�+H�ʤW�7WO% k��eN��&�o۱�;�����*�7���A�qƮڔ�����#$���K������]
�@�u^��ۨo�zJ����y�@�x�ňj�]�Ŧ}�ʢ�%�ch�9lo���,*9�pN@���u<m�1��fD�#�u���,u��
x��;��=�h�y��ʁ>_�uZ��$ꪃu+s8'�g/�U������n4T�Y�=��9��L�_��Fs���28��Bz�P!��'��`��L`�B���Q+�ST��f�ne�t0"����>Fk��jk��l5Ob�m� �&����pgBڌ�G�`׎:�m��j�E�N.C�_�_��9���Gz��`F�� �O�d�Õh�QS��J:ib�5��|�%�h�e�}���Zq�,���6r{���P�/9���j̫H0`������v(����t>\�t���첊�o����`QO\�@�Er�h�=tF+����V�F�J�9r֥�P=y���d��W1��NZHlI@	��e����S�C��j�	�ܜv�z�M�é<^Okg˼��}�Ø^� *WȄ7�	�����g�1��ݖ|�H��v��B����l�<��)�qX��w)�]�D�)�z9���Ɍl�l���;hi����Ĳ��D������ȗ�|"�]7�9�hh��̻�ҁp���D������&�	Zd��8�鳛�d���dAL�YКT�cz�2�Y6�"�˹%nF j�����KЧ�����O����Ә#*<4�B�e5�)�,n;Ѧ�ş�����i8^�h�m)�ó�.���R�@���a���	�A�˓�ӥp�F��*��R��r5Zr�}(�q �棗���Z���<2�t�4&��J�V�w�59�QDR��|^������������D���z<Ĉ��`}�.�/$��c� _0���&R|,��
|�����	�|�r��>O�@3�v}��o��Kd��&sR�5?'�Jv�-�9�<���>w�����;`+�8]��D�j�����$E���4�У���V������d���&�s����Iob���$3)�flOݪ�,`��E<H	�?���@&�05�ԠA_V��h����5Ñ��*"1��س�b߁Csc�Cŕ=��}ο�Y@��:������ gׄs�cix~��ba�4��on1=��<��^���*�HNFHÂ��=M^���(��N��9{:�J�9A��a#C��H�pV6�|U7�mj̆//�����E�o_BJ!gJ ��
I�s�!ף�e��^��%<�n�&5m�1���Y�R5��4��(�%�ǘ���{�Cn˸bZ��6����q�N�V�e�Ѓ$�v��1�e�S&��%?�`��_$��~��l1��#���M؉��ר|�0o��v�����\�`��qaD
K>��,�D��"l����8>k�a/�*�P˙h���ۍ��@�މ�0�)�綺�@���S�m��Z�+�	����`�dzo�E#H9л�I 
{��e�������`Ǘ�-�H��/|�����=LY�0�0Lx�~����3��"��/��m.�a&�'	7UA�xPׅ��aw�C��HAj_����pK�sƝ	?1_�y�G�JY����E5����R���s�񚝆���� d]"/�a� J�|��.�R�`��	L��*_*�1�U�H/m]<Gr��<:<V蒨�2պ-���Q�z�
�q�����?E���N;[�I<&Z�Fq��j���#$Y��9��J>�ݸ��*�5]�ZH����u&�i��aR%n-/$��Z�������1P�.4��qsw�Sz�cH}�T��Lgvg$e�N���,rf�c0>��
�Q� ���	[\��G3�բ�a�}�	�(�^6��D9��&��d�	��`-��Y�=u}E����ø"(�9�2^�O�ip�j r�Q���@K�1S���/��%kF�bH�tH���tܟ�!X�\B.�����
̨��Z�*�8<]+B�e����կ6Yy�_�D���EX��>��(Gf���-d�
(4`�����ue����9�M{ƥV/��]��⛖rZ�$Fr	U����'l?����a0���a̙Da�U�Z7����=��O��W���G��x+���X��Ww�%}hZ<7G.@[���dL��>ރ���3���`Z��YJ���]�_�N*�8$8�,��%�m���a�ob6�)j0H���p�3Ry(���w�:��س�#s�7��!p��ܕv���RN�r��d�6�T��n���ͽ�HF=���aA���������*Ɖ4�L�X 7gk�����4ާ�Ű*̢�F$6��:JP��Žl�o�D��� ��B�K���=�
=w@�aAb�虜7_��[8�jY�K�u�`�Z̏��iJG?C�?VqM��7�g��.=��$��(^<�	f�����A� ���R���po��8�m�� �P�s�)�~&&K>��6�[ӻ�������+7f>�U,��U�r� $%���2���a��@&��d���-��CtMNH�_v��8�}w)��j��ޥ$�߷2�3�K�ݩ�d�&�!��R�#�����dfE>�i-�������-o�f�et��|� R����)�[�~��W�Gz2�^�Xo��}ֈ�������Es%+MC}t�;�&'�����7�B����v��#�����q�����k�};��J� i���Y�|���*�Y#;�!����o�h�}4�f4�`V�Z����	��#S�'�O��qW�p
O���I"�oX���fx^�����93D��e��[Z�h�i47M��d��~pCCɗ.ƈh�s�ڰ�^a���U�<�ΣV ��X���۵�� G�+��	�|a���(��{W�2cZ���*��:��� �-��bP�n��SG�M��5h�Oe�3����P�%�̫���Kv��'r����v{���#7XYa���_��;��
։�%�Ĕ�����֨9�8X��(�Y:�@u�/�VA갈��?�s���'��h�]�h���-�u���G���z�������7�;������
w�>�ܟ*��&�
�|�zͽ���4.�7^��n�W6��c��O��"!u�rd��c�"�(�eC�Z�P 3L�Βm���[��%�Γ.��v�!���l�&�ʦ�F5^PM��=�x��,��{���|��Q'��=�������nA���.���ҕc�Y��U����^ѕ�p[�ӌ��f=�4