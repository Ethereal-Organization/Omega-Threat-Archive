MZ@       ��         @  �    �������������������@   PE  L ?/yF        �       @   �  �         @                      `    ��                                ` x      x                                                                                                          �hk0    �                        `  ��hk1    @     d4                 `  ��hk2      @                    `  �                 0  $                          .text   �                                        �                  0  �               	  H   X              4   V S _ V E R S I O N _ I N F O     ���                                           ~   S t r i n g F i l e I n f o   Z   0 4 0 9 0 4 E 4   L   C o m p a n y N a m e     M i c r o s o f t   C o r p o r a t i o n   � 0  L e g a l C o p y r i g h t   ( C )   M i c r o s o f t   C o r p o r a t i o n .   A l l   r i g h t s   r e s e r v e d .   r )  P r o d u c t N a m e     M i c r o s o f t ( R )   W i n d o w s ( R )   O p e r a t i n g   S y s t e m     D    V a r F i l e I n f o     $    T r a n s l a t i o n     	�	       �      �                                                    >                                      �    �  �                 �&              x               # 4 E T b     p     }     �     �                 � $             � @             � H             � P              X                     KERNEL32.DLL MSVCRT.DLL USER32.DLL ADVAPI32.DLL SHELL32.DLL   LoadLibraryA   GetProcAddress   VirtualProtect   VirtualAlloc   VirtualFree   ExitProcess   _controlfp   CharUpperA   OpenProcessToken   ShellExecuteA       �        �   0  ��]y��d.��`�   ����a�\�������`j@�<��$��������  �   �Ջ�����+Љ������������,����6�����h   h   j ��`�����'묐��������    [�T  �PS�  a������`a`��   e]��   ��������뾋߃��    WQRS��d�����`����֋ϋ������  ��[ZY_�� t����h �  j ��������d����������N�V�6���� t?�G,�<w���z t�8u�_f�������
�_������+�Ɖ���������*  �������A�� ��   ��+qtz�q��,����6�^����t
��y�I���y�I3��G�t <�w���$��f����u�����3ۇ���� t��t�f��3�����t�f�󍽸������������uBVVRVjh   R��\���_^��B�a�^����   ������V�v�h   W��\����݁�!   3Ɋ�� t(C�������VQSRV�3�s�C�P��\���Z[Y^����e� �����������   �������> u�~ u�~ u�z�^�SRV�����~��W��T���_Z[�� tY������>��3Ɋ�� uF볋��RSP�8�u@� %����� QP��������X���YZ[Z�� t��F��v����F����   U��u�}�����m   s�3��d   s3��[   s!��R   �s�uA����P   I����D   �.���tO�����"�H������)   = }  s=   s��wAAV��+��^��u�F��3�A�����������r��]� j ��h���Ë ;Qu
�A8`�ÊB���D$�8agV <ЃI�j�X^��s��� ����N�|Au�^ SV�q3ۅ�W y~,U��9���;�r+Ѓ�:����s��5腉A� �Mu�]��b_�z^�9�[g��.��W�9����x<�� ~;�s@�cF��f�4п=��+��� �f�9�~�P\��)�*�N��:quf�r��B+О��V���ޏ�
���ꡞ¿�F���>@_^���QSv}�(����~�]���U�4��>1�?���M�u�^�B����_[	�*:3v���90W��B9}����P�~ V�xB�
�GϠ��	E�G;H$|�6�H�a��2���@�n���Ϩ��p=��(|�V[�jP�3��(RC�7u���e����F��L�vG7�s���;�u��C@��dW�E�vEY��3���Å�V������A��&u*�W�j�L0aZ�܏1�;�N���2P$Wu�K$D��"N����j���B���,�|�8�&T��M�H3G���HRzQ��יM���Q����f4K�M� �@����6Z
2�JO�89M`U�.�sjX�ᄘv�u���n��^@���f�
�u@�M����G�} �p�]�$#�3 ؃����fG��� ���N�U�dD��vĂ�#�G��*M�A��!�G���@ 	;���l}e��${
u=�r�
���`t ��s+`���y�U�Ae�l������T)j�C�~�i3���bF�;�����d-:�F�/��/uEIG%���
F��uX9��j�U�(�>���+#��D�	����r�f3�Jc��J�HX�DF1u�H��'+VȊ�.���	uv���p;�m��Q�E���h
�2�UՄ���#~H���ϲ#魄����[���ڄ�,�dR2"
7�P���H�|�}IX�(Q�zI�&`K�t(��!|I��я�##�J��a��1>�*]}HQ�;+�^N^�:�]p�!�����H>�E�Pj�"�DZ���i��	b�����I40L�y<w:~sI��8B�Ǌ�@9A@J��C�~;� r�����������+�n�u�xâ��]r��������Hr�D閕�U.X-.]_ r2�����]��T����Hu�<	uM�9��-�����a��h�$��L��SR�㝚wA��!zC��(�� 䈤���$e:@3I��Fn�j�.�@��
�_�=��0     ]    v&   �   *�و7�d����3T����8�R�Ǩg@�_`t{EOp�䁜O5ȃz�^Hѝ׬��:�[b:?G<cΣ��ո1���L���g�h����d���Y�@���D[� $4fs�Qh��4���>@�'����}[���Q�%��o�a)�ȗ#�v����BX&R�pCA��	� 5�wdı4��m�~�{��6��=�)kt� B Y�5���M?�
s��Lp;W�u��f��oet���Yu/NϬ�kh�9����{������`Y�Ϡ���_-��6դu�"��[^�)�[_����:�[cvB""0n��nh�!���5�x�
��h�c���cw"0�1ҫ�����5m�em w�i���غ�a`
�Lr-o2��v�G/�C7[��|کY�>)���g���P��,S�M�~cC��y�碛ȯ���B���?�����T�[��_�n���>���r��>��6-�LY���U[E����H��y���ӎ-Y�l(ZyC��-� ��P��g+���LYXS9TuT&�k$�F�&���e�+9R,����躳{�Q
K��0��X�ML�jC�?����e7�Aŭ���1i���/�����͸�n Ы��an�XCRA�z��]EP��YN�H>�,ǂ'n���Bl+������Y)�U�^���)hsѱ�Z��d�!����H#Vu#�og��1��ia	=ZWsJo������(�)AT	�.B]���	���W����uB���6��Y3e����S�?oP��������>z�eD<����G΃;ٛ7���t�����x��r7Cd������
���r�ޮ�	rh�`b�������XWz0	=��9�n��϶�JU���t��]�Y=�ĦrM.Qy���c����<;�<�(=y����L�V�-"��n&#?�Φ��'�~���A\��.��N�B@Nxi�����Fo3���V�<υ�e�^&P��b�~�ӌ�j���뭋Os�KC�e3[�W�KM���QHc�����V��5DJH�_�Z�s�v�}j}'|�U6u�z�����Q����[z� >D����+j,��"Ό�71��3�j6�n�×+�E�H Ï�:Y�W7��)�������A��:�7ƏS�e���Akmb#�La�_K�/EH�IR�!6vye�;Lߘ�$��-���;�Ѿ
����D�ň�gI�@�2˴a!�xl��cKel*d!-* ��㎺Q��/�槍�WX{����P�6��@�ć�V��/�'��Q6��؜��1z�2G:`q�ѩ���_JtI��)ՁA�"엯���ind�`�-��	��9Ӣ[,!�c�ϴ;fX|��I�2jt��&����e���%#�=��0$9�W0z����ֻDIF<�(��^!Z��n�B�i���>�QV���������G��POs��?qa�:��<�H���^�3���u��K�P��x?��������K�F�<>�Iz��1�[�X��(f.<�2�M�,��2�� �e�N��P�X�ңB0���BO��H�ss�J��u�� �I�9
C 
q�����!�hV�>�C	3�{U|�e���	F��j[��s�h����T^1�g�Ş �/��{���2����'?��MA���9ʞ�9x̑��@D��z"�Z�^�#����/�]�RsdrJ�R���1��~ ^��v�&��xh�.gp�X��TuQ��K��?;�&u��s����`��j}u�H ҫ9�2jC����u�͠����gQl݇ 2���렌�P��= �"Y)ֆ�Uv���̛6�e�,n��{�J�)��ReW;�kWH��DB[�q���k �q}Hu�,/	=��R�4zlA�i�GH���%�6��c�H[�L�������Ӓ�nT�vH^��^:�S�Y�P��o����w�{�68ߴB��7�v!٘}�����5ǼJ��࢏����������\�T
Yg#R�s�������dC�;B�2�(�*�^qk���{�AAW(���९���Q2k��E��(bý\l����X�bc�<��̔���1B2"y�΄G`�:O�U����'�;�
�L2*���/ې���@��h�^�J	>�m�gE��z^�K2S��l���C�Nd��!�} �Yڦ�,�\�����R��"��d7u�!i�Vn)\�ٮ��C}2��n�>�uD��(l5��QwA(R0:�@~�~KsNk
&�rĹ���?�L�9T��� �(���A�=�Sek�J|M�	�q���Iw����N3>�`��	�ZR
K�sZ��/�FH�&�4c$"j��}זR�+�Ifw��a���sQ�1��׿���?������G>rE���`�{,@���_��c��U�����
��ZL�קÍ����7���m�7E��v]�J�4a{[Yq֕��g���0Nv:�����dA��hk�h����aǦ$::����OSsE�4nl�F_۟�|����}T��]�{('ؖ(�ɫ�}�L���H�#�%�F-����(��F�3$�����O˽��>q*���8��P������O�"�\�FG�#�E����E#�FߥvӅs���zn�n�V�}Hx�C5)/G﷋�e��XѬ�x[�8K�覠�]��s.y��ZÕE�Z�7��6_ OI9ʑp��B��u@�������|�e8�5Ժ�BNR�ք���?2iH�~���L9ph*u�a� N��1��� �>��U�(��Y)g,��R��`[n�:4[8b�馘0�1J��.'�?Ht��a�dD7U�|�ެ�x�����D�ȧ�H��E\A�$]�s�n�B:7�>��sM���ּ�sd��
T�*zy]�h�߮0�9�&\��[�ՙr�>��X��/����H!:X�Oz�>j3��)v�E��m��w`�b�Q+��C��@$��c�R/ȑ�v��ΰ�U�V�l�;?o�(`QێN�>vb�n�:�R��c���\�9�Z����e����`XyQ�L$mV�	��_�ũ=��<��#9' غ�H�r���/�g�̓6�b�t��W��s�(��]i�e��"��W���+2Ϡ&e�A�a��A��0��ŭ�S���N�����a,-ۭqy\��y���Ӟk�<po�di��X	�����7_�
�h~�h{��7�f9A_nβ3q��(Uޏ���=��nǲbLz8��I���9qݲ���y��WO��mV�E�,x���ñ����bұ�|�J+�o�k*x�u{��Ҍ����&����H���?�.�"��5M�C���~$%�m~'�2��_� B{�"+<���g��j�*S�*�zv��^Azh�{Sb�`nޮ
��D�
Qu)��B7��H�lÈ��ȃ�����3��l�A���T�b������C�<^$���ܢi���Td��XT4�~�w}D܉��Rs��&Qk��|Vz�c�P��lȯ�]��������%m�p��� )g*���a���� ��Wb�}����w���<J����Ey۴�m�gR�:5�D�Zӫ���8U��*��{����L��)5�g^�W��M$��{]�}Wʅ�\$��.���+�\��Pk95JA�vX`0Ę�>�J}j:������}�]��)f���q���Ql�Ԏ�a�-��2�Fy͢0�݀�����!���$!X弇�ht*��>W#��I�!6��絤⡯�jzwyo��}�����^xD="�h4�K��ή�Ŀ�ݽ�<n5N_9�yJF���f,)��{h)�%EMS3��`vp�7�i��%!K�(�{6,`\#�@�4��s��"2��w*c�p���/>*��v�ɸߝ�-����
�E[ET @Cm�E�ˈm\��b ������4��r^���0���&�Z�l��k}��qѤ���Л���t�����W���}�s���=�{	|1�@^#��g���9j_��O��j˜�O��7���K�V��ajYU��ǃҕ
d��k4�U�!2?H���fj3�oF����M�����	R/�������p����[TUѼ]�!�
e,;T�6�Q�mA�2��H�}��iF�8߄<f���;�7Vq�ڱҜ�7Ǖ��ПۦyB�s���^J�XQr��`��r�o�0L�K@�����a��9��o�,�3���kҙ��"D��lY��ur������#����uiZ�UR���މدNOT
Y=o��ǡ����-đ܋9��݆g���Ɠ�T���xKTv���j��s��_��^�
�f��������= !�}�� |t�K5��I6X3�Hk�/�h�E�b9,�Y�$�jp�[I3C3f��DF�?�@��S��H���
۠�<����7�y�M�~ˣ�2��O�����ܲ�)s�N�b�P_�{��%�(��7�Ca~�P�	ZPR�y���p�X�q����H�骏Ğ�4X:�{�<��S���t�:��[K�����_�.	:@a��S�����)��|vm�~w��D�<ಔ���]y��n�қ��)��v?�mJu�B�7���3?��h�Y>��O��.��P��/����އQ\���L(������C���c��CN���Eܾ�;�����ޅ��A������}qИ6�{�U,�, ?��V��
W�`�R�n��i�5@���y�l8~m�\۫S��K?��H��i(�U�S�,;yvz�wY�`h~�X2�
I�q��ݟ�u���Y���Q Z��d3`��y�M�떃��}{Z�Ŀ�󮔊��D8����W�h������ҽفpA&���/�J����j�w�W����z���v2 )��`Mߪ����x��>��Y�kP�������nU,�9]�)��±;��seJ�� ��2El�ʑ����51�<w��0��� O|�Ts�<DA�����PX�=J�mь �[fDQ�QH�-�������̰�d]�.ˑ�}�ժsA�'(�3
q9�_�u~��62U�_̈́�(��c#MN���ײ'���t/͞��mA��<�盎\ZH��ņg�0Y1�H�m[5cJ�kfx\;zT4{S5o��-�	��g���t�� H�5G�z! !�j�'�{W�aQ1y�_^�r� ���xm�0"���}�ƹV9l�=���\���A��o�0n9�N̈�`!C�\
kf���x�P��ShSiPͻ�;��F�&�?�u�V����`F�m���������S-ӷ�v�MR7�#� p��̬%q
e�T�ƗRم�6�5���,L�'M/3<c��"4y��B��d�\��;
�0K�@�>���'�j|$,�aeBӔ!x�|�R�[�B�����kc�t��'%��S�5���y���#M$'�"�U�@��ąqT���W���*|��#�D$�nnY�j��q��!kN�j�g�xb��.y)ء<��d�l�#���sh��7��
en�=K�r�S���neB��/�3�h7o��@f��0�����D��4��bO��M�W�B�Z�4� ��c�1�_����g�~j0�0��y�I�r����i��9�>~-��j����H��v�ߓ�co�@B��/�y���E�NYS�5�kE2N����q���Co�zaޮ�7f��Z_��4L�۞��g��6O�lT��ҭȺCp1Ɗ�P,n��퍨�����CQ�r_T�*� 3<;� ڿ�Bs�0��睑���}(����2��k���.1k����pۂ?%b��Q�V���Je0_��;��A�ڬzl#K��=l��Co���!�Ƭ��i�
L����PY�% ù��G���|:���Pt�j�c�h�
nk@�mv^�Gw	:�I�z`���eiѭ�dU�<h����Uu�2$}� +�c�s�
���4���ם��T&���JuO��#��Y��x�����W�v�L�����-?�9O�,K>�Б�-YMc�Ô��cvR8��j'* �P���o�1������"� 2kF�כ�p�S{�t�J-de�u�`���f����{�;Ɵ��z�=
�f���(�K#�]l��`��v#����\���؊Z��0�V�/y4��Bʛ��_�fāɵ%f�G�xT���n��c�Df��*ޘ��j�����#a���6��r�lm���jSvkM9F��63?��$�G*�n����+�GQ��&����&�|짨�xժ�)y?�8��f'�!�خ�1c_q����L�P�!]L�u$�f<_���@tnU��C��ܬ���M�U"o�K! �k��"�d�$	Lh�|Ĳ�����&2�
S�D0��������f�����97lZ���P��S���\��댅ǝ�ƺ+��ޢ?�͸5)��H�}�!�� �}Q�{�����=K�/��JP4)�"�#�������!�*�>^ԡ�T�⊾��L��[�]ܙP~H�]X�(ո�Ȓ<���-0)R��f��&Q*֡�e)��uVhDs� Nv�� Q��}��CM���p2��zx�+0D4c�hzIU&�Z]0���y�}mn���0�9y(���)m�E�2 \k�֧�p�61wY~YO�lGj@����Q���Q�e�X3��P�J��{ӨSf�]/��eͱb�7�^��!:��:�\�;ѱ;�4U�98��ɋ�,��9ʌ3�":\͊�%֣ն:�ɣ��ςx�'@�r^�V8/؝у3%�B���M��;h����V�����E�U�;�J�k�y��J�O�w��OH.���:bc� \���1��/�]y𦤍Lވ��h�u�F!�3]�X�0M{b78@θ�8��ma_4�S�fn㹈�F��דaqF\쇉�����#3$n�j
?�Ң�	X�:���U�ˡ��2y{4��w̧"�}�X�]���I`	�)���������YŎ���	FS���ԩ<��ʙG	�u��31�x36���P�̓|��L���e�@��ZF�=�8���<�Z�l%]�L>��5z�iP�����/��BL���UH6O�׹�2�i��!��8}PQ{Q��cH��4�\�V_�V��I%��Uh2]Mas>m��{	�����G�v�c���c���� ��.dq��lf��b��`���wT�3��ZЖ<=駐��&l;�Mu%پo|or����<�]N�u�סęE���^�y�����x`�c�z;�+*�4�+�--^	E`/F�H�-�����6�P�~n|�<�S���JIj^aȋ )�Z)c��Rx-���Fz�ԁ�D��?N+gm���P���5vB��}d�j��FǧhF�N3_Q�����D)v݋JÜʮ�؞@o���
?�u�cv@�;w���nI�|Z`�T�TL˱+��q2���$��6�a�j��p�c�A\�o�&3{O~�/l�K���f,�=_7�[P9qo�ZOk���-�V�н��	�� ���<��~N��3���4XJ��u��7�n�
�و�@��2�����o'�?LM-�U�6���ڋ??^U���I�8��c�i�J<DOՅ:�V�\��r_7��}�z���Zן�f��sw�����3�$Uw����Gy��>�U���X3������$��E2J$K�S�ܖo���m�L���5�D�\�b#�����t�օa��\�~d�T?��5����LD?�`�}tF6����	Ж-�'�	4MrA=���U8Uoh��G��v��m��<�"����@��OU�-N]j�4Ai P���B,[����l�E��g�U��[ke�����`�9�se�c��q7Ecٛ�|�����f&y��[-~�����gE	Ԥ�c�ax��z\��7������{摝����� �!w:#��?[�"C�JK7zϼ��t0s�Q�@�!�q�b�E����ܻ����g�C[>	�ZO'C�r
�s
1��]ǽ<������HE|9u\��Z[|c��`��.yt�vc�������4�&8�(_��.��Ӱ�ԩ�R��0��q�a� ����b��\yq:��gOq�ֳze0t�q?�=��x���d�A���3~�����e��K�N���8z2%��t3��>�rW1i���Wq�I�7�?9y���c����
�4V2�Lc���@���2��s�\ݤ�¿�!�
�כS^G|���Ry笄�K~ѥ���q,m���N�g1�ҒoE�RHeml�\�2�v¦�� ��^R���p��d@MoS�+�>T6� �Θ��SX���t��4 Y�K��P�;�6�KQ��X>��(g����97�����y�*�D=�XR7�^(φ�s,��B'�2�"�?�!R�5U$�W���-�2��V�A4γ���rE,�%ڳp�;���kB�b1�Q�!Y,OY�\�\���L��ܝ$opwX��q���1Goh��cn�>�	i�m�4�܄#��߈d��ha��V-���r���y��]tЧV�+?��M ��֐\,6:���2jk���)�&�?��R��ӱ.hI�+k�{)���-�Ԗ�Ĵf��˻�t�L	����<��Z
����	l;K�|�[��br��ӯz]��;�p4�z6۔�(G�Y<i��%�U�߅���&��?��NiYJ���Cz�:�T�f~"j�K�=�5b&W�xE�r�/F6��r6�����rk���<�c�X@���a0$���8�o�9,ڃ���e�Ƕ� ���a1�Y��H�{�5�kx6�b�5����5#�E��DG��c�%��lB��5K�0�wZǨ-̓z�/"_lGBϦ� @Xk�U=<n�/�E�Rk`*&�t������(b��h�
e�nO��.���ܼ��"G�j�U�q>��ٳ@2�TT�r�́)V���c��(ʿ��(�؇Ax�����e�ʧ���N��M�OgO�t5@�����}O��Qv����&ѨC(jx�����&.b�j�Ç=?�V ۿ^x �����$�b*^�Q>*�V���KBj�����Z��a��q��%�}���C!�+���������} �u�D�Fu�G1�A���h;�H��/x�(T�#�U�!��%D���<lb���� �n�"zU��u�an���}�|�v_ߴ�.Ǻ��i���~f�^E5�z�������?Lð�?�U�'y�h���U{W��������h;��ZI�qGh����|�QB�<�w+N�	�����);��W���v�[�g��5�G�|"������M�s���H#ԗ�^�O!0v/�8�KK/�Ke��K�^O��-U��|��[O�P*⪍lUn4xlpY�����i��c����7��q��F+��Hն����[U8Z�"d�\�eH�$ͮsQ%	{~D�nV�T,:t�Q�"N+��OS��9�S���끾N�*ဥ��<�����R�N��Ԟ#۷Q�.9zbw�[F�(�O�Om_�F�P��t�1�Y�)1H���.?�Ů�L����t�wg�V�/Ѭ���JX�8P���c�v*Ή- +�������$��_d��|{�j� ��g�d1�솞���G�ѝ����x�^	3�| �Hb������������ �@tZ��>|�70;j~²�K�)��%�tr?�B�Mɤ�E��lP��C�Ϛ�7ʮ�?D���w�[������$� D7iHYIYdQ!eiX]N'epcbe.<=h!;<ugh'ki)vkev.