MZ�      ��  @      @                                   �   � �	�!�L�!This program cannot be run in DOS mode.
$        PE  L ?��G        �  C                         @                      0     �N                                                                                                                                                       .flat                                �                                                                                                U����    [����  P�i  ��'  }�1���'  P�  ��t�ǃ�GP��'  ����U����    [��R���  ��+  P�y   ���  P�  �P4�U�PP�U��ƋV(U�U��u���  �u��u��  ��t>����  �}�+  �h �  ��'  S�u����  P�u��  �u��J  ��  U��`�U�M�3�/  �BI�σ���t��a��    ��[�,�&ɠ���SXu��4�e4�           z��VU���`�u�C   	�t(�Ht;Mr �@x�U��ЋM	�t�P�� 	�tE�� 1�d�I0V�I�q��@^�U���`1��E��E���MZ  u@<���PE  u�E�a�E��� U���`1��E��E�}j@h 0  WP��  ��t�E�a�E��� U��`�u������t(���J�Bt�Rx���Q�z}�ru�J��(Y��a�� U���`�E�Pj�u�����	�ta�Ƌ~	�tX}VW��  ��tC�ǋ	�u�VU�vu���t)��s%��  �E��RPW��  Z��������^���a�� U���`1��E�����hu��4P�K   �E��}���<.u���)���    )ĉ���PW��DLL �U�Y	�t̖P��   PV�   �E�a�E��� U���`1��E��}�U�RPW�����ƋH�F �1҉ǋEP�   ;Et��B���1�}�F$��P� �N���� ��E�9�ru�9�w	P�+����E�a�E��� U��`������ǋu��	�t(�6��  �ǃ�����	�t	PW�R����������a�� U���`1�@�}�	�t����5��B8G��E�a�E���     7�����T����5�X�5@|}g4df{sfuy4wuzz{`4vq4faz4}z4P[G4y{pq:0DQX���S�#4T�vDdT�d�ADL$T��ADL%4DT�ADL&dT�&:$$ADL5=D�&\q�r�U�4:2�����%�T�X0�U`�P0�@0����c��GBCD~�|Tp�!��ɭ�14�L;d���`4/`k���00`� b��@\h�a�c���@���p�!��KJO�A��HA~���z|�N�a�	�I��I��o���4��7�I�Q��$1�	���)��T����Q�	�����Q���W�g%o��;�ɐ�6�b��`iBA�:��������$;�A� V�j{��,dE�  )(!�m���)M��ZO�jcIJ��`<l xG��b�&�9tBm�`k����W$1 ��	���:n�e�~�9���b�tj~W
(v�g�a5��֑�/�3��>D�0��ߒ
0�<��WI�)8*������f��L�p����M|#�|��D���8��q�D�(0r�0���8w�<:04j�x�)	�� 0�s�\ ��%ݝY�D�;����p�w�4p�T$B�
��d�J on맩���7��:�i�h���~P�i�C\[��-�x��:9� �7��(*��V�9�F�e"���_�%���A��y�=��O�y�>��u��^U�˖�!-h�6D݂��O���$RG�5�����럅�����c(����T��wkl 䂅�yh����/xT4&�ӑ��y/�`C�7�=��`�{�(����/Q/p��"�^0�KM� �Du4ϫ4�(jN�������--���H���U"瓞���{X�$��+a�*��)����Ʌ:aSӐ)�PXX�b	���1C�#�<�����6�`
BÝ�n�L�:�V��`�7��� �c��_-»���y�g�O�K_
�����ci�/()�'g�����p�� � ���g?���;	������xwW���W�#��ϱ���4p-h����8��h�� |����{ED����`@� �!�y�Q�� ъ*��	:���/`'$r��a�e�C-�f�×!�����M�?���Hl�����3�D䭧y��C@�x7�9�2��\�r�	�m.jCx` ��$�0�r�FC1<I�O��� ้��/8��r�O��������k9���c�8���ߢ��Xf���^��~��`AK��5��8��L7>�����l��Kv�R�J{�b�z�nD%�J�qy̗�-������% ��#�Sb�8�-)�ȗ��uCE`�M��$n��U���2ia|�/`٢�G����	�xrм$��j�p`	E�arX�a�/�a����)8��Kn,��[������r���ҕ�|���{�,R�2��
��-�["�
�,��Y�:��9���G
H㢧a��a��< �7�����k����b<h~�	���"�~�H��L�-=�Co�gI�$��#��zѡ�tW"ց}�D?ûV;�U.�C��_Ґ�6�c�W$J��^0m����&T�,z�i�)�>��\�l���X��Lc��
��S�h���r�/$��zҝ�K�9u.IA֝ ��s\-s`�,����`�T�b85 �](��k��-�`�	���=�-�`��MxԦ��<@����a �3^�?���Xw���h��a�h٬T�.�:uN:Mߘ��6�2��Cr�
������8)�x�����w"'��D\�$����¦���H����(��Ł�'D,������-�I�S$D�'�!t"6.?����i��\�ݤ�	�-��J�j�W�X`�B�#!�(|iJ���UxF?�1#��ut�$L"T���^'~S��������-�p ��H���9�������}���[�����x6>M/D��rC�OR�p��J\�f@<@��a�Ht�0��0�8��+씋�!�=��bb{C|���
,u��|`Q� b�]U`�>� �a�
�u��X�c�Lpu��T�P�"�2ם�����p��6�����*���)v$Ckh�G3/j:��p��|��p
��	��}џx�+i}�4!(������Cr��\|�4���m1�#M(�?�����>��ςro�hiH2]���xtǏ0aJ���F;�d�>�\O̫�h*�:/���ѯ��xr)�|��z�ʗ1�hrg�	!��hO�.	}t&C,tb�2$� l<ML�Oqtb��#L�W9M%"@�=�t/φt2j_�� )�B:�DN��ML�=�q�3t��3�T��(��Ml��	|���Ws��=�k��bj�T�a��p,��5S�&y��=x�����a$t�j$T6@fM	)s�řR/����q&�:St��5���
��Ԧ����f f��O��wg��l5�E`0�ti���3x�#��g�����;���|�@�M[�x��<��)�4Ɣ�R+�Ha<�a�y�O�B��=��2Sq�>��p���7x��RN���<�/(����X�Cd�COpo a�(Ė]ģ_8�B�r�r/i�9�Κ��43[������	B�h%:���9��@��W<�Hb�$����M���0&�E��JL�1��o��|4��3���T7!�.���8�6a��Ez��$�F��%X~�W��wH�$]�3���J��:��;V)U� I��X��kՆq'-����$';.�\�|o�M|i"�q�Q��A����,R2�_l5|l=��,!RT��ђ�8mf��-�����2qv���r���5�1�c��nS&f����.L�\��5�<�����1�1B�I��_?�I��U��(̆�����ru�0lL�&���<�)J�\���Uo|�
�4e+ow�0�=`!|g��7�\8�V�|zP+�?�0hࠇ$Xh�o�������d�&BL��0,�j��e�v�O�Ж�`�>(hu�1\�c������:�a�Ô7�?l���h6��yi,ͫ����ç�QK|>���y��
2��T��\���p��u���]�T��f��GP�ȴ-(Cz���ܻ�a<|n��b��_�75_��Ҵ�����[5��������
���-܍og����,�܁�f
��)o���;�����l4`Yommm:`\8`W$h-j-���3c`9C`<D`7d`����
@``` 9`T9b���ce&v�i�-ch��	�7�GpJ�\��
`��z�ӳ	"a�IB���gY��5[������#A�aS�Q[l�)>v�CR�n�b���M��|�x^��f�{ d��D�P��w��� O���O. & e4��|0����o�d��59��\f������������f�)��Nc���N�p��q���# ~���$OP��$���p,:�L]b���	�����`��ڑ�`���͘����%��	��V��/&f�܈��"�C�m4��sx"�VJ�����u��8��� �}��6+g�{.(������c����g� 0���00�h0r���#��r��x�(0�H��xLSM��kϣ9�)g�=���	NoW{�1�TO&4����&4����x&4���E7���|~:�?��8��H@&�k� Y����E����������}w��Oz(\�-@<P��-�W+�3�PR���M��^��gk�[3�[���2������Jfx����T%:��$�#��|Τ�03(������S�)�˒��|6hLue��o�	-,��������0��^l�Vh��;*��C;0	�;$��h	1�	;6��{�";5	g���j; ���1�����7�*S'r<N�$��Ͳ���f��Hd�CE�6�4�����Ldw,���ߩ� 1 %t��|c�*�+l�����(]���� �$J���h�� ���0�$� I���8��Y� Y�� �� I�`����� YǬ����Y� Y����P\`�� TX�G���J��ԛUPBUD]'&:⌯ WF@FUG��
K.;;�����57#����D-7F.F!7'M7*7'OMDO13D4=-.g�k�TUg�{�.9$I%�}�5bmj_^^STV��H�WVVgW_SfL^*/W8T&DU͹�VP_UurTS�d�{g'�'l?�y�c!_(~W�p�xS�/
Eu�H��T;�$upgx��_Y�G�}gpzy{pqy�>�I ��U�UA��k6-��PiLUa�q;�T�k�"Y�<$,U;���TT�V�� z��K"L�$F`x�[��Azc}zpq�KKSq`Yuwk� Ufsgql}`yqywdmgk���q`fu}.g}szux�km�DQX���S���4/�#4��8�$jxbr
�D"�'�
 ]$_��D,:`<�zuw�
�7�$"��t:pu`u��0�yLL]�:}<�'"��83td�O0�t�DT������C�����������R�S�a�
����f���a�
������g�a�
����g�%ݗ�f���R���``���a�
������a�
�����a4U�a�
������g�a�
����g��������� ;���b�V�S]a��w��넟�������c���X���J��L�S8�(c�+a��Kr������=���������͙�T��`(�K��$t�D���(t��S�`ȝ�C\�A�Tt�`������\t��Pt�����D@~GC������4k�t<kLD@DGC��Lu�P0�~-�a����͹��Ld(dqdDdddjd�d�d�d_QFZQX'&:PXXWF@PXX:PXXX{upX}vfufmUSq`Df{wUppfqggB}f`auxDf{`qw`Ql}`Df{wqggql}`44$$n�V                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                           