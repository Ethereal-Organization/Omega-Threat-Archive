MZP      ��  �       @                                     � �	�!�L�!��This program must be run under Win32
$7                                                                                                                                        PE  L ^B*        � �� �         ��      �    @                      0                                  �    �  `                          �	                                                                                  CODE    �      �                    `DATA    �    �      �              @  �BSS     �   �       �                 �.idata  `   �      �              @  �.edata  �          �              @  P.reloc  �	     
   �              @  P.rsrc             �              @  P                                                                                                                                                                                                                                                �%��@ ���%��@ ���%��@ ���%��@ ���%��@ ���%��@ ���% �@ ���%��@ ���%��@ ���%��@ ���%��@ ���%��@ ���%��@ ���%�@ ���%�@ ���%�@ ���%�@ ���%�@ ���%��@ ���%��@ ��S�ļ�
   T�����D$,t�\$0�Ã�D[Ë��%��@ ���%��@ ���%��@ ���%��@ ���%��@ ���%��@ ���%��@ ���%��@ ��SV���@ �> u:hD  j �����ȅ�u3�^[á��@ ����@ 3ҋ���D����B��du���^[Ð� �@Ë�SV���������u3�^[Ë�P�V�P���X�B��^[ËP��
�Q���@ ����@ �SVWUQ��$��] �$���P�V�;��SS;�u�������C��CF�F;Cu�������CF��;�uË֋��V�����u3��Z]_^[�SVWU����؋��2�C;�rp��J��k;�wb;�u�BC�B)C�{ uH���9����?�΋zϋ�k;�u){�*�
J�$�{{+��|$+��s�ԋ��������u3�����;�u�3�YZ]_^[ÐSVW�ڋ���   }�   �����  ��  ���sjh    Vj ��������;��t#�Ӹ��@ �l�����uh �  j �P�����3��_^[ÐSVWU�ً���C   jh    h   U�������;��u����  ��  ���sjh    VU������; t#�Ӹ��@ �������uh �  j �P�b���3��]_^[ÐSVWU���L$�$�D$����3҉T$��$ŉD$���@ �Q�;�s;�wF��C;D$w;;t$s�t$��C;D$v�D$h �  j V�������u
���@    �������߁���@ u��D$3҉�|$ t�D$�T$��D$+D$�T$�B��]_^[�SVWU���L$�$�Ћ�� ���$���  �� ����T$�D$�(�D$+ŋT$�B�5��@ �<�^�~�;�v��;|$v�|$;�vjh   +�WS�&�����u
�D$3҉�
�6����@ u���]_^[Ë�SVWUQ�؋���  �� ����4$���� ����$���+$�A�5��@ �8�^�~�;$s�$;�s��;�vh @  +�WS������u
���@    �6����@ u�Z]_^[Í@ SVWU���������@ ���?  �� ����] �3;{,�΋׋C�����> tP�FC�F)C�{ u>��������5�;�uɋ֋�������> t!�̋֋�������<$ u��̋V�����3��YZ]_^[Ë�SVWU���$������@ ���?  �� ����] ��;�t;su�;suW;{��   �L$��+S�CC������|$ t3�L$�T$���]����|$ u��L$�T$�D$�%����$3҉�   �L$�׋������|$ t4�L$�T$�������|$ �f����L$�T$�D$������$3҉�H�k;�u:;{5�$�׋��q����$�8 t(�$�@C�$�@)C�{ u��������$3҉��]_^[ÐSVW�����$���?  �� ����4$��� ���;�s[�ϋ�+Ӌ������L$�׸��@ �]����\$��t�L$�T$���&����D$�D$�D$�D$�|$ t�T$���@ �����3����_^[�U��3�UhF@ d�2d�"h��@ �9����=5�@  t
h��@ �.������@ �������@ ������@ �x���h�  j �������@ �=�@  t/�   ��@ 3ɉL��@=  u���@ �@� � �@ ���@ 3�ZYYd�hM@ �=5�@  t
h��@ �������  �堬�@ ]�U��S�=��@  ��   3�Uh*@ d�2d�"�=5�@  t
h��@ �f������@  ��@ P�4���3���@ ���@ �h �  j �CP�%��������@ u���@ �������@ ������@ �u������@ ��t����@ P��������@ ��u�3�ZYYd�h1@ �=5�@  t
h��@ �����h��@ ��������  ��[]�S; �@ u	�P� �@ �P�H��   8;�u��y������@ 3҉T���$��y������@ �T�� ��P[Ë ��P[Í@ ��@ ��J;�rJ;�r����@ u����@    3ҋ�ÐS�ʃ����|�  ����  [Ã�|�ʁ�  ���[����@ �Ѓ�����������@ ��  Ë���|����������Ã�|
�ʁ�  �� ��SV�Ѓ���ʁ�  ���  �t
���@    �ځ����+Ë�3������t
���@    �t �Ѓ��r+�;pt
���@    ����ދ�^[Í@ SVW��3���   �t%����؋�u����X����F�؃#���_^[�SVWU�������$ �������؅���   �k��C�Ѝ7+у���+���+Ń�}�L$��+S׋��������L$�׃��F�����l$��t4��+֋��c�����D$�SS;�s
�7+������T$�������$�$��]_^[Í@ SVW����߉s��ƃ��p��   7�օ�y������@ �D���u��@ �\��[��:��C���Z�,�� <  |�֋��������u� �@ � �@ ��C���Z_^[Í@ �=�@  ~@�=�@ }���@    �+��@ ����@ ���@ ������3���@ 3���@ Ë�SVW������<$���������L$�׸�@ �����\$��u3��R�;�s
����)G�G��t$;�s�����G�G;�u���   ������o���@ �G��@ ���_^[Í@ S����؋ԍC�D����<$ t���W�����u3���YZ[ÐSV�����؋̍V�������<$ t���&�����u3���YZ^[Í@ 3҅�y����=   ��@ �T���u@=  u���SVWU�� �@ ��@ ���@ ;s��   ��C;�~{�s�[;s���B;t��c��   �������؅�uN��������u3��   ;u �)u �} }u 3��E ��@ 5�@ �փ�������@ ��5��@ �L�������S��+ƃ�|��֒�T������;u�C���ƃ ��Ëփ�������@ ��5��@ ]_^[�U����SVW�؀=��@  u	�������t�����~
3��E��T  3�Uh�@ d�1d�!�=5�@  t
h��@ � ����������}�   ��   ��   �Å�y������@ �T���ty���Ã ��B;�u�Å�y������@ 3��|���&�˅�y�����=�@ �D��
�M��M��A�M���ƋR������E����@ ����@ �V  �   ;�@ J)�@ �=�@ }�@ 3���@ ��@ �@ �Ӄ�����E����@ ����@ �  �2�������E�3�ZYYd�h�@ �=5�@  t
h��@ �������
  ��E�_^[YY]Í@ U��QSVW��3����@ �=��@  u�f�����u���@    �E�   �a  3�Uh�!@ d�1d�!�=5�@  t
h��@ ����������u���@ 	   ��   ���@ ��%�����)��@ ��tE�ƃ��P��|��  �t���@ 
   �   ��+�;Pt���@ 
   �   ڋ��T����������Ë�;=�@ u,)�@ �@ �=�@  <  ~����3��E��	  �   ���t�������}���@    �7��)�ǃx t�8 t�x}���@    ��P�������Ӌ��'������@ �E�3�ZYYd�h�!@ �=5�@  t
h��@ �W�����m  ��E�_^[Y]Ë�SVWU�����������}�   ����} �������ǋ�;�u��  ;���   ��+։$;�@ u8�$)�@ �$�@ �=�@ �L  �$�@ �$)�@ ���3  ���u�ËP$������<$|��ދ$����Ã�������   ����   ��+ǉD$;�@ ug��@ ;D$|S�D$)�@ �D$�@ �=�@ }��@ �@ 5�@ 3���@ ��+���@ �E %  ���u ��   �>�������uM�ӋH�$�$;L$}$�ڋ$)D$�,�����D$)$�<$|��Ƌ$�n����:4$��ރ#��.��   �t!%���Ë؋T$���������t	�������3����+���@ �E %  ���u �YZ]_^[Ë�U��QSVW��؀=��@  u�������u
3��E��   3�Uh=$@ d�2d�"�=5�@  t
h��@ �����֋��������t�]��6���������Ã�� %�����;�}�ƅ�t�׋ˑ�B  ��������}�3�ZYYd�hD$@ �=5�@  t
h��@ �������  ��E�_^[Y]Í@ S��~�$�@ �؅�u���   �3ۋ�[�S��t�(�@ �؅�t��   �3ۋ�[Ë��t2��tP���,�@ Y	�t�ð�   ����(�@ 	�u�ð�p   ��tP���$�@ Y	�t�Í@ ��@ ��
  �SV��؀��=�@  t
�֋���@ ��u�?  ��   ���w
3��Ê�0�@ 3��Ë�����^[Ë����$�����S���  ��   [�VW�Ɖ׉�9�wt/��x*�����_^Ít1��|9���x�����������_^�SV��3�f�Cf=��r/f=��w)f%��f=��u���S����u���S$����t���s������8�@ t
�g   �_�����^[Ë�W�ǈ͉���f�ȉ���x	�у��_ÐSVW��P��tl1�1ۿ����F�� t�� ��-tb��+t_��$t_��xtZ��XtU��0u�F��xtH��XtC��t ���t-��0��	w%9�w!���؊F��u���t	��}T�	F���~KxI[)��G�ŊF뜿����F��t߀�ar�� ��0��	v����wЀ�
9�w���؊F��u���u��Y1��2_^[Í@ �%��@ ��S3�j �������uj�����% �  =   t=   u���[ÐU������@ �E��E�Pjj h�'@ h  ��1�����uM3�Uh�'@ d�0d� �E�   �E�P�E�Pj j h�'@ �E�P����3�ZYYd�h�'@ �E�P�������  ��f��@ f%��f�U�f��?f�f��@ ��]� SOFTWARE\Borland\Delphi\RTL FPUMaskValue    ���-�@ Ë���t���Q�À=�@ vj j j h�����@ Ð�=�@  tPPRTjj h�����@ ��XÍ@ Tjj h�����@ ��XÍ@ �=�@ vPS�����Í@ ��t�A�9�t�9�u��AA����Ë��=�@ vPRQ�����QTjj h�����@ YYZXÐ�=�@ vRTjj h�����@ Z�PR�=�@ vTjj h�����@ ZXË��D$�@   �  �8����P�Htn��������@ ����   �҅���   �T$�L$�9���t7������=�@  v)�=�@  w �L$PQ������� X��   �D$�H�0�D$�H�=�@ v�=�@  wP�D$RQP������ YZXtp�HS1�VWUd�SPRQ�T$(j Ph�)@ R��@ �|$(�  ��    ��    �o�_�G�)@ ���f������#   �^  ��    ���    �A������   Ë��D$�T$�@   t�J�B@*@ SVWU�j���F�����]_^[�   Ë��D$0�@�*@ ��  ��    �
��    �B�`��8���t�B�k����r���1���d�Y��]_^[�   Í@ �  ��    �
��    �B�1���Z�d$,1�Yd�X]��������1ҋL$�D$��d���� Ë�U��U�=�  �,t\=�  �tW-  �t\-�   t=HtN�`q��?��r6t0�R=�  �t=-�  �t.HtHt$�:-�  �t/��=t&�,���*���&���"������������������
��������%�   �R�`���]� �D$�@   ��   �=�@  w�D$P�p����� tq�D$��%����T$j Ph�+@ R��@ �\$�;����S�Ct��@ ����������҅�������S�������@ ��t�ыL$��   �Q�$��  1�Í@ 1ҍE�d�
d���@�+@ �h�$�@ Í@ 1ҡ$�@ ��td�
9�u� d�Ë	���t9u�� ��U��SVW� �@ �G��tH�_�p3�Uh�,@ d�2d�"��~K�_�D���t�Ѕ��3�ZYYd���-����������������_^[]ÐU��SVW�(�@ ��tK�03ۋx3�Uh-@ d�2d�";�~��C�,�@ ��t��;��3�ZYYd��������P����'����v���_^[]ÐQVW� �@ �}Ĺ   �@�@ �<�@ �-4�@ �8�@ �(�@ �0�@ �Mĉ �@ 1Ƀ} u��,�@ �@ ��@ �@ ��@ �����E@�H�@ HY��D�@ t<}��Q�L$��t�E�U��Y�E<|���=�@  u�$�@ �=�@ �EH�!  ������ �SVW�T�@ �� �@ �ÿ
   �����03�����û
   �����I��u۱��@ �Ѓ���t�@ 3ۊو��I��u�_^[Ë�1�� �@ ���@� �@ �_�o�w�w �7�   �_^�� Ë�Q�=4�@  tWf�=�@ ��u�=�@  v��@ � �@ j �D$PjhT�@ j��B���P�\���j �D$Pjh/@ j��'���P�A���ZÀ=�@  uj hL�@ hT�@ j �3���Z� ����   
  SVWU� �@ � �@ �0�@ �{( u�? t���3҉���Ճ? u�=�@  t�����2���3���@ �{(u
�> u3��C�����{(v�> t!�C��t��  �S�B;Bt
��tP���������{(u�S$�{( t�����; u�=�@  t��@ �P�]����V�����   �^�v���]_^[ã �@ ����Ð��@ �����Ë��t�     �J�I|��J�u
P�B��S���XÐSV�É֋��t�    �J�I|��J�u�B��*�����Nu�^[Ð��t$�J�APR�B��\   ��XR�H������ZX���B����t�J�I|��J�u�B������Ð��t
�J�A~��B����t�J�I|��J�u�B�����Í@ ��~$P��
���P����Zf�D�  ��Z�P��@�   �1�ÐSVW�É։ω���������ǅ�t	���G�����������;_^[Ë�U��RP�EPQj ���@ P�-���]� �R��   ����ZÐ1Ʌ�t!R:
t:Jt:Jt:Jt����BBB��Z)��x���Í@ WPQ��1��u��X�X_�]���Å�t�@�Å�t?��������SVW�É֋y��V��9�t�V  ���N�������_^[��?  �����Å�ta���h���;t\;tPQ�Y���ZX����SVW�Ӊ�P�C�F������ǉ؋K��5��������N�S��&���X����t�O�����_^[É��������I����SVWRP��1��L���t9u�ϋA�J�1��L���t	A�9�u1�Ju��t�$�w��  �<$�77K�����P�ƋD����t
�H������Ku�ZX��u��t�J�����Z_^[X�$���Ë�SVW�Ɖ�9���   ��th��tk�F��W�)�w�R��t&��9�uXJt�N�_9�uK����Ju������Z��t"��8�uAJt8�u:Jt��  � ��  � 9�u'��#�W�)���F�)��Z8�u8�u����8�u8�_^[Ë���t
�P�B~��@�Ð��t� ��3@ Ë��t8�J�It2S�ËB�������P�H�����X�H�I|��H�u�@������[��Í@ ����Ë�S��t-�X���t&J|9�})Ӆ�|9�D$������1������D$�����[� �SVW�É։��������t0�J�N|*9�}&��~")�9�~��)���������؋R�)��   _^[Å�tVSVWU�É։ϋR��t�R�O}1�9�~�׋k�����u   X9�u���/�H�)��������؋�������]_^[Ð��t@��t1SVW�Ɖ׋O�W�V�Jx�F)�~�u��VW���_^t����Z1��1��Z��)�_^[Í@ SVW�É�1���~H���t#�x�u����	P���U���X����p�� �(���o����ǋ��t���H�9�|��������������;_^[Ë������Å�tPj ������������Í@ ���tR�����Í@ ���t�     PR�����XÍ@ SVWU�����P�����$����	��������]�n���  }(V�D$�L$��  �����؅�~�T$�ǋ��9   �*�݋ǋ��l   V��L$��������؅�}3ۋǋ��M   ��  ]_^[Ë����T���PQR�$���������Z�2�����Ð1Ʌ�t�J��B���Ð��t�@���Ë�SVW���3ۅ�~'��������؋�������~;�}�Ƌ�ɋӋ�����ǋ������_^[Í@ ��a����U����SVW�E�� �@ �E��}� t93�Uh7@ d�0d� �]��E��S3�ZYYd��
����������E�� �E��}� u�_^[YY]Ë���@ ���@ Ë�U��Q�E�3�Uh�7@ d�2d�"�E��@�t���3�ZYYd�h�7@ �E�;�@ u�E�� ��@ ���@ ��t�;U�u	�U����� ��u���c�����Y]Ë�U����S3҉U�3�Uh8@ d�2d�"j�U�Rh  P�i����E��U��   �����E��U������؃}� t3�3�ZYYd�h!8@ �E����������������[��]�U��3�Uhr8@ d�0d� ���@ u#�8�@ �I�����@ �?������@ �5��������3�ZYYd�hy8@ �������]Ð�-��@ ��   ��@ ��@ @ ��@ @ �6�@ � �@ �6@ �.�����t�U�������f�<�@ ��f��@ ��f���@ ���X����,�@ �����(�@ ����%   �=   �t-����%�   f��v���@    � �/����������@ ������u������@ �G���� �@ Ð�%8�@ ���%4�@ ���%0�@ ���%,�@ ���%(�@ ���%$�@ ��Pj@�����Í@ �   Ë�S������؅�t6�=��@ �u
��   �=������������u��   �(����P���@ P����[ø   ��t�z������@ �������@ P�u����\�@ Í@ �   ��t�=��@ �t���@ P�O�����tP�-���ø   ��t������=��@ �t���@ P����Ð�L�@ ���@ ��u&d�,   ����%������@ P�������tá\�@ �P�������t�ø��@ ����Ð���@ �}u*PR�L�@ �M�P�@ �J�B    �B    �����ZX�5T�@ ���@ �K���Ë�U��3�Uh	;@ d�0d� �X�@ 3�ZYYd�h;@ �������]Ë��-X�@ �U��3�UhA;@ d�0d� �`�@ 3�ZYYd�hH;@ ��������]Ë��-`�@ ��%d�@ ���%`�@ ���%\�@ ���%X�@ ���%T�@ ���%P�@ ���%L�@ ���%H�@ ���%D�@ ���%@�@ ���%��@ ���%��@ ���%��@ ���%��@ ���%��@ ���%��@ ���%��@ ���%��@ ���%��@ ���%��@ ���%��@ ���%��@ ���%��@ ���%��@ ���%|�@ ���%x�@ ���%t�@ ���%p�@ ���%l�@ ��3������U��3�Uhi<@ d�0d� �d�@ 3�ZYYd�hp<@ �������]Ë��-d�@ �SV��؋Ƌ�����^[Ë�WV�Ɖ׹����2���щ��։ʉ����у��^_�SVWU������������   �C;�|�|� v�;�}
�������N�|7� v�U��+�A�Ӌ������]_^[Í@ SVW�������z����؋ǋ�������֋7��t�<ar<zw, �BFK��u�_^[Ë�U��j SVW��3�Uh�=@ d�2d�"�؋�������t3�ù
   ������ù
   ����؍E��W0�����U�����D�����u�3�ZYYd�h�=@ �E��K�����Y�����_^[Y]Ð��l����$�   T�����|$���Ĕ   Ë�U��3�QQQQQQQSV���3�Uh�@@ d�0d� ��������)rH��)r��E���@@ �o�����E���@@ �`�����	�����)rH��)rH��)r �+�E�� A@ �9�����E��A@ �*�����E�� A@ �����������)rH��)rH��)r&H��)r/�:�E��0A@ ������+�E��@A@ �������E��PA@ �������E��`A@ �������=6  }H�����)r&H��)r/H��)r8�p������)r;H��)rDH��)rM�X�E�pA@ �{����I�E�A@ �l����:�E�A@ �]����+�E�A@ �N�����E�A@ �?�����E��A@ �0�����6  }"��s�����*r6K��)r?K��)rHK��)rQ�   ��������)rPK��)rYK��)rbK��)rk�v�E��A@ ������g�E��A@ ������X�E��A@ �����I�E� B@ �����:�E�B@ �����+�E� B@ ������E�0B@ ������E�@B@ �q����u��u��u��u��u�E�   �����E�P�E��E����й   �E������E�PB@ �u���u�E������ЍE�   �����}� u�ƺ\B@ �����hpB@ �u�h|B@ �ƺ   ����3�ZYYd�h�@@ �E�   �Y�����C�����^[��]�   ����   1/2,    ����   2/2,    ����   1/3,    ����   2/3,    ����   3/3,    ����   1/4,    ����   2/4,    ����   3/4,    ����   4/4,    ����   1/6,    ����   2/6,    ����   3/6,    ����   4/6,    ����   5/6,    ����   6/6,    ����   1/8,    ����   2/8,    ����   3/8,    ����   4/8,    ����   5/8,    ����   6/8,    ����   7/8,    ����   8/8,    ����   ,   ����   ��δ֪��    ����   ��  ����   ��  U��QSV��ډE��E������3�UhF�@ d�0d� �E��\�@ �,���t�E��p�@ �����  ���   ~���   }�ƺ��@ �o����J=  ���   ~���   }�ƺ��@ �N����)=  ���   ~��  }�ƺ��@ �-����=  ��  ~��5  }�ƺȀ@ ������<  ��5  ~��_  }�ƺ܀@ �������<  ��_  ~���  }�ƺ��@ ������<  ���  ~���  }�ƺ�@ �����<  ���  ~���  }�ƺ�@ �����c<  �ƺ,�@ �w����R<  �E��<�@ �����t�E��P�@ ������  ���   ~���   }�ƺ��@ �4����<  ���   ~���   }�ƺ��@ ������;  ���   ~��  }�ƺ��@ �������;  ��  ~��5  }�ƺl�@ ������;  ��5  ~��_  }�ƺ��@ �����;  ��_  ~���  }�ƺ��@ �����j;  ���  ~���  }�ƺ��@ �n����I;  ���  ~���  }�ƺ��@ �M����(;  �ƺ,�@ �<����;  �E��ԁ@ ����t"�E���@ ����t�E���@ �����  ���   ~���   }�ƺ �@ �������:  ���   ~���   }�ƺ4�@ ������:  ���   ~��  }�ƺH�@ �����:  ��  ~��5  }�ƺ\�@ �����b:  ��5  ~��_  }�ƺp�@ �f����A:  ��_  ~���  }�ƺl�@ �E���� :  ���  ~���  }�ƺ��@ �$�����9  ���  ~���  }�ƺ��@ ������9  �ƺ,�@ �������9  �E����@ �l���t�E��Ђ@ �]����  ���   ~���   }�ƺ�@ �����9  ���   ~���   }�ƺ �@ �����i9  ���   ~��  }�ƺ�@ �m����H9  ��  ~��5  }�ƺ(�@ �L����'9  ��5  ~��_  }�ƺ<�@ �+����9  ��_  ~���  }�ƺT�@ �
�����8  ���  ~���  }�ƺl�@ �������8  ���  ~���  }�ƺ��@ ������8  �ƺ,�@ �����8  �E����@ �1���t�E����@ �"����  ���   ~���   }�ƺЃ@ �t����O8  ���   ~���   }�ƺ�@ �S����.8  ���   ~��  }�ƺ��@ �2����8  ��  ~��5  }�ƺ�@ ������7  ��5  ~��_  }�ƺ �@ �������7  ��_  ~���  }�ƺ8�@ ������7  ���  ~���  }�ƺP�@ �����7  ���  ~���  }�ƺh�@ �����h7  �ƺ,�@ �|����W7  �E����@ ������  ���   ~���   }�ƺ��@ �H����#7  ���   ~���   }�ƺ��@ �'����7  ���   ~��  }�ƺ��@ ������6  ��  ~��5  }�ƺЄ@ �������6  ��5  ~��_  }�ƺ�@ ������6  ��_  ~���  }�ƺ��@ �����~6  ���  ~���  }�ƺ�@ �����]6  ���  ~���  }�ƺ,�@ �a����<6  �ƺ,�@ �P����+6  �E��D�@ ������  ���   ~���   }�ƺX�@ ������5  ���   ~���   }�ƺl�@ �������5  ���   ~��  }�ƺ��@ ������5  ��  ~��5  }�ƺ��@ �����5  ��5  ~��_  }�ƺ��@ �����s5  ��_  ~���  }�ƺ��@ �w����R5  ���  ~���  }�ƺ؅@ �V����15  ���  ~���  }�ƺ��@ �5����5  �ƺ,�@ �$�����4  �E���@ �����  ���   ~���   }�ƺ �@ �������4  ���   ~���   }�ƺ4�@ ������4  ���   ~��  }�ƺH�@ �����4  ��  ~��5  }�ƺ\�@ �����h4  ��5  ~��_  }�ƺp�@ �l����G4  ��_  ~���  }�ƺ��@ �K����&4  ���  ~���  }�ƺ��@ �*����4  ���  ~���  }�ƺ��@ �	�����3  �ƺ,�@ �������3  �E����@ �r����  ���   ~���   }�ƺ؆@ ������3  ���   ~���   }�ƺ�@ �����~3  ���   ~��  }�ƺ �@ �����]3  ��  ~��5  }�ƺ�@ �a����<3  ��5  ~��_  }�ƺ(�@ �@����3  ��_  ~���  }�ƺ@�@ ������2  ���  ~���  }�ƺT�@ �������2  ���  ~���  }�ƺh�@ ������2  �ƺ,�@ ������2  �E����@ �F���ut���   ~��   }�ƺ��@ �����w2  ��   ~��J  }�ƺ��@ �{����V2  ��J  ~��t  }�ƺ��@ �Z����52  �ƺ,�@ �I����$2  �E��ԇ@ �����uS��  ~��5  }�ƺ�@ ������1  ��5  ~��_  }�ƺ �@ �������1  �ƺ,�@ �������1  �E���@ �a�����   ���   ~��  }�ƺ,�@ �����1  ��  ~��5  }�ƺ@�@ �����m1  ��5  ~��_  }�ƺT�@ �q����L1  ��_  ~���  }�ƺl�@ �P����+1  �ƺ,�@ �?����1  �E����@ ������   ���   ~��  }�ƺ��@ ������0  ��  ~��5  }�ƺ��@ �������0  ��5  ~��_  }�ƺЈ@ ������0  ��_  ~���  }�ƺ�@ �����0  �ƺ,�@ �����r0  �E����@ ������   ���   ~��  }�ƺ�@ �c����>0  ��  ~��5  }�ƺ(�@ �B����0  ��5  ~��_  }�ƺ<�@ �!�����/  ��_  ~���  }�ƺP�@ � �����/  �ƺ,�@ �������/  �E��d�@ �i�����   ���   ~��  }�ƺ|�@ �����/  ��  ~��5  }�ƺ��@ �����u/  ��5  ~��_  }�ƺ��@ �y����T/  ��_  ~���  }�ƺ��@ �X����3/  �ƺ,�@ �G����"/  �E����@ �������   ���   ~��  }�ƺԉ@ ������.  ��  ~��5  }�ƺ�@ �������.  ��5  ~��_  }�ƺ�@ ������.  ��_  ~���  }�ƺ�@ �����.  �ƺ,�@ �����z.  �E���@ ������   ���   ~��  }�ƺ,�@ �k����F.  ��  ~��5  }�ƺ<�@ �J����%.  ��5  ~��_  }�ƺL�@ �)����.  ��_  ~���  }�ƺ\�@ ������-  �ƺ,�@ �������-  �E��l�@ �q�����   ���   ~��  }�ƺ��@ ������-  ��  ~��5  }�ƺ��@ �����}-  ��5  ~��_  }�ƺ��@ �����\-  ��_  ~���  }�ƺ��@ �`����;-  �ƺ,�@ �O����*-  �E��Ԋ@ �������   ���   ~��  }�ƺ��@ ������,  ��  ~��5  }�ƺ�@ �������,  ��5  ~��_  }�ƺ�@ ������,  ��_  ~���  }�ƺ,�@ �����,  �ƺ,�@ �����,  �E��@�@ �!�����   ���   ~��  }�ƺX�@ �s����N,  ��  ~��5  }�ƺh�@ �R����-,  ��5  ~��_  }�ƺx�@ �1����,  ��_  ~���  }�ƺ��@ ������+  �ƺ,�@ �������+  �E����@ �y�����   ���   ~��  }�ƺ��@ ������+  ��  ~��5  }�ƺċ@ �����+  ��5  ~��_  }�ƺ؋@ �����d+  ��_  ~���  }�ƺ�@ �h����C+  �ƺ,�@ �W����2+  �E�� �@ ������  ���   ~���   }�ƺ�@ �#�����*  ���   ~���   }�ƺ0�@ ������*  ���   ~��  }�ƺD�@ ������*  ��  ~��5  }�ƺX�@ ������*  ��5  ~��_  }�ƺl�@ �����z*  ��_  ~���  }�ƺ��@ �~����Y*  ���  ~���  }�ƺ��@ �]����8*  ���  ~���  }�ƺ��@ �<����*  �ƺ,�@ �+����*  �E����@ ������   ���   ~��  }�ƺ،@ �������)  ��  ~��5  }�ƺ�@ ������)  ��5  ~��_  }�ƺ �@ �����)  ��_  ~���  }�ƺ�@ �����o)  �ƺ,�@ �����^)  �E��(�@ �������   ���   ~��  }�ƺ@�@ �O����*)  ��  ~��5  }�ƺT�@ �.����	)  ��5  ~��_  }�ƺh�@ ������(  ��_  ~���  }�ƺ|�@ �������(  �ƺ,�@ ������(  �E����@ �U���uS��  ~��5  }�ƺ��@ �����(  ��5  ~��_  }�ƺ��@ �����e(  �ƺ,�@ �y����T(  �E��Ѝ@ �������   ���   ~��  }�ƺ�@ �E���� (  ��  ~��5  }�ƺ��@ �$�����'  ��5  ~��_  }�ƺ�@ ������'  ��_  ~���  }�ƺ$�@ ������'  �ƺ,�@ ������'  �E��8�@ �K�����   ���   ~��  }�ƺP�@ �����x'  ��  ~��5  }�ƺ`�@ �|����W'  ��5  ~��_  }�ƺp�@ �[����6'  ��_  ~���  }�ƺ��@ �:����'  �ƺ,�@ �)����'  �E����@ �����  ���   ~���   }�ƺ��@ �������&  ���   ~���   }�ƺ��@ ������&  ���   ~��  }�ƺ̎@ �����&  ��  ~��5  }�ƺ܎@ �����m&  ��5  ~��_  }�ƺ�@ �q����L&  ��_  ~���  }�ƺ��@ �P����+&  ���  ~���  }�ƺ�@ �/����
&  ���  ~���  }�ƺ�@ ������%  �ƺ,�@ �������%  �E��,�@ �w�����   ���   ~��  }�ƺD�@ ������%  ��  ~��5  }�ƺT�@ �����%  ��5  ~��_  }�ƺd�@ �����b%  ��_  ~���  }�ƺt�@ �f����A%  �ƺ,�@ �U����0%  �E����@ �������   ���   ~��  }�ƺ��@ �!�����$  ��  ~��5  }�ƺ��@ � �����$  ��5  ~��_  }�ƺď@ ������$  ��_  ~���  }�ƺ؏@ �����$  �ƺ,�@ �����$  �E���@ �'����  ���   ~���   }�ƺ�@ �y����T$  ���   ~���   }�ƺ�@ �X����3$  ���   ~��  }�ƺ0�@ �7����$  ��  ~��5  }�ƺD�@ ������#  ��5  ~��_  }�ƺX�@ �������#  ��_  ~���  }�ƺp�@ ������#  ���  ~���  }�ƺ��@ �����#  ���  ~���  }�ƺ��@ �����m#  �ƺ,�@ �����\#  �E����@ �������   ���   ~��  }�ƺА@ �M����(#  ��  ~��5  }�ƺ�@ �,����#  ��5  ~��_  }�ƺ��@ ������"  ��_  ~���  }�ƺ�@ �������"  �ƺ,�@ ������"  �E�� �@ �S�����   ���   ~��  }�ƺ8�@ �����"  ��  ~��5  }�ƺP�@ �����_"  ��5  ~��_  }�ƺh�@ �c����>"  ��_  ~���  }�ƺ��@ �B����"  �ƺ,�@ �1����"  �E����@ ������   ���   ~��  }�ƺ��@ �������!  ��  ~��5  }�ƺđ@ ������!  ��5  ~��_  }�ƺؑ@ �����!  ��_  ~���  }�ƺ�@ �����u!  �ƺ,�@ �����d!  �E�� �@ ������   ���   ~��  }�ƺ�@ �U����0!  ��  ~��5  }�ƺ,�@ �4����!  ��5  ~��_  }�ƺ@�@ ������   ��_  ~���  }�ƺX�@ �������   �ƺ,�@ ������   �E��l�@ �[����  ���   ~���   }�ƺ��@ �����   ���   ~���   }�ƺ��@ �����g   ���   ~��  }�ƺ��@ �k����F   ��  ~��5  }�ƺ��@ �J����%   ��5  ~��_  }�ƺВ@ �)����   ��_  ~���  }�ƺ�@ ������  ���  ~���  }�ƺ��@ �������  ���  ~���  }�ƺ�@ ������  �ƺ,�@ �����  �E�� �@ �/�����   ���   ~��  }�ƺ8�@ �����\  ��  ~��5  }�ƺP�@ �`����;  ��5  ~��_  }�ƺh�@ �?����  ��_  ~���  }�ƺ��@ ������  �ƺ,�@ ������  �E����@ ������   ���   ~��  }�ƺ��@ ������  ��  ~��5  }�ƺē@ �����  ��5  ~��_  }�ƺؓ@ �����r  ��_  ~���  }�ƺ�@ �v����Q  �ƺ,�@ �e����@  �E�� �@ �������   ���   ~��  }�ƺ�@ �1����  ��  ~��5  }�ƺ,�@ ������  ��5  ~��_  }�ƺ@�@ �������  ��_  ~���  }�ƺT�@ ������  �ƺ,�@ �����  �E��h�@ �7����  ���   ~���   }�ƺ��@ �����d  ���   ~���   }�ƺ��@ �h����C  ���   ~��  }�ƺ��@ �G����"  ��  ~��5  }�ƺ��@ �&����  ��5  ~��_  }�ƺД@ ������  ��_  ~���  }�ƺ�@ ������  ���  ~���  }�ƺ��@ ������  ���  ~���  }�ƺ�@ �����}  �ƺ,�@ �����l  �E��$�@ �����  ���   ~���   }�ƺ@�@ �]����8  ���   ~���   }�ƺT�@ �<����  ���   ~��  }�ƺh�@ ������  ��  ~��5  }�ƺ|�@ �������  ��5  ~��_  }�ƺ��@ ������  ��_  ~���  }�ƺ��@ �����  ���  ~���  }�ƺ��@ �����r  ���  ~���  }�ƺ̕@ �v����Q  �ƺ,�@ �e����@  �E����@ �������   ���   ~���   }�ƺ��@ �1����  ���   ~��  }�ƺ�@ ������  ��  ~��5  }�ƺ,�@ �������  ��5  ~��_  }�ƺD�@ ������  ��_  ~���  }�ƺ\�@ �����  ���  ~���  }�ƺt�@ �����g  �ƺ,�@ �{����V  �E����@ �����ut���   ~��   }�ƺ��@ �K����&  ��   ~��J  }�ƺ��@ �*����  ��J  ~��t  }�ƺ̖@ �	�����  �ƺ,�@ �������  �E���@ �r�����   ���   ~��  }�ƺ��@ ������  ��  ~��5  }�ƺ�@ �����~  ��5  ~��_  }�ƺ$�@ �����]  ��_  ~���  }�ƺ8�@ �a����<  �ƺ,�@ �P����+  �E��L�@ �������   ���   ~��  }�ƺh�@ ������  ��  ~��5  }�ƺ|�@ �������  ��5  ~��_  }�ƺ��@ ������  ��_  ~���  }�ƺ��@ �����  �ƺ,�@ �����  �E����@ �"�����   ���   ~��  }�ƺԗ@ �t����O  ��  ~��5  }�ƺ�@ �S����.  ��5  ~��_  }�ƺ��@ �2����  ��_  ~���  }�ƺ�@ ������  �ƺ,�@ � �����  �E��$�@ �z����  ���   ~���   }�ƺ<�@ ������  ���   ~���   }�ƺP�@ �����  ���   ~��  }�ƺd�@ �����e  ��  ~��5  }�ƺx�@ �i����D  ��5  ~��_  }�ƺ��@ �H����#  ��_  ~���  }�ƺ��@ �'����  ���  ~���  }�ƺ��@ ������  ���  ~���  }�ƺȘ@ �������  �ƺ,�@ ������  �E��ܘ@ �N�����   ���   ~��  }�ƺ��@ �����{  ��  ~��5  }�ƺ�@ �����Z  ��5  ~��_  }�ƺ$�@ �^����9  ��_  ~���  }�ƺ<�@ �=����  �ƺ,�@ �,����  �E��T�@ ������   ���   ~��  }�ƺl�@ �������  ��  ~��5  }�ƺ��@ ������  ��5  ~��_  }�ƺ��@ �����  ��_  ~���  }�ƺ��@ �����p  �ƺ,�@ �����_  �E����@ �������   ���   ~���   }�ƺԙ@ �P����+  ���   ~��  }�ƺ�@ �/����
  ��  ~��5  }�ƺ��@ ������  ��5  ~��_  }�ƺ�@ �������  ��_  ~���  }�ƺ$�@ ������  ���  ~���  }�ƺ8�@ �����  �ƺ,�@ �����u  �E��P�@ ����ut���   ~��   }�ƺh�@ �j����E  ��   ~��J  }�ƺ|�@ �I����$  ��J  ~��t  }�ƺ��@ �(����  �ƺ,�@ ������  �E����@ ������   ���   ~��  }�ƺ��@ ������  ��  ~��5  }�ƺК@ ������  ��5  ~��_  }�ƺ�@ �����|  ��_  ~���  }�ƺ��@ �����[  �ƺ,�@ �o����J  �E���@ �����uS��  ~��5  }�ƺ �@ �?����  ��5  ~��_  }�ƺ8�@ ������  �ƺ,�@ ������  �E��P�@ ����t�E��d�@ �x����  ���   ~���   }�ƺx�@ ������  ���   ~���   }�ƺ��@ �����  ���   ~��  }�ƺ��@ �����c  ��  ~��5  }�ƺ��@ �g����B  ��5  ~��_  }�ƺț@ �F����!  ��_  ~���  }�ƺܛ@ �%����   ���  ~���  }�ƺ�@ ������  ���  ~���  }�ƺ�@ ������  �ƺ,�@ ������  �E���@ �L���uS��  ~��5  }�ƺ,�@ �����}  ��5  ~��_  }�ƺ@�@ �����\  �ƺ,�@ �p����K  �E��T�@ �������   ���   ~��  }�ƺh�@ �<����  ��  ~��5  }�ƺ��@ ������  ��5  ~��_  }�ƺ��@ �������  ��_  ~���  }�ƺ��@ ������  �ƺ,�@ ������  �E��Ȝ@ �B�����   ���   ~��  }�ƺܜ@ �����o  ��  ~��5  }�ƺ�@ �s����N  ��5  ~��_  }�ƺ�@ �R����-  ��_  ~���  }�ƺ�@ �1����  �ƺ,�@ � �����  �E��,�@ ������   ���   ~��  }�ƺ@�@ ������  ��  ~��5  }�ƺT�@ �˿���  ��5  ~��_  }�ƺh�@ 調���  ��_  ~���  }�ƺ|�@ 艿���d  �ƺ,�@ �x����S  �E����@ �������   ���   ~��  }�ƺ��@ �D����  ��  ~��5  }�ƺ��@ �#�����  ��5  ~��_  }�ƺ̝@ ������  ��_  ~���  }�ƺ��@ �����  �ƺ,�@ �о���  �E����@ �J�����   ���   ~��  }�ƺ�@ 蜾���w  ��  ~��5  }�ƺ�@ �{����V  ��5  ~��_  }�ƺ0�@ �Z����5  ��_  ~���  }�ƺD�@ �9����  �ƺ,�@ �(����  �E��X�@ ������   ���   ~��  }�ƺl�@ �������  ��  ~��5  }�ƺ��@ �ӽ���  ��5  ~��_  }�ƺ��@ 貽���  ��_  ~���  }�ƺ��@ 葽���l  �ƺ,�@ 耽���[  �E����@ �������   ���   ~��  }�ƺО@ �L����'  ��  ~��5  }�ƺ�@ �+����  ��5  ~��_  }�ƺ��@ �
�����  ��_  ~���  }�ƺ�@ ������  �ƺ,�@ �ؼ���  �E�� �@ �R�����   ���   ~��  }�ƺ4�@ 褼���  ��  ~��5  }�ƺH�@ 胼���^  ��5  ~��_  }�ƺ\�@ �b����=  ��_  ~���  }�ƺp�@ �A����  �ƺ,�@ �0����  �E����@ 誾����   ���   ~��  }�ƺ��@ �������  ��  ~��5  }�ƺ��@ �ۻ���  ��5  ~��_  }�ƺ��@ 躻���  ��_  ~���  }�ƺԟ@ 虻���t  �ƺ,�@ 舻���c  �E���@ ������   ���   ~��  }�ƺ��@ �T����/  ��  ~��5  }�ƺ�@ �3����  ��5  ~��_  }�ƺ$�@ ������
  ��_  ~���  }�ƺ8�@ ������
  �ƺ,�@ �����
  �E��L�@ �Z����  ���   ~���   }�ƺ`�@ 謺���
  ���   ~���   }�ƺt�@ 苺���f
  ���   ~��  }�ƺ��@ �j����E
  ��  ~��5  }�ƺ��@ �I����$
  ��5  ~��_  }�ƺ��@ �(����
  ��_  ~���  }�ƺĠ@ ������	  ���  ~���  }�ƺؠ@ ������	  ���  ~���  }�ƺ�@ �Ź���	  �ƺ,�@ 费���	  �E�� �@ �.�����   ���   ~��  }�ƺ�@ 耹���[	  ��  ~��5  }�ƺ,�@ �_����:	  ��5  ~��_  }�ƺD�@ �>����	  ��_  ~���  }�ƺ\�@ ������  �ƺ,�@ ������  �E��t�@ 膻����   ���   ~��  }�ƺ��@ �ظ���  ��  ~��5  }�ƺ��@ 跸���  ��5  ~��_  }�ƺ��@ 薸���q  ��_  ~���  }�ƺġ@ �u����P  �ƺ,�@ �d����?  �E��ء@ �޺����   ���   ~��  }�ƺ�@ �0����  ��  ~��5  }�ƺ�@ ������  ��5  ~��_  }�ƺ�@ ������  ��_  ~���  }�ƺ4�@ �ͷ���  �ƺ,�@ 輷���  �E��L�@ �6�����   ���   ~��  }�ƺd�@ 舷���c  ��  ~��5  }�ƺt�@ �g����B  ��5  ~��_  }�ƺ��@ �F����!  ��_  ~���  }�ƺ��@ �%����   �ƺ,�@ ������  �E����@ 莹����   ���   ~��  }�ƺ��@ �����  ��  ~��5  }�ƺТ@ 迶���  ��5  ~��_  }�ƺ�@ 螶���y  ��_  ~���  }�ƺ��@ �}����X  �ƺ,�@ �l����G  �E���@ ������   ���   ~��  }�ƺ$�@ �8����  ��  ~��5  }�ƺ8�@ ������  ��5  ~��_  }�ƺL�@ �������  ��_  ~���  }�ƺ`�@ �յ���  �ƺ,�@ �ĵ���  �E��t�@ �>�����   ���   ~��  }�ƺ��@ 萵���k  ��  ~��5  }�ƺ��@ �o����J  ��5  ~��_  }�ƺ��@ �N����)  ��_  ~���  }�ƺԣ@ �-����  �ƺ,�@ ������  �E���@ 薷����   ���   ~��  }�ƺ�@ ������  ��  ~��5  }�ƺ �@ �Ǵ���  ��5  ~��_  }�ƺ8�@ 覴���  ��_  ~���  }�ƺP�@ 腴���`  �ƺ,�@ �t����O  �E��h�@ ����uS��  ~��5  }�ƺ��@ �D����  ��5  ~��_  }�ƺ��@ �#�����  �ƺ,�@ ������  �E����@ 茶����   ���   ~��  }�ƺ��@ �޳���  ��  ~��5  }�ƺؤ@ 轳���  ��5  ~��_  }�ƺ�@ 蜳���w  ��_  ~���  }�ƺ�@ �{����V  �ƺ,�@ �j����E  �E�� �@ ������   ���   ~��  }�ƺ8�@ �6����  ��  ~��5  }�ƺL�@ ������  ��5  ~��_  }�ƺ`�@ �������  ��_  ~���  }�ƺt�@ �Ӳ���  �ƺ,�@ �²���  �E����@ �<�����   ���   ~��  }�ƺ��@ 莲���i  ��  ~��5  }�ƺ��@ �m����H  ��5  ~��_  }�ƺȥ@ �L����'  ��_  ~���  }�ƺܥ@ �+����  �ƺ,�@ ������  �E���@ 蔴����   ���   ~��  }�ƺ�@ ������  ��  ~��5  }�ƺ�@ �ű���  ��5  ~��_  }�ƺ0�@ 褱���  ��_  ~���  }�ƺD�@ 胱���^  �ƺ,�@ �r����M  �E��X�@ ������   ���   ~��  }�ƺp�@ �>����  ��  ~��5  }�ƺ��@ ������   ��5  ~��_  }�ƺ��@ �������   ��_  ~���  }�ƺ��@ �۰���   �ƺ,�@ �ʰ���   �E��Ц@ �D�����   ���   ~��  }�ƺ�@ 薰���t��  ~��5  }�ƺ �@ �x����V��5  ~��_  }�ƺ�@ �Z����8��_  ~���  }�ƺ0�@ �<�����ƺ,�@ �.�����ƺ,�@ � ���3�ZYYd�hM�@ �E�路����ũ����^[Y]�  ����   �� �� һ �� ����   �������(һ��ת��)  ����
   ����(�Ϻ�)  ����
   ��â(�Ϻ�)  ����
   ����(�Ϻ�)  ����
   ����(����)  ����
   ����(����)  ����
   ����(����)  ����
   ��ͨ(�Ͼ�)  ����
   ��ɽ(����)  ����   δ֪    ����   �� �� �� �� ����   ����ʮ��(����ת��)  ����   ������(�Ϻ�)    ����
   ����(����)  ����
   ����(�ɶ�)  ����
   ����(����)  ����
   ��ͨ(�Ϻ�)  ����   �� �� �� �� ����   �������(����ת��)  ����   Ӣ��֮��(����ת��)  ����
   �ɺ�(����)  ����
   ����(�㶫)  ����
   ��ʨ(����)  ����
   �츮(����)  ����
   ����(�ɶ�)  ����   ��â��(�Ϻ�)    ����   �����(�Ϻ�)    ����   ��ա�����(����)    ����   ���ߴ�½(����ת��)  ����
   ���(�Ϻ�)  ����
   ����(�Ϻ�)  ����
   ���(�Ϻ�)  ����
   ��ϼ(�Ϻ�)  ����   ��ȶ�(�Ϻ�)    ����   ���Ķ�(�Ϻ�)    ����   ����(�Ϻ�)    ����   ��ϼ��(�Ϻ�)    ����   �� �� �� �� ����   ������ʮ��(����ת��)    ����
   ��Ȼ(�Ϻ�)  ����
   ���(�Ϻ�)  ����
   ����(�Ϻ�)  ����
   ����(�Ϻ�)  ����   ��Ȼ��(�Ϻ�)    ����   ��ض�(�Ϻ�)    ����   ������(�Ϻ�)    ����   �����(�Ϻ�)    ����   �� �� �� �� ����
   ��Ͽ(��ͨ)  ����
   ���(�ɶ�)  ����
   ���(����)  ����
   ����(����)  ����   ��Ͽ��(��ͨ)    ����   ��Ƕ�(�ɶ�)    ����   ��ض�(����)    ����   ���׶�(����)    ����   �� �� �� �� ����
   �漣(�Ϻ�)  ����
   ����(�人)  ����
   ����(�Ϻ�)  ����
   ���(�Ϻ�)  ����   �漣��(�Ϻ�)    ����   ��¶�(�Ϻ�)    ����   �����(�Ϻ�)    ����   ���Ƕ�(�Ϻ�)    ����   ����֮��(11��)  ����
   ����(�Ϻ�)  ����
   ����(�Ϻ�)  ����
   ˮ�(�Ϻ�)  ����
   ��¥(�Ϻ�)  ����
   ����(�Ϻ�)  ����
   ��ի(�Ϻ�)  ����
   ����(�Ϻ�)  ����
   ս��(�Ϻ�)  ����   ����ʥ��(12��)  ����
   ��ɽ(�츮)  ����
   ѩ��(�츮)  ����
   �ػ�(�츮)  ����
   ��կ(�츮)  ����   ��ɽ(�ػ�ת��)  ����
   ����(�츮)  ����
   ����(�츮)  ����   ����(��կת��)  ����   �ƶ�����(15��)  ����
   ����(�ƶ�)  ����
   ����(�ƶ�)  ����
   �ĺ�(�ƶ�)  ����   ���ǵ���(16��)  ����
   ����(��ͨ)  ����
   ����(��ͨ)  ����   ����ר��(17��)  ����
   ����(��ͨ)  ����
   ����(��ͨ)  ����   ���(NEW!��ͨ)  ����   ����ɽ(NEW!��ͨ)    ����   ���¡�����ǿ�(18��)    ����
   �ٵ�(�°�)  ����
   ����(�°�)  ����
   ��ҵ(�°�)  ����
   �Ի�(�°�)  ����   ����ʥ��II(19��)    ����
   ����(�츮)  ����
   ����(�츮)  ����
   ��ɽ(�츮)  ����
   �ų�(�츮)  ����   ��������(20��)  ����   ���    ����   �̲�    ����   ��ɽ    ����   ��Ұ    ����   ��ɽ�续(21��)  ����   ��ˮ    ����   ����    ����   �׺�    ����   ɣ��    ����   ��ͨ���(22��)  ����   ��    ����   �Ͻ�    ����   ����    ����   ����    ����   Ⱥ����¹(23��)  ����
   ���(�Ϻ�)  ����
   ����(�Ϻ�)  ����
   ����(�Ϻ�)  ����
   �޵�(�Ϻ�)  ����   ����ʥ��III(24��)   ����
   ����(����)  ����
   ����(üɽ)  ����
   ����(�츮)  ����
   ����(�츮)  ����   ����II(25��)    ����   Խ��    ����   ����    ����   �齭    ����   ��ӡ    ����   ��Ů��(26��)    ����
   ����(����)  ����
   ����(����)  ����
   ����(����)  ����
   ����(����)  ����   ��ͨ���II(27��)    ����
   ����(�人)  ����
   ����(�人)  ����
   ����(����)  ����
   ����(����)  ����   ����(�ػʵ�)    ����
   ȡ��(��̨)  ����
   �Ǻ�(����)  ����
   ����(�Ͳ�)  ����   ���δ���(28��)  ����
   Ǭ��(����)  ����
   ����(����)  ����
   ����(����)  ����
   �ݼ�(����)  ����   �����籩(29��)  ����
   ����(̨��)  ����
   ����(̨��)  ����
   ����(̨��)  ����
   ն��(̨��)  ����   ��������(30��)  ����
   ��ң(�Ϸ�)  ����
   ����(�Ϸ�)  ����   ������(31��)    ����
   ���(����)  ����
   ����(����)  ����
   ����(�Ϻ�)  ����
   ��˫(�Ϻ�)  ����   Ӣ�����(32��)  ����   ��ɽ    ����   ����    ����   ����    ����   ����    ����   ����ʥ��IV(33��)    ����   ����    ����   �ٶ�    ����   ����    ����   ���    ����   ��Դ    ����   �׵�    ����   ����    ����   ��ˮ    ����   �����(34��)    ����   ����    ����   ��Ծ    ����   ����    ����   ӥ��    ����   ���յ���(35��)  ����
   ����(����)  ����
   ����(����)  ����
   ���(�Ϻ�)  ����
   ����(�Ϻ�)  ����   ��ͨ���III(36��)   ����
   ��ԭ(�Ͼ�)  ����
   ���(�Ͼ�)  ����
   �ػ�(�Ͼ�)  ����
   ��©(�Ͼ�)  ����   �о�(ʯ��ׯ)    ����   �峯(ʯ��ׯ)    ����   ��Į(ʯ��ׯ)    ����   ���(ʯ��ׯ)    ����   �ų�����(37��)  ����   ��(����)    ����   ��(����)    ����   ��(����)    ����   ��(����)    ����   ����III(38��)   ����   �ƺ�¥(�Ϻ�)    ����   �紨��(�Ϻ�)    ����   ���ݳ�(�Ϻ�)    ����   �䵱ɽ(�Ϻ�)    ����   ����IV(39��)    ����
   ̫��(�Ϻ�)  ����
   ��ɽ(�Ϻ�)  ����
   ����(�Ϻ�)  ����
   ����(�Ϻ�)  ����   �����޵�(41��)  ����
   ����(����)  ����
   ����(�ϲ�)  ����   ��ˮ(������)    ����
   �ǳ�(��ɳ)  ����   ����V(42��) ����
   ����(�Ϻ�)  ����
   �ص�(�Ϻ�)  ����
   ���(�Ϻ�)  ����
   ����(�Ϻ�)  ����
   ����(�Ϻ�)  ����
   ��Դ(�Ϻ�)  ����
   �A��(�Ϻ�)  ����
   ��ϼ(�Ϻ�)  ����   ������(43��)    ����   ɽ����(����)    ����   ���ܴ�(����)    ����   ս����(����)    ����   ����Ե(����)    ����   ����ʥ��(44��)  ����
   �潭(����)  ����
   ��ͥ(����)  ����
   ��ɽ(����)  ����
   ����(����)  ����   ����ʥ��V(45��) ����
   ����(�ɶ�)  ����
   ���(�ɶ�)  ����
   ǭ��(����)  ����
   ��Ϫ(����)  ����   ��¹��ԭ(46��)  ����
   Ӣ��(֣��)  ����
   ��ɷ(֣��)  ����
   ����(����)  ����
   ���(����)  ����
   �ݺ�(�Ϻ�)  ����   Ӣ��(����Ͽ)    ����
   ս��(�Ϻ�)  ����
   ����(�Ϻ�)  ����   ����ʥ��VI(47��)    ����
   ����(����)  ����
   ��(��ɽ)  ����
   ��(�˱�)  ����
   �Ƴ�(®��)  ����
   ����(�ϳ�)  ����
   ���(�ڽ�)  ����
   ���(�Ű�)  ����
   ����(����)  ����   ��ͨ���IV(48��)    ����   �Ǻ���(����)    ����   ǧɽһ(��ɽ)    ����   ǧɽ��(����)    ����   ʢ��һ(����)    ����   ʢ����(����)    ����
   ����(����)  ����   ����ǿ�II(49��)    ����
   ���(��ɽ)  ����
   ���(���)  ����   �����(���)    ����   �����(50��)  ����
   ����(���)  ����
   ����(���)  ����
   �н�(���)  ����
   ��ѩ(���)  ����   ����ͨ��ר��(51��)  ����
   ����(����)  ����
   ����(����)  ����
   ����(�Ϻ�)  ����
   ����(�Ϻ�)  ����   �㽭����ר��(52��)  ����
   ����(����)  ����
   ����(����)  ����
   ����(����)  ����
   ˫��(����)  ����   ��ʹ֮��(53��)  ����
   ����(����)  ����
   ܽ��(��ɳ)  ����
   ����(��ɳ)  ����
   ��ɳ(��ɳ)  ����
   ��ɽ(��ɳ)  ����
   ��ɽ(��ɽ)  ����
   �ŵ�(̫ԭ)  ����
   ����(̫ԭ)  ����   ���´���(54��)  ����   ����(ԭ����)    ����   ����(ԭ����)    ����   ����(ԭ�׹�)    ����   �޵�(ԭ���)    ����   ��³����(55��)  ����
   ���(��̨)  ����
   ���(��̨)  ����
   �ٵ�(�ൺ)  ����
   ����(����)  ����   ���ǿ��(56��)  ����
   ����(�Ϻ�)  ����
   ����(����)  ����
   ��ˮ(�Ϻ�)  ����
   ����(�Ϻ�)  ����
   ����(�Ϻ�)  ����   �׻�(�Ϻ�����)  ����   �½�����(57��)  ����
   ˿·(�½�)  ����
   ����(�½�)  ����
   �ŵ�(�½�)  ����   ��ͨר��(58��)  ����
   ��ɽ(�½�)  ����
   ɳĮ(�½�)  ����
   ����(�Ϻ�)  ����
   ����(�Ϻ�)  ����
   ����(59��)  ����   ̩��(������)    ����   ����(������)    ����
   ����(60��)  ����   �������˸�) ����
   ��Ӱ(�ɶ�)  ����
   ����(�ɶ�)  ����
   ����(�ɶ�)  ����
   ����(�ɶ�)  ����
   �ƿ�(����)  ����
   ����(����)  ����
   ����(����)  ����	   ����(����   ����
   ����(61��)  ����
   ����(����)  ����
   ����(����)  ����
   ����(62��)  ����   ����(����ͨ��)  ����   ����(����ͨ��)  ����   ����(���ͨ��)  ����   ̫ԭ(̫ԭͨ��)  ����
   ����(63��)  ����
   ����(����)  ����
   ����(����)  ����
   ����(����)  ����
   ����(����)  ����
   ����(64��)  ����
   ����(����)  ����
   ����(����)  ����
   �ļ�(�Ϻ�)  ����
   ƽ��(�Ϻ�)  ����
   ����(65��)  ����
   ��¥(����)  ����
   ��ɽ(����)  ����
   ̨��(����)  ����
   ����(����)  ����
   ����(66��)  ����
   ����(����)  ����
   ��˵(����)  ����
   ʧ��(����)  ����
   ħ��(����)  ����
   ����(67��)  ����
   �ɽ�(����)  ����
   Īа(����)  ����
   տ¬(����)  ����
   ����(����)  ����
   ����(68��)  ����
   ��ѧ(����)  ����
   ��ӹ(����)  ����
   ����(����)  ����
   ����(����)  ����
   ����(69��)  ����
   ��ɽ(����)  ����
   ��ˮ(����)  ����
   Ȫ��(����)  ����
   ����(�Ϻ�)  ����
   ����(70��)  ����
   ��ʩ(����)  ����
   ����(����)  ����
   ��(����)  ����
   �Ѿ�(����)  ����
   ����(71��)  ����
   ����(��)  ����
   ��ȸ(����)  ����
   ����(����)  ����
   ¹��(����)  ����
   ����(72��)  ����
   ����(��ɳ)  ����
   ����(��ɳ)  ����
   ��´(��ɳ)  ����
   �껨(��ɳ)  ����
   ����(��ɳ)  ����
   ����(��ɳ)  ����
   ����(����)  ����
   ��Դ(����)  ����
   ����(75��)  ����   ������(�Ϻ�)    ����   ��ū��(�Ϻ�)    ����   ������(�Ϻ�)    ����   ̤ɯ��(�Ϻ�)    ����
   ����(76��)  ����
   ����(�ɺ�)  ����
   ����(�ɺ�)  ����
   ��Ӱ(����)  ����
   ����(����)  ����
   ����(77��)  ����   ������(�Ϻ�)    ����   ���կ(�Ϻ�)    ����   ʮ����(�Ϻ�)    ����   Ұ����(�Ϻ�)    ����   ��������(78��)  ����   ��Ǯ��  ����   ��ķ��  ����   ��ɽ��  ����   ����̶  ����   ��Ѫ����(79��)  ����
   ����(����)  ����
   ����(����)  ����
   Ҭ��(����)  ����
   ����(����)  ����   ��˿·(80��)    ����
   �߲�(�½�)  ����
   ����(�½�)  ����
   ����(�½�)  ����
   ����(�½�)  ����   ���¹��(81��)  ����   ���ͨ(����)    ����   ����ͨ(����)    ����   ����ͨ(����)    ����   ����쳵(����)  ����   ˮ����ɽII(82��)    ����   �׻���(����)    ����   ������(����)    ����   �����(����)    ����   �����(����)    ����   Ӣ��֮��(83��)  ����
   �ĺ�(�㽭)  ����
   ����(�㽭)  ����   ��������(84��)  ����   �Ӷ�ʨ��(̫ԭ)  ����   ��������(̫ԭ)  ����   ̫�йŷ�(̫ԭ)  ����   ���Ų�ѩ(̫ԭ)  ����   ���۷���(85��)  ����
   ����(�人)  ����
   ��Ͽ(�人)  ����
   ��̨(�人)  ����
   ���(�人)  ����   ���e��(86��)   ����
   ��̩(��Ӫ)  ����
   ����(��Ӫ)  ����
   ��ͨ(��Ӫ)  ����
   ���(��Ӫ)  ����   Ц������(87��)  ����
   �齣(��ɽ)  ����
   ���(��ɽ)  ����
   ����(��ɽ)  ����
   ����(��ɽ)  ����   ������(88��)  ����   ��ɳ�ӣ����ڣ�  ����   ����ɽ�����ڣ�  ����   ˮ���������ڣ�  ����   �����ţ����ڣ�  ����   ��Ƚ��(89��)  ����   ��ѩ����������  ����   ���ӣ���������  ����   �ʳ���������    ����   �����������    U�������SVW3��������������������E�3�Uht�@ d�0d� 3�j �b���P�d����؅���   h�   ������PS�P�������   j h��@ ����������   h�   ������PV� ����U�������袔���E����@ �����tO������P�   �   �E����������������������������P���������@ �ޔ��������X覊��u���jS蠓���؅��<���3�ZYYd�h{�@ �������   赇���E�艇���闁������_^[��]�TFRMMAIN    ����
   ����ͻ���  ����   legend of mir   S�� �����h�   �T$RP�����Ӌ�螓����   [Ë�S�� �����h�   �T$RP�˒���Ӌ��r�����   [Ë�U�������SV3��������u3�Uh��@ d�0d� �h�   �� ���PV耒���������� ��������������ȩ@ �o���u&���@ �=��@ u�5��@ ��=��@ u�5��@ 3�ZYYd�h��@ �������O�����]������^[��]�  ����   TEdit   U��3�QQQQ3�Uhê@ d�2d�"3҉��@ j h�@ P谑���=��@ ��   ���@ P��������   ���@ P�Ց����t}�U����@ �����E�U��u����U��@ �l����E��U��]����}� tG�}� tA�E��!����Сp�@   �����E������Сp�@   ������p�@ ǀ4     3�ZYYd�hʪ@ �E�   �^�����H�����]Ë�U��ĔSVW3ɉM܉U���3�Uhѭ@ d�0d� �E� �E������Sj h  �z����E�}� ��  �E�P�D����E��E��E��E�3�Uh��@ d�2d�"j�E�P�E�P�E�P�O����E��E�}�   �!  �E܋U�詉���E�P�E�P�E�����P�E�P�E�P����3��E��E��
��
��  @�EԾ
   �E܀|0�/�}  �E܊0<0�o  <2�g  �E܀|00�Y  �E܀|09�K  �E܀|0/�=  �������3�RP���$T$���U܊\���/t��*t�� rI���uу���   �L9�M؍~3ɋ�3�RP���$T$���U܀|�/t*��3�RP���$T$���U܊\���0r��9wA��u���3�RP���$T$���U܀|�/��   A�3ɋ�3�RP���$T$���U܀|�/t*��3�RP���$T$���U܊\���0r��9wA��u���3�RP���$T$���U܀|�/u#A��E܊D8�<0t<1u�E܀<8/u�E؉E��
F�M��k����}� v@�M�I�Eܺ   �ֆ���E�P�M����   �   �E��|����E�� ������
|�E���E�E�;E�s�E�����3�ZYYd��
�A{����|���E�3��b����E�P虍��3�ZYYd�hح@ �E��,�����:|�����E�_^[��]Ë�U��   j j Iu�SVW��p�@ 3�Uh�@ d�0d� j h�@ 蝍���؅�u�ƺ�@ �'����  �U��������E�P�   �   �E�蚅���Eغ8�@ 聄��u�E�PS荍����ƺ�@ �ہ���^  �U�E��K�����u�ƺP�@ 軁���>  �  �   葍���  �   耍���  �   �o����   �   �^����$  �   �M����(  �   �<����,  �   �+����0  �   �����E��Ҁ���E��ʀ���E�����E�躀���E�8*u�E��   �   �̄���U��|�@ �c����؍E�P��I�   �E��i����E�˺   蚄���E� <0u�Eຈ�@ ������(<1u�Eຘ�@ �݀���<2�  �Eຨ�@ �ƀ���E��   �   �H����U��|�@ �߄���؍E�˺   �*����U��|�@ ������؍E�P��I�   �E��ǃ���E�˺   ������E� <0u�E亸�@ �N����<1��  �E�ĳ@ �7����E��+����Ћ  �����E������Ћ  �����E�������Ћ$  �����EԹг@ �U��-����E��ق���Ћ,  �ˋ���u�hܳ@ �u�h�@ �u�hг@ �u��E�   �c����6h��@ �u��ƺ   �M����E���~���E���~���E���~���E���~���E��   �   �����U��|�@ 芃���؍E�P��I�   �E�萂���E�˺   ������E� <0u�Eຈ�@ ����(<1u�Eຘ�@ ����<2�>  �Eຨ�@ ��~���E��   �   �o����U��|�@ �����؍E�˺   �Q����U��|�@ �����؍E�P��I�   �E������E�˺   �����E� <0u�E亸�@ �u~���<1u�E�ĳ@ �b~���E��V����Ћ  �H����E��@����Ћ   �2����E��*����Ћ(  �����Eйг@ �U��X���E������Ћ0  ������u�hܳ@ �u�h�@ �u�hг@ �u��E�   ����6h�@ �u�ƺ   �x��3�ZYYd�h��@ �Eк   �.}����w����_^[��]�   TFRMMAIN    ����   û�з������е� Mir2 ��  ����   legend of mir   ����    ȡ Mir2 ��ɫ��Ϣʧ�ܣ�
�����ԡ�    ����   /   ����   ��ʿ    ����   ħ��ʦ  ����   ��ʿ    ����   ��  ����   Ů  ����   ��  ����   (   ����   )   ����   ����A-  ����   
����B-    U��ĨSVW3ɉM�U���3�UhR�@ d�0d� �E� �E��{��Sj h  �:����E�}� ��   �E�P�����]̋EЉE�3�Uh�@ d�2d�"j�E�PS�E�P�����u��}�   ur�E���w����E�PV�E���~��PS�E�P�׆��������t�U�l�@ ��������U踀�@ ��������v��  ��v�E�P��$  �׋E���~���E�����;E�s���b���3�ZYYd��
��s���su���E�3������E�P����3�ZYYd�hY�@ �E��z����t�����E�_^[��]� ����   On Win95    ����   WinSock 2.0 U��3�QQQQQQQSVW��E�3�Uh7�@ d�0d� �E���{���E�8  �E�   ���,z���E��D������   ��t��~��4�  �E�P�S�ϋE���}���U��P�@ �~������   ���$  ��   �E��f{�����E�U��9����E��A�����+Ѓ�|	�+ǃ�~��4�   ��E��i~������~z�E�P��I��   �l}���ƋϺ   �}����d�@ �6~�����O�ƺ   �}���E��u��U�E�茆���u�hd�@ �E��   �{���u��u��6�ƺ   �o{����E�   �6�u�hd�@ �ƺ   �P{����4;]������3�ZYYd�h>�@ �E���x���E��~���E��   ��x�����r����_^[��]�   ����   {���q���{�� ����   
  U�������SV3҉������U��U��3�Uhf�@ d�0d� j ht�@ �����؅�u�ƺ��@ �x���   h�   ������PS�&����U�������訄��������P�   �   �E���{�����������@ ��z��u�E�PS������ƺ��@ �9x���'�U�E��������u�ƺ��@ �x���
�֋E��P���3�ZYYd�hm�@ �������w���E��   �w����q����^[��]� TFRMMAIN    ����   û�з������е� Mir2 ��  ����   legend of mir   ����    ȡ Mir2 ������Ʒʧ�ܣ�
�����ԡ�    U��3�QQQQSVW�}�]�E3�Uh��@ d�2d�"3���}WSP�x�@ P艂������   �uf��ua蕂���؍U��������U����w����U�E�踃���E����@ �y��u,�E�P�   �   �E��sz���E�Թ@ �Zy��u���E���3�ZYYd�h��@ �E�   �{v����ep�����_^[��]� ����   TFRMMAIN    ����   legend of mir   U����SV3ɉM���E��E��y��3�Uh��@ d�0d� ����u���U����@ �z���؅�~:�6�E�P��I�   �E��y���u�hȺ@ �ƺ   � x���K�E��   ��y�������%w����|�/u��w���Ћƹ   �y��3�ZYYd�h��@ �E��   �}u����go����^[YY]�   ����   
  ����   /   U��j j 3�UhO�@ d�0d� ���@ Pj �����E��r����E��U�������E��x���Сp�@   �v����p�@ � ��tj j h�  P�؀��3�ZYYd�hV�@ �E��   ��t����n����YY]� U�������SV3��������������������������������������E��E��E�]�E3�UhC�@ d�2d�"3���}�URSP�|�@ P��������  �A  �l����؅��2  �U���� ����U���������������E������������\�@ ��v����  �E��p�@ �v��u~j h|�@ j S���ƅ���� ������Rj$jP���������� ��  �������p�@ ���$����O�����t�p�@ � ��tj j h�  P�}���p�@ ǀ4     �m  ������P�   �   �E��,w�����������@ �v���>  �p�@ ��4  HtHtjH�O  H��  �  ǅ�����  ǅ����Q  ǅ�����  ǅ����m  �E�P�~���u��u�������P��~������  ��������  �n�����t�p�@ � ��tj j h�  P�~��ǅ����4  ǅ�����   ǅ�����  ǅ�����  �E�P�3~���u��u�������P�a~�����U  �������p�@ ���   �s���������������U�蘄��������P�������E������������E�Z��s���E��|u���Сp�@   �k~���p�@ ǀ4     ��   ǅ�����  ǅ�����  ǅ�����  ǅ�����  �E�P�j}���u��u�������P�}������   �������U����p�@ ǀ4     �pǅ����h  ǅ�����  ǅ�����  ǅ�����  �E�P�}���u��u�������P�1}����t)�p�@ 3҉�4  h̺@ h N  ���@ Pj �}�����@ 3�ZYYd�hJ�@ �������   ��p���E���p���E��   ��p�����j���Ӌ�^[��]� ����   TFRMMAIN    ����
   ����ͻ���  TComboBox   ����   legend of mir   VW�l�@ �p�@ �x�H�@ �   �p�@ 3҉�4  �=|�@  uj �P�@ Ph\�@ j�E|���|�@ ��}����t�=|�@  �����_^Ã=x�@  uj �P�@ Ph�@ j�	|���x�@ �=|�@  t	�=x�@  u3������_^�                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                 �=x�@  t�x�@ P��w����t3��x�@ �=|�@  t�|�@ P�w����t3��|�@ �=|�@  u	�=x�@  t3������ÐU��j S3�Uh%�@ d�0d� �=x�@  u@�E��<�@ ��k���U��   �|�@ �o���E��k��j �P�@ Ph�@ j�0w���x�@ �=x�@  �����3�ZYYd�h,�@ �E���j�����d������[Y]�  ����5   SOFTWARE\Microsoft\Windows NT\CurrentVersion\Winlogon   ����   huanqi  �=x�@  t�x�@ P�v����t3��x�@ �=|�@  �����Ë�U��3�Uh��@ d�0d� �h�@ u$�=l�@  t�m����p�@ P�u���t�@ P�cu��3�ZYYd�h�@ ��d����]Ã-h�@ sn�l�@  h��@ j j�Vu���t�@ �=t�@  uh��@ h4  j jj j��u���t�@ �=t�@  tj j j j�t�@ P�u���p�@ 3��|�@ 3��x�@ �My_Mir2_MapFile U��3�Uh��@ d�0d� 3�ZYYd�h��@ ��\c����]�   ��@ ;@ �:@ |8@ (8@ L;@ ;@ t<@ D<@ �@ ��@     ��@ U���ĸ��@ �s���h���@                                                                                                                                                                                                                                                                 �@ 2�� �@  �@  �@         |@  @ �#@  ��������������������� ��@ Error ��Runtime error     at 00000000 ��0123456789ABCDEF����                        ,:@ �9@ �9@ :@                                                                                                                                                                                                                                                                                                                                                            ��  @�              ��  $�              ��  ��              ��  �              ��  �              ��  l�              �  ��                      �  �  2�  H�  d�  r�  ��  ��  ��  ��  ��  ��  ��  ��  �  �  "�  0�  <�  V�  b�  r�      �  �      ��  ��  ��      ��  ��      ��  ��  ��  ��  ��  ��      �  $�  6�  J�  X�  j�  z�  ��  ��  ��      ��  ��  ��  �  �   �  .�  :�  L�  f�  v�  ��  ��  ��  ��  ��  ��  ��  ��      KERNEL32.DLL KERNEL32.DLL KERNEL32.DLL advapi32.dll oleaut32.dll user32.dll user32.dll    VirtualQueryEx  UnmapViewOfFile   ReadProcessMemory   OpenProcess   OpenFileMappingA  MapViewOfFile   GetVersionExA   GetSystemInfo   CreateFileMappingA  CloseHandle   TlsSetValue   TlsGetValue   TlsFree   TlsAlloc  LocalFree   LocalAlloc  DeleteCriticalSection   LeaveCriticalSection  EnterCriticalSection  InitializeCriticalSection   VirtualFree   VirtualAlloc  LocalFree   LocalAlloc  GetVersion  GetCurrentThreadId  MultiByteToWideChar   GetThreadLocale   GetStartupInfoA   GetLocaleInfoA  GetCommandLineA   FreeLibrary   ExitProcess   WriteFile   UnhandledExceptionFilter  RtlUnwind   RaiseException  GetStdHandle  RegQueryValueExA  RegOpenKeyExA   RegCloseKey   SysFreeString   SysAllocStringLen   UnhookWindowsHookEx   SetWindowsHookExA   SetTimer  SendMessageA  PtInRect  PostMessageA  KillTimer   IsWindowVisible   GetWindowThreadProcessId  GetWindowTextA  GetWindow   GetForegroundWindow   GetCursorPos  GetClassNameA   GetActiveWindow   FindWindowExA   FindWindowA   EnumChildWindows  CallNextHookEx  GetKeyboardType   MessageBoxA                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                     P           (  8  H  H�  ��  ��  ��  \  r  �  �       Mir2Dll.dll DisableKeyboardHook9X EnableKeyBoardHook9X StartHook StopHook                                                                                                                                                                                                                                                                                                                                                                          $  0
000"0*020:0B0J0R0Z0b0j0r0z0�0�0�0�0�0�0�0�0�0�0�0�01(101�1�1�2^3�3�34|4�4555A5\5�5>7z7�7�7�7�7�7�7�7�7�7�788 8.848<8N8Z8i8u8}8�8�8�8�8�8�8�8�8�8�8�8999 979B9c9{9�9�9�9�9:_::�:�;�;<<&</<8<C<L<S<b<i<�<�<�<q=�=�=�=>>>%>j>s>�>�>�>�>�> ?:?d?m?}?�?�?�?�?�?�?�?�?�?�?�?      $  0000H0T0\0s0�0�0�0�0�0�0�0141X1v1�1�1�1�1222#2,2}2�2�2�2�2�2�2�2�2�2p3�3�3�3�3%4+434W4w4�4�4�4�4�45$5�5�6!717G7e7{7�7�7�7�7
88(8@8N8�8�8�8�8�8�8989A9s9|9�9�9�9':O:�;�;�;�; <4<<<G<s<�<�<�<�<0=@=F=L=R=W=]=f=v={=�=�=�=�=�=�=�=�=�= >,>7>T>^>�>�>�>�>�>�>�>�>�>�>???=?Q?�?�?�?�? 0    )1�3�6�667=7O7m7v7�7�7�78/8;8B8L8V8m8~8�8�8�8�8�8�8�8�8�8�8�8�8�89/9@9J9R9Z9b9j9r9z9�9�9�9�9�9::<:D:R:W:p:�:�:�:�:�:�:�:�:�:;;#;/;<;N;V;^;f;n;v;~;�;�;�;�;�;�;�;�;�;�;�;�;�;�;�;�;<<<<&<.<6<K<W<d<v<R=�=�=>+>R>a>p>�>�>�>�>??.?=?L?[?�?�?�?�?�?�?   @    00^0�0�0�0�0�2�2�2�2�23;3\3}3�3�3�3�3�3444U4v4�4�4�4�455,5;5]5~5�5�5�56#6D6U6g6v6�6�6�6�67=7^77�7�7�7�7�7868W8x8�8�8�8�8�8 9A9b9�9�9�9�9�9	:+:L:m:�:�:�:�:;#;5;W;x;�;�;�;�;<><O<a<�<�<�<�<=(=I=j={=�=�=�=�=�=>.>O>`>r>�>�>�>�>??<?]?~?�?�?�?�?   P  ,  0&0G0X0j0�0�0�0�0 1141U1v1�1�1�1�1�12?2P2b2�2�2�2�2�2
3,3M3n3�3�3�3�3�3474H4Z4|4�4�4�4�45$5E5f5�5�5�5�566.6P6q6�6�6�6�6�67:7[7l7~7�7�7�7�78#8D8e8v8�8�8�8�89909R9s9�9�9�9�9:9:J:\:~:�:�:�:�:;&;G;h;�;�;�;�;�;<1<R<s<�<�<�<�<�<=<=]=n=�=�=�=�=>>(>J>k>�>�>�>�>�>?4?U?f?x?�?�?�?�?   `  (  0?0`0�0�0�0�0�01)1:1L1n1�1�1�1�1�1272X2y2�2�2�2�2 3!3B3c3�3�3�3�3�34,4M4n4�4�4�4�4�4575X5y5�5�5�5�5�56>6O6a6�6�6�6�6�6	7+7L7m7�7�7�7�7�7868G8Y8{8�8�8�8�8 9A9b9s9�9�9�9�9
::-:O:p:�:�:�:�:�:;9;Z;{;�;�;�;�;�;<0<B<d<�<�<�<�<�<=)=:=L=[=}=�=�=�=>">C>d>u>�>�>�>�>�>?,?M?n??�?�?�?�? p  ,  0'090[0|0�0�0�0�01$1E1f1w1�1�1�1�12212S2t2�2�2�2�2�23=3^3o3�3�3�3�344)4K4l4�4�4�4�4�4555V5g5y5�5�5�5�56@6a6�6�6�6�6�6	7*7;7M7o7�7�7�7�7�7888Y8z8�8�8�8�89"939E9g9�9�9�9�9�9:0:Q:r:�:�:�:�:�:;+;=;_;�;�;�;�;�;<$<5<G<i<�<�<�<�<�<=2=S=t=�=�=�=�=�=>->?>a>�>�>�>�>�>	?*?K?l?}?�?�?�?�? �     00'090 �  X   g7�7�7!8W8.9d9q9w9�9�9�9�9�9�9�9�9
::/:G:r:�:�:�:�:0;�=�=>> >R>l>�>`?�?�?�?�? �  �   0=0T0�0�0�0�0�091t1�1�1�1�12)2x2�2�2�2�2�2'4m4�4�4E5�56�6�6�67�7�7�7�78+8I8�89T9y9�9::@:�:�:�:;;=;�;�;<<(<`<v<�<�<�<W=�=>&>�>�>�>�>??�?�?�?�?�?�?�?�?�?   �  �   000$0*030J4R4c4i4q4�4�4�4�4�4�4�4�4�4�455�5�5�5�5�5�5�5�5�5�5
666'6-656L6R6b6m6t6{6�6�6�6�6�6�6�6�6�6�6�6�6�6�6�6 �     $0(0,0�0�0�0�0                                                                                                                              vh�0       
     �    vh�0       �  �8  ��  �`  �    vh�0           P   �                 vh�0           x   �  L            D V C L A L  P A C K A G E I N F O   &=O87��$B�:�  �       Mir2Dll KWindows  �System  �SysInit UTypes  Unit_DllMain                                                                                                                                                                                                                                                       