MZ�       ��  �       @                                   �   � �	�!�L�!This program cannot be run in DOS mode.
$       ��ù����������������������������퐺���Q�������Rich����                        PE  L *1�F        � �E  @        �  @D                          �T  �  8                               `N  (                           �R  �  �D  T                                           @D  �                           .text   �A  �  �A  �                 h.rdata  \  @D  `  @D              @  H.data   �  �E  �  �E              @  �INIT      `N     `N                 �.reloc    �R     �R              @  B                U��QSVW�e� ��E�@�E��E�;Es�E��M�A��y�M��Uf�J���   P1��   3��   �   Y�   �����XQ������E��Mf�$A _^[�� U���t  SVW�   P1��   3��   �   Y�   �����XQ�����Q�   Ǆ Y�   ��
Q��5�%�YS�   ��S��[����[Q�   Ǆ Y�   ��
Q��5�%�YQ�   Ǆ Y�   ��
Q��5�%�Y��l���Pj	h�E �����hLF ��l���P�u�'  �   P1��   3��   �   Y�   �����XQ������   P1��   3��   �   Y�   �����XQ�����hLN hLF �  �PN Q�   Ǆ Y�   ��
Q��5�%�Y�=LN  t,hXN �5LN �e  �TN �   �   ������  ���E�0F Q�   Ǆ Y�   ��
Q��5�%�Y�  ����u=3��'  Q�   Ǆ Y�   ��
Q��5�%�YQ�   Ǆ Y�   ��
Q��5�%�Y��!  ����u=3���  Q�   Ǆ Y�   ��
Q��5�%�YQ�   Ǆ Y�   ��
Q��5�%�Y�E�@4d( Q�   Ǆ Y�   ��
Q��5�%�Y�   �   ������  ��S�   ��S��[����[Q�   Ǆ Y�   ��
Q��5�%�Y������Pjh�E �����Q�   Ǆ Y�   ��
Q��5�%�Y�   �   ������  ��������P������P�PD ��4���Pjj h �  ������Pj �u�LD ������P�
   ǃ���   X�   � ���   �P��XS�   ��S��[����[������ }"3��k  Q�   Ǆ Y�   ��
Q��5�%�Y��8���Pjh�E �����Q�   Ǆ Y�   ��
Q��5�%�Y�   �   ������  ����8���P������P�PD ������P������P�HD ������������ ��   ��4��� t:��4����DD �   �   ������  ���   �   ������  ��3��  Q�   Ǆ Y�   ��
Q��5�%�YP�
   ǃ���   X�   � ���   �P��X�E�@8Z* �E�@@Z* Q�   Ǆ Y�   ��
Q��5�%�Y�E�@pB+ �   P1��   3��   �   Y�   �����XQ������   �   ������  ���=TN  t�5XN �5TN ��  �   �   ������  ���   P1��   3��   �   Y�   �����XQ������50F h�= j j j j ������P�@D ������S�   ��S��[����[3��%P�
   ǃ���   X�   � ���   �P��X_^[�� �U���8SVWP�
   ǃ���   X�   � ���   �P��XS�   ��S��[����[�   �   ������  ���e� �   P1��   3��   �   Y�   �����XQ������E�   Q�   Ǆ Y�   ��
Q��5�%�Y�E���E��   P1��   3��   �   Y�   �����XQ������   �   ������  ���e� Q�   Ǆ Y�   ��
Q��5�%�YhDdk �u�j�dD �E��}� u
�"  ��{  Q�   Ǆ Y�   ��
Q��5�%�YP�
   ǃ���   X�   � ���   �P��X�u�E�P�PD �E�   �e� �E�@   �E�Eԃe� �e� P�
   ǃ���   X�   � ���   �P��X�E�Ph?  �E�P�`D �E�}� }�E���  �M�3��}������ʃ��E�P�u��u�j�E�P�u��\D �E��   �   ������  ���E�Eȁ}�  �t'�}� ��   �#  S�   ��S��[����[�u��XD Q�   Ǆ Y�   ��
Q��5�%�Y�   �   ������  ���E���E�hDdk �u�j�dD �E��E�P�u��u�j�E�P�u��\D �E�Q�   Ǆ Y�   ��
Q��5�%�Y�}� }1�uS�   ��S��[����[�   �   ������  ���E��M�HQ�u�TD YY�/�   P1��   3��   �   Y�   �����XQ������u��XD 3��.�   �   ������  ���   �   ������  ��_^[�� �U���LSVW�e� Q�   Ǆ Y�   ��
Q��5�%�YQ�   Ǆ Y�   ��
Q��5�%�YQ�   Ǆ Y�   ��
Q��5�%�YQ�   Ǆ Y�   ��
Q��5�%�Y�e� Q�   Ǆ Y�   ��
Q��5�%�Y�   �   ������  ���u�E�P�PD �E�   �e� �E�@   �E��E�e� �e� h`  j�E�P�E�Ph�  �E�P�tD �E�Q�   Ǆ Y�   ��
Q��5�%�Y�}� },3��B  P�
   ǃ���   X�   � ���   �P��Xjj�E�P�E�P�u��pD �E��   �   ������  ��P�
   ǃ���   X�   � ���   �P��X�}� }x�u��lD Q�   Ǆ Y�   ��
Q��5�%�YQ�   Ǆ Y�   ��
Q��5�%�Y3��}  �   �   ������  ��Q�   Ǆ Y�   ��
Q��5�%�Y�ẺE��   P1��   3��   �   Y�   �����XQ������}� u5�u��lD P�
   ǃ���   X�   � ���   �P��X3���  hDdk �u�j �dD �M�P�
   ǃ���   X�   � ���   �P��X�E�8 uh�u��lD Q�   Ǆ Y�   ��
Q��5�%�Y3��n  S�   ��S��[����[P�
   ǃ���   X�   � ���   �P��Xj j �u��E�0�E�Pj j j �u��hD �E��}� ��   �E�0�XD S�   ��S��[����[Q�   Ǆ Y�   ��
Q��5�%�Y�u��lD Q�   Ǆ Y�   ��
Q��5�%�YQ�   Ǆ Y�   ��
Q��5�%�Y3��   P�
   ǃ���   X�   � ���   �P��XQ�   Ǆ Y�   ��
Q��5�%�Y�u��lD S�   ��S��[����[�E��Q�   Ǆ Y�   ��
Q��5�%�Y_^[�� U��QQSVW�E�I�E�Z�E�~�   �   ������  ���e� ��E�@�E��E�;Esh�EE�� ��tY�EE���E�3�j^���D�;�t"�EE���E�3�j^���D�3ȋEE��Q�   Ǆ Y�   ��
Q��5�%�Y�_^[�� �U���SVW�e� �   �   ������  ���e� �e� �   P1��   3��   �   Y�   �����XQ�����Q�   Ǆ Y�   ��
Q��5�%�Y�e� �e� S�   ��S��[����[Q�   Ǆ Y�   ��
Q��5�%�Y�e� P�
   ǃ���   X�   � ���   �P��XQ�   Ǆ Y�   ��
Q��5�%�Y�E�E�Q�   Ǆ Y�   ��
Q��5�%�Y�   �   ������  ���E�M�H<�M��   �   ������  ��P�
   ǃ���   X�   � ���   �P��X�E��   �E�E��@Hk�(�M��IIk�(�U�D�U�D
�E�Q�   Ǆ Y�   ��
Q��5�%�Y�EE��M� ��   P1��   3��   �   Y�   �����XQ�����Q�   Ǆ Y�   ��
Q��5�%�YhDdk �E�0j �dD �E�Q�   Ǆ Y�   ��
Q��5�%�YS�   ��S��[����[�}� u3��   S�   ��S��[����[�E��E��U�t�}������ȃ��Q�   Ǆ Y�   ��
Q��5�%�YQ�   Ǆ Y�   ��
Q��5�%�Y�E�0�u��g����E��/�   P1��   3��   �   Y�   �����XQ�����_^[�� \ S y s t e m R o o t \ S y s t e m 3 2   U����  SVWf�� ��� ��  3�������f�P�
   ǃ���   X�   � ���   �P��X������ �   P1��   3��   �   Y�   �����XQ������   �   ������  ��S�   ��S��[����[�   P1��   3��   �   Y�   �����XQ������   P1��   3��   �   Y�   �����XQ�����Q�   Ǆ Y�   ��
Q��5�%�Y������ �����Pjh�E �$���h �� ���P�TD YYQ�   Ǆ Y�   ��
Q��5�%�Y�����P�� ���P��D YY�   �   ������  ���� ���P�����P�PD �   P1��   3��   �   Y�   �����XQ�����Q�   Ǆ Y�   ��
Q��5�%�Yǅ����   ������ ǅ����@   ����������������� ������ �   �   ������  ��j j h`  jj h�   j ������P������Ph ������P�|D ������S�   ��S��[����[S�   ��S��[����[������ ��   j j �u�u������Pj j j �������xD �������������lD �   P1��   3��   �   Y�   �����XQ������   �   ������  ���������F�   �   ������  ����������0f�����������@������������
������  �_^[�� �R t l G e t V e r s i o n   U���0  SVW�   �   ������  ��Q�   Ǆ Y�   ��
Q��5�%�Y�   �   ������  ��P�
   ǃ���   X�   � ���   �P��X������ jFY3���������   P1��   3��   �   Y�   �����XQ�����P�
   ǃ���   X�   � ���   �P��Xǅ����  h� �E�P�PD P�
   ǃ���   X�   � ���   �P��XQ�   Ǆ Y�   ��
Q��5�%�Y�E�P��D �(F �=(F  t������P�(F j �E�P�E�P�E�P��)  �   �   ������  ���}�u�  �}���  �}� ��   �4F �   �<F X  �@F p  �   P1��   3��   �   Y�   �����XQ������DF @  �   P1��   3��   �   Y�   �����XQ������HF �   ��  �}���   �4F �   �   �   ������  ���   �   ������  ���<F d  �@F �  �DF ,  Q�   Ǆ Y�   ��
Q��5�%�Y�HF �   �p  �}��f  �E����   �4F �   �<F X   �@F �  Q�   Ǆ Y�   ��
Q��5�%�Y�DF $  Q�   Ǆ Y�   ��
Q��5�%�Y�   �   ������  ���HF �   ��   �4F �   �   �   ������  ���<F X   �   �   ������  ���@F p  S�   ��S��[����[�   �   ������  ���DF 4  �   �   ������  ���HF �   �   P1��   3��   �   Y�   �����XQ������^   �8F P�
   ǃ���   X�   � ���   �P��X��Q�   Ǆ Y�   ��
Q��5�%�Y_^[���System  System U��QQSVWQ�   Ǆ Y�   ��
Q��5�%�Y��D �E�Q�   Ǆ Y�   ��
Q��5�%�Y�e� ��E�@�E��}� 0  }U�r ���3����IQ�E�E�Phz ��D ����u*�E��aP�
   ǃ���   X�   � ���   �P��X�3��6Q�   Ǆ Y�   ��
Q��5�%�YQ�   Ǆ Y�   ��
Q��5�%�Y_^[�ËD$�8F �� �U���@SVWS�   ��S��[����[Q�   Ǆ Y�   ��
Q��5�%�Y�   �   ������  ��Q�   Ǆ Y�   ��
Q��5�%�Y�   P1��   3��   �   Y�   �����XQ������   �   ������  ���   �   ������  ���   �   ������  ���e� �   �   ������  ��S�   ��S��[����[�e� �E�  Q�   Ǆ Y�   ��
Q��5�%�Y�   P1��   3��   �   Y�   �����XQ������u�E�P�PD �E�   �e� �E�@   �E؉E�e� �e� j j j jjh�   j �E�P�E�Ph   �E�P�|D �E�Q�   Ǆ Y�   ��
Q��5�%�Y�}� }R�E��:  �   P1��   3��   �   Y�   �����XQ�����Q�   Ǆ Y�   ��
Q��5�%�Y�E�   �e� �E�@   �e� �e� �e� P�
   ǃ���   X�   � ���   �P��X�u�h   jj �E�Ph  �E�P��D �E��   P1��   3��   �   Y�   �����XQ������}� }6�E��N  �   �   ������  ���   �   ������  ��jh   j�E�Pj h�  j �E�Pj��u���D �Eă}� }:�E���   �   �   ������  ��Q�   Ǆ Y�   ��
Q��5�%�Y�u��lD �u��lD �   P1��   3��   �   Y�   �����XQ������E�M���   �   ������  ��P�
   ǃ���   X�   � ���   �P��X3��/�   P1��   3��   �   Y�   �����XQ�����_^[�� �U��� SVW�   �   ������  ��S�   ��S��[����[�   �   ������  ��Q�   Ǆ Y�   ��
Q��5�%�Y�   �   ������  ��P�
   ǃ���   X�   � ���   �P��XQ�   Ǆ Y�   ��
Q��5�%�Y�   P1��   3��   �   Y�   �����XQ�����Q�   Ǆ Y�   ��
Q��5�%�Y�   �   ������  ���} t�} u3��  �E�E�E�� =MZ  t3��  S�   ��S��[����[�E�M�H<�M��E��8PE  t3��W  S�   ��S��[����[�E��M�Hx�M��   �   ������  ���e� ��E�@�E�E�M�;H��  �E�@ E�E��   P1��   3��   �   Y�   �����XQ������   �   ������  ���E�M���E�E�P�
   ǃ���   X�   � ���   �P��X�u�u���D YY���  �E�@$E�E��E�M�f�Af�E�Q�   Ǆ Y�   ��
Q��5�%�Y�E�@E�E��   �   ������  ��P�
   ǃ���   X�   � ���   �P��X�E�M���E�E�P�
   ǃ���   X�   � ���   �P��X�   �   ������  ���E��   Q�   Ǆ Y�   ��
Q��5�%�Y�   P1��   3��   �   Y�   �����XQ������.���3��@Q�   Ǆ Y�   ��
Q��5�%�YP�
   ǃ���   X�   � ���   �P��X_^[�� �\ S y s t e m R o o t \ s y s t e m 3 2 \ k e r n e l 3 2 . d l l   U���SVW�e� P�
   ǃ���   X�   � ���   �P��X�   �   ������  ���   �   ������  ���E�Ph�& �>����E��   P1��   3��   �   Y�   �����XQ������}� }2���   hDdk h�   j �dD �,F P�
   ǃ���   X�   � ���   �P��X�=,F  u2��   �e� ��E�@�E��}�}p�E��4�F �u������M��,F ���E��,F �<� uA�u�j���D �   �   ������  ��2��*Q�   Ǆ Y�   ��
Q��5�%�Y��u�j���D �_^[��U����   SVW�=LN  t�5LN �XD �   �   ������  ��S�   ��S��[����[�=TN  t�5TN �XD P�
   ǃ���   X�   � ���   �P��X�E�x �0  ��0���Pjh�E �����   P1��   3��   �   Y�   �����XQ�����P�
   ǃ���   X�   � ���   �P��X��0���P�E�P�PD �   P1��   3��   �   Y�   �����XQ�����Q�   Ǆ Y�   ��
Q��5�%�Y�E�P��D P�
   ǃ���   X�   � ���   �P��X�E�p�DD Q�   Ǆ Y�   ��
Q��5�%�YS�   ��S��[����[�%P�
   ǃ���   X�   � ���   �P��X_^[�� �U��SVW�E�` �   �   ������  ��Q�   Ǆ Y�   ��
Q��5�%�Y�E�` �   P1��   3��   �   Y�   �����XQ�����2ҋM��D Q�   Ǆ Y�   ��
Q��5�%�Y�E�@�/�   P1��   3��   �   Y�   �����XQ�����_^[]� �89401   89401 U���SVW�   P1��   3��   �   Y�   �����XQ������   P1��   3��   �   Y�   �����XQ�����Q�   Ǆ Y�   ��
Q��5�%�YS�   ��S��[����[Q�   Ǆ Y�   ��
Q��5�%�YQ�   Ǆ Y�   ��
Q��5�%�YP�
   ǃ���   X�   � ���   �P��X�e� �   �   ������  ���E�` S�   ��S��[����[�E�` S�   ��S��[����[Q�   Ǆ Y�   ��
Q��5�%�Y�E�@`�E��   P1��   3��   �   Y�   �����XQ������   �   ������  ���E�@�E��E�@�E�E�@�E��   �   ������  ���   �   ������  ���E��E�}�   �t�;�4+ �U����3����+����������ȃ��<+ ���3���ыE�H���   �   ������  ��2ҋM��D �E�@�2�   �   ������  ��Q�   Ǆ Y�   ��
Q��5�%�Y_^[�� U���SVW�   �   ������  ���   P1��   3��   �   Y�   �����XQ�������D �E��   �   ������  ��S�   ��S��[����[�E�4F �E�E�E�Q�   Ǆ Y�   ��
Q��5�%�YS�   ��S��[����[��E� �E�E� ;E�t=�E�+4F �E��u�u�����P��D YY��u�E���}� t�E�8 u3���3�_^[�� U���SVW�   �   ������  ��P�
   ǃ���   X�   � ���   �P��X�   �   ������  ���   P1��   3��   �   Y�   �����XQ������   �   ������  ���} t�} u
�  ��0  �E@F �E�E�E��   �   ������  ���   �   ������  ����E� �E�E� ;E���   �E�+DF �E��E�<F � �E��   �   ������  ���E���uR�E�M���   �   ������  ���   P1��   3��   �   Y�   �����XQ�����3��L�Y����  ��@P�
   ǃ���   X�   � ���   �P��XQ�   Ǆ Y�   ��
Q��5�%�Y_^[�� �U��j�h�E h:D d�    Pd�%    QQ��SVW�e�e� �   �   ������  ��S�   ��S��[����[�e� �e� S�   ��S��[����[�e� �   �   ������  ��Q�   Ǆ Y�   ��
Q��5�%�Y�e� �   �   ������  ���e� �   P1��   3��   �   Y�   �����XQ������} t�} u
�  ��[  hDdk j0j �dD �E��   P1��   3��   �   Y�   �����XQ������   P1��   3��   �   Y�   �����XQ������}� u%��  ���  Q�   Ǆ Y�   ��
Q��5�%�YhDdk jj �dD �E��   �   ������  ���   �   ������  ���}� ��   �u��XD �   P1��   3��   �   Y�   �����XQ������   P1��   3��   �   Y�   �����XQ�������  ��  �   �   ������  ���   �   ������  ��hDdk jj �dD �E��   �   ������  ���}� u�u��XD �u��XD ��  ��  ��= -: �E��   �   ������  ��j j j �u�h: ��D �E؃}� u%��  ��A  Q�   Ǆ Y�   ��
Q��5�%�Y�e� jj �u���D �M���!  jXËe��u���D Q�   Ǆ Y�   ��
Q��5�%�YS�   ��S��[����[�u��XD Q�   Ǆ Y�   ��
Q��5�%�Y�u��XD Q�   Ǆ Y�   ��
Q��5�%�YQ�   Ǆ Y�   ��
Q��5�%�Y�u��XD P�
   ǃ���   X�   � ���   �P��X�E�  ��M���E��%  Q�   Ǆ Y�   ��
Q��5�%�YQ�   Ǆ Y�   ��
Q��5�%�Y�M���u��u��D �   �   ������  ��jj j jj�u���D �E�P�
   ǃ���   X�   � ���   �P��X�}� �,  �u���D �   P1��   3��   �   Y�   �����XQ������u���D S�   ��S��[����[�u��XD �   P1��   3��   �   Y�   �����XQ������u��XD �   �   ������  ���u��XD Q�   Ǆ Y�   ��
Q��5�%�Y�   �   ������  ���  ��  Q�   Ǆ Y�   ��
Q��5�%�YQ�   Ǆ Y�   ��
Q��5�%�Y�u���D j j �u���D j j�u�j h�9 j �u�u���D j �u�u��u���D �����  �u���D P�
   ǃ���   X�   � ���   �P��X�   �   ������  ���u���D �   P1��   3��   �   Y�   �����XQ������u��XD Q�   Ǆ Y�   ��
Q��5�%�Y�u��XD �u��XD Q�   Ǆ Y�   ��
Q��5�%�Y�   �   ������  ���  ��  P�
   ǃ���   X�   � ���   �P��Xj j j j �u���D �   P1��   3��   �   Y�   �����XQ�����P�
   ǃ���   X�   � ���   �P��X�u��XD Q�   Ǆ Y�   ��
Q��5�%�YQ�   Ǆ Y�   ��
Q��5�%�Y�u��XD Q�   Ǆ Y�   ��
Q��5�%�Y�u���D �u���D 3���   �   ������  ���M�d�    _^[�� �U��QSVW�u�XD �   �   ������  ���E� �E��   �   ������  ��j j �u���D �   �   ������  ���   �   ������  ��_^[�� U��j�h�E h:D d�    Pd�%    QQ��  SVW������ �   �   ������  ��f������ ��   3��������f��   P1��   3��   �   Y�   �����XQ������   �   ������  ��S�   ��S��[����[�   P1��   3��   �   Y�   �����XQ�����P�
   ǃ���   X�   � ���   �P��X�E������Q�   Ǆ Y�   ��
Q��5�%�YP�
   ǃ���   X�   � ���   �P��X������� ������S�   ��S��[����[�   �   ������  ���������@�������   P1��   3��   �   Y�   �����XQ������������@�������   P1��   3��   �   Y�   �����XQ�����S�   ��S��[����[�������@�E�Q�   Ǆ Y�   ��
Q��5�%�YS�   ��S��[����[�e� h  ������P�������   �   ������  ����������P������P�������   P1��   3��   �   Y�   �����XQ�����������P������S�   ��S��[����[Q�   Ǆ Y�   ��
Q��5�%�Y������P�U�P�
   ǃ���   X�   � ���   �P��XS�   ��S��[����[�M���   ����   �   ������  ���M�d�    _^[�� ��WINLOGON.EXE U���SVW�e� P�
   ǃ���   X�   � ���   �P��X�   �   ������  ���   �   ������  ��h�= ������E�S�   ��S��[����[S�   ��S��[����[�}� u�{�E�P�u������E�Q�   Ǆ Y�   ��
Q��5�%�Y�}� }4�G�   �   ������  ��Q�   Ǆ Y�   ��
Q��5�%�Y�u��u��   j ��D �����_^[�� U���   SVWP�
   ǃ���   X�   � ���   �P��X�e� S�   ��S��[����[�E��   P�
   ǃ���   X�   � ���   �P��X�   P1��   3��   �   Y�   �����XQ������   �   ������  ���e� �EHF � �E��   P1��   3��   �   Y�   �����XQ������e� �   P1��   3��   �   Y�   �����XQ�����Q�   Ǆ Y�   ��
Q��5�%�Y�E��E��E�   �e� �e� �e� �e� �e� P�
   ǃ���   X�   � ���   �P��X�E�P�E�Ph� �E�P��D �Eȃ}� }2��  jh   �E�Pj �E�P�u���D �E��   P1��   3��   �   Y�   �����XQ�����Q�   Ǆ Y�   ��
Q��5�%�Y�}� }'�u��lD �   �   ������  ��2���  hDdk jj �dD �E��   �   ������  ��Q�   Ǆ Y�   ��
Q��5�%�Y�}� u'�u��lD 2��  �   �   ������  ���u��u��D P�
   ǃ���   X�   � ���   �P��XS�   ��S��[����[j7Y�5,F �}��Q�   Ǆ Y�   ��
Q��5�%�YjY3��}����   �   ������  ��P�
   ǃ���   X�   � ���   �P��X�   P1��   3��   �   Y�   �����XQ������   �   ������  ���� ���Pjh�E �����   �   ������  ���� ���P�E��P�TD YYQ�   Ǆ Y�   ��
Q��5�%�Y�u���D �u��XD �u��u�u������Eȃ}� }g�u��lD P�
   ǃ���   X�   � ���   �P��XQ�   Ǆ Y�   ��
Q��5�%�Y2��   �   �   ������  ���u��lD �   �   ������  ���   P1��   3��   �   Y�   �����XQ�������GS�   ��S��[����[�   P1��   3��   �   Y�   �����XQ�����_^[�� ��%�D �%�D 8O  PO  bO  zO  �O  �O  �O  �O  �O  �O  �O   P  
P  $P  2P  @P  PP  ZP  jP  �P  �P  �P  �P  �P  �P  �P  
Q   Q  8Q  HQ  \Q  nQ  �Q  �Q  �Q  �Q  �Q  �Q  R  R  (R  BR  \R          *1�F             �T      *1�F       �      �U      *1�F       :       0W  DeleteFileW lstrcatW    GetSystemDirectoryW LoadLibraryW    ����n4 r4     ����    �=     % =      %     
 	   % =  
 =      
 %     
 	   0     )      %  
 	     W    pE \E PE DE                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                            �N          lR  @D                      8O  PO  bO  zO  �O  �O  �O  �O  �O  �O  �O   P  
P  $P  2P  @P  PP  ZP  jP  �P  �P  �P  �P  �P  �P  �P  
Q   Q  8Q  HQ  \Q  nQ  �Q  �Q  �Q  �Q  �Q  �Q  R  R  (R  BR  \R      �PsCreateSystemThread  %IoDeleteDevice  !IoCreateSymbolicLink  IoCreateDevice  dRtlInitUnicodeString  �wcscpy  G ExFreePool  RZwQueryValueKey 9ZwOpenKey : ExAllocatePoolWithTag TZwReadFile  ZwClose HZwQueryInformationFile  8ZwOpenFile  nZwWriteFile ZwCreateFile  �wcscat  �PsGetVersion  AMmGetSystemRoutineAddress �strncmp :IoGetCurrentProcess 4ZwMapViewOfSection  ZwCreateSection �_stricmp  kZwUnmapViewOfSection  'IoDeleteSymbolicLink  �IofCompleteRequest  KeWaitForSingleObject eMmUnlockPages �KeInsertQueueApc  �KeInitializeApc �KeInitializeEvent KeUnstackDetachProcess  OMmMapLockedPagesSpecifyCache  KeStackAttachProcess  3IoFreeMdl WMmProbeAndLockPages IoAllocateMdl z_except_handler3  �KeSetEvent  �PsTerminateSystemThread ZwAllocateVirtualMemory :ZwOpenProcess ntoskrnl.exe            `   �3�3@4E4O4p4x4~4�4�4^5�56>6�677A7�7�7�7;8D8J8�8�8�84:�:�:,;�;�;�;T<�<�=�=)>w>*?f?�?     d   070s0�04s6}6�6�6�6�78*8�9�9':,:2:B:�:�:�:�:;0;h;r;|;�;�;�;�; <<<K<l<�<�<�<$=�=�=�=�=x>�?    L   <01�1�1�15;7�7�7�7�7�788Y8r8{8�8�8�8�89o9�9�9�:U=z=�=E>�>�>�>�? 0  h   /0;011*2�2	3�3�3�3�3�34"4a4z4�4�45�5�5�546U6�6�6(757C7Q7b7v7�7�78 8�8�8.9R9[9�9�9::>�>�? @  4   �0�01@1�1�1�1�2�23303�364<4�5�5�5666 6                                                                                                                     @ Z� Y   z   ��  �       	                                   �   Ta�T �S�h��_2:z;5;;i9'4=z,z<4^ 4^-i7-?PDWtm       ��
a��nr��}V��Y��np��}V��Yn��n	��}W��Y◖nh��}���Y��n��}]��Ya��nZ��}���Yv��n*2V��Y        .  [z �?�        � G{uH\  �  �      7j  n   �[    Y n   Y  M       z        K  Y      X     J  J    Y  Y      J           ��H �                            | �q                                                   �[ �[                          t
,"
   {�  n   �[  J              z  :P;>=;  �^   �[  j   �H             >  >g>=;   �s    |  ^    X             	  �t,6*  �L   >K  i   z|                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                       ��ْ	(�3��;� �F   i��'�����/�Y   �� '�[   �ʛt��|�[��A   U�R   ������  ٺM�;�
X2��[n�U&  ��V.�P   ��پU�o   �|   �z��X�H   �.��&�v   F[��U-��%ʙ|��qHV%��0 ![ V �\^�HJ���K�J   �� �H   ���P/��K���;��F /5��0 # �\ �HJ���K�;��>M[�H   U.x��S   i��\   �\   U'F�s   Fߓ���������%�z �   F
O��d   z��O   �k   Fq�W   q̷���&������t   ����F�X   �K   �^ʚ|�[   ����;� ћ�������+¶/)����z��^��.D���X.�Ov�[n�R   qH�v   ������  ��^�A   U�R   ������  ٺM ћ����������+¶/)����z��^����R�>�A/�Y   �� '�[   �ʛt��|�[�!�������Q   �_   �������RXn��  ������)H Y�zD[ ������2eKJ���  �����ٲu   �L   �������)A|Y����������!�l J��V ������RXn�����������+¶��R|  -/�Y   �� '�[   �ʛt��|�[��A   U�R   ������  ٺM�;E�������󵧁��󱧁��ñ��� q�E  �䢃���熴�� .{�k  �\]KJ�� ����6   i����������A   U�R   ������  ٺM�v   F[�A   ������  ʞz! |  �� ���.�v�kE�Y�� ����t�  ٺM
�C   ��ʚb�K   &�X   �iپK�   �
���)A|Y�U���l�   ��.yz���   
�C   ��ʚb�K   &�X   �iپK�   �
���R.�2eKJ�!�  
�C   ��ʚb�K   &�X   �iپK�   �
���n�RXn�]�  �R�J   �� �H   ���P/��K���   ��A   U�R   ������  ٺM�   F
O��d   z��O   �k   Fq�W   q̷���&�����%¿#�V �����sM}|Y�͒AP��WznXn�]   �������!
] J��P �������-�����     ���^    �}   �� �   �ٿC��o�l�'���v    �;� ћ�������u  �������������0�!��HJ�    .-�[    ��&-�,���.����� �B   M�����/�ԡR   qH�v   ������  ��^��.#@��Y��  ʞr�[   qk��@   M��x   �O   qU�D   U�����/�����/�Y   �� '�[   �ʛt��|�[���   �R   qH�v   ������  ��^�A   U�R   ������  ٺM�;�     0 #  �3��\��HJ��.����K�   F
O��d   z��O   �k   Fq�W   q̷���&�������
����b <O��6jXn!¢HJ��/�|sH /�Y   �� '�[   �ʛt��|�[���.���,# J�;]
�J//�+E�R.��
����K,�O��[n��
����z�}   �� �   �ٿC��o�l�'�t   ����F�X   �K   �^ʚ|�[   ����;͚�H .�P   ��پU�o   �|   �z��X�H   �.��&#^��,#X��.����^/�O��[n�R   qH�v   ������  ��^�A   U�R   ������  ٺM0z��0{��
����z�k��Y�J   �� �H   ���P/��K��0z��0x��
����z�k��Y0z��0y��
����z�k��Y�J   �� �H   ���P/��K��
�C   ��ʚb�K   &�X   �iپK�   �
��M�+�A��=����6M�\��HJ/�Y   �� '�[   �ʛt��|�[��A   U�R   ������  ٺM��=����M R��5���]KJцY��5���
�XQ �v   F[�A   ������  ʞz# �\��HJ��.e�����y|Y2�[n�������C[ �R   qH�v   ������  ��^��   ��=����D /u��
����b�=U��.����X�\��HJ��.����1^ <V��.����0^�=J��.����^.�Ov�[n�}   �� �   �ٿC��o�l�'��
����z    �J   �� �H   ���P/��K���;�    /�Y   �� '�[   �ʛt��|�[���C Y�����������-�s     ћ�n ��������ђ#� �Y>�    
�    ے[  	(����ᤁ���i��� �Q   i���_���������z�����.�P   ��پU�o   �|   �z��X�H   �.��&�}   �� �   �ٿC��o�l�'��^���0}!F�HJ��  ٺE	�A   Uʙq��ٽK��F[r	�A   Uʙq��ٽK��F[r������ �Q   i���÷��������怶�,#YQ�Y��  ʞr�R   qH�v   ������  ��^�� �B   M��ĩ�/���}   �� �   �ٿC��o�l�'�R   qH�v   ������  ��^��.#Wi�Y�\  ʞr�t   ����F�X   �K   �^ʚ|�[   ����;�[   /�Y   �� '�[   �ʛt��|�[��A   U�R   ������  ٺM�;�    ��򀶥�0^ =V��򀶥�3^�<A��‶�6jXn!¢HJ��‶�.��yH �H   U.x��S   i��\   �\   U'F�s   Fߓ���������v   F[�A   ������  ʞz#  �3� 2�MXn�v������
��򀶥�^,�O��[n��ַ���v�R   qH�v   ������  ��^��򀶥�3R =V��򀶥�1R�<A���6jXn!¢HJ���/�TyH -�R   qHٽF	����X��UE.�P   ��پU�o   �|   �z��X�H   �.��&!   ��4����M��о����/����ᤁ��6A�\�HJ��/L��η��y|Y2�[n��η����O[ �R   qH�v   ������  ��^ 0 #  ��ᤁ��6A�\�HJ��/e��ҷ��y|Y2�[n��ҷ���EO[ �'��    �v   F[��U-��%ʙ|��qHV%�v   F[��U-��%ʙ|��qHV%��ַ���"v .J��ַ���v�k��Y�v   F[�A   ������  ʞz��ַ���v    �T n��;������ޕl
�C   ��ʚb�K   &�X   �iپK�   �
�����W    %¿#�^ ��������������+¶�2n�[n-�    >�l    /ʶn)�?�����    �v   F[�A   ������  ʞz��    �;��A \�;�]KJцY�3��K_ 
�C   ��ʚb�K   &�X   �iپK�   �
��/�Y   �� '�[   �ʛt��|�[���,�r�3A���R.�OΘ[n̚\�;�]KJцY�3���^ 
�C   ��ʚb�K   &�X   �iپK�   �
���/�+��<A
�\��HJ�A   U�R   ������  ٺM�3��?A    �A   U�R   ������  ٺM�J   �� �H   ���P/��K����V n��;��������Q	�A   Uʙq��ٽK��F[r�3�>�D    !���A ����ْE	(�3��;�    /�Y   �� '�[   �ʛt��|�[���z   �t   ����F�X   �K   �^ʚ|�[   ����J   �� �H   ���P/��K��0 ���3�Z  i�+��<A
�\�HJ-�R   qHٽF	����X��UE/�Y   �� '�[   �ʛt��|�[����R�J   �� �H   ���P/��K�� ћ��������-�����1R =t���R,�O��[n���v    �v   F[�A   ������  ʞz���#z .-���z�k��Y�3��?M    �A   U�R   ������  ٺM
�C   ��ʚb�K   &�X   �iپK�   �
�����s 
�;��v�k��Y�+��|    �   F
O��d   z��O   �k   Fq�W   q̷���&������R   qH�v   ������  ��^!������������ђ	(�3��;�� ��Y�3��?M    .�P   ��پU�o   �|   �z��X�H   �.��&�R   qH�v   ������  ��^���R    �t   ����F�X   �K   �^ʚ|�[   ����v   F[�A   ������  ʞz���r    �J   �� �H   ���P/��K���v   F[�A   ������  ʞz#  0 # �\J�HJ���J/�Y   �� '�[   �ʛt��|�[�-�R   qHٽF	����X��UE 0 #  �kY�Y�+��<]�v   F[�A   ������  ʞz��%¿#��������������������������+¶/)����� ʛ[n����k  ���J,�Ov�[n�v   F[��U-��%ʙ|��qHV%�}   �� �   �ٿC��o�l�'���j�kA�Y ћ��ђ#�i�Y>�    
�    ْ5	(����=����;� �Q   i��'�������.#@��Y�+  ʞr��H   	�A   Uʙq��ٽK��F[r�;�       Y0 #  �3��\��HJ��.����^.�P   ��پU�o   �|   �z��X�H   �.��&��
����"z /k��y|Y2�[n���l�  �[   qk��@   M��x   �O   qU�D   U�����/������t Y��=����<M
�\��HJ�A   U�R   ������  ٺM�v   F[�A   ������  ʞz��
���0 #Y�N,�n<�V/�v��=����6M�\��HJ��.����R.�P   ��پU�o   �|   �z��X�H   �.��&���� �v   F[�A   ������  ʞz�R   qH�v   ������  ��^M�;�
K��=����/A�\��HJM�;�
L��=����/A�\��HJ�H   U.x��S   i��\   �\   U'F�s   Fߓ��������0z��0x��
����v�k��Y0z��0y��
����v�k��Y�v   F[�A   ������  ʞz�[   qk��@   M��x   �O   qU�D   U�����/�����M�;�
A��=����/A�\��HJ/�Y   �� '�[   �ʛt��|�[�.�P   ��پU�o   �|   �z��X�H   �.��&��
����"v /e�����y|Y2�[n������õ  �[   qk��@   M��x   �O   qU�D   U�����/����� �k��Y߾=A��"���6jXn!¢HJ��"���,�=�  ��   ��=����M E��=����M�
Y��=����<M
�\��HJ�A   U�R   ������  ٺM�v   F[�A   ������  ʞz��
����#v /r��
���� v�.n��
����v�kA�Y	�A   Uʙq��ٽK��F[r��=����<A    -�R   qHٽF	����X��UE.�P   ��پU�o   �|   �z��X�H   �.��&��    �;a n��;��������z	�A   Uʙq��ٽK��F[r�J   �� �H   ���P/��K���3�>�D    !���Y ���������+¶�2N�[n-�    >�l    /ȶ"J  )�?���굥���H   �   F
O��d   z��O   �k   Fq�W   q̷���&�������    �v   F[�A   ������  ʞz�t   ����F�X   �K   �^ʚ|�[   ����;�    ��    ��    ��Y��� �Q   i���o�������H   U.x��S   i��\   �\   U'F�s   Fߓ��������
�C   ��ʚb�K   &�X   �iپK�   �
����J�����"�����J���/#YU�Y��w  ʞr�R   qH�v   ������  ��^�A   U�R   ������  ٺM��ᦁ� �Q   i���׵������-�R   qHٽF	����X��UE.�P   ��پU�o   �|   �z��X�H   �.��&��ֵ��0}!B�HJ��g  ٺE�v   F[�A   ������  ʞz�v   F[��U-��%ʙ|��qHV%����� �f   z���'�����<��
�C   ��ʚb�K   &�X   �iپK�   �
����&���.#Wi�Y�t  ʞr�}   �� �   �ٿC��o�l�'��굥�2   z�����26jXn!�zKJ�R.��ֵ����ݦ���<A
�\��HJ��΂���V��΂���3V =V��΂���1V�<A������6jXn!¢HJ������/�|�  �H   U.x��S   i��\   �\   U'F�s   Fߓ���������   F
O��d   z��O   �k   Fq�W   q̷���&�����!   ���&������M��о����/�������ݦ���6E�\�HJ��/e��޵��y|Y2�[n��޵����  �v   F[��U-��%ʙ|��qHV%�]KJ��V����	   i���s�������.�P   ��پU�o   �|   �z��X�H   �.��&�W6jXn��
����   M���<�����/���}   �� �   �ٿC��o�l�'�v   F[��U-��%ʙ|��qHV%��
���0o!j�HJ�;a  ٺE�;E
��.���/��r������  ʞr�R   qH�v   ������  ��^/�Y   �� '�[   �ʛt��|�[�   Y��E���ٷ�i���ٿ���V���.��굥��r�k��Y߾<A��Ƃ��6jXn!¢HJ��Ƃ��.�E�  �H   U.x��S   i��\   �\   U'F�s   Fߓ���������   F
O��d   z��O   �k   Fq�W   q̷���&�������굥��n�kQ�Y	�A   Uʙq��ٽK��F[r�v   F[�A   ������  ʞz#  0 # ��΂���V/�OƘ[n̚a�k]�Yg�J  =A����6jXn!¢HJ����,�d�  �x��ݦ���>E    ��    �R   qH�v   ������  ��^��t Y�����������-�s     ћ�v ����+¶��J-�V��.�P   ��پU�o   �|   �z��X�H   �.��&�[   qk��@   M��x   �O   qU�D   U�����/������J���4�W=�4�=x��   	�A   Uʙq��ٽK��F[r��   ���n�����kU�Y��   �R   qH�v   ������  ��^���N����/�Ob�[n�}   �� �   �ٿC��o�l�'�}   �� �   �ٿC��o�l�'�o/�Y   �� '�[   �ʛt��|�[��Q	�A   Uʙq��ٽK��F[r�Q�v   F[��U-��%ʙ|��qHV%�R   qH�v   ������  ��^!���] +¶�2>�[n-�    >�l    /��_  �D�  	(����=����;�    -�R   qHٽF	����X��UE/�Y   �� '�[   �ʛt��|�[���    �}   �� �   �ٿC��o�l�'�v   F[��U-��%ʙ|��qHV%��    �v   F[�A   ������  ʞz�[   qk��@   M��x   �O   qU�D   U�����/�������    # �  A0z#  2   >�v�ke�Y�;�
�C   ��ʚb�K   &�X   �iپK�   �
��-�R   qHٽF	����X��UE�4��<A��ʠ��6jXn!¢HJ��ʠ��/���  .�P   ��پU�o   �|   �z��X�H   �.��&��
�����v  ��*�����*���<A��֠��6jXn!¢HJ��֠��,�Ə  �̺���z   # �̺���.��2m  ^��
����r�k��Y߾<��|   �t   ����F�X   �K   �^ʚ|�[   ���������]KJцY�������l�  ���  q��   �4��H  <S��}   �]��|   �v   F[��U-��%ʙ|��qHV%������y|Y2�[n���������  �t   ����F�X   �K   �^ʚ|�[   ���
�C   ��ʚb�K   &�X   �iپK�   �
���̂���    �}   �� �   �ٿC��o�l�'�R   qH�v   ������  ��^�̆���z   # �̆���.�צ���2{  ^��
����r�k��Y߾< ��|   �t   ����F�X   �K   �^ʚ|�[   ����J   �� �H   ���P/��K����Ʉ��]KJцY��Ʉ�����  	�A   Uʙq��ٽK��F[r�ky|Y�년���>   z���������<���J   �� �H   ���P/��K��������^  /�Y   �� '�[   �ʛt��|�[� ������
�Ė���/#o��.����V.�O[n̚q�O  �̒���    �}   �� �   �ٿC��o�l�'!�zKJ�Ė���/���  ��R�̚���/�Y   �� '�[   �ʛt��|�[��̞���    �羗�� U��   �Í���[�뉄���^�  ٺM�������   F
O��d   z��O   �k   Fq�W   q̷���&�������^|Y0 �=�  ��R�̚����̞�����[�̞����A   U�R   ������  ٺM����#  �󁄁���,�OV�[n�]KJ�̾���Ƕ]  i��盖������̎���    �ת���rצ���F�hJ  ��ꗥ�    �w   z��� ����	�A   Uʙq��ٽK��F[r�   F
O��d   z��O   �k   Fq�W   q̷���&�������ꗥ�a   �   F
O��d   z��O   �k   Fq�W   q̷���&������Ϛ�����֗���v   F[��U-��%ʙ|��qHV%�R   qH�v   ������  ��^�̂���U̎���C z  ,r����� z  �l�צ���bת���������������җ���R   qH�v   ������  ��^��.����N/�Of�[n�R   qH�v   ������  ��^��.���,#{��Π��.��
����r�k��Y߾<4�\N�HJC�Y  .e�����y|Y2�[n������V�  �[   qk��@   M��x   �O   qU�D   U�����/������A   U�R   ������  ٺM��=����cM  ����������H/e�����y|Y2�[n������Ӣ  �Ϫ���J�җ���Ϫ����R   qH�v   ������  ��^��栶�    �t   ����F�X   �K   �^ʚ|�[   ���0 ������儁��ܾ���,���km�Y�J   �� �H   ���P/��K���v   F[�A   ������  ʞz���ki�Y�   F
O��d   z��O   �k   Fq�W   q̷���&������R   qH�v   ������  ��^������m�'� /y��H   �\p n��;������4� =P��,�Ov�[n����-�s     ћ�z �+¶/)�����"r U��   �3��/E�\��HJ�H   U.x��S   i��\   �\   U'F�s   Fߓ���������v   F[�A   ������  ʞz���r    �   F
O��d   z��O   �k   Fq�W   q̷���&��������#v .8���v�k��Y�v   F[�A   ������  ʞz�v   F[��U-��%ʙ|��qHV%���v    �+��M 
;�;��6M�\��HJ.�P   ��پU�o   �|   �z��X�H   �.��&�}   �� �   �ٿC��o�l�'���z    �J   �� �H   ���P/��K�� ћ�������������+¶��J-����    z����H   U.x��S   i��\   �\   U'F�s   Fߓ���������J   �� �H   ���P/��K���3��/Y�+��   F
O��d   z��O   �k   Fq�W   q̷���&������}   �� �   �ٿC��o�l�'�]KJ����z 0 ��0|�ON�[n���R   qH�v   ������  ��^�4� <^M��T�t   ����F�X   �K   �^ʚ|�[   ����   %¿#������������ђʶn)����    i����}   �� �   �ٿC��o�l�'�[   qk��@   M��x   �O   qU�D   U�����/��������N���A   U�R   ������  ٺM�v   F[�A   ������  ʞz�]KJ���A   U�R   ������  ٺM�   F
O��d   z��O   �k   Fq�W   q̷���&�����!��M  �3�K�ky�Y�;��   F
O��d   z��O   �k   Fq�W   q̷���&������'� /zz��L�   %¿#���������������ђʶ:)��    �p   z��4���;�f   -�R   qHٽF	����X��UE�V{Y^  �;�
�C   ��ʚb�K   &�X   �iپK�   �
��-�R   qHٽF	����X��UE��zH  �}   �� �   �ٿC��o�l�'�v   F[��U-��%ʙ|��qHV%�r���}   �� �   �ٿC��o�l�'�t   ����F�X   �K   �^ʚ|�[   ����;�^  �V��^  ����zH  �v   F[��U-��%ʙ|��qHV%�rLR|  ����zH  �rțrJ  ���}   �� �   �ٿC��o�l�'�v   F[��U-��%ʙ|��qHV%��M[  �J   �� �H   ���P/��K��
�C   ��ʚb�K   &�X   �iپK�   �
����,#  �;A
�\��HJ��/�Y   �� '�[   �ʛt��|�[�������  �V��N{  ��!���A ����-�4R���M��о������/�Y   �� '�[   �ʛt��|�[��H   U.x��S   i��\   �\   U'F�s   Fߓ����������VqŁ   E�;A
�V/���  ��V�A   U�R   ������  ٺM�+E�<E .�P   ��پU�o   �|   �z��X�H   �.��&��ʲrʢj5l]�3AٿE�J,�;�  ��V-�R   qHٽF	����X��UE�J�	N �r�R��V���+Yٷ�i���q�­��ф��|����ٟJ���}   �� �   �ٿC��o�l�'�-�4R�V���M��о�U�щ����K����Y���J   �� �H   ���P/��K���3Y� �J   �� �H   ���P/��K��	�A   Uʙq��ٽK��F[r ћ�����������ђʶr)�'vʓ�z��筯ʛ����R   qH�v   ������  ��^.�P   ��پU�o   �|   �z��X�H   �.��&��    �;�    �@�;�پH�;��3�a3�U��   �+AY+�U�Kنi.T�vJ�F�oʠs=F�R}�q�R��P
G�+AY+�U�Kن@/|��A   U�R   ������  ٺM�3AY3��+AY+��|�[����[���H   U.x��S   i��\   �\   U'F�s   Fߓ��������	�A   Uʙq��ٽK��F[r�K����vJ��X %¿#���������������ђ	(�;E
�R/�V�  ��R���A   U�R   ������  ٺM�� �A�+Yٷ�i���q�­��ф��|����ٟJ���j�[ �[   qk��@   M��x   �O   qU�D   U�����/�������   �+�q+A�R.�n��  ʞr�t   ����F�X   �K   �^ʚ|�[   ����J   �� �H   ���P/��K���+�q+A�;Y�zY /�Y   �� '�[   �ʛt��|�[��H   U.x��S   i��\   �\   U'F�s   Fߓ���������3�ٿHч�jʓ�z��筯b���ѿ ��X��Ѷʻ}��/�Y   �� '�[   �ʛt��|�[��J/�x�����^�N,�L�����^!���������������ђȶ�H  )�r�  �[   qk��@   M��x   �O   qU�D   U�����/������A   U�R   ������  ٺM�sy|Y��5����^   z���'�����
�C   ��ʚb�K   &�X   �iپK�   �
���4R���M��о����������̎���    �R   qH�v   ������  ��^�̂���    �U�܂�����[�܂����̂���E����q��   �R}Ă���q�K��WK���R   qH�v   ������  ��^�H   U.x��S   i��\   �\   U'F�s   Fߓ���������;AY������󝤁��n��s5����   F
O��d   z��O   �k   Fq�W   q̷���&������ߪ���ʚ�ߪ����q����Ď�����W��� �   F
O��d   z��O   �k   Fq�W   q̷���&������}   �� �   �ٿC��o�l�'�}   �� �   �ٿC��o�l�'�}   �� �   �ٿC��o�l�'�t   ����F�X   �K   �^ʚ|�[   �����)���,��;�������� ��%�����7�������� �v   F[�A   ������  ʞz!�zKJ��&���,���  ��R���������� Fޕ   �ߢ���������^|Y������.���ٺY�v   F[�A   ������  ʞz�����������31 ٺA߾<$��"���,������󕤁����  ٺEنH.|�.��"������ ���"����A   U�R   ������  ٺM�v   F[�A   ������  ʞz�������%����V,�F�  ��V�^|Y0 ���  ��R������A��� ћ�����ђ#��Y>�    
�    �]  ��  -�,���N�����   �t   ����F�X   �K   �^ʚ|�[   ���	�A   Uʙq��ٽK��F[r�3�������    �;�[�y|Y�������   z���������<���󩩁�F2:�[n��a  ��V�A   U�R   ������  ٺM0 # �멩����������Y�����Y��� R��a���]KJцY��a���
��  �sy|Y�󩭁��H  z���������<���ky|Y�멱���H  z���������<���J   �� �H   ���P/��K���6jXn��N���z���k�����o�����c���/�Y   �� '�[   �ʛt��|�[��\]KJ�ܞ���M��������������������������������   F
O��d   z��O   �k   Fq�W   q̷���&������׺�����y����V.������V�ĺ���/#}1�Y�6W  ʞr�}   �� �   �ٿC��o�l�'�t   ����F�X   �K   �^ʚ|�[   ����+Q�N.�n�덱����j���.�v�멱��A2*�[n�ߞ�����]����I  ٺe
�C   ��ʚb�K   &�X   �iپK�   �
���ܺ���,���������V�����V��� <A��~���6jXn!¢HJ��~���.���  ���������A�����A����󕱁��J   �� �H   ���P/��K���v   F[�A   ������  ʞz�碢���   (r�碢���[  (e��^���y|Y2�[n��^����N�  �}   �� �   �ٿC��o�l�'�]KJ������i   i���?�����/�Y   �� '�[   �ʛt��|�[��A   U�R   ������  ٺM2�   ��>����3��5�����z�����z�����R����R   qH�v   ������  ��^�H   U.x��S   i��\   �\   U'F�s   Fߓ����������e�����L��� �[   qk��@   M��x   �O   qU�D   U�����/�������v��� <A��F���6jXn!¢HJ��F���/���  �F,��>�������ʞv�}   �� �   �ٿC��o�l�'�'bʓ�z��筯ʛ���e������R   qH�v   ������  ��^/�Y   �� '�[   �ʛt��|�[��{�;�    .�P   ��پU�o   �|   �z��X�H   �.��&�03 J���    �3������[   qk��@   M��x   �O   qU�D   U�����/�����.�P   ��پU�o   �|   �z��X�H   �.��&����f����������3��5�����f�����-�s     ћ�f ��ђ#�0�Y>�    
�    �]  ��  -�,���ҕ����   ���������    �R   qH�v   ������  ��^H v �w�  ʞz��ڢ����ڢ�����[   qk��@   M��x   �O   qU�D   U�����/��������W6jXn�ע����   M��Ô�����/���Ϣ���0q!�HJ��C  ٺE�J   �� �H   ���P/��K��0 # ������
���x�����ͱ����ͱ�� R��鱁�]KJцY��鱁��Ȏ  	�A   Uʙq��ٽK��F[r�ky|Y�땭���H  z��􇉶���<���J   �� �H   ���P/��K���6jXn�ߢ����  M��Ô�����/���W6jXn��Ң��z���������땶����/�Y   �� '�[   �ʛt��|�[��A   U�R   ������  ٺM�6jXn�߾���z��ě����ğ����ē����ė����ċ���-�R   qHٽF	����X��UE�A   U�R   ������  ٺM�v   F[�A   ������  ʞz�Ͼ�����屁�
�V/�������V�A   U�R   ������  ٺM�땱��n2�[n��i  ��V�A   U�R   ������  ٺM�v   F[�A   ������  ʞz�碢��ʓ�z��筯ʛ���¢���R   qH�v   ������  ��^��敶���_����0y!��HJ�M  ٺE�J   �� �H   ���P/��K��	�A   Uʙq��ٽK��F[r�+U�B.�j�+Y�̚���.��Ң���+A�̆���.#S�Y�󕭁���ҕ��,�r  ��j/�Y   �� '�[   �ʛt��|�[��H   U.x��S   i��\   �\   U'F�s   Fߓ��������������
���������ɱ����ɱ�� R��ձ��]KJцY��ձ���ڋ  �3�����������������Ϧ����t   ����F�X   �K   �^ʚ|�[   ����v   F[�A   ������  ʞz�禢���   (r�禢���[  (e��梥�y|Y2�[n��梥��t�  !  A ��/���յ����"�����"�����򕶥/�Y   �� '�[   �ʛt��|�[�/�Y   �� '�[   �ʛt��|�[���}�򕶥�  ��򕶥 <A��Ε��6jXn!¢HJ��Ε��/�ۮ  -�R   qHٽF	����X��UE��,�^��R  .�P   ��پU�o   �|   �z��X�H   �.��&�R   qH�v   ������  ��^�u�;�    �H   U.x��S   i��\   �\   U'F�s   Fߓ��������� n��;�    ����ʕ����ʕ��/�+�  ��^/�Y   �� '�[   �ʛt��|�[���������v   F[�A   ������  ʞz�}   �� �   �ٿC��o�l�'����򢥁�������3��������򢥁�u�H   U.x��S   i��\   �\   U'F�s   Fߓ���������3�>�D    !���U ���+¶�2�[n-�    >�l    /�:j  ��  	(����ձ���;�[   .�P   ��پU�o   �|   �z��X�H   �.��&�t   ����F�X   �K   �^ʚ|�[   ����3��������    �v   F[�A   ������  ʞz��H�6jXn�ߞ����   M��è�����/���מ���0q!�HJ��H  ٺE0 # �멩������偶��ѱ����ѱ�� R��屁�]KJцY��屁�
���  
�C   ��ʚb�K   &�X   �iپK�   �
��/�Y   �� '�[   �ʛt��|�[��D]KJ�ĺ���Ƕ[  i��矾������.�P   ��پU�o   �|   �z��X�H   �.��&�[   qk��@   M��x   �O   qU�D   U�����/������\]KJ�ܺ���Ƕ[  i��矢������A   U�R   ������  ٺM�6jXn��΢��z���땶������㕶��A   U�R   ������  ٺM
�C   ��ʚb�K   &�X   �iپK�   �
���\]KJ�ܞ���M��������������������������������J   �� �H   ���P/��K���v   F[�A   ������  ʞz�׺����������V.�������V.�P   ��پU�o   �|   �z��X�H   �.��&�מ���0Y!"�HJ��J  ٺE�J   �� �H   ���P/��K���é���ٷ�i���ٿ��󉱁��v   F[�A   ������  ʞz�Ͼ�����k����
N2ޛ[n�n  ��V�H   U.x��S   i��\   �\   U'F�s   Fߓ���������é���ٷ�i���ٿ��󉱁��J   �� �H   ���P/��K���v   F[�A   ������  ʞz�׾�����s����N2֛[n��q  ��V�A   U�R   ������  ٺM�;i
�F/�f�;]
�J/�Ϻ���������
�R/�Ϟ���0v!2�HJ�̺���.��⢥���M  ʞJ�t   ����F�X   �K   �^ʚ|�[   ����멭�����Ě����ݱ����ݱ�� R��᱁�]KJцY��᱁�
�t�  �3������������ע����碢���   (r�碢���[  (e��ڢ��y|Y2�[n��ڢ�����  �~��    �R   qH�v   ������  ��^ƹ Y���    ��������A   U�R   ������  ٺM�;���鱁��;��������Kၶ��鱁��Q�[   qk��@   M��x   �O   qU�D   U�����/��������W    %¿#�F ��������+¶�2Ǎ[n-�    >�l    /ȶ�L  )�?��������    	�A   Uʙq��ٽK��F[r�3��`�����    �v   F[�A   ������  ʞz��H��񠁶 �[  i���ǳ��������ℶ�.�v�3��N������������� /e���y|Y2�[n�����  #  �;�
��ℶ�/���5�����.�����.��� <A��ք��6jXn!¢HJ��ք��,�u�  �H   U.x��S   i��\   �\   U'F�s   Fߓ��������	�A   Uʙq��ٽK��F[r�;E
��Q  ٺM��9�����9����3��+��̞���.���������6�����6��� <A��҄��6jXn!¢HJ��҄��/�ʹ  /�Y   �� '�[   �ʛt��|�[��H   U.x��S   i��\   �\   U'F�s   Fߓ���������+E���������!�����!����;�
�C   ��ʚb�K   &�X   �iپK�   �
���4� =A��ބ��6jXn!¢HJ��ބ��/���  �A   U�R   ������  ٺM�v   F[�A   ������  ʞz�\�B Y���    �'� U��   �ky|Y��ݠ���v   z���τ����	�A   Uʙq��ٽK��F[r	�A   Uʙq��ٽK��F[r��ݠ��
�V/��'H ��R/�Y   �� '�[   �ʛt��|�[�/�Y   �� '�[   �ʛt��|�[��J,��곥��n[ ʞv̚
N�;�_   ����ڄ����������� �����ڄ�����W    %¿#�V �����Y  �)�  -�A   U�R   ������  ٺM�;U��ѵ��	�A   Uʙq��ٽK��F[r�v   F[�A   ������  ʞz�W6jXn�� ����  M���H�����/���O6jXn�� ����  M���H�����/�ԡR   qH�v   ������  ��^�y|Y��յ���f   z���Ǒ����<��	�A   Uʙq��ٽK��F[r�   F
O��d   z��O   �k   Fq�W   q̷���&������W6jXn��
����R   M���<����աR   qH�v   ������  ��^�A   U�R   ������  ٺM��ѵ���B.�� ����y�  ʞr�t   ����F�X   �K   �^ʚ|�[   ����v   F[�A   ������  ʞz�� ���0z!�HJ��R  ٺE
�C   ��ʚb�K   &�X   �iپK�   �
���� ����� ������M��о�U�щ��ٷ�i����������K����Y���J   �� �H   ���P/��K��	�A   Uʙq��ٽK��F[r��=���
�� ������M��о����/�� �����[ ʞr�[   qk��@   M��x   �O   qU�D   U�����/������� ���,�j�3Y��]  ٺE�J   �� �H   ���P/��K���� ����+Eٷ�i���q�­��ф��|����ٟJ���v   F[��U-��%ʙ|��qHV%�[   qk��@   M��x   �O   qU�D   U�����/�������Ƒ��/#]9�Y�pN  ʞr��
�����յ��
�� ���/�/�  ��V�A   U�R   ������  ٺM�v   F[�A   ������  ʞz�� ����rʓ�z��筯b���ѧ ���M���ʝ���X��ѵʻ}���A   U�R   ������  ٺM�   F
O��d   z��O   �k   Fq�W   q̷���&������� ����rʓ�z��筯b���ѧ ���M���ʝ���X��ѵʻ}��-�R   qHٽF	����X��UE.�P   ��پU�o   �|   �z��X�H   �.��&��榥�    �v   F[�A   ������  ʞz�R   qH�v   ������  ��^!���������������ے=[  	(
�C   ��ʚb�K   &�X   �iپK�   �
��/�Y   �� '�[   �ʛt��|�[�����.#Q��Y�OL  ʞr�v   F[��U-��%ʙ|��qHV%�}   �� �   �ٿC��o�l�'�W6jXn�ׂ����   M��ô�����/���}   �� �   �ٿC��o�l�'�'v�ς���ʓ�z��筯b���ѿ ��X��Ѷʻ}��.�P   ��پU�o   �|   �z��X�H   �.��&�炷��ʓ�z��筯ʛ�����}   �� �   �ٿC��o�l�'�}   �� �   �ٿC��o�l�'���F��D������
0��٤��U��_����ʣQ=<��^|Y�뵤��ٷ�i���q�­��фʓ�z���ٹ�ѵ��|����ٟJ���}   �� �   �ٿC��o�l�'�R   qH�v   ������  ��^ �]�  ʞz���  ʞz�[   qk��@   M��x   �O   qU�D   U�����/�������΀��    �[   qk��@   M��x   �O   qU�D   U�����/�������΀����΀����[��΀��C�Y  $yz���   �+E�(�  
��  
�̦���.��淥��+Y��  ٺQ�J   �� �H   ���P/��K���;Y
�\n�HJ�����v   F[�A   ������  ʞz�t   ����F�X   �K   �^ʚ|�[   ����] 
0 !�   K0 #    	�3Y�\v�HJ��ր��.�P   ��پU�o   �|   �z��X�H   �.��&��򷥁�.s��򷥁�kA�Y�   %¿#���ْE	(0 �'�  ��^.��  ��^-�R   qHٽF	����X��UE�{�  �;��;��sq�Y�Ky�Y�;Eq;A�;��;�����  ���A   U�R   ������  ٺM�� N�;�     ��  ʞzJvJ��.�P   ��پU�o   �|   �z��X�H   �.��&�t   ����F�X   �K   �^ʚ|�[   ��� ћ�����������ْE	(�;�    �R.�OJ�[nʢ�F��   # �   0z#  2   ��v�ke�Y�;����q��   ��    �t   ����F�X   �K   �^ʚ|�[   ����+���.�OF�[n���}   �� �   �ٿC��o�l�'�t   ����F�X   �K   �^ʚ|�[   ����3��\R�HJ�Lٶ��^���A/�Y   �� '�[   �ʛt��|�[�!������������������ђ	(
�C   ��ʚb�K   &�X   �iپK�   �
����    �S����[����EV^�+AY+�i��X��#�J}��H���v   F[��U-��%ʙ|��qHV%�}   �� �   �ٿC��o�l�'�nJ��X %¿#����R[  �9�  -�̢��� �e   M��ð�����/���}   �� �   �ٿC��o�l�'�߆���0r!��HJ�@���ٺE�v   F[�A   ������  ʞz�R   qH�v   ������  ��^��B���/#W��Y�����ʞr�[   qk��@   M��x   �O   qU�D   U�����/�����/�Y   �� '�[   �ʛt��|�[���b���,#Q��Y����ʞr�t   ����F�X   �K   �^ʚ|�[   ��������
B2��[n�p�����V��"���/#W��Y�j���ʞr��淥�0t!V�HJ�����ٺE�   F
O��d   z��O   �k   Fq�W   q̷���&�������Ʒ��0u!B�HJ�𧁶ٺE�v   F[�A   ������  ʞz�צ���0v!~�HJ�ŧ��ٺE�   F
O��d   z��O   �k   Fq�W   q̷���&������R   qH�v   ������  ��^�̺���v   �v   F[��U-��%ʙ|��qHV%�[   qk��@   M��x   �O   qU�D   U�����/�����.�P   ��پU�o   �|   �z��X�H   �.��&�R   qH�v   ������  ��^��,! n  �̾���.��)H ��/b�ת����/�  )�Y�󝷁����  �v   F[�A   ������  ʞz�t   ����F�X   �K   �^ʚ|�[   ����+���K�롧���v   F[�A   ������  ʞz�R   qH�v   ������  ��^�A   U�R   ������  ٺM�   F
O��d   z��O   �k   Fq�W   q̷���&������ߊ���    �   F
O��d   z��O   �k   Fq�W   q̷���&������}   �� �   �ٿC��o�l�'�ߒ���    �q�ߒ���ʚ�ߒ����ג���rז���Fٛ   �ϒ�����뭷��
 2nM  �OB�[n�ߎ����玴�� U��   2zH  �׆���0 �ώ����J[ ̚
5������    �F������پH�������󭧁�a󩷁�)-�Ϛ�����{��k����
�Ģ���/�H;H ��R��A�	�������ý��� 
K�c�}   �� �   �ٿC��o�l�'���ܪ���,�Ov�[n�犴�� .|�_����������� ћ����sM}|Y�͒AP��WznXn�]   �������!
] J�]�  �����0�!��HJ�    .-�[    ْA�:mY(«�=~v��6O  z���x  ��
x  ��x  H�:mB�ao  �2mV���W    ʞj���������ْ	(�;A�6A�3��+��+�	�A   Uʙq��ٽK��F[r�v   F[�A   ������  ʞz�'� /{��z  �A   U�R   ������  ٺM�   F
O��d   z��O   �k   Fq�W   q̷���&�������ʚ�e�  ʞz��������ʛz��4�����K����Y���;A�M @�;�"�HJ�@�3A�/M�+����+�ٷ�i���q�­��ф��|����ٟJ��������    �v   F[�A   ������  ʞz�v   F[��U-��%ʙ|��qHV%��ʰ���S����[���4� F��   ��J�F�oʠ^=p��}�q�R��W
U�+�Y+�U�KنC.p��J�F�oʠw<d��}��  /�Y   �� '�[   �ʛt��|�[�-�R   qHٽF	����X��UE�P�b�R   qH�v   ������  ��^�����   ̓
�+�U�Kنi._��F�oʠs=L��q�R��P
B�+�U�Kن@/]��ʛ���v   F[��U-��%ʙ|��qHV%�X�K���'�ʓ�z��筯ʛ����������� A�+��+��y��H   �;��;���X	@�;�[   �@�3�ٗK�3��+�a+�){�L:H �R�1^ Fބ   �v�zz�����U��   �3A�/Mi���t�   q͋   �4� F��   �v�zʰ�����R��[���Ci�̚
@�3A�M K��v�zz�����.m�v�zz������   o�+A�<EپK�;��3A�/MٔH�+��;�
��  ٺM�g�v�zʰ�����R��[���C�;A�>M    �R�R    �v�r    �;� ��   �;�
�R�A`  �;�[��   �� g�   ̓
E0�v�K  �Z�+A�M 
C0 �v��F  �� ��H   ߾=v�R�0Va>Q�R�VE�Q0�v�NK  ��/�v��G  �i�   ̈^�;A�6Ea3�)r���3A�p  ��H�;��   ̚
�3A�/M�+��3�����ѿ��|����ٟJ�ڏ� �3A�+��/A�;A�6MY3��3��+��;��|�[   qk��@   M��x   �O   qU�D   U�����/�����.�P   ��پU�o   �|   �z��X�H   �.��&%¿#�����������+¶���   --�R   qHٽF	����X��UE�A   U�R   ������  ٺM�CY\|Y q�|  �^|Y0}!�HJ�>���ٺE2rLXn#Y�Y����ʞr!z{KJK2.�[n������V�A   U�R   ������  ٺM2JLXn#X�Y�Z���ʞr�R   qH�v   ������  ��^/�Y   �� '�[   �ʛt��|�[�_|Y0|!�HJ�����ٺE2"LXn#Y�Y�����ʞr�[   qk��@   M��x   �O   qU�D   U�����/������A   U�R   ������  ٺM2LXn#Y�Y����ʞr!�{KJK2�[n������V-�R   qHٽF	����X��UE�_|Y0}!�HJ�y���ٺE�J   �� �H   ���P/��K���v   F[�A   ������  ʞz!�{KJJ2�[n�������V�_|Y0}!6�HJ�����ٺE2�LXn#Y9�Y�����ʞr�[   qk��@   M��x   �O   qU�D   U�����/������_|Y0}!>�HJ�6���ٺE�J   �� �H   ���P/��K��2�LXn#Y=�Y�.���ʞr�_nOXn    �v   F[�A   ������  ʞz�]KJ���F   i��'������4R���M��о�������    �R   qH�v   ������  ��^�A   U�R   ������  ٺM�;�    �H   U.x��S   i��\   �\   U'F�s   Fߓ���������J   �� �H   ���P/��K���;�    �@�3�ٿH�3��+�a+�U�[  ��q�`  �R}�q�R��g:�;�[   -�R   qHٽF	����X��UE�A[  �J   �� �H   ���P/��K���   F
O��d   z��O   �k   Fq�W   q̷���&�������   �R}�q�X��z
G�3AY3�U�Xل@/`�e����A   U�R   ������  ٺM��vJ����J�W��[   qk��@   M��x   �O   qU�D   U�����/�����-�R   qHٽF	����X��UE����[��/�Y   �� '�[   �ʛt��|�[����3��:D� �v   F[��U-��%ʙ|��qHV%�r�X    �'� U��Y  �;��3A�*H[��.����V��^��"�����.������M��о������&����������'� ,u��������P��*���   ��������'�K-r�����H   �r��ʲ|����������r����:_�f ��1����M q�m  ��"����^M��/�߬F�_H  ������zz������   q�]  ��&��� Fߡ   ������zʳ�����������XRH��!����z���.r������"z /|�-��"����^M��<�߾=O��"����^M��<�g�   <v��"����V��X����"����^��[����,�#�  ��^�m��1����6MٗH��-�����-����|e[��>����H��1����<M    ��"����	R    ������r    �;� ��   ��5�����"����Ch  �;�[��   ��5��� �   ̚
F0������S  �s��1����M 
g�;�    �� ��������v������zJ��������R�� �-�H   ߬=d��"����1Va>K��"����VE�&���h0�������R  ��&���.������O  �e�   ̓j��1����<Ea�5���)l�������1����Sx  ��H�+�ۜ�   ߬=��"����^����&�����.����4�����K����Y��;� ��"�����&����R��"����^}�&����������X
�C   ��ʚb�K   &�X   �iپK�   �
��-�R   qHٽF	����X��UE��    �S����[���4�pF��   ���+�1�]ۼ�^|Y��l ٺA߾<4���N�V��R{KJ�X
�C   ��ʚb�K   &�X   �iپK�   �
��/�Y   �� '�[   �ʛt��|�[��i�J   �� �H   ���P/��K���#���F�;�نn/w�r�[   �r�`<R�V�q 
�3EٿM�����ٺM
�C   ��ʚb�K   &�X   �iپK�   �
��/�Y   �� '�[   �ʛt��|�[�!��������+¶�2��[n-�    >�l    ��F-���S+  �;�    -�R   qHٽF	����X��UE�H   U.x��S   i��\   �\   U'F�s   Fߓ���������Aٷ�i���ٿ��3��   F
O��d   z��O   �k   Fq�W   q̷���&��������L;  ʞz���}   �� �   �ٿC��o�l�'�R   qH�v   ������  ��^����[GJW�;�    ����������  ����   �+E��.�v�3���8  ���[   qk��@   M��x   �O   qU�D   U�����/������V}��K ��   �������3��"8  ���A/�Y   �� '�[   �ʛt��|�[����W    %¿#������������ђ	(0Q�v� �  ʞv���}   �� �   �ٿC��o�l�'�R   qH�v   ������  ��^�4� F��   �'�ʝʓ�z��筯ʛ�ʣ^F��   ��ʛ£�V���M��о�U�щ����K����Y��v   F[�A   ������  ʞz�=.�P   ��پU�o   �|   �z��X�H   �.��&�t   ����F�X   �K   �^ʚ|�[   ����3E� �v   F[�A   ������  ʞz%¿#���ђ#�-�Y>�    
�    �2�  �7�  	(��'��0 �צ4����]  �A   U�R   ������  ٺM�v   F[�A   ������  ʞz�߲6��    ���%��    .�P   ��پU�o   �|   �z��X�H   �.��&�R   qH�v   ������  ��^�̶��    �R   qH�v   ������  ��^-�R   qHٽF	����X��UE�̞��    �ߎ6��    �v   F[�A   ������  ʞz�R   qH�v   ������  ��^�̊��    �v   F[��U-��%ʙ|��qHV%�v   F[��U-��%ʙ|��qHV%�ߞ6��    ���%��    -�R   qHٽF	����X��UE�y|Y���%���V  z��������<��v   F[�A   ������  ʞz�[   qk��@   M��x   �O   qU�D   U�����/������4R���M��о�����Ď���̂��    �}   �� �   �ٿC��o�l�'�ߢ6��    �q�ע6��ʛ�ע6���Ϣ6��rϪ6��4+�R}̆��q�R��WK���vJϢ6���ߦ6���P��_�6���R   qH�v   ������  ��^/�Y   �� '�[   �ʛt��|�[��܂����[�܂���;������%����L��� �R   qH�v   ������  ��^�^|Y��%�����  ٺA���%��	�A   Uʙq��ٽK��F[r	�A   Uʙq��ٽK��F[r�Á%�� q͢o  ���������������������H0 ���6���%Z  ��    �R   qH�v   ������  ��^�����,�߶6���`���ʞv�v   F[��U-��%ʙ|��qHV%�}   �� �   �ٿC��o�l�'���6�� /r�ߪ4��1�Y�r���6���ת4���Ϫ4�����6���R   qH�v   ������  ��^�A   U�R   ������  ٺM���%�����'����'��ٗK��'���Ù'��Wq��n  �܊���mω� n���6����  ʞz�צ4���z�[   qk��@   M��x   �O   qU�D   U�����/������xJ  
�C   ��ʚb�K   &�X   �iپK�   �
�� ^  ��'��ټA�����.�v�����V.�P   ��پU�o   �|   �z��X�H   �.��&�t   ����F�X   �K   �^ʚ|�[   �����'��ۿA^  �܂����R,�ه����R��U  ���%��
���  ٺM��'����y\  	�A   Uʙq��ٽK��F[r�6F  ���6���6�  ʞz"�B�צ4����BO  �}   �� �   �ٿC��o�l�'�v   F[��U-��%ʙ|��qHV%��p  .�P   ��پU�o   �|   �z��X�H   �.��&�[   qk��@   M��x   �O   qU�D   U�����/����������,���  ��^�f�Ă����x  �A   U�R   ������  ٺM	�A   Uʙq��ٽK��F[r�2G  ���6�����  ʞz�צ4����RO  �R   qH�v   ������  ��^�\T  �v   F[�A   ������  ʞz�}   �� �   �ٿC��o�l�'���6�����  ʞz"�B�צ4����:O  �R   qH�v   ������  ��^��W  �v   F[�A   ������  ʞz�ϲ6��ʘ�ϲ6���t   ����F�X   �K   �^ʚ|�[   ����v   F[�A   ������  ʞz�ߦ4��Lx  �����������0^ <V�̖��    �x�����������RU^����\  ���߲4���ϲ4��rϲ6��:j�Ă����O  
�C   ��ʚb�K   &�X   �iپK�   �
���̂��{\  ���%����%��ٗH���%�����%���M E���'��    �i���%�����%���>Aq?M��\  ���߶4���϶4��r��6��>Q�������E  ���%���6M���%��2 M  ���6�� �6O  ���6��J�.���6���-���ʞr�ϲ6��ʰ���6���ߦ4��Lx  �����������0^ <V�̞��    �x�����������RU^����\  ���ߺ4���Ϻ4��r��6��>Q������DE  ���%���6M���%����'��ۼ\  ��5%�����%��ٖH��1%����5%���M E���'��    �k��5%����5%���4Aq6Mѿ��6O  ���̚���ܚ��E�"��	B��5%����W  ��6���z���6�����6�� �6O  ���6����n ^  ��"���x  �����}�
�����ٺA��C  �v   F[��U-��%ʙ|��qHV%�ז6��ʛ�ז6���Ϧ4��Ș6O  ��
6����
6���"z /r���4��    �^��
6����
6���vbz��6O  ������������Eܲ��B��'����[  �ߦ4��Lx  ��f���Ĳ����[��b����f���3^ <V�����    �z��f����f���	RU^��x  �����'�����'��a�q%��-@��:6��2&OXn��66����e  ����66����%����G  !J�HJ����,���  ��f���^���������,���  ��^��b���x  ������PZM  �[   qk��@   M��x   �O   qU�D   U�����/������rS  
�C   ��ʚb�K   &�X   �iپK�   �
���̶����[�̶��/�Y   �� '�[   �ʛt��|�[��Ă����x  ��n����n���3^ <V�����    �z��n����n���	RU^��x  �����'�����'��a�%��)]�צ4���no  -�R   qHٽF	����X��UE�̂��{\  ���$����%��ٗH��$����$���M E���'��    �i���$����$���>Aq?M��\  �����4�����4��rφ7��>d��^��.!xKJ��R����C  �;�X��R��/��f6����r  Y�Y��Q%�����  ���$���6M�� %�����%���z�  ٺM��$��3�\  �� %����Cvx  �A   U�R   ������  ٺM�N  �}   �� �   �ٿC��o�l�'�t   ����F�X   �K   �^ʚ|�[   ������%��پH���%����'��ۿ\  ��$����$���M E���'��    �i���$����$���>Aq?M��\  �����4�����4��rϺ6��:Q�Ă���:U  ���'��_6O  ���7���׺6��ʳ���7�����7��� z /r���4��    �^���7�����7���vbz��6O  ������������E��~��	w���$��
\|Y��$���XQ  ��J��$���Ă~���	Q  2n�[n�Ϧ7���g�  ���7���z�׾7�����6�����  ʞz"�B���7�� �6O  �Ͼ7����ty\  �v   F[�A   ������  ʞz�}   �� �   �ٿC��o�l�'��{  �̪����[�̪���A   U�R   ������  ٺM��'��ۿ\  ���$�����$���M E���'��    �i���$�����$���>Aq?M��\  �����4�����4��rώ6��:Q�Ă����W  ���'��_6O  ��7���׎6��ʳ��7����7��� z /r���4��    �^��7����7���vbz��6O  ������������E�"~��	w���$��
\|Y���$����_  ��M���$�����~����S  2n�[n���7����  ��7���z���7�����6�����  ʞz"�B��7�� �6O  ���7����t}\  
�C   ��ʚb�K   &�X   �iپK�   �
���k^  �J   �� �H   ���P/��K���v   F[�A   ������  ʞz�߮6��ʚ�߮6���}   �� �   �ٿC��o�l�'�[   qk��@   M��x   �O   qU�D   U�����/������Ă����x  ��.~����.~���3^ <V�����    �z��.~����.~���	RU^��x  �����'�����'��a�%��)/�צ4����u  �H   U.x��S   i��\   �\   U'F�s   Fߓ���������v   F[�A   ������  ʞz�ߦ4��Lx  ��f~���Ċ����[��b~����f~���3^ <V�����    �z��f~����f~���	RU^��x  �����'�����'��a�q$��-@��:7��2&OXn��67���j  ��{��67����$���N  !J�HJ��~��,�e�  ��f~���^��~�������,���  ��^��b~���x  ��~����PVO  �R   qH�v   ������  ��^��[  ���%��پH���%���J   �� �H   ���P/��K����'��ۿ\  ��}$����}$���M E���'��    �i��}$����}$���>Aq?M��\  �����4�����4��rϞ6��:j�Ă���\P  
�C   ��ʚb�K   &�X   �iپK�   �
���̂��{\  ���'����%��ٗH��'����'���M E���'��    �i���'����'���>Aq?M��\  �����4�����4��rφ4��>d��^~��.!xKJ��R~����H  �;�\��R~��/��f7����{  Y�Y��Q$�����  ���'���6M�� $�����%���N�  ٺM1�u��'��3�\  �� $����Cbx  /�Y   �� '�[   �ʛt��|�[���   F
O��d   z��O   �k   Fq�W   q̷���&������}   �� �   �ٿC��o�l�'!�zKJ �u�  ʞv�߶6���[   qk��@   M��x   �O   qU�D   U�����/�����������#[�������H  ������ߦ4����2O  ���6���[   qk��@   M��x   �O   qU�D   U�����/������[���%��ۼ\  ���%�����'����\  ��'�����%��a�'��U�
[  ���%��ٷ�i���ٿ�߷=z������� z  ���M��о������U�A[  ���'��_6O  �ߞ4���מ4���v�ώ4�����6���ߖ4�����6��ț6O  �ג4���y�ܲ����x  �ܲ���̶��{\  ���'����'��a�'��.k��4����  ���������Ϟ4���vdx  �̾���[��'��ۿ\  ��'����'�����'��a<A.|���ĺ���R��x  �̺���R�A   U�R   ������  ٺM	�A   Uʙq��ٽK��F[r������צ4���#z ,��4��ʝvʓ�z��筯ʛ�̓(�Ñ'��۹A^  ٷ�i���ٿ�߷?�܂���KV�צ4���[-�R   qHٽF	����X��UE/�Y   �� '�[   �ʛt��|�[��܂����x  �܆���̆���1^ <V�����    �z�Ć���܆���RU^��x  �����'�����'�� d��'���|EX�Ă���H�J   �� �H   ���P/��K���3�>�D    !���M 6� n�� Y'� JY� n� Y#� J�� nz� YS� J�� n�� YH� J�� n�� Y��2�[n-�    >�l    /(�.Zi���5~j�9�  �V��V�&VM��*mF� �^�R�V�R�D&�HJ��a�:X��a�</E�я?_�nD ѳ��j  �RU�a�:X��߈?j�^U�Y��jz-���  �R��VU�ѳ# -�;l  ��.vѳ�ol  ����]  �]�[n!%�ZM>�D    ��J�M E�,:r�	�8Ma�<_�1�Y���g0��T  �8M߾<_�1�Y�;M�0A�3A�(E�+E�6�������H	����X  ͚
��M߈<_�1�Y�Mѵ��X��Ѷ�ZYٟJ���z�v�MC �ZE� ـY%-�s    ٺY�z ����?Y߾<_�1�Y������F/�ZM�����Z 2Ψ[n���  ����0�!»HJ�    .-�[    ْA	+�~n£.�&ZQ�:mN6jXn�&�  �=~V�rz��G�-M�u�	v�	r�v�W�[n²E��*mzKїr�<a�«L�~U[ �bI  �=Aq�r�Kю̬y�-Mq�J�.�^P���  �AٺEq� ��J  ޾=R+��J  ѵ��l  �N��HJ���2mB!%-�s    ٺ]�z a�?E�/>�zr�L��[n�"��)P#[���{D  �z̚L��[n�z�v�v�r�	r��������0ѵ�ln  ��.��,z̬L��[n�!z����X��Ѷʻ}������F  �Z]� �Y�!���������������я�\�[n�n̚
T�6��>�޾=PB�.x���H�w���  ʞz�J    �j    �8Q    �7�  ��������F/�ZM�M   �Z 2n�[n�p�  ������������ZA[
@���  ٺMѸ�z ��#��Y>�    
�    	+�
mz)£(�&Z]���  �rʜr�rz��~b�Y�^�R�V�R�D&�HJ��a�:X��a�</E�я?_��@ ѵ�oo  �
RU�a�:X��߈?j�^U�Y��jg+�^�  �"R��VU�ѵ# +��p  ��.vѵ��p  ����Y  �]ޓ[n�~j#>�D    ��J�M E�,:r�	�8Ma�<_�1�Y���g0�FQ  �8M߾<_�1�Y�=M�0A�5A�(E�-E�6�������H���>G  ͚
��M߈<_�1�Y�Mѳ+��|����ٟJ����W  �:mJ� ��HJ�������������8A߾=G���	���.tu�
O���[�@�Y�  ٺM�8A    �V    �n    ���+¶���x  -��6�����⇶� ��  M���𣁶��/�Ԏ�L   �v   F[�A   ������  ʞz�[   qk��@   M��x   �O   qU�D   U�����/�������    �R   qH�v   ������  ��^��    �[   qk��@   M��x   �O   qU�D   U�����/������A   U�R   ������  ٺM��%���_6O  �����������v��ʰ��������z��Ұ����ʰ��b�Ұ����6O  ����ꇶ���*�����*����VUR����\  ��ʢFټK  ������ z /r�����    �^�����������vbz��6O  ����2�����2���?��*����3^ <V��>���    �z��*�����*����	RU^��x  ����-�����-�����)����t�����H   ��9����M E�����    �i��9�����9����?Aq<M��\  ����"�����"���J������ް����ް����Ⱕ���Ⱕ� 't��Ⱕ�    ��գ��3�\  ���  ٺM����������ݣ����9����6M��ѣ���]��갥�Ș6O  ��갥���氥�Lx  ��������E��
Q��ѣ����·��.��p  ��R����ݣ����ᣁ���񣁶H��ᣁ�
��*����TT  �    �6O  ��ְ��J�,������v��������*�����W  ��9����6A��*����^.������4y  ��*�����*����VU^��x  ����ţ����9����<M��٣����٣���>�  ٺM��飁�3�\  ����Y�������r������ z /r��&���    �^�����������vbz��6O  �������������x  ������}��    �6O  J���*����R��*����������^�jX  ��9����<Aq�������\  ��ʢFٟ   �[   �x  ���}�
��*����R,��ʰ����9����E  ��ư����9����<Aq�������\  ���[   U���*����R/������(r  ��*����R��އ�������҇���[������ۼ\  ������������a�ͣ��.k��  ��⇶���҇���챵�[   �x  ��*����R}���9����?A�\H  z���[q�M  ��*����R/������v�    �6O  ������vb�.������!u  ��*����R��&����H   3�\  ��9����/Aq���������ʰ��r�����=c��ڇ����x  ��ڇ����ڇ����&�����x  ��&�����[  ��5����ۢ������"����[��1���ۿ\  ��1����    �6O  ��ʰ��J�G�"���
\��H  ��ư������������    �6O  ������vJ���*����R��*����^��.���!���������ْy	(�3��A q��   �4���sz  ���M��о������.q��Lsz  .�O>�[n�[   qk��@   M��x   �O   qU�D   U�����/���������x  ���B�;�_6O  ������.O  ����r�=q�4���rz  ���M��о������.n��țVM  �k	�Y�����X    �[   qk��@   M��x   �O   qU�D   U�����/�������[  i��'�ʝz��/�Y   �� '�[   �ʛt��|�[�����jx  {   �}   �� �   �ٿC��o�l�'����BO      �v   F[�A   ������  ʞz�R   qH�v   ������  ��^����x      ����&O      �   F
O��d   z��O   �k   Fq�W   q̷���&������R   qH�v   ������  ��^����x      ����O      �;�_6O  �����v�����z�����v�����������M��{\  �;��3�ۿ\  �3��+�a+�.q�/���  �4��챬�������v�������V����x  ����E�
K�������v�[   qk��@   M��x   �O   qU�D   U�����/�����!���M �������������~v���v�5~j� z����M��M�A�E�о�7���L��G[ �zr�
l�?�޾=DB�.dr����?�ѳ��   ! �A E�/l#[����   ѻ%�R �rʢa>^E�)o#[����   ѳ�w{  �=~j�'z����K����Y���;M�#A �^f ѻ�A ���(«�^��.c����͚
Cf�=\����S/��  ��^�^    �v    �8E     ������8M
�~v��  ��^M��8M�8A�8E'����������������ZM��я=~�^��.c����͚
Cf�=\����S/�2  ��^�^    �v    �8E     �^ �������ʼA �������������#���Y>�    
�    ʶJ�ZJ	+�:mN�\|Yٷ�i�z�H�о�7�ZUї�ZQ�~Z�Za��K  ͚
o�mB��ѯ�&OXn��|����ٟJ���ZU�mz �FV�ZY�"m/�Za�:mN6jXn���  �~j�2mn�~2H�*mn�������[n�Z]
-�2mf�k   �*m~Y�Y�~.�Ze��HJ��   #����-�=~j�mN��c	A){��sH �R�~bU�a�:X��a�F��   �v�g�[nJ�E�){�=sH ���jM  �vb�E�)|¢��,H�zb�}�
�]c,���  �/vʞrb���0 ��H  ͚
C�;M�A�zO �=~f����J  �vr�Kц̥q�  �^U�
�]c,���  �/vʞrb���0 �-H  ͚q�x  (�j[  ��#�r i�r�8a�<7�^E�/{�"�HJ�1��:�^E�.a����͚
Cf�=\����Q/�k  ��^M��+M�+A�+E�9Ma�<_�1�Y�;M�1A�3A�)E�+E�6����6�ѻ%�V ��[  a�:_��P �3M߷=����.`u�
Sߥ<��	�����N���ѻ%�V ́[0�S�����#�r �;EنV-zr�X0�����	����H  �z̚L��[n�'z}�ѿ��|����ٟJ���z�v�^u ��#�r �:m^�R�I^�M[ �^ ���������������)�&ZYف�я?_�dP �8Mi�r�
c�6�`�=y���
Wa�Fߤ   ��!���z�v�rh��v �2mNE�/(s�
a�=v���	�D�.gu�
\����z�v�rh��v ��!  ٺM� M� A� E {�%�R r�
L� A�fL��A D�.#�rʣa>^E�) r�
}�6��>�`�={B�.c��)�[��� M� A� E�+   �H�A /�  ��^)�^�R�V�z    �[%�R p$r:R)�W    �[%�R ������񧁶��������������0�!��HJ�    .-�[    ْE�;A	(ª��E)����,����<�L�;�ю�|��    ߾4XM�
��   ٺM�;A�Y�v��ʚ|̚Ki���3  �vʞz�� J����/��v̚ka�?X���MѶ�v��X�1[��Ѵʻ}���<��
^�2R��.c����͚
Cf�=\����S/�m  ��^�R�
R    	a��z�� �E-|­�^�:R!�^O �3��W    ћ�z ����������i��^E�U��   �?�޾F��   u�q��   ��я��¤���M��+M�+A�+E�о�7���N��N[ z��^E�._��͚
Sf�=LE�/G��,������� �r�G0����� ��rʢa>^E�)o#[�������ѳ�����4^��ѿ��|����ٟJ���z�v�^u  ���������*m^-�ZEa�=p�~n��.u��  ��ц����x  {\  a�<�!�E �~n�r ��~v̚n	�~nѮ�ZE��.u��  ��ц��{\  � �r ���������������mR��.s�
mJ��[  �����������+¶��-����.�¡�  /�Y   �� '�[   �ʛt��|�[��A   U�R   ������  ٺM�3���M[      �A   U�R   ������  ٺM�v   z��4���R  ���M��;�_WH  �J�^�R�V/�Y   �� '�[   �ʛt��|�[�/�Y   �� '�[   �ʛt��|�[��O   i��'�ȝHH  ��ԡR   qH�v   ������  ��^���
      ��0l!֭HJ�4⁶ٺE�v   F[�A   ������  ʞz��0 # �\ �HJ�A   U�R   ������  ٺM�v   F[�A   ������  ʞz��0 ![ V �\^�HJ����  /�Y   �� '�[   �ʛt��|�[�-�R   qHٽF	����X��UE��!���ђȶrH  )�׊���!^  �R.�O:�[n�'vʓ�z��筯ʛ��׆����vJ׆���F�/�ل.$�vJ߆���F�6�هf.6�vJφ����X"�[   qk��@   M��x   �O   qU�D   U�����/������R}̢����	[ �߂��� �>   z���������<���J   �� �H   ���P/��K���󵤁�B2��[n��ȶ���V�A   U�R   ������  ٺM�õ����+Aٷ�i���q�­��фʓ�z���ٹ�ѵ��|����ٟJ��%¿#�^ ����^  ����������ђ	(�3��;�_vH  �A/�Y   �� '�[   �ʛt��|�[�!���������������-���p �C�t   ����F�X   �K   �^ʚ|�[   ���	�A   Uʙq��ٽK��F[r ћ��������������`[  ����������+¶/)����Ll  �z�J   �� �H   ���P/��K��	�A   Uʙq��ٽK��F[r ћ�����-���4R���M��о������B10f�v�3�ۿ[  ��(  ٺE�+���[   .�P   ��پU�o   �|   �z��X�H   �.��&�[   qk��@   M��x   �O   qU�D   U�����/������c�A�;�_HH  ���M��о�U�щ����K����Y�� ћ�z �������+¶/)���'�ȝHH  ʓ�z��筯ʛ���A����z�J   �� �H   ���P/��K��	�A   Uʙq��ٽK��F[r ћ��������������ђ	(�3��;���[  �L�}   �� �   �ٿC��o�l�'�R   qH�v   ������  ��^!�����+¶��r-���y|Y�+Aٷ�i���q�­��ф��|����ٟJ�ڡR   qH�v   ������  ��^�H   U.x��S   i��\   �\   U'F�s   Fߓ���������;�    .�P   ��پU�o   �|   �z��X�H   �.��&���kыY�;��� }�+���.�O�[n̚
i�xH  �}   �� �   �ٿC��o�l�'�_��   ��ٷ�i���ٿ��3��;�    ��    �S����[����E�q��   ��}�M��vʣS<X���v   F[�A   ������  ʞz�}   �� �   �ٿC��o�l�'�vJ���J��R�C�v   F[�A   ������  ʞz��ʘ���v   F[��U-��%ʙ|��qHV%�����R�J   �� �H   ���P/��K�� ћ�z ����+¶��-�4R���M��о������H   U.x��S   i��\   �\   U'F�s   Fߓ����������VL�rH  �v   F[��U-��%ʙ|��qHV%�[   qk��@   M��x   �O   qU�D   U�����/�������v   ��B   �;�\   ��t   ��H   �;�^   ��w   ��K   �;�    ��}   ��L   �;�]   �A   U�R   ������  ٺM�;�    �@�;�پH�;���V_�3��*Ğ���R�]K�_����R���A�+��.M�3��6A	�A   Uʙq��ٽK��F[r ћ�����������ےQ^  	(�󡡁��6jXn�vʓ�z��筯b���ѿ ��X��Ѷʻ}��.�P   ��پU�o   �|   �z��X�H   �.��&�R   qH�v   ������  ��^�A   U�R   ������  ٺM�v   F[�A   ������  ʞz�t   ����F�X   �K   �^ʚ|�[   ���
�C   ��ʚb�K   &�X   �iپK�   �
���A   U�R   ������  ٺM�J   �� �H   ���P/��K���v   F[�A   ������  ʞz�}   �� �   �ٿC��o�l�'�J   M��ñ������v   F[��U-��%ʙ|��qHV%�e   M���q�����/�ԏ߆���~�   F
O��d   z��O   �k   Fq�W   q̷���&������[   qk��@   M��x   �O   qU�D   U�����/�������b����Ħ���/�Y   �� '�[   �ʛt��|�[�.�P   ��پU�o   �|   �z��X�H   �.��&/�� ���� �R   qH�v   ������  ��^�ܢ���,�%wH �̪���.�P   ��پU�o   �|   �z��X�H   �.��&�ߎ���l�   ��.@�ߎ���l�   �^  �v   F[�A   ������  ʞz�R   qH�v   ������  ��^�̶���    �U�Ķ�����[�Ķ�����b������   Gܶ���8������h�̶�����_G�����V����v   F[��U-��%ʙ|��qHV%�φ�����A[ �ߎ����R   qH�v   ������  ��^�̪���[�   ߾<X�L�����׎���Ȼ�   ̓
�������   �Z}  /�Y   �� '�[   �ʛt��|�[�/�Y   �� '�[   �ʛt��|�[��Y   i��熲����/�Y   �� '�[   �ʛt��|�[��H   U.x��S   i��\   �\   U'F�s   Fߓ��������������i�A   U�R   ������  ٺM�J   �� �H   ���P/��K����p�����a����
OXn��|���ʓ�z��筯b���ѿ ��X��Ѷʻ}����ƃ���Ħ���/�Y   �� '�[   �ʛt��|�[�-�R   qHٽF	����X��UE�� ���X�ܢ���,��xH �̪����A   U�R   ������  ٺM�������   ̚
b�������   ��  /�Y   �� '�[   �ʛt��|�[���b��� �B   M���p�����/����0z!��HJ�z�ٺE�   F
O��d   z��O   �k   Fq�W   q̷���&������ߊ���    �q�ϊ���ʘ�ϊ����犲��O'J�'���F���ʓ�z��筯b���ѧ ���M���ʝ���X��ѵʻ}������见��   ��駁�۟�   ��Ń�����   ,��ഥ�l�   .��㴥�Ȼ�   ��է��ۜ�   ��b���.�v��,  ʞ^�v   F[��U-��%ʙ|��qHV%�[   qk��@   M��x   �O   qU�D   U�����/������R,�������^�A   U�R   ������  ٺMi��i-�R   qHٽF	����X��UE/�Y   �� '�[   �ʛt��|�[�!���M +¶��R-��ݏ���;�ȖA   U�R   ������  ٺM	�A   Uʙq��ٽK��F[r�;�    �@�;�پH�;��3�a3E'�vJ�z��K߾=9�R}�M��o����Y   ��i��k�a�=}�R}�M��o����Y   ��i��k�i��vJ��P/�Y   �� '�[   �ʛt��|�[��0��� ћ��������-���   �8�[   qk��@   M��x   �O   qU�D   U�����/������A   U�R   ������  ٺM ћ�����ْU	(�3���۹A[  ٷ�i���ٿ�هi.o��LR  .���c����4���s  ���M��о������V
[�3�ۿ`[  �������v   F[�A   ������  ʞz# �%=  ٺM�+�c�[  %r����.H   /m# �=  ٺM�3���[  
�C   ��ʚb�K   &�X   �iپK�   �
���A   U�R   ������  ٺM�3��з�������/  ʞz�������R   qH�v   ������  ��^�A   U�R   ������  ٺM�3��3�
�C   ��ʚb�K   &�X   �iپK�   �
��������^  �C�J   �� �H   ���P/��K���+�ټM�+��J   �� �H   ���P/��K����۸A[  �v   �'������ʚ_���}   �� �   �ٿC��o�l�'�R   qH�v   ������  ��^����s  ���H�|�z�z�v�v�r�r�[   qk��@   M��x   �O   qU�D   U�����/������A   U�R   ������  ٺM�+�ټD�+���۸[  �x   �'�����t   ����F�X   �K   �^ʚ|�[   ����;�پP�;�
�C   ��ʚb�K   &�X   �iپK�   �
��������
  �H�J   �� �H   ���P/��K��
�C   ��ʚb�K   &�X   �iپK�   �
����/���𲥁ʞv�v   F[��U-��%ʙ|��qHV%�}   �� �   �ٿC��o�l�'��    �v   F[�A   ������  ʞz�R   qH�v   ������  ��^ �;�
��/���;A
�\~�HJ�H   U.x��S   i��\   �\   U'F�s   Fߓ���������v   F[�A   ������  ʞz�������4*  ʞz%¿#�^ ������������-���4���R  ���M��о������z
C�   ��   �4���s  ���M��о������V
C�   ��   .�P   ��پU�o   �|   �z��X�H   �.��&�}   �� �   �ٿC��o�l�'# �}9  ٺM�3�c�[  %r����.H   /y�[   ��v   F[�A   ������  ʞzz��f	�A   Uʙq��ٽK��F[r�v   F[�A   ������  ʞz%¿#������ђʶZ)��#�����  /�O.�[n�t   ����F�X   �K   �^ʚ|�[   ����   F
O��d   z��O   �k   Fq�W   q̷���&�����# �   0}#  2   ����ke�Y�;��J   �� �H   ���P/��K���v   F[�A   ������  ʞz�'��/# �   0|#  2   >���ke�Y�;�
�C   ��ʚb�K   &�X   �iپK�   �
���4��=L��/���뇶���,�Ov�[n��}  ���s����;�
�C   ��ʚb�K   &�X   �iپK�   �
�� �;�
�\b�HJ���A   U�R   ������  ٺM�J   �� �H   ���P/��K���3�a3�)o���3��c�����|  ��.�4  ��^��������    �R   qH�v   ������  ��^ �+���.���+��\�HJ��U�LX  �;�
��/�"�����R�A   U�R   ������  ٺM�+��+��;��3��o��zH  �R   qH�v   ������  ��^����^���4���R  �A   ������3�ٿh�3��+���a[   �H   U.x��S   i��\   �\   U'F�s   Fߓ���������J   �� �H   ���P/��K���;�_WH  ���K�Y�/M�.M�/A�.A�7E�6E
�C   ��ʚb�K   &�X   �iپK�   �
��-�R   qHٽF	����X��UE����W������o   �R   qH�v   ������  ��^/�Y   �� '�[   �ʛt��|�[��4���l  �O   �����v   F[�A   ������  ʞz��ʛg���[   qk��@   M��x   �O   qU�D   U�����/�����/�Y   �� '�[   �ʛt��|�[�����   �����K��
  �������߾= 0 # ��.�OV�[nʢ�=V��/���Ɉ��-�R   qHٽF	����X��UE.�P   ��پU�o   �|   �z��X�H   �.��&��������  ʞz�}   �� �   �ٿC��o�l�'���kA�Y�J   �� �H   ���P/��K���v   F[�A   ������  ʞz����*H  �k�Y�   F
O��d   z��O   �k   Fq�W   q̷���&������}   �� �   �ٿC��o�l�'%¿#���������������ْA	(�3�0�����*H  �k�Y	�A   Uʙq��ٽK��F[r�J   �� �H   ���P/��K��0 !�   J0 #    	�+��\v�HJ���4��Fߑ   # �   0|#  2   >���ke�Y�;��J   �� �H   ���P/��K���   F
O��d   z��O   �k   Fq�W   q̷���&������'��.~���3�������}   �� �   �ٿC��o�l�'�}   �� �   �ٿC��o�l�'���kA�Y�J   �� �H   ���P/��K���v   F[�A   ������  ʞz���.���Q����A   U�R   ������  ٺM�3��\R�HJ�A   U�R   ������  ٺM�v   F[�A   ������  ʞz����*H  �k�Y�v   F[�A   ������  ʞz�}   �� �   �ٿC��o�l�'%¿#������0�!V�HJ�    .-�[    ْA	(�3��;�پE�;��3��    �+��<M    ����N�!����;�    ����&x  ������;��     �J   �� �H   ���P/��K���3��?A    /�Y   �� '�[   �ʛt��|�[��H   U.x��S   i��\   �\   U'F�s   Fߓ���������+��<M    ���ɂy      �t   ����F�X   �K   �^ʚ|�[   ����   F
O��d   z��O   �k   Fq�W   q̷���&��������ۢN      �;����������W    %¿#�������������\  
�~v�'  ��^M���\  ��\  ��\  '�������)\  
�~v�J'  ��^M���)\  ��-\  ��!\  '���ђ	(�3��;��3A���]  0 #  0 �On�[n�]KJ�A   U�R   ������  ٺM	�A   Uʙq��ٽK��F[r0 #  0 �On�[n���z�R   qH�v   ������  ��^�A   U�R   ������  ٺM�;�پA
M�3��� Y0 # �\�HJ���K�;��v�k�Y ћ�z ��-���y|Y
�\F�HJ�A   U�R   ������  ٺM0 # [�3��/A�\�HJ�H   U.x��S   i��\   �\   U'F�s   Fߓ���������v   F[�A   ������  ʞz# ���^/�O.�[ntX  G0 ���X.�O"�[n�W2jXn�kA�Y�v   F[�A   ������  ʞz�t   ����F�X   �K   �^ʚ|�[   ����+��|�kA�Y�v   F[�A   ������  ʞz�}   �� �   �ٿC��o�l�'���z�kA�Y�v   F[�A   ������  ʞz�}   �� �   �ٿC��o�l�'%¿#������������0�!z�HJ�    .-�[    ��~-�,��R��/�Y   �� '�[   �ʛt��|�[�/�Y   �� '�[   �ʛt��|�[���    �\   M������v   F[��U-��%ʙ|��qHV%��țO  �����/�Y   �� '�[   �ʛt��|�[�����&x  ������3����]  �v   F[�A   ������  ʞz�R   qH�v   ������  ��^�H   ߬F��   ��    �3��CH  �}   �� �   �ٿC��o�l�'�\ƿ� Y�������!:�  �y|Y
�\
�HJ���H   U.x��S   i��\   �\   U'F�s   Fߓ���������� K�M�R   qH�v   ������  ��^�A   U�R   ������  ٺM�B������z�kU�Y�   F
O��d   z��O   �k   Fq�W   q̷���&�����# �\:�HJ.�P   ��پU�o   �|   �z��X�H   �.��&�R   qH�v   ������  ��^M��3�>�D    !���M +¶��J-����ρ�߾=_��X  �3���Q  ̚L��K  �t   ����F�X   �K   �^ʚ|�[   ����3���O  �t   ����F�X   �K   �^ʚ|�[   ����J   �� �H   ���P/��K���3�ۿ5\  �t���̚L��H  �붥��.{��  ����]  	�A   Uʙq��ٽK��F[r
�C   ��ʚb�K   &�X   �iپK�   �
����΁�߾=_��[  	�A   Uʙq��ٽK��F[r�   F
O��d   z��O   �k   Fq�W   q̷���&��������j���v   F[��U-��%ʙ|��qHV%��ʸ̈q��   ��[ [  ߾F��   ��    �J   �� �H   ���P/��K���3�����B,���w  ��.:��ɖ���R   qH�v   ������  ��^/�Y   �� '�[   �ʛt��|�[������N�4� =_��   �v   F[�A   ������  ʞz�����.|�7�H   U.x��S   i��\   �\   U'F�s   Fߓ���������;�ٞK߾=n��    ���+�ۼ\  ���SU  �v   F[�A   ������  ʞz%¿#���������������0�!j�HJ�    .-�[    ��-�,����A   U�R   ������  ٺM�J   �� �H   ���P/��K���q   z��4��v   F[�A   ������  ʞz��u   �   F
O��d   z��O   �k   Fq�W   q̷���&�������	^  	�A   Uʙq��ٽK��F[r�   F
O��d   z��O   �k   Fq�W   q̷���&��������\|Y�J   �� �H   ���P/��K���;A�;��3E�3��J   �� �H   ���P/��K���;�    ��,�Oޘ[n̚Ni��h  �A   U�R   ������  ٺM�   F
O��d   z��O   �k   Fq�W   q̷���&����������W2jXn���}   �� �   �ٿC��o�l�'!��M  �+�K�ky�Y�;��v   F[�A   ������  ʞz��    ��X  E0���k-�Y
�C   ��ʚb�K   &�X   �iپK�   �
���H   U.x��S   i��\   �\   U'F�s   Fߓ���������3��\R�HJ�O�,� n��;�����M���X  qܚ���W    %¿#�R ��������+¶/)�[   qk��@   M��x   �O   qU�D   U�����/������H   U.x��S   i��\   �\   U'F�s   Fߓ���������A^@�;�^   �O�;A�;��3��z�"xKJ�^�v   F[�A   ������  ʞz%¿#���������������ْA	(�v   F[�A   ������  ʞz�v�B  ʞz���[   qk��@   M��x   �O   qU�D   U�����/������A   U�R   ������  ٺM�3��/A1�u1�u�;��6M1�uY���JJ��-�R   qHٽF	����X��UE���Q	�A   Uʙq��ٽK��F[r ћ�+¶��j-�� ��  ʞz���R   qH�v   ������  ��^/�Y   �� '�[   �ʛt��|�[�����&x  �.���߾F�H  ���n���t   ����F�X   �K   �^ʚ|�[   ����+�a+�'{�q  ��.�������ʞz�3�ۿ5\  ������3�ۿ5\  �����3�ۿ5\  �i����3�ۿ5\  ������3�ۿ1\  �w$��̚
.�+�����&x  ������v   F[�A   ������  ʞz��țO  �����A   U�R   ������  ٺM�v   F[�A   ������  ʞz�?���V��/�Y   �� '�[   �ʛt��|�[���,�������^��}��3��+��;��<Y�3�ٿH�+��4E	�A   Uʙq��ٽK��F[r ћ�����ْU	(�3�0 �@2  ��^�����[ �R   qH�v   ������  ��^����6x  ���4� =O����U˂y  E�qǿ  ����.x  ���A   U�R   ������  ٺM�;�a;�'{��  /�Y   �� '�[   �ʛt��|�[��H   U.x��S   i��\   �\   U'F�s   Fߓ���������3�ٿ]����&x  �����
��,�3�����^.��țO  ���.��țO  ����.��țO  �����.��țO  �����.��țO  ������.����O  H   
�C   ��ʚb�K   &�X   �iپK�   �
�� ��  ʞz���ۦN  �R   qH�v   ������  ��^-�R   qHٽF	����X��UE��   �+���9\  �;��3������ٺM�+�Y���������
O  ��ʘ����O  �R   qH�v   ������  ��^�H   U.x��S   i��\   �\   U'F�s   Fߓ�������� ћ�������+¶��B}  -�Ĳ����V�     �Ĳ����R�Ȇy  EK(t�[   �\  	�A   Uʙq��ٽK��F[r
�C   ��ʚb�K   &�X   �iپK�   �
���R�R��jx  E�vx  C�   �Yx  �H   U.x��S   i��\   �\   U'F�s   Fߓ���������AٹMٷ�i���ٿ�߷=@�4R��^z  ���M��о������z
C�   ��{  �A   U�R   ������  ٺM�3A��}\   l�+A��u\  
�R��bx  ,�B�����R�R��nx   ��  ʞz���}   �� �   �ٿC��o�l�'�v��r�JO  4]M��kL  �t   ����F�X   �K   �^ʚ|�[   ����J   �� �H   ���P/��K���󡦁�ۿ5\  �@����vJ�>O  p�4]M���M  �v   F[��U-��%ʙ|��qHV%�}   �� �   �ٿC��o�l�'�'vȝ[M  ʓ�z��筯ʛ�̓q��   �\]KJ�ܮ����	   i��狷�������̮���.!^  �\*�HJH�3Aۿl^  �\|Y�뽤���u؁�ٺY�   F
O��d   z��O   �k   Fq�W   q̷���&������}   �� �   �ٿC��o�l�'�vL^z  .�vț[M  �+AټM�Ĳ�����"x  �-#���;�	�A   Uʙq��ٽK��F[r�J   �� �H   ���P/��K���� q�F|  �y|Y�������>   z���������<��	�A   Uʙq��ٽK��F[r�J   �� �H   ���P/��K���sy|Y�󥦁��>   z���������<��v   F[�A   ������  ʞz�ώ���2zH  �O�[n�R   qH�v   ������  ��^H������
�\|Y�󹧁���ځ�ٺY0 �ϒ����;A_[M  �k%�Y�v   F[�A   ������  ʞz�vț[M  �k	�Y�v   F[�A   ������  ʞz�[   qk��@   M��x   �O   qU�D   U�����/������R��z   �R   qH�v   ������  ��^/�Y   �� '�[   �ʛt��|�[��R��rx   =KH�󥦁��\2�HJ�h0 �ϒ����󡦁��ɻ���ߒ����k	�Y�󡦁��+A�|�ۢN  �R   qH�v   ������  ��^.�P   ��پU�o   �|   �z��X�H   �.��&��    �~  ʞzª�R��jx  ,�������^}��;A��}\  �3A��y\  ټH�;A��y\  	�A   Uʙq��ٽK��F[r�3Aۿl^  ��ف�ٺM߾=\�4�{<>�R��z  ,�O>�[n�v   F[��U-��%ʙ|��qHV%�R   qH�v   ������  ��^�R��z   �}   �� �   �ٿC��o�l�'�'�H/B�r�[   �}   �� �   �ٿC��o�l�'�v   F[��U-��%ʙ|��qHV%z��4� Fξ�A/�Y   �� '�[   �ʛt��|�[�!���A �ђȶ^J  )�מ����r�     �}   �� �   �ٿC��o�l�'�R   qH�v   ������  ��^�R�^��-�R   qHٽF	����X��UE/�Y   �� '�[   �ʛt��|�[��B�;�_6O  ���v�v�Ϛ�����rߚ���F��O  ������BO  r�RO  4V����x   =X��
�C   ��ʚb�K   &�X   �iپK�   �
��-�R   qHٽF	����X��UE�4����M��о������.d�'�ȝ M  ʓ�z��筯ʛ�ʣ^=_�I���
�C   ��ʚb�K   &�X   �iپK�   �
���H   U.x��S   i��\   �\   U'F�s   Fߓ���������+���	\   l�;���}\  ����jx  .������R����x  �A   U�R   ������  ٺM�v   F[�A   ������  ʞz# �  ٺM�;�
�C   ��ʚb�K   &�X   �iپK�   �
������E�x  L�/����מ���țO  ������}�bx  G�L�S����'�ȝVM  ʓ�z��筯ʛ�̓q��   �\]KJ�ܪ����	   i��珷������/�Y   �� '�[   �ʛt��|�[��̪���.!^  �\*�HJH�3�ۿa^  �\|Y�빤���t!��ٺY�J   �� �H   ���P/��K���   F
O��d   z��O   �k   Fq�W   q̷���&�������L z  .��țVM  �+��ĺ�����"x  �!(���;�	�A   Uʙq��ٽK��F[r�� q��|  �y|Y�������>   z���������<���J   �� �H   ���P/��K���sy|Y�󡦁��>   z���������<��	�A   Uʙq��ٽK��F[r�륧��M[  �k9�Y
�C   ��ʚb�K   &�X   �iپK�   �
��H������
�\|Y�󥧁���#��ٺY�v   F[�A   ������  ʞz# �ܲ���,��Lrz  .�O�[n��țVM  �k	�Y	�A   Uʙq��ٽK��F[r�+���a^   .�P   ��پU�o   �|   �z��X�H   �.��&����VO   .o#[�Ĳ���/�O�[n�f �롦���ĺ����S���������
�\�HJ/�Y   �� '�[   �ʛt��|�[�����~z  ,�מ���țO  �����.# ��g  ٺM
�o���ٺM
�ĺ�����&x  �8���
�ĺ�����&x  �����
�ĺ�����&x  �䝁�
�ĺ�����&x  ���
�ĺ�����"x  �I0��
�C   ��ʚb�K   &�X   �iپK�   �
������x     �t   ����F�X   �K   �^ʚ|�[   �����   # �zg  ٺMю����BO  �ܤ��ʞzJ�����x  .�P   ��پU�o   �|   �z��X�H   �.��&�t   ����F�X   �K   �^ʚ|�[   ����3���u\  ټH�;���u\  �3�ۿa^  �O&��ٺM߾=\�4�{<����rz  ,�O>�[n�R   qH�v   ������  ��^����rz   �v   F[��U-��%ʙ|��qHV%�'�H.w�����.+�r�[   �}   �� �   �ٿC��o�l�'�[   qk��@   M��x   �O   qU�D   U�����/������L�L���%¿#�R ��������������+¶��N  -�Ķ����̮���   �R   qH�v   ������  ��^�̢���    �v   F[��U-��%ʙ|��qHV%�]KJ�� ����v   i����������.�P   ��پU�o   �|   �z��X�H   �.��&!�xKJ�\&�HJ�̦����A   U�R   ������  ٺM�õ��� q�O  �̪���    �v   F[��U-��%ʙ|��qHV%�t   ����F�X   �K   �^ʚ|�[   ���2�OXn�ׂ����k1�Y�������v   F[�A   ������  ʞz�}   �� �   �ٿC��o�l�'�玷�� .-#  [  �� ����̢���.�ώ����ߊ����R   qH�v   ������  ��^/�Y   �� '�[   �ʛt��|�[��Ħ���/�O
�[n�}   �� �   �ٿC��o�l�'�ߊ����M�A   U�R   ������  ٺM ћ����������+¶��R-����� ��HJ�A   U�R   ������  ٺM
�C   ��ʚb�K   &�X   �iپK�   �
�����^֚[n�[   qk��@   M��x   �O   qU�D   U�����/�����/�Y   �� '�[   �ʛt��|�[�/�Y   �� '�[   �ʛt��|�[���    �S����[���4� H  4J���M߶OXn�   ���[   qk��@   M��x   �O   qU�D   U�����/�������    �S����[���4�>4E�����   ���^��q�V�N�\|Y���t   ����F�X   �K   �^ʚ|�[   ����;� ћ�(«�Q   �:mR=S(��I  ��^���M �ٝ��Y�����������~zʚ}�ٜJY���|�^>���������������ْa	(�3��A 
E�Y 
O�E 	Ni���z  �A   U�R   ������  ٺM�J   �� �H   ���P/��K���v   F[�A   ������  ʞz�[   qk��@   M��x   �O   qU�D   U�����/������H   U.x��S   i��\   �\   U'F�s   Fߓ���������;�    ��z   �v���}   �� �   �ٿC��o�l�'��Jr���}   �� �   �ٿC��o�l�'�n���R   qH�v   ������  ��^��E�qͧ  ��q�K�M϶OXn���R   qH�v   ������  ��^����[��/�Y   �� '�[   �ʛt��|�[��4��   <X�ײv   F[�A   ������  ʞz�}   �� �   �ٿC��o�l�'����x���t   ����F�X   �K   �^ʚ|�[   ����;�Q;��;��J   �� �H   ���P/��K���3�ٗH�3��J   �� �H   ���P/��K���v   F[�A   ������  ʞz�'� .{����������X/�Y   �� '�[   �ʛt��|�[�/�Y   �� '�[   �ʛt��|�[�����R�������[-�R   qHٽF	����X��UE����R���H   U.x��S   i��\   �\   U'F�s   Fߓ��������	�A   Uʙq��ٽK��F[r�+��;��|��ʛ}����    �;�^   ������+�q+Y�+��;��;��3��3���[�4� =I�$��'� U��   �2H  ����|���R   qH�v   ������  ��^�����[�A   U�R   ������  ٺM�+���A�+��v   F[�A   ������  ʞz�����R����X�{[  
�C   ��ʚb�K   &�X   �iپK�   �
������^���A   U�R   ������  ٺM
�C   ��ʚb�K   &�X   �iپK�   �
�������A�   F
O��d   z��O   �k   Fq�W   q̷���&������v   F[��U-��%ʙ|��qHV%��ʚ�+-�R   qHٽF	����X��UE���
�C   ��ʚb�K   &�X   �iپK�   �
���H   U.x��S   i��\   �\   U'F�s   Fߓ�������� ћ�r �����������ђ#�-�Y>�    
�    ے\  	(���A Ni��dk  /�Y   �� '�[   �ʛt��|�[���    �}   �� �   �ٿC��o�l�'�v   F[��U-��%ʙ|��qHV%�O�[n���'�   �(h��l�   ��^@�;�[   �N�;�    �4� F�7]  �t   ����F�X   �K   �^ʚ|�[   ����v   F[�A   ������  ʞz�}   �� �   �ٿC��o�l�'�t   ����F�X   �K   �^ʚ|�[   ���	�A   Uʙq��ٽK��F[r�J   �� �H   ���P/��K���J   �� �H   ���P/��K��2zH  �מ����+A�\®HJ�A   U�R   ������  ٺM�E 
Q2zH  �ߚ����3E�\®HJ�a�CXn�Ϛ���ʓ�z��筯b���ѿ ��X��Ѷʻ}��/�Y   �� '�[   �ʛt��|�[�-�R   qHٽF	����X��UEM[  �󝠁��\ήHJ�A   U�R   ������  ٺM�둡�� 2�CXn�ߪ����kيY߾<]M���[  �v   F[��U-��%ʙ|��qHV%�ת����kŊYU��_����ʠ"=H�^|Y������
�\ҮHJ�H   U.x��S   i��\   �\   U'F�s   Fߓ��������2�CXn�ת����k��Y	�A   Uʙq��ٽK��F[r������W�̋���t�߬��� 
�C   ��ʚb�K   &�X   �iپK�   �
���H   U.x��S   i��\   �\   U'F�s   Fߓ���������띠���\n�HJ���q��|  �P|Y2�CXn�ߢ����}b  ʞr�}   �� �   �ٿC��o�l�'��    0 !�   K0 #    	�󝠁��\v�HJ�̒���/�Y   �� '�[   �ʛt��|�[�/�Y   �� '�[   �ʛt��|�[��������<A��2���6jXn!¢HJ��2���,�T  K0 # �̒���.�OV�[n�}   �� �   �ٿC��o�l�'�߲���    0 �ײ����Õ���ٷ�i���ٿ��܆���,�߶����km�Y
�C   ��ʚb�K   &�X   �iپK�   �
�� �󅠁��􊄶����M��о����/�Ϯ���������
�\~�HJ/�Y   �� '�[   �ʛt��|�[��ĺ���/�Ϛ���2�CXn�ߢ����`  ʞn# �Ė���/�碵��ʓ�z��筯ʛ��땦���̒���.�OZ�[n# �Ė���/�箳��ʓ�z��筯ʛ��뙠���̒���.�OZ�[n�[   qk��@   M��x   �O   qU�D   U�����/������Ē���/�Ov�[n�}   �� �   �ٿC��o�l�'�A��>���    �� J�������q  ��������p  �܂���,�O>�[n�R   qH�v   ������  ��^�̞���    �}   �� �   �ٿC��o�l�'��K   0 !�   J0 #    �������
�\v�HJ���.�P   ��پU�o   �|   �z��X�H   �.��&��ʳ���/e�����y|Y2�[n�������n  �}   �� �   �ٿC��o�l�'# �   0|#  2   >�Ϧ����ke�Y�������J   �� �H   ���P/��K���v   F[�A   ������  ʞz��³���/e��"���y|Y2�[n��"�����o  �}   �� �   �ٿC��o�l�'�}   �� �   �ٿC��o�l�'��泥�    ��񠁶    ��ʄ��    �[   qk��@   M��x   �O   qU�D   U�����/�����/�Y   �� '�[   �ʛt��|�[���ʄ��/��ʳ���kq�Y�������v   F[�A   ������  ʞz�t   ����F�X   �K   �^ʚ|�[   ���������
��s  ٺM�������󝣁�������������ՠ���v   F[�A   ������  ʞz# ��ℶ�.�׾�����ՠ�����.�O2�[n��*�����޳��z���.w��ڳ�� /|�+������M��6�߷=H������M��<�g�   <u��������X��j�����������[��n�����n���.��V  ��^�h����ٗH�󙣁��뙣���|e[�Ċ����H����    ��򄶥    ��ҳ��    ��ՠ��ٷ�i���ٿ���Ƅ��,��޳��� `  ��}��.���������z���.w������ /|�)��ބ��M��<�߾=I��ބ��M��/�ۄ�   /Q��򳥁ʚ|��V���������ʳ��R�����R����ya  ʞz�x��ބ����[�̖����Ė����XڔH�������n������    ������    ��ք��    ��M�Ù���ٷ�i���ٿ���]����s5�Yq�᠁�a�]���-{���  ��N��� F��   ��ֳ��J�j�����Z���# ��~���.��޳���|ն��̒����Ē������   ��.��ڳ��J�ֳ����^�����j����﮳����^�����X��Ѷʻ}����F��� ��Z�����ֳ����ڳ��J�Z�����f�����f�����b����R.�P   ��پU�o   �|   �z��X�H   �.��&��γ��    ��ݠ��    �A   U�R   ������  ٺM�É��� q�1{  �􊄶����M��о������^�����^��� <E��ꄶ�E�򄶥	X�������� ����bH  ��γ��r�ֳ��Fف   ��ֳ��b�γ����n�����z���r�n���Fݥ   ��z���ʳ��n���b���J���������}�ꄶ���R����e��E���q�A���ٿH��Y���q���n�����r���ʚ��v�����n���U�܊���,��v����Hd  ʞr��r�����r��� .)��z����箳����r���z��ܞ�����.uR�����̞����Ğ����Ě��������� <N��V���U������� ����Y�.����&�HJ�� ����� �����΄����΄��E\&�HJqͫ}  �̚�����[G�ꄶ�L��J  �v   F[��U-��%ʙ|��qHV%��곥�b�γ����������*���.��޳����f  ��懶���{�t   ����F�X   �K   �^ʚ|�[   �����9��������,��m  ��R�H   ߾=S����� <X�:�����i���̈
Z�����i���ȣ�   <u�������X�ܮ����������[�̢����Ģ���/�UZ  ��^�k�����ٔH��񣁶��񣁶�vɳ��ư���P�����    ��6���    �����    -�R   qHٽF	����X��UE��"����̪�����.��� <V����[n�V��.������ ��񠁶�̪���.��ʰ���������\~�HJ ��񠁶
�􊄶����M��о����/�׮����������\~�HJ��.��� <V��ꇶ��[n�V��.�����ꇶ��P|Y�������"�  ٺA߾Fߓ   ��泥�H   �v   F[�A   ������  ʞz�Ϟ���������
�P|Y�󕦁��E  ٺY�   F
O��d   z��O   �k   Fq�W   q̷���&�����# ��ℶ�,�碵��ʓ�z��筯ʛ�������
��愶�/�OZ�[n�}   �� �   �ٿC��o�l�'# ��ℶ�,�箳��ʓ�z��筯ʛ�������
��愶�/�OZ�[n��곥�ʘ��γ���}   �� �   �ٿC��o�l�'�v   F[��U-��%ʙ|��qHV%��M�   ̚
@��=��� K���
���z�����.m��
���z������   f��5���ټK�롣����=���ٖH�������󥣁��({  ٺM�\��
���ʰ��Ұ����Ұ���R��[�������C��=���    ��"���    �����    �������泥� U��[  ��%���    �A   U�R   ������  ٺM2�CXn!�tKJ�̆���.�9c  ��V-�R   qHٽF	����X��UE�A   U�R   ������  ٺM0 ������Õ���ٷ�i���ٿ��܆���,��³���km�Y�J   �� �H   ���P/��K��0 ������Ù���ٷ�i���ٿ��܊���,��³���km�Y�󩧁��ܾ���,!�tKJ�̆���.��b  ��J ��%����􆂶����M��о����/�Ϣ���������
�\~�HJ ��%����􊄶����M��о����/�Ϯ���������
�\~�HJ/�Y   �� '�[   �ʛt��|�[��A   U�R   ������  ٺM�������\R�HJ��愶�,�Ov�[n�ߪ����k	�Y�J   �� �H   ���P/��K���󝠁��܂���,�O��[n��J�   ̚
@��͠�� K�������z�����.m������z������   f��Š��ټK�멣����͠��ٖH�������󭣁���D  ٺM�\������ʰ��ְ����ְ���R��[��򇶥�C��͠��    ��҄��    ��򳥁    �;�X�H   ߾=S������ <X�:����i���̈
Z����i���ȣ�   <u��������X�܂�����������[�̆����Ć���/�U`  ��^�k����ٔH���������vɳ��ڰ���P������    ��ֳ��    ��堁�    ��   �Í��� 
R��������u�����u�����G  ٺM	�A   Uʙq��ٽK��F[r��q���    ƢSY���b�����   �J   �� �H   ���P/��K���   F
O��d   z��O   �k   Fq�W   q̷���&������������#_�V,�v�kɊY߾<^M��1�t   ����F�X   �K   �^ʚ|�[   ���
�C   ��ʚb�K   &�X   �iپK�   �
���H   �3�>�D    !������������������ђ#�ݜY>�    
�    ȶ�J  )�v�k}�Yن�/t�[   �]  �������󉦁�0 �׾�����ⶥ�4R���M��о����/�v�󉦁���X  ��    
�C   ��ʚb�K   &�X   �iپK�   �
��.�P   ��پU�o   �|   �z��X�H   �.��&�纵�� /r������1�Y�r�ߺ���������#z��҂��/�Oޙ[n�R   qH�v   ������  ��^������ <V��ނ���[n�V�ܞ�����ނ����ނ��.�O>�[n̚
`��񦁶[   ������#[�Ě����������񦁶�NO  �[   qk��@   M��x   �O   qU�D   U�����/������A   U�R   ������  ٺM�������󝧁�0 �ת����f嶥����ε���Ϛ���# �ľ����V����;�X�̾���.�ת����뉦����_  ٺE�   F
O��d   z��O   �k   Fq�W   q̷���&������]KJ�̮����6   i��狴������.�P   ��پU�o   �|   �z��X�H   �.��&�׊���2 K  �O�[n�Ϯ���0 !�tKJ�̮���.�O�[n̚��妁�    ��#[�ľ��������;� H�󝧁��Nӥ�������0�׾����F䶥��������^  �   F
O��d   z��O   �k   Fq�W   q̷���&������}   �� �   �ٿC��o�l�'�׮����k	�Y߾<��򂶥    ��H0�ך�����綥�� #[�Ď�����Á��;�����H�󉦁��Х���ֵ��� z  �H   U.x��S   i��\   �\   U'F�s   Fߓ���������J   �� �H   ���P/��K���Í��� E��ɦ��"�HJ�E�덦����ɦ��������
��ڂ��/�O��[n̚q��   ������ <V��&����[n�V�ܞ�����&��� ��5���
�l���ٺA
�C   ��ʚb�K   &�X   �iپK�   �
��.�P   ��پU�o   �|   �z��X�H   �.��&��   ������ <V��"����[n�V�Ğ�����"�����"���,�OJ�[nʢ�<L ������
�ۿ��ٺA��   �׮����k	�Y�J   �� �H   ���P/��K��	�A   Uʙq��ٽK��F[r�Í��� E��=���"�HJ�E�덦����=���0 ��
����e���ʞv�[   qk��@   M��x   �O   qU�D   U�����/�����������    ��H�   ̓
@�á��� K��ϖ���z�����.m�ז���z������   f������پK��զ���󡧁�ٗH��馁���馁���L  ٺM�\�ߖ���ʲ�����������K��[��*����Y������    �̶���    �ߎ���    �;� �H   ߷=S�􂃶� <X�:�둧��i���̚
Z�󑧁�i���Ƞ�   <u�̺�����X��΂���Ă�����[��������,��k  ��^�k������ٖH��%�����%����oɰ������J�̂���    �ߢ���    ������    �������[   ��.w�纵�� /|�)�ܞ���M��<�߾=I�Ğ���M��/�ۄ�   /Q�߲���ʚ|��򵥁�׺���ʳ�������4\  ʞz�x�̞�����[��2�����2����XڔH��!����n�ߺ���    ������    �̖���    ��ڵ����-�s     ћ�����������ђ#���Y>�    
�    ȶ�   )�v�"z /r�����1�Y�r�v�z�������������'�ʓ�z��筯ʛ����S����[���4�|FԲJ  ��J�F�|ʢ"=H��}�q�K��uq��}  ��.# ��/�v�fv  ��6�����6�������    �&�HJ.# ��/�r��붥���������[   ��.x�'� /|���M��6�߷=U��M��<�g�   <z����X������[����.��m  ��^�W�3�ٗH��!�����!����|e[��2����H�;�    ��    ��    �+A�<A�;��3�ٿH�+�q��;�پH
��/�v�;y  ��>�����>�����&�����   �&�HJ�ڹ�    ������v����r�:_�5�  ��5����/A�+��;�q;��;��3�a3�)x�����nr����<s�D&�HJ/��J��3Y�r@  ��0 �n��v  �>[  �� qϲ   ��&����R����E�q̊   ��&����0^ <S���[n�V��&����^����M��/�ۄ�   U��   �   ̚q��   H�3Y��ۥ�������#z /r�����1�Y�q������z������n������z������v���n���v������r���n���r�n�zʲ��"�����"����K��[������Y��   #[��/�n��붥[�   ߾=4��&����3^ <V������[n�U��&����^������J�^���������}<��4�����K����Y��;� �J���R�J�^}��������X�;������H   ߾=\�4� <X�-�3�i���̈
Y�;�i���ȣ�   <s����X��.�������[��"�����"���/��n  ��^�V�+�ٔH�����������vɳ��*����P��    ��    �;�    -�R   qHٽF	����X��UE�L�_�����-�s     ћ��ђȶZM  )�ߎ���    �6jXn�� ����   M���H�����/���t   ����F�X   �K   �^ʚ|�[   ����J   �� �H   ���P/��K���3E�/A�륡���������������J   �� �H   ���P/��K���J   �� �H   ���P/��K��������    �̢���    �U�Ħ�����[�Ħ����ܦ���Eܮ���q�4|  �V�REĦ���	L���  �r� z .M�r�zz�����.Z�r�zz������   
X0 �r�v�3E�gڥ��r� z .t�r�z����+E�<M�󵡁�U�]R��zqʹ  �V�REĦ���	L��  �r� z .M�r�zz�����.Z�r�zz������   
X0 �r�v�3E��ۥ��r� z .t�r�z����+E�<M�󵡁�U�]R��Wq�)  �V�REĦ���	L���  �r� z .M�r�zz�����.Z�r�zz������   
X0 �r�v�3E�]ۥ��r� z .t�r�z����+E�<M�󵡁�U�]R��Pq͢   �V�REĦ���	L��  �r� z .M�r�zz�����.Z�r�zz������   
X0 �r�v�3E��إ��r� z .t�r�z����+E�<M�󱡁��뵡���zY��D ����A   U�R   ������  ٺM
�C   ��ʚb�K   &�X   �iپK�   �
���Ģ�����[�Ģ����H   U.x��S   i��\   �\   U'F�s   Fߓ�������������φ�����k ��� /�Y   �� '�[   �ʛt��|�[��� ������M��о�����Ć���H������
�V��ʁ��   ̚
�3E�/M�롡���󕡁��� ����á���ѿ��|����ٟJ�ڏߚ��� �3E�땡���/A�;E�6MY󕡁��󩡁��멡���������|�[   qk��@   M��x   �O   qU�D   U�����/������V�X�;A�n# �R��ց��s5�Y �+E�R��ׁ�������V�ߎ����v%¿#�-�mJ(«M��2mN)�&ZU�:mJ� �^�R�VG7RL�S�  �v�ZiѦb�E�)|E�U��   �;A�K5�YY�r�L� �  ��ˁ��;Aq�r�Kю̬x�+Mq��rS�zx
/�!p  �R��VU�ѳ# -�c���.vѳ�W���ѡ�>ﶥ�RE�)|��U��   �3Mq��jP/�ip  �<R��VU�ѳ# (�����U��   ����ǥ�ѻ%�r ߥ?E�/6�z̚L��[n�"��)H#[���*¥��z̚L��[n�z�v�v�r�r����!�� '�V #[-�4ԁ�޾=v�^��/{�"�HJ���Jq�Mѿ��|����ٟJ���z�v�^g ��#�E ���-�ZE�����,{�4�  �^M�a�=~����.cu�
Pa�<d���?��+M�+A�+Eѻ�A E�/n#[����å�#�v �;EنV-zr�X0�1Ё�	��� ƥ�(�.ZYѿ�M��K����ٟJ���z�#A�MQ �A �������~n�;Aa�:_�_�  �Mi�r�
�8�޾=B�.9�����8�ٷ�i��z�v�r��Hѧ-�
���.e�'z��	��X��Ѵʻ}�����oĥ�z��R�~j�&ZQq�r�Kцr�q��   �^�~jJ�U�
�Mc.�PE  �/vʞrb����L�R�  �zr�
l�?�޾=DB�.dr�{���?�ѳ�3���! �A E�/mr�
o�R��#�[ �v cE)vѳ����^�<R�MT ѻ%�R ����������WznXn�[��/vC��D^YKJ�N   �������y Y��   ������$Z  �o�sXn��j  �\�DKJ'�W�sXn«U�ٸMa�:g,��j  ��J.�o�sXn�m  ��V��/zz��e�s�`|Yqs�`|Y��sXn��|�V��W�sXn�ZA��_�sXnMю��l  ����.ZM������e����!�   �&N  ߾��sXn<WQ��X  ��DKJ'�z ��DKJ��`|Y�(«R�x��Y�%\  �,z߈=](��k  '#A��O   ���������ZA[
N��]  ���M +¶/)�rʚr��-�c    �}-�    �v�r�9��7���!��R �M~��'�^Z��+¶/	(>�    �;��;�^HJ �E���A���  �r�zm��V�^�    ���J>�T    !��R ђʶz)��;�i�
.�/��/j�/n�/r�/v��k  ��z�N!�N���ђʶj�r�?� �3A�;��;]�;��^HJ>����-�    ���ߒ���-�    �/f�Y��T  ���    ����ђ��;E0 �Y�A0 �/n�*r�/v�ok  ��z#���ْ}	(�� ���h[n�f���r���b���^���?� �� �,� �?� �;��_HJ�,��$��    ���̂����    ��   �v���n�����;A�N��c  �2'�� �4� =M�G    �Y���J>�T    �@�;�>�    �;� ��ђ)��;A�>Mٞ/߾=U�V�	~   #[&�H�;E�]�;E�Y�;E�A0 �/n�r�*r�/v�jj  ��z�V�1~ <Q�<R�<V������#E�U�i�Q0 �ђ	(�'r �4R�>V�J���A�;�&Gʤ�<_�{D  �3Y�M�G�z�^�4_ER~Lـ�/r�v�r���/v�'r '����j�O�f�[EV	Ma�?_��G  �z� �^�����+¶-+#  2�k[n�/v���  #%¿#��2m^�^x   �[   
F�:mR�~n�X�J   �-�~n0�!�\HJ�o    -�[    �:mz�R�9V���
ga
m~
a�J?�r��2mR�V�5�z /l![  ��v�   ��v���_    ʞr%�i�-�s    �M�\HJY�/E�,Ec/A/{�[   ��YQ|Y�t�YQ|Y�3A�5A�=M�E%�^ ђʶ^�vA���Y�������r�����������k��Y ��v ��ْi�;A�����J��<   �;��E�;����%.�`  ��V����"v���z �W��.# �mG  ' ��-)�&Z]�CT|Y[~FU�N0v�]o  �FU�N�s	V|Y�zٞA߾=Y9��q�m9ʤS´
Lـb/zF�Ii��g2GXnH$r#^(��[  '�u�rKJ�M*��^��.s�^��8�U�~��كdѽ<X�� ��.ZM�����+¶��z-�E�@  0v�ri��'�#]���_�F�]���J���{�Rfެ<��R��/x�r�
f�XHUȹѰy�����Y�o�̓
N޾=Y<�����|͚
WUȹѰ#[]�����J�2|���/}���x �;E �
fU���R�]���C J  �2mR]ۗ J  w Y  �[C J  )�b����»�A�>M
���2mV)̓
3-�=~j��}   �&ZY/y��|<5�h�x�y
l޾=s��Y   �ѧ��|<��Y
D�x�y޾=u5<��~n!���J   .l�]9IU��   ��J   /���X%�y� �ZA��M��^7=�Ķ��7�xJ����M��hʜz� H�
�ެ=v��.`��  � =V��   ���i�B����  �^�pȸ�   �M�Mi��M��^M�
Ci��]��^7<���Y��:mJ%����~v	(�K�5~n͈
 �Hވ=���2mN�NF�.k͚
B�xb�=P��/�!z���\8q���~��Kޚ=r�OٸKb�<��Y��.f�<�ʛ|q�
���z� �Mm  ��!�ѹ!���ْi�;A�;�   .�����.Q  ���J.���/r��m  ʞn���=~z�Ip  '�0�.ZA��E  �ђʶ^�v�Y�;��;��;��E�;�   �������S  ʞr��ªA�;��^ �s��0 ��g  'Ѹ���4i  �~z�j��^  �j ��
Y ț��| �j��J[�%  �+¶���   ��.�O��[n���k��Y<��r_jXn<a��/a{)y|Y/P/�;�<EL]KJh<��r_$jXn<N��/a{y|Y/y�
]KJ���}���
�\��HJ���
RنK/l/�� 
B�� 
L0�yz��Jٶ�)�/��]KJ�����.jXn
q��U��.F�;�
q��U��.F�;�
�9t  �3AٺU߷=X�H���I   �#u  �jXn�JQ  �����|"HJ�L.pKJ�[n�*pKJ�L"pKJH[n�_GXn?Y�{�T|YD'HJ��T|Y����+¶����'��<����V���7��'��7����������M �)R � b�[n�����   �ZA[
N��������M (�mV���xU�Y�I�qS  >������8M߾.t�m.��L  '�8A[   �� �^ �5~r«�OF�HJ�R���8A.[�-z��R  >������8M߾.m�-z��{  �O�9M�8MѸ�M �0R �[b�[n=S�8^�I�����z̚L�Z�[n����������4RM�ٷ������;E���FN.zz��Kѹ��������������(�/r�n�'v��Y�r�Aa�F�H  ��}   <N��X��Y��R`�۶~��qYѹ�Y   ��^EٞJY��~��pY�Z��UHJ�~�uqYʮc[n�pYzUHJ]��x�]�[�[�X��X�X��Y��Y��R��۶~��qY�7 y��\�N�8H��K�9HٸKٹKهA(غ��m��b[n�y��\�N��X9ʣv;֍�Z��UHJ�I �b[n�qY�UHJb[n=qY6UHJb[nqY�:Ǿ�՚���:Ʋ�Ԓ���:Ǫ�Վ���:Ʈ�Ԇ���:Ǧ�Ղ�^�    Y�J��m��b[n¥�b[n�qY�UHJ�b[n�v����O�y�v����O�y���v���7 �x�]�[�[�X�X�R ����
x��5c���}   <~��X��Y��RD��즁m�>d[n¥���ZĪRHJ�I ���}   ʣz;V��YU��Z�RHJ�m�>d[n�RHJe[n�vY�8Jy��}��K��R���즁m�>d[n� �}j��Y�X��X�X��X��X��Rŧ�즁m�>d[n��8Jy��}�|�|���|�ʴ}ʵ}ʣvF�$�����۵�Z�SHJ�I �e[n�vY^SHJrd[n]wYFSHJZd[n~wY�:�F��b��Q�:�B��j��]�:�J��n��E�:�V��v��A�:�^��z�^�    Y�J��m�>d[n¥.d[nwY2SHJd[n�v����Y�Y�R ��� �}�}�|�|�v����Y�Y�X�X�[�[�R ��ђ�A�@ 'yz��[[  ��f  �\Cɮ} $&t%u�%q{�T|Y�;A�;A
��o  �C�T|Y 'ªq̓   (�:L  ��q͐   ��T|Ys;A�;A
�o  ю�8i[   ��   �wo  ю�W{  ߾�\'=\UL�pKJUL�pKJ)#f�R'�ч�����h4]}��h`v�v£羥}^�R羥!̈�^@ټu�(Ms3A�;A0fЭ�Y8A�;AÉ�߬�v4R}��(As3A�;A0f���Ѷ̓�R~V�8Q0yJ�'Э��f�vHr�vHb ���8Q0y�vN羣�B�RV�V��%�ʚa�j�r�b%[  �8YQ   ��������������ZE	��.4�ZAi��ZE��J   .l�P<{�
%
g��J   /�ʲz;H)¡��R}�х��nJ��^��^
C�th�=d6<�%�ٖM(��PM�偷�~J����M�ټM۟ [�.���{�
jh�=C��JL�.r{�
K���<������������ZAنHU��   �kՊY0��]KJ��`  ߾.B��]KJM��s�y|Y�   �w�jXnY��jXn�W�jXn��vJ���y|Y��G  ̚@��s  z��;�k��Y��sXn�G  �=y|Y�G}  ��H  �vl  �bH  �_jXn�dM�a�<vGD*]KJ~��s9y|Ycs�y|Y/{�k  ��o  ��G  �,D  �EنJ/y�OF  0�r ��	�R(�/r�Y߈<S�t*]KJ �|��[
LـK/\��DKJ��.w-����.r-�������/zz��(�����ʤ�r<V��/I
-�������.{ʤ}<|)	�����߾<Y_V�4V =K��`|Y߾=R)	���;E�;E �E �5y|YنH.s̚G�C�y|Y[L�`s  �.ZM�0s  !�   �\
uKJ'��qQ|Y߾=X��2J Xn!z KJ��   2b Xn!  KJ��   ٺY� 0�.ZE�m   ʞr�0#  �z   ʞr���   0cC�y|Y/o�.ZA�k �Y
�\>�HJ�5~r 	�~j�g�jXn�G�jXn<f��`|Y߾=x�D�DKJ(�+�r�Z�x̚
K��ʴzro�sXn:� ! KJq |Y�=    |Y2: Xn�h   'ߥ.y�G   !��
mR�t�]KJ�\��HJ!�0s��|  '�0s�A}  '��=~vr.ZE)s�\��.|����^���ђ�#A)́G�E�H  �fH  �/r̬G	��X  M��}H  z����q΃   @�"K  ��s  �;E߾U��   aK J|Y-<	.�.<  ��V��.z¡�b��g  ц߁=x�
�6r�KѸ	)�;  -�/r�;D  ��N��/>̬J0ٸF٘� �K5c|Y�kA�Yц̥
W�=�E�(|.�H  	�<V�T`  ٺ]0w�C|  '�}@�qK  ̬'<YH��U���(0 �opXn�Oz�[n¢��/c�gZoXn .j�,p  ̚'F�z���������� �0w�  �=~r��p  ߾.n�,�#S��S��[  �P0w��  '0 �opXn�Or�[nª����oZoXn�.ZA�}   ��&ZM�	k�
m^�U   ߾/hpZA.n�.ZM��q  ̚'<�M��(�.ZAaK J|Y	h0w��   (�B  @ц�z  ��V��.z�U߈<YH��U���(# �|&GKJ�\R�HJ!�(�on�[n�o�BXn���|�uKJ���K1Q|Y���o&BXn�� �)�gj�[n�uKJ�O߾=q���uKJ
jۀ�Q|Y.eȤBXn=I��uKJ
B
���H��   'ʜzȤjEXn5��|"uKJ���K�Q|Y���o�BXn���|uKJ�� ����;A�u�*BXn �J�uKJwQ�����¢'̥A0o�����'#K������@ )<P�\J�HJ�w�x�p   '#K�D   !�l�\B�HJ �+¶�R�}�*BXn�Ob�[n�(�.ZA߈=g@������~  ߾.m
��m  0w�������V �0w��'0 �opXn�O^�[n����������*m^�~v��}   <f�K`<tt�.Xs;<t�.c��ns|<Ct�.os;}<J��^��^t�/�¥M���R����¥��[   
]�|`<�?C�
���K   .�/�|ʘ|s[�P�=�D([�P�=���X�����<B)�z{�CGw.{�et  �R�	^=E�7^ =5�4F <3��<N�<V�UY  ٺY�(�$r ..�b:7�<vG1Nn�6U�7A߷=Gq�Z�i�U�<N�<J�<V.����z�V�i�U�m�<N�<J�<V.�P   ��zH!�ђʶf�r�?� �>Aن��;�&v�frz5_��S  	(�/v�9$�)�z{�CGWU�[  �~YY+c~]/#�$b /)��y  �16 F�XH  ��y  �96��]  �>90�;Y�;�[�C  ��L�M@  pDq̣   �7J}<JG7NB�~U L�k@  pDq́   �7J}F߯   p$jF߶   �'����;�
)�/^�/f�Ӕ����N���;�a;�U��   cE6&E2^>�=Y�;A�=E߾��7>�F�	V�1^� ߾��7E�?F�~�A�CH  ʞr̚S�3�ٹMc;�%����vY�� ��Z�/��/Z�/^�I�/v�/f�/j�/n�/r�rK  ʞR�'���ʙj�3����4F =PH�8_  '%���4F <z�<~�<z�<��<B�<N�<J�<V(�P   ��z����N  ђ(��O  �" ._�/Z�/^�/f�/j�/n�/r�/v������F��/�'b���;�
)�/^�/f�9�����N���;�a;�)1rd
a~M%@�r�n��zJ�����.x�#v /X#[����<~�<z(# .�/f�/j�/n�/r�/v�z  ��v����N�� ��(�mV�^��.4�"v �.A.?�.ZY�0Ma�=J��R/�'���߾/\�\|=_�NR
Q�:mN� �=_�N[
@�|=S�NXMi��YH!�+¶�2F�[n!�HJ�    .-�[    ْE	(���#A�A���Ya].+ʤ�7_E>^L��O  �?� �9A�:�^��.r!Y  -�M  ����d�/��u   '����3���4J�R�<��R�}��<����A�3�>�D    !���:m^� �F*)�.}z����{  +¶�4z �#U)�'r=J�<z-�A��H  ʞn�'R �A/}�}�/R�ɛ���<~��Q�]�L����8M2 H  �/V	�9A�E�Q�Y�<R�Z   ٺe߾=])�o���%�+¶�26�[n!�HJ�    .-�[    ْU	(���#Q�#��� �<V�����b^  �>%�;��^M  ����Oz  �4R�16�C^  �3Y�69�� ��   �/^�/b�]����ٺ]�;��� ����`   �����W    %���<��'   ��?��?� 0�������M����/r�'v������}  ���6��Y  �3��69�A*)�/W�%nJ/]�%ji_�P/d�'� /j�'� .p�י��.��H  ��ZM� �b:7�<C�1J}<I�1N^L�g<P�1F <^H�z��ђ#�)�Y2�2[n-�    >�l    ��V-�,��J�^��U�<[  �A q�1  �R��U�)[  �+E�YV�,� �[v=�<RH�Q��w  ��U�y[  0��w  ��U�W[  �8Q�y�jʛv
��[  '�]�A[  �]�xH.,�v#[�:B��d  '̚q;   H��d  '̚q͈   �?N�:B)�3�����V�7NzF��   �]��U��   ٸA���~Q �RH�Q/D�@  '߾F��   #[)�@  '߾=$�?N��R(�)f��   '
)�S�����V�/�jw  ��.(#[)�x@  '߾=�?B�yd  ��.E�\z=FH�8A
�:B��   '�Q�7����a�v�Q��   .�,f�#����_��X  �3�����W    %��H��?��=|  +¶�2�[n!�HJ�    .-�[    /)�?��v̚
R�6U�7M߷=K�,� �Q���������3�>�D    !��i�qrFϾ���� K  �ZA�=~v�[�^}�߬5W�}h�IR�ET}�Y���������ْM	/�rʚr���v�Y�3Y���x����� #�nѕȣ H  <_�K   �����'��E (�鋶��\v�HJ����yV|Y.D#.H��t  ª'̬'=s(�oNEXn�OV�[n̚
Q�}   �\~�HJ�^�#[�O �i��������NEXnʢ�=T.�ON�[n�WNEXn���~z�.YJ|Y�>][   ��\N�HJ�|jrKJ���kq�Yю̬v0
#[�g  ю߈.X�KyV|Y�ka�Y߾=O(�󁶥'�OZ�[n�z��x�RY������\n�HJ�� ��NEXnʢ�F��   �
mR��/s�kq�Yю̬
%�8m߾=].�����'�V̚
N
�Я���j��.y������8q߾=].�'���'�>̚
N
�&������.y�����8gnYXn=].�
���'�7���0 �oNEXn�OV�[n�+¶�2��[n!�HJ�    .-�[    /)�?�z��<������c).a��H   �Ƿ���
�/��QH��?��?� �3���    ��u  ђ#�юY2�2[n-�    >�l    /	(���� �}V|Y߾=L��   ���N0��,��,� ����    ����(�.ZA�x�b:7�<N�1J}<T�1N^L�g<_�o����VmXn̚
]
�5`  ߾.w�ka~|Y�|z� �^ !�>HJ�\f�HJ�a~|Y��|rZKJ�\f�HJ�ђ�<V�V�J��U��   �>Fߐ   �[
_�M �YU��   �0A~��T�V�V�/^ �?r ~�EX�V�r<x���nKJ
Aۀ�J|Y/u��w  ̚'<](�@  '/�8ER.�v�dU��6H�p�fI߁�z7J)	�nf  ٺE�;E�Hʡ�=C��ѽ��{ʺa�V��c|Y�z��zȱ{�qKJ�	^^=WK0 �jr  ʞr�v�v�R�]0�v.��r  ʞr�rp'r.x�ri�q�vl�   �AV^�rʒ�#���ےX  	(�Ei��E9́�<��<��4Vqͮx  ��M��v���/�z�G�qņx  ��zZڅ1%pF����[nʺq�XM�U�͜Ν[n��zʢy��F��O  �~��Y�3���������������1\  U��ٖi.Eʲ}=w��R
V6=H��Yq�x  ��v�
x  ��z�x  ���dx  ����ox  ��|�vx  ��pj�;Y
��\  ߾�;�U�[\  �3�^���;��zO  ��F��^��?�������{  ��pW�;Y
��\  ߾�;�U�_  �3����_  �z�U���:�����_  څI.Pɡ=z��6
[څ>U��_  �3�R��_  �3�J��_  �3�z��_  �A/j�%}/p����'r�6{  ���DrKJ��q����.g���AU��
�6_  �aʞr�E�;�
�<Rq��.�<{  ��V�l_  U��ن.U�UX  ن,U��   نU�   U�1X  ٖ
U��   6=*6.ʲrFߗJ  /�;�jv<^��v�/�ʤ�<_����6�;Y
��_  <��nA���3�U��[  ߷<S�DfrKJ����   ����U��[  <�q q͐  >	����H   ڽi�3���⃶�E���U�   �;�\   ��   <��NA/z��A<��nA�;Y

r�NL  ��񧁶
��f  ٺE�;�߾4h��   �s��Z
{ٖ@.�U��[  �vJ  ��z  '��ƴ����H   ��񧁶�;���K  �n��M  ̚'=i�^��.R��A.iF� ��������   ��|  �,� ��F� ��|  �qV|Y�;�
��   /rɡ<]��   �n�/�ʚv�n�/���������F���񧁶
��.�OGXn�/�ʞjȼ�   =N�4� <T��⃶�.�OGXnڅ./l̬G��񧁶
�\.pKJ'��ƴ��d/s��H��𧁶���	J  ��[  ٖ U��   ٖLU��   q��   6=��Yqͧ���6U��   ٖJU��[  �;�}   �uq�����[  ߷<S�DbrKJ����Ѩ߬=R�q 
J��q���  ��v   ��N   �;�ڹ�n   =����NM��|   ��������A   .E��K�K�n�eJ  ��i
@<���R�L�3��v��H   �]K  ��	�;�P   ���=V�J.��|  '���^={��>�n.r��|  'F�б[��|  'F����>�n.v��|  '����X  M��;�
R߬6MM߾:K��٬ ю���� �Mю ���<Y�� �4� 4S��   �^�,��u�/z�?� �;��;��;��3�߾6\��Q�=a���
)�;��+���s  �/���j�<�)�s  ʡGª��$}J������B���;�q;��;��;�X��
P�3��Gy/z̚D�3����Hj���4� Fߊ   ����>=|��[
O�;�w�]��H.x��b�w��|=Q��^��H   ��q�q���E/l���Ai�iH  ʞn���;��A��
�{[  ٺY��A.i��z<H��.�/v0N��   ��J�4� =�4� 7a�����1��Y=�;�
=��F  '̚'7h��/�/v�;�
��   ٺYѹ߾<��\�;�
�<R�<��<���   ٺY�;�^
[�;�
�<R(#z�8   ٺY�E�aޥ�'rF�m�����%��d[n�YQ=HJ)
[n�Y�=HJ�
[nY���3E�7M"p�K�R�K�F쾢Q/�/v�߉��'ن��;Y/{�R��� ��5~n1̚~h�
mB(�.ZQ�
mN�奁�ٺE�@�.y1̚� �	�~r5��$X�&ZU�
mJq�\)�
mF.�/�����V�v�
Nѽ߾6�!��ZM� M� ����:m^� R�A�?��/���~z� z� ������R�[��   	E�s	V|YU�M�Ѷ�K	V|Y��AUȘ�:[�.p�?� �3��;�0|�S�,� ��#[&�t#[ 0 
��.#[��b  ٺU߾<X��U�P]V���������:mR�~nB��~r<S�~z���Y -�����:mR�-~jJ��~v��}��Y ��������������%���m    �-~ z��~vѦ��v�ZA��J   .m�P<q�
�޷=��Y   �Q�ѽ��nQ��P����7ѿ­M�Y�J�������M�i�ʘzȻ H[�<F[ [�.�l H[Aۘ   �/�%z����q�
޾=�F�.Y;
���Yb�=O��.�q�
Oޚ=���!����� ���%��<�!�+¶���  �,� �<VM��O�#�޾��Fޟ@  �'v�_�4RM��CT|Y[~FUȉ0v�H����F�s	V|YUȉ�zٞAa�=l��)��
�lP  '�xC  F�8H.��G  ��V��.pF�8H.��G  '���wq̃v  �,� �?� �� �,� �?� �� M��� ����������F� H�tpKJ7Uq��M
�Ч��'�U�DrKJq���M��^��.l�����^��=��;��ʡ06d
مc.Lʡ8=��
Cم/I����7[H<v�7XJ�|<y���,� �?� ю�}���kم!.iʡ=P��-
A�;��p�����\�����4� F�1����'� �E/l�n��ʚz�n�����?� �� ]�xu	
Cf==\����^���rF�Mʔ^ʤ�/�=r��9
]ـ2.q�/v����A  �u�/v���,v  '��z�G�
@c;�U��]  ـ&U�X  U�C_  ـ*U�eX  ـ-U��^  U�#X  ـ.$Fʤ=A��4q�|  �4� �'�F� N  �{y  -����wq�$|  ��� |  ����f�����wG��u�����t����{ʡU<M�4R����)��y  �����J�A�� 
@��  ~N�;�  �tpKJ7VM	�𡁶'�Q�	V|Y�zٞM߾={������.i���D8���N  '����FT
pKJ/�;��3�߾=��)�y  ���.GXn�\'���CT|Y[~E0z�5����B�>EXn�^&ʺz̚
h�;��3�߾=M���W��)�Xy  �������� q��   ��?
@مU��   �;��3�߾=,�O?8����O  'ʡS��<_�O�Lمb/`����̚L{;��q����O  '���g2GXnH$r#^-�����'�u�rKJ�M��^��.l����̚
A�;��`�Ŷ�	�;\  �� 'U��_  �� q�{  ���o ��f���.F�;���.�OGXnʞr�s{  G�C�;��;�[   �4� 7^���2pKJ�B[  ѸʲF��K  ʲ}Fޖ   q��|  ��Yq͙�����Y
mU�Ja;�U�v_  �3��� q̙z  ���J��^  �� ~M�;�[�4V9�'r�e F��   �1[��   مb/\��<V�4� =\���K�<R���!_  Ѧ�#�مyU�X  �A�;��0L  'ɡ��=u��
cـ1�;�[   
A0�hK  �/v���FL  y��[  �A�;��wL  Ѧ��#"���� ~M�;�[�)T|Y�3��i�;�0 ��}  ʞr�'�2/p�e#<S���^�Y���Nf#=9uwެ=g�Fڇ.H`�:^�zØ��`�>{q��q��U���Ѽʻy�[��Y���:L�vQ0<�L���F�Ê��ٟN���}���_�AB���A U�H^  ��!J�E�A���3��<��<��^  '�'� .p����̚q��   ��)�@z  ���'��=$��0ʻyU����Ѷ��}F�2D�M�߯=:�4� <�4� =�DrKJ��q����.s����J  �;��KT|Y�;�
��.�pL  ��ʞr/�x�J�x��������������)��J  G<�q�r}  �4� F�K  ���'�*U�;X  �� ��
@<�i �)X  �^ �&K  ��H�#�مd/x��H�{ʡU<x��E�� 
O�;�[�X�A�;��dJ  Ѧ���'� U�F[  �� q̹   ��"�CT|Y[~F2�   �z����D�>EXn�^&l�   ��U��   �;��+�0z��{  �;��+��K  '���	�tpKJ7VM	�񬁶'�Q�	V|Y�zٞM߾=��5\مq'-����#Y'��L  �F0 #P�<��<�������;��+��;��=���o��4� =_��
m�A�;��HK  '���q����<R��-�c|  '�� q͆   ������ٯ �;�������   �4� F��   ʤ=e��*
s�CT|Y[~E0z������B�>EXn�^&ʺz̚
?ـ&/tʡF46��Y�v�B����b�tpKJ7U�   	�����'�W�	V|Y�z�   ̚
~	��^�[  Ѧ�#��;��� �5E�=_��
m�A�;��&H  '�������<R��-�  '�� 
K��ʤ8<^�,� �'� U��   �� `�;��� 
Y�;��3��v���z�J�4� ��=^�q�}/�F���r�/r���)��   ��q�\8r����<V�s	V|YUȊ�:[�=B��)��   'F�pa��/r<d���4��<J�w�;E�H4ю�\��U�����N�/v���/��_��)��   �^�3�.�'   ��)�   ʞn�'��/o��̚Db;�/vʒ��Y��!���CT|Y[(7J�=~v#^(�d���'�q�.ZA�>EXn�^ʺz̚O٘�ِNѸ��~z�z1S�CU�H�C�,�uN  '��m^�=U�=~v�.ZA��y  ��
mR)�.ZY�x�䁶�����u  ���ѹ�����ZM��J   .j�[?͚
	��J   /�L    �H����~J����M�ٿM� H[�=�����.L;
m�  � =I�   �.|�����~zb�����ZMq���?��2m^U�����~zb��ђʶZ�#Aە%]  مU��   ۅ�   U��   )�'r�n�I|YYY��J/xʥ|7[8�Kx  ���5�3�$[  ��KѨ�/�J���}��+U�r	�;]�;��r�1�uY3Q1�uYs�T|Y�4z�'���K���v=z�4z�<z�t�pKJ =M��.�:v  '�v̚
OYs�T|Yѿ�Y���%��  } 2  [ �xN  '�+¶��B�Lj�HJ���Lr�HJ�����<����$������Tb�HJ���L0��z���2*�[n�O>�[n̚
\2F�[n�k1�Y߾=_ ����綥��
mRq�\.��N  ��?'=v8�g2GXnH$qF�x#^.�����'�qF�x�W>EXn�^?ʺz̚��sT|Y�x�T8�T�Oп�T8͓���ZM�kT|Y�v͓
E`�=R�[>͓��v	޷=p�A޷=W��?
Aڇ.}	��6�bN=�FY/�o	���n<���ZM� �G�[n���;^H�z��ђ�4R �/n=A��.��J  �V'�3��v���z���J.��J  �V'�3Y�v��+¶��r��(�;�
�R/� �FZ�0K  �<J��.�r�i��'�dU�i�̬q֛}�Y���}  ��# .�/j�E�w   �rʞN��ђi�qf�]�4R
Ri�prFži��dSFξJ�.�,|  '�@dѹ<\�Nw�[GV~[�.H�6H�n�D
pKJ�Ai�qf!2�HJqݛ}�Y3E�(X  c#Y'
J��8E�qj
u� ML���[Sم-&o-� �� HѽЭ�?ʡt5K��0t��� 群�� 'Hѹ%�+¶��r��(�;�
�R/� �FZ�J  �<J��.��J�.z��4�SFξJr��z  ��# .�E�w   �rʞR��ђ�<J�R)�z�] 
Sa;E/kz��wwqݛ}�Y�� j�)[ �dS¡O�}d�H�8M߾6JH�v[  �Nj'�|J��4V 7H�n[  �.GXn�y�,z��'U�'j .z���N��p/r5Y�<V�<V)��   �<Vy��p  ٺ]��%�+¶��r-�;�.���;A/� �U~�Ii  �;��#Y��i��'�dU�Y;Eц��	)��L  ����F6r�q՛���oa�4x��.t�]9͚�z9��;�0	�<V�����ٺY�k��#[.�/j�E�ɴ��ʞj%��+¶�4J=h�4J;=v�4J<I�<N�<V�<R����ٺE��/f�/j�/r�/v�n����X�Q�]�E�A�|���ʞn�)�&ZE߁=@(�.ZE�|���.Y������ʞn������5~v�0��~    ¥�~z��J   .q�[?͚
r��J   /��[Ķ��7Y�ʪ�z���^� [�.���͚
jޚ=@�  � .p�   �
K���#��W�0��A���}�#��ZE��J   .g�K?͈
-�i��J   /��_�^ٹM����~�[}�َ�i��K��^� [�.�͈
}ވ=}��  � 
[��   �.|���^�:mR!�<�^�:mR�X ��M�~v��^�:mR!��C�~|Y m0u�0����t�ZKJ /u�U   �L�ZKJB�ў���+¶/	(0ri��#��H����WFFXn��saU|Y��TjZKJ�M~Μ[n�yL  ��E�U��   �/����zmbZKJ�\��HJ���q�|  �q~|Y�s�~|Y1�u<GT$ZKJHZ��T|Y�ky~|Y.r«�f}���GXn/cc�~|Y.e�ZKJE�.lb��\�pKJ�f��T|Y�r�G�GXn�G�GXn���o:�[n	v�^K  �obFXn#�u~|Y�|XKJ��߾=JG�B�bFXn�:A �v�FqKJ�i ��.0A�o^FXn#��~|Y�|XKJ��߾F�4H  p�F�?H  �zqKJ�)e �  �w q�n  ߭~|Ya�=K.�ş��߾U�S[  �K�~|Y�(�����	
�����ٺEa��ZKJqͨ   (�,����i���#Y(�obFXn�����UU|YٸJٺQ�J �wwA�;�[   8������N�Jp  �D�pKJ�OfU=RD�&yucJ���@s/0�ݞ��1�u�D�pKJ}��s�T|Y�xs�NfG6Y8���w`j(�3���'�W�GXnJ��D�pKJ�O`�5]Bp%}���'� .v���D�pKJq�\����GXn=FJ�|zqKJ�Ɵ���^FXnʞr�:} �o�zqKJ�i �N�e���!��B�Ý���.ZE�n   #Q���r���ʞr �	(i�pg�GXn<]M��2H  �.ZY0�8]a{aU|Y/rr_FFXnF�|H  pgNmXnF޲   F�s�~|Ypg�mXnF�s�~|Yq�W�mXnU�D�ZKJ/<Gq�W�mXnq�W�mXnU�D�ZKJ/	�]U�D�ZKJ/U�D�ZKJ)
)�pH  F�{�~|Yٺe<Gt&ZKJ.F�{�~|Y
q�_�mXnU�L�ZKJ.<rq�_�mXn
q�_�mXnU�L$ZKJ.�,j��   ٺe�<F�{�~|Y
)F�{7~|Y.�,j��)#X)	M
-��   )#X)0{#P�?N-�   ʞ&�ORFXn�fqKJ�FE�'`r�q�倶�E�U�����a�7DE�'d!�r��a�6�E�$vr�q�π���R�f}^�f}O3��Y  a�<UM�a{yU|YU�ѿ��M�a{	U|YU∱�ђ�'rH	�J(F��   �j�n�?nJю<Q��X��FmKJ�@��K��I|Yѭ� �H  ����Kч#]}���sⶥ!Э��fa+U'p"�yb�}F�[��P�]U�Y;UY��'fL/F�'n /v��^ZXn�\��mKJE�$^ʳy�A�N��Y@�r�FmKJ�N�r�
mKJ}z�4R<q�~�DvqKJ�f}r�TrqKJ�f}v��}  }j�yU|Y�+�Z�WBFXn"�BJV"�BJ_�GXnJR ��J  JN�qKJD_ |{I�>FXn�K� XLa�5TU��	U|Y�suU|Y�cqU|Y%��~z)�jM������̬��'yz���   �	 ]0Z�7���'�>̚ǹ~|Y.}�>��E�NÉ�Ѯ ���#�J��]�8   ��M�[E�&eb�<r�]q�� ��[<r�LU��}#[%�N���/H ���^ZXn�b ��礁J���/{�mKJ�FH�^GZ'x	ٽM���b�?Y0ybN��Z]��[ �r� 羥!#f��^羥���nG  �fЭ��?A3�����Y�羥�^�fU��i �xѿ%���ْ	(2�M  � �������/v#A�ז���|�GKJ�L�DKJ^   ���M  r�W�M �G��/R �{C��pXnʜZL�z  ���;�
�\�HJ�'� U��   �;�߾F޸   �b�^�Ma��� R  a�5X��cC�`|Y'(��GKJ�^  �����̚'=f�L�DKJ^�\���z  E�)b�:z �v��A �	_t�T��~���z  ��ٸMcC�`|Y&ɢ\�t�DKJM�߁7���Aه�.F�Y�H.L�RB�\
�HJ��.]����LٞV�r��GKJ�M��M����@�v�Q�^��zE�&�z��D�GKJ�M��uہ�n�<���8M�L0��t6��e�پ�
�\�HJ��ف�.i�k�Y߾=V[�   �@ʢ|<\�^>�U��YC�0MR�M�0M�=ʡ}5́|�DKJ�\�HJ!��	(��pXn�\��.I¢{�^  a�:{�V�2� =]-�Oj�[n�\��~{�^  ٽma�;���Y����| ٸMۀ�`|Y&�%�	M�cc�`|Y)<_��w  �K=y|Yi��\D�.lug
H(�s���'�.xH���^�M   
�w���юa��o�jXn<R@�"����C=y|Yba=c+�����²'�At.\�w���r�'�\A0w�w���'�H�󋶥'ʜzY�qE��|.]KJ�;����T.]KJ�W �_�sXnH   �ђ-z�GT�DKJ(/{�jS  �]|Y2zH  	�\V�HJ��`|Y�K�y|YрqB
Kц���;�
-�   �;��3��z�
� ���юʞfr�A0v�ѷ��'���;�
���M�.�^   �;�ٺ]�|�]KJ!��jXn��ђ�f�j�h �<J)�'r�    �v̥
A�Iʝz�'r�b\<�[>ɠ\=s��.[F쬿�?aXnM.r�[��.x�J�_>�[��.��J�_���̬
M�X �qx�
�̬
L�n�L8�J>F줿�?aXnM.r�[��.{�B�W>ɠ^=S��.wɠw<���/}�v̬
M�� �,B �b Fޞ   �J��z
Lڄ@/}	���b F޶   ̥
A�Iʝz�'r�j�X�R   z��qM=���qxe��H/[z�G4B
D�Hx�[MѼ�Y�4R�4VM�c+QU��+Q��5̈
G��.z�\"�/��J��.4�'f /tɠ^=e��S
s�A 
g߈=Cq����VKJz=\�_>�[�Y�h�qF쬿�?aXnM.}	��[>������.z�| ��M�����.}�} �j%� #�/�BXKJ-�S-�Y)z�M�i�r�z��ªE�.r�_foXnH   �V�O�[n¢E�U��   �{Q||YX   ��   نHU��   a�<V��юr�q͘   pD��.p	pB�>/cf<�U��C�Y��	>	.	-�Z}��²E�.L�����r�'�ZY.]	+�
m~(	��߾<T�=~n����'�ZY�"mJ(�O"�[n�نK/2r�E�k)�Yцr�
uba
CFQ/�	bf<�U����&���юa�<^M��u(��s  ��V)�O&�[n�Ki�#'�i�# G~v! n  qݚ.�O�[n̚�5c|Y.k�i|  ��/q�opXn�O�[nz��#[&�	M�cc=c|Y�dz�HJ~�pXn�t*�HJ�9V   2  J �l��2 �  # ����,z# �|&GKJ��ٸ]ET.GKJ� �opXn# �|&GKJ���K5c|Y�k!�Y%��jXnʢ=W��/T�g�jXnH/_!�   �Q   �boXn߾=X��2�   �X   '���ے�[  �+Ai��*qKJEY.uʚvg YXn5�(«��YE�*qKJq�F  �5y|YنHU��   ߾<W�t�]KJFީ   Ƞ�   Fޏ   ��"���!^  .# �\V�HJ��/m��"���!֦HJ.�Ў��'�����.��"����ϔ��>نu,W��"��������¢�������aJY�!ҦHJ)�Ƕ���J��:���%�Y
�}�����)���.�m�����:���!�Y
�o�����=U|Y��)���
�]���2ni[ �����!�HJ.��Y  ��v!�|�R��.qKJ 
������
�0��O2�[n�km�Y���^oXn̚
F�
m^��߾.z#[&�i��2>H  # �|&GKJ�\R�HJ���pXn<[��pXn �[=c|Y H�pXn�_pXnY   ��.GKJ�E��1c|Y�r�a�:N�~zb
rȠ  J ;]��N��i����ْ]�+E�3A	(�n¨U8V�����)��q�3��^|  5�'���[  �#��3��rZ��H�3�/��z#e7�3Ea�?Y�4V�IzrmA/6�rʣ^:F�   ɉ��M��h&��w<q�R_p�Zʛ��   ڭ��3E�2H^��{���   �@/x�vh#z�mA�Z^�0^�Iz�&mAY#��A�#�х��zفv,}#e!��ʻ��F��   b�����z#e��7a��r?_�V��Y#�х����za�?X��a�=1���^ER�3Eهi)b�   ڭ��2H^��{*��@/U�vhK�mٿ��   ����V�[z��_��   �SO�3A{/M�3��/A�7M�4M�3��/M�7A�4A�+��� @cEU��   �3��r��7M�4M�3��r��4A�/M�4M�/A�4Ma4A/�yMفi�3F���yM)[�'q /p�   ������v@C�   �ѱ����:@B�`�F Y�1��   ����Rw^���   ɉ���΍   SF�����@�I��Rq̠   �9c|Y߾Fޡ   �WpXn�g�[n��qJr� �     	/���D2GKJ�9c|Y�   ���wR�9c|Y�s!c|Y�>Y����    �*GKJ�	J��9c|Y�6Y�
 @�M��9c|Y�A�%	 �E���*GKJ�9J �K5c|Y�ki�Y�
pXn�OpXn�^���|�9c|Yq��o��N/�v��vʞr�W
pXnr_pXn?Y��N�D"GKJ�D6GKJ�J�;A�pXn�opXn%��+¶��N�=c|Y�k1c|Y	(�^��B��;A���6^ٟ��3���M��zGٰ���������nʛ�ʒ�z������;��pXnE��#A)g�z�a]�]�Q�<Q��NE��R�a#�/E��#A)k�z�a]�]�Q�<_��N��a�<E�X�A Aٽ]�#A��r�<|��a��v:W�2R <_��N��a�<T�qX  Ѧ́�R
]	��X  �J�H�=Y�F�/yz��FX  �c%c|Y�=Y�nʠ���=N��ʺ   �&�y3�y�B�~��   �y+�y��� �u���/i���   ��j�ʛz¤]pQ�=�����i� �zK  ��[  �3��2�]�/s���   0^j�߷5_�����3��*�^�Cq3�я����zـv$}#e r�q�W  �^ER(فi'U�   ��������&FM����j��"��F/F�v��hQ�x�1��   ������5bz����   ��hC�F�#�/u�v��hz�Y�R�R�3^�4� �#z�z� v�#vF��   ���&�M�r��M�4A�/M�4M�/A�4Ma4A/�xMـi�3B'W���4Q �xM/u�   �����@a�   �Ѱ����w5�:�u���B �\z<W���   ɉ�@!z������   �0��   ���w~�3�߷=Q�C�2X��J�3���Y���P�h��/��T���H�@<@ET*GKJ[�3�as!c|Y/y�pXn �3��v�z%���=c|Y�s-c|Y)z�E�/N����K
�|"GKJ)�opXn�Oz�[nr�
(�{-c|YJ�1c|Y�
pXn�WpXn!�?  A�zɥK5c|Y�JȥkA�Ya��n=pM2 i  !  Y )�O
�[nr��V]�Y�|&GKJ�\z�HJM��i�v��@�$z�_
pXn�n�R�!�+¶/�v)�+n�vz���&{��=����0A �zK  ��y  ���	R�	^��R4<���0z��qJ#r! n   �  �\.�HJ��/vʒ���   ��   E�-B�n������U  ����q  �	��F  �R�������^�ɲq  �F  L n  ��E�,����rL�  H�^�R�V�R�^�-�: ��מ   �􁤿͚�R�JSM�   �����h
v!����ْE�3A�;Y	(�Eѩ�*ibr�nʼ���q�^|  ��[:H  ����Ia��n�G��p���q�  ��[q�  }�a�F�;H  ����zIهv�3�,x#e'���zrv<��zV�   ������[z��_�:�Sb�3A{g�~����   ɉ����M��h��   �w<\�R_^�R�^�^�^�6R�0R�JU�[3��� q��   �4��V��^1�O�فv,}#e!���F��n�z�z�n�v�z�z�v�zrv<�]zʥ^�m���]z:{�4I <T�   �ѱ���RwP�:��   �ѱ��4I <J���   ɉ��v@z���   �1��   ���wY�+E�3��:{��A�2H��J�+E�8H�<��:{��[  i��  q�`  �VW<J�[���i��/n�r��z�5�ـv,}#e ��HU��   ����M��eJ0A�1Ma1A/9ʤ^:D�   �Ѱ���=\z��_�:�Ta�3A{g�{���   ɉ��xM��h��   �w<\�R_^�V�R�>^�8^�^�>R�8R�<J}<��<J��^0ʤA?Yv���5�z�V��!z�v�z�z�v�zrv<�\zʤ^�q���\z:{�4U <T�   �Ѱ���Rwp�:��   �Ѱ��4U <J���   ɉ��v@#z���   �0��   ���wY�;Y�}�f�0 �������+¶)�E�3Y�Aѿ}�a�?RE�U�1[  ��J   /j��|ʸ}ʣv;s��Z��HJ���}   ʳz;V��Y}��Z��HJ�m��0[n٥Z�FHJ��"Y�HJ 0[nj��O�y���|��|�|ʜ}ʝ}ʣv;���Z��HJ�I ]��x�]�[��X�[��X��X��R�۶~��#Y�]��x�]8��|هA(���m��0[n� 6#Y6HJ0[n#YHJ20[n#YfHJ�Ԛ���:ǲ�Ֆ���:ƶ�Ԏ���:Ǯ�Պ���:Ƣ�Ԃ���z�    }�Y��~��#Yс�#Y�HJ�0[n�#Y�;A!����\�N�;A!����\�N�8H�9H�;A!���I �O�y���|�|�v����=k��&G���J   /Z��|ʸ}ʣv;W�����~�i!Yс���m׮3[n� �J   هM(rʺ}b��m�V3[n�~�i!Y�F3[n Y�HJ�Y]��9J��X1ʣv;샺���~�i!Y�7 �8Jy��}�|��|�|ʴ|ʵ|ʣv;փ����~�i!Y��Y]��9J�8K�9K�8H��K�9HِJّJهAU������즁m�^2[n� � Y�HJ�3[n� Y�HJ�3[nM!YMHJ��b��U�:�B��f��]�:�N��n��Y�:�V��r��A�:�R��z��M�z�    }�Y��~�i!Yсy!YbHJ62[n!Y�;A!����}�}�v���7 �8J�9J�8K�9K�;A!����}�}�|�|���v��H�=~r�.ZE�k��Y߾=XM�Ѹ�(#[ �.ZE�
mV�\"�HJ��.|z����0�
mR�\��HJ��.|z�������Ly=yj+¶��R-+��#E�;A�>M\   q��   ���J�����
��:V�2R���
(�r?��^ =(�Y�*�^#�#EQ�=iu�A	�����ٺM�Y-��ض���R�E,H�:�R�����z��=E�*�R�2R�E,�}Օ��    �F�H   �k�Y0���論ʞv�    ћ�+�ZA�W�b�?Q
�$���ٺA�M -�
mV)F�
mN�����-s̬J0ٸF٘�i�ʤ�>`ET nKJ	T0w�vƶ�-�����@ц�$ƶ���V��/U0v�opXn�Ov�[n¢��/\�gZoXn .g�����̚'=N��	 ��R  ٺEѹ%�i���C�,���#L��M  '#Y�f�=~vro�sXn:��Ѹ��{ʺa�V��c|Y�z��:�^=)��S  �.ZQ�
mB(�r   (¢��@  ٺ]ѹ���g  � S   ��C  �^ ٶ���
mR)�iS  ʢ�/s�!g  � S   �d�
mN �
mB.�OV�[n¢���A�k]�Y�|z���.r��Q  ٶ��a��E��_���r��GKJ�M��-�z��:�^�� ��=~vro�sXn:��Ѹ��{ʺa�V��c|Y�z��:�^=)��P  �.ZQ�
mB(�r   (¢�E@  ٺ]ѹ���f  � S   ��B  �^ ٶ��ђȶjM  )z�G4J�4��4�Ni��<  �R��_�U��pXn�vʺa�n��Y��X�jzi.p#X)�/v�������V�JY��z�U��   �;EcY�;��AU��   �������3�q3Ea3Y)W�����S��PN�;�� D�A���륡��q�ȣ M  5���������q���# .�ߒ���
�J�Jy�km�Y߾=���E�&u��brrn;�M��;�a�F��   p'v=8LG<R��^  � w   ��i  �y�?�Oj�[n�v����)�Y�E�N�OZ�[n̚
B�;��A�;��ٶOj�[n�v�Ɓ<R��L  ����e�}�NM
E�;E�FSU�㤁��8^  � b   �i  �q��b�%���LrXKJ J  ������2m^���?A.s�rA�?Q n  �X�7E^�N�R�B|   �v�;z ���:m^EL�DKJJi��Ѷʺa��{�^��V��c|Y�:�^����:GKJ(#N��N� K  �\E�'y�)c|Y0z� ����6`Xn̚'<{M�|:GKJ������s|Y߾/v#@�ꁶM���YXn�O6`Xn�^oʚ^ʛztBmKJ�i���nKJ��ѿ��{ʺa�n��c|Y�z��z�ن�.z̚J�t�ټi��RoKJ���.f  �t�]KJ =_�M  ��~z��nKJE�(it�lKJ	Yq���{ʚb��������z.�Of�[n��:m^��NBپU
��遶��ZAپi
�\B�HJ��ZM��YXnr�^g�[Xn>JU���LپU
��遶�ʚ^�kU�Y��~zʢj4Q��F.��Ͷ�'��:mR��z.�Ob�[n���	(�VYKJ)�k��Y�C��Yi�pGvnXn=T(��Z�����0�E�A�`   �;Eߥ.t#I�v遶�J���;E �ђ�v̚K��gFoXn /l/�3E<��� >cH�v��v�?v  �KT|Y
�VH
iX  �K||Y�k�Y߾=\�4R =T��N  � c   ٶ���������������	(�ZQQ�<B�~j�ZYi������:mV��ѭ����"mN�~n�ZE��������B����ª�-~f�~j��}�(prZY-v;]E~r?[0z���%�J ��������-�Z]Q�<B�~n�ZEi����~v����i��
���"mJ�~r�ZA��������B�����-~jحmJ}�(prZE-v;TE~v?RU~nRZ]q:mRe~r����٤ �Y +¶�2Α[n!�HJ�    .-�[    ْQ	(���RoXnz�E�/@��0�Y�\��HJ��.z�T�;�
(!��HJ(�k��Y߾Fް   #X&�vXKJ��Xm�;Ua�<_�q||Y�]�Y�E�A
�\��HJ��   نHU��   c#Q/v�XKJ�B-�Y�E�;i��R���R>�Q�k��Y�;�a�=9���u ��پJ~��]߶��,�����-��H  ʞr�QH��?�z�M��3��E�.W�/��Y�E0�/f�O��[nr�
Y�]
(�/v�O��[n�XM����3�>�D    !����	(�VYKJ)�k��Y�C��Yi�pGvnXn=T(��Z� ���0�Y�E�A�a   ʞr�ń
C0m�dζ�'�Y(���J!#���	(�/rz�E�.kpn=J�O`�<J�RE�.}/�fz� �pGFoXn<I�RE�.y/Uȉ<�H0���W>EXnF쾿?H�
�2GXnʢ7pGJfi�pvFϿ�A
(#S�|XKJ�\��HJ���2GXn<�GJLb H/�+o  � p   �����i�pvFϾ�A00w�o6oXn�O��[n̚q�"������������������*mV�~z̈
i��ZA��لM(S����Y
Aq��]9I/���R}�Ѷ��nJ���ٜJ��K.x����.x�]9/��ZA��ZM��tpKJ7TA�
mR�@���'��:m^�DrKJ�M��R�ɣ>:O��zOUۋ���Ѯz���E���M�i���=~v�r��q͝   �	U��   �|=Pri�8E��   E[�V�r<S(�t���'�_�R�O�Q�A�Y�-Z  ʞr�z̚
&ن�.�r���<m�J)ʣ�=M����LٟV�B��GKJ�E��uՕL�6FXn�zڟ�ڇ�/xɔ^�r�$f X  /j�r��v=V��^N�8Q n  �G�^q�[?�T ���R���J��JwV�/^ ʒ��-�ZAم�
�
mJ�V�H/v��
{�|<t�7R <](����'�\ER@�~M ]�O�8E
X�p�\FQ.q	�xʒ���T�O�f�r�zm�rH�8Eѽl�   ����(҃����D   ª�V��y��vjrB�(��   '�r�EѸ���ZA�����
mR�񥁶'�	�~vz�+��.}#J&��z=XrA��A.|E^��J
KV|��^=XrH��K.{D  A q��(� V  � J  j�� X  .aȠ M  =N�� v  
Aa�<Qu��yB��JڲHy�.ur�EW  [ �_s  | #��n.{D  M ��"mRM���J
J0��A.|E^��^
KVv��|=XrY��H.|Ez��  A 
KV|� Y  y�� |  
Tۇ [  .lr�
@a�<W��V�AڲA�}ɖz��  J 
Eۇ   /xB��KQ���  z 
JڲY�-z�GTbXKJZ�:mR��ن%*ʚ^�(�VYKJ)�k��YccA}|Y�C��Y.p��#I�.�H�=~n�D   ���~n=PZ��⥁�}���ZY �+¶/�gFoXn 	(/c�vʢ?F��   ʢ$F��   ʚ^��   �R� [  0r� 4G|pKJ~B-�6���'�t�rKJ�M]�߾<^����O>EXn��Rq����.q�?t 0|�v�w�w�?w �#AѸ0 ��#Y/�;A
)�oFoXn�Ml  ��z��.�r�OU���DU��q����vB�!���:mR(#z���#E���:mJ羣'�ZAq�ʐ������j�/bـJ'o�^��b <T8ʚzʤ}5�H �i���~v)#z�~j���ю�Z]É��B�VHU����I��m  ��V01F�u���.k0�m��I  ٺE��^��'�%���/�r)�"�#z'�?� �!H0^ Э�#E��ѽЭ��v0���^��rb�$���n={=�A�j���߾/p�A�0����;��V�������#Y'hJ��>r�E�+Aq��f�z����;� ���ZA�2m^(#YU�Z�y�JHپM���mRM������ZMi��b <W?ʚzʣ}5�H�z��ђʶr�r)#z�4R%ʔ��ѵ��J   �����rЭ��?r Ѵ��U����]��y�����Q;E�y����^���3��;E/��'�#X%­A��XE�&q�vU��zY�zX�y�v�~ ��^� ��ђʶf�v)F�6CѧȻ �  �v�x���|F� �'nȹ�6  ȱ�v  ����nȡ�����<|��M�
�O���߾U��   �;�
�����K��   �;�
��.�퀶��>R��.�E�����J��.
�9MѶbvr�E�;�
�ँ��ua�6eU�ю���;�
�?����;�.�􀶥�>R��.������V>�;�
�ݤ��ٺii��&���EV&V���(����-r����;�
�$����	]ٺEYI#[�����	E�	]��%��.J��I���'z�VUV�6J���3A��R���   �u�Q�ف	/s�r���+z�K�Cفi/{�r�k!��2�ZXn�.ZE�
mV�ˤ��ٺE��I|Y�
mV�=~r�6�����V�ђʶrz�.
.�/r�r�;�
�H  �A�;�
�奁�ٺm��ђʶrz�.
.�/r�r�;�
�@H  �A�;�
�ܥ��ٺm��ђ�n�#E�<R�V)�$�\Ń��$a�vz��Xެ=\q��?�YyZ�Y�R��+Y�^ ߥ5H�poD�qcL� y��� �wkL�<M�l�����	
)�ҥ�ʞn%�+¶��r(�v
��.�   '����
 0oʶr¦��<ۡxh  �<J�4N�Rq���\q���z������ٺi�~EѸ�����V-�x��y  �� �  ��zj��V�^�[Uɐ�   �l��F ����.mr�
A�� f  �V��  �hi�r�[a�<T�R�^�Q<�R���Hf  �#�Ѵ��k��uB��Ru���Q�^�Y߰<G�YY���Eu��r[�v�zȝ��  ���3EQ�/�6A ��#X�O�����g�sXn 	(�o�jXn.̬RcK�y|Y.'��i  ��/.�o�jXn̬
�"mJ��.@����ц�\��.Q�%���r�'?M�O�BqgF-�^  ʞr̚
LٸM���\�b�XM� �+¶��B-P���/v��  ��ETJYKJ'�v<]M��H  ́q�  M��ZXnpB
=پyC�N|Y&���	�\��HJHE�U�h[  0>�:`Xn M��>aXnp/�����GnnXnFܕ   �'� U��   �3��o͈q��   q��F�r�q��   ��VKJz	���?� 0>i��VKJ�}�⛘M��׊mKJ�r ��.R�͈
lU�HUȳa�>N�����mKJv�VKJ>r��?�c <�����R�4�z;��R�LvYKJ   �nnXn��   ���mKJ�i}|Y���:`Xn�,�0� F�9�����VKJv	g�   ;�-��   '�WKJ�|vYKJ�N�[e}|Y M��^nXn��բT�t
XKJ =U��   ��   �ր�����P�LꥁѸ%���~z�.oXn ن�/n�_.oXnH   �[��Yن�/n�_.oXnH   �[��Yن�/q�XKJ�L
XKJ   ��:m^S�Y  .\ʲz=M��W
E
Ji���zM  ��lM  ��zA  ��oM  �	M��>aXn���z��i}|Y�nnXn�vYKJ�s|Y����ђȶjL  ��
�|JYKJ�\��HJ��[q�L  M�� H  ��{����E�(����ߒ���i޾=m-�+�U�CUȉa�>GU���L����?�z^iz����K����Y��<��͚�%# �̶����|WKJ�|JYKJ.�ߒ���
H�q���# �̶����|JYKJ(������.�Ks|Y��A  # �̶����|JYKJ(������.! |  �|WKJ��R  ٺi��ג���/�o��=L��VKJn��{������	}|Y�b��|=J��VKJ^��{��������>nXn ?a�;�Ii��   ��Pن-j��?aXnYжɛ^��>nXn�E��;Zن3-p��?aXniжɳ^����YKJ 	a�;� ���t�DKJ <H��f����{�`|Y[   �i�pG*oXn2��[n�O�[n¢E�.�o�[n!��HJ)�����*oXn=
��Y��2[n�&oXn���||Y�&oXn̚
_����.p�XKJ��.{���=~f�.ZQ�
mB-�O*oXn%�i���+¶��V�R�,� 	(
.6=��^
ٖJ.Bʲz=p��\
Q
Aٶ��8H  �GoXn�2XKJ��c-||Y�oXn�o�T6XKJ�%||Y�V��׶�����A�lH  ¢'ʝv�a�G�T:XKJ�)||Y0��H   �֥��/vمH/h�'� U��   	��Ł���   i�r�]c3�.v#[��Ł�J��ҥ��vʢv=P��Q
LنM/e�*ʢv���*<���   ��ʢv<m�D�nKJ��J|YY�r�a�zI��K�(پE�K� �O�YXn�g�YXnY�r���|�U�4� =RH�k֥��ARB�0v��'�l�/v���4Ru.x�'vM/l���'vA�8/x���&z�!���*mR�D�nKJ(�.ZAcM��.l�f7�f�ʚrr�LcM/��V7�V�r�LcM.|z�!�(�,   �~vz��A��]XnrR
kپACQL|Y&�ʣm;x��~	T�<   � s   ��|   �r��jKJ �R�ȣ�   ;O���   	D�k   � v   ��A   � _   ���ٶ���R���ٶ���V��ZMED�DKJ):����L�B��GKJ��ٞV�J��y��|J��	^=m�q�
{�C�y|Y[Vi�b�
Y
AZ
��v0��Y.#��\�HJ�N�ry�M��h�ف��� S   �ȥ���^ ٶ� ��:m^EL�DKJVѶʺa��{�^��V��c|Y�:�^�^�=Y� ��v���� @   �C����z ʒ���:m^-��E��_(�J��GKJ�U��pXn�f���|J��7R <yX��ե��$v D�8E
�\J�HJ�RX�vԥ��}�FE
�\B�HJ!��ZMѶʺa��{�^��V��c|Y�:�V.�Ob�[n�	)#XM��ե�0}cC)c|Y$#�6`Xn­��X�M\��.?�r�.s��F  ʢ�.
ف]&W�WKJ�M\��z.�Oj�[n�WKJ�}\��Ɓ��6`Xn�ZO 9rgpXn5� #X�Ɓ���%��=~v�]   ̚'=_��� ��8D
F�Y��F  ��'A��i��-�
mVM��V��ٟJڇK/I/�vH.O�v�dU�߁7|)�Y�ӭ��ʞrr�G�8E��=TZ��8E�y�riٵ��8A�M �O��%�0�X   '�	(0|z�M��/ҥ�z�'popXn7.�s|Y�z�߾=�	V�=.�񮥁�WKJ'�z��6E���.N�&ZY[F
�U���ن�
T�S�mJ <I��X
G
�H���ن�KQ��WKJ�}�(�˙��'E|:GKJ�0|�v嶥�5~jH��.|!��
mRE|�DKJ	Ѱ��_��E�E��pXn�^���M[
l(����=~f�.ZQ�a   �������ʞj!��릁�� @   �޵���z ʒ��+¶��V�,� �'n 	�V(ѭF��H  �v��E��_�}��M��pXn�f��c|Y��KY��z��|F��H  ��6=G�	_BC.h�n�Y�N�-H�;�[   �j{C�;�0 �y�/n�Jy�k�Y߾<c�\N�HJLE�/j������ S   ������N�J��7q�~  .�2���'ʒ��M  �N�+�[+��2y^�jz��q͢   ��.w�at<^rM�|m��H�;E�3��;YY�r���qʑ   �J� fdF��   uW
B�}
�;Y��   Ic3Y)f�n	�FC/x�nK� �Ys
�;Y���# .�n��#[.�]�}j�\�HJ��/t�Oj�[n̚�� 
�y�NM
Z�;�ft=M�JW�F�k{�sEVB��PL�}C�f#[��A����ʞr�'�C.z�Ys
�3�c3YU�����n�]�=jz�\�	/zEX�Oq#E�#��;��|z�!����0�!��HJ�!Y>�    
�    ʶb)�?�z�Gt�XKJ)#[%2֑[n�   (�k��Y߾=R�T�XKJ�k)2ڑ[n�\�HJ��U�k[  �{�||YX   G4N~Y�]�Y��H  �N��||YنK/c�/b�/f�/j�/n�/r�/v�Oʙ[n��   ��[q̉   G4zA�6oXn�^�<N�<J�~��A�ʺv	
�<z�\��HJ���#�a�F��   �'��^eʚ}m���݁���Ѻ������m#[&���i��'�����#�c�.���]�Y0�/^�O��[n̚
)���E�A�k��Yю�/�r�
{�;D^
	cUU��   aU%`�/b�/f���E�A�k��Y߾F��   z��,����W    %����   �^Hʚ}m��t݁���Ѣ������l#[&���i�z�����/�r�
�-�/��/��/r�/v�OΙ[n̚
�cU)<^)�x�/b�/f	iX  �i�k�Yюr�q�+����������ZA�:m^����
D�F .v	яI߈<��q  <_U~z�Ѽ��*m^(�.ZEi��VLr�Ma�:YH�~n�t��=~v�mJ(�m������ʞr̚
^�8M
H�N�큶���V��.}�v�z�	M�N�Ł����V��.}�v�v�	A�N�݁����V!��~z�y�MѰJ��y�Jv��VQ��v�9^��E��Q��6A��ZM)�
v�z¨����V��B��^�A��V����u��R�A�ђʶn�r�#Yi�r�(��  �m�	z�	v?)�n©�4���	ۡ*���-�0�����.�|����$����v�?� �� q� ����.�����ʞb�v�n<�M�GRa�5Mѿ��n�v�Y����Y��YQ���n����  �M�}��� �  �A/n���������  ��<�� /�=C����ْ	(�Y�;�0��z�$�����������������������'n�U��z
Fڇ@.tɣt=_��WJ��0z�aنBU�>X  �Z�D�HJ��kEڅp%y#Y�TX  `cT|Y/y#_�X  U��ٖb.`
GٖJU��X  ��   #X�� �  ���?� 0|��ɡO��5_��c~�`cT|YU��   څb.OɡS=v��j
څ
U��X  څ$lɡF�K  ɡF�K  #\��[  B��H  ɡO5S��cq����DT
pKJq������jq��  ���c�����pO2GXn7Kq��(��᥁HZ�G�s	V|YUȊ�zy�̚
W��CY�;��;�ڕy�;��f�Y���V��`cT|Y/������� ����Dڅy/v���E9��G\pKJ~XUȊ.�ֶ�'0�p�W>EXnF��^?j���.b�'�P)o����ɱN�����B�V��څbU�C���څdU�H��������pO2GXn��7Kq��(��HZ�G�s	V|YUȊ�zy�̚q��   ���)��ɡO�n5_��c~U��ٖb.

-ٖJU�F[  0v�?����jL�a��ɡOF֌   ɡGF՗   �P��kGڅp%w#S&�ƴ��ɡN<���i 
cU���1�ٖb�3Y.jq��   ���#]&�Ӄ��N�ȧ��0t��Pq��   �&����Y��   ��H   i��g2GXnH$qF�#^.��ض�'�q�W>EXnF��^?ʺz̚
UU���z��
���
j  L�a���j  �<��tpKJ7Uq��M
�����'�U�DrKJq���M��^��.{�E9��1�X���;E�� �qU��   0fc;�,k�'�L&}�������;��}���'� U��   �q A�3��;������;��
�#����;�i�ʞrp�4X��Y;�c3�/}Jfp�<YUFCN  $N��H   �#Y�Y�;Y�+Y�� 
)i��  �   �i���K   � tꕶ�@�;�[   ���]
��.��y  �����<�����V��i�z�M�i���M�i�z�M��;�^   �\�� 
Fi�z�M�i���H   �3AQ;��8\�X�t��<�X����HJH�[n��Y��HJl�[n��Y��HJw�[n��Y7�HJ)�[nj�Y��ْU�;Y	�F(��%  ۟ �  y�/߷�;���������;���������;���������;�������v�;�[   ��.x�|d�z�|i�E<��/`̥ScA/k/�] �=Kz�
Y�zy��H  /a�< �   �<�J[ r�O�A 
F��   	/y!r�HJ�<��.kȥ   �<W�4R <ti�Y�qr�j�A T2f�[n�z�����=J_'�?� �H  !J�HJ�
^.�ȶ�'�}O��Uɋѱª��B�J3  ��R�?� 0�V0/�+�1�����HV����R��J��q����
��.��{  ��V�'��eY�;�.����J  �B/�M=K�4Nq��}�߁6R������]ف\$}#O!F��ې�e  <�,� �bA   �;�
�����3U�߈4M��ۘ�   $s��������1H�=M߷�b7
�N�<��4R���;�
ۡ@�����.�K����R.���ؾ������������b�?� ٺ]^N�b�j�[��;U�6�6ɣK�z5jE�(q�bG<\� j6��E�)z	<�J� c�RJ�=JU���Q^ ��%��E�(r�bN<Y6��E�)�/�] �=Kz�
Y�[N�9{ 0��ђ�'n /zz�#��KY}|Y�Y�E�Y�A0�o:`Xn��z  ��F��/y񥁶%#�پ��	+�K�y|YM��xr�
�c�Y)�
)#[��іr�
w��с�a��:mJ
f)
��H0����.`�
mN��\  �8MٸME��i�#�ʒ���(�.ZA����V>=\�/V �M(�Φ��(�J   (¢�����ٺEѹ��
mR)ʕ��r�.J����ц��w  �?J��R  ٺE߾4_����[�8U߾=Q.����/F �E �� �	�~vrG�sXn;ѽ��{�f��c|Yѽʺa�n��]��X�jzH.,������]'�NM[
`	�ʹ��.�O^�[n̚C�k]�Yю�XM�߈=O������N������ S   ���-�����'�G�̤��� w   ʒ�%���ђi�
.
.
�V�I �KP�=]<F�zm���/vʓ���OP�=]8F�zm)���z ������(�3Y�X�4R��i���Y�¤�<V���8�i�s�>^
M7���� ����������+¶(z�.
.
.�+E�7 �|C�
Nq�^Z���<R�OP�=P8F�zm)���ʞ^��ђʶZ�#E�<R�tz�)��������/�8Cч�  M�y�j��� �  t��N�vF��H  /ۇ�%q��  Ƞ��U��[  <���A>^M��D/߾󥁶%Q�;A�(A/nz�G^Bcx<]�&[  i�/a�<D�R�R_c=M/opYD�8A�8M�x�1  �������V{   ��J��4V 7}��5A�;��;E�3��;��;��3�U� U�@Uш�3�ٿ�.�k�����ٺE߾=\��� ��|�7�K�3�/���K�;��3E�E ��;AX�  �'v $[���/f��������v��  �'v %�/�A p�;A��  �'v 'UF�;A��Hv��=Y����.�����5/��'� .z��H<�4� �-q��l��H C � /K�'��/R�?� ���T�� �'���B�;A<�� ɱp/�;��v���Y���Rt�:A��B��T���X���\�t�A��e��M ��   ��� ��%�o �7R!����ْE	�yB|Yi�ʱpr=9Y�;E��PXn���V��:GJO�;A<�Ac3E.?�V���4V}ʺyr�
n�z	<�u� ��J�(r�'���۶��/��A����M�c3E/�%��+¶�2N�[n!�HJ�    .-�[    ْy	(��i�pG�oXn#[!<)��HJ.
-�k�Y߾=R�t�XKJ�j��Y
)	-�Oҙ[n̚q� |  �L�XKJ|   �/jr�~Y�<J�q���'ª�<NGF~Y�U�Q�_����Fߡ||YنK/e�/b�/f�Y�E�A�k�Y��H  r�q��  GzA�6oXn�^r�
@c#UU��   aU/v#X&�"  G4F~Nѹ�6  E�%?���i�k��Y߾F�/H  r�~e��Xk�;�b#�.d�
s�
Z�3Y�wsRM`�?�>	bf<�J��pb7k�4�|;���F�
��.H`�=��B�@`v;RD�U�1���>qB�����	(�/n#S�<z�\��HJ��E�U��   �#�Y�ʚ}m���,����Ѻ������h#[&���i�������]0c#�U��   �����<J)�/^�o��[n����.	�<F�<B@�i��ª�<�E�.�'��^Hʚ}m��;,����т�'�����l#[&���i�z�����/�r�
d)�/b�/f#[�<z�\��HJ��.h�<��<��<V�<R�\�HJ�Ki��?���-�s     ��ђ-M�cA.+#g�<R�\_  юa���.>p/v=a��y|Yi�qFνr_�jXn<V.��  '��]KJE�/*p'r=CGt�]KJ
X�3���̚
wٶ� ��r�q�V  M��ʥ�r�'��]KJ
��Fpg�jXn<IM��ʥ�r�'��]KJ
��Fb/v�g�jXn�'��A��   ª'̬'5�v 
wߥ=h�}��u�s߁��v 
B�9M�NٹM����X.�/��]���'̚'=f�|�;A�z��Ĺ3߈4X���z�R   .��ȥ�߾U�	����3A�r���^ ��]KJ�4V =�<R�B���>�Rʥ�ª'̬'=t�<R(��ն���UR'J��z 	��R���y��\��HJ(�����'z�������|�]KJ)�\��.S�&ZY.�.Z]�����ʞr̚D�x�^Fug
W޾=@�^��^��/�UL�]KJ��X�� �Ѹb_�jXn��|��)�&ZAi�̥Mi���v �^
C�nپM߬<�-�z�^   (�˥�ª'̬��/v#S��%���Nѡ̚
Z
��^��Y  �x�Y'ʜz���o ��#��
mRE|�DKJqѰ��_��E�E��pXn�^���M[
T(�t���(�r   (¢�6���ٺEѹ������ S   �w����^ ٶ���
mR)�̬��ʢ�.Bʤ=_��X_0|�����Hц�ț��'r�'=F(�ܛ��'�kA�Y߾<P�\N�HJ���|z�(�������٘V��L�M��pXn�V��>�M ��.r�<���ٶ��|z�!�(�.ZA�8E��=G�A.g�,v������<r��M��O�8A�8M�������������ђ-�/r�'v�_NoXn�"v /E����P�=t�O�nF�.�eBS@�ɻ^K�zܞeBS@�ɻ^K�zb�=�d�F�F侢"��_rnXn�gvnXn %z# �\��DVYKJZ��ȥ��^ZH   �   z��C�
n�x�ab�=�.������^����ٺMb�=�e�٦�ѦQ�<S��WrnXn�PZ��ȥ�ʞz%����(�3YQ�Fޗ   �/v�'r�_NoXn�"v /0���^� �|t��y={t�.cF�(xq�	KX�q�Ob�>X|�b�<W7<�M�b�F��   𥁶�q��   ����   ��{E}|Y�CA}|Y M0 �C��WrnXnZ��ɥ��^ZH   ѵz�M�с�\u��a=yu�.a/	�=���Ѧʞz�0�����^'r�@�i�r�
@ぶ��;X��u�/w��sE}|Y�pZ��ɥ�ʞz�� ��ђ�gRnXn 	(<U�<V�<R��́�'�,P�;ɥ��/v<q�D́
UȊ��r|Y^
S�8H��.cF�F쾈�vB�GV
P�vF�pr=F8��P�ɥ�i��P�+ɥ��8��f#C�ځ��;Eq��U���R���y�#��=~v̬
W�0���.��~��'̚'=Q(�; �i����������������HJ�T  ْy�;� �3��;��<����&�HJ(�}߶�'���=���� ��.���L   ���Y
���[n���� �HJ��W  /��)«.�/���y|Y��:���v�?� �~E0 �Y���y������|&�HJ��0 ��������\�[n!�W    ��z ⒏[n��s  /я�/��\�[n�?� 0�r�'��������)���3��W    ��+¶��F/���p   ���Y
�{7�����ඥ��ZA[
N��*�����M («�=~v�ڟ���O*�HJ���M � �Y��E  ʶN��0 �����������Y��Ł�.�3�� /���?� �;�
��������;�2n�[n�;���HJ��6���L^YKJ<]�D^YKJ�O   �L�DKJ<]�D�DKJ�V   y Y�j!����Y�v!�����N�HJ�V  ے-^  	(i��?�2�   #Y-2   ��/v�OR�[nʢ���F��   �����Ct  �|�HJ�R-� M  ���
�<����v��GRm�A��١���3�
�dQ  �;A	.���
�<����E�3ٲ7C  �/��Ov�[n#[&�K�<��\R�HJ�\�Y�M��3� -�s    �����Y��~zH���x��Y.y�_&��Ѹ�z �V�[n�2u  ���S  �E�� �<R��P  �Y�3Ѳ�@  ��-�s    ���&ZE w�*mR�~z��<KU�U�1�M��H�nʚz��vB�q�"���vB��X�jOٿMa*mN� �V ђʶ.��	�8�A�;��8�;��8�;��8�;��;�
�Υ�����#�ѹ��y;�y�u��3�Y;���H"�#�����P��NQ�J���y���]�Q���J���t�Ѵ��j��rB�}�ѯ��]�чj�u�Y+���Z�i~��ф��q��oB�}�ѩj���y��'�B���}���I�����L��Pu�Y�]���j�u�Y#���Q�q5�����P��NQ�}���y;���j'�B�}4���cT��9��N��Vu�Y;�Ѷ¢]4�����j�u���Y3���FI8y�����F��XQ�J���y���]4�u�ѧJ'���DH�8�ф��h��tB�}�ѩj���y��'�B���}���I�����C��]u�Y�]���j�u�Y#���Q�������]��EQ�J���ѡ��]�]�Q�J������ѧ��q��oB���Y�]���j���u��3�Y;���H������_��CQ�J���y���]�Q�J���tkK�"Ѵ��g��yB���Y���j���]�u�Y3���F�ѧ����]��EQ�J��v£�R�R]4�]�ѧB��4�}���M�
#���U��Ku�Y���j����4�]4�u�ѧJ'���FhR�Iц��h��tB��R}�y�j�u��#�Y;���J8[W�����R��LQ���j�}��;AѼj������;AQ�J���	�>�ѿ��i��wB���Y;���j�]�Q�J���tZ oѴ��l��pB���}��3�y3���j���u�Y+���^�����ѱ��j��rB���Y���]�y�B��4�}���M#Yu� ��A��_u�ѭJ��4���y���j�u�Y+���Y	jX����^��@Q�}���y;�фj�u�Y;���Jۘ�����[��GQ��'�J���y#���j�u�ѤJ'���G����ч��j��rB���Y���]�y�B���}��4���Q���_��A��_u�Ѧ��}�y�¢]�Q�J���d�]I�ф��i��wB���}�ѡj���]�Q�J���n�W��Ѯ��l��pB���Y�����y�j�u��#�Y;���J�j����]��EQ�}��#���]�y#�Q�J���L���ѿ��e��{B���Y;��;�y3�Ѽ����]�u��3�Y;�j���]�굂��M��Su�Y�¢]4�u�Y3���C�|&=����[��GQ�}���£]�y�B��4�}���M�p���N��Vu�цJ�M�i�J'���Ec��х��b��zB���Y�z�M�Y#���Qۈ8�����\��BQ�J���i�z�}���[\(���J��Ju�ѵJ�M��;�ѿz�}���Xrq����M��Su�Y;�i�J���q���ѱ��b��zB��4���Y�z�M�Y+���Z�����\��BQ�J����+Ai�z�}���E�¡��J��Ju�Y�x'v�vz�}���B�����M��Su��#AY�z�}���C�7�V��F��^u�ѡJ�M�i�J���d�}ߣѤ��k��uB�}�ѭz�M�Y+���^�N������Y��YQ��vJ�O4R�RM�Y+���Y_c�^����^��@Q��vJ�M�Y+���Xc�������U��MQ�}�i�z�}���I�Ё���O��Qu�Y�M�i�J���a�&�Vх��n��nB���Y�z�M�Y#���Q?(�����^��@Q�}���B���M�Y#���P\`�����S��OQ�}���B���M�Y3�����tޥT
Ѵ��h��tB�}�Q���z�}�p��0k��y�y�����<���K��Uu�	}���,Ѱ����  �%,0x�/����<��<��<�.�<  ۖr�0t�/����<��<��<�.�  4���0q�/����<��<��<�.�p  ����<�����������
�D[  217�#\�<�����������
��   2��v�#P�<�����������
��   2j
[�#U�<�����������
��   2�XR0���;�Ѱ�/��/��/���   !�~�O���;�Ѱ�/��/��/��   !o�s�C���;�Ѱ�/��/��/��$   !ᬞpF���;�Ѱ�/��/��/��B   !˭ϱ)�/����<��<��<�.�E   ��!H2��H.��H*��H&��^ ђ�j�v��uV(#zMJ}B}zA�nьbb���F��Q�J/r�j �b ��0># �^�O��HJ.�����/ �<: ٺE�8[]=�
�◑�*���ѝ8,*{J����&ZE t�*m^�~vٰ��<Hq��K���X��A�n�K��J�[�X��Q�.KپMٿM�jOa*mJ��E +¶��r-я0v���$:
�֥���y#b��Y��e'r�J0q�2nRXn��   �;�0vѰ�%   �Y
��.�)����#A�] i��]KJ�4���M����<���:|���/l��!eKJ.�s��'�^uUq��.>]A|Y�{!
eKJ��.�R����V��.��Х���J'5�!��^ ђ���4V���ѿ��}�V�ʺA��}r��J�80>%��cH6b�E�(<�:y^�<R.��ʶ���V�^��
�:����#Eٽva�:B�R���:Q�.�Z����V>ʙ>��M��z�?r �3E�+Aq�J�)�NM.��ʶ���V!#�R ��[ŋY�[��Y�[ɋY��#�.-�    �:mV�    �6ZE�mV.���l��HJ���������������֕[n�!"��������� �Y�����������HJ����������Δ[n�"���������A�Y�E���������:�HJ�b���������3�������Ɨ[n�H"�������������������.����B�HJ���������������������
����1�Y������������������3������⦖[n��%�����������������ț6O  ������9�Y����������������p����ѺY�������������������%���k������%���G������A%���S������$���_�������$���k������$���w������A$���������^�[n�]%�����3���-���"�HJ��Z�������������������5��Ɖ�Y���������������������>��▨[n��$�����������������3���������}���Y�Y������������HJ�2Z���������3�ٿ]�{A�����[n�$�������������HJ�Z���������f�[n�a$���������������\������ڄ���@������*����������9�Y�y�����Ě����������Ď����������ľ����������Y�Y���������񺀶����満����Y�������ƞ����Y���������f9��➭[n��'�����3��e*���R�HJ�6�������:����y�Y������ʗ[����&�[n�'�����3ѳ������HJ�
��                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �[ 1� ܖH �[ � ��H ��[ �� ��H ��[ M� L�H Z�[ w� �H �[ 9� $�H �[ � �H ��[ �� ��H ��[ O� @�H Z�[ y� �H 0�[ )� *�H ~�[ ð ̔H ܣ[ �� ��H ��[ �� ĎH �[ 3� 0�H $�[ � d�H J�[ a� L�H z�[ �� ��H ��[ � đH ��[ �� R�H \�[ {� �H *�[ +� ,�H ��[ ٷ ƓH Ƥ[ �� ��H  �[ E� x�H N�[ u� �H (�[ -� ؐH �[ � �H ��[ �� ��H v�[ k� `�H *�[ +� *�H ~�[ ǵ     ��[     ԒH �[     �H ƥ[     l�H     ]�      �[ �� �H j�[ ӱ ޕH �[ � |�H <�[ � �H ��[     wEvg4IfAIn3	fAv?   }L}YOkQ3'@h]SfDJe\F<
  dBd -	 q@dUSs
-	
:   qF~dB
A DFtc.   GTpSu_UsUQ)SLj d^@)TL8GfDF)TL8   JiYc_eR@:P! LjrSu_"CbHW:P!DJirAnD"CcR"E !\Pst jYP:V XBR
] J.j nPi\[)P XWs@Oh_H)U[bGJuUPoQQlFU   PiYEaUQ)U[b Tn^Gr]S)U[b FoCMnVEbBbHF   bDKbBG)U[b  iUWBB FU nBJtFU        ���	      �ACJi Wn] cQW SP  @c  kC  BFj SuU cT  XVe @kC bBM \V KpT     ����NtDBdYN)CJ` ?tfCD33rg4t  5h.   '#)$*9)2!t7+?K+?x5<.~},<"M#;"h+dZN&q -l -G�� Y��HJ�V[n    9$�           }   i_�P        	�Y>WHJcc[n4'5	'z199.&4   ����Y`Y@DHJ    ����    �r[n    'EHJ�r[n�����CHJ�t[n    ����Iw[n	dY    ����    �>HJ    �Y�>HJ����    �>HJ    �Y�>HJx  x [  J J\ OXnM;_{L_{|j     ^ab.]v mNy.N  izv    R!:):  *1"1RyA  N vAR  R A yA   r '  6 % W     V'/%s         �7[.   ځ�?I).;5,)&(8,;
<((:?=   ;;iL            ,qNyj   -<43&4*<?),>*!/8;3-(.   4(48,83((?9(3(#4<44<6?<=-,*1*.0&,:,9    Z  ('.$?^,(&(^  sC  1	^,(&(sC   	7^,(&(sC    :?I^,(&(sC  lN{bsCw^<4+6i.i3 .(63?^!?9Wt    HyhIDPSi4=z'5.2^:**?^/5i6>3i3 .(63;
 5DP    lN{lsCw^'5
i?&/!z9;,z&(^:. 5^ 4=3%3(.&4sC    ,jL|Wtdz<(i,;.(6^//*.&4^*;%Wt   lN{nsCw^'5
i?&/!z9;,z&(^5,"=u=? .^=;%?sC    ,jOpWtdz';%?^=5^&*'z&4&6i>?3,Wt    HykFDPSi/,",9
,>^!?9z;(;Wt    HykIDPSi/,",9
,>^$/=3
!((>^%5"z;(;Wt    HykHDPSi4=z'5.2^:**?^/5i.;?-z(.DP DP+4;7%z;5;;i.;7';
 5DP    lNycsCw^'5
i?&/!z9;,z&(^,4 ('7'.sC ,jNqWtdz&.^,4<=i)(9i<;z;=$?=)sC   HyjLDPSi<&;
 4i* 4
i4=z&;,>sC    3 9&)/.^3<;iUbz,<4
 7i+(;#    CP  '.$?^(&(_CP.;5;;sz   Pgt u*&=(7^';,z'1&-w              ������HJ��[n?
;==3,
9/  9,.?*.??) 4&- ?:;,1 <);iLg>%  ������HJ��[n�����HJ+�[nxy/0  Oj0   k]I:   xy-0  ������Y��HJ����U�Yz�HJ6s7s) >->Ri3^->Ri#0# uf#  .    *?+?    ??+?    =5,( ?=?+?   /<)
  4<6    '?    * 6   3((!   +(((    '/;# ? ? 1*. ? . 4<6 / 0 ?9( ; + 4(4 ;
<((#    (-;  *!/:>0    ),>,)(#   *<?-; '>0  /-;  -(. ( < ),> / ' -<4 �Y��HJ�� n"�Y)
;3.z
&5^%5. ��[n�� Y�� J�� ny�Y�� J�� n�� Y3?; >^:. 4i*:3
 5 w�HJ�CXn        ����        ��[n            H   ��HJ            �CXn��Y    �MXn        ����        n�[n            H   r�HJ            �MXny�Y    fOXnH       ����        �SXnK       ����        �[n�YJ�HJ            }   ��Y            �dKJ�[n    �HJn�[n                X   ��[n            Q\|Y��HJ    q\|YX       ����        ��Y�HJn�[n            J   J�HJ            FOXni�Y       �^|Y    ����    ^           [   �MXn    ����    M           K   2�HJ6�[n                ҢHJ^L�gK   ��HJ   ��Y            ����    ����            [      ��Y                }P ni_�PX   ^�[nH   j�HJ            ����    ����               H   �HJ                �G Yz{�C|   1�Y[   ��[n            ����    ����            H   [   ޔ[n                a J^L�gK   ��HJ   ��Y            ����    ����            [      ��Y                &n ni_�PX   V�[nH   b�HJ            ����    ����               H   
�HJ                7t Yz{�C|   ɄY[   �[n            ����    ����            H   [   ֗[n                UG J^L�gJ   ��HJ   ��Y            ����.�[n                [      K   [   v�[n                b3 J^L�gJ   b�HJ   �Y            �����[n                [      K   [   �[n                �- J^L�gJ   ¡HJ   ��Y            �����[n                [      K   [   ��[n                �' J^L�gJ   ��HJ   Y�Y            ����΍[n                [      K   [   V�[n                _# J    �^|Y    ����    V   �`[n    [   F�[n    ]THJ    �Yz{�C   ٺY                    ������HJ^L�gH   �HJ                    ������[n    BxKJ    ����    b   y� Y        q\|Y    ����    F   �� n    Y   ��[n��Yb�HJ    	� Y     �[ni_�P]   >�[n                    ����Y�Y    b�[n    r�HJ    }�Y    >�[n    �HJ    �Yz{�C   ѻY                    ����*�HJ|   ��Yb�HJ        � J    �Yz{�C   ��Y                    ����ʻHJ^L�gH   R�HJ                    ����Ό[ni_�PX   N�[n                    ������Y    ��[ni_�PX   �[nH   *�HJ            ����    ����               H   ҜHJ                �� Yz{�C   �Y                    ���� �HJ^L�gK   ��HJ   ��Y            ����    ����            [      A�Y                �� ni_�PX   F�[nH   �HJ            ����    ����               H   :�HJ                � Yz{�Cy   ٹYX   ��[n            ����    ����    ����    K   �HJ}   �Y^   &�[n����            [      ��YX   {   O   [    �[n            � Y            �wHJ^L�gJ   j�HJ                    �����[n    &�HJ   ��Yz{�C|   !�Y                    ������HJ������Y    �SXn    ����    U   ��HJ    J   "�HJ��[nq�Y    P�[n    HJ^L�gH   ��HJ                    ����[ni_�P[    �[n                    ������Yz{�C   a�Y                    ������HJ^L�gH   
�HJ                    ������[ni_�PY   �[nH   ʛHJ            ����        r�[n����        H   X      �Y                x�[ni_�P[   ��[n                    ����i�YژH         \�H  �[ a�         c� �H ^�[         6�[ � j�H         6�H Θ[ A�         ׶ үH j�[         ��[ ݋  �H         ��H ��[                     �[ 1� ܖH �[ � ��H ��[ �� ��H ��[ M� L�H Z�[ w� �H �[ 9� $�H �[ � �H ��[ �� ��H ��[ O� @�H Z�[ y� �H 0�[ )� *�H ~�[ ð ̔H ܣ[ �� ��H ��[ �� ĎH �[ 3� 0�H $�[ � d�H J�[ a� L�H z�[ �� ��H ��[ � đH ��[ �� R�H \�[ {� �H *�[ +� ,�H ��[ ٷ ƓH Ƥ[ �� ��H  �[ E� x�H N�[ u� �H (�[ -� ؐH �[ � �H ��[ �� ��H v�[ k� `�H *�[ +� *�H ~�[ ǵ     ��[     ԒH �[     �H ƥ[     l�H     ]�      �[ �� �H j�[ ӱ ޕH �[ � |�H <�[ � �H ��[     e 
((./
,"?  �H,43<.1  A 
6:?6(4%? m[9,.3&>%?8 6;,  k 
((.,'.?  dH=:.;;(;  bX,,)=,4
  K	=,4
  � <)3,/<;)  �|(=?8 6 0|?
3,
 4
,(  n 
((.3, �X)(3
5/=3%?1+0*.  sH=%??=. 8=?  [[9,.8 63, �H,4.;5,)  ?,.3, [9,.-0)
,7: (*.;#? |?,;,=?  fK(>8 6  �K .8&(- 4%?1+0*. eX,,)$?*!((>   
((.2,;  �K;7';
,;?- ~  .*!((>  �|?$3(.(*?:  �X) 4;1? r 
50%?? ??
?9
=2?  � ,?2 8(( d?
(*-(:)  �5-+(;#?  �H??8 6"? �5,%?? �|%)
;9=  R}%)
;6'  9?
?9%?0(7  4[9,.) 4&-3,9
&(  [9,.-!5=
=20(7 
H=;)&4  2|?
3,
=(+/
,)?  50M{t%6  �5=;?-:).??  +,zhP-6  
 	,6"*/
, -2iLg>% ( =?'?

6:?6(4%?  7'.;4=
=?9.=&4,9
   =?'?
?
*
 5   7'.;4='4*.?   =?'?
*' I 6=.?-8/:.?  ? 
=*?->,,+,)
?-?:   .
9,4,,+,)
  > 7'.;4=(>8 6  9 
=*/<?0/5?  � =?'?
?
.=/
;%8*1 1 7'.;4=(>8 6"?  I4
,(,.=;;"% 0I;t%6 E 9,.3&>%?<();,  _ 4$
&9:): ..It: �[+<35-=('=? �/-,;
,  
=Jg>%  � 0,. 5 ;.IiLg>%  fX,=6+'-'> BX,(3,*?=3'  9[9,.* 75,/5$;
 5  #H=	:.$$? R[9,.2&9%$?  � ?

5$;-'?? ' "=
&9:) � 9,.=<(,4
(*?: �H(*,,%5 �?9%5 �?9	3?  �I4=3%3, .*;?=3' + %?
, .*;?=3'  =?
(=3(6-,9
 5  �H(,
(=3(6-,9
 5  �H(*8;?  � =;('.*!((>7-  �X*%)-,.((6, �K:%5  �K:,? 8X-,.2()
(&(  �|6?
;<? �X-,.+'2'>,>;199.&48 6
,( o[9,.3&>%?6(4%??  �K-?=!;53<6
 =? $X-,.6(4%?=&/=  [9,.-=>6(4%?  O?
3,9? [9,.-=;=/I4& � 8;?4 ('7'.-=('= � ,?;',;5$?=	
;3.)) \?
4 ('7'.-=('= R?
4 ('7'.-=('=  �[6,;?=(0 �H(*=;?=?  �|3=/%,? �X( (
<;6&9  �I)<(>);3
,

; �H;?-

;  �[7:--?.=(  �I4
,(&9,>:,9,7'.  �I4
,(&9,>7'9,7'.  �/=3<0.5) >
2; -H=	
;3.9??  (H=	
;3.9?)  � =.I4& � ==  x[9,.1=  5X-,.-=>6(4%?  �3(*-=('=?  �H=;. 4  h =&7((. 4  k =&7((. 4  +X-,.;',;5$?=;3+6                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                             yH Y*l J�] ni4 Y�`HJh�[n        V[n��Y6�HJ;[n        W�[n        ([n    A�$d*,>@�1����A�68Aߖ�@�M+��'�jb��
�����Y���G�p��q���:�h���dpd���̋K(rz��6TƬ
�>��j�J������-3RV$�+?I->�����utR�.~H��9�W*�yH����������l�=&���P]p&�0ޅV���At�)^��ދ=��䉰��Iƞ�X
'eD�_�p3R�����)�=h�R >kEo�ڣ	���)Vw>��B��ӗ�QB��L^j~�Th[�3C̩�wqN�	�v���Ҏ�>X�W��m���U��k�7� \;#0[�^��҆���"���M�v��H��������(G״�� �EMW��_a@¯�JC��C7�QF�}���０W��s�f���X�Y�>ᾶ����m9g%�6�S��?�tQkC��棲�����Q��s����s�&��>u�Qc�2��V.g{�Q,�H�G����E���k��}��{�8eŹ���ah-�g@�V�5��G�T�9�g����������>�.�.c��r�M�'"���;G{M�kh���_� Ë�]_����k)->nLΝ�>16��7k��e��s����X1R���t~w�T�x�EG�H��b�Т���n<D!��W��nׅ�шw��j��0�*K�;��T���1L�È�w~^��,gr�6� f�����%@�F��uX2F��mG�9�Z�I�����/>7e�z�l�O��'������M��MWh\�����.-�
\�����Z2p�hZ�J��;d:j�1�1�T�umvx
��H��=4�����+�r{N9�r���B������ŝ
;�����5�j��H>,�m���~,	kU% ��k3岢�����L���b!��,)}N#6<��=�2��%��yz.k�g_�OT�޺��|�K~G��1��h"��P�jv��Tjْͫ�yL:О�)����9��x��x�&�ܖa^���p��@n���e䞅�Y�򑭍�
�1���%v�����l̠�t����ѐ�����ԣ4�}��f���f2QS��q}�k:4SE�	9</�g>	�8�S9���n��HJ    g
?    ��[n    t.    *uOgj    iwQs    C   C      ��[n    tA199.&4>	                 K                   }                   ^                   L                   x                   ]                   A                   w                   P                   B                   r                   W                   G                   q   H       ��[n    tA&=*;(;=>>	   ��HJ    ge?5=/(4,=>>	   4(6-z,9
&(Bd^:/:9 *
 p   �H  �^  �t  f\  �t  5,4    ," .9 7'.;4=='4*.-	
(."?    -'3,.P-6 �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                               [:g[:     %;?(7    )I7*g0I ~>3 '/ $0 ��[n    tA
0*3/5>	 ^L�g            �Y            /�  �  �rY�VHJ�a[n            2kY    �jXn                            �]KJ            nmXn            �y|Y                                                                                                                                    �>HJ            ����YF�HJr�[nV|YrKJ  z i ^ z i ^ z i ^ r a V r a ^ z i ^ z i ^ z i ^ z i ^ z i ^ z i 6 J Y n J Y n J Y n J Y n J Y n � � � � � � � � � � Y n J Y n J Y � � � � � �  [ H  [ H  [ H  [ H  [ H  [ H  [ Y n J Y n J � � � � � � K | X K | X K | X K | X K | X K | X K | J Y n J i                                                                                                                                                                                                                                                                      g   [           zwdW#          p�[nG�YT�HJp�[nG�YT�HJ        �     ����
-                                                             .                                                             �T|Y�pKJ    ����            ����            ���� P                              n   K   B�HJv   ��YS   ��[nC   ƩHJn   9�YK   >�[n[   F�HJm   ��YB   Ɵ[nP   ʨHJd   �YA   ^�[nU   ��HJ   ��Y#   ��[n3   ��HJ�   ��Y�   ʜ[n�Y              _  �u       G  �z       �  �z       �  �v       �  �v       �  �v       �  �v       �  �v       �  �v       �  �v       Y   y   1   P   `Xn    :WKJH           Y                  X                              K   X                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                       ����W   a   $   1   �   �   �   �   oH  y[    H  ����D   D      -   �   �   �   �   Y[  u  3H  %[   z  ���|   Q   >   �Y  �   ����Q   R   ^   6   [|MR    �Y  :�0�_       ��      ��      �ֺ�    ~ɦ    �Y  �ݓ�^                       ��      �      �Y  �ݓ�^                       ��      �      �Y  �ܭ�d �ܡ�%                 ��      ~�    _  ��^ �#�L                 ������  k~Ȥ    H   L   |   K   Y   |   M   B   {   D   \   w   N   V   v   E   S   r   C   ]   u   A   V   h   D   L   q   K   J   s   X   H   l   K   {   s   |   X   ?   D      |      K   ,   D   	   s      L   '   B   6   s   $   z      U   (   w   O   L   �   C   �   t   �   S   �   _   �   s   �   s   �   D   �   |   �   Q   �   D   �   o   �   X   �   B   By  r   
                                                                                                                                                                                                                                                                                     biKJ    !�Y>�HJ�[n�Y�HJ*�[n�Y�HJ>�[nq�Yv�HJ^�[nQ�YV�HJv�[nM�Y �HJ��[n��Y��HJ��[n��Y��HJ��[n��Y��HJ��[n��Y��HJƐ[n��Y�HJ֐[n�YΧHJ�[nɃY.�HJ�[n%�Y>�HJ.�[n�Y    P       �iKJ�oXn�||Y�XKJ�oXn�||Y�XKJ�oXn�||Y�XKJ6%6%6�iKJ                     �K         �L         �A        �E        
�F        ~�[       ���_       i��P     ^��A�}   ߤ��R��^���9q��� ��[�@�C��ߍ�
T{�s�����:��l�����u�؆�7V"�����ڷ�����1+nc�*�5Ԡ�ǅ�$�߯,���Wf��oVYMԱ�n�������� ����G���C��s,Mr<��<,�&���cE|�̤	3�#t�#r���Z����z���~;���$[Ӈ�=�ܢ�n�܁��42���i�|:�l/    �����������A8gt��tP��A>E���4lʯA��R,C�Mɘ�A�U]�e���A	�� 6�L�IϱAzg� ������A����;�X-��Af%����믓A۞-r/:�N���A�=��c;�Dφ�Amy����rk� A('�$�&l�A��Q�\���k�Ame۠c�n��pA4�߭�5��@*!x�y*>ف��CؠDP lO��Bhӯq�9�� ��E��&AAϡ���YE��;]��/I�tDz+b�y�{�7�ZG����������L�2�X�,�'�JRl�dlJ	Ї1[�z횠�'���`׽��u�.�xf+����x�'o�w�֔��^��t    ��HJ    ge?6'=
!;(;=>>	  �                                                                 Nl" yj                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                       n  �   j�y�N�k?{L(h�{�L�hYz�M�i�zjJ�n�}�Jo�|cH�l��H*m�~�I�m2q�F�b�q�F�bZpG�c�p-D�`;r�E�aDuB�f�uTCUg_tC#gt�C�g(w�@�dsvBATe$v�A   i  5   'N�jMx�O�k�{FM&i�z�M�il}J�n�}�J�n<|�K�obnH�l��Hym@~I5m�~F�b�p,D�`JrcEar�ETfUujBf�u�B1g�t�CLd2w@.dw�@?e�v   j     (yO�k�xSLGh8{�L�h�{�L�i�z�Mjn�}�J#o�|�Kbm~6I4m�~�I�m�q�FTcKp*GL`*s�E�a�u�Bge   >  6   �n�CI�mxq�F�b�q�FXcQp=G�cas�D�`�s/E3a�r�B�ft\@�d�w~A`e-v�A�e�v .     �jax�O[hi{�L�hZzsM�i�}K�o�|�KGl��HYm�~FF�b{p2G$c�p�G�c�soEsar!E\fdu�B�fxtDC(dw�@Qe�v   :   kHz-M'n�|EH)l��H?m�~�Ifb p�GK`Cs	D `�s�D�a=t�CkdNw@d�v   *  
   �z�M�i�z^JXnf}fJ
n�}�J�n�}�J�nz|QKyoI|,K4o�|�K�o�|�K�onMHll;�ERfxt�A   �  U   "O�h�zJ�`qr�B�fw�@ �  2   wyuNh{�M]n�}�I�m�~YFNbuqUFZbiqAFVb]q}FbbMq F�bqppGc�p�G�c�p�GV`�s�D�`xrqEa�r�EPf�u�B�f�u{C   �  a   �M6nMqF�b�q�F�b pGA`7s�D/f�u�A �  F   iyN�j�x�J`o>|�IfJt �  :   �i$|�Khl�Hvmp�Gf`�s�Dka�rxB)f�u�@�d�wBAkeMvAev�A�e�v�A �  v   Ey N�j�xYLCh�{�L�o�~I�m�~�Ib3q G   �     N�j�yO�k�xNLrh{�Lki�zgI�m�~dF>b�q�FccDp�G�cr�B�f�uCg�t@�d_v�A�e   �  *   (k8|�K�lq~LI7m�~�I�m�~�Izb>q�F�b�qkG�c�p�G�c0s&D�`�s}Ear�EQfcu9B�f�u+CRd�v  H &   }h,{�M�iQ}Jn�}TKo�H�lD~I�m�~�IAbkqF�c+s�D�`�r�E�azuXCg!t6C[d�w�@�dv�A�e Y[    _N�h�{aMPn}�J^o�|�H|a�r3B�f�u�@�d�w�@�d�wOAbeOvlAe0v$A�e�v�A�e i[ �   `N�jJx9O�hgz�M�i�z�M�i.}1J�n�}VF_b_qtFrb6qFbq�F�b�q�F�b�q[GNcupKG\cepEGmc!p�G�cssD�`�s�D�`�s�D�`�sAE|aBrEa6rEa*rE�a�r�E�a�r@Blf>uBf.uB8f�u�B�f�u�B�f�u�B�f�u`C	g:tCg�t�C�gXwv@�e�v�A�e�v�A�e�v NH �   Bjny@N}j<yNj�y�NHkbxqOk1xZOkx4O�k�x�O�k�x�O�k�x[LOhl{ML}hD{�LTi]z*M?i�z�M�i�ztJ!n}"J7n�}�J�n�}�J�n�}�J�n�}�J�n�}[K]ob|K-o
| K�o�|�G�c�s�DjfVu�C�g�w�@�d�w�@_e\vrA|e;vAev-A�e�v�A�e 	[ 9   ~Nuj<yNj�y�N�j]xcOk2xOk x�O�ki{~L�h�{�LUn�}�Knl6H�l�p�G�c�p�G�c�p�G�`�sgBf�u�B�d�wXAWeUveA�e�v   
 �   @y>N=k�{�L&i�z�M�i�}�J�n�}�Kzl.2I�m�~�I^b^qaFb*qF-b�q�F�b�q|Gh`SsE�g�t�C�g�t�C�gvwT@Ud\wv@}dDw@d(w8@#dw"@�d�w�@�d�w�@�d�w�@�dxv{Ate'v9A�e�v�A�e�v H JH  JjsyBNkjNy7N�j�y�N�j�y�N�j�y�N�j�y�N�jyxKOPk_xsOzkBxOkx�O�k�xSL~h<{�L�h�{�L�h�{�L�hszDMbi@zMi�z�M�i�}�J�n�}�J�nt|fKo|&K�o�|�K@lqFHtl+H�l��HLmo~AIfmC~Im+~�I�m�~Fnc>p/G4c�p�G�c�pD`�s�D�`�s�D�`�s�D�`\rtEqa>rEa(r?E>a�r�E�a�r�E�aruB+f�u�B�f�u�B�f�u_CBgltACkgTtjCrg=t�A�e�v�A�e�v�A�e�v   * �   yy@NljUyjNj=y:N/jy-N�j�y�N�j�y�O=iz�M�i�z�M�i�z�M�i�z�M�i�zKJknV}aJ�nq�F�b�q�F�b�q�F�bkpFGicZprGecNpnGqc�p�G�c�p�G�c{szDn`RsjD}`/s!D�`�s�D�`�s�D�`�s�DSa^r~EaaRr�E�a�r�B�f�uQCgt�C�gqwq@wd�wA�e�v�A   �[ �   LNjy�N�j�y�N�j�y�N�j�y_OhkNxOkx�O�k�x�O�k�x�O�k�xL$h{�L�i�z�M�i�z�M�i }KJmnB}J�n�}�J�n�}�J/o�|�K�o�|�K�o�|0H�lY~nI-cp�G�c�p�GE``skD$` wL@   �[ Q[  CNkjQyN�j�y�N�j�yYOFk?x	O+k�x�O�k�x�O�k�x�O�k�x\LGhg{Lh#{2L;h{�L�h�{�L�h�{�L�hz(M�i�z�M�i�z�MKnl}iJvn/}J'n}�J�n�}�J�n�}�J�n�}�J�n�}_Ko1|Ko|3K�o�|HH^lJ`H�l��HXm"~1I�m�~�I�mVquFbq�F�b�q�F�b�q�F�bzp�G�c�pzD{`(s3D�`�sjEsa uPB�f�u�B�f�u�B�f�u�BPgHtC'g�t�CFd	w�@ � �   �y�Nk�x�O�k{{wLh�{�L1i�z�M�i`|xKooT|tK{oH|`Kwo<|Ko�|LHnl:�IMbXqoF[c\pGc�u�B�ftzCbgHtCg-t;C�g�t�CKd�w�@e'v�A�e�v�A�e�v �H    Djdy�N�j�ycOIk�x�Oh"{"L�hXzvMsi�z�M]nd}rJ�n�}�J8o�|�K�o�|�KNlduHl~�H�l�^IEmf~{IdmH~Im$~�I�m�~QFYbVqmFb   �H &   �k{�L�h�{�L�i�z�M�i�z[JXn_}kJn$} J�n�}�J�n|#K�o�|�K�os{Hxl�H�l��H�l~OI`m �[  [  �L�h�z�M�if}FJinB}Jn&}J-n}.J1n�}�J�n�}�J�n�q�F�b pRGEcJpbG	c:p6D9`
s"D�`�s�D�`�s�D�`�s�D�`�s�DMavrJEaaBrEa&r*E�a�r�E�a�r�E�a�r�E�a�r�EYfjuBBefBuBfu�B�f�u�B�f�u�BAgntCgt2C�g�t�C�g�t^@Ydfw@dw*@�d�w�@�d�w A]e^vrAuev.A�e�v�A�e�v�A�e�v   � �   ^ynNuj.yN-jy"N�j�y�N�j�y�N�jzxROEkjxFOak:xOk"x>O%k
x�O�k�x�O�k�x�O�k�xVLQhJ{fLh.{�L�h�{�L�h�{ M]i^zrMiz"M�i�z�M�i�z�M�ir}BJ}nB}Jn}.J5n�}�J�n�}�J�n�}�J�nz|JKeoF|K)o|�K�o�|�K�o    K �   MjvyVNYjjyBNmjVyvNyjByN�n�}�JQlF�DiaFrfE	a.rE1a�r�EifJubBuf>uB9d
w"@5d�w�@Ue^v.A5e�v�A�e�v�A�e�v�A�e�v�A�e�v�A�e�v   J| &   �y�NymF~fI	m:~Im.~Im"~:I-m~6I9m
~"I5m�~�I�m�~�I�m�~�I�m�~�I�m�~�I�m�~�I�m�~�I�m�~�I�m�~�I�m�~�I bzqRFEbnqNFib�s                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                