MZ�       ��  �       @                                   �   � �	�!�L�!This program cannot be run in DOS mode.
$       ᱇����ӥ��ӥ������Ӧ���&��ӿ���M������ӥ��Ӽ��ӥ���5������Ӷ���M�������Rich����                PE  L             �    P  �      �P     `   @                     ��                                       P <                                                                                                                @  PEPACK!! P     �                 @  �PEPACK!! P   `     �              @  �PEPACK!! �   �     �              @  �PEPACK!!�H   P  J   �              @  �                                                                                                                                                                                                                                                                                                                                                                                                        ��K��ӣ厘j����0�T/<�
֚��N�v��)�M¹W��fD�y�q�\S��ZX�m[��Z����pM�^��P���;S�'�"�xU�!��G=�WԂ<��`NZ�?��X�̑ܻp�� Z}I+�n$ ���U���������2��uzA!��*%m�$�v��+c�u��ۣ�q��Y��c�[�� g���̧��' ��35QewAٙ�p(�}1n�ɻ�����꽁�c
߉G�s�ϛ�1Bg�{�z>=#���Q@ ��v�@��u;�⺑e8z��zǮ*��g��80~�a��R�X�$�:��m���t�:��>PG���2�3b����{v��aˊ"�R�a���g������V2�`��d����#��d�o^z$P���,���n��y���h��VlG�	�Td�~y������X���*�I.p$p���x�i�{��no��|86��j�Ӂ&;J�R�_�TshG�����(Y�-�cb볮�|e�҃�T�ͤ/�Q.3a�g�TXQ��(>�������t!��M�|/�27H�_�~-S ����Ք��#����R����]���ka��&�@e�j(�ҩk��=WlNDQ^v?��	��&�ʇ �{��]i:OV���m=� �>��
�Oϯ� �o��A�����{5I,�B��*خ�5Z����}ч@_�:�d��$b�PZ�=8�f<��s$d��$��:I��XvV�~%���ࢗ��7C l�=u���U�08i{��۝v\� ���q������)�!���o�- ����yj21�	^ա�.��VT�=��NX7G:Bit̳g��V�����������0͏Ә6v�s
k�66Ҟ�����&�[��$V �M�_���K'�C%�%kU*T��d��~~#� k�XT����,.�,˥��e	�Ý ����~�\�߬�n�.>���'����_S�UCo��,'��z�$����F��T(�k���onW*�|�2�f��t�Gk�>&hFc�"��3�m#���*D���f�yj]�ӼELWQ��$ji�/ldʛ���D��AW��/i�s�=��&G?��`$y�Չ���4��Wύ��z�$;h�U�Y�E�%?��� ����9�N�@�o �����q��������V[A�j����.�<���#~4�$�o1f����v���n�tm�O�M2X�b����ڡ�c���'�	a���}��?�=u�/v��<�f��E��P���L�Ϣ��R#�U۽���g�r�*��#�X��`{On�
�"ͳ�:�e|G���7�ځ[�0G���8�R����|CY�㣚��-���IsPF��.�I��7`/A�EJ��E�f�DX�H�6SrV�>☯ �W�g�V��0p��r?|�;�/����0�4ż�~���a*��;/2~W� u*_�ݟ@I�eZ�{����۩�Fl��Cx�\�i�~^n�l�ǔ�i{'�e�X5�x�����D��Л��}7�:!0���R���ɓK�4)�d���i��8���&P7�9�q;�w��gX���M{2�йr�5#�Hw�٭p<۹
�5l��=#�jb k$ٶy���ZlI�s �T0���f@��8(= �u�LqG~ K�&#;�Klx5�tO��A��&H�e[!h	�����z��~�gfh�x�
ca��gYKAJj�Δ/rM�%�2_��{-MT�֫.�$������͐��3�&���2����wK/�>i�k���<7�f���C%����t�yu/l��G}��*4���-�`�Ws�[�-p��v0��[cN),��P��9w�>�qvAW�,[\Nó�t�����6r�v�0�=�Qy��L��죊�c�r�N<�_"��"�Z��b�����Dn�b�r�EaD��G3�a.���������UZ��ϰ�T�"z��p\�]Kfioe(��h���{����6o����Z2��AY���k����m??�@/5�N���B�DV(���0�)΁L{�J�M~"�$���?n
��,a�� ,����m���aJ�N�&�1n���8���p� ���!"x9]�R��f���.s����:KRui�?j��b�P��˃�2��4�rk��	�t��Da�i�c9
ͭ]Q/�Ь&������v��b7���9��R��^�<�7.��{�(8���Z.E�
�3���$��1�������l��Ա|�4w[
ah�9jq�L;��L��	}���u�����PH#��θa��kpe$7�}l�I|o���W/����I�@d���P+��>k͙ 7�*i?c<U�Yh���U�b%�cru�8�X��&?F����v�e�bn��I��6���#<�A~�,���b��J�'�N6�&~��"�Q�5E���
Q�5\�o����d�
s��{�C� lE'V�v�@9����:�0��j|/A~�����X�B���F�:(��膞.:����v�c�5�ٲ�R�@�.��&]�N�]�����K�~�'����H��ڿ�A��l$ b���2j�v�~K���^Ώg76+y��R ?��u3��?|���zړ��ή�S��
����gA;�\�a�����K(K�ڲ􌰾 &�s��Vk�N. �L��A0gyT���m%N���͟���F���f}#-a�����"�/h{�4���E�m)��w(��E�)"Zs3���s@��l'�?D<T�mC�X%n��b^�*u�g҈-�����j ��z� ���W8��,��_�@�����ҍˑ%v�{Z���Rd|���/C2�%��p.�^Ng�xH�3fI?}��Az���1��0.&�͇`}����J\��IlD{����~��(o�?�|�r}.��cr܅�M�1ȅ�AU�̖�@�
0!t���G'7�ŗ�	��\�=�M����e�[��z��"h;�F�� ��)}"{V�����9#���|j�̖�L}}��ihoh-�����kE�`
?���D1�������������M5�_ta$�Zi}#�j�A�(t��mQ	��9�A�&��rZ�����V6�opG�/2Z�m�3���2�	Xv��nE�$��9��׹X���cԛ���JW��g_��) ��&h���N��5�w�2��� ��&sm��bl�aYT\���X��qa\U�3qB'8%�C�V����b�o
h-�!�HpV�'��M������}��m)��' �� ��%4ri����t�Z���AE����\kR��){���0�ǟ5�9sI�$a2^�l�E�'�TQ�~hu}����[�#�z7{��8��t�����S[^���P�TS�Y�M\�n�o��|x�����(sv"���s��;�ݞ[���N^�v�0(�_�kq�뙻@u�Z�n0�����
$��9hb��x;���%����lz�Hr2��T�hb�r�ū�8�v� #x����u4[����{���$<jZi�RUa *�)>���21}�It���A(=�������r�:��+/�S_�@��+ح���;<��d��8/�[V��ʕοcڠ�y��\Ey$��I��f�����e?O}FM���]v�0�aA	Ѻ��E&���6��� �u�؈��1�����J,ɑ��=g@X�l���߽���lzZ���(z���0v�t��eH�^(h��\���٭#��yrǋx]N��~���Vʠ&�H���
��GJ� #��Ne������� �{����օp}���@2S��@7ҩ�q���BeI:.S��u����	�;�ʅd�\�=��0\❕�;��3��@�S���A�ڳ�่����[?'��TgK�2I�ަ�W|'d�H���  ��b�����@j���$�(�m�Ҡ'�Rb�,>�P�w�I5��F%��e!V�-��6H�?��Ҹ����H�����)JF��*?��l�L�Z��3��?�P����Tz@?S�����J ON�z	A\�}o1t`���eֹF0攨"��o6�-�k���udh�AZ�mr!Q�-���-g1���y�I�,�$vѩ�I{<n���Z�|�(d���J-�Y/����?0%��M�H�R ӭ�j*�{��-�a������
�Yu���|���/z�
݃n�T>��k~����י��p,/��<�����?�7�0�	Q��2�ܕk=2���1�o=�8�Q^F/x� -��<���&c�"�0���/����	�>6���7����XZ��Q��@2^���i��UŹH���?�[5l:�hC��&!��w�� *A���יI�}E��� #�sVl�>��+��ŉ���vUA�\�	�ȭ�(�BA��L5;���7H/�x@�nǁc3�VW�;��9[�_#C�?�
����ɭ��?��߉`9��=���	L���,�I��d!��Np  I�|M�n�x>~sg�m����M$��0m2��r2$k8C+�C�������2�f���q���*���6<�L�&"��)��]%�h�k�A(=��R��w����-��"��L=N�Jv����V�;E�
KH)����-JE77�I�UU6��в�u��>���4�^B��B���!x����E�/ÖN�uy.E���#��t��&�Z����M�1�)�d�{k�B'rЌ.셫]��#�hSXL�A%��H�?c�<y^^�%���J���Y��fX�����א�*�m�����hRɠ���F��)euUfx��ov� �:�Xrm��r�4�"��_m�u�4Z+��B��OZ+��՗�_�$4H�?�Ц�w˖�@·�̀���fw���믃�Vy��IS#�r�v�V���sh������՘��ܩ���"T6w%d�+�L�_��_ᨡ��C�����b�Dl��mq|���Td��J�[��΃7���dy�pC(�V?@S������<)ͬ�Ly,O�3ZSw�`}m;.��������I����� �\|<��ɳL�~���JN�a�X|�%��t�!��b���yZ�O���Ӣdb�4�~��W\��u-ǖ�C������oGc��=��Ów�Eg�L�Kԅ���t�:����K|M�s9��e���<Ż4Dyb]�b��T~GG���Ʋg]�G��W�g�����ow;	�����ҕ�z`ȥ*��h랬�R���(<���zJv!}w8�Ⱥ]stK�*��S�5s0h
ƋM�^�^�##�&�í��e1���bpg,����O%Y_Jx�� R�3�rtY0��~��{��Mr���ٞ�x��Q��׻3G�Đ	4@w]\�ݪ'��v|*{��4X)yh��r s9���P}�2��}�~sv��R� mt��V��"����fl�-EX8�N����4�^��L�#l7СR�>c�c�b��e���C?on�z�>Bn��nj�C��C��ʭ*�����OB�F�s�\b��%)3Eږ2��lz��Ŝ.����o=j�O��(�<���5�d"���_S_ȟ�B(Z�
��/�>R�>���!��o��m"d������&dv%ӧOw�@!*B��o,G}Myt��H�n[���,et�,'v���%w��>u�N
\��s\�O�-�P���c&^+�����<d�vk���h��;ﵫ�D��-z�p�=��*4>-�(OԨ�ŋֳ��u�N��g�L	��Q5=��g]1�+��ؽV���%�n��K7W��P��2�u����a��u�&�:ZG�Ge�7��Zvq�4��M�_��[�=3��I�*Ф��K�{��|����]�������ѹ?�A��;�֜my���F37ᖓ̝��v�����������"�iֆ4q)Q��:����xe⓾���k탦�r�l�@j�;�M���ҟ<J�#�a:�	v��'�d�Id��g2g�'���"o�Rl����ˋ���+�{zW3;f�H�I`1� �f��g�2K���D��?1V�t�s(!c�	�].��̽칻�'��w1+"S@�s�>�L�t[�m���ռa�3^�@%�Κ��ǔ�������c������bzЅ}�%+�%�<�_����w�@P��:$�Y,s�w�Q9+��)u�*�Wi�>�0�N%>�BgF���o�6
��%]��k��dI3fk�y�j�#�~������#b"П*���{�8�����$�EROE�$�M(�Ś�n����܇��`e1�ho7ĕ�rMq�) J�z㷒BV�H(�}�t\�]r��9�%�hw�՜o+�4'���̚*2g����=�h.��&��������.�N[�`@O'h�,%8"X��/�6Ӊu����D�c���~ �B��i��,�Q'R!N#BG��SF��K�M���s��{̱�K jJ��o	i��.�ޑ@���Cw;88k>B��s0'�P�p��XN��i�ö�B�_��wH�l�@,%�B k1R,�&�N����H��K��o�B����駍H�Q�(3�+k�x@SF����z��.>��4� �:��.1�D�uB�֌���<� .��ǘS{��VKUЧ��'o��:_�hL�V��A�"Y/��/�h	�bS5�EN����&�%3�ԋ������p5�%r�7�6,�YiR'�dZ��R��ռ���<Ƃ�a�B��ct��&�Qz��;��9_q��ᬋ߿�*f�%�h~z��tA�&�%4Y�2�a΁7
�Qȏ����W��EsQ��:|_RdN��P�b~���r��
���a�>�iG.�xYĹ�%@��!��.y)����D�su�ޠ��1�G f�sݯ�M
� )���⑕�M[qh���l0�S
�m3w��)�i&K�h�BaF(С���*��D�I����e��*����O�}�q�Z��b*n�J)�H��ơ��N���������g��9�6�.�L�w�@���9`�?w)�z�Pa�ˤ����*�L�i��T@�H16����껋13��\�_��!���i��nG~S�T�Z�yzjc��	YD;�. hph����e;u�#�&��u�U:�>�*�=�S�EV� ���o;p[��ƾY�vM�M�p��pª9+q͠nZ��:�v�?��|����i����Xu�����+ހ���9����)��ct�8~L���߳r%gs0}�72���_M�a<2�Iǵ��G��=����%�?��#�S�@�eY�>w�._,?�V2��R��<�`CnEE�&����лx�~׋?��#庯<\�Þn��`�
�_��诶<A!)!9��]�
���P��0�e�Gq�3>>.1�F����1��w��D����㍃.�~�#"����P|�A��f�;��f��=뮃���ݾf�'�P�����B��MTn�=P^�e�/�Y�ϫT<��m3��c*�|����(O�oY8wӔ�SU�4�"��K(D匥,\����eA��9jfC����}f�9\`��Ct���˝p�d"�)E���հ����`{�m��v�~g��'w.y��{|�U���afT������(=N4���J�]��Γ��M4n
�x'��7�F�ĵ���S��^��p��E��\(;��k�4��N\�z6V��j$�
��S��F������!�˶��pi��u�M$)��>c�z�L����B6�v��%��$P�(4ܥ��\�3��Af4�e��+ɥe�C���J��<�Ƣ�� ���X+c̅fY��{`.]�b�}�eW�{�j�R�!�%f��.�l�K���4��0x��L��L�F��>c��W�H�DZu�ԈK�CIp������o���f�mUxgi�����R���ų�a1��e�S�7@�I�=�?�nXLa���JE�b�ۼU�A@?�R�_L�x��h��6����HK{gdw�Qt��VK�7���fz����T�,�S�ϥ�hT/�瓨�Z2���1���򜅹-�-��/N:�DIέC�(��&���`��<�g�?��k8����w�1��踬�dK�c`�E2-Ŷy�8�2�	=G3K�;�>K�*�C�s<0<si���DWLhF��ko��1P}NGa� ��d��ؘ�e�]����}4�}��%��LB��&��}��w��]��V�#��s
���K�
 �>�Ïb���j��ʾ+��K;O�
��||��ֵ��Ã	V�q5����F�Ps��O7�:�cL�ز�4-NES������-�ye����C��?�b�4<-\g��kTB�_�jB���K�t��y��V�OX/�d;Ѝ/��a�'Ƀ�{D[%�']��&{�!��]���s���ҵ�-+��;+>��W��v̐!S�u��O1�Q�?%�$��p̱@\�d�H(�k�'ev�5�"[�"�}���f"�S�4����M�{Ե6O���o ]��`��߼cWf�tu�`D�MX�*�O���)���T+��D�����0d��[C�Wˌ��H>��L�����2����;�*�Ic'GW#B������Lt���x�Di�q +3�vX"+�_ݢŔ/�G�� ���aIb�����n��?��또����N�^Y�1�4�Q�h�կ��9C[u[�-�Eq�y��s��н�o_*?�{C68R����t�$�ڹ\�a�`�L���I(��s^��s�(�a�[R�:����>PV�]���&IF�W��m��#<�C�O���ۅ�[�Wo����#CYn|
�@��X�i��oZ���"�i�՗��(zX��N��/w����8m��d����IPZ�*���%���=�s�G�V"I_?�|1��.����eU�F���E`D���Yл�'hܩ�'��x�Ox��R���^ǻ�V!���6�f�к�K]e�-P�\��$`��H�<j;L^g�C�>�C� ��+�]���&��r͖�;Y��ۄ͇ǜ֧+� �Xz�*9a�c�`ò}��|��[�h�"w�v�Kz��'����v�r�,M���<�N<�![���Ȍ2Wg�&�8Ui&f$u �t��ɍ\aU��զ�aL*���i>����Kh�^(B�c�:���uDí�4W�C�E!i��W�!�?j|��?ry����(��v��q�/#��k��,�������*,����*���N=���$����ZӺ�Ze�ÅH�Y�=i�\`_�IE��!��u�6����.�{��R����&����ȃwa���:v �@�-Xukbs^*�]"�1�=@.5 �?�˧y&O�=+*��{Gz'�C�L$ ����||�;�]c1� ���]�)����
��[����y'�W���h�LV$��o���}��]P�)�q�"7Q�J��뽼%B�\Yܽ�-@�Hi0HQq �'��p˿ҋ]mN�V��'��M����h��ln��qg_�Z:�c>��V�U�U:�f2P�$�����`̶�sB_#�ȷ�vwB����|٨�/�3u`���+��lՄ��t39~vG7�u�]+.�)�MI|�0]_�E8<�L!w'�3�o���`�v	�} ������EZ���w��j�{�sR���f���x�u}#�����cnђ��?���
&Ht��,��1W�z�r��Iۛ\p=8l�@�����t�sm�e�Lب!2�Zx��%�!U���I��w���HON����v	����Q�|�2ZM-����� p��0�y��g��H$��)�1�m=���D W�AB��6A��="V�:� {՘��QYE//��������;2͂.Ͼt&�Z���3�Q��emN�̤��|��ˀ�����'���j.�kM] ���J�$�i�y������Ml��V�1b��a7.h��^fL�/�F���O@w���|�*��o����F������t��db�{S��Z�V�EU�U����[&$�d�3󆻭��e���W8��-�ů�9=��ʻD��F�lLlq����H�>�Ub1���ځ:���6��؛맜�~b<X� \*��M	0~�^k0o�P������L�z�@c{x�w`���Xt[A=�jx�L��C�?֙���_I�����T���H�9��G"�o^!&F�\�Юt �� �@�Sہ;��qJ�	�_8F��A0Q6��g�$��A�{!���ծ�2&�!�� �K�G�5B�ɘ��~/��],"/��(���Y� �}w�"��� ��
ց�"̖5 廠�n@��E�!�D�ҙ3�o%�N��9d�-���j}���K"ΗH?��D��}�t+�y�h��ӫ���AP7�����P>����%��3Kǔ�NC�Y��������$J�o{;X���ÖI)(�D����i|{Atw/@��Ҿ��3X2
Qc��<"mH�v�cI�X9G�S5��)^'FH�QE*9�[j����1��� #z'�=�OD��^rG�ގ�pA4V>(����#�>�F��l8�t��c�!)"��2�Y����w��{S�H�4FY�E����[�v�N��)�:�F�.�e����&ƭ\Y�#!��_���#�@2p$�H*[s �ϙw�,�������Fć���Jc��W$T[(c U�E�$묇gH�p�ix*V��soY#e�WI��X��)�7hBXM��p��eQp�����O�r	��X=�_j�nx]�����H�u��X��2�Դė�7u3�ʪa�Vi�K��� �#����<��"`gй9c�Ig-�%�g���۟}���7�&2_B��I�'	��*䏘�6m����;ǥ�P�:��c�� �w�8�	�rt�ס�ǘ�.�W� �/UV��i`ɋ:q�3}A��6�t� �+Ӧ44�h?���	`,̃��\�-6�ƺ���規�����^s%~Zy	�/�~���T�RI
[���H��k�hE � �E��|s,|�L�=�%��/s�EW����#
�qåZ��
�������:�Jc韛\��~�r���c���	�h�I�gs�� v��Q��s$�T�ڢ��e*��w�b*�OB�5~ao��Hm�F|�(�+��J�tE�-�����q��蜶�	<�R�%B�,[�xT�;�dM:)-�3M}V���x��5m�x=�gE�-��k"S��}��TF�h�h�^ĳ�w��b��O|�O� UoFU�Qc7�*n�=ZZ���=U�+��ɣ�m��IV�@�I�2Q#n�QA�Y��)\ܴf�B�"��K���B4�VUzcDk~c�:����r�ۡ�ܲ���[0��>D"F�� ��N�:�vd��n��A�������~�ʤP���䧦a-��q�'�X�%&�g���m���z!M<m�4��-�}�R��,��\ �#�J���5�Zy��?�%�P�,�����7�MZ�2�Z�ΩVz>�;�VZ���F����R-��RIƃ ��[�^ۆ����4J+��A��X���U�Ы������ ����[Bv�	;� �Ԛ��.����*slB�������!^�@'��K_i����^��J��#�)����] ����Ψ�[��K!�m�$����+����%/�y�"0��c�7s'���
oX�Q���K�+�T�f+!��}�$N��z�_x7�k���V�Ij	MF-Sf�$��hUt��Z	 0�X������cWf�-� YG)A��B�>9��"�5 ���|ݙ��j ��
uL��@or[��GK�7�c��J�Wn�!L���Ք��q`ª�
v�%�6�����ά�����
O����:ޢkQ.o���y� ���]Y�K��Q�]�FE������n߰z�~t�:��m���l����{s�
�P�-T:@|����jn��}�p�9p�z�R}{Er
Ťcd�_8(,��^Xu�U����}���O�A/�l-)�W�Q�)���9�UV���/&����rC�43�J��w?��Ѵ�=@~���r���4e+�Y�56[\��zltT���\~,�����*�@t�Z��S�H��u�5x�K���H�Z}$StקW��Nr"5���ۊ�ɿ2���7�d�`k�]7�b>y_�@�d�w�ĺm�f�Q8�5�7�Ҭ>���Z޻S��=�{[��v��Y�+[��R��7I=Z�r���<�����m2.��H�&-z�.��X���pb֓�E���ESP��^��6���]M�\n}Ř����j�61x����yUVM�&���u�e���w��8�tm�p4��<�Ї�pwRrZOZ� ����SUe~E>YC@���4�ѷ5an�U�b��"<�N����Xf��^�^S��c���M!U4��m�ݝ��S��#� �{�[��:Oy� *l���4�]'=���$�#��:*�������b�9��jb�
fQէ�g��l�C%M��p����[�ܣ���HNsld�y����Z�1�4��r�nn仁�����@�=��=���1 ���8�Fچ�sv��fS����5�%^57���W�ـ賱������Q*T�u�5�BɡU,�3�6�׮�ҡo��Bh)0jl�L����8qB�� N�h��G�������:Z&�$�R�����n0<���Ś�FC��_����ה�"@lz��%wS���CJ�T:'f�=�8?��؄#Q<9��[J�nU��ꦯ�~9�/�m��S�V���jUUz�y�V]����m�ܟ���h7ߐ�쓼��R�	FMJ���B��w9��I7�r�f����O&tM�*�c�_R, �V݇
��d��X����>	�_wwC>����|A�.���؈���pn{Z|
G����[���]br�8��<�A���J���y��/9ӄs%1N�7�YO�?��a�X,�����h�C����Sڇȸp6���+�v��)�~�k�cgr$�}>w��k���=��xT����tI���-��f�8O�SC�s'�p���W����>?�����񊝋�ImboIKݛ��L�����ZUs��U���X�Qn�������Umװٲ�YA�[����!��9E��q�E��y��eB�되%��ܭ��{a�Y=
Cw$&R�`��[�a�Mk|s�P��y�]6�yȚ�ܰ��(om_+��X	����ʄ@��	c&v*݈,�	�<�z)Z1�I��hֱ��Q�0φ�_*�Y��/^��b˺)�<�j��Q��j:�F|�&dF���V�\��j�d�Κ�[�N��kH�����P]3��V�s�Up3�:�p;�b�(Kƍ�Qأ��}:���ċ���1� U��f'�{}���O�z>�IH0 �L��a�t�Cq��90�=���B��(J��;�kQԢ��Xv*���&[���\��0I�wn�K�o*8	j5�����˂M\f�u8;�B��^@���uSfr-[���fK"z@���,�;�c$Fi��Yɲ�S�5s��/��~�;�Wz,ʧ#�Yp���Ym�������Qt���A:�Ku6����Y�p��y~�?�ڡ�XG��p�3W��Rh/��p߀:G�>�n.�q� ɹ�*�Ԣv-��ܐ��5���]Zy�b r�dA�<�+�OK#<���:Ĕ'��6PB!���Z<"�����~���*OВ���1/����-�tU�E*HH�3߫!�(x��c�}}M�7ﳹ{{l�c��jq䴥o�w�0��:�dM��*��:&�.�T L���I�ad
�����a����,س@������5(�W4)���M�-�(ki<�)IdR��5����]l��]�����!���<D#	eG�k+����y�V2�JT�CS䤶�`�j@x�����i�a�_4��a�#����-�5.�%1Z���D!W�\B��E�k��w{l�HH�2��c�4z'N�����b��mͫ��9�F����D��]����F�z�ª��!,�=�j���_�鰇nf���z�T��y	�K#��m$Q��a�q_�P�[o1�x��c��><�)�%Q�W�+��7��ȼI4�GE�C��y�[iȭ�.T��X`�H0� C��]'���,�v��gp��`����(�-XІip�j,�ұ,;_�ſ{��ʽ9���.y��,�d(�y��|�xC� G��C�bX�dY^�ѹ�};I 
���ہԠ��7¦�}��5�X|��?7#=���+k7Ky6&V�U���=��C�O�P@~ڍ�y�T%*;�r�>��x��|`#�eh����NH�\/��\=���N��v�];Ԯ�А�C�ڰ>�q��e+��DZaQ��ԩ%3�M�<�غ%�c���_:���_���0��y�|�w�-}a��������m��Rc��s
-CܝG�l�"���4�+?)㫘&��e�*������`� �F��mՔ�g؇ifl�Q�5u�����Y���^�e�I<�kN���|����]~M�6���zqK�owj����,J��[�a�6��7���T,�ƥ�1�c�?b�'1�� (Q�W�RT��<|T��(-���I{�[�k��i��f�))%��@�B��3~���^�c.%o��"�ڌ|s�
+MrY�?~�q�P�w�вw�a*��A~>/F+�F:��?��`w�JؤEưvj.�\a��a�Q9�mK�\g�ɀ݈���9s��s��zO�&�Ӿ��;�
���ʂ���{~3��$��U1mzH�6����m�NR=`���BN�8[�*?]t#瑯�0 >i 7d��b��kZ"Hհ��L�2<��-��&~�-�H
���q��&��Gė�$%p[M�zVm8�e%��.���6�(�T�'���:^z�%���x�`��n���tͯ���}[�vx�\�����$� O�x�@�-�;���_���m)�(�k%	��x���/�y��{\��r.�����Nr�C���#9���$m^�;��퀤/����D�m��9t��e����XLҕ��U�m�,Lҙ�Y�|��E~.S��0�u�Ї��+� }&~��j*�YXf9�k>"g	Qd�{�j�����jy�
XU0E��Ĕs3\\���Z�5�K�w1,��v�9�22��.�GD�:��Y;���J�΢�B����H.*�)9��|�3e!1H��n��[*w_=��ΕEY!M�1���N��'(׆���5wT|g��=V�ÜR�~��#���b�%;��*]7�	aZ��Gmf�� ��f#�։�F-�����l��y�0f��A��M��Y��ݠ��`<K?y�Fڢ.����f�͏Z�ps߰���~�^�,a7r����j�
�*,���!����E�N�1��;�׿Q捀P�CP�σi+���Q&�3Bd�;C��͒���l�®<��(��j7���T�Ӓ(�,熴�Ji�$�֮��$�7R9W�x��l�Q�������א�]�
+4f�,$6w�(���Ff�9�Q�YnZ쌃o��/��}�=^�ҍ���*���(z�.��ٟ�����O���9~��6�$��e�2&r��ucqp!Ҁ�����"��y%p1X�`\d����+1Om�p�y�_�F�( �ځ�{�kuv�v����J'����X7��f(n�[�@�Ӊ;�u�B��~`y�4g���Iz��;@�
e&�^��Q6Z�06Y%<jG\��}w,HTKA�j��*~�?�%�[c�k�)�+d���'R~-�z�:�Rg~M��o��l_Q�`M�7��<J���6)ć�g����� �Ceʌ{�����_W�<�Ʋ:����?�ķR� e���F�Bs�[Å�.�,]��X��C�~7Q��<�!��*y�/�������Q
�����nG�,������Lz�}2;`T�*�	��B0���Ny��
�O��"�<�4��G��Z3B-�r#6��%�L������2EI?I���P�t����I7
t�|nh켊�M��bv�:qřU��F_[�,�9۾ɼ��3�PawʽQ�mb0���a�����b�U➸�uu
Gb�O[���v�"���~v�;4:��p����᠌���Z�~�Q?���8P�a�+��5I�A�E�u�闸�,E�.0�W)�9��yg ����<v5XEo��h��W����n�kL7�ei��aiЈNYD^+����&U�(/����\����77�;уG�L����ǀ�jc�@�����ںV�-�����g��NZI�S�sZ�,�(�u-HP���x|:̱��(�T��U͌�q��'�D	]��V�aY	 ������H��S�ъ|�% ���d�[Μ5���.�hB~�ٙ�5@=/�z����x�yI,�v���׉�¿sq*��e�b�蕴/��M��|�Ӯ��h��v�V?p~^
l������e�K��=2˃�of���J�wgl�^XkB�?�2u.�4vm1(�V˃���X@	�W���vnr��%��6*u��eʠj�W�N���t�2,Ŵ�I��>����D��`^`��C�<�G��j�����֎�D}0S�����s�������$t��v��)G�K�d�)�
TD�깔v��F�;�͜��$�����ޒ�يږU�
M��\�~m5�7&ϛ�(�@���x� �S�Cɮ4s-���I�6�	Zp��y���g��
f�+�xtZ=K��y��cC����٪��漭I������N�	�+Ơ4SA�Ӡ�:��P0!y�� 3�A";�����1�I�`C�	P^��J!Lh <	\z��6<�ef�L3?��������a��%��]
�W��P���[�d�(�/�1�{�+	��7QFT<��7���g,��I9���&�k��_߼X�!W<䙦2���Zlq⫬80'����u�@����i������y!ƛ��'��*v��{�/������2��8��*��5)�/��ǂ�.Mb;�/��F��b���Wq̵NeM^X#��f<�gkO�	�t������Ҹ�'u�y����!�{�����W!xwqVrJq�k��H��F���q/p+��p2��we#ܳĄ�
����I[��h��h�9&���v��CHn友5�q��2Y_GݝP!���¬�zI��V������G�bjrr���e�дl��I��m煀�tS�g̣��ܯ� ��a���6��UT#��ֻʊ]�q���vت��[H?�����ѣ!�ya�8�*���:m]v�-����mF�X�
,,����,ܑ L�5�����=��%ӌ������HŶ¸	��Z#�`�^���7}gA�{5�t�e1��t��
�c4��N�"f�:��t�0:��F"j��f���S\��pm#Y�Rg����Wg�����f�!���ތ��	ׂ��f�H�V���Zn�},V	Z4
�7j�����LF������{tk�މSd
!A%$���Xy���Q?|(�Cs�ɗ���Ib!#U{~^�*�[�b�V�H��O�e����t��*6g���Y��������_�����?I+��_�$��b)B����A,��Q�"�+,��IS�Yj�%y�5N�C�n=�E=��K�&xDQt�
6+g��\l��㝰w"ÕIq�7e���(�&`���<�����xZ��l�n�:@�Bk�Z��/��"[+wVj�i����!��7lK��Q;�R-V�J3�B�=X�v�N�2��xCW[�$l��J��.�w��$����H��~�d?~�r��]�ަ�^M�+b��[0�Hg��­8
�?�	����Y?�+*�i=�YuD�*�]fNX��s��u��Ѕ��ȵ{*�{09YΗ�l\`��f������Uy��lx�i9R��u�7��>ԷA��	����U�	�iJ�����}a4��*��ɂ�#��R�ҙ��LqW8E(��_>��v�+�s��@>|
H#�S��O�Am�s������ܓ0]�zy�*A0R|
�w���U*(~�d>����,��0c����֟��c�IEg�� �ShA��on�;zz%�<��Ƌ����'B{3�|���3V1�
�����wr���J+�l3pF�g�ػ8 Qb-�B��:XO-�@�BgCK���$������M� ??cŝ���{�cC�i������\���#��X�j�EӀ�zGx��;�Q}�h�$V����)��]���VQ��u2b��؞���gQ)�]7g͝\g�<�^�T���X���IުQ��pf%�a,�$y���'iQ����%�u�횏�����r1I���>,���(�p�(:fw��{-)������P�����p���x&��蚝M���ܩo����3����!c�������I�w<hgH�1�Sַ 9/����R=~
V���P��Kv
Ρ̋ 	4	��N�:�'!����F5Ã�A,[����(����H`�.2�	X�^-�Рڽ {�þ�����7���v��2An��y�}?i"��A��&E N�0����&���`Z���ih'0��WXɲ0�����#�D��y2i]��sFe�g	6��c,�Qqx��x��z��{����X@�'��������$��	�®��b�/�����RdH��*h4E�'刋��!@��x���ߣ��ق���p���޻0��%�ݚ2ǸZ˪�t�.r)�VƭKH%�Ҁ8w�.�c��YZ^rC߱��C�T��MX�� ]EBԈ��R۲&���s�2.�����W������3Ƃ��b��[w��;�粴��>|f�.5}	�,@Ѱ��h+,\b<�$0�~��UH��e4w�;*|���oo�4�U���	���]8�~���/�"|�qb����G�HH��n�}>��in��`��<��u�IT�M��'k��ɿw��Q����1���B������r�<_ �.a��;�"���Я2�?8��>���2o��^QwaN��V.d� ���F��8�w��n�DL�����yv�Q�:� w��C�?-�����{���3�R�`�}GcC�B��i3ۅ��QC�e�7��q���L[H�ИE�򠺡.<�t��I�OF�% I�?�6�}�AZ�c濖s�4�{/C	R%�w��[F��|��H�'�	i�� =��\�5c����9*�&6�c6��f����m��l�ɋ�zCQ=�����v��v��#�;l�r�E�$�|�q�].g�RI��XB��]mf%΅��([�NQmڞ_ȣ-qc.��ڦ.�Ě,���D��s�_���ޝ��˸R��洕�ǵO�+?1��h����u�$�1��q6�kE%�1�j��C|��C%��<�fT۩����H.^�)�1���atSMph]<>����u��W�1��P�����O���J�:l�⬮\��"�TP&O'd�0�Y�YxU����^�*?�&�,^T���&��-��7㺜�)�W��(�(YG�9i[�Z+Vb͂N���wO����ş ?�x{����mx(l'�I6������,���{��]B[¬)�6!ѩ��yZR���P~�T+"��_i�KKFO�ۦ�V�H8�XJﮄ�h^�A���6��Q�<)�ȀM�kIg'�:�4�t[�D��l��~��!�H~9� ���/�R(�5)E�9pJ؃� pg��K7N6Y��ߔ�oE���x�t��Ƃ��)B� emu��>�2ϓ��T�8����� `t���_+�ZmIQZ\�?��e�4Ђ�6���P|�m�d�w]N�$ ��� �+n}de16n�)r"��T�RG�B%j�+K�4O �y��#��尩_^� �L8Sin�n�XB��x�(�V�=�M�M���3?��XH���2��֨�W�� ����a7	���9�nW(>-enj���MJl&�]�p0��i��oGr w9W�mp�Y_�����̎�֊MTxǕ�(��5st�9��m�*�r���r�+�P��&ı��c&����ʽ��D�VTy�'�����s�O:�*��=-դ.�'�y�{?v��U�D{�����U=��k��4�Z�ڪ�Ft�%qk�����Z��x����J���x`�d`���!���9���h&�MU�R��酉�Hى���`L���V����?r�%��Ә��A x��'K�>Hlo�ψ4Ρ��v�_ؿ����5����?R�K��3^�NCm��m�??��:]�ҽl�������3UmZ�T��>X6�y������}���W�p�o%���y��a0�^H"�ج��r�Ј~|+�Zq���s�z��pb��2�Dk/W���O��<�ʻ��[��]z/�[>Ds���R��ek����F2���/�k�{e�n���I��3!����뇊�%6JHĄ���|{ї #����5�!�C;����Ѣ8}֭��>�5,��ټ^�c�8C*� x�sGL�j�(TS��Yt�<b�5�=�1���D�l�[���L|ʢ�x}�R��R=qP����W-�'+��U�mkDf��#
5��oR@�J��F�^�sg:�}��.�oih�/��Vb_!�E��/>�'��[�CD��&N���s���*��L0��~�C��H��D��@q|�ί4v�:��%Ӫ�z oA�t!���pl���K�y.tf�\P��F� oZ�`�����Je�*�S��-7Z��F٬;e��_��x����F0 SL"nq�~et�i���*\�a9a��=K�c��ߎr��l����`0UG�0�����A�b�DU	� �N6�Q{�,�x��5���#-�0ѿ.�j��q^���G���d&MI��aq$�$��z�f�RY���L��o<�K)�E��zO�k�}ػ8M���,���M�N��S-(����۳�Ɗ�n�a/F1����H���8�|�������&�����f�y׬���Q)~3QP�u5z�>��6�f\"�.56x�e���c��r�=/ �,ҍ�_��KX/A�&�[#��I��#�w̧��_���^��6��DT].2�-��n��y���1ծ�	�*:�ѹ� {K��5�xp�m�&>p����$̩�y���PH���Xp�d��ɧ�ÞŜJz
�G��G�#�E���8�,K�r@2�����*�@|m�i�W[!D�24���# �;��l�ʒ����B�4�RD l�+	����'E���ioi{���Y���d9�MUV�!�H�P�!�Lg]O��zs�+��(����i�	�{z� �P[h��MZ���@3���ꨄ&F���H��M=����W\4~�z`ksQr��	.z��`��]��}5�����W�u
�[UKnS�>Q�x��&<v��\���H������:}���ބVf���y�N�f�^w�}�_��4�#���
�KL@Y��\�7p���(�>�kZ�J pä���e+j��'���W�q���0M���!ְPV�dx3ђk���A �UVbA�q����HT�qtܲ'昒�L+#���I�e�a�|5Ɛ�!�&5�s���[a��l��2 U%3��_��;7I���=`�=�إ�[��zf��:�n�*m���<�r߆H��v��@cp	�#X&�ܼȑ��l��b[,2�v]�\���8W� �n��h�W������Ѿ�;m�^��r��Hf��B=�f
�p�$+a4���7��j<6wnJk'�GnUS� �W�{�J�9��!N��73%M��աu��:z�Hа��ԩA}h���o.����ۋ�,4��;ak�h��
�x����f�kE��|��o��W���f5�˛-=6#����B�`9�\>5�����XB]�2N	 T)n��݊MFI�H�S�S)_��5�gP��P����}~:$1S��Y*ft]����Xʅ�A�u�����I����T�-4�+������}y
�Г���$��f%�f�q�N�-�@����>�fr;	QTX���B}�|�X�z���Њ�;�%��iYj; ���9YJ������P�j�߂2��~�x�ҹa7/'\�,��W<���QLdb����� �C������&�Ki:I��<�-3�M@<�)��ѩ7S?��t�_��iӢa�1&y _�yS��lο������i��Y���{x=�޿�@��7��)���.�2b��[zS��;�w��t[:<�\��c�Eg>�2�c���o%eO�U���5�)��J��9ԟ��8E���?�N��ϴ����KV>��P��
5��gߒٛ�vd�)��);�F��ܷ�/Qk�3�t�t� j5:B��p�� 6@8s3Fv��A��������IM��$��߀�]�јw<}#�ON�BT� !vw�Bf�j�R��19���Ǜ���3�#���8�%���j����}3���_IN��\~��MFH Q��wZb��2/0�A�)�#�+�N�޵\�(�p^���&��{���<��Q0b����Hr�k�i��	鉆^� 8�����7�t�,d������k��!����4�Ib/"DB(��O�´k����L�}v/��1:���1� �޺j���Q��9�����C�s��f���ά���}���z!������v���j15 �����s�KK�d��41#�%>�:y�T���gӤ�:��@Y�߭�����;�OHV $	���X���X\*ץT��^���1I�k���ԕ���i�W������c�DP�K�tY�T&{K(�^ۏM�aGc�ʚ*ΜM\V6���[̜��z�f�"=�3��W�*�ͪ�K�}�!&*[`�r�����e�a[To/��H_z�xsz�jR��j���	o�s�_�pCU�U�p��,��K���%��=l�bϺ�I"{7�/b��6��ߠ�!}���;�ЪahU*"��rP흷R����I�I�wdq�m�N�n���	��0/)4�R�9�(�h���ݠe_$h�?�c���## ���T���ʯ%�7P�XϦ��ޥ���b�R�g��/���HFW��I��#}Mgu�u���0�"Eh��� LA�0�
e�T6 � 4Ym����sF�)��8P�@��E�%�5���[-	<v��A�k�G�Bk��W	���� g��w�殺�=�n-2t�3��f8=���r�;���� 'S���XKJb�h����~D�w�pB@��KB�9y7خ�/�h1��2��h�8���۠� �d��\G� ���X]5N Ťi_:-��
�J��ӏ#,*��8_�
���4�IŠNem��Rh�!�k�����-�ISjJ��Vi�$R\������+T:3��y|��r#��r�aPJɜ��dE�`Ȉ�ġ!��zʴl����Y%���^q0���z�nw7��:�Vq�ϕ���'J���)w���tl�E���ny���ln���A0C��K�`���M4�Mn��`W&g��?x�h�Z�g��Nk�4����oU���`�����B2��o%�a���fo6P�"cjwn��ܡ�i-y�D��p V�(�4?xTHA����C��;�W�J8��H��)��~^��N�B��K��8�i���\�U8��'�����VM����d��R��O�\��G�쎐9l�:�Ȭ[#3hUN������+�� K�Om�U�B�Ukt�N�����v��7Q���CdEbf����w����߳h�*br1���gȧ�ᯫ;6�H L\˩4�r8�B�b��U�kQ=�ȳM)jl��R"4�t���YY��?P?|������ԕq%���d=��Ʉ���ΏwLO�$<�m�B���"��B�+���Q^�Ụ�C�;�2��WC�߻�lv���k�;O�ڝY�=;|������� 8N?ч���@�3J����͖��*Fz^c�g��/�5L�i!~+���&��xsS)Cw����� ��a;�_Dn���n�;�B[.~�p�]3�5�e�=$������+�ju�-�q~��d��핔��o���55�ɸ���#A.-�G��q����WEW%�r�|0ʟ>w��V=f,;�d���JҭL9��-�=����a��ś�T?�e�*˰e"X������h �{wA-H��(	EF� �}kB��!w��,-B��95b��}į�͈�N�ǝõ0�R�"��������u�X�li�JISa��0	�9�6ȶ�	�XO8,�z���|�,'��-�+��1�G^��F�)H
��+���շd�)R3�4�	�,BnP�M�8�qc�����೏�u��9����ܞ����q���\����t��v�m�x3>#^��{G��=?]�1�?m�G#6+����=��QQ!Qӗ<���븬�.��\/"���a��!�Q�����n|�H�j^Mז�P��a��Œ������ʭ8�,t�[z�(�)"�ES����·FUB7��$(As����P�����O_cN�mЂ[��r�Iz=̾��R�j��qA�;�a�l�4O��6�
^E��N����~J���s*P�..{��V��Y��L�V�Ąۅ!�C��LQ����aX=W�V���▫�u�7w!���$��
��(-�Xf��Ӣ���̸?5·|��V�ރRN"_+������\�
B������@ԩ��<��e���9�u�L���i�:'�x��6�I��Z���.O,��.	��)����|'�}"*d�UI�p�E�����~�摾�hW"J�e�,G�&�T�t����kLuQ�pA�	�i6�����݉����d���Mt���ǐ�z�s��b>ȳ�y-��A3G�镤�Fk�D�B`�f�S��V ���r
���;:�x-*x _d��,6B�z���w�ڙ3Sc�I�
j*]_�e�3l���t,_��Ǘj�^���y�7��K���� 0�>h;: ����� վ��+��֕���ϭ��\������x�z��>�Y�2j�+����G�&��>=0˥��$i��%�~�����>wU�OO\����;NE��B��c�-�e#%:��b�����E>�{�q��D���	=05; ��[�Ek��^���X[�]���1"TF���q!���I^�#}�a������b�U'tL������l���,�C�o�c�HHdK�Ȕv�|��ٓC\�� g�2૗�e�i�ϝC^mc�^���@�$
�Iz��D��&R��ӳ6� ���}^��7�t�Z�_����:���̶��Q�U�k�GIO�O�A�������n|���pi�j��� ���/A���?�r+_�ڃ�zh�<��X�?3����Z͜�K|�Pz ��t��i����I��&���' {I��o��ij��ĢqY��f�u	�Ib�`M7�-��g��C2�1�q� :\��.R��� ס������*y&B쾝CXă8C�1�O��������t�ٟ�D��a��:�/��0���M}m�cȒɠ�عN���C�aHS���Ԙ�<l�"5or��8KW��-gm�man�c���`�x��8�A�i�YW9�����Q�li-]�QH����*� �%t�Rm�7��<����C�C+�M��i((��ӜB{�@di�� b����Y��P7I��Q���.�c)��J��1�VxQʀ�d�T�-�kH
&�T O�	bbm��O3;��wIy���^�DHn��Mp����'� ��w%	��V�*�!���@C�<���2и@����?�)���fMcPHt[������Z�(�LY�{� h`�.D�AnW���tf����y ���7ad�%�_������T	�1�x`v�0��j*g��� <0�5�FG���S+k[D�!;�����k�1��Ê��ס�~�]������0 pr�(?ץ��-���^_A�vāRn�.[>^�s��d�
9��t��J����U��2��"�`B��ʐ���ܥ:�Z�k��YH}�Vhp&�l�˿��*sC�.Y��Z�.��� �$�q�lrѺ0���&�/��j�O�Mo�xn�N�F�Rb �L�3g�Q�� Up�V�=�!}ϐ�d�� 
U-�H�1�M�ȝ�tP	u�7��@����q���mPm"\/l���Nbs�(�=F���G3���#0��ɛ�L�hi�Y�����PC���A���O45�S�j��mpZ(\�Tx��Q���\cL��h�s�QSI⮴�X������I�`�cU���!�vS�".�u1����V[�ҡƪ[�wn���{ ��H� �ykbG��n�ƨK�������ߙ��ih�m�ɩI��UVb��+��ح�;39�2	zC�Ie��Sc�=�Cud����'����o�v5�@�#��3$��<-X�\��N���W6�#���cߚ��t����*��������>��?j��v��x����a��]�ފ�؂4q������~�7�H ��X�q"�}᱖l
����J�r�D6#�]s�������%��G�t����i�
,#��Af�͒�^�6�X���E�Q���v�| �c{<�*�쟞R:KBtA�(��vm�h(,Zl�?F�V��^�k`�,K�@�5�@_�Z�H���YWh�5ؿ��Z����1��ml�m�)���k����i�-��+�HcY]A*s}q�x�|"j�p�t�@����h��}�X�VO��}����\xx��R#$n��u����$���yJR[.{AW�EF\�%㏆�|�m���O��P#���hԈ���3?�*G29�_m�l���$��;Ҏ��YN�L���a�AnDM��e�uX��6�9KSba
�t�c8�Y,���?�h��9�����B�oP�1ć���h)�W֥Ez�Kc��fΗH0If��!V�L�a��k�0Gk��r����;���e��؆�)�8��a~la���0M���Q��"�ԷTB[���MrX��!Z�I�Q��LJ�����QJ�(O�S��_���@5�H(��5�I���fU�<g�h��y�T�����D���pu���ˮT�pU1 �P�]$���r�5+�t��/@^2G���8�atGT��d��[1}���a�:[ �OA7��b��:'����]<Xa�h(��9�`8��� ����Q[�����£��eϱ�W'S���Y����HT�]�,�I���ߌ�;���ƴ?B=�lw���)������鵄"ya.�\nG��3bo�=��W�5����M�&hɕ��R����1�l&�A�e ,� _��P�?�����+���w��YV�l�"�x�Y��'��P�h��O�ɷV�Ӑ��F�Uȓ"��ƿ�MDa���U� IJw����c��P�L=K�A{��S� >Ӈ�[����]�s�+�h�7 �v(�3dz�*/"=1B[��{`����F�am��t?77�)cL�J*�M�P��&���|�j���
5�*E;�j�h]�ߎ�(x�@��Yv���.����Uti�b
��˚)���u{�{4���Q9���7RomH#V��x�%>Ad�jH!��+.��¾�$�
�џ�4��]��j��x��^��o��T��=�t_����Y7nR�Z|0^��fJ��R��?�_�d��^7f4��/��}X��7łMk� �ƍ��#��� ,�*.>����U����:h:�$���J��W�N�� +�@[�+_��$FH�z�=�D�Z�;��uvG��2���Ǭ� �(vU�9x��`�
V�2K����kj	�:��V�׆Q�B8�IDwL($�{G�$(0yI*k;��3���l*À�H+���S�Y��0���+�f��ݔ�1m����9k�p��pQ��G+�u�%Y;@R%+��:P�r�V�9�/\���� "�El��Cm&��R_�����nEb�����H{��ޠʵ>Z3�F)�eW�=�WUMk/-,�Y����e"�U{���~rj����<_@��)�lᠷg�[B��x��W؜�<��Ѡ�}_���s������٘���~�����Y<�
vPB�PP��DJZ�������������ʮ��h;oU:N;Ņe��C�1a�mg7��%a��[ �k�=���Z��(����q{���?���dQ���su�=��$yoÕY%�~:��޶��j����P�M�U!��d��;4�Û5+Dm� ,ϜB?���E��F����"4^ռ"�~p=��͒A5+�$�Sb��%r�]K�}�� ;CY�.w�IM�'Q�>N�#�k꣮H$�"�\�J��^칽ͅ�Z�V����Q�C~F�R�bȫtoT�SC]$�Ш��⧠�ew�ʒ����lǠ���H'���p 0,�.A����T4�|�'�Xv�w����U��e��rr��<�b�ώZ��g=�5`�����J���*�s2t�l?�av�+��X;A��������Q�O���M,�CcnĖ�a�� �nK.�x�պ�<��&°�H%y<�tX.��WI*�ً@��B�更��X�zT����a��r�5 aE�@q&�^��Wk��Њk	T��!�oX7ϴ0:x�[N��E��|����>�K�0D�V��W�!Hĳ�����+�?of?�頞�T~��nbA}�Z{H�h.4L��K#�oP�ζ�U�Q��" ����>�09Λ�l��!�+���wt�u�)�:Ղ-�A#��D��_�^H?c�Q`N���߄Z�w�;��{ip��oK�hŉ1�r��W�|�Ut�>�i�JQQg��)Q*xfI�Vj�R\\eiO��X㵰2�[8�a�(� !����������=�d��Tc��K;+��c��9;��>X��|eg4��z�0�qa{E��sf�6(�GǊ�Iujdn(�9�5A�	���!I���~�F�V�С9�I��^�T	��+rn��n�L���F��19=��e��6���
�88`i����5B�v�Q�)�������-ժ^����gD�A;�/��2i�`M�^�6���
���~:oB7?,Z��嶆/�R���j�?��y`Y=~�2���xy%޷���c�0�qS�[xSn��S�X	��ԕ�8�#�3���R�"��7����{R���P��*{�o3�"؃�sK҆��8��YA�(�j�:��p� +�B4sҊ� ���P۫��$6�'5o���]LEȕ�B��
Λk�{�N��7�P���s��&>cm����`M�	,ݭ���]�t�چ��np;�Y�*�a��^&��������"-~\�d��F����d����D���DY�|8&���+� &y����ʺ��������hl$�N�����ӻ��Ϥ���y\��SWa��SN #;��3�ņ�� S����uv7t��}�\��;�3� ~)��XGY�8��Ȑ��_�����%*��K���܆n��L��:�Zm�)�����N�n��K�=Jf�R���l�RO:�vR(�Rk5�#��Ă�J.���Y0z�B3W��-���%���P�a��,�3�e �X������bk���E~F������]{^fZ��p�(2�I9�R�KP�`K���n����0��V.Л����܏$�i���ۍ/W'�?U�W�G�`�7���O�_�t���pL�>GL�-H]r�=���D �*����u�SF�����Q[��J�t�����U�uS�
U`�����b�L^�3�fhqh����"��2l��F����:���eډk5��ž��R���,]d��=}�2<hZ���J	�o�P���ntgT3S������Ye���$����@����\T�����YLߺR�0q�F ��z���A#��,J8�%��n~SՁ�<]+���������da���(G�=5NS0��Y��xTM����&��>�z�8��)'�n��f�GS��������:��w�n��g+�^�B�ODu��H2i�4�f��A�>�HE�cZ�")ds�k���9qc$���g��,v���\����򋛡� )[i�̜6�*a�)�tct`dIp��n���L�2���\�n^� ����)p�c���n�ېs��ܾ@f�q�J�d,�{�����������)!SM��{2�ʦ��?z�_r����R�&�.��?�8��mI?�d�Z�/�z����!��'��W(��r"�gЯ���0��{��SK�q�B�3-��ո�p��r]���Tx��A7���E��%(۳����@`�W�U��9E���g�̺ �꾏V�t��!wWfV����	���/��I/�IF���r�]�n�����bO�������#HX��}w��/��*Ќ�0V�;�3��qT����Ts� ��`�0(�΂��5�Z|�m���Ys�U{ZUfTQ����߅
�E�qme2��۽@���0��I�]&���3S�[�?8���H�{{I�8��'�Do�]&;���4�_�|D"�+c�c����-�S�?.ZuԵ�'{�����%(��Bi�;��e9.6]ۻ�|����t�$�`��1�+�`��6]�rcWi�	
��>�O�#E|Hm��]�e$�c�0���uúI&-@�%�zp/V����Ɇ��
���T��礷�,:mD����鷰�l�(��,
�Y�"+)��	Ћ#���Ty/I|G�݊�m\������F����+��� ��%��{ʜ`�K��h��ia���B1����< �;�hT��W%���.|]�q�p�)˥����^R=����>�������ۢ5bq���;�\w�]����\�jj*z�v��؛�:��rKd���-���A\�Y1g}�C�������<���QK�#��6�[�0�4{��O�M��ȉ�7�cC#��/�8gܡg�A-����|�U���Wh�ҲΟ����T�Ar|T��������=�x���?ڂ����wS�"^��<aɯyĒ��ٔ����� � �%�-s�0���ϊ1��(� ������hn�4����������\�������bKuɟϾ3�¿��UOaD���}~Q�:u�O�[!�����y��G�$	d����#�U�-5������-wXv<�iP� nPD�|�7T�}� ����p�N�5<M�(u+��JGUxd��MJ�'�SRc���?nn��sttY�V�f㷡B1�N��`��¯��xB�"m� $�6��}�����Nժ����繹k�<��M�q2L)��# �jj:IV�<���ϱ�,�X��5p��e�Ηd�|=]�?a'Ÿ��×�����d$���B�	���9�k��0fD��Qi�A?V78J�vC���*Sͫ�.��YA�����W�"������*����l�!��ҹ����~��Vk�~<g�MՕ>a;�UfqF��@�"Z)oo���C�%(�/�W�!�e<:�i�'n���~D�=Tw��~��������7����@c��@\����w�YV0�]��
�)�ll������G$�n��h�#d����ZU��jxRB!<�t��Wd��FA51:xR��`.����ؕ���ƂV�������� d� �K���k�麐�%��z��?�{�"������lz(BU�|���UR_RRm��Me���UMr�J����	<��JŌC@�R����T��(��B���:dmH|�S�Η������䡁�6�l�P�F���5���@��%{fr8���_R�s�.۰��=�i�tmI9^L�<9���� �6�9��%J�r[�%,��&b*3F�<)�q&;eb����h���ʦ��S� =9E��[S��ќ�2�^%r�oy��#�wљ\���p�.���If{���SiU����r@��n�у��MIb����M2�+Up)F8oX( �}F��N���H��+�&sS}l/����#Lf�����b�.m��Z�F��N������]L#v�8W�S�a�iX�ً}�N��w���{�������[L��F�:2�M�׏n�E�,X�,�؆�d����'��T�ߝ��~鴝-
���MӨp��qS"pb��Q��-"��m���Mq�#�~=p�X�S��M�s���VfF�>hڥA����=�bhs�'�_��@��
MHBy_��R��/lX�FXԩ#�xN����٧�:�rޘ1�����Ė9��o���T���F��4��{%[5��5����x ���1�44�v�.F�q oy�8�h~`��hP��Fh��X�mBNf�>qy�._�|%$.��wމ`V�����tVg������%X�l43T�5����(-K�~qP�9�Ҵ�_y��*�f�I� Z��CZ̚� �W(=E�LY�����0���X�>�N5�����۶�$$�J��ҾϚ��)��y������שp�C�x�sCu'Ď�3��.�V�g�a~.���T><��諏/�h;l�{<��]L��F��~�:"`�z�̩AT �6߁`�H�׉	<!��_F.}su�  I�'_!&��1x^$����Z/P' �$Bg��jK��Nc{Ȭ�;l.��s�"���D�kL �f���7#-���e|?��P],$#e��K��I��������#��S�h�+2N�!!o3p_9�Y��"���F�PܘS�;��1u35�)j�2��'!l���1�;}d�ܼVU-xCh�@��MlNuG]�0@�.�����Z9ϱ�绵�k[����+�W|W�� �.R(;j}hד ?���~ҕ9Ӓx�vh�b�>�%� �$Z�5ک�Tm^����;�5ާ�(Q7���'I�3�˖0�`��31od ��M�z�sz�$�BR�P���F!
ЛβZ	bz��K�-��w/��������s�R	v\qcb!"��0�j@��r�f�ɕ ��|s_���r'�NI	��<�W"+��Ih�iܸ��@�(P�n�ԵUw?�c5�&��O����+xQX�ڔ��m�~e�8�u�j���U���R;��*
���'	�f�,r��)JL�{C_]���,�w�2��V �S����Y��B!g��m<D-OL�"����đ犰\�73�'���Rfeo�\�ӿ�ܷ�<��D�jL㇪��ƿ��z(G��Q�ЋBc�S�.s`�\�^�f�[I�(;v�{aO���xr#���n���J�,%O�? �Ub��N�Qe�<j�=XN��o]ͭ���;�{V�I�U�F��cD��zh�Q��-��щ�62�~�K������=��삫ѳ�]i|�%�<8���s:5n�VQ�暇+-D ���VI��ѽ��1�x�*W5=���n_�#׶�֠C��f����F
�
����D_ѥ�S/��8ɑ�Naqqw���#8�����(!� ��̢\�鶪�o��`�W�q!A�`��ǅ�9|���Yuؚ���6�B���r[K�c�+A�!`�7( ɱM���
l�,rWh���l+/Wd�'r�{�ʡ�T�}�չ��'*���Zq
l;�E}�$�C	EǨ�AyC_����w��ĒrQw�m����"do�>��3.���� ��?&0�����5�@��L����Ot��/��I�D
cV�3���oR:;�}UN8����W����&�5�>�-b�V�z��JU)(��������YNE�����ư2\� �✈�Ą��d9ˁB��X�����^�V�@�j�� .J,�θA;e�˜#�r����CfٿKѣ��v�y�x�[��F��>��>Xo�<e���Y���bD�(P^�|��o�]����y�Va �Ϧ6� ��G	�bE�g�Xё�I$���ȃ��c��k]{��+�=��z�_m�΅/��?��I��� ���dr%!!G�ǹ߂EM���qZ�=�l�P˷ܑbF��~�	B��w��j!8�L��{�J�);����WT�S�Pu������?��ߘj&�L��!f���Ղ`�ˉi����_�v��P�S��V�ˏ����x����D CAr/l��ܤcI��.�J|sN\�����$5�����j�+�<l�N
J���P��Y�� �3l��W�)��s25�M��L2�C;��xb9:��?g|Gf��p]2P��CȜ��@~�w"d�Z#��`��W�6�7���_���Y�����	��7۷B�쉭�Id>x.v�S�ϫgJ'�:(���a�������U�nM3��]��z��J��Y(�߃�ų������.�w�ߓ���6g%�2�9
S0몾�X ��j2W�m&��$I�<Kp �?�Ey�H M4�r�BtWH�٨\`+��z��o �S@�dZ�Qb�2Q�$��LO���b��h�t��t�����h4rc�3�x_�\�b�O��:Iӝ��L�Q��2E�,���E8�U4�<|V��AM6��5��%�.E!�v��W�)�$C�~���'hT��}f_�P$�"u qv��팛�t�.MƴpA��L��l�*{HŘ�w�b��s7�83�Y�}��%��p	�����Zc|���{ S�k�DbZ�����U�X��݇�VC�r����1�I�QB�������#�P�QUĪ��P2��usw�*��ܑ8��b�ՔY�0g�Fh�i�ƅ.��[����^Yu����8��]�ᎉ.�.
��Y׃�����_�8_�y��r�Tߜg��lv�^9��~}�2]?�E�(�A&R`0Pܢ�z���Q�l�.�[��w�?Nf1M���K�hW��P͛���(��L�<�VY��n[��*��6$>̒6���o�<͖�\1 ����W���}F �j�3�*3��b��ک����e�����(�/my��G6X]y4��٤m-d��1x��d��Z�K(����T4���������y��8b̡d��3Q�bu�s�ͪ��J���%9#@Uie<$yl�	�x>I�`ƨ��X>�6�z6T\�8��d�-���	g��9���c�uZ��Sj�}~�Mqh	��`�U���$�2�;��a�2�6��u&=���b	$A�U�J$+��\�8�I5�y�onS]Vr�vX�� [e�"��X������?�΄�oe�Ws�R�+�}p�Ѣ�u�\��Ƶ���؀�j6���$�Å�B]���S>�o�ؤ�P�bt��
���[k�B3� �=���\ߎ&�q�@����p���h��Z�>�1�|��J�1��#�w���%0ۤ� Y�G<���Sr|�}|�T�t)z&�c�ܮ�����*����2�{R^,%�`Q���7��4�{&Z"� Ŧ�c�Dꐈ޻��ы���VWw�|�^Z��ԤƬwf��!B�U�.jލ��&�% �$J9�w������N�Z�����jRIX�S~�vz�+?#�A6ѶgD���岳�|m9Ƽ��Gmzp���|��T�=���^�7��~bWNp�i��<`��I��1���p�̛�q������h��u�� ������� Vr��>y�fR�1{V���SK�,�������y'��j���;�te�@lE ��X�挖��c';z�cܢ�U1�����b��(�3�'E�.�fa�J/?�Q�2Ry�|Z�BGI|s:���~"K��0�T<x�S�`0+�t�3�Z�4�u��u�B�4o!Rr��"��!��])��NÌ����o#afy9L!3��}ɷ^`&��1e��\�V%w���8`b�J2��+ex���O�0��νC�f��d�>etbH!+k���H�/L����e�M/�!�B��e�`&.��a����2�N�����
�$��0�h�kL�TD�	LWmh*�R�P.ɂ�\�//��x��¯�`�z-B�P)�^��ˠ��h$��?����ro�b��B���i����,x�M�ͩ����9&��;�YB��J`�r�E��. x�'z�ob=t���>���ɺ��#r���a�i�%t34Vo�RQ^.��?�|�z�%-6"���OUy��O"�a��h��V�_��o�v�� ���y'99:�P��,�8������r�P�j���cpZ�	���-6�/�.R#��fx��OCG�`� ���Q�;z��{��r1�oZ����\GA��Ҥ�s����`a�����s$��ħ9/Ԣ��Z9@�$��R@b���m��J?�!��n�=��M�	��F�f�w6��1D�����`{
[\������4P?��2�/ɸCF6�T�߁cgUF��2�A�_\�����޺�U�~���c�K�ǟ<�(6[˚����Ӏ�J9~q�ȄL�/��*hs��ܙ��74�v��O>ϭ�M9hS6���c�M��&+?��,����чs��6�Ļg"��kp��X���	W8����v��X�F�Y�X�i�{��ݠRNi�"z�y*f�i"���� ������S*pI�܉�(�P%E��@��ҸE�hHz#�/z�o"\_��I��j��8�>��q)�wW�\<Q��P��X�:�8��iA�?	�,�@��` ]�������PA�#DR[����B�'*�x��:�������I�2+( �hM�DWK�;����#7�X�D��BI~_�3.7�.�=�5yQ��N'xIvX��O5�_�.�M�j��hP�WȹU�0п=��]h�~�-7���0y��Z4��h�#�0��(���uWL�Ƽ?x���X*0��p��2�*���T�S��j�j�/��)�6AO7V���Jٮ�E�a�t�8�M�z�@&��
��Ԯ#}>rW��&XŪ��S����0s&^f.	
0�tsMo���.�'7}߲��c��2KɊ@�?�iV�����ct��Ǜ��u��19+�`��ݿ&Q3��I^���_4�;(��[К�z�����rY�"5� sFZY�%jR�l]�6g���Es��Q�DԳ�	/,(��e>���H}<��E6�fMe�Q�sfy�u��ߜ�G\�}T(�P��0��'������4OOd�JHۆ��S�|���s��?���N����a�W�B�I��>�%/�f�����Y�3��:���9W�|͒�2�B�i�Ś)��F~��y���A���`��V�����+P�`����/�]ޭ�ڈq��0v0 ��7z�)�}�N�73 S��r<���T���üH�����[G!�����C�6�^�)S��1<���Ι��5nR�t4w	S>=�a(�"0�D�����;����������0����୶��9-&߄m�F�4�$6Юі�B��"e�A�U�F;B��s>�U��s����Ȋ[�o�Z���L�L�6VRf=!�3F-��`�	�.z*��-zM�}�}e�MaٷiW��_�N��7��BY�5��1#���3�]Lr���B�c�"����[=8�B���l�����֭SP��za�W+����S����v��rN���l�u9g������U�Y;��KG�.���cm]�톢�p��ϣ��!#�j�;�L�!D�Z�Lz�p� �_�G%ƒ���#l ��K�B��ړ��e�O,�������7��shҽ�- �o
Ճ3q�����Xò��`5�F�:���qW �ɸ��u��|iᶏ\�7��8-@��t�Y�0��E+���/L�p�'�U#t�%#C�t�tY~ŧD4V~A�|S��=@6߸|�v�k^������"�ɸ��	\���? �7|��{Lg��� �O�g/�v��_�q��ΧHX�e홇�p��+�'�n��F��Ł)'��aa�����%����K��U/`1[@_Q��e�a5�E$w�ܔO������U�>`
W�O�>�g�I��X	m3�w,�!��m�k�2�=2lTz�P�s㰤�	�OV`�t1Y�85�ƞf؝+���Noq��hp؊tu�>�eď�0���[��/ɕ��DC�o�����a���d)t��T��ṵXٞ���l-��' ��-w���"��\�w�2�����v�Y�[s�a�-q]C*mT5�LlI@�g�	 o�+u*Bd�ڼ�5x���*tԵ�!~$� ����[*BP����_���P�2w�

AC��o�O�� �"��C��U��H0mԁ�d^�֤ta��#�6~�R�"W�ͳ�>�����b2�p�#i;'�����U��Tt�3�>�x�4W�$G�rO��ߺ6L�x��<�WV�#�,C��'� L
+�^�&⑝�vP� ��wgK�� ��7YI�aU��&��U,�'��%x\R0�v[�����l�(�˫�Vz�#I֦��m�c�ܿ}?3)��E��"T@�`�zv�j �;�w�����ˍ���a�Y�-����q��𦥐/v���>[�����O���*Q�'��� �-}Ћ�S���;!�u��m�)[	w7�F��̔j����=��[���DA��3�s.��v ��Q� �ٰ��] h/���\ �X�^���Za}�?I��)�DH��`�q���u}�\�6��
�ϣ*d	�;ǥQ���?̎���YVI&��@<ە�sy	���eU��B8��j���b�F�+�;�3xs*R�>j��I�∰V��!�pN0��"I�ȵ��^�����I�0�9�[<�G�'Y�y\8�� 1��0���2�p%��ީ�SU/�-{6mg���OC}H�ø�0����ۢ�s��W������ޗ�띴�*aL`���)�է�ag:Q�|���ze�����{U���֝��*��h�'�L$�dr���מ�������c'J,�>�f�e�a[!/�����k)Z�,��a�u�:����@�T&�H�V�Bo$�� �GJp*$B&|�l�'�Jeؚ����Z͂�����F��ٸc�C��z��|�[
}�b��!����UPN{]խc�H���)w��4�i��Q��,�)�۸t��239[􄦷H!^��	Mp��ΐH�����ȕ�_:�y��[�z���L��y����F�
ZP9�L7%��SX�j�_ƌ���Ҭ�~>�c����3�#�_�|c��?M1|�r؝�-ZH���-�y�b�� N�4����^�~��������J��/�o�t��e�8��~�v�P˼1���Q��$epGo&_��Xmh����Q�BOPx���+8m}�.Jt��f���i��M��1��X�L��o�Ǹޠ��-CL"E`}���~JX�Vv-��2Xٕ�#2ݟP���d��,b�
�x� Pk�V�
�:�0ޒR�C�e�2۰��\�ksD4܄�^v����%��Ks.Y\��AِG��:0W��G��b

C<��V�DkCh>�S�U������4d	R�Ӗ���2���uZc�Nq^)T��F�`tV1*K�^�X9j%���t���N�S��||R@��p�x���}(-��d?��f���*�����9��	�gĎ�w�;�s�M��,�s9��R(�8����3�)V7+�_�_M�)Ѷ�q0�A�5N���l����N,���庘�t�F�J����c�a�-X@�@��T3f�A��ݟ���i�\7�[�b��׏1�h� �y)��&2�<�гOI�7�Ey������(d�����P�������B��L���;�}Me'|�%}:E��.0C�T�L!0L9P�t�y Υ&��'�x/�psX�DG ;�1�H�nzG�̰�Z�㯡E��́�w�Kl]qW�Pa����-/)UW��D�>t�*)_g��&A��"�/#��7��A'���z������ЊvJ}m��'Jʓ'
=�+d�;�捄iC�o-�.��
�i��E���}M_Le��C��m�|��^k����q��M�o�I �¬�h�t(GON�TX�TI	�q�|�_�"Ef)X�#63Mg��

1�Ah�W���o1��p��۲�%v���ß�&��E�j�B��"�˵��F��]S�
�Ӳ5��ȘʉrM��H_��cXf�1(`�5AK��s�]qPag�	o/����P����C}G�Q����Z�`-�[���I��N�+��[J%�%R�H�6�d�ァ����T��Olw`���i93����������ҎЍ�����Q	g(���n!�F���
�,m7h��"%�qp9u'q��QTV����������)3�����g6a �:D�6���nb�:d��˦�r�߼@؅Vo`%>ĉ^�t6��G��W,i��mC���l�Y�dm?��!C��0�&O����p�$б,�+�I�C��2�����K�쪛���yD�!:��'��� �V7�7��	,�
���P\Y��E=-*f�����ӏ�(����'��,C�r0�ī����'c���8h��f��~�+Sq���-Rus&R�0�S���<��T./�V�ۄE�eT�1��s�������JrD���� ��|>u� ��I������_��)p%�$QJyE���2�bh��'�g�
ؾ�6�"�k�^�4$o��!1\�:��3$���Q�@4LdP�5M��ݗCnӗvQ1�T.�h�b���j�K�,T���=q���4/*�塑��*\_��N���}h�3��U�4A]m²?����kM���#.����|�A�<�@d��խ��&I�C����C�_a�:��`����+V%�*��Br�'?���o���e�X�������Ѹ� �q.+������9u�uv'U܃Hi�:��=��G�v)t���4m��b�Ta���L�|���R	N��NԽ��h:V���ɼ$�:Z�x	�c��������^��p��ؔڬd~�)[摯H�'���~�m|;8���
�����1�?@*o��/���Ûim�_���v�?ē/{� .�{�������Z����؁�,8%��6�DfE����j>_�;���0@�*Ww�C;��	�F�1˓�i���3y,�|\熊��$͟���_ ;�SL�$���aO\�g��`�:�eʧw@h#������Z�����|�3C���Ьg�r��*�� �V �+4���h7a��pΊ3���ai�����w'��a��oL���4�T��6jH���u ��i�H��p`�.k�
W�k���eZQ�]-$՗E!�+ډ~�����CR)�;*�C��a���X�Ѕm�W	T�u�!B���W�61���E(�J���L+���3_��k�nb#_*�������u���|�Tm���dpH���~}-�#�~(�:j.��<m�uѧ���׷g���{T���[^���6x�?��c5���7&Q��q2W0��(`?a��j�Arwn�0�`3&i��FҨgK����j0ɑdb߂�w� "7i�d�<X�?��~�,��OP�qtL-Lp�tȔA��s�nAb��?!�'
^���Kf�`s�#hI�JP�iF@�_"l���s`)YD��ё�rm�Q���	>��g�'Dr���jzc���]e ��e�	Fxd�9&��r��nk
y�]�{A_��$	x_J�ȐY�"�N������ó�z��~���p ���"�/_��L���i�2a���R�m�Z(Q�}sx���U!g���h.�9�^��,�8����2bȁd�o+���:��S��e���S�7ܕ;�c��׶�)��XE0�3��6��C5�-��÷(�	#�]]z�x���߇�8�-���SՃ�c~��f"�Vy�u�<�y�~�P�w��Vxο(@Eb�@���w��e��G明��!3w�p^P<j>��ㆽ�mI���EZWڻJ�
�lOI�s�dT�k�Lݣ3
�MA1]�Ge�4��ijO��	�e���}`BH��?Մy���TֶI�D^��Y����:����P��[�{r����\�I���ﹷm�lTP���JqӝL��c���!�J���ub]����	�TrC*݅�z��.�Z�E��1@��Pd�����[�g��	ɛT��$	#������C�60j�k�ICn�%'}P���@��0r��[s㣬�d]j̻:�������:F`����L�|֢Rd��9�fcۈ-T�Mِ��;Gm?jkT=вDy�����K�s�Kŀ�� �Z{�����eU)�(�T�BZ�攮E�t#�꘾@�3;� q}]N��/�3�F�=jG��
�mq����\��JU�Ƞ��C6���*`�I����J����(�q�Oq�yM���+�'/z�y����l`��cߊ@}A�#�A�ʭ��p|81� �[H%7%�SH��ku�2�l�f�j���?��;��}��_��{�R�G�Dُ��V�_
y!c���M���sj�o�����WS�� �-�T���$�����q_�pY�6�I /����Hj�c�IJ��#��܈*ƾ$C��0�|���K_��\��P"�R�x^�q��l��ik>����^7y�*�]HjR��X�MIM�[<HX?��XҚ/�w�뢱�q��8sz]��*�#����1�����6�H� ���I*u�jRQ�������7�Xy�&��_+�|�AZg�.z0d�npXCK��G�h��p���{����h������L��<��?�^���&jH/!R�6/d�rVOp��*�K���}e�N�,#cj5-4s�؂�õ��pix^>�3Ū��X�M���)܉B��C����W�V��|d�L؛��Һ	h�"}u1�h����h�S����s�m+���6A�[��y0J[rZ����L�u�0A]B�b1 s��[��M �O3����1��l�^Czkе�;�w(�J|��T) �$����t�V�!*a��̫'V�� �(6�qC�>���BѠ&b�J̗��M��;���y�Y�������<��le&���"og����W���5�,r�1ӿW+ :�3>���x��`,�
������{pyǄ�y�&j̈�
	Z��k��&T����|�')y�D������H�l�c��q@���m����+8_�3���)q����'�E*�0M��8�Et���Hab͌�;��}~q��5���[�gCbe�'���v4���SPA�-�-k�ۨ���Lwз"I�@����p4�P��,$̴	�ἆ\��ͭΔ�{n�w�@Ǒ}?H�_ܞ�Ws�$��v(_"M���<� ���!8S������Β��b���؟Ď���L��p	2#:����w�ÖC�Rbm[�����Ua�����N�.�{O)�@������ړ�}u\��mzT���D�ّ�8���pRB�p%����	{�p|ti�?㾐��-n[�5��`�����d	��Y6��x�BY�''���E����	/Jشc]���L�.$�WKŪ��0�a<����u�?`,\)�2�%��F���T��|Z7Kv-S�`�Dt����T'DJ|֌k��U	��4`.W��#y��M�X���B3����&�[��.`٬'��:�UU�GN(��>���;$�
M��Q�����.��eGlg��]���Ԉ��*ά��u�ʽ�H:�"��$�w�}��	}��!tt�Ӈ����Ƣ�v�󱰇��Öi`5����o��y4�|�O�ɢdtwI5�q�͗��IZD�I�E���d�K2U��Ax���{	��hݰ�BG��Y�ZQ�+���4rNkA�xd��|���>�UGtVJ
��\J5�.���ųK��w����5[��q3;�OhC�y�l���i��r�\��O���9�zԗ�;A�3a�U��SnH�a��<�$�!�ޝ]/�v���&K���,��`����T��j��|y~���zc'R�ON��Fk��Z��q�=�6F���������9���z#�L�ok���' 2�ds���\��Bnp�y���X5uG�^�im���0�?���;�Au�"�!�xǮ�#�u�z�eO�e&!�o3��k��^!�s�f�3t��nN	5����v��&c�T1�x��Ј��7	N�f���Kht&���}�v-[L5MLeW����8&���M��c2���(�ί�l�=��t*	I����Ld�9C6�����	������ETGf
�� ^FZ���W𘻷DC�3�8ܥC�
2�
@x����A����d�����/���h��OM2�bMd�%�L��Y�$p�O��|��{E��iN�֯�4��"�=��H���]dS�u���-|.��o K����U3X�u�-�yCc�k��Ba��0�~E�QKdM
c�ĖX����j�����0A��-j��u}Z����FK�q ���4�(8bso"��e�Oتʛ&ͱ��3���#�2GB��+��i���$qnضB!��li^#b�ы��7���f��:sc�N��WV^eo/�7��F��Xf>8�0�z�q�!�7�Le����:	����J�L?��1bOc]��nSHi&cd�y$��Y���iac���)΁�Q��*���Wk���l�S-��dp��x|����^��?���'Μ_�bj`򊐹��8�AqY@_	�����8;���u�X��ޣ���\�b������oCd�!�-����O����b��#`C+m=j-������>��b����ʈ7���$��÷2���̽�:���t]!3~KSyv����9�bۯ�� 6�v$Oo�\��-?͇���k���Ha̹Vj��3��H9.W�պsM ���m��'B��Ǖ8�/���|��-���kg��[�;, s����K��c�Yä��ȓ+.`��=G�#��oI�l|0S�׉��o���+� N&�P�˜!r�40�(���_gH��`FX=��7��������c����� x
ky*�c%N^~�����g���,��� ���U��*EZ9�R>jB�S�����ԕ�E�����H� [�6��T��UjxpB�� �Sy��k�V�#� I�YЫe�8<�12����X�Oߙ�/u�/�����X�����������̈́X��������3��ϬL�ò�_��ұ��8�X��͕o���Ul���^�b���R�/�	)ްC���'+��>�(��H&�sJ�.����o[��H���/�{@�fl]=��� �QG%�|fw��V]$�<�����J�5��vE&I��Q�/�d^�.%����!z�'�qt4����	����?� nO�)�<��K��ҟ_X���2,�	dN��O.ӵI�0��h� �YV>�a~��2�˥U���i#?n��O����I5�dj��?Mj.��H[ĺ����D�� �ʰK,�T4�l�#;&Y���&�igy�/��|�e��In�Tk��y�������jߣ�"�Eq_�z��%�wY�k:Tze�n�d
�J𭟺��.u�y�w?����0 Kɍ�	M���i�:��Y��:Jn�hF��;/*�
L.	��\>�;Xqf�c�;����p_:G�*Bo|�N?�i�,˜B��Ģ��!������*�]?���NJH�f
�+$ToL�a���daF�st�pY,F��'�J�,Ҷn�&%�.�5������v�92�� �<�-�h	�tG|N�C�BVK��ܳ5vf���'g�$10$�Cڄ��Ӱ�;j���Ĝ5/���^y�^~�hpJ�)�Ϟo��@]IpX8D��Y}2؁���>�_W�y���� ���s��[��cQ ,hv��L�{n��E�՟潍�N9��PaT{>��[T���vԐeֈ���#�M��.����UJ7��^՜7�u��fp��K��b�X�^p6�frq*��O��>܍/��F��~-C�&6�]�3#�3[=W~#��El/�����}kvѓ �Mi�Ӷz��4ݩ>L�\�d�� M��Cǈ�x�Vq�ʹw�9�M&�"��:���'Q�.�L�a�)9�L�$�1$�	#[S���&�̀e�`��0z��������}�#y[4m�U��V�L�S������r|I�	{_U�a˸;�9�	�HI�N�.:��F�i�
���T���~�q!��I��g�53 a,��|�QlKTW�C���g�R���_].��Ύ�v��7"�E��w_�nE7��DC&� ����i�Lc��!|䡅S3���UclD�)��"?O�7��88��R��QƐCM�ƂC��;[��������5��Iڔ@�{~��%i����Y�BT��p0�8��rF$Qf�\{�;��;E#H�ݫ��3�ϥ��A�]��}�W-�~+�o/�����X�t5���:��)��][8��Bl���APYo���>#�@��5.Pp�����L��d��p���Sq���)@f�N�T �/	���F��D牸�pʭ��8�My�_�o8�D
�)fOa��2 �2�)u���	 ��](Y�dU�ӆ�`U��F4��Yb���쳣��,�3���jifp�XV��2_��X��4t~�K�	�U���&�f�^n��1tZD��g����՛�u8h3����P���a\1�m��p�!���P|4|�
	b�a^̞�7d���E<ve5�S*��?Yw`4����S�B�񕆹Zض�?�7�r�Wھ��>���N��W8������i
HT�-wE+/�gɇ�]�.mE6N��B��h�s��K�}Ds6R+*�����=IԂyW�=������ rN�P�WA�e���#)��u;~(!LxC�2�yy�@���Km��9�5�P�1�G������x7������h�pd�gV(�A�xJ~�p�~I!9iBA����=��W'���� ��ƫ�H\a�%o��t�H�dѾ�����1�>Z
IJ(����Ƥ�i8��F�5��P�����	��o��I����Z&x|�q@�I �Q	�aO;|Uo[֭un"�=�X��5c���kCd��`fs=ƽV��z@C�-�n��<���Fy�O���~]>�/
���ҤƼ���v	�rc�G�!�*@w�{>�$��S��^��Ҽ��Vެ��=�§�ޠ��2;T�s��6�&K>4gD7����@Sڕֽ��)�O<~��j��u�,5?߱Qk2��Q�����:��/�@�ّc�?�/��X=d{�!�	s�uQ���ښ9\p:�����M�D�f��g3�t)�4�:vOKީw�Ӝ�Li�-e�΍v%dƂ��π����P�hm��k�O��͙L��+o�����U�$�ñn0U�)ił��6"����ج�����#�;�^ar���P�b�`�/Ӂ�#�:^ɘ�����̩Y�rp�f2��e�4È�ܓ�J_g��3Ք9o~��Xd�u�j�^(�����'c��3��^h6h���0�8O�:�&@X)�;h"�n���ڟr��s��.��r^z̑�/������R^D|��j8WZ�Z�{C��5{]$G``Ƌr��>�|K����b�����'=���em�MnP�6�DR�R�U��o�}����Ad�F`#_�7^��Ϣ���g�m�eQ�i���'���h�e���=�����8le ��<��ǳ��ʀ_K�;���&��o�NS�פ�ّґߣ�G;b�6'=�7K��~�ӷ�`$�k>o�d~۝��^�,m��@�o ����=�*�!�-"�X~mEHn�>P��2�~	���h��U	B�XA{�V�ڪ�GޒhV�t�X�K�DzR�H("��r�Fc�F�����Q�G�	��������(V�h�0(�`)��l(���Y�Q�H��ɋ8�sE[Y���ȱ�v(����������+���V�A�H	��A�E��'}^����X_]�IGx�Մ̓����E��|F��һ'�8�.+۴���g|��&�
�����|��I��$�x2hqqNqܐ��[8�!Ul��V	�{ζE��d	uA�e�U�[��Łg@DԜ �z���I�6�<�F��Q�tbi�W�3���)�2"�p,�c\s��>�֯�I�(��;z0E�!����v�a7]�b�J�fIR.�~�7&'��X���0���4�%ieSB��-��=I�������a�-X6�`��A�,2�/R�[�;6/� � �P���Z��ů���Ut�)$]�Z+��+��9�yFY!�IDذqƈ��D�2��w���a���&���gk+��`�P��Kl�>l*x�b�Cc�t��ǉ)�F7�2ir�e�-�Ali��p�����M&���>g�_&�.��7ܝQ�-sB����A��m�Yy��W�v�8}�	�9?�����꺜��`9�
����*o�f����W�����tD��.n7=�)�©�T��<�Tb������nR�坫�ȹÄ\"X�N����ٌ��w�R'R�HZ�m6�r2�XDU=+��l��L&�|��A0��5�-\[UY���!�8���.�Y��Vs������me��K��zv�c�_ ����*㐢ga4J1�Q��+�;�AT̾�w��,��fs��7ќ;y��3����9Z-+��%��D�^O�@Y��!z�F�|o@-���3R&�K��
��_=��&#�}�Ax[]8�"�fC۔�0?�~&J2<"M�wt�:f�({6< p��~{���7Q����R~"�u3����9���%�%n&x$�M��-Z�x���!�vq�X.�-����s��'�������d8B�w���务2�108�S"��P�����ws�s���� ��RM �ç��?( �,����rY�]�e�WN46�CNm���M�����t��}p7a�����8��J#D�(
$��}�PX$Q ���ٖ��9e�<�Ҍ܆y�+�� D&~0�[I\�ԶP�Km��wJ�"Z��ޭ�3�v*Q����g���	0mM˃w=�6�un���TP�3[#��x��Ky�$u�Z�����+Y�,��r�9�>��K���ƪ��◜���޷m����L��*]��?���!N��o�#��Є/̙�4Ԣ��əi��w/�����3�)��j��w:tc�Ѕ����8&�KF���,�8��o-�'�S|T��G�^>L�o�n���C�c\�gJ��=.�R���%K���E��o񮉎��nu�/��<lx"��Y�����"�jf��j%�魻贯���8��S=VƉGCz�Vi1��@w���u��د�����X�-���
�||��o�{�30�?�t�b���S-��y�c�&�Q&�|xz���[2}j0ߥ�{9� ��o6ƕ�H�z���BChRZ��t�L]�f�jc��#lǨ��ڨť]HO`�$*��u��ѝ�|4���S�]{���c���|� ۬�J��]��������,EH������L����Q����ᥥ�)S�Ė��Q]���8��ٳbvJ��Q�� 'Ru&���R;cx�!���yz����L�Y�L�`K�VB�hN���P�4�zKc�Y�h��5׀�P��/����#���>'O�L�������7Ty���u��X����*�Ɩ�d�b���@��xy�MF�OK8��1�q2h	]���k1��j`�Ӣ�O����{{���d�@[.6�t����x�٧<���Q��-�,޶�cga��FR�~!O=kl��3	a;����}�b�m�?�㞉�9L�ݔ+C*�!�G�����^0���4!)
A'xK�ǿJC��`{�	5mv»]$�WK��r� �,�F��N�3í�g��o
����i b;m��:T�P��ǅx��M�Z6$o.�eU�vC�K<W�.j��u#�H��k]z�C	�S���+,[n}v�2���&��S"�P��.Ob$�Z}�a�F��e�n�E���A젣^F4�	�&�(�Y+��bP��
&J���}����.8� �I@�B��oA��Q��T<�{��`%7 ʱјza$���ʚ�b����c��P_���Z�:�SV?��&P:F�7l�>�� �5p�"ۉ�&y�/�����)H����nF�<�3�����1���H����M�t�(�a��#��o�AI�r��`֩�I�I���5�O���E|�#��rB�~�T}	�v��E~bU}���Oc��d�>�,i��Q�:.��.��/d�H5ց�:�! c���w��(\4<AUk��!`Mb�|#�EM"Y�۬��vBR�%q��K5�I&��hS��G���K`h[��Ŕ�^	N�0�X��=���a��z0���_�T.��&Ɩzy@��������T�4�'˒���_��9BM+Mt��Q(d-�$����3X�<�j��I�Ih@�8��<�֡J��՟��-᫛��d�v�G�0)}����)S��kQx)"& <��nDr��ܯF���V�>ў���{��
jy!�Aӿ-�M1��&��d�T����Φ	��>��~1�J�pp[��)iɧ���d0iK������XYkB�6�鮾��ٙ�Ҟj/��8�7�xg<x*��߅#�-��5��Ww	��7����y�m�T)��a0lY��)Q��M�cjФ�g���o?"��)l�	�NցZǈ곩�S� �w���t�5(�l%f1�Bil5��K�&�Xc��`W�'��%�NM�@����r��3�d���VX������UlKC�D�?|�7��o�K7�6��v���w����aj�;+cR��߉m2��ؔ�n.�Ee�(ٱ,ѥ$~PU�k�2��?/c�u��Թ���3z�g��S����q�'TD:�%��
���Z�u������
�r�H�Z������`�f�4W���N��Y��?ޣ*��	�ED*�^Dި�4��-� 8S=7��gV;=��!��@��ZCa-�z�[���ZG�
�:�	h�����f����?��M��F�8�S����vV�����y:)%���'S���^�O�ρd:;�ͳkS�ٺr7�N�c���/ �v�o����$��YV��'�k#����� ��b�����厊��+d���j{�:���ݱ�CqN��c���F��|Ɔ0���F�|1�Ԇ7�s/Li�5����k%hXZǓ�a
t3+?P �s�f{NADV���,�2	���m�
���.� J�v�֐Q��#Y]���9":��.�X��6]�p�I��'2�mcNN�,^�a��r(?�&2E�FQ��$xܯH�	����HPgj��MU���h)i�Ӛ5ɩw@(lX�)���N> ���ި�{�,��l^��,�@i����
�e�
��4���o�������a��\�[��ѵ+���rk5h R����~glm���xvV<7���
���iT8h�ܳ�G
,[{�R��(5�_��ݱ|B�C�����El�2*�_�7��&�L�"���v��#L�I!/�I�w �+�SK���X^�MP�[.;0�(������3��C%�{��U����ł4��Ģ�����?�R)�eK2�#��\Ŭ�Ҏt[#>�O ����7�m�l��@���Oe4s`�uS�̯duDU=r�Tߥ�{s�g�pZ�~�l�Ow�a��!e�&���w�z�J@Z͙J؇�@�[�`"�B��)��4�e����A ��,��3kX��%{��J4�k9ܳ.l/ 5��N��o�*�������}��!���%Ή��uj�W��^b�Hՙ� ݕ3�9�^ИU(��H`��u�qg��"�{����W��|g�<��7�u���,��/��߅Y�n�y�~&�x�H�CE��_N��<��6鐯��k8���-� �2���#=�f���5���c[����`���H�����9�gN����/�%uw2/Ӻ-S�*�ƝM���3n6��-�T�}"7<��f�����Bshn�� &��2��:�ǋ�@����.9Gst6ˆ~�LQ����>w���f�����B�m(:��a�-���4��5�H���Iڨ��5�7z�r���޷�;ᅳ��+D���ne�_4���[@�u��� ٧���o�4o��A�C|�^�D=�d��鎿�%�I����~v7�L����ݽ�0F��!�h�����
Ih�^���|�J= f;��������u@��z�tr,V?�7�q�����d�+n�B8���~��`N����v7Q�u�X�l���z���&Egm�r��b�[BY[�?xcɄK����;J���ٛx�s����;:Fi���\7�;Y�ّ"ee9��'�pkl��:�p�;��D�9���#VB>��`����J���׎c�V�/�l��.D������N�����\f���_�-�(����?^�;�AsM�V�f,�{�8?=�d=�т�� �9�*�e�4�%u�Aҋ���ɣ��<��h�5zMm��:Y]�С�s��s)���O�mx����z����`>6RX�򙝲�,�c7-M��(�\bh+�B���[��FJ�Ї��,ղ�NZMp,ѢXh�>��ө!T��T�����	���:�<�ݞ���s��i�$c1E�$^������%����W�q#��e�bl�*������-E ·����2ȈR�v�y���o����Bd�����e�6`))A� ��4��S�Xp0�GS,;+(��9�� o��� Fe3����|�߰��w�?�"�<�h�Ǜ��E�@����v"��`�)(�����\��$����o���;W����� �ɏ��ظ��(J�|��<��h?j(U�(0������� �_	�h6p�f� k�)�^NXxM�d�EY�B-�v�<��֙Sm�R�䢾Q�&p�q#���y.�4���̃,�A}��C��|�$������i8R��jwv)H������cu&2s��H�;�h�:<4sg�<�k��`�n�`�o�����Z2%1S#�����$W�,<.��Fs�����	X�=f�4d���%+���8���Ԙ���:�OlO�}~�f��}��d��D�x��;]�}uJ�i�v|�?�">肎�ό��p�g�g�)�Y�)o@���n�T���DO��! ��4���e�	\p��F�)FzEp��`��;��.I8׉Ёz����-�WW�@`a���j���3��]�Zx�5���u+���8h�,�n���eI+Qڋ9k,����
�~�٥N&�.I�!��鸚XVR��!\��� &#J�.�x��o���W�U�`�1��\��+p�2�F��O�܄&�O�v�>�-]b�<]��	�<�:�t�Q��.�S�G��u��ttj^[A[���q�1�[�{�zP���"��(¡T����\%�_�Ŀ|�x�(�ܴL^��.����Bmy��.�ϛh누��vQ�b�p����g���a�O�KZ^w�%�V�mY����gH�8_��/��RM+o�hL�u�"ʀ��nJ�U�ʴ�,eA��"7�'={d�/P�� ڠYl���'�L����ܒ��H�do����I:����-��U g���t>�����F��į�ޒ�����N�+�@b� 	�~���b�GG��'f!{h��zf�Z6>�L�F"��R� v�*Z�)Đ:®�{�F�� 7s��I�%}�no���E=������l�aZ��Ob.�����Z.�w� Jp�6������)ڵf��-�
$��-ۡ�n&ǹ�,2s >{�;j�qb�W�6DS|[.zޛ��	���
��G[��X�$kd�R�9By=�;a4}9�����aT �y�̕�w^g�;��e��[���T�B=�X`Mx"c�a�_��}�oB2eF5��VWN��{���م����xF���k��"�U�t4�v0j��"Hĳ[d��F�� ��w��sR.�O�+M���y�Y��4��(�ڗ?�Q�G��%�]�/T�E�J� ���+�4[P�$Zeuv���q���)��)tĭ�(w8O
,��F��|�p�UCԞ-���+E$$��a����h�	h�sM��%9�`��t��mF˰���\s��T�b�Z;̊�Jc��ͩ�%c�T��*�8����R�2U��-��s�����/p�6���NL��|��S�"�F$|Z�V�U���S��]r���/|x�0�B=�v
�􍅯3TP%	�`ފ��$������p��j�@$|�Q�'�ĠW� #�6�����n�
��e��!݃B'��l����^��А���G�i9�35�h={��������C�!���6��B�A�X�fNH�bRa-�K�b0u���a\>�	]�?�]�>S���Q�3Ѕ�9�7�S�ij�Q����mu�t�g��q���!�A��u�!Ul�Y����Ԉ����]��s�]zr�1G���3��l�^[Ei�<��0(�eٺO���k��*l��h��y%%*T�h���h�<�:���p�F]�hx�Q�Tv(_~~4�RM|�c����$��J*�*XK6aJ���Ρ��ଡ{B��mĆ+%ݏ%�wq�>A34���
�`��&P眿�d� �2�?��t���~U&����7m�0�r���~�H=�vP:~Oe���d��5���~_I����:S���]�m� ��b���y��f�^�	�b�7���n�Fy�'�Z��3�B� ��q�?��}�4Dew���8Ƽ_������%�ᰁ��wzS@�b�h�YS5a�{1Ak�C�~ǉ܍⑛�s��Oe�0Ng|V8˯WBf��+�;�������\`߻8��;�Q��v	#���`��ן�$e�{��G�2� �'Cc����\3o� ʦ���YC���d���_\���o�;&m1��$�y/�����D0�_Q �9�d,�I��M���#��%�~��f�_6����,�XA�I�FM8v|�(YX��-hZ�h��\bN�4l�t9X��C�%�}��> D	�~��E@$*�9���5�Ls�l�����1Qg�w'x�kF��I@���#*营5����Fk_�(��l�b���n�� D;�
�(�ݨ�Wc�j$!,2����Ũo�=���@�-S�긍�C���'��ӯ����\Evl��i�W���u%��]�	�E�v�M��g\��鼹'�XE�����@����;�堟��
j�oT�n�ڍ����0�@J_�g��=�;CĠ{�3ʞ���(S��եQ�u7.&Ӓ-H�n���C�����4��]t<jҖ��8�A� 2~}:m]�;���S�,_���y�..w����aw}O�Eń�qhCG�qpf�"cf}1�ɿ��)0BF��-��*8��C�$>ҥ�ܫ�{4(��@+vV�P�i���O6|Į�;%�Z!��
�U�#�U��<�^pq闵e�לhfL�q����Y08�S#��#�q��J���G��i�W��ʭ.OG_��
�F�f�J6)����"��QGMl� C���F�|Q�f�5��S!�g"��ȗ�	�@�k��o���oDx>�����X�S�DaB�Z��)�2E��*�����c�̓f�
>�U���ԣj�\�b���4�nס?�C֫_Joc��D8�Ow����֤hH@K5��� J!����PR5�@�X��+��l�����Ԣ�~��O�H�92A;���ѝǍH4І�+�r�(�ւXZ}�QqX�~c�O�^�6m��_���W��%c�`R��;Ȼ�!�?�î�;��24=��o=��*�2�i�=I��_q#O�_H&?���1�3�F��������26��[.x��X�-ۙ�wX0�.�H����;����?d�m�괠��6����/<E�',R�[�*V��I�fBMk�L�Q���iR����+� �<�r�tH�ɋ,H�'_h\N�zm�(�Z%��R���OAl�1���YQ���ĳ�j`vp��n}�~up���T�D���.pW' n�q�/����=�������e�	X���F�r��ߺP~��z>7����zJS(��K�";5A��#Ek���McǍ�-�\Qd����G~�[z欻)Z��s�a��A�@�o.Q`##|�����_�F��c(3�p���#��X�܌tՄ�jYb��^��x����2�����r�ڢZ�Q�r^�YnY�Z�م�v�#>\+�kbl� 1��F���W����P��%�弰�|
^�`�.9d�&(!�à�j_���	���(��v�_��'{�D���J=��T֡���>�����$^Ҟ��-�3�b3�K�N�A����>8�b��	N�{�qDU�3�pP/b�Ua��be���L�;<���y����Z����_1��k�2�T��)[�P!��"���ʀ!�l�{�4���'�0_�٣;0J�W���`z,�c������+J^
�z<�c�Wd^g�����Đ`7��9��_��������X� �����=k��C+��Q����ϧX���w��܇�#vW��ҭ��̄�Ku�4�'>+���m����U�N���N������4�UjIb^	�d��k:T��m���%C�!��W��G6B,��֎��.���;aU"��)���do��Vf�%{6��==�c�/��J��f�Gw��ݼq3h�� ���r�ŕCw��q���~Ėr܈����Z����`�c~��*M���9з��X���J��S�k:�Ob]��]����m��lx[�@F�K�a�b�(�C�{�r�P*~�\ֈt�x�F��ߵc�`�mβ��!�0�x9�+�H�%�	���Ky�*A?���+�U¤�6��{�:,j��Lj+oP˞E�8�rZ�H	Yt��T�s=����	/ߡ����5H�_�o�"kޤ���ƒ��hq`��5�r�fwEk�t�[%�����U�,O�>����&�(��R���ԕݛ4
��FD��� ~a�`��z�]y!Y(�"��N�ɫ��b��Jx���>N���z�7�ve`�W_�Ӿ�Z��#��X6�+��k��w��eCԧ>��Ȯ��1G���x�`
��!	BM&���������J�`w��g��:U�-��{�Ҿ�rv�`v2v�5�FG��OFC��,��3�`�o,]�H�+q�[��62��j���>�)��f~������������[��������!zE�����|���Mo@^���mK���F���>�^�_\�D�m��u�#k�$'H�k�E��i���b��/)�����3�O��`넓��BL������*����afW�w��8��${:�X{Զq T2x�-�l l�u	�k�\�W��Pɝ(�5`(�S�c6	Q�0��b���H�?�s����p�����6������z-n�6ñ�=6���J0ȏ�Cx$��������5��)�فvz��+���b?�8��j�*?�w�e��)���\r[����Y��o��@X;e݇����g%JD�K����
���X�I��޺��@�p�͵V�q� j�~�	Ȓ��EHk�@�W���8�+�T�Y�nΠW��@Lu��oo�Z�-� ��Q\a0���P6��|ux����(��L�+<���}���:�i� />:����5N^2J���R�O�����'�#��q��P�Ț̢�寀�CT�Wòȥ�U�3-#(�D�E�m?O7}�T�x�ͫp����*�:�ŚU]t�p�O6�����E��b���\�ǃ�˫��xE9ś����t�!��/�xM��ܧ�1�z������U�pO^T'�,�;u�L
uZ��
�8�#fu�T�t�$Uy_�2��Q@�~�ƃ	�|��O�T\��M?;�XG��K����d��)B��BB�]yصJ˺:�'J�ĉ�d�����5#O�����(c�NR�Ŋ�GbR�g���� �~�wE�*���%:��x�
J(X_��
��۞ �F��~:7d�t���r��~��s?���5��l��v�CV��L�xN�5�ױ�^�z%�ȨȀ�U'�~�?Őr���R?~��Dx=�)����$)�'?Ʀ�e���K�0a�O�����S��D��2��Y�3D����bWJV���cw�K�5�O��$mrY�ܟ�;�yy�{E��o�Y�?�1�O��~'�?�eZQ���$n���oC��H�e�^e�]��0�����f�C�.FK���%�|���=�^�u���#I4�����8r���5���Jj�	��K! +����L� U����31�P�u@����\��sN%}��nAʩ���ql����ƈչ][e9��<�ƫ��Ʈ�h闵ݍ[�(fv�����o�ê��L������h�p�}�_[��2f�z׹�s�B&��1�4N?�ߚ��e͏Ê��_	���� �����Eaxg�ߞU�\����A�UɎк��:6fAF��!,M��}h==Ԣ�7�KX�n���#���ة��|���Wf�f�#.�2n����Y3�ӈ��is�t�`@���/	L{�YJ���?�Z�zH��� �
ژ��u���.t���:F����.`� Y�t���7`�"���.a�ey�s�H�:�7�%��T����P�;������<Z�q��O�����I�����RTt���<W�pYzbP�^�(
��I�j�����,2��'q����:s�ڧn��,�g!�pi�j<�����4����S�nS��A�'v�
���:�V���կ�!��'<��U���7��\X�O�ho�7��]��R�&4z��6.�c[q]i�0�=�Z#�M�����$�5!-����=�x�Y9��XRyݭ�#��^S��N�ϭP.���xguB[r�����9鹎jv2�u�o�����xZ�8
��i�)��2���2���A0Z"�_�-pZ��z��z�dFwC�S(�Ix��~�=�@$��5���m��2� J�e�-��0�u=����<(����cM>�=���*2��j��xҙ%z�X�L�$��@�����x�������۹3̏�燫<"�C*�$s���y%'Z������~��J���O$��Q���>.��,A?_�ɄM���Z˯��Z<���vT��\bO\�����M�'�FM"nE7._��)�ʼHܡ%�.��E��ݒ��m"jQ�kܨs��yU��;Y���D�k����f27I����aT�X�c��Q�oâ��7���RG ��G	?l~�_;��{#+��3�	"�u��1?\��Y$,�:���`"�&�
Yֳ*[���[`�&�~zFb����ɹ�NL@�߬��ZA��L����1�BM�!߮�MHY6���7���k�k&�8
�(��=�8'h�E@�y�Jͱ���������U\�U��eb{�@�D)�¿_9���':/�2�������-'tn�W4�ᱠV�g�&��J�Ƕچ���t�>�*zGD+����=Q��#�8l�l�9��*@7Pt5���$�ZX��<򘞃�ҧ�2E�ŠT��ht��q	�t�\��v�e���Ma�W��B�VΠ� 
� �iBt�-M�25�y?{�}���CB!� ��̶'`��3Ԩ�C �$��?�cؐ���Z��Oi1�V���X�# .&0��xj;�+��
cM|	;�bNH��g����dB����]���F1�i��w6K�����k�� ,`C��q��j��_"獷J�c]��z�r緁��;�{�E������	z�����;�0E��t�`����?�W�b ���1�]�=K]x�G�y��Vj��B�W*�~<1�9�����:�&����9v����r���G�+��wkD뱕�R�ق��c���|/<t�4��.0�?�H5~M�Nk�@�_�?vU����J��Я� �ݪ?L&o���\��*�](�J�����~�<��y	�0e	�˒�ɓ_6��ల ڒ\�>R�wͲ��x�s#�����)�G��o5
��V���H���9�@n�$ԟ��|�$s5�|��3�������&����}�WO�g�Y�1��ֽ~�F�?d\˯��g83,ب���_~�uԥ�ȋGb�$%��'���u���x�Pn1
g@��&
)k&���[J�23�����}8�#��}�V��Z��?O{~������e�DD�ŉݪٕ�o�`�m��Ô�
�f;l&�)T��V�&��ih܇����𥉉>�0����k���	\~����5������O޿YV��>���}$x�_��&�[��,_WQ��0���Lv��qU���W
]6����;��6f�=2�q�Ի��/{�T����6b��/p
K��aJ��?�f!�WS{��|�hI�lR`��+g�G�"|q��s�1G��[�2w��"�[k��Rc�K�O����.^�.�m]��פ�r;[5��Kѝ �ɹ�,[���ײ�as58�l�������ڪ=��đ� ~ۗ�"X��4|��h]���@H��׼�K��-���<��=Y���̈́�I�P}Z(�j/N
�%Vk`h>������ʁ=��./�r�N琍?��hW�%2\r��B� �V^ݒ�s��w��y���%��^<Y��U�=�d��j��x��Ȗ�MFrB���������K�CS߭[ڮ�
Os�;�W=�/�ǽ�s�k]�%k��\e$��]�P�^��wn�e�S�~6vF\"�J�n�(��o�� �h.�X��/�W��^+�i5���<�28�e�$�<TN���Y���0�O<>8*dl�ۦ#W�GIJ�v(A�A~\o!gC4�r���&�ssawO���YC�tg�����lr�7n{�C	��@��q�'���\0�;�ߊ��б�._߬����')�̵DV�M����좊�+e��X�NXʝC���y��s�`X/�_s��^e�l��1灄��2��Z�H�g t	�G�����ޢ��Y�X���-nC=���fk.�#�f�, Q֖���V���PP         lP PP XP         wP XP `P         �P `P                     �P     �P     �P �P     USER32.DLL COMCTL32.DLL KERNEL32.dll   MessageBoxA   InitCommonControls   LoadLibraryA   GetProcAddress �h`�    �$���+� �K��,$��F �t�uǁs�z�/�sw C���k�  ����� �hr�]3�A��������   �Z������� ������N@ �B<��N@ �w�rs��$��   �s��r���r�r�h��$��4$�A�����   ���� �$�;�Yڋ���N@ S���L@ ��������i�Y8ڋ;���O@ �[����O@ �    Xhh�e�w�/�5s�/���؁,7���d$��%�!   ��  ���O@ O��������i09��I������+�,$�$�$$PR�y��DM#��d$��( /@ �D$ZX�d$�d$�������   hX�H��  u��p�h��!�@��@ ��2h�   Y��~a@ �   ����h�$Í�9I��   ������$ã�,$�$�$$PR�a��DM#��d$��(�/@ �D$ZX�d$�d$��� �   �Z���tV �T ��+����   h�   �4(�   3���   +ɀ�%��6�F����H#�I���� ���,$�$�$$PR��Rvଉ��d$��(70@ �D$ZX�d$�d$���ݠ-�p��E��s���x���ᣰ���xP����C���}�hj  Y��r�봇e��0GI��,$���$�$$PR�%���-p����d$��(�0@ �D$ZX�d$�d$�&�F���H�и�0x+Ƀ�����   ���N@ �ֹ   ���t�N����    Y��   RQ��#����O@ ��?
  ����O@ QP��n�E -p� �����  ���H@ +�+���A2�H(D9����  u���t�@ ^��������
   �    H@th�   �X[Q���2�c�Y\�   %�X�   �h���$�ٍ��W@ P�,$�   X���1@ S���   ��tCu�R)��,}!����|J%�����H)���h=By\��{��mm;��1� �_x8g:���M	o�c�]W6���������Y;]�X��dk��u$��1Y�V��Rb>��De��������ɃQ��
�FL��P���fC3�b��������۳Y���A�ܖ)NY�
�|�Z�X����c��mt��x	cJ�#�^��%S) �+>3�l6�r��]�����<t�w���;ܸ�1�!�-T�`��<�F[����m�nL)�Ђt��2�}�X��|K����W�9�T���Z-ݤh.�cW�>pǄ�̙����&�[�O0�f��O�� \M�Z\��8�"���*~*\�1���A�,6d�����i(w��d6��.�E�6�Yg�B�d�8v����ea$��5�+�ف�-sd�'P�]�	?2#�5_=��Q�3��.� {��[����P��v�3m�J����:���Ճ�|U��X��]���a�Y��Q����"$g�]�@�D����~s�\.,_��'AXl}����R+�&߇�ϡ\وEs_�0�0Զ[ ���r�R)��@����CT�׮�ҬǺ�:>����f�6��B8�p�W��_c��3%�i�@K��_!H�p��u�^�V�����3hI0"�/R��(R��u$`���B���x�B��`�q��q��%)XPk�Y�`G��M��'�=(�ʣ��$�NsO����`B�JLW9�(%Y&�}���	�J�;Yo�[S�g�t��]G�h8E$w���x/Gm�%{čC�o�B;�&���2-$�-�����<6�C��O��e�y�I��2aZ����q3Z�@x#ִo����Q���~�g=���1zH�H$�n����F"��%j���歔�
!���
��u�Ǧe��bW9�2
k�"D��N^J�S���OX��/�.I�k��ۙ�͗!�oBY�A`��Rx�֏	��庀�����a������j2���k��VV�cn@�=l�Y!� a�ٶ9�������-	����}�,v��B��=�f�l��\}�Y,1��@K��u�/�q[��k����3�L��	'pV@s:�#���j+;�E*���~�(\�^��yI����2��G-�K���fo|Q�
��h�@�d�f�.�F�.C �-���}�PBm��[bc�AOJ���L�@7�ɜ�n|�m�����WD������[;x	59A�
���l���g��'��z���3xAY�N��ȇ.?�����g���V�i�[tLҋ9�RtC�7M�W�qHjt�ġT(��1��,(\{�E���W�Ce�9�����������y��6��(�4@b{��j��ڞ"�`��	��f+_ `5f�������d/i 2�`2ꏻ[�$u8���-9G����+G�s��Ы���?��W[c�J����ئ$ԩU�ɚ"��Nb���
�������]�+AfS�j��B�B��|�دu[�GU�e'�ڷ~Щ�sN�fC�6����;t$K�(������
wdU"�a4{d�Sl�l����wrm=*k_r�={�*��gJ��� G�
��~�U%چ�e4p1ك���%���m��N���L��2�~sX�#�z�A��t��ý���j��G�L[�H�� ��_�j(I�� �Mld�
�F�-.m�`?�.:0c�L��|vիC�4���W�"S2s,�������$����:�4�CP���Y8zQ��)>vh�F�}J4f����U�nd�y��d�޲1�p�sE�n�����L,*.���P\0X� 3yQ����4G�C��I�߿e��dy8ɶ�C����i����U]W(�����z�[�8�6�2ۢ$e��.b��;�.Y��QÒ�G��@:v�6͔@g�9�q^���bk�K��\����o�ܔ6��N�a<�0� ��*:t�6�1QlОYcw^`���$Z±8��6�"G ��Ь+��)5�W���{�L1���ݳoW16��ay�PmjG�ѥ�by��� �IW���`���\��� 9��(��G[&�'<���Ba��q	|��&�4=����V��[UU\�?�2�#d��������4�<0"���Sc��R��y��㸑9��m����I�k+����7��^�B�=l��L�6��F9	�����Ĵ�}�k�(f�C#DѨ�1I�U`�l.�4v
�?�eꋞ�DE��o�x�2E�<�1Y����y�ȑ�����@S�{��y)�^�#5�� ��.�|�1�_��w)e����u����H]��w���fd��.ܣ�����������ʿO��R��Eͮ�$φƽ�|�P���o�	jv���bUP� �*�?5�-[Ud�^�x	����0_��:�@�$�z�"����n�zm[��Ip%�D��x�`a�
�݋�Ă�=��`Q�p_�(�_�y��"�̅��f�
v�#>��W@�S2؆�J!��b���?v�	9�7=Y�t�DY��X3r�!�/�Ie�3n��|���8g��d�$�2V����E���X��O�ً̨�}�B��Yc���(b�Z0������ݛ���)�S�~�Y��UC����ͳw֠rWk�5g3B�q|
���hm�}�I��uZ�x�jIզy��j/�I��+���=�kE���z�%�0�R��ϭ�X~�L�7�R7�&��n���U���Ρ�(���Z�T�V�. ��/�X�����s{��Έ�gR�3�ee"���7�+���ߗ�-w.��Ӈ�7�Ϡ<�u�v���0
bN�D�7�nJ&FF���i	J&}+yvd�8�4D1X���;B0�pӋZTy!���bEng����<ۭ�����[��]�S�MW��!��m�|7���\�+	�	l�� 7�I�D5�& �T>�_&����gl��#t��1�`����B��|��m�a
<O$�����K]�Φ������~�wK�I�`~�Q߇������Io��%��:�&��ۮ�?!��n1R���F�%����(��~XcԕV�9H���~�z�m����Wbp|wf����L��s��0>9r�2�aÖ�? ���x�]�Oc�"p�:��w[�M���ֽ�80?�i�1�}x'��.g�x�2#�V�Z
��� G@ ��~��e���s,M_�jz���Ā�О��S4:�`��t5��L���~���!P�ښ��{PYt :z	�Z�ERkL����h��<rŴ��

"�*��W��9(W�7�A�E��l�7=_'M5�t!���C�b�ɡ�V\)6m�R4���q�|�fh�G��Y���:b8��D7�Ō��O��l�.%�4������C�S˨��°6�E	����<����d��b��nyB$y��[��J`��K[׆��m����z�P�ΎB"GnkF��UOC��*��D�tM�ps�OO����d�K�xM58~�^�Lȼ68�Q���t�J]�4����Q=�c_N��uu�y�����T��]�)��x~�nTfo�yt�dX���C#�zV-~�!f	�9v�2l�si���}Bs��wU�T����/ԯH�qV+.�`Y���oTW	�L�2���q���7�|=��%R�𬣬\ N�:`G�L6�L�iM~��I7���H�bo���O���a�̺�c�����A?ӋOٿ�r�X4(w^�c��=2���WP!}��퇬p��k��������h���#�ت��4��$����S���� C�(�����l��rH��5)���r�ط�`5�^�p70���v���c?�{ 	�C ۗ���+�)��"�Yl���AYWx#Ms�I�v�O�[��f8.x'�Ϧε��ŵ�Oi�b$�| !��;D��O`E�9ԫ}�QDG��m1
��$_���{G8lX��$ߏ��P��it�dH}n�oy|B����lK���i��zc�ܻ��.}[0:��+Gt���U�?.d�"7�7�'��:���o�����bJ1���Q����Z�y��G]�@R-�,��>Xu3�o}�&�3��ܳ6�-S�J��&rp��aﾩ�i�@�P�v�-l�s����u��4[��ܚROP��ҙ��R͆�"FF^PYߦ���OND�X����K���Ω(������y��~4�9���ᥫt%���3�\���KL�ܽVC�������ڙ=ᆤ:�/ž��)�3T���� BIɨ܀3L�p\J]y˜����m�5���'u�5-�gv�,���Kc�9gLB& ^�t�]�E�r�2���1U'	D �%9��
��L��>m�+�y�����X�J�J  hzL� &~T�h� 21{�S��E8*�pq����}��Sx�5�`*"-r��nc�K 
������fH���EjJT����1�e�-D���Չ�+�2Z�7L��+V�*	?eg����y�8�Y��]Նm�[>s��0��~)����ШC�Yp9�pl������T�1m�*�D�1kD������~����˚9iW��ռ?1�ѩ!��N#]�x�
}��5���bH����������2F<>y�?$��ֹG'�%vn�Ez�x�м19�=�ͷ �%�OSӵ�x��=����k�_�u|�Mx�{f�C^��"h�:WxgYNq�d@xw��d5�Lj̠,�.�6���x~�E�`����x��S�%�z�X�P0�;6������o��.,�<Js�U�ϓ�/�O	s�>Y}���D�eO^�b������*���[�fȂ���j�:SɸuC3�ly.��S�������tH�_��:���~���k�}-�
��%���1���I�u����d��Ю{�7�ߋVpjʒ��l1���+`��.,y��W����).�߉��$������D��A|� ����hy1E�(HFo��	4��, ȹ�O��S"�� �Ju$Y��6=���xѯ˨d���}�`,Gb�����)U�3ۚ��6�*G�yWi�k@,o�Ei4ݕ`ϦE��V�Ц@Q0`-���h��Xyn���i`����ID1�౏@Ǝi������>��P�X^Ω$���h��y���^�/��`8Fz��@�Q�S�`r!����9����y�]�D�X:�����.~q!����_	�����dX)�n�
c!��8є����t��f��s��N>lD֟��U���t}�,�ϱ���lv���*�c	 �-�O��|O��($�r�W;��D�챋aC�+�z��O����.	����e�����8ĳ�ͺ�N��}�Ok�5u'�x�����I��=G��7=�,���!�9�"`�C�IUf�H��H�!�������������c��娎���y���C�i�?*AS'�m��7Z��`����2��#T\��<v��2;�d�9O�fi���ȸ3�(��F�$f�Ϸ���Y��}K_��u4ߵ��$�ZY�>��|�K֔�|ۂA͛+A[9��e�|�M���p������Z`gp��_��/�!��N����=h$h&�:�=�w�:a��]��ܒn�r����nR^�0p�������>�H8X	�9�2�U�|=�W�7n�L��>�H�c��lvg�%��P�%bO`-G5��o��/�ymڗ��_�?�m�`��SrA!I�U9�oC�&L����ϲb�\�ͽ�H�W��M�P�����F)���7�첇\D ���۝%�+j�)��K�#QP��^X����rЊ�I������G   �h������������������������������������������������������������������������������������������������������������������������������|�}�x�y�t�u�p�q�l�m�h�i�d�e�`�a�\�]�X�Y�T�U�P�Q�L�M�H�I�D�E�@�A�<�=�}�9�4�5�0�1�,�-�(�)�$�%� �!������������	��� ��������������������������������j�QF��)�i#$=ж���Z�6F	���-����P&�M��qL����%�C��=��6��D���S����0X�CK�fK���cJ��	������U����=�y�������vy %ɷ=d���SI^�]=۾�V6܈��Q@L���H�E�ￚ�,O�S��=���B@9E�0����=qb9:�$��:K�\w���в\<���Y=�Y.�A5��Q1���R�r���L4� �0��g����6<��bhz�aV0i��E�A~���S:`�r��d�<ɂ�p�������[~��=�L�r��H��<�(hZXm�����������������������������������|�}�x�y�t�u�p�q�l�m�h�i�d�e�`�a�\�]�X�Y�T�U�P�Q�L�M�H�I�D�E�@�A�<�=�8�9�4�5�0�1�,�-�(�)�$�%� �!������������	��� ���������������������������������������������������������������������������������������������������������������Q��/M����=.�Er{���Ű���r��y?�pf�p6o~�G��H���}G����zH��ݵqG��J��ԩ�DQ�頺�Sp�z@��	g�h�[�/�. ^�D-�9T�A-�8R��} ���0/EWF��m���jX�������������ih   h~a@ ,$h�a@ ,$P���N@ ��h�   �h�������@�����$ h   Sh�a@ ,$P���N@ ������w�rs��$��   �s��r���r�r�h��$��4$Ë��0@ ��sj ���N@ ���,@ Wh�   Wj ��JO@ _���3�����\�GG���-@ ���W� tF����_�� h0   W���a@ Pj ���N@ ���N@ ��������ŉD$a�$h0   h�a@ $h�a@ $j Q�������w�rs�$��   ��s��r����r�r�h��$��4$Ë|$ ��  ���   �h����$�N�$k�!��i1�!f9u������:f�� �u;|:4t��   ����   �h����$��h�N@ P���N@ l$��A��덀����������Ѕ���,$�$$PR��<�����d$��(�/@ �D$ZX�d$�d$��%  @                                  ��*���q#cc i3h��rА��o�lOr��1�r"
�2e��Īa/���t潤t��yNeO��oeW1t�K�e��� rr@�Tt��Xt_@�e��S&e�&�Wt:N��tH�-t>Fa�t'4w�r���i^|Tin��'a�Q8i�h��r�y�     arB>�t ��6tj4RsFA��s�S�Be�-uVt�3Gt�'��a�i�d�d�     v0�y�+��&C����F�0�~ƿ4RHG��S����?"I��͢H˒q��K�$�)9�D����2�17�!4���n����bk���x���1�v��� p!Y ��v���[L�4K��e
Nד��M^��'�� �(&�8--.�7���du6�O8���m~?h��A/�H��H�����iP��)U ,�^]^_�a:� A�bKijk�iJ�����XCJ,�*�G�
J�C�s[:&���Ƃ9�Qq��kji��]w�\��#Z��Q��k����p�6>�����M�|��A w�������Fq��G�^�����ޚv6+�����O��dW���Vb��������f�e��莹�xN��u�K��b9��J�$�[=C� ��#(��ĕ����<@5�9�|=�����I��D��ʀ��JQ�Q˹W�����^P�(o�\`ab�`썜��nO`��(B��{�t�|��|���Qk�w�0dtC�keG�ny�K~�Ps�epd�t��WZ֭թQ*���nF�����AƧ\�#�V�V�J��7�</-+K���92���\Qa���2�DQ@���of6����*cn�ܮ��h���Yqx�@R��UG���|M_��@T��i��3����l��-��ڽ��}t5f��i{<���B��^I��,|Oa��d=��f�w^\]*s�c��`hieN45�~u��W[x/+�QZ��b��D�y�� ��8�ΏS�o.�ט�XL�B�]6D��ݮA�Ć|D�Y�s���S�E���T�>��Į�H4����B����YՂ��������	������솇���7�4��د����9�wjm[TH	R����]P�����<T2�"L��()*+��*�tΰ�$^�\2�<|��(�C� �D�ϸ�^O �~w2�Wk�>�l9��p&��5��Ak��6���B����87x��#& ��J}9�ǈ�c�����mzĖ�gq����u�)JYJ'���kV'.���74����=
u����6}B����>~����'�&$�9(�[R��ی����lW�����[�u��V!rx:�8���u�B�	
���w�'��T�I���P_ 
�� ��#��ъ�)./0�234o�%mk^�Y�(���Ժ�#�KɏD�
d��6w\1�T�ohijާ�bcd�Ydդ$+l�Bs��qstu�sђ���yZsCz�Ƈ1����r��Ie@�M��L��������ǧ*�M���6j���X��1����� �g�����,5���KC�����D��؋�^���(��&A#�&�#	���`1� ������O�H�|%���a����g��o������#�G�3��t�����@.C�*qv�gJ�U���6Sz
B'W>��fD�<O�<A��JT�X�V}��^��]��[Ê���%j�(e�o��j`��8}-V�� "�Z{h����vyf��[tn�M0�ђ[�Ֆ�ķ����۟���������©����=�����P�|U�"*�`/=�ȣˡϧΥй���U�(M���ܝ�����l��i��f1 �q���o��������e��LD_����o�ȏ�"%7U�Y���VU���%%&'�q�c3"��212F5��G;ѢS־�����DG�9J��|P�֬W��v]�Ҭ7"c��-1(iY�??<>"#��$��~79z�+�q��j����l�!ap���Rye��}r�Zq�v����\̢6��B�����1\e���;����T�����K�έ�-�ɢ��-��(���+����03���߽�������) �l秱�aù�������� ��8KE���
��
���{yE�XVZ�(U)|�)&O����/F�512j���x9��<>?��1EŶr�z�zTҎ|uT�@q�s|X
	�*�pd&.G��La��D�9/p�6W|/.�]~�Y��~�������Ju� U&�咡SW���sc��t����J�MO^�$���h���}:���d�fR˼:N�����x!̶�G.74�$��C�^���(��&�5�z
��g鲶ah�ذ�������CPꆧ/s��6�E�8JB��"+�7�12HK�r���jln�A/��Xtm.�4��7���ر}3fe�[dE�'`�ܸH��fb\NO��6�QUVWXh�ܲ_pab�YB=%��Jmba�������?Xy�3��	����~b�u��	���-�������v���&Օѩ'&������[��;3 :;����K@z�������5̍��*�>���
 ����`+���'��-��L��2x8'=e�����_�����}ܙPV���y9���¢,�f߭��0�$2�ש�K����;g� �تk��
�X�7����%�t�N)6BR�s���_GA��6�:��W�����1�j�:����'�������d�#�}�A�1�&�EV��g؜���ml'Қ�)��܌oԒ��O�kB˷��>,�X�d.�|�����RT��Gy��B�r���x��e�b]���]@`�ӯ�v��%�]�Jd
�W�1�Wd�\Q8�?*�.S��5(Jg���l4�dY��I�k�۽l��r[�Z�	U�����?jNpٛ���(!�� ���P&�#�Պv��|u����L��s��AW͹��<�oj�=yR� �iW\���v�ζ	W�o�����T�6py�~�xsbp�ڻ�*�.ܡ/ی�'�Z,G�s��MI<���iW�TT�>)�=.>��T	�'�
S;�-�_���S�W��T���`��  ��	
�~�\��+�����b�����������M�_��j!��S';Oª�
�m�Ēq03�F6�E	�9@�BN��EEF�KIJK�IԤ���WpY�ͰXZ[\�ޣJbcdghi3�h��k���rqwHyz*}-�%��Ä��y<~�̍O(����e3&�mW'Ō액Q����;���s��v�w}��'}���7��@��Ǘ�qK��?ˏUA�$���Z\�χ��W��鸻i������T����Fꮶ�]�� �������	
���TP��NV���{��$%&�I)*+F)F/ 12b^5eȝ7u{<2?����E�̗�lKLM��V��U��S���3�� aa֢>&g�B�fmnoʥ;ҏ�<t�;�|���k�{h|�E�H@�'�d�{y��~mxY���k���������2Y��	ȡXԕ�>0�B���3�����M���;��;gD�ru����\g3���$|Jc����T] ����[!���h+�D�����	���(�����>͚\=����<%�,qv�o�u#}H�ww�2�S�zr�;���[�Bo��F�/˥�N�ͥGp�zs^�~]���a i�Od��G�,2s�1R"!�Xy��}jÄ���H�6�sf��Q�Rt����q�X�~\%a��IYw�ݛ�G�E�O�i�?�=�S�P�3����>�5/��Db�P���R��Յ�od�"ٝ�����hb�ͷ��e��窩���	���vcNA�W9ԃ[r߆|�HRp��M\~��ز'�"�P4��AB��-�vhn44��{��;�,eJ�GEFG�Mà���Kt]��W��Ҙ-n.�Z��e�����v����KpqrY��������~�y�*��Qo�ll�wa�ufv�Soo��Aar�qw�`t�XI[���/S���Ǩ.A�I_�4O�m�lθB^��)����9�I
���ͦ���Ҋ?�L<�"1 ݷڷ���㵏�L䤬���|Gv���`s&C���������
�	*��*iij���#g7� !"�?�U�c)�n�)��0��0���Q
�q��6����RDEF���L��SQRS�QY��Y�_xQ�R��hcde��S6*kG�.00q�؟r��y������h�����y��������~�s[��dK⡤Eէ�B�TG�ADKY�JKJI_����W��T;�A����7)!�V&�$;*-^Q����Z�ۨ�6���⋼���m~����jp��m�{9�{�]@�7��ŀ��	�������qKpt. pH#۰(hh)�q�-./0��34u6aoі��¯���E�.GIJ��\R�U��S��^[�����#d�^gg�klm�/
prpvGxy+|��q���
l�ǈb�(�:^�ђB�טXc���$�����e�L�BA�6FUo�q����<µ�q���~��9{��/�54]&�$;��8/�%s�����^���~"�����i��쾽H�@/������s{(@cC�B# SR�h)
�t5���������`!���Ef'#�^&D-n/0`d̡&yw8�;�Y;���.fDk}�J���O'QQRSU����[Q����������������릕qΡ�������������P?
Y,72��7^X+%^Q$S!Ji43$(#4x*(?/��/y��
=(/r<�wv}��QLZU\K]XZ] GBP��riLZVa
!0wr`�ΦY|o&ym':Iqws-P?"5MwZipSO�У���ϒ���ډ���������צ���ʹ��� �Z��<f� �T����}.$##C��d��'p����J�!�z���3EǠ?�{n�(�A�Yj80�e+�W�5E�?��{n윲A��j8�0�e+�W�5E�?��{n윲A��j8�0�e+�	�r�?Q��{n윲A��j8�0�e+�W�5E�?��{n윲A��j8�0�e+�W�5E�?��{n윲A��j8�0�e+�W�5E�?��{n윲A��j8�0�e+�W�5E�?��{n윲A��j8�0�e+�W�5E�?��{n윲A��j8�0�e+�W�5E�?��{n윲A��j8�0�e+�W�5E�?��{n윲A��j8�0�e+�W�5E�?��{n윲A��j8�0�e+�W�5E�?��{n윲A��j8�0�e+�W�5E�?��{n윲A��j8�0�e+�W�5E�?��{n윲A��j8�0�e+�W�5E�?��{n윲A��j8�0�e+�W�5E�?��{n윲A��j8�0�e+�W�5E�?��{n윲A��j8�0�e+�W�5E�?��{n윲A��j8�0�e+�W�5E�?��{n윲A��j8�0�e+�W�5E�?��{n윲A��j8�0�e+�W�5E�?��{n윲A��j8�0�e+�W�5E�?��{n윲A��j8�0�e+�W�5E�?��{n윲A��j8�0�e+�W�5E�?��{n윲A��j8�0�e+�W�5E�?��{n윲A��j8�0�e+�W�5E�?��{n윲A��j8�0�e+�W�5E�?��{n윲A��j8�0�e+�W�5E�?��{n윲A��j8�0�e+�W�5E�?��{n윲A��j8�0�e+�W�5E�?��{n윲A��j8�0�e+�W�5E�?��{n윲A��j8�0�e+�W�5E�?��{n윲A��j8�0�e+�W�5E�?��{n윲A��j8�0�e+�W�5E�?��{n윲A��j8�0�e+�W�5E�?��{n윲A��j8�0�e+�W�5E�?��{n윲A��j8�0�e+�W�5E�?��{n윲A��j8�0�e+�W�5E�?��{n윲A��j8H4�e;�W5���?�h9ĺaK���G��0�e+ħ��>���~����.�o�%�m�8�H��== ��&�BȚ/e��:j�*C�(r�h)�K,�q���*Ȕ�X�N<��-+�s����k��#d��1xX~�ZR�`�eEĦ���	f�N`%p񝝽#h�4����C��J�5=���Wh�����i`7[�}�`��[�����B.�|�=��mh��p�X�)�/�(c@�Wm�t�?�����0���z;�r�^ ������A�9+�V�M�W����?(��a/E����Zp Z⡦��E�?}ŋ{^��'�v�5[�0,u�?��uE��N��b���u����j8������(������K֡���W��z���d����qE�̐��;n�a��+p��+�C���9�?�c9��Ċn���ܲ�>���p�Մ�<�9���D?B��{�t�A��<�d�p�'�Ss�+�n@}�wC�b�.�盀�p�e��W�5ʏ�
�_�l��BMz9�X7�����̬iDA!�p�o����5��3�eCM܆TǼQhy�H{�#L*NRYR��fQN�W9��Q�)(��|nN^~VYR�r�\D�1�El�T�{� ��P��M����P�9�9:�c���Qs��|u��>����)�?{�uE>�u�わa�p^N�ZR��^�M�W;�}�D?���j�uG���$�G88`�-XG�A��@s5e��j�vՍ.�W��AD��@�Wb-s9�A�*8��0�e�O��qH�K��ς�}%� �ַ��S�����5E��C�(��踾�v?@,�p�?��W;1TD��u�㼮�ghy�0��0�e��ZeȣDD��;�O�+T���?�F4g���W5é6?p6=%p[�e�xN�biQ���v7��o�����c��r.�h^����H�? �3�Y�Lmn5�d3Q�Xڒc������n��6������G���l7J���ί�n�v��r�E�W�02ׅ���w�z��eԩ8���v�J���!�̏�� Fr��O;f�|6�j��G�[GQa3����fWJ�tA����e�B��^5޷�(���܂�,�.���l�6�/�3�4>jR�4Wf_����j�V�8�=��{��!����*����A�n��t�PaȚ]� �̐��b{��x�����"��h�)��$Hp�.^�a�Ɨ�v�ƻF���V5�o�N���H����o��uخ�s�/�� @C�[rC�k�m *d�v�8^��2�5΋ GM�hJ�a�e'����XZ�*E��Ȭ���Z{>��	A��j��0ь'K�K��� K�":�gu��>�����VD��J�E��$����A�n��t�PaȚU�ھ��y� ���>l:ť�Q�e�ok�uEDPR-cP252�3<�;���8a"-�G��mf�<����K��*8�
:�%+����D�?��l��`�e�8���%@b�
�ں�hB���K�AA��p�QwR�W51?�?y#�9=�q�(�h�>���1�y�����g�]P������]�=�3�ߩD?���N��bv���22�%+m�c��g�/�F#m<���y�������8�	%����B�{Y��AT�l�08`�-XG�A*�y����J�<�壣���GM��ı��{�gv�OJփ���1�S,Z�5E" ��8h�jȐo�^~RYR��n�M�W��өD?�H`?���Pgx��V�	�P�(����J���b��A^v�ZR��V]N�W9)v�3@!s��ŵ>��ƏG8Pʽ��=�-��eh�'4�n?�E7�m�iٰ�ř-�-	���оk��X}B�z�0Z!��9Qa��#/=l9��aa��jŅ�}�e���[6r" ��98�����A*nauR�Zј�9�5�����g�3u���c8����Jz�Z�NN���&�	uQ">��d�8��:��L�8��Wd�l�Q�Яq�d� �f�U5�b@c?� 漫�5`�%��ߝf3,[�5Ej��>�fs�l�����~����1��W�5�!\D���{��G h��4
����?J c���O�GF���<����� �uE@@c���
ȘK%����"��Ἡ?���{��d�A���{�@�e�Ok�uE��4m�U�)�]12Wg8�����=�31a�ŠsNx|��Z@��j���(���{��H6��O������y�*�c���cX��(cj��6��z���S�^�>��p�Մ�</o��eF�{��/��<�d�,�.�W��AJ�@�Wb-aف>���p�Մ�<0Έ'�C�{�W
��<���0ь'�K��� K�'F�讜ڕQ�jL5�S#+�j]���C>(ߺ���Q�jP�rј��:�5�� ���!^F�ZR�Zь*E��8��������^��A9���0ь'G�K��� K�"&r��Ҩ��7�d40���	�#�)��+�W���v튯���VwҰG%�������]7)�Q�z.�Z#+Hǎ��J7����{n�n�._�<6����B�]�MF?�v�.�5b������;�G                                       =�2/        a����Fx���8n���Bd�����y����m����e���|Y���rQ���hE��؞�zx"��pn��fd��\Z�v�RP�l�HF�b�><�u42��m*(�a yYqM
eE ���䑱��։����}����u��άi��Ħa}��Еu��ҍi����a���yU���mM���eA�~���vt���lj���b`�}�XV�q�NL�i�DB��}:8b�q0.��i&$��]puUrmItaA�������x���肅���\y���Vq���Pe���2�y��$�q���e��}]��"uQ��,iI��&a�|zЕ�rpҍ�hf���^\�y�TR�m�JH�e�@>��y64��m,*��e" �}Y�qQ�iE؝���"�������������u����m����a����u����m���a���|Y���rM���dE��r��xvd��nlV��dbX|�ZXbr�PN,l�FD&b}<:P�u20R�i(&4�aFzU8lM
BbA ����������간����z��֤t��̖j���}��b�q����i����]��ptU��rjI��tdA~|���trx��jhfȄ�^\�z�TR�l�JH�b�@>Ȝy64��m,*��e" �zY�tQ�jE̜���&������������t����j����d����u���m����a��|Y���rM���dE��~��xvx��nlr��dbl{�ZXfs�PNXk�FDZc}<:�u20N�i(&H�a2{U,kM
6cA �ț�������꼃����{��֘s��̒k���}��f�q��X�i��Z�]��\sU��nkI��hcA~|���tr���jhv��`^�{�VTzs�LJ|c�B@��y86��q.,��e$"�{]�sQ�kI�c���\����N����H����2{���,k���6c���H�y��:�m��<�e���{Y���sQ���kE��̛�zx&��pn��fd��\Zs�RP�k�HF�c�><�u42�m*(��a VxUHnM
RdA ����������꠆���|���tr���fh���h�}����q��|�i��v�]���vU���lI��bA~|���tr莭jh�`^�z�VT�p�LJ�f�B@��y86Ԓq.,ƈe$"�~]�tQ�jE                                                                                                                                                                                                                                                                                                                                                                                                                                               