MZ�       ��  �       @                                   �   � �	�!�L�!This program cannot be run in DOS mode.
$       �h3�~`�~`�~`�,�`�~`�,�`�~`��k`�~`��}`�~`�~`j~`�,�`�~`�,�`�~`�,�`�~`�,�`�~`Rich�~`        PE  L <��H        � !	  �  �                                     �    J]  @                    �\ �   tN �    � p                   � �                                  8+ @              �                          .text   >�     �                   `.rdata  l]      ^   �             @  @.data   �0   `     J             @  �.rsrc   p   �     `             @  @.reloc  6%   �  &   d             @  B                                                                                                                                                                                                                                                                                                                                                        j�h��d�    P��$  �b3ĉ�$   SUVW�b3�P��$8  d�    ��$H  �L$�Y  �D$Ph�� V��D$$�L$ +���3ۅ���   ��$L  ;�r	�d�  �L$ ��h  �T$0RP�p�D$,�Pf���f��u��}+���;�s ��;�r���}r�U��U�L$,��v&���    f�*f;)��   ������u鋬$L  ;�r3�;�������   �D$$�L$ +�C��;��`���3�;�t	Q�F�  ���D$P�t$$�t$(�t$,�-�  ��3���$8  d�    Y_^][��$   3����  ��0  �f��f;Ƀ�����j�����$L  �p����L$$�D$ +���;�r	�8�  �D$ �4�3�;�t	P��  ���T$R�|$$�|$(�|$,��  �����l��������������QV��F��t�L$Q�N�VRQP�rD  �VR�b�  ���P�F    �F    �F    �B�  ��^Y����V��L$3�j�PQ�F   �F    ��f�F�n  ��^� ����U��j�h�d�    P��SVW�b3�P�E�d�    �e��u�}3ۉu�]���$    ;�vd�u�u��E�;�t�Mj�S3�Q�F   �^��f�F� n  O���]��u�ċu�};�t�]��$    V�����  ��;�u�3�SS��  �M�d�    Y_^[��]�������V��F��t	P�9�  ���P�F    �F    �F    ��  ��^������������j�h�d�    P��@SVW�b3�P�D$Pd�    ���wVhxj3�Sh����;�u2��L$Pd�    Y_^[��LË���   SP�ҋ����   SP�ҋ����   SP�ҋ���  SP�ҋ����   SP�ҋPj���U  �6����   �L$QV�ҋL$�D$PQ�\$�<�D$���   ;�tPSh   �t ���   �T$4hP R�N>  P�D$$P�\$h��  ��j�SP�OT�D$d�kl  �   9t$0r�L$Q���  ��3��D$0   �\$,f�T$9t$Lr�D$8P��  ���5p SSSS��SSSS�G|�։��   ���   ��  Ƈ  ��L$Pd�    Y_^[��L�����������j�h��d�    P���   SUVW�b3�P��$�   d�    ��$�   h@3�P�l$8�K�  ���   ��$�   9Xr�H��H3ҋ��D$,   �l$(f�T$�p��$    f���f;�u�+���PQ�L$���  ��$�   h,PƄ$�   �ܨ  ���L$XhP QƄ$�   ��<  ���T$$R��$�   PƄ$�   �7�  WP�L$TQƄ$  �s�  h$P��$�   RƄ$  �82  ��$  VPWƄ$   �A�  ��<9�$�   r�D$pP��  ��3ɾ   ��$�   ��$�   f�L$p9\$Lr�T$8R���  ��3��t$L�l$Hf�D$89�$�   r��$�   Q��  ��3҉�$�   ��$�   f��$�   9\$hr�D$TP��  ��3ɉt$h�l$df�L$T9�$�   r��$�   R�l�  ��3���$�   ��$�   f��$�   9\$,r�L$Q�A�  ��3҉t$,�l$(f�T$9�$�   r��$�   P��  ���ǋ�$�   d�    Y_^][���   �́�   �b3ĉ�$�   V��$�   W��$�   j�D$tVP�;  ��Ah3Ƀ��L$��t���L$QhxP�ҋL$�G;�t$��t�Q�H�у�$�   �1  �T$tR�  ��   U�   �b  �D$Xh0P苦  ��9hr�@����L$x9�$�   s�L$xSPQ������9l$tr�L$`Q��  ����[t��B�   f����    �}  Ƈ�    ��Bh�D$    ���a  ��T$RhxP��Ѓ|$ �E  ��Q�5��   �L$8f��Q�֍T$HR�֍D$(P�֋D$x�   f�L$�D$    9�$�   s�D$x�7�T$8R�L$LQ�T$0R�L$$QP�L$l�$5  ���   PW�ҋ5��D$XP�֍L$Q�֍T$(R�֍D$HP�֍L$8Q�֋D$����   �P�B���   ��   ��   ��t~��T$RP���   �Ѕ�|f�L$hQ�@��t;U�[�  ����t�Wx��L$�H�3��T$Rj Phs j j �l P�P �D$hP�`Ƈ  �L$��t��BQ��9�$�   ]r�L$tQ�R�  ����$�   _^3�3��!�  �Ĉ   � �����������V�����~$r�FP��  ��3��F$   �F �F��^��  �������������̋D$��Pw"��� �$�� h ��z  hW ��z  h@ ���y  Ë�� � � �   �������j�hT�d�    P���   SUVW�b3�P��$�   d�    �D$$hP�T�  ���L$dh�3�Q��$�   �:�  �   ��9~r�v���9xr�@���3�P�l$�� �D$;�tVP�\ ��l$9|$tr�T$`R��  ���   �t$t�\$p�D$` Ƅ$�   9|$<r�D$(P�q�  ���L$@h�Q�t$D�\$@�D$0 虁  ����$�   h�RƄ$�   �}�  ��9~r�^��^9xr�@���3�P�|$$�� ���t$��tSV�\ ���|$ ��$�   r�D$|P���  ���   ��$�   Ǆ$�       �D$| �|$XƄ$�   r�L$DQ��  ���\$X�D$T    �D$D ����   ����   ��$�   R��$�   P�f�  ���xƄ$�   r�@���jj ��$�   Qj P�Ճ��Ã�$�   Ƅ$�   r��$�   R� �  ����t&��$�   P�׋=� ��tV�׋D$��tP�װ��=� ��tV�׋D$��tP��2���$�   d�    Y_^][���   ������̃�SUV��nW9nv��  �~�;~v��  �USWP�D$ P���y�  _^][���̋D$��u� �L$�QRP�N  ���   � ������������U��j�h��d�    P��SVW�b3�P�E�d�    �e��u�}3ۉu�]���$    ;}tE�u�u��E�;�tW����  ��D�]��u��D�׋u�};�t�����  ��D;�u�3�SS��  �ƋM�d�    Y_^[��]�����:  �����������QV�t$�~E W�L$��uqS�   U�k��I �G�L$P������?9^@r�N,Q�\�  ��3҉n@�F<    f�V,9^$r�FP�;�  ��3ɉn$�F     Vf�N�"�  ���E ��t�][_^Y� �����̃�SUVW���o��u3���O+͸�$I�����������_��+͸�$I�����������;�s3�T$�D$ �L$Q�L$ R�GPQjS���������__^][��� ;�v���  �T$�RSP�D$P����8  _^][��� �����������j�h�d�    P��D�b3ĉD$@VW�b3�P�D$Pd�    �����    ��   �L$,�8.  j�D$P�L$4�D$`    �#  ���   V�L$�D$\苚  � �L$Qj�L$4��O  V�O<�����j h������  j j�L$4�$  @Pj�L$4�H�  �L$�D$X ��8  �L$,�D$X�����90  �L$Pd�    Y_^�L$@3��M�  ��P�������������U����j�hd�d�    P��  �b3ĉ�$�  SVW�b3�P��$�  d�    ��$(  �t$|�.-  j3�3��   hD�L$D��$�  �\$\�|$Xf�D$H��  �L$<Q�V$R��$P  PƄ$�  ��g  ���|$TƄ$�  r�L$@Q��  ��j3�3�hD�L$d�\$\�|$Xf�T$H�\$|�|$xf�D$h��  �L$\Q��<��$h  VRƄ$�  �hg  ���|$tƄ$�  r�D$`P�5�  ����3�f�L$|�̉d$,W3҉Y�yh���$�   ��$�   f�Q�4�  j	��$�  P��$L  �k  �L$<h0QƄ$�  ��  ���xƄ$�  r�p��p���̉Y3ҋƉy�d$,f�Q�X�d$ f���f;�u�+���PV��  j��$�  P��$L  �Dk  �|$TƄ$�  
r�L$@Q�T�  ����$�   3�h�P�D$\   �D$X    f�T$H�_�  �D$��$8  hQƄ$�  �A�  �D$,��$�  hRƄ$�  �#�  ��$�   ��$�  P��$�  QƄ$�  �>  ��$�   ��$P  h�
RƄ$�  �ޚ  ��$�   ��$   PƄ$�  �B*  �D$D��$�  h�
QƄ$�  褚  �؍�$�  h�
RƄ$  舚  ����$�  h�
PƄ$  �l�  ��D����$�  h�
QƄ$�  �M�  ���xƄ$�  r�P��P3�f�D$`�H�D$t   �D$p    �L$�d$ f���f��u�+D$�L$\��PR���  ��$H  R�D$`P��$�  QƄ$�  貸  ���~Ƅ$�  r�v���VP��$�  R�j#  ��$p  QP��$\  RƄ$�  �l�  ���   Ƅ$�  9wr����WP��$�  P� #  ��$�   ��TQP��$$  RƄ$�  ��  ��Ƅ$�  9sr�K��KQP��$T  P��"  �L$$QP��$�  RƄ$�  �ݷ  ����$�   Ƅ$�  9qr�I���QP��$  P�"  ��$�   QP��$�  RƄ$�  葷  ����$�   Ƅ$�  9qr�I���QP��$�  P�C"  ��$�  QP��$@  RƄ$�  �E�  ���L$Ƅ$�   9qr�I���QP��$�  P��!  ���L$Ƅ$�  !9qr�I���QP��$  Q��!  ��9�$�  r��$�  R��  ���   3�3���$�  ��$�  f��$�  9�$D  r��$0  Q��  ��3҉�$D  ��$@  f��$0  9�$�  r��$�  P�V�  ��3ɉ�$�  ��$�  f��$�  9�$�  r��$�  R�%�  ��3���$�  ��$�  f��$�  9�$,  r��$  Q���  ��3҉�$,  ��$(  f��$  9�$�  r��$p  P���  ��3ɉ�$�  ��$�  f��$p  9�$d  r��$P  R��  ��3���$d  ��$`  f��$P  9�$(  r��$  Q�a�  ��3҉�$(  ��$$  f��$  9�$�  r��$�  P�0�  ��3ɉ�$�  ��$�  f��$�  9�$`  r��$L  R���  ��3���$`  ��$\  f��$L  9�$�  r��$�  Q���  ��3҉�$�  ��$�  f��$�  9�$�  r��$�  P��  ��3ɉ�$�  ��$�  f��$�  9t$tr�T$`R�r�  ��3��\$t�|$pf�D$`9�$  r��$�  Q�J�  ��3҉�$  ��$  f��$�  9�$|  r��$h  P��  ��3ɉ�$|  ��$x  f��$h  9�$�  r��$�  R���  ��3���$�  ��$�  f��$�  9�$�  r��$�  Q��  ��3҉�$�  ��$�  f��$�  9�$  r��$�  P��  ��3ɉ�$  ��$  f��$�  9�$H  r��$4  R�U�  ��3���$H  ��$D  f��$4  9�$�  r��$l  Q�$�  ��3҉�$�  ��$|  f��$l  9�$�  r��$�  P���  ��3ɉ�$�  ��$�  f��$�  9�$H  r��$4  R���  ��3���$H  ��$D  f��$4  Ƅ$�  99�$�   r��$�   Q��  ��W3�j��$0  ��$�   ��$�   f��$�   �V  �D$;���  j��$�  P��$0  �T  �L$<Ƅ$�  :�>  ��$�  ���$�  Ƅ$�  ;�\$ �t$�I ��$�  ��t	;�$�  t�^�  ;�tY��uM�Q�  3�;Xu�E�  �T$9S(r ��u3�3�  ;^u�)�  ��S�L$@�����L$�(  �\$ �t$뒋붋6��j3��   3�hD��$�   ��$�   ��$�   f��$�   ��  ��$�   Q�T$@R��$�   PƄ$�  <�V]  ����$  h�
QƄ$�  =�Z�  ���xƄ$�  >r�P��P3�f�D$ �t$4�\$0�pf���f;�u�+���PR�L$$��  W�L$ Q��$�   RƄ$�  ?�ذ  ��j�SP��$  Ƅ$�  @�}B  �   9�$�   r��$�   P��  ��3ɿ   ��$�   ��$�   f��$�   9t$4r�T$ R�[�  ��3��|$4�\$0f�D$ 9�$  r��$   Q�3�  ��3҉�$  ��$  f��$   9�$�   r��$�   P��  ��3ɉ�$�   ��$�   f��$�   9�$�   r��$�   R���  ���D$H;�t"�L$Q�L$P�T$HRQP�p  �T$XR��  ���D$<P�\$L�\$P�\$T��  ����$�  Ƅ$�  9�+  3�j��  ��;�t��$  ��3���$  ��$$  ��$(  ��$,  j��$�  R��$0  Ƅ$�  B�7  j��$P  P��$0  Ƅ$�  C�  Ƅ$�  D9�$h  ��  ��$�   ��  ��$d  ���$L  �T$ �t$��$d  �   ��t	;�$L  t��  9|$ ��   ����   � �  3��L$ ;Hu���  �D$ ��P��$�   R��$�  �D$��s  �0�X��$�  ��t	;�$�  t��  ;�tj��u��  ;^u��  �D$��ul��  3��L$ ;Hu�~�  �S(�D$ ;P(|.�D$��uG�e�  3��L$ ;Hu�U�  �T$R��$  ������L$��$  �t$�������-����6낋 뗋 뼋�$(  +�$$  ��$I�������������  hD��$4  �pW  ��$0  Q��$  R��$�   PƄ$�  E�kY  ����$�   h|
QƄ$�  F�o�  ��Ƅ$�  G9Xr�@���P��$   �
W  VP��$�   RƄ$�  H��  ��j�3�VP��$  Ƅ$�  I�>  9�$�   r��$�   P���  ��3ɿ   ��$�   ��$�   f��$�   9�$  r��$   R��  ��3���$  ��$  f��$   9�$�   r��$�   Q�b�  ��3҉�$�   ��$�   f��$�   9�$�   r��$�   P�1�  ��3ɉ�$�   ��$�   f��$�   Ƅ$�  D9�$H  r��$4  R���  ����$  P��$�  Q��s  ����$  Rj j����3�9�$  �t$�D$~B�=���$    ��$  ��$�  s��$�  �Q�D$PV�׋D$@;�$  �D$|˹    f��$�  ��$�  �D$    ��$�   h
RƄ$�  K�u�  �   ��9Xr�x��x�5L W��PW�L$�  9�$�   r��$�   P���  ��h
��Ph
�L$�m  �L$|�q�\$S�L$@�  ����$�   R���   f�D$�D$$   ��$�   h0QƄ$�  N�̋  ���xƄ$�  Or�@���P�L$`�I  ����   W��$�  Q��$�   Q�L$(QPVƄ$�  P�ҋ5��D$\P�փ�$�   r��$�   Q�$�  ���D$3�3�PǄ$�      ��$�   f��$�   �֍�$�   Q�֍T$<R�֋D$P��S����$  r��$�  Q���  ����$L  Ǆ$     ��$  Ƅ$�   Ƅ$�  C��%  ��$�  Ƅ$�  B��%  ��$  ��  �   9�$$  r��$  R�V�  ��3��   ��$$  ��$   f��$  9�$�  r��$�  Q� �  ��3҉�$�  ��$�  f��$�  9�$�  r��$�  P���  ��3ɉ�$�  ��$�  f��$�  9�$|  r��$h  R��  ��3���$|  ��$x  f��$h  9�$`  r��$L  Q��  ��3ҍ�$(  ��$`  ��$\  f��$L  Ǆ$�  �����  ��$�  d�    Y_^[��$�  3���  ��]���������������Q�T$V�t$W�|$�D$ �D$P�D$R��QPVW���������    +΍�_^Y� �j�h��d�    P��DSUVW�b3�P�D$Xd�    ���\$hS�D$ �X�  ��3�;���  ����  ����  S�D$,P���}P  �D$`   �l$�D$(��T$RP�A �D$h�ЋD$;��Z  ��T$$RP�A$��3�9l$$�=  �l$h�   f�L$H�ωL$P�   f�T$,�׉T$4�l$H�t$��D$hP���ĉ(�l$`�h�H�L$h�H�L$@���ĉ�L$T�H�P�T$\�P�C,VƄ$�   �Ћ5��L$,Q�֍T$H�R�\$d�֋L$h3�3��D$;�t�� �T$Rh�Q�ЋL$h�D$;�tQ�l$ ��T$ RP�A8�D$h	�ЋL$ h�Q����t�D$�P��  ���D$�L$ Q���L$h�D$�\$`;�t�P�B�ЋL$h�D$`;�t��BQ��G;|$$������D$�D$`;�t��QP�ҋD$(�D$`����;�t��QP�ҊD$�L$Xd�    Y_^][��P� �l$(�l$`�l$$�����   �L$hQW�D$h��j3�hH�L$4�D$L   �l$Hf�D$8��  �T$h�L$,QR�D$h��������|$D�D$h�D$`r�D$0P�C�  ���L$hQ�D$L<   �D$P   �D$Tn   �D$XU   �0�=4���5x u7�T$hhn U jh  R��h�   jd�,�  ��P�֋D$hhn U Uh  P�׋t�
   ���$    �L$HQ�fG  �L$l���������Rj h   Q��jj
�П  ��P�փ�uŋT$hhn U jh  R��h�   jd覟  ��P�֋D$hhn U Uh  P�׋5�U��U�ְ�c��������������j�h��d�    P��   SVW�b3�P��$�   d�    ��$�   3��   �   ��$�   �D$�D$��D$   �D$h�D$    �D$$P�D$(   �D$,D�|$0�D$44�D$8   �D$<�\$@�D$D��D$H   �D$L��D$P   �D$T��D$X	   �D$\��D$`
   �D$d��D$h   �D$l|�D$p   �D$td�D$x   �D$|LǄ$�      ��$�   �L$;�t9�A����u�$�   3҉X�xf�P��$�   d�    Y_^[�Ĥ   � �AP��$�   Q��  ���x��$�   r�P��P��$�   3��^�~f�F�X��f���f;�u�+���PR����  ��$�   r��$�   Q�J�  �����i����������Q�D$��u	�W �Y� �V�T$RhP��D$    �D$    �Ћ���|/�D$��T$R�T$RP�A�Ћ���|�D$�T$�RP�A�Ћ��D$��t��QP�ҋD$��t��QP�ҋ�^Y� ��(  �b3ĉ�$$  SU��$4  VW��$@  �L$�D$�\-  �D$Ph�� U3��97tR�-�� ���$    �L$$�D$ +���;�s0��h  �T$0RP�Ջ�Q�T$0R�Ӆ�uF9�u���D$ �D$ 3�;�t	P���  ���D$P�t$$�t$(�t$,���  ��$8  �D$��_^][3���  ��(  �����������j�h��d�    P��$  �b3ĉ�$   SUVW�b3�P��$8  d�    ��$H  �L$�U,  �D$Ph�� V��D$$�L$ +���3ۅ���   ��$L  ;�r	��  �L$ ��h  �T$0RP��D$,�Pf���f��u��}+���;�s ��;�r���}r�U��U�L$,��v&���    f�*f;)��   ������u鋬$L  ;�r3�;�������   �D$$�L$ +�C��;��`���3�;�t	Q��  ���D$P�t$$�t$(�t$,�m�  ��3���$8  d�    Y_^][��$   3��+�  ��0  �f��f;Ƀ�����j�����$L  �p����L$$�D$ +���;�r	�x�  �D$ �4�3�;�t	P���  ���T$R�|$$�|$(�|$,���  �����l�������������̃�<V���������Z  j���^  �F|�Nx���   S�D$���   U�L$ �T$$�D$(W����؋�Ɔ�    �������R  ��h�  j �|$袙  ���D$�D$��}���5��|$���%��D$��}�����\$��D  3�9��   �D$����'	 ������I ��D  h�   Wj �T$,RU���d;�uhjj j j �D$@P�x��t7���$    ��L$0Q�\�T$0R�hjj j j �D$@P�x��u��^D  +�i��  ;�v��+��y���=  ���������   �1D  ��+|$h�  ���  ����   ���    t!�NQj ����(  ���j  �VRj���(  ���|$�D$��}���D$�\$�D$��}���D$�D$�������P����|$�D$��   �D$�l$�|$�L$�l$i��  Q���k   ����������X  _][^��<Ã�t"��u,��蓐  ��������F�P���   �Ћ��X  _][^��<Ã���������X  _][^��<������̃�$�Ax���   SU�-\V�t$4W�=x�D$�L$��B  h�   Vj �T$Rj���d��uSjj j j �D$(P�ׅ�t)�d$ �L$Q�ՍT$R�hjj j j �D$(P�ׅ�u��B  +�i��  ;�v��+��_^=  ]��[��$� �̋L$��)t-�D$�@��t"��RV�t$V�t$V�t$VQ�L$QP��^� 3�� �����3�� �����������j�hX�d�    PV�b3�P�D$d�    �D$����   ��T$Rh�P��D$(    �ЋD$�D$    ��tR�t$��VRhxhhP�A��j���Z  ���D$�D$������t��QP�ҋƋL$d�    Y^��� 3��L$d�    Y^��� �L$j �hZ  �L$d�    Y^��� ����̋D$�@��t��D$�A4��3�� �����V�����~$r�FP�!�  ��3��F$   �F �ΈF���  �D$t	V���  ����^� ���������j�hQ�d�    P��8�b3ĉD$4SUVW�b3�P�D$Ld�    �l$\���D$P�L$3�Q�͉\$\�l$0�\$(�y  �T$`R�D$0P�ω\$\�D$(   �L����   9pr�@����L$QS�T$,RSP�P� ���D$9t$Dr�L$0Q�6�  ��8\$��   �T$Rj@�� �D$���D$`P�L$0Q��������xr�@����L$�T$RQ�T$,RSP�P� �|$Dr�L$0Q�̾  ��9\$��   ��    3ҋ�f�T$0�D$D   �\$@�P���    f���f;�u�+���PV�L$4趹  �D$@�|F�tF�L$,Q���D$X   ���v  �8�|$D�\$Tr�T$0R�E�  ����+D$;D$�y����ŋL$Ld�    Y_^][�L$43����  ��D� �����̃�,�b3ĉD$(�D$0V��P�L$Q���D$   �����|$(�D$s�D$�T$R�L$Q�T$Rj P�P� �t$��t�t$8�|$(r�L$Q蘽  ���L$,��^3��k�  ��,� �������̃��T$S�\$V�t$W�|$ 2��D$�L$�D$�D$PQRWVS�}�  +�yxxx�������������ȋ��_�^+�[����j�h��d�    PQV�b3�P�D$d�    ��t$j��  ����t�0�3�����D$    ��  �F�@-�F�@�F� �F�@�F    �ƋL$d�    Y^��� ���������������Q����������̃|$ U����   �E ��t�|$ ��   SWP�����D$�;�}_[� �]� VSj ������u^_[� �]� �M Q����v�E �?RP�QV�c�  ���D$�T$�PRP�~P��  P�����3�f�^�U ��R���u ^_[3�]� 3�]� ���������������j�h��d�    P��$V�b3�P�D$,d�    �t$<V�D$8    �t$�D$    ��L  �D$VP�D$@    �D$   ��-  ��j�j P���D$@   �8  �|$(r�L$Q�$�  ���ƋL$,d�    Y^��0������j�hh�d�    P�� VW�b3�P�D$,d�    �L$@3�j�W3�Q�L$�|$�D$4   �|$0f�D$ �A8  �T$D�|$4�p�d$ f���f;�u�+���PR�L$�  �t$<j�W3��F   �~P��f�V��7  �|$(r�D$P�_�  ���ƋL$,d�    Y_^��,���������������̃�S�\$(U��EV�p�~- �аW�l$$�T$�D$��   �C�S�ȉD$�L$�T$ ��L$�~$�n �t$r�F��F�|$;�s����;�r�Ճ|$ r�K��K��vf�f;u������u�\$4;�s����f��f;������t�\$4�3�;��������D$��t�6��v�~- �g����l$$�T$�M ����t$(�|$$��tU�E�0��t;�t	螾  �T$�L$$;�u*SRjQ���  _�ȋ�D$,�I^]��H�@[��� ��E  �t$(�|$$�{�S�Nr�C��CR�QPRj 蓳  ��}�D$�L$SPQ�T$0R뗋D$0�8_�p^]�@ [��� ���������������������̃l$��S  ������UV��NW��u3���n+����|$���L  S�^��+�������?+�;�s�1�  �8;���   �������?+�;�s3���;�s��j U�6  �N���؋D$SPQ���~  �T$ RWP����  �L$P�FPQ���~  �F�V+������t	P���  �������^[_�F�N^]� �D$�L$ ��+���;׋�,�    �T$ sK�(QSP���A~  �F��+L$�T$ ��R+�WP���e�  n�v�D$�T$ R+�VP�mV  ��[_^]� S��S+�W����}  S�F�D$WP�n  �D$$�L$,Q�UP�4V  ��[_^]� ����������j0苼  ����t�     �H��t�    �H��t�    �@,�@- ����������j�h��d�    P��LVW�b3�P�D$Xd�    ���G�T$�D$    �RP���   �ЋL$����   ����   j h,  h,  j j j�Q�,����   �G����   j�P��jd�x �D$P��  ������   �L$<h|Q�=q  ���x�D$`    r�@���P�L$$��9  �D$�T$ RP�D$h�V������L$ �D$�f�  �L$<�D$`�����U�  �T$�L$QR�Xj
j �܊  �L$j
j �tU�ˊ  �T$ �DnVP��P  ���G����   j P�Ұ�L$Xd�    Y_^��X������QV�t$V�D$    ��������^Y�����V��W3�Vf����|$�   Wf����F��u��t�
   h �f��F ��)F  _��^� ��j�h��d�    P���   �b3ĉ�$�   SUVW�b3�P��$�   d�    ��   3�3��^�~�t$f�F�L$8h4Q��$�   �o  ��T$$h�RƄ$�   �o  UP��$�   PƄ$�   �V�  ���   9l$4r�L$ Q�'�  ��3҉\$4�|$0f�T$ Ƅ$�   9l$Pr�D$<P���  ����$�   R��3ɉd$8f�L$\��j�W��$�   3��Y�yR�\$|�|$xf�A�E1  �0�  ��$�   P��$�   Q�k�  ��T$|hRƄ$  ��n  UP��$�   P��$  茍  ��<�   9l$lr�L$XQ�]�  ��3҉\$l�|$hf�T$XƄ$�   
9�$�   r�D$tP�0�  ��3ɉ�$�   ��$�   f�L$t�  ��$�   �苄$�   s��$�   VPU�  ;�t��  �tU�0 �   9�$�   r��$�   R�²  ��3���$�   ��$�   f��$�   9�$�   r��$�   Q葲  ���Ƌ�$�   d�    Y_^][��$�   3��O�  ���   �����������̋P���������V��P�0 �~r�NQ�.�  ���F   �F    3�f�V^�������������U��j�h��d�    P��SVW�b3�P�E�d�    �e�jH�p�  �����u��E�    �u��E���t'�E�M�U��E�NP�N�V�'�  �M�ND�FE �ƋM�d�    Y_^[��]� �U�R�w�  ��j j �ó  �́�   �b3ĉ�$�   ��$�   V��$�   j
j@�D$PQ�D$    �g�  ��3��F   �F    �D$f�V�P���    f���f��u�+���P�D$P���$�  ��$�   ��^3����  �Ĉ   ������������̃l$�6L  �����́�,  �b3ĉ�$(  ��$4  V��$4  j�L$QP�D$    �� ��t=�D$h  �T$(RP�| ��t$�L$$Q���N4  ��^��$(  3��*�  ��,  Ë�$,  3��F   �F    f�V��^3����  ��,  �����������j�h8�d�    P��V�b3�P�D$d�    �D$4�L$03��t$9A��   �	���f�8u"�P�t$,R���3  �ƋL$d�    Y^�� Ë@P�T$3�Rf�L$��;�}�
   Pf�L$�D$�@  jV�T$R��P�t$4���L$�t$,Q���C3  �T$R���ƋL$d�    Y^�� ËD$,3��@   �pf�H�L$d�    Y^�� Ãl$�x  ������V��> u�Z�  �F�x- t^�K�  �H�y- u��x- u�I �ȋ�x- t��N^Ë@�x- u�N;Hu�F�ЋB�x- t�F^�������������̋D$�H�y- u�I ���H�y- t�����̃l$�3  �����̋D$�@��t��D$�A@��3�� ����̃y$r�AÍA���j�h��d�    P��\�b3ĉD$XSV�b3�P�D$hd�    �D$,h�P�!i  �   ��9pr�@����L$Qh  j Ph  ��( ����9t$Dr�T$0R設  ������   �D$HP�:����L$Q�D$x    �(l  �L$T��9t$`s�L$L9pr�@����T$\�RQjj P�D$ P�, 9t$(r�L$Q�;�  ���T$R�0 9t$`r�D$LP��  ���L$hd�    Y^[�L$X3���  ��h�����U�l$W�|$;�tUSV�w43ۃ>r�F�P�֬  ��3��   �^�f�N�~�r�V�R赬  ��3��F�   �^�f�FЃ�D��D;�u�^[_]�����������j�h��d�    P��VW�b3�P�D$d�    3�hL�|$�� ���t$��thXV�\ ���|$�D$     ��t<�D$P�D$  ��ׅ�|)�D$��t!����tV�� �ǋL$d�    Y_^��Å�tV�� �  ��L$d�    Y_^������̋D$V�5� W��P��hDt���֋�_^� �������������̃�SV��^W�~��+ϸyxxx���������u3��3;�v�հ  �L$���t;�t�°  �L$ +ϸyxxx����������L$$�T$ �D$QjRP���̈  �^;^v膰  �6W�L$�t$�\$�k�  �D$�L$�T$_^��P[��� ̋D$��SV��P�L$Q�������L$,�y�Qr�I����xr�@����RQjj P�P�, ���Ã|$ r�L$Q膪  ��^��[��� ��SV��^W�~��+ϸ�$I�����������u3��5;�v賯  �L$���t;�t蠯  �L$ +ϸ�$I������������L$$�T$ �D$QjRP���x  �^;^v�b�  �6W�L$�t$�\$觢  �D$�L$�T$_^��P[��� �������������j�h��d�    P��V�b3�P�D$d�    ��t$�F��PQRQ�D$P���D$0    �  �NQ�g�  �R�F    �F    �Q�  ���L$d�    Y^�������S�� VW�|$�GP�Ӌ���u��t��Bj����hDt��_��^[� ���������j�h��d�    P��X  �b3ĉ�$T  SUVW�b3�P��$l  d�    ��$|  �D$<h�3�P�\$��B  ���L$(h�Q��$�  ��B  �   ��9Or	�W�T$����|$9Hr�@���3�P�|$ �� ��l$;�t�D$PU�\ ���|$�|$8r�L$$Q�&�  ���D$8   �\$4�\$$�|$TƄ$t  r�T$@R���  ���D$T   �\$P�\$@;�t5�D$Ph<�ׅ�|%�D$;�tPh  �L$`Q�B�  �T$R���h  �D$\Pht�� ��$`  Q�� Phl�T$dR�� �F   �^��t-3�f�F��$`  �P�I f���f;�u�+���P��$d  Q�3�Sf�Vh����c�  ;�tU�� �Ƌ�$l  d�    Y_^][��$T  3���  ��d  ���������������S�\$U�l$VW��9ks莦  �{�D$+�;�s��;�uj��W����0  Uj ����0  _��^][� ���v��  �F;�s�FPW���M  ��vf�{r/�S�-��u�~��r�F_�  ��^][� �F_�  ��^][� �S�N�^��r����W�RQP�5�  ���~�~r��; _��^][� �����̋D$�    3�� �Q�T$V�t$W�|$�D$ �D$P�D$R��QPVW�  �΃���΍�_^Y� ��̃�V�t$$Wh�V�@������   S�\$0U�l$8��uQ��u3�D$h�P�`  ���xr�@���PV��:  ���L$��v  �L$<QUSVW� ][_^��� ��u�Wj�V�$h�V�`][_3�^��� _3�^��� Q�V��u9D$us�^Y� �t$��tdS�T$R�D$    �D$    �h�P��Ћ��T$Rh�V�ЋD$�L$;��Å�t��QP�ҋL$��t�Q�H�ъ�[^Y� 2�^Y� �������̃�V��NW��u3���F+����~��+���;�s�D$�����~_^��� ;�v蠩  �T$�RWP�D$P���Ԙ  _^��� �����������̋D$VP���  ����^� ������̃l$�m  �����̋T$V���W�F   �F    �F �x��@��u�+�PR���]  _��^� �������j�h(�d�    P��DSUVW�b3�P�D$Xd�    ������rLj3�h��L$�D$4   �t$0�D$  �+]  �D$P�L$4�t$d��  h�5�L$4Q�D$8��s�  �T$t�G�t$pj RPVP�,  ��G�   _;�u�h�G�(�O�i�"�|$l t�.�G;0u�(��n�G;pu�h�U�z, �E����   ��$    ��Q;
uQ�R�z, u�Y,�Z,��J�A, ��r�   ;qu
��V���  �F�X,�N�Q�B, �F�HQ���)  �{��z, u�Y,�Z,��J�A, ��r�];1u
��V���z)  �F�X,�N�Q�B, �F�@�H��P��z- u�B�P�Q�W;Bu�J��P;u�
��J��H�N�y, �F�����W�B�X,�D$h��h��L$Xd�    Y_^][��P� �V��> u���  �F�xE t�@�F�xE te^�ߦ  ��yE u �A�xE u��$    �ȋA�xE t��N^Ë@�xE u��$    �N;u�F�ЋB�xE t�N�yE t^郦  �F^��������QSV�t$�D$    �FW�|$�@�D Pj@�D$�� �~ ��t �~r�v���h    �D$PSV�3ɋ��G   �G    f�O�P�d$ f���f��u�+���PS��踛  S�� ��_^[Y����������̋T$�BV�0�r�0�~- u�V�r�p�I^;Qu�A��B� �J;u
���B� �A��B� �̃��AW�x�E �D$��   �L$�ASU�i��V�D$�L$��L$�   9D$r�	�_ ��;�s ��;�r��9G$r�W��W��v%f�f;u������u��f��f;Ƀ����u;�r3�;�����}���|$�?�E t��D$^][_��� ��������j�h��d�    PQV�b3�P�D$d�    ��t$��  3��N��j��A�A   P�D$�A�D$$P�����ƋL$d�    Y^��� �����SV��L$W��tI�~�F��r����;�r4��r���Ћ^�Z;�v��r� �T$+�R��QV���p
  _^[� �F���U�l$+�;�v�(;�s���  ����   �~������v��  �F;�s�FPW���n  ��vl�F�^��r2��0��u�~��r�F]3�_f���^[� �F]3�_f���^[� �ӋN�U�l$+�U�P�JR���  ���~�~r�3�f�{]_��^[� ������̋D$�@��t��D$�A8��3�� �����V�5� hDt�֋D$��P��^� ����U��j�h0�d�    P��T�b3ŉE�SVWP�E�d�    �e��E��E��F�u���u3���N+ȸ�$I����������ڋ}���~  �N+N��$I����������¹I�$	+�;�s��n  �8;��  ����I�$	+�;�s3���;�s��j S��  �N�E� �U�R�U�R�VRP�E��E��EPQ�E�    �@  �M��� QWP�ΉE��d����N�E� �U�R�U�R�VRP�E��EQP��?  �F�N+ȸ�$I���F�������ʃ����t�U�R�NQ�NQP�7  �VR�*�  ���E���    +ˍ���    +ωV���V�F�Z  �E��u��M�PV�!  V��  ��j j �4�  �N+M��$I�����������;���   �U�R�M��v����E�V��    +��ۍQRP���E�   �/�  �N+M�E�P��$I���F��������+�WP���E��0���^�v�E�U�R+�VP�E�   �#  ���M��   �M��    +��M��Q���R�U�P��   j j �\�  �E�P�M�迩���F��    +��P���P+�W���E�   �E��w�  �M��UQWR�F�S  �E�P�E�SP�  ���M��Kl  �M�d�    Y_^[�M�3��p�  ��]� ������������̋D$�@��t��D$�AD��3�� �����V�t$��t'�|$ j t�P��QX��
PV��^� ��HXV��^� ������������j�h��d�    PQV�b3�P�D$d�    ��j臟  3Ƀ�;�t�0�3���N�N�N�ƋL$d�    Y^�����������Q�T$�$ �$P�D$R�T$��Q�L$PQR�J������ ����S�\$V�t$;�t!W�|$j�j V����  ����;�u��_^[ËD$^[����������̃��D$�$Qh  �D$    �D$�L3�9$�������U��j�h1�d�    P��SVW�b3�P�E�d�    �e��u�}3ۉu�]���$    ;�vF�u�u��E�;�t�EP���ӆ  O��D�]��u�׋u�};�t����8  ��D;�u�3�SS��  �M�d�    Y_^[��]�����j�h��d�    P��\SUVW�b3�P�D$pd�    �ً�$�   U�*�������u覝  �;�C�D$��t;�t萝  ;t$t$�~$�N r�F��FQ�MPQj ���Ò  ��}x3�3��D$4   �D$0f�T$ �D$x�D$PU�L$@�71  PVW�L$ Q��Ƅ$�   ��&  �8�p�L$8��7  �|$4r�T$ R蚗  ��3��D$4   �D$0    f�D$ ��u(��  ;wu�ۜ  �F(�L$pd�    Y_^][��h� �?��������̃�LVj<�D$j P�Κ  �D$`�t$d��;���   �L$QP�T��ux�T$RV�X�D$<te�D$8�   tZ�   uS�L$�T$���ĉ�L$0�P�T$4�H�L$�P�T$���ĉ�L$,�P�T$0�H�P�Q  �� ��t�^��L�2�^��L�����������̃�S�\$(U��EV�p�~E �аW�l$$�T$�D$��   �C�S�ȉD$�L$�T$ ��L$�~$�n �t$r�F��F�|$;�s����;�r�Ճ|$ r�K��K��vf�f;u������u�\$4;�s����f��f;������t�\$4�3�;��������D$��t�6��v�~E �g����l$$�T$�M ����t$(�|$$��tU�E�0��t;�t	��  �T$�L$$;�u*SRjQ���/l  _�ȋ�D$,�I^]��H�@[��� �����t$(�|$$�{�S�Nr�C��CR�QPRj ��  ��}�D$�L$SPQ�T$0R뗋D$0�8_�p^]�@ [��� �����̋D$�@��t��D$�A,��3�� �����Q�b3ĉ$���L$;�tP�PS�XU�iV�pW�x�h�i�h�i�h�i�h�Q�q�q�y�Y�P�p�q�Q�P_�p^]�Q[�$3��>�  Y� ������������̋D$�@��t��D$�A$��3�� �����SU�l$VW�|$��9}s�Γ  �E�\$+�;�s�؋F���+�;�v�;�s�o�  ����   �~������v�U�  �F;�s�FPW���d  ����   �}r3�m�1��u�~��r�F3�_f���^][� �F3�_f���^][� ���F��r�V��V�N�S�\$+��\] S�P�JR�W�  ���~�~r�F3�f�x_��^][� �F3�f�x_��^][� ���V�t$W�|$;�tS�\$j�j S���  ��;�u�[_^������̃�4SU�l$D�E�V�u W�L$�D$    �\$�t$�}�E ��t;�t��  ;�t9��u1��  ;^u��  �K �T$�DJ�L$�D$�����\$�t$봋6�ЋL$Qj@�� �U�:�u �D$�D$L�|$$�t$ �d$ �]�E ��t;�t褗  ;���   ��u8蓗  3�;xu臗  �_ �\��u �w�  3�;xu�k�  �$r�G���ˋ��GSP�D$TP�R�  \$X����u5�9�  ;~u�/�  �O(�D$L����L$ �D$L�����|$$�t$ �R����6�̋T$H�|$R�D$,P���Y����   9Xr�@����L$�t$�QVjj PR�, 9\$@r�D$,P�H�  ��V�� _^]�[��4� ��������̋D$V���    ��t��Vh�P�ҋ�^� �����������̋�3�� ��@��H�H��������̃|$r�D$��uP�Đ  ��3�ÍD$VP�8�  ���|$ ��r�D$P蝐  ����^�������������̋D$�@��t��D$�A��3�� ����̃�V�t$$�W�=h h�   P��=  u\SU�-H�   �I �L$h�Q�aK  ��9Xr�@����VPR��9\$(r�D$P��  ���h�   Q��=  t�][j �d _^���������̃��AW�x�- �D$��   �L$�ASU�i��V�D$�L$��L$�   9D$r�	�_ ��;�s ��;�r��9G$r�W��W��v%f�f;u������u��f��f;Ƀ����u;�r3�;�����}���|$�?�- t��D$^][_��� ��������j�h?�d�    PQV�b3�P�D$d�    ��t$�`	�F@	�F(	�F��FxP�D$   �P ��  r���   P诎  ��3�ǆ     ǆ      f���   ���   �.  ���   �\  �~lr�FXP�j�  ��3��Fl   �Fh    �N<f�VX��T  �N$�T  �F �D$��t��QP�ҋF�D$ ��t��QP�ҋ��D$�����  �L$d�    Y^����̋D$VP���R�  �h��^� �������V�t$h�V�0�  ����uh�V��  ����u	�@ �^� �D$�L$��P�B��3�^� ������j�h��d�    P��<�b3ĉD$8V�b3�P�D$Dd�    �t$T�D$X�D$    3��F   �F    �t$f�N�T$,RP�L$T�D$   ��U  ����t<j�D$0P�L$Q�  ��j�j P���D$X   �s
  �|$(r�T$R�ی  ���ƋL$Dd�    Y^�L$83�袖  ��H�̃�SV��F��W�|$��t;�t	��  �|$9\$ uf�L$$�^���t;�t	��  �|$9\$(uF�N�QR���84  �F�@�F�F    � �F�@�F���D$_^�H�[��� ��$    ��t;|$$t	舑  �|$�\$ ;\$(t�L$�
���SW�D$P���U  �|$�Ƌ6�D$_�0^�X[��� �̋��tP�� ��̋D$VP���c�������^� �������j�h��d�    P��SUVW�b3�P�D$,d�    �L$(3ۉ\$$�|$@3��D$;�t���L$Qh�W�ҋD$�\$4;��E  �\$��T$RjP�A�D$@�Љ\$@�D$��T$$R�T$DRjP�A�D$D3��Ѕ���   �l$D;���   �\$�D$@��T$RhxP��D$@��;�|]�\$D�D$��T$DRP�AH�D$<�ЋD$D;�t*�T$ R�\$$�hpP��ЋD$ �D$4;���   �D$D�D$4;�t��QP�ҋD$�D$4;�t��QP�ҋD$@;�t�\$@��QP�ҋD$��T$$R�T$DRjP�AF�Ѕ��/����D$@�D$4;�t��QP�ҋD$�\$4;�t��QP�ҋD$�t$<�>;�t��HW�ыD$�D$4����;�t�P�B�ЋƋL$,d�    Y_^][��$� �t$<�L$(SPV�	����D$ �D$4;�t��QP�ҋD$D�D$4;�t��QP�ҋD$�D$4;�t��QP�ҋD$@�D$4;�t��QP�ҋD$�\$4;�t��QP�ҋD$�D$4����;��\�����QP���O����D$�@��t��D$�Q��3�� �����j�h	�d�    P��   SUVW�b3�P��$�   d�    �鋴$�   �F�HQ���,����F�@�F3ۉ^� �F�@�\$�E��RH�L$QP��$�   ��;���  �D$;���  �T$R�\$�hpP��ЋD$;�tL�\$��T$RP�A Ƅ$�   ��;�}Q�D$Ƅ$�   ;�t��QP�ҋD$��$�   ;�t��QP�ҋD$Ǆ$�   ����;�t��QP��2��  �\$$�D$hP���   f�L$T�   �L$\�|$h�T$�2�D$$P���ĉ8��$�   �x��$�   �x��$�   �x�|$h���ĉ8�|$|�x�H��$�   R�V,Ƅ$�   �H�ҋ=����D$TP�׍L$hQ��;�D$$}Ƅ$�   ;�������P�B�������P�L$D�4l  �D$@;�tA�\$D��T$DRP���   Ƅ$�   ��9\$Du@S���D$@Ƅ$�   ;�t��QP�ҋD$$Ƅ$�   ;��������QP���}����\$0�E��T$0RP�AHƄ$�   �ЋD$0;���  P�L$L�q  �D$H;��R  �\$,��T$,RP�A Ƅ$�   
�ЋD$,;��  ��T$PRP�A$��3�9\$P�L$d��  �\$4�   f�T$T�L$\��f�D$h�T$p�l$T�t$,�>�D$4P���ĉ(�l$l�h�H�L$t�H�L$|���ĉ��$�   �H�P��$�   �P�G,VƄ$�   �Ћ5��L$hQ�֍T$TR�֋D$4P�L$,�j  �L$4Q�L$|��	  �D$(;���   �\$L��R8�L$LQPƄ$�   �ҋD$Lh�	P� ����   �\$8�\$<�D$(��T$<RP���   Ƅ$�   �ЋD$(��T$8RP�A4�ЋL$8�5�Q�օ�tM�T$<R�օ�tB�D$8P��$�   ��  �L$<Q��$�   ��$�   RƄ$�   �d������t  �L$|�tV  �D$<�5�P�֋L$8Q�֋T$LR���D$(�L$xƄ$�   ;�t�Q�H�ыD$(Ƅ$�   ;�t�P�B�ЋD$4Ƅ$�   
;�t��QP�ҋL$dA;L$P�L$d�����D$,Ƅ$�   	;�t��QP�ҋD$HƄ$�   ;�t��QP�ҋD$0Ƅ$�   ;�t��QP�ҋD$DP���D$@Ƅ$�   ;�t��QP�ҋD$$Ƅ$�   ;�t��QP�ҋD$Ƅ$�   ;�t��QP�ҋD$��$�   ;�t��QP�ҋ�$�   �D$9^Ǆ$�   �����D$#;�t��QP�ҊD$#��$�   d�    Y_^][�Đ   � ����������V�t$�F�WPQ�~X  �V���FRP�oX  ���Ћ�_^�����̋P��  Y������̋D$�@��t��D$�Q��3�� ����̃|$ hDtt�� 3�� �� 3�� ��������������jH�K�  ����t�     �H��t�    �H��t�    �@D�@E ����������S�\$U�l$VW��9]s��  �}�D$+�;�s��;�uj��W����"  Sj ���"  _��^][� �����v见  �F;�s�FPW���fR  ��vz�}r3�M�1��u�~��r�F3�_f���^][� �F3�_f���^][� �M�~�nr�E ��ŋT$�Q�?SQ�N�	RP豁  ���~�~r�m 3�f�+_��^][� ��������������̋��t��QP���̋L$����w3ɍ�    R��  ����Ã��3����s��D$P�L$�D$    ��  h|2�L$Q�D$h�g�  ���������A��I��t�Q�H������j�h)�d�    P���b3ĉD$SUVW�b3�P�D$(d�    �|$8�l$<3��t$3��G   �w�|$f�G�\$@�t$0�D$   ;�vI���    �.QhX�T$$jR��R  �D$,���Pf���f��u�+���P�D$ P���T���F;�r��ǋL$(d�    Y_^][�L$3����  �� ���������������V��~r�FP��  ��3��F   �F�F^����������̃� V�D$h�P��:  �   ��9pr�@���S�L$Qh  j Ph  ��( ����9t$$r�T$R�  ����[tD�D$P�>  ��9pr�@����L$PQ�$ 9t$ r�T$R�E  ���D$P�0 ^�� ���������̃�V�D$P�� �L$Q�T$R�� �T$�L$3�3���V ��*h��� ��!Nb�QP��  ^������̋T$SVW���tF�~�F��r����;�r1��r���ȋ^�;�v��r� �L$Q+�RV���C  _^[� �F���U�l$+�;�v�(;�s��}  ����   �~����v��}  �F;�s�VRW����$  ��va�F�^��r.��,��u�~��r�F]_�  ��^[� �F]_�  ��^[� �ӋNU�l$+�UP�Q��}  ���~�~r��; ]_��^[� �������̋D$V���    ��t��Vh�P�ҋ�^� ������������VW�|$�P��������u2���u_3�^� �>�    ��t��Vh�P�҅�t��HW�ы_^� ���V��N+N�yxxx��������W�|$�;�r菂  �V�����_��^� ������j�h��d�    P��SVW�b3�P�D$d�    ��3ۉ\$�\$�F��T$RP�AH�\$(��;�|�D$;�t{�T$R�\$�hpP��ЋD$�D$ ;�tU�L$,�|$(QPW��������D$�\$ ;�t�P�B�ЋD$�D$ ����;�t��QP�ҋǋL$d�    Y_^[��� �D$�t$(��D$ ����;�t��QP�ҋƋL$d�    Y_^[��� �̋T$V��3��F   �F    f�F��W�xf���f��u�+���PR���w  _��^� �D$V���    ��t��Vh�P�ҋ�^� �����������̋T$�BV�0�r�0�~E u�V�r�p�I^;Qu�A��B� �J;u
���B� �A��B� ��V�t$h�V�w  ����t�D$�L$��P�B��3�^� h�V�vw  ����t5�D$��t�T$�H�
��QP��3�^� �T$3ɉ
��QP��3�^� h�V�/w  ����u�h�V�w  ����t�D$��t��T$�H�
��QP��3�^� h�V��v  ����t�D$��t��T$�H�
��QP��3�^� �@ �^� ������������̋D$�T$P��Q�L$QR�  ��� ��VW�|$j����   j W������j�j �GP�N�����O8�N8�W<�V<�G@_�F@^� �j�h��d�    P��(SUVW�b3�P�D$<d�    �|$L�D$T�t$P3ۉ\$3��G   �_�|$�D$f�O�N+N��$I����������\$D�D$   ��   ;�vs3�;�r��~  �F�T$�RP�D$(P�`S  ��j�j P���D$P   �	����|$8�D$D r�L$$Q�y  ���N+N��$I����������C�;�r�3ۋO�T$�R��+�;�wj�P���a  �+�SP����1  �ǋL$<d�    Y_^][��4��������������̋T$�V�p�2�p�~- u�V�r�p�I^;Qu�A�P�B� �J;Qu�A�P�B� ��P�B� ��������������SU�l$VW�|$��9}s��w  �E�\$+�;�s�؋F���+�;�v�;�s�w  ����   �~����v�xw  �F;�s�FPW���w  ����   �}r/�m�-��u�~��r�F_�  ��^][� �F_�  ��^][� ���F��r�V��V�NS�\$�+�UP�Q�w  ���~�~r�F�8 _��^][� �F�8 _��^][� �����V���(����D$t	V�4w  ����^� ��j�h��d�    PQV�b3�P�D$d�    ��t$j�|  ����t�0�3�����D$    �#����F�@E�F�@�F� �F�@�F    �ƋL$d�    Y^��� ��������������̋D$VP���-  ����^� �������U��j�h��d�    P��SVW�b3�P�E�d�    �e�j0��{  �����u��E�    �u��E���t�E�M�UP�EQ�MRPQ���`  �ƋM�d�    Y_^[��]� �U�R��u  ��j j �?x  �������������̃l$�?  ������S�\$V��W9^s�su  �F�|$+�;�s����vU�NU�n��r	�U �T$��l$��r�U ���+�P�D$��P+�Q�R��u  �F+ǃ��~�Fr�m �( ]_��^[� ��������������h��v  �����j�h �d�    P��H�b3ĉD$DSUVW�b3�P�D$\d�    �t$l3ۋ�\$�D$pP�L$@Q�͉\$l譪���   9xr�@����T$R�U S�L$$QSPR� ���D$9|$Tr�D$@P�t  ��8\$��   �D$��Pj@�D$ �� �L$pQ�T$$R�͋��9����xr�@����L$QW�T$$RSP�E P� �|$8r�L$$Q�,t  ��3ҽ   ��f�T$@�l$T�\$P�P��$    f���f;�u�+���PW�L$D�&o  W�D$h�� j�S�L$D3�Q�n�^��f�F�O����   9|$Tr�T$@R�s  ��3��l$T�\$Pf�D$@�j�S�D$|3��F   �^P��f�V����9�$�   r�L$xQ�ms  ���ƋL$\d�    Y_^][�L$D3��1}  ��T�$ �������������̃l$����������̃l$�  ������V��> u�zx  �F�x- t�@�F�x- te^�_x  ��y- u �A�x- u��$    �ȋA�x- t��N^Ë@�x- u��$    �N;u�F�ЋB�x- t�N�y- t^�x  �F^��������Q�L$�T$�$ �$P�D$Q�L$R�T$PQR������������j�hH�d�    P��`�b3ĉD$\SUVW�b3�P�D$td�    �D$4h�	P���M-  ��3��x�|$|r�H��H�   3ҋ��l$,�|$(f�T$�pf���f;�u�+���PQ�L$�m  �D$P���   Ƅ$�   �;������̉d$Lj�W3҉i�yPf�Q���������   ����9\$,r�D$P�wq  ���l$,3Ƀ���|$(f�L$�l$|9\$Lr�T$8R�Nq  ��;�u2�L$P�e���h�  W�L$XǄ$�      �����L$P���l$|�̾���x   ��xr�ƋL$td�    Y_^][�L$\3���z  ��l�̃�V��~ Wu!�D$,�N�|$ PQjW���G  ��_^��� �D$$�V�:���t;�t	�v  �D$$�L$(SU;�u9�|$4��QW�N�;_  ����  �D$0W�|$,PjW���/G  ][��_^��� �~���t;�t	�u  �L$0;ϋ|$4u=�N�A��WP�N��^  ���B  �V�BW�|$,Pj W����F  ][��_^��� ��Q�^W���^  ��tk�L$,�T$0�L$�L$�T$�<����l$W�EP���|^  ��t>�M�yE W�|$,��tUj W�oF  ][��_^��� �T$4RjW�VF  ][��_^��� �D$0W��P���*^  ����   �L$,�T$0�F�L$��L$�L$�T$�D$�  �T$R�L$�N<  �l$��u�EPW����]  ��t>�D$0�H�yE W�|$,��tPj W��E  ][��_^��� UjW�E  ][��_^��� W�T$R���K�����L$(][��@_�A��^��� ̋D$hH2�L$Q�D$��p  ���������j�h��d�    P��D  �b3ĉ�$@  SUVW�b3�P��$X  d�    ��$h  ��$�   3�P�t$�� ��$�   Q�T$`R�Ǽ������$�   P�L$LQ��$p  諼��hTP�T$<RƄ$|  ����WP��$  PƄ$�  ��G  ��(�   9\$<r�L$(Q��m  ���   3҉|$<�t$8f�T$(9\$Xr�D$DP�m  ��3ɉ|$X�t$Tf�L$DƄ$`  9\$tr�T$`R�|m  ��3�j3�f��$�   hL��$�   �|$|�t$xf�D$h��$�   ��$�   �vh  h  ��$R  3�VPƄ$l  f��$X  �p  ��h  ��$P  Q�� f9�$L  �   ��$L  �P�I f���f;�u�+���P��$P  R��$�   ��g  jV�D$$P��$�   �D$(\   � X  ���t-��$�   @;�wj�P��$�   �  �+�VP��$�   �%  3ɉt$�t$�t$ ��$�   ��$�   f��$�   ��$�   ��$`  9�$�   s��$�   VV�T$(R�L$ Q�T$(RVVP�� ����   �D$PhD��$  h�   Q�m>  ��3ҍ�$  f�T$(�|$<�t$8�P�f���f;�u�+���P��$  P�L$,��f  j�V�L$,Q��$�   Ƅ$l  	�#�����$`  9\$<r�T$(R�k  ��hT��$�   P��$�   Q�_�����$�   RPUƄ$x  
�hE  ��9�$�   r�D$|P�;k  ��9�$�   r��$�   Q�"k  ��3҉�$�   ��$�   f��$�   9�$�   r��$�   P��j  ��3ɉ�$�   ��$�   f��$�   9�$  r��$�   R��j  ���ŋ�$X  d�    Y_^][��$@  3��~t  ��P  �����������V�5� hDt�֋D$��P��^� ���́�0  �b3ĉ�$,  S�tU��$@  VW��$D  j j h  W��3��D$��vJ�L$QVhs  �D$HW�D$,    �D$<�   �D$8�ӍT$<RU� ��t	F;t$r��j Vh  W�Ӌ�$<  _^][3��s  ��0  ������������V��F|W�=P P�׋��   Q�׋��   R��_^������������V��> u��n  �F�xE t^��n  �H�yE u��xE u�I �ȋ�xE t��N^Ë@�xE u�N;Hu�F�ЋB�xE t�F^��������������j�hX�d�    P��4SUVW�b3�P�D$Hd�    �D$X3�;���  9\$\��  �\$��T$RP�A �\$X�ЋD$;���  ��T$$RP�A$��3�9\$$�r  �\$X�   f�L$8�ωL$@�   f�T$(�׉T$0�l$8�t$��D$XP���ĉ(�l$P�h�H�L$X�H�L$<���ĉ�L$P�H�P�T$X�P�C,V�D$x�Ћ5��L$(Q�֍T$8R�D$T�֋D$X3�3ɉL$;�t��T$Rh�P��ЋD$X�L$3��D$P�T$ ;�t��T$ Rh�P��ЋD$X�L$�T$ ;�tE�\$��D$PQ�J8�D$X�ыT$\�D$RP������   �L$Q���D$X�L$�T$ �D$P;�t��HR�ыD$X�L$�D$P;�t��BQ�ЋD$X�\$P;�t��QP��G;|$$������D$�D$P����;�t��QP��2��L$Hd�    Y_^][��@� �D$P���D$ �D$P;�t��QP�ҋD$�D$P;�t��QP�ҋD$X�\$P;�t��QP�ҋD$�D$P����;�t��QP�Ұ�j�hx�d�    PQV�b3�P�D$d�    ��t$�L$3�j�PQ�F   �F    ��f�F������D$ 3�j��NR�A   �A    P�D$     f�Q�����ƋL$d�    Y^��� ���̋A�T$��t4��t�Q��Qh�RP�^?  � ��t��u�IQh�P蔝��� �@ �� ���������j�h	�d�    P��SVW�b3�P�D$d�    �|$,�t$03ۉ\$�G   �_�|$�_�\$$�D$   ;�t/�:�u8^t$�N2Ȁ�2Ȁ� j�T$�L$R���a������ыǋL$d�    Y_^[����������V�t$W�|$;�t/���~r�FP��d  ��3��F   �F    f�N��;�u�_^�V���h�f  �D$t	V�d  ����^� ������������3�� ����������̋��tP�d  Y������������������̃�\VW�D$P�l�5P3��D$,�D$<�D$H�D$X�D$P�D$4�D$8�D$<�D$D�D$H�D$P�D$T�D$X�D$`�D$d�D$�D$�D$ �D$$�D$(�D$,�D$L�D$0�D$�D$@   �D$\   ��j���֋ȸ��  ����5Dj�D$$�  �D$l�D$���  ����L$Qj�D$x�D$$��j�T$0Rj��j�D$LPj��j�L$0Qj��h�   jd��8  ��P�x j�T$LRj�֋D$�L$PQ�8_^��\����������̋T$�V�p�2�p�~E u�V�r�p�I^;Qu�A�P�B� �J;Qu�A�P�B� ��P�B� ��������������j�hV�d�    P��t  �b3ĉ�$p  SUVW�b3�P��$�  d�    �D$lP�L$h�Q��  ��3۽   ��$�  9hr�p��p����3ҋ��A   �Y�d$4f�Q�x��I f���f;�u�+���PV�z]  �[  �� ����Ǆ$�  ����9l$0r�D$P�b  ����t
�@ ���   �L$lQ�T$TR��<  �D$ h�PǄ$�     �  �L$d��9l$hs�L$T9hr�@���QP��$�   h  Q�&4  ��9l$0r�T$R�a  ���5�D$|Ph   ��֍L$4h�Q�  �L$\��9l$hs�L$T9hr�@���QP��$�   h  R�3  ��9l$Lr�D$8P�3a  ���L$|Qh  ���9l$hr�T$TR�a  ��3���$�  d�    Y_^][��$p  3���j  �Ā  ��������������̋D$�L$;�t�T$V�2�0��;�u�^��̋L$�D$P�2����   � ���������̋D$V���u���^� P�����u�h ����������̃�U�l$VWU���~������|$��u�e  �S�^�D$��t;�t�e  ;�[t*�$�G r����P�EWPj ����Z  ��|�L$��N��L$�T$�L$��D$ �I_^��H]��� �V��~4r�F P��_  ��3��F4   �F0    f�N �~r�VR�_  ���F   �F    3�f�F^����������������S�\$V��W9^s�#_  �F�|$+�;�s����vi�NU�n��r	�U �T$��l$��r	�U �T$��l$�T$+��P�;�B+�P�Q�L$$�YR�_  �F+ǃ��~�Fr�m 3�f�LE ]_��^[� ��������̋L$����w3ɍ	R�\d  ����Ã��3����s�D$P�L$�D$    �_  h|2�L$Q�D$h��`  ���������̋L$3���t�����v�W ���|FSVW�|$�q��L$�D$PQVW3��a  ����|;�wu3�f�w_^��[�3�f�w�z �_^��[���������������j�h��d�    PQSUVW�b3�P�D$d�    �l$,�E�x3�W�\$��]  �����t$,�}�\$ r�m���SSWVj�USS�� �|$(���G   �_�_�P��I �@:�u�+�PV���^  ;�t	V�m]  ���ǋL$d�    Y_^][�������������̋L$����w3ɋ������R��b  ����Ã��3����Ds܍D$P�L$�D$    ��]  h|2�L$Q�D$h�C_  ��SUV�t$�l$W�|$��+ϸ�$I�����������    +��ɋ�+�;�t+����V�.�����;�u�_^]��[����������U��j�hi�d�    P��4�b3ŉE�SVWP�E�d�    �e��u�}3�3��ủu��E�   �]�f�Eԉ]��E�;}th�uĉu��E�;�tj�3��F   �^S�U�f�NR������W���E��0������ũ�븋uȋ}�;�t�]V���0A  ��;�u�3�SS�!^  �}�r�E�P�[  ���ƋM�d�    Y_^[�M�3��e  ��]Ã�V��~ Wu!�D$,�N�|$ PQjW���ܷ����_^��� �D$$�V�:���t;�t	��`  �D$$�L$(SU;�u9�|$4��QW�N��I  ����  �D$0W�|$,PjW������][��_^��� �~���t;�t	�h`  �L$0;ϋ|$4u=�N�A��WP�N�I  ���B  �V�BW�|$,Pj W���$���][��_^��� ��Q�^W���YI  ��tk�L$,�T$0�L$�L$�T$�l����l$W�EP���,I  ��t>�M�y- W�|$,��tUj W迶��][��_^��� �T$4RjW覶��][��_^��� �D$0W��P����H  ����   �L$,�T$0�F�L$��L$�L$�T$�D$������T$R�L$��&  �l$��u�EPW���H  ��t>�D$0�H�y- W�|$,��tPj W����][��_^��� UjW����][��_^��� W�T$R���K�����L$(][��@_�A��^��� �U��j�h��d�    P��SVW�b3�P�E�d�    �e����}�E�������v���"�_������������;�s�����+�;�w�4�Nj Q�E�    �%  ���E�(�E�e��E�@j P�E��%  �E����� Ë}�u�]��v �r�G��GSP�E�VRP�X  ���r�OQ�X  ���M�G�  ��w�_��r��� �M�d�    Y_^[��]� �u�~r�VR�IX  ��j �F   �F    j �F �Z  ��UV�t$�~- W���uD�GP��������~$�?r�NQ��W  ��3��F$   �F     Vf�V��W  ���- ��t�_^]� �����U����j�h��d�    P��  �b3ĉ�$�  SVW�b3�P��$�  d�    ��$�   ��3�P�t$P�\$H�� ��$8  芢��Sj��$@  ��$�  �D�����$�   ;�tOj��$<  �
8  j��$<  ��7  j��$<  ��7  j��$<  ��7  ��$�   Rj��$@  �;  ���   �H���   Q���Br���G�@�G�_� �GW�Ή@�������e  ��$  h�R��  ���xƄ$�  r�P��P3�f�D$���D$(   �\$$�xf���f;�u�+���PR�L$�Q  �L$Q���   Ƅ$�  �ɽ��j�SP���   �����|$(r�T$R�"V  ��3���$4  �D$(   �\$$f�D$��$�  r��$   Q��U  ��9�  t?Sj
��$@  �˗��������+�=0*  v ����Pj
��$@  �W:  ���   R�V  ��$  h�	P��  ���xƄ$�  r�H��H3ҋ��D$(   �\$$f�T$�x���    f���f;�u�+���PQ�L$�vP  �D$P���   Ƅ$�  讼�����̉d$dj�S3��A   �YPf�Q�����'������|$(��r�D$P��T  ��3Ƀ�$4  �D$(   �\$$f�L$��$�  r��$   R�T  ��;�tWS��$@  �H9  ��$  h�P��  ���xƄ$�  r�H��H3ҋ��D$(   �\$$f�T$�x��I f���f;�u�+���PQ�L$�vO  �D$P���   Ƅ$�  讻�����̉d$dj�S3��A   �YPf�Q�����'������|$(��r�D$P��S  ��3Ƀ�$4  �D$(   �\$$f�L$��$�  r��$   R�S  ��;�vWj��$@  �G8  ��$  h�P��  ���xƄ$�  r�P��P3ɋ��D$(   �\$$f�L$�x�d$ f���f;�u�+���PR�L$�vN  �T$R���   Ƅ$�  论��j�3�Sf��$d  �   P��$d  ��$|  ��$x  �����|$(r�T$R��R  ��3��|$(�\$$f�D$��$4  Ƅ$�  r��$   Q�R  ��3҉�$4  ��$0  f��$   9�$l  t��$X  Pj	��$@  蕧����$t  hlQ�  ���xƄ$�  r�H��H3ҋ��|$p�\$lf�T$\�x��    f���f;�u�+���PQ�L$`�VM  �D$XP���   Ƅ$�  莹�����̉d$dj�S3��A   �YPf�Q�l����������|$p���|$xr�D$\P��Q  ��3Ƀ�$�  �D$p   �\$lf�L$\Ƅ$�  r��$x  R�Q  ����  s�D$x  �D$,P��ǆ�   �����O  ��$�   Ƅ$�  �;���j��$�   Q��$@  Ƅ$�  �M���j��$�   R��$@  Ƅ$�  �/���j��$   P��$@  Ƅ$�  �����L$<+L$8�yxxx��������3��Ƅ$�  ��  3ۍ�    �L$LV�f9  ���A  �L$<+L$8�yxxx���������;�r�V  �L$8�T�L$LR��$�vl���L$<+L$8�yxxx���������;�r��U  �L$8�TR��$   ��  � �L$<�|$8+ϸyxxx���������;�r	�U  �|$8�|8 t
�L$L���   �D$<+ǋȸyxxx���������;�r	�YU  �|$8�P��$�   �~  � �L$<�|$8��+׸yxxx���������;�r�U  �L$<�|$8�|@ tk��+׸yxxx���������;�r��T  �L$<�|$8�+ωT$H�yxxx���������;�r	��T  �|$8�P��$�   ��  �L$H�Q@���   ��$�   �T$|�D$T+ωT$P�yxxx���������;�r	�tT  �|$8�P��$�   Q��$�   ���������t;D$Pt�ET  �T$T9WtY�L$<+L$8�yxxx���������;�r�T  �L$8�P��$�   R��$�   �'����H�QR��$�   P��$�   �<  �L$<+L$8�yxxx��������Fʃ�D;��������$�   Rj��$@  �Q����D$|Pj��$@  �>�����$�   Qj��$@  �(���j j��$@  �������$t  hHR�D$P�"	  ���xƄ$�  r�P��P3�f�D$���D$(   �D$$    �pf���f��u�+���PR�L$��H  �t$L���   ���   ���   �D$�T$TP��$�   RƄ$�  �3  �����t;�t��R  �D$T9G��   ��$  hHQ�o  ���xƄ$�  �D$D   r�H��H3�3ҋ��D$p   �\$lf�T$\�x�d$ f���f;�u�+���PQ�L$`�H  �D$XP���   Ǆ$�     �D$H   �C������̉d$lj�S3��A   �YPf�Q�!���輻��������   3��D$Dt,�d$D��|$pr�D$\P�jL  ��3��D$p   �\$lf�L$\�D$DǄ$�     t6��$4  r��$   R�+L  ��3�Ǆ$4     ��$0  f��$   �|$(r�L$Q��K  ��3҃�$�  �D$(   �\$$f�T$Ƅ$�  r��$x  P��K  ���L$<+L$8�yxxx����������c  ���   ��V  9|$H�L  �_���+�  ;D$x�7  j�T$\R��$@  �|������   P�L$0Ƅ$�  ������P��$   �Z�����   Q�L$0Ƅ$�  �����P��$x  ��Y����$  R�L$\Ƅ$�  �  ���   P�L$0�������   Q�L$0������$  R�L$\�x<�r  � ;s[���  h@  h�  ��  ��P�x ���   Q���>3  ���   R�L$0Ɔ�   �7���P���O������   P���|����$t  �  ��$  ��  �L$XƄ$�  舠����$�   Ƅ$�  �t����L$|Ƅ$�  �c�����$�   Ƅ$�  �O�����$�   ;�t	P��I  ����$�   Q��$�   ��$�   ��$�   ��I  �D$<��;�t"�T$PR�T$@�L$8QRP蹜���D$HP�I  ���L$,Q�\$<�\$@�\$D�I  ����$p  r��$\  R�uI  ���t$L3�Ǆ$p     ��$l  f��$\  �N|Q�T ��$8  Ǆ$�  ����������$�  d�    Y_^[��$�  3���R  ��]�����j�h�d�    PQVW�b3�P�D$d�    ��t$�|$ W�<J  3�j��N���GR�A   �QP�T$$�Q�š���ƋL$d�    Y_^��� ��������������̋D$�T$+���V�t$��    +��~QRQV��H  ����^��j�h��d�    P��(SUVW�b3�P�D$<d�    �ًl$LU�M�������u�M  �;�C�D$��t;�t�sM  ;t$t$�~$�N r�F��FQ�MPQj ���B  ��}o3�j�RU�L$(�D$@   �D$<    f�T$,�>���3�l$8�D$PVW�L$ Q�ˉl$T�����|$4�8�pr�T$ R�G  ��3��D$4   �l$0f�D$ �3�;�u*��L  3�;wu��L  �F(�L$<d�    Y_^][��4� �?�����������������Q�L$�T$�$ �$P�D$Q�L$R�T$PQR�����������̋D$�@��t��D$�A ��3�� �����S�\$V�����+F;�w�GF  ����   W�~������v�,F  �F;�s;�NQW����  ��v`�D$�NPSQ���2  �~�~r=�F3�f�x_��^[� ��uω~��r�F3�_f���^[� �F3�_f���^[� �F3�f�x_��^[� ���������������U�l$VW���tF�V�F��r����;�r1��r���ȋ~�;�v��r� �L$Q+�UV������_^]� �|$���v�=E  �F;�s �VRW���<�����vV�NS�^��r,��*��u�~��r�F_�  ��^]� �F_�  ��^]� ��WUQP�iE  ���~�~r��; [_��^]� ���������̸@ �� �������̃l$����������̋D$�L$;��T$|;�~�D$;�|';�#�D$�L$;��T$ |;�~�D$;�|;���2������������j�h��d�    P��VW�b3�P�D$d�    �|$(�D$,�D$    3��G   �G    �|$f�O�L$ �D$   ��t;�p�F���u8t-�����%�   Ѓ� ��j�T$�L$R���M������ȋǋL$d�    Y_^������́�   �b3ĉ�$�   ��$�   U��$�   �D$���  VW�L$ h�Q�����   ��9xr�@���Pjj �� ��9|$8r�T$$R�C  ��Sh�  3�V�D$D   �D$@    f�D$0�h �P =  ��   ��$�   Q�	U��jD�T$Hj R��F  3����D$�D$�D$�D$ ��$�   �D$@D   9�$�   s��$�   �L$Q�T$DRj j j j j j Pj �X ��t�D$P�ӋL$Q��9�$�   r��$�   R��B  ����tV��[_^�D$UP舁����$�   ]3��L  �Ĕ   � ���T$S�\$V�t$W�|$ 2��D$�L$�D$�D$PQRWVS����+�$I�������������    +ȍ�_^[����̋D$��yE u�d$ ����yE t������̃� W�D$h@P�M����   ��9xr�@���S�L$Qh  j Ph  ��( ����9|$$r�T$R��A  ����[tbV�D$h,P�������9xr�p��ph$�L �L$�Ph$jj VQ�, ^9|$ r�T$R�wA  ���D$P�0 _�� ������������j�h��d�    P��l�b3ĉD$hSVW�b3�P�D$|d�    ��$�   �D$0h�3�P�t$�C����؍L$h�Q��$�   �+���SP�T$dRƄ$�   ��  ���|$,r�D$P��@  ���   3ɉ\$,�t$(f�L$�|$HƄ$�   r�T$4R�@  ���L$hQ���̉d$03�j�f�D$XV�D$t3҉Y�qP�\$t�t$pf�Q������9  ��$�   QW�  ��(�|$dr�T$PR�<@  ���ǋL$|d�    Y_^[�L$h3��J  ��x�j�h��d�    P��  �b3ĉ�$  SUVW�b3�P��$(  d�    ��$8  3ۋ�ω�$0  �|$@�\$褥���   �D$�\$(��$0  �F��T$(RP�AH��;���  �D$(;���  �T$0R�\$4�hpP��Љ\$ �D$0��T$ RP�A Ƅ$8  �ЋD$ ;��D  ��T$<RP�A$��3�9\$<�L$D�#  ��\$�   f�T$X�L$`��f�D$H�T$P�l$X�t$ �>�D$P���ĉ(�l$p�h�H�L$x�H�L$\���ĉ�L$p�H�P�T$x�P�G,VƄ$X  �Ћ5��L$HQ�֍T$XRƄ$4  �֋D$3ɉL$;�t��T$Rh�P��ЋD$�L$3�Ƅ$0  �T$,;�t��T$,Rh�P��ЋD$�L$�T$,;���  �\$4��D$4PQ�J8Ƅ$8  	�ыT$4h 
R� ����  �\$8�5���$�   P�֍�$�   Q�֍�$�   R�֍�$�   P�֋D$��T$8RP�A,Ƅ$8  �Ћ-��|$h�	�Ջ��t$$;��  ��A ��$�   RjVWƄ$@  ��VƄ$4  ���|$h�	�Ջ��t$$;���  ��A ��$�   RjVWƄ$@  ��VƄ$4  ���|$h�	�Ջ��t$$;���  ��A ��$�   RjVWƄ$@  ��VƄ$4  ���|$h�	�Ջ��t$$;��G  ��A ��$�   RjVWƄ$@  �Ћ-�V�վ   3�3҉�$�   ��$�   f��$�   ��$  ��$  f��$   ��$�   Ƅ$0  ;�tP��$�   �Y����L$Ƅ$0  �&3���$�   �\$|f�D$l�L$�D$hǄ$0     j�SP��$  褹���D$t�d$��L$h�  �D$�   ��$0  t�d$���$�   �  ��$�   ;�tP��$�   �ÿ���L$Ƅ$0  �&3ɉ�$�   �\$|f�L$l�L$�D$hǄ$0     j�SP��$�   �����D$t�d$�L$h�  �D$��$0  t�d$���$�   ��  �T$8h�	R� ������$  ��$�   ;�t ���̉d$@P�����?�������$  ���$  ��$�   ;�t ���̉d$@P������������$   ���$   ��$�   Q�L$D�)*  ��$�   ������5���$�   R�֍�$�   P�֍�$�   Q�֍�$�   R�֋D$8P����-��L$4Q�ՋD$�L$�T$,Ƅ$0  ;�t��HR�ыD$�L$Ƅ$0  ;�t��BQ�ЋD$Ƅ$0  ;�t��QP�ҋL$DA;L$<�L$D������|$@�D$ Ƅ$0  ;�t��QP�ҋD$0Ƅ$0  ;�t��QP�ҋD$(��$0  ;�t��QP�ҋǋ�$(  d�    Y_^][��$  3��C  ��   � h �������QV��F��t�L$Q�N�VRQP�R����VR�b9  ���P�F    �F    �F    �B9  ��^Y���̋D$�T$+�V��W�|$��    �49��vQRQW�9  ��_��^� ������������j�h(�d�    P��@SVW�b3�P�D$Pd�    �\$`h�S�@�����<  ���D$$�D$(�D$d�D$|�D$l�D$P�D$4�D$ �D$,�D$0    ����   �t$l�D$PV�p��������   h��L$�6����L$QV�D$`    �sq�����L$���D$X�����	  ��tNh�] j�V�$Ph�V�(�T$4h�R�������xr�@���PV�g������L$4�k	  �D$l�L$h�T$dPQRSW� �L$Pd�    Y_^[��L� ��u�Wj�S�$h�S�`3��L$Pd�    Y_^[��L� ������������̃�0�b3ĉD$,�D$4V�t$<P�D$P�D$    �D$    �D$   �D$ ������h@  �jj j �L$Q�  ��ta�D$�T$Rj j h�  P� ��tD�|$,�D$s�D$�L$(�T$j QPR� ��t�L$j �D$PVjQ� ��t�D$�D$^��tP� �D$��t	j P� �|$(r�T$R�j6  ���L$,�D$3��<@  ��0���������������������������j�h8�d�    P��HSUVW�b3�P�D$\d�    �ى\$�D$t�x- tLj3�h��L$ �D$8   �t$4�D$$ ������D$P�L$8�t$h�t���h,6�L$8Q�D$<��8  �L$p��貆���M �y- t�}��U�z- t����D$t�x�P;�ug�- �uu�w�C9hu�x�9.u�>��~�[9+u�- t���	W�n
  ����D$�X9kux�- t�ƉC�kW蚆�����C�]�A�M �;Eu����- �pu�w�>�M�
�U�B�K9iu�A��M9)u���A�M�H�M,��,;�t�����8],��   �L$�Q;z��   8_,��   �;�ug�F�x, u�X,V�F, �����F�L$�x- uv�8Z,u�P8Z,tc�P8Z,u��Z,P�@, 袻���F�L$�V,�P,�^,�@V�X,�Ɠ���v�x, u�X,V�F, �q�����L$�x- u�P8Z,u�8Z,u�@, �A���v;x�G����1�8Z,u�P�Z,P�@, �h�����L$�V,�P,�^,� V�X,�����_,�}$r�MQ�3  ��3��E$   �E     Uf�U�3  �T$�B����vH�B�D$l�L$t���H�L$\d�    Y_^][��T� �������̋L$����w3�Q��8  ����Ã��3����s�D$P�L$�D$    �4  h|2�L$Q�D$h�N5  �������������V��W�|$��t;t�@8  �F3�;G_����^� ������̋D$�@��t��D$�A��3�� ����̋D$�L$�T$P�D$QRP�2  P�I������������������j�h��d�    P��V�b3�P�D$d�    ��t$�F��PQRQ�D$P���D$0    ��  �NQ�2  �R�F    �F    �2  ���L$d�    Y^�������j�h8�d�    P��   �b3ĉ�$�   SUV�b3�P��$�   d�    ��$�   P��览���L$h�QǄ$�       �����   ��9Xr�@���P�` ��9\$(r�T$R�X1  ��3��D$(   �D$$    f�D$��u9�$�   �Y  ��$�   Q�D  �T$,h�R�X������xr�@���PV�\ �|$D��r�D$0P��0  ����$�   �D$D   �D$@    �D$0 9�$�   s��$�   9�  r���   ����   j j QPj �օ���   ��$�   Q�8H��������   jD�T$Lj R��3  3����D$�D$�D$�D$��$�   �D$HD   9�$�   s��$�   �L$Q�T$LRj j j j j j Pj �X ��t$�D$�5P P�֋L$Q�֍�$�   �  ��9�$�   r��$�   R��/  ��2���$�   d�    Y^][��$�   3��9  �Ĩ   ���U��j�h �d�    P��SVW�b3�P�E�d�    �e����}�E���������v���"�_������������;�s����+�;�w�4�Nj Q�E�    �X��������+�E�e��E@j P�E��;����E���q� Ë}�u�]�M��v$�r�G��G�	RP�D6PS��.  �M���r�OQ��.  �M���G3҉�w�O��r��3�f�H�M�d�    Y_^[��]� �u�~r�FP�.  ��3�Q�F   �F    Qf�N�0  ��������V��~r�FP�G.  ���F   �F    3�f�N^�����̋D$VP����������^� �������j�h��d�    P��D�b3�P�D$Hd�    jh��L$�D$$   �D$     �D$ �����D$P�L$$�D$T    �R���h�5�L$$Q�D$(���/  ����������̋L$��    t�����v�W ���|FSVW�|$�q��L$�D$PQVW3���0  ����|;�wu3�f�w_^��[�3�f�w�z �_^��[�����������̋D$�@��t��D$�A��3�� ����̃�DSU�l$P��   VW��  ���    u�D$\��Q���f��@ �_^][��D� �L$XQhxj3�Vh��t$l���D$X;���  �h   P�Bp�ЋD$X��Qhh   P�ҋD$X����   VP�ҋD$X���  VP�ҋD$X����   VP�ҋD$X����   VP�ҋD$X��T$RP���   �Ѕ�|�L$jhQ�(�D$X�L$�t$��R<QP�ҋD$\��A;�t�T$��D$;�t��QP�ҋ��pH���L$,�T$4�|$X�   f�D$(�\$(�   �D$0�D$ �D$8h�Pƅ�    �L$$�T$,�������xr�@���;�tP������u
h �蟼���T$����ĉ�P�T$0�P�T$4V�P���   W��V���L$8������L$(Q��������  �D$��t�P�B�ЋD$X��t��QP��_^]3�[��D� ����̋D$��y- u�d$ ����y- t������̃�j jj j �D$P�D$    �  ��t�$�L$QjR� �$j P� �L$�D$A3����D$�������������j�h��d�    P��SVW�b3�P�D$d�    ��t$�/���3��`	�F@	�F(	�F��\$ �^�^ �N$�D$ �ۏ���N<�D$ �Ώ���   3��~l�^hf�FX�L$Q�T$R���   �D$(蓲�����   ���   S3�f���   ���   ���   S3�f���   ��  ��  3�Sf���   S���   �p �Fx�^|���   ��  ���   ��  �ƋL$d�    Y_^[����j�h(�d�    P��DSUVW�b3�P�D$Xd�    ���#I�rLj3�h��L$�D$4   �t$0�D$  ������D$P�L$4�t$d�y���h�5�L$4Q�D$8��+  �T$t�G�t$pj RPVP�v����G�   _;�u�h�G�(�O�i�"�|$l t�.�G;0u�(��n�G;pu�h�U�zD �E����   ��$    ��Q;
uQ�R�zD u�YD�ZD��J�AD ��r�   ;qu
��V���v����F�XD�N�Q�BD �F�HQ�������{��zD u�YD�ZD��J�AD ��r�];1u
��V���z����F�XD�N�Q�BD �F�@�H��P��zE u�B�P�Q�W;Bu�J��P;u�
��J��H�N�yD �F�����W�B�XD�D$h��h��L$Xd�    Y_^][��P� ̸  �F6  �b3ĉ�$  ��$  �xV��$  �D$    r�@���h �  �L$QP�\3��F   �F    �D$f�V�P��$    f���f��u�+���P�D$P����!  ��$  ��^3��0  ��  �������������Q�D$��u	�W �Y� �V�T$RhP��D$    �D$    �Ћ���|4�D$��T$R�T$RP�A�Ћ���|�T$�D$�R�T$RP�A�Ћ��D$��t��QP�ҋD$��t��QP�ҋ�^Y� �����������j�hh�d�    P�� VW�b3�P�D$,d�    �L$@3�j�W3�Q�L$�|$�D$4   �|$0f�D$ �!����T$Dj�WR�L$�|$@�\����t$<j�3��F   �~Wf�NP�������|$(r�T$R�U%  ���ƋL$,d�    Y_^��,������j�h�d�    P��|SUVW�b3�P��$�   d�    ��$�   ��$�   3ۉ\$�   3ɉ~�^�t$pf�N�T$RP��$�   �D$    �\$���k��uM�D$;�tEP�L$<襨��j�SP��Ǆ$�      ������$�   9l$Pr�D$<P�$  ���L$Q��j3�h@�L$\�|$t�\$pf�T$`�  j3�h<�L$$Ǆ$�      �|$<�\$8f�D$(�a  V�L$ Q�T$@RƄ$�   �)����L$`QP��$�   RƄ$�   ������j�SP��Ƅ$�   �h���9�$�   r�D$xP��#  ��3ɉ�$�   ��$�   f�L$x9l$Pr�T$<R�#  ��3��|$P�\$Lf�D$<9l$4r�L$ Q�#  ��3҉|$4�\$0f�T$ 9l$lr�D$XP�b#  ���Ƌ�$�   d�    Y_^][�Ĉ   ����������̃�SV��F��W�|$��t;�t	�(  �|$9\$ uf�L$$�^���t;�t	�g(  �|$9\$(uF�N�QR���H>���F�@�F�F    � �F�@�F���D$_^�H�[��� ��$    ��t;|$$t	�(  �|$�\$ ;\$(t�L$�����SW�D$P���  �|$�Ƌ6�D$_�0^�X[��� ��U��$t�����   j�hp�d�    P���b3ŉ��   SVWP�E�d�    �e����   ��E�F�u���u3���N+ȸyxxx��������ڋ��   ����  �N��+V�yxxx��������º���+�;�s�����;��  �������+�;�s3���;�s��j S�A����N�E� �U�R�U�R�VRP�E܉E苅�   PQ�E�    �<���M�� QWP�ΉE��P{���N�E� �U�R�U�R�VRP�E苅�   QP��;���N�V+Ѹyxxx������������t�U�R�FP�FPQ��s���NQ��   ���E܋���Ӎ�����׉N���N�F�d  �U�u܋M�RV��  V�   ��j j ��"  +��   �yxxx���������;���   �M�Q�MD�  ���   �N������ۍRQP���E�   蒆���N�UDR��+��   �yxxx���������+�WQ���E��#z��^�v���   �MDQ+�VR�E�   �c  ���MD�   ���   ������M��Q���R���   �P�   j j �"  �E�P�M ��  �F������P���P+�W���E�   �E��Յ���M싕�   QWR�F�����E P���   �SP��  ���M 胿���M�d�    Y_^[���   3��%)  �Ō   ��]� �����������̋D$��SV��P�L$Q����T���xr�@����PR�$ ���Ã|$ r�D$P��  ��^��[��� �������������S�\$V�t$;�tCW�|$j�j ��D��DV���+���j�j �FP�O�����N8�O8�V<�W<�F@�G@;�uȋ�_^[ËD$^[���������j�h8�d�    P��HSUVW�b3�P�D$\d�    �ى\$�|$t�E tLj3�h��L$ �D$8   �t$4�D$$ ������D$P�L$8�t$h�~��h,6�L$8Q�D$<��>   �L$p�T�����yE t�o��W�zE t����D$t�h�P;�ug�}E �wu�u�C9xu�h�9>u�.��n�[9;u�}E t���	U�1�������D$�X9{uw�}E t�ƉC�jU�M  ���C�\�A��;Gu����}E �pu�u�.�O�
�W�B�K9yu�A��O99u���A�O�H�OD��D;�t�����8_D��   �L$�Q;j��   8]D��   �;�ug�F�xD u�XDV�FD �����F�L$�xE uv�8ZDu�P8ZDtc�P8ZDu��ZDP�@D �6����F�L$�VD�PD�^D�@V�XD�ʠ���v�xD u�XDV�FD ������L$�xE u�P8ZDu�8ZDu�@D �A��v;h�G����1�8ZDu�P�ZDP�@D �l�����L$�VD�PD�^D� V�XD袸���]D�   9o@r�O,Q��  ��3��   3҉_@�w<f�W,9o$r�GP�  ��3ɉ_$�w Wf�O�  �T$�B��;�vH�B�D$l�L$t���H�L$\d�    Y_^][��T� �����������̋D$��SV��P�L$Q���Q���xr�@���j�T$0Rjj P�P�, ���Ã|$ r�L$Q�  ��^��[��� �̋D$V���    ��t��Vh�P�ҋ�^� �����������̋D$�@��t��D$�A<��3�� �����V�t$�~r�FP�  ���F   �F    3�f�N^� ̋T$��    t�����v�W ���|d�L$SV3�W���tE�|$����+�+���    �3��t'�f��tf�����u�_��3�^�z �f�[� ��u���z �_3�^f�[� ����������̃�U�l$VWU���y�����|$��u�6  �S�^�D$��t;�t�  ;�[t*�$�G r����P�EWPj ���S  ��|�L$��N��L$�T$�L$��D$ �I_^��H]��� �j�h��d�    P��  �b3ĉ�$  SUVW�b3�P��$0  d�    ��$@  ��$D  3��D$$3��E   �E�l$(f�M��$8  �D$$   9F��   �~�^r���ÍT$RP�C  ��3�;���   Wj@�D$�D$ �� �~�D$ r�P�D$ WPS�  �t$ �L$Q�T$Rh8V��  ��tF�|$ t?�D$��t7�H�PQ�HR�P
QRh �D$@h�   P��������L$,Q���b  V�� �ŋ�$0  d�    Y_^][��$  3���!  ��(  ��V�t$W�|$�Ƌυ�v�T$S��H����w�[��_^� ���̋L$����w3ɍ�    +���R�B  ����Ã��3����sڍD$P�L$�D$    �v  h|2�L$Q�D$h��  ����������������j�h�d�    PVW�b3�P�D$d�    ��D$P�L$ Q�ο   �����D$�D$    ��t`hP��������t3��K�T$hR���Э����u1�D$h P��軭����u�L$h�Q��覭����t�   ��   �D$�D$������t�P�B�ЋǋL$d�    Y_^��� �������̋D$�@��t��D$�A(��3�� �����Q�T$�$ �$P�D$R�T$��Q�L$PQR誹����� ����V�������D$t	V�  ����^� ��SVW�|$���    ��t�D$9Fw;Fv	�Q  �D$�\$ ���G9^w;^v	�3  �\$ ����t;�t�  �O;�t:�F�D$ �T$R�T$R�T$RQPS������V�؋D$(P�NQRS�\�����(�^��_^[� �������������̋D$�T$U�l$V��L$W�3�j��N�~�VP�G   �G    U��f�G衒���M�T$ �O_�V,�F- ��^]� �������̋D$V���    ��t��VhpP�ҋ�^� �����������̋D$�T$P��Q�L$QR�g����� ��Q�D$V�t$��u;Av`�QSUW;�sP+Ћ�;�wH�   +���Q���T$�L$��r�	�l$�A��    �ǋ��v�M �d$ f9t����u�_]���[^Y� ��t�D$ PUV�H  ����t��+������+���^믃|$r�D$�_��]+�[��^Y� �L$_��]+�[��^Y� �̋��L$��u,�xr�@�L$f�T$f�H� �L$f�T$��f�H� �xr�@����T$W�<P��v�D$�Ћ��������f�_� ����j�h��d�    PVW�b3�P�D$d�    �|$(3��79t$ t���L$d�    Y_^��� h  �  ���D$(�t$;�t	����������HV�D$�����ыD$$��
WPV�ы���BV�ЋǋL$d�    Y_^��� ��������V�t$h�V�@��u#��th�� j�V�$Ph�V�(�^�2�^�����j�h��d�    PQVW�b3�P�D$d�    ��t$�|$ 3�j�P�F   �F    Wf�F趏��3�j��N�GR�A   �A    P�D$$    f�Q苏���ƋL$d�    Y_^��� �����j�h��d�    PQVW�b3�P�D$d�    ��t$�|$ 3�j�P�F   �F    Wf�F�&���3�j��N�GR�A   �A    P�D$$    f�Q������G8�F8�O<�N<�W@�V@�ƋL$d�    Y_^��� ��̋D$�x�Hr�@���Q�L$P�APj ��  3Ʌ������ �������������̋D$�H�yE u�I ���H�yE t�����̋D$�@��t��D$�A0��3�� �����V�t$��W�x��I f���f��u�+���PV��  _^� ����̃�SV��^W��u3���N+˸yxxx��������ʋ~��+Ӹyxxx���������;�s2�T$�D$ �L$Q�L$R�FPQjW�w������D�~_^[��� ;�v�  �T$�RWP�D$P���kd��_^[��� �̋D$��u�W ��$ �L$�������	wd��� �$�� �L$�Q����P�BQ���$ �L$�Q����P�BQ���$ �L$�Q����P�B Q���$ V�t$�NtQ�T j �N��n���^3��$ �� �� �� �� �  ����������j�h�d�    P��  �b3ĉ�$�  SUVW�b3�P��$�  d�    ��$�  h  ��$�  PV�| ���   ���  ��$�   Q�T$Th�R�������   Ǆ$�      9hr�@������̉d$4P蔒���  �� ����Ǆ$�  ����9l$hr�D$TP�u  ������  ��$�   Q�T$pR�����D$Xh�PǄ$�     �u�����Ƅ$�  9hr�@���P��$�   �����   �L$P��$�  �����L$4h�Q�,����L$x��9�$�   s�L$p9hr�@���QP��$�   h  R�7������L$4�[�����$�   9�$�   s��$�   ��$�   �=�	RPjh���$�   Ph   ��׍L$4h�Q�����L$x��9�$�   s�L$p9hr�@���QP��$�   h  R�������L$4�������$�  �P��f���f��u�+����D P��$�  Qjh���$�   Rh   ��׍D$h�P�������L$<hlQƄ$�  �������9nr�v���9hr�@���jVjP��$�   Rh   ��׍L$4�+����L$��$�  �����D$h�P�����L$x��9�$�   s�L$p9hr�@���QP��$�   h  Q�������L$������T$h�R�L�����9hr�@���Sh�jP��$�   Ph  ��׍L$������$�   �����L$l�v���3���@ ���$�  d�    Y_^][��$�  3��  ���  ������U�l$V�t$;�t=SW�|$�_j�j W�������j�j S�N������G8�F8�O<�N<�W@�V@��D;�u�_[^]��̃�SUV��FW�~��+�������u3��%;�v�  �L$ ���t;�t�|  �\$$+����T$(�D$$�L$ RjPQ���tR���~;~v�N  �6��|$��u�=  3��<�;xw��t�6����3�;~s�  �D$�x_^�(][��� ̃�dSUV�t$t��   �FW�9  �T$R3��|$�h�P��ЋF�L$;���   �T$|�9J��   �T$x�|$x�RP�AH�ЋD$x;���   P�L$��x���D$;���   ��NQP�B�ЋL$xQ�L$�3����D$;�tQ�L$|�|$|��RQP��9|$|t*�D$|P�N �7����L$|Q�N��  �D$|;�t�P�B�ЋD$;�t��QP�ҋD$;�t��QP�ҍN$��#���N<��#����賱���D$x;�t��QP�ҋD$;��  ;���  �Q�H��3�_^][��d� �D$x    ���O  ���L$xQh�P�҃~ �D$x�`  �L$|�9B�Q  �D$HP���~�L$,h�Q�!������xr�@���P��$�   �3���� ��L$HQ���   PW�ыT$|R���L$,�L����|$P��   �L$(�\$ �~�   f�D$�l$3��T$Xh�R�D$,�D$<�L$@�������xr�@���P��$�   譧��� ����̉)�Y�\$D�Y�\$HP�Y���   W�ыT$|R���L$X�����D$P���F����   j�P�ҍD$HP���v�L$�D$    ����   QV�ҋD$��t	P�������D$x��t��QP��_^]3�[��d� �����VW�����u��  ���t��3ҋD$������G���;Bw��t�	�3�;As�  w��_^� ��������������VW�����u�  ���t��3ҋD$�4�    +��G���;Bw��t�	�3�;As�]  w��_^� ������������VW�|$�P����a����u2���u_3�^� �>�    ��t��Vh�P�҅�t��HW�ы_^� ���j�h��d�    P��4�b3ĉD$0V�b3�P�D$<d�    �t$h�D$P�D$H    諗����jhT�L$�D$L�Cg��j�j �L$TQ�L$��q���T$$R�D$P��������ta�L$$�T$(�D$,��L$0�V�F�N�   9t$ r�T$R��  ��3��D$    �D$    f�D$9t$dr�L$PQ�  ����D�   9t$ r�T$R�  ��3��D$    �D$    f�D$9t$dr�L$PQ�d  ��2��L$<d�    Y^�L$03��+  ��@�����������SU�l$VW��9os��  �G�t$+�;�s���\$ ��;�r�Ãr����P�D$ P�oQ�  ����u;�s
_^]���[� 3�;���_^][� �SV��L$W��tI�~�F��r����;�r4��r���Ћ^�Z;�v��r� �T$+�R��QV��� ���_^[� �|$�����v��  �F;�s!�FPW��������vg�NU�n��r1�E �.��u�~��r�F3�_f���^[� �F3�_f���^[� �ŋT$�?SR�QP�  ���~�~r�m 3�f�+]_��^[� ��̋T$V��v�L$�D$f�0f;1u������u�3�^�� f;^����@����������̋L$�T$�   V���2;1u��������s�3�3҅���^�����1+�u"�B�q+�u�B�q+�u
�B�I+�����3҅���^����̃��$h�P�O������xr�@���VPjj �� �|$��r�L$Q��  ��h�  3�V�D$$   �D$     f�T$�h =  t<�T��jj ����|)h  �7  ����t���7�����t���=������tV�P 3�^�������3�9Dt������̡@tP�������T��3�������������K����V���3����̸   9D$u
�L$�@t� �������̃�<�b3ĉD$8�Pt�D$DS�\$D�D$�D$LVW�D$�D$    u�Pt�Ht��Lt    �L$h�Q�     �ڼ�����xr�p��p�T$4R����3��A   �A    f�A�Ɖd$,�x��f���f��u�+���PV����������� ��t�L$4QS��������t��2ۃ|$0r�T$R�  ����tq�t$h�V�o�������u+h�V�]�������u�@ �_^[�L$83���
  ��<� �D$� Ht�Ht�QhHt��3�_^[�L$83��
  ��<� �L$D_^[3̸��w
  ��<� �%��%��%�jD����  h��M��\���e� �E�P�M��I\��h�5�E�P�  �jD����y  h�M��Q\���e� �E�P�M��Qt��h,6�E�P�d  ̋�U��]�  ��U��]�  ��U��V�uW3�;�u3��e9}u�R  j^�0WWWWW�  �����E9}t9urV�u�u�"
  �����uW�u�1  ��9}t�9us�  j"Y����jX_^]Ë�U��EVW3�;�tG9}u��  j^�0WWWWW�  �����)9}t�9Es�  j"Y�����P�u�u��  ��3�_^]Ë��` �` � $Ë�U��S�]VW���$���t&P�  ��FV��  YY�G��t�3VP��  ����g �G   ��_^[]� ��U����M� $�	�` �H]� ��U��S�]V���$�C�F���CWt1��t'P�'  ��GW�J  YY�F��t�sWP�  ���	�f ��F_��^[]� �y �$t	�q��  YËA��u�,Ë�U��V��������EtV����Y��^]� ��Q�D�  YË�U��V��������EtV�����Y��^]� ��U��E��	Q��	P��  ��Y�Y@]� ��U��� �EVWjY�H�}��E��E_�E�^��t� t�E� @��E�P�u��u��u����� ��U��� S3�9]u ��  SSSSS�    �  ������   �EV�u;�t!;�u�  SSSSS�    �P  ������t�E�B   �u�u�=���?v	�E�������E�W�u�E��u�uP�  ����;�t5�M�x
�E���E���E�PS�X  YY�M�x�E����E�PS�@  YY��_^[�Ë�U���uj �u�u�u������]��̋T$�L$��ti3��D$��u��   r�=x� t��$  W����r1�ك�t+ш����u������������ʃ���t��t
�����u��D$_ËD$Ë�U��E�Tt]Ë�U���(  �b3ŉE������� SjL������j P�J�����������(�����0�������,���������������������������������������f������f������f������f������f������f��������������E�Mǅ0���  �������������I�������ǅ���� �ǅ����   ��������j ������(���P����u��uj��$  Yh ���P���M�3�[�  �Ë�U���5Tt�#%  Y��t]��j�$  Y]����3�PPPPP�������Ë�Vjh b�������h��^Ë�U�����u�+  Y��t�u�+  Y��t����dt�Xtu�dt������h*��P+  YV�M��l��h|2�E�P�[���̋�U��QS�E���E�d�    �d�    �E�]�m��c���[�� XY�$����U��QQSVWd�5    �u��E��	j �u�u��u���  �E�@����M�Ad�=    �]��;d�    _^[�� U���SVW��E�3�PPP�u��u�u�u�u�6  �� �E�_^[�E���]Ë�U��V��u�N3��  j V�v�vj �u�v�u�h6  �� ^]Ë�U���8S�}#  u��M�3�@�   �e� �E�D�b�M�3��E��E�E�E�E�E�E�E �E��e� �e� �e� �e�m�d�    �E؍E�d�    �E�   �E�E̋E�E��F%  ���   �EԍE�P�E�0�U�YY�e� �}� td�    ��]؉d�    �	�E�d�    �E�[�Ë�U��QS��E�H3M�  �E�@��ft�E�@$   3�@�l�jj�E�p�E�p�E�pj �u�E�p�u�25  �� �E�x$ u�u�u�����j j j j j �E�Ph#  �������E��]�c�k ��3�@[�Ë�U��QSVW�}�G�w�E����-���u��5  �M�N��k���M9H};H~���u	�M�]�u�} }ʋEF�0�E�;_w;�v�5  ��k�E�_^[�Ë�U��EV�u���#  ���   �F��#  ���   ��^]Ë�U���#  ���   �
�;Mt
�@��u�@]�3�]Ë�U��V�#  �u;��   u�}#  �N���   ^]��l#  ���   �	�H;�t���x u�^]�5  �N�H�ҋ�U����b�e� �M�3��M�E��E�E�E@�E�:
�M��E�d�    �E�E�d�    �uQ�u�5  �ȋE�d�    ����;bu���05  øZN��c��cAE��c�D��c.E��c�D��c��c�M��c�D��cD��c�CË�U�������+A  �} �ltt�@  ��]�U��WV�u�M�}�����;�v;���  ��   r�=x� tWV����;�^_u^_]�A  ��   u������r*��$�d��Ǻ   ��r����$�x�$�t��$������#ъ��F�G�F���G������r���$�d�I #ъ��F���G������r���$�d�#ъ���������r���$�d�I [H@80( �D��D��D��D��D��D��D���D���D��D��D���D���D���D����    ���$�d��t|���E^_�Ð���E^_�Ð���F�G�E^_�ÍI ���F�G�F�G�E^_�Ð�t1��|9���   u$������r����$� �����$���I �Ǻ   ��r��+��$��$� �8`�F#шG��������r�����$� �I �F#шG�F���G������r�����$� ��F#шG�F�G�F���G�������V�������$� �I ���������D��D��D��D��D��D��D��D��D��D��D��D��D��D���    ���$� ��(<�E^_�Ð�F�G�E^_�ÍI �F�G�F�G�E^_�Ð�F�G�F�G�F�G�E^_���5�z�  Y��t��j�d@  jj �:@  ���?  �SV�D$�u�L$�D$3���؋D$����A�ȋ\$�T$�D$���������u�����d$�ȋD$���r;T$wr;D$vN3ҋ�^[� ��U��j
j �u��C  ��]Ë�U��]�������U��EV���F ��uc�"  �F�Hl��Hh�N�;�jt��i�Hpu�3M  ��F;�ht�F��i�Hpu�E  �F�F�@pu�Hp�F�
���@�F��^]� Q�L$+����#ȋ�% ���;�r
��Y�� �$�-   � ���U��QSV��3�;�u�$  j^SSSSS�0�����������   W9]w�   j^SSSSS�0���������   3�9]f���@9Ew	��  j"�ϋE�����"w��]���9]t�]j-Xf��N�E�   ���E3��u�E��	v��W���0�E�f�AA@3ۉE�9]v;Er�;Er3�f��3�f�IIf��f�If�IGG;�r�3�_^[�� ��U��}
u�} }jj
�j �u�u�E�u�����]Ë�U��EVW��u|P�mX  Y��u3��  ��  ��u�X  ��� X  ���|��V  �tt��P  ��}�m  ����U  ��| �cS  ��|j �N  Y��u�pt�   ��R  ��3�;�u19=pt~��pt9=`{u�!P  9}u{��R  �  ��W  �j��uY��  h  j�L  ��YY;��6���V�5�c�5�t�!  Y�Ѕ�tWV��  YY���N���V�-  Y�������uW�  Y3�@_^]� jh@I�fY  ����]3�@�E��u9pt��   �e� ;�t��u.�t��tWVS�ЉE�}� ��   WVS�r����E����   WVS������E��u$��u WPS����Wj S�B����t��tWj S�Ѕ�t��u&WVS�"�����u!E�}� t�t��tWVS�ЉE��E������E���E��	PQ�pX  YYËe��E�����3���X  Ë�U��}u�TZ  �u�M�U�����Y]� ����̋L$��   t$�����tN��   u�    ��$    ��$    �����~Ѓ��3�� �t�A���t2��t$�  � t�   �t�͍A��L$+�ÍA��L$+�ÍA��L$+�ÍA��L$+��Pd�5    �D$+d$SVW�(��b3�P�u��E������E�d�    �Pd�5    �D$+d$SVW�(��b3�P�e��u��E������E�d�    �jh`I�TW  �u��tu�=<�uCj�7[  Y�e� V�_[  Y�E��t	VP�[  YY�E������   �}� u7�u�
j�#Z  Y�Vj �5t|����u�Y   ����P�	   �Y�W  Ë�U��E3�;� btA��-r�H��wjX]Ë�$b]�D���jY;��#���]���  ��u��cÃ���  ��u��cÃ�Ë�U��V������MQ�����Y�������0^]����U��WV�u�M�}�����;�v;���  ��   r�=x� tWV����;�^_u^_]�07  ��   u������r*��$����Ǻ   ��r����$���$����$�H��(#ъ��F�G�F���G������r���$���I #ъ��F���G������r���$���#ъ���������r���$���I �����xph�D��D��D��D��D��D��D���D���D��D��D���D���D���D����    ���$���������E^_�Ð���E^_�Ð���F�G�E^_�ÍI ���F�G�F�G�E^_�Ð�t1��|9���   u$������r����$�P�����$� �I �Ǻ   ��r��+��$�T�$�P�d���F#шG��������r�����$�P�I �F#шG�F���G������r�����$�P��F#шG�F�G�F���G�������V�������$�P�I $,4G�D��D��D��D��D��D��D��D��D��D��D��D��D��D���    ���$�P��`hx��E^_�Ð�F�G�E^_�ÍI �F�G�F�G�E^_�Ð�F�G�F�G�F�G�E^_�Ë�U��MS3�VW;�t�};�w�2���j^�0SSSSS����������0�u;�u��ڋъ�BF:�tOu�;�u������j"Y�����3�_^[]�jh�I�kR  �e� �u;5,�w"j�OV  Y�e� V�V^  Y�E��E������	   �E��wR  �j�JU  YË�U��V�u�����   SW�=��=t| u��6  j�G5  h�   ��E  YY�<���u��t���3�@P���uV�S���Y��u��uF�����Vj �5t|�׋؅�u.j^9�}t�u��  Y��t�u�{���������0������0_��[�V�  Y������    3�^]�jh�I�RQ  j�EU  Y�e� �u�N��t/��t��t�E��t9u,�H�JP����Y�v����Y�f �E������
   �AQ  Ë���j�T  Y����������̋T$�L$��   u<�:u.
�t&:au%
�t��:Au
�t:au����
�uҋ�3�Ð��������   t���:u��
�t���   t�f���:u�
�t�:au�
�t���눋�U��QV�uV�l  �E�FY��u����� 	   �N ����/  �@t����� "   ��S3ۨt�^���   �N�����F�F�����F�^�]��  u,�j  �� ;�t�sj  ��@;�u�u� j  Y��uV�i  Y�F  W��   �F�>�H��N+�I;��N~WP�u�h  ���E��M�� �F����y�M���t���t�����������`����j�@ tjSSQ�	`  #����t%�F�M��3�GW�EP�u�1h  ���E�9}�t	�N �����E%�   _[^�Ë�U���@@t�x tP�u�fk  YY���  f;�u��]��]Ë�U��V����u�E�M�����>�Yt�} �^]Ë�U���G@SV����t7� u1�E�0��MP���~���CC�>�Yu������8*uj?���c���Y�} �^[]Ë�U���t  �b3ŉE��ES�]V�uW�u3��������������������������������������������������������������n���9�����u3�L���WWWW�    W�	����������� t
�������`p������
  ;�t��3ɉ�����������������������f;���
  j_������� �������i
  �B�f��Xw����H ���3����h j��Y������;���	  �$��+3���������������������������������������������	  �� tJ��t6��t%+�t����	  �������	  �������	  �������y	  �������   �j	  	������_	  f��*u,���������[����������?	  �������������-	  ������k�
�ʍDЉ������	  ������ �	  f��*u&���������[�����������  ���������  ������k�
�ʍDЉ������  ��ItW��htF��lt��w��  ������   �  f�>lu�������   �������x  �������l  ������ �`  �f��6uf�~4u�������� �  �������8  f��3uf�~2u������������������  f��d�	  f��i��  f��o��  f��u��  f��x��  f��X��  ������ ������R������ǅ����   ������  ��d�/  ��  ��S�  t~��At+�tY+�t+���  �� ǅ����   ������������@������ �������   ��������������  ǅ����   ��  ������0  ��   ������ �   ������0  u������ ���������u������������ �������[��������  ��u��n������������ ���������   ����  ��������QP�+i  YY��tFF������9�����|���  ��X��  +���   +������+���  ���3�F������ ������������������tB������������P������ƅ���� ���   ������P������P�gg  ����}�������f�������������������������F  �����������t:�H��t3������   � ������t�+�ǅ����   �  ������ ��  ��n������P�g���Y��  ��p��  ��  ��e��  ��g�������itq��nt(��o��  �������ǅ����   ta������   �U�3���������af  ���0  ������ tf������f���������ǅ����   ��  ������@ǅ����
   ������ �  ��  ��S����  uf��gucǅ����   �W9�����~�������������   ~=��������]  W�A:  ������Y��������t���������������
ǅ�����   ����������C�������������P��������������������P������������VP�5�c�  Y�Ћ���������   t!������ u������PV�5�c�{  Y��YYf������gu��u������PV�5�c�U  Y��YY�>-u������   F������V����ǅ����   �������$��s�g���+����������  ǅ����'   �������ǅ����   �j���j0Xf��������������Qf�������������E���������   �E����������� t������@������t�C���C���������@�C�t��3҉�����������@t��|��s�؃� �ځ�����   ������ �  �ڋ�u3ۃ����� }ǅ����   ���������   9�����~���������u!����������������������������t-�������RPSW�b7  ��0��9����������~������N뽍�����+�F������   ������������tY��t�΀90tN�������������0@�6��u��n������������ǅ����   �	Of�8 t@@��u�+������������������� �e  �������@t+�   tj-��tj+��tj Xf������ǅ����   ������������+�+�����������u������������Sj ����������������������������������������Yt������uWSj0�������Q����������� uu��~q������������������������P���������   ������WP��a  ����������~)��������������������������������� Y����������������V�����������Y������ | ������t������������Sj ������������ t����������������� Y�������������f��t*�����������������������    3�PPPPP�2��������� t
�������`p��������M�_^3�[�����ÍI s#U!�!�!1"="�"�#U����}��}�M��f�����$    �ffGfG fG0fG@fGPfG`fGp���   IuЋ}���]�U����}��E���3�+���3�+���u<�M�у��U�;�t+�QP�s������E�U��tEE+E�3��}��M��E�.�߃��}�3��}�M��E��M�U�+�Rj Q�~������E�}���]�jh�I��A  �e� f(��E�   �#�E� � =  �t
=  �t3��3�@Ëe�e� �E������E���A  Ë�U���3�S�E��E�E�S�X��5    P��Z+�tQ�3���E�]�U�M�   ��U��E�[�E�   t�\�����t3�@�3�[�������x�3�Ã%t� Ë�U��V�5�c�5��օ�t!��c���tP�5�c���Ѕ�t���  �'��V����uV�,4  Y��thxP�\ ��t�u�ЉE�E^]�j ����YË�U��V�5�c�5��օ�t!��c���tP�5�c���Ѕ�t���  �'��V����uV�3  Y��th�P�\ ��t�u�ЉE�E^]���� ��V�5�c������u�5�t�e���Y��V�5�c�|��^á�c���tP�5�t�;���Y�Ѓ�c���c���tP�x��c��mB  jh�I�?  ��V����uV��2  Y�E�u�F\�3�G�~��t$hxP�\ �Ӊ��  h��u��Ӊ��  �~pƆ�   CƆK  C�Fh�dj�!C  Y�e� �vh�� �E������>   j� C  Y�}��E�Fl��u��j�Fl�vl�z.  Y�E������   �?  �3�G�uj��A  Y�j��A  Y���̋�VW���5�c�������Ћ���uNh  j�e1  ��YY��t:V�5�c�5�t�����Y�Ѕ�tj V�����YY���N���	V�����Y3�W�t_��^Ë�V��������uj��1  Y��^�jhJ�>  �u����   �F$��tP����Y�F,��tP����Y�F4��tP����Y�F<��tP�y���Y�F@��tP�k���Y�FD��tP�]���Y�FH��tP�O���Y�F\=�tP�>���Yj�A  Y�e� �~h��tW�� ��u���dtW����Y�E������W   j�WA  Y�E�   �~l��t#W�i-  Y;=�jt���it�? uW�u+  Y�E������   V����Y�X=  � �uj�&@  YËuj�@  YË�U��=�c�tK�} u'V�5�c�5��օ�t�5�c�5�c���ЉE^j �5�c�5�t����Y���u�x�����c���t	j P�|]Ë�VW��V����uV��/  Y�����^  �5\ h�W��h�W��t��h�W��t��h�W��t�փ=�t �5|��tt�=�t t�=�t t��u$����t�x��tf.�5�t��t����c�����   �5�tP�օ���   ��1  �5�t�����5�t��t�����5�t��t�����5�t��t�r�������t��=  ��teh]0�5�t�����Y�У�c���tHh  j�.  ��YY��t4V�5�c�5�t����Y�Ѕ�tj V�v���YY���N��3�@��!���3�_^Ë�U��QSVW�5h��Y����5d����}��I�����YY;���   ��+ߍC��rwW�\Z  ���CY;�sH�   ;�s���;�rP�u��-  YY��u�G;�r@P�u��-  YY��t1��P�4��d���Y�h��u�V������V�K���Y�d��EY�3�_^[�Ë�Vjj �-  ��V�$������h��d���ujX^Ã& 3�^�jh0J�:  �.  �e� �u�����Y�E��E������	   �E��":  ���-  Ë�U���u���������YH]Ë�U��E��t]Ë�U���5�t����Y��t�u��Y��t3�@]�3�]Ë�U��V�EP���b�������^]� ��������U��V���������EtV�5���Y��^]� ��U��VW�}�G��tG�P�: t?�u�N;�t��QR�'���YY��t3��$�t�t�E� �t�t�t�t�3�@_^]Ë�U��E� � =MOC�t=csm�u+�y������    ��  �h������    ~�Z����   �3�]�jhPJ�8  �}�]��   �s��s�u��#����   � �e� ;ute���~;w|��  �����Oȋ1�u��E�   �y t�sh  S�O�t��  �e� ��u��-���YËe�e� �}�]�u��u���E������   ;ut�V  �s�8  Ë]�u��������    ~�v����   �Ë �8csm�u8�xu2�H�� �t��!�t��"�u�x u�8���3�A��  ���3��jhxJ�^7  �M��t*�9csm�u"�A��t�@��t�e� P�q�Y����E������m7  �3�8E��Ëe��G
  ̋�U��M�V�uƃy |�Q�I�42���^]Ë�U�����u
�X
  �
  �e� �? �E� ~SSV�E�@�@��p��~3�E����E�M�q�P�GE�P�_�������u
K�������E��E��E�;|�^[�E���j��������������    t��	  �e� �	  �M���q	  ������Mj j ���   �v����j,h�J�6  �ً}�u�]�e� �G��E��v�E�P�����YY�E��������   �E��������   �E��������   �����M���   �e� 3�@�E�E��u�uS�uW�������E�e� �o�E������Ëe��F�����   �u�}�~�   �O��O�^�e� �E�;Fsk�ËP;�~@;H;�F�L�QVj W�������e� �e� �u�E������E    �   �E��S5  ��E�맋}�u�E܉G��u�����Y�����Mԉ��   �����MЉ��   �>csm�uB�~u<�F= �t=!�t="�u$�}� u�}� t�v����Y��t�uV�%���YY�jhK�4  3҉U�E�H;��X  8Q�O  �H;�u�    ��<  � �u��x�t1�U�3�CS�tA�}�w�rT  YY����   SV�aT  YY����   �G��M��QP�����YY���   �}�E�p�tH�*T  YY����   SV�T  YY����   �w�E�pV�x��������   ���t|��W�9Wu8��S  YY��taSV��S  YY��tT�w��W�E�p�_���YYPV�'������9�S  YY��t)SV�S  YY��t�w�S  Y��t�j X��@�E���  �E������E��3�@Ëe��F  3��S3  �jh8K�3  �E�    �t�]�
�H�U�\�e� �uVP�u�}W�F�����HtHu4j�FP�w����YYP�vS�������FP�w����YYP�vS�����E�������2  �3�@Ëe��  ̋�U��} t�uSV�u�V������}  �uuV��u �x����7�u�uV�����Gh   �u@�u�F�u�KV�u�������(��tVP����]Ë�U��QQV�u�>  ���   W�������    t?�������   �>���9t+�>MOC�t#�u$�u �u�u�u�uV����������   �}� u�  �u�E�P�E�PV�u W��������E���;E�s[S;7|G;wB�G�O����H��t�y u*�X��@u"�u$�u�u j �u�u�u�u�����u���E��E���;E�r�[_^�Ë�U���,�MS�]�C=�   VW�E� �I��I����M�|;�|�]  �u�csm�9>��  �~� ��  �F;�t=!�t="���   �~ ��   �X������    ��  �F������   �u�8������   jV�E�P  YY��u��  9>u&�~u �F;�t=!�t="�u�~ u�  ��������    t|��������   ������u3����   ����Y��uO3�9~�G�Lh�c������uF��;7|��	  j�u�d���YYh��M��7���hTK�E�P������u�csm�9>��  �~�~  �F;�t=!�t="��e  �}� ��   �E�P�E�P�u��u W���������E�;E���   �E�9��   ;G|�G�E�G�E��~l�F�@�X� �E��~#�v�P�u�E����������u�M��9E���M�E��}� ��(�u$�]��u �E��u��u�u�uV�u�K����u���E����]����}�} t
jV�:���YY�}� ��   �%���=!���   �����   V����Y����   �&����!����������   �����}$ �M���   Vu�u��u$�a����uj�V�u�u�������v�����]�{ v&�} �)����u$�u �u�S�u�u�uV������� �������    t�T  _^[�Ë�U��V�u����������^]� ��U��SVW�g�����   �E�M�csm�����"�u �;�t��&  �t�#�;�r
�@ ��   �Aft#�x ��   �} u}j�P�u�u�������j�x u�#ց�!�rX�x tR99u2�yr,9Yv'�Q�R��t�u$V�u �uP�u�u�uQ�҃� ��u �u�u$P�u�u�uQ������� 3�@_^[]�jh�K��,  �}����@x��t�e� ���3�@Ëe��E������  ��,  ��P����@|��t������jh�K�w,  �5�t�����Y��t�e� ���3�@Ëe��E������}����h�A�6���Y��t�������U���SQ�E���E��EU�u�M�m��uM  VW��_^��]�MU���   u�   Q�SM  ]Y[�� ��U���(  ��u��u��u��u�5�u�=�uf��uf��uf��uf��uf�%�uf�-�u���u�E ��u�E��u�E��u������� u  ��u��t��t	 ���t   �b�������b����������tj����Yj ��h ���=�t uj�����Yh	 ���P���Ë�U���V�u�M��S����u�P�N  ��e�F�P��L  ��Yu��P�N  Y��xuFF�M����   �	��	�F�����F��u�^8M�t�E��`p��Ë�U���V�u�M�������E��u���t���   ��:�t@���u��@��t6���et��Et@���u��H�80t����   �	S�:[uH�
@B���u��}� ^t�E��`p��Ë�U����E�����Az3�@]�3�]Ë�U��QQ�} �u�ut�E�P�>M  �M��E��M��H��EP��M  �E�M����Ë�U��j �u�u�u������]Ë�V����tV����@PV�V������^Ë�U��j �u�e���YY]Ë�U��j �u�����YY]Ë�U���SVW�u�M�������3�;�u+�}���j_VVVVV�8�;������}� t�E��`p����!  9uv�9u~�E�3���	9Ew	�9���j"뺀} t�U3�9u��3Ƀ:-����ˋ��,����}�?-��u�-�s�} ~�F�����E����   � � �3�8E��E��}�u����+�]hSV�k�����3ۅ�tSSSSS�L������N9]t�E�GF�80t.�GHy���-F��d|
�jd_�� ��F��
|
�j
_�� �� F�~t�90uj�APQ�������}� t�E��`p�3�_^[�Ë�U���,�b3ŉE��ESVW�}j^V�M�Q�M�Q�p�0��M  3ۃ�;�u�����SSSSS�0���������o�E;�v�u���u����3Ƀ}�-��+�3�;���+��M�Q�NQP3��}�-��3�;�����Q��K  ��;�t���u�E�SP�u��V�u��������M�_^3�[������Ë�U��j �u�u�u�u�u������]Ë�U���$VW�u�M��E��  3��E�0   �1���9}}�}�u;�u+����j^WWWWW�0��������}� t�E�`p����  9}vЋE��� 9Ew	�����j"���}��E�G������  S#�3�;���   ����   �E���u�����j �u�^PSW��������t�}� � ��  �M�ap��  �;-u�-F�0F�} je����$�x�FV�dG  YY���L  �} ���ɀ����p��@ �2  %   �3��t�-F�]�0F������$�x��OF��ۃ����  �3���'3��u!�0�O����� F�u�U���E��  ��1F��F�E9Uu���M܋��   �	�	��O����� �M�w;���   �U��E�   �} ~M�W#U���M�#E���� �L  f��0��f��9vËM��m���E�����F�Mf�}� �E�M�}�f�}� |Q�W#U���M�#E���� �XL  f��v1�F����ft��Fu� 0H��;Et���9u��:��	�����@��} ~�uj0V�м����u�E�8 u���} �4����$�p���WF��K  3�%�  #�+E�SY�x;�r�+F�
�-F�����;Ӌ��0|$��  ;�rSQRP�J  0�F�U�����;�u��|��drj jdRP�J  0��U�F����;�u��|��
rj j
RP�sJ  0��U�F���]�0��F �}� t�E�`p�3�[_^�Ë�U���SVW�u�؋s���M�N�������u-����j^�03�PPPPP�c������}� t�E��`p����   �} v̀} t;uu3��;-����� 0�@ �;-��u�-�w�C3�G�����X����0F���} ~D���C����E����   � � ��[F��}&�ۀ} u9]|�]�}������Wj0V�
������}� t�E��`p�3�_^[�Ë�U���,�b3ŉE��ESVW�}j^V�M�Q�M�Q�p�0�H  3ۃ�;�u����SSSSS�0�Y��������Z�E;�v���u��3Ƀ}�-��+��u�M�Q�M��QP3��}�-���P�F  ��;�t���u�E�SV�u���`������M�_^3�[�����Ë�U���0�b3ŉE��ESV�uWj_W�M�Q�M�Q�p�0��G  3ۃ�;�u�����SSSSS�8螻�������   �M;�vދE�H�E�3��}�-���<0���u��+ȍE�P�uQW��E  ��;�t��X�E�H9E������|-;E}(:�t
�G��u��_��u�E�j�u���u��������u�E�jP�u���u�u�������M�_^3�[荿���Ë�U��E��et_��EtZ��fu�u �u�u�u�u� �����]Ã�at��At�u �u�u�u�u�u�����0�u �u�u�u�u�u�w�����u �u�u�u�u�u�n�����]Ë�U��j �u�u�u�u�u�u�Z�����]Ë�VW3����c�6�������Y���(r�_^Ë�Vh   h   3�V��G  ����tVVVVV�ո����^Ë�U�����]���]��E��u��M��m��]����]�����z3�@��3���h<�p��th P�\ ��tj �������U����}��u��u�}�M�����    fofoNfoV fo^0ffOfW f_0fof@fonPfov`fo~pfg@foPfw`fp���   ���   Iu��u��}���]�U����}�u��]��]�Ù�ȋE3�+ʃ�3�+ʙ��3�+���3�+����uJ�u�΃��M�;�t+�VSP�'������E�M��tw�]�U�+щU��+ى]��u�}��M��E�S;�u5�ك��M�u�}�M��MM�UU�E+E�PRQ�L������E��u�}�M�����ʃ��E�]��u��}��]Ë�U���(  �b3ŉE���cVtj
�  Y�sF  ��tj�uF  Y��c��   ������������������������������������f������f������f������f������f������f��������������u�E������ǅ0���  �������@�jP������������j P觵������������(�����0���j ǅ����  @��������,�������(���P��j��  ̋�U��M��c�U#U��#�ʉ�c]Ë�U��QQS�]VW3�3��}�;� dt	G�}���r���w  j�I  Y���4  j�oI  Y��u�=�t�  ���   �A  h��  S��wW�X�������tVVVVV�;�����h  ��wVj ��x �d��u&h�h�  V��������t3�PPPPP�������V����@Y��<v8V�x�����;�j��zh�+�QP�H  ����t3�VVVVV贴�����3�h�SW�gG  ����tVVVVV萴�����E��4�dSW�BG  ����tVVVVV�k�����h  h�W�E  ���2j��h��;�t$���tj �E�P�4�d�6�����YP�6S�l_^[��j�H  Y��tj��G  Y��u�=�tuh�   �)���h�   ����YYË�U��E��z]Ë�U���SW�u�M��/����E�}3�;�t�8;�u+����SSSSS�    �������8]�t�E��`p�3��  9]t�}|ʃ}$�V�7�]�����7GG�E�PjV�  ����u�f��-u�M�f��+u�7GG9]u3V�G  Y��t	�E
   �F�f��xtf��Xt	�E   �.�E   �}u!V�LG  Y��u�f��xtf��XuGG�7GG���3��u�U���V�G  Y���u)jAXf;�wf��Zv	�F�f��w1�F�f����w�� ���;Es�M9]�r)u;E�v"�M�} u$�EOO�u"�} t�}�e� �]�M��MȉM��7GG끾����u�u=��t	�}�   �w	��u+9u�v&�}����E� "   t�M����Ej X��ƉE��E^��t�8�Et�]��}� t�E��`p��E�_[�Ë�U��3�P�u�u�u9{uh�j�P�������]�-�  t"��t��tHt3�ø  ø  ø  ø  Ë�VW��h  3��FWP����3��ȋ��~�~�~����~�����d���F+ο  ��@Ou���  �   ��@Nu�_^Ë�U���  �b3ŉE�SW������P�v�`�   ����   3�������@;�r�����ƅ���� ��t.���������;�w+�@P������j R������C�C��u�j �v�������vPW������Pjj �L  3�S�v������WPW������PW�vS�kJ  ��DS�v������WPW������Ph   �vS�FJ  ��$3���E������t�L���������t�L ��������  �Ƅ   @;�r��V��  ǅ��������3�)�������������  ЍZ ��w�L�р� ���w�L �р� ���  A;�rM�_3�[�O�����jh�K�h  �"�������i�Gpt�l t�wh��uj ��	  Y���  �j�-  Y�e� �wh�u�;5�ht6��tV�� ��u���dtV裾��Y��h�Gh�5�h�u�V�� �E������   뎋u�j��  YË�U���S3�S�M��A�����z���u��z   �88]�tE�M��ap��<���u��z   �<�ۃ��u�E��@��z   ��8]�t�E��`p���[�Ë�U��� �b3ŉE�S�]V�uW�d�����3��};�u������3��  �u�3�9��h��   �E��0=�   r����  �p  ����  �d  ��P�4���R  �E�PW�`���3  h  �CVP�=���3�B���{�s9U���   �}� ��   �u�����   �F����   h  �CVP������M��k�0�u����h�u��*�F��t(�>����E����hD;�FG;�v�}FF�> uыu��E����}��u�r�ǉ{�C   �g���j�C�C���hZf�1Af�0A@@Ju������������L@;�v�FF�~� �4����C��   �@Iu��C�����C�S��s3��ȋ�����{����95�z�X�������M�_^3�[�J�����jh�K�c  �M���������}�������_h�u�u����E;C�W  h   ��  Y�؅��F  ��   �wh���# S�u����YY�E�����   �u��vh�� ��u�Fh=�dtP����Y�^hS�=� ���Fp��   ��i��   j�  Y�e� �C� {�C�{�C�{3��E��}f�LCf�E�z@��3��E�=  }�L���f@��3��E�=   }��  ���g@���5�h�� ��u��h=�dtP�ƺ��Y��hS���E������   �0j�'  Y��%���u ���dtS萺��Y�Z����    ��e� �E��  Ã=l� uj��V���Y�l�   3�Ë�U��SV�u���   3�W;�to=�oth���   ;�t^9uZ���   ;�t9uP�������   �H  YY���   ;�t9uP��������   �FH  YY���   �޹�����   �ӹ��YY���   ;�tD9u@���   -�   P貹�����   ��   +�P蟹�����   +�P葹�����   膹�������   �=�nt9��   uP�,F  �7�_���YY�~P�E   ���it�;�t9uP�:���Y9_�t�G;�t9uP�#���Y���Mu�V����Y_^[]Ë�U��SV�5� W�}W�֋��   ��tP�֋��   ��tP�֋��   ��tP�֋��   ��tP�֍_P�E   �{��it	���tP�փ{� t
�C��tP�փ��Mu֋��   �   P��_^[]Ë�U��W�}����   SV�5� W�֋��   ��tP�֋��   ��tP�֋��   ��tP�֋��   ��tP�֍_P�E   �{��it	���tP�փ{� t
�C��tP�փ��Mu֋��   �   P��^[��_]Å�t7��t3V�0;�t(W�8�����Y��tV�E����> Yu���itV�Y���Y��^�3��jhL��  �������i�Fpt"�~l t�����pl��uj �r  Y���  �j�  Y�e� �Fl�=�j�i����E��E������   ��j�  Y�u�Ë�U����  ��f9Eu�e� �e�   f9Es�E��nf�Af#E���E��@�u�M��α���E��p�p�E�Pj�EP�E�jP�F  ����u!E��}� t�E�`p��E��M#�������V�D$�u(�L$�D$3���؋D$������d$�ȋ��d$��G�ȋ\$�T$�D$���������u�����d$�ȋD$���r;T$wr;D$v	N+D$T$3�+D$T$���؃� �ʋӋًȋ�^� ��U��VW3��u�6�����Y��u'90{vV�x ���  ;0{v��������uʋ�_^]Ë�U��VW3�j �u�u�E  ������u'90{vV�x ���  ;0{v��������uË�_^]Ë�U��VW3��u�u�F  ��YY��u,9Et'90{vV�x ���  ;0{v��������u���_^]Ë�U��W��  W�x �u�����  ��`�  w��t�_]Ë�U���O����u�����5�j����h�   �Ѓ�]Ë�U��h�����th�P�\ ��t�u��]Ë�U���u�����Y�u�,�j��  Y�j�  YË�U��V������t�Ѓ�;ur�^]Ë�U��V�u3����u���t�у�;ur�^]Ë�U��=h thh�H  Y��t
�u�hY�n���h�h�����YY��uBh9l�������$��c����=p� Ythp��G  Y��tj jj �p�3�]�jh0L�  j�  Y�e� 3�C9d{��   �`{�E�\{�} ��   �5h��B���Y���}؅�tx�5d��-���Y���u܉}�u����u�;�rW�	���9t�;�rJ�6���������������5h���������5d��������9}�u9E�t�}�}؉E����u܋}��h����_���Yh����O���Y�E������   �} u(�d{j�1  Y�u�����3�C�} tj�  Y��6
  Ë�U��j j�u�������]�jj j ������Ë�V�*�����V�����V��F  V赢��V�����V��F  V��1  V����V�F���h�d�|�����$��j^�jThPL�q	  3��}��E�P� �E�����j@j ^V�&���YY;��  �`��5@���   �0�@ ���@
�x�@$ �@%
�@&
�x8�@4 ��@�`���   ;�r�f9}��
  �E�;���   �8�X�;�E�   ;�|���E�   �[j@j ����YY��tV�M���`���@� ��   �*�@ ���@
�` �`$��@%
�@&
�`8 �@4 ��@��;�r��E�9=@�|���=@��e� ��~m�E����tV���tQ��tK�uQ�$��t<�u���������4�`��E� ���Fh�  �FP�\E  YY����   �F�E�C�E�9}�|�3ۋ���5`�����t���t�N��r�F���uj�X�
��H������P�h�����tC��t?W�$��t4�>%�   ��u�N@�	��u�Nh�  �FP��D  YY��t7�F�
�N@�����C���g����5@��(3��3�@Ëe��E���������o  Ë�VW�`��>��t1��   �� t
�GP����@   ;�r��6药���& Y����`�|�_^Ã=l� u�����V�5ttW3���u����   <=tGV�X���Y�t���u�jGW�n�����YY�=D{��tˋ5ttS�BV�'�����C�>=Yt1jS�@���YY���tNVSP�{�������t3�PPPPP�\��������> u��5tt�Ϯ���%tt �' �`�   3�Y[_^��5D{詮���%D{ ������U��Q�MS3�V���U�   9Et	�]�E��E��>"u3�9E��"��F�E��<���t��B�U���PF�C  Y��t��} t
�M��E�F�U�M��t2�}� u��� t��	u���t�B� �e� �> ��   �< t<	uF��N��> ��   �} t	�E�E��3�C3��FA�>\t��>"u&��u�}� t�F�8"u���3�3�9E����E����tI��t�\B���u�U���tU�}� u< tK<	tG��t=��P��t#��B  Y��t��M�E�F��M��E���B  Y��tF���UF�V�����t� B�U��M�����E^[��t�  ��Ë�U���S3�VW9l�u�t���h  �h{VS�l|�d�|��5T{;�t�E�8u�u��U��E�PSS�}��
����E���=���?sJ�M���sB�����;�r6P�q�����Y;�t)�U��E�P�WV�}�������E���H�8{�5<{3�����_^[�Ë�U��p|��SV�5W3�3�;�u.�֋�;�t�p|   �#����xu
jX�p|��p|����   ;�u�֋�;�u3���   ��f9t@@f9u�@@f9u�5� SSS+�S��@PWSS�E��։E�;�t/P����Y�E�;�t!SS�u�P�u�WSS�օ�u�u�脫��Y�]��]�W����\��t;�u����;��r���8t
@8u�@8u�+�@P�E��0�����Y;�uV��E����u�VW������V���_^[�Ë�V�82�82W��;�s���t�Ѓ�;�r�_^Ë�V�@2�@2W��;�s���t�Ѓ�;�r�_^Ë�U��3�9Ej ��h   P��t|��u]�3�@�<�]Ã=<�uWS3�9$�W�=�~3V�5(���h �  j �v�� �6j �5t|�׃�C;$�|�^�5(�j �5t|��_[�5t|��%t| Ë�U��QQV���������F  �V\�(kW�}��S99t��k����;�r�k��;�s99u���3���t
�X�]���u3���   ��u�` 3�@��   ����   �N`�M��M�N`�H����   �k�= k���;�}$k��~\�d9 �=k� kB߃�;�|�]�� �~d=�  �u	�Fd�   �^=�  �u	�Fd�   �N=�  �u	�Fd�   �>=�  �u	�Fd�   �.=�  �u	�Fd�   �=�  �u	�Fd�   �=�  �u�Fd�   �vdj��Y�~d��` Q�ӋE�Y�F`���[_^�Ë�U��csm�9Eu�uP����YY]�3�]��h�nd�5    �D$�l$�l$+�SVW�b1E�3�P�e��u��E��E������E��E�d�    ËM�d�    Y__^[��]Q���̋�U���S�]V�s35bW��E� �E�   �{���t�N�38�D����N�F�38�4����E�@f�  �M�U�S��[�E�M���t_�I �[�L��D��E�� �E���t����  �E���|@G�E��؃��u΀}� t$����t�N�38������N�V�3:豝���E�_^[��]��E�    �ɋM�9csm�u)�=� t h��#;  ����t�UjR�����M�  �E9XthbW�Ӌ��  �E�M��H����t�N�38�.����N�V�3:�����E��H���5  �����9S�R���hbW���M  ������U����b�e� �e� SW�N�@��  ��;�t��t	�Уb�`V�E�P�� �u�3u��� 3���3��� 3��E�P�� �E�3E�3�;�u�O�@����u������5b�։5b^_[�Ë�VW3��x|�<�4ku��0k�8h�  �0���:  YY��tF��$|�3�@_^Ã$�0k 3����S�V�0kW�>��t�~tW��W貥���& Y����Pl|ܾ0k_���t	�~uP�Ӄ���Pl|�^[Ë�U��E�4�0k�� ]�jhpL����3�G�}�3�9t|u����j�����h�   ����YY�u�4�0k9t���nj����Y��;�u�����    3��Qj
�Y   Y�]�9u,h�  W�9  YY��uW����Y誥���    �]���>�W�Ť��Y�E������	   �E��U����j
�(���YË�U��EV�4�0k�> uP�"���Y��uj����Y�6�� ^]Ë�U��$��(�k����U+P��   r	��;�r�3�]Ë�U����M�AV�uW��+y�������i�  ��D  �M��I�M�����  S�1��U�V��U��U�]��ut��J��?vj?Z�K;KuB�   ��� s����L��!\�D�	u#�M!��J���L��!���   �	u�M!Y�]�S�[�M�M�Z�U�Z�R�S�M�����J��?vj?Z�]����]���   +u��]���j?�uK^;�v��M�����J�M�;�v��;�t^�M�q;qu;�   ��� s������!t�D�Lu!�M!1��K�����!���   �Lu�M!q�M�q�I�N�M�q�I�N�u��]�}� u;���   �M��ыY�N�^�q�N�q�N;Nu`�L�M���L�� s%�} u�ʻ   ���M	�   �����D�D	�)�} u�J�   ���M	Y�J�   ��ꍄ��   	�E���D0��E����   ��}����   �8��5 h @  ��H� �  SQ�֋8���}�   ���	P��}�@�8�����    ��}�@�HC��}�H�yC u	�`���}�x�ueSj �p�֡�}�pj �5t|���$���}k��(�+ȍL�Q�HQP�~����E���$�;�}v�m�(��0��E��}�=8�[_^�á4�V�5$�W3�;�u4��k�P�5(�W�5t|�� ;�u3��x�4��5$��(�k�5(�h�A  j�5t|���F;�t�jh    h   W�� �F;�u�vW�5t|��뛃N��>�~�$��F����_^Ë�U��QQ�M�ASV�qW3���C��}���i�  ��0D  j?�E�Z�@�@��Ju�j��h   ��yh �  W�� ��u����   �� p  �U�;�wC��+����GA�H�����  ����  ��������@��  �Pǀ�  �     IuˋU��E��  �O�H�A�J�H�A�d�D 3�G����   �FC�������E�NCu	x�   �������!P��_^[�Ë�U����M�ASV�uW�}��+Q������i�  ��D  �M�O����I;�|9���M�]��U  ���E  �;��;  �M���I�M���?vj?Y�M��_;_uC�   ��� s��M��L��!\�D�	u&�M!������M��L��!���   �	u�M!Y�O�_�Y�O��y�M+�M��}� ��   �}��M��O�L1���?vj?_�]���]�[�Y�]�Y�K�Y�K�Y;YuW�L�M���L�� s�} u�ϻ   ���M	�D�D��� �} u�O�   ���M	Y����   �O�   ���	�U�M��D2���L���U�F�B��D2��<  3��8  �/  �])u�N�K��\3��u��N�]�K���?vj?^�E���   �u���N��?vj?^�O;OuB�   ��� s����t��!\�D�u#�M!��N���L��!���   �	u�M!Y�]�O�w�q�w�O�q�uu��u��N��?vj?^�M��y�K�{�Y�K�Y�K;KuW�L�M���L�� s�} u�ο   ���M	9�D�D��� �} u�N�   ���M	y����   �N�   ���	�E��D�3�@_^[�Ë�U����$��Mk�(�������M���SI�� VW}�����M���������3���U��0�����S�;#U�#��u
���];�r�;�u�(���S�;#U�#��u
���];�r�;�u[��{ u
���];�r�;�u1�(��	�{ u
���];�r�;�u�����؉]��u3��	  S�:���Y�K��C�8�t�0��C��U����t����   �|�D#M�#��u)�e� ���   �HD�9#U�#��u�E����   ����U���i�  ��D  �M�L�D3�#�u����   #M�j _��G��}��M�T��
+M�����N��?�M�~j?^;��  �J;Ju\�� �   �}&����M��|8�Ӊ]�#\�D�\�D�u3�M�]!�,�O���M�����   �|8��!��]�u�]�M�!K��]�}� �J�z�y�J�z�y��   �M��y�J�z�Q�J�Q�J;Ju^�L�M���� �L}#�} u�   �����	;�ο   ���M�	|�D�)�} u�N�   ���	{�M�����   �N�   ���	7�M���t�
�L���M��u�эN�
�L2��u��y�>��u;�}u�M�;8�u�%�} �M���B_^[�����SVW�T$�D$�L$URPQQh~d�5    �b3ĉD$d�%    �D$0�X�L$,3�p���t;�T$4���t;�v.�4v�\���H�{ u�h  �C�  �   �C�  �d�    ��_^[ËL$�A   �   t3�D$�H3��5���U�h�p�p�p�>�����]�D$�T$��   �U�L$�)�q�q�q(������]� UVWS��3�3�3�3�3���[_^]Ë���j�c  3�3�3�3�3���U��SVWj j h�~Q�a  _^[]�U�l$RQ�t$������]� ��U��QQ�EV�u�E��EWV�E��Y.  ���Y;�u������ 	   �ǋ��J�u�M�Q�u�P�� �E�;�u����t	P����Y�ϋ�����`������D0� ��E��U�_^��jh�L�(�������u܉u��E���u蕘���  �z���� 	   �Ƌ���   3�;�|;@�r!�k����8�Q���� 	   WWWWW�������ȋ�����`���������L1��u&�*����8����� 	   WWWWW�͈����������[P�-  Y�}���D0t�u�u�u�u�������E܉U������ 	   �ʗ���8�M���M���E������   �E܋U��k�����u��-  YË�U���  �����b3ŉE��EV3���4�����8�����0���9uu3���  ;�u'�X����0�>���VVVVV�    �����������  SW�}�����4�`������ǊX$�����(�����'�����t��u0�M����u&����3��0�Ӗ��VVVVV�    萇�����C  �@ tjj j �u�~������u�i  Y����  ��D���  �Ю���@l3�9H�������P��4�� ����� ���`  3�9� ���t���P  �� ��4��������3���<���9E�B  ��D�����'������g  ���(���3���
���� ����ǃx8 t�P4�U�M��`8 j�E�P�K��P��  Y��t:��4���+�M3�@;���  j��@���SP�q  �������  C��D����jS��@���P�M  �������  3�PPj�M�Qj��@���QP�����C��D����� �����\  j ��<���PV�E�P��(���� �4�l���)  ��D�����0����9�<�����8����  �� ��� ��   j ��<���Pj�E�P��(���� �E��4�l����  ��<�����  ��0�����8����   <t<u!�33�f��
��CC��D�����@����� ���<t<uR��@�����*  Yf;�@����h  ��8����� ��� t)jXP��@�����*  Yf;�@����;  ��8�����0����E9�D���������'  ����8����T4��D8�  3ɋ��@���  ��4�����@�������   ��<���9M�   ���(�����<�����D��� +�4�����H���;Ms9��<�����<����A��
u��0���� @��D����@��D�����D����  r؍�H���+�j ��,���PS��H���P��4�l���B  ��,����8���;��:  ��<���+�4���;E�L����   ��D�������   9M�M  ���(�����D�����<��� +�4�����H���;MsF��D�����D����AAf��
u��0���j[f�@@��<�����<���f�@@��<����  r��؍�H���+�j ��,���PS��H���P��4�l���b  ��,����8���;��Z  ��D���+�4���;E�?����@  9M�|  ��D�����<��� +�4���j��H���^;Ms<��D�����D����f��
uj[f���<����<���f�Ɓ�<����  r�3�VVhU  ������Q��H���+��+���P��PVh��  �� ��;���   j ��,���P��+�P��5����P��(���� �4�l��t�,���;�������@���;�\��D���+�4�����8���;E�
����?j ��,���Q�u��4����0�l��t��,�����@��� ��8��������@�����8��� ul��@��� t-j^9�@���u�Ɛ��� 	   �ΐ���0�?��@����Ґ��Y�1��(�����D@t��4����8u3��$膐���    莐���  ������8���+�0���_[�M�3�^�Å����jh�L������E���u�R����  �7���� 	   ����   3�;�|;@�r!�)����8����� 	   WWWWW�̀�����ɋ�����`���������L1��t�P�%  Y�}���D0t�u�u�u�.������E��謏��� 	   贏���8�M���E������	   �E��\�����u��%  YË�U���~h   ����Y�M�A��t�I�A   ��I�A�A�A   �A�a �]Ë�U��E���u�!���� 	   3�]�V3�;�|;@�r����VVVVV� 	   ������3���ȃ�����`����D��@^]øPlá �Vj^��u�   �;�}�ƣ �jP����YY���ujV�5 ������YY���ujX^�3ҹPl����� �����n|�j�^3ҹ`lW������`�����������t;�t��u�1�� B���l|�_3�^��'  �=\{ t�V%  �5�*���YË�U��V�u�Pl;�r"���nw��+�����Q�X����N �  Y�
�� V�� ^]Ë�U��E��}��P�+����E�H �  Y]ËE�� P�� ]Ë�U��E�Pl;�r=�nw�`���+�����P����Y]Ã� P�� ]Ë�U��M���E}�`�����Q�����Y]Ã� P�� ]Ë�U��EV3�;�u����VVVVV�    ��}���������@^]Ë�U����b3ŉE�SV�u�F@W�6  V����Y��j���t.V����Y���t"V������V�<�`��y�����Y��Y��Ê@$$<��   V�X���Y���t.V�L���Y���t"V�@�����V�<�`��0�����Y��Y��Ê@$$<��   V����Y���t.V����Y���t"V�������V�<�`��������Y��Y����@�t]�u�E�jP�E�P�>(  ����t���  �]3�9}�~0�Nx��L=���A���D=�VP�ב��YY���t�G;}�|�f�E� �F�x��Ef����EVP��$  YY�M�_^3�[�̀���áb��3�9~����Ë�U���SV�u3�;�t9]t8u�E;�t3�f�3�^[���u�M��'����E�9Xu�E;�tf�f�8]�t�E��`p�3�@�ʍE�P�P��   YY��t}�E����   ��~%9M| 3�9]��R�uQVj	�p�� ���E�u�M;��   r 8^t���   8]��e����M��ap��Y����u���� *   8]�t�E��`p�����:���3�9]��P�u�E�jVj	�p�� ���:���뺋�U��j �u�u�u�������]Ë�U����u�M������E�M����   �A% �  �}� t�M��ap��Ë�U��j �u����YY]�jh�L�S���3��]3�;���;�u讉���    WWWWW�kz��������S�=<�u8j����Y�}�S�9���Y�E�;�t�s���	�u���u��E������%   9}�uSW�5t|�H ���������3��]�u�j�����YË�U��3�@�} u3�]���U��SVWUj j h��u��P  ]_^[��]ËL$�A   �   t2�D$�H�3��A~��U�h�P(R�P$R�   ��]�D$�T$��   �SVW�D$UPj�h��d�5    �b3�P�D$d�    �D$(�X�p���t:�|$,�t;t$,v-�4v���L$�H�|� uh  �D��I   �D��_   뷋L$d�    ��_^[�3�d�    �y��u�Q�R9Qu�   �SQ��n�SQ��n�L$�K�C�kUQPXY]Y[� ����������������U��W�}3�������ك��E���8t3�����_�Ë�U����u�M�詁���E����   ~�E�Pj�u��#  ������   �M�H���}� t�M��ap��Ë�U��={ u�E��j�A��]�j �u����YY]Ë�U���SV�u�M��(����]�   ;�sT�M胹�   ~�E�PjS�o#  �M������   �X����t���   ��   �}� t�E��`p����   �E胸�   ~1�]�}�E�P�E%�   P�t���YY��t�Ej�E��]��E� Y��q���� *   3Ɉ]��E� A�E�j�p�U�jRQ�M�QV�p�E�P��  ��$���o������E�t	�M�����}� t�M��ap�^[�Ë�U��={ u�E�H���w�� ]�j �u�����YY]Ë�U���(�b3ŉE�SV�uW�u�}�M������E�P3�SSSSW�E�P�E�P�i-  �E�E�VP��"  ��(�E�u+��u8]�t�E�`p�jX�/��u8]�t�E�`p�j���E�u��E�u�8]�t�E�`p�3��M�_^3�[�z���Ë�U���(�b3ŉE�SV�uW�u�}�M��.���E�P3�SSSSW�E�P�E�P��,  �E�E�VP�p'  ��(�E�u+��u8]�t�E�`p�jX�/��u8]�t�E�`p�j���E�u��E�u�8]�t�E�`p�3��M�_^3�[�z���Ë�U��MSV�u3�W�y;�u�{���j^�0SSSSS�9u�������   9]v݋U;ӈ~���3�@9Ew�C���j"Y�����;��0�F~�:�t��G�j0Y�@J;��M;ӈ|�?5|�� 0H�89t�� �>1u�A��~W�'���@PWV�.�����3�_^[]Ë�U��Q�U�BS��VW��% �  ��  #ωE�B��پ   �%�� �u���t;�t�� <  �(��  �$3�;�u;�u�Ef�M�X��L��<  �]����������M��E���H���u��P������Ɂ���  �P���t�M�_^f�H[�Ë�U���0�b3ŉE��ES�]V�E�W�EP�E�P����YY�E�Pj j���u�����f��1  �uЉC�E։�EԉC�E�P�uV�f�����$��t3�PPPPP�Gr�����M�_�s^��3�[��w�����������WVU3�3�D$�}GE�T$���ڃ� �D$�T$�D$�}G�T$���ڃ� �D$�T$�u(�L$�D$3���؋D$������d$�ȋ��d$��G�؋L$�T$�D$���������u�����d$�ȋD$���r;T$wr;D$v	N+D$T$3�+D$T$My���؃� �ʋӋًȋ�Ou���؃� ]^_� ̀�@s�� s����Ë�3Ҁ����3�3��j����YË�U��E�M%����#�V������t1W�}3�;�tVV�Z:  YY��G���j_VVVVV�8�r������_��uP�u��t	�*:  ���!:  YY3�^]Ë�U��E�~�~� ~�$~]Ë�U��E�(kV9Pt��k�u��;�r�k�M^;�s9Pt3�]��5 ~谖��Y�j h�L�2���3��}�}؋]��Lt��jY+�t"+�t+�td+�uD�L������}؅�u����a  �~�~�`�w\���]���������Z�Ã�t<��t+Ht�2����    3�PPPPP��p����뮾 ~� ~��~�~�
�$~�$~�E�   P�����E�Y3��}���   9E�uj�p���9E�tP�O���Y3��E���t
��t��u�O`�MԉG`��u@�Od�M��Gd�   ��u.�k�M܋ k�k�9M�}�M�k��W\�D�E����T�����E������   ��u�wdS�U�Y��]�}؃}� tj �����Y�S�U�Y��t
��t��u�EԉG`��u�EЉGd3������Ë�U���SVW�����e� �=,~ ����   h(!�� �����*  �5\ h!W�օ��  P�/����$!W�,~��P�����$� W�0~��P�����$� W�4~��P����Y�<~��th� W��P�ؓ��Y�8~�8~;�tO9<~tGP�6����5<~���)���YY����t,��t(�օ�t�M�Qj�M�QjP�ׅ�t�E�u	�M    �9�0~;�t0P����Y��t%�ЉE���t�4~;�tP�ɓ��Y��t�u��ЉE��5,~豓��Y��t�u�u�u�u����3�_^[�Ë�U��ES3�VW;�t�};�w�x}��j^�0SSSSS�6n�������<�u;�u��ڋ�8tBOu�;�t��
BF:�tOu�;�u��1}��j"Y����3�_^[]Ë�U��SV�u3�W9]u;�u9]u3�_^[]�;�t�};�w��|��j^�0SSSSS�m��������9]u��ʋU;�u��у}���u�
�@B:�tOu���
�@B:�tOt�Mu�9]u�;�u��}�u�EjP�\�X�x�����u|��j"Y���낋�U��MV3�;�|��~��u�|t�(�|t�|t��:|��VVVVV�    ��l�������^]Ë�U��E��t���8��  uP�4{��Y]Ë�U��f�Ef��0s�����]�f��:s����0]ù�  ��f;���  �`  ��f;���  ��
f;�s��+�]ù�  ��f;��s  ��
f;�r�f	  ��f;��[  ��
f;�rɹ�	  ��f;��C  ��
f;�r��f
  ��f;��+  ��
f;�r���
  ��f;��  ��
f;�r��f  ��f;���   ��
f;��e����f  ��f;���   ��
f;��I�����  ��f;���   ��
f;��-����f  ��f;���   ��
f;������P  ��f;���   ��
f;��������  ��f;�rs��
f;��������P��f;�r]�*  f;�������@  ��f;�rC��
f;��������  ��f;�r+��
f;��������0��f;�r�  ���  f;��v������]��̋D$�L$ȋL$u	�D$��� S��؋D$�d$؋D$���[� ��U����b3ŉE�SV3�W��9@~u8SS3�GWh4!h   S�0��t�=@~�����xu
�@~   9]~"�M�EI8t@;�u�����E+�H;E}@�E�@~����  ;���  ����  �]�9] u��@�E �5� 3�9]$SS�u���u��   P�u �֋�;���  ~Cj�3�X����r7�D?=   w�5  ��;�t� ��  �P�J}��Y;�t	� ��  ���E���]�9]��>  W�u��u�uj�u �օ���   �50SSW�u��u�u�֋ȉM�;���   �E   t)9]��   ;M��   �u�uW�u��u�u���   ;�~Ej�3�X���r9�D	=   w�S4  ��;�tj���  ���P�|��Y;�t	� ��  �����3�;�tA�u�VW�u��u�u�0��t"SS9]uSS��u�u�u�VS�u �� �E�V����Y�u������E�Y�Y  �]�]�9]u��@�E9] u��@�E �u��3  Y�E���u3��!  ;E ��   SS�MQ�uP�u ��3  ���E�;�tԋ5@ SS�uP�u�u�։E�;�u3��   ~=���w8��=   w�=3  ��;�t����  ���P�r{��Y;�t	� ��  �����3�;�t��u�SW�f�����u�W�u�u��u�u�։E�;�u3��%�u�E��uPW�u �u��C3  ���u������#u�W�|���Y��u�u�u�u�u�u�@ ��9]�t	�u��u��Y�E�;�t9EtP�u��Y�ƍe�_^[�M�3��k���Ë�U����u�M��Mp���u(�M��u$�u �u�u�u�u�u�(����� �}� t�M��ap��Ë�U��QQ�b3ŉE��D~SV3�W��;�u:�E�P3�FVh4!V�8 ��t�5D~�4����xu
jX�D~��D~����   ;���   ����   �]�9]u��@�E�5� 3�9] SS�u���u��   P�u�֋�;���   ~<�����w4�D?=   w�V1  ��;�t� ��  �P�y��Y;�t	� ��  ���؅�ti�?Pj S�"d����WS�u�uj�u�օ�t�uPS�u�8 �E�S�����E�Y�u3�9]u��@�E9]u��@�E�u��0  Y���u3��G;EtSS�MQ�uP�u�1  ����;�t܉u�u�u�u�u�u�< ��;�tV�s��Y�Ǎe�_^[�M�3��i���Ë�U����u�M��Nn���u$�M��u �u�u�u�u�u�������}� t�M��ap��Ë�U��V�u����  �v�!s���v�s���v�s���v�	s���v�s���v��r���6��r���v ��r���v$��r���v(��r���v,��r���v0��r���v4��r���v�r���v8�r���v<�r����@�v@�r���vD�r���vH�r���vL�r���vP�r���vT�wr���vX�or���v\�gr���v`�_r���vd�Wr���vh�Or���vl�Gr���vp�?r���vt�7r���vx�/r���v|�'r����@���   �r�����   �r�����   �r�����   ��q�����   ��q�����   ��q�����   ��q�����   ��q�����   ��q�����   �q�����   �q����,^]Ë�U��V�u��t5�;�otP�q��Y�F;�otP�vq��Y�v;5�otV�dq��Y^]Ë�U��V�u��t~�F;�otP�Bq��Y�F;�otP�0q��Y�F;�otP�q��Y�F;�otP�q��Y�F;�otP��p��Y�F ;�otP��p��Y�v$;5�otV��p��Y^]���������������U��V3�PPPPPPPP�U�I �
�t	���$��u����I ���
�t	���$s���� ^������������U��V3�PPPPPPPP�U�I �
�t	���$��u���
�t���$s�F��� ^�Ë�U����u�M��k���}�}3���u�u�u�u�8 �}� t�M��ap���jhM�J����M3�;�v.j�X3���;E�@u�p���    WWWWW�Za����3���   �M��u;�u3�F3ۉ]���wi�=<�uK������u�E;,�w7j�����Y�}��u�����Y�E��E������_   �]�;�t�uWS�4_����;�uaVj�5t|����;�uL9=�}t3V�Ό��Y���r����E;��P����    �E���3��uj�s���Y�;�u�E;�t�    ���~����jh0M�,����]��u�u��s��Y��  �u��uS�n��Y�  �=<���  3��}�����  j�����Y�}�S����Y�E�;���   ;5,�wIVSP���������t�]��5V����Y�E�;�t'�C�H;�r��PS�u���d��S�����E�SP�������9}�uH;�u3�F�u������uVW�5t|���E�;�t �C�H;�r��PS�u��d��S�u��������E������.   �}� u1��uF������uVSj �5t|�� ����u�]j����YË}����   9=�}t,V�"���Y��������4n��9}�ul����P��m��Y��_����   �n��9}�th�    �q��uFVSj �5t|�� ����uV9�}t4V蹊��Y��t���v�V詊��Y��m���    3�������m���|�����u�m������P�Rm���Y������������̋�U��M�MZ  f9t3�]ËA<��8PE  u�3ҹ  f9H��]�����������̋�U��E�H<��ASV�q3�W�D��v�}�H;�r	�X�;�r
B��(;�r�3�_^[]������������̋�U��j�hPMh�nd�    P��SVW�b1E�3�P�E�d�    �e��E�    h   �*�������tU�E-   Ph   �P�������t;�@$���Ѓ��E������M�d�    Y_^[��]ËE��3�=  ���Ëe��E�����3��M�d�    Y_^[��]Ë�U��E�L~]Ë�U��E�P~]�jhpM�����e� �u�u�@�E��/�E� � �E�3�=  �����Ëe�}�  �uj�t�e� �E������E�����Ë�U����u�M��e���E�M�U�Tu�} t�M����   �A#E�3���t3�@�}� t�M��ap��Ë�U��jj �uj ������]Ë�U��j
j �u�+  ��]Ë�U��MS3�;�VW|[;@�sS������<�`��������@t5�8�t0�=�tu+�tItIuSj��Sj��Sj��D���3����j��� 	   ��j������_^[]Ë�U��E���u�j���  �j��� 	   ���]�V3�;�|";@�s�ȃ�����`�����@u$�rj���0�Xj��VVVVV� 	   �[��������� ^]�jh�M�����}����������4�`��E�   3�9^u6j
����Y�]�9^uh�  �FP�����YY��u�]��F�E������0   9]�t����������`��D8P�� �E������3ۋ}j
�M���YË�U��E�ȃ�����`����DP�� ]Ë�U����b3ŉE�V3�95 ptO�=�p�u��)  ��p���u���  �pV�M�Qj�MQP�P��ug�= pu�����xuω5 pVVj�E�Pj�EPV�LP�� ��p���t�V�U�RP�E�PQ�H��t�f�E�M�3�^�&^����� p   ��jh�M�3���3ۉ]�j�!���Y�]�j_�}�;= �}W������9tD� �@�tP��)  Y���t�E��|(���� P���4�jg��Y��G��E������	   �E������j�����YË�U��SV�u�F�Ȁ�3ۀ�u@�  t9�FW�>+���~,WPV�����YP�}�����;�u�F��y����F��N ���_�F�f �^��[]Ë�U��V�u��u	V�5   Y�/V�|���Y��t�����F @  tV�Y���P�K)  Y��Y��3�^]�jh�M����3��}�}�j�����Y�}�3��u�;5 ���   ���98t^� �@�tVPV�^���YY3�B�U�����H���t/9UuP�J���Y���t�E��9}u��tP�/���Y���u	E܉}��   F�3��u��4�V�g���YY��E������   �}�E�t�E��e����j�8���Y�j����YË�U��QV�uV�S����E�FY��u�]f��� 	   �N ���  �=  �@t�@f��� "   ��t�f ���   �N�����F�F�f �e� Sj���[ÉF�  u,�+����� ;�t������@;�u�u����Y��uV�X���Y�F  W��   �F�>�H��N+�+ˉN��~WP�u�K������E��N�� �F�=����M���t���t�����������`����j�@ tSj j Q����#����t-�F�]f��j�E�P�u���]f�]���������E�9}�t�N ���  ���%��  _[^�Ë�U���SV�u3�W�};�u;�v�E;�t�3��   �E;�t�������v��d��j^SSSSS�0�U�������V�u�M��^���E�9X��   f�E��   f;�v6;�t;�vWSV�S�����td��� *   �id��� 8]�t�M��ap�_^[��;�t2;�w,�Id��j"^SSSSS�0�U����8]��y����E��`p��m�����E;�t�    8]��%����E��`p������MQSWVj�MQS�]�p�� ;�t9]�^����M;�t�������z�D���;��g���;��_���WSV��R�����O�����U��j �u�u�u�u�|�����]Ë�U���S�u�M��]���]�C=   w�E苀�   �X�u�]�}�E�P�E%�   P����YY��t�Ej�E��]��E� Y�
3Ɉ]��E� A�E�j�p�p�E�PQ�E�P�E�jP������ ��u8E�t�E��`p�3���E�#E�}� t�M��ap�[�Ë�U���,�E�H
S�ف� �  �M�H�M��H� ���  ���?  ��W�M�E�����u'3�3�9\��u@��|�3��  3��}૫j�X�  �e V�u��}ԥ���5pN�N���������с�  ��]��E�yJ���B�|��j3�Y+�@���M����   �E������҅T����|�� u@��|��n�ƙjY#������  �yN���F�e� +�3�B��L���1�u�19ur"9U���t+�e� �L����r�u;�r��s�E�   H�U��M�yщM�M������!�E�@��}jY�|��+�3��} tC�p��+p;�}3��}૫��  ;��  +E��uԋȍ}ख़��¥������  ��yJ���B�e� �e ��������E�    )U��׋]�\���3��#ωM�����M�u�3�u����E�}�u�|Ӌ�j���M�Z+�;�|�1�t����d�� J����}�5pN�N���������с�  ��E�yJ���BjY+�3�B��\���M����   ������҅T����|�� u@��|��f�ƙjY#������  �yN���F�e 3�+�B��L���1�<;�r;�s�E   �9�M���t�L����r3�;�r��s3�G�1��HyދM������!�E�@��}jY�|��+�3��pA����������  �yJ���B�e� �e ��������E�    )U��׋]�\���3��#ωM�����M�u�3�u����E�}�u�|Ӌ�j���M�Z+�;�|�1�t����d�� J����}�j3�X�Z  ;p�p��   3��}૫��M�   �����������  �yJ���B�e� �e ��������E�    )U��׋]�\���3��#ωM�����M�u�3�u����E�}�u�|Ӌ�j���M�Z+�;�|�1�t����d�� J����}�p�p�3�@�   �p�e����؋���������  �yJ���B�e� �e ��������E�    )U��֋M�|����#ΉM�����M}�|���}��M����E�}�}�|Ћ�j���M�Z+�;�|�1�t����d�� J����}�3�^jY+p��M���Ɂ�   �ًp]���@u�M�U�Y��
�� u�M�_[�Ë�U���,�E�H
S�ف� �  �M�H�M��H� ���  ���?  ��W�M�E�����u'3�3�9\��u@��|�3��  3��}૫j�X�  �e V�u��}ԥ���5$pN�N���������с�  ��]��E�yJ���B�|��j3�Y+�@���M����   �E������҅T����|�� u@��|��n�ƙjY#������  �yN���F�e� +�3�B��L���1�u�19ur"9U���t+�e� �L����r�u;�r��s�E�   H�U��M�yщM�M������!�E�@��}jY�|��+�3��} tC� p��+$p;�}3��}૫��  ;��  +E��uԋȍ}ख़��¥������  ��yJ���B�e� �e ��������E�    )U��׋]�\���3��#ωM�����M�u�3�u����E�}�u�|Ӌ�j���M�Z+�;�|�1�t����d�� J����}�5$pN�N���������с�  ��E�yJ���BjY+�3�B��\���M����   ������҅T����|�� u@��|��f�ƙjY#������  �yN���F�e 3�+�B��L���1�<;�r;�s�E   �9�M���t�L����r3�;�r��s3�G�1��HyދM������!�E�@��}jY�|��+�3��(pA����������  �yJ���B�e� �e ��������E�    )U��׋]�\���3��#ωM�����M�u�3�u����E�}�u�|Ӌ�j���M�Z+�;�|�1�t����d�� J����}�j3�X�Z  ;p�(p��   3��}૫��M�   �����������  �yJ���B�e� �e ��������E�    )U��׋]�\���3��#ωM�����M�u�3�u����E�}�u�|Ӌ�j���M�Z+�;�|�1�t����d�� J����}�p�0p�3�@�   �0p�e����؋���������  �yJ���B�e� �e ��������E�    )U��֋M�|����#ΉM�����M}�|���}��M����E�}�}�|Ћ�j���M�Z+�;�|�1�t����d�� J����}�3�^jY+(p��M���Ɂ�   �ً,p]���@u�M�U�Y��
�� u�M�_[�Ë�U���|�b3ŉE��ES3�V3��E��EF3�W�E��}��]��u��]��]��]��]��]��]��]�9]$u��W��SSSSS�    �H����3��N  �U�U��< t<	t<
t<uB��0�B���/  �$�|��Ȁ�1��wjYJ�݋M$�	���   �	:ujY������+tHHt����  ���jY�E� �  뢃e� jY뙊Ȁ�1�u���v��M$�	���   �	:uj�<+t(<-t$:�t�<C�<  <E~<c�0  <e�(  j�Jj�y����Ȁ�1���R����M$�	���   �	:�T���:��f����U��  �u��<9�}�s
�E�*ÈG��E��B:�}�M$�	���   �	:�]���<+t�<-t��`����}� �u��u�u&��M��B:�t��<9Ճ}�s�E�*ÈG�M��B:�}��*Éu�<	�n���j�����J��M��Ȁ�1��wj	��������+t HHt���;���j�����M��jY�@���j�o����u���B:�t�,1<v�J�(�Ȁ�1��v�:�뽃}  tG����+�J��M�t�HHt��у}� �E����  jX9E�v�}�|�E�O�E��E��}� ��  �Yj
YJ��
�����뾉u�3��<9 k�
���L1Ё�P  	�B:�}���Q  �M��<9�[����B:�}��O����M��E�O�? t�E�P�u��E�P��  �E�3҃�9U�}��E�9U�uE9U�u+E=P  �"  =�����.  ��p��`�E�;���  }�عXr�E���`9Uu3�f�E�9U���  ��M�3ҋE��}���T���M�;���  k���ظ �  f9r��}�����M��]��K
3��E��EԉE؉E܋E΋��  3�#�#ʁ� �  ��  ��u���f;��!  f;��  ���  f;��
  ��?  f;�w3��EȉE��  3�f;�uB�E����u9u�u9u�u3�f�E���  f;�u!B�C���u9su93u�ủuȉu���  �u��}��E�   �E��M���M���~R�DĉE��C�E��E��M��	� �e� ���O��4;�r;�s�E�   �}� �w�tf��E��m��M��}� �GG�E��M��}� ����  f��~7�}܅�x+�u؋E��e����������?�����  �u؉E�f���f��M����  f��}B��������E�t�E��E܋}؋M��m�������E������N�}؉E�u�9u�tf�M�� �  ��f9M�w�Mԁ��� �� � u4�}��u+�e� �}��u�e� ���  f9M�uf�E�B�f�E���E���Eָ�  f;�r#3�3�f9E��E����E�I��   ��� ���M��;f�E�U�f�EċE؉EƋE܉E�f�U��3�f�����e� H%   � ���e� �Ẽ}� �<����E��MċuƋU����/�E�   �3���  �   �3��E�   ��E�   3�3�3�3��}�E�f�f�G
�E��w�W�M�_^3�[��F���ÐN�����+�p���������v�%���U���t�b3ŉE�S�]VW�u�}�f��U��ʸ �  #ȁ��  �]��E���E���E���E���E���E���E���E���E���E���E���E�?�E�   �M�f��t�C-��C �u�}�f��u/��u+��u'3�f;�����$ f��C�C�C0�S3�@�  ��  f;���   3�@f��   �;�u��t��   @uh�*�Qf��t��   �u��u;h|*�;�u0��u,ht*�CjP��S����3���tVVVVV��?�����C�*hl*�CjP�S����3���tVVVVV�?�����C3��q  �ʋ�i�M  �������Ck�M��������3���f�M��p�ۃ�`�E�f�U�u�}�M�����  }�Xr�ۃ�`�E�����  �E�T�˃������g  k�M����M�� �  f9r���}ĥ��Eĥ�MƉE��P
3ɉM��M��M�M��M��3�� �  �u���  #�#֍4
����  f;���  f;���  ���  f;���  ��?  f;�w3��u�u�u���  3�f;�uG�E����u9u�u9u�u3�f�E��  f;�uG�@���u	9pu90t�!u��u��E�   �M��U�ɉU���~U�L����M��E��E���E�� �V��ȃe� �
;�r;�s�E�   �}� �F�tf��E��m��M��}� ��E�FF�E��M��}� ����  f��~;�E�   �u-�E�M��e��������E�E�������  �E�f���f��M����  f��}B��������E�t�E��M��u�U��m������M������H�u�M�u�9E�tf�M�� �  ��f9M�w�M����� �� � u4�}��u+�e� �}��u�e� ���  f9M�uf�E�G�f�E���E���E��  f;���   3�3�f9E��E����E�I��   ��� ���M�3�;��{����M�����?  ��  f;���  �E�3҉U��U��U�U��U��ɋ�3�#�#Ё� �  ���4
�]���f;��L  f;��C  ���  f;��5  ��?  f;�wK3��E�E��9  f�E�}�f�E��E�E�E��E�f�}��V���3�3�f9u���H%   � ���E��\���3�f;�uF�E����u9E�u9E�u	f�E���  f;�uF�E����u9E�u	9E��v����E��}��E�   �E��M���M���~J�M؉M��D��M���	�e� �ʋW��
;�r;�s�E�   �}� �_�tf��m�@@�M��}� �GG�E��M��}� ����  f��~7�}���x+�E�M��e��������E����?���  �E�f���f��M����  f��}B��������E�t�E��M��}�U��m�������M������H�}�M�u�9E�tf�M�� �  ��f9M�w�M����� �� � u4�}��u+�e� �}��u�e� ���  f9M�uf�E�F�f�E���E���E��  f;�r#3�3�f9E��E����E�I��   ��� ���M��;f�E�u�f�E��E�E�E��E�f�u��3�f�����e� H%   � ���e� �E��E�U��E��}f�t2����+3�f�� �  f9E��B����$ �B�B0�B �^�����~j_�u������?  3�f�E��E�   �E��]�M��e����؋E������M��]�E�u؅�}2�ށ��   ~(�E�]�M��m�����؋E������N�]�E���؍G�Z�]��E�����   �U��E�u��}ĥ���e��}��e���� ʋU�����֋��4	����U���ȋE���<;�r;�s�F3�;�r��s3�B����tA�Eȍ0�U�;�r;�sAM����ʍ4?�u��u��M������0������C�M��}� �u��E� �K���K�K<5}�M��D�;9u	�0K;]�s�E�;]�sCf� �*؀��ˈX�D �E��M�_^3�[��=���À;0uK;�s��E�;�s�3�f�� �  f9U��@���ʀ��� �P�0�@ ����3���t@��t����t����t����t�� ��   t���˺   #�V�   t#��   t;�t;�u   �   �   �ˁ�   t��   u���^��   t   �3���t��   SVW�   ��t���t   ��t   ��t   �   ��   tǋʾ   #�t;�t;�t;�u `  � @  �    �   _#�^[��   t��   t
;�u �  Ã�@�@�  Ë�U���SVW��}��]�3���tjZ��t����t����t���� t����t��   �ˋ��   #ƿ   t$=   t=   t;�u����   ���   #�t��   u��   ���   ��   t��   �}�M����#�#���E;���   ���
������E��m���}��]�3���tjZ��t����t����t���� t����t��   �ˋ�#�t(=   t=   t;�u��   ���   ���   ��   t��   u��   ���   ��   t��   �U��3�95x���  ���}��]��E���yj^�   t���   t���   t���   t���   t��   �Ȼ `  #�t*��    t�� @  t;�u��   ���   ���   �@�  #ǃ�@t-�  t��@u��   ���   ���   �E��#E��#��;�u���   ����P�E��0	  Y�]�M�3҄�yjZ��   t����   t����   t����   t���   ��t��   ��#�t$=    t= @  t;�u��   �
��   ��#σ�@t���  t��@u��   ���   ���   ��3ME�� t   �_^[�����Q�L$+ȃ����Y�j>��Q�L$+ȃ����Y�T>����U����b3ŉE�j�E�Ph  �u�E� �D ��u����
�E�P�.���Y�M�3���8���Ë�U���4�b3ŉE��E�M�E؋ES�EЋ V�E܋EW3��M̉}��}�;E�_  �5`�M�QP�֋� ��t^�}�uX�E�P�u�օ�tK�}�uE�u��E�   ���u�u��$A����YF;�~[�����wS�D6=   w/�������;�t8� ��  �-WW�u��u�j�u�Ӌ�;�u�3���   P� G��Y;�t	� ��  ���E���}�9}�t؍6PW�u��1����V�u��u��u�j�u�Ӆ�t�]�;�tWW�uSV�u�W�u�� ��t`�]��[�� 9}�uWWWWV�u�W�u�Ӌ�;�t<Vj�s���YY�E�;�t+WWVPV�u�W�u��;�u�u��A��Y�}���}��t�MЉ�u�����Y�E��e�_^[�M�3��&7���Ë�U���VW�u�M��;���E�u3�;�t�0;�u,�A��WWWWW�    �L2�����}� t�E�`p�3���  9}t�}|Ƀ}$ËM�S��}��~���   ~�E�P��jP�����M������   ���B����t�G�ǀ�-u�M���+u�G�E���K  ���B  ��$�9  ��u*��0t	�E
   �4�<xt<Xt	�E   �!�E   �
��u��0u�<xt<XuG�G���   �����3��u���N��t�˃�0���  t1�ˀ�a����w�� ���;Ms�M9E�r'u;�v!�M�} u#�EO�u �} t�}�e� �[�]��]ى]��G닾����u�u=��t	�}�   �w	��u+9u�v&��?���E� "   t�M����Ej X��ƉE��E��t�8�Et�]��}� t�E�`p��E���E��t�0�}� t�E�`p�3�[_^�Ë�U��3�P�u�u�u9{uh�j�P������]�3�PPjPjh   @h�*�T��pá�pV�5P ���t���tP�֡�p���t���tP��^Ë�U��SV�uW3����;�u��>��WWWWW�    �/������B�F�t7V�����V���  V豱��P��  ����}�����F;�t
P��=��Y�~�~��_^[]�jh�M�"����M��3��u3�;���;�u�y>���    WWWWW�6/���������F@t�~�E��%����V�Q���Y�}�V�*���Y�E��E������   �ՋuV蟰��Y�jhN覔���E���u�	>��� 	   ����   3�;�|;@�r��=��� 	   SSSSS�.�����Ћ����<�`���������L��t�P�r���Y�]���Dt1�u�����YP�X��u���E���]�9]�t�=���M��j=��� 	   �M���E������	   �E��!�����u����YË�U����b3ŉE��ESV3�W�E�N@  �0�p�p9u�F  ��X���}𥥥�����<�ыH�����Ή}���e� �������ˋ]���׍<�0�P�H;�r;�s�E�   3ۉ89]�t�r;�r��s3�C�p��tA�H�H�U�3�;�r;�s3�F�X��t�@�M�H�e� �?�����<��P������Uމ�x�X��4�U�;�r;�s�E�   �}� �0t�O3�;�r��s3�B�H��tC�X�M�E�} �����3��&�H�����P�����������E���  �H�9ptջ �  �Xu0�0�x�E���  ������0�4?�H�����ʉp�H��t�f�M�f�H
�M�_^3�[��0����jh8N�����3�9x�tV�E@tH9�st@�E��U�.�E� � =  �t
=  �t3��3�@Ëe�%�s �e��U�E�������e��U�ב����������������U��WVS�M�tM�u�}�A�Z� �I �&
�t'
�t#����:�r:�w�:�r:�w�:�u��u�3�:�t	�����r�ً�[^_�Ë�U��V�uWV�����Y���tP�`���u	���   u��u�@Dtj����j������YY;�tV����YP�P ��u
�����3�V�����������`�����Y�D0 ��tW�):��Y����3�_^]�jhXN�{����E���u��9���  ��9��� 	   ����   3�;�|;@�r!��9���8�9��� 	   WWWWW�k*�����ɋ�����`���������L1��t�P�8���Y�}���D0t�u�����Y�E���S9��� 	   �M���E������	   �E��
�����u����YË�U��V�u�F��t�t�v�>8���f����3�Y��F�F^]�����̍B�[Í�$    �d$ 3��D$S�����T$��   t�
��:�tτ�tQ��   u��W����V؋
����~����3���������3�3ƃ��� �u% �t�% u��   �u�^_[3�ËB�:�t6��t�:�t'��t���:�t��t�:�t��t��^_�B�[ÍB�^_[ÍB�^_[ÍB�^_[��%������������̋T$�B�J�3��l-���3�	*������̋T$�B�J�3��L-����3��)������̍M��ء���M�С���M��f���M��f���M�鸡���M�鰡���M���p���T$�B��J�3���,����3�)��������������̍M��x����M��p����M�h����M��`����M�X����M��P����T$�B؋J�3��,���D4�9)������̍M��(����M�� ����T$�B�J�3��l,����4�	)������̍M������T$�B��J�3��D,����4��(��������������̍M�������T$��X�����T���3��,�����J�3��,��� 5�(�����������̋M������T$�B��J�3���+���,5�q(��������������̋M��x����T$�B�J�3��+���X5�A(��������������̋M��d#���T$�B��J�3��t+����5�(��������������̋M��4#���T$�B�J�3��D+���6��'��������������̍M��8����T$�B��J�3��+���D6�'��������������̍M������T$�B؋J�3���*����6�'��������������̋EP�M�Q�Ch����ËT$�B�J�3��*����6�H'�����̍M��X����M��P����M��H����T$�B��J�3��t*�����J�3��g*��� 7�'���M������M������T$�B��J�3��<*���|7��&������̍M��Ȟ���M�������M鸞���M��c���M��c���M�頞���M��m���M��m���M��m���M������T$�B��J�3���)����7�i&������̍M��x����M��p����T$�B��J�3��)���$8�9&������̍�|����E����������:�����|����/����������$�����D��������T$��<�����8���3��?)�����J�3��2)���H8��%������������̍����������������������T$��|�����x���3���(�����J�3���(����8�%�������������̋E�P�M�Q�Cf����ËT$�B�J�3��(���9�H%�����̋E�P�M�Q�f����ËT$�B�J�3��{(���l9�%�����̋EP�M�Q��e����ËT$�B�J�3��K(����9��$�����̋EP�M�Q�e����ËT$�B�J�3��(���,:�$�����̍M��������,��������M�������h��������M�������L��������M������T$��(�����$���3��'���P:�R$���������������̍M��X����T$�B��J�3��'�����J�3��w'����:�$���M��h����T$�B��J�3��T'����:��#��������������̍M��H����T$�B��J�3��$'���;��#��������������̍M�������E�P�M�Q�{d����ËT$�B�J�3���&���J�3���&���t;�v#���̋M��ș���T$�B��J�3��&����;�Q#��������������̍M��X����M��м���T$�B��J�3��|&����;�#������̍M��(����T$�BȋJ�3��T&��� <��"��������������̍M�������M�������T$�B�J�3��&���J�3��&���D<�"������������̍MD�8����M �0����T$�B�J�3���%�����   3���%����<�l"���������̋M��Ț���M����M����M��� �B����M���$�'����M���<�����M���T�A����T$�B�J�3��m%���\=�
"�������̋M��h����M��������M��� �����M���$������M���<�����M���T������T$�B��J�3��%����=�!�������̍�p���镙����t���銙����x��������M��w����M��_^���M��W^���M��_����M��wh���M��O����M��G����M��?����M��7����M��^���M��^���M������M������M��/h���M��'h���M��h���M������T$��l�����h���3��=$���>�� �������̍M�������M�������M���g���T$�B��J�3��$�����J�3���#����>� �����������   �������������_(��Í������c����������X����������M����������B�����$����']��������]���������!��������������� ����+g�������� g���M���\����p�����\����P�����\����`�����\����������f����������f����������f����������f���M��C������������   ��������M�����Ë��������   ���������4�������Ë��������   ��������M��d���Ë��������   ������4����B���ËT$������������3��g"�����J�3��Z"���?������̍�\����f����p����������|��������������������M�������M��������p���������M������������������d�����������������������������d���������,��������������t����������i����������^�����(����S����������H����������=����������2�����|����'���������������D������������������������������H������������������������������`���������������������@�������������^2����p����s�������������������������0���������P����w���������l�����L���顓����L����&�����������1����������1����d����5����������*��������������0��������������	�����$����N�����H�����c����p����Y���������Y����P����Y��������������������Y���T$��D�����@���3��������J�3�������?�r���������������̍M��c����x����m�����l����b�����x����W�����l����L�����x����A�����l����6�����x����+�����l���� ����M������M�����������������������#����������$����8����0���������0����X����~0���M��������l����������������   ���������x�������Ë��������   ��������������x���Í������0����x����a����M��Y����T$��l�����h���3�������J�3��r����B�������������̍M��(b���M���/���T$�B��J�3��<�����J�3��/����C�����������̋�0������������T����������8��������M������M�������p��������M������T$��,�����(���3�������J�3������C�O������������̍M��X����T$��\�����X���3��~���@D���������̍M�(����M�� ����T$�B��J�3��L�����J�3��?���tD�����������̋Eȃ��   �e���M��.��ÍM�������T$�B��J�3��������J�3�������D���������̋EP����YËT$�B��J�3�������D�^�����������̍M�鸒���T$�B��J�3����� E�1��������������̍������E"���T$������������3��[�����J�3��N���,E����������̍M�������T$�B��J�3��$���XE����������������̍M騐���T$�B��J�3�������E���������������̍M������T$�B�J�3�������E�a��������������̋E���   �e���M��X���ËT$�B�J�3������E� �������������̋E���   �e���M��h���ËT$�B�J�3��C���F���������������̍M��T���T$�B�J�3�����4F���������������̋EЃ��   �e���M�����ÍM������T$�BȋJ�3������hF�h�����̍M�8����T$�B�J�3������F�A��������������̍�����镐��������麄���T$������������3��`�����J�3��S����F���������������̍�8����E�����(����j�����T����/�����0����T����M������T$��$����� ���3�������F�������������̋��������   �����������������ËT$������������3�������J�3�����XG�4����|������   ��|�����M��2���ÍM��)����M��!����M������M������M��	����T$��t�����p���3��/���|G�����������̍�������������������������������������������T���������p���������������������������T$������������3�������J�3������G�>�����������̍M�H����M��@����T$�BȋJ�3��l�����J�3��_���\H�����������̋E����   �e���M������ËT$�B܋J�3��#�����J�3������H�����������������̋E����   �e���M�����ÍM������T$�B��J�3��������J�3������H�[��������̋EЃ��   �e���M��X���ÍM��O����T$�B؋J�3��{����H����M��|����T$�B�J�3��X���I�����T$�B�J�3��=����J�����Xth�Xt����                                                                                                                                                                                                                                                                                                                                                                                                                                                                  �W �W �W �W �W nW XW DW 4W "W W  W �V     \ �[ �[ �[ �[ �R �R �R �R �R �R �R  S S &S 6S DS LS bS rS �S �S �S �S �S �S �S �S T T ,T VT lT �T �T �T �T �T �T  U �[ �[ �[ �[ v[ ^[ F[ ,[ [ �Z �Z �Z �Z �Z �Z �Z lZ TZ BZ 4Z "Z Z Z �Y �Y �Y \ B\ R\ b\ x\ �\ �\ :T �Y �Y �Y �Y �Y zY pY bY VY HY 4Y (Y Y Y �X �X PX bX vX �X �X �X �X       �
  �� �  �  �  �	  �  �  �  �  �    �Q �Q     HR rR bR TR ~R     �V �V nV \V JV >V .V V V �V �U �U �V �U �U �U �U rU ^U �U 2U U �V �V �U NU     R "R �Q     X �W X (X                 d-A4�\+�        ��܉                D e l e t e     N o R e m o v e     F o r c e R e m o v e   V a l   B   D   M   S   bad allocation  0,($���+�� R%D,3�&��� �O�        �      F��P0����� � ��4�P0����� � ��      �      F��P0����� � ��      �      F˼"�hN�� � @Gp ,@C @U A   E M B E D   O B J E C T     I M G   n o     9�E�R�]�R�#]E�P�    ?cFKY�S@AZ�Fe3<+�ANC\LVD?N�]�5�*)O�]M�Y"INL�Q��'%ShX�G�L�Z�N%Y�=� �A�]�7GE�O�H�EOP'^C    1%4�/�/tCOS�O~JlE�C�E�:�E/*�G�A�E�4�    PeR2I,MOF��H�HH�    /Ft]�`S�GEQ�Y�A�A�FrR��DAJwB�H4L_K�    I s R o t a t o r P o p u p     I\�^4P�� �BAB�^s	�MAD�DAF�K�@�>A"F)Q��O�@�	qB�N�I�I��Y�C�W�      L,@C @U �,@C @U vector<T> too long  invalid map/set<T> iterator EM�K�F�E?C    6�E1SYL�^2P�@�    93'/*V6$0�)�8�)e9,(m@A3Z�A/Q�F�K�W�?�5J�A�A�N�X�W�2�$�Z�Y"QR@5H�Yd1fNEQ2\�IyO�E�<�4BU5JN      I n t e r n e t   E x p l o r e r _ S e r v e r     )HNZFu^�F.GeT�
@ UXxZKM�T�I�R�5O53DES�X�K�Ub    " "     +.D�,�Z�^�D�H/XBN�SB    >s+�&�6>�*�=R':\"�L	N3P�J[�J_@�Z�40�AB�H�H/ZwS9.cZETr^C�A�_42I�U"Q3E9J�N�=�)�Q�Y�JG�_�IQ28�(bQ�@�\TL�Y2�/hEEC�]�H�_2�-�EROjEeD3^�\�>�E^    8�N�Q�A�NAE�@�N�K�)�G�A�FeI�    (�U L�YRX�G]JUC�P4      -�.�4�)'�6��S�9� 	B�4 R"L�N4�C�[�WBS32          -�*�<C*�!�<<�Q�    I!N�AaF�B�I��I�S�K?W^�DU]�G�CM�C�K�OJuY2      "       "C|N4�T�T�Ir      	�2w*y(�#�&�:"52�6T�Y�_�N�Mc�>,=�RONG�OEl#��L�V8H���     wF�BOB�NqI�=LD�DAF�K�@�R2Q"F/Q�A�_�@�Y9]C\�N�Y�Y�R�Y�    map/set<T> too long     �/U �R �� �r �� `� p� Pz �� 0o  � �n ��  C �e ��  U  i �/P� �J pT �r �A t/@� P� �_ p] О 0B �� �,0� � 0� `� @� 0� �� �� � X M L   V"G�JVVRL�\�J�9?U�J	G�A�    c l i c k   f e e d _ c a p     c l i c k l i m i t     p r o v i d e r     n a m e     I F R A M E      
     !�I�A�QM�F~R��4DZyR�H5Z�BSp^ D�D�D�IqU�B)D�O� /X�}V�]'U�-H�GO^R@m]�[EK5BHsB�DTN�E4      vOv\p<�O�]HJSD%JEKT]      
�Je[8I�D�B%N��    V�H�B�^�C%JT�      �JcO�G9A�MKBeI��       6Q&N�RB]�N�HoL.-      O)@�    �]�D��    
�CANA64?C)L��    �D>L�X�0AiDt]    I"�QcF�B�Y�A�I�    ,   L'EI?J�<oNsM\C�IJK6?FFC�M�W$    F3B�DYMcKk=�L�Dn\$B�Y�_@�D    [tL�G�KeSCWDC1B�T�      H�DRH8?DIOMT _�I�VW      ^�[@E�H1R�H�=�Y%QRJ�          �A�������?�������?     @�@  �O^�K_�@1ULWr3OP�B�[�VE[�      3�+?'>�4W-6�'�3      =�S�K�_ZtI9EM�[�      I�HULJ$=_N�D�[�W�      I�DAM�;\cZ$OQV$US    D�LvO�3�F)A    I<Ha]�Z�2?]UPL�GQ[�I�:oC�]T[�J�DmR�U�      V�IyB]B�ZW�F!@]S0      E�@QV�RT1�OY[      J}N�]x8�HSILO�O�D{]s    E�@�^cP�@qBLGl6�A�MT    C#CEH#L+;�N�L�ZMnT4Bu_�      H�CA�@aV�      C�Aq]      ICDL@9E�B�2�]#VL�X$    A�L�P�ZBM�W�PS?�\#S$OQYT    @]K�QH9/J�I�W�QBAe]�^�      0,($���/�u �e �W � �� a f x _ c p c x d R t   F o l d e r V i e w     C o m b o B o x     S y s H e a d e r 3 2   S y s L i s t V i e w 3 2   S y s A n i m a t e 3 2     W o r k e r W   S H E L L D L L _ D e f V i e w     S t a t i c     0,($��L0UUUp] О 0B U80UUU@B @� P� �������� � 40,($���$5�3QB��`��ϝieframe.dll IEGetWriteableHKCU  a x 1   T E M P     LiO�B6_�D�I�A%^N4C�M�      '�.%'F�_$0�ZB�_�AEA�G�@�D�-�B/O�N�ET�=�J�UT@�    4�MN$G_`$QEnMD*F�D�C�     �E�K�N�@�C�J,Z��I�KFL    "�AqW�$AI�It.,M�K�C4    % d . % d . % d . % d   \   {   }   % x     C : \       % 0 2 . 2 x     �     �      Faӯ���> �O��n��4�e��J  �ǬM�     �      F�#?�>���; � ���H��+��) � =sR      �      F       �      F�@Qm6t��4 � `	�string too long invalid string position `0_RUnknown exception   t0�csm�               �        �ll    EncodePointer   K E R N E L 3 2 . D L L     DecodePointer   FlsFree FlsSetValue FlsGetValue FlsAlloc    7�0%5Rbad exception   �t ue+000      �~PA   ���GAIsProcessorFeaturePresent   KERNEL32    runtime error   
  TLOSS error
   SING error
    DOMAIN error
      R6034
An application has made an attempt to load the C runtime library incorrectly.
Please contact the application's support team for more information.
      R6033
- Attempt to use MSIL code from this assembly during native code initialization
This indicates a bug in your application. It is most likely the result of calling an MSIL-compiled (/clr) function from a native constructor or from DllMain.
  R6032
- not enough space for locale information
      R6031
- Attempt to initialize the CRT more than once.
This indicates a bug in your application.
  R6030
- CRT not initialized
  R6028
- unable to initialize heap
    R6027
- not enough space for lowio initialization
    R6026
- not enough space for stdio initialization
    R6025
- pure virtual function call
   R6024
- not enough space for _onexit/atexit table
    R6019
- unable to open console device
    R6018
- unexpected heap error
    R6017
- unexpected multithread lock error
    R6016
- not enough space for thread data
 
This application has requested the Runtime to terminate it in an unusual way.
Please contact the application's support team for more information.
   R6009
- not enough space for environment
 R6008
- not enough space for arguments
   R6002
- floating point support not loaded
    Microsoft Visual C++ Runtime Library    

  ... <program name unknown>  Runtime Error!

Program:        	
 !"#$%&'()*+,-./0123456789:;<=>?@ABCDEFGHIJKLMNOPQRSTUVWXYZ[\]^_`abcdefghijklmnopqrstuvwxyz{|}~ =   CorExitProcess  m s c o r e e . d l l         �         �       �  �       �  �       �  �       �  �       �  �       �  �       �  �       �  �        Complete Object Locator'    Class Hierarchy Descriptor'     Base Class Array'   Base Class Descriptor at (  Type Descriptor'   `local static thread guard' `managed vector copy constructor iterator'  `vector vbase copy constructor iterator'    `vector copy constructor iterator'  `dynamic atexit destructor for '    `dynamic initializer for '  `eh vector vbase copy constructor iterator' `eh vector copy constructor iterator'   `managed vector destructor iterator'    `managed vector constructor iterator'   `placement delete[] closure'    `placement delete closure'  `omni callsig'   delete[]    new[]  `local vftable constructor closure' `local vftable' `RTTI   `EH `udt returning' `copy constructor closure'  `eh vector vbase constructor iterator'  `eh vector destructor iterator' `eh vector constructor iterator'    `virtual displacement map'  `vector vbase constructor iterator' `vector destructor iterator'    `vector constructor iterator'   `scalar deleting destructor'    `default constructor closure'   `vector deleting destructor'    `vbase destructor'  `string'    `local static guard'    `typeof'    `vcall' `vbtable'   `vftable'   ^=  |=  &=  <<= >>= %=  /=  -=  +=  *=  ||  &&  |   ^   ~   ()  ,   >=  >   <=  <   %   /   ->* &   +   -   --  ++  *   ->  operator    []  !=  ==  !   <<  >>   delete  new    __unaligned __restrict  __ptr64 __clrcall   __fastcall  __thiscall  __stdcall   __pascal    __cdecl __based(    �������xl`���tT8XP�LHD@<8,($  ������������������������l`L,����lH( ��������pT4���tP, ���( n u l l )     (null)         EEE50 P    ( 8PX 700WP        `h````  xpxxxx          GetProcessWindowStation GetUserObjectInformationA   GetLastActivePopup  GetActiveWindow MessageBoxA USER32.DLL                                                                                                                                                                                                                                                                                        ( ( ( ( (                                     H                � � � � � � � � � �        � � � � � �                           � � � � � �                                                                                                                                                                                                                                                                                                               h ( ( ( (                                     H                � � � � � � � � � �        ������      ������                                                                      H                                      �������������������������������������������������������������������������������������������������������������������������������� 	
 !"#$%&'()*+,-./0123456789:;<=>?@abcdefghijklmnopqrstuvwxyz[\]^_`abcdefghijklmnopqrstuvwxyz{|}~���������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������� 	
 !"#$%&'()*+,-./0123456789:;<=>?@ABCDEFGHIJKLMNOPQRSTUVWXYZ[\]^_`ABCDEFGHIJKLMNOPQRSTUVWXYZ{|}~��������������������������������������������������������������������������������������������������������������������������������HH:mm:ss    dddd, MMMM dd, yyyy MM/dd/yy    PM  AM  December    November    October September   August  July    June    April   March   February    January Dec Nov Oct Sep Aug Jul Jun May Apr Mar Feb Jan Saturday    Friday  Thursday    Wednesday   Tuesday Monday  Sunday  Sat Fri Thu Wed Tue Mon Sun 1#QNAN  1#INF   1#IND   1#SNAN  SunMonTueWedThuFriSat   JanFebMarAprMayJunJulAugSepOctNovDec    CONOUT$     ������  �����EEE���  00�P��  ('8PW�  700PP�    (����   `h`hhhxppwpp           H                                                           b1I               `�+           �+�+�+    `       ����    @   �+ `        ����    @   �+           �+�+                \`,           $,0,�+    \`       ����    @   ,            |``,           p,�,0,�+    |`       ����    @   `,            �`�,           �,�,0,�+    �`       ����    @   �,            �` -       
   -<-X-�-.$.x.�.�./X/    �`	       ����    @    -�`       ����    @   t-          �-X-�-.$.x.    �`       ����    @   �-           �-�-�-    a        ����    @   �-            .�-    a        ����    B   �-,a      ����    @   @.           P.\.�-    ,a       ����    @   @.a       ����    B   �-Da      ����    @   �.           �.�.�-    Da       ����    @   �.a       ����    B   �-da      ����    @    /           0/</�-    da       ����    @    /a       ����    B   �-           �` -           �` -           �` -            �a�/           �/�/ 0�-    �a       ����    @   �/�a       ����    @   0           ,0 0�-                �`t-           �`t-             `�+            �a�0           �0�0    �a        ����    @   �0            �c�0           �0�0�+    �c       ����    @   �0        :
 D �n ~ �� ��  � X� �� �� � 8� x� �� �� � 8� h� �� �� � �� �� � V� �� �� � 1� �� �� �� (� i� �� �� �� 0� p� �� ?� 	� H� �� d� �� � �� ��  � Q� �� �� �� (� X� �� �� 	� 8� �� �� �� T� �� � �� �� )� �� �� �� �                                 X2   `2    <`    ����               @�     �2   �2�2    `    ����       �u      `    ����       �@           �� @           � ����    ����                  "�   �2   43                           �2              �2@           O� @           �� ����    ����                  "�   |3   �3                           l3              \3"�   4                       ���� �    (�   0�   8�   @�   H�   P�"�   h4                       ������    ��   ��   ��   ��   ��������    ��"�   �4                       ���� �"�   �4                       ����0�"�   �4                       ����p�"�   $5                       ������"�   P5                       ������"�   |5                           P     �5   �5�5�2    |`    ����    (   P�     \`    ����    (   p� ���� �"�    6                           P     h6����0�"�   <6                          x6�5�2    �`    ����    (   �� ����`�"�   �6                       @           �              �6����        ������    "�   �6   �6               "�   D7                       ������    ��   ��    ������������ �    �"�   l7                       "�
   �7                       ����h�    p�   x�����0�   8�   @�   H�   P�   X�   `�������    ��"�   8                       "�   l8                       ������������   ��   ��   ��   ������@�����K�"�   �8                       @           �Q              �8����        ������    "�   �8   �8               @           }�              09����        ������    "�   T9   @9               @           �              �9����        ������    "�   �9   �9               @           �j              �9����         �����    "�   :    :               "�   t:                       ����P�    X�   c�   k�   v�   ~�   ��������"�   �:                       ������"�   �:                       ���� �"�   ;                       @           ��             0;����P�           X�        "�   T;   @;               ������"�   �;                       ������    ��"�   �;                       ������"�   �;                       @           Hh @           {g "�   �<   h<                             4<            $<����    ����    ���� �              ����(�@           �� @           �� "�   ,=   =                             �<            �<����    ����    ����`�              ����h�"�   �=                       ������    ��   ��   ��   ��   ��"�   �=                       ���� �    �   �   �   )�   4�"�   (>                       ����`�    k�   v�   ��   ��   ��   ��   ��   ��   ��	   ��
   ��   ��   ��   ��   ��   ��   ��   ��   �����0�    8�����@�"�   �>                       "�   (?                       ����p�    ��   ��   ��   ��   ��   ��   ��   ��   ��	   ��
    �   �   �   �   )�   4�   ?�   J�   U�   ]�   |�   ��   ��"�Q   @                       �����    �   &�    &�   1�   <�   <�   D�   L�   W�   W�
   _�   j�   u�   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   �   �   �   %�   0�   ;�   F�    Q�!   \�    \�   \�   \�   \�   \�   \�   \�   \�   \�   \�   \�   \�   \�   \�   \�   \�   \�   \�   \�   \�   \�   \�
   \�9   g�:   r�;   }�<   ��=   ��>   ��?   ��9   ��9   ��B   ��C   ��D   ��E   ��F   ��G   �H   �D   �J   "�K   -�L   8�M   C�N   N�O   Y�"�   �B                       ������    ��   ��    ��   ��    ��   ��    ��   ��    �    �     �   �   �   �   &�   1�   <�   G�   R�   Z�   e�   ��   ��   ��   ������ �    �"�   �C                       "�   �C                       ����@�    N�   Y�   d�   d�    d�   l�   t�   �   �   �������"�   8D                       ������    ��"�   dD                       ����0�    I�"�   �D                       ������"�   �D                       ������"�   �D                       ������"�   $E                       ���� �"�   PE                       ����P�"�   |E                       ������"�   �E                       ������"�   �E                       ������"�    F                       ����0�"�   ,F                       ����`�    y�"�   XF                       ������"�   �F                       ������    ��������"�   �F                       "�   G                       ���� �    +�����+�   6�   A�   A�   L�������"�   PG                       "�   �G                       ������    ��    ��   ��   �   �"�   �G                       ����@�    K�   V�   a�   a�    a�����a�   l�   w�   ��   ��������    ��"�   LH                       �����"�   �H                       ����`�    y�"�   �H                       ������    ��"�   �H                       ������"�   I                       ����    ����    ������    ����    ����    ����    z    ����    ����    ����    S    ����    ����    ����    �    ����    ����    �����,�,    ����    ����    ����    �/����    �/����    ����    ����    t1����    �1����    ����    ����    �4    ����    ����    ����    �6    v6�6����    ����    ����]7f7@           D8����    ����                  �J"�   �J   �J                   ����    ����    ����    |9    �8�8����    ����    ����c;g;    ����    ����    �����; <    5    dK   pK�2    �c    ����       �@    ����    ����    �����A�A    ����    ����    ����%B)B    ����    ����    ����    �X    ����    ����    ����    v\    ����    ����    ����    �_    ����    ����    ����    |d    ����    ����    ����DgHg    ����    ����    ����    ur    ����    ����    ����    _�    ����    ����    ����    n�    ����    ����    ����    ��    ����    ����    ����    ��    ����    ����    ����    %�    ����    ����    ����    ��    ����    ����    ��������    ����    ����    �������    ����    ����    ����    K�    ����    ����    ����    ۯ    ����    ����    ����    e�        1�����    ����    ����    ��    ����    ����    ����    ��    ����    ����    ��������    ����    ����    ����    ��Q         �Q � �Q         <R � $Q         �R � `O         U 8  <Q         �V  (O         �W    �Q         8X � �P         BX �                     �W �W �W �W �W nW XW DW 4W "W W  W �V     \ �[ �[ �[ �[ �R �R �R �R �R �R �R  S S &S 6S DS LS bS rS �S �S �S �S �S �S �S �S T T ,T VT lT �T �T �T �T �T �T  U �[ �[ �[ �[ v[ ^[ F[ ,[ [ �Z �Z �Z �Z �Z �Z �Z lZ TZ BZ 4Z "Z Z Z �Y �Y �Y \ B\ R\ b\ x\ �\ �\ :T �Y �Y �Y �Y �Y zY pY bY VY HY 4Y (Y Y Y �X �X PX bX vX �X �X �X �X       �
  �� �  �  �  �	  �  �  �  �  �    �Q �Q     HR rR bR TR ~R     �V �V nV \V JV >V .V V V �V �U �U �V �U �U �U �U rU ^U �U 2U U �V �V �U NU     R "R �Q     X �W X (X     �RpcStringFreeW  �UuidToStringW RPCRT4.dll   VerQueryValueW   GetFileVersionInfoW  GetFileVersionInfoSizeW VERSION.dll BStrStrIW  � SHSetValueW � SHDeleteKeyW  StrCmpIW  YUrlEscapeW  SHLWAPI.dll �lstrlenW  C CloseHandle �SetEvent  � CreateProcessW   GetProcAddress  �LoadLibraryW  ExitThread  dWaitForSingleObject � CreateThread  u CreateEventW  3OpenProcess !Sleep �GetModuleFileNameW  � CreateMutexW  MGetSystemTime �GlobalFree  �GlobalAlloc �LocalFree �LocalAlloc  �InterlockedIncrement  �InterlockedDecrement  �lstrcmpW  *SystemTimeToFileTime  �GetLocalTime  �LoadLibraryA  LFreeLibrary ExpandEnvironmentStringsW zWideCharToMultiByte MultiByteToWideChar YGetTempFileNameW  fGetTickCount  �GetEnvironmentVariableW \VirtualQuery  yGetVolumeInformationW �GetWindowsDirectoryW  IGetSystemInfo KERNEL32.dll  � DispatchMessageW  MsgWaitForMultipleObjects PeekMessageW  �TranslateMessage  �GetWindowRect �GetWindowInfo oGetSystemMetrics  � EnumWindows �SetWindowTextW  PRemovePropW \GetPropW  �GetWindowThreadProcessId  cSendMessageW  PostMessageW  fSetActiveWindow �SetWindowPos  �SetPropW  �SetWindowLongW   CallWindowProcW .RealGetWindowClassW � EnumChildWindows  �GetWindowTextW  rSetCursorPos  ]SendInput GetCursorPos  GetClassNameW USER32.dll  *RegCloseKey xRegSetValueExW  [RegOpenKeyExW BRegDeleteValueW 6RegCreateKeyW hRegQueryValueExW  � CryptReleaseContext � CryptGenRandom  � CryptAcquireContextW  � CryptDestroyHash  � CryptGetHashParam � CryptHashData � CryptCreateHash ADVAPI32.dll   CoCreateInstance  k CoUninitialize  > CoInitializeEx  g CoTaskMemFree ole32.dll OLEAUT32.dll  ZRaiseException  -TerminateProcess  �GetCurrentProcess >UnhandledExceptionFilter  SetUnhandledExceptionFilter �IsDebuggerPresent �RtlUnwind �GetCurrentThreadId  oGetCommandLineA �GetLastError  �HeapFree  �HeapAlloc �GetModuleHandleW  4TlsGetValue 2TlsAlloc  5TlsSetValue 3TlsFree �SetLastError  �GetModuleHandleA  �WriteFile ;GetStdHandle  �GetModuleFileNameA  [GetCPInfo RGetACP  GetOEMCP  �IsValidCodePage �LCMapStringW  ExitProcess �SetHandleCount  �GetFileType 9GetStartupInfoA � DeleteCriticalSection JFreeEnvironmentStringsA �GetEnvironmentStrings KFreeEnvironmentStringsW �GetEnvironmentStringsW  �HeapCreate  �HeapDestroy WVirtualFree TQueryPerformanceCounter �GetCurrentProcessId OGetSystemTimeAsFileTime �LeaveCriticalSection  � EnterCriticalSection  TVirtualAlloc  �HeapReAlloc �SetFilePointer  �GetConsoleCP  �GetConsoleMode  �HeapSize  �GetLocaleInfoA  �LCMapStringA  =GetStringTypeA  @GetStringTypeW  �InitializeCriticalSectionAndSpinCount �SetStdHandle  �WriteConsoleA �GetConsoleOutputCP  �WriteConsoleW x CreateFileA AFlushFileBuffers            <��H    
]          �\ �\  ]   @  P  p ] ,] >] P] X]       BannerRotator.DLL DllCanUnloadNow DllGetClassObject DllRegisterServer DllStub DllUnregisterServer                                                                                                                                                     4D    .?AVbad_alloc@std@@ D    .?AVexception@std@@ D    .?AVCAtlException@ATL@@ D    .?AVlogic_error@std@@   D    .?AVlength_error@std@@  D    .?AVout_of_range@std@@  D    .?AVCBannerRotator@@    D    .?AVCLiteBHO@@  D    .?AUIObjectWithSite@@   D    .?AUIUnknown@@  D    .?AUIDispatch@@ D    .?AUIOleCommandTarget@@ D    .?AUIDocHostUIHandler@@ 44D    .?AVMyClassFactory@@    D    .?AUIClassFactory@@ 4444444D    .?AVtype_info@@     4N�@���Du�  s�                                               	               	      
                                                !      5      A      C      P      R      S      W      Y      l      m       p      r   	         �   
   �   
   �   	   �      �      �   )   �      �      �      �      �      �      �                 4            ��������4D    .?AVbad_exception@std@@     o�o�o�o�o�o�o�o�o�o�          x   L	    
   �   \   ,      �   �   |   D      �   �   `    (!   0"   �x   |y   lz   \�   X�   H                                                                                                                                                                                                                                                                                                                                    abcdefghijklmnopqrstuvwxyz      ABCDEFGHIJKLMNOPQRSTUVWXYZ                                                                                                                                                                                                                                                                                                                                                                                                                                                       abcdefghijklmnopqrstuvwxyz      ABCDEFGHIJKLMNOPQRSTUVWXYZ                                                                                                                                     �d�  `�y�!       ��      ��      ����    @~��    �  ��ڣ                        ��      @�      �  ��ڣ                        ��      A�      �  Ϣ� ��[                 ��      @~��    Q  Q�^�  _�j�2                 ������  1~��    <$����C                                                                                              �i            �i            �i            �i            �i                              �o        8"�&@(�n�i   �i�d�d    �����
                                                                   x   
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                            ` P  �                    8":$h*d*`*\*X*T*P*H*@*8*,* ***** *�)�)�)�)�)�)�)�)�)�)�)�)�)�)�)�)�)�)�)�)t)p)l)`)L)@)	         �n.   �oH~H~H~H~H~H~H~H~H~�o   .                    ���5      @   �  �   ����                         �p     ����    PST                                                             PDT                                                             Pp�p����        ����        ��������         �@         �@         �@        @�@        P�@        $�@       ���@        ��@     ���4@   ������N@ �p+��ŝi@�]�%��O�@q�וC�)��@���D�����@�<զ��Ix��@o�����G���A��kU'9��p�|B�ݎ�����~�QC��v���)/��&D(�������D������Jz��Ee�Ǒ����Feu��uv�HMXB䧓9;5���SM��]=�];���Z�]�� �T��7a���Z��%]���g����'���]݀nLɛ� �R`�%u    �����������?q=
ףp=
ף�?Zd;�O��n��?��,e�X���?�#�GG�ŧ�?@��il��7��?3=�Bz�Ք���?����a�w̫�?/L[�Mľ����?��S;uD����?�g��9E��ϔ?$#�⼺;1a�z?aUY�~�S|�_?��/�����D?$?��9�'��*?}���d|F��U>c{�#Tw����=��:zc%C1��<!��8�G�� ��;܈X��ㆦ;ƄEB��u7�.:3q�#�2�I�Z9����Wڥ����2�h��R�DY�,%I�-64OS��k%�Y����}�����ZW�<�P�"NKeb�����}�-ޟ���ݦ�
       �D        � 0     ����   ;   Z   x   �   �   �   �     0  N  m  ����   :   Y   w   �   �   �   �     /  M  l                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �   8  �                 P  �                 h  �                  �                 	  �   �� t  �      � Z  �      t4   V S _ V E R S I O N _ I N F O     ���             ?                        �    S t r i n g F i l e I n f o   �    0 0 0 0 0 4 b 0   $   C o m p a n y N a m e         6   F i l e V e r s i o n     2 ,   1 ,   1 ,   0     :   P r o d u c t V e r s i o n   2 ,   1 ,   1 ,   0     D    V a r F i l e I n f o     $    T r a n s l a t i o n       �<assembly xmlns="urn:schemas-microsoft-com:asm.v1" manifestVersion="1.0">
  <trustInfo xmlns="urn:schemas-microsoft-com:asm.v3">
    <security>
      <requestedPrivileges>
        <requestedExecutionLevel level="asInvoker" uiAccess="false"></requestedExecutionLevel>
      </requestedPrivileges>
    </security>
  </trustInfo>
</assembly>PAPADDINGXXPADDINGPADDINGXXPADDINGPADDINGXXPADDINGPADDINGXXPADDINGPADDINGXXPADDINGPADDINGXXPADDINGPADDINGXXPADDINGPADDINGXXPADDINGPADDINGXXPADDING   |   00'0Q0X0�0v2�2s3�3�3�3�3>4Y4h4�4#595U5�5�56�7�78K8�8�889�9�9�9�9�9�9�9U:�:�:�:�:�:�:3;I;b;s;�;�;<1<i<{<l=�=6>H>    4   #020?0�0)1;1L1~1�1a2�223]3{3�3�3424Q4�;D<�? 0  �   /0�1�1)2R2~2�2�2�233�3�3�5�5�6�677;7�7`8f8o8�849S9h9�9�9�9�9�9�9�9::&:6:F:V:f:[;�;
<<<#<�<�<�<==W=/?5???E?S?�?�?�?�?�?   @  d   t0�0P1\1�1�1C2P2u2�2�2E3�3�3�3(4Y4�4t5�5c6q6�6%7G7c7�7�7�7s8�8�<�<+=K=i=�=\>o>�>�>�>�>?�?   P  �   �0�0%181v1�12�2�23s3�3�3444S5b5o5�5�5*6H6�677"71787r7�7�7�7�8�9�9C:i:�:�:�:�:�:";8;�;�;�;�;�;�;�;B<T<�=�=�=1>J>O>V>�>�>?�?�?   `  <   0H0U0�2�2�2#414T4�5�5�5649c9q9<:N:f:x:;;]<n<�>   p  `   1272g2�2�2343E3�3c4q4�4�4�4�4�4�5�5�5�566�7�7�7�78�8�8s:�:;�;	<y<�=>>T>�>�>y?   �  `   �0�0�0T2a2r2y2�2�2�23�3�3 4>4[4k4�56s6�6�6�768`8�8�8�8�9�9S<a<�<==B>S>b>q>�> ?8?�?   �  X   #121A1W1�4�4�4525f56q6Z7m7�7�8�89'9�9�9c:v:M;|;�;�;�;�<�<�<�=�=�=�=�>??�?   �  D   00�0�0�0�0�1�1�1�2�4�4s5�5�5x6�6�67:(:�:�;�;�;<�<�=�>�? �  ,   1�576�8-:s:�:�:#;6;�>�>g?�?�?�?�?   �  �   t0Y1�1�1�1�1�1�12#222@2]2t2c3u3�3 4�4�45X5_5q5�5�5�56>6G6�6�6�6+828�8�8�:�:�:�:�:�:�:�:�:�:�:-;h;q;w;~;�;�;�;�;�;$<t<�<�<�<�<�<C=V=|=�=�= �  |   m0z01#1�1�1�1�12^2}2`3n3�3�3l4_5s5�5�5�5�5�6�6�6f7m7�78L8`8�8�8�8#959U9\9c9j9:C:V:w:�:�:K<�<=�=�=C>V>�>??*?   �  <   11@1|45&5L5}5�5W8�8#:5:G:�:�:,;Q;�;<#<1<k<�<�<�<�> �  l   0!0�0�0�0�0�0�011�1�1�3�3�34444434E4W4�4�4&5z5�5�5	66�6�6
7Z7v7	9N:y:�:�:�:`;t;�;�<�<==;=   �   W0z0�0�0�011!1a1t1�1�1�1�1�1�1g2y2�2�2�2�2�2�233(393C3`3j4~4�4�4B5Z5�5�5607�7�7w8�8�8�8�8�8�8
9:9@9H9U9i9�9�:�:�:=&=_=n=s=y=}=�=�=�=�=�=�=�=�=�=�=�=�=�=�=�=�=>O>h>o>w>|>�>�>�>�>�>�>�> ??????^?d?h?l?p?�?�?�?    �   000010[0�0�0�0�0�0�0�0�0�0�0 1111W132;2P2[244$4X4p4x4~4�4�4�4515I5�5�5�67'797�7�7�7�7�7�78j8�8�8�8�8�8�8�8�8#9A9H9L9P9T9X9\9`9d9�9�9�9�9�9&:1:L:S:X:\:`:�:�:�:�:�:�:�:�:�:�: ;J;P;T;X;\;<"<r<x<�<�<�<)=I=N=,?3?   �   @0'161Q1v4�5@7p7�7~9�;�;�;�;�;�;�;�;�<j=s=�=�=�=�=�=�=�=�=�=>>>.>5>I>P>h>t>z>�>�>�>�>�>�>�>�>�>�>�>�>??"?/?R?g?�?�?�?   0 �    00"0:0`0�0�01?1G1�1�1�1�1�1�1�1�1�1�12!2&2.242;2A2H2N2V2]2b2j2s22�2�2�2�2�2�2�2�2�2�2�2�2�2�2�2�2333,3L3R3n3�3�3404Y4^4u4�4�455/5�578_8�9z;�>�>�>   @ l   �0�122:2E2�2�2�2�2�2�2�2�2�2�2�2�2�2�2333$3)3/393B3M3Y3^3n3s3y33�3�3/6�6�6&<�<�>�>�>????   P �   �0�0�0�1�1�1�1�1 282C2g2p2w2�2�2�2�2373J3b3t3�3�3�5�5L6�6�68$8^8k8u8�8�8�8�8�8�8�89999p9�9�9(:E:�:�:;�;�;�;�;�;�;�; <<5<><D<M<R<a<�<�<�<�<�=�=>k>�>?h??�?�? ` �   0/181D1{1�1�1�1�1�12282S2Y2b2i2�2�2�2333%3/363A3J3`3k3�3�3�3�3�3�3454:4E4J4h4�45
55?5E5w5�5�56 6H6a6�6�6�667<7`7~7�7�7�7�7�7L8W8a8r8}80:A:I:O:T:Z:�:�:�:�:;;;$;[;�;�;�;<<<=<B<v<{<�<�<�<�<�<�<�<�<�<�<�<�<�<=�=�=�=�=�>�>�>�?�?�?   p �   0[0u0�0�0�0�0�0�0�0�0	111D1R1X1{1�1�1�1�1�1�1�1�2�2�2�2 555.535B5K5X5c5u5�5�5�5�5�5�5�5�5�5�5�5�5�5�566 6.656:6C6P6V6p6�6�6�6�6�:�:�:�:8;};P=[=c=�=�=�>??5?S?�?�?   � �   y0�0�1�1�2�2$3�4�5[6�6�6�67�7�788�89&9,9F9U9b9n9~9�9�9�9�9�9�9�9::6:i:x:�:�:�:;6;X;�;�;�<�<D=�=(>`>�>�>�>M?Y?�?�?�?   � |   �0�0�12�2�4�6�6�6�67;7I7�7�7�7�7�7�7�7�7f8o8u899 90959M9S9b9h9w9}9�9�9�9�9�9�9 ::::�;�;�;>>,>8>B>J>U>�>�>L?�? � �   0�0n1�1 222)212>2E2u23�3�5�5�5�5�5�56606B6717�7�7�7�7�7O8�8�8%9+9|9�9�9�9�9::V:;;;=;Q;W;�;�;�;�;#<�<�<�<=p=�=�=�=3>>>l>z>�>�>�>�>�>�>�>�>�>?
? ?;?H?i?u?�?�?�?�?   � L   �0�0�0�071�2�24*4�5�6�6Y7;8�8�8|9�9�92:I:�:�;�;�<=>>�>�>�>v?�?�? � 4   J0313|6�6�6�6�6�6�6�6�6�6�6�6�6�7�7�7�7C8g8 � P   q2E4b4�4�4�4�5�5{8�8�8�8�8�8�8�8Y9�9:):`:j:�:�<�<�<�<x=�=�=�= >4>c>�?�? � `   0j0�0�01]1�1�1�12J2z2�2�2"3�3�3,4{4�4�45C5�5�5
6:6�6�6�6
7L7�7�7Q8!9g9;�=�>/?�?�?   � @   0p0�0�01:1j1�1�12J2�2�23l3�3/4�4�4H5�5�56!6,60656     �   �2�2�2�2�2�2D3H3L3P3T3X3\3`3d3h3l3�3�3�3|5�5�5�5�5�5�8�8�8�8�8�8�8�8�8�8 99999999 9$9(9,9094989<9@9D9H9L9P9T9X9\9`9d9h9l9p9t9x9|9�9�=�=�=�=�=�=�=�=�=�=�=�=�=�=�>�>�>�>�>�>�>�>�>�>�>�>�>�>�>�>�>�>�>�> ???? ?$?(?,?0?4?8?  �    1$1(1@1D1h1l1p1�1�1�1�1 22�>�>�>�>�>�>�>�>�>�>�>�> ???????? ?$?(?,?0?4?8?<?@?D?H?L?P?T?X?\?`?d?h?l?p?t?x?|?�?�?�?�?�?�?�?�?�?�?�?�?�?�?�?�?�?�?�?�?�?�?�?�?�?�?�?�?�?�?�?�?      00000000 0$0(0,0004080<0@0D0H0L0t;x;�;�;�;�;�;�;�;�;�;�;�;<< <$<(<0<H<X<\<l<p<t<x<�<�<�<�<�<�<�<�<�<�<�<�<===== =$=(=,=0=4=<=T=X=p=�=�=�=�=�=�=�=�=�=�=�=�=�=�= >> >$><>L>P>T>\>t>x>�>�>�>�>�>�>�>�>�> ???,?0?4?<?T?X?p?�?�?�?�?�?�?�?�?�?�?�?�?�?�?   0    00(0,000D0H0X0\0l0p0�0�0�0�0�0�0�0�0�0�0�0�01T2\2d2�2�2�2�2�2�2�2�2�2�23 3D3X3h3x3�3�3�3�3�344 4(40484@4L4l4t4|4�4�4�4�4�4�4�4�4�45(545T5`5�5�5�5�5�5�5�5�5�5�5�5660686@6L6l6p6t6|6�6�6�6�6�6�677(7H7P7X7`7h7p7x7�7�7�7�7�7�7�7�7�7 8888 8,8P8p8x8�8�8�8�8�8�8�8�8�8 999<9P9`9t9|9�9�9�9�9�9�9: :4:<:X:x:�:�:�:�:�:�:�:�:�:�:;;<;P;X;h;|;�;�;�;�;�;�;�;<0<@<L<T<x<�<�<�<�<�<�<�<=(=@=X=d=�=�=�=�=�=�=�=�=�=�=�=�= >>,>4><>D>L>T>\>d>l>t>|>�>�>�>�>�>�>�>�>�>�>�>�>�>?,?4?<?D?L?T?\?d?l?t?|?�?�?�?�?�?�?�?�?�?�?�?�?�?�?   @   00 0(00080@0H0P0X0`0h0p0x0�0�0�0�0�0�0�0�0�0�0�0�0�0�0�0�0 1111 1(10181@1H1P1X1`1h1p1x1�1�1�1�1�1�1�1�1�1�1�1�1�1�1�1�1 2222 2(20282@2H2P2X2`2h2p2x2�2�2�2�2�2�2�2�2�2�2�2�2�23333$3,343<3D3L3T3\3d3l3t3|3�3�3�3�3�3�3�3�3�34444$4,444<4H4h4p4|4�4�4�4�4�4�45(545T5`5�5�5�5�5�5�56606<6\6d6p6�6�6�6�6�6�6�67$7,747<7D7L7T7`7�7�7�7�7�7�7�7�7�7 8888 8(80888@8H8P8X8d8�8�8�8�8�8�8�8�89$9T9X9x9�9�9�9�9�9: :,:H:h:p:t:�:�:�:�:�:�:;;;,;0;L;P;X;`;h;l;t;�;�;�;�;�;�;<(<H<d<h<�<�<�<�<=(=H=d=h=�=�=�=�=�=�=>0>L>P>p> `     00 0<0\0|0�0�0�0�01,1D1d1�1�1�1�1�1�1�1�1�1�1�1�1 2�3�3�3�3�3�3�3�3�3�3�3�3�34444$4,444<4D4L4T4\4d4l4t4|4�4�4�4�4�4�4�4�8�9@:P:`:p:�:�:�:�:�:�:�:�:�:�:P<X<�>�>�>�>�>�> ???????? ?$?(?,?0?4?8?<?@?D?H?L?P?T?X?\?`?d?h?l?p?t?x?|?�?�?�?�?�?�?�?�?�?�?�?�?�?�?�?�?�?�?�?�?�? p    �0�0                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    