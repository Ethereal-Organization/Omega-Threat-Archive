MZ�       ��  �       @                                      � �	�!�L�!This program cannot be run in DOS mode.
$       �IW��(9��(9��(9��45��(9��72��(9�C47��(9��73��(9��7=��(9�(73��(9��(8��)9�'d��(9��2��(9�.?��(9�?=��(9�Rich�(9�                PE  L ��.H        � !    �      �                               @                              PW ^   P�     � �(                  ��                                                                                                 �                 @  �         @      8   �              @  �         0   `  
   �              @  �.rsrc    0   �     �              @  �             �     �              @  �.data    P  �  D  �              @  �.adata      0      >             @  �                                                                                                                                                                                                                                                (;����H��T�g�y8Y.�ֈ�����3׀����_5��� �j9��s	,��6���f�̲8>~��j�Q��dP�Wxj���:[�{%��S�"�vQ�=iъ>4�Up����h[	�Sz�z�f��6�:�ic�Aԛ�A��V��b<M�~g;���������"߸m�M4���>���<��&Hh�G��H�ƅ.��DQeZ1�N�SL�tf�}�N�
�TVG�PyƁe�+�	��1��6J��ɪ��9��_�5���m(�/��T����(������A����q��g0���;�J��ߝ������{�xzq�'C����!jr�۰��>�V�N��b!���)�Ѕ�&O@�� �QWò4 ���!ƛ�\5B�S���{�z	|;�6��ȑk�������C��Zf�2s-����)�&��j��"{�F�:E�]�4~���_�\ٜS��n�;ov�TA5-Pچ�@m밠���љ�1�I����<�n=AB����h��$�?�k�##��2�F/�q�y�8-&���$���J$۸!dNC�5�5f�ޢHK5���j��uE�i��Kh,�#�58P%��A�jw�?U�Q���4f2V��{����u��j7��[��	�q�ى�����b$[>� %��HJ��+)����=�6c5�
d�(����Y���J�3ʅkI:�q!C�}s�.]܁���<�x��X�L#��ʹ/���\6@�����/��n�����5[S����x���"��:+ ����Ύn��L��H=K�p��Q�q����~��FF�hI"a�i~۟0W��|*�DHu�kF�Bz�P��J&�����׵��������9��0)�ƕ���?�Y�^���� �u8	_����C���%8���@�i�z�ny 0 C��e������ ��,b�C�����[�h�=j�(`����3"�ߢ[=!��D���"���^nʶxE��7I��΋�f�X�@?���L��@��pQ"�g�Y�B<��� �r\B��}�|p��BU�>D�%٘��Ʈ�;FC@b��v��Z�����D0��|%��E�7A�˘��Q2?�]�Ƒ�$�?��et�KU�r��|n&o<T����Wp��V��׻�� ��������S��P8;�:h�ھ�x!>�Cm���Wr�%Y�f1�a�@ѫ��u i��;V���N���	@j(qS<���S�a�MH��-|�SHMǛ�U��%g��bh�;*3��x�C�7.�K�������햾/��@vNT+)�Y�dA��܀ڸ�������^n^���xQˋ�t}��ѻ�h�ec�z�bU��>�7�����!UԀ8��O8�o���q290Z���Ӗ,+k���CM���J��YA%���L1D�p<�\�/�)�%� G�gm��	�A#@$X׽�Z�!L����'���S��ډA����;v)}��3�v~���x�[��Y?G	q�m�Z�"�|�Wm�?�r�9CVA�t��{Cg>~�O�J�N'g������8��۾ oh�X�+kX�~C�c���$�G$�B:��ֆ�����nAޑ
����:Hf1�\���h{�G)[]#���!�c�����l�#���۔�=	?Tq�G��80͒U�W>�^�2M{Q��/���'$�35�,�~���ؘ�rt>Ad�@i3dU�v�ɍ�q��x
�^����q\:¬v؎&��:��g%�v�E@��]�� �MS
U �h���a�쨒���6�>o�5�D�9)?w}�qK$��q$�3a[J#��=aU �����0Mm��B</�R��:4�R��ӑ�7e�ϴ,p��+��cu@�zy�j���28D���u�%*�Lu<��1E�@��Χ;VY��B_��:��dE2�BB]��"��	��M"�U��&&�ؠm3��9���8+f�ng+�%�y:-�sI�/��_�T�E��V`��Qu��K�É
��wl��j7�'.`1&�??$�Y�ӳ.�`�G+\v[^���{��[ _�O�;��,���9������))��g�tX���A!�����\2{y}�����BE�d��tT�zh�C3��E��'x���=A����q����5iDRP��辇޳:�{m��+�N�(��.��9�3���LB�j�}�ɹ�zƼ�|M��u��d�tӔ%��oX���	�X�}�����3�t������v�t
5/���x�M�tR�.�1�i� B}��˟˙���dB�~��`F�fܱK�1��	bQ;=iC�?����ZJ��֔$�v5k�ԧ�`��C���z��q-ˢ0O�Yc��i���s�HFu��Y�%�K�@W�J�W��ʰ��Tf��A�Y�N-�pj����7Q��2�YV����;��@�K$�+IM� {N
�y�&��Rh[_tv�O�/��L����d��c�'�Bq��42/4ij�����Z��Y|w6�oj����t�9��q��Qzt�[ a�Mˋ�u�� `���蜮�	���4�0Z���&B�hkP�ȇ�f��&���
�f��eL�����8SЊ`�[���1λS�\�eg4o-�Jiy��s�GS��2�<ߌ�)*����S�����N�ɟ���^rlY����jz������@��5-���S\:�1afYlܚh)AO�ce�H��?�=�J��" xǪI�J�6��� N�	=����om8�Q�q�v�+��C�z�Օ��!��Pߦ; Ǌ2��_7m�g�Ys���@g��E,�q�6��U�q������_(��
ߋ�.:�[e��i��٣p��_��˙�6)��3���˅߃8qf�x4�Y*ӓݲtܛkn�d84�.�>���AqS;�E�T~E�.����1�`�*�A׸S�c��W-"am�)CnRB��κ�$g��F�����X	N��1P7���.�f߁@v��_9I�ɑ� ���硏�U�~<�������R9��@���w�
�m�?����n
����
.Ƴ��`���2��0`M)	� ��cv���B_��$mQ'��uRNY,:m.f�[늃G�~�\�oE�k��=Bf+�}�����)6��0��O
���>	-���]�J2|���0��xŨ�:++>"ih*j~�<��m\��G$c�r�/�[	�W�w�c!�����j�55���=5s)������ґ�%8��(l��#�ή�b�g�S�V�I�����D	!NĘh�`�|X�)X���ma���p��(�ZA�(��g|m�d
g���eD�t!&LdF��}㪪��{��- �!�
��5`���!	�nNud�hrN��>��R��PuN�D=P;�!�90X-U�oڿh�н��;%�0ua��|܄M!�Qb��vm�߬b+��A���M�e)g��(��W��"�DAwޖ�8� n����:C�u�&������1c��f�H���/�ay����NX6ݐ�<���� d��FK²�IYQM��IÌ2����#�&�$���D��!R>n�]!�nJ��%C��$z�*�:���<RIV��b�lK��ⳛ%v��b|词)�-M&�n���'���1iLi�P�\.�	��LعwO��Sb�}�g�Z����Z<.G��> gƀ3���ܖ�O�ۜ"0��W���Y��C�֖D�U�l��k5���S>7�X�~X.q|"7����~�^���s�l�V=M��c�Q5H�G�v�ՈJAEnW�2���N��8Ϸ��`�!-�s�{v3�n~�^���jH1��{�h��	E�tA&6��Y��Vʭ����#�T��9���P���Hj���kc����
ɤc�K�*�|\I�<����M��~3�r���rgL�s��Ta��c��JZ��8c�����%��
�;�f|p�����>Te����C��heR�%"_�ɠܓ�ui�o�Z��%b_��F{�rPΪ�+��*q�U�)�m��k%M�(�ָ�.�$��l�~L(?A�2m4+X��X����ƺ�#V��d��M�l�j݀uZ�hs(Ӻ��a��u��m�<���������Mv+�MJ��{��/\��/,	0�%��f�k�(���,��Ֆ�.�慈ǡ�SoZ%�G�נ�*�t���RPV��w��x���"F���Y����"﷙!K�'M�]e�����p���������K�N[Lc�P��B#��Ϡ�ꓧC�_m�]#YT�����eq�v�J��Ek@�0la� Ad�r{\�:P�RM*ҍD�L\,2ԠX\�/$��!�4��1�,X�f�*�r�7�$����ZzG�U�B�t�:+��*!\�
����L�F�!gz�wktɰa�([���cc��/=R�-b��E�?d;�B�g��aL�h��t����L�B�=h^5��$��G�7U��}U���`�E�7�b���+n�~�&MAJ�'J��X�Y�S��`�֔��g��F0���@����,�Εv8�����U���?�N��9�����6�P^~��x��B���:�|�k�|bI_����'�;%_�w2��������3�[�B~M~��ө��9j���j=ѡ�g��?!|��l)=�R�`����*p]/Gy���m~��$ ��X�E�u�U/�<*0n۪�������s}��+�+�~�7���f�)�@L��+t�^�i	LZ��n��N��Tr��5Oގ��V�k�� ���{��++
�U��x6��&�D^��O�2���y�����f/-�d0���z+�����@9�2KersV��R��x=�٩��ە>�m�E�}hT�)�F��p��, �$��z��#�r�&��r���z�:�ԟ��N�/T�k���H'?��\5�;���K�UܾY&�!��^����4�\��v �&\(���
�9�ɢ�g�1���7~�)$��/͂�AԎ8D�:e�c�G}��P-kH��P�I.�U���aQ�ߴpc�'�o�AD}�*;��̦xA�US�ɥ�:,��c'�iM���x�&���F6��bC����΂�!z%H�@z�Wټe�5,!�Y�L�sj&,�Tŏ��g���/r(�L�˥b[�����qΟ����)3�e_��߾�kt�q���DF:�� �"M����4���D
[�=�&�����ݰ#�P�:[o�(�K�2~�JK�����"�3��|����ę�3�z��p�� �il���������ҵ3��P.���@j��{�k��^�A�e��X�b��X�A5sّ2���=��[	<p���u��ޢ�&�� P���Zq�e�P6���5ad�������?}��4��9~x���Bɦ�>��mȣ������T
+��V�+�Y�E�L҇���ef*�oj��P�|�p�6��6���^˩��;���h.$:a� �BiX�\���(�\��	�t�F�섹��uHy \���%e�0�y�*`c�v͘�G�)�uI�tr`)��c��V�8�����*�Z��>'f�����l��������"�<g��NF��~n$�I^m8����ƾ�-J� �!�>Y{jd��w��L�o�1@��g'��@怸�ܘ���z��[�b���z.��t�z2K���o]ݚ�1n"�O�����f�I�ID|��^e6��D�/������	�b|��U�<��U�r��=�B�$_l��Rr���Sk^�7�Ѵ���a�3C{��K�8�qƩ5��p����T���nxӬGM)�-J��,m�(�7��%��CQ�_�L����:�h-�'��u��(^粃,�*1Jy�?&�s�;��$b�R{2C촴O%�Zl�<dT�b��c�a�HJ��_o��a�&Sv����V�Tĳ��X԰cZ�q�~��X�� �˃��V+�`��^9*��埉�&-����螡�ޅu�p�{���3�F�gZJ�<l�4��e��I���굥8�W�f|�\f��n����-Q1��]֌]i���z|���7Is3���
�³��17��ڷ2��~�0Oe��ǥ-'6�����OB�g����QR�!��"*���U�L� g��!�0�W���4ާ�;r�L�m��h*�C͎mfc*�td8hHE���"T��� ]�ws(�4��2�f�k�=/���߮� "���bRr;~2P1�����,e���eF�p�f[�- Ԟ��*��0צ�32��WM���#U�¯]�7����
��E�����k1	8�/pl�%�܈�x�%P�!�릨�z��1����o�}&���gib��d�+T��F�3Ә�%ɔ��]B=��G�)��5�i%�x�K5&a�kk�� ?m�b��/��`���`œ��˩���;Z���N}��@áR�YMy�v�c47�Ғ�;9�@D�*>ϧ����;O*Y-�hd�L[�����%
ډ�_l�ӹ��v���3����帰z��8�����dx��1P9���]��M��Y�_��Gg:���y��P�oe���Z�0�(5(c��NO�6oa�FB�>X*+}u��~Z�u���yr�R^b��F���I3A������L���l�t*C��cE�]0r���Wp��RC���w}y.����T'x�ۓ� �bG=�	�NX�iA`����7@��]���}�5�x��ɵ�uDkt5e/��S�^�pd\Ǣ���]i��J�K9�����w��.ʧȽ�)�0$���J-�*�P.`����*�C��{�qU��b�����f�s�'�n���Ç�4��_4�zq��6�Pa�`���dO�����s���7���ɭZ�3��v���Ze�MZJ7\�@j&�%�07�@⎏ۇM�{?�W����	M���
����p�	��&�&@<Uװ>��ȸ���{��>ǘN����O*\r��{w�؈0��m�h���?��8Y_~�CZ1��/���!�M�}����aL3n�2�?��Tҙ|`s�Vl�X�BL���n�Ɓ�q�fXDΤ"hz)�S*�G]Y�햂yP]k���& V��IB<4�����,d&r�K�fVX��jS�����U ���f����H'���ޅ�O4��F���*��j�%H��ʏ9���i8�G=�OR�˘
��+���ً��':ޣ���XB<����B�� -fTM��Y����3NO>�RN�~��ꠒd�����b�UR>.�_�SN�(�sty�߱�\v�3�B�ۿ�a���T��:[�d?�;;�
_� <ͳu˰=Z��@پzL�o`?YڇC��x�YQarҸ
9v� P_�9V*��Vy3DMgzu�YҴ�{K��9k�anDrC
��.�6e� �G�����Ģ��[���_hfb����:P�i:J�%�;�G?�`B���@J؅�!in�n{��h�-��h=���?8T8���T�s:c��_"]Pv�rVE���G����ۄ���#�)�z1?a�Ҩ��Fi�
V�&��$���L�:�l�gFu�9�ɩH�z\Qb���G��dx���"#�j@�5F{�a0�'9|�t\���r��|��Rٓ�"̝�6̼]���z���WO���Ls�����C�M�(�J���>���Ug�I���G�aɸ���:�����v��uJ
ê��'����0N�[�w_�w������gy��x��R���7�+aB��9�^H+K=�4G]�7<z�b:~�ZN�zc#`K�@e��ֽ�-;bD{U=�8~�����8P��]���ݳ	�#�����?[�f�}.H$Z�.�����ٖ|t&=�I��@��if/�3 �Yng~�\���ǈ��ŷ�;���gS���H��;���0�?W��	��c����F�%�7�U"��֭������9E,XKL��u���RZyNΔB1����
�,�E�}�T���/�n
��Q����k��{)U��5�����X��?��w0���#-����K���\��Ei/�f�y�;���p8i]��s�����:T�YF����9,X tn}��u�~��Wc��k�r�E�{|+�1#������`S`H�kqd<�37�Tjy ���{�U.#b�}�q'���g�b�h�LT��RuT"a{S�A&W����&�%m�ȧ��uBЧ~�瘍/�c6�{�	��])ѷ��B�bC.Y�^W�i%�8������e�KV�_B�����L�1���e�ik�#,(^YP&�~C�|�,h�&�Z� �wF�>4�(Mh��6Gex����h�G����k�����-u i+���ù���0�vt���������a�#�����4ۂ'#�`Q�`��#�����2���R��iB_����v�+[qK"�t9�G��n�e�Z%�x>�#4�r����@}�"��i�C�� 8�����/�ӺÛ�`�~<+���IЕ��X���'�r�0�������O��m�v�t�6�'���a���=Z�9x>z�*�*c�����U^��u�8�Aҩ1
�r_(e�� 5�dE���׏�ѩ����ec����������˱ԿH_֦KU�I�O� 7t�{��#;K�B��|�+v�� GU��R|^�ՙC�+�����`���%��V4�A�2hEJj,�0�z&ǝdm�ny�z�j.���m]�j��
��`&��#�E!���ߧ�.��a�aJ�hj�Set�!ʹb�h-�C��E�t�)]�n�!n#��SM%���-*�{L[K�F�%MG�s���m� 9�X��wv�3H��]�S���qܥT�Ix�Ǖ�s�gF�G)LFX>_���E��(�~�P�C�1�Z#=��r��d@�Ó��-��,ͅ����ߖ�5#s	��"�;�n6xzOz����*^�?�~�#Ě͠n�
d�hF$��?��/i�������)Ƀ���:�G4���ab��0��?'7�FO�$�E9T6�n̉������z���'-�E�����(�YN�:�&�'T��"{�����ux�bg��
��D�0���:B$�e���X+��4�Z�A�Y��=�/ƻ�ouf+C�#H���������8��:ȟ�%ץ��~�o��<ܓ���mU�M��|�S��z�[֓���,ec��)���53��H�O:�,�C21���T��X�(q�3�xEv�0a�Q�@���
�xX�@�A�m2հ
� ?4�0��w;���i�£���u� ؖ�v{�'�������/���uR5x�@�'1�s��i&:\h�w�����M�yTS�$~���4.?uŁ�T��=�ڻ���eK�]���o/��孀�-�W��IF���/N�K���������v�&B�K
r���BDS��q	�C�lR(�}�����n�K%�Q+ m�oo>Ec�su����.�B	�JH��״�8 �,�^�M:F��O�~��Tr1���	n%ҽ2��t)�"LC]P�Nf۰M�
��^��$R�p���rPҳI�q�'`}E��2��V~�}E���ۭ�DF5����eI~��q����h�_��� �'�]��m���q�I���i{Dk���/��80�HV��󀊾���
�"^�F� ��Z�|l��q�&��-��,�� �h��9Z��tĐ���J�p�"q4�YU�l&�M��I��N��*T��N t�ѻ?3�w�+hM�+"�J+�/��}�)ͮ�5<�\��ǜ��X�a�'��h��(����8<!,5\���
�w)�LZA���i���娄���ʻ��U�,<]�%K���4HkF�_�ȭ�x�>+����c��tfLk[��M����������>G]N�;uč���P	][�}l���c��R��_I��g����N�������E]W�)�4uݓ:0����4�a�&d�O�ۻ�zq�j�b�D�/��@�O���V�L{�D߆QD��9�ʆ0Ԅ���.���f��N�4�T��b�⭎�aq���t�e��4���A��|���� A�"+�
l"��n����H�W�6F�"� ��6c��-1)-�>�K��M8�����$�}E2]*��	d�XK>
K�
|��ZuV:�;qE?	�s���
D�X������A����6��f�xZl��R��\�5�3���mϻ�F'�_�˾��$�iE�x��m�p�CA�ZR.q�{�jL�f{��ag�b>�8��s]�B
���
��_����A�%cޮ��!��{:���)#�	p���׬��0� 		?�!�M�>�&i'v�����+�4:����3H�}����T	�����Z�z&!�v�m�x��Y5_�6N0��`Ewb�AS1 ��D;u��_���^���T�U��NJd���9)���o��vh��_"E�pM_q�Y��*�=�<������V!���3qI�nF�9(e!�:Z�2�n!/�F�V^�t4�n5t�D|Dzw��!)��_�8&�(HƘoMB�@��ޚ *;W���l1M�Y��58���I�����,@�� v�`@����pA�:�QI���׻0D��q�	�Sy4���ܦ9w@k���d�T	�e���qv�����B`����w����<�c�7��i	z�Lk~	�1VV��)������b�W���Ov]��e�.3�U�)�SM�����UWx�:lS�fH�v��@Cjɢ�m���*���-:�mWL��:܉��Q���]�(��{�4�ORO�$)�ܞ���'�/�c�>����N����'�HY=fG�����~9����+	�K�Ӑm,�H�{MMh|hQc=�k6��!�D��8��@KN����Уe�:�F<�p�����H�k��=� 5t�	5�	����O��5~\&�L������q71Pb����j�>��S�T@]������1�*k;�C��u�د�A��1țM³`��
A��&���F�[^il����7?dzg8Q{|��X+B�{���W4 ����*#�y�e�}4�vW��� ܲA�5�V����ڱ�҂>MJa���PO}�gGl,�no�(�Ґs��8�O�{�@��JPh�J9;u�� ~	8L��s��{9oYQ�J��:v��\��.Q�[z��^�o;_Ի�������`���=��f�tb,���/���G8L�B�MX"m���kT�]�0��U�5���PL�,[��t�bn�z�0�b�ҭ�j����j��j%����z��;;K���]&O����3���u��AX0�`���?��2{���z0@{��AY�����t�o�^gu��L;i�Bd��#T�^�@+�jlyw_�\8㙣�`�/��B3ǆ�>�'~��F~#z��	�����'�ɱ���m���බakN*m�W�O,B���{Ҍ1���Cn/�كG1giIF#�<{��r� ̊�Z�f�+��_��ܯ���xYz�4�D����"\?�+�Z�����^���pM��w�v�*��Z�a�W�F9F:I�0L���{�m����E�`�WV`|`������1�v��0���3��p��E� �t[Xs�WJ����5��=(0�l8����*�7�B@x�88<�����Ez��E����;�j���$ɕ�����b�Vꐎ3V��gjj[���I|,�tΏ�T��Ϧ�AZ(���2SS�Í��8���x:eᲢ�`-!3��%ۏuE?�����@X��O�L�Y���n�Z=��k�z�W"�%<��������y �`0����ؘ"7j�����2ͽ����􇳩����}��2g܁A�6�!�*n7z*�
����&-f�I/��wh�(z/<�,����H�0䲵�����z�a�R�d����]0���GS�"Y:����-.�a�͍�:�]��y����YX�O�Zz,)~yj&���!�
�&�5��Hw���i^�x��?��v��e:�s��S&�k�����5��Ҽ��1�)����ғ�$D
t~�������2�rXR�dP¼�F�>K���Z�y�_��n6��X�	 ��\ගC��BŹJ����r}�P�E�5��jS4tXZ���H�x�.t��o��&�b�$X�qw�A%G�Mf���[���#m�Hl����n�#>�]i� �*w�;|�#k��i`����.����&l.�_Bs�Õ�a�P�ˋ�`�й���=8���a���k�"�����{�� l��F �����F}�2�]]�O�vw)H(�>�?
ȿ��P,*l��,t �e9*ԟ!=�_# >{I֪�yٱ�ZI"@�0�S���A��cy�N�L$yZ�(N�ۏd�����C���Io��'��;ʕ�/g�O�d1�^�[��<��Q�E��׊�4[�?�(\5f�Fͱ�=�o�ö����xv���Ş��+����);�L`?S�� p�K���
�F����������Ve�����qyԳ踲�Z���Q�(�,�O��z�)	v�o$�W���M~����'���f8
�\"�V�1�0��#�D׻F/�9�c7�
��n���M�y��RZ�-�v�MT�F�q]�cnl��Bq^j�v>QL���ټey�iR9^�o��@i���9�fV��'��G��B���	���u�[�*Z��c��~�\��#M�AO��wz)��3RryG��������s��1�� �F^�|!l���t(pN���I�`��T8���f&���G!E3I2bc�ۆÏ�|��/ҌZ�jn�&wg��]� ��>��>+T�KB���Ĵp݊T֚�*�ʙ]�cu�ŲW�d$}W�[�����BY�=��k��(pd%ne�th�PA��P����!ϐ��vr�b�;�TBnn��\��ƚc���
�"���:��
�Z;-yIviW��
��I�8�*�c��ڏٚ3ay����2�e�G�-�Q�U%�^kA��������ɮi��$��(ȝrޖ�H�'����K��B�*�E���
�kP�r�7	�	��\t�� =�a/t�p0V;��}t�ô�2���7B������R�7��o�_j�զ��Z��KH���DF��|���\?��sqSs1�)(�~��~�����K>R�#�X��iI�ݘ����B�����4���+�9�9�D����~�k3	�������y#�-�����L���� J�s�a�t�P�y�Q�h�����"KdAXILEfO��]�� fvje�$�%칉q��5�&�B�+��
3�~�.=b�+�`es�A� ����HZ0˚XG<��`��k ��!��I ��
Bp��(j�#=��^xƚJTaf�V+�����j�`�E�_�⚠̚y�E��=��wY�b��A(�NK,�ͪ�$�4���`~ʕ�A3��<�x4����U��[�~;��m(��M���mqۢm2"��/��](V�% ���z�
4g48��UvZ=�_.{���2*l�%p��M��ɓނM������}�K�X��;x�YQz#1���:{�U%�|>M�B����Oe׬oS��!:N�h����2k�ԋ��5��r�����%7#Z�L�xzne_��>��G{\�$��J��و8�2G�L���	���ڧqi���bpۈ�挡��3�8p&��c��V����.Gq�N�Yg�")���M�.j�?3��Uр_3*"�
�#6x���M�(���(X��C1�B"�>�9���Q�aI�����F���{r���T&���n���H6��XL���2V�r��������mOj �o�u�ag���)����]�d ��ax��C�j�z��6Z��ʋ��76���k�ύ��I�XT�	�D%�F��X�ɂM:�o͈�)sT\�����eU����W~�����$)5����:�r�@YQ3go���<�X�� �w"�5��*�E����%Q��\?�jD�K�VO@|�m�Q�1lP����ClkO4�f�ʅ��Vm�/m�E-�"�/��I�q`����6��uXK.s�=��6�%�`���;���eZ�w�2��z��wX_;\�N"Ɡ�r�d�s̚�#�{�����?k�a�<�ۑ!F܎+���R���+3�7��I���A��xW�K���o�+{}> �@ﹰ�$3��v��W�	�����pV#�|;z��k�����ݖ���xP�@��V,�l�}fR@4�	x�l��,���u��;�,�=�i�}4^�b��x����x��f�7�y�}����*����^W��oO�f�&�����m#{v�8�icr �cc�C�������h3:�3r׉�|N��� ��'�p�}a�.�WVu(ɧ|H�L�\0�'�3wh��;n�Mr���{�!�[��%�v���K�6��pq��u���M�v{�*)�棆��u"�h��t�'U��a��P��	O�x"2O�A.o�9E-��1�:% t;C��)˨��/.�5�.�R�5{�Ψ����7�c5{�t���9��z�m3v�ـ�m("
 ���K�V�.h
n���&>�{WOs�Ív �8��9��^�%&�IK��ٰt ����Mx��4�����`�������h��z�Y(��jswJ�a��U��d���G�����w�m��ł���v�
�-����������a��mL�KW�AQ*A��@܎�D.+�]3��CL	�� �$���!�@jƜ2p�ؤ�Бl��.�ѧ�o7�<�p�)�h��BX�_E��Tl���[�i���L��qGZ����kի�д�'�T�\p��м���ĈM+ԡ�I�Q��|&^2�Hl��]^ ���<<u8)��Xe��AYO���oZ��}p5��}�Yaյ��C"/!ڀ�ԫ+�]�P��K�$4$� �+���D���U��H��z�^t���ba���mMb�*8,�Ѡ��]*��'����n#9���cyE�w9y&�iU^n,}x7�b
�-����p�d��f�h�ҿ��r�޹Q��H
��|B�k�"�U��=r��C��2�AR��s9/_%e���.�zc?����ڀ� �c���5�ڝ����4�yK3Ұ��w��b��$���2�O�F�I��ݼ��G<�	(�>_�m��7�Ҫf:k.�3����H�̮�-K�lq��ˆ���zw5��������fnZ���.�$����5B��������M��G;��vt���xi1�p4R�L*Ī8Mz�妺T}FCt۾~�j�+j}�9P��ؠ�9u����)�Т�mE���n���(	G'��n��y�d\#�9 6l���<,Δ�/��������V�O�"�~r�#>���66T)��L^͖�ċO��e<1j��vX����9�������!q��3�U���U̴�:�$[�W�A��^w�
��.����xC�����L��RP|l��6�X9�������|=n��i]\�a��d������c�מKQ�S0GEKh��LNT$NA�	��;�4�UWo����3Gk��wV���,?��+tҒ���3���t�:5��N�a|0�)�AM�/0������>e�H���mk�?>�S�	퀒˰���U��-,�,u�*�5;4���q�yK5��״�m, ���0�������B3f�"ܸ��_|���J�UXZo%f�+��-�V�F~����~.!�S�m���%3?FP���&��GNb���ε>��]�BZuK�ʷ�pߴ���Ju�;@�[+C���P�Z�O泴�j}:�i���N�*�������78iF���[�KK�W���˅��ۻ �a%\Z�J�._I�T���Q3.���xM ޒȑ�Q�Y���64���@|^̋��c��&����[qG4ش�hbW��V��-��u��q�f���1 � �	��vZ�z�Q�\�¡��6G�j}����+J���4c��8�����Az���ڻq*�,�:���R>��~�K��/-��c?�� TX��(����8��1mVg�c�0^���J��~��A�P�	����na8h�$CLh��V���_�Z`T�nf9a褉l⒕���Ϗc�w�R�ơ��PJ����x�����6sm��lP���N5V�4��,V���ɱ]#�-(&s�F��:b|��e���������gm54	��o
�#�Q��$�L��d!~�AT]T��g���W.ڿ�A���p��ʮiN�ouZ�e�H6�`�$�@f2�~`P���
����Uw:j*i%kAY��"Н��nH)8C�T������5�Q���l!�}�n��d'%�ka@c/����J8:��p��#��I��X�8�枦��ÄM��M]Ї�(�$�/'t?����mв�!��E=8-��؎��CDd�~����$םyl�
Df���Zx�Jfq��ͨ?��7��.ޯ�4~�\��%�
e���{7m�z��m[-���5m,#�����I��q�o(r�X��u�Yz���'�)�:γ�~:���G^�3�	�f��~�{\qs)�͓��#���l��XO��IR��_�Y��a,�vm�p�w��uϥcq����
���0���˃c�H	�o>���\�k��=[�sk��7U�C	��x\z
F�~#�*Ks�g}p��z��#�)P�O��,��*>�$��~~��}���� 	�X&q����;�o�=��� Z�n ��qv/D��6�H٤��D�[�'�,����Z��*���dP}L
h==���Er⪖���3���r,�s��+<u��3�6�����V�� d����j�v�b��fs�����ᯊ�Ѩ5*CGQn���ؘ�Y�
F�FuZ�ռ���P�L5=�b���gP.�7g�a; �|��a��s�gl�A��י��c�g9Ȃ�΋�v`n�31���	gK��9��VS�J��s%�$�U .[�C/%�g`@�pkxK�e&�'e[i����̓�L�`|9ۘ���x�ϥ\i(� K��W�F���+�r�
5��̵w��W�6�d>����]l���ֳ/=��"��BXE���c�������!��Ec@�V�L���:8j� eO��&�N�mM�O$;��V��t�e� �Y&x`�5"�ȃM��K�:1�R�����t�{�<��ڃ�Հ���F T�̋��J.?��?q���h�h���s��M+�m�������.��ا� p�ҽl������"��g^�o~��\��DI�DE&z��ƖX��2����9OJ��Ʊ�YZ��o�^���gi3~��'b�Y���)������� ����ձa�Jf�c�	˧�c�A�eݸ���b53_�*f�i���c!Gx�m-*a�����J�(�ꈮOjv"g,���yΫ^��O�)O���n�m
ty��޾�@���n!�Y��	�N�zQ̓ �������I~��sJ�:���r��2�L=P�`�I F�`�yn�܈�ι��P�./Wf�-�����)9�g��-��4d�Ƒ`����&)�,�*= �X6$G7�%KPJ�*1NJo�4�}�H�̥"��)�K���#�I��.��M�][����j����߂=�y/�����Q�����=}���f� �{&.W���	[cp��<c�C)���:�5:��g��aɸ���{����"���H�I���m-As�.�u�	�HQfǹ����TeX���t��q<��a�owL]ѷq�'��{:����L��]0�u���7qɉ27}\uc�v����>ӂ�YjVu8�IVxu�?<�Ex����t�d$y��U7��Ѽ�<�Z�Y��W��Ǻ�V�g#�i�Į���'�D�Bk��:ڹ%�Ep�'�G�?����W�?�C���o�K����u��Df�3lD��4 0n��w��Xw������s��|�l�D���uw��j�zʲ񧻇�mJ!�({�]`� [�V��ג��~!� ZR���xF5j�&���zqC�ĚI�� von��������eQ��3&�+���Ս��}���yks[W��8}�"�*XL�I�j�N;��;=A=�cR2�A��l�C�������Xѹ��7��_=+
���R�Iۉ)�E��qI.�ڼ=:O�J�T�U�B�'�\!����-�V���ԧV�Z�K�[�c��Am�9�2�G��=a[By��D�@4hx�b�s�Nk�_�A�{.�/D�r�
C����>�d4��D��]�.��4N6����Rs�ÓKj�ٺ>�HYR��$\�F�K1y`B�q�w�VC絇�i�NT$'��f�v�3EO؇G��)d�y�q�GFvI\Il���
9��Z�VeKUT��ʁډ��y}u��_W+<�;����D��Y̜�s�U�bov���:3QFf3��E�C�(EK�o��Y���~]���
*^Z�K�:VvF����DΎ3-H	 �	��˃ h���t��]!�-h̴�f#☱�_�M��l��Uu�u�;剧3�'���8̡�V@��:��:J�^/��G��;l|���kƢ��I%��]�Ĕ/#JS�z��jw����~Y���\������E�����h��[�K�^=n��~L�H$rW�ĮXq���l^#�f���{t�`�fbV���:��¼��޾���|&8V\i:܋lv���qR�K�fB����\���0�ڈ�mʊ'��7�u���"�Pw/~�v���esfncF�I(4j�+�xA�s��	�G��ʡٹ��N�U�~'x�w/�2]U���ÎR��n�+"�aM@_#�,h+,ʌk^�(��K��~}	�6���<S�ɩ�g-ώf��~X��û6r�7y��e2�)������y��3��V�d0�;�G�êF)����e�L���tJ��&���`"�XI��)x�j9`zDn^Xq{�_����m�/���$Xy�9Rx������`);��jX��wz��������ŧ�M�D
�s���nZȊ�[k���UĆ�= �L��JZ�@��#-�Y�M+�
_3��W�G��D-O�Ƙ�Vk�̄�W�kH��������X5�ҵ�^�E�ڦW���~zE�h�u�%��)@��j,����o�p�찿@�aC�J�$X ,n�gz>�=iKT��V�L�v?�x��D�`��U�\���>ץ�7�#m��/���׳&u��_L���  �{�ż�y� >���ȓh0F�x�k%j}\��[��O���JӥJ8�*��t��cut!��y3���[��S�g�%�5���Zzt��@Ӡ:����Z�1��@�X���2T�_� ���3/F
��+l����Gy3N�&U���9"h]����~��,,��+����)�q�a2��i�v�,�!�G�A �6�ͯ67#߱U�M�ډ.��\�ʱ�?}�-��� ���C��&� �л�q�Hv��+#�Q���s�v��Rt+Yas]���aX��i��,p���HC̹��e��_Z�����c��`� b�k{���%�6NO�@�{i2ue�������=ɉJ�wv�r-��Ⳓ��5(�R� �ȩ��&^-0JK��Y�,�V�����x����P�HR;���W��or�S�c��6X	ro��p�d!}� @�W��HY�^P��	�9��`��$�np�k�=��nRt�H:�p"N�OD���@,[Q�V2�Ԭ�%��I�F��H4����7@q�o���j��˝�H.1�Y#��=V����G���9�:���T3��rJ�@����wC� 9`���~�R���B"��X���M�a�8�.�K־v�{��!`�
�w��q�[SDLp>MS$ې�( ��w�Wd�yz'�>V���<9ڍ*�L �89�^����v�o{��̃��T��*�z���҄Z�,�R -Jf�u˲��B�_
��8
gz�!� ����f ��?��Դݘ,�.�K��P�(�C͌�;7(��-�UPpbo�����"Z�,���F���+0�5Ĥ� �	�]d�I#�W�Y�=����R����ȸ�r�[��]��N_L� ����rՐx�{:����ٴ�d����Tm w�o�^�%<�a��/�	
X�`V�d��� � �~#ͱ?l�Ǌ0�뉦a,���,x��T��S��*V[��߅��7�L���=!����on����h_ O��&�������]&���m��r���o��^ɾ~����ύ�����e ��m�����m��T�>�Vot�p�͋gj^���
��v��u�����UFTb(��xɲQ4�!��ِ�� ݟs3��o�@�	d|��c� y
�E���e0����6��X��>ޔ%��s�oU�ZiZI	""���k�mS|���Yql��7X�9U
�$t$B�/"�Gu��#X�,�)�b*��U�W͎݂[��I���_1Q���M�a����� ���<]?��n�!q$��%�HHA��7p��5�B�C�&X���7h����+;1�&����
��~:�j�����	�7�)+.��Eyw���q��%��lY'�K�ya��۠uɮ�uƘ�q ���OE���u�*X�[�
mUW�8Q�b��ǲ��6�\�s����A��\�����@�;��^��t�e`Ŕ�<U����D�Ɣ�>��qP�؄E�v�v_����o+k��e����/ ���2�����A�j� �7��Z��Ts&^V���w R� 9�ru��h���� Iӵ��%�>T���e��J~B2H�+7V&A|��	qfC�3pޮ��Њ4�PҮ]+�i���k+\�Iㄕ(j�햯-ݮ��շڸ#�N�<�L�ʺ�&tJ){][$�?Lz�L�ﵒ�ҧ��~BB�Z�6�) 趼&��G��x8����\�JN����%�����O��8،��]s��������b����.Q���v�*��k�u�OV4?`�K�C�c�3�h;b�`��s�^Mx I"�Wـt<f�-�B��ַZ�j4`���Yg�@��aI���7�zs���H�*MX�E��B<ˋ_�l�����k|����CI�|,���7٨���b���!ʕ�@��rM�\ZS�4E-~rP�;@N9�Ok��Ek�?Ds�r�7+�fBv�u4zg�g�l�~�@*h�+��a�y,��Q��<"� -:GP�7r�\��
}��c���<����_��pP��D�/�?��Am���A���V0���ϯ�^���Ui$��@�04��]��6`vHT�䜡��*P�T�[�x�dV8���i�FIsD�gp�(�O�@�n�<� ��(�\{̊�;�v`��֛�ﹹH��o��nv���k�c3t*��huP;���Gn��Cc�B����l�O##��k o�O�8�Λr�:袉��ɖ��
:���g b�Vb��)v�ny9�0�N��=@:Nv��Ss��& -W[<���T⨺���9��MuE)S�j��H�;��.����МG�Xղ"w�ߤhPx�H�%�S#����1���)����l��Oh'r|ғ�V�I3��4Kz��la9���/�`4��ۑ��Pbt�]&���щ^����&	B~�0�!o�]��7�u��;jFc���$�}kA��>]Lv��P��ʤv�GZ���u�A��`����������W%��y4"�����y V�X�$��9HВ�H� o�^���1�4�#'�n�]���o�-
.{����.�!L��I3:�k9fL�Ύ�m��$%�^�����?�zt�m2x�.����ud�D�lLdM�xo6�t���.˜���wYI��}��3V%�E�~�����9ű �`�0��\�[#nf�F�ƥ���0әL��[�sy��y*���}�\ˀ�<���b�$56��F���!�i��b-���*f��lꠞ��p���1χ?d��I���U�}�)U�� �_�$<�""��O͆B��w���AQi�(;��:��p\|3���>P� ��i�h���Q:YQ�<�O8�]!�=��f�s����O�"}�p�?9[���������Ϸ�=;?	C���t��t=���DZ ��<--����Q�{�k��e;q����曙hA��8V	���Z/��?���c�ݒ������,�:��7�o�'���^�5�;�rd�u�j��DƆ�eT���>��C������}�lH��{/�/F�"FL��?���*�����hۂ�@F��`�J�;j���E�?����y��>,��cU�8Pr��>�C�hׂ�4�Ѳs��9����xpP�+[�K�\�Մm[���k�G����ܔ�p�KA��>�
n:��so��\n��8�	�hSf�Y31�n(dx��U��������&X�C�d�Y�G��}�b�#_s�7�`�|g�������jؖ��=}#k/��t��3�"VY�Al*� �d1j\�f����u]b��/�����P�$�bT���'FGf�-�6����9�ݒ` MR�`��R+f�����3{y�Ms��ͪ[dPq�ç����x�vZ���ܻ�������
f���>:0!��^%�K�N&*H ��Ņ��x�׃���uP~z(����k8(w\GӮ�5��)�l�5�H�36H�i#ePؔ*	X��3I�>�ۇw�,D%zT��A�?���[��r�|�~b��ŕ�P���k {d�;ѣAoO�U�B@N^X6 -HWI? 0(-���%X�i��Ġt�qj񇙡�}���}b��8F�����&]��Ԥ/lܳ�{�	{J��d�~���c�O�\)����ƾh5����K�׼3Vڶ���[,�6 N�G̮
�(��x��e�X�V��B��(���U���%ȼ�1��I[�O(.�H��;�gy�Y/I��6�ք�	=�:i�&��e���5 ���^�~��u&�ҭ�P�X���*� )C�ZW����q���3���z����#���V�o80��h���k���P
�y>tm��D��s'��H%:C�;�$�,���8c���`�5��XFp;o�*8�⸑?�#�l��jZ(�DW��F�H�``����D�Of����x�G�|Y[7m4o"�A0+ת	Z�Ⱥ��c��~��9B��9�2������8���Pv?�=��L|��+��\��+ �p�]av��'|F2ބ�T�>�L��r"Q��_k��?CF�q�K�M!��9�{N>�����>µ|�	6�Wʧ��f���^�����/nQ�ݸ�4��ڙ|�蟪u�!���e\~�4nN��.���"_V�O�������3aM3��L�AQin����9�T�ۃ\*,1E-�u\+��O����*�e���ChX�P���NC�1(�H���>R���#]$V�(=���>�[�
 �z����`qI�0�јGkX�V�>�+� ޼ÁE爆vE� ��g�;j���L4�#/�����i�����} �!H)Nb�n���%� ������~JXR\��d��_����He��04��XF�n]�؂�g3� �ѓ�JW#d���! ��0�"�up���pFw��	��
/�͞(1�oh�:���w��*8�(兎<��^�v���W�^�k����sV�8�����c 8�����Aң�-]2�?���j�>ϰ���J}�D��U� =���h��i1�);O��J����x�
�Ѡ����r������m����j=>�,��G'uk�Bt]�jM�%4!��g�'`�b~��L �ֺu;7��0�ai�7���$ճ�]���U�V��.�Ei��-&�#?+/��$�`1��^,�����g�uL2�ɱ��=��u��_�/e�����[4����#V��"�X%-�ֈsD�_aOY ���i������{j��Z$�$������U��y&�r:�Zpő���z̿5��L�.����&�N�b )�yY������t��26�ד���CR2E
�du���t�=X)
����{�u^xt�W�3l�Y��8np���-��g��c� �:��� ���[��G������=�4�BiVr�U�0s����҂�5��Nu�Bh�{�-0��e}�ŉ�7��dc���ގ�jN���ǡW>X�s�<�$e�.���H�#����>�jxY�p=UĖ X��,��/�F*�c=Ƨ���f`�.��$J��X:~ٖ�Q��
J>�����ktLQw@������s�W�5��J�h�@w�sk;]_�\Xo_=�4S�-��ڍ%n^��G��L��z��S+~���\m;�~<����j�����Ĩ�`/��G�RX���~2"~|�Ux�u&�_����Y�JF�[= ���[�}�[�x��o�b ~>�y�z����l�K˅�X�< 7��tn��c7��U��Ł%���� ,*'2�zl�������ԤԲ�aFC��ѷ�U6׫Y�mw����(m}�H ���S/.�0Ӆ"���bSb��(��rs��E�j��տ��?�<�M-�u��`�6j�
X�[���]@V�m,��Q±H)���	�uz�8z�oթ+��k/
��ْ�|��{� �����n@�����4@���$���$���◓��T�!	�1M�E�B� AWd��22���)PR<��l{`�����(�.8Q��,���_����%(��r��&�_��X����tF���=�"9~/�ߝK��_�W�U�ܯ
[Sbk"[��1X�S�:��3���}M�7�������f�5��P-eh�� ev:tˇ��p���H�Ȋ~��{��H��M���ɜ�qR��I=DC�ZyQ����5+tz������� RVX!�t	!+l���ፘ�[� �0����{&���O1T��I��/%��߆��ۉ9"�;�^@dbʉql���T�b��؅L	��sP+�3�D�wM�|[�_T?��z@�@TyS��Ӣ0�l�~IX��c�%X�!�t�ʲtI	�[2�Yxb��1���^	ڟ�����`H.���Fm(=���y�IBd��*O�}����o��޵hRz��X�����lB�(����i��n��FB��1�|��F"�x���$
�G��H
o�����z�C�.⠔Jl�O`�ivPo깝 x���:2t��*�{��b�f;'�5]%���ӣ�>1���c�mQ�=���ڬh�Cx�G�	�@?���"K �YF��W/jWW�(�A�+�]�Ibȓ��20<�#-_��ȩ���#��1ly�7_��>L��
��X�����a��Z�x�,{�1]a�f(��:���)+<� ��"1�>�#ʺ
����0"�t���%4ע�(�/��\Wa����gy������k�+�^���(�u�h|� #(Sz���gN">+ci�8���Å"�A'c�pv�C���<Λ-
���9�V
�D��<��1:υ���gR;c����+���	��N|�U��`}FQ�@wg�zI���m�$W�[��(�pn��LG_#����Ʀ�u!`>��).�I�ρX�?]28_;��U8Uo�twZy"�mG��$H�5n�;b��'��X�V��u8Ë�ସ����$��	&�^(������/;�y�������ڀ{�� ���b�̦�VXE�Mj}���\��:q�����U.k-~�K]���_ȃ	�C���t���>����ٚ&}���3������v��]`FM60��8��Tt��n3��6�[Kz�?���)�|�0A�#�����.v9Y��<�ɧ��u`����nW�1��Sw�:�Y��տ~�����y�x�z��!����D��Ft]�d�2�i���9Q�nSz�Y�̄��4���
��&呜�&�M~R�_ࠃ�����4C!k�co�I�E;����|���8r#�9V�6���X��X��d��$ʎol�^� 'AՉa]����˼�|������x�0-����$�^�ٝ��n�|��zEh�J�.(�����H�5���?Mc7>�Æ�2t���!���B�՝�ϡ����֘y�YU!VK*�P�lg�Ռ�|٢�p��c����T�#Jc9a�|��eը��ƮXy]�i0q?j�*���l�TUE��ɒ�#݇n��	
�{ǏmH��%7�O�#�sL/���έ�=�;q�Ab"��x.�
E���l�s�x��nRS"�s�s�1UQ=���sYsE�S��D�i^w�濴�b0��V�v�4Y�pZ(����)�E�R%���9cOǴ6]�,��+=,8i����u���cΘ���� �7�e�ӑ�5c�e���F��`���hH�!��)2������,��\|�cab��X*t��(�$Z��a�=��z��l}����zUV<��#���[�c3jiN��.��O�x�"�u�q��Z���a2�i+ңrJE��,�	$QG��0cLL�7��@��˓{.�9������N&��n+YV1��.T�S�W��?�;!�7�X�=���cf0Z,Bߚ�O�ʠMO5DbR[k���*��
L(q�a�B�m��xo)��h���|#����,;ۡ�K��"ɑ�~��X����.��mL=跬c�M������h�=&z"�)�H>'�P���B�޶P^[�T���@�hw�*Q!K������[�	��!����������-p���`O�R����.Xvy]�>Z��{��n�C�B��f%������#�S��m���C�h�ߙBMS�;l�u"�oz	�~؅K���?58�R����y�f��*��z--�̎�3&��E�Ջ%����˾���6[�����VH�,���'���Xpل�{	q�iâT��ߏu��y:(����/s�(@#5X>5�@��%�1��&�^��g�6[J�u�n�d��%�i7��#VTZ2�_�/8���r���S�/��lq��E���� H�L[��	��ò�k���3�(;fU��8�âٲsqUd�0sl�9���_f���Ȫ�i��I�b��/���!4w�߶ۙ|Hb��5~Sy�4��<�۲�f�Ɩ�:����ڬ���8k\CO�x�C	 8+T��J�㍞�i}p�+dlx�&$'�ݭ4m�=r���/�T=n�RSM��!�k�8��0z�ysC@N�#0�����q���+]�A�����A�;#2̙Iu���pY#GnV�1���pJ�7�h�h-Ot�$f̯�"�s/�����J�B6Mc�?(/8T	�1uT�௖�g(�仙�O�1�^��x�:=�yN��֫[�i��wu�h*&N.��������%�'z0W�I[?���|���6�:�֦t�=�ۃ�vXVhQ��H_���\5�G����2����o��i�!YN���|��"9*w�����1b�(���棧`�P����UV���Y���g�I�����XֳN�s�d�崵��s��y��"�3N�C��U�=��GV���*n��s��c���*�tw���9����U�Wl�p��J y�)s/��D�v�����)�bW�C���$���A�SZU�������z���f?ov�u���m�(��7,��SpP�x�Q�E*?�D̗�ȑ�@H�u)$!sPL��N,a9��4�C@���\w��ګ
M&�j��tu�A�,x��](ӉH}l�k���v���Z|$%�oԞ0#�9jyBߩ^\���m*y�n`N��	���o��r�5��N⸿��B����ߜ	���cX�!�nJ�9�IҐLv��5��ݾG
\�M�_�ւ�T?/<M�zB�y�L)$�a��*z���t�j�[��������� �o	! ��	��0��3�7r�tL<�/��ԕ����-����3���L_�f�Bpຝ��s_)���ر����h�[yE�Q�N$�Ǥ>��4����e��z��x����=��1��dj;t��4��v�&���w�v�XWj�#u,p��Չ�*X�Z��Ϟ֫�}95Fk�8fWؙ�p�%o}�R(6�=�&���S�.�)���z\%�ƾκ�_W����L͇`9����,���֒��I;,��kJGqd6�C��sǋ�� ��e`�y�D_!�����b��`'���kmGN���7H}.�7�Q�5I�S*;og-�T3GƖ�E`?�56���Y��7��:��.:���J�sٰ�."�{�:�`x|���(����J��i�����PH��C� }�HxB�R���sj���Q��dF�N���c�O�$k��Q�˄J�Rɷ�A`���d!0M�3�2�`.%����^��Y�l��"�(�� <��b��P1I���y���%F[�Q�ǡn��i�NAe�c��QcG��W����ïr�Ѧ���nC��!�)�[�ڦ����q�)�}"w�7#bm�RO�Jxl"�x[��U5����q��c���٨r������ڒ$���
=Z%@mͬ��Yt�BV2��gm/��r}ť��wI��݂z;�JDS��*� \����,�H5�$�v���9
��U-ID#���h�Q��gn6�߽K�jԱyV��3=� Y�6"�ީ�T�wг��+i�N���ۘua�@�y�.J�j�%uyI1d�w��g�-n��JI"���Z��W��0��
)�QʢQ�<�;�t~���y �0� �M��Q�}k��*��y��1�O2Y��K;G��@6��+Ԝ��-v���B�p��H ~o�[y�w�!���@+.�`�fL����!��B��W&�?�x{�go��+�-ki��l�&O�ɇ���^Pv���m�p��AiB��p�����8����5���Th�<�k�`�ʴz׵��d	H�R�KA#,G9p��Td�F �fK �!�1���!h��XM�E�o�p��J��o���_��ǺeFK���6ݿ�hk	x?/�M�G+�W���"���,}P+��@���CG0���J�'�a�lK ��J�OC/2�řV������vC	�F�z���T���=�X�X�(�Sp���,�A��G�b�&�ihG*�� �V���U=�Z1�E�Be����O�^�=�����)r���o����{�`�7Ë������yVGe`�k�k��TflR�t�{|�U\��!�t6��(˪��j�~���W��;9Ikz�@Ș�b7����7�S�������e������a��*��4�,���z��2�5O���V��M���]�V��A>�S��N��啡bګ����ȅ`���Ӝεp�+�Z�|�<\�n��� 8[�<�z����'bU ~a=�I�kUE���WI�40"��9� ߌ�u�{��&��L�\\֤ⱼ�(A2F�P*��}%X�%��2��>��8|�Dl�예*H�63	U�ѽ*4{ُ?hH`�ۋz;��unX��e
B"�mk�8����p�pP;���n/$��Joc*�����e�C����&�u��	r�����!N���Z���9���DW ;M�9d����g劊b,��Z�
�qش�_�q��oC�)
j����F�>Բ�=\�Xrdg$�kq��4u���7y�L^b͝��HZ =�Yƃq]I��0�x�g���/�إ�?oC�%������%�՞��{4zP�Ƀ ڬ�U�\�z���덉Vq@.hj	�P͛X�5�6���h�ڇ^g�	��U��鵕E��z,���L�*K܄T�PS=dr��m�VՁ���ڳSPO�mH��JO��Oͼ3�S����$�z{4�T(@Ô:�->�DIH1(�_�{�%�;mNf����{�q���M�3��X%,���z:FnI�1�/��Ɇߡ��Z~�$]���ru�c�ҥ�T��m��tV�a��mjM${\��kw7���C�%�dD��͡���s���jl;� �@���%�)Fs��Y5��&& ����k(Gn�x��p7l����&�|�^�g�j+ `��`�z�L�ď�?����7@�0�4߷�d�\KxE�.�14]��MF3Wk`�T�Xܔ�|�Ք�����x��O_�V����P�$�L���5�O�3��Â��)��u�u�wy01;�7n|�d��5�_H�[ĥ@e����腍����q�[�A ��)��g�1�\��O@�Z��r���Z�
�-f�xQq��mjy��r����P�̑u����NQ?�~�=i�Pϒ�s�{G~�/�,� 7a$	��l�/�g����B��ְ�QY���w6Ǎ�rE^\l��jI:�Ł�_�w�����>�%
��8?��̿��8�t�Z,��t�h�9���Y�y����lo��Wފ!�sʦŮ^LT%O�RH4?�z�Ϩ�/�x�XШ�9"�}-�=�յR,G�@+�g$��M"��#Y���䦻���KBEg����ZO��W[F�}A	�U��KY)���]��o]�].^bT�qcB������5������>0v�e�~Z�4�.t��yӡ��e(�x�T�/D�2/뢢>�W���E.�VoOA�4)�@[RҲۛϷ/H���O:�S:�>���^�&3��:�30�y�Ty��e���ܠ���d{��0G��t-u��:���3�b���@��h�1��Ȫk�� ݺ�E�M�_�H?�ZJ*9C�q;�z��5]zB�V���}�@�}ÿ��A@�]ܜ�n�Z9$h+�d~�B�\�Ɔ��n�� 1eݨV��w��X���_ !�O�S��c�}������5%5��	g�#�B�����b zH��2��1��%��`��w�2����ڋc�O��%0|��n�[��mO&�/�k��y;��b�-QhL�F1��۔%~`L�l��
�̰�*�8��/��qPF��\̥�b6����O�z������8��Q �?����h.��ʤ%M�^�ۋ�bGn��F3�Z�s��,z�1~H��c,��L$��s���^,#zѮ����瑁W�B��aV�Df��tȱ;Kx}�i��V3��P����{H:��%�x��BF(���b�v$�����h��^hy'���X�$�!d4���œ�F��7{���q(����z�+��ӟ�T_�U�{�C������s�c-d��<~�%�l���,���}�=�t������d!�^E_<h�'d5h�-���4]:+ݢc4a:h�\T¬_�u��|��Z;�0��/��d��0.n_Dv)KIyw�W�)�$��\����[YY�f����>,64aZ�z2�M�B�:�北��@]��v���18��+y�B�eP���ZHh[�0m�GfgH~��F�R<u+�m�d"�/��9ti���W��Z����c��b)1f:g�$ۜXb�|�!�;A�]�D�n�	@(\�$�g���
����A�/�5��w��^7�
�v�%>���^gS$/���E��T�x
Y��ᔅp4�����D����򲖟������T`<췉پh�m�>���+N�M��̻���DBU"� HC>ޒ��֊Ԛ7��bM���؞U��B?�}�~��s~��r ��l�X���z�`D��0����ߕЈ�k�g�l@
!���������K�n�#�}&��'�]�\����W?+VX�!;���~��
�������ļZٹ�G$�D0�xm��ǼP��/'����J:O��h�k�������*�;xuwL�f0�c��5se�����U�s\�r��7R<4»Q5S3C��(��6�H�V�ag���͊�`�6���N�OM�n�~=E���֣��rO�ջu��6�d.�aP����bң�R=���Yy\��3�|���<n�� |��;��oE����'�����ߍ��O��fc��gW�:�Uyj�~.7E}uv��>����k�G��5�B!ot�Q^�4i!���V%%^�[��z��ṈU�.��;�7�"�ޢ�c���u�Pq���"u^䃘qθb�l1�wΠ@��ɜxP/���>>�٪H��Kֶϊɕ�2��)	<�I�B����Di����k�e����C�?T����WY�{l��
�i
:q�m��_�=���Ƞ���Ƚ�X����y/�ܥ�ߡ}TxD���k��xm%4�^6l�9Rٴ�'R�������fT�J�]��\Cֱ�E�f�	E/c�->P�U�д�'eׇ�A�@6�=���\���W�(��v?�.E2#��=םJ����ø���M?��(����d���?Y]���+lU3I��j�p�UW�:�>(�G�5{�IM���l1�[���ldU����.��L��S�gdur#x�Z0t� �	��)Vr�K2�	$#��Q��7���¤=�����F�v��6iF�&��F��=�t�ᣂ$屁����[�E� �p�a�����f��[�z������d�̭����g��'6�\��G��nV(?� �P���q��A�$U=+{�e��2��;Ҿ����N[��-މ���'�Ʋ��MF��6��1b�����}X��V��%��^��+Fw�nr��i�淁d���93�n���8`;o���H���%�����0zbq�<V���~3��$�c��������"9fwSIo�p�؃��������x9�M��J<�HD[]N�8:�PC#Os��r�yS@�s�+{rB'$G��(��h)���2������6���V�Wh)��WH�� zߴ_��՞B�(I��z���At�ȉ�1*�-n-v��g������3JG��qb����$�������px ��&JiW��37��1�e�ٻ�7���}����.xq|�؆�.��mˋV���Kx�a��# XP���r7NA-�K�Cϫ��~=(�̠<��3�k`�7��ALzv�p/9hK��O'2��R�I��m��{�����S,-���؀��ϵ���s�A�e�����!R��qevN��d�2v�@>bX��%n�o�cw�G_�҅Z��ɬ�q�vU� ��]@����j���TeycV�~q�a.�G^�|,���(�{��qf���=&@S�I�����v������Q=���ެMq�"M*.W���~�o�`��3H�PT��a)y��ޗ�H�������w�-�m\����8UZ �:�nЯb�Y�O���e
o��D:8u��8����Q����:,�IJr��e�'觅�#���s'%'��n�lḾ���L?�L�V�2�*�p���W���l��кi&�}��{KP����Pä��1��R6�=�G�:b��n��Zr,�FԪ��4+������T���*^�(`mu2����f���`#a�꽨�B�Ax�N��S��	uM�S_n[g��w��_�;O�r�X������V�u��3��ܵ�
��bw{�,7�Ҵ����g}��&�j��s�h��;��/���J��9JcE��u>e�u���~0  �j�*���<��<�P K�| �f�k2xȘ����y�O�<��)�;��6�p�!eu�[x�o
��ˡ
��mfӕ}�t*&��K2'Np�^w23f�wbZ7*)�ŉf�s3�g�	�!:�����S�ǋ,�;exwZN��2��eJ4{%�pk+C %o%��C��ievj/O7WdK�l§x���[�'�5?��ǢOq���+���+o(���3Iu�g���R0��<��������p1_��w�j�D�%ؖ_��~%kV��,���A��X�?CQ3m�����Z�"��Z,��F�vWDLu�`�~���Y��IO��d�����o_b����m����?�IVv���B��A^���x����p �O�M������<ce�ݩR�F��c��.�����������񑩓?�G^p��2	:&ܵ5�VrO���a�xAmS �dǥ����},�P|�<�奭=�Gj�:Z�!	RG?.Rĉ�4`�p����萢n\ߏ�ǋ򖰗K 2��c]��]_�L (��5��[�?�C��;f3�M)�(�E�ҍ��Rf�`�V�&m���[cz��=���֬����[�A��������SAg�e������C=�5�< ��)F��$LL��`,���c�T)_e���i�8� �n����U�;�<���A$�ٵ�Tl�:&���'�@G^�
CzIݞ,�N�=�֘�
� ��_����k[�lk��
�?{��	)�o�q0U�j��xx��� �g.l��Q�.��t�����IƧ�ْ>H�G��,J{d^l��������w����Be��@f�ᠬ��SF9�O�.���Lez�o�dH�-��W]�M]�).Fs��g�2�!�FJ�Hk?v���9�g�#�s��΋�c��KS��s/8�*ȅ�[��V7Z�ay	�6��0��M�6$���cWa��o/��)�Xg"-MP���&L8��[^0�ɤQ`?I��'I�F�h���&������� ��������x�`�}Qx��d���N�7{I�V����y����ǲ���4���	j�"�/͸����Y�`���7<np.	ڛ�;ɚDϦ�#��E��kD���&��a�ͬ�N������)Ѩ���(]΄��&ے��3����4��V����N^�����m	$1�靲u�_6	<�e���y�
��_Ƿ���p͹���֔Me��^BA	�9�{�Ԅ�`��u�T���a��*}`��1�`�W�q�(k�	Am�t(�Խ�����%Qd���/-�Bi�j�d��(����yõ�Y�)p�E��,&��x��c�ج�Z�Z�����2�
�&�j�'q�5H6�%(�]�9BnV�?`�k�l�%��RY�w�w��F���i�fY	YD.<#��$��5�ql�PH�W�Vg\B�A��TX�'�����D@G�t̕*R��	Vj�.G�Mxq$d�U�Z�h                                                                                                                                                                                                                                                                                                                                                                                                                                           @p{��q�T���S�w�M]�y{�F�m92�bF`�PL&tp{њ����am4�̨�lA�=�My.�u�0�B��t&��z�ː{9�a����V,� �h��A�m_�p4Lk���}B��mGB�!=Az�8|$�v@���x�����M"��.]��ڃ�U\�$�    &В9
���    s}e/��4����;p6s*d�����3ͮQ    5zDO�Y�|J�    W���'�\� �������409�:�)�:7p�`ͅ�G��FS=���ӀD�ľ4�A�o+ƣ1�����J�����&x '_�y=T��W�.:.��3��&� ژ���\���p������Y3��)�
	ڻ��'�o�G�u�;�ޥ�O�eہ���(��0+�q��H�*�������܂+*H[���u����{��6��g������!��KPy�Νp+L'�k�CXY�ʎ�5�_�qY>T���ڡQ|����g��c-_��'�ˬ���Fzj��u��OW���1����5�K�X7��� l)+K���|<iɂ�E'��dE���|&�H-5��3j��cE<cJ-3}���_�d�j�����d�n",��9UjA��"*�"t.�
Z�H6    ��֪��])����uS�� 9��lcI��dӃ�"��&.o��    U*w�3�l�qJa��A��k$C�~�P'�3uw�evO�'�Y�'d�?<�%����bj2`?�	�m}b�3�mjx�۸��.����ݿ�jt7�r���    m�7���1�@b��!yґ0>�!�`:    ǲ<�O{    ��a˷#��    @3�*    �ʹքC���x�������+�/+����O��t���pTy�p��N�FL0kh�=�2~"a�7�Ǖ�c�+REĮ(����7a��=r�������s1w:l��ۉ�+��J��.�#���0-�˶�ف��	E���O�"0�]�-�qAI&yN��&.34 9J������z��>0���(S��j�4���O��*    mˉ ����R.�Z8    BrCۭ��"mޯ�e�t��cZkBg"߮������96x���c>�^(�n,v�?_.�
�r    ڹ�p���~�`�ޜ���Z��`�\�ԡ�3�&v�p��ic#��O�$a    ����jW�    � � @ �       P?@           (@j�t��?�( p5 �6 �7 ����7: =:     ����    �M  ` �` �d ph 0k ����    k  n `n     ����    _s     ����    Ku pw �y 0w P� �� �� �� ��     ����    � p� � @� `�   �� deflate 1.1.4 Copyright 1995-2002 Jean-loup Gailly             ��     ��     ��       ��     ��       ��   � � ��    �  ��   �  ��    ��                    	      
                                                                                                                                                                                                 	   	   
   
                                                                                               	
   �  L  �  ,  �  l  �    �  \  �  <  �  |  �    �  B  �  "  �  b  �    �  R  �  2  �  r  �  
  �  J  �  *  �  j  �    �  Z  �  :  �  z  �    �  F  �  &  �  f  �    �  V  �  6  �  v  �    �  N  �  .  �  n  �    �  ^  �  >  �  ~  �    �  A  �  !  �  a  �    �  Q  �  1  �  q  �  	  �  I  �  )  �  i  �    �  Y  �  9  �  y  �    �  E  �  %  �  e  �    �  U  �  5  �  u  �    �  M  �  -  �  m  �    �  ]  �  =  �  }  �   	 	 � 	 �	 S 	 S	 � 	 �	 3 	 3	 � 	 �	 s 	 s	 � 	 �	  	 	 � 	 �	 K 	 K	 � 	 �	 + 	 +	 � 	 �	 k 	 k	 � 	 �	  	 	 � 	 �	 [ 	 [	 � 	 �	 ; 	 ;	 � 	 �	 { 	 {	 � 	 �	  	 	 � 	 �	 G 	 G	 � 	 �	 ' 	 '	 � 	 �	 g 	 g	 � 	 �	  	 	 � 	 �	 W 	 W	 � 	 �	 7 	 7	 � 	 �	 w 	 w	 � 	 �	  	 	 � 	 �	 O 	 O	 � 	 �	 / 	 /	 � 	 �	 o 	 o	 � 	 �	  	 	 � 	 �	 _ 	 _	 � 	 �	 ? 	 ?	 � 	 �	  	 	 � 	 �	    @     `    P  0  p    H  (  h    X  8  x    D  $  d    T  4  t    �  C  �  #  �  c  �                       
                	                         								















   		

                            
                         (   0   8   @   P   `   p   �   �   �   �                                          0   @   `   �   �      �                               0   @   `   inflate 1.1.4 Copyright 1995-2002 Mark Adler                     	   
                           #   +   3   ;   C   S   c   s   �   �   �   �                                                                                                             p   p                     	            !   1   A   a   �   �     �                     0  @  `                                                                  	   	   
   
                     (3�    Pz        ����        �2               3            Pz3     �   `3                    ����� �   �3                    ����  �   �3                    ����  �   �3                    ����@    N   \ �   4                    �����    �   �   �   (`    ����                  8`    ����                  P404                p4 �   �4   �4            ����    ����                  �4                �$  �   5                    �����    � �   85                    �����    � �   h5                    ���� �   �5                    ����0 �   �5                    ����P �   �5   �5            ����    ����                  6        8`�����P  �   86   H6            ����    ����                  `6                �Q  �   �6                    �����    � �   �6                    �����    � �   �6                    �����    � �    7                    �����    � �   P7                    ����     �   �7                    ����0    ; �   �7                    ����P    [ �   �7                    ����p �   8                    ����� �   08   @8            ����    ����                  X8                �n  �   �8                    �����    �   � �   �8                    �����    � �   �8                    ������������& �   (9   89            ����    ����                  P9                {  �   �9   �9            ����    ����                  �9                }  �   �9                    ����` �    :                    ����� �   (:                    ����� �   P:                    �����    � �   �:                    ����� �   �:                    ����  �   �:   �:            ����    ����                  �:                R�  �   (;                    ����0 �   P;                    ����P�=         8H �  �?         �K P# d=         VL �  �<         |O    �?         �O <# �?         �O H# T?         �P �" �@         2R 4$ $A         <R x$ (?         6U |" �=         �U �  �@         �U  $ X=         �V �  �?         �V # �?         �V 0# `A         W �$                     y5-�|�n��!8�ͷ��?�g($�jz���p�"pK<?����x�%�ٺ��(�3������E~;C\�l�~�����-v]�<�䣆kr�F��a%�]x�\#�g��u\��z�ܝV5wlo>a((�F�Z�P%�F��ڤW�5/�AI;0�1I�ѯ    ���4)�    "[��,��A"�5�w���.axo�*c�%ޫ�    t��I�j�p�K"5    ����ͦLڏ�Y�\ϔ���,B��r>(͂m_���1ͬjv���PP ��B�DxH�PIEa�h��X/9l����6I��Ge�=d=/�1�s�<��NF���bug-c�Uo��dQ`�ГM��:
������.��Hެ�s%�_:*���_�M����R�F�T<�&cC(��Fq��Ò�G]�,�oa̪���K�����q4�'j;}�a�4۠�6��n�
T�4)�R}ȧy�c��Ob��aBlY��6M��+yuOA��@l.m�O�I�f'�k�d���;��=�H���l������;�a��� ,,����L"�{����usj?�H�� 姑"�2_P&�:c�l.qw.�WR	4���#�̥��!�&h����lPv����Fb�    Sw�ޱ�����	Cz���gT�O4)��`��3gd�E�    |�ի��1��m1����%���#Et���{wSpu����U��}�x'�l}�\:�1�g��ȥ�F�B8x��ȗV<���8ST�M�]r��gh1`2�    �^ce��9�a�������H�i�rf    W��5n��Q    ��d�F|    ��c�    껹��#���I �Cx�����;:��{��[�%ʋ�2=�y�\����Z��c����s^��}�V}�`gH*Rx3k�p.ߏƓ�?�HD���8Y�0FK���S���N��-&+���0IO
C�-)N�A��5�<;�K;o���y��\�B|�l�=���-�UP�W��b"�:���[OKYPMU-0�+\G��    <�U����0����    ��# �[R�*�l��L��S�P�!��(�Dd^��\V帣u��5��~�a�ܖ�,��N�j�,u5��    Y�a8�����l�+���K���畕��!�B]� g�$Xt�a�*MB(��f4�i�    NG?�;}�%    K tYo��T�/�m�  1 )?�u�!��� G�.���W�7ʜ%^ z���ܓ�|%��&��*i�� ��LB��=F  �jėֽ���  l �Me�k���X���  �2��L��ǵ�<
����6�l,B�  �A*�ChKp�z��G�)��� m��W;"Jݘ7t� @)�ɇ�i#�W��	\������  � �O ��J�n	_Y�WX�+甑  j-�@"���QNi  �, ���]W��  ���l�Η�  �h�<Q��  �E����F�TP�n�Q� f� ' 	䔼�T�J  >q�zE ��v�-��?*  ���6Rz�J�m�Ԙ���0���f�$�P�f�  �/��h��  �����dq���m�7[$J�b  � c!�gm3��Q ��-�2��I��7*u  A���6WY[�>���  d��kVx _��{��{�l�Z� ~�\���Pn�!6��_�3w ��g0%�]<1  ��d��	/V����g34�. [  �תi^�.�rs�� � T�<)�#A@-F h��r�)��>{  G =�Y9:3v	:}���>  V�qDL�w[=���ѥ�4�{  b y͠�1}��(���r  Ky/��kv$��@��� FQ��M���=E���<I��i �dg�S��@`�@Ϋ�Gá�L� mO7Q9���2�+�b�����x�v�� � ~+�C����� K/C���-�p � ��r0��~N_
 N%��j�������  � अD'Ҝ��^Z�t^  G+]/����_/  ����]gq�wfV��H�  ['�dUa̕��e� O �<��S^���m ���z<��{  �����3��G��D  ����l�乁 ](��j�נ s��w7:<znK�r W��T  ��O��?��  �0�l������r���� � ;ʅ5���QiΒ��&K� g ��m�����y���p�C��i  �e%���v���Q�I�7��  k}*�T�"�Y�
��.1  t=��� ���-� ^qHg����l5$ j��Wn�=�Κ  �&��l%tK  ������Kt�a�  W��Xh'�N�,�+b P [�f���K��[�A!x.  ��TEl�$�� Z�>8I�#b��ёC ���O�_�<��  ��ssk��;&]�P  ���#G�
_�
  �!}k)F̄�:� �:P,���,M^  �/9J]�Z��u�d�N� a �.��8�_64  � S^Ϥtы��G"�uh�*� Fï����d�;�����X  �$�8$[�jLu,4 x0؛�`�����TD�����  =� q~Ky�D�BX���  F�k)(�
3�D�  � w�ҟ�lz�k�?g � �d��p.Cģ�ؐ� BZX�C��,f�g�5;  u�� �x�6�����8  ȋ������Z���dCI��  �M��m&�(I����  k�Cp���I�   @EYY�ҍV��  \ �(2�tP��W�O�  2�T��Aa{O��s��SbRw�.��h � GT�v�1d籡 P��;"��5 ���1�֘�N�4 ����3	�˦pn@Ko  o ̜�{�c��Rn-�ʀe|�o�SH  ���θ�,�R� >�������K� ��ov(  tM�F]c�"i��#  � ����q� q�d��s  ��LA�2�^nq�w�-��  :ЇO�z�=�] �(<z��u)e * ux��GŹg w���i�;Qk}���  � �G=q߆:i��F��$ �H���-�\V�Q~�  -ܞ�3���׼ď�  ��:c�Z �֚���N ���1\�s��G� �`�n7� �!pƲ7W�y� � ��E^YJ��e���  �[���K�>~  ����N�	/���Q~0�)]�r ;,X�Ơ[$��%  �u�|p���� ����U��`^��QQ��  D��?�f�x��}  �e�7("V�`Oic� OK<=Ĝ'Y�fO��  ���Bf�j��B�� B �DM�^��w�ظ�|o  J���;	� � up���  � {�`���%��H��  ��=��I��I�l'V Ú����?y���d��  ]���}����Pd�����  lz̩!Nu� ��A� /!�^k���&T���j  *s��� 
���f!�f�2-� ��A�&���c  hI�V�[  g��N�IY�N�C�,~> ��"�II �FM�J���  Hx�Si��WG((�c�XȻɺ� � �n���ozЊS {T�-,O>8�R����U�i�'v'  �ڙ��y�|��bB;E � u�	b�{��!� C �>���7�j8�  y�C~�R ���{F�v�F$  �=��%��?�����K�  f���*��C/ط:�:6}V��mqbݽ a��1��C����/HQ  ��ْz=:��Ƙ~  �R"z��h~d�}�  ` -����Ȯ�-�g%m D w#��x��I�� ��WtN�L w  �H����,�  �< l��qeB"�  2 ��.4������\6W0  - �l���)_����pa�  � �9Qa��Bx   � /U�P>�   � �tD�  j���z�C��5 , ���V�L�V3����
-  ����� >
�b5�O4�  E��C=��_{1�u����*  Ty�߫���"  � �6�>����E�∉��  s��]^�=P��\ b���mqF�㘣1 ��-�%���i �3�rVBM_���z	�  �=:�1�cC,Tہ$ > ��<&;��������|�  � Gg*�k,Q&I��iO B ek��m���'C�  �J5�;N(�����'�  ��{=�.�ʢߎ  ���`�&�QS��i�  �dAdO�/"�5�R  ���%�0˺?`u� �wl��o�M�|��1K  ��X�4_�ja8� = q����
�s:ۛ� 9 ��)䞏���.��  ���=�ͽ�Z�V��  %��\���0�yDE�,�<y� M0���z#b�Z�DXQ�+˾�P� �g���!-�m�u����i�  � ����� 0
 q�g�D��FOQ���u&���  s����zH�(��*��yɺv 1�wH�O���%fe � 5	Ö����'q�M   �|E*�Kh�u�5�kly5*���o{  2g����ić�b�'mq�� �!A�T,�)Z  ��?����\�`0 �Ow�@����OgĢ �f��r�����}�O�J �Qnœ��� (�Q� ������pǻ�|��x� ?�8�g����̀�h �ܬ)�HhA��{�O�c\)�i��J'/x :3A��# �����L.u�  G���H�L��lTI��	_ uz5��s�|�P��۟� ���zYԓ^��M  � ��>�D�R ϋ�Q�T���'��O_ � �����9V�%���  H�9}�Δ� 5 � pi��^�  ���p�:�m0�  ����ƤjWy���   Q��:��Ǐ  I �m1� ܀v~OS�_A� ��vkTyo� A؛UY  � 2#�: �s�=  A fb��:��֗����  �(�U�  ��/2�JE  ^�  � �?}M��;/���љ�U  ���1\d�{ �����џ� ���+�L� ��)��� =j8��  ��|��;�N�  � �����D��a�zM  @ӊ��%  (~�_24��dt   l�.|Ali�]5a���gI���  k�/�&0�� � o�%�ZU�H�  � �(N[�/>WP��  � b-���6�F8Mfl���1\�A�B  � ��({%�X�vx  � Ԓ�@,��c*�c � �l$���[@��Cz����T � �m�WAr�2, � �NT3#�| ^  � p��f.~�/V~�  � ���_�|���b � ��0�Qax���*��Q � ���.����In�ס|� � �5c��1+�  � �e8�R�^�~����sw}  � ���C#G�N�*`� Q'  � ��(�+�W�{8 � U�)N$#�u�P�Q��J� ������	 Y@��>0E�!  ���
�+d��%�ׯ���1�m �Ys�Ŷ6�e���5c�Y�้sKc���T�M�gw���rc����Պ��s�B  -�+���H����X<;���G� Ѽ���o�$^��D�[� L�K�d�y�ۖ���g�00���	�pZ�֝ ���_���z� a*u� � X����y�^�Aƙv@����w�]c󾖤c�DL�=��Yn�AL�>:�He_�<�ߐ(;'�ث��3�=�   ]P	�waMC��%+㕬��q�5��հ�W����(C���v, ���Ŀ��vM��iD�����*`�y��{Yev��_`eFS  ������(d��Nc�$Pk���~]EE�Ӿ]��Q����}qx�?Uvq3����"d�0,j�J�¤��)�0v�  ��A��%�|Tt�a��%0M ���Mz��|��7"�B�.fGɓ;�F�]��+��P.�a�����W�%�R��<�U9��gz JJ�l�'Q����աے�^�0=L�[G�	���f��w��"�t$!Ro�䥝Y\��ZbB2#Y��  �A]�"&����xH�ܸLS;"e7��v^U��X.����w���e5/h�1��v]��1���i�\�$r6;� ��B ��.�F�ŀ&�-� af��ێ�<`rX:,����S�����Zc��k�s/,/\�ėt���}�6�M1��T�rL����I���F  ��6t%��� f J*~!y/
�+�-�o�Æ� 2 ���6�ɬz���.>F��O=��  5 �������~tR, ����aFk�% i ���* 2$���X���53	u � ���0��툇��iy�  � `�nkk� *�U��<  � 	�<�>'ֳE�� �~�s�&Z�x  ��hZ����}i�4��D�7n�5(   ��P�M���}��u��'�:v & �����5G�x�����x  ( �+hi���S�G�����ֲ�uB�D % Zx �����P�� " z=���   ��e3u�+  �B��_8��F�z�x  ' ���Z���'�A�H�bm�q�� ;MU~l��my�4  :�+9@f��  s����)�Uc��X~;�v�   �;��� j�t1P�\�  �-�R�7�   ��P�VT��yVr  �^��G�%k{X�J��n���-�s�ʁ_ #�K��Z/��o  �	6b�4��t5 ��<�wY]@                    ��.H    �W          xW �W �W @�  P�  �W �W    svchost.dll ResetSSDT ServiceMain                                                                                   ��*�  �_���܈z\)��=��	�.7I�A�`�jQ���"�+*�F
��Ҫ?���{����?>��Ś�;�PKD]��G2��0��X�-쬯!E3V�_�RP��~�r�+Y��v�nOW"���D��M4�v��J6+�v�eY�\�H�L��I�t�e���لM΄�b��r���V{Y��n]�cl���j�2%��/�e����� 6^�a�p�����ɶ�H�0B�`�]I >=���I�L���L��n�nJ�����������>3_��&�2��e�,��ٕ �xb����T���`p���X_��*9l³B��I/�F��6#�Ck]�tŕQ8���%�� ���>����!���"kٻ�a�%ʱZ3�y�=����«�e!������IG@����3�/��^S�O���J
�6.E�����VM{H����[Fy�6-��^�c�� ���w��-b��K���<�O��J]��u�+��T�Y��+⨠��b���U�؎���k�b����ݬ��7�[��+J�i��
�����Yq�h�+mA��U�cR�ືvQ*��]�D�+�B����T;����Q�Ga��z����y����Q��l�+���ȳ�cJ����pJ's�����[5���wF���å��K�O�S�cٿ���kB>b�����=V��U~|�8�ete=�Ui�U��/�폋ޒ	��7�[ѥ����7G�L@�67SHͰKjO� �r��쾲�4��%�}�6E#��b�Y��b��T���O�P���(����/?�,��s}���}۷?{^��Q�
�'��u��� �n������6 zY�]����(Z�-��/�:�������ya��¾�SD%X�|����qo=~R��j/a��R��]�!8��C�ځ�OMy���˨?�v�]�.G��j>��mH�R�V��,T��n��;PP,Rd�Yv�j�'���3����ז�
♫n���#*����_�ݶ̅�cq��zjt����
,��<��I>�E��.d�����Mzü.\���w96��8���4�m
�)�jHlD�Zi���~O�9������Wu��R�yhjO��U^�R�f*
��/�ϏF<*���T1'�aNͿl�	�Ǝ��=j�������4�Թ�X��mW͓����85�"�QI�7�T�VHpx��OfW�$��q�dI��U��� ��̹��d�9b �@����-g"��`��a��j(C�jiE��0d\zy׬�`
��x$N=� 7y��4�>ɧG۪GU��^y�yB����k�P���AG�/<�7X4��JPo���V`s��ʕ�hl�ݴ�?ŚtyaP���6�8�ɺ�����ֶ6(U����u^L��g��_�2�:;Z��Y�U��G�	��S�c�0<CK�H���ьɋq��{%�Z9�"��tphf0[ܵ�>ם��XOTLG^-��������-0f�/3?A��pL��sn�w�H�4浖n�v�݆��b���ý�y/�ڊNdO$�����;˶�� ]!�(So
C;Vh�is�E�������O�Ԧ���:�˭'�Ut�I��Rđ�QD�;�3 �p���_�<t�ѨE��$��=P�O=��&U�Ⲯ�,�$���r�I�ut"�_�<�K�^@����C7�i�+�v����Ÿ�?���w�$��_��U����M,�~tJ���,� >j�m������}�͔���= ���I:d`���UI]_~��%4y�,����kk�!!-CǇ�r����6�4���rKs�{@�$ԙ�Q��~�U�%������<�Ā`��������曤���O�ލ���G��^K���W3L@���&P����̤���g���Q>�X�r�����zU��x�g#����]r�y�W��;Fu��I��!wT"�y��U�S���o��ͷz��u��'5�+��>�U7%:�ɛHח��H�Hu�(���܌	\�zwS�R'0�gZ������|�U�)��qt                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                  �  �   �   8  �               f   P  �                  h  �                 �                    �   ��  $          p�            B I N  ;�;" �8;k�}kk"��jL��.�%/ҡ�7�`�͔��7��$P���!���"(��Q�QB�t����Ыhg��݂؍"p��?;�JzO�?�i��]D:)�5�*�4����%NB��)�&���{R����
�OY_" R|���j�]V��=s�A&��Ϋ,� ��	�D��g@�����˱���}>:C��Tk�ý�|�1Q�	��9�m+�F�j�f:��h�^I��&h|-�N����~�e��r���x}$S釦'^J�M��}�H�%+vN���\���0H-B�	t� �*I��g����Ey=�]x˧�<��-H��:��Y�V�x���Ax�/�3�� i/J�3NsSM����{W'O������rA�>�J�f.�E�:F��γK wM��k0�s�d)��z�gXkp>x��"l"6�ؓa4O2G��\s�}T��v@�2T猅\ wu�Ưո������.;-?=<D_&I�!�U�[�H�3�zy�vs`���qr��=Aq��(GK��%pO`v�i��ϸ��I�i�O1������fJ�fca��#+ʩ^-�����2�P�}O1���C�c#�~q��,qGn{����˙|i�lKgн�a�����[ߤ�h,N7�F	x}�0�<�z3!Y�=��M}@ 9d8P2��_���Idyg,�#<4���1��F��.|�<�ڤĻ톷�<��K��eE�*J�&��[�R�B��j�E��̛?�ӑ���ꞛ����
��7�q"���Ǉ���.�У��	�-F+>��}(5��Z�[$$��sJ�v���%��"�D��s�a_���@ˇ��?t��+��'ъV��b`�+^K:K!�9*cC�4bT%����:*���l���C�`"��ge��%D�+k~��S{�Ma(���Z�a^y��c���n��,.w�"�9�پS�d12M4�޶Ak3��(Nӳ�T�\A�V�����p�����ZrM�N.dv�����`U��څ�t��2����@dg���A�Du������cW��#�e�\M%��A��z��wP��
��I��[Z����N�\�]eAv#�s{yI�_ ����H��e�k�V��VH��?�����V���l�?m�xuW�o�c���E�n���M�RD��y����R�޻=�?�W�$��&�1���f=8l1���1K��e��q�O��zAcg�S�4�C\�/h\TP�:��1"����\xp�,�/�s��G��|e�w�Ȉ�)���?�@�{�=_K�V�5�5D/�I���Ӗ--7M��x g�qe^p]	|b�Ů���Q���Q�� �CЕ�S�u
9����q��%�Bȹؒ��DR�iw%������c6;�6򙎺�����iJ�m=g�3��5L�x�b1w����!5X��Isd>��#ꋻsC��g�P2��ôE�_�o������9� Ƒo:aI�����O�'W\�X@�Ж_!9,����"a�A4�.�N#*f'����'�Qă��ޯ+8�^LCk�\�Pr��Tto��u���A}�`��&��QsZ��,٨��S�+u�R ]Xi��7�1O���O�,��/j�J��"æ���.3�-'�g�Y���G@3��F����O��J���^��D�&��;dā�5��!��+�|�ލvۉQz���ƈâ}F�|���=I_�}�YD�v̝�J�9�EjFR+`RF{\\<"٧.}	�4���7T��8�Рg˂ӿGC���)b'���B�Cزaoԗ��f��$:t�(ެ�5�|R.����<:�Y��J|>��?��}L���u���ѿE�>�(��k�3.�H�3tR���e��P��%���PU#��#�a�k��Ex]Ul�ξ�����~���|\ �N	a������*���8��d����2c�:HLlM��>\���(���' ������th�<j��7�8m(�d�?AF����W��Ӊ3�ټE� �$�)�_?ոŜ����^��F�8�x�&^�'{�Y�{�\w���ʹow�bn�V�-;R�x�i_�;]zp?	�˩D���]P ��]]���Z>�ъ��.@���a���qM�b�,a��T\-��͆�-���4yI�P �Y�ab ,QH�F�����A�l�a�+J�� ��T��������z����)���d�ރ4z
e�1�{Um$<�:D+��,a��
�E���e��ZMA���,K����c���M����_��8���7R6g]�gӳ�r�*'#�H�D��5w���X-�92�6\b����`� ���-B�6��"�6ɵ)�z�&�G՞�Z∯O����&���<�q�mB��Be��0GѸ��Oi�j���<���������.���O��{����Jz�<r����[\��o��`�P�%~�$-%��c�۶"��(ш���x������F�鈯��xE�~�x6�����N�G{tk�+.��}-��4�o�#�I疡1n]V�!�d��M�sb� D�r�+J��[~����t4};�ѩ]�S�jN#8sF@Qv�(y��m�o"�?Mu�� �����V�S����ë++�@AC|b����23��U��������
v�~o)'r<�%���x��/s����W�&���4�6`�k3V��'DM�ϔlu��"wlC}�J9S[C\���M9��i2��h��i�r#jt�ݠ1��p�b��e�G�'W{@l<u%�M�v��������Ћ�Gu�u���
yc/���8�7첢ՠ��&�jWu��=
�hImq`�)����tLv��S��1��F3,���~@�A����u��pun�n�#�M<n���$�I�D�׾��>
�-S��A���\�;h��`Sg"6�����r\F���ۃɿ�H
]�m�L�D�U��ei�â1�L�_uC^�^x�8���Ӄ����6S��*�%jCM�p�_�y��Gi�zc ���˅�}$��g�W��Ѹ�bl��/��65��3_��ɪ�)P�M�ƒc�α';�Վܫc�`�'9����"��~tc�AB�������9���L�D�\��D�
����|L�#�!��U;*Dށ��ۀ�X������On֊��4�����"Z��P~�V[L�.Ww_L�Fd}��[oJ���Ҿ��}9qq����5y��CR$r��X���¥h/'u�Xb� 糜T�1���-�YB�$�Wl�Y3��FZ���
��M"CʼU�B��f7����_?lFKa���s7J��4DlFfBa`�Hs�vSaK+8�	���>1�'�LڻޥO'_����yTa�^	��L�&S�i=�i�&��MBdÕU  
3s�����Q�k["If1�G��8�Kl/_='��w�K-�[C���}�e�mԽ�Dr;v3�k�T`�ϫ

*�t�@�9��J���V���GAG����}��"��R�F������'�XRՔ��3��r+3��F��׎Pe�VO#$��#�AJ�В���c�UU�aP�X:��y���1P)���*�W��w�����,r�|	�qAr���sMD��;�L,!��7Ȉ��E���a�� �Wn���_0����a�&�����c�}��o*g�H��	%��98_�I��d:Q�"���H��\�+�����4'9�碲+�{u���bu}Y�XnD��Bj�y�հ�tU��U$Wq���Gfk�M����)�#KC�˺�������C�
�:Sd��A~���|���;D�=0+ LT��CSo�-sDr鰕H�_�|�ً����F��KK�A��o�q��ߺ��ю�\�暦X7��C�+�y �2RH(��8�>a]q��˗ ��V,J��U�xx�/�<g�,��Ó��[rR��f/ؾ>��T^��]��x1�[�%��|�#�D*<R����~P�p
>� ��=W:gAa��X��^��^j<^�<����JM���i��]MF��^t�B�L� {$}՚�T=876x\��)�w@�
Q�3�%��O� 4q�B踝��N��s<R��t��A�z�`o5��O\�W(�%���؍L4�g�o��.,޿��[ �+��/�d_���T�;m��e����Q&�rع�s-+�R�n�/��W	>Ҽ�p�/="c`�R_��L�� ��J�CcCR�Oq����Q�������a�4�V����H���l
����)���Ĺ��4�6�ޘ_f��1�!���iI�D�Y��u=ė�Iq/>���4\b�h���r������_"�K��`��[�N���e�]����W	k�4�zj
���0���2��_P%0eBZ���)�����5[ݥ*�_p�K��8/CT����U5��A���41T�r2\ސ���$tk�w��
X(�!{l���'B'�D$R�͖���Q��c"wr~o���&�_�,v]o�n��>�?;��V�MP|n�[�#sg�5��v@F(g�V�ZP�x0PP�º�Xl9s�^>m�9;6��7+�9��Q�(q�؇a����[xsF���l��"8���َP�(�t�_o��(��P�D�н�
o��%�J#�V��*`���54��1F�?M�C����G^�]L%I�Y"����E�$�:ג_��װ{LN5Q0׮~�$W�+�&�k"]`�MYG���s�N��=�/v]6���ApTfY�}v1���ʍ�~�Řh�>q �_]KI���d�zj�&��wݫ;#�̎�р����[��J�x�w���Vlf�[,��8��B�]���h"�"��;��p"de",�Ǹ��S���a�,>ڈGp��ti�ڋPg��Wcdc�A��?���{�/!��
��űJ�<m���5�VZ�g��*�����I� JI�����E	�n+ǰ�P�x8DZ)a����;�#/�d�M^ ����{C�؋��l2�<]U�-��i5E.�*HF�)��ۭ����H8��H�팗#G��U�s�'�
�J{���-G"N���Cnf�qX�'S!�3wI-w��Ky�Ls�yL�&/f$�fq�rIp��	�O�x�A�^�'��%��j�b�OES&�÷�R�l7��K�eѫ�`��{Wm6ύy��C9� ��F�@���ݡ�uR�I��Ie&�/���:5(^�l���x�3���Kf��2�<�/(zQБ��&5��"+�=��Q���I|ǳ@>gӞ}��&J�i�n�����B�x�!�*.ht���]�}L��aa3�y���wE->�7������`E�*qS������C8��'Z��m�!���hQ�7�2K:y�����BIz?s�v�x�U�������@c����I�Te�}B6���t�U ��l��{��'�)P�J�U�>[���u��sR.N�D�nF�&t��P*�D�V��8%���v��o�]��`��q�B~p��R�x���b�M�\=�-��it%��d�����*���x��}���d�]a?��*�nF��4��r�H|Y_�k�?�^�@�<��������K8�P̐�|�����Pe4�[�u=�ʙq�-�.�\Sc�rE��"y�GGhJ�#���E��m�	��,�ƅ���-Yְ S�_��Y��)�痕��q�L��Fi
�ԉn��t��)�� E`�_���Y֗�w�N2Ko@��)C�k�	qJ-�S�d�=��g��؊��	�c.�Ϋ�)�0���I�17�'g�,m+ǜ5���k�����x`hD�<�F���s���|Y��q��'����嵥$la���%��\�1��Faa��p9��)O�ٷ@��
��٣oNovE=��z�^OX�v��ʹ�z�$m���꺁���<���]c�r\&T�UЈ/�Ē�S�2`c�[�Ko��%�l���cwv:�\��jj"�D�"��'R�$����8Q�� Xb��� ���$�3���Uj8a�@ �H:�/`x�'�1/�6���pz�2�r.��ϾL����mɖ�����_?�C����+I��i��<�V0��9#��w�z-�o�}�zx��Ea���'����W'��
�6nCN�@���h/�0�65j�P��J:n��9��r)j���t �dhϏZ�	�7/��ܥ�O�2�KI�=K�D*��V��i�P��s��`�H�fΣCs�D��Qh��]�X��j������Ab�?x��ρQ�ԭ6��}���{���|�
̻���fWI���!��fҭ��h�l�/�?������0�>�oB��!I��Q����ȸ`�*���Tk5x��G���V�e���>��
�o�#�V)���v1���p��W1����l�K�y�ޣn������.�=�p�{V�'i1|��������ĉ�L��	\�����xY�{Yy1��R@6��x
��gw|��0T�@��1\aؘ�
^�+	~����	5�AV�sx��S��f� ��i"����4]�0�k#L����|�>=bLHIޟ��>����s��h/UzF�g7õct<�����v?�AizS~\��-z�{�_�Y2}=VRSO/=R_�hAh��#f��<�>|j�K!C\����H��"�                                                                                                                                                                                                                                      44;�� [}�s������n6��N�MP4��r�S�?�dl�b�}�-�p�0�C��ț��.y��G@������C���u�{JJI����-�� ťMb����ٰ��nA~/9�:��8�A'�J��}|����uk��Д��(ƨ!` c��$�#(�q�+Y^���w��%�2�Ӥ˘�Sg��k��(T�1��E�k�D�<6�]`���j���<�t@E,�;�JjD�,.��Jڷ1�@{)E;ܗi�lO.�w%
jBa9�I��`4����U�|[�%_U~s�$�O�:c�q����?GS6x_���G&�?o�B�E1<�
��h� ����a��z��^զ?���\��3~Y�v�k�u2(�YH��k�mQm}�q�׈���A�AU��T�<?\�q̃U+����axKSᲠ:�u�PQ	�kIMQ^9J�N�E*�Ga~�1�I���_b����
��Gz�M�6�'��{l�y-� ������N�RF���_��Yl�\�a����B���9�����;�o�^s,�ϵ- ��@j��蚜Z��3G����jV@؟�=>��湊��4�5�z��P��3�q�pW�SF�J����i��U�+S����IH���ۏ���H�)קlB<�V�&E)�&o���1��G�G��u�бb��T���O���(뜾�v$X�gt�����wR�|�
����i�������E�+��|�u�[F�=	��L.��k�T���-%ڼ����tB���m|���yXU��4����P-���Ncʍh�q�-�I���p�;9��W�r�FAtsQJ��'�+�v4�0��N�ffܕF���C��$kf��H�߸{q�p�����~2��Ν�?x�"����z��#�l�w;wU�����
؍���������?��*�����B��0�;�X~3s
�"{H4�Ġ�n��O������h؝�ƹ`�)T�v/! 0#����H�������՘a&�׬z�W�A�Yc9�X{]'�`�[S�LJ�D4[ z+�ұ"7����{u�?��ݑ5�~���KH��/��;7G�O.4�?�y�c�s���ş���}@��E�d�e��j�����!xvW3I�2���2�,�T�[�n	�H�?��Ծ��{ŵs�7�@��^��a��(.��'�:�~��%�9g��*��?��]�ӯ�g��Ƹ��I���q��0dV�g���(#Κ+�;qGj菋h|?1���ʈ�E���i8F
��'�	E��2�(qx'O��rD���+��rs�Q|-��A�ǷX��Q��6u`(��,<�j�����o�|`h���:���79�	Ϊ�p%8�����K��xuԶ�Q��/]�ؙTY���ˣ�菲<quPR���o���@��_
���^��ʭ�(��o�39%�Т.�ڪ+�1ι���t�����[f!WiR;�簃��>Z�y���T)|�G����T�w>� t*ɏ}<]�5B/II)9�{�kw|1of>Ho!,<%A��׉�V���h�A׹�ߩǽ6�h�9��U*rWZ��{�8�����d�tv����I�L�F �H�2 ����|����Q&����Ia��<��:�� 0�Ù7� �D�԰���N��E��V��ł��}Ԇ��ƞg���ӓP>�ݥ^hS/�}��o������؄!Z�]*�}X�}��&Z~�s+>��	��1�6'ev�d�O��8PD��u��T~�枓�=U�Q��r�N��!�t�j�{�2f�o$����?�ML�Z�sU�1ףto[�P���a�@ࠛJ%�L=����O^�e�o�֢h��k�����b1��;�s`$�	��˻]l���#�q.0�A�3l'X�.���C��sk�������)�q�Uwb2����-U�Wy�#G���n4������]�e�`�Ǹs��<��+������M��$�z�b	G�ڭ��[���O5�t�bsL(�3Br��Q>ߢ:�V}�}��F�WX:�'Q���eD�=�;�v6�f(c��u�����~�Ҽ�}��m�����o�6��!P@?�I�t=�F�����N�WF������������	(fn�y�mq��aM ,��5��t�7K�k,.-�[q;)cg�}��Q~Ig���[��q����ł�ƭc�=Y��R_?6�ܼ���o�搡풚�~0����/��T�] �᚟�m%�ä;�{Ѣ�3����A��D	:X�E����Wiܲ��5��[�p�)E��ݍ�p�R���C+��S�����X�U���Q�~����YM`�q�F�zL��LP��|G�T�t0\��]��%��:�0�M�\q�![��#kv�"�g�`w�D��י+����+�J���G��V�2�?%�Wk�
�u���Zy/o���U��eЋh�B�g�HK�}�d�u�9��]��$��J�,��5efVᑗL�(�I�z��?T�����o�gf�;�^ҋvS �����\�wy�I�1z`+�rG�A1X�������I�:����ԙ^�g[T=�69���g{����;�u���W����Ɓ�~ �����&i2c�U���clP�����A��0g���1g�Cv��uSW�{���E���Ze3@�piӉ��up������}�$�Q3_~s㓠Y�[����;b��°ꖏ��l�9`�CѦL�KM$7B��K��}�5�ЂMEm��,5-�U�U�����������	�3���X@�R.yG�ճ�ݱA�x��ӛH"3��P���-�<��o��2Ԁc*T��S]'�ȅ	���G�kC:w�*�$\�*����7���9�&�38���/�7��be;�vW�����{                                                                                                                                              �`�   ��]EU��   �]�����݁� � �}Mu�t$(���]Nu1�ESPS���	  �E5P�                               ����#PPEN[��t������#t53�Vj V�uN��^�� u$3ҋEA��tRR�u5�ЋE5��th �  j �u5�U=[�aujX� 3����@� �   _�u
{���WD-b�)�O����Y�   ���^?Uj[��67����   /<�K(A�'�}r�@y�l5f���I_^��9  V�   �!F4]ң�Y��*��[Y��  f�ދ��[zq��yq�    9~�,�����&rQf�ө�_��gyC��c���Ճ��Í��;��   �   �1   �E�˨�f�T��C��>��J�����F�����3�i�%���Ƈ��R#��~ %�E�q|;4��]�-2B�!ƞ%�J�Y'	�
����4�&�pmr�z��L�'g&��3�'4���5��"�5����ˆ��<��4c��`��.������
>wd�� ����4�&�?H��D��ǐ��n��W���C��?+��?�4�&~M[�bH6/�&s����Z���z��en]�u�,��E/���!mm�]4y"�ݏ�E&��m��ѼQ0�P�[�m-�tLP\)�#��E���m��A�^�f	���M^��enX�Ģ���m��A����m-�E*�vkއ"�;N1�rOQ\6����|t�k�u���É����{��C��'��m �t/ǈ��T�yC���",�����mF��m-���Ë��_��G�������P\)����ݑxJ
D����m��'/��D�ym�P�{�v�y�%��	*.0�Nw�y���n�
M��y�$Sձ]H@K$��"��7C�R�ð�m�y��K�Q8�q�Cl�y�1ٙ��sݿxUM�[xV�pm����ٳu&r�D~�	�DÆ�H�E���]U�fy�� �@'�WЛ�oIN�HNT�ɏ�oH�l�Q��o�{(6�KF���E�]��h�o����������o��s%b� �pSh˗o������o��{��oЛ�oЛ���m����G"�wyph	�o��(&T��o)��c��(ԛ�os1�Л�oЛ�oЛ�oЛ�o]0�sЛ0蛥o���wܛ����0a���Qٔo�:qܛ�vY��o�KfXܞ�o�[}p����A��oЅ��a�o�&""ܛ��Q͔o�o��Л����o[�n�Q͔o�&��Q��o�&UtI<pЛ1!'Ux[�vЛ7�"Y���F����o��o��Ԙ�c�W����cՐؿ���̕�vv܌us0�����Qٔo�K���o�vn&"U���"Y���C��t��o]^�Rat�����o[�n�QҔo�&U|I�sЛf�Ѕ����Ȑ�F�qЅ�Iw@�vЛ}pЛ��Л�oЛ�o!��!z[h��6#{$�:�w^�c��n
w�����Q���eF��w^�c����Л�u�����Q���ۗ����熐��d�%�9�ͦ��w^�c����c҄��^�z��T��8��oН�d�%�9�ͦ��w^�c��o��h���oН�d�%�9�ͦ��w^�c��o�I["��s1{Y����w^�c�h4�oЛ�����熝��d�%�9��X��rР��В�o��TJ["�_s1{Y����e�u"�����}���w'�9���W�����Y"�����}��wH�l�&�%K�wЛ�o�o���ow�oО�Л�o�[=�]�vЛ�[Ֆ/Đmh]�vЛ(���oI(�vЛ ]`	qЛ�~Л���ޱ���X%�u�Y��o�`�"��"Л�2��a���!w�ܱ^}�^���XYQw���x���v���[���]YQ�%�g.J�N4��c������f��s2�񈠇^om�/N�*��\����ӭe���8Л�oЛ�oЛ�oЛ�oЛ�oЛ�oЛ�o���o\�o̔oЫ�oЛ�oЛ�o���oЛ�oЛ�p�SNqО�oЛ�oЛ�oЛ�oЛ�oЛ�p��U,�@XB�㼧M/�t��?Iީ�7��4R�ɂ���l!D�淭�LS�Ka:�� ��G��� D�!y@��)ed%2-��@�a�?�}g��:�DFB{/R����oS�;��7u
i["��,-V����#!�Y`ېخ�$� [jA����Л����ݝ��?�R�O�w[�S�2:���O�i�K�d���랝[V����[c�q�                                                                                                                                                                                                                  � .� A�         kernel32.dll   GetProcAddress   GetModuleHandleA   LoadLibraryA             � ��             �� ��             �� ��             �� ��             �� ��             �� ��             � ��             � ��             � ��             &� ��             2� ��             <� ��             H� ��             U� ��             a� ��             k� �             x� 
�             �� �                     user32.dll gdi32.dll advapi32.dll shell32.dll shlwapi.dll msvcrt.dll winmm.dll ws2_32.dll msvcp60.dll imm32.dll wininet.dll avicap32.dll msvfw32.dll psapi.dll wtsapi32.dll oleaut32.dll kernel32.dll �     '�     0�     ;�     U�     d�     p�       �    �     ��     ��     ��     �      �     7�     G�     ]�       SetCapture   BitBlt   LsaClose   SHGetSpecialFolderPathA   SHDeleteKeyA   _strnicmp   waveOutClose   ?_Eos@?$basic_string@DU?$char_traits@D@std@@V?$allocator@D@2@@std@@AAEXI@Z   ImmReleaseContext   InternetOpenA   capGetDriverDescriptionA   ICSeqCompressFrame   GetModuleFileNameExA   WTSFreeMemory   VariantChangeTypeEx   RaiseException   4   V S _ V E R S I O N _ I N F O   4 ���               ?                        t    S t r i n g F i l e I n f o   P    0 8 0 4 0 4 B 0      C o m m e n t s       L ,  C o m p a n y N a m e     M i c r o s o f t   C o r p o r a t i o n   x P  F i l e D e s c r i p t i o n     . N e t   F r a m e w o r k   S e r v i c e   P a c k   A p p l i c a t i o n   8   F i l e V e r s i o n     3 ,   5 ,   0 ,   0     t R  I n t e r n a l N a m e   M i c r o s o f t ( R )   W i n d o w s ( R )   O p e r a t i n g   S y s t e m     H "  L e g a l C o p y r i g h t   C o p y r i g h t   ?   2 0 0 8     ,   L e g a l T r a d e m a r k s         @   O r i g i n a l F i l e n a m e   s v c h o s t . d l l   $   P r i v a t e B u i l d       t R  P r o d u c t N a m e     M i c r o s o f t ( R )   W i n d o w s ( R )   O p e r a t i n g   S y s t e m     <   P r o d u c t V e r s i o n   3 ,   5 ,   0 ,   0     $   S p e c i a l B u i l d       D     V a r F i l e I n f o     $    T r a n s l a t i o n     ��8pa,�W\80C���I ��x�%o�P$0�Y�|(�D�@�L��P�D��(Y�$�o"0D� ��^P�3�
+�(� '&���p8$@ Strin5gX�P ��3�, �"	�D�Ȉ�+���	T Object� %��C���� �Ȱ�r� 9���G�# ���Ȑ�r�9��"�#��|Lx�p9lh"d #`�\�X�Tr�9PL H#D� �����r@9<� �#����� ��{E� S�	ļ�
  �T�#�� D$,�t �\0��8�[�B,��<4L��x #(�$� �| SV�1LD� >�u:yhg�j�� ۋȅ �u31�^� �H�C�J�}�����<� @B��d>u�x� �Y��T@�GX��`�� 'ϖ��I� ��P�Vg8���bX� B(�g P��
�Q R�e>�ÐWU����v$ �b`C��j]���;������PS� uH�� Q'��
F�P iN;�uWQ�������ֆ� �+P��� 
jZ]_����tH (�����2 ��;�rl��aJ� ]n���w^P$� м��)� ��{r
@De��<�=a�����} 0P��)ws6 �&*�y�$+�]|������� ��j��$� :a�;����Y������C ���8N
}9� 7T���� ����s jh V��B� ��;�� t#��$�PH �dJ�"�9�} ��UO��d��I�?�HTa<j�P�:��,S� y��)%1$�� �w��ZI l��L!$�ǘ�4��f�T��W	0���*{P�O�IQ �$s��wF��C�5��tPj����v�k� ueVSsA�
 �,��	� ߁�Yu��`���|pB����6" *+��% �
��j�� �tǅ!�� ��C�yw �I 8�� Q�L�(�+�F�T5��<�s^ ~��v ��m����c �DX@+�WHSZ��R���6���P�>����t�,&� �����e 4��u�? ����+)A�D8,;��}�
 ��U��� �@t�B!)�E��8�X/�`7���?��簾�]��;,�J�אU�_��rwH �F7IhY>
,5ϟݠ�A��� �H/!�̱>�� �<$\��<#C�觬�Y� �7G�\K t��
?�vP=bX��U(u��TW� *���I��P�+����hV� /ӽ]�g3 7I*ɆRd�T�`��Ԍ��m ��@N��� G�4�&�f ��K��H�k�� �$I�[ئHz�T!�f 8�(�@�O:�	RD��J�� ��i"#��h.ōk ���6 ��;� s[�� t+b Ӌ���H�uO ��\ ��)t�e� ��9� �G���� �%�!<;�RzU�@�p�� ���hn�K d�2ω"j 0(ɀ=6 A@~R
"�aw����(h%����1��-�= F�5/��
�3ɀ��� @=T�u� �p'X��b |�(��ZYh��u� R��#��w!�堅.]��S| L�����u�R)KȐh��,��'�Q��� �<H�J4=ų����q�,�	t�2c�^��u�+Y�ڼ���
 N��[�S��0|	Ƀ F�H��!�8m`��y� �����Ք ͼ
��$R	��7�.`��Ƃ8���	�H��D0���LJ��r�v ~�� u�ȅ �z����������������0��a����(|�B�L�F`�9&���Ѓ� �����  2�� <n:|�� _+,�*RJ
�� 
��M� 3�	%t1*�ڰT� d+���3����� �0*;����F� r+�;p�X��� �	UEd=��3���
g�% Z>����$� uvx�U� 2�F��# z�K�,��� 	�E�\fM�?]�g��A7+�R���`�d��� ���})k�S ��f'���% ��F�W� ,���y�0��+@��	���
Msh��:�
���� ?5��,�` �YZ�H�k 0�߉s�9 ƃ�ɕ@���7��Қ5��� �L.M	��� �D�\ [��:i�C� ÒZ��, @<|K!9<�����3��K.�e��� ~�	��Rb �!�+�A�� 0�B�Q�D�Y������xi	kgA�`����� �J"5���ЂF;|RP�&� g�{)G  ��It$�?Ɓ�׫3�-�=z�$��2YHm �^o�57�} >M�!]�� ��l���t� 	�s�3�6 >�Ė{�u �8!ƾ�^̍� R!�aJZ1�P`ւ�]�  �=!� (\݉T� ��u)^�� 	���A�"�轀 2�t)�w� X�(��l& ~{I�1���B�(p�� ��crhqg$�� AN�� ���(�= ;cH�)
�}S����E	 �5�(�� )�v
~y��L2K�L�,>�ܼ��� �<��֒�&MXj (�;u�= &�k�O N�]lԒU�����@�S�) 
����r ��Uh�!-& 1�Ã���Fe�� �\� ��A��l\͚�&}cty������HBP
�pA* y	pK�| ���Q�� =7D�
�M�m.k��ap��)�U�r��!�*,'S�;� �J)��T�c*�b@�^U �R2D��	Aq�B�=��VK�t& ]�I$�Q�< d�,R(��qg�ؽj��� ���F"���\���@u��C	 �x�y�dh J�%����:v.���tE�;���P �gU���� L?
�0H+� ;�F�V &�ifW��: 	�;=Hu, �q�V�.� ��@~�� �pi*���� ��t���\���7�: �)���xA� m]1O $��Q�f 2(ӈ�%��=M��"]���Ԃu L�� �D�����U=��x�LS��� �;��P��-����� ��u8��)LS� ��g}�|��� %2)�� �b`3����̚s����@���pS] P�y��>�� I5M< �Ƕ ꫄�g�.� #|S��6h=֌<r� 5��P 4,�%� ��u�� �{���j��?߱ M%x¡}�e;���J����&@�$�,�ʇM�L��@� ��Hc�:�4�$��) .=V� !��+��z3 �t	@w�P �J
��� ����t�nt� ;�"9F%� ��A�� �]��6�l ��3�XH �,b��O� }�8��*�ˑ�S������ }g�@%_.8/ �
�Y0 �b�I��<U�?܁�duH ���%t2 |P�q� B �Yu��$v��:����e �Щ�2��O I����� ��Z��H ���P�y� �L���z ��&��������� ���� ������� ���XPR Q�.���ż|Z D�1�f�TP�B�Q��ҋ���2�Ȁ��_�� �9�	wt /`)x*?� ���Ҥ81t���:|PS�X�f i�C�@�/	�P��?�@��@�v� �;"uS{q�@�� ��4_%�� �C�� P����!����p X��6(� '="|��_H����։ {���w8�x�4hK1�$v�"��2�� wƣ:��� ��[m=��� h�/@|K�����Lc�P��X�� As�g�E�k<f���!@�U���ic������$< ʽ��]x��,ߎ��XZ�l ��ٺ:- I�%��(? ,�Y	=��1B��"��)��r@ ����ڎpF �r8�?w �с�G�#�z��*v�H`� ��1I�d� 
�hAb@�� �	(���P��$Q�ΰ��&��?� 9�uEN��Y��Z�;\8� H9¼N��X�� ��^�� t6�:
u0�TO>NJ~�����1 R��8�z� ��ޥ����e1PE��� C��fQ�24	��M`m_ @i�+�.B�; ���L� HR0>&ϋ �1�)��r� ې(��L>0 C���� }��-����G�HL���a�O�A)��, � �Ҋ DĐ+Ku���H�@�c����L�L�P%�s�ƿ�� �F�� t���-�i�
 +�f$�x� aX�\.0�*(��OBJ�`?  �g4�� 0$	w,9� �(���� ذU4u��\p�`�|Y1 �2s��� j��~�=x� �)�����Q� J��;�2t ��ar� >�T vw���
ɿ��Z`]���P���* B��t@� (��u�Z!<�4 �9swI Q5D�B�E �6R؄Z�?&W?J	��Q�� �V a� ��Xe_�	Ð|؀��LY	�K� ��R �"���%��hb3��pYX�Xu��-�%$ ���Q�| >�����\,�S�0� O����P�j�h\�����`�Ok ̔M�-Uhu5 d�s0� � E���`�P�� "ixk�� �g,�<� c��
�f �q;P���� ~���?��*f�p�SOFTWARE�\Bo rland�Dw ephi�RTpL FPUMask V�lueRi, ��ӸEf�;p� p�1ɊA�.l�Pt����Gp��X����� �u�6���� v�X� -Ep��	u� ����2�xJ�H*5��n��&Od�xe0����� ��yG��ŸOڲ 1Q�K��׫���A��!��e`zY���c92 �,�Xl<Q$4[�g����9�?y�������{���48 �Iu �;�pg� n9��ِ'u �ð,ąW��hd������ �Q��f���
YVd@�X;)� \G�ޑ[��` �Q<XS��sP	`�|�(��g`��:��zX�[����a���R(QS�
���A� .tdn9� i�% -|����	 
[YZ�c �,� $t��P�X� 10]!�`� �RN�TD	 �X���� ����u� �=I�vj	�k߁����#� RL�Pb Tjd=�) �ɘ����J�(�P��s��U�`�d
~SI��o �A�z9 0a*
�u��� �� �v|hNM��kڑn�8Y�Z�(�R D�����v �X��4� 8B;��?�dE�0�ި�P\� tn��9jI;���2��Q ��"�^���W� ����t07����	�v)��w kJ mP��e�9 C�"x��0� {.��+�;(�VPP� ����=���t��H S1۾j&�d��Q(��h?�/ � ӛ��k| $D8��Pmq� �o��_>�G�kQ1�`W� ���6���P'���A8] /�jmEH,�s tH&�8R �u
�� 1�!M",' D=���Y� q	���O �C�%Z?��� BA@�;sO 3ud��W� iq�	DB� /��tƌ�Li�uЃ@K��y&�R' ���bA �F���6�;�Y�����'"��l�����٘V���0�[M�I���F�V �H���c� ���I�� �GT�B�L1��o�j�����V�D$�9�(ZTUW�S� �J�j"/{ )�TC0�5���u�!�
�X��=:` �����R�ub %1���$Y��� oS�I�#:Z �d�Kt�D]�' ��� �,M/f1�� (4�)��t% �/�F���H��� ��[t\*� �DW-[ ��~�=�X�?�` q��?�� M�6�0�R= ��*8(-��� .F$�: ��0/P�� &�,���*����G��"'�@>!������������
���'��C�4����LRs"�]��$ )�&@S��L=�tpE�8%�26�@��=�;��S`�C. t�q�| ��c��lD �C��%F b�7��
��I	Q#=�m�`�R$�
�[�wM���h ���j4��\�- G9�Huep �S.	���tC9��;"@��� Eh������L>VpW�@K���(��~��3D�j I��$�����Y����#� �zi��>� X�`�����T03t�Tx^B@4�;�~@ ߸>)�'6�(��`\b Q��� �}� ����l�! ���-B��������M�� �7���}�L�h� ���O�� RE���,HY��Đt. ��%�}�o A�ă=�{	u�C$!��h��6H0, F��ӕE�D���S�F�I�' ���O ���NH�Ȑ�`<�˶ǀݿ�8�� \�ZD�JK��<8� ��)�P����DYp��@�� �PW�� ��Ѩ$�� ���3w  �7N>�V �]T�s�=�	wXɁ���(��P��b4 �{U���?�^�����S v��1��#u	� 8tG�7%� 4���(P	��B �D�� �-�>0� ��H�r& ���o"�8�Pl�K 
��$�Cf�+v·%P����_-X�� ;�t�"��o�-0� S(��� ��;�Ao `�ˋ�V {	��8^�� Porti�ns yC=p@�?gh z(c)�19 83,ӯ��m �S���0�黭��#�|K� ��.8�J -��I|���@�P�B��� Xx�`A֋ �U�,� V)[�N� �l3Q$EA9��Bpu�^'&��H;O�Zi�x��n�|��L�R D
~_*��;p�P�U	� aZ���po�����F��^�2��\���� �����	G���5�E�s�n%;�i��]��?٘? ��	�Ǩ#>�g ��Hx},� �N	� PSU��{H �b�~t  ǓΣ"-3��S&��L�U�D�� �F��I���R����U, �hq$!,R:� �E1���&�%� ��kB��Z)�A�@�$T0 -Rf;b � 
[L�2��4�� h�:bv�!v\)<��B J�WPQ��ރ�����X�� ��_*`J�� p3���G� �w��5?�  �����4 p��y����9Pΰ�$',z�N&�؏j�J�� �(�7a>��B�;��\ �ZPG�0O�5W)�X����_ �F�u��B�؋Kl� ��c�X � C\�3O� ���q��� jQ�T�R P�@�L�O �KA�Jq �VZ0ƋD �o���4�TΦ� u颂��J1ZX��^��ඈ O�9�BǏ�� ihQ�k�G�7W0 yw �R���O99" XJ@N_�K���ǡ����ZX�* ", 8@A
��4:� ���� ��s'
 ��#a��5�Z�b�ۡ
J��Pr� ,�BxK	Cq�.�;�r,�Ć ��S��cے I�-�k ��R@�[�XS�g�-���\�&Ju| 9�	})�x �P�Q�l����1Ҡ�� ��l[- �X���+� W��0�N|v*=}H&C��")� ��fB�� �:4��R����G2�y� @yI1�ËO ��ЃJx�F�~�� ���;�`;tT
��H� u]Ax���:�E��`1�� H���#�x�o3u�N�&�	�w�U׋� p�A�0B9�(�n��2$�z� �9�|�.� t�P�,$ �����]� ��)���>C�Y ��[��BA<(����=���� �����Ar��)�<
$C�1���j ��Y^�8�
��M�X1t �K�[-� ə��4P �B2AXL�٩�����;� 迈���S ���*��� �QRN��� bj�!`BP �#���Ӕ (Z"|.� �BS���D�L����:|'� ��$�� �.y�O��� 'J��rݤ��FkP� ���
|��F�X�b���f�@����X� �̠�H
"��ې��?@'�Rxp}f-j/P 	a�(�$�6 ���RU �ՋT.
�, \��YJ���T;� �5=IqY��P�]��Cʰ PD��� ��8E�$� ��(�J�  �/�%���Y�2�B<!F_Ip@�z
i wB듈� +��nX��Fy- _���Ptz<�H<=3�Ǵr�a[ \��!�8 ��+�>�.'�=�ʀ�|t�o����Q�)�~���G�.� �v��i=����=���I���eU� _����~�>� �]�X�O��K� ��} Bc-!l��W3� �[�FB� _��	��L;$�\d  �0X�;�b 1Q‐� /�R"[?>,�N, �8���K M�d"Y��
�����9�G�$�πl�� ���C�RDa "}�
#��|A M�%�,��u	��e1�Y� �z%� 4��(�f��O�Q ���w��&7B���EtS� I�G9F��:��((�f�Z4 A�c
)E�$��7���q ���u�� a��!W��s�E�� nǫ��ͣ�UêZ@/�J&.�!K��$*�g�	�+T�}ΨjX {O%(l���x1)�#R	P=��+ �w��PbV3z5q �W��	Z�/dQ�S P�7c���
��U�q�lh �(�� ������u(���r# ���tn �u�%�C�� �|`�&���竦���� :f�8�*PRԁ �֖��� '@���H�LN�1�Z X�`:�s� ��;��VH A�Ùp: �~u'� 3X��w �	�9R�-�u�ī���	X?�*����4��' r�}�Q�* "^Yh1؍. E�k�,!T DM-B��/) U+���w4�  j[Q8� ^��JX��DЬ�Q��U� �Մ��d# �qsT-�\�L �3L�,� ���_�xQ oʴ��h�:V���"��v Z�d� ?2��
�SC �0�4J�q} V'W�Q�S iN]�+ɘD	��$� \Q��a=2\lf���%:{�4؄Q�Z2� �M'1i:Ī�w�6S@\CJ �٨;�uo ��02�Z6�Y=��L���K5)# U�T ���!vI-�� ��'��_Fa3^�S�i�̩�v�v�\BI+ Ac���� �L��NF@6�[e� �HD�4 ���L�_%g��	�5��5�t����k[�
;y ��L$�PY��D`��p�  Q�3� ��k�ZP��Δ�'�#O�4� ��2T�|� ���X�H���] ����8�0�|} �K�&�9z �I�v	�h8 �e�� bic�l( �HFD?��a ��}�lc80 ��3\�Y� m��|乊� ��;<�>�LWb	$��H�5� ]�{zIP�K�,@����U �M�+� ��� Z��U ^�%W�����;K����؀WHin �|���
�* �V�C^c�� 3���H�� jP.�c� �ǭ�m� U���X� &��N$4çL1Q�;& �+��P�} =���T`z� �(~.�Hs� I$O7|"G�J@�L����e��� �� O ub�ˉ�T�!��������@ �E3�X\e I�D݉���T
�t�3�Gl4v�� �܄�X� �Cs�I,Z3�K~�j�� �Č�Z|X%[ ڕ�_  (��j��\ P��|�,.ѷ kR-V�`�0߹� 0�H�;B�
 �� u���>� ���;�"%��u�\a���İ ������� h�iJ���3�t�A��ya�Lpq< �CS�t,] �l���wPm ӹU�R�� 0�CE��: ����8�΃xA�íR`��;9�2��� ꉍ�j�� T�M�H�\� �+u	��� ]�h�`(dEy�9 �ǵ���
�B����| ��@PS!3�I5����\H��Et����g���!���G ��,:V��@=�NH	Ƅ5��W�CAL9�@�7`�^�: ǀ_��*d ���ker n0l32.ud~� �>G�tLon gPa�q��m �AD���B�I��}��pR���E�� �~�� �/�L@
+�Pt���>%ur"��K�$��p�>ā�y�)o	�O* dŷ��s#X !K�Ch�i�=^�����x���ͫ$@C�j ̔��+�&�W�� -!H
���}������� -#mH�R'P� Ku,. )%���`
tmC�=��QJ�SuG�s�3�ހFi��V&����j $rI���Softwa�e�\���c���s�ؾ �Lx�#�Z �l�D���58��	�9��MB�'`�TL "-��
� �!�oΰ9u ǟ�A�8LV ���xQ�� �Y�BM�������<&ӈ�A�;t�P(��E �����Kt	A;U� �(ԕ�<�-����? �l�'�[� �t=�{ >}*�FƋC 	bx�d{ ����
����(��O3�N�~H�%�q�����Q�Y ��=�? �x|��4/�H�ki����R�t��D\J5Y] �����$�����V��@�k��N�ZQ� �3��YH 4�k�,�q]?���[ �uRv ��DL�2F^�-���9H� �. �e_���K� �i��:@�� FtN�.�'#��)`� X$І" �(���N���@�QXR�F�T����< 눉
�~ ������ N��P�6�{t2D�#-��s���	P09�����9�5 Da���_�t	 6GZ{� �n�SL�� BA[@q,!b�+�J��+�H�*�]�"��U�`��X?j�^��V��0�; �ȱ��ok L~a6u R��,�^i��|H$�ĸ�A�� .�&�"��� )���$� I�;�z�~�$�� q�����`L$fz� b����� }���
	�̀�(U,h؀��1S� dj� �a ��g���+��%F��Xء*�P D��w T���SJ$����,�&H�W��?Z�� ��x�%�u ��;��s��9������� B5���ä3� �hTF�b��B�A�t� ��P�v)X Lr��� �@��f� X�R|BK��Z�
��ML��C����� ��HТJ\&� �K+�� | �(B<�tX���z��J f+0�FwY[�����OR�7 ���b�)��}�i�t���T�� 6=�@uV� $
�0'� Ki�TlD� ��v�sB� \
��P���^ �VT�Ji* �+�fv�� o;����~�B�%�j��Gf �=u.�> Q�p�+�E �G�����_3�X� ��z�"n= U'u[R�T ��X)ZYI�t���w���q����`@����~!A 鐓Q��& Z��GK�u [ս̏`��s^3��D(,�"�=�+�~�W� ���Z!��[H�kཊ~T� ��R�ۉ| E;�}	 `����ՄӀ'Z
��Ÿ��J�!@���� X`6�QU�ztp �Vl*Z�� ��LH�-�;�� \���I ;Z+H�[� ����7)�}��1�`mE =DՍW ������ �,U�T@�� ��
�x�$ =�*V>a���"�E��� ��QH}B^D  ���ๅ;1��,��z�7-�es ���
A��;\�?��@� �(�Gw# ��P�p$����� �� ��`(k���������C�#�P��� B�*焑Jp �� �-�
�1 �_�0@��!�4�(���7��v:k!�D�= J#Ǌ> b��7x�Arz �&��@D� �n2x��H� W
?h�K� �����N ����aQY �R�ȥ�t� o�U�: �'���X؄	��x9�?�\���6=����_`�Ng��r�zb�܁E �|o�e螵 p+��ŝi�� ���Ix�&��� �����p= A����H���L���+���&BkX 9��p�|@0�<����R��I������~RQC �/j\�& һ@v���)� |�}D
�� '��o@� �������Y��� ��dE �����Jz���b��܀�>� 9FǑ�� ���u 9���v�HM䧓> ;5���S� ]=����� �Z�� �T��7a����%8]� ��g��'��{� ݀n�� ���R `�%u�Y�� b5��{� ?�Ә��N��� �o�	8ќL� )#VJU� ��'\X�tL �uC��� ��FX	y
���� �N��4�9ـۺA���� Z�-�u��� r�t�v��=;� w���+��@`��[� È�tSFK�����3��BV���#���� u���y�(�[�{�  ����7�Oe��W9�����/�%�!�Ћ� �{��d]HY VGb�J���k�r������sN �X�n"3A/ Չ
��V�r� � |8�X05 ��p��b8����*���w ���:̙ �f�8�H��v�`}~�Y�9�԰K�
 Z�:�$�E '7�5q,%� Ħ
�wb	 D+R����X(셙qx��B`�]h��<,�������0�z�{2 <!�B��bD`f��� l���B� 	�G
�(����=���pZ)�_��� ڍW���8ˀ�N��i" ��[=;qW&�R� ����,G �2 zP(
gXDU ���#[I L�x�B�dr9Q�`�! �Sg�� �=U���}
 2��%�w� hj@�K���J�>�S �1?P07=� ����XO�2 �/��"N Tuj?1(QLw|S�"/� y��)(� ���-G*'L�� �� �0�({d5,m�Â�Vn4�[�@"���s �/�SQ:��2 b�Ԥ4R�&	Q �P��A0$� ����� �	�O=Zni{%�ż�~^ u�9�P'�� �Mw�
S;O ��D��A�GL��5ذ�P� NWZ$��2� ]84܊e	�A�L`�!�=H�$ @��<289 4#0�,�(�$|F������r�9����l�;��e�R�9��D�����r�;�L960�"�#�L�� ��r�9�0�"�#� ��Ȅ�r|9xtp#�h �d�`r\9X0T"P#L �H��b98���P9LH�D# @�<�8�4r 09,(�C$�������`��Т_�>���]�͟�ܗ��XNEkn׈�sp� {�c+��P `���hxBv�y wj����|�T���1���#0D� ����r�9������*�#����@%r� 9��!�Q�����2ș�0�B�#�H����r�;נ�9� � �#ّ�����9�� �#��� ����r�9� ��#H�Su ���r�9�H�A����ȳ,䴸9�� "�#���Ȼ �r�9����# ���ȣ�r �)���b��/:�8�Bc��N�\s���o�>����\)$>�;����2D�:	�Excep�O���{lP  ���h�# ؜�EHeap\[�+ d�� �Bx�E Out`fMem o'ryA�|^���� ��" �EI<n��8r��{Xt!ސf�^t��al��V+X�,eÒ��B�8lѯ`��;�	)2���#��x� p
EDivByZ��o�<f�X��
�6RangCe �Xs�.�M (Ov�	flo �t�{\#褸� $M�L���Hg�� ֤ft��v0 idOp�����Ñ�$������?��x aI�(h^��X@� �UnRdY?��9쀎��tH` �Po�͓��z\ �0~V��:C�stJp`���@�E�o����W�\��)� �@EAc��?qs�V�la%�.D�; ~k@,B Prhyle��+�t�s$�LS	@ack���$�\ٝ��DpHtk;9l�(���@�}	Var��+��B� ��Ȃ�eߐ�Fa�oId�+`4��nb� rBs���@Wl\��@���f�9��G��@��(a e�´qp��v R�$��ֽ'�� ��f���] v��� �^�x��\,� P�胻Z�O!/Y ij�w� s�#�BmSN ,�ߋ^��	wzM��U���= 4Ig��e� ���Y]?� �N�8�O)3 ������� 7+���L <I:zw , ��BFK� *u���R�< �A ZB�v [S��	��{ ���R���9�v��װ�� t*�^���qi
�_��r ?��r��8� t�����)�[���$�J��P!+�@� #	j^WO� kM�D�Q�� �@z�<�� �𻉲.�� ;�|�` � v��}
 ��?̔dN *7L�l�+ �A�gsW�� DZ]�j	&5�O �S�� ��n@�ۥ�V '��dD%vK ��if�� �ƃ��M,��x �1�]�
�4 �(b��)�T=d� $�ǆ�<uU�;�i"`� .*Kx�L�? :E�����w �|Yy�� ^@N�L$�i�vO�C�Q��I=�\�0֬� ��6�Ѕ���� C�b�L`} Qj�r7�5d�Z���1� ��?0%� ����� L1�P&��$ =��@G�; {M�,Q� $j��Z�;�%�N�����R� n|�Z�2�� ,����cKHȹ'� @|��e� 	�Q�JM� p24�%�Bu�]D��Ȣ ,��3e��  �@�M�p�*�i~(�V�0�`�@����������v ���`(	�-\>�M0ԃ��cGR��� �`�<uNO�3 ������ ,�"��pq D��`L�&� O��:��+���(�pe�4�����Kb5�aU�Ih	��`������ R��"�N�$��� >���m~K �f��g3��>�8�v�0�A�M�j�>1�L����O���}����=�I ��0{���� �)ȉg
� �;7�4�ʿ ��t+��IU������"���;!� ��< �Jn4�?�.ɫ ��睛ʙ�D���^k_|Q
ԣ�K� S�Tu A)��-��Z�xg����{ ��5�w� ����YD�b��M�SƠ#1? �J�"$�Fy 'X@�;�W��	�� ����!Q�e|��2 *�S�D� +��WP\� �_�I�cp� u.�H�h}AD(�%@܄0FT -+It.�� �߸)�1v �^�A� $'�Ȑ�Pَ_�����G���9 3�K�Z�(&�������`�����4G
!� ��>zĬ����p�} ���v� &�B�J�/��K~p0���3Ab/�t� H ��¼ ��`1�� ˜(�<���o�6��*�'�& 3�%T�� -�]z*�s`	� �}��Je��H!U�����t�%H?<�?+� Pt�1���L�]��E�-u` 1ڬ�}^e��:�
�4�����b��=DW8.�2)��&9p*� u�QR��4 Z�J��s@V ۀ3}�
���ю ��� ��T3���E�
R� ��dƇY��6���*t"	
0 r��9w7k{�`8�t���À0�f�X� �S��n;`� w5���| C�:&�t� �Oܬ�$߈ �\�w��9;<�R� u��4�	���N$��� ��v"6 9Mw�xf}�	?D� Cv��!��� I\�d�J R}�x��U�^M�)��#� ��]	f� ���S���D _t��U�*
Xuй��#�C�0��t��pH�[��0 �f"�-A	N ��]C�u�� ̋�뀒I:Y WBR�=:r���)N>�H'���	 �uʍM�� ������v B9Cx�
� 0L�?�ҏ!"	��=*� ���ay� 
��g�TJ ��͔{�X2u���=S����� "�+^�%�	@��{� ���B1ɤ!	E�pM����5��8w �~�9 R�;q� �j_]�� �|4	�t� ���;M�_w ���PC`Y *\0d)�7?O(���_AP @��E���# ���$8fn���Gt?��Ew�� F��N��MNA�����s�9�v%�-�b�u ����d�c ���-�� �)��SP�����|� ��O�!b� �P���t�x� u,x�%~ �o���)�c-bQ"`�H΁9׃.�dgD �es|2iQ�$	���1�h݀�N)�I�� d��C���� ��=EO 2��:�� +�;�}$�P�� uMn� 5��E{� u@���8;P�0 /�sk5� �SK���UG9-}v����?��c�u��t 2�JS�	 -��C<�3 �#M��� U�R0(@S�\\�� b�U���=��V��k�ɡ� �,$j�qP;�� ݩ	�hB�we~�`%tm��5l��� 
�S��6=��$`�� �]V|�E� ��=�sM �v<@G��A�`l� z�:��ri ��63��% `���@\� �j��
P� `��5�z� H�1����@^�ƀ� �LpI�%W�	&�� k{(f� y�'���� !OBju� >�H7��T�k"��\p�p0{ �F���_&��� eM-���,u� 5H�UR�>���u� �ҳ
�� E!<�fd�'�� ��.�B��\ 9�0�4���=Z��!١�� 5.E����� ���¹�T �to�4[� ^�X��Ll��f��K���2�v�k�� ��@g4 ��+�H�}�`h���!���'w~& argx���3� l?�ǁ;\F� ��H� ~0�f\�N?�A u�P,�I) �������i�m?�X #�q�+��@��`���b��
���5u��$ �Q�K\Hi?)`���|RG��!k��0}�"<��h��)� ��$D���P������� �^��Y�S !��z��4 Dn%�2^�I@����:| �'� !q`k�2 }��R�	�� ��4��� u
��M�: �.�k>d t\خ�7 x���-��s� �^H�RK �,�P]�#m�9�O?t Ȋ�LJ��]�� �;�r��	�@ ��^z38  �m�&� �L���DQ���K4%`�T @�m,^�k� ���g�8+ ���.$�� @3�'J�V �P
�M�GL<������+�$e l(����6P !=�迩���� ���� !m�
�TLa${ˎ�S�����+��vӓ �	�X�� ��FC ������>*�L��K ��S�[Z�(t� �@nYt� �x��!&j 1��a��l U?藵��`(@p1bC� �r��f� �H��FS�& �����={H��	��:K�tQ ��!;P��B��x�W���u*�>@_��a �H�AP�R L�n0�� @�jt8�� 1�X�P? !��ɵW�7k2��)Ə��@pTV\� ��a�MJ<�� ���B���r� sf��t��D����PY1��m�,0bh.�A���`3lXD�V�;nN OM��T���p�� +��f#)�N0��3���,EC ���#	<�{W���p@q Ȭ�#��^ F=�aui T0��G�\�[?�o��3;��.� N�]pq%��D Y�j� -c}��' <��E��P��� [��?xd�:%ga�@�oHuS �8f�F��� ��$|�k�����)#z�tH3v�u�$ �80�S�A�I 6c� b���\V� ��yg�D� ��I� ҉��ܫ� V 	B��� }����F
��5������O��E��~ ,��A��~��L������  ��Y�s�}���`A�r-iO������ Zs���@ <Mu|:�H��N��J�5 �98�C?���� ������� -����3��0j\P�:,B	 
Ɖz��� X��"�y �������QH����MPi�	 y&U�o2Y�V���#$�� J��z�����?(_��n #+�J Oҏ&i�	�=Ȑ p��?z.-!d �qo���XH� ��t� 0��K�����,����G�@@y��u^%�
t�� , g�y�{)w� kSJa/�o�U��u��!� p��bD)�r 6G��,Ep0���Lu��j�{l� @F�>M��'��|��}Ht{:���c 
u	@^#�3�_ q�>
�` S�}�uML�d C�w�+�Q�*� ���B$:# u�J�X �4و
 F�����i�;��g7p�Q�>���
|�g�:a ��4�~�z�@PUR��ml� �|S�0�`� �g̀��� 1�)�b{	U�� �E�� X��yf� C��T�*I� N"l�u(h� �r]*@,�)'�߃pa�a*zH �z�=C#t�9"��4��s��`2���\��l� �,���4:����\D�Kʕ��� �����qĨ ��Z�`����K� .0��D �5I��Ÿ8T�O����( �DC��u� �X�_%��f��bJYĊtxuE �"�:��u� ��U��R8�8�*�D� ��5> �l:�?� ��f䊄PJ��'8k��AM /P�x;� ���%  \@��4�w 
���e�.�Q F�& � ͸��'.�7 �M���1y ���C\� �!�#�7zj?ppE�B3 ҺU9P{��;� j� @t��w( �v��[;�%=��ǿ��W�(3 ���~�� a�ȊT>��0C�dȺ�=( �D2�, 
s��`$� ͉�;~�w�O*\^���+u���:�0���pZU�� ��k��$�� ��4��B :�֓��\ 	EǦYyQ iVf��-,�^ Ce0!� �2	��"�,�o�-���`ܗ��6��F �N�|��`�R�:$ uϷ���xZ �)��e���x� F>�$�,� t���
�wc����g:� 3	LR� ox�G`Y�~��߈_��$�1kY4;B��V5i|�Ձe���� =� ��H1���75�� ��})��	�l�T �Z�b%\YQ ��d�	�Os�!�u����,�Q�p��C u:��c $��Rw�=*  1��39�+� ��:0�k ���؇9�xK���X ���H 3�����l �I��2� �	䫞��!\�N ���E�] �A�0I� �CF�a�S;|m %�޸J� -gu4��z ��7�s�I ��,	&�U�J^`c۵ MyŤ���a �����"	 ~�@d=� �n*�W �z�q�1a �ӊ)b/>|�^D��������� N����h; �,�rE"I M:w���}�(�&�>�� _�Y�� ��6�Cmz# ����A�@	&�j+ �� �,��Uv�&=� ��p�� �-�j踵	 �,�[� f+��HQ�yY�L p����v<� v�~5w"�u/6!����p8J�R� ��'���{�=t� ݙ&�!� �+L0��y:�>, d���l �%��1 	yuu� {�tӳ��:>T�;N�e��Y�,BU�� �[2t*T�x��ቡ �u�� ;N�U� ��H�.��9X����d*J(	$��/ �e�� 	Dd׀NbT����a���\�%��"����{?#!�&���@x(tX ��*)! Y���8.��	�]�Fx�r=��4���"wE ��6�]֐��IXI���4�
� �n���>�b 1�������}S��$ f��FP,w> u�<A�,��Z|��
P
������O[����%]�@⇄`kP y費�� /̍�Uo*} �d���;A |���!P7b�0�@���ǀ| �6��䡏 �	$� �� �T)A�|:�u���n�"��	�@p�:)����ip ����r��#�ͥ d�1�( [~�h�����m��	���� ��M�~:ҙ�{1�``; "�G��r_� X��j��  A�£�x{ /^��Ҵ�M�?	���&�� �A�j�$E��'v��Ӊ� �od7l�yNQ� �D4�);$�������M ��DUjtK �F�>t1_����DH���Y:�� �M�R#� �(8���T��C�؞@1��u� �at��-^ n෌X� ���2P=���N+�q�K��>�!*O�CM>錀�l�su ��E�c��ğ��1�� �~t�%<��\_A@gV
 �OȻ��'mz&�j��Y���)�L! ,�"���� H�����_ 
����� ᠖�v/Y ��wC� �aHP�ƹX )-��=f �ףQn�H�<9�#��
�j �0�Ph��~ ِM�S� =�.�\lV�) u�ja)4�K����o�z�$(�� Äˈ_e �!��
H/=֮�[8�4D�	�j �`���=Z ο&�l30� ���en� 5�#�D �,GN� ����T���(��W)%�>�~����I�g�U ��6kX$!� ٌ8��� MiՃK��?m� �5�wR)��1L�D�3x��~$�H <�X
a��V�`ON�lq0L`Y t2u7xT���� �B��K�� %���� 7�4�qg�|�|���`��e� Zά*�=�����-�0�����5��:����uअ� �$T$�N����/u�?[�������!%��q�#rUL�"�Nw9� ����Q��(+�y3�\'@�@��c� E�B ��H�"��/l �(�r�	��B�sYp�!s� F�\�صS b�K�'�,.�,oq/���H&8�] @�%�u�[Oo����(� -���g��+8<2& ��}K� Ҹ��O���HğԽ�d�"��Jx��7�� �Ϭ���ht�j�I qvJ�.	A���9L�$D� !4��7*\@-ST$`B�6�G'�%��@�j������O�h��U��H עacO�n@ӗ2h�ǧ��� a�Gg�L��ۮ*�i0Y�Ej :A\rɜG, �1nMdǝD�m���{< �%J�.�S~ �Yt|ʀ+� y�O����s�=V� ����;+�b���b�T�,f ��i��|�	T��kRec ���UY� 3��;-+Nt� ��	�4 �2�u� �?"�����^ R���4-$ ƥ�T�� �6J?� �pYZF�0h�&
� �ť��S�) �Jtg` ��r�#9����!@�D�w �,���Zc ǒ}����- S�yד��)�D ȼ2��t/X d��'��9{� ��ߐs%�� �,o�	�x:F�v��~  }�I���tP�U�+8�M j��k�L��,� B�%��mF>	�Q`�H��8}�
�����a�c�Ѓ��� -op��<l� '�W��h Ȍ#�k�� F!j����� ��S�Ub<O���4� 7�GQ5(� �/�%^ ����Û� @��	��  H�L�:/� yI����� �B�Z�
9���iO��ء��|HXt �{���dG8I���Xs 'jD�:C K1&}�-#��t��Y�H�?�� ���df��R�Hh����Е.?�J�o)`��H� 5a#r���:�I�������'ص�,� WdB�Ȋbٖ�-Q�XpLiH��Z������T\�� �!�����
q� 8N��ˤ"�Q ��d����\?c�߷Ջg� �����U�c�r��L���� ��X��'a �d�
,s" �^��;U�[� Y�0��*��t���T �`6����B dҠ]�� �Y?��_,��Z���q������5� ��H� �B��"l����cw�.��MB(ء� 7�b!\hD�_�l�p��� �Vb��� �P�����,L�� *,#T7 9��\���� �K�>ZԷ�=�� @W	�&� r��+��(�� �"549�%�B����
!�E�r72°��l:�� ��B�T� K�a�X��� �0C�T�	 �(���� F���R;���;ni��� �2�ėf� <�z`�����M֒L�n�H�uN ߘ��|� 0��  r�fc,�&@� yI����l\�� ���v[ 8�F`���_ ^�� �'�sg t�C��J �6����3� �T��)�<I{���.	���1�o���\ O"���~; �<�V�X>&%�mB�,|@��+ ���@ F4}��pEu% '��K�AS��M����L$ �!ڋHxit�> h|�2u �'��: �Y���4�s� ^��!�R�J�bY?>�6~7��.T� (�!п� /K;P�+�7 z�CD���� |)i�:�d�F��	���h &MgJ`}ʉ����3��9N{�l\�R[��H.f� Ђ�+� Gi�uϼ���0{ ���U� bt|��Gx �}K�rT�� ���W
|`��+�c��?���ַ l;Y�#'�� tn�V�� �P��(*' �a^C�#�� �����+�� ���;�v�8�.����5�� ��Ԗ��(���@��D�yI��S� `ewW��U���K�[�fta0�G�!I�bu �W�(��� ;��l�����ȉ	���F�⏑�~�;�}�af܋�9�i���V+�b�h�z�YNj _KOq��9߈ 	�*��� ^E�@U�4�AM ��D5�r\ *�rC��d�9�я���@�%u�p���O
*G���B� ��Y�m�JA?�I��S)��� ��7��~-� ��k/G�� �eǯ�P�~�Yߥ�}��DC�G'	�ױ ��K"i*� ���S�H�Q�Di��j �-��$��A �,�Hk���L� { C��J��n��G
"�6�� 7Y�܁�����W� ����� �B�#]F�ZG�x!� �@�:��m��E���(�U��W�b �P")����8��S�<�2ȹG%#c�J�w"�: ��4�V,e�2?#nCΈ�:Ӄ���� b��8���ZH��� ��hX!� ���N�W�*#d� Ւ�% �E��q�U�O��S��^�:�%m?/d��PX�� �,���"a�G pPLh�$�}�D ��U����{8� :�΄��s�S��]z��) ���/~BkX��
븄h� @]N��9�5�!��$#-� <ҋQ=�Z 
��q@In V��.�Di skFr��Sp a~cExA�$?���<��04" 𥎨��6 H�4f�!�p���V�d��Hș�1�$ �L8!�=�D �&`E��$$�� ��,8" �D ��Lx&�A�p��h�T1`<"#Xd�PHG�?`4D@����d��LtQ(�̑@ 2<1&�aD�}�M�)C d6�"# �7�1�LH����:�:�<t �J<a�y���L��1)${� #l���C�"0��\ԉ��4Я�G<̦�Pȭc�0��T?�.Ћ��@��J�>g$���8���GD�(W$P�8���0��h�T�����C9��!N�:"|7�4�Gxd�`�t@��� �����<Q
 �	�Ӟ��'�S �p0?I9N F:A[\&� ��E��y{�J<�T�e}���z̰~ ��XHP� ���}rN �`�舤?	���ń-��0s���0 ���I�N�8����#�u��]� �t�w	�0��� ����Xn�VE��ϙ�: ̲%d��r� �
�u0J� `á��!� -�Umd�M��;� �� �|y�eN���@S�^����  ��o��BǑt�����Q#f�`�?(H�*�X�/3�R �+�b�� �%#)�*�I Ƈ�+a �r�Z�E �]��U�J �
�u� ���}���?��� 䀱�Ī� P��2�5I�_�ςC ���@ ���*�>; ��Xs��b��r��V� oI���(3H��{��� H��� �C��It Ku��=|�2��J����	1?s�Ap�'+�&�Î��]`^2� FRd"�!p :�v��� �	��V�� ��<�t;,QS )=(*�� ��'?��= ��[YC�ܮ�\5� /��*\N|r^�$=� �m� �u�(��)�-}�GjH��5���.?Q8� ���lgX3 )�u5�Б@��^ٽ�ubi T��G� ��OP����L�~*�� O�(�W �L�-��� �6�%�Y���rL�J /ұK�� 3�f}N�=	�Jt����@��u  �R~K9ޗix�o3�� ��! 4�^�����t�;�� ��w�g�~��p� u��<':�$�" & ��0V���2��E�@�`��:z �Y�
����2�������fP�����U�0 �#t&�9%�.@,���3"�5|1'EG:`eo6� �F���@B �����y��'�� Uwc `���" q���-� =+��|�p����X�kJP"�x��+���N�z���9�f�E[� �*!��)�u ����� �!�bV�+ t2�܀؅ ���c�]�_ �(����� ��E'�$�H�"D� �S�O������&ͬ �n�+�?�&&����
-u0�� �y;A�e ������ S���Tύ�t�3[.��e�
 �،	|�� C�>�M�u� �wE{�4���~�A`p��*Kg��1�f�"rl������ `$E�U~ ����% u����I& �d^6�8K ��`��cm��,.��F� �H%��
=p�"f�F��4�> 	�J~�h�@��C�����.�[p? i����� �@���J�>����K��w��� -خ��I�� �����A t	�s�P����Luz{���k��D��#��%�f 0h�b	�L2|��`�y*� ��;�,<` 
��s����5�%�D�Ox ��9w� �fǦ(1 b�_R��S%�!��P�V�w: 0��։�LSf �j��. ����k �i��y��~a �����z `�|����-d(� ڳ��s� I!�$	�x��m�׸�*+�@y�4܅� ���Z�� ����!� :���$u �I`��9�� 0� �Z� "�!d1D��捰�X��Ѐ? �*������������W�H��E�Aћ�`��=�� -�W���� 2���>��a��
�FՆ,�=�:�:�f` +F�@;� 1tJ,$�a p�FR�Y+��U�C8$ Z�'��	�\|� �jP��v> �?���� �f��L�.p�\	* ���Qm�6�ì2�p��&N�� �,:�
s �L)��� �pS�&����:�Q��*��k�ځ�@��8� r�(��	\߸\�ˇ �3�?U �F	��<J?�ϒ)D2� N�d�gz�"��!�.�� m�J�?�jE��K8�t�BD#�:y��s \
����D !�d�, �B0��RV P͸�Y�x8 ���E�s@�*F]�$�1�% �=��˄ 3��iLlqvp ��;s� ���r�?�U �<�� 0x�"��u�8JF��|\��x�"�C��\W�+�� &]�`r\N:�M�1 ���(Њ�<������ �s5Aq,�� ���8d� a-�稭Y@=���9ض���0��S� 3��9��uM���k��Z��v\cdO�)�� ���uN��f@�7�&zK ��;�wZ! �����s�|$����' ��QM%P�) �!br�y0 �Nu�����@zJ._� o��c)��W�/��+��eU�ڍ*�� �{��Y�7 '�C��K ���{w�U��PɅ�v�<�3 ��p]�@� r'���q>�րtP�������2��) 8��/�Hud�P��Q�mv T��}B�{ )W�����Ǵi�q�&�p�*!�I �X�үJ@ �=%�r ��SV�'��ܬ�J��m��x PUȊ��-� Bm�4V� �1�yJù lՊaC GF~���pu �"��A	�LR� ^:H>2� ����C$�1j=��G@Ku� �f2c�9� �b�O�� :��ñ��� "5��qHNv�X�/���:��|}%���/L�7A���̕�� zU�
�� �]H�V�P�0<*����.�$j!��<� ��2*��u��4��7��,�� �b>����M�ˀߜ|����q ٨؆� �W�R��� �;\Z��� L(�t��`:�7��R'� V�K<�%_t�r@����'Y*/����z ;W����1 �}���'F� y�q?�f B%�v�� ��b8�}o �!����mD{��8"���_� 35��� }��E�� e¬S���V�|�@C�v� ��^9;!� �ѳ�',��0��%:)�����=�W�/|`�K�" P*�ǥ���T��|��b��d�b݋u@Fwf<H���s[�9~u ���ތ� يK���l �@oIuf"�� ME�F�Ļ� ��)I�;B�vݪ�j�Mu'E����o���`6鹪�0�T Z��D��Ƥ ��d V�G�R���|P\��ZTg.@�x '}��E� �X�|�� ��yk�@t�+�1l������j 6��M�;��c�XB��� �PŒ4�t]O0J�9r$0r��p���Ϸ@��z��~��#M�;����/�`Y5��£� (C`�� &��\!r� �L�vdz�q^ ��S|��k %yO��u0j ��eR �,Y�'��PTF���q�.�� K��Q`�r� �1�I�S ��ڬ0Ȉ鼇��f� ��sx	58 � ����� u�1�G�Op�[�ҝ`W}�K$��� 	�a��Y� �X.��%��J (�Z`.V׉qFp��+�� �W߀T�� �|���	 P�D��+8T��,�N����$!��w��;� �G��J�)�f� � �	�ȗ� /��+,J� r�VX�(��`&:����F B�=����^��DR�X���M ����� �������|�g������A�3�>��R
D ���6� �F_�u� K�!ڧ֑^ �� �I��� �z1dk�Z [<|���p� q8�}���z� �����P�s4�D�n��q��_0>�@�� CID��+�� ��/}O�% 1�8v�N�� ���ͨ�*�=��u�Y�R �'�)\ ���[�"L� ��3�$� .�Cg�9~=p ů����T=4〡�/�X����@�	'���Ŏ2H�=,i�p,A (5P��%�\O&rJ����Ф# HY4��Q�wL (�[w�L�;��T=�����K	� �m'���� rNh�:��!���
 S�>}R�^���$��<��,��ʀsV��N5 �a�Թ��% m<ܤ��C ;���	g9 fJ���� r~��w�Y�v Dÿ��f ~ּ�p � @������} �ZBDt!z �Ā��(�� H�^L�~E�*�bH�r� KY��&�2�[�� ��=��׈ �1gE�A�����S4K��z�� �3�:�h�H�0 &Nre�� �)k�<���� A�P�{�c���p�Da�[ �&�x�%�� ��C�!�'�o�໪g $9D�-"7 �Ȥ���4;��� E�LQ� B���OM��G A2>�?� R4#�oѦ:,E�? ����P�����^,a�D0�I�S�;� +��>���oy(��PK} �X�$�HrQ�-��/!�!��� 
{k�	�a G�(W��u�phQ���0��$�P ι�`�’0�5N�)�����T�hEdt ��/�b�ɠ��B ן�8J���{Y-�}T���i�8���� ыϺ/P���.���ש S&�Fp ��]|��3�i�EB������� �C�xY���~� �G��
v�H� Kȣ+���x� F�Z]�4�W���d@˳�� ���ƺ|1� _�iu!�� q�;�{xNs��|�@a/�)o�k�Et�~�p`Ty0�L-ibq@@X*Su ���v�y�M��� 7p4� �����{����v�
�s�^?V�L&���w�l�N�j|йy ��@�CLS�� \+�=ѡH�t����p��I ,4��u{�*?�k#Rn�͸zG��䱹$(���#�Z �����p 0��or�����M��Jcu/� �Z��A�P �-T��s +k*C��� V2�aĔ� ���� ��I����� �.�9<:�,Y� k��� �	������ M��D�"#;�5u}� ����������=�Y �ۉ��qvT���!���"2]����	� ������7Q.�My$Y��Bo ���i�� ��K�~8?M#/�Ⱦ���6h\ g,�an*�0H� :N3�MB ����-��, ��>�#�E� ) ޡ�h� b�v��B� ;�O�r�1) ��G|e��BP��˒h��U�pF�� eM�xЊ �&��Z��S j�b'�q	��*��l 
�5Rtc�o�X�I�d���l�2 ��.$/�� �P�\�( C�#J�, �����؟s>��0r+� �n�}�I	u�������J3� ��(�O��!R68�)�F�ArT4C��%t<c ��>�P� 'Z�~�b�� V��Q�п,� 
��}-��P�=� �UD�.<��@��~"i� ,�L�W�=���N$uޚ`�� �Q�ZU�x��R�	z'�aCl�:�9��.V�e�u0�!��x �;}4�� H�|Ҏ���u��-�]�R���l� :���Y{�E  �}$L�6F ӳ�I�V���'�{�EXe����^@ (F3���%���H�S� ���
~<��$Gc��� %�̱=�	 0��o� <�.��:Ș� ���#��% �g�	S�� �B�*��� ���Ž ����jN� {²|�L8P ��"��oR�(��4³`��V�`�I�$��J� u����Yx�9Hס��T�- yǽ�f�i+]�^���LU�-�ަP-�}Rԋ��I{z��T���}Q�ӇYf:� DEu�t��ՎqN��Φ ���{�� �Ã�&"� ��U�lXZ e��&Ώ ���)ؤ�x��;E@v��$a��?���� ��U;!G�� �Aj����H��Z�qB i%�����W ���X��� ��<?tF�' "ksp��S �����W� H�_�mT�N ����y�(P��}E-��ף�݄��h�y�!Y���܋��I��"��vE� �gu�h�Nd:�G�Z�s� ˩&���9�p�غK��)�� �\�@ƃR�1�yo]�9&�+��r����8N��x��40:�ڀ&�_;(?��Ǡs�� ���'}F�~X �����mZɍt�Bg�2��x,؈�n����h$S�� 2����̐�ѐ�͖ �L�T�.� �$��2� ��j�N#}�ǣ=�p	�Ck�e��H� ���
g�P Cf#�u ��XAQ�>bN���K�� ��	�R�� w�ݏ���*F�q��R ���q� �"\���)������sl=mB���`�� M'\�vɁ�f�xt 	Q����=� Rִ(��h�U��\�
��+<�E@�� �\��P�� �'^���G� w(���.&�Y�@�;H _u	�ӰZX s=`��}� (�C+�� f�t�� ה� ���� ��]Q:rW BU<t��0� ����6��[d��@ɖ?�'M�(��T�f�����`rd2�wB s
�v��=�� !wOR�i���L�`�D� E*Q�Y��	��U .�ú5�:>]ĠZ*� ��k�gS �'��$�3(��	�� C0w��o��v1@���Ϳ! (�Z�k�Sq �F;�ri �eL�| 3+�DS�;�tZ�p���jL�J*d)��`7C �FHL	R4> ;�v��� +7�@�{�� :C���%L~� �ܗy�ᦛ �,Ge��`w�� �r.|(�ي�@Q 
�s "}��D�Ϊ�R�WД!����^���� N��)���B�X��VW>&1�`�M$� �E�e�� �ɡ&��<�+ �M7t�� �$F2�9���!tZ+�H<4uA3`n '��/_ ���T���<����!�U��`��MBy� �qF�� h<;0�	Zȇ���p�,� W5�!�ϩ 1i�C '�Y��P޸ Fu�H3���N��׀W��Kؑ�-���qP��������*x!��z^�10�@��2B )+���� '����|���8��7d l�q	�@�D�変�9 h)<M���TC ustomIni^F��������	��S�ϸ���+���g\���q ��	�T� 䔐�n�\�=
_ �t>�� ��-u��	 �C��� ��;ҍ /�yf='�~ �,CN�<��
r�u`S�����$co����]o�ؒ�Ƅ[_����򯉒]��0�j �67n���>� X����~ >�V��6 �a�?�}0	
xu&�.�� l_�mW�X0 ��x�6� 1gJКGtE�� z�#�/~ ����ȼ ��]_�}�^ |������ Srp�U �/젭\�( �@v��r��<�Z`�/�~$Qwy���i�S�� �Ȗ,��d�� �	�#���3N�
'��p�I�1�O��B�� ��]�<a� %�A"�_����`���y�:'����p���f ���+�Y����[��F�5� ;�#��!y���>�B�i=�{^:�Y�~?�t !1��F���{N���8Bܭg lʓ�Z�n��G,@zk�#��~R �0�`�� ���?��� 聜��o� A@�iZd�^�?�����F�<� `�����z�Y�]�ȝP<�}�U[.p�S�_ ���4�� (���J��� WM&<dN �
}�'%)� ݩ�����ZMQN �덅�z� ��r6���J)��e���+�/{Z _0�UmT �ܴ��D~� �$�%�	 ��ܚ`9�p ،�S(%� ��,A�~=e EB&�8�F�Q ��w2�J �GB���q����g�ΰ� ���'SM� ).�GƇ8� ����n� MZ�U� �z�,'BX� �c1��� :R��y�� �N���@� �uL�W� �BU٘*��>>9��bv
'^ x@��ف�>H�� �Q�����V �б�-��� �Xt'���$�����h�<�� a�nò��҄}¸� �)T=\�k� |
֫y8 fj-��@��ɦ��"�X� ��l�Z�Vn��|4[��q�� �x _��(#P��d�h��й�<(�B�� �� p�$�A�(������2�	,�0ଁuT �t^dȌ�p ���] �����	�w�u� 8��2�� �x(���> L��3D�?:\_�-`2Ap ��h1�?�� "tB�����0 A,<| �4>�(�@�F���1ͨ��3G��0	�`_XO~ RM6�+�l�?��G��i�.���CqESt��1"rs�g�� �L
�X�px=g�S�轟�0��� ���2��� �Iu=�[�8H��ˤ`���Z�S�ȉ�+�Kn��� 3�X�*	� ���Έ� ��~4Ge �7j�\再���DX'p�d�qH��L�!pP@T�\���,�հ l�: �������� ߗ����#��p� l�z���v g�:1��t�1��9ٍ�����۔ �3���X�/�8��;z�lߖ:� �7��sS �;Wt!���r��b�v1 �6��e S; qts� X���d�8 u�F(��$, j"�B0�!��r4 y���� 8� �B<��O�1��U� *���y�Z ��f�a9݌���j �)��� �CÊbR>�j )�	�?( �t��b�3j0'�� ��!�
��V~����rB<�1�.@�4�#$�mH�4s� ��B�}��VF�P�Y
 ����؉(L�! s8�B:�@?��
�R�<M���V�.��v G|h,赆C�!< L� =ǡ��n�3ې���R���� )�:��W��  	���0�4��+�;�<��Ѡ�b{5Ŕ8|B���Mg�F�������d}8a�
h����$p�ґ��`J(̵C��GC���! :�b_�,#�Bx
!��R @�� �3���r׸�9�* �|�,�$JH��ALr.P�?T@����i��� H�|�O�$/ �@�Y�� �H#Eg�L����P�� n�9Tv2 X����\��"�`_����d� ͫ@�hgE&#b -<3_���ٵЈJ��8C��?�D�9@� �~�o+� i�$�Ly�S�x �~�Qv�1������N�l���eS@X�� ��~�hNEW��4`��!�/ x�=~w�n� �?^�_�J5�t��;�}� ah.$~���O���d�V�@+�)�<j(��� F��A_t|�L�Pǰ�� ��}�M5�to\Q��� *�C�x��:?�$�D~���� ��|��3� -V�w!�4 �+��2H��� �?X�� �p $2i� �8L�����7����tz� y$�N��3�  @
|���~����4���)+� �*ƇGj �[�#I �F0�	!l��p�p��1sX� �ؘ�}i�2�B�`� �D���i�@(�8[��0��p,��\�)B���y0�">��kLS�]��C�a}��q������a�98��CyB��u�<�! =�I�����?� b%*�i!��)���
 @�%� i��5�x)� �J��QZ^& �$�O�� ��:i��ȶ�	�����D� ��@��v> ]/քg� <\G� (SD��6#{� �� ��S�LB�Ș����� �$��FJ���� ��!1�~�8�7�����������5� �� �ZEAX�.B��@��' �C���t&�z��!�� 
�H�)~L��og��@��0��L *�C��{�B9 ��,����g<h���\Ѕ�q<�!�*�2j	��+"a�m�I�еA`Δ8�� �	j��#�<& �xD�+�� �_�b��9 ���K�y���`����T?�p �����4��~#��������� '�ꃄ1� < L���0 �@�P�O����q�$�9 ���af�# ���@�����F���Q<�|�Ԙ�eV��� ���D"0 )�@�����n�@W��  ��*C����)<� E
,�8 ɧ#��iG Њ���X�p 9����
�B ���T����(U��Y[AeϽ|�� ���Q���Ѹ
��}���ΰ��9�]ᄅC�!�xy�O~�@o��G%x� <��,�TC��D������X�w�ע4 ��NZ�l�
�~S�_}�!�D,�5�	:��DТ���&�*� �yR0� ��ӆ�� ׋&3�na�z���mc�o�p��u�"{�E @.῔ZTx RX�|J�?h����r�q� �d��~*�H��4�>׮����,*� \��xB R+%���� �y���L���m?:ȻH ��}� ��L�r��+h�> #�T��%�����g\z+�����R�?�۽	Y���`��zl$�� !���	;ُ�F���� BOם#�8��(�!>�D=*�4=,�gT��ؿЅ�0���l�B��4 �15� 	�j;!<��{ H� �3�ǟ�l om.-�#��J�� ����
N�7!��ଁ B�'�l��� �7K4� R��@v���� �9{md� r.'�h��Ȅ�H(��  $�~!��x	�僎]��a��< �#g�� ٘L7��7��
�0  !����ɇ8G�)� t%��Q�	>�p �t����b��Mـ�7�<���Ed8+ 
!�� ˇ,�;�>��� <@�����'N��	x���������I�� \�$��Z�KO�,��1�5 �N��g<4�C��Ӑq�Q�<D!<����vw����%� 3�Ɋ��Y <
w̄�� d�ŵ,� ���W9��y�}�=�P,�<�O���CL͡#b��R?��u�!���5�<��B����� D4> |��,hNB�@�C8��#A�Ie5G ��B0�t�8����*�r �u��J$ <�����|��5랰 �����s�#��y.�z�7e�KE\�#�� y��[��-h�7ҎŘz<%:a��$�(��4t7 ��
���8� %�1$VG0��&
W���^ 7�n'鐾I�DB�� ����q��n,�C_O�b]<c��@HW�8�qF������z �?Ĵ�,�C�Ļ��9o��X{א� �����N �S]�o��".Hz|�?2�n`���q��t�;T3� �$�� غ�;n�3������� �7v!�e 13���n� L��:�0���~�G Kk8V��Z�Hb�?uȢ (���
O*6�@�8��#��I����[�(�}F �z�!�KA�j	 x�F��!s�� ,�����B!B�%4@w����d<(�F��?Nu8:�!G
Y�o��z^�$t�� \%�" /+�#���>�P1��)b O�
� 83����IGH��`1S?3	���4!�gT~��� ���N0�hj3i�/p�7.+ �B���-����\/���RqY̊���
��{.p�4���Is�y��� u~G<������b� �@��.�!��nt���� N*A�Hc* إ���0�-���&o�0x�F��'��75z���s �M\�H��	�؀�7�m� &�5Pه>W�Z�[�v�'�0�H����y�I�����	�[�4ׁGT$�� ���G�+3,�Cڈ&(�0~H8���B\�8�� �F# ��V�&�r��qp;N���Fϋ��2��<�]|��L^�D��+���xx� o����<b"�\�x��cpm!�)p/U ��3V��}�>�;�9��K��Ĩ?)�� 6���q`0��o֨3��KܞW�֣h�`G��(X�*��T��"�[�mg�ҟ$8%?ͼjp�����ѵ:����ѺhL6J����!�('�9BSW�ז�d�a�(�}/����Q�}|� �P�ޗ��Y4J0�߄%?wQ���zU �y|�v{����ow`æ�|����2��:{C ��'����v �oq�>?-�Z ��	1�� 4�n�K�d&�h7�,H�>i�Y� D<Bx�s�~ -��m��M n:8��H��C����xZ/\�X��D�f0�` Ҋ"�w�{��|i�nSt��� 4D)y,	 �������`� �� �	���o��S���W�b("�y���Њ6S�7�8z{����	Z�� ���_x� ���8�K ���5B�4�=3�w_�-[?� ����ܰϗ ���l
K �y�U����� ���� �����=Ó+�8�ˋa}PDC���Y���+���`�s�y=4^Y� ��8�H�=� �?�����X�>×����4�H�2V��W,��a\�<�L�&bL P>"� %�W�?RTK�3F���JP"XtB�=�K�`�� /c��pQX���%�{�	�� aSQ��1 ��=d�~<}�� -���6� �^@A��u�?�/�*J- ���Z��� t �Cf�v� @��rѪ$~� �S�����N� B��F@��H p�"5�WB����΄�
I`.=([�@4vNX�- �A���I9 .�S$]�3 �E���a4��~J�$� �c�� ��!�2*|4B�3�A��p�F�j&ެ� �[��� 0�I.���6wh���ΫV9Td��L�� ��Q4�t ��R8:�� �h�<z��`�N���#F��2�fB��P� =+��Y � �1�#(VC,�0�@�� 87�<j�@} �D�!H�FL �P�YT
�U ���X/���j��C�\2���Mw� �`�.��r���Yd�6_��9�h@.K�l5 dp>ܣvCx ��b�$U�����!j��]�b�����r��}�}2}� ��є��5 D�z���� �_A�d% |T5����{k�ߐ��s� H;���� �o�Dr#� �������VA��
j��C �n^�@� �h�+%����!��#�sV`�b��=|G��!>������̢ �FЭ1 �\�ԑ!�#;4�� ��w� ��Y����,�X�k�OB�.9�������x ˈ����J, �����b�w��5ҋ��t1���ڔ9��]W¥.��^kv?����!�F ��B�(,0�t F8�<�Q@�D5�	��ts�  P���XT=�f ,��/�H~�r�������?�1�XT+ ��u��� �2H�$ʯAt�`3���� �fǾ�*�/�� o��� 2	BIu�� ��0���
 �t&g�T#! S1ۊ0��P ��/3�]� +�X�_�[0 M�����~8	����A�/�<���`��C)�~ ���Apy�	�ρ��a
�����8����A���������ہ��v�ހ߀����8A��ԁ �@ ���A����� ��с�>��0��8p� 3���@2�6���7 ��5�4A��< ����@ =��?�>A���N:�;���9����@8
(� 2B)��+��*Au�w�y./� -���X8@V ��$�%A��'��f� @&	"����#��! A�נ�`�a��c� ���8@bH)9<�8� g��e�d8A� l����@Pm���o�nA��`.j�k� �i����@h�xø ��yP��{�zA���~�Ͽ�}�����@|��t� uA��w�����v9<r:�8� s��q�p���P����@Q ��S�RA��NV�W�U@	���@T� \�]A��_(����@^Z'�G� [��@YX?A����H�I� K�����J<rNL��pO��M�L�Ό D����@@E� �G�FA����B�C������1����R�@���^LX� 5&]P� 1Z��m������� KS�AL�� �a6�[�� �ZYݜdHi}��)�����|$�s =��#�O�� ����~� d\���BD`Ј뱤�� ��w8l�0 �4!���� 2��Ac0�V���f J�_��ƿ pxRVQ�� �$;���*M �0°� s`��� ����u�I	 ���~_Z �)�`XN� �,�]��E�C�Ҁ���U�a�������� ]\��U�;zsf�`� ;+�& F�%�\P
 r����3?H& Jƹe�s ���vj�� ފtҖ֯  W�u��w ���_ʕ 3z�UBp� =���G]� v��>� �<UeT�Wg J�8ыE� ̆�k�R�)�.A����q��2�a��`��ߌHGX�l �\E= J�ހ���# �I"���g uP��%� �\׆��8 J��н97� �YM�?UĀd�q�X�9����ʿ���\�\�F�9[������Ou;b٘X��to�!���JЈ%7\�@A*�?�R�� ���$	W��
(����,�p���0ȁ��4%�.  8�qy)�<��rK��w��j�S�X=}3A�c���V��!	0,�\����c��N�йV
� ��E�bo2��N$(HG�<"@D9(!�7�$��1�(�8�B* A#� R� 4!�;ӌ�@W�0A0	U �� $M%V�A�3 ���Bi ��� �)(�cI�ҫ&�b��`28��d�}� ��W�*�<�V{cr�J�ҩ�ΐ�?�A(,�`�%�if½�-@��Y}B�q��|0�f�̢<K[�P �ԫ $E��(^�YB ��:�1�b�[(
�<#/�e��]D!��$�P���_f�<���)�W鈄T�����UD��<���K@D�4*��$�����^� ,�Q�+���%�x�$@�D��� ^.��N �V��0ODh�<8(��رTN��X&�	�?�>�p�/<��j\$%!�tFU�6/�����I ��2i
�� ;'��8�� If�:N�3�����.� �� �� �����w2�����`� �+�������R�.� s
�p�5�`��W�<Z�#� ��Y�I> A
k"B}X *l��8 �W�(R���P�5����+9R�
� -���� �P>Yh[_�v��������� ��Ӣ��� Z.�N�h;�s+�V��� fx$-N91 �*r�&��y� �O� H�TB?��ɀh"�D��[��\�S����ׇ؞��܊w�-]�h��p32 ��0��"� �1���m�;�� RA���� Vf_/�K ���(�uYd�n� �!��� ;�r� u�Q,�O� 4��_Y�� щ�k�L��}�4��@���x ��'@A�9� �[�]��0 *홒@|� T��K�:�y���|�;�u ��:WeCNz' ��`\m�ǅ;z���� �C@�����D %��d~[� �}b�#��0L`� ��@5�� �,�)��� ���!4���.� �,s ��2�# �� �_�[X����Y U�F�7W3 )�5ې�A 9�t�BHe_�!���W�@�CDpE FGHIJKLM�N OPQRSTU��XY Zabcde8fg hijklmnpo pqrstuvw�xyz01234�56 789+/=	  $()�Z{},p;:-_ "'	4
���z�񸍨 �XB��}��ͽqO���6 ��	�-�t�r au�q��ob�O� Z�\�L� S-��;
�|��� 
nj��_��<�Luz�� �|a�$~� �;ӷ��~���}I	��g1x�B,*�D`;�M��^����Ѓ/(7-' ܻn� �V�{�k]�|�~XO�K���2�� Wp�G KHu�.f�LT�I ��C /�S�aQ?kLDU L�v'9�� �H��*�VƟ)�hk��~�YZ]���C A���%u�3�������i���J� �|B��pup����J�V�d[��/�lŝW�U�ȴD ��E�?�c� �F�4�0�;�(<�؏ <á`8 :���_ A�i���H7�/f��S���BhI���G�� ���RT�L ⋫w� �����Y(� ���U	�E����"1!� ��|� �qE�$� �ۂ���lF �ܞ �� f��=@�����- �^K��P�>�Z �9�,� �`���1߱ʠ���1e0���~wHh�,����-l�V�҄ ���%��`�68�wAFX 'c�N���a�h0T׎���pF)Y��� �vT ����G|}j	Vň��!���n:�Uϰ� ���CuZL{�3 �S�� q���'�&�dp �D"O^9� �M�UA�� ����W��l:��?XN\.aScs i���<:)> B�C���gK
,�MA�CvV�r��'ZQ!�h�p�� �a:t�=�� |c@DJ� �4̮��bi�G��@UJ�I0�q	 �g�XP.�� �k�E����85u��mM ��94��G #�NHT� .������@��)N{H�g���1 ���@�ZǶ-�q��D� k��'p$d �:\���� ���w�m�� ȥu�#�t�8Gf��C��;C�?�5���6܏ "�jL+���`,	�EL�@f� L �s4��<���� ˋ��|��(t � 9�8u�`C�&�8=K�W�]��YVd T 	�I�k%:> uq���z����W�J A"�(���H	 lz��!S�O ����I+� o�TDV	�y��cal�vr�e 0�TC:ʄ)J��4!��Q�3���� -�8��Eo� 	�C�X@<�\��:���r Ň��_�R ������ L�y�Zu�_�s �+����5`��N%?.��F �?�	��9�۩�x��E�u �	ࠊ�� Te��X�E� 5���0�� [�@�x�B K���~��b^� y(�� 	uQ~�/� �D]N�<�J���:��M�@�+� _PL�V.Z# j����X {�	�� l-�K(��t������,��B�L  ��;7u��bW9|  :���rt$��?0P8�^%$A<����[ �:�R1f? _��ֻ
� ��+7�Z�&�Wv��E �L?'\ %���H�� ��8!G��(~�>�c TModeI nf�rmz�= 2(��L�S�� {�T����� ������ ta���=�2 ��	�H��>{%ղd����J @A>���v-Ҡ�� C�2@�5��uy��L{��QC;]>��BN��n�p7� j�e��8�:�M�b)>C�S�N�4, ��TV��%j }vW�B*��M���N���� h���>y�� N�%}6a��z��| R�ұ8:�J�4������.Ɇ� �z�uj ��$�]�KS��R0 Wtf'[ �!X�g_�,V\�& {? .��SP����( �OpG����B�3H1(�#d|�P\�,P�ѥ yZp��@tN
�vd �P��� �u	�H �4R��� ��$%UN@�?��@�d��_��N�K�1�
	 ��PC�S�kX�K �W�{GF px����?�	��*�<� �ţS`R ���� D�(��& FOuف� ��Pz�]��LU��(�c7�%@$ �l��y�����N[�@�C% ;��o�bs  �������C J��׉*$^У@T`����u;��F��H2�|�� �S$��[pH50��4��� ^t�}�1�98�v R��~B�x|�@�
hI<�H�*>�7 ;�}_~η sK=��� �ǳ��_ �����D){=��� @120
3J� �;P }�@�I �`�åx)t ~!�iʣHY���Hl�T�IsVr�=�<�uJt@���CP� �(\�HA���X ���շB M��4 ~��p�N� ��|Z�M�s? ��7E�-���l ��Bߡ	(^��`�Q0f� $3N;&@r����
(^�::� ���* �@�K�Tf��L{ �tЊU�0�h1�(��:?� ���K�%�� ����+ե �����G Ҏ��.��p ��~�ŗ 3���Ec%� >6$ٚC KZ�,����H�� �5��i�� ��[$B	@ g(��5c! �pJI0> v�UR�5 ��n�C�$HJ| �}+eҖI�b/�w)���������s0->�&���/� �B�M �u��_� (����\��N~P�/�(�>��.�ф���ELT ���!ǨS �:�U��t} ��e�ZC� PY�]#� �U�xH� m� B�FS �6&k�� ���+�*� �5�0G�� �
u�C�j�z}�'�m@v�t`^ %~K�Y ��i��-'! �әSZTaH�8�u ��_Q�rw K����Ps�)��h0B=U����DR.eg �:KX�F�Ȑ� �W�8qQ R0KE�1�L9 t�	S� ,[���
�� 0�W�A���<b�t�Q6��:9v��o5)�=
+�%�aH�����--=�����'��h �Yk(�Q	 �}_I�븢d��TU��$���WH ,i;^��Nf`!G��� �� ���ؙ� ��u t3r�/c }����I U$�(&*t ��X�Ԉ� h���	3��� ���J���V�.�~a��>���^��@J�5Ģ�a9�:�2�&dF@���tU ��{L�a/�$�Z���$+V_Mt%���G� ������ ���F�`� Mu�|�� ��/�T�*��$�S�� 
���XA�G��t?*L�ѨB�5`N1�A$�Q�\f���3E��)�� ����@	DC�H�!����˫��eȭ����ى �^��x|� ܜ
�h>�����.�Q�W)��_u@�ER�&�X����t�z ��v� m�@Z���RW*1�����d��Z�����:+�	��!�(�$j�`��)����ʊ�ѯ��`"@���V�����7ID�{��V @.tg���aH�_[jU��<P��>Y5�-S^p��0<f� �̈��j,�W �C�H5}�?�� %yf��� ��>0 �8���
���SRi�(��M�^����Q�K2E(@P��?�JІZ� d�	�YX ��p�:f1� �D)h�^ �~%�}��8�����H��� �.���a� �8�q���K�H)[��	EN$]�q�f�� B�U��d�2� �_@Ī6�$y@�3��&.pldej�ͻ��#���.^ ETܣ�� �W�׾��� �H���x5�j (���X�a��*��HC �:��/4�� ��2cL
�����ȴ�B����~�?�� жz�� �<`jl* �F����J� ���f �FD��z�U 4t����� ����k L&(<0X��
��f�Z�o/H �WТ�!�\;A���� v�i F�.wХ+Qx �P�EAM��y�(0 8# +3R^�T���؂ ���jpŘC]���ո�)� h`3�+��7?�]Ts�0fD$��vIx�zu Og��N&^&���Lb��0�$�[R�N��@�&�Vy� ��J�T<�(�C���U6ȧA ��W-r�">�X>3Ylb B�)^�����$���kb�B�G��2n |\���H ���B-�� =O0���Mp C1�	]�  蛐��j�m��M����wЕ� }��9\)c� :q��Nb ,�Ӵ:�t=�O��
�1��`��#@ \`�d��0����m�0'� �V�4�{!�s�5�1@���t 4Qס��	 ��a$"- �h�����	f.�\�Pj	�X��X���];`��� ���O�K P�hQ�(���m�.����5�e �^�j�d�	�H��@������X��R��$� B���Lś�wS 24$ ���+_�� ��
H �K�����fb�q�F���c���8 ��&�R,�Pp�
ȧd ���H��'����]	��\r`N�OZ) {���� �^��PDXV �dv�.e= I��j��u�| �EPU��! (�O�i� ������" ĜSgc� �b�p>��� Ok+$U��� t���^o� '=PT ���d���
 D_\�@^�|� �"�eg�zb� o��ny��:�ȟW)���YLA �SO��~U ��2eT	} !+�,@�M��B�`;>�} ]":�a�D A6OFI�|� z;T��&3���o��HG�qXl� ��p�D�E�������! �jڔ��H<.u$� 2��� �[���, &�V�K	8���*���(f?b���)�R/B�`�4��0�h �^G3�W� {H(��79� /�_'��^� "S�,���t��H{Xjr8M�hW�g4E	�����$�o ���q�OK�� �#M^ ��>���� t��y�1w;7���$����ͨ @X��h�C D���2���Wi�53�j��"�
9�����피�� �"�T���� 	+gS״�?��L�S �)��$ � ����ePO ���Ymi�6%�� �1��vj�0�����\��&Z"��%�V F@��Y#-� ʘ�֮�D ׄ���	���s ����?W&ڢ���qZ ���#:�?D~) ���]Z� ��N�j>�� �E�� ��[:�� �e�� ��]�<ڈ$����y�)��� %��9Mu+��b5[7��ߨ��ZքY\9l 	.�D� ����� ��v��ְT��D�H����zO@M�e�~����<�I>`J�$�Os� ?m��+	v� o�/���� �ޜ�t ^}f.�˼ ��R�w����� [��� t���P�� �sO�|$X��P}�v ��d�Dyn �	L���� ��R��I�rj �K7��Nw� o�`�9�%ux ��_"o D	��ڗt y���( X���n=� �'���ܙ`b�@;3��� �.c���a<Ik �Ew)v� @7R�?�.;T�j@�ZMi���b�`��pG��z� ]������� ���N�_�� �I��J�w�|��a�qF	`� ����3�5� '8�;LS�� I$b����? ^Q5ּ�'O r �M��	g� �12����: )�O6i]� �KbU�m� �-wr��P�� @��6Z�N� _Q�[3J��G�@c�r��%d�N��\x� �o�|�[Csc�Ї������% o��hv �d D���	t"y'-?^g a$uV�j Xy�N_���;��{� If~S�� �%T��3�#h��_�����G +�k�� �"D}ȓ (�V@�� t&�
	7�� X����0� �x ��," ����f� ����^HWg 俽�t�re�@@ ����p�5h`lt��eT��� r�m���ԑq�1�	��"c�9;L 	 �e^���\S8
�vAy�*���Yj~�[�d�@��n�?2	���������L&6� y���� ���d$�� C���j���Q�n{ %s$�wq>�!�Q�;8)s��7X�����ƈ�VK �`�
�O �m.wbjp�p��?Pc�"aA}�vsn�g���DJ�uqfG A|@`vrn� �L�z�k� dti�$T@ SawH}W|� F�N�n�{g~�b�p�C�?�ol�eq;` P�s}i_D ��dy� Cz pf*R�qszJ�eވU��r~cUma�J`� bd|�fpg�DF`vRq�E \a�9cs�n���M��fOj� vdwG�� *�rT.s KcCo�b XGhlfQ� wkp1ecF8@H�r<�gQa�'U�t(�To�J�p@nk %���B�H0Kejaic��(���!�|4|` �h�8nHR	0�ʎ��tFg avc�`wV9�b 
mf}�z��tQ p!�0:o)kb�WhOv� �Egi e`�0Bvw Hcl��rAt q:aki�� m{zD���>C��} ��3�9�WM��]�E�I��!zQ�6���dY�L8���Kz�D:�Ȁ��{�'�<C���| qTHashs� �x2@Ad%X|�� �f��1�v� Ĉx�ܘ{��y�SH�1��� ^�.5���� �Ӿ�!� ��U4)3��s��Q��A �U�?�3R� �(o��}�B���@/��ý��uO�����>�@���Ц�%P �NDwZ�;xp ����:�!���?�=�_�36�%y�6�:�ZP����^�`�NꃐV� ��~�ω9 ���� 1�!�N� <�P
�z2�� J��� 1�!�kBU 	u�>������nsq�eD�^� �R� �#��1�!��,\��C���<�;�7� �mj�T U�
�V �P���d{ #� �c�u( �,�G0�4=�8�<�d@�4D�H* LT�P�fd����)��
:����J� X�����	⍧(�ҝ�54��`�Uv:L#�;h��l�Fp�t7x�|������Z ������� ��%�j�'��pOA�q՚���� �~!��	0� �������9�CN�oVp�	�����F�J��C�$U%~ &	��] ��J����$<�	������թJ����%S`�	m=��F�j�B�U$[���]�@��t�� �ąy���D�.��.د!� �����;xs Y��,z����M�s�������jg��tC��cG��pN��w��L����@ �? ���
(�,��0~#4 �8�<�ŋ�"@�� �s>��F �����~ ��$�'� !�<��� D�:�؜� C��~� ��P�75�8k_Ƚ@�����)�z��[��KJ��o�6�?�`�8~T1+4э%���{�|�uR #(���w~��n0��ؓ �Q���� ��W�g�� �z�VΙ#I��7u�0Z��t	{y���?� ��ٖ��aY	Z^{� ���� �>F2�s��x-��/y�e{� ��?]@
����L�!�;U0��EsD��}@ ��ύT;��j� FZ�/� �8�B���z)�b��S�9�w�<~E R,*>�V�w��)���Uo9g ;��^`� �m�]N�9 G�lsTˣ Ǯ�v@~gj�r���� �P��.� �Bt��Ȭ � ~������ 0��#�F3�͏���8ǌ�PVC��=�� �A�u�L��Q eBitsJ ���3�! z/����` ��A|*VNÊ�j � ndex�ou yf�r.� Ԩ�;_Р�����e�CM�s� 4�m��}��� �y�F z� ��a���Ӂ�lC����`�;�tO ����W� ���48�! ׂ��t&W�Ʋ@��*��E� ��DCN�P�>
_ eb�ѐ o�L;{P� �@q(�t�H��|c�؃�����WüRQ�B*� bX��ÆY�� KaD� ���o�<;�� ��4�!8�Q�6 �iY��p
�����ĺkW ׉Zp�y�8( L�R���9TM�ol���^� ʬ��؉H� �bCK������;�,sR� =f��q>��$��� O���=/ 4w�׆Z����J �'o��N� r��dT/� �����$gG�N u�;ksF` �
�A�{ot����e���#�c$}�+Hb��	 J��_M�"�']�@�E\�. Cache: �� 7��p��� ��P;�X��tIk��`�_aH>6� �]Ԡ��
d�3P��Zb�Wt@@w�D)�� ���N� �\	�ղI� �
3]}&?{��Nň s����V}���X�԰/�qg��&>y�j�t e-M�U@�۴�<TS�#��$#D�Ⱦ̩��)2�_��.'V�y�C��� ~�G�Q�>/u��z��tr ,�Ř7 |nM��GX~��Ҥ�����'	�zY� WG�� _���C��+ �;��<^ sq�K$) ��ьb� n��F�\Q 2���Bra @3�0`;� �F�C�t�u���f3�(�G� �zs :��I�{��D=	;@�c�:>� BuS~ 1�<��* ������$�P�	�$�f�C�Obta1{ȉ� QA�m��,�t_ ����K>� ���"��W�Zh�; 8;� X(��*�@��� ���_H ���u ; �sE��v'�L�@J!����?+Ȅ. ����ˏ 
lY�M޾$O �+�|Tyr?4B>,����1 �k'�S< �@�+ ��v�L���8���%����<����溜�I
 )���M�� +!�#� ���ˮ� '5� � ���	�� ��w�v[2 �7-\;)�D��� ��� ���Ε�A�\И BS2|�3 �l����� ja6[��P �s�C��
&�cz�T�$Z�d�hp�e{��>� ��*% �|$���F�RL��?�X� ����L .�&�%,�#�;;� ~zPD�� H��!B�0�ᷜ��O�9�jd�%b��� tx��D��Pw� ���0��� �;t~�� ��֙���# �	}j� D��<J� 1f,�@Y2�o�O;�̊0	u��] ~<O��X�)R� Q�uoӢ�|Dˀ�/4�� �f;g�l� ���~�>�� ��A��LH7�s���;��� 0�.�@)� uŃ� ��D�B��:K���@�+� ����Ss ��'[w�W ����Y�z�v���X��G q֟�<jNd |y�O�H�.�KG&L�� �st�% �ǔ���(� �I�T��� Q�A�� ��H�u��g�n���)Q\�0~ x�WVU�r� J֬ApXP< ��� ��߇�1����"pU��� W����G\�� _x���� �ݝ�~� /u� ]^_eԲJ[$	�Y��:��I�M��P��kn��-��>����)$o�X���4 f���%]ꮥMGR��6� #��vSP� ���8~e,V�<�RQ�$�� B#tTCX�*��>K9�wA.�x@	 t�R�(ӈ ׄ��1ҽ \��Љ z0��uk�w(
�!��ՀF?��4 �aXZ� ��[�tdJ� �|T���K�)����;cZk���D��P�E6� �>��
kO �Qe%h@� ��K�\�Ǡ� ��:�9{ e��E�� ���%�Za�<�.�RA&/�'|l�ݠ��IM��Ơ	0�n�=�;������� 6چ($̐ @j���{8�3 ���;� s����k �rg��� E��+�DP��� �>�a	-H<�;�v�M���#6,���l>���Ҭ� ��T{� �\cD<�X/Q�C` �JP� j(L����
 ya���Q�\ ҃P~�uv9f{�d鑇9 �!�B���L�؃�,�p� �U�e���i>u!}��I=� �¤���� B4�����}� @��A��^u��Rc�_����tS N\����B ��� �ǥ��x>�~��Ï`k��
��t� �:�ڻ������p�t )��J_���HL��P��}�4� ���9�t �BL���? �݉���i 1�@������e ̨����Y �!r^�� �F�S|A�0;"���G��0������@PH`�gG��
� �*�`_�1���$�Q߰�� �5��0�)7P@iՙ�� ��ߖ*�0� �Bv�H+��;��|��4�x'�g��8 U�/���� ��Ȟ�p��*�&`�M�
��s�A�;�@�e}��̺��b �)r1=�� v ��L�����+Oǂ�3�b� �G��ʍ $���'s� e�;��u:
�RZ��VOJ �Np���<�� �V�`��� �0��jɕ%R�b� ���F�D �鲎M3AL%u�7 �˃){H����$8OW9Ҹ��͎Qk��wz�&�v' �R`�. $�:�S�� G���%CqQ
����� D��=�rK�0v4� �w{�Q )1BU�D���î
��<�W�+���v�'@�����[ 	�d�eY �;�-� ��Ф���	J�I��6�U��O"y�# ��2FBV.i ��}�
�hrGU�Qp;u������cK�D� ��N���� �3O��5������I�D n)�6&����+� ����"^Ԡ��}\E� �@؍F��� ~&�H���� ���F��
�u�E���`g� �猝 p� $��JbE�;2�I��S V� g������ ;�٤�����_���
į �Ah��w� �;ޘ��su��w�ǟ���ش� ���H	.�<�� ���LW  �$t;�y��� ��YkZ!�� l&r�奼, ��HəE5�����#�O� 	̆،����upa��~e0�� "*��+�#;�� ��d%� �,�FoӔ Eqt������ D��@�� ;�w]b�9�_8V�S��*�=շ ly��"'s^�b�cze����{< La=g�3.� ��Q��y�k���$xj���K��� ��J/Z� �T�Ԑ-\� ?���6J� 3mM��s�C>�U�;��T�A.3���OL��Ԙdк�Z��� ��9�'%� �pO _�� �&wU;( t~�c� ��ׇy8& Є�=ԋW?e���} ��R*
�:�:�[�2��_�� -�r+�` ���/�6���r�4�+:�:",�<72�	�$�SE�I��O�����ģ�X�@��@8i �vqk	� 
�J���F� ��5b� ~Ap��<�ua̬Ü�M��Y��H=b�^�����J*�G`�bˁ�ud�aB0)9s����X�|D� -��3uN�s ���=���� ٨�ܳ]O��]"�d��/�m܃�;�u�`/��t� ��W�����at>���6[3�r�G ��(��~.t@�_$������6�v*5� O��JN��)Ų�_(��`Ѷ�.�I l%o��� �w��up&��ҕ�N�w�� ��yR)v�PX�u<Y����T���F �H0���]�$ \�{�E��� ��?��^��?s:���e�{O<؛��g SZ1S#-��z��~PR]�UK�b ��|:@����s@$��QZ�� �*	� VP���G�T�ҊU����� ��y�-�zn�/H#|��uD��������� �;�c름��ph>H TBF)J�0 ��W]�� ;�w�5#� �M2��;��!���j�-�XD0B ase256To MPInt:  L��g�h? O�S�r�Nx c}ds�Ma���SOz��[ �0I�;_| ���� �1=��P�~���l� �	;+�<>u�m� X�CBH{ ���_���k �Q��r������s�$��b�`;]� �tW���L�  ��$D�=� @��TcH����\�NK:�<| �}��#&���|�5�K 1��l+�>� ��鸄-�8��u�	" U��f�4� ����s- �J���� O?�HA�|裢Dwl�%�S�����r 
v	�E���ՙI����#� }��!Gv� �-�xa(� ����;;u���i���|�
� �@2"�I�rU�0�X� �/18 �A(�^�=	 »Yϔ� !�j褧 h������� ��QHI}� N�W���z� �k�g܈J ��6@���	 ��'تh ����l�&� �U�MT��^6�s[�0?J������s�Yب�������B�!�lu< �v$�I�kVa7�0� G�M)؊�DY@$,�S�b?!ԝy� mUP���(.;i`@\?o܀�@C�� ��R���� �3��	;)g��?����Q_ԍ�� 	�\��?KT I��Ps`�x����y c�}Yv�$� 942+�KP= s(��� �B6$�^� _!Y�1�"��F㛬�c�0=
 �+����Gǩ D�2� ���|C�!� �������� (��O[�� ���A\� ��U�!H�Q�*�;ɀ���Y��J�I$���> Őۋ��V ��o�X���|n�ǚ���T 2��g���K]��d��G��Z;���8� �f���� ��Z�|(hdq)���U~��	o 0����y� �%���@nu���P"f�`� B�׀�6X�R@��)�b P�ruJ��� ��"�#�C������n�疠p�-  	��|!����h�B΢�U'����Z?3���K� ��x� ����8�.R� �0P���� ˟:dR�	��3���Ŵ~%�[� "t\lq �H�!�9~�� 87�Cc�J���NG ���X�Q T9����X�� 0�	��5@ �)%�&���@�G���4��˓�L M*�� +��r[�����i!�]�� ��~�d��9�&PY` ���O� XG��k��x< #|Y1[����o�-�Z���	��Xi��~��X�ɀMk���U���q�Y� GZ2f���F��Ķ9� ���{+< $9� ��F����8N"�
�ub:[aN��j� ���A�=���h��@���u���F�/���H��������`����@C�q�[ �S#�"ZK� '!+G���|ˉ��P��� ձ��.�F-�uj���m�<�#�%�Ɵ��b �����0u jV#�>�Y�6��˸ G4���Ũr��\�۸�bl 1�Dti� ����L�&{/�`�Ҡ���|�&[����G��>w. ����O �k���F$PC%�|&ɋЉ\ '�+�� %Z]��Vë�|�P�3+�9,S-�fs�Ȃ.&� g5 tVq}���� L��]���F:0x��jA-=O{_�
@�2�'�`3�Fu�Y4�9����!6NVt���	7(u8ݖ��� �tb| �{:���	%i��W�kDk& �el��T\G�<΍���+�� ��5�� T{�()8! �k��F�K��[�4����`�y;�9ٝ�@�+� ���z�0�ٰ8��cB�q%�� {Xi@ܐ]��Q^ �y� J��fU� א�<��Ο��%�`F���ƺ���^j� ��R���n ;��ֻ!Du�PB� ����� ��TQR�����@H��>,ɀ|��-�{�����ㄐ���a: �"�U͂0 7��HΖS<�{ ����B��- �3�+60 .�V��\:- ٚ�O_&C˭�ŷ)���yR�9;�" ǑK�`� 2��;�(T N	t�����A�Jw)�u�&*,��u hʯ��� #�B�R ɥ2LU$�v� >1�B� �A.u� k} `��-T��� @&������\�#���XC<5 ���/
¥@�J�"O `L��PQ#(��@8
�w����� ���@P`�p� ���x2s$H �RQCn��.	�
������* yQ�� V� �W9J r5S���7 ��@���5�$|��`�� ���z:��/����� [�r�H', +��ܼ�� &�%��4 �a�>^Y�W*�����`}�� �� �� ����/)�f�SUV�.W+Ū��g�, `��[�� �; -v�P 8�\�(��� C@;� �r ���( ��Dh3c��� �8�]0j ('�4,�}���H�@n��7 �1~`} ]<���X@�$l|�M�u6�ރ,����� (�%>+�X�$� �jl'c� H�9f��; ��T�� ��� {���ꄢJ U%@I�Ů�5	��� � �b�B����`�]2&�[�� DKH��� a�;�#	�1v�"ϐ��� ���h��� ;�7�0�!}G8�<A��r̭����JW�� � �r��@�A�MT�}�H���� ��ʫI� �1�x�4s�''c�L+� �� 8�%�i�\� "d��)�� P�܊� ��;�F,0sq
\(�ޒ?����s� �� "4B��D8�@<�a#;p9y������ �(�qf�=�_�)�D�1�
���� Y��Za�4@�Nh ���� 8�A_���C z���@�� :rH拇�O1Phцe� �B�j�����0!;d'��\ i`kN �&[�� ѾK�WC� g�my~ � ႣTj�� (D�����P�T?�X�A�`R&\R �ʪ脺�X_'��E�ف) �k��jG��%����
�6*S�j�4C��0�p F��r퍻 �x�K�P_� �]��M��Y ��l1٥�@s|��R������ 4$F�` u(j�Y�V �0�~N�"�p�`}HL4#H[��,��e6��j(-�~W2w8ơ. �FH�q��A �se< O ��RN��� �$�)�WPK"Ì�4@QF��J�� ƃdsf
� �+9�uw �r� ���`��eCҊ��n���@ ANu�)CQ G� (��^ ��$��T�]r�:\��8�p��� zW∋�bg P,�CR<N�h�=H�s��n�֋ ��#���5��O���%A� �谙	���� E�A�N���ͬ݇B�?�� �|�鲛2r� ��� Z��YͣV�!N��p��O~,�f�.����g����4m��ה S�`�P� ʰwb� ��D-��� h�a�blH����tv ��'rq�� �o�"Z31 ����HkL,J�/�4�'� 1̽���SuW ��8s��y�~�����81F.���H?C0ɯ ��� [Q��Jl� �� jx�FB���Z��ҳR��ظv ���s� ��'���t0 q�c�*�? ����JI �����X� �1ݎP��A� 8;�p�sJ�@���� P���$1{r{� ���� ��4���` ;n(�ý���,G,� l��s�f(���Ј��p�H�w�sT!,�^���j2� I@�l��o�̵ 	��B ��}^(lEC���p.LǅDs1\� Man�g>2 �� �0��* ��ؔ�h�@p� u�ㄡ� XD觮ϲ) �z��^x� F<}j��3 O�>icw{P�t�b1V���  á8P��;<@��0 tV !}[��uj ��M�e �a1�S�[HU� RG�6�: CbqVWA�`�Ȁ 5p�<������@�1� 0�t[`�)of�b�`.�[��TӇ�E�� +��I�219!*��"/ =eA�sЩ�E	��?�Qxsb�!D��X��B� ���+2�)(ݕ�A�����q��T�v@�Gz& �I��}�B �@
_�CH)g UÐ�|� �_��#�� �Ϯ��G ����7C�\���@���Hհu�>L�w���,�ʮ  
�$�u ��/�&U���G����Y]@o}�%D����������?� � ��$��3(�%�m1��-� �ӎ[��}� ��6�/V ��N.�S��L�� ���1 ";a���Y �m(bo~�|���x����� �A���!��Œ <��(Pw0 �'Y+-�LK �J�|�u&G��� hߐ)�Q�E�A�ٮ4ȿ}�b��@�p����)ɐ�p���9 �6K�� �_���2� ~��Ħ�"� �p�K��H Pthe#3 ��,)�u/����@�j*#eW ��PN�� �=hD¯d k��4%�Hc�p��A������k` ��e�r37* ��[�� ��_�5 8үˈJ�� �����=b k������ ��O���] $�.�XK �j�;�u�� y5�%@sUB�^�K¡��0�RQ��a��𮎦 I�A��Y"�p$C�� �,ִ� �%�7��� 4B�X@���� Aj�W4q�0X�� ����^=�� ��]�6� �N��� �@*�B��l� ��8�;K ,��}X�9�?B Pܽ�Ե}�8L�3�Ÿ���j>W6S(� Rt
X �/�8�w$*�l _G�D��M.�:H� �1s��� Qk!����� P�u<a���Y��\��&�� À~,H�� C!.���F "��:�n �[�j!� 
fp�.���-�bo�� 8 Q/�jr p�Pu&?G 
�fQ�7m� n�Z�P-�Dc��0���>���)�.�=|- F}�X���P��	���B� {�d>����� ��${p Vf����	��N�֝�CZ �a�	��܁ R���w+K'�O �t�r�7 .�:4�^� }�R�! u]��	J� 1��ɪo0��Z��� �����}"9Ӏ/��0����� ����\�_ d=w�)0��n�<P���y���~�D0�k N��d*��C ����	Bx��Ԁ�WL�� _Ӓ���� Ou�Z�� �[�dT�";� V��#�&7�E�ŀ���h �d��J.7� �0�>D�L \��x�7�	�+� ׾U!�$V� A��[� ւ*y\�E3U�,Y@OO ��ZEՕPC���({<��~\�� ��]k�< p�Nq	�o �*�Ч-� e���`�Unr�gist\d4 V���/y�D���k�l�Ʃ� P_����Do�@@1�J>��"�@�/i��a H�I���dz�N!up�| ���i;�� �$���z a7Y�nL� ;�uM��{��D��	��8q :i�Pdj.5 ]�"�����9�M�A���z� *�O�XD n���@^� �:�����)sC �.�
�E�x�������D� ���#�x�>�7���g�;Kh�ɀ�ǿ�FaCMu`0?�L�H ���	��tC �q�I�y�s Xij��ݒ8��,PjA921���!��x% ����qt��z`�6�:����x�B<�� A��#�v>p&�(f��	� �;,$���0OD�H;���S~�$0# ���5/#i���u@��9��x� �k����� n������,�� ���H�� �5�
S+U�� �2�`F��GtV��Yd (�\;��J S��%2*,$E^�� ��D���m� *w������0G�/ e	Ry�~� ���VbOW	���lL�d�qd ��Q {8��$T�w�Ŵ�[�f Rz:�%��}�;
B��Q� �+3�E�� ��H�KA�1@�m� m�P�f6 �s�Dd���	�b�g {3W!|�N$��>7�ʙ�3`�%���[�=�t|�c2 Iby�� '_K����+��� /����[(R�D@oÊ�@�u�� ��{!��2�X	�pi&�M����
�͞���@!�	 0!��=��X-��nP�@�ȱl c��N�T4��� ��AX�uI�� 1� ]݆�s�.<�O' ~t��m�#�ZDЇ ʪ���3�`���2p ��4N���S	/�=� �`ꨉ��� �!�F+j �Ad�x � @����?氰.
�� ú�0�}�� �^#��OJ����D�:gH�b ��
-� �c��~�	OԻ��ו{�IWـ��K�v,�� u
�~e��<�,�X�tJ�rU�s��P��j�1��8b�v� H&\C�9 %;��Y�� +_�gj	 q(a~�A<=��,�r� �G$:5�= �̫> �1<�/vy� ��}|��d	K�^���X�& �
h%��U29�� ����@�"X�� lL�E��}� ;S��:Ii �Q�kV�% _8;�bFi	t���gu��,& �����ǒ;	� |174
 �K�AB� �V��	� �~%��7�x ���w|,K)�0 Ggо�r^':�]�XW|�	U CЍM��+ �ג�V�t ;|�QU_-z�������� P��-ٱ9'u����GzK R���n�"� ���E����O�ү��!�\b�.�� �����N8�δ��|�4hZ�}0JT�P�@��%C�ϥ�� PS�> `�O�|:P��H���z s�p:�_f�6L ��S ����?B��ݢ�JI� G��	l9� �B�m����M(݀���7T �i�U�\
: ���J^�= ���tT[8 ��i/z~� ,��C}"  ���]Ә1x!M�O��</�B6sC�}��t.$�m��0��I��:�8 fv����� }e_��� i�.-�~��o ���4�>p [����r�.��� ���;�"<� 0�b��`� ��Q-�	j��EH��ȧ� �(�M����&����G0ӳW ��e8ܥ6��h �t}�@$��:�(�� fR�JT� 5�Z�L w̻��=��e�؀0^t�X�!��S%�]���F j�6��,� �5� �3A! �'n^y�(O ��MJK��� �2eS d�-l4J	.q� �h�t�����3 ����ɳ�S	�w�`h G�J��%<�9 �#�s� �,u�	�� e���G�� w;�~8� ��t3Rd�+:�D��Y���'� "x�3)W� E̅�.p�� �J����܈U�� ! ������&�V3	�֎w�u��#� �-_S�\�w��y���� ��}�2K�	 ���p�w ��o/�,G ���W� �l!�_N*MUS<�@� �.W٠O�2�YJ�#R�u`�N� T�X�ַ�| ���!�˲uP��ɏ�O
_@7Zʎ&'����\H�p 交�۞8
�Ě��F�V r� �u�;^��� �KM<��(9+���G�����Ǚ;��{ XQ,�f0� "�:1I��#Ouc������CA|� =�ϋ�OytL��=X�0�� J�i� ����(�K �Mt��3X)�CH�۽s�<` � ;���k|��J����['�} F0�ʟR�� ��&B�$+� ������cu(�F��I�<~�&�?Q ����� , 8�� ��^�ԧ� �|�b"��1���KBdy�3����O�@�$X �ه抖����2,�&�`�� ��O���� Jb^oK@~d����H@�PCuA�|�� :�D%IĄ�Y� ���� ��B��wQ �L�	)�j ��i��
CO %u�|Tx3� �q�м:
 �~1�H� �`i�� !:P���Ҡ� F@I-u�x&�!x N��"�o �2m�Ds�f� un�&�� �^��3H� -���xJ ���}���HFKu�EȈ�k͗�����K� d�ڀPx�� =[�ŉ��i dw��$Jw> �(Kj���@�����\� ˨VN� X�ԃ�]�)j��`���z�5 $����!�7�+�Kd� ོ�!�*1�-A� @S��B� 6���m�yL�\�5��j�}���= �CS�) (*�oI� =D�uH���08�@r#˔EIb��
�ڻ �&��*� �9Fw��� J�'��a�L��{�`����QH ��\4� +;�K� 	G2l&i$�L-y�O`9�� %f�,�.� e
!_j9����5�R�� ��̶<�� TX�0�|� � /��	�
 N^�����;�+�y�!�u� FuS�É%B;��)��
� �"GW�#<� %^ M
4�Q��!�%`�I\P��<H���AF��� � ����i%vE,�s�� X$�f�=��T=uN��<" ��D�+U�K/Zs*v>��眄�8 ��;���� ���t�� �Si���� �Y)��߲$��\�kH1]�����蟚��� �6X��&$c �]kYK��_��� u�,iDm�wz� W?�NU;*�s�~���T�B� ,Fk ���^�심 ��\y�O��S�a!� �-)�\��l�k��ķ�?�� �v�Z���)�6ߠVuw��XM\ j��E�"�(Τ� K;��$��C���-���� )�����	!_s�J`B#��6�ʝW"0T��{� ���*,�k<��$TL �\���F J����P�bp9��� ��K ��k��d� ҧ��[�^W��{C�Ȱ#�x�vd�c��F  }eP��) ,�L��C� �ߢ�v�3� hJ)t$8�D ��æ7��F \��u�W S)h/Ѡ�*�;Xq$��Հ����Keys�.8�N
a{m�Ldk<P���orEږ�=V�lue��@�t�|�����x������.�Do �Q��ݿ� 2��Ԣ��UH��>,�$����!���G�S�\�3 Wn�<� ��?��H � 8��J��� ��LN�ADG !�+
� RE]����;z���K�@3H� ���rMhi =�S�(�� �Et	��;����
h$ �q�e��3��#�����,
j���K��S� ���V��I��J4 ��P� ��j�u��][s�if G.��WVx;Ծ Zu|�I�G �r���	(��zP��*ctX�BUS%�^�'����)��WĦ �c' 5"Ӏ �=�;J�:�P �M_A� ��%����Iw�	2S}���M� g��t���~O�h����� �"��v�_O A;B�&�� s�z}Q�f� �a�_�
� ����윖2 �d��l�I�?�#9� ^ģ[8i� bxG����1 t\�Ɩ�Iۥ� �@�� ���}D!~��Lh��oô�pм�' ���_��,��Љ�<0\����<L��D��aX������-�8英�xc�����O ��ݍ=l?  .w�5h �`���z[	��*���@�\ $N�
%�V,Ff�@��� <���>t�/���3�&�8�Lr ;�w��r� �q4
�9b��)��0��Y~��З� �(����� ��E�%��q�y�~�$`ٿ2� �]���jN� ���"쀸��z�R؀�N���y�@��ȼRk#��x y��j`��S �Ce	�X��} �@OǲtR�B�ܽ�9�A���PV� 0K��R7���^�-� �68�P�'��.H/E�&@� ����Ge"� u(�����
%+�
� �\�jb �4�hC�S`5�8�̍<�T��0\K %t#x��V�".!�: 0d(L	�*�:�بi) �+�� �.���� �A���������0�U�!�A�����ЯW�]U�A�6R��sSy?r��0:E���`��"� H�Z�<j�� �3Jm7U{� �C�+�R��j?EJ �����N�d����e�v�\��~ �5T��j iC�I�� &�X�����k�����<��9� �l�r�?���|\?�q c���� db����� ��������\����}�� �� �䳥Nu�]��I��� ����q� �������Џ|�~8\d� mpPi�Lkn Ij�K��� �h{U�Q<l=i� R����w������GV�܇'cH��r�m��a�RP�^��q�lf����� g��`��T@UVX	3Y�b`W�T���|A�#yS�'@B��������s� ���iu5z �X�����8����N���648OR PU\Y����� Nw��[�� ] �\�z�� �gZW�� R��n��� ��f� *. ��������ڥ��g�S�);�K�M��[& r�|�4����n}j ���=�����N =[��4�� �;��<� ����8ٚ07+������w��\���3`��� ����\ T��{���I��G>ywvq1$�� ![\���8��Ԏ HI`pDR� �T�ZU��S8Q�����H�� >��[�Dp�p� X��24�� L��*큤��� �RE����d�8���� @���946yF AT�|�=�� x��\d`f^�v]��[�� �S��F�@_ ��8����(��V� ��� ��F���XT�r
��}<�8��`� ֩bf8gy ~}�����8��JI�R^c� s��yY�X ��]�U�0E_��s�@׋�34����d�� �\�=�u�$eI7P&�P ra����pn.�R�� S�����
���� HG~ �da@n��yN[����c�;�Jz� ���u��VD�* `�쐌�&��J� ��'������`������� <927;���*w���IHz��b�!���g:c^8e��i�L�L�o 4_��,]��$ �&����W�<�b��{ ��j
�Pm �~��Ƌ� ��@���m hj��8�ȜlvN  ���e ��X��T� ��QZ�%�� ��I�Hg�������14����*����� ������� I/�����|�u�:�׎�q� ���Vo[s�~ r�'3�����H@ ���<� 5#�O>�� ���c��"3$6��P� ���fL��^������
�㉵�ǆ d������؂�@���΀�� MQ;��8u� �_��`��d���eU�����\ ����a��-U0 ���t� �	)��f'��0����y� ��ꢿ�� +;�?"�9�?��X: %*o�� v�Cw��x�M���|���t|� a��f�� �$����� ��Zm� �;�S������.�g���Ȳ� �CHF��\�� �쪣� #<Z_K{}|B "9pm@wtCus��$EG�оV�@& 9<�,��� �Z�Q��w { jU���� ,�����,��� ��&+)z�&�5� 2��N�� ��B�x<y4 v,zs-}�;k�Ü�;QP�L ~|���������v퐔�_'P*� ��3LI������0�$0�W U6;9c��z�8tu�%'/2�� �y��p ��gs�J���ź��Hvw X�T���� �|N)�O�� ����b�ǩ���̓�.� NLK���	��1�%`c`i:C]�ol*�%DG���``�8x�����g��{��� 25����q� ֤"��� yF|�S^�5�*j0��:,π&���� �USR��� ���jl⬘p� 10:BhmL��$��7��� �Q�с�����p �u��� 13�ǒ��� ������8� g�%<��wV,��� ����� ���	ʀ 񿽼yzx;v������ 8���>L� ��<? ��l�����/Je�z�)
 21���� �~��'��|?��Z�*�jq��:������w`��p����GIJ��� ��@L��_�v� |W�ć����}��@Ϳ��	��+ ,���� ���bI��H����RV��� ;5���� ��P(DEI1A�B�������� ߨ�d üj�p�8[X&'`0@K��\�1"GEu���j�s� J��q���~���E`ޟ Z)�uV6pJ����`:(� ���q�en�8�� �|��S�� O�vR�lqp�g��97̀��4l��5mw!�Jȕ't�����TVȓ% F_���|� �̯C����9��n�� ���x� �U��W �n��8����	d ͒pL�S��M
��`���w . a����� ^Bg��!� ��pfJ�� ��L�R ���"��� ���B���� I>��z�� ��%��n�� �is/(D��!���`��x���mb�ȓ3�� (.��o�0 Q��_O'� H~�f-�X���@��.���� u��GW�pR������l/
�HJ{��"�S�� ���T#� ��x"�� �kE$[YHsl����ƕ�M�"b �%qJ�����+ 0��5�Ϸ��ڵV�� �b���)���R҄������]Z��� &��!���~�F���j�B��P���S�rsБ�Z���!M;*^��J�m�4�,�]�Y`. f�6tϻ�� &*7���.~V�K�Y��Ώ�
 r��9�h��_�� ����� ��-�e:!��G��&"@ƀh2�r-+eJ�'8M6S�pa nUs
 ��rif� \��P6� �p�j<t�"E*a�,�h�o>�d�P"�sfw%r)R:F` �1�Pt�.;�H𲬕 ���Plp��?(��$Z����P�� 2O��u���� ��c�ed6 '����@b0���;3<ְ�� H�p�6�U2	/���0�E� ѵZs�� ��\}
� 1Gq�-� ��A�; �u��~����{�?�� ��.I� ��/T)w���Op�fu' ���i�*���O��o(�=�vW !�UP$n� �[�ш	� R^�x����HD� ��j7V;� ��8���Q vd<�,T� S��R�7 P�0hr&W �Es>�,�� �D��?�M� aBuv%Z]�;��GK�� Tg�]� c��i���{�<������� _�q�� C�hx1���c�������* �uP�EN� �ʞJ���������j.Z��dI�ho�'�] }礒"����  ���Acti vZ��D��l�g.�[ 8h�E��� ?u�8x-|`tWH�wf�}� jU��
+���e�&�� �� �uS7��q) �:hDJB� �S�#0��@uGhd��)��'o�ä Q�,�In}c r*e� �� �!
�4�C 2&S��Ϗ �v�$���=C&�G�2yM1" @trP[ ���_lo �#�Z�٪!r�/��㡴2�F� �g��֕��\��L��;�s Β
àM�� 4j�^�0c8B��Њu~I U	�w��j�$��x� -.1�H� 0�C8�) �$ ��- t��5� S0g����2 &cW�?� bŋ΀$�V�% ��\�B��� ��D� �돯p�EF%� �'��7� ?��do�� 9jN��k� ;�J���_ ��t��4��uw Q��n�׊O �CiG����R�� 4A���W��	,_� �.�j?]� �����B{� 9�:��X# ����>�=΍)��J�7�y�#j@֨4�� ��U�NC�F 5�+�O7��-�n��GE-��v� ��Ke wD�T7�* ����X�� �:45��� ���
%����F*�E(�^�
�O�`��u ��R_e� B,�J��l1��>����x�Win �ws��t � 95�{�� �OSRk�P� �8}ӄ �E��M�<NT �3.%u
V!4� �20�`���% t�C��Nr�=�1����@Ҙ�y�y� ��J�a&v͒�D8'z���?�� ��)��3 c��h	T B'�*OK~ �4&u��\;B(����� %Y�mf> �Z���4�\ �tX���������Sq� HΤ�W�J�L ���; �-k�Ɠ��҂?��uB |�E��V� ��N��w)<C0 	���w� :�*�[��N �����
B���} ^jʝ԰p��:�>�Q�f mJ
�aN!� ��pb����F B�����Ss� &�}r��~?�� 9t�g��:�� ��Q:(�  m
k�5 tUg/��0��6(�	�B}����]%���,=̦� Z4��� dzx�y����D#�X��Tpʡ��>@~�o
�' �(�<u�X�.�og���_A�&��"C����	�K��m0t8� _
��#e ����|� fB��A���4�`#��y ��~e�J� oU�=X�r�2�� @P��|(� /��}K��W
��'���RpA= ��dv \2G�1/tj P�<u(f �S��G�� �
�IHP�M� 3���� Rn?��;<� I7Z23�`9* }QO�% G��=��� kj\�[ � �P�T��i��Z��3���� ���]��� j�,p�Vԇ
�p�;� 4�����?�h��w@Edu�_�'$�	/�ǲ�< m\Cuhy=n\w�J {S�\� �L5O[pIRsE�WpNT�&؁�?�V&���LANM Γ'��9@� ݔr�B�? $wv��?}�
��W�|E��	����H�y}2>Ie�z��t4�E�p�uD�&�� *Cx�|���� �S�{4G ���)�R� $��3N���Ih�2dg��*#@q1B~�<�� G����ԥٻ!�{���b$�����w���qp� ��	w+"9� �X�OG[��l��|��6F���қ�˴ WorkŢ��O)t0��iv}�� Ad�anc_pB:��s��om� �F iT=��0�C�f es�-+alq7Dξ *��VJ]� �٥4��\���r���2��>���9v@�E�]>�� �!��ǧ��[�E�ړ�� Dr�7�V�;����K���� ���ǩ��:�U6��d`�C.SD�*(n�\9�YTE M�	��&x��ސ@F��iJ ��p/%~��^GS�F�\J2�ߣ M6�W\�{ �SP�L$� ln�^3�= ����%D� 1�C�; z &����A �u{���6\#� &�K�
=� =� �Cݒ�Z,tW_Q����
��K�����>;0} 8��J���� ����+�������<����l;ߘ������ ���	B:C ��su�
��Zn B1VHŘ��)@��� �1������Fv� �#�)0�?ԝ'� �� �M� �z��_@N ���ע �v��� �x�D�s��] ���N�g �$>I�� ���*Ca� �}�Hct j"���\Q���< �J���K _Pj�Uo�Z �+I�@x2r d��� 4�-=i!z����X:ب5�&r� Yc�� F�P��� ��"��2|+� �ȁ��]� �a�ià� b-Q��D ��m3V�(�A���51 ���07�v �]���/� d�H� ��NR@�,�9�u��[��{� ���s �?�[+� �3¯*�12 ���f,F@��d�|k��KV���'���_��z�~� �!ad�c�� �7��b�+Ѓ�?��6�$D �U0/�L� ��X�	������+å q�)�@1 U�PR	�W{yC�������[��� A�} ����( �7��C, !Ќ0f� ��X4�{:� �n_�� h���Om+|� ��0�wQo	��|&ڔ�D������XV�@�h� |gz�<�"HD��χ���6�� ���� �C|,t ��O?� 	.?�q
�d�C����p�i �7�6�� �	1"EDYm{�L�@��{6* ���.��c �T�B�8�h��q� �) �Pv#(��� >�"� �\)� �R��	~�Tty�&�X����|�� ���Wz-~^ ��;ȩ��* �<
,�@V �Jk�.Rh�z�_��}� (�_Ÿ/��� 	E!O ��H��m|t) .�>�์� H�ej<���֙ �٬c��[M%����6��brd���� $�3|��P ]�C�LD �<;�"*� �2�6�!�Ieh��
b#i�]E�l� 2\� 486;DX[pc��� Z�0�S}2���.�`�����/��Wri&� Back E�n hW��+ 4`�-P�]i um�0jX^� �qI��C��Y�nZ���� X��p0֥1;Җu ��u�P(r����%R)H�4�_�� ֵ9 �P��^�X3{�H��.���� ��F����:	��{�̽��2N@q�%^b�psA
�&��T�Q �~`�C� i�F,t 	�\B4�P Kd��:�� y)w�.�2�����F��� ʢ׿(�C Xy1&xLR��`M@�aGX�|t�06���Rw ���>u(Z$ MX�H�>V��� �!��2P, ��' �@�x���P }H�%	� "��X�xvz !� �^(�WP��	`���z.�; c�w�$�H��@���"�QP"�`��8��u�d�"�SPC@ޡ�p�1�! ����# �"	�AMD�\�m��	( S or� �5*��y-<KXԢ0��@��1 ?�2�3�R�L|���aw��  ��d 3.�Unk�ow� �EWl� 1Chip��\<#�l�Q��Lv�t� Transmev �C�uo��;4��� !T%��FHM{\�`J���B(��Wk� Fp#o1rz�u���.x� |(ER�~�׈� ���/dWSsQ2RVv`%�� (��HX]�zN��?��)|h���' U��M��}� Genu[�iǧI��	��:�ˇ!pq�i�A�t@�N%	$c*�A�����Xub<Ix@C\�3c�� ad�*�$� R� �J�� 	��n�� ���/*��O ?M��8�:V ��x�]���}��� �����6��%> �;s1��G h��$ �Sj���9� ���,M�v� Ry�	 �g�QY �2�������u"�f�Q�:�����*ځ	u�Y G0�g�@m�� ���~ HۀU9�� �ap���(	��B��w��� �<, �&)Q�K["J̀E]P�� ����R�\+m��G��y����4��fL�H����)�Z�<����G���xwB�|V`걨EZ�z�*k� �޴�  ��^Z_Y[ �X�v.U� Qa�#)kpN��(�����t ����<
� \5�0�B���!Xq���
#؈���^T�2D�"(�+ ��N8)#E�!<���^@`A� ��D��}��;����J%���рz��e��/w]��4E %��~��e<�]7\2� ��xrs�n�1HTM<K98¼��_ �Ĥ�(P�B*�� ɺ$ �~i|�-D���d���� hS� �l+�N��D� �[��: ��$���J��PH�2u"���S��jI��%��Z�(� ���� �ѯ�S�Xǃ QDZc�l$u$����"���� ��v�0� �m�C d�8�[�<�R���I�P�$L< 9YP)��T�X��҃\" �`	2��*	�.OM��ker��o��f�+�ȧ/���4WN �
!�d�,a����|�At Yp
R�Ċ+�l @���	 Jx��V���<(躯p�/�P�:����@��.�ʀ�����}��� u�, &r�6ð� :� �����v@O�w��9����i)�@��#�NQ��Р��9,� F�u.� ������� ��z9+ ��@j����|���Yf �')S� ֹ��:H}x [z����p�$�z to��I( ���/�2� �>,r|	j ��R��D� ؛�Ю��ZU����,B~$�A
��"b���:�?D!��H	{�P ���o� �Q/T̗ �^N$��Y4���������\K FB��d c֬���G =�՗v8 ]�����uF:i� od	�������5K���� P��u2�� Y@X��$v diBn.�T0��!pV6)=�DE ��Ҥ��N�,PH� �+��S}y��i ����I�� Vn�
'r� TRhU��� ���Ү�� ���YNZ��V'ar���D{� xe�:-t�LP��@U�Q�����ct�p� ?�f<7� �ο��H_$Ո��F/�)p�� �P�\�!�:�,!��sx����`ۉ�{ ��ɻ^"�0�a ��{Q�eh�1��,���^�T�h��Wz�<�����ŕ�|�̀,:� $��C� ���4֖B��c]�pm�_ �[>�~�� "\Str g-��'}���i���Ȼ��J]��Co mg�s
,q����p�	y_����1�dT$��C sc	�p�7w�4��T�� >�_�c2.�Ԅ /+�#��?"Lp O����TW:���B �Ԉ �r�Э�� ���0L egZB�px��hRt0���|��� d�m�ks{J��t��O�@U�I�ޖ���h25�G� ��ĥy�J.�Y������2;DSpec���Bu	�d6� �0����i<eK0P���z�� �p���C�/T���p ��� �]�d3?f� ��v�&p%�V .Osx��8 ԟ�����Q� h`��#Ͻ�oU�o�16�~P����]��? C������� q�z��� �
P�ݮ�w�U��A�4����Q���\��������`a��r����� ն��.U� �S�l6P��5�@֨���GS��{�ܤj���O?�� ������)u<� `�dJ���ǂ����~1۷�$���a�	��6]^�Z VU� K���bz3s��R@CrW�M�DC1�%L&�� �f�� c�� �K`X
�o .��~�A1C��� H��P&y*%�,tL(1��	 ���Ap����u�<�47��x3 ���>&�B;���uR
�@gs� �T�`\��+D�z���,����G$�� @�8vu� ���
��93=V��꼂`�������'u������� ����!� ����}gs� ֟$��}�v0&�s{ f(%�KX�� {���)/C ��x90� 2@t�
��k�� ��W�I� ��`��z� 5t�*�YH3�����a\6�ا� >�x��F��}\ .�</ yu�H��4NC�[@�����T3�d �=��p<��} v�BN+�
 h/�	ۋ�����N����7�+KT8P�Q[R �Ji&�2dX ��8�VW/9w�����u�6�HCs���q �X_4�%g ���8���9V��B�v��a'�GL��"�M  	@p<|�Cw{�R�N�H� ��&4cC ��X���G�x� >!���" jCtsw �)*�� �N;�G>�$��~[B8��5
6��E+�����o��N�;�t2 ��}iˠ� �X*�wSV�)�T���d� ��^�0 ����9�	@f��� z�D��r Fv�	 �\ Y������: �wu�Uq 	+��d�A ����`.V��> 鲱@B ���,�* %^�S�9p� �<�u����$~ ,�p� !���2<��~g Q'j>� �����(���w��TCg��M�<0$.�s|� V f�ب��2 �,.�~mK�� ��v��t; 2�dne�jI�S>� �=9ps� �ҡ�o�|al�$7 @�5�d� �꣖!�P���3�JP%��&�����n�� �Ήl|JG� A/'�������Oz ���+� ($-,�!�{ Q);�1o� ��T�tP~�������E�p���;�� ��$R(B�uM8>@��2 ���n��Q �������� E/
�Qw% D��$�w���!5�`�tg��w�} �4�����@ԞKN �� w�J�� :�W��؞� �9`��y<��! ��1	�q�>���ȓ� (�/�Z�� [+�5*)7D �A ~�S>	��~ ��+N� �����"6 h�f�.�CE�q� ��j�U� *3�I��0��6`��"�!r=F�ԯm��<D�[��)�׷Ш��';o�Q�ě�z���!2��N�0��C� �"	�4?S�`]�$st7ѤM_�@G������E�i��C�z�>�>ۀ�i�,��w P�-E%��� ���R�` lhap��kb q%ei8uwN��Z쐴�>�s� ,Æ�"bx _دElۙh ��I���;��5k���)� bM���� i*'� J�l�T;�.FO� ��Ģ>$$��%. Ԭ'� �LEW !��?
J	����%��U� 閯'���=\v�0�N�� >��r�=��'􎠱$� \W�0��4� 8h3u�U���m<n� qŸs�]�@u6zF� H`t/hTnx��Pp�'��� �(�����+zG���̻�� ��%�Ѿ�->>����*R�ڏ ?��q��� ~W�ހY-� i���HB��4@
��� �%�����G�@	U�(�M��XAR�F� ��}	;Uy �@Є�v_��p�]��� |�.u��� D9}�tL� ?�����	�0�������) 
$u�q�\ 5�Q�˃v�Y���A��`L ,@��uo�� �E#�_A n�@�ʼQS�������v �bu�eV�{)Ђ[���:rk�<����x S_�gs&�������P���s�`y+}� d���:T/$���9�Q� �(C\ Thfa��n��@ڸ�!�2���|ߟ���K��%k��� ~r�|=K{�<��5��Z d���BH�� ��K�Vu� ��ϒ�EPSXG� ��"�`'7� � >2�P� �i.W�� @�x ��Tu��� H@�g8� �a����Q`�AF$�#[���O* �C����X}��� �tB� ���f�9��ƨಊ~�c1��=�j��Uڿ�O�K��ƃ����`�l�t�<x( ^����R� w2��a� ��J *��������胆 �8`����Q �,d��&� cp>��� g�S;�^�R`�4J��ȅ� =�i�;0�yo��[ sL�tD8\ E��N#4)� f{@��<�"\�isP���� �L�h�'�� ���,R[���ܷ|@A�x�-t�� �]�IU:XQ���)�4� yݹ^�iZ��b%E ��)Xf d�KiP'��45��B�?�`ac� �pѩ��s ���h�ҵ	=5QT�R�Pp_F�$�a�t�z ��f��R) 3�0�B���4x	��z<2u�� 6sDt� ��Y���� ��Q+�fF��'�d�ǥ n ot��� @HELO 0Us> �i:th�t� �IA���0���<G�0���� 5�P/�L89�~3��I�<u�b�+ {\)���2',_p�D��g C�\��W��<��>Ǐ|����Z �L}�6��f�GBr�{��Z��]A+���8�MA IL FRO�: �[��NHntd&�U���RCPT �O:V����-k�����" ��U^p��E ���-�}X ��O�ue�D�M�»I`�X�;�0�
�0�Q� �~����� r�h���� %"zV�
m�~9��H�6B�? ��n���D AT���"L��$m�� ���~�8	�Su�C)e*�",�����-��l2x�/��ain;�churP$�=ISO8-@�59U1L�!�r��f0eK E��3dpg�8b V�=�"} ����|J#���r*�1�k8 ,��y.�:6&�J��� ��d�;~� �8��Y�i���`QЉ.\�yX J�<"�]
�[|��Bӡd�8� ��-^��i�=@}��J��02
,�d�Z����a�P�6|	�;J\��T_m�Ok$�0<H��}�o py�Tx} \t+4��]bG�P�u�$m��t�q R2p�r�<@<� P��ٿ���Hu�V ��� ��A�ws�M(�=��Vo�,Di�Z�;�;_�h"��� P��
�<�,=�@O��W� ��P_�z �}|Y� ^6I�B�ȃ �XM��7 ݗY��S� �d��,��!���M��:�h�����\ȬN�<���g3}'Ȉ U ���~N�C�����Z�� ��T�lhԄ ���km�~ U�H"�,���B���(���@�E� ���0��v2	��  Ut� p��Ji�M�?I��(��!� �<k��.f3Oi4D�t��û����" e^ŵh@xO �E���N��� �_�`a }CPUq�/8  ,�JN��xWZ��[a��(���u��d) �gMX<q>@�Q�O��HzJ �p���d ��E>(�� @�o��-��<��	L�XvPy>hp*�@��)�]���e$ ����� K����E �ܸ���Y-��n � [O�z ��+=�H��P ��ZE��J||�:�Yx����On" Qfqrm@` VgdKl,�OCS�i@&��� �ȴ,h�b' �l�-�QO�u	 ��ic��a(��Qb���
� �.��ƻ !���"� C� �DȨ� @�Љ�ԁ ����$�2� �8̅C� �d�5Đ�`������ݲ�ȫmG��Q\�q�f�uE ip)%x��aZ	dc(̅b�six<?��	n��� ��R|u�� $SN=%��_ rj2V��Y ʓ��+�3���MS���hn0���� Hy۵b� _������n�h��.�/ �pw3u� TSv��� &z�Wh`�u�0 Q�D��� �I���-1q
 P	D�<mq @k`?ϰ� \�L,���~�4.�x�[�ڄ Z��*�
K�x9z!.����T��pD �(/�K �7��}����6t!�G�������$@V�R_�Tܵ�`�F�l!�A �$8D|���� �*�v�tL,� iA��"�h�@7��,� ��Ȅ!�A(�p� �cwzV�
� �E�t�� $�.�W��o ܥ�&��LA ǃ=� ?� <h.�F� 7(P��f~� v!�ة% �j���N La��D7� ��̟'����٨�`��2��ԆA�#��� ȼoД�ω��~}�d�2�)��m��r6���e� ����S㍋�>9Z�2Q�;�&� �7B�1�z9��ol^�DV 8B ��Hĺ�����5T��Wd pqjlR��g$�x�H�cef A�w�P�G� 'v�=�[%;�]�����)Lx�ud-_s�Љ���[�Vy��� m�BW�j��?t S
LO�c��J@� _[&68CX�
 �	?Q;���I0̪D�+�Hd& C�;5-��#�bG��A ��%�hmK<��	EW�� ԗ�Y?�z� t��l$s�8Ap� 8ߙEd��:]����� XGB~J�D� Yu!��5?�j ��)���X8���(+O�[7ɝ]*��;��q�J#}�� C�f��Z`�JX$O��Ԙ�%S�
��W�ks؄- �9�JHA�ڠ@�6�. D���X �8�C��H<�0�:�,5�*6=(4�;�H�tr gpCbw�d fm(
he�c��+��@pn j`He�uh:&B�zg{�`M���Y S�V�d� \G��%� �Z�,��� �����B� #j��*%��xD���i�R] S\zWTZw�0�d$q�~�sv��P |)�ox�$���kޘu (q {�P*V�-�Xp&/�"��dَ� j�S}�f~\�I	�V� qJ��H����40eosV �L�ǡ�� ���5�2 'k�Q& s ��{�#+x�<�邤)4����� �U�n�X�r� `��O]�[��tdc
���� I��GJ'uS{� d
�b>B}�~�@�/!�&� W�d H� @�gI���F�XF�]�S ���K��+���y��}�Li `nh[B� �'�1RW V95�Ȉ��_�\�8Tไ��F3�Aɀ�-������2�p0�\��:� � vELP7�Y�P��6
 �B*p�<\ ��X>�|��Gu�-����D� +�\��	e5aW���[� mh��P��p o�C��� �z½}Ǵ� ]q੢nBx ��T^���[=���D:�[��3�a���6	u-��f�8MyZa$�x<�6 �p`�h�� �VX#	�> PE�Rr%�.����+��������Z@�KM�? �e����O��b��
�[H �9xI|<��;� -y&�( ^�A{�*�b�g #LGMc�� �p;�s�3�� 	� }��if����L�����}�U���@� ]^<��- я
�G���1HVB<�-�`,� t2��{��k���V�0�[�-%��@o`�4��!�>���G� W�|���Y *t@:� �`U�wE� (~%ה�=����2 t���X�_ �<Z*�΄� ��L֠1 ��q�Y���[r@ܱ�_;�ƥ�<PІ�`��¾�\�_�� �!��a&�s� P�jɍr Q�}�*� EZ�w'�:g �	ԭj4�q !��p��� ��u�C� ���?�
���T@�%H:���-Ϯ`�_���p���0�?Ѿ�6!�a�HX T_ƹ��� -�D��S1�|]�Ԕ  $�Df9�e P�(�3M� ��?��+` ~C��J\N� �
)	UOt T�g��^=�� �����\�� �Bj�, �y=&�� �Z�Ru�M[T�Ǥ���8\ �d� �Ļ;�K���(�� �Whob�� �'YED�Ʈ򌒟@R�ԈG{�=�� ]*�N��?�	 �����; �u��҅ x���}i� ^�et�dB,�C��Ш���9��S�] ��;3.5R ����� b%T�kh $e���	S ���qD!�� �yL�8lQCe���XS�D�1�R@���� �I�ʻ8<�۬��H�+��"���s	�#�����Iu �1r�-ڀ�w �[��Cщ���U`�ȇ������<�>� \�y�˗כ ��T ��^�`�\3'SYҭ�	�h(k�7�R�܅$�#��@��K� :
.�BIu 𰖦�>+E�F��@�A���� 9B$�2f�?	%���d"[ �� Z���p�� 8rU�&��P<����@x� jX�7�} �0��VԺ� ��fB�	� �UK̘�_��:; �u4@Se���[����>��/��=A�H+������� LC��?�?�sO�F�;X���W��]��I<V|K�D��wHT��_з\�t v�W�h@#$ ��"�Y�}�y; ȹ	���s �.��� �[�2dQ��}����-oax� %Ð��R%y�j �s�I ����1-�U u,��j�,A� �(��e�, �' ����M]D'�N�@�� C&4���$y�PTϨZ,��Q���?�X DgH �s0 �F�*ӌ� O%�L<�� $�y	�"�+��uz�/ C(����  �0I���'"�]�і/��i��w������x��� �Y�^�kP��E\�t
���,��(S��X �bx� ���C�*�HJ�B�Gj@;�
W \�A����% D�;�$vs
HP E���� �N�eu��a��S� ����H Y�$� �F"��@� �2w����;�r�l$E `�vF���/���t�- Ҹ�Sw�����}���͈� ���WU	 ��+Qϋ�~i f�����u	h\ Js� U�k,ru�M��D�܍> Ƿ);ؤ�����Ee� �R}8Z� n���l��b��6���´Lu�`�J; EKԿ.#-� G/m��� |ի%�t �l��m"n���(���Vp  ��\�Bl� �Dk��� ?'�v�뱛 "�_��r4XI1 �jd���q[Z����
�)r����^C�n Si!�׀8 �u@�. tf��Z�"J ���%uP�	��� "ĉ� S��C�;uk t�ϊ �Ɉ1�]X�-��I��h�=��^	b����~��LY 8Ġ253� %ݖ<��	� m�Ky�"�yg ��d>���6�s��`4��0��`���r[ j���lNu�W��y���ݵr�8Rﰹ/Y� �n�;��� ����j �4��
�ֆ!�uLK h%� :���.�X� ��$�pBZI =���|�8:��� �'^@bÁ�: ,��KX�5�m�&##"l �~[�� KCYL��`�D ����5X �H�P9=<U��O�"��`� ���x]Y�9	0W1�����d`�6�IB�5�>fN�D�% w^ư��
u��0����X�=�t����� ��n(����h�ջ�� ����p/G q���&�� ��<x�C � �%gN�GJ lH�9 W�3��D���LhS`z�;,�@�BD8uL�Ww�$@:�c� mH���2}�3$ݏ��@/�7��6� �\1�`pD�ah�qy��x N�[p��� �K�c�Lv �D{B}jT gA�V2PoI�aGet���d ޜsp Rai ��Ex}c�y?�	�V�����Sm�6�1b�� yA|�W�ռ '���.zC𸅔��g�J�b��x��u��B�r����#����) 0�vpI�l 	}�"LEd.�=r��2���� OC	f�?��96�)�J8 �a%��:� ����=�r�"�@2�OtR&�� v�,[� �T��+ �=��SvH 
�R�m�� ����'P S]�r(t
 h�sn	�+���C R����t� Ή���8q ��^�}h�GB�clx,�
�F���s�6�8� �O�B����V��K] ��"�P�h R����=��ע%�����]}� ��ʴu�/�{� kw�����&?86���2@V��3��@���/t �
\���B�;:��L�T��^��p z�]d3 !u`��c�PsO��@%�� �0'�f� ��<����� �{u��*A �$RSW/�rJ ��Ԏ{<� |;x\ �CK
�_�4 JD�Fh8{�ی���/@��� kF|�,t^�g���h��г��> E*�4j�5 otG��[� ��i-p��~ ��G�����u� z�i� >��<һpD The��Jd �+x�E2�coul� ������a��~N��c�y^m��f. k �Y�1}LOq �����{V�) d�pY��u	�O�V]w�哭 p���IV%� ��W���-��p�t`�K & ߐ�	C ,vP{�� }����u^� ��݄�� ��aR`�}�����p?�(ȳ� ��Tk8W��&Xj� K�х� .*�7�6P�z��c>�`s�og��@5��t	"	6�Έ7��9&�]g
���"� 	�uԘ�  M���&U|,<�i��k��TW$��(����dB(��Rk��b�v�� f8�B�� h:Ҳ��; tU^�a�S �H*�e u��J��p ��� �;�tZ�5��`zQ�N����(% �Y��|~�[]!��w
90Q� ��\�ٗ ���#x �����'�e������0@ohE W�%� MԞ�neFP�� 0R�IxK O��	j2� �bY��4����^ Ã���� O�L�גp�jS2��nY�� '4-@t�	@��Q͒����`6FH�p�<
+�L 菩hW� .�G4@��;D T��Ʊ� e�:^7u	��[t������e�.��a�8 |��nE�D9u&�����3��� �c�By��[G�a�R� ��S�d�4���H`�
��^���;8��Cy���̧�En�����8േ�zTC5�q�!<Y�N������0e�q� �Q	�Ĵ�4 ����k�xX�� O�'c8�} i{��ok*M���b~lth��؂a���������TZ�+�F|���$����Ovw	GĀ�~��?|B /��9�� @���DNi��;`��W ��a3��;�
�	_T��,����v %�!Z�? ���Bx�� W.N֦�#	t~ <KRB�%� ��ι��(�jH���"_� �Vz����5)S���e?0�� �^$�v��� ����KC�V #h	��i&;2 *��j�� R|�A_'G�F	� �����I����+$h 7/kԣ�J �w��n$�{��wb ü�C %���/�` SR ��C���V(ݡ���:��H�-M Xξ l�sZ(�O�*>��֯!�p���;� U�:�б53�˰��\ !�}��x�ݨ܆#~�����Q�>�K�_`%W<'�Y| ����@ B��
u��͏��D@>� Y�I�v�n���ӊ���!C �CR��� ��\��$�4� �X���B ��溵.4� �M�a&��r e�k}�x+^'�j�?K������"֩�@��-�PЦ �p�wGHbq���ư JP�3�!W������c�x� �	]{@�� K����sOj ����[ z��U
$I9dS�_W�e�p ���
w����������/ R�ߔ��j�.�JG�]i�X�� ��:hZ��\+0TR�ͤ�B��, �OZ'��� �j�-ޜ4 C ��?^ �B�;�(�j�Wl��)[Xr�"�B���_�@��O�
K�%� b3cG��ê�P�q+�z �hЁtY� �l��;�0r� 9?-�s�7��������
����@�Y���I��X$��;� ���m�y�7��`좇(^|F M��]\���e� 4)�%�.O� �bJ'H� �!�B����X,>�1���Q�� �x&~C�ra�4�
�� �+�3��D=���U $׈G~�H���� F�����	E�+� ��n�`ԕ�����-=R�&wf��� �t�@�O u�2�Ejl9 h����u��v��퀑��l: ��z��q���u0�0�Z]_|p��7������ �>�#�� ṵ����T ��M1��Z�@����8سC5A	�˂4 _\t� ����|��c ���K5�� ��C��' �-�dp	 �H���"�D ���� $3H\��"�D�튂Hj� $�aG� gw|%i�� ���ǊR' ��vX�ܦ��w2�|*�ܛ)�NSvۭ��%�'P<����R����@a+AY o�7") ��f�SF8!��>t+��gI z:�������d��� R(�? �;��b-� t��� 0�Q�*m��27	��E��� /;�#�&X�-�:��RNԍsK���ǨF��T�@A��Ҕ`
! OЀ�ua7�������L�� 	z��~(y k+R<�! ��)z�\T ��'
� ��	Y@j;��wN���(�D0?�K �*��� m5�|�� RH&��EP� 0��)� $A��QT�e� 3w���〒d���\�\	�x N�_�XT$�ԀC�"�|� �����{Bt �C�T3� &\�n��Q�-?��	t=� ��a��y3 Ln�gPho� ���A� zk�B��j�E���A �Sokد����&`<e 1S@XHh, �{K���ܨ'�M�;G w��nB-�9��`@郿���ݶ� �,NA4߀<���Q`@�t ���%w��?c� E?逥I ��^̛�cN l���D� ���]Sx��;0���z�mH?�2��R�t!s0�{���4)EW�7+���hw�$@炅�v8j���@;��� �h-f�t *���">1��x Os`l pw�h�M�d��� @�XNP� S���?��* Ń�s�c@( �v+#;{�8 ����K}|J='���\�A0��tc��{lvd] W Q@K��E�� k��Xm`�Uꬅ �t��֟� s2h��ʵr.'F��M�� Vw�S��|�"Ct�� ������Z���	� ج�e���~ �����g��=�,�S�� ���t$�x+��X@��;�{| ��w"��{� ����^� �蒴؅C���?�3�`~P �J�ر���	��Ђ��;�V������c �9Htf
{����ú T����Sd �tل!�� e$K��)D 5}�B0 48	h��� ��\2��1 .�} qCa n'txe�d�X�V ��X�S�6�B(T��!�� R���\�h�� D��8;����2#��P�D�p� _ذ�0� ����/�  )��T�� G�cǾb�2�D H���% �W7�f1U 2N*&� ��m^; x�)HA ��pP ${��~�?.�R�^�$�����=� ����! ,0�4I�D ��J�Ut��L�U 6+�@��� ��铀��� �K��G� 5	���L4 ,���0�u���	8 ���`��	���J��K)���͵� 7,"04�8$�2�U��A�:� #��«?� 3M*HW��1�V�@D0�� N�I:� *�b���>q݁)�hP���C T��U~�A� ��*��"��,a�$��,��}`��X �L�CZ@Rt �mk��u/ ��=	l�h`Kn��� ���c�\-�8k, +�n;� t4�l� �p%(3 "N�ޕ�$�_���,�`<�&��w�Y��L�� W�}��%~#�E��� ���˴�ҵd��a��+����w�� Z� ��� ��]ȇU� �oМ���r9V�K���%�שׁ  �e�}�=������t��)(�R���D �c��'�7�_t�zʁ�������$)�x�IЪA i[{d��Z�	+�Tz��D0(� \F�:�W�� �=�����<�ʀ[伪�; Xs
hL�/ y�.���10���kQh���V��IԮ����|�`#
�Z=�u��p� l�\�!%�v� ��,`�j� be������ 
})��cY�j�H��zH���|��p�5 ��2����1�L~�@��� ����*�����ۄ���$�E����I5ؐ�V%����"� �+����& ��X���v�P��!t�G⤜N`x��J@ �Ё�p5Cj ���V$�6Z�� W`�G\��~����/��W@�� E!��w�h�C �觌8=�F����R<�D�l�Lji�J������C�� �pX.t�h �Muԑ'JsQ�� �Ơ��G  bF����A� K����` ���%G\TL�)*����O���G������o4n>з �_�=J�. ]�oQ:Bz�w}T����%� ��,X� 4�����W�3H ]����#<1S�0���D:�R4���y 8!�1�(���� � ��a;�<��C7N�@׶��� .��B)^� ���M���ک�C����Q`xn%@|*'ޓ� ����������S ���P�:�T �B)yZ�#����`?��0 V���%�M 떮"u�+ 1Ѐ�;�w2�  ��?u� t�#y��L�<�p* ��A)�٢ G8JY+~�9�dF��Z� (�Qz�p� �X_�l�jA <��&a�z|��8�7���% �wΡ[��� �(��Z�5	u��'T� �qP�ҋ|}΄���T�J X]�;�w ^?��}�s ��+Э�4 �f�܊
�  arR�zS��W!q ��w� �u�+{K��m t$I���;��	W���@���	ّ�p?��'<$NHc�u"�D����:�_�W@W���B��i@���`�1~�y�<7t�/=�$�
1�W�<z����B"���~����<�)����P�>�dp:`X�C.�"���8����| P��С� ���RH!�c��pKL���.� [��]-w� A�Bs @_ӱ��֕���I KETW N1!��P��U��۝QþX	��Pj�WFSU�`D?# ��m���� ���u ��J�� Dw��]� �_=��$� ��Iw�� Gʤ
�H �v��!��	s�  7��� 36,��:$�z !2��D��q��Cj ���BH��/�q�(�15 o��%2&�| ���H�w\� lY�<) �$�eu ���h�K� ���bL`8P���@��� ��[�� ��Z�wlu�P�� �5�xZj� ����hJ��$X��I�P4 -���7M =�x<�3��
>���'2 A� �)� �����]V ��;s�P B�����y	CXt 2N�-��T���u���XM@��9����a&'FU>`|�* ����V� +CIT�e2�i~����]�^)��6��	�l� �T��i(j$u�P�����by��C����1���J�s�?�@&���E�
I��ٻ�P�� B9+lD 
��"R,��|�S_��fsN�AM�@�>� a��ώ~�� �v
��&Gg 1ɿ�(�{��Q�`bLE ���G����ي@J:�� S��$�[&����X7	�σ�P"�xW�g|���`!�;WA� ؟,� �u��.���D���H4N��!\��Р��l�;�� ���ѱR @��*�S«;"K�u~����$�� /��-�K���^��m��>�����w����. ��4A�	#rv ʪ�y?�>; tH-�{s'��Y\���[��Z���h� �-�u���t3v #4����� ���׺5� ��~ɖp_�L� B�e�'� Ѳ"�S�� ����D}��;�ȸ�J0���=V �6c���P �Y�����.aq �k�:�Q�Ԉ¹����v=���B0�}t� ���b�Z�L�g �T��� �!Q�$k�^Z��2`�DBJ tTK%u> y�7<[�]	�����%I�� ��m�n��X���]3@� m%�P)Ouo��R�i�
肈�j��H��u�t!�M� �#�,���P�E���']�w�p}qR����0Puc5 賕�� s��o���p �k�Qub^�\
�v!�`z�ܓ X�5�?f$ Rq��4r�j���z��+�����܉ ��LuPg� �E��[��sWl�	_�|abO�/�MșV L�X�|Z�1 ��{�F�oMu@o �h��_�9�pF�� B7#˯S'�4�o.�Ǭ��`F� u���G������$l��P� ;���}��K[�̱���UYXO��i�� �d�2��fp�����Ӈ�C���=	�Q�)�r��p<� �6Dί�X$q	������ :�{i�Z�g�qf ��;A�t��� -�! �Q���A�;��`C���� ��:��F���e(J�ڔ�;V΀��:^5t@
6�	L9 �xA]�D� ���4kG@��'/� �_���<� ��C^�y-�W��p��IO��� �H� J��8Y��?.] ��צ,�N9&��O�}�� ~P�%V@��E=�c�	���� ����DOP��U �X�e:S!���� Ϣb�
� �ʮI1�;� ���./��r��*��I !��7%�)?�> =�� h�*4B�K ��_
$s9 \�V���� W(�<�CԞ �Њ���{� �Sw�$WHu� ��I2��� �5�\'�T ��F~�}w "ud�NSR� ��9B�۽ �w�Y�j�h0�Q7�k\U Gi3�㾄 ~a!��
����ȍ�C��W�]Yt�e )�	�@�HZ \ V�8�? b���Ĉ �s�ѵQ�%�p��̟� S����y�k��a���BY� Ľ/���y������gvB(����9�/�0�r z$!�Kg� �ș	�� �.�n��.��j`�_a /�IA�������,��G��s��Z nS$���'�ŀ���� �W�S@� ��@:O��� 2_)���� dx�3j}
�� 9��(� �CT��v,%�6 �t�N&� �;9u�c� �)*<K@�k`A�"u'@�B(�2� �����
զ�1�_��$� S�)�ǞМ�RZ���'�^ -@D<7C haB;�+�m xG�e���� �&@HJ�� �8U�u\�~ ��G�f��!0M�@� ��%����M�b���`�o���l��C��i�1Y&�\ �M���/��T.S�$>��qD��t�\/��:�~�y��H�q����,`�ؗ�8ir��\�z^�Q�q.�`,胨ꗈg=���/�@���r�HwU�سKʲ�ـ����� �_�n.� �g���*AB �P/(��9�)��E�!#�{*_�:Yސi��� ���D��� EWj� @<��: �.m="�(RzO �U߁j%� 
��m].- Ŗ�K�+��� 3X�B�T� �2��S	 ����N��u8 +�����x�:�� �F��0];ܵ��@Tbl�gR�� ��
=�B��Q�� �\����D!�� {@�<�g���j��b�n� '&�W����� �<Ғ��= �o25+Q T�G%Zݰw3 �?��J �B+@� � l=k� ;�&�PM�<7� ��QSuG3 �\Ɨ��� ���+ t��Bd�x;Wz�ń��L�� M�L~�{����	�p:$� ���&�R��� |+	C<�� ���T&!Ñd �	�����n ʎ�C,w��	;��d� �F�Tw��' $џ��b�~U�p�z ?�ܰ��?$쀥�}\�Jr�#4�|� P�j�: ���80C�S �g�-+]<�B�����s[��, 4����� y8!�oP� STNL.F}Jǈ�a�PW1	 pRQ(e� *��^����� ������ ��%,�:�� (2Th�	��@��u%҃��6��ӕ� 6��
 +`B@�7X0�2X�Q� ,ψ���[ E�����u��f�b� �6)�����:CKu�O���� j�=��;�
 �����T�-OJ��1�S�$� !�� ��d�9U�?>5�����b�7|t�����U�>�>;�r���s��*�� ������֎ ��[ `��bLJ�N�@�웭��-���P�i� �_�(!��3����P������H~J� t����� WDu{۔�( ��7�.t}��5���p�o 4���b%P���G��tI��w�n� ���4;!�;Q�G��@�t� ]���� `2$��E��I�G�㥘�/� ;�J����xp �!�{�Q ����	�[>wH}ߟ{إ~� U'�"S- yI�%um�^e_Z��j�]�' ��RB�W� FEI�U��~ �'na��s���#�`Z�{/ �?1[�Xһ �.$�Z�V` �OX�����`o~$!zK N"��V5 �	��\�I��}�<q�Yf�'* ��CG��#��U��ऌ} ;�%�p ��~�v�� ��o�xu �5k(lQ�j /}U?����d�)��; u ��R�� �I��b�W\P��<�}��<ѐ��%ȋ� hB��Y��5 C�QFN�x�� ;
u��P�Bn � �t�����ӫ��k�}H �%Ufup�� ��3��� ���;�{ 2�CVN��t"#����� }B%3n�ms�"�X�eIQ쩿 Y!i� �B{ p^��J�P�w�h�@��V����^W��kE �r���ݤ guW^xe _�3��� h����/@�S�c!xy��H�*K 0���_� Q�ݧz *���I7� ��ĝq �e���2Q ��щPW�X�@藲y�[�(d�Z�0�OH�X��Q�/����8Y������ޠ�D 7� =���(we 	0���6�$9�����Q���!P�q o�-��:O �m��Z��
D��&�N+O0@�!� Tk"w�� #�O�3K�}����P��h�j�3�t�q� �+���A� X�$�sH�� YS[�Ҩ� �T|��%� ��§H!5���h<B����� �N�*�6? ��T�EX �S��Jut� (�7�P ���2.?����$���	�6Z������1�t5��8IH��6�@�����
 �4�#� lŞ���:+�*���=It�'րʄL:�,*� ~���R,� �j�_W�&`NT!����h�Bg�ee� �:K)I� rԵ%���f9�ȴ���d �vpi��uG x�^�zH���Z�ǦX1@+h��T��f���AP-_t�� K�=� ����f�G F�MJ� H�i��� "{t͈@l� 
��d����� �^��@z 1b������Kҿ^'�@�Bi �PQ��و=���U�V�s=M(�YZ@u��H� �oҲU�c1�L�WP�׮� �	\�.�SICE
t�)�WV�D �]�0�{��mC�)�9�f�
BG"Ƞ�� ���K^�)xp;X��$�ǘ����Q�� �:�l�߷��wu"�p�),��� e��[.=:���Vh�K����"�te�ש�� 8�V�R�&�H\��g�@�yTJ'��b�j]�=�*�`�:�6� \I<�	u %���S�A �E�W���X��	C .-�Qܧ� ��k�Jɯ (\P���f� Lg��G}p���q�| nɄ� ���̈�|��_�� !���l�uE�$J������ B�����. p�_0# $�(m� �������[��u���n�Җ �,z
A�=(�� ���\�߮��?K+�%���,1G>�Դ�<|7�;U z,-��X 8�^�BL6��z�S|ajNSm9����J� z�_E� ������M����4,6��k�L�Q��"�o� D�
�8O�� J4�`�� �3P<N�	�u�5��@��� �y3;�	(�.��U��H���߁��@�l6�	��@��4 +��t%� ��]�m���8zV oPR����&8�Iu ;�j ��C�%�p~qf����0�}`'��A��	8	�V�J &T�r�R�+�#�Z� ���BD 2XtP���^��5W����i���FZ +�C�������8��	�밀-��� ���(7)S6�T��V�{�Z�`�H%�+C<� =0�f:� oe U�X �9�W�Ks� 	D����� ��=�E��@ ��)�.��� >J;��\B� �}�?�����`��2�u�w� >G�8D Q���e����1�n�C��� E�Y�I$8b�<�����</6�0X٠�� D���"��� &_3��:� ��$}ʟ M��U��Z `c|hfP>	 _��8m�� HJ�^�&P�� $�k�A�F���0���D�^��Y� `���sw=ؽ�_���%�a A���' 3�1S�݋U \��2Q;�:@ۃ@�[��d �TE�Q B��2� ��hd��3� �(��@��8 �P�V���LrG *Y��!Q |@���7xH ��ǰ���o��+���
蹺8�� Y���J$}_����z�G	 ^ ��'P 0�j������ ���+�4>�� ��1�!��A����I�[���O�g&v`$�� T�}Uӗ����+פ��,]��K���|�u9�� �i0�M�y(�� F�gY[VP`�;��h���>�����6|XIP ��5{e����\ ���zC: $NɥcW� X������ Τ�p�d@ �|DNV� ��:a,�X ��3|�C ߉_�(�S[��0����T"� `ơ�]0� R-�Hs�2 8��Q���7�
RFW�c- TC�A�� ?�߄�:��Lx�$ٳ��� Qϕ���B ����`G@��� bw�>�[���y]> ���@��~ v�S�D� �Ux%o�������D "`aqMW� �S���3�����"��Y� ��l~r��X D�ċ���K ��U[�z ?*�+�d ��׸�_Z��< :MG|� B\5Rh`��	 ������d&V�K�q �Jl?��e ��4E�g�t ĥ�1�X�� ��ca����`�I3�H�[ta���aK��
��X�`�� �Z����� k_S���Ad �Tw^�%� L�+8���8M� \{.���0����aT�J��	S8߻ �;�+ڐӰ�/[���8�(�b�pFM�]�b?��0P- ��)#é @86k��Z y0w�I��EW�'�JG`[
��PQ� ߡ�_ ��؜��[	(����^I=V���0~2+���`	�w�)����VU W��n��^ AQ�����,8��@TW�� d[���MF� OU�^`� ��>NIƆ y�$�_�` 3�R���&} K�+^F�H<���0� YX��$g%s��Hۆ� �	���� �_�7a��E 3���c� >Vh%A̾� �7�͏���� (���b� P���m&� R{���6��$q�|�����v�� ]��[�~J�X �ړ�Z�)��|�gWH`��l /�����\����Y��|$ �Q8h���ޠ{H���qP�S�T t���`C�;�	���?
�R� Kx��3�I��� ��h�)� j{��	ڕ� H��-�+R,�@0~���| �s��Z ���d��P ���1�ކKs�+�������(i	 t׍��g 5
�4� ���� ZpL����� �X�^�F�� 9�p`Q�G�X��Z�؈mY ��Q+�%� .���-��p��<��J�>� x[�5�;�|5���o�� ��BW�|i=Đ�r��U`To ��	�' ��z$κ����@�P��5 �+ְ!� @�R��	����S��U3?�[��Bใ� ��5��������=p ā�V�{(]�:\� ��,[��� +zZ�@3A &�J����a�ؠs���-����km��7 '@/&3g ��Z�X��� �=C�"	�p(���@��&FD�%�>�b~ �r���$ �X��"$p�@��N�� ��֟(�U �{�P 9R/�� 1��(���z�jRA�:�Ӵ���;Pc�OV쒝 H���F��G��U �vJ��n��uX SPWh ��g��l� �+�ү�D rW$>�%FZ�H� )
�)��P�@	FBID:�3@ßq��+ �r�X[^j�ݢ����8����鸒� �XEZ�58� :G���� R�EB�� �(����7�<�w�� � :�!�A O�&(�tK.�FD0~B͋ "#W�c ��ο�� �[)�qy �S.�Ÿ�� ��-k�c 2~ ���_(y� A�~�������C�y� Ln��ξ�� ~퐓�5� ���S�u�� [%��@�?U����I
	h`خ�s"*[� �O��H�}�<�( X���2����!C��  k�|VSW� ���x�1 �	�t9�7� <�ւ}B=u ��EI� ���}Zt� �:U�u����o�)��� ����O�� a�Y{8�� 4k����v !T��C�Jw��B�E`� U#� ��lu *���$4 (W1�%�|�>��x ?(]�m ��=6�� �"V[WA�� ��Db4%� ͠�cV�J���^B ���I�� �`o��G��x��������� ,c������]�UX���a�h+� 锎�<�� %節�� ��/�6] L�[�y8�� �^����5 �m��+� �YМ�NA�0_p�?b' DJ��	G}&X^S>��;��07�z91%��>U����g�H$�
���FǾ+�&�"��C��΁d�Q ��W@�6>A� è�+�� Y��?2l_ 0���^+�Ⱂ�
]��i�rB �V�$د �K��}� Z���� &��S_�H��L}� ��ݮ`nE�I����`o�a� AW���65 .PR`{) A
+Օ�L,�� }���B� �JA_j�H 3�P��qD��5Z�`+���M �#nk�� r�Hm).(�*\�z&�p��h��,�x��~� >uV��	+s8�� �Q��eJ@�k&�|z �����o��HP� Z�Y�k� �(&�3#� ;����n� ��|Cu� ��Lk��?2�[>�`���\�4 7��l� r]�hֵ�}��G��d��� V@��,3�6B����^�v ��F�L)?#��5�@ًƚ�S�.�PT#�� L6��9 �<�>��v, #+�X��ޯ ̶�S9�w �JϹ� ���*�2k�S$�Q��>����~ J�(��D�P��v=s@. �X�a^�H���H�*�� �<߇z}{� e?��L'js5 �N�`t� =�����Gq��އ���BF �+�j_�Q �����N�,ж`@#�h�k���
D�0�B$ t���Nb?,/�	��;��*��ikɪe%p�~x� �" ��7�� ���Z� �-����.� �R���<�s/ޓ!�ׅ� �9��2 ��ֽ� �- ʞ#�B��7	z�D�2^�}�a ϵ,�W�#��T�a7��0� ̑.V�> ӀI9����@�ʘ�� _
Ip�B�x�u� ���w`ٹ� H	���Y ��,�ID�ZQ6֡�aA�e�� R"�ski �
KO/� �@^���}R%���U ��=/��&�^b���� ����7��$k% &i ��&�L���\?N .���V�� �/v��S�����G� �R�^�N$ �&�*~c�� �d[��XG �`.!2� �^zT��'��]`��ǠM[�o� �,Z}eQ@ �Ck��r�?암�0_� U�ֿ�Y����	�g� K�iuH ��'}�. ��݂�# 4��R̐Si	�p� 
��ԅ~D�� vnX�.eI�� 7�0��	�ACF�/6����&WV���� �~��:� �2��"< D�^�uX�f~��������SnH�  t�,<v�h\p_���Qo�89J��;�& 1���+A�r C����\$�wY�( �:�_�� �%��`BG��bW�uZ(k��� +K����; 6�
���< (���B�,y� ������"FTd �� ��N�B@�t!�׌?5(��=����&`�8��?� ��:R�� �)�,����� �
�&� c!��B[a	�Z N�HDt�<' F�D!m ������� ��۹�7G ���x��� �-�S���� �
������ԕx� A�T�h �@ģ�LS�>�Z��@��( @�j&���.Qa�  ��h ��"���t:^���O_��HT f�vu�� ����z�LT:%���v�݇YS �����_ ���`A�+<�v ��7��2�S� 	���{�H�� D��H��8M� e�v[��Q0�+rpZ@s�?�J�שe}��v �A0B
�:+ C�YV,|b� ��@D?�� 2�Cê*�! %[d��V� ��W�Q��{ �	�\E[ ���o@� م���-� �UT�	t^ >*$H�=J���`�ۊ_�V �5նIW��&]n� ���8�XK(���E�n���_�.��� ���wh.PV� �2�?��� 	�-xlR $�<�W�æ�>�����~ `Y�&j� M �޽� ��%�N��� ���R�y �x�]b|& �X�L +�ȫGl?�� |��X��, �$�iyE Un% �ǿ �(巇߁���� �����Q-�zB��aJG�pc@��=l����Rf�`	i�4A Tl?��EZ� o�r	��~�B\/R ZN���q �st��d�9���n]�$� �k�{Z�� �X�<��sF�� ��P]V�����6�����q^ ��k�yR�HJ��J�a ��>���l w��}�.�X \�U�-��<o }Q���	R�W%�`�*Ϯ �7#Y H�2G��L�� I~�q�v�9�� ��.�y&� ��W��pAZɱ�"� �8D����M�}G��Q��WO�J �q�G��V;�F Y��_ԋ�n�X�0Z��WPf x-�ɍ�0!|<�-��AW�p�� �N|P��� ,��o�< �Ҹ:>��x \�����B>7� �*=���Y �X%x� ���V�E>?0Ԁ+Ө�B' P�c�`�X�i��*�J �fjz��%�&� \8�� �>�J�Y�`0LK�_6 ��[�%ӈ� ���M�|C� ��˹��h=���.�;��ų� zdG�`���� �J�wtR��� �*�pG�0L~ �'�+�| V#�k	�rFu�;�އ偃� ��U8�? �W�v{��+ƀ� i��_���yQ�<�Ů0r�bIjX0� @l��LP�?�,�9�&��! ?k��:K�� (�%�5A|`�WNF��_��o�A����Z�8��$�KU�\Ƚ�����u �v��G� �=a],3  ��/ĹZ tv���4 �h۸i��� /z��B ���ϭ� @�eV��,_�[�.���JKl��� ��d0�� &\�<��� 3P���y� a^Ⱦ6�;{bg(�O�7d `���������� �����sQ� �8}IZ�(c=T;� ��ſ�S ��Q�?�V-��\I �kc���&d����( JW���w��x��*�	pMR@ �N,͊r��H�ڀH�;(X�� 	BC9�X`f�d����.у�?�B2� ����#�] _�ڠe��PE$�2���Z �!�X�0 �އI�W�& 	��Q� �Ƹ�X�O� B�*��������@a�� 4(I��r� EPt��ٝY��(\�_Ӑ2�	 ]dR �� ����L�=6ƻd��0�my� �����	F \j�v�Ie �,^*.� 
) ��]p I�v'�XQ�5�$ �� ����jYA �C���� h��}G�:� xJ���^o '�>�!��8T� W��k��` �4^���/��m����@�	ֿLf�&��	�_ +ޚ���	PBm���kp� KZ�Jh�e 6�|�]� �X��0��c #ު�k�  u�F�KI ���(:�ŤiG
�Y�R�B���;�Xt9� � ���� �;��G�u!	��n��6��@I�r�%u 	w#���O4 ����פ�*{� xw�M�t1�I~N #	�C:'� &�8V;�A�<$��o�f�^��� �*b� �E�hL� �d4%� "�j*C�}� ���n�[�Z ����M ��	 Â��� r��I3�v;���Y$���VzJ�0� �d��MDb0�S� ���ߪ�#� +�6A&��TB��s�}���� ���KA��> ��M�+ �R�� �w ��� 6�,�Q���
�I��=�E���_��+�Ԃ=B (M�4 �$����� m�SX&<���v��P� �u@���� W���/]T<+��*IVP������eh� �������_� �X��� �@��  ����_#B� ����QiT� J8�+��Rf/%���X�e����^P9a	(���� b�GK�0�� �J?�@:� ���� �^%cE
w���@ j�U��nY �[-�	g�$� �aQL oqP -��&��<� z
��A�f D��[�n� -Zah�Y�k &/�4'`� P���hQoK XW��E}{N0�*�?��/ 3/�� �5��8�ʸ� �;}/��G� unQ�t�R��@b����*| �Q�Rp	�BH
�,T�� P��+�Zf敡�-�ɻ ��w[&���ۀO0I�Y W�<�� 	&B�q�f �V4�� �Wi-�&���~ ���+�	� U`.Ð!�'��ϣ��)\�� �5bk��^�x�Ɲ� �+|�,^�R��G�.A�s�x�����n��.� R&3�� �N�H��+��}Z�]�� ��KL�Q�ؤb �:��Zw�Yj��� ��?I~ �\4&������P�^��8�_N��� İxV�� ���aG�Z���^`�l �QVh�� '��i�8x���V���c ���_��� %�-��r�6L�V�Q����mY���C�Ё2�s]�� LU�cƑ����.N#~ �ȂVC	� `l^9��Z �Ä�����@O� ���p X+�k�ghX����w���,�_����$�y�8�= �\:+����D���m�� 6yK��L�N ����h�s�H[5_���p� ��a�,�	 ��l�%�� ̎��![�<� ܿ<.�Q��� o��XH��h�UCY���p<� �e�3��� <;UO=QmX� �	�����D��I����+� ���E_S ��&=[�X� ��G5����X���w r�+�� �k��9X�@�@�� �+d��(�x �Չ5h�� I�%p��Ǘ :�r�	�� �;��-O �3��ύ�vH�օ���t�����4�(��< �85��` �7�60 *A�h�!;�Ѐ�p�߸ ��P5�N D�ϩ�*1�i(@}[ ԯV�t�J ����÷r_ �v�Y*�� ��8J�� �H���_)RVE�f�[� |s���� 8�@�h6v2�B"P�8�wsF&
�fZVT����R��M� W&�|`e�	��7� �	���~�8�;�/��I�����~����o�}����B�=DKk`z���];^�3݃�����w��)h*=�0R��I e��\T�Zp?������x�<7��o�n] �b�%9���	E ���A=)��}v�ؽuD T�*��?���K@Z0���u���N�<��|	Ge� ��Q�\~2>����kMs ���1��Vv��n�B���x j�Π���q F���a� ��>�Q�ֻ�h܁7�� �F �`޳�Y�& _���W�Q AN�(U�,T ��Z@6�D� ><�ђ^ ��u	x'����;Dr$`�{ �]o�-3$;l thD� z�Y�R76:� U=o�q]%��8��\a "����P ��uAR�v8f������ N�(�#�H\����p]i3�����T�kv Nu�n;�� /�\�%U�� D4�L�3���Z���ۄ�=�7���?� _m�� ���3 �:��!(	B p8+���T� $����GH 
�A��u*���+ �M�Jv�S%��H���9�}��js���� i���Py�t*'�kCp��x� ��)��r��Aj��Z��[ ��_����h�.���N�(����\�`�b�}, )h��#6p�: ~�&�fl ��	^�P��x�����]U� ?��w�V%� LG�'�u�0 $]I���L�� 	 *���� q�>���s �G�+�=( �p'%h�n���X@��� �]�˜sCE0�| ��:s� j����A�� WQ�_/2� ��I,k� �PӍ�_� :�Ր)ރ� F*@RfDo ���+�!�' �c�;�Ţ _����,\�9CZx �n�KHX�� h3>��N� <�'xL"K �u�T/��߅ ���N��< +������ �=�k�I� ��<� z��
���� $���%.��[�p+� p���ە",xq�/FN >m�| �&����)�2�A� �O�&#�"9�i������р+jD� 4*5|	��" �L)�(, ϐƣ��b�WYXia��E
��C�����J�����뤮 ���=TgB� NX�܉�):Hz �j��_�� L���D~H,˳I<0~�J u�Q��������	 ���rf�\[�|z�:gQVP	<�R��` U����9 �P���� �@�^�� �w��� �J�z%�@��e�N�4���Y~ ��ڵ��K $��|,2L�j�z���7b +�`i�>���rn,|�� ������� ����AZ�	�n����a�� Fp �ǔB4��I d��
�� �Y�1'ZzX �NhI�/��L�+� �f�B@�� (�'ZY�=��H� �,�X�8 	�YSf�� @t�l<a#�� cR�.��8yMY�o@E%�9��aJp��>yPO�wrP�QszO���	_�>���c* ��4�U. vIQ
m�H� עB('� ��e��+ ^SY.s� lE/�	'y# �K�"����� 7.���t���$# �) m�ʇ���,� c@�' us�+��0� ��҉�t���R���� ߱UV���� �S��"8$;ˣ�-v�JRQ' ��P���1�k *��R�\ l��̫Q� G�0�<P�T ]�Z�� ځ�7�2=�N �yGQ�F� \��3��KCi�����и6 	3�Yq�I�� )=�a�`B ˳�}mU[z/ �V1ݐ����F�j�n��0�8<� �?��`Q� ��Zw!p&�H�J�E 'Q%���Gb����F�J:0����)d�@! h��W��� ��Sڧ�=�<;��m4�`��|� 
+���f=w� D}dWL��h5xGg��v�&��D P�	�Lu�Xӂ>ɀэp{��~�����! ��֓���; 5��$���i�+ ��ݛyҕ� ��2O�% V��~�G~� ,���>c�[ �S�Q�� ��`�^ 5kE�6�v ����� ��tC�=�`Y�eMO�W�� Vtd~K� ����a_n �3���]� �,m0
��� ���rB#^F8S� �č�� Z/��N�&��`w�o_`��� ������2k���=E��%� ��e�4` _�ۃ�Cd�M�R?b��V��� D��>��O�S�;N����� 	����|�� d�q�$wY5 ��b�(�h�� ��x�!Qt� 5H@���ZK���tG�`'�ϵ�х�8Q� (��x]�\�	��� % ��lU�rp0�=r?� ���'���� ~����� �R�F����y2 <�]��Y ��R@����PLj��u�'H9 D	(^�U }%.gi~R�����}@�r� ����,�� *"����B��ݎi����/M �H�#S'+� Xcv��E0z� �]x�� � ��B�uJ�� ��!�I
\�D S6�, �A��ێk�������
: j J�q �wP#��Lx& !H�S�/
����3� N��\	��WD"F���+ ޸sTO�wt b����^2�l?����w���n("{H���G E-���� 3�#� ���:��,�O� �X�	�;�+�QMA(��h��-e�����q�#�l������,^��&�y� T�)|� RkN��[��=$D� ML\U h��/X} c�����D�;2�H� h�C �>)}I�i R��������ö���. ��_�+r�� /����A` ~f��� jL��T�^ �cC�[N� ��z��� �#�P�,�2 -�tO�هF~:N��z�Њ�w/ �p���� @n}t\ �D��>Ek �Z���P �c��h���, X��%��a;P���@f�]	�?���!��  9�Z�ڰ((}��� 0��Cе���%��Z�~�l�? u���D�W�V�b��w��y��A󖣝�|���U �-��@�h� N����> \���jX;v ����� ����" �h�
��ow O�&�'\,T H5ܴ��< ���'�q{ �@�n��Z�3�Dޚ��J 	R<��u[ �5*�#͔ �]ٝiX{+�3C�ذ�� R��e�+�A����̺@����p� �O@��� /ً�[zkZ &�t�;�� �e�������[�b�X�y����Z�>���b�vh �	����^�JLg��-Q� �3�Y�'<\Uz8_�F\P7%�e��"�I��� ��W�
��� 	�<7U�Ī��������@�k/ 屐��$� .��A)Pݥތ(դ
�XΉ.0�<�J��u# �R-	�(@�F�$0�w K�,��M1� 0t"�	���G|wD��t1? 7�߄+��f�@ t��iI�	�X�:���� /L�D"�G�����rA����zJ�,���p� �_�\����� E�<��d �A��H�(i]�W�Y���t� [ܗN�_ə  
&V��8"S ��\	�b d�2~�$ _3G"A�.�F� ��X*�� 5���oR ��y|cK� ����\I� "��D %d�0ڵ�8�Q�X1@�*M�� A����� �P��a	�:(O\�L�k1��� Z��0,� g *_7�^6�������� V�9
�^� �:���I�~ ��T�HXf� �Z�V�a\ ;rE����#�h�X��j N�uZ���(��4�h���tX /�v��� �I7Ë�� �qS��� s��C�� `V8!+�� X�_��Qp -���ߺ �|e
��Q��-��V�OJ� ����!�\��Yפ� ��CL�Hbt���GT���̊ŀ,��8
g  �þR'� @�D�X�G*h;��O�`��C �S()r�8��n�J	^��ľ��=�n�� G��� ٲA�2J '��R�w�SV#�h��� ��ε�♘r �����i���\�@�:��~� �KS��O� a��V>� L���$��Sq� �R)�PΗ �f`Ɂ�[ �$�p�:� �B�ɉ;�w�&�����q}s|bLI3�p)� RPNV -�����^�(pz.�%{�Ϥ��& ^!��F
�* �8���kY7�` �Z	�֌>"w, ���_T��� GB^���a �Asnؚ�[V�� ��m#�@ �|5e~?R�=�.r �&�� '��R�n�08Ѓ ��[��E�gO��qɨ��N�쀀&�\RQ KbY�9+P����4�~ h�5��[� ]Z����� �֤��O:ws ��o��e�Z��DM� ��'я� �1]�Yj����.��7� @3�5�ˡ�� �蓀� N��i�<�.�e�����R|� �'[0fހ^=\��Vh�� ��
Ͻ�CUSpr�7�_�x���H 	h��u� ?�`^��� l����� O�k��� �h�f��/-��9�`����L�. ��^��g�
�l��  !�x�b
����=��Q '��!6��� mP�+��C a|~�9����=`��������ܧ\6�?�� �g�p��w<;�C߿~�P��G��
Џ��_ ���dxah C�����/�L�
�8�����]G���\�)ê@� �F�P��=L�� ��C!�� I�l�0V�-�s<�����yu ��1H�� �κB�އ Rw~ C> s�c��4 P|���F���!�0=S����4hԅd
C���_�D�7@�2�>�R iH�%�X �\@Z��Yv <`�_�?c؟b�ϸ�緀�P�t ��D$���1 �\މ"	�Dd�Ä<м� !t4A�p	�� �"=�D�������>�C��H0�G4=J 	�L"��M<��$N��4OA��6U�3X�W}"w@v\��,�;�dz�y��l:�"�&�+�*P�, ���3�pl6<"8���?��Ds��J�4\9�!�-͘�0A^:�i�P� ������T�*$�<�t�D@���L�Y������`�0 �"�3l�,��|6P��&D�:0����d�?8��\e�aPLg��y�%@0�� �_I� c}	z3(�1@� ~�}�"��(`��� �p��"��KO�@� �<v�:@�(���d#�ɢ�@����8V �"� jL�qu ��<&u0XVL�� �%���:U8�R�2@<�@�ƌ��! $2�H Runti me �r�o�ڃa��0;�@QE���X�567 ^A� #FW �U
�Np��[$��<&!>�*2�p� ��
qK ���Wlp����D�� �'6`(	��&�L� &%.*d��!��G�$	�HБ �D����b���� (�08=/���PX�`�h$p�x���������������������;��S#��d�erj8
C@ <f���Hg 1���#Phiļq�j��G t(k�#�� ,�ߑl�� ��2��u�G^H�NP�� WX ZV�AEIO bcdfg8hj^���tw xzv aeiLo; ё��� "�&L�� �ȦDU Ai��� �����\w �	ԑ� x"<DXt���$�H$X�G*y�{4�|$�ਏ��ɍ��?p/8�� zk>KI�Q8�� 9���lp� �x\;U���6��"�J���	��S��$��{D J�*��M/�
I��(�T���B� ��H�j���(��ELC�`�!�i�\��P&�Z��+$t6��� x�p^�	 $8_k hA`a���b	"���cDp��0d���h��f y$b�	�l �m An1Pi `kqtD:�s���$|�x���`��	
���Q���8�ȩ�����1�|"T$���D\��X���!@��!B`�H���q�������.R�.S ��l2�X�� &T����H,�� B��\�"��?$���P�� C7�苀`���|��68:pn\.�̴ �p.`�hqb�c��> 0G\��,�XF��1A�	�r��&D 9 �4fq(u��hIn��%�蠑  )��>J5 ���0��	�1� �!p�P`����4�s�Q���8)�Ļ���1X�(}�x8 ��$�49� ��b)P`Q��x�!f�Idp�0��"���L����y �5P�lH�,�9 )�`F�x ؔ�c$�*( �Q�d�	��y� ��R��{S$X3� 	x1IHA �0�l�L��dTf��I� -T�dH`2 R�|X%� �x������d1���L��%@�3)< "�f�!lYD�����I���-Ѝ$QZ��
������C�SІ|�  V����ǀ�>D�G���Ȱ���H� ��# ��B�|^��X� �#l�Ht.�ԛ>�f�1�pC�l���8�FV	$bHp@��D	����A���� ?� ,�BT$dHv��;'���M�������zz"��B�R nT3�\�R�S�`�D��.�\�d&�qH�X"hE~ࡠ2.�s$ �ґ�)� �Ƞ�2F$ZHj�z���� ��	��$ �\�"D&�:A��|�������?���� �	4"qD Td�v�$�H����������q	6B$Tq���D�������nUML��	,*���j�\|x~�$�Hr���D��@f��8 $RH^�p"�����NĎD���	� [�&".�6 @�N\$hH%r�^�e9n�Ux�<d� >G�tCur���Tha dI�mDF0 �Crui�c{ a~S�on�LDv��@�� YI�o'$�z5V]@rfu"F� �J(A�$oc<m@]�j *gQL�y� Wicd�ha� ToM1ul�B yҊ4�.Y!�-�stz�n$A�cpy����$z��ibr���Ex�N��)$��[ 9S{��p@�foA��7Pr >�dRs�L 6Mo���Han���Fi�N�mu%ZeMJҔ��r��Ә=8m ꓚ:U5"}WQ�,d��԰LjW $C2s�� ��5�b�WJ ���
Unh��{ �<p�M3�atAS�&Po�� �E\)Of =��?�͂w�D�`�:��R��0�o	� j-Sz(N y���mTi����Bp� z�8)�M�L Iu�r��sK$yb�
�d:i}P��n�g@M��a� �Box�HiN��tg`��p����{�H3� V�4�����n�� �!M��#w ��auRt@�pP������/��f�o���d9(�^�
 ��e��9%�&���'�=-[�X�T��� )ΩG��d�|W �t�@{I�>�bAM@���) V5v<�$um��f���EI ��P�
�� of��g, ��b�ܩ�kqr�4����YS ��,<˲D��o��y4�M] PG�{+� ;�q�&yJ �Eu:�� ��ƆIsB"�WPt�8(�Sb���=�R�L�z ��)�25y �m�B���� �FA(V�is��G,���@ET$��  ��hj��� Jn%^��� �z�������D�׫��� k�paWc \��2&Aqdxz�PX]� ��(��t�f�S �DV ��%6�3 C�i��&�QD�v �>�LJ���Rl�f�b�\>&T �x$v��:YJ��΀1=47Qt"?)�{$,g� =X�D(IB��\p@���SWHowyT�) �P��DlgI5�Y#�%��ip�K��& f�'� �*.kJ+�e0ImL�h��� �?(b�$�΋ �ec)�_ �PC��hHUV�@�ԟZ>6g��X���)*Ֆ�&5 -OP2�М�3�,䚸�>s�\G�d��<�=w�]�*Ț6xH&W� C��lB� T$�[�R\}Vn!��hG,�C� �af��� Y���Qv�zq���Rp��U�I�]n�hu�0f8 ��2Zg~
��
��p�L n0',G8g<��w�H�L'PGTgb�j�r�z�������������������������1
���"�*�2�:�B'JGRgZ�b�j�r�z�����������������2 rtvx&z/|P~X���� 4���5. '�G�a)6] �iф�7 f8���ʞ�ݟ����� 9'%O��BH�V\Gdgv����ǝ�ǰ��������������:'G0g6�>�H�_�:�(�ʤ� �";8ɇѧ ����<r�=�60?�HS�\cGrgy������>�� �a?�, �5�z�����J�� �ID � �(0rBtl vux�z�|�9~�:�;��I�4?�����  1&N8�P� \dI{$� ��F2 
�<`�~����@��3
'G g)�z��Ǒ�'�G�g��������m4 �ɳѿ��� !5r't/vRxjI�8?����� �7�NΎ���8�CA:ȓͣ ݳ��;'� >�S��C� n�������>.�w .���$��� ��]E�
 �0���&A �YO���� �31w��2�9���d�x�z� |�4�*��p�z��|v����觕��?�N���g�D']Gh�p�{�����I@ŧ>ϧ����6��(�-�;�&�� �3�@H<�N�4. �G��5��# 16AX9j�z �-;rKtav�x�= �V]�o� ������ >?C'JEQ�P�X0K?�� 1x��; 23FN����l4�I������� N9r�t�v�x�z�|�:�'5 �<C�IP�WO:h�q�yуه����������J��֒�� ��;� &�.D˓j P�Il���������&�
P t*��^0�s���r�t�v�g�=�������= ��"�*�2�:�8 4�z����~�T�⪼|~�v�}ʰ r��������>
�pvx"z*L2�~���R�Z/boj�r�zς͊|��M��?�N������Oڏ��������
N�:"a*O2���Br'R�Z ��r���N��� �d�@` ,A�0 Z" �1��8I>H�.X�`�h�p�x�������堓��1d��������������1�� ��(���@�H�X�`Nh�p$���r�t�v�x�z�|�~�~�~�~�~�~�~�H�<��2P;�>� �(�0�8�@�H�J�Dh�p�x��im�����`��Ob��Гߣ���#Z���8��b@�D�HNL�P�T X�fi����4 �d�㴇ZUp�sԣ��� 4rtvxz|~�0��M\�?d�h,l�t �xI��V��������`����
�5 ��� ��� �$�(�@�d3l��t�x�|��Äӈ��?��?�?�2��M�� !1�x6 �� �$d0,���4T�;H<h=p>t?x?|��0
�靤��̟�ԟ؟ܟ�����F7z$z(z,0�4�8�<$$D�T�z;|I�`$�b��Jd��̒�I^�$`�b�Id��988$�,�;<4g��@�D�'�\�|��$ٌ��H��~|�~�~�~�M��?�?�?�?�?�?� ��9'4G<g@�D��L�`P�X��Hp�Μʠ������ƴ	�Ɏ�	�:���(�>%��L��X�`�d��l�p���������ɔ���'�G�ğ�v�x;N�� O� �$&A�NDd�PlcR�t�x�|��帹7�dj��{�d�9<: ;$�(=,:>0�4���P1L �O�Ac�Ȉ�v�x�z�|� ��=�5� ��T$?rct �v��p���� 0J91~n4 �5����� ��6�
� ����"�&'*G.`2��7 �$O�,:��GBe�2��� ��<�'�@	>� �����, r`��*1��2"᪚̘� r�t�v�x�z�|�~ٓݣ�������������� 4�L�5c �����Y^ �7�LWBw��˱8(�9�Qف����r>9*���R;h<�= �'l@�C����������=t��� ��$9>).7 r��~?V' �G�g��ť �"���\,':������1�,�̽���
 ����JP�t ��4��5 /�_�d ~���6 �?�[�z�� |�~�H�<M�P�p��z�%z8�iv��̟�Ғ�Ȳ:`�,� V�g�%; 3��Y��� <d䞜�� J+j@�QdO|���O����>, �;�OP$��Y?����� q0�'� G�g�?1k t����ڒ v]!�;:<B=Q.[�;f'kDq�.|����Й��'�G�g��է������3 	��$-�6�]e�n�w c���KhHa� ϯ�B5 \�
��M%� �G�U�p�	y�f������hJ i9'NF �^�g{K�A���'�G�c!��N� ^�f�{,�$ ��?n;�Ns�`���I�b�A�0',�L�&�^~@�D�HM��9?T X�\$`>�h�lK�t��h<=����ϼ���.��0��������"��� ~,�9:;<&�
>?r(t04LK-@��e琄�`�Y��.�������������$��;�(��ĤC�5�A� ��N>' Gg� ����0�8'<IBsQq\�`�h��t�x��Ռ�������܀�Z� ��M?y��`�����ӛ��Y�O�7` ��������`�c �B5&�� p�O7�' �G�g͠|�2�)8'+�5�.���M_�?s�}���������Î���%�(� G3gW�c� ��p�K|;��Xv�<�=,$&� >�˅�M���0^1p��Z���I j��\�P>% p� #��� 5U'�J���7[.^8>�G�-�0ֲ�J�L� (q:r�;  іٱ��� ��4$�g�;�����C��t� v�x�z�>!N.�� ��܅��0S����~� ���,���2%������Ѽ<�t�|��4K��<<v�5��F�0�@u�w7 �^��Q� <�=���' ؐ��K�^�k�w$����'����N̎���A��)Ͱ��� ���� ����  �$�(��:�	�t�|�������	�ɠA��)�~~���鑊��%�c��=�	�lQ W�� /1K�b���2}�-�g���P����蓼 ���^ب��S< 
=�>�.�� ���V���;��� 6J��N�	 �/���bqP x�K�� ahOt���s���X������� ������ ��X��;�ʜ�Ht�T��\�Џ�� �ɰaּ,ظ�?� ��?`,���YȀ!��2 ���X��  %�4��\hc�,�e��؀����i Ik&�TF0 D\���$LLRZ�ʃ0�Ӓ�H���\~�ɲ���� �<�NZ��� c�*�Vx� z�^�" �� ~���<bS,&G@�ȸ���i��$ځ�~�Ϫ�93�-��`���x���Б$ ���_96�XuB ~:�-�8'(�4i��n�� ���%:�l6�j����xβOI2���\�$�/� �?]�~��� ��t&��N�a�s���ߗp�?M�;6<=H>L�P�tmO0"x2���kz��R �Tv6s�u�w �y��jr�tX�C 8�4�a�eT-X���,9z ~J��� ���!�% �f�z�6e =��
/>�� �8�:�?.7��,��2�` ��!0oɿ ��������t��91�&F;��=���2bB _3cp�v��4�<R;��=� [w�I���� �����$.� ��t:x'|G�d*�$Ձ@6��L�|�஺� q>u�h9) �p"�- 01�5] ����o2r st�W3��X�� ��ϟ� וۈ�4P 5���x.rf?Oj $7�&� 3�?�L�^� k�w��~��9 ϝ����� ��pk@�R��x�DRJ� T�$� ��X��Z?�,�~Y$�4�b0-4��8( ��Dt������+7���? |&�<���� ���J��:;��v>�\��崋�� �jNq���5 X"M�L9�: �%A��hl��$0X�A�/	p� ��� `0�B[2� P�J˃��h��:�B�I$>Z��C�6�=�Mˀ���� 7-�U��X�� 98O:l;� '��|����#9/Z�N@m�7:� .,���s;��X��7>N	xb� t{낰��� I��J�G�e}��8�� �%$a ,+4×2��� ��6(9�!:1��;T���Az�<`& '�3K�R��u�}@�䛰� ���ʗIpMкL��K��^�d��s��`���D�2�������l��I���� 1���t~L2h:��B$&���Ct�� ���� 4<���%�� �ڨ�L�:�;�<�&Rd�48���t�L4� ԥz��d� �q��2��� h$Z�P:��1�C]2�!�`��@�3�y�;�	 5EN����&�6r� )7��t�( 8c�uȇ9$J�/����x{@H���Ih�� ̬������� ��"�O�� ߋ�� %l ��5|��� �I�dt� v�3'�H(�\� a̾����i<�A<v �P�#6Z�_� -���N��7l���/�r��tӕ�8��?��a �>	��Kgf����V2 �&�֟� �
�"#�0� μI��!�1��� ��),�:p �zK|S^�	9�'nL����2� �>������� PN�3�? �FLO^�n �tq.��>	�,X� �R8o� ,���'9���:;�j ��"p�u� ��O��	>]a�� �=r)M80<b �5>SN W�[�_cI g�|o(�&w�������������Ű�������Nn0�8A(L�i�o�~ �?�/ӄ������� ���T �����C0� �.�h ��1A' FE��,-9 &����3AX4� +T�@J�Ѓ	7�I� ��!�%�?)d5��:];q���~���[� p����8 �
��I�|4?"�&��B�nӂ����-�N��z0 Ռ���Õ�������`r6JG	iA��x>�t%^/�6z+��\�� *?��� � ��07�� ���C�G|b O�S�,[�r_tg {�t��� 0���� ��3��G�WL�Q �7r�'8 YN2|ɆP��T�����+ ������0O ��i2'�+�/(�\�P;��CyOK�Sp�~e�nJ w	��A��( �%���������	;A�&(�g jD�N�b� ~���<�-��v� �ªy� (�,�z8�.|An ��-l:u� �B��Y>�?����iN������2�ʭ�7��P�t�v�Z��F"5C96 �\;n%�a��"7�p� �9��R� ;NL���� �`"t����^ ��r��x��� ���E I�lpB~�Ys� Lh?�'��$�
�=<�I��_ �m>��φ��X~@ݐ^  �0���:��>J?R-Z��D���1 :�\�d �*����z ��3r!N� F�P�tO v[Zo�ĕ� �Ը�I�2��v�N���� ���6���Rg��Χ�� 7/�yѕٴ |�'�z����XL eKv ,:b�|�� �Ϡ"����t �J����� ��\=i������>4��[�rz �Kiʯ�`9�� P�@
&r0 L�ҏv1�2 $4�j<O- T������|� }3����� ����^@� �4/���>Tؒ|i �Zs
�}ڟ������J��T,� *�-�\<x���� �R3/�u� �98) �Z�~��Ԣ���� zஎ� �즺�K˂~` x[��D�\tP �����ᝁ 0
<)�Ex>�Q:=W�c?o*v�K�����D�z "8��?|�:X*j���Z��� �Ԋ
��D�� _{���� h�H"  0$KlyPZz �Nƈ�7�C �Q�c�h� �����,�NIi���$t���.�V�Q�  "�𜷇>��4:Ԭ Z$������ ����%X:RV~6#N�<����t�L�
��b�{`$� Cq9��_��:t������O��pr�1vw��� V�>�F�������� K��R�]� l֜G��I��' �������?3�M���b��t\�������G���0a���� \���$( 	Ð��'PhI4�J.�� �f�n��� ���Z���� 1:N���@� O�
$�a i�|X&������(��rG ���@8f �9�%����vV����'H.�~� �֭�:` *�����( �VUE��F/�������%�K�Ȭ����̔�s�b1r��i[���) 5-���x9 N=�EA�M�Q.@�Y�J~a�5iT��%: $��!�P��` p��f;g <s�t�� ��,$�>2����^l���А�( ��1*�7Y䦀���^�	 �xT-���DE��aÞŸ�������';l���n��pK���v �ܮ�3�� |�4�NΉҧfڥ���9 5�:�06w%I~�T����0�=-�� x":]/�C ����\��. }E���T�e �z?['u�����`��I�@��ì���N� c�q�y�0_ �	�'��� 4~&6 K����_��ϲcx�t�[	H-�� �K��������wp��������h\d��� 2)�D�Y���҈�~��H:��<_�g��� �K����� t���$ "�Z7���v JU����5#�dB������ �Ѡj��� �6�a �k9��JIj\� ',�䖠 t��ˉ< ;X�$r8���W�@z�N��F$9U�F� �@�����-�<��: !K-XFx@[ J�2`�k�r p8^���PN� ���]��?���-��,^ɨ �/�8C�M�]����|�Ӣ�ԁo��0�� \���$��pJ�x��"P�Ю]�R(�+��Ngy�����`RH~�9� :�nz��9� ՟��i��t"��^�k �\��!�0 �ɹ�2rI6p<�=z-�AJ���$�ʻ�LH�8/�34A���% �ה�rLX ;C<o.H��� �d9n��� ࢡ���x�!c;�:���8��<����J_T��d�Rv�N �2�=p�i� �"~�����v ���0&��{�(��E�pd� 92�%��8� {	,�X�� 4���:5H� �^f�҂ӊ������[|�V���������{�.� ��4�I��(82�H'�t(1�� f�k�y� �_�Ȓ��������`��x5Iʼ��$�݀&��Rt-v7N��Go�}����ȫ8�~��[��'< 2�vIxZzsen���^� ���p&'1`@G�\� x��|���� l�?�/��N%4��<U,e�����LE�s��l���� ���~�^� е�d2m� t����3�.��8�U�r�LG�� %7�aD�ٳ ��:N�� (h&*�I� �-��t�� '�������H��m�t RܑU�=>�� ?�,J�z������	4 l6��T8�, �'�~(�� ��C�bQ�ra w���j��� �~�Y�' ��tlb;2 7D��L�P� )����{Oh�π��$F���'���I{"e@��B�L|� ��P�IOؒ�C��O����� ��s�w,� ߥ�D@����|�X��`�8pn1���Jt��|��W �����}�L�� ܨ�%��� ���+��� �X�r]-L�,� �nlO|����t 6G��� � �]�"%�a���U}�Zh�� �^�	��T����Ę�����ԥQ��ڀ�䈶6������ �����X�O �,	5T�rU�A(�?4�8%<<P ]D'LAVT�X�\*��?�.� 俒�  �%���� �	��T�\~�^�$��I ��� <�(?D/H��P1sv,��`%d�J	l���$��x? ���������%�}(q�~��hp97 :;'�F �� *�> �H�Z[P,X�\O`����~��{txe<ŠӀ��p�]�?����Ā�XhJвj�����8���K�d� ��H$�(���?s�p�d �hv�8R�p��_��`�@b�D���V�.�[MûD)��+�q���0�}�0/.�>g�f�'P���1��������S�-�fyy�(�DW(}��ڍI@Vjh��u�oF��6Lh�&uQ:E*��S�t7?�Ȩ����V#vQ�6��W��Q,w��
� @!c� � <�R�	��:!0�
�V (�, p&����� U*��t 
A��Y��І �q8�>��GH��Fj�h#�Pǘ��U��V�(�� 4QS�� ��p-�uL(0����>���7���׏��bVS���`��?3�� �tx�<w��{p� CI��)� 9���nL� A�[^YX�b H)6��� �����^ ��j��P���} zR��E�,�=�<*�K�� +�tu�x�t( �̸]#��:��t��N�� �u}��f@ �����3 t��  ,�/�����#���@ A����⸻�)p�� b�@`�H�qS} �T��� A1�&uS E� nM��G �h5(����z �j���~:� �(3�ۤ �,Y��@�u8�C�S@�� ��P*��g [uo%�WZ ��LҸ+�1{� �E�I9 6�;�7 �cu$Zӕ��B���{<�|;xt\��� #_+�QD�v0 K�)��� �2���J�AX��$��� ��e�P=�[	�/�au�D I�e�c����QP� �V����%I B}!�'0 r��L<������_j00�FL� ��(,�G��[0 pCk� q�Q.��ϱ@8{�D���� ���M�=e78��<	�^(T� �"�h�s BR#N����\�tG,3� ��<u��.�O� om��_E ����f�| ��:�h�S Z}p"abu ҃�еRv��qD��� �:��`� n*��j�� R��Ɋ��/^x�@��
)L��Bڀw��{� �p̡�� �ZX�Ho0����� ���"X�� c��{OG�e�R)M�������O`wN�8 -��(�
��j!Q~�`��":�� S�-�qd� t�}#��
��Cm��H{ ��ڐ<Aa ��$��:�'?��րLD���f #���Kg�& }�����-� ��?d2I��SH� �Ql�gM�j�u�	��< �vf�>��P8q��)1(�*�:�]�"ڜ��EcY\�H.���� :+��$�>M �v���6� "*�{X^� Q�i���<hz�p�t0?�ku ���х�(>B �F <�#~o; =��{�� -V���A �x�i�" G'u��-y  �Y�W!w7��0� t��9�����p�ҁ`�5��wK�� q�1~�= ��h��b�\ }���ǅ'ӕ|
_"���� �ýu^�8�~�<� 5��k� �	/=6<�e?w� 5#��ݍ�8ᓀa�i	�^�̀����D;dY;u���?���[U�6�˧��c�ʪ�wV�n� ��y�cH�=+�Ř
|� o�c�$Z�� D�2缐�4 �E�\Q]�(
�P3zO vʕ�4 ���H��1�,$��K�O�{U5�`�5p}�� ��F�G�u���s�PJ3W�	��b?����tW+|�0_�렸S>�r�}��(V� ��xV� �+��^�X`�H������1g=}62s�A@�D@��w��W}� �3���t�������]�A&���a��Ny"�kern;v	N��ViGtua�A+ocF�ekPo�=cpExi���sƧEu��LCM�)ag�^�Aw�printf�LO�DER �<��T=he(p>7du���B�y �S%s�c#uld����b�8�ma��8w�k^y?�m6c. ckbr�u�hQ>o�d,�uZC��pd�	�R+gG��gA����1#MoC�l��xF�A'Lo�t�S�=���5���� ��    J_  ^�!��(�G 単T���"ٗ�x�>�K��N��5b�w�v5hr���M�_[�� �MA_`}Á��<�fVR�3?:�پh�Vcn�4ɣ��M��Ո���3�PAJ@�@��z�v��2��%8��$����!�c����
���p�؅���ߤ�%1g�[jŚ#{�0�����F'��NU��jx*�\H��'���ӎI�K�S�J}�J������f3&�!�'�fw�~��U�/�[t�>A�z�
��+��I7�>f�|��M�u˕�I8c�f^ɻ�<��>���	��A���92�6&�LC;6�X���|�/Zi��xP Eq�����Qn>���L�r�ba������ {ߞ�a���t����ae�wO'*#~��c��-W����$��b�?-������	�n!Y�jLYZ�7���'.�=��0
�v/�$8��U;��s'���H�>�LNg����m�-�Ӓ�'k��*��?*�LS�~ڞ�Zu� ����M�M��� �7H�;nnG���7Hd��l���nep0O�o�b$�|�mI*G��_N4��e��y�ۉhcA��Vw�O6����$3�h�+M���2�<�,�����uZb=0E�q�P��;��3{�v$��C�������Y�N���PbT��77فC(U�=}�Y��ԪI��V-q�*�<�
���R�������kGԅ�'@�7����jT�E�Bn4�c�����8�u"N��C4��M�f���*����[ܐ��1�+v��SH����_�--�*���p������>��P�y���Zm0/;<V����~�lm�>�C�av(�D�Y�+R���i��7���~MV���W�����k��f<,�*��G��%Xy���ͷ�j)��\֒���3�V����{�c?���+��f��m"�Y�DK��!����7�A����գ/�$("�g�ؓϝ
���ͯ�+�S�B�A�x{�!;an���`Zy;4�jxcQp�,�������O p��w��z���œV�r_�伃iJD��R�UE��P�D|5i�����0Ȉ����܊}D���(�������|8<TGԝ$7\�f��qah�|6iYQ�6�;h�@�MvWײg���ji���"p��P�3L�0���i�
ID���	��Mۚe����ޛ{Uk�^:��1�c*	�70z6X��?6<��bѣ��?.XT� ��Z�«��^2�V�v����:ό`�,��!�˪���e���Xj65<1r�c�?ި,�+���
����-���9a.��b���c[�@��K@�@�P�}>��=k�Q��#^P �Kd�o&DH�L%3�M��q�߷����d�6��ߞ�zZR�ِ�鮚M��WB
;�����}��%4���H�(��xW;����,���p��������y�X��AB��ӢH�FZ��+����z�����U=��J�E5|D��[q�rs�T�a�.΄������������*�ÐŃGg>U�u븛��a(
� �
��Ϋ���
h� d��X�oa��;�(<��G�����b��g�ul�9�t�Ǎ�OwW��t^�@Pm���p6���ђ����E��!d�L5���H5�*NU�:�ל!J}S.�>H�%x��0����L#��2q�N�D�o�g� ���J�>���(zi�檪�*�O�	e�9��?W������&:>L���X>e��j��Kɑ#�j�Yc
��7(�NB(�bc�{��kC�h{�iN��|�����/d��Z��vsU��Լ�f���J��-��dGfo��0�\QP��d5�C��f,�XȂlM����4ŷ��H:���C�f�@j�_*�dSt�튒�A�
�݃��ҿ��s��@9짞�7�R�o���vsL�4��z� %M�)��龽p�=��X�,�~_�C�N�&�����B�eymC\��!3ఋ�/# �s\��9���琅1	���}h��.F/$�z�\��Ѭ{�,}�nɗ�p
���3�fEh8U8r��300/��%b{�@!�F3͒�um���P�o��V_�Ka˷�ܯR�O_��ma��3�u)�ʃ�^�\>��  m�k�>W�K�%���8KC�(��&]&F�P�yQ��P�(��?���hkMS�G��ᗕ�c����:���AM���c��p�IB�G�*��,��vW�2~���C���(:�2[>�M�n.�w�5"7	��Q�R��P�敶������^����5��)[T��5���cM�EUΆ���K�؏���l9_�>����r��Cg�j5��!jֻ�v�嘈��#�6Z6s���.���O\��]A�;���yl��!fԲ����E�,seS:/�_��K�o��
p�������s�s��ݖG&�,�s�����fL�r��m#N�qyUS���fQgpc��L^?���A���Nz�K\o��733$h�ѥ��r�ܡ%���	�o��&h]D���{z��aO�&@��h<.X� {{^o1� � �(zcT^�Eqo��;�@��+azq�0�U����l,�#G}8�S����Ә�����B�Z��˾v(�֣'�G�e� B�3z`��l��CC�k6�ރ��ĝ��<L�-��u�i��������VV�Y66hJ	M���}��R�,�)�JTd_�釴'y�KH�x-��+@qB�j)<�]�јڊ�!S�=�z��r���'`�(����j��L�w�T��W��e�*����ЎV�(�� �f?��dNl����[�l,����G˘	['��tKɿ�%<10���xI�F<*�8Zd���_��8�	�5_a�����ϸ[�\�j�@!ٸ5��q��%��k�zr�=�C�1V��|@���/F|6���&U�x܈���kx9�1�;��X��֙�"�SZȻ�x銂�<m�&������(�N�{��ݾv�-9�N�)�'���;���b�S����4&�dRB|���?s�) 6��t��j	{���f2��*�OB���;�L�'^`��g�|�+
�q��Q	���ƕ�P��҂`�`B"*�=I\��$F'`��[p����ӂlI��'au�[��I&��Qn��{i����vj�`Ï������Ɋ��:�y&@8�K�؁��s����!�Ԃ��%Y��5����](U��=������&��7X���h����#�WJ8.j�9�����c�B���ή���ēV Д��A���wO�K���ן�,ք��'�wFqK��}�T��mT����$���M4%�N3b݅��$�~X��t!��~�G��D܅!��}ُ
n��'Lџ�}�|�@��g�I��~��lW��)9t��&�S�[��b��?�ð��at&������o�㭒pۜ|��fY�*����"t�}�aU�+�w.N��-�	ݩ���>\t�h�Ý/)����:�>"6_�q������1W4N���R�+=��}=�c�y̞N�?��м�p�B&F4*"�vC�n�p��3��e̳�|��ܞ��p�̲��Iu���] �Ş̗X>F��~*�r��Lf�՜F3N2mh����wB����f�11��ȶ7���9���1�3^�Z���A&u���B�W�#}��ޜ}��<S���h5g���MKh�F�>1���_�y&�yC����3G�E���Zw?��M~���i9nܥ������|΄�r\64�@�`����E�����;�S�µ��y�&�#۱b-	KAtrک���]w��׆�����um;��AG(����aҹ��0n�*�I>d�Q�+wPz�SU���ϣd�!<�A�2�6��:��䶥�l���7�
O�0�Z�!�A��4_�fݤ�o���`m,e�vQy�.��v�po]�j�Ut�.��ؠb�5�s�vi؎���e����t(��p[������3 �ay�]������Y����pz���cQ�g:��	1^#D<6�Ng�G��O\�#Y�lmQ�pk~�)��[uBt���ݬR*0͕O('#�P9�ޝ������__��7�H[�u�OΟ����s\��"1���'�q8[���b���>#���.6���l�ᘐ^��R��kg�?v��aͲ�w�����I@���V<_�d�j��˳ `����'^ ��`�-6�AY��f�}^/+�ЈIl����?1�Vg{���w�HV٘�eL���&����d��K)ƟFQ�1&�VR��V���C�m�눽0'4;�w�0���e�uk������-�^d���J���q�XMK��0F��Pt0��ReT�%�)��('������;S�c�lݗ����`�%�
P�]l_"�bv���;��}Z�fS蛏�a��۾g۬J��ۀVtɧ�h;,"�v	�����W�3��E�D{��M�nsW�wEl���ʮ�Ƣ҃u��9Xp�}�Od��AP^���5����i�ma�P��ub�6Q�����t+�Q זּ��"��"SPN�)���j-.��	������f�+���^S��7;��]���uyH�	�X�/�Uh��P�I	�{�'zw����Ŵ3�8�\0�j��gu�|�ɸ�`�;rd�.MO1����R�9u��x=�l�$*�[g�[�Q"�hU[`|��?��r��s�\�~.���1�}�[Ck�z���ZdM���4;�`�*��4waT͕D���-=�g&}A�h/�%e�V:�Ġ�D����$��um���!�[��K
�Y�a~�{�YP^���V����z+fx�v�����t�XsȈ�[����/Y�d��Z'����Q�gE����m!l�j��QOG��(,c=��O��lM��%���K1�X�d�(��Ǧip?�ElN�n�^j�w˛s���dw�����3�P�M��ۧT�� ~\�M��h��@�1�<߹���a�֏�`;�oU�<��!�2�Y��/� �B��|�z9���%�������k�Ԫ?����T!����`i-C"9E��T���9���_��!�Z�!<�5����R��p��m��$�(�W�����[R��f��0߄a��[R��긿(Aĭ�ȝ�,|ƛ|���"Q�:��2un����8����Ke��ؠ����>%E/��btx����8�B��4v�rر��z�����	�Ef1�jι{$����o	lw�S��\Sa��䣲�����9�rɏl�"��Y�o���+T�:�wl����<  i�z�4��V<lW!�Z�RqS����0w�JV�����!�,�Ha���S�>?�,�"Ӵ��a�ifoV��9���(A[�	�C����q��Vx�E�J��xt�U��aX����m�+��78���p'���pq�����4ڸ��}A�J�����6��������h�TL��~�FE�S�T�;���N7r��:7��},�!)i���A��/C����k�2���lױ����XQͣ7���%��#Ɇ��T��p.��ݺ�Y�F��(*q�F/_�A�a�!���_�r$��G4�S'f�/���đ~�Ww��+��1`�ap��b�N���᣷�׏���E9p���ӟQ<�iJ�
Af�WYe�wd��"�������x��}�9�R4qOR�F��Q��b�*����;����A�����?'\"���̸�����;�8?��G�2L���庲�#dG[G&�yE�I�rJ���>Qw��� ��T1�`�a\��z�>D�JxZw���yՋ$1���AUlWl-K�ga-8?�]�p�j۝}��ߩ��8�kh1`U�Ջ�sB�
V";���	�'�>�⥹+Y�I�C��������\��z�2�Mf�m��,�R���A�ٮ��I�Ç+��'�����ڸnW��A�y�e>P��kq8��(��6�t�F#��&�q��)yg����`4/!tzt� Z)"8��}����䈑��㱜[�Iɞk�Z��Y���W��;l���ч
�2-�7P��-8L5^i6Y�S̜��X������)�#?�^ �F��(��D��8b}~�d��	bm6��~���c�o��&�ȾjL���-�:害b�I������:zȥzM7�+ r-����ߑ�u�q�	��cԶ��h�Yvm Lz_���)"�@�k�v�z�`뇍�8�VZ�������`��\F�9��GȌF��g��C��b�D��J������p�y�"Q�Ѧ��%��y�W(�3��״����~��i�᪳[�C�z�iM'���?�h���<��qY�� �9�$fQ��w�B�����h߮�+���'F=���,(3��z��%]�Ջ��Ψ�̷��Ү�y��%��Z  u�+p4��<r�q݆�!�z�� Қ+����
��͛`-�9z8$�� �_�o�q�8,R�Zb�k����З<7�d���!��W���ݥC�v
�_G"���Q�/L�~�+!�d]�;7b*ؼR��㍭�0� w���lh��Ꭰ�c�{�b@r����~��L�<a��N���I�����'���U�o��+-�J�M�Z_��."�C����J�ƕ��|��+10q��gK�Ү�]���`�LDS�'���	�D�K���>��V"���!�ۘ&6u���L��J��2����#:���!����~�4@�{�r�e�{�����eEܲ�],���9z/�*F�ؒ�!K��Z??S���N8}W�x�Ւ�ݢ���Qw��; �{&���\�N_�r��vU�iخ��F���ڜ6�d����k{��?�\֔�W�����)o����BMZ_��z���\�E�z���b)�2�dF�9�;���6(��O�Q��w���^,�\��g���2�P�o̺�N.2���JJ����d#���)g%h������h�5s�]Ŝo�	Y&Fj��<r�'zr������哇������ROWP��O�(�'���EN��E�!_���1�ա�+��Y�4o5��~ۅu�2�`�0Y�``>�B�ZC����ʂ;tl�R�,qd�t0�Isf����Ss@K��7�̢Od�z2Ȃhr���9u���7��e7(gZk�XE�sʫj�m,c�j�ζq�\3]
�x
�RHL	S�T��vN�	oϐ�<|�?�J��^&��R�WM�RHP� `��%�E�_f�
�G���O��>=��7 Gw������}�=�b�,�W��.�I_��ȗ�<��}�8�
�6�Z�|8��#��6��밗�H4��h�հ!���w�6�H{}�Q��Yw���J�T�N�WwzD
lU�~�k���m}��,��|��V/d;�#[���>%i�J$���W��w��Sr��(�����޵z|[�|���q/�J�W���EYÐ���3��x�Y�82x��>HX�U�N-�C>'��4.b�SD�����腛�|���2n{ݡUR^���xu34!G�&2J+��k��H�L[�gEɎn��;������%x(�9*�=[H`(1��ɍ6��m��8�P�)�ꢤ��`��.[PFӾc��d�<�{1 g�A� �bU�>�s����;3HUjPڧ�k������
������]����h1jF�\���B���A }kK;��׃<�����"����X�|~�YԽ �����.��Ri+	c��#��k!"5�?�ܽ�P�V�:�a�Y�2�&�(y.4�Y��z��8?���0�
�#p�~}�}fa���x"�gKY�p�k�B\c���Y7q���o�n)
�_R'+�g�}$C����1�A<3:�t��Y,HA������5����W\�N)؇�zb�N��6�d-ʛb]v� H���[����^�F��tx�0u�;b-,<N�o+De���t.;�J�3�LY���2\	�����P�,½�L~��!�˪6�I�T�Gجl�s}�!*fi6���t�?-ߞ�H/��dj�7���/ j��~��2�꧵�&b�U��l��~��ל�}�bԣȗf��&0dw3L���p�t�E���jz#7ɨ~X�xݳb��&\vR�6Ѭ�{�3h�7mmL�:M�����������G�^" ����Q�}G;�{�c.���8+���؛`�C�ǆ�(,wߠ�=C�ad!�[��� Zp:}�04L��c�S�g�Q���é����d"IIgQk��E�j�8����l#� "�QvΧ~����:s6�e��I��:��hsޛ�
�\E5)�|<Q���^�ߏ��R����bX�1�K�"A���<�E�2����T��h���`���9^8�_�^ �5�L��4��24>f݀����z����A���GF���ʇ�<����2�+F��H}��=T�)H0R.N�T�K��za'<�|C���Ù�'����%�;g=ǝm,������+��;��{��p�,�����Bg'�nO揕jA5��S?7���Y U;X�D����``�_Z{TAA����E(�y�3���a�J������;��2�%4���&O�P�	����Hd�?�|�R�\�6���G2�8���j���� ��-���m�.��e�4T<�5W8����s?�zr�1BtA�7T<˵m\jn�X�)K��팩_�),���N�Ξc�d�ޓ'[��Ơ.h)��&2� �Ci��9it�.��"l8�C�/�%ϔU.�ls�n#����t����֚u�$0RɬF8	��n��B?^�� %9��2��������(� ���mƞ�b;?�C�B��.A-�D�0��A�h������	(��4s�і�ˡ�'u2/����p``�RE"��Pq��3��0��ɶ4��?=�2���%����Qu� ���)j
�Te�!h�6��ٷ	�w�:�f� �׮d$2ۃQ��b�-�q:��&��>��v��3�l���26�f߅E	���w����T���8������>�o1"DB||k�S�,h�[���-��Ψ��m����~}�@:h����@�;��V�����]-*��[�6�ȽP��G����i��j���ўNo�^L�tP�h�ȭ.�������(�+d��5�7�ͻ�F	|]��gpgb�=/c��Q1��Z��� z�߮M���He�kZI�w`(IwyB��/���( Ul�ጠ��1�;���
p�f�E��\u�_���Yake���\ذ����N�5��K�����[��{j��r��l�6<�6o�����#n���TN=�T�ߠ��+>��K�����C� �_Y ��y?QY2K�3���^�zǸץܒ6{��+@���W�(��n�Ҹn�+�i�N��`��F _Fm��wyѠ�~/O-��B=��czk�$q�i�CiЃ��P�K�>�{�{�H�Ej�W��=�Q����5a���1D��G�U�a�)m�ź��X��ʔ���S�!mp9�7����h���������iڏ��w�$��R��h�x� 4uI�ݯ�5Պ�v�%a�$��&�B㓠��Rǹ=Yrr�q=}�I�����.�x"���(ə��h�)���7�Z�.sP��WV�<�3��u򓞍 ����>Қ�S��TQ2
��S���l�m<�_M�Hq��?��w�U��=���J�M�4Rl���.����*cb������8I�W5LZN�!�^)mh�\��}�`�U�*[�$�Ȳ�pi/?�h��%�ڵs�x��6��$��
���mΪgZ*�V����ƞ��d���(,�_r���KZ�4�^[�U41_��7�yM�~E�^�C��8�9��>�ͬր����;���~ V����k �#6����Pi�~�7Tq��Z��Q�_J����
���Ɲld�pK�/X���F��qO�������N���#d^��n:�PcB� �e��9-���S)��W�y�7�|x�`�.oS�R�k�y��1��=��W�O�'��Q��*�����.Êә�{�̬��1/�Zܐ-@m�p��N��-||��wa�&, #Ɓ��	}�k|h	�}��؎@quNg�'���<���o��A1�D�Q��:�'[AO4�кJ*)p����h����ܿDa.�(6��a��53�(z��:
t,���n~x��:���Hꡯ?��'k��@=�Wk�#�	Y&�o'-�E�%��%�n�$�i�H��K�#��T1p���[n����Q1��B.��]?�S���	�ukBt�L(x�bde"�:y�
�w�&��V���O�
SHR�^x��1R��ՁÌ���Ҥ�_����Qu��� <�W���MO6�Ζ�YA��LL>\��\��-%j �bb��-_Hh�Z����D�:]x�썂p?�)W#BيLY���ȸNf�q5'� ���}Pޤ7�y���م�JwmN�,�Ü��&U��Q69�=��d�.�T��(ӑ��z����?=�.��[F��r�@��G��|V
��l��9�1��ݷM��޻�6�P]a�������P�;�oʦ&�O���^�k�����4��؉�)�z��V��,�F|��w���?H<�6$<�B-o^�Z@�u7��+Q!3���r�����|�⠟�m)�'�\r�)�۝xH&?$�X={mr�Nb*��I���7G��­u����r�����6���P��og���C�ЩJ���f�}�n��k�P�jz;S�>8�Y�PH"�ǆ8�S�m7��]O������^W�����ߘ��1G0:��j�!x��Pr������KUQ}�i�8p����{ʰ�L&h�/2�ň7�[F[��=_\��yMی�ҰiP����A*��O���yL��s�G�Y��mi�+�/����a4s2%(�<�e0�x�.�e�$~od�j���yyȈz1G�>?"e��|�n!Ss��Y�G���gޞO@=���
��HdK�g�L�?��\<n�%��Od�Fb�j�B��[H/�]}\�_�ӳ��	;[01�3&��ԨS�V��
��.�{��v�xs�P�8�'��}����#|� �L�f�=��A�H�d^�U!>y�#NPa0�3�x�nA^&H"������_�S���W"R�_��3�X?6xY��#���:=xy(��C:&�p;T��(�l�.A呶���%��%G{��w.���X�]p[��{���?3f(O�����W�"o)o���[���a啁ǂ�+gI��8�-k`���1(ݑpI�7�-q���r�d�}��[�%����1���ܢ1/lwUw�&P�7 )�5��3/xt;�s`l!�p��y�zb	�B2���Ź��������<���c��(y��.j���a��\v���DÐ���-�g�,a�W�Iuns��2miq&@�s0���QDf��Auؼ�����'좴v �9�7�p��2�j���ݖC�k�������^���-���j�wRd��-~�r�b�fV*<�e�ҁ%���፴�{���:4�?p�ܜ<�xR"��+_��&Q�M�����uN��H>%�����0DӤ3j�g���M�vV��95ɥL{�Z�E3�p��e�B6��|�Ugn+���(GV"4��ę%ݖV2v �ƹ��>Q�3�_�ZYN��ؕ*η�p	I%gҿЀ�C\�blc&���v�]�2��\�ct�[\6!���m#��� �)#�{�`_ʾ�j;k�|����#HTؗ\�es��	O��m�ʹ�y:�/�� A�t�0WB��a��l��Dp,�ng\"�%,Ћ�����[i�Z9�Nu�:=�U���ң�闙l'��P��q��Ϋ8�WX�ch����"��8�D s�p���B�*�g����Hi])�ԨA�`ޫ)'��سB_B$V��#o9��!�r/�O�J�ޞ���u6���������!eh���B<h����Zh�o�!3�\lX7��\K��=�m�VGN�u0�S"8kٮ������"��uwk�&�L�T��V	�;�u��\����5�1�.�ioM���mR)��gw/ޅK�QC3��B�b*L�('���v�t��`�rҚ��vr�
A4�i� ��â�S�,h��s��G��>y�v���l~i�w���*!��Ubn܍xx4�YW��`��&;E�1�i���ݼ,*�{" �V���M���Ip:Ŵ ihh���N�0`��d�	����-�1k��y������AvZch4�q���;}�.�w(���-��n���"�P�?I@�y�������S~��u��YS`� c���!���>maù�U�eg����%��g�j�����5��=Qh(	��BV	)�����ݘ�2����Eg�ԣ�*M}���M��a@7~��h��0���(�ȟ���3\[f2mvU��fdv.�>1ӗ�hX�aS(��Ma�	:�l@ڣ���F+�}1������	��L�x߆$�b�+w(�xe~��-���qE|Xv,qiǈ��?��	Uy�v����8��<s�����Me��toL!V���U`��������-�\��v�ۯ�q����$�$�܆���`�4k�V>���E9e�HOA���Ǉ<�I�\$�̠&I��6^&���̛2��#K�����E?f��|�����Ԫh͞�.���+�����ٌ#��tL��;hM ���E��$���l�}i!}�;�H�7���=�!�*���@�<�"��T�����Ӊ�ME��!pX������j)�KUV�O-~��Eٚ?g3���{8����PJ{S`�"s;y$t�������{T�ž�ݠK�Ę�l��mB���(��h����3�Nn0�TvWh�F���y��P!���2���E���G���|ٷ���c[�Ӳa�J�,ۯ��D�u�]|�T�#�������u��xPՓ�����ˣS�4�vn�T��gl���jj�NN���~�\o8AC�=t���'���f��.TԒ�
I�IBI�-x+�НjkǮ���.H�7˼'��W�?!�ɰS��X�T�N'����#�6�� �+8_�V xո�K̌���[�ߵ]�e���H�X�;+��˖2�D�C	Ņ���#�����m�^��;K�4�2��ҫ����H�����B�
��9\
 �����$ј��@�b�'E��p�:V'���r�;�nq���?�.W��|��K�4oq�Lڜ�(�W�k��Q�}����.d�U���$��Ə��T=����d��3;��n���\�o6
���B��"��D+k�XΓ�HT�׎��������R���117d�Р��U�}1�)�0�4��o���A4�\��䐯R�J��\��4������������]ά\�Ks��tM� ������i{4�cA�fAж(B�������|�_��(ږg&�E�����Y��3� �(�C
�(�G����t���\��0�3��d�B��r�f��r�86�v�� g���R��&v?���	NR�����l�5�ݥ������VcK�����?����.��P,/p�_1�C�����`U碸�����J�dǪ���c�ƭu���@�%y�nKcU� �ʢ���:7_�Y��ܤ��J�6�-gu]���͝����p4ׁ%P�����	�{ۺ�3��Ȑ�ZA���q���:�$o�2��43��h��㑫j'�sߤӶf>�я��´Ƣ��GZ/^��.$[���l1�Yةs�Yǻ����L�}67[���j{	9������q 5����(o"w`t�������1ϰ���b�:�`��6����K�;)nM�t��M�]@�� *��K�b�0<
�L�X#۩�WR�"2����y@
��^�2�a��k��;.ݱE|�F��M��S;ޯ��p���xt	����b����R1�lھw�\i5
��^>��n�j���5>���괲�dN�m� ��Dpղ��e�F�6��
�Y���&7e�/q��:����֕l��w�y9�x�\�q=ץ@Tp&\<C�����x�̲��{�Z�\sq�%20/7�m���ÆҖb��.7��C��֛Ǖ��%�G ��>:ч�t��F/s�ik���4�ư]�2��&�����8�:C��<�%5�$��e��jwM#9M���dY�7��"/�%���5�Mma�����b`�$>����_��r"�͙���Up)�7t�o�i���I����S,��[濎��ʱB� ��w?DW��������'Z�omA�}�h��ՎΫ}F�������T�ʔ�7���ǐ<��Q6I���)dPo�7P��W�����Ƕ}�p/Ĺ:�\ڄ��y7J���d��8�2�b��j�z���w]��
�&�d�>|���H�J}Y��W>d��Y�6��'��bx�B��S��Ko�$��S[��)W?�������W�H�Nw���=�Uj����u�ح�����0���w�@ͪ'�l8��Di���^P�2 �����:��7�gW���b�̾@Ȥ��D��(��W�	H#��vޠ�S�4]�F��� Gth��pi��ͳ�5�$�p��/'�ב=Rl�y���	C�d#̉�MGQT͋Z�h�a�3cZ�F$��q*{� �(��aQ O4e�Z��N��ִY�M�L6t{A����m��t>:�J?)�8��C>�{nک�؊f(��5�V;����{1��lȱ��e��?�a�̀lrr���N���E��(��� wq�n;�>6#6�]	t�I�@��]�Ӊ�i�5_#5*9[V��zn$u�����5��;_�I���*��Pc��K�=i��5�h�Øl��ٌϫd����1���z��7U89�P����*?-�-�}�Pה�q�i�vʔ_��xym�� ��'�D����(�p%��dv9|�Q�L��PO�a+��:	f�#5��s?�Y���Z+�߳���wt�8�FǪDs��,>������*��v,�[.Ϧ�<��E�8@��E� |�g������>��g�>w�F�
�c��b�E��f��s0���`�	xaS֌A�fCր e���o�S��J����?$+#䫉�x�G���c��V7����"ze�O]��?�UK��S;���Z�uN�p�H�!��e��M"��fز���� j��w!^���v�9�
� )�Gi���Ǟx<D��pi����@D��	��0�=��]�NFB��`��`w�t:���$�{�1F.@�m��H�qc:ַ{��M���K?�F��ab��G!�P{M$V_��uwʔ���,P�� ���8�Ʌ2M�µd����K��J�~����T��F�kl� ���N�F��j�q���#�$��pF~��VvS���4��M�[ހV�q��>�ƭ�Q�'�
���3�^� 	"b���?�LK�\������f��s[}ZU�ջ�o
����{v7#`���sti-�vr���>�������g�-p�; �7�UukM1'�L�b�����	i��4��*>2��m9�'L��wy�g�k�LVum�e�����̶d�Zr��k�X�I����k�~�ys�8�Ɵ������m�!�����]�U}�YR��g�F�z��,�= �+'�������7x���Ai;7����#����,�����Ezd{�⃠j6�U��E^#�֤2:\YwT�_�`B�x��I^fJy.nt#��h�&�31�n�L�� �Nx���؎KZ.a��`f��3.d�I_��E�_ʋ;Y��{��x\E���\`�SSJũ��=>g�ͼ�P��L��R� QM�m����*��({��T����a$y��XWwȫ���ټ(WbdёN��h�?#��?�?A��j�-���k�$�^E�mvN�hD�V��X'&�ԝqPs���
����/[�0����]p!В��r�"rP�� �F��<}5ˊ-Pڷ�}\�Z.��ȇ���	I%��w<P-��ec1�[`�	��ԣ_y� E��~�Q!~!^t�F���,� �|�=���<{�~ݛy]ڙjZ9E�'8ԭ"W����BJ�+�x��� �{������<��)Y���|yFs@āG��!��'m}p�H������{i��z�q���N�_89Ahj��{��V^��A�&s�	B[��aI[�>���Xk�[QL����	>���ob��2ǽTC��3~B���
���7\J 0��ؼ.�$��J2`��ZnƎ;��}�G�6V��]�V�������+�q�_�y4�'��'�t��&�����Hbyq�q��6�3f�S��ϑ�~ФC���YǼ��,���w�?��a%�w^��"\�U�����/(��� O%���^�h"�>!�/7���n�p�ii<fk
$J�Q��C�"$�H���>�aa���%��QrU���QB;�2z�	X0"ǁw\����	�qv0��Y�0�s?y~�r�ߴ� 8K�4*�~���%���2Tʃ��O�	n{C���6��$�hҵK���6]��o���{]Qa^�Rզ[�>�&��`�VTT���H�k�
j`���9��" 3��y��ғn�,"�d]Q��ע"P���n���BK���~!��a�\4<��3�wA�"q<G*�͹/�L&/=zB@O��\��=�*�.�*�9�^
ⰹc0q�k�W�����=�n��m3D)$l �y�{��`�?����\���3[��/�?��8e��x.Βg��Ԏkh�ᢏ��0����zx��qD�0[�=6vpLJ�+��夎s���c�)/1Ҭ*�6�W���,��nɹ<μ��n��B��W��竀=$Qຟ�n��(e�� 陞g� z��-��Y��*�Z�
�� !=�e�u��E�&m��[��s{ǯ;-,y(�2���jt�V�s�d�@��g�����9`�8$���yl��y�>o����\`�l��!!f�SV��e�H���V����z�]#�S��:0ɚ9�l�2��h��4�=�-�r�t%E�]��6-	������ۯ��������aܠ���Yi5�S�b�p�C0V�����8<u�o�z[ 2	L0�|/G��j��ˀ9���-���S�jՎ� %:��.��چ�-����V��G�B�^(� ��fB�hq�/)wٶO���PJ��֚xOg`� mW�U�]���S�{D����e���+�cu#���%�k�J�M�̲U�ՠ��u��d���KW��>�x@Uc7w�Lw>�y#(�]�����ڦ�e�W��|�w�c?;��2:RƑ1�6ɡ�iN��r�=}V� !4����٪5�%Ɂ���Ɍ���ɩ��W6�ۧ)|���A����KF��t���������j�gfe�r^����߃�Uڊ���Ϧ�+%j��]��a�gH)���P�G>��Z�~�	�N㡜z��j-f-6����U g�7����&.�p���[5l����X�jN�Š��M�j����g��4�pd�gFa�l:�����!���^�#Mr[g�U"F�1C�_J�K;�(�[S�Be�8�������>���v�����?���tf��Ge�RG*�.�h	w�����J�&�n�4��ﻰ^����dĩ����ev�F���GD;�L�P hg��[M��TD_K$r=���ϳqB8x}<�v���6�� 9|� �t恓/�X�&�Q�ʅ𓁟�a�[_��ɩ;��z�R_L���LK�I�sI�{���x¾e��0�4��M #����c��@��
J51�n��bK�2��G����7��77K������8��/��Ŗ�����R�޾�-����ğ3f�\	8f��>g�n��'6i�_�KJ_W ��;AWّ�N\���*�)u��6R=�&����P��Ri���N������w:���m����0y?V��	C���Uu�`��z�P�	E�#G���=�Q�;��o��p�}��+�X���E��\�*b���W�D	��ܹ���!� 
�b�5 +�7'[U<,��g_��(�T���tY�w�eY��]x⚔ �<��*O�2�u<���WQ��%z d����*��nX:�]��70~���>A߰m������q�}�.'&l�>p۾o(�vU���fi'7%[-X�E�S�l�8�����%L��%eמ���Ji3O��L�F��%ډ#W�K*�!F��[�]���Iw���j{g�ӯ\�>uhn�����2�=�q!�2_"�G�bڛVU>��)J�ܦ�K�D���l����?^�z�+����9����/������Xێ��?�3J0�ӫ$�U���W��t�B�'��MQ����p�8�d~v�>�,f"���}3P$�e	J�᪁��և���x0��2�ı�4�z¸������q2����� ���j����A�z����׽ί'�#uKQ7��>��I�oh,	���2����_e&>���?V��$�a�%-�yIʠ� ��-2鉽�NI�s�^`��7��e�n�|����{N��%��H������Ʊ<��CU�!�r+�C	���ςP���8�|P�V��=���,G;z�,rJଢ� U��飐|5ի�^�ߺ��Ĉ)��T��(��K���J�������r+��t}av۱��>,y��t�Z�'[U���cAg^Fi+sw�`e>�u�/����Vx�D�}��v������+Wg}[�Fe��e�j���xX��ٖ,�=j��BH(��,J�{��pb���:hE]����;��{~�u�>�������
U��ж�7s�S��G�S�]���QGᒃN r`�r��L�Ws E �ݪ��H��ʶ�ǬN�|�KbͣB@i�Ȇ�\���x��y,	����h	\��L�j��{"�^�"�#4���=���L���;
+���k���yE^6�V}�c���e]e�OBS��lm]f����CDl��3{��;?��@Fa�Y���eV���\�`�l�j��=��ܗ�f;$3UT�uO�}�!'�pA�<�]%�a��%,�|욫�_�-�[��z1X�'�w��&��_*	Qc}�����7~e��&���^,��軋r�9w���]��짞��W)c��K�Dm�G��n��|V�=������q���%��BRy\���C��o��}��=^S��A��˸�h�)Mӗ��i�+�F��,�0�[[��Wr��[��m���|�z�B}J�۸Ŏ�)�㥯��'��	ƏH�$f�pϠ�㱞�H��"_6��A��M��_"�)��AlB��H/���P�jcL4��\4z�n��'��{{�ouD��r��Օ�]7X�KQK�!�����	��DD���,<��u-,wy�B���<G!u˶��>�_�Yj(=�#���������B1C�w��c���p|Ta̮�A�J6�G���g��Gv��6 ��<AL���� 7���jT'��Fr욣�"
����q��#B��Դ�4k�ɠրIx��w�N`�����U~!럺�K4�H6x��(��RD� ��-#w�e�%i�a��&�aŌ^w�1���~�v���,ٷ�p�9�n���haX�	��L_�H�zA���:�WK��T�VTg����rn~���솶n&L'1�v��ӽ*h%t{^z��>Rpì����(Y�
�팙�9����d��
EBټ������b���>���T����&�9ܸ���C_|��1řD��b����S���S��18�s��D�)���]�Ŗ�Bps�6��[�3�uY���O[C���!\%�}&]RG�&�����7ڣ�JW/�,U.��d�$�4Șo���ri�}d�SJg Q=xO�?��7�7�2�gP?{�Ǒ������\�s�6���{J,�amU�e%\t,�Ͷ;�8��T��:���V\��r��g�ŋ�)s�.��)��?o��1��Cd�c�ܪ:����IQ�Oң� ���.F��3y��@|�������Y����@�|�s��x�Mn�W�"H��1�Dz��
EQ��Y�Ol�(t�N���{C�����Q��ݏ�lE��
�������4��"cH�NT��pS��%`?�N�[m���l
�2 ��n��"��b����\V�t�oV������rK�ے���y�@q�X��%EM1�]�p�s�j�q��2V��?Z���U$�@'v'�% r	�ޖ�1�e!p�3@F�RԘ}�OC��7uaP/����x3g�<�����{A,�]}�D�F�ɖ��V�O8�
�B�)��pG�Jk]J��UA^�]Iz�/i�+w��90�\��Yի1�ܿ8����H����-�(|z�ޢ�d���9�9��ѣhh4����fd��{qS���z������HPe���R��d'��o�)*��i?Aͷu�>N�:�7�=�Tv�!�g[�t�����xU��ߊbk�W��ɤ0t�5��b��EJ��{4�qr�w���mY������#�EB~�S��c�
}؎B H�|���O�}/��7��n�bq@/��'�z���c$){ڑcU,v�/jA�Ok��������+��9ձ|@Y��v��$���}J�9�3���"�7��:�4�N�}
DwwO-�>�IMT�}{v��"��bj2���˕ˠ+��#��Q���@W./Q�b���s�\T��C$w�w~Q��l���"����@R#r����`BO�P�7BB9X�c��墸H��F��j7� ��r��U�^�����
��4L���pR��L��C�i?Q�|�.�Kî������݅�:F�\����j�,���df�~}��oa��᾽ѕѡp�g])����k�2�o�4!)+��<�l�s|f��d����^�&���nbM��;>�d�*�� m���ŕ�C=#Q��KJl��|��I�A�k��Iι��2tM���}I=�p�G}7�G8:vIF%ql�v�������cr��Qw�z��Yb��1��k��j���x�]=�֠ݫL0s3�"�j��cp]:��+`��I#��eǭ��d(�.c�F�se��&s�@���W����@Bu;K����\���
���G׺���JĆn�u����j��N��l�g�L]l鯏��I��ϩ��=�EV�m�N]�����5r��t'^]�Fݳl���5��)�}	=��y�����M���k���~��pT����=a������x`�9�DY��-.�tsAM':�?
�;5����L-L��������qb�@˓�`ώ?m�\`������8���;suvp�`����0����Qf��:��D���Ϳ@|��Y:����	�	��
Qwɷ�"P��1q;��u�{��4�[���v8�nµb!�=~=k;�>]y����8BSǬ�?֒��xH�e��)��P�ih�)��{����.ıB�k'H=�-���t��qb=Z�Kh���V
ڭ_�C% �(������6or8��m֟��մ!ly�X����]w��ӎ��j�L��C�w-�� ���	����H�esy$.\�X6r�+�1���$��d@�8�L����
1�(��i2�Z�1T<��G����ҥ.�B��Ϯ.�ά�����H�V�:)�w�?]��>�g ����4��go"��u�=�c�S����չf�X�l[FC���n!��9�e XT{&(��?[a',.���bQ�%��w�(ݐ��^���S0uP��G>���>B�zC.q͟�Q��v������5=�wj+��9W�d���^���@��Bj��1�;�G����������Ab��]iW��q�u����g�]��M0U��lM�����-�;�u���2�+���2:*�Y�t2��Q�X��� �g���D�v���U�x�g`�9�V��`�qr�:&�px��*���>�[e��̤j �m	-q��J8d�}�ԯӠ́d_oƳO�����?/�!�(��hǠ�6� �=���Aҩ�/̀�����#���p�-�4pㆾ]:�S�&3���-�r�B���<-�Caw����/�<��ON#I��3��Ƽъ8T��;�ݙ<�mxqX���6D0�RFH�3��8�OȤ�$���K& �b�X�Pm�ǩ$���~9bp�w��E[Q��c�{=Hy�<#]���k��_q[��y�y�:`WP�@l�LAWy��xGux�(d�=be&O�ƍ��y�I���Q�e�B=���f�o���Q(���{j��ؒF(KV�y-S�e He�������hhy�E�Ff4yΰ��k:�lB��5_��}s�q��5����M�!���� |����);�J�Evׂ���+pJ7	��� Vs�ٝ�����Tk��c�6���!���8)�ќӇ��G��YV�(,-f�A��/69�;�j�*�@=�"·�=�T�Be�����.$���@U��G/�6*}��A\��e�f�
�۰��%�i���2S��7����}���;"�<˫���)�v����^�3/A�(T�lK��%��Sa�q����,5�59���.�O�)B]��­	!��iJ[0t����J���������!؂J%gpN� �
�U]Q蕛M���� 1T=�q��_o��,m /+F�I��c�l���=�S��+��G�������_��'�+>v3��VEʹ��`��vX���mOx��=�:����˶��^`oK�~FU6ݏ�AIIIʳk�O�˶�uG�\%�h\���V��wP�MJ\+^}d�b�$��PF�]*�������)�j����d�+[��Y�}����L-8{���Y��7�Z�!`�InV	�W���D<��n�乑a�ي �ݩ�[����R��z�'�*���h_������� _i���˽���N�놡SN
�r�DL� �4]��|÷V̌9=��)��w[�7�h4|G��]��a����rb8�T���O֜�g�/��N5�l�d]�b\����!�7�0��A]��DS���}�H�����8��{��(!��:��^���\����z#�K?�V�_�B��4!�VܕSзq��o��2��r
��У8߇꺕k��@�z@�IY�0��GUT�h׾��K��&}n��I�|ᡀ��!�p�9�����r\��X����G����<0�x5�Ky1u�o�� �t����y�(��f�4(;un9�Rff�rF�GR!0)�o�Fm��:�͏e�GN&F�x"[��LZ\t����C��:����x*C�yet�, >�g����O�]�E��%�4��E�� mu~��.s3��[�D|�4 mD��M�r�I�d���<(��P@��(f=8Y��J�4�|:�Ѝ|�n��b��yyc��P��!Zi��5����)5l޲��3��V��&B�٨!I�o��`�i������6{�N��,
K��ϊ�v�ȃo�e�9���c-�B��V�f����a�)y@M[rPʣ�m���v3������eb� �ԕ���>�AA�����̿yeL�ko:$�a��Ȱz���y���\~��n�.�\:��\F2�u�J�M�}��Z%�0�6$� 6Ǣ�%#�{K��sN����!gJ65��|�mL��!��_O�d�aΑ�,����]�u[A�Į ]�b�ˢأ�o�D��D	l�YV�A$`_�$������_c^����]\B��h��ֻ����=�?����f��m}Z Ӟ�|�/I��j��L�vT3פ��a�wZ���'3��$O�sj�Ip�A�3�C"%I)fm�t��."
��EZe�J��IssT�%��NK:�FQ��U�G�K�5����5�a��˳���%[�=s��56m��'!�N���7�vN1�����+w�3C_  �AC�                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                        