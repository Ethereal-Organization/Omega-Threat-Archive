MZ�       ��  �       @       �                           �   � �	�!�L�!This program cannot be run in DOS mode.
$       ]e��������������$����Rich��        �4:��p��F�fk��PE  L ��SH        �             �  �       @                      �    �H                               ϶ (                                                           �                                                    .packed                             �.RLPack  �    A�                    �8149og4q P   � �G   �                 �l0u15g4l �        �              �  �=K
�Ս<q�U��*}�[���B�#��+���j~�d��ݢH�T������yb�����]���t¸�-&c�4&"13�<[i ���
�\s�Z�u"������z/��S�<㛈4va�hj�{��+Yhq�/p��Ď���,iY�ԘX�1ز����$����Βp@��gE���^���V��7�D}j�a�X�B/�+��R�D�^�h�ҷ2_3�8t��0�'�$�냨 U4G��--B���n �r���H}�75|�hX�����L����H���P���d�R%u��v�^K	�T���8����n-~km����~����Ӫ�O̩OO�_]��Kj�e�P��[��1�9�;�L�N�*N��&���׽D�L<��qA0���R���"hk��<]�.���<m|ү *�و���@��?
�p�6��zq��0���5�~jB<�IN�\u���N�c�0K�/��8�fR�T
V�r"���M�&��f�=��9�/5y�����nU�bhF~祊�06�����%�J.|��f�����#Ör��$ն�R�v�U��	_�Ey�*N5��u�Oױ�-4�����RǱi�����~���F�����Sn#�������{��vف}�Vky�q�|�!���znL�K)8�r����x���[<5Q�������>��R�خ94�}|!���3�0;&�v� ^��nĢ���W���0�;@�
�s�qv�7��������}Ԝ���)W&�W�Fd$�C�����>f��T���ҡB���oo��/c\��5 �����6��+^�E�
�X�� /���	����*����0�t��1iՑ�׉d�Ѿ�m~ﯸ�����N@*���fAU)7:(j{A�������i�d.�Q�3�i\i�{�Cl��2t�%3�k�À0���^g���4��KC�Z%�_)`�6C�:-Y�١����E�@d�����������[b�&�Q�?��h�K-/��;�]��zߠ���� n8��-*�e.���iA<��<���#�U�^0��mA=mb�v�6 ]ǻ ����'T�C'4�+�=�\��=^h繙�_��n�j)���
��N�Nx������8�M$E���j�G��J0��f����p�y�n&=+�[s�_��j�=\,�|�Q����a��s
V>��-����M���^�19�:���)�Z��� �W��/�)ؗh�x�n��g�.�?��9��n�m���/�Ѷa�S�{�������d3_��ɥ]�䛚����@R�S��4��ˢ���&���(8�C�?z�H�.L��={����
"��Z,e���'"^Qp^=\��0%(�c����4�����ʵ�m���㹯��A��]�3n��E�KY����M�bTI�
Q��2�B��ݶ���vp��yڨ� �8�����}me��|�F�����<�h���M��w����
A]�qi2v�������Q�;��{�7 ꪴ�,[AZ���=�P~�Wk͂��l��5�#-��F�3��
���D����О���Sxs"���;
��脱3��l�rAx4�B���ey���>b/���,ⓘ�/.'a�����JD@�I�5��rm�aX@s�����P��r���ת���!KA9�F�Л�F� �X�G%���1dR�Ѵ�ˆ����H{n�����M��K����ٹ7�W�_��a��Ix�l�|ܐ+�������h�Ib]�|f=�g�+��9\'��(VB�)ib`�s��q��t��D��+jZy��_3��.�a��	�*�i�����b<[) �'�s�/��AV?(�-�n?�e&j97/�&��Wڥl!�������^9�Q���`y���D���	��ko�8Ir�g\{�Ӝ��.���Ik'�Ksm"��#���y����oڧ�P��&)��8��Flz� �t��p3�w��\Non�O��bL{���Ynf��z0�T���\TE �%�	���������l�I�ˁ��]erڋW��$��Y��'��m�z���:V-bCLE8�n��O�i T��"�"R�1b��X�8���q�	��c@����U��	�k9�d����)����pj�b�^!ft �p�Ƙ���֐���Lq�hj��u#].��	�e�c�T��/R֜�-_>��sIu�<n#�@���Z�ӱh����*�o�r=15d�wb7�A����>H�I�m�0��L�Y٨���,
A�(BޚΕ׽���z�\�zB����y�2}+8��Ulg�Ӛ6F��e
�Ȫ;G� �XW�-�H�O{�)�B�1��j��d��"�1�؁�e_�)�0��熯�AЎ�N�L��	�2X�Yl���L{ߥ��g��{ĭH�� Ixű���d�{q[�X����L��6�s%:Glg,p�Hg�n��3"��t̊��"3��	�I��X��u�AH>�@�/Ӕ�k��S��ݺ,܁~��F�D�q @��h:^1��/�@��2��/|=��1��6ay}���c��^��u�a!�^44=����+V��F�aOd��nq���ņ�qj���9_���r��y�TX�B��\'W��� �a� �����D[Y�D�p�YG�77r���$�ApAG�ܕdN��n�Ϡ}������o�4�-��+4hN��0���،�U����t��ya������Ʉ�b;I�Flxc�f��?�\l�w��C�\�\@�$����/�����Xrm�R}�d�G���X�Mxe�@�f���e N��������B�C{�*�@-���ID��.�#V�!�]k�E�4Hew��4��½�O�@o l	���!\}�1�6ډ8��|K�w-���ٴJ�_n���I��*��-n=�ao�8����^��(�	�Xf��%ɶm�W�ɔ	�T��&�X��	~��d���ε�Lk�����!������}=���*i=z���&@am���S���h3fsi�D��ht�	
�g�lF4�b����^�qí���M����7��)jSa=B�<Q��o f�z���U�Ƨz�Z���Q����� �8�WYGmĪ:f�h7s��Ym�ylS��%5woz���8�a�޷(�*|�X��_��5�g���֘d��E/�L���J��'��7��[�$h���*��_ش�W*�J�d���Cf?T�ϒY"K��ޟ&�xi댮K_�&\�_Z�����0kS��\��A8��]�3k�<��!~=4$|��p��e�z�B�	�[߄������aP�Plt3���z�hGT�jS�/ܷ9�k" �Q�9�+`��X��t�2�4����As5�u�-����m��ز���ǘ���Ed�r�<-1�������n�i2�����QrZx�j���ԍ۟$F������1}=^�ҕ-c�]n�rܾ �K8e���^k���9�9*-H�
$�G����v"_'rIx{�6�#�}�$e���yй�0�&W� f��o��+�hU�$�� />yD2D?h���I�:���Cx�#���I�(��c�C.��8Ge'�(�vb=���G������6�xv�}�'ֱr�$��ޘ���g��Fm���By���)9Kt	�y�������lj�f���V��jP�� �J&�M��5_~ �_��q(�Q��Z6B,qy��ȥ05M�(��.髪͸9���
9��G��c�9��M��ȧ���:Zu��&�g����,-3���\KW�>�A�z��x�2"1Nrt��g�'�휒��W�$��}��ݱ��|��d��I-t����8�3q�>�4ZU�
��݉8L���լ��:N���X�����;nt�r����Ҹ�c[(L�g�9B���S�+f���F�5�T�hW��ڍ��yk��M��}5m5&.e;���J�|�
7�F�t�ɏ�ILj^�&�U����Sd�G������Ñ��ͷ��ޜ�j!�n�0A0�L[��amz.s��>�����<��^7B_�T"���� �LUR��v9 ���9��ν�zd�FD�/��N8���Ĉ��|(��]����J��-� ����888j������sʈ�Yzc�Ʉ��i'bbV�'�A'�t4<��$t�&�HxK"���D��%R�l��끓3o%��Ѵ��8�H��/�^��<S�LA7�]#�2��#�\Nj�<�R�s�3�����օ�
�	�sb�),	I6*U�Hu
�6��n*�c�N���1<�ۛ�k�����ǯ��3 3�Lȭ���t��D�+Q:�������<4o�q���Ʃ����,�*�6J
]A�]��9GJM�:#���~�0��m!����Hr���Һ�48/09K��F�>����M?aJGe��Evȥ4ıB�<�g�W��I�����l(�x��t����G1֣�0O<?/�{H_R����^F^�}��E;-�D��x"R�;���A�X��,��T�{����-�J�Biҿ�����]�����w(� {��a;?�F�ګ��'6ɝ��L�mi��{� �P܃���l)#�j�Ԕ.{Z�b����R�c2%�dQp��4��S_3�_��~�Z�� �̺n D��	�Y[ok��d�D�jW�5)Mū��H#���C7��	l���3E�X�G-���N�D�7*����A�d���OC�n������R�d1� $�Í,8���/���Q˼�i˨r�Z�n-L����e��Yc�{p�R����l�I��V��`[�q�9& Gu?G(`��8���쪘��й��e[ ���)���YnJ�Ց5[X���k�B�)H���|���
)b@�e�l	쵭K ��"�?*�ljRҎ�;g�n����D?� ��;�l�j��!��� J��[��/+���ED�;o�M�PX����@����������[��NE^L)J��D����_����a�!�<�c4��!�	<���C{����F�X�A��$B���N�Ϳ%���=(E3I�ϐȦ��$�?���7|6W���T���sEíՑ��m�Q)��0#�_-3�<��
؉��;�aRg���*����l`�8����E�hz	GD%_��>��h(F�ؔ [��U�m~�1�}��l�e���~��f��̟B��":�TĄ��>+^�>�	]���b%�,�����g6Q��1B���JXR��+ s �S��~B���7EHEל� �G%ܔVY�*lxeְ���nս��Ph�\7D�H����1��O�l���>Bl4W���x�G��`DpG�|1���=M�U����9�CmW�~���ց��<d�//���tS���<������*OF����Jp�������>���	|7�?m�+���[���>��۸Ji��u�/����Y$�V�[.�f[�	���3���Uݙ��&�lݴK��a�fW����6���E�PD�.��'[;�Ezݪ{�'�M�#��L��Z'.��c�>���!ʭ�����VoT(��;3���%;����,0��k�@ᐐc�)//\o�r1�ׁ*`S�$(P���2
�?�wB�������؀2SLɓ�����L����|S�X�8�/�i��׃�Ԏb�9�����z�9�����!���U$��JU��Kۜ�x'��U�#�9C|�?^���&�-9�*���W(���J���T*�g��v&�O,��e�3��f����� 'E.��\��ȴ7V�e[��,����!�d�i���lc��`�)P\���V�8����Lt��:���]>�)As�����Fiט��}�Y�+ꤳGc#�:�M��.e{�V�@���K�O���w�X�M�������m%���v�Y�|�\��%'��	nX��[�����l��K��A��Q_�I|�)�
�d:iŎ�+�0GN�J�kK*�KX�=�U�w��W�<��4qc]+\<��4/���~����P��Xc��0	A��h��2N�P�N�J{3���Xn ô5q����ӽ�p�#���x�T�Ԋ�+ �i��Z�]k`"����e^���V-[�y⨄��h&Bd ��Ī7U��soN�6��5�	dwwV�G�4�-�}N���0ޚ#
��L���nHC�w@��'eyY0��z���~�W=�s���,�Ѐ�
�z�Wr~4(�I�yz��+��Q  �`�=�̚N���m�#���'sݗ��=[�ĺSϱ��P����>9J�C�Œ�s��h��k+��d]We�<q�g�AݦQ�ҟW���Ѻ���W P.us���Mi�O��(׳=U:PG�NW��9FOx�yw���0A=��d�w"�������i���V�H�z��_� �
�f���S�
���?�p�bA�<r3V��]��x�+��f�d}���a'|'aّ�R)}�F� Z©�9�=��:L�ZO˽�$�}��)�)����Ԅ��`�}�{ۊ	��0Z�ǒ��^��*�!���
�^��Aop���rʄ�90�Þ����PT]j���6ByjA�L��;4O�ImдE���M�TN�"FL�c��f���`u'�E�?��VX�I���J�G�)Hrk�MG�5?���	yW��6n^s>���$8�s��[�P���jP�9�r!�&Wn�p�z{I� �I����ߞ����ԀBZ� ��%h������f��"�+� N�8ԻեB�;��E�?M�P(��������%�.���3�ՙ����`�g�GWH���+��ra�&���X����̹�	F�:�I��{�.`�kp}Sq�/�6��O%uU �����)�~�'�mP�� Q��{�H�
�L�0�M1�h>�0Vuq�do���j���������fB��z$)��CR��S�L���g�%7:c�2��'�������^����<��Ê�ت�9}��v"����JBVO:��g7�H�
�+p�����5�լ1�;��vZ�X#�G���[��k��ӂ���L2���ld�pATH띯������u�=�x�C[����#��d���d�>�����0���prn¯i���J7g��i@f�~1�
���
���ﰅ鍼<>Gɇ�\�0G���o�FZ�j��V��#9�����י��H4�U�]~T�J���c[�y\>J3�H�8S��͍~/V�:�q(�@���?���	m5��S�����Y0_�(y��{�-b��C3R p[����xZ��@Tb�O�a�Y�6(�*)��{n�a�{��d _�[ZAG�vTo!Z"���Z�M�vU�K����Ba�Q�&Ө�):χ����_:��"z��r���Мޗ婒���l�"kͱ��=�h�z��D�*�z����3��Y��C.�w+����6)M�:�
�*�H�
�N(��հ���ҚχwݮT�<�g&*o�r�ݵ��|E�ຳ�s���f�2���tx����j۱r��:�R��J��&�.�j/�v��b�C�O��'p�?�-"o�e� ��<^4W�p��,�o��3:����(&m�7JW��Y֜�p|Cx�9%���4��S��^+e��o��h�+7b�Z͡f�͆E����x��l6w�7K�T&L��4.n���amB���K�(I`�@�m���jr!��IW&�+
���?��K�<��:����O�r��٬�Eo�^�.k�A<���ľJ�3�������(�K���kX�T�~޿��8
0����a�H��],@�4����&f2�-<)�Zmbb��1k�J�q�����W�2GC��~�<
���|�/�b�r1(�L�0�$]�*{�W�+x�Td~r9��O��;�-XF��o5ϑ�G�����yYx��W�I%�u���rX(��+1\Y�j>z>6
��B%:b"Av]%��RT�����,�x+����{���2��(��)*��SV��~�+��R�Ȃ������8�	����q+�r�xٜv��K�ᇜ:��<���F�����D�=lC�h")쁒P��c��K&���"�߽Rv4����'��̐�����x��� �o���a`��l��/���?��e��(Ē��b!��]��Q9ͩӄ�=�JH�p�Ƒ��d#(�sI%d�i��'.5�Em7^���� Bw�������5Y<�-_S"�Y�"��0!���a���),a�Θ���#`�P������t��"��/q� ��b���+�������cQ���k~�bQ���ZW~����	fAP�K��![�����_�SIT�L��&&�~ZE4S��[6��d���W�_��y�����6lb��q�L���t	��G�׎�s�{&��6G��n��돈�+'l.�ny�]�e �B�Ϋ�@���,v����'��Z7���������ˉ��n��ʏ���'�[<������z�+֊� gO#���x?P�(Ks ��K�-|���nt�8���r7��3�l�<^*��D�CP s����]D%�`�����O��sT�k�Zh�����u�u�M{��UN^O/z�(��!_g����-���ỳ�*-���>��HJQ�x���+�PqQvK��U3 �/th���=�=`?����^9}O�`�@�Z���"@I3�������io�>M�pnݭCT�<�൅|����]�=(�$!����m����>��u@�Eߜ�����&��L��eoW����R��n����|!_���z~���˼<�2d�u���a臑�n�����)ct���66�[ɜ�g˘��RYY_Óh0��<Z��%��UP����:���*h\�N7��bǢ�g�l]�����g���Ч�w�A��=T4M�\��7�"{wD&�%��.�������!ۇS䙈𽝂�s?��?[�,��Bq�d娟�D>�2Sv�����`�VG��+����צ-��;B����q���w�@
+O�צ�S+tw O�߉F�Z`{�	���X9���T��D�xХp*��WS/���K�8ʄU���Z"�٨�D}�>sqY��/���!;���\��Յ�����:�Nq����6��㦿ܹe��<�}ֱ�h�@���r+�� 9<��Ig����ۜGu��z�%�U�;���*_L�%A^y���W%3�����1�Gh/B�g*��g����;������>���]����nmsz�&;�G��t1vs�С�J��w�ηW;��� ���˅�]�}w���k�\���4�X�_X��s�=��H�����e/�����e�/3 7�����αrL��F�/N>�8��Y*T�����k�A�r�i�i��K�>Yg�e]���pG�8�2�1}�6��9Q�8ﺈ|�&SnK����������E����"�.���&#T~/��d�ێ�Fv�V㲤�#�w�i�u���{�R�Sn��$����'Cy�t�S[Z�X/�9�W����V�Q�{�߿���e���|v�6�	���<�ʟ�����]�ż�x��4Pd��xڸӁp�[^�\�g�:�
���]\����t�	75`���πӰd?|
k��ۚ�f��2a�����i�ځ28�ō����f\��ʮP߰׶���r9&��Κ`�JdET����r({X�ؒǒF���؀�����J�Gx-t�en�+�Z�����]���M�/�4�'4��On���_~Ъ֛M�O��8�u�eޙ��q�M�'1Z�J���?�L��GuoIÔU�>�p3ṙL�0_l`����u�R?�%�B�p�*�s�h*�s�4��nL��g��n���~��7nf2�
�PG��_�{E���N}<ռlH�=Q��p����A����]��"�5BK+L^�Gw�JN8���X�=)���� !)�w�%x$� ��1�G�5-����S�����=��]?ȋ���H�{�I�4��v�DI=n��������P
 K�}���� Nam�,4�L�f�{,T�6�.3i���p�#�b��V���j��#tG���1�g�'6h��Ĥ�w��l�������9P-�5�/��������;!͇�p���9JV�Y&qG/�dQT\�3�P�Z�R����")�Cl��1�*���/�}�Eq��� �oW�@�H	��U���pw;+�w_����F��}Qc���!�{ջϔA�|9����ʶС�<�l1׉n���q�[!�C���3��[P��_W��Oϔ+:Ji(�������&*�����	\�1+t�X�jI��D�{]��{©x;�׉Κ�10���g�c��Al�v[68�\�[�����	E�%�ŵ59_�ʔG���D˨r���i-s�D�,���i2��4h\꛸��
!�@���|��ţK����Q2�S{�`2�|��7p�:�+:������M]��y"{*Q���ܜ��~G��*�"t��$�Ũ�M @c�̉d���o�;��~F��::��4 ��.��"Հ�蟘i\WED�ׂU����3{�<��%��h6�l��Y�������c@�����[��	�U���`I�V��AO�>�W��*��(�t�֐���u���������������P��7Q���9���A�zj�<3/��Z3�o2���#K�J����&�����#�Ix����r��Ub�����<�.A=^�$r�1����wL��5s\�G�S"����e��X���1�g'�U��j+�	\tn�F�@�Hs~�����io��RlR.�L/���nQD>�e�e��H��WT"i��4V��d�U'���֦t��V:w�6}P���"�/�U+����J�#�F�aq!2�{��8G�����J����މDsD/Ƶ=�N�E���a��n5�����j��z6��8x5ܑ?0�Z+��j2B1o�V�o]r%n:����	{m'����1����cݘ����M �Tm�4��q�i��V�fK}@��]o�ؕ55�-XC`�w�
f�Н�f+���p=�p��A�!�e��uq��*Ǖ���n�~~��h��Q��O�l���1hy�Ƌ��H~t���<;��X+n����H1r�m�����!���f��|si��l�G4v:�9SE��i'/��q�c*�VH�I�T�.��R�!��<�y`ｆ�7s_��?�"��ߑ�Һ,��z%�uZ��᧕A��X� L�ԍB����=����#�(��M��/@��b�Zǝܾ��A���C�'���B�P� �� T݂��� �m�CY�������#���Q���,2���}V�ρ"C"9/Ѫ���j����1h�p{�53@o����	,���,���8ř��@���v���XQ	�Ps5#/�M���2N^�'��^#mAtw�Snz�X[h��-����4��X �3:C�A���dup�>�Ɠr�uPf�I#����Y�v��iD���fa�{J*pǨk�[��pyLII�3X�w\��X)&���/B�����E*MV��;k�S���u�ݯ%ϙ^NY:W� �ԗb�/�>�q���'�ƛ�։��1�6�^��8G�]�lĉ�>v�=�$9�[�>!��� +�8�!��������$��`ƿ�ήM��\W���#���>|��C��^��3oz����f%�Σ�` ]�\��)���mr&��t܂d�tt���q��d6��|��:��.^r�A����mN��l/m2�5רW:+�`��%�ª�"�����~=z߷����Tl��c�-J p:�^���6�G�����p�X�S�������m՗��;"P�����x���Y�%G	#�"����H��݋u��^D�� o�G��2M�h}P|i���f��V��}nM+��@|ڰɋ+�v��W��R�ߒ�x�5|x�2�AG	��P�l�D]7:�A�/�y��6����a��R��	n	�-�Hq�*���-�⽐4�}I����ƚ%���oB�M�?��Ւ����bG�usU��R{&�#�)ܵ7�{P��W��R�	>�c��$D�r	��g��8d&J��lY�㦇�%Si Q�v�t7�h��*�N�.���"�1�%��)���4�����=��6��F5��)����Ǎ�+�L0sx�c�tt�r�ל�%j�;_�>e�_] �|�H�j) t��,�EGn&Z�� `r���"i:g�(�`�vmOޤ��}��tPi�d���p��`�Oj����P� �������"���j/=������W j&�y/��V��<P��#P,�/�P�b�p�\���������)�w���r"�d��8#�әp���9�#Hԯm[�\�2uin]	����g�h���~Xd�����Xh��9�a��(0<HC]ٚ!�95��(��nN̿k�~se��D�h��)|6��V�&MAO�4 �Y+�&Y`k��<�W���������G����ʼ����6���k!P*����	�5eR=#��4�g�*�4��&�6�jʆ�ˆr�`B�N����@�Ђxgebkg�Z��9�M��^�LApE�ꑛ�-WG"e�l�M�ֈ��} zztE��m�R�B4C�����*Lv�b�~��mh���+����7�fǩ�צ7��6���Z�Θ�JI�p�Y8,�;��5�)5^�����O�|sV[_L9�hY�!u����10�j��my�|�)0�E�i0쁢�p꡻S�8`��:Tҧ8����.�uw �7ـF/&a�����K߆q��= k)�rgըz&���+	�ϴ�峽Ñi�$��	�ts��U�~�H8Լ;�*3jJ�ܰ��h���U�a��AQ�@FM׵�����M��jm��8��/F]G���C'pf��7��M�k�5��}U���5�C��evI����qN`��Ax�&���q��:�J��n�1cȪT�����xE�쀎��H������{�Q���+mV��OO�=+��BO �|:�_�����Ŵu���=)�'
J����� ��a��|@.h1;{�j��I2��儖��@7e^*�|ۑ�sN��3�Z���AyA���N�ACp~Ҙ���'HJ �����.�8��,f]r�3�"D��sn���b�����2>�c��������t#� �%5�`�m���O�� 22д]n�D	m����3շ�|�c^�I#�MV�Cp�|UP��']�u���:���
U�x^BQ'�w]�
�Y��P���)����y���h3]�pf]�*����ouiƌ��QZ�1�� �=]%>���{-ߣ��>^;#O�p�)E�qTܴo��<ۃ]���RX.�&�sq{XuT>U@�ڍ���O
��sC"i�[����cW��C2��T���O��[���-��ӕP�V&���`�j�8� ��ڑcb�a�=�I�O}���f�I�6T8�fJ�}����׷���sU��N sb�A �M���(�����\�W�������~�=�n��@+$��<�z#�1�Ī!�.��+�D>F� �H9W����s	8R��d�X7h��VEV�m�t��FR����b|��Q���樬��)�m0ܖ�zQ���͹���/��e@��ұ�X�/��װ���w�1hs�&y�-̞�d3領ߔ�f3x��*q�.P���������ó|M�=���t���A�N��<��w7
�t<�1��G�N����ػ��^h2�ax�?��H���K��t����r}��*���<�.ke�c��D3S�ȗ[�C՝�dz#�U�P��_k㙄��q�l��]\ݐ걼)<�#�>�q��:�����X6��h}�tO�*��!�jb;�e^3�����l'o�`�s�A!�H��xc�}������Rg�7Ȳ�1��	H�m���UJ(�1s����L
�Shq�͝�
���y��S7���^P)6�����j���b�#Գ"�^0b���5�،�R�A2�'.��U�v�֏C��Ns�8��~�`�H�HiA< 9$���~�'������"A�t�k��n��iv@,�z���ˬ���/,Fo̳�i=��<��MZ��zz��߽J�����δ�.?!>����G�ME%�ۭ�f�%��3����� ����p�%x�:*z_+d�\�C���ot��q��8 ��];�����vwuI;�L��g��5#6��mNA^�:G೒����q�_D���6J4A���
G�R�An�ﱷ\N�$F����z��������45�2i�L��EE{�xi��l(�(s-�[K���&��;BA��%����E�,�S��6|la�`LH��D�p{����Gf�jX~ϗ����.'��E�;l����`�����bĳ��aӉ�L���J����W1��Yw,F��˫��}F|��q�ЃY9j厷|	J�,�$4�����W痚���U�z�,rc.@�`Xq�D�/~���p�ݙ"C��m'��,�a�j����Q��+��L%b�c���$����(p�$"����;!&�aG�K%4��@�d��,|4��+��DDಢ�%�`�tGRՙ2?@���l;���2���OMl�
&��R�j]%?כs7�
�k�i�����F<��Z��4pI��J��i�,� M��fJbj����1�C��u0���qpG̹���+:1��(	�����6��2rf9a˵2��UkYd$.nEh���������ď f��?�	�;��!���*�LE�L������7rDH�l/�#����70zq3�>�������	3����"��k�D"U�5�`Z��� ���o�R�TD�b��0��i|�Ɣ��P%�PE��`���ۈ�7��-�t0�;3i��0ئ�Ƿ_��0�Eo��A5��&>�@W������V�ϭ��0�}�ї�b�5�|�q)Z��Mb�Vͳ��j��i_	y3�v'�?��tA��ӌi�	a����k������i(��ٟ>6��F]����sc��1�W� ��d%H�G2U�Uɟef��F�I����g��!"vD�m�|٧罩a�����=N��Lrq��@���/(����Q�;cr�y�+�dB����7G"E���������D-?	|�w� �ь��R��KӢ�c�r
oe��������A}3�O2��9�+n��L��#��`�CUHďo ��k�1�~���8P��	JA�)��o�"��S��rR��"�T�d1�yǬ��� ߐ�N*������Y��Qq�jHdXI��:��a�
�8u'�J�)�������f6�X������dpE�U�U>�O����~�Q|���&��x֞���g��n���y��'].��*y�M�=t�k^��
i�ץۺؕ#�VW3|���<4�TODUP#(�T�ԤA�
���m��Q4�}��Ѵ\=2��'�?�@�)�e9s}���=�1Ox@�y"����0ʢ��"}5f@�E����oE:
֪�/h�/��­�x:MD�����I��]�d��ۻL��a`��t�<qO4쨌�l�ѩ*z����5A%�R"���5z��Xõڐ��>&���LfgV�2V!�JK��'{ ��r8V�K*������{|�E�ޘ�seG��z��-eU�(Tܮ�1U��0�0����0�VI����zc;O�@kME�8���sjM��N={)������(�vA�)���"fD�=*/�~@�Mz��yO��j;�x��m5I���[:Y_t�Ui��,A���}ĝ����Q�M^��1gn9�q!g-s��}{��>j�����S�H���x��04�0(��9�Bx���̽y����&��Z=NXFRn�F��|/ݷ���Z!	me��|u����iCK�^+�����H�x�Y+�{�ږ��ؕ��+Sw��ГN�鑌��Q�j�@Lh�@S�� 8�Ve�B/�1weH|�=�#�=J�SU �5FإsMߟNkj�wc}i������$��#�D-���PRJ������_ea��#�t��ov��M��JE���i�?w��F�nDC��[0�m�WR *V�c`���b'ۖy�J7&7&��:��zh��A�JR�:'3{h_s]v�������+�܈{y�<O��X�-�~�~o~���G��p@�!U浜Ă����
�1���9��=��9����*��Z�T��ǉ�iy͞`c�XI�,�)@̵6��C%�PFn����߿��� ��C�zǊ�6�[��x2���hmV��qm���]?G���mf�������K��
6|��c�{d�#�FbxC�PၝtHcش�h�)t@]B�r(CׯN��)�*�킧e��40Dy��5
v��	�f���'�'����c��F�!xSf��?�3$�m^�y�O�A��׳6��q��?qA����.~��g.X�����d!B�`<tO�ڲ��6O<��L�5�*�~1�;Qj���	��z'�A���fڶ����9�R�L�<0��P�(�̄qf�L�'�oE�C�'��e�{�E�:G�;4�Q6�8��2��E�� fi����'6ށ���`vW`��b~nt̢a-7��CV��)l÷\)�./�X������א��R��f�J
"�|�����S�*�U�D���D:'�B���^&���`��v������f�>ܾ䀝��)��$��[��1}�󙅌�>����~�_�Lġr"[�����V$%P2�y��춒���|:�ܔPW�`ɒ��q��>_���M ��=&�?���#e�[���B���$<A��/,���~�ټ�  �h�>�{La"읞q�������iA�l4�փ~?���P9��.X��(�{q6������Fpi���E�p\�!O�x�F�!u�jqC�q�K����h�%�<2=���ѱ7�ִ�О��qL�i�]�z'�g!
��j���nQ�a � [����GD��k��!/.���rIO�<͜	-<:�7S*k�`
��U� �V���f���:��� #-���0j��E&�@�7�}{0��
+�./�.�f!�VJ�# m���R�� %�w��[�u�j=�Q5)_�r�^�Q��g�@7���!�,VM��QȒ9R�A,��ķ��c��i.��r�K��.s�����y�'0D�H��4F��p3�ܵ'�Hq��7�/)�H�}�P��~r#���g�e ���橐M��P\x6IN�i� W�R|j�_�b[�̠c��;�+�� �g��]���6�$�I�j�4�O޺�?�S��k;�P7u� 1������n�Uv���t��,ӳw�pl�� �X9�^�8
�����WQ��FX�e��ME�6w�?��vl Y?E,2rb2�q���O7%,���ro7$1�O�bM���ԩ�����x!��LdST%Aa*Ai�m�"�T[m`@gwy��^|���H��'�������뜓`�3pD>'�"H8�����!�6iMs)ii�Kq2�1[�� Y#��^�%
�A��v�Sm�̎��?4GԖ�W�2ʪDڣ�[})�.&\��	꾢܉�/s�/=��A�9*/��Ryl<J����>�~��lp�bjx;X�_��H\9ѡ��`J��W��݊Y.f,�"�(�:�ҴT�e�b�y ���<�
��u��83�U3Eڝ5���ҥ}d����I����d	�~N)�%��ya`"Sy�F�qR��{�wՔY�J&wX�!�	�_��韁���5�֕E�4Mo��H�����N��S�A_��~@F�|xE����D��ml��H���t�^�����Dy��\�6��i��eǫGs�G��1ܒ/�'|��~o�n�;x>e����a�K�[E�ʤ���	����F�d �{f����Q,��Pb���#����m�w��1W�a��E�:ψ�C�e�q���OVwEH�!R�"�䳳�����i| ���.���'��}�3f��@!�H�cQ�ɨS\(w_k��I8\]�Vl�b1��0�#kϨ�,�,?�v���]��(/��E���L��6�I���0�ͪv-»��d.�)����m�;0SK��f3޴'Li�������	ۑ��؄%�դ&�~�����J�``��P� _�O�2����Z)<��~��A��?q����R4g���N�u]h�Y\�-���1)pNWϾ{�r��"$6ˉ������w��C<g�)$c�lP��8��M�*�����0حm6p#װ�d�'˺�n߮�3m�6$�&/�NnW@LA�����d�@��O;���+�=Gz�,�'Ȁ���7]� v{�'���}����^���s8�
�ǩ�b}cŲ�/�$&d�l%�j�dj)F���W���ng�mk���.����3.�V���\����(B[eu�$��
�u�n���{�����b��c
�&@'��4��	�%��Bh����b_=}�`5��O�~t�E��x��K?�Vl9'&�b>9�m�b	
�Cʮ>��U?�WX� $����Ć�>K�$�;��X����gb�/��Oܣ^�Z]�����4��G1'��W�n��ӡXYR. �:{�HB$A�!|��
�d��(Ȍ��Zs�B�@��R/��A1��]3��N�"ʐe�w�d�������1>�"�=��_q�:��D�#���k�e ��ru��@�úC7!�Ǡ#��s&b�L�8�~���9����� x�@^��FK��(JÔ��i�v_�I6�����u���1�|
�h��bsd��L(/�뼃�-"	�Dh�(��}�Ԗ�������C�sQ/���0��
c -��\�S�<�x�t�@/��Xa��D[�a,u���_؏���D� I���'��B�L�3��C��BV4�ѭQ����m	Bst	�Z�y�~ؽ�Ԝ�"������^J�v�ԛ�Z�~�ݤ����-��n����D0�>���6���d����ߗ�ζ'�e�s���Vs �7�~=���N.�����4Ȏ���GA_��V�v"�&y3r:�����j�l��ww�knkFO����۞D���}�3��MB���ǩ�Ȃ������7�73�
���J^�+��#���9 1���ۨ7��8��1:fH�8\�ޙ�N�>"�ο����[5]FRb��MH畩�_���xI;:�ھ��H�sǼ@q�D>��		=�d:�Ԙo�cjA����r�1@�!���� �E�&Yt:ˋm�R���;�,��9�ʸ��п�F�?��y�{C�#v�D��*:|R���Ń�ܝ�qI�[�ΐ�E�W6f�a5vl(�����P��t9��؉n]��K��ߑ_@EeH�������(p&���@Z�rghYO�v̈`1������ٰBG�kX�Y��W9�����������5�V�vM�ݩhːO��r9g�X�l�B�h�[�l���,����#a������)r2LK��#��(� �����-����٤��J���o_ЏcG�M��e��wD5���I�'�Ň1���=S�sU.O��|��6M�7an�C�n��x�U���._s�,2c�!7M?��їg7�Y����k��V��z?`y����I���^���|:x��@CV�ՖAG�z�qP�`��D|{wi+�k��~���	�I!�O�P��T@FoB��?�%]�2������S�Ka{a��!��v�
�s �D���O�6@B{r���=7K���#O��l�i�h�.�3>:̓�4ϋ�#K��l��fS^�}TQB	���w��8�����ߌ�p�T��GΒ6Uw�>k���gO1镝�6�ٵ�sɊ��ܖ�!M�b͠������x��� Ɠn@��Q��2�8x�����AkaBz*?�  d���������-�=T�$Pv6RV�/8�}9L�wF���2E�4!/�����ɏ���L�5�{>���%n��_���Fbl�"�d�5��VV��{0�#K�leY �T�!����y>��.#��9֖�!�w�փ+��!#��(�U���ݣ��iC%S7;�H?�"�+�KJ^��<�������0-���{��(CTrQ�&��5h�T�!Wf�.���9�uW�(���!�<;n�HC�	W|7�)�Mъ��O�Z�������|��ʓ�IM2Չ�K��%C�ž�"��[ƭ�m�mY��'Ƹݘ�S���7
�CLs~Tϳ�e����s�OT!�����I��j����ϋ+�V�U�m�F�qñ��ֆ���2��=k�/��xaO����4Y�fA	\H�����!]�y�m�1�--���h�J��<A=����J&i6����2����G:�$�k�ʺ��
�z�F����������F)}ug}rۛq�Sa� FE����R9Ʊa*
�1?����Z���op&�1P@u��T�$�z��D��ͩ]�W>6��KGN���;l"��tmF��9�ЖK���3�s�>A\f�����,T�$� ���+z䨋�����n��)�n�d2(�~u�_R�&ߢ�ֲ%bUaJ��fC��ض2%|�D���B��u5j�p-6��{g�v�;���U�Q�h,~�çLc^IdP���vͤ�yk��\K���R�i�7pS<d���/�Gd(�}�P81�"Ưuf���C�y������>�-oW���bJ�k�MS�K/����qLN�^�����M-��ɒ��f����S��Oȋ��s���Y_B��T�|b��c*�4D%.���Y��N�;I���߃2V����!���#�#P��?`boHxV�̛�%r$܍���,&!��@�M5�Pa�$��ѹ7�������<�	���\G=\9㌗Gs`�?i��O�7h��"a�d��Ѩ�$��5� /�u�>\��)\�=�N�"*�!Ps���R�·�����_re2���=.z��rL��ʷ�B�J��y�� ^d���7&�Va�`���eb�Ḽ���T�Ji�_+�w�W���t��%A�"�6+���99F�~	���>��X�;��Q)ab��H1G6�$�t��dFW�5
�ڿA5U��a�a��M�?c�$ۓ�g&҄Q���	}��<��ujʡ�k���������U�M,p!3(�8$�4��a���AM�n�HiX��}6)ׇ6��vh4����}�g����'#ֈ]���H��� ��।]m���'�*z-��U���)e��e�����*��-O�
��Ť$4m��qF���ߗ(��N 0Ӥu���=Ȏ]���P���{��h@�	^K���C�2߳���|yw}��@�-R�i�cv7sZW/t�����%.�/���T��ғ��cz�gL�ǳ���!�O쁛 ��o����>�ߘ�w/~��pCFO��_DwHg�>��C��~����κ���%/-���V�z���-�8e�ևB�[�e�6�;�=jl5d��e�ͬ�x��}��y�O�^�>���Ң��8�Oeǋ��oͭϓ  8G]y+�r�댗���ΡH%��w� �Q�l�'H,&L�_!�ق��"օҝ�������(���
���m�~2B!4���:5p�(H{|8w#=5ۨʋ����,�Gv��Αm�Y{���)��� ��`E��xQ��e�oa��2�fK�z+q������5�$<o��G���ݞ�,F��.?(�
��KO�wg�5˅�ގ�<k�i�{��2�!�5Ȇg����; �R�8�MZ��7,�Ϻ��>�jT�_ވՐ>����ukhv��_̷>�Qb+p�
�q�C����kI���!cy*��ww��<3qB��+<̒�h1J�{�4�E��+���X+S�r.��
X�	�)�'��e��&��>�V$:.U�;��ҿ��mIb�e0MI���κ����i�<�ȼ���J�ѽ�/r�tOkh���i�[n3�P?�_�Jsʟ���08���Ŗ�U�>ڻ.3#���T���ɗ��}�Ѷ�fm	�$5�GNw��Q�}R��[���CԼ
�=̅���2�ȡ��ϊ�d�ɳҵ�>Q:*����^m���C���F[ �,��|Z�q�H�"����n}�I�|Y��+"�W��@��d��a�<$�z�~�F����&��
R��m�E6���#؟a�Nkyp�I��G�l�Ԇc�VW)��r�*�5�Zٸ��:`�E��3P;}��|����봖�^�G�Ty��Qd�f5dFRnn��|��h:H�,=��|{�p�NO�ē��N�1��GNx���I��Nle�y�TuE(����1 ��J��^0�q.���
ȍ]�+E�)o�C�D���_���dF尺_J�x�ǚt�/�,慟l��g�^���{��e���qB�NtQ��Fx���X���k�_��N��>�懶�i�L!�I�Ba��OU�R���U������bSGv��*��Q�Wc6�C#��b�ƺK����?�NdrEh�љ�m�)jaz0�ve�u!�RYz��$����I�$E�??�/I��
�Z��~��)^&��T1٣)蛛(y��	�F�=��wp����{H!Ɠ�lW�az]�!����C;V��3�S�����j�1��j�'�D��GdP�#
���l���a��/�W=�1�ĳ����|h�1b�}l�{��"�z���'��Z�b:?�]�k��A�"Rք�E"��!�y������u7/��n�p���ٍf��\ CN��J@�S8��xߎ�[���@e��~�4�F`��U��d�0�Lm�y�GU��O$�����y�g&%PG���GOS4/R�Jյz�t%��N�d�Q�7
�l�0ӤA�z�i�S�U�Tnu� K�~Q�U�9t�"�SO��wbPЙ��ը@�H�bb�����vx`A���DY2X�b���L�?���(�g�P&0M�d�E�U�~�ح��Q�&A�= �uP��9]�_[���ᰵ{v�ޏ1V�9%��ջ�?��C��������J,���y6�4�!tw:��ƹ� �����)K�k�-�d�VO]C�+��e3��C�;����FA+���ŹɈb�#�=y��W��\/��s�u�t���ר�"���T�q7\ďԶ׷�I�	t{�� C�¸���~溧��`x,�j猪��Ө��Z�����G��n�{����x���C��\%K��7DV���&?{���/C$�ti���k����*��%8?\�0�s�gYu�~~���n�p�҂ )h��_���/i� B��H����	����� ˜�'9λ�K���R��oU��]/U& :"�
�S0�΢S�Te� �I��xq�!XOG,������n�	mpl��J۩jbyH䯜�ޓ_���k�VA֢�@f.&��z�*)�K o�b�BH����yͿ�sS�{���w&���+Wޙ����'�Io�A�G�r��6�O^-o$��G-�g�E�@���H���L&}1�/�R3 .Ng�oE�r��f�n�5��Z��Nr�,>����6X�z�� "���O�MM�m%��0H�^�2��f3=S<G�.�Jֲ�5�3U-��Q��o8U�R:=ī2������$i�����~`�Z	!a��juf�;DXl.
�57��]<�α	9G���Vc��I2�4�N�_n�������Z�t��1��3���2�f@'0G��O.b�R�ֹ[}�}w�̤˛�yŞ5F3~-�Ȧ�5��掐9͘&z�������
�mJ�W,�o�(Մ\���|h|L�"���E�)�mp����f�� �i��:�6P��bD��j�����d�M�� ��¾��?S7C��q��ו�|�"!��z���A��:���jԼ&Evm�� ��ϣUd۷�{i/�vk�xҕs;��a� jvF��,D#4(�Z<:	.�����/+ f0=��Ҟ	(�
�+�׃KPKl�$���p��:����pEn>��$�3"J����}�_=z^z����	�Pe���BY�k��4"`���_��*j=;#�b���:�lXG�"���P�Sq�%�(++I��;�2��h�����n�(�`z��l�K�J|��!���J�Ī����I3p�m�Щ��� <�X�m�Gi���;�F�R�<}�]Q'�j�V����1xk���;�# �-��r��J����Y�/�x��"�){�[�v�^���{X
�w� X��։k1ϣ*���u=�VK���˩Vc.J�6 X�T�a e�֠���B�[��G�L���ߕ��<��F���z��Xn��(�k�G$y�-f�Z�t���!� ����]Y<�Nu�rU3;a��DS�C���c���H�˚��� s1��'��1�{ü�
+����v��?��S!)�}��"c�������ݶ��膎H�N=��g��Ǿ�Xt��t����C�x��|SP��F��%	κ�T�z��z��O(���M>�Zw��a�M:����=�j^���s:�܎�PL����{0��v���s�U䆐4�s.�3�ۓTB��F�u�G�L�W�"�Q50,b��o(J@�_�5($���=$��K5����x?��������d�8���|�gj�Š��֞��/��cX�h�}�e���R�b���zr���@��8�v���*��1�֧wE߼��N�6D�C����7/���:tk�,0��-D�ⱻ�	�WQ	Y'��Q�%�P�����j���?���b����l��5.y7+ż�7��G��}����f�Z�7N6ҭ=c7��&�!�hG����tԌ<�3�YS�M��[�(.	�c{�^�rI;�
f�W^�l���w@va��PD�~�����66�;/�]����B�V�]�mn�ni��I"9\�*_�ׅs��7.�VW�/�Q�d�~2xHʀ�B��Ft��L�"�K��'_�g��������|J�>�;��v��wps��H����`L;p���>;���~aS�S�ML��ŉ�u�r����9�a�����l�E�1o�.��0
!u�sn\�'��R���ʟ�7�x47i�./�]��D<�}K��Z5N>;!�bآ&�H�'=3S�'p~L��?F|�N��Jy[@0%�� �_��>ܦV�s�y���~�+=�g
l}���x�(t�߰�L?���m6��tr��	n]T�������6�,7��z�	\��߈� ������w���� �I��H@N�DK�9)С4뚦���{եZ,i|:6E�6� �&bA>�a�2c���b�E�J_��� ���j�"��f�3��я�������Ĺ�̈́���j�>��42�g�e��r ���*V";) һ�8�_rM۷�v�T�h�vw%�~vA���J�D��D����Y�.9x�{%�J/ym�ٯ�޸�xjH"�s�B�da�� �����p�JK���#�#��o㐃xM��?��^��ʧn���X�QI��G��������A#>��Ό,9�l����^}�c��Ro��8&���]N����y1���*7��z$�a��/�#䶿���i��Qd�D
�P~�j��y��.X���b�El�	�i�Q��@��o�I���&l���uX_�z���PR���Ͼ���N	V��{�2�%G�F��Y��Wnt����LԞ\,���C�m��-w����U�mH%,�МɢOG*�؛{�4�@M�B���㸢����]I֌�����\�q� 
�2{l�c�I�� >��#ޣ�N�XPnRn�JϬ����J^2ɵ�:��!����H�PK^iRv��&�H"�V'��Q��i����)�B��+��iN#5��G�z��߄��kK�<1[���3>�0��|f����ЃB2;(��O�o5Qs�6#p2Q��QV�1�<�X�c��$�����&��":�	�R{��}	�Y���la��l���a��h��
�Q⹜ڻ������F`c����g/�V�[~����L�l��b\D5�x5Ւ��!�@<ʨA�
pUBW+��D��2(}�3�ԓZ���L+�O�^��|���4�t��{�ӹyJgE�Iz�b��E��(�yG��^m����(����GN@�j8̤5pD�#�����>R�][�*���F5��ʣ	G��1č"��;�$I��1ܥ�x��Bd��)n1��"���	fR�y�gg��� K�~]-g
��2s��V��7Z_}��x�|�#}�,!�O"�ݱA�=_�~[�'�b�JP�s+k�T*���q�FAcUۣ�Q6��!�kB;�f)`/&���*�Km��x6#tf�o�'a<�/8ʋ'����ܖ�s���y�t��z��|(,R�b�PG�����)C��/�����g�"�J2���MyGd8�u�Z�4��+bK�S3	ChK(u,��ɋ�� u�K@��8�eK+�	�q�V�"p�Ro�9�)�e���j'���z|�p#1��F���׭vث���
�ܚ��Z���oU�)�3z�/9� ��h ���D�p*oǑ}'�E�B�닒�Y���ӷ�-�]�+������� :.+���Q��L'4g�,�3#�\��$H�ע0�������I9c�g@.	$UX.��bY#�W��{ �xb�*��
t�]�lF2n� F' �1������'�a���rB5��-e�M�-6�,��tn���y�a�8V������x���b�����_�ܾ����*;�vPb)�����n9)}��̇{'}���s��1�P��(H,�{��c&Ɂci\P5T��9�SeL,��M5�Cs1`��a�'	m�7��@|t�`J�NK������\ߺ�f!���e'Pŏ�BiRR�������G��j�{#�7�C�s�ە0����k����!_wE����]LSA�k��D?3����k�`�:��V<�]�7��@YR^CTmw�9��$c�\�&�j/Fc&h�:IV#?[�!4.�|t_�@ֈx�_�I�1�D/S��qvⲟi�����^P�P�if�:����!��0�����9�3)�$%���@���w���`?k�!�V�I߽��\�9������DXTDdًȢ�1�ʡ�lB�� ,����"��%�cLo�4y �R����wWk+4c_����RkF��n�˗;�����ᅝNc��|}K�B�{PZ��nC:����߁/L9�5��,��n2I��\�Ԑ](����Z�}B����qL�ߩ㏔�)95�R_=Q��_o�}��� �D�ټ�I�xm3�Kz���AjLތ���f��?������٨��M�����/.�N-��4�9)����
U:����6�aAz�Kw�({d���D����ܒ���d�T{!� [wK���f=#�Q,����`�7��ML�~��ˑz�Fn�N�"|(�K��=�QX_1N '7w�@�(�㼺
��(�$9��+q�7>�\�Ltܡ�0�p���jb���'I�q��+ثjx���%�s@פ�u�9���x犒D���ze}�`o�Dr�����
�'����a9>Ǎ)���}�:$�	5f������������+�Oax��H����r�GAEƾ���&9����H>&�w ��������e���9�"�m�0ie�
b�&y63�/n�!�E���/��U��ɗər�o�(�yw�������Wb��V�����W�)K��T�LP��\B	�//J� �@�=�l�?�)�4wN���F�L� ��]���$��랻�T�����^�[�3�W	31&�æO��я��̿=��?��Ϙ�a��<,�IO��D,��>��^��vZMw�|#�  J�]g�p�+A�0�mV�rD���c\ʨ�w0��Y����:J&Ʀ ���[n2UK�ţҒ�����w,�~��oܓ�I�Y��fre��f�o!�u^-,YO{�lwz�}�2P�:�9��?]���u\wɮ��G����]����9�g�u��>"Ĳ ��
1���fat�ة/R�X;������?��*q��������r)�=7�$��x�
M=�s$R�e�����sCW�!�?��B���i&;$g,��e����^��l�ۥ]�Uw�*�q#�>��})�#K�@�$��+cE�b��*=]�{br��t.�nO{u���hu��|#���<��@�r��m��V�&J�CfEЙIϥ���o]�jBE�d��(ZGj��M<����QG�V�'6e�]l�F`�c����
z9@i���d 8-�eS��&��(���{o���Ȩ�������=kĳɣ4�#�?�L�|�hD)��Xv�F�w�.�����'�H`E���6Ǟ�?U�T/��g�=�fb)s�4���dɂ�%42����ɉX&Z1��eBif���6^��&V����p5���c���;N�漏��+��ezϱ����۫�8�����D>h����HWW���E$MD7���1U)��Q�'�ԧ�s~��8�`G�D���a��:�@
(�#GH��R�+E�F�B��{��+�G���Z!>�-ܪznt˲EWY�u��X��E���=�Ϩ$ ��og}����&,� Ȁ�8LV���+��dw�cS�&M�LZNzrN�T�n�2���	� �^]��dv�O�5q��LǲG��(�y�?���f�w�t����E�q��ܥ�nw��O��Hl�EJ�e�G�q]A�8��M	�P�����}9��aS����.6����6����3ӗ�N�u��~ S��0�%�����jO�±��tf:˗��	R��荴�uثd��&	�7��{nϤ~��u�(���Q�x������P���?�@���ۀ�1lx��_�e�x{��U���A��-n5'Uzn�z-��mF�Fϕr��s�?�<o��ǘ��5,&!�D�Yn����um��({���v`A<���f����*9���I��V)�4HY���.��O*����u�b6Z	���s��Ue����&헥�-��*1�6�U
�m�a�Q�Tm<;�Ʉ���Y�
������Ɲ6��z���l~XX����ȟ4��ҭ�(�����ǆ��VA�����8y`B�m��'�E��@~
�#]���Z�x?6��B���p�?�c��'���Ј�s���V�qMXF]�3B�'^�X�� �X�#3�]<�I�ߴ�&�r\l,br a�]�%anXiۼ�q�G�[]���Y�����=��V_��E7'6�j�_�+;���]�9��w_��ZŹ�p���No`stө��0)�h�QԀ1�ܣ�Y�w��qEb����L�*�� 3�� ��Eq/B�/@�8�C���]���_Z���1�����֟�_XT��1����h����
��6�@�3��4��q?����\�>ԛ�!m4+0�"�mö���(�!E�����F�tqx����܆F��B_�è�~�0�J6s?!���a�u������7���@g�/7n<.�r�vdu���*��M|��9%����|h��Ig]xsa�a���3��Q���:�#K=]Np8��*�ߖ�8��.��o%���9����vx�!�kiQ!������h�M
�9g�!�b*
��:ό�@��	���f�� 8�%6���ؙ۳kWe_�����?Ӭ�Ѵ����7u��'Ӱ�A���r< ���|�������8��[Y�@�D(�*%^��<�׎��wc��.u����o���wa��~9�!(��>�j'%\���U�L�G�I��T�)�����1if6i0��|�W�b�C�/X噀�8Ng�T(1l��9�1݄�E�_���5���B�ŝ�٩�(�Kg}o�E_}��:(.�~` Xg��n5��ނ(6�|���,,?��(6]����
5��� 2Ы���sֺI��ͽ�-Dh��|mΞ[�Rlp��f�oя��bR��w�1\<,�V��k��=�}e�^�c��E!�YX��^v������s�G]ʎ5�fk�[ʊ��و�%�<xO7��\�l0��b{�j3~!����߿�zI]|�ZZ94T� �ȧ��ZG�i�:�����F��o�c� Ή����kZO� K@�/n{�OZ����L�:%M$$z �_A�`:-����z�XA+]�;��v���d�h� y���i�O�z��R��~�`
}ұE ��PUI��x�����s\����`A +�^-Ǜ�q����>�Pa�]��9�L�Jܯ���X�N����l{�B� �e��H�7?Ei]
G�`;^O�R�����M'B~v��\����꘭�H�{�c����O��      L  �sN�t&�u[E"͊�;B�$�Taj��n6D�߮w@�R]l^�����I'1N���Z����f�g�#\�a�O�xq�$�L����8&��Z����0�D��bi��Ũ�~�^D1ջ�w�7}�X���z���F����Rk$��g�I��g�R}�ҵS��@?�vh֙�"}\^���!r���тls��B9<�1�S��5��N�&@΋ꚇ�:�an鲗X�k�\9���S���d��ǽ�00�ST�ᑐOcħ~:����ׁ0�� V"�6�#�FKo�� _8���}UB��������u�%pq��bO[`G��y4��"��Q�#��6V���'$ouQ9��j :=��5?��{�A͗�U>��$�`�{C���:;E����Pn��4�1����a�MX��	��V��lf�ś�xҷZm���uD=�z��S��a���Ee>w"VKnӱ?�]�Ѐ`�*}j��+V����*J��
Rb5�<v�m��U{D���4��?6��|M$��{P��v ������'5�vf���M���%H�{�&a2�'��\J�a��L��t��z�5y�ԅ�R2�!
��S&�����fv��['q'6Oj1�-�Qz���N �.0T���b*��s#�r�[��
�x��U4�QE��H�C٭�Ox ��HAҬ�A�#vHRiҍM9@��ۧ�&����)b l՛$��AT��$�P�/�ԧ�A��=�7�F���c�e8*Q4U��J�@�+Ө��G�7:����a��V����c�W��❑�nD���03l&U���Љ���n��N$ғ��<O,}���I�>���e�-��^�*Iգ�{do�W c"�sHf�K�է�B_�b	���*ZT�# �����Q=����{�&���L�p�����&H�ѧ��]���WR��n$w�"(��R�oS8>!X<c�2#�9`�2qP������l�l�v�j �D���K�'K�\�2����#J�������ѢvВ�<`�Gdh�l7N>7��S6u�LFL�:x��6�p.��|�ӽd��:M�']Eg�}��=�S'��YH������g;ᩰw��G@�řE߆�V�B0s���=^�w�޺�f���49h�d.�����d���I��Z�kzl���vJ�����Ub��ӫq�4Ԃuu�Z5e��e��f�󊦜�#�z�3��i	� m�'����l��9[�9��F��;9�
~��4���
A�_�m��b�!5X	N�!�N�i�L9��<�>m�FLB�(�Y�n;@��v�"B�+x ��y6c�M�w�
��1��=���J���b�l?�
m�i�6�ȃjVM����y�T�G@��S�JK��X3P��G1�6x>Þ�e��Z]��loE��*�B������K9����Cė��u����!��N��88���>�E�򱈚���͍���|Pn�&X��2Q� u�_x���ZX�ވ�n^pHa�Q9�`��	7 �3��e�����9���n�Rv�hQp�,-ߜ��2�"�g�N��#R1Y���A�_�d<X}x��5��(,˦�_I�w~4�w^���H�Zq�:$�OA����W�l3)RW����^D��i]{|�M�,�Q�_m�yU��:&S�U�R���j��t�6�����L��s�q�*�?�J�m�H{�I����}O	�R)���"Ѹ^-/�l��5�#��A��Z#�o���#�_��_�dD�\0��4U�=5���ٔ|�J&Cm���\�V���RZ`\L��1�4ËF����|��)�y� /��UA>wwgP�ߑ7�3Fu�xf���A��[ߏRB�8�/�3� �ppr���}8Vsh�l&l��g�&�l��4(|Z�U�( U�+t!{S �y�8egc[O�Jҹ� ֌�̹=):,OL��IiK�5%�]ĝF|a����Ѿ�&�Wai��=��מ&+t�2,γ�p���x��������B5Q���D�����W.�w=6:�����������b
�]_��� �>�<-���Ӥ�����e-��)��~㉱?�8<���	z)��\`A��(��4����st ���v�8�O�!�Za�� ӌ��a_W&ߝz��Kl&���R�.쪈�Q,�,�/c�k�3Z��b�pw�/��j�����l�J_�+8����O��D�Ol?�2��T�(^��������T�d�c�k!�r�ъ�`��i�>w�1Z�<��)�ـ
b���p��w�/<��ɂ[f�|"�տƗ�'�b�f8�V������n�q���*���sӶ�w`��Cɉ�7�չ�Z��V���ø���Z)ɂ1˘�q�:�š�Z�d�����\��|CA�ǠV�\���sF���2�`^P�Wu4�M�-NSt]c!����M��������9ޗ��_�jH3`~z8$͟@�d�W��4�[��?2W�G���:f'���b{%� ]@11YW�8t��K�'�9�T>��P0A*�Z7��.d���e/�� >���GCI�x����2
��� ��I�Ot��ˏrlĮ���h�s�{x�]@"h+"��r���f|��^������cOo^�-q2K�@�m���/�N�����Q����.��y6iD���~�a�����S���˅BO�� �C_��[ُ<�KZ4��K��E����V&���t���&��NL���INp<a;�AGO�G��δ�=5i�y�ͼf�׆�2ʨ��r��lW��
��q�SJk#��`ǂ�Ֆ׏>�K�E|��4�y�y�C�����fib82W�=a���pjÂv��$�+\bH� �|Ydw���g���V�|��%*sp���^G�QW%�	�"t���s�吗/��	E��&���3;�����"��r�� -9A�zyVJ{�2����fT>��5}�!����>�4Hc�T�-k���K��f� X��H��{�Ԍ|�]H�������R�N���y����5��A�:$o�=a �6y�$�h��/v��qtE�%@E����>Ǧ��Й ���>���>H��� ������˪~�a����ҭ4u� 	dq�x��=&�zl�/�N?Qd������6	�L-�\�CC�eAF�X/�y��Q�� 5($!��L�l�v�!���C�"K/�v��]
e"���g6�Z>�_i�+	z�I�{�R!.��_�H��l瑖�1���݈�:���}`ğ��' ;��Xzx`o��j�r ��0�C��C.��x�PZD[*��������<�ۍk;9(cx��>���M�G�4u�u����ReQ����j��y���d�${�.�v ����nn���И�g����V��QOD�d0����
����E��}ʣ�����4�S��C���;Jh��HCa��2GOO���\�O_s͓��`�4,��G�+<�LN��U���a��Dssw���SL�B�kP��:^׌.]���7�W��&�b��g1��ֻ��.{e
�ayR'PE�N=������ܰr��È@�R{�,Y�/&
�D{�m	���x��fX�F�"��\���50Z��7f%W@ ��{a�in��Ry5XϞߖ�~���������WR�T�m㞈�|%��8߇��ef%�kl;:x�{eA�q%��i�٠8������^��҇�-���9�];���kd�T5��E��^Д�*�ī;v-�A1��g��mw�1�Sz!g��2�3� ,AY
8:y��ӗ������n� ��\� x.Ov3�g��u��Oӌ�^6;�����r�p:5"��� bRYǸ����h:�D�9����t���Q�����O#GM����2���U��;3��?�(~w&�SeN��#̑���>�@VZ�O0�a����0N��V�s[���!�A��:��q^��w����d�L*w�d�����L��~c
1�ک��K�e���-�^$p���2�bں}
�h��'����Zb�4+��6,� �z��������!:X�V�k���fať�u�>W谛A߅���P~#z ���%W�=,��A4/����,�W��qQ؋<�o����k�^Ue1c�&U�<HR9�[�a�jy�>��c��\/���ׂ�������+��)���P�T�X�/;Z���mAe'hxi҆պ�`���y��zJ�2�oD�̀�J�<z�CU.��-O�W�R�I�F#8/쯲g�T;g#4�-��.&�O�<����$U���9�#�"�#�?JSE�^����N�>��Y[��Aƶ{�`�$�pY��HT�4+*=5��%�/����D�HجSp�Yf�-aدi�<K�3�8%��=�QGA�:|��/���낢f�D���:-+�2*�/zO�}`%��Ί�2�>~��� �6?����e#��
���[mHw_��
�҈x
_�4qNi�~C�~W�a>stq���n�ڧ}5.TF*�� UT��H�2^�q���R�;�Qa�8eN7��N�v�������12�n���T�I|��l ��Gkf�OHI.�R�5
�"[�*�~�y�<�Ξ�Efҋj.�\4�MhU�=R`C}0y�$"w�Nr�_�������Nq�'������	���?�$���P�S#���	o�$�}:����2U^xU&�2���o5!��tR��:�E&�R�"������!�}��
_B耮��ǑX���� w�;��������CN��RsG��H�7���[��Ṣ2����ԑ^֗�7+;Y�?�7=֥�v�VxR	SDAL�=;K+���S��9�/=/�{�ooa����ݲ�%Oxe�#u½�p���TL��.oe.��zl_=�&7%�Fx���>R�B�8shA=S8��\��s)��d�ĐdKr`W���c9����͕+ȴ��K,��RAr��w_����n��K\ԐYv�i@X��v̝���Rg��v������#3r��-Oi�[l�f�1�L��Ǩ��"+�"�鱇��[��({�.��=�F���Ƣ���;�	+5-�$�>� ���7XӲah=�և["S�Ц�}��o��,R0~S�q��J����jg�w��[2$�̖���G���?U����Y�u�q�(�fu�ho��X�c.�jzWَ�\�r��8��`��Ƶ����F����ڱ00l��ޑ/�]�NA��n��W���� `��lɵ�%',RMYzu�^���B#m&�W�'e�MӬ= ^FsH��x�|R>6�_YN挟���U���"��"����F>���h�?<}�؂�������e�B�"�P����a(z^�z��k���������{`����'��֖sz��.�M�2mԹ�c��AS%fg�GL�zV�@Z��xo'!/^LMOv��,y��\v����ւ���D�� ���'u+�o��u�u��Tg�������n�?�y���5:ʫ�3դ�2@���)��$�SY�,3b."F���Ϙj��Ye�6M��E!��I 6�5�~^w����E���ģ�6x�������7�"J��~�7��ُ��,��NF�$.H=����:: =,�(GCD�}��*H*�@��>,�_���7�œ�<X���k�a�t�4鎟(@�Y�
�7�Z'��6��� 6�% W9Q�?@���B��g��$��f;ÃY��q�"(*��z����A=|�����9��vd���oI@<���E:�����1���i���U'���V��k�ig
Ό� s�.�-˨	�����Z�V��i�����Z'�:�;�DC���*=<U�;P��=�hb�w��Ơ�<]�u	�����xH�,o؆8}����*7��ޯ�2�J~��b����_�sA&�nI ��l���^���㚇��j��\��h����#>�'3r��}y͐~T�Ɩ�ݚ$ئ�.�:�pC��S`?E��r�e)������aǸ�ɣ���ۉ� ��V��V��m�7�,�#�t4w��xɍ p�<g�/ �|�E�����6�7k��&�4�t8�q��6��*��f;ٞS���������r;O@J�G�7��ꀊ�G*��^w	�ï�f�]v��v�@��������u�|��p$�Z#�77��h�p��f��[u�$z#�+��E3�^�y"��w���P+˷���%��Z�!mї�)����=W�g.y��;\������=����/�[�@�'�Q|E���#�Mߧ��?�F�E��;d&w
*�Ӯ��/)� ����J�[^�Gn	��i�>?3�⺙�)�p�����̡��3��U�}��G|� �1a+�դG���+#p��*�;��}fP�X97Y�����DF�1U�g̎�t%�!�q�2�u�#����ɸv�j��JbH
������(����	�n�����`X�h�]���0>�.U+���9T;�3�	̓\L�R���0(;V*�]�#�j�-a�B���8�%� 0�?�����,\��� ����{�:���)ʌ��s�b����(�:�ڞn�wh�+Y)��n���,\;�Qrʿ�#���=���(c�mm�k���V�~��6ߎ}䘑�u��#����i��gE� m�X�gQ�G�6�����Y�ޅ��Ei��u96�~u�X\�g�LҮ�Sf0=A#2I�������N���G��x�!����G<���|0^�0�m�^�G}�Ȁ��x@
�;)������= u��YY�+�2�1}�>����SV�%�������)����ZT����5�nMӢ���:����@b�f�s�9;�ZkA��Fv����]�äLg!0N�>g���&��Ǜk�6g,��6��GcL��O��n�i�ZV�b�%U��Gp
! ��x�?��l��q�.l��4�J�V�-hk[=4��>&�y�mwC�����������,�z_�ؼ�xka�"��E} (!��2̨�\�V����\4!5=C�Je��p	#�L�����v����vƐ
��F� �#J[�*����S��$i����-S4 y��m}E���/Q�������㶷M��
�3@�i�vf(|��m�s��f<��JRm��_��]_�$��@�|�6#3o&�&Դ75��9Hr��wĹ<��Vy���S]�68��
�Tͬ �c�V:��7U�L��O�V2|��\;gC
�rr.[zI8�'�5�3�#�ʳ�� 꽭�3���ٶ�d�[f���j~���CƖ�'��k_%_P����Ӈ�Sz秭$�ӷIN.����虼i�,x�cVL��ꗋr�cY)�/����ߪ�],�z���RݢP@&��҄�Z���H���61�w4\l��8�%���dڠ�_T&;���M�V�#R}��tv٥�1{i������m��.I�w*�vs>|�O{�6��&�ZnkfF�*���Y�����o0��8�`G���
a`=��e���)���Ğh�nBRT�<]#+�y&��܉r�	]�B�A�@Y񖃌��d��Z&�a}6.�?�5�7�ch'��+s���~�����ѭ_�	1�T��8#ctL�Џ�n4I�Q�ј�tRsl�u"���"�e?�j-`���'�e��-� ���㷁89�����	RxaM��rF;�����V�r��"P�#�ϬI�Ȟ����n_0�K�@���,^�������[�uI�	þFb4("e����q&�AG�=�.��~�[�T:+7����#T�}x*+�TA���l|�1?�Q����6F�}+tm�@C$晅Qn%y�}��XQ
0�}>�?�;is�_�� \�׊t��6�M��Ty�#@��.ғ
TJ)'�weit�$5*�G�}3s�;��ژ��; ��jȍ ���e*����]��+H@a�ѫ�PJ�;[� ����z�x��iĪ���(Y�տs���q0o��%�s*����hga��"���ݎ���j��쐖@r��NɋN�i���NJ��G���7y����T��.!���0v$C0ֹ8JޖQx��:��U�>7��Zi��^x9%����mMWO�y{�č<2���c �t�3M�w���A_L����
�*��2(x�A|[t��#���r�<Y�ț��)T,�D9��_X�.��V��������˥���k]��F��'@e�X�l.0�x+B7��QցYl��'Q���Y;�Ņt���dj�j���0�O��e��o&�ӑ�'8��ZM�bϠ�̶Z՞��`�U���&?��4u����R��rotK5�	��4�Dx@"H���*�R��CA�w�䆑S�Fp�My��|4{���������)^;8��"e^�ȩM�؆�����M �T7D���T���ԳB��x-'5�NΓu�c�����DW=#�QN�`�$�?��?>�L"5#��N��qJ���c�4��o�5�H5��
k6[ï#:��l�ߍ�v����������Љ"�>$��f�sq���>9��xZL�۵b�:<l���`)}�� ~����B"�>P��B M:��gZ�|]y3�x�H���Y��󠂿uJ1B�bH��zu�2�2�N��_�����K(����|
W"�$)V~�3EIǾ�*]�i���3C�����b����K�V5x[���z�<7��1�<!U�]�G �	}`�v�)	 ±��q�<q�����Wl��!jjZ�km�~�E+.T�"8�|atF�Y?b�E4M9�!�~=<:O�.����4�E�����>Jb��NOՌ�5��Qu������jxZ� ��a���?��,=b�Fn���a�/����D������,|��]�9m��d�%�t��}	��WY�L������45�\�<-I�b�͈˚=ܒ̰�x,)~ђMҤM�"�l��y�i�����j��T��������m    `�    �,$���|$(u�D$$���  ����  ���  �  ��  ���  3�j@h   h   j ��q  ���  �  � `���  ���  �47$�t7$��a���<7 uڃ��   t���   t�1  �t7Sj@h   h�  j ��q  ��  [`���  V��  ��a��  ���@�8u�@�8��  ����   �rV��i  �u�%  ����   ���  ���.��   � P���  �m  ����   ���   ����   �8 u��F�> u�F���8��  ����   �>u�h @  h�  ��  ��u  h �  j ��  ��u  h �  j ���  ��u  �   �  a騻���a�`���  @<���   ��  �@��  �   ��i  �������I�� w�a�`���  Pj@h   ���  ��y  ǅ�   ���  @<f@���X��  �H���  Pj@QS��y  a�`���  �tw���  ���  ;�tg��^��F���  ��  ���  3Ƀ��8�<�sP���$��)8F����f- �P���$��)8��;��  r��> u�a�`���  ��  �����  ���   t4�+�>�t�>�u�F:��  u� ȃ��+ƉF����FI�� w��(�� B�>�t�>�u�F�+F������FI�� w�a�`���  ���  v<���   �t/��  ���6�t ��V�8 tj j���  ��^����u�aÍD$`���F��<�u��5   �=   v5   �P�6�    ����v�6�   P�6��m  �D$a� `�\$$��[<�[xً{ �3�����3���2B�: u�;D$(tF;sr����щT$a� `��\  P��i  h�CwP�U�����j@h   h  j ��q  ���  h  ���  ���   t���  ����  �׋��  �@�8 u���  H�8\u�@���F@�> u����  ��i  �D$h �  j ���  ��u  a�U���03�@�}�E�E�E�Eظ   3ҹ6 �Ej�E��U��U��U�U���Y�u��U�6����E�I�Uu�u��M�U�����=   �<�s�U��M�������E��M�������9]�j  �   +�����M�i�   3҉7�uB�}����  �ÉM���   �M�+M�u��M��e܋u܋}���   =   �2���   �M�s�]��}�������E��}�	������9}s�ǿ   +�����M�҅��9��   �)}+ǋ���+υ��}ԉ�Ttg��   �s����a=   �M��<�s�u��M�6������E��M�������9us�ƾ   +����7��)u+Ƌ���+Ή�T��   |��u��M�E��}��U��1}	�e� �i����}�
}	�m��Z����m��Q���)]����+ʋU�+�=   ��M���   s�}��M�?������E��M�
������9}sC�ǿ   +�����}��M�M؋M�M�M�:�M�}�e� ��E�   �M���  ��  )}+ǋ���+�=   �
�M�U���0  s�U��M�������E��M�������9U��   �   +���ًM������}΁�   �<�s�M���U������E��M�������9Us=�u��º   +����3Ƀ}���U���L		�M�M�+M��E��
�M��2�����)U+���+ʉ��   )U+���+�=   �U��M􍔊`  s�}��M�?������E��M�
������9}s�ǿ   +�����M�:�z)}+ǋ���+�=   �
�M�U����  s�}��M�?������E��M�
������9}s�ǿ   +�����M�:�)}+ǋ���+ω
�U�M؉U؋U�U�U�U�M�3Ƀ}���I������M�M���  =   s�}��U�?������E��U�������9}s�ǿ   +�������e� �9�L1�^)}+ǋ���+�=   �s�}��U�?������E��U�Q������9}s+�ǿ   +�������y��1  �E�   �E�   �#)}����+�+ǉQ��  �E�   �E�   �U�3ۉU�C=   s�u��U�6������E��U��������9us�ƾ   +����4���)u+Ƌ���+։��\�M�u��M�3�B����M�+�ك}��]���  �E���}���jY�u�����  �E�   =   s�u��M�6������E��M��������9us�ƾ   +����4���)u+Ƌ���+Ή��T�M�u���@������   ������I�����M�}���+ʋU����
  �F��=   s�u��U�6������E��U���9Er)E��IuЋ]�È  ���E�   3�A�]��M�=   s�u��U�6������E��U��������9us�ƾ   +����4���)u�]�+Ƌ���+�}܉��L	�e��M�u�G�}�t.�]ЋM�C+�CM��u��}K�E�A�ۈU��7u�������}��ՋE���             �� �                     kernel32.dll � *� :� H� U�       LoadLibraryA  GetProcAddress  VirtualAlloc  VirtualFree  VirtualProtect               @                 `                         Ɇ  �      &���2��VWHc��#���zgݾ&�p�|.��_��t��،lIcx6�F��Uam�@�YN����c�k1���o��2<̤��b�rrh�WP"�	ZG���C����3���i�uS�Kt�@)k(�%]�
g	Y���ᕧ����%[� X��u�:Y_"��B_�����fL�F�I��sYAK(���z	�G�vԇ�	G�>�|�'�DS�)��ߗ�A_�leq�
Lm+겳F���_�=�el�|�fO6��MЩ���~���R�����p�TN��m��HDˎ>�8�B�6��i�;�-���p�h�p��P��Х��\���9��C��@��. <�$��m� �͊t��q����8@�\)�3��_.�M����B�3!3�����Z��WB�"�r൨u��=��fR���VLO�#SQ��ƥ����X��J�r��T�|tGr�h�_"��C�Yq�Gd��I��ͼ�O��9B�!&�G��s @����]X3"e�e���#��~�2(�M�A��q`�N$�RAT���V��0��gy�*�/mE���3���N�t�k �:�����DQ�pg�A�.��r�Q-�/�8� ~[�?'��v���No�QJ�DԠ?q�:�S�H_G7U���N�    �^X
�/��"^�Wt���C%�����Y���4�ڜ�l�%�u��R�4�N|���#���^��+'� �Y2�D�ϼC�2�$�� I8�ݺ6�����2� T�*�!Q���{T��sŜnm�?1ɹkr�
�M)C�F=m�}5����O]��W���_�lyhS1MqUH���:I���|W��``�	Ah�m�C$8n$���w���gŔ<��PW��z"���jX���� iP������q�N�Og(]��B�v��b�00"���T����C Ȯ?��D2��PU�.�;޳_��J>�s��t�>X:"՚��[��Q̈́�:�u��V�:t"�N�o���4���H�]�E?ص�jZI��%�)��~v�ao���ަ�����{�|k+��U���<@kU�w�C.��w��Lc7<�K�V`���$Z�`0  �E��E���E  PQh�d�Y�5  �$Zh8�ԩ^�~  �[3  Uh{�B �Q   �<$SQ��j ��  ��  �m  ��89  ��!  �	  ���  �	  �$��2�B h.�B �?  ��B  ÜhP�����B �$Á�?�v���  �:�E  ��[h�B ��  ���B � ��58  ��  �  ����E��@Qh�p����!  X�x  ��'(��F!  P�����B ���P�  �<$_�����  ��[��!  P�����B �����(  ��  �E��/  �E��}� �9A  �.  �������N�m���   h"��h�B �  Z����E ���|��$�@  �E�x��   ���N+  Y���-  �-  �D  ���L�hCC �   �?$  3���1  �O'  �E  �5  ��  �� E}���  ���1  ��  �Znr��2   h�C �)  �U�l�B �M  �E�P�&  �:  �����  ���y   Z��  �  hfmZ��o1�������$ZVh��s�$��[�Ɛ`]��  ���  �/  ���  �L	���  �3T�L  ��h94H Z��V=A�Ձ�i�vo��T1  ]���B 	���.  �  Ph�=>�X��
�J��  ��,$h��B �P  ��Z���B 	��"  ��2  ���t(  �E��E��B  ���B ��  �Y�E��@E��  �E�@����E��  ��   �D%  ���]�|�B 	���"  ��>  �&  ���`B  �	?  �E��8���   �4  �U�DC h��B ��  �)����@  �%  �q  ]#���  h�C �9B  �}� ��	  �EP�}���h��B �   ��]�5H�B ��
)  � B  ���A  ���w4  �4  ���"  �  X����n�Ł���l���!  d�    ZY[���  �D  d�5    d�%    �  �  �ǟׯ��~/  �	  �E�@������U��  ��  �  ��2%  �1  �  h��B �?  +��k+  ��
  ���SA  ������P�  �E��0  ����=  �E��8��e  �E�@��#  ���Y��`�a���M� �l  �E��E��8  �$   ���  �M-  �Ƈ4$^�E��
  �,$�,$h:#�5X���g-  �  �v>  ��U-  ��  �"3  Rh��cZ���2?�m  ���[  �������r  �$Z���B 	���   �U/  �E��a����  @�E��E�    �E��r@  ����`*��6   �1E��E���E���  ����0  ���F  É$Y��  �<t�<��������
  h��
ZhJ�B �?  �	���   j j j�h���  3��Q'  �0  hG?}�X�����W�$�~  ���B ��0  �{  �  �b�����P�c  �x��	   �E���+  �E��j  U����E��;  ]� ��1  �  �$���1����  �4$^]�5��B ��/  �'  �E� ��  �  ��  h8%�Z��H�g��C  P�  U�
(  hV�dX�����H�6� 	��>  �$[h$�K�$�=  ]�U�����V%  �E�E䍅�����E�h�B ������ E��E�E���   �4$^	��������  ����n�  ��  �$XZ�E��E��M��)  Ç$[�E���]��B���U��Q�=<�B  �3+  �����E���  �E��(  �:  �	���+  �)  h�B �;  ÈE��}� ��/  �E�   �E��/  �$�B �  ������%  �0�B �  �  �����  P�����B �;��$  �$Z�E��#  U��  �$�j  ���B ��@����n  �#  ��P��L  ����   ���hT�B ��;  ��]�5$�B ��F�������  h�~��X�v  ����[  ��	�(  ������  �1���  �E��E�h�B �N;  +���  ��   �E��W  U�E��  �I!  ��V���  �������h��B ��*  ��  � E��7=  ���U��E���'  ��.  �  ��  �;��R  ]���B 	���  ��+  ��   h��B ��$  ��m:  ���6  �⭺@�*  h�B �   �,$�,$��Q��]��B 	��8  ��Q��]h�_��X��$���}  �$�$�F  ���l  ��	a|��-  �X�K<�Lx	��]
  �L�9
  �@������X�K<�Lx	��  �E�@��  U�E��(  ;��6����$X�  P�=  R� ����$��]h�B �.  U����$  ����q*  � �<�<�B  �N%  �k'  �,  �x&  X��o����xLD	��J  ��}���   �K<�Lx	��)  �L	��  ��8  �)
  ��"  h`�pZ���^�R�6  �H�B � ,��  �}��   �E�H��  �  d�    �   �8��X� �������  �8��R  �h� I����_
  �?����t  ��  ���  ��   �����  ���B ���   Y1��1�d�    �B,  �*  �������:  U��Qh��B ��(  �E�E�@H����-  @�E��:  ���J��7��mN�́�>���  �����E  ���B ���B �s-  ���  �E�x��   �  �E�x��   �C#  ��  �A!  � h��B �  �]  ��  ������  �}�������E�H��`  ���,  ������E��   �  ���f  �}8  �  U�E�����Y�E��
&  h;�B �$  ��  P�,  ��,  h2F��$j �p   P��  Ý�  �E��8 ��*  �E��  ���I!  �8  ��"  h��B �5  #���9  R����������t  �$�B R�+  Y��8  �E���   U�E��l,  ���B �s+  ��	  ���+��+  ������v  Y���U	B��8  �}���  ��r�O)�j  Ã�<� E���  3��E���  �E�x��	   �E���*  �E���  �E� �   �  ����  �U���I  R���  ��B ���PW�������  �8�����	  3��$ZRh�}��
  U����E��E��  hb�ء_�R  �������P�T"���  �$Y�=@C  �,&  �U�h��B �:���Q��]���B 	���)  �  j ��Rj ��  �4$^��h�C �%  ����E��E��E��E��  ���  h��B �  ���}  ���  �   ������E�h���B�#  �$T$hB�B �.  X��;=,�Ł��ڴ�6  �$X����$� �<���� 	���  �
����5$�B ��������B 	��T����o���+���  1E��E��G���h��B ��	  ��  �S<���   	��7  �������$����X� ������������o  SQd�0   �@�����$[������   ]���B 	��������)  �����  ��  �F  �D����E�E�� �E��E��E���  �C  �������U��E�3��5  �$Z]� ������  U�w���PRhP��Z��j�9ׁʯ����  ������
  �8����<$_3��E��E��l   �l����E���  U�E������Y�E��  ���Q  �w���Y�E��E�������$�p  �$X���$T$��&  �E��}� �(  ������  �M   ���S�����5�́ó^:?�$�:���P������E��}� �I  ������  QYhI��X��^@:����'  YY]����$  �/  ��'  � ��������#��u�u�uh�B ���������t%  Ë��   �t����   +E�E��3  �}�f��%  �   h�C �@  VhS
�^��&�8\�4$�  ����]�  	�h��B �����$Z��<�B �E��}� �N2  �	  �$R��e�O  1$P���s���RP�E��$�  �h��.��,$��Q�A  �$Y�M  �`�B �E��  �E�3��E��  �E���  �������$X]��  �Eh��B ������Lx	��`  �L	��T  ��"  �I  ��"  �$[�	   Y�E��k  U������4$^��  ������P�g  �<$_�  �E�   h�����~"  ;���  �E������  $T$��� �   	������C�������3z����E������;E�h��B �  �p�uShbڇ4$�	  3�R�#  ��� �  �B���  �}�hw�B ��  �$[�}��!  �E�H��K   �%����g  � l�E��E��  �E��3  �E������E��M��%  �<$_�T�B �
  �����e    ��
  �Wl        ��  �ʚ    �H�����3  Pj �C3  X�  h=�B �2  ������$�  �U�Phu��,�B �
  	��   �3T��	a|�  ��  �/  3��ښ4hQ�2  ��  �G����8��B  �E��8��6  �
  ���  �q  �<$_E����t  �E��!  �h   E�3��E���0E��(����U�l�B �����E���  ��   �������Q�����$z�Gh�C �)	  P�����B ��W  ��P��  �8 �7  �E���E��E��������2#  �	
  �$[��]��B 	��R"  �0  �/  ������P���  �}� ��#  �E���<� E����  P�����B ��  ��  �q  �$Y�E��E��  �E��E�%�   ��<�B �E�������   ���f=���j����E�h�(=X���+���Tx^���8����  P�E�x��   ���D  �?  �g  ����������h@�B �M  ]� �B 	��  �(  ���B ��������  U��Q�  RP�E���r���������$Z� l�E��E�h��B �+  �E��E������  U���������>!  X��`����DIg�Ł�YPv� �������(�������.  �  �<$_�/���;E�������E�������T�B �  �=`�B  � ����������  �윉$��]h]s��X��G|{"�����f=���  ��	  h1�B �l�����W����  �"  ������1�������؁�PpB�<  �6�B��
  P����U�l   �4$^�E��������l���������P������U��h��B �  �<�B �  U��Q��  �E�Pj(�E�P�   h��n������É<$_�E�� d�E�h��B ��  �U  �EPh��B �q  ������������  �$Z���ˑOhg�B �������o���Sh�b[��O�<�$�E  ÁоT[y�$Y�@$E�����������$��X�E�   �E���   ��������  �#  U��Q��]�  �S���#�������ߐm>����Z>�;��C  ;E��  �E��@dE�;E��  � �V���	��   ����   � �Q���1������hT�B �  h����+�������	  Q�ȇ$�����B ËU�B��Z  �.���ÉE�������E��f���U�E�����������$�
  �������  U����E��� ���Ph��3+�,$��3+j(�E�R�$�������  �,  Yh��B �K���������k  ��A�ղ�$�E�P�  Vh�x��^��`��^�E��E��  ��$V�$hS�5+���  �$[�E��x< ������  ��������#��|�
�  �$X�E��t  U���j����P  ��
�4$^�<$���$����)  �E��@<�$T$�����E�8 ��  �E��  ��f}2������Iw݁�Z#���  ��  ���c������  �������  �e����$[�E�@����E�}��!�����   ��  h��B �1   ��Rh.X[�$�ѧ�P��B �  ��0  ������������  ��:  �d	  �〙HdZ��������*  ��  3�Sh�Λ�[��y�#�ö0�$�N  h+�B �h���P�}����Y  ��������	  ������P��  �E�������������U�����  ��<� E����E��E��!  �  ���G  �:���P�E������$T$��� �����������  �$X�   �E��E�������E��.  ������2�����  h˲9����(���������ӷ��<��|��R�Շ$V������]ËE�� E��  �E���h��B �a�����������.  ��  ]��  �}�������E�@������*  ���������U����  ���T�B �  �=`�B  ��  ��I  �E������E���  U�E��C���Y�q  ��^���������$�_���h��B ����P�8  �4$^�E�S��  �,$��Q������(  ��)  �z����U��Q��]h�fC��  ��  �+'  ���E��E��8PE  ��  �I  � E���;$�B ��$  �E���  R�$[�$h]�0���  �<$_��P��h      �)  ��  ��  Ã��8���0�  � 	�������x  ����������B ���B � ���  �g����-����{    ��  �/=    �d  ��    �T	  ���    �  @�����Vl3#.2� �/  �%  h�l�@������$  �     ��/�����x  �   ���P  �C  Y���U	B��(  hk�B �����E�@� ��������v#���  ����~�������[�����1E��E���������E��!'  �������
  �����U��Q��$�  ��!  ��������׆�K��&  �=  �׀���
hq�Ӿ����������   �;   �  ������$[�U�����  RhN�B �m  E�����h��B ������݂���E�3�RP������E��E��e��A����Y  3��E��   +�3��E����M��d"  �6����E��}� ��  h��B �V���ËE�8 ������������.  ^�1  �6����  �E�   �E�h��B �:&  Ł�$t�<��  �	��������������`�B �E��`  ���h�B �z��������E��}� �K  h��B �
  �L�	��2  �   ������L��4����j����$Z�$�|  h	�B ��  h��걺��B �$�������O�Κ�W  P��������8���+��#  �E�3�RP�����E��8  �E��X  �x��   �   �E�x��   �B  �G  hK�B ��  ��	  �E�   �    �  �  ÉE�PhP�B �!  ���&����E�3��E�}� ��  �  ����3��  +��  �}�h��B �Q  �$��  �@�������E��E�Y� %  #�������������i  �����k  SQ�U����d$1��M����@���E�}� �
���������e  ���  h��B �  �������  �����U���#  �������������)���;��M���h��B �����E�}� ��  �E�h��B �w  ������E��E��  �,  ������4$^�H�B �*<��9����  Y����   ��������  PWh�b5�_��`�y���������nFO�S  ���yi������$����  ��)�����a  �n  ������$[� �,$�ͽ��B �,$�[����4$^��)4`K�_�����3D=	a|�f1ہ�   ��������h9�B ������E������E�����U��Q��   P�B�B ��  �9  ������RU� E��E�E��%����}����$X��B �  ����$�f   ��U��P�	  h��B �^���������������s  ����/����3�h�B ����h��B �K�������������Y]���  ������������;�����hB�B �v  ��F��������.�������  �}� �  �E�3��������=  ���`X���������C�	�$Y��fj^�<$��  �f����TC �@C ��  U����=@C  �  �1�a����������/�������w����L�����������������$[h����hy�B ��  �"���h �B �������l  ������m  h4�B �����#���������h��B �����;����}�f�  h��B �*  �$[��h��B �e���X�����U����w�@� 	����������Sh�[��[��H?��3�/���B8��$�h���hvF�D�����Qh3yfZY�髒�/������[  ����  ��  �}  ��\  �4$^�������]1�������   �$�B ����������   �0�B �����U�l  �U��E�3��E�}� ������E���<��  �$��[���h6�#Չ$�@
  ht.rX��fpŁ����������   �  ���B �k  ��YCA�$�����윉$����B �,$��  �=������B �>���j��U  Wh=�B ������  ������Znr��4���P��
�|�B �  U�)���Ph����4$���j �Q  Zh�&���$�  �E�@�8h��B ����0�	��   �W���	��t��������������=  �  ��  �$ZU���  ��   �E�@$h��B �u  �K��������$YP�_����`�B �E�3����������h��I�Z��Vz�����U����$�$Z0��S���������>���P��� ����  �<$_�E��E��������,$���B�E�Ph��sX���ap�����������������]��E��M��b���� ���f%�8f=� �n  �����$  �<$_�s  � ����E�@�8h'�B �'  ��	  ��;��m+���  �����������  �&��������E�h{C �_���P������U��Q�W  �  ��m����1����!  �����X  [��P�����P�r  ��C���WhS�B ������4$�����������  ���������ݺ������Y�����3�;��|  ���  ��je�������<�B � �H�B 3��<�B �  ���·$X�E��  U�E������E�@ E�3�RP�E������E��E��@`E��  �����E���  �E���  �$X�E�� �����}���  Y���D�w�$��������������]:Ɖ�1���h��B �������  �E��E��M��g�������������6  ]�����h$�B �������  ���<$_� ������8 �����E��E��e��;����E�8 ������ ����������������  ������D���Rh�8Z����&�������9  �������������������J����DC �����E�P�S���ËE�Y]� �v���ú��1��1���P�����B �����h Y�������������  ���9  �u�u�u�ЉE����B h��B �*�����^���������O����E�h��B ��	  ���  ��  É�Y[��7����r����j  h�B ��  ��������j������   �U��Q������hNe����  ������������E�P�3����TC �@C �E�3��r����  �$Z�E��E�YY]�%  �}� �k����Eh��B �  ��
����J  ��]hL�B ��  �$Zhp��[���I��Ìow���c��������  +���      �����2�    ����n        �  �z�    �A  ��&���h��Z�ʗ�߁��F��������������=��B  �/��������������e����.  ����]�h1�B �}  ���������������Ł�Z�΋ ������$Á���<��sۚ=��	  ��<$_��]�������8�������U��Q��������_���������  �  ��P�U�#	  ����c�$[�E�����$[�U���U���E�������  �I������~����K<�����V�F��������������h@�B �D	  �}� ������EP�}����������ho�B �����j j �y   P����X�������M�
�1���Z���[	u���¬����1������  ����"�$������4$^]��T�������������E��8 �i  ����������P�  �������P  �u  ������E����U��E��&���É$X�E��8��  h�C ��������������h��B �����E�h��B �����=<�B  �  hr�B �O  �<$_�@`h��B ����������E�PPhJ�B ������U��E��}� ������E��E���������U��l������  �	  �  ��E�#������U�R���@U�B��E������E��`$����E�P�Y����0�                    ��  �n    �����<C �
�����Y͢�u���h�B �7�����d����E�������  Q�L$�  h��B �U����4����}�p�/��`	  �E��S	  �������������W�$������T$���E��^���U�������}� ������  �E��E��<�B �E��}� �������  Vh�&R^��8��4$��  �������[  h T_������U�B 3�RP��  ��D����}���XPSh�@�[[� ����$Z�8 ���������hSC ����������Eh(�B ��  �Uhr�B �$  h��B �7����������  �K  �������?��$X��E��E����������B �����������h��B ��������F  ��
��������R�+h&�	����������a����B��E��Eh	�B ��  ��]h~���X��I�&��ȴf�,��+�H�� �   @� E���;0�B ��  �k���������0���	������f���Ü�����Ç$Y�E��8�������E��8����������P�E�@�������P���������U�������y���	�����Qh'�Y�������<$_	�������  ��3���E�3�Rh��B �W�����9������(�����҇$�������������Y���&���e����������0  ���������������������  ����  �  �   �<�B � �H�B 3��-����(��  ËE���
E��E�����  ����������h��B �  #��9�����  h��m�X��� M��VD~��   �	������7�<$_�@��?����G  �E�   �V  U����������
P��  ��+��������������}� �\�����  �y�����#��Q��������4$^�E�}� �{����E������\�����#  �����hK�/^�"ȁ�c�O��4$�E���Zh   �E�������������E��E��E��E�@����  �����I����u�����  1�������U��A������  ������  �x���������U�j����E�E�E�������TC �E��E���]��x�������������h�C �  [�E�f�8MZ��  ����J    �  ���������\    �.����p  �\���f�`P�� hT�  j �P���N����E�� ����  �e��������P��������H����r�������7����h5N_\Z����hE�B ������$XU��Q���f���������"����E��	���������������  ������hR�B � ����,$�,$��Q��]����ËE���$T$��� ���Y���f�8�.�   �0���������E��   �������$ZWh5\q�����������������  �=H�B  �t���������!�������}���ËE�x��	   �E�����������������N���  �?  �   +E��E������U����� P�����,   �E�Ph��B �������Q��4$��^���B 	��"���X1�V�&��������;������h$r��Z�Vq�$�s�����;E�������E�@$E�3�RP�����
����$[��f������E�������_����b����,$Ë��B h��B ������� ���U�R����E������;E�������E�@$E�3�����������E�H������}�g�C�������������]ËE�� �E��E�$�-  Z�§�Z������@  �������P��  YY]�3��"������=  �� �������y���d�5    d�%    � h��B �=��������"���������$[���]�|�B 	��/  �P�����������������P��
���B ��}�����
�����X��;��K�����>߇$�  h��B �-������v!r� ������]��Y����0���������}�{J#��7��������E��E��E��Eh-�B �"����E��E�YY]��=����4$^	���������������h��B �2���锱���Q���U��������̍�B � ��M������E��   ���R����E�����1������U�윉$������O������m����������������l-s���G��j����   �E��]������U�G����������IF%������H�B �J����=H�B  ������  �%   �<�������Y�E�������E�@������������������d�O���P�'����J����<C �������Y͢�����7���� ���N    �i���
Bb    �������            �   @                     �   @                     �   @                     �   @                     �   @                      �   @                      �   @                     �   @                                                                                                                                      @   B   �   �                                                               �   B   �   �                                                                     `                                          �   @                     �   �   �   �   �   �   �   �   @   @   @   @   @   @   @   @   �  �               �   B   �               �                     �   �                                             �   �   �   �       
  `                                                                                                                                                                                                                                                                                                                                                                                                        �   �   �                                                                                                                                   �                       �                                         �                                                                                                                                                                                                                      �A2�2��6 ������    �����,����E�� �U�B��E������������4����������a���Ä������YY�����7���h%?*�Z��vhށ�	܁�#����F  W�$X�E��E��  ����T~�����������P�,$���)����$[�V����H�B ����������E�H��E�� �U�C���#������$Z� ������p�/�����������x��c����E�x��V����������3��������������$h�B �m����E�E�@H��������'�������6�����R\k(�<$����������P��
�|�B ������Q��������x|�	��������������U�h��B ��������$Y�{������ E�������>���P��ShHl�3[��d�k̉�����$[	��������������������������+�������������B����A����K����}��)����E����H  �)����_��������������������魽�������@�����B���[�-���+E�E�E�� �E��=����E������ڌ���K���� �<�<�B  �����E�����+E؉E܋E܋��-���� ÉE�j�E�P�=��������;��K���3�������$X�r���Y������������������������E�}� �*����T���������������U��[����$�$������Z�������4$^�4$����������E�� $�<��A����E�f� ����� 3��u��U�E��]�U����$Y�E��E��a�������1������1�������$Z��<�B �E��a����E�    h��B �����������������w����4$^3��E��E�Y�������������������s���	�������X����H����L�	��s���������蜽���IF%��v���������V����Q����������ÁƛnVh*�B �����U���E��E�8.�����[���������$Z�U��E��D�����{���Y����������E��  ��������/����������ٸ�  V����������ha��w��iH}&V������\ū�����{��������+��� ���PhP�B �����Pj �   X�8 �������������������U��Q��������B �8���        �C �C             vC     ��d�[����2�|�\��
ʟ��{�׏�F�Y�٦^;m^?��t�.7n�[y�ڽ���/�
8�CG���y^�{_����We�W���IҢ�e�}U+�����aͪ�1--�fx�3Hl��o��GuRH���œV6�����Nkb��3(��65v5�ҜV;v��to�%���$RX�����N'I�j�5QH�&]?����ρ��F�QW�����Z��a�Le�2.5\�`W����� �sѭ�Y^�l�*L�I��H���"�2��?���"�g���ʴy6
��N{��V��<R���ѽ�ן��H�5��S�.s@\ҜmP(����y��Uf�������c��P�Ǜ���_�F��K�^F�]��-���o�A����Y���_Hr�=���������@���Ǥˑ�m�ɮ�0Q! Z�]����лG�7�n�}�䦬�+T����o�g}j:3��c�Ц��)1A�n0Dkn_֜I�Q ,c'��8q�B�!�ߡǊ���`��yh�u�Q�W�4?A�1˓4��ck���Gc i�i^ϗ�>�|�]|*����q��C�s�D΁�y���,)э�