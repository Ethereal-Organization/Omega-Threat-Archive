MZ�       ��  �       @                                   �   � �	�!�L�!This program cannot be run in DOS mode.
$       M��'	��t	��t	��t��t��t	��t��t	��tz��t���t ��t��t��t��t��t��t��tRich	��t        PE  L �HE        � 
 `      �   �   �      @                      0                                      p P                           �                                                                                    UPX0     �                        �  `UPX1     `   �   T                 @  `UPX2              X              @  @                                                                                                                                                                                                                                                                                                                                                                                                                   2.02 UPX!	�< �=���  �Q   �  & Sv [`P�WSP��}�} ��ȜXR�Z~ [_Xn���A ~ �өV��P����X���w��S�OK3v��&a��[��8>¸�MgƁ��ǁ�;&ƹ �w�����Ń�i���	!7�� C���N���n.�C�q�΄��m0(��	�*N�L=�~n&�����}U�o�J����I�׿�0ԧ�O�G �����XR�\��?^_���s�ښ��HY����C`Y�О{y��N�Q��]�l?Z(v�{����dFU[�Si�Z�Ԓ����@���1�`|�����qbɥi�+q�6��"A�zhH3�~�7i$�w-�<��D4lE�Ca� �����[�(��4����� Ue#����G���,����\g^��A�	���D��&(�0ƽYt�����]]E������a'�@`�I��<>���:�J�/�=0+���\Y�[e��\MK��.Dt�<�'%�s(s��pC^�uJ�㰽n;��)��,��"�����Z5��i��a�UG��QՂHD$_D�?u���\�ș�b�y8�
�q�����p4V�d+�k2�-�xy�jw�x���m��F���=d=��x��������h
M��z���+8y�si�ȑ����WC��� D�n(��ts�t��[_m�B4J?Fq��	�֋����S���I4ܦ��\�4��'�i 9�t��D�Dr��-x�0�԰hИυ��!l�����#�ŕԠ���o���+��ɹ��k�&�ՙgX*)K�H���N�����H�]�����^1TUM��u�K�Y��R�<��q$tw#]r��S���&��)�0'�������)�u�+��(C��!��7�\�0��N�U�IL��pwt/i�oi�k�e�Β;.ĺ������͍�zep�bԀ=��Y09�	�	�,��b�}r?����j��7[W�Fæ5�%ѝD�Cq�D$�2P~ -ɮ��
	���Pn�	-�$�>8�	/ٚ���?���`Z��XY���h}��O
c�<�i
�E��F������e�=O�
ܦ"�s�2o5I^��*t#H&e�G���yyD�d�>r������DGA��W�|vhl���Aa1�Q�Zv�����,���?��e�S�q���trKWQ1w�z�*t@��DJ:ڪ����ԍd�:�+�l�7ͶG���]܀��^��Y$�m��ܻ�����ц��8�;QH�1�r�x�ɨ�Yۜ˽�ػ �/[����v:��)�|�_Q׏��.C%�&#��[ؙ�█c#I�~��R�MxGs/�PH�
�#�%�w?�)�c*�א�
�)^N�-�y*}�pE�<�S��8τRDaU��!�0�FlbLT�1�6��%�N������%U�'X,e�DÙ��8�%�27L���x��"� �'e$L.��SV�$X���j@j�\�~�=nW<�F�����5�l�×��N��k����y�>u��7�$#��jo�����ή�#�ܺ�>���;DK/��W��8�S�Q�%1V���l*��r��������t��>�Ɋ�a��Hu�o�j�ڃ:`��ג�����th/z�u ̌��Ұ����"��-��������J�56s�9��y�K�>��L�\� ��� H�m�ES�1x�z�1��-ȏ�J$�*��G�V�A"
�ri�AX�b��͓j�F7,鹩�Æ&O�4^��ҍ��*r,5y9��w�]��_�.�?u�P�&�(U"��;�+�K��Z,�T��F�=9@�/@���d5����B*s�7���T�]*��SVY���:�1_�_��e^�c+�	��{�=�'� ̸��ٲ��ү@�����{��L/�Ѩa|uU�V{�62/�R�4tL��v�6k�a0��~�aS�$h?��4��fs]Q������tmq�}˳&E�1��9�A���Qov�lNg~_���f��f\1z ��'�8��Z������n.$
�&��遈��f6;RoR��x��=|�@�$t	 �R�JK��a�q3q����]���k�XVm՗ޡ�$^�]��yT�v\E�C�!Ε>E�^��Rt���KIbv)iX� &�&�7bڢ��goq�Q��s�
>���\��|ݙ[g�$� N�v�}�q���P�!<����� ���v��}�� �1\���F�
\m�F��D���ހ�xWhL������3��	� ��� 	\r*F\���ی�΂�RÀ���#�R�kП��!��۽z�`�c�D�v�$]�Q#D�Y��|4���&!W�ꯍ51���OH{Wr��i�,TU�������b�%*A���f���	L�>:X���J�����<��Zʢ�"$k��b8�ͷi��X���+�Q�$:���pC�>p$H��w.P���@�9m�m.�V�d `�A"ρ�N�+��,Mt�:�'���=��3_�m΅إ`���='Z4|�	o��ۯg��2.���Z������7�9iw���{�)����W��RL��I�+����'�2�U˿�1�H�\Ex�;����i�'D����O���>l���~0����]B� ����Z�F�}e�^�I��� �#q��Q�/Ƒv�)y=Sz/��r$܏+��Y��6_44�OkC��J��j~m"�H'L_�Y��UU��'#�x��u��F�C1�D}Ͼ�Gi$qVJT��3����w��#tn�d[���n#�V�����-� %�B�_�Z�5ٴ;}ո�/���g�떏u)5�j6;�AȊ�p�˝�8�5z'�؅v�{2�C^�#m��׫��&;  F�N��7����L�g]�u@fcה���u��H��W�N�BA	�΋P.�%wA|Su)���fW�O���gA��l���5
Cm����3%5I���~�v��
��W�K��u�
��D��vR�FvnRPvbR��˃����0�	=2��;�EhHvC��"*Q���y(��mAp�hx0��k[>	Ty��y\��	H�-�\�����?Y	i�NJ����q�����,$K�18^�B�ZW6����d_G/�Q�S���o����,N��_�e�K{�f=-���貔�horb��%�K��Q��'/��G���r�~7u;�B�j������Ӂ�4ʑ�5/�彝S*\1-t�	M䆱���&���1$W�.� 0��Y�����͑|�KK&�V0��#0J��ku�9����Y+�S}�I���	�U ޲�����%Cv� ���.�{#{�@u�oG�xh	w���(n|*�e�$`h���=zn��*��E5CWt����b�0���x�!�p=Q�W�o��.��?���-�DG�(��MI�?��}�O ا���E�.��h vÅb/yM5��^i����F�7J�x�fN'�T.�"[��D�/��<�.3���7Ͱ�_�J.BSXo��i�5!��w�mi<��)��.��R� �~�ߴy�y=Xۙ��šo�����B��|T3�4�ە_r�7� �o���k5Q�{s���q�����0��<TD,���5!�o�9��z�U���! 9�"�ۥz@��D���B�~�BeF���ߝ�j��2���_��_择ѳb��B��*G*
sY��PD�{=��a�Z�� �4���ų2�}/�q-!}���z�	CH=I�X��
Ȗ|x��+EJ��lɞ7E�1DK��ع��ZKQևO�c��9iV̢��lǅ�y�
�>��>JϽ��t[�R�w,DB=7�2u��e5�Z^�j�D�ƚ�=�Lqj�'!�u�9\�[.R�S]'� ��%�3����@�{78��):���N5;��&�������W��Yx�p�7�L����(�˃n��s����h��B��(0�Z��Q.a<��dDLՀ=���R�c��i�~�����[eRd�u������s��n�:� �s�el�|�&D>�G���9ҥ�D�
fƿږ%ݑ;��/��:]�T玙�!H�Х��F�0Vn�����X_�x���>�`S�Nw�.��&�_��ډ v����7$lŤR ��mp;O�8�e�DL�g����P �w��~���J��E�t����F�o*�[�'�Fw	U`�!�Av�&a��S	(���d�҃�6!�yS��-���Ch���������)�3p(�i�o���UPBt+���,��&L��實�5���.mbb��yc��l��RS%��to/�<,j"��X F�ߘ���d��>��e0d���0��&����
�0��0�����^1
w\�~���k5��I��'*�"˖�w~r�)2�7�Z�T�xW��J���u�o�����Ɲ�Q]$F�!y��i$e�ׄ,`d$�5i��N
c��S-_�!_���!��h_��ԣx�
���|P�^�&����`ۓl�#׎�/���QGݥ��B"ďb����׿ʠ���+Ӛ?�%3�� 4eo��=I��)w5@rz��:|��?��N�&�H'e+gYn��I�'i	�)�a��_���8��!̶�BT�I�v{��x��Ʋ�4�8o�e��*�\�ó�4�jB��U��u�(8�p9v�)=d1��G�8���B�2�L�j|Wq��̵ ��-{Z��6ҹ�����x�)�E��.ԕ��w��,M�&���j��㱃���P���g0D��>r��R����ҿn?te�����
L͍4��.�>�L?�.���k�7��9�qԿ蓩5�<a{�ר܄�l�n"�Ι����:�r;Q�Ň��n9H��8��hx��<@�z	���Y��Pʔ4���� ��z5�oP�ptj���8����R������A{b���'�_ј��t_}C0жm+�H�|<��UNVn�h�<�;��BOwRp*6��@�U�s�v��T� c�1#�3���<�*�
^b������{�`��p)tQK0С.Q1��9`$�,�]�n�_UI�NO<S���1��&b�d{�қ8�TO��Nn[E��uO�G+�9�:��MJ��{�	�Jw=Jr�Y�1&I�m ��]����*�d%�?fH��JXe]�}��L5HA�3�س���yd����˦�7g���<k�s3/g-�y�Ċ��CZKe��#����4���<Pt<�1���{q5�Ĳ�(��x�~���I����8>�s%�/���J�'*7F�۝̀5?�@�yO}�ط X��&��zl�\�]Q���3���m oS'��@y�C���l /��>�_�{i���k�A>aZ��=��>���j�8n0rQ�]Z�C K���ڔ�KD5$u��*�p��;���)�¾�����%[
���M�Y�&Զx���W͈�[M�}})�-�_�M!cmB�&y.�����=�N7��ey�p�k!d�R���`�r\���������n�3�!W���#}x��.n��\��J�8�}��ˍ�BJ]�k*�<�A������4Niʌx�"���U=#�BߩOl\x�
S�<\G$�J��X��*b֯\�>��B�;���Eq_��eb����?o$�#ک\��{r�H\��T�d�N����F��H�lЕ��[f~.p7lR�Ŵd����,/�����}���\(����p��AK� 
AVhm7��0����f����t�Nb��'!i��o�&�h@�����/�]��|H�6ڿ��5�i� ����j.�#_��V���-\����"7�:��!������[����Ìm���j�����L�"�n%��oONH���`��L�=<�UQ�a2zy-N������q�.Ǫ��;�0K.Q>T�i0������8�6�Уs$��I��@<s@�M�HbI�٥��SJ8V���ͭl�O��U`Q��,h`�;�;�$�@|�@����bX�x
6&�J͆�F�.�L�b���i��t�����1[�
>�$�L�$��n��v�פs#C���6c�Ӡ�	��x}�ܐ�&bq2.SBo��^��3��VQ��
�/˷��q#p��p�Wb�F���UI��i�F;.a:ؘ_��S���KɄ%��Y��O����&I�Yg�U��8"�� �!*\�C�Y)��!X���NL��&M���e��c�U�wӍ��:�:~Vބ-gL��,�dCl��X.R*[��J^^�j�1�I.������厬��?"6�Շ+���N���������a�P7�� ~���a� ��>��X7��Á�.�t(g�ƻ$��>�J�\gl�?L�K�D�4�Np��,���1�׷D�km2Յ
�F���
(;n�k��s�s�
�up#<�ɔ�K��=�i�?h@l�1ר�TT�Q6��C��{k�8����]Z2V�v�����=V�^W ��n�
Ѽ����������XC�4`=����n��3�:�LsKj�m;,Q;�l��:B��=N��e�6��R�v(_�1<	' �D�r�A�7 �k�X�~CV=�"�i��]}���Jȣ
���TqdD��<��CXM_��M9m��䡒��8�u��e�D�0?2�cg��Yg��꘤t���&k���4��[�NN*�5��ธ��z���d��X*����kq�b�H��_ɻ"�o;�6�YY��ޘ�
%	-�গ�-��W�s�Kt�b��X=�.b�>9Ș�[o�`ˑ��r�����ɞӷ�`E�[��s䉺��m�+-|6{0)��THi��H��ې�D ,����W":�D23|ߍ�\6
������-��D��I����T�ǡ_�@Q�Y��9��Ybܫ)�O��|�m��c9G�kt`5v���78����P/�/"���l˾�hřHT�'��7����'kG�E��s�f�QW\@ꋰ��Z���E'=:nEɃ��� G=e��-�Yd�\$E�Í��~`�d�)Sl�g��e�_j�"�뒳PU0S�"��bDF^ʳ�o0660֟Z�I5���U?�Ǻ��Ƨ��@���Pu_��4���^�\~?ƌ�-y��b�����}`�v"��R��Z�\�h�n�o�>ʨi�eUt�Цk�ҩպT�r��I�xM��C����'��������q�t1�su�3��Ha3��jgH�� ��q�n��w��r��R���.�}AZ-��7��B嬠)���1͸p*��:�7�&�s����@vK��B�&�;5���Y���������a�lbv�h�C���@�����$�����J�d�AZ�)`��v����z�Q� X^Y]E�&�e��-�;��T���e�&���m����>�T��*I�t2<X���=j9:O&�t���VX�Q^������1���Eǵ���k�P�Z���>��2�����Xt�\��i��x7�*��w��BPY��ڼdb��+d���j�C�����uOz�P���0ph�2��1c6�����X��:�ř��P���b�C�q�cu/M��S��_��r�����jL��ۻ ��̤�9S���V[H�o�7꥓w8	����˘��ĶؒI�PU�H��^k��ë9��n~k�Y�	��~Lj��ֻ+��6�*>����4z�ꨵ����9�xBhiz�T }��MVI��E���*�(�İ:P�ʍ��@�(����d��I��4��
�k<���0E�ʿ��y
]j9���܍Ʈ���Qtٸ>��[Qc�$���|;"��m��}���#�P�A	�@G�3b~b��R�w������ș��<��n.�Ow�-��3h��@��=>�XQ�?'��ՙ��Ws{����&���q�A5l_��a�5���L�IϏ���Bf[0���e/�h����Y���{|�@�)���X>��5m�s"Q�c�K/Q�erU��N�y2�U3R��p�#F�-oo%d�Ag�j��FY�pL�I@c��fmO�͛m���66r�c�=���wzؠ�%F�s�l&?]�D�w�JL���b%T��Vs��C���i���j�g��$���rN~J�埕� �۾^�5V�Ȳ؎��q{ڔ 9G��uo"�ء�jNX��~9�,���� �D�j�|�Uxm��mƁ��w�������#^2��{���0���U��,�����J5P}���Ek�	0Q�]&[5�̙�.�����̘�X�&1ݏи���N�;JM��@�j�B�Ȁ�P~��_3Q��<��I��x�`yc7Ǳ����� ����ȶk�u$�MZ���7c��.0=iZ׵�'�b�:�h\�7KNm`�<s$��2��qt�����v�m�?#X�����)��S��5`I��.��Y���g�2��
���4��:�����|�`[(@<���ŕ86p�,�CFE�ս�!ߒ����^�Nw�8 ��ǒԋ�qZ�uc��s픨�~2�h�m��QL����놭lk�疠��<�	�����#@'����E� �Lȇ'
␬D�^$]��Vݡ��4�K�e 6	W�.6]K�9�0{ה�ZP_�)��;�*�������m�(L�rJ�Cy��ɻ�����X��z����E.�2�~e�u��B�5���
�^�l��Fqv��'�+W�o�!RP��՘H�8�5����~v���x� G� ߳���F�@�pRW�PE�0���em���FMق6��詫�Y�q��v�˱h&⇭j��G�=C=e!���ؗ��]��#�ۡ]��Ȥ�{���°5���/,�_9@#Fm1C�Lr��V�X%s]�y(��nY��"�bէ
@p��!�sѰ��I��w?��#q����I.Ӷ`����{��Wd��-Ҩ���a���c{���y�T��js+jy`�2���uM�wn/*q�
��84[��߯&!�L�aƾ�� ���2{��j�Nd�U��C���A��w�Z:
��'��K��]�DG�!��Z>��0�;����"����G��˗1<SQ`1"������m~��b��WQ�93"c*���f�<��eAN���:|�{⌥�~�Cs0�v��^�1H95y�>��D���l\vO/�Ι�B�;�8���z7�W�?�E��-�y�{엺��hD���|AIH-�8�����(ɛT'�g۹�P�9j��`�MbV@Bd��?>����<o�/T��֦.Oa��mX��� �A���˂o��a���G`ѡ�v�m�\��[�83�^�rП�d#�g4�v/Ӽ-*3�._�S����s�b��CbI20�>�n���~(�b�����?K��_S�k��
�����uB]2��i� �c�v2P܎~<޹��)�|�G�4Z�7�e��e�Px�#�Hޓ�sJ�l�^$5�O�uj̥���̈́۴L3y�b�:�+�"����FY��S���,:�[F�d�U֭\��^��\J�1*�s���"�!�=]�$\�F3��ς�oYC�Ti��,]��0�0�i�!-}b���2%FBReP��/���u��X���o��3���+y���9Vפ��	�O�-֡�{h빲w�ϩ^�H�n�)�����|�~�1�*�0���Yoj��}䃎�
���~��:s�:�"�uئ���s{������˵��2��O��b�A��~��Q.�,Ԗ;����͗������4�Vp17�h���ox�������2���!0߇Uv�f�V���*q�$���E���I
�*�t�g��7�p|h��1�S����(J-p��]��O~\�J�%(�|x���V{��U�ܯц;�{�X ��f>���N~i�<cFZ�H}/��/,x~������^��O#:>���a�g��^AY�����a�������,�=I�Jy+A�h�w��δT1y"E
 �c�����4����Hy�f�H�_���mV3�a�8�R�5��g�TTK@�2�gw�1���`�Lg&v|F�\˘�X���姞|���A2�=#�F)	&����[WpR0��9ìn���%�w�|��S��h��;R\lg�<�E}�g�y�{��9�׉��Y���G���[	^o��Z Y���ؠ,��
�09�;��3����~�:�O�� �7v��Vy���n�K ���׀L�T�/xr�z��
e�	��ۍ�<�jC����Gէ!��'��?������(��S��Ҙm�1M�l��?w�5���/[TwG%�m�Ǟ�?��i��g�t<�¯�b`4���`}�x�gJ�d���	t�f�v�Y�t(R~��w�@�|7�N�����ݮ����q9�~�xW���w1/���f/^��%'H�?a�X=����*���#�>�� � <Xɖ#J��afKe���!�&��fK�r%�Vz%v�P�SE1�w�Q�]cE7��6�))a7���xD{��-�����Ax�sv���'�Oj!�e�aW4�1:3;�!�6�|��t�}(�8c�G=����2��W����c��N�Ǩe6
2"�-9����H��Ǚqh��E��2�D�_�)'( �	3`�U\y%m_�lr�gN~�f��&�nxUN߸���$5�[��_�|������9�bx��8Յ���2S�uEAV��%�œm��@zFX&�Zi���=>�_W�������N�1<Ư�Ł��M8-{Gd�W�㗟�Ҷ-r��4�M��W{�,|RC ���A���$,��'��,��֎yM��E�wC*��@��-�¢���c=`9����r4����7�p� *h#�k�AA3e*�5�u$�,
�|���qÏN�ζ{8w~��F�,w�RSk�
z	�Ho�.�ĸO',���(�&9Nm�K��+8���x!��J���^h�RE��eeg�Z�h��|���4���d����U=���.P�M��sZ�bd($��/*�,`"��(���8�tm��y�.g�ׂ�}�/s�d��h��6�gq�6��fr�f��y���-��!By�3l�	1"{b"ɋrg�a�-z������#��١�����\P�<G����«� 6�=�J
{�dB�e>�s�_�H���4��{E��a����
H|�a��(��2���Vh���E��	����'�UO�,/=���5�3�?���b�*v����<�h��UN�e���]"���3�	wy~J�m}a��?�AQi� ��%A�;Np���vS�tdw����7��𖍚���\�����������
A��8=a�&�p��=��g����@�<9����  o�ޛ�R�j��iP���tupB��XL�������ߎ�h�����o�j�>�y�	s���bRB��T���ߞuP�]�?�y��������i���Z�Z��2�,� ����&�m����Tqo'�a��a7ln?�Ծ���������tcG$U֧HXw2�$Ҹ�G���m4�N��M�q��2�G�VN�ۖ4�:�0��1~aɯ����u�W[x*z+"̓Mw�wQm7"��ĆO������6͂;F�x��kk��V��M>K���:P�r���{e$�_��v#o��X� �a:��$�pR����E�dF���Y&vVm�"p�]��	5����%d��9E��S�UޛN��>�us5��\.Pͬ+(G��#�������!�S�.���zbAŨT��]F�ɶ�4�'\�����P<��0�S�'�ee����v��^�k.�ݍs�̏t�6�5lQ\2�����i���#�T�"��C�0�5��h*(�τU6�;�&�c��SD	�n�	&�Q��I\��"�NuO� /~�\g����S	3�란>)���k����lǮ���׵�m�b}ig(Y���a}�ߪv&��DI����`�J��T�%�,U]�z4i��q6-�U�	r�>���L�,�:{k�g�C6�V�v ��$P7Lj3�;���U��ѡ�.ѓW��S8a�´f�T���kk"�/�ˎ /��v|�[ҷ��^��E�t�ǀ�
p�.�%!X�d���c�]�W\�� h
QAA]����=�N�G;*�d�#Ѻ��y�ٟ%/��*��B��}Y:h�S�2z��ϙ7A�1���rB.E�P�}pH�$s���x+P�][Bh�A��J�`�C�W`��
��aە�g�Xu8�H���?�g���I���,^���3�����Qcη�̿j��1H��[;�#.T��ԕq�����������/�h�@��p��c��eQ�����i�,n`7.�O_~�D�B������v��ۑ��	��fv'�5^�l/$��d$(o����j���Օ��/ɺ
^%��>(e��N"�i􄋽��L_��$�]�f::Q{�9�Դ#�N�Q�������N9��bR�� ���5��8Z2$���wN5��%
{�k���b�Mr7V�CN|p6B|���9_5��$��i{r
ȗ�G�W�� K��)%���K�a,r����S3�BX�U!b�� �$�X�0�W��wA��9����Q���70�2}�	�%����2_�u'�-C׋!'��y%�0i�C�=Zy#������0@G{1�ȼ�p��*��_m]H��&�MŲ0�7*�Lk�E��:��#��3�+���	1H��x���6D-���U�B�'�#!�,��.�ߣ�I�.`�ih���+���;4W��[ݭ���V��̨��'�O�&��i"�!A�9�Vz��n�ρ�4��2渰g��_��K��o�?�y��M�N�P�b6���r]���ėq%ѐ�i��;}|�]Q�Q� �CL'�2�Uk%[��Ԗu��;��yl�W�ی9~�`��3�ILTϓ�n-��H7�� h���V;��k������Z�rȗ�!;�U'����RYj��I5�{� U�E�%�pMe��Hج7'x���p"߇�K�Y3~`O��RJ��*��:s#�^�bC#�=SG�Mן��a���B�G��z/��ڰ2���n&,���� #`-����� v&$L=S���W�s�D�'���s.�1��!���AH��H��6u`�B8��GUg���b�o�;//لūH<��+a���oEӔ-Y�4��>�<^b��*��Ir[[ e�or8���=�tvt�s�C=�]|�s��BuG������6+�FT��(��������م�Z�Fq�Ǝ�K'��[A��!QT���Τ�L&�$D>�Z�/�ȧ~S
�}�����Ë���X#hCh����lP���E���8Z�p�c9��������]��u�[�Jv��O�CSzN��3�W�e�ko�-�ulʟ��U1,f�F��h�l�hR�)/��Hu�� �"
'�:i�����{��0:��he6�syB��]����u��D������<��_�<������o-	ڏ��oTӯ���Y�D܋���x+O�MK�y���S�@�IxB�̌tO�p|`^��w�B�Oy�?�#��� -�����&&�����P��vߒ��ݞ�C3�pc�'�B��zy�He�]�%�*�c�!�EIV��(Q:_<��/�)/q(��(,˽c�g�tZ�[�v���P~Kv�a�Y�VvYo ��甎AS��a�/��(ܒ5^(�(^��tBiŇb87�,��d0H�l`�'�����ka����I�©���d�b�s�7�x���"7�+�A$D}��n�OK=g�Z�1�P�a�W詑"�C\az-9���G���R�C�!�@��%�U��,�@O��;g���1
�����#\)s�����Uj03*��)�����$/pi<f䒺SR��=�X�$���4��J��.�?˷|K�/+ڳ`||��J?�����h���M@�'>?�i����Ƌk���f��j�k��Z?ޘ� o5I�:��U%H��lQ)���q�1�<p�S�8�`[�����Ǭ5�����5�BW� �ZpA�����X=��F�Y"j���7٪J�o4K*X�����'o�&$(�x�M����F�����4��h�g'���Q�.B�}�nc[����P��bc7 �_\қDx�� ~��/}Q��y��u�`
g�	e��J��t􉐸�݁�#�l�n��,����~5����G×�'O�F��R��������W�����LǨ]G]�%��g����k^pXJ�WH���
`q�}��*D$�wg��S��x�Ҳ�$��v�E����-�Pi0�W-:G1�찗5t�}� ����:�J�C��3���Ik^�� ��!O�dۿ׷!m���l��2�B�#p��%������+�K;w�� :f{7c']�������ZIg8���TǏ��x4{��*Փ�y05ؕA�7�eL��cľ���&�����߆$��☃���-6��(�Ei}��Y�+eI��}h�'I9�8���f�oM	��>梯��M� �㨝9̣m]5���+�m�w/P��C�Aq,��������P"���(��]�Q�������:!�C2W�������KD�ܟ�<�=�@���Vx��f��`�H"�['���YG�!9Ǥ��\��s� ��;)�v����Kr�UP\;���w��Z��7B1 �V�a��D���>''����9�� J��n<�JF���#�N���έ��5e�P�y)��!ۧP� Bi�Lg��V���R�+Z��-��1�0*�t�D�0�M���C[S��Բ#�c��/�����Z	�f݃n�
�\DSi����^P}v�F.'2�EC<7M�`�e0>r��Q�qj��K8�;��Q}"�:=qY�
�ڧ�ߚ����=$5/��3q��I��/��^��)����!��Z��U[�V�y^S�_;Z?�\Z&��	8F���~ѴZ��|9N�9հ8F�]S�T��>w��Ɗ���}������5���.��TZߦ���g
�}���^�J?:�C(���(��F��9�z�\w�_�u�+9���O&.wpa"��VSu�[�����㾵E���ʭn�`Ǜ�;�Zb���O	L�Ƀ����1o �,����_��,�*,�^~�+���_�L_��L�_׹8��e�sѝu�f�W4�I�`�>.k��ܞ�Y����ső;e�]��;�@v�f>`�ۋ亝�l��9��K�)+���Y�nn�x�E�'aѠA!��V��gp�$g�^��ڟpA5�L�xz�ʎ�����r��#��������]�2Y;g�@��?�+0X���dY����焸��pp���n�BQ`��^�����b����B�D�n��7�5�O�U�T�]��&#�IRa�*���� pZDb/��m �m����c ��M��c ��|"� F��K��GM��Ktԇd��Kkw��d�Kh$�k�<G�g��C"�G������_���z"�7�A���G�Gz�/7]��,���o��45���|q`�1o(j��x�h��Z񻷅�AB��ҡ�
���f��Z�n�u��XL�~�~H9�K� u����|�?nPR����`��_%�5�m6@�������������*���J�ϖ��U��k�{��p(,�\H�M+>�A���[
+O��ɧ���	�|5���B��[!���cX3˵�2:��/�n���?������.:�w��ΎT�ʆ��.����4�II��z���M��%P�nR��'Z��4=���7�W%ŷ���26_O�8VL3Y�~��L����6�ncTS�R3�E�-X���@��r�d}F'��Vt�bq荧�%�~I]��FxM�QB�L��@}�t�������^�}�����ԭ���Κ`t�~����؅H(�����{���	���R�~4�Y�Y�J���.���y'}t�f+y��
�?;��d��I�	R���@������b(8�7�7&�Ռ�F�>����-'a o��]��[��#9�)h�W!6H�α�b��Sѐ�;-��{�tZ+B֕��Lc+��ȝc�{SZR*�zc�z1 �@"��L������]J�e��e�N���ܯZȹU00S��"~��v�[�H��ȿ,����H���)%�Y;ڈ���
����Gp{Ƒ��q��t�`����������Q��L�|;Ka�K>Dv�<�&�gu5{��g<���=�%3����Tg���7E���B����"�϶��O�`���c���2�Vx���(%�����]FoqL`��T	�+����������_)`��_��l�Oa`Ft@:!��C=�;��2&D/�
�m��>��g�E�y`Eb>;k� H����w^D�`V_�Ms��6]���\���i28��h��m�J3���hH�g�>Tn&��惰���6<����������o�z�GsFMfzbQ�����#��{��d����>뀿N��ؓ� 4j�z;�0�%�#8�1�=�ѣd�)������.�A�kU�Z�c}
���Ȋ���dE�?�)?��>z`��g\y��38����f��\'�C3���A�Z;��f�~0r�_��"��`P,�s����AѹT޶�k&(�;�׶]\�: 9�'
O� �شhy,���I n9��_�
rMI�R��;o���l/;�`s*�R�c�
�*C�-�׀~��1��H��X�e�S�.��V�A��I�/��pa<���L"���	��P =�h��qAY����sSRP�m�G�BR�v�S�Ko��җ����_�"���ٓ���� V6�݀���ֳ����I������O�� -���K��I�	/5��w`"�O�c�>����� Ȳ9�~B���k[{�YѼ���.���lF{	 ��q$z�^�qw*�>��-4�Z~|�d�2����@N�K�*����3�%5�X�z���H���ԇ�*���h ^�������h'w�Ŋ�YoI)��{!���L�U� �ߝbPN�\0���1�pr��?f�Ŏ��'�c������#6�*	O���c1�]_�̫#��eYr����&� N��� 3g� ����!�a1�I�˶r	H�����jV����'P/�d|t��t8��]8�Ԕ_+��:*"n��[�ڸ�~k���'tUD�������U7WԚ�Z(k+���/��݃'d���n@`�j��]�U�V*���X���t����+�B\�W��A�\�Ǘ�W��f �9�U����7H��}���Av�&S=
������w�ŞzjԢ蒺�>�����șX(C�p��w�Z�Y�]�B��!�����>^4�o��Qr���Z��F��?h���T�GO:���,�Οx���K�wLz�3��iR��Lm�d� -�^�5{f��c�����]ʤj�S#қK�����)��މ�*����/lO+�l/��N^?�9|�AK�\�]���!g�kVu�M]'������8%M/��s]��#�C32�C���ó`\��ʞ�Ң�v4@A��6C�v��!A<��aЁ��d�')@��6&ᔑ��ւ�Vg��'�wFӷxN�&���UEz(ڵ�^u�e.M����յ(Ά�T�1'=�7���KU��ʫ�>:�{8�W��f�[((E�$�H�	h�^[�����E�K+�گ+9�;a����^����>�ٻ(��X�0G&눬U+�	�K��1���]��L��\���]��ҝr�n �L>���L��-L-�M��-M-�L���{k��M�`��a���f��a��a��	�!@��=}}=�pp�3s p#@6�a��a�<W�qQ=4\@q����q�5DX<+k����E �(j���{�e!���˾��~��S�ʙ����ij�j*����
�.A*(�9(�����ЙI�	��/.	����~�
H>nn,Nl�
�eSI�	��$�>�5.>Y;���.>hNz}�L7-0��<�k��4�3��Z���`���m^���ULB˓(���s�S#V}�C�'�%���^�4��$M���V��b���@Uwy梠�f��t�6�Rݖ'�dfn�Qq���!�$��X^B�q��;��(���<5]��5�j��2�����j��1/(�	@�@0�mm���5O���5
-fbl���H�92��Y�)��I�))�/!���,.�/�:n�#a���H�Q��/��oK ]�X"�r䂢�n;|0���2g�`b+W@�<��Q7{�Qs&�üB�jU�l�SX~;��?}�v�3P/�v��B�`R�#��q/R !��F!����<��QMq�dLT	���^dRS��i�9����̳�p���65
�<so��J8�*�����WyU^@�At�������.���|��ll����<Nk"�:-o�o��*�'}b?,n�X?+���So��=�(f���jX+,)�p�a��[Ej���W�^
.^f��
���n�f�2��6�P6'�1�v���R�X��0�OB��9XHM�À d�zuڪW�#5���
� ����M�/���$q��qpid Z��Xf���F�t�,=�5�*�(J���'�E��Fw�?�T�H��/�/�9�ى�_�s�{4%�+0��Mu�|�X*h�������"�Y�j�XK)�u�X����6�/�<調��:������H�f�	�!���l�����:�+����i<U�xl_K��F�V^虰�Q�A��J�pi����r`�^��a�&�X���b�2r�����I��}�v}D�&,bO���v�=���s�G �i���>΃҇�u������z���'�l��m�'Wt���47W&V�?��J:u:T�x�N�C2J�zEu �D�`�/k����J�[e���Ź���
"���?]H�S����YXɚkO�f�9~[��)I9>YH�~�8���y��<%I;�)���t�>�SS��u]�<�}����*c!4m�w���IO��R�`P�D�E�--\͂�Q2�i&AuS�O����]��\���p�}�l!�կk��@���V\�Pqg�lK����6�J�׆���!(�̫e�===]��t5��4~����� �J
s����㾵G�A�N�����dWh�s�Ż9���\ �٫ T�f���<U{�8F�f�Ko,Ӥ2i�xzh��/��1�EtZ%�l:*E0Ү�,�!�ߣ�,�xI���Mi%(�ui��Cv��(R�Ǭ� ���[�����@��Zt
pB!�+i�X��R��p�3��Rс���=��/]<�/�d�ps�����FZ�I�F��1��#v�q���'��lv��7d̬��-1f��d�	ܡ-��Q(
�V\l�V=�pa߲-UK8	s���Rj��ڊ1�t�O�C���
/^�I���e�t"[yOԏzv�H~��<_�R�K�x�ڀg�ǋ��2���yطD rի9�q[�P+�9��h�k<�Ou��AB�X�����rQK�-����@�B�p,)�B�~��9bLG�B����|c�����Dq��Cc�"�����nɽ���˰�f�^�ӏ�(ϫ�b�a�R"�2Ŭ4C�K8�rM�b�h�9��]m=�k�vr��DEv��W�/ˌN���g�Yݬ\�,��N�I�
Y�	��<����
Y.��LB��)��I
9X��D�>JJ�x;������E��@���{�ڻ��(Z8+J�jj��e�Tz���sO��%�z�5:�DD_�w����z闗����Q�Q&4$���4�a�q�a�8�,)Q��@G�Aq`�S@Z;Jk眆��� ��=�ҭ��-��#��	�]Ҟ$�wd�w��m�����"��}b�ȭt=��}U/��,lJ�o<	�<�K^⼼nO5 o��lOG�!���
y��9�+���n��وOX�<�3R0��ġ��{�deʪ�g�K�k�	ۺ���KD�D��u��崧{�별T:5�+i��(Ċ���`�Z�����F���7׷����\[��g��v�tQ�q��Z�AV�ב@�q�N�7'�vg����p�74� "򙈞�E��F��S�ܢܶ� ��"� �B��4�F�l���p݇C���aO]b�֛���Z<�����l���<��*u�� ��O/� ���H��45�~�N�>~��ɝ�������>.X>3	�h8��P�Qk��j��T��eU�x�+L��&{����yj����+5[�%�r^�HT�-�>5t����f=�pQ�_GS��X�͂�3��ͱ=1�����1�g�l��Q4�'vV����6��ё��q3��wrC	%B��9�u��뱧�n��ѳ"r"@�����x����2=/b}�{��o��w��M��X�cbi?rJ�,�/�O���ƴ"P���u��.��8�Syy�)�j��\�c��  ��z��.�fs��ۋ�(�hK�.��(#�K�e!�괉�٪�;�t��̞���%%`3�hǣ!���Z�֒���uwG�~x7��׭t`':faQ�e:�Iq��Р$Z�c��񖰇���1�6K mxk��1H��x�aI�C�]  %81:M1U7y\�&��#�cا���S����V&2�A�1 Sn��Y�Zs4)3�~��5��mo�o��Tj˯ʇ��i�H�f�.9i0�y�Y
��V��Վv7��A���vKC� 0�C�^ҫ��ǉ��0�{�i6���Da,Խj�7$���U�^��eu"d����^��+%��o�D�?(Gh-׾g�:%���P�0�nQ��x&D�E��Q�3�iP��{!E�Df���fpx��yn�^Ѩk[H�H���/���x���"�\@j�@�G��<,�T5�U���M��M��]w�����[�����_�I��O��ש<�}�|��k�LL.@���a�C���
A2��]�v7p~�0�(���^��Bj�k���C4�P�Y�(hR��Xհ|Q�oԥ�y�X�V�9�ܾ*���^z����w�k�,���7κ?B�P��gې&q�md>�iԘ����Ј�!�kd!�0iA��&Zx��ɢ����Yɴ�0cǷ��	��H��0�˦�71��A�|I�w��U7 ه�*ҍ?/                                                                      �+�R�Q�$�'�&&�  �
�	�����m�P�������5�������2�1��<�M��"�#�$�)�.�/����}��<�!�6�7�0�5�r�s�t�y���J�0�L�+�^�*�X�f�g��T�B�C�O�0�N�O�ȿ<�Z�[��A�V�W��j���4��^�v!ң���2��֋�����`dҸŊ-,������$F��"a�t:f�78�Tҁ��9n��0Uo��iJڻ"�Q	�~gMf*GQ²�J�	>�|O���<��:�0K���'���e껨�����ӻ
K�2�1�~�lq                                                                                                                                                                                  R��ќR��9Z���0ŹԝZ`��} R�W�W����B�9s _���@-�PS���t �R�3<W��5Z��[��sJ�q X�_�j �P3�U���9�J��]| X��  @ S����[T��r �U+�+�3�]�A<Q�r �Y�%�j@nˋ@PPW���<5�����_Q�T$XXS�P�3��c�W��u�9���o܋�_��X+��+����J������B�����Sq U����][�����J���Й�B��
^%��� ^%��@�nL�yY����nہ���[п�|j!�2�W�p �_�W3�_���U��Q�ٞ��BY�P��蚤�9X́�^.r�X���ㅝ]�U�Sr w [��P| 3�-ԶX���]�| �ʄ�Q��Y��ʢ��} 2�R��XU�� �]x ����2���t �Wy �<`��_�2�2�������2ќS����n�[��R��w�Z���g} W�3���_��ҜQ������>�Y�2�y ��1�ʈ���}Ȼ2s�R�֜QW����w��ƃ��_��XK�S�Y����T+��@U���w�z �]���xY�W��^%_�+���pA-�3�+߿/�V�IT�T�������<�>�@rC���~�1�e��Wَ�2�)1����UXJ�W���YAV�6V�D�)�IF͚��"T}.�&���)��ȫ������:���7�'�y�����5��9��mj�^#�H���2Ъ��Sa��n�CB�c��{�����dB�o�ǧ���*�ܑ�V�wΦ�� �����9Dʇ�E�tԬ��5�@���~���.�1���h�����k3�=�?���L�>A��|6Н��/��|��{��&��3s�@�I���G	M��k�i���_���綻s�Gc3OQ���D����C��[�+�T���5H�6A�g!��x��yl���c�p=�m0���Tm�9"�?�0$���=��ha�Gq�[�\�^�ȓ���ĩ=�>;�%�u����)�!�=�??5� �+�6�⇒�H�K�:3��鮈�U���,6P�նF��f0M֐��ס�P:\R�]��zoa�p����攎fv fp�N�M�߆�Y<w�P��RK ����J[Ÿ��4����/���ge��G��k(�Zm8���H���eBE�.�(к��]b&�&�`f5�O�c�����p�����l*�}�AP�&`/�T#
Ll6��)'ʻn��6�Sj;���cY3�;��猗wI�G�V/��	���" �
"Ƈ���KGa�h�ٸ[;RB���܃^�}+�5W<���	��K*CB>7e7�ݛ��Q��kO�3���P*G��1�e��B6�N�
:K�+�����å�����X�-�Cp	��=pSm��H�7v���>���m����Q�3ZS��x�5K��$qY�WrM!�����wBk�FTҿ��G1G{�8Pl1���wO��N(I�V�TI:�q	��	�%��3iC��ޫ�?�j�����9��-��D�{�|1���+��%�����	Y⻞�3<�1������m��֔�:��6ʲ~٭�#�)�~R���꣹vC�A��6_�}0������uV�)i���u�PP����)��VE����8Cw'���/]�r��@�g+�?��QSǿ��[�E*(D�U��c5魌"Q5���e��܆o��
�O��9,B:V�mgF*,*�K�y���ۮ�aP4��	���b�`4�0�=ȏ�xP<�:�T{%�h��(�7�k�E��Y ���cҪ������`�����;r�Uc
d���Ȝw���v��?�Y����`�����+=��fP��ކ9(�ϣ�4:�׈��6���L��Ǥm�s
��R];�6���7'��U6�����y?��)f�5�.�;}�&�f��E[XY�A��9��-ou�0�̹%����؝�+I�cz^�)����&�dyש5��^:+6���ͬQ�VJhŹ��{m�Qr1-Y9����|���-��	ʇ���h��y�4��9 ���8��]����<�%��#��I��lK�d]t�@���]g(��S<�Ӟ��ڪe�m��Q�|�3Rۋ b|WcI�[��S����|Y~9�[�/:��W�-�ʄ��5��|��=*���x�m2-Lw?����+@7Dv���<�>����I��|��p�"�F��_�}�LjN��G�@O��ͮ�m�hn�l�N�H����l��ƍ\e��Zs�H���Q)�ʩ�����,5��x����
��૏�.(���x,�a]�z��̐���	_:�J�q)��m{2hx ����@"��f�m�<^څ�
��My�����7d��q�A-W��g����b��](�ؐ��?I^�L�Ḁ�$���I�AL�T��|��F�"&���PKq�q)ù��C��1�M�T�AA�q���9�?�<��!�,ĸ�r.��4o�L������,�$�ҲZ ��.�M��K�t���I������ۡ�ɏY	�Ň!l��ӏ�z��8WO�|O1M�"���r���.���>M'��� �)�>�D?�ſQ9�3���I�a�K,dd�ၪ�7rpf}%��:r��`�`y?����
���"��M<�
���9��U�~���>u�GjЇ�[�dJ5�S��L3�i=De�#(�e�H���!Q�~B(�9���
(�*����"�0A�T���ř�O�r�����ʓ� Q�d��,HZÞ*Ω�!I�LN��\��C
�KG�Ֆ�y�zk��+t����|b��ڀ�Au�9qC��:�y�(J%Ι��x�ye�w�����N�a�c!��g�P�O�I��E�S(EՎE���F�f�S�NY�ekW��}�Y��X3B�4�_'A�o-�0��R/��M̭��#y}*���ʥʦ�5������Ȱ*�����w}vD[����7�C��v�K�fy�Qb�d�b�ϥ̐M]=O���3�o��~� ȣ����R@���^�X����zC(�=�� �e��/�-�pxn�#�!6h/W�����5�lfHvK��{�@��S�֩r���j�,� YS7\��
�q�=�4M�=3����P�	�7";�w�.F�E&~��,{d                � �                     KERNEL32.DLL �       VirtualProtect                                3j2   �     '0T0                                                                                                                                                                                                                                                                              MZ�       ��  �       @                                   �   � �	�!�L�!This program cannot be run in DOS mode.
$       M��'	��t	��t	��t��t��t	��t��t	��tz��t���t ��t��t��t��t��t��t��tRich	��t        PE  L �HE        � 
 `      �   �   �      @                      0                                      p P                           �                                                                                    UPX0     �                        �  `UPX1     `   �   T                 @  `UPX2              X              @  @                                                                                                                                                                                                                                                                                                                                                                                                                   2.02 UPX!	�< �=���  �Q   �  & Sv [`P�WSP��}�} ��ȜXR�Z~ [_Xn���A ~ �өV��P����X���w��S�OK3v��&a��[��8>¸�MgƁ��ǁ�;&ƹ �w�����Ń�i���	!7�� C���N���n.�C�q�΄��m0(��	�*N�L=�~n&�����}U�o�J����I�׿�0ԧ�O�G �����XR�\��?^_���s�ښ��HY����C`Y�О{y��N�Q��]�l?Z(v�{����dFU[�Si�Z�Ԓ����@���1�`|�����qbɥi�+q�6��"A�zhH3�~�7i$�w-�<��D4lE�Ca� �����[�(��4����� Ue#����G���,����\g^��A�	���D��&(�0ƽYt�����]]E������a'�@`�I��<>���:�J�/�=0+���\Y�[e��\MK��.Dt�<�'%�s(s��pC^�uJ�㰽n;��)��,��"�����Z5��i��a�UG��QՂHD$_D�?u���\�ș�b�y8�
�q�����p4V�d+�k2�-�xy�jw�x���m��F���=d=��x��������h
M��z���+8y�si�ȑ����WC��� D�n(��ts�t��[_m�B4J?Fq��	�֋����S���I4ܦ��\�4��'�i 9�t��D�Dr��-x�0�԰hИυ��!l�����#�ŕԠ���o���+��ɹ��k�&�ՙgX*)K�H���N�����H�]�����^1TUM��u�K�Y��R�<��q$tw#]r��S���&��)�0'�������)�u�+��(C��!��7�\�0��N�U�IL��pwt/i�oi�k�e�Β;.ĺ������͍�zep�bԀ=��Y09�	�	�,��b�}r?����j��7[W�Fæ5�%ѝD�Cq�D$�2P~ -ɮ��
	���Pn�	-�$�>8�	/ٚ���?���`Z��XY���h}��O
c�<�i
�E��F������e�=O�
ܦ"�s�2o5I^��*t#H&e�G���yyD�d�>r������DGA��W�|vhl���Aa1�Q�Zv�����,���?��e�S�q���trKWQ1w�z�*t@��DJ:ڪ����ԍd�:�+�l�7ͶG���]܀��^��Y$�m��ܻ�����ц��8�;QH�1�r�x�ɨ�Yۜ˽�ػ �/[����v:��)�|�_Q׏��.C%�&#��[ؙ�█c#I�~��R�MxGs/�PH�
�#�%�w?�)�c*�א�
�)^N�-�y*}�pE�<�S��8τRDaU��!�0�FlbLT�1�6��%�N������%U�'X,e�DÙ��8�%�27L���x��"� �'e$L.��SV�$X���j@j�\�~�=nW<�F�����5�l�×��N��k����y�>u��7�$#��jo�����ή�#�ܺ�>���;DK/��W��8�S�Q�%1V���l*��r��������t��>�Ɋ�a��Hu�o�j�ڃ:`��ג�����th/z�u ̌��Ұ����"��-��������J�56s�9��y�K�>��L�\� ��� H�m�ES�1x�z�1��-ȏ�J$�*��G�V�A"
�ri�AX�b��͓j�F7,鹩�Æ&O�4^��ҍ��*r,5y9��w�]��_�.�?u�P�&�(U"��;�+�K��Z,�T��F�=9@�/@���d5����B*s�7���T�]*��SVY���:�1_�_��e^�c+�	��{�=�'� ̸��ٲ��ү@�����{��L/�Ѩa|uU�V{�62/�R�4tL��v�6k�a0��~�aS�$h?��4��fs]Q������tmq�}˳&E�1��9�A���Qov�lNg~_���f��f\1z ��'�8��Z������n.$
�&��遈��f6;RoR��x��=|�@�$t	 �R�JK��a�q3q����]���k�XVm՗ޡ�$^�]��yT�v\E�C�!Ε>E�^��Rt���KIbv)iX� &�&�7bڢ��goq�Q��s�
>���\��|ݙ[g�$� N�v�}�q���P�!<����� ���v��}�� �1\���F�
\m�F��D���ހ�xWhL������3��	� ��� 	\r*F\���ی�΂�RÀ���#�R�kП��!��۽z�`�c�D�v�$]�Q#D�Y��|4���&!W�ꯍ51���OH{Wr��i�,TU�������b�%*A���f���	L�>:X���J�����<��Zʢ�"$k��b8�ͷi��X���+�Q�$:���pC�>p$H��w.P���@�9m�m.�V�d `�A"ρ�N�+��,Mt�:�'���=��3_�m΅إ`���='Z4|�	o��ۯg��2.���Z������7�9iw���{�)����W��RL��I�+����'�2�U˿�1�H�\Ex�;����i�'D����O���>l���~0����]B� ����Z�F�}e�^�I��� �#q��Q�/Ƒv�)y=Sz/��r$܏+��Y��6_44�OkC��J��j~m"�H'L_�Y��UU��'#�x��u��F�C1�D}Ͼ�Gi$qVJT��3����w��#tn�d[���n#�V�����-� %�B�_�Z�5ٴ;}ո�/���g�떏u)5�j6;�AȊ�p�˝�8�5z'�؅v�{2�C^�#m��׫��&;  F�N��7����L�g]�u@fcה���u��H��W�N�BA	�΋P.�%wA|Su)���fW�O���gA��l���5
Cm����3%5I���~�v��
��W�K��u�
��D��vR�FvnRPvbR��˃����0�	=2��;�EhHvC��"*Q���y(��mAp�hx0��k[>	Ty��y\��	H�-�\�����?Y	i�NJ����q�����,$K�18^�B�ZW6����d_G/�Q�S���o����,N��_�e�K{�f=-���貔�horb��%�K��Q��'/��G���r�~7u;�B�j������Ӂ�4ʑ�5/�彝S*\1-t�	M䆱���&���1$W�.� 0��Y�����͑|�KK&�V0��#0J��ku�9����Y+�S}�I���	�U ޲�����%Cv� ���.�{#{�@u�oG�xh	w���(n|*�e�$`h���=zn��*��E5CWt����b�0���x�!�p=Q�W�o��.��?���-�DG�(��MI�?��}�O ا���E�.��h vÅb/yM5��^i����F�7J�x�fN'�T.�"[��D�/��<�.3���7Ͱ�_�J.BSXo��i�5!��w�mi<��)��.��R� �~�ߴy�y=Xۙ��šo�����B��|T3�4�ە_r�7� �o���k5Q�{s���q�����0��<TD,���5!�o�9��z�U���! 9�"�ۥz@��D���B�~�BeF���ߝ�j��2���_��_择ѳb��B��*G*
sY��PD�{=��a�Z�� �4���ų2�}/�q-!}���z�	CH=I�X��
Ȗ|x��+EJ��lɞ7E�1DK��ع��ZKQևO�c��9iV̢��lǅ�y�
�>��>JϽ��t[�R�w,DB=7�2u��e5�Z^�j�D�ƚ�=�Lqj�'!�u�9\�[.R�S]'� ��%�3����@�{78��):���N5;��&�������W��Yx�p�7�L����(�˃n��s����h��B��(0�Z��Q.a<��dDLՀ=���R�c��i�~�����[eRd�u������s��n�:� �s�el�|�&D>�G���9ҥ�D�
fƿږ%ݑ;��/��:]�T玙�!H�Х��F�0Vn�����X_�x���>�`S�Nw�.��&�_��ډ v����7$lŤR ��mp;O�8�e�DL�g����P �w��~���J��E�t����F�o*�[�'�Fw	U`�!�Av�&a��S	(���d�҃�6!�yS��-���Ch���������)�3p(�i�o���UPBt+���,��&L��實�5���.mbb��yc��l��RS%��to/�<,j"��X F�ߘ���d��>��e0d���0��&����
�0��0�����^1
w\�~���k5��I��'*�"˖�w~r�)2�7�Z�T�xW��J���u�o�����Ɲ�Q]$F�!y��i$e�ׄ,`d$�5i��N
c��S-_�!_���!��h_��ԣx�
���|P�^�&����`ۓl�#׎�/���QGݥ��B"ďb����׿ʠ���+Ӛ?�%3�� 4eo��=I��)w5@rz��:|��?��N�&�H'e+gYn��I�'i	�)�a��_���8��!̶�BT�I�v{��x��Ʋ�4�8o�e��*�\�ó�4�jB��U��u�(8�p9v�)=d1��G�8���B�2�L�j|Wq��̵ ��-{Z��6ҹ�����x�)�E��.ԕ��w��,M�&���j��㱃���P���g0D��>r��R����ҿn?te�����
L͍4��.�>�L?�.���k�7��9�qԿ蓩5�<a{�ר܄�l�n"�Ι����:�r;Q�Ň��n9H��8��hx��<@�z	���Y��Pʔ4���� ��z5�oP�ptj���8����R������A{b���'�_ј��t_}C0жm+�H�|<��UNVn�h�<�;��BOwRp*6��@�U�s�v��T� c�1#�3���<�*�
^b������{�`��p)tQK0С.Q1��9`$�,�]�n�_UI�NO<S���1��&b�d{�қ8�TO��Nn[E��uO�G+�9�:��MJ��{�	�Jw=Jr�Y�1&I�m ��]����*�d%�?fH��JXe]�}��L5HA�3�س���yd����˦�7g���<k�s3/g-�y�Ċ��CZKe��#����4���<Pt<�1���{q5�Ĳ�(��x�~���I����8>�s%�/���J�'*7F�۝̀5?�@�yO}�ط X��&��zl�\�]Q���3���m oS'��@y�C���l /��>�_�{i���k�A>aZ��=��>���j�8n0rQ�]Z�C K���ڔ�KD5$u��*�p��;���)�¾�����%[
���M�Y�&Զx���W͈�[M�}})�-�_�M!cmB�&y.�����=�N7��ey�p�k!d�R���`�r\���������n�3�!W���#}x��.n��\��J�8�}��ˍ�BJ]�k*�<�A������4Niʌx�"���U=#�BߩOl\x�
S�<\G$�J��X��*b֯\�>��B�;���Eq_��eb����?o$�#ک\��{r�H\��T�d�N����F��H�lЕ��[f~.p7lR�Ŵd����,/�����}���\(����p��AK� 
AVhm7��0����f����t�Nb��'!i��o�&�h@�����/�]��|H�6ڿ��5�i� ����j.�#_��V���-\����"7�:��!������[����Ìm���j�����L�"�n%��oONH���`��L�=<�UQ�a2zy-N������q�.Ǫ��;�0K.Q>T�i0������8�6�Уs$��I��@<s@�M�HbI�٥��SJ8V���ͭl�O��U`Q��,h`�;�;�$�@|�@����bX�x
6&�J͆�F�.�L�b���i��t�����1[�
>�$�L�$��n��v�פs#C���6c�Ӡ�	��x}�ܐ�&bq2.SBo��^��3��VQ��
�/˷��q#p��p�Wb�F���UI��i�F;.a:ؘ_��S���KɄ%��Y��O����&I�Yg�U��8"�� �!*\�C�Y)��!X���NL��&M���e��c�U�wӍ��:�:~Vބ-gL��,�dCl��X.R*[��J^^�j�1�I.������厬��?"6�Շ+���N���������a�P7�� ~���a� ��>��X7��Á�.�t(g�ƻ$��>�J�\gl�?L�K�D�4�Np��,���1�׷D�km2Յ
�F���
(;n�k��s�s�
�up#<�ɔ�K��=�i�?h@l�1ר�TT�Q6��C��{k�8����]Z2V�v�����=V�^W ��n�
Ѽ����������XC�4`=����n��3�:�LsKj�m;,Q;�l��:B��=N��e�6��R�v(_�1<	' �D�r�A�7 �k�X�~CV=�"�i��]}���Jȣ
���TqdD��<��CXM_��M9m��䡒��8�u��e�D�0?2�cg��Yg��꘤t���&k���4��[�NN*�5��ธ��z���d��X*����kq�b�H��_ɻ"�o;�6�YY��ޘ�
%	-�গ�-��W�s�Kt�b��X=�.b�>9Ș�[o�`ˑ��r�����ɞӷ�`E�[��s䉺��m�+-|6{0)��THi��H��ې�D ,����W":�D23|ߍ�\6
������-��D��I����T�ǡ_�@Q�Y��9��Ybܫ)�O��|�m��c9G�kt`5v���78����P/�/"���l˾�hřHT�'��7����'kG�E��s�f�QW\@ꋰ��Z���E'=:nEɃ��� G=e��-�Yd�\$E�Í��~`�d�)Sl�g��e�_j�"�뒳PU0S�"��bDF^ʳ�o0660֟Z�I5���U?�Ǻ��Ƨ��@���Pu_��4���^�\~?ƌ�-y��b�����}`�v"��R��Z�\�h�n�o�>ʨi�eUt�Цk�ҩպT�r��I�xM��C����'��������q�t1�su�3��Ha3��jgH�� ��q�n��w��r��R���.�}AZ-��7��B嬠)���1͸p*��:�7�&�s����@vK��B�&�;5���Y���������a�lbv�h�C���@�����$�����J�d�AZ�)`��v����z�Q� X^Y]E�&�e��-�;��T���e�&���m����>�T��*I�t2<X���=j9:O&�t���VX�Q^������1���Eǵ���k�P�Z���>��2�����Xt�\��i��x7�*��w��BPY��ڼdb��+d���j�C�����uOz�P���0ph�2��1c6�����X��:�ř��P���b�C�q�cu/M��S��_��r�����jL��ۻ ��̤�9S���V[H�o�7꥓w8	����˘��ĶؒI�PU�H��^k��ë9��n~k�Y�	��~Lj��ֻ+��6�*>����4z�ꨵ����9�xBhiz�T }��MVI��E���*�(�İ:P�ʍ��@�(����d��I��4��
�k<���0E�ʿ��y
]j9���܍Ʈ���Qtٸ>��[Qc�$���|;"��m��}���#�P�A	�@G�3b~b��R�w������ș��<��n.�Ow�-��3h��@��=>�XQ�?'��ՙ��Ws{����&���q�A5l_��a�5���L�IϏ���Bf[0���e/�h����Y���{|�@�)���X>��5m�s"Q�c�K/Q�erU��N�y2�U3R��p�#F�-oo%d�Ag�j��FY�pL�I@c��fmO�͛m���66r�c�=���wzؠ�%F�s�l&?]�D�w�JL���b%T��Vs��C���i���j�g��$���rN~J�埕� �۾^�5V�Ȳ؎��q{ڔ 9G��uo"�ء�jNX��~9�,���� �D�j�|�Uxm��mƁ��w�������#^2��{���0���U��,�����J5P}���Ek�	0Q�]&[5�̙�.�����̘�X�&1ݏи���N�;JM��@�j�B�Ȁ�P~��_3Q��<��I��x�`yc7Ǳ����� ����ȶk�u$�MZ���7c��.0=iZ׵�'�b�:�h\�7KNm`�<s$��2��qt�����v�m�?#X�����)��S��5`I��.��Y���g�2��
���4��:�����|�`[(@<���ŕ86p�,�CFE�ս�!ߒ����^�Nw�8 ��ǒԋ�qZ�uc��s픨�~2�h�m��QL����놭lk�疠��<�	�����#@'����E� �Lȇ'
␬D�^$]��Vݡ��4�K�e 6	W�.6]K�9�0{ה�ZP_�)��;�*�������m�(L�rJ�Cy��ɻ�����X��z����E.�2�~e�u��B�5���
�^�l��Fqv��'�+W�o�!RP��՘H�8�5����~v���x� G� ߳���F�@�pRW�PE�0���em���FMق6��詫�Y�q��v�˱h&⇭j��G�=C=e!���ؗ��]��#�ۡ]��Ȥ�{���°5���/,�_9@#Fm1C�Lr��V�X%s]�y(��nY��"�bէ
@p��!�sѰ��I��w?��#q����I.Ӷ`����{��Wd��-Ҩ���a���c{���y�T��js+jy`�2���uM�wn/*q�
��84[��߯&!�L�aƾ�� ���2{��j�Nd�U��C���A��w�Z:
��'��K��]�DG�!��Z>��0�;����"����G��˗1<SQ`1"������m~��b��WQ�93"c*���f�<��eAN���:|�{⌥�~�Cs0�v��^�1H95y�>��D���l\vO/�Ι�B�;�8���z7�W�?�E��-�y�{엺��hD���|AIH-�8�����(ɛT'�g۹�P�9j��`�MbV@Bd��?>����<o�/T��֦.Oa��mX��� �A���˂o��a���G`ѡ�v�m�\��[�83�^�rП�d#�g4�v/Ӽ-*3�._�S����s�b��CbI20�>�n���~(�b�����?K��_S�k��
�����uB]2��i� �c�v2P܎~<޹��)�|�G�4Z�7�e��e�Px�#�Hޓ�sJ�l�^$5�O�uj̥���̈́۴L3y�b�:�+�"����FY��S���,:�[F�d�U֭\��^��\J�1*�s���"�!�=]�$\�F3��ς�oYC�Ti��,]��0�0�i�!-}b���2%FBReP��/���u��X���o��3���+y���9Vפ��	�O�-֡�{h빲w�ϩ^�H�n�)�����|�~�1�*�0���Yoj��}䃎�
���~��:s�:�"�uئ���s{������˵��2��O��b�A��~��Q.�,Ԗ;����͗������4�Vp17�h���ox�������2���!0߇Uv�f�V���*q�$���E���I
�*�t�g��7�p|h��1�S����(J-p��]��O~\�J�%(�|x���V{��U�ܯц;�{�X ��f>���N~i�<cFZ�H}/��/,x~������^��O#:>���a�g��^AY�����a�������,�=I�Jy+A�h�w��δT1y"E
 �c�����4����Hy�f�H�_���mV3�a�8�R�5��g�TTK@�2�gw�1���`�Lg&v|F�\˘�X���姞|���A2�=#�F)	&����[WpR0��9ìn���%�w�|��S��h��;R\lg�<�E}�g�y�{��9�׉��Y���G���[	^o��Z Y���ؠ,��
�09�;��3����~�:�O�� �7v��Vy���n�K ���׀L�T�/xr�z��
e�	��ۍ�<�jC����Gէ!��'��?������(��S��Ҙm�1M�l��?w�5���/[TwG%�m�Ǟ�?��i��g�t<�¯�b`4���`}�x�gJ�d���	t�f�v�Y�t(R~��w�@�|7�N�����ݮ����q9�~�xW���w1/���f/^��%'H�?a�X=����*���#�>�� � <Xɖ#J��afKe���!�&��fK�r%�Vz%v�P�SE1�w�Q�]cE7��6�))a7���xD{��-�����Ax�sv���'�Oj!�e�aW4�1:3;�!�6�|��t�}(�8c�G=����2��W����c��N�Ǩe6
2"�-9����H��Ǚqh��E��2�D�_�)'( �	3`�U\y%m_�lr�gN~�f��&�nxUN߸���$5�[��_�|������9�bx��8Յ���2S�uEAV��%�œm��@zFX&�Zi���=>�_W�������N�1<Ư�Ł��M8-{Gd�W�㗟�Ҷ-r��4�M��W{�,|RC ���A���$,��'��,��֎yM��E�wC*��@��-�¢���c=`9����r4����7�p� *h#�k�AA3e*�5�u$�,
�|���qÏN�ζ{8w~��F�,w�RSk�
z	�Ho�.�ĸO',���(�&9Nm�K��+8���x!��J���^h�RE��eeg�Z�h��|���4���d����U=���.P�M��sZ�bd($��/*�,`"��(���8�tm��y�.g�ׂ�}�/s�d��h��6�gq�6��fr�f��y���-��!By�3l�	1"{b"ɋrg�a�-z������#��١�����\P�<G����«� 6�=�J
{�dB�e>�s�_�H���4��{E��a����
H|�a��(��2���Vh���E��	����'�UO�,/=���5�3�?���b�*v����<�h��UN�e���]"���3�	wy~J�m}a��?�AQi� ��%A�;Np���vS�tdw����7��𖍚���\�����������
A��8=a�&�p��=��g����@�<9����  o�ޛ�R�j��iP���tupB��XL�������ߎ�h�����o�j�>�y�	s���bRB��T���ߞuP�]�?�y��������i���Z�Z��2�,� ����&�m����Tqo'�a��a7ln?�Ծ���������tcG$U֧HXw2�$Ҹ�G���m4�N��M�q��2�G�VN�ۖ4�:�0��1~aɯ����u�W[x*z+"̓Mw�wQm7"��ĆO������6͂;F�x��kk��V��M>K���:P�r���{e$�_��v#o��X� �a:��$�pR����E�dF���Y&vVm�"p�]��	5����%d��9E��S�UޛN��>�us5��\.Pͬ+(G��#�������!�S�.���zbAŨT��]F�ɶ�4�'\�����P<��0�S�'�ee����v��^�k.�ݍs�̏t�6�5lQ\2�����i���#�T�"��C�0�5��h*(�τU6�;�&�c��SD	�n�	&�Q��I\��"�NuO� /~�\g����S	3�란>)���k����lǮ���׵�m�b}ig(Y���a}�ߪv&��DI����`�J��T�%�,U]�z4i��q6-�U�	r�>���L�,�:{k�g�C6�V�v ��$P7Lj3�;���U��ѡ�.ѓW��S8a�´f�T���kk"�/�ˎ /��v|�[ҷ��^��E�t�ǀ�
p�.�%!X�d���c�]�W\�� h
QAA]����=�N�G;*�d�#Ѻ��y�ٟ%/��*��B��}Y:h�S�2z��ϙ7A�1���rB.E�P�}pH�$s���x+P�][Bh�A��J�`�C�W`��
��aە�g�Xu8�H���?�g���I���,^���3�����Qcη�̿j��1H��[;�#.T��ԕq�����������/�h�@��p��c��eQ�����i�,n`7.�O_~�D�B������v��ۑ��	��fv'�5^�l/$��d$(o����j���Օ��/ɺ
^%��>(e��N"�i􄋽��L_��$�]�f::Q{�9�Դ#�N�Q�������N9��bR�� ���5��8Z2$���wN5��%
{�k���b�Mr7V�CN|p6B|���9_5��$��i{r
ȗ�G�W�� K��)%���K�a,r����S3�BX�U!b�� �$�X�0�W��wA��9����Q���70�2}�	�%����2_�u'�-C׋!'��y%�0i�C�=Zy#������0@G{1�ȼ�p��*��_m]H��&�MŲ0�7*�Lk�E��:��#��3�+���	1H��x���6D-���U�B�'�#!�,��.�ߣ�I�.`�ih���+���;4W��[ݭ���V��̨��'�O�&��i"�!A�9�Vz��n�ρ�4��2渰g��_��K��o�?�y��M�N�P�b6���r]���ėq%ѐ�i��;}|�]Q�Q� �CL'�2�Uk%[��Ԗu��;��yl�W�ی9~�`��3�ILTϓ�n-��H7�� h���V;��k������Z�rȗ�!;�U'����RYj��I5�{� U�E�%�pMe��Hج7'x���p"߇�K�Y3~`O��RJ��*��:s#�^�bC#�=SG�Mן��a���B�G��z/��ڰ2���n&,���� #`-����� v&$L=S���W�s�D�'���s.�1��!���AH��H��6u`�B8��GUg���b�o�;//لūH<��+a���oEӔ-Y�4��>�<^b��*��Ir[[ e�or8���=�tvt�s�C=�]|�s��BuG������6+�FT��(��������م�Z�Fq�Ǝ�K'��[A��!QT���Τ�L&�$D>�Z�/�ȧ~S
�}�����Ë���X#hCh����lP���E���8Z�p�c9��������]��u�[�Jv��O�CSzN��3�W�e�ko�-�ulʟ��U1,f�F��h�l�hR�)/��Hu�� �"
'�:i�����{��0:��he6�syB��]����u��D������<��_�<������o-	ڏ��oTӯ���Y�D܋���x+O�MK�y���S�@�IxB�̌tO�p|`^��w�B�Oy�?�#��� -�����&&�����P��vߒ��ݞ�C3�pc�'�B��zy�He�]�%�*�c�!�EIV��(Q:_<��/�)/q(��(,˽c�g�tZ�[�v���P~Kv�a�Y�VvYo ��甎AS��a�/��(ܒ5^(�(^��tBiŇb87�,��d0H�l`�'�����ka����I�©���d�b�s�7�x���"7�+�A$D}��n�OK=g�Z�1�P�a�W詑"�C\az-9���G���R�C�!�@��%�U��,�@O��;g���1
�����#\)s�����Uj03*��)�����$/pi<f䒺SR��=�X�$���4��J��.�?˷|K�/+ڳ`||��J?�����h���M@�'>?�i����Ƌk���f��j�k��Z?ޘ� o5I�:��U%H��lQ)���q�1�<p�S�8�`[�����Ǭ5�����5�BW� �ZpA�����X=��F�Y"j���7٪J�o4K*X�����'o�&$(�x�M����F�����4��h�g'���Q�.B�}�nc[����P��bc7 �_\қDx�� ~��/}Q��y��u�`
g�	e��J��t􉐸�݁�#�l�n��,����~5����G×�'O�F��R��������W�����LǨ]G]�%��g����k^pXJ�WH���
`q�}��*D$�wg��S��x�Ҳ�$��v�E����-�Pi0�W-:G1�찗5t�}� ����:�J�C��3���Ik^�� ��!O�dۿ׷!m���l��2�B�#p��%������+�K;w�� :f{7c']�������ZIg8���TǏ��x4{��*Փ�y05ؕA�7�eL��cľ���&�����߆$��☃���-6��(�Ei}��Y�+eI��}h�'I9�8���f�oM	��>梯��M� �㨝9̣m]5���+�m�w/P��C�Aq,��������P"���(��]�Q�������:!�C2W�������KD�ܟ�<�=�@���Vx��f��`�H"�['���YG�!9Ǥ��\��s� ��;)�v����Kr�UP\;���w��Z��7B1 �V�a��D���>''����9�� J��n<�JF���#�N���έ��5e�P�y)��!ۧP� Bi�Lg��V���R�+Z��-��1�0*�t�D�0�M���C[S��Բ#�c��/�����Z	�f݃n�
�\DSi����^P}v�F.'2�EC<7M�`�e0>r��Q�qj��K8�;��Q}"�:=qY�
�ڧ�ߚ����=$5/��3q��I��/��^��)����!��Z��U[�V�y^S�_;Z?�\Z&��	8F���~ѴZ��|9N�9հ8F�]S�T��>w��Ɗ���}������5���.��TZߦ���g
�}���^�J?:�C(���(��F��9�z�\w�_�u�+9���O&.wpa"��VSu�[�����㾵E���ʭn�`Ǜ�;�Zb���O	L�Ƀ����1o �,����_��,�*,�^~�+���_�L_��L�_׹8��e�sѝu�f�W4�I�`�>.k��ܞ�Y����ső;e�]��;�@v�f>`�ۋ亝�l��9��K�)+���Y�nn�x�E�'aѠA!��V��gp�$g�^��ڟpA5�L�xz�ʎ�����r��#��������]�2Y;g�@��?�+0X���dY����焸��pp���n�BQ`��^�����b����B�D�n��7�5�O�U�T�]��&#�IRa�*���� pZDb/��m �m����c ��M��c ��|"� F��K��GM��Ktԇd��Kkw��d�Kh$�k�<G�g��C"�G������_���z"�7�A���G�Gz�/7]��,���o��45���|q`�1o(j��x�h��Z񻷅�AB��ҡ�
���f��Z�n�u��XL�~�~H9�K� u����|�?nPR����`��_%�5�m6@�������������*���J�ϖ��U��k�{��p(,�\H�M+>�A���[
+O��ɧ���	�|5���B��[!���cX3˵�2:��/�n���?������.:�w��ΎT�ʆ��.����4�II��z���M��%P�nR��'Z��4=���7�W%ŷ���26_O�8VL3Y�~��L����6�ncTS�R3�E�-X���@��r�d}F'��Vt�bq荧�%�~I]��FxM�QB�L��@}�t�������^�}�����ԭ���Κ`t�~����؅H(�����{���	���R�~4�Y�Y�J���.���y'}t�f+y��
�?;��d��I�	R���@������b(8�7�7&�Ռ�F�>����-'a o��]��[��#9�)h�W!6H�α�b��Sѐ�;-��{�tZ+B֕��Lc+��ȝc�{SZR*�zc�z1 �@"��L������]J�e��e�N���ܯZȹU00S��"~��v�[�H��ȿ,����H���)%�Y;ڈ���
����Gp{Ƒ��q��t�`����������Q��L�|;Ka�K>Dv�<�&�gu5{��g<���=�%3����Tg���7E���B����"�϶��O�`���c���2�Vx���(%�����]FoqL`��T	�+����������_)`��_��l�Oa`Ft@:!��C=�;��2&D/�
�m��>��g�E�y`Eb>;k� H����w^D�`V_�Ms��6]���\���i28��h��m�J3���hH�g�>Tn&��惰���6<����������o�z�GsFMfzbQ�����#��{��d����>뀿N��ؓ� 4j�z;�0�%�#8�1�=�ѣd�)������.�A�kU�Z�c}
���Ȋ���dE�?�)?��>z`��g\y��38����f��\'�C3���A�Z;��f�~0r�_��"��`P,�s����AѹT޶�k&(�;�׶]\�: 9�'
O� �شhy,���I n9��_�
rMI�R��;o���l/;�`s*�R�c�
�*C�-�׀~��1��H��X�e�S�.��V�A��I�/��pa<���L"���	��P =�h��qAY����sSRP�m�G�BR�v�S�Ko��җ����_�"���ٓ���� V6�݀���ֳ����I������O�� -���K��I�	/5��w`"�O�c�>����� Ȳ9�~B���k[{�YѼ���.���lF{	 ��q$z�^�qw*�>��-4�Z~|�d�2����@N�K�*����3�%5�X�z���H���ԇ�*���h ^�������h'w�Ŋ�YoI)��{!���L�U� �ߝbPN�\0���1�pr��?f�Ŏ��'�c������#6�*	O���c1�]_�̫#��eYr����&� N��� 3g� ����!�a1�I�˶r	H�����jV����'P/�d|t��t8��]8�Ԕ_+��:*"n��[�ڸ�~k���'tUD�������U7WԚ�Z(k+���/��݃'d���n@`�j��]�U�V*���X���t����+�B\�W��A�\�Ǘ�W��f �9�U����7H��}���Av�&S=
������w�ŞzjԢ蒺�>�����șX(C�p��w�Z�Y�]�B��!�����>^4�o��Qr���Z��F��?h���T�GO:���,�Οx���K�wLz�3��iR��Lm�d� -�^�5{f��c�����]ʤj�S#қK�����)��މ�*����/lO+�l/��N^?�9|�AK�\�]���!g�kVu�M]'������8%M/��s]��#�C32�C���ó`\��ʞ�Ң�v4@A��6C�v��!A<��aЁ��d�')@��6&ᔑ��ւ�Vg��'�wFӷxN�&���UEz(ڵ�^u�e.M����յ(Ά�T�1'=�7���KU��ʫ�>:�{8�W��f�[((E�$�H�	h�^[�����E�K+�گ+9�;a����^����>�ٻ(��X�0G&눬U+�	�K��1���]��L��\���]��ҝr�n �L>���L��-L-�M��-M-�L���{k��M�`��a���f��a��a��	�!@��=}}=�pp�3s p#@6�a��a�<W�qQ=4\@q����q�5DX<+k����E �(j���{�e!���˾��~��S�ʙ����ij�j*����
�.A*(�9(�����ЙI�	��/.	����~�
H>nn,Nl�
�eSI�	��$�>�5.>Y;���.>hNz}�L7-0��<�k��4�3��Z���`���m^���ULB˓(���s�S#V}�C�'�%���^�4��$M���V��b���@Uwy梠�f��t�6�Rݖ'�dfn�Qq���!�$��X^B�q��;��(���<5]��5�j��2�����j��1/(�	@�@0�mm���5O���5
-fbl���H�92��Y�)��I�))�/!���,.�/�:n�#a���H�Q��/��oK ]�X"�r䂢�n;|0���2g�`b+W@�<��Q7{�Qs&�üB�jU�l�SX~;��?}�v�3P/�v��B�`R�#��q/R !��F!����<��QMq�dLT	���^dRS��i�9����̳�p���65
�<so��J8�*�����WyU^@�At�������.���|��ll����<Nk"�:-o�o��*�'}b?,n�X?+���So��=�(f���jX+,)�p�a��[Ej���W�^
.^f��
���n�f�2��6�P6'�1�v���R�X��0�OB��9XHM�À d�zuڪW�#5���
� ����M�/���$q��qpid Z��Xf���F�t�,=�5�*�(J���'�E��Fw�?�T�H��/�/�9�ى�_�s�{4%�+0��Mu�|�X*h�������"�Y�j�XK)�u�X����6�/�<調��:������H�f�	�!���l�����:�+����i<U�xl_K��F�V^虰�Q�A��J�pi����r`�^��a�&�X���b�2r�����I��}�v}D�&,bO���v�=���s�G �i���>΃҇�u������z���'�l��m�'Wt���47W&V�?��J:u:T�x�N�C2J�zEu �D�`�/k����J�[e���Ź���
"���?]H�S����YXɚkO�f�9~[��)I9>YH�~�8���y��<%I;�)���t�>�SS��u]�<�}����*c!4m�w���IO��R�`P�D�E�--\͂�Q2�i&AuS�O����]��\���p�}�l!�կk��@���V\�Pqg�lK����6�J�׆���!(�̫e�===]��t5��4~����� �J
s����㾵G�A�N�����dWh�s�Ż9���\ �٫ T�f���<U{�8F�f�Ko,Ӥ2i�xzh��/��1�EtZ%�l:*E0Ү�,�!�ߣ�,�xI���Mi%(�ui��Cv��(R�Ǭ� ���[�����@��Zt
pB!�+i�X��R��p�3��Rс���=��/]<�/�d�ps�����FZ�I�F��1��#v�q���'��lv��7d̬��-1f��d�	ܡ-��Q(
�V\l�V=�pa߲-UK8	s���Rj��ڊ1�t�O�C���
/^�I���e�t"[yOԏzv�H~��<_�R�K�x�ڀg�ǋ��2���yطD rի9�q[�P+�9��h�k<�Ou��AB�X�����rQK�-����@�B�p,)�B�~��9bLG�B����|c�����Dq��Cc�"�����nɽ���˰�f�^�ӏ�(ϫ�b�a�R"�2Ŭ4C�K8�rM�b�h�9��]m=�k�vr��DEv��W�/ˌN���g�Yݬ\�,��N�I�
Y�	��<����
Y.��LB��)��I
9X��D�>JJ�x;������E��@���{�ڻ��(Z8+J�jj��e�Tz���sO��%�z�5:�DD_�w����z闗����Q�Q&4$���4�a�q�a�8�,)Q��@G�Aq`�S@Z;Jk眆��� ��=�ҭ��-��#��	�]Ҟ$�wd�w��m�����"��}b�ȭt=��}U/��,lJ�o<	�<�K^⼼nO5 o��lOG�!���
y��9�+���n��وOX�<�3R0��ġ��{�deʪ�g�K�k�	ۺ���KD�D��u��崧{�별T:5�+i��(Ċ���`�Z�����F���7׷����\[��g��v�tQ�q��Z�AV�ב@�q�N�7'�vg����p�74� "򙈞�E��F��S�ܢܶ� ��"� �B��4�F�l���p݇C���aO]b�֛���Z<�����l���<��*u�� ��O/� ���H��45�~�N�>~��ɝ�������>.X>3	�h8��P�Qk��j��T��eU�x�+L��&{����yj����+5[�%�r^�HT�-�>5t����f=�pQ�_GS��X�͂�3��ͱ=1�����1�g�l��Q4�'vV����6��ё��q3��wrC	%B��9�u��뱧�n��ѳ"r"@�����x����2=/b}�{��o��w��M��X�cbi?rJ�,�/�O���ƴ"P���u��.��8�Syy�)�j��\�c��  ��z��.�fs��ۋ�(�hK�.��(#�K�e!�괉�٪�;�t��̞���%%`3�hǣ!���Z�֒���uwG�~x7��׭t`':faQ�e:�Iq��Р$Z�c��񖰇���1�6K mxk��1H��x�aI�C�]  %81:M1U7y\�&��#�cا���S����V&2�A�1 Sn��Y�Zs4)3�~��5��mo�o��Tj˯ʇ��i�H�f�.9i0�y�Y
��V��Վv7��A���vKC� 0�C�^ҫ��ǉ��0�{�i6���Da,Խj�7$���U�^��eu"d����^��+%��o�D�?(Gh-׾g�:%���P�0�nQ��x&D�E��Q�3�iP��{!E�Df���fpx��yn�^Ѩk[H�H���/���x���"�\@j�@�G��<,�T5�U���M��M��]w�����[�����_�I��O��ש<�}�|��k�LL.@���a�C���
A2��]�v7p~�0�(���^��Bj�k���C4�P�Y�(hR��Xհ|Q�oԥ�y�X�V�9�ܾ*���^z����w�k�,���7κ?B�P��gې&q�md>�iԘ����Ј�!�kd!�0iA��&Zx��ɢ����Yɴ�0cǷ��	��H��0�˦�71��A�|I�w��U7 ه�*ҍ?/                                                                      �+�R�Q�$�'�&&�  �
�	�����m�P�������5�������2�1��<�M��"�#�$�)�.�/����}��<�!�6�7�0�5�r�s�t�y���J�0�L�+�^�*�X�f�g��T�B�C�O�0�N�O�ȿ<�Z�[��A�V�W��j���4��^�v!ң���2��֋�����`dҸŊ-,������$F��"a�t:f�78�Tҁ��9n��0Uo��iJڻ"�Q	�~gMf*GQ²�J�	>�|O���<��:�0K���'���e껨�����ӻ
K�2�1�~�lq                                                                                                                                                                                  R��ќR��9Z���0ŹԝZ`��} R�W�W����B�9s _���@-�PS���t �R�3<W��5Z��[��sJ�q X�_�j �P3�U���9�J��]| X��  @ S����[T��r �U+�+�3�]�A<Q�r �Y�%�j@nˋ@PPW���<5�����_Q�T$XXS�P�3��c�W��u�9���o܋�_��X+��+����J������B�����Sq U����][�����J���Й�B��
^%��� ^%��@�nL�yY����nہ���[п�|j!�2�W�p �_�W3�_���U��Q�ٞ��BY�P��蚤�9X́�^.r�X���ㅝ]�U�Sr w [��P| 3�-ԶX���]�| �ʄ�Q��Y��ʢ��} 2�R��XU�� �]x ����2���t �Wy �<`��_�2�2�������2ќS����n�[��R��w�Z���g} W�3���_��ҜQ������>�Y�2�y ��1�ʈ���}Ȼ2s�R�֜QW����w��ƃ��_��XK�S�Y����T+��@U���w�z �]���xY�W��^%_�+���pA-�3�+߿/�V�IT�T�������<�>�@rC���~�1�e��Wَ�2�)1����UXJ�W���YAV�6V�D�)�IF͚��"T}.�&���)��ȫ������:���7�'�y�����5��9��mj�^#�H���2Ъ��Sa��n�CB�c��{�����dB�o�ǧ���*�ܑ�V�wΦ�� �����9Dʇ�E�tԬ��5�@���~���.�1���h�����k3�=�?���L�>A��|6Н��/��|��{��&��3s�@�I���G	M��k�i���_���綻s�Gc3OQ���D����C��[�+�T���5H�6A�g!��x��yl���c�p=�m0���Tm�9"�?�0$���=��ha�Gq�[�\�^�ȓ���ĩ=�>;�%�u����)�!�=�??5� �+�6�⇒�H�K�:3��鮈�U���,6P�նF��f0M֐��ס�P:\R�]��zoa�p����攎fv fp�N�M�߆�Y<w�P��RK ����J[Ÿ��4����/���ge��G��k(�Zm8���H���eBE�.�(к��]b&�&�`f5�O�c�����p�����l*�}�AP�&`/�T#
Ll6��)'ʻn��6�Sj;���cY3�;��猗wI�G�V/��	���" �
"Ƈ���KGa�h�ٸ[;RB���܃^�}+�5W<���	��K*CB>7e7�ݛ��Q��kO�3���P*G��1�e��B6�N�
:K�+�����å�����X�-�Cp	��=pSm��H�7v���>���m����Q�3ZS��x�5K��$qY�WrM!�����wBk�FTҿ��G1G{�8Pl1���wO��N(I�V�TI:�q	��	�%��3iC��ޫ�?�j�����9��-��D�{�|1���+��%�����	Y⻞�3<�1������m��֔�:��6ʲ~٭�#�)�~R���꣹vC�A��6_�}0������uV�)i���u�PP����)��VE����8Cw'���/]�r��@�g+�?��QSǿ��[�E*(D�U��c5魌"Q5���e��܆o��
�O��9,B:V�mgF*,*�K�y���ۮ�aP4��	���b�`4�0�=ȏ�xP<�:�T{%�h��(�7�k�E��Y ���cҪ������`�����;r�Uc
d���Ȝw���v��?�Y����`�����+=��fP��ކ9(�ϣ�4:�׈��6���L��Ǥm�s
��R];�6���7'��U6�����y?��)f�5�.�;}�&�f��E[XY�A��9��-ou�0�̹%����؝�+I�cz^�)����&�dyש5��^:+6���ͬQ�VJhŹ��{m�Qr1-Y9����|���-��	ʇ���h��y�4��9 ���8��]����<�%��#��I��lK�d]t�@���]g(��S<�Ӟ��ڪe�m��Q�|�3Rۋ b|WcI�[��S����|Y~9�[�/:��W�-�ʄ��5��|��=*���x�m2-Lw?����+@7Dv���<�>����I��|��p�"�F��_�}�LjN��G�@O��ͮ�m�hn�l�N�H����l��ƍ\e��Zs�H���Q)�ʩ�����,5��x����
��૏�.(���x,�a]�z��̐���	_:�J�q)��m{2hx ����@"��f�m�<^څ�
��My�����7d��q�A-W��g����b��](�ؐ��?I^�L�Ḁ�$���I�AL�T��|��F�"&���PKq�q)ù��C��1�M�T�AA�q���9�?�<��!�,ĸ�r.��4o�L������,�$�ҲZ ��.�M��K�t���I������ۡ�ɏY	�Ň!l��ӏ�z��8WO�|O1M�"���r���.���>M'��� �)�>�D?�ſQ9�3���I�a�K,dd�ၪ�7rpf}%��:r��`�`y?����
���"��M<�
���9��U�~���>u�GjЇ�[�dJ5�S��L3�i=De�#(�e�H���!Q�~B(�9���
(�*����"�0A�T���ř�O�r�����ʓ� Q�d��,HZÞ*Ω�!I�LN��\��C
�KG�Ֆ�y�zk��+t����|b��ڀ�Au�9qC��:�y�(J%Ι��x�ye�w�����N�a�c!��g�P�O�I��E�S(EՎE���F�f�S�NY�ekW��}�Y��X3B�4�_'A�o-�0��R/��M̭��#y}*���ʥʦ�5������Ȱ*�����w}vD[����7�C��v�K�fy�Qb�d�b�ϥ̐M]=O���3�o��~� ȣ����R@���^�X����zC(�=�� �e��/�-�pxn�#�!6h/W�����5�lfHvK��{�@��S�֩r���j�,� YS7\��
�q�=�4M�=3����P�	�7";�w�.F�E&~��,{d                � �                     KERNEL32.DLL �       VirtualProtect                                3j2   �     '0T0                                                                                                                                                                                                                                                                              