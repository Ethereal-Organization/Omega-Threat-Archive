MZ�       ��  �       @                                   �   � �	�!�L�!This program cannot be run in DOS mode.
$       � ��A���A���A���I���A���M���A���M���A���I���A��JI���A���A��\A���M���A���M���A��Rich�A��        PE  L �U'F        � 
 �   `      �k      �    @                      @                                      � �                                                                   ��  H                                           .text   *�      �                    `.rdata  �,   �   0   �              @  @.data   �#                     @  �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                ��  �hA SU��$�  V3�W��$�  �<   h   V�t$$�t$�t$(�D$ �D$<x�@ �D$@p�@ �D$Dh�@ �D$H`�@ �D$L   �D$P   �D$T   �D$X�D$\�   �D$`  �D$d   �D$h�t$l�t$,�E   ���@ ��;�uǅ�      ��  3��   ��V�E$jP�  �����D$t��tǅ�   �  �  ���E��  j ���@ �M$j jQ��  �������uǅ�   �  �Z  ��t%�U$j jR�  �������  ��u�D$NuۊD$j j��C�M$SQ���@ ��tǅ�   �  �  �D$���  �U$j jR�C  ����tǅ�   �  ��  �E$j jP�  �������uǅ�   �  �  ��t%�M$jj WSQ�c  ��;�tǅ�   �  �  �; �E`��uS�,�  ���E`�U$j jR�  �������uǅ�   �  �H  ��t%�E$jj WSP��  ��;�tǅ�   �  �  �; �Ed��uS���  ���Edj j��C �M$SQ���@ ��tǅ�   �  ��  �U$j jR�)  ��<tǅ�   �  �  �E$j jP�  ��<�D$��  <��  �|$j ju2�M$Q��  �����uǅ�   �  �l  �U$j jR�  ���[�E$P�  �����uǅ�   �  �:  j ��M$jQ�  �����uǅ�   �  �  �C3�f�f���   �D$ ���H��   ��tǅ�   �  ��  �U$j jR�,  �������uǅ�   �  �  3���v6j ���@ �E$j jP��  �������   �;���   GA;����   r��; �E\��tP���@ �ÍP�@��u�+�@Pj ���@ �5��@ j �E\�֋}\�Ê@�G��u�S�  ���6�5��@ 3�j �֋M$j jQ�m  �����t]�;G��rދ�5��@ �D$$���   �|$ub�U$j jR�6  �����uǅ�   �  ��  j ��E$jP�  �����uǅ�   �  �  �C3�f�f���   �D$ �   �M$jj h�  SQ�>  ������C t�E`��uS��  ���E`���   ���j   P���@ =   s\�U$jj h�  SR�E   ��  �C �E\����tP���@ j �֋ÍP�@��u�+�@Pj ���@ �E\�ˋ��A�G��u��D$H��@ ���   f� ��   HtYHtǅ�   �  �  3�f�ERf��u�D$ jf���   �ELjj���   �у���E(uǅ�      �n  �E8   �N�UL3�f�ERf�����   uf�Erjjjf���   �у���E(uǅ�      �'  �E8   ��E8   U�U����t���   �  �|$��   j �֋E(�5��@ jWP�օ�t%�M(jWQfǅ�     �օ�tǅ�      �   �E(�T$RWP�D$$   ��@ �|$�t   �M$jjj�M,��@ ����E$uǅ�      �n   �UH�}pj f� �Ut���@ jf�Er�E$WP�օ�tǅ�      �;�U$�L$QWR�D$$   ��@ ǅ�       �j ���@ �D$ ǅ�   �  �}$���  ���$    ��I �|$�D$��$l  P�D$   Qt�U(��U$R��@ �|$�
   uY����   ����C �C�S��$p  �Sf��$n  f�C�|$u�E,�5��@ j QSP���T�E$�5��@ j j
SP���A� ���   ����5��@ j jS��Z�Sf��$z  f�S��$|  �C�M$Q��j ���@ ���   ����  �D$H��  H�9  H��  �T$$f�D$ S�Utf�Er���@ h� j ���@ �؅�uǅ�      �r  �}(�u$�   �|$l�L$h3�9t�lt@��r��u�   �t$p�L$h3���v�U,��9T�lt@;�r�;�u��@s�M,�L�l�D$h��;�v�ǋM,;�v���T$(Rj j �L$tQ@P�D$<  �D$@    ���@ ����  �E,�T$hRP�dC  ����  �U$�L$hQR�NC  ���  �Et���D$   tf�}r ��$|  u�Ep�U$�L$QPj h��  SR���@ ����
�t$0��  �; ��  �C����  �C����  �CHt9���*  �S�ҍC�   t�s�ʋ��t$0�z�; PG�5  ����C�   ���   f�;��;�f���   �D$   ~6j���   R�U(j ��+�P�;QR��@ ���  ���   +�Ɖ��   �M(�D$hPQ�4B  �������T$R��$�  Pj h��  �K
�C �C � �C�U(QR�D$,   ���@ ������   ��$�  �T$f��$~  R�C�EpPf�K�U$j �O
QSR��@ ����   ��   ����ǅ�   �  �}$��R����  ǅ�   �  �  ǅ�   �  ��  ǅ�       ��  ǅ�   �  ��  ǅ�   �  ��  ǅ�   �  ��  ǅ�   �  �  ǅ�   �  �  �E(jP���@ �U(�M$�T$l�D$h   3���I 9L�lt@��r��u�L$p�D$h   �D$$�����;ыD�D�D$(�D$,    v�ʍT$(Rj j �D$tPAQ���@ ���#  �U$�L$hQR�@  ���  �U(�D$P���   QR�D$$   ���@ ���E(jP���@ j ���@ �M(Q���@ ����}(uǅ�   �  �   �D$$��t;��   tǅ�   �  �   �|$j u$���   �Sf���   j
f�C�M$SQ��h�   �]f���   f�S���   j�C�M$SQ��j ���@ h�   �1�E��t%S���@ U�U��_^][��$|  �@  �Ā  �h  U��  �����   �|$v�D$ ����   �T$�D�4Ph\�@ S�M?  �U\���ҋ�t�p�@��u�R+��hT�@ P�'?  ���b�P�@��u�+T$$�QR�B  ��j ���@ �Íp���@��u�+Ƌ��D$ P���@ ��QhL�@ �V��>  SU�U��S���@ U�$   ��$�  ��_^]3�[�.?  �Ā  ���������V�t$���   ��   ���   SUWP���@ �F ����   Q���@ �F\���=��@ tP�׋F`��tP�׋Fd��tP�׋Fh��tP�׋Fl��tP�׋F(����=��@ ���@ tjP�׋V(R�ӋF$���tjP�׋F$P�ӋF,����-��@ tjP��j �ՋN,Q��V���@ j ��_][^������Q�D$P���@ �ȁ��   Q����R�T$����Q�D$��Ph��@ R�=  �����̃��hA V�t$���D$t~Wjjj��@ ���D$$Pf�D$ �t$���@ �T$(f�D$
�p�@��u�+�=�  ~��  Ƃ�  
���  3Ʌ�~	�4A;�|�j�L$Qj PRW��@ W���@ _�L$^�r=  �����������������̋T$3Ɋ<a|<z~<A|<Z~<0|<9~<.t<-uA��  |ԃ��ÍA�������̋T$V�t$�N��d$ ��  ~�������3�;�|/�<a|<z~<A|<Z~<0|<9~<.t<_t<-uI���A^Ã��^������̃�U�l$VWj@U3���<  ��������  S�D$$���e  d�D$     �k  ��+�+�Q�/R�U�����߃�����,  ��+�FV������t8������t$ �  ��  �  ��+Ã���   j.�W�C<  ������   +�;���   �.<.��   �|.�.��   <-��   �|$$���e  ���D$    ~\+�V�T$���ƍH�L$��    �@��u�+D$;�uR�+RV�=  ����tf�T$�D$���e  @��  ;��D$|��t$ ���e  i�  ��+�@P�+Q�R�@<  ���e  i�  +���D8 ���e  ��@���e  ��t$ �~�/j@Q�G;  �������|���[_^]�����SU�l$VW�|$���Ǌ���:�u��t�P�^��:�u������u�3��������tUW�=  ������tRj
W��:  ������t�	8^u%j
W� �:  ������u�ǍP�@��u�+48�D$�PW� �������_^][��������̸Dk  �>  �hA SUV��$Tk  ��$Lk  ��W�P�@��u�+�@P3�U���@ �؊����$�e  t��+��I ��P��<  ���7�FEF��u�L$Qh��@ S�+ ������T$Rh��@ S������D$(Ph��@ S�����L$4Qh��@ S������$�e  ��0��tx3�3��~M�|$�ǍP��I �@��u�+T0���  s*W��4�e  h��@ P��8  ���$�e  ��E��  ;�|���$�e  QhN  Ƅ4�e   �W8  P�!�����S���@ ��$Pk  _^][�9  ��Dk  Á�  V3�h   V�t$�t$�t$�t$ ���@ ;ƉD$u�   ^��  Ë�$(  ��$$  SU�D$W����   3Ʌ��L$(u���   ��u�N$�L$,�   �L$(���   ��u+3���v�V(�I 9T�,t@;�r�;�u��@s�V(�T�,�D$(�F(�N$;�v@��A�L$ Qj j �T$4RP���@ �؅��8  �9  �N(�D$(PQ�7  ����   �L$�T$R�V(���   Pj h   Q�   R�|$(���@ �����   �F��t-UV�Ѓ���t"��$4  i��  ;���  i��  P���@ �|$3���$    �T$�L$R�V$�FpPj ��+�P�QR��@ �؅���  �;�|ϋ��   �T$���   �Յ����   �T$t9��;�3�b   �+  �Y  ��}�=�A 3'  t�]   �  �����   ���   ���F����N$�D$(PQ�h6  ����   �L$�T$R�V$�FpPj h�  Q�   R�l$(���@ ����~}�\$S� �T������l$3�D$P���   P�F(j ��+�Q�+RP��@ ����   �;�|ы��   �T$���   �ׅ����   �T$�������;�������c   �3��   ���w����=�A 3'  �g����]   �����W����^   �T$R���@ _][��^��  þa   ��[   �ھ_   �Ӿ\   �̋N(jQ���@ �V(R���@ �F(����3�뫋F$jP���@ �N$Q���@ �F$����3�������������́�  ��$  ��$  V��$  �T$Rj �D$j �D$�L$P�NQ�t$(�D$$   ���@ ��uj P�T$RV���@ ��t���^��  ��D$^��  �������̋L$�A��tQ��YÃ�V�t$��W3��P�@��u�+�=�   v���   �3Ʉ�t��<.uG���<0r<9w	�D1A��u�<1 u^��uY�D$P�L$Q�T$R�D$P�L$,Qh��@ V�:  ������|+�T$�L$��3ыL$��3ыL$��3�R���@ ��t!�= �@ V�ׅ�uV�ׅ�u_^��Ë@��_^�����������U�l$V3���}^3�]ËD$W�|$ j WP�l����ȃ����u_^3�]ËǙ���S�؋�i��  �����  ������|$ ����I �T$�F���t;�t;t$}�D$USP�����ȃ����u�[_��^]������������̃��hA V�t$ �D$�~(�W�D$   �.  �F\��t1���   ��u'P�E����������   u_�d   ^�L$�'3  ���jjj��@ ����F(u_�   ^�L$��2  ���f�NR�VLf�L$j�L$QPf�D$ �T$���@ ���u_�   ^�L$��2  ��ËF8=   ���   f� }-�u)�F(�T$RWP��@ ���ub_�   ^�L$�2  ��ËN(jWQ��@ ��t_�   ^�L$�Z2  ��ËF(�T$RWP��@ ���u_�   ^�L$�12  ��ËL$_3�^� 2  ����������������U��j�h��@ d�    Pd�%    ���ESVW�e�h   3�PW�}����@ P� 1  W�����@ ;�t��   rh �@ �M�Q�}��<<  �U� ��+@ ËM�E_^d�    [��]���������������U��j�h��@ d�    Pd�%    ���   �hA �M�USVW�E�E�e�PQ3�R�]����@ ��;�P����C  �5��@ �փ�th �@ ��$���P��$����;  3��$   ��\���󫍍X���QǅX����   ���@ ��uh �@ �� ���R�� ����V;  ��h����   ;�th �@ �����P������0;  3�3ҍ�T���P��,��������S��0��������j(��(�����4�������������ǅ8���   ��T������@ P� �@ ��uQ��=�  th �@ ��@���Q��@����:  ��T���Rj(���@ P��@ ��uh �@ ��L���P��L����:  ��,���Qh��@ Sǅ(���   ��4�����@ �=@�@ ��8���R��T��������Pj��(���QSR�ׅ�u$��T���P���@ h �@ ��H���Q��H����:  ��=  u$��T���R���@ h �@ ��D���P��D�����9  �M�U�EQRP���@ ��T���SSj�����QS��R��P����׋�T���P���@ ;�u)h �@ ��<���Q��<����9  ���@ ��.@ Ë�P����M�d�    �M����.  _^[��]����������������U��j�h��@ d�    Pd�%    ��  �hA SVW�E�3�ƅ���� �?   �������Mf��e�h�   ������P3�Q��}����@ ��t>�u������VR�0  ����t'h �@ ������P� �������8  �E �Q/@ Ê]�M�d�    �M����.  _^[��]� ��������������V�t$W�=��@ j jjV��j j h  V��j j h  V��_^�U��j�h��@ d�    Pd�%    ��  �hA S�E�VW3�ƅ|��� �?   ��}����f��3��e�ƅ{���3�����@ ��|���@��u���@ ���@ �M�M�E��u���|�����A�B��u��]��|���Rh�.@ S���@ ��|�����th �@ ��p���P��p����7  ��|���QVV�5��@ S�֍U�Rj j S���֋؅�u$��t���h �@ ��t���P�Q7  ƅ{��� �1@ Å��5��@ t!j jjW��j j h  W��j j h  W��j jjS��j j h  S��j j h  S�֋M���{���d�    �M��P,  _^[��]�����������U��j�h �@ d�    Pd�%    ��  �hA S�E�V�uW3�ƅ���� �?   �������f��3��ɉe��E�u!������h �@ ������P�b6  �E ��1@ Ë}h�   ������QW���@ ��u������Qh   jW���@ ������R芣  ������VP��-  ����t
� 2���]�M�d�    �M����[+  _^[��]� ���U��j�h�@ d�    Pd�%    ��  �hA S�E�V�uW3�ƅ���� �?   �������f���3����e��}�u!h �@ ������P�������r5  �E ��2@ �j.V��*  ��;�t�  �}h�   ������QW���@ ��t
V������R�������Ph   jW���@ V������Q��,  ����t
� 2���]�M�d�    �M����[*  _^[��]� ���U��j�h �@ d�    Pd�%    ��  �hA S�E�VW3�3ۈ�t����?   ��u����f��e�hH�@ 3�h@�@ ��H�����t�����L���h8�@ Q��D�����P�����l�����p����?)  �(�@ �,�@ �0�@ �}���U؊4�@ j�W�E܉M��U�]����@ S�����@ ��   uh �@ ��d���P��d�����3  �M8uh �@ ��X���R��X�����3  h�   ��t���PW���@ ��uh �@ ��\���Q��\����3  ��t���R��  ����t�����t�����I ���:u:�t�P��:Vu����:�u�3������;�th �@ ��T���P��T����J3  �uVh01@ W���@ 8th �@ ��`���Q��`����3  ���@ h�  ���@ �U�RSSW���@ ;�u#h �@ ��h���P��h�����2  ���@ �|5@ Í�D���QP���@ ��D�����H�����l���BQ@W��l�����p������@ ��p�����l������Rjh  W���@ �M�d�    �M�   ��'  _^[��]� ����U��j�h0�@ d�    Pd�%    ��`  �hA �E�SVW�e�3�3ۈ������?   ���������@ f�����@ �   �h�@ �}����@ �E؋Ef��M�8��U��]�uh �@ ������Q��������1  �5��@ S�֋}h�   ������RW���@ S�֍������E������:u:�t�P��:Vu����:�u�3������;�th �@ ������P�������Z1  �uVh 2@ W���@ 8th �@ ������Q�������/1  �U�RSSW���@ ;�u#h �@ ������P�������1  ���@ �7@ �P�w������M�d�    �M�   �L&  _^[��]� ����U��j�h@�@ d�    Pd�%    ��<  �hA SVW�E�3�3��������?   �������f���   ���@ �}��e�h�   ��������uPV�U����@ ��t$�M�Q������R�(  ����t�EPV��������M�d�    �M�   �%  _^[��]� ���@ ��7@ ��������������U��j�hP�@ d�    Pd�%    ��   �hA �E�SVW�e�3�ƅ���� �?   �������f��3�ƅ���� �?   �������f���Eƅ���� ��  �>  �E�    ��������@�A��u�������P�Н  �}��V�5��@ W�օ�uh �@ ������Q�������=/  ������Rh�   jP���@ ������P������Q��&  ����uh �@ ������R��������.  SW�օ�������u������h �@ ������P��.  ��  PW�֋؅�u$h �@ ������Q�������.  ƅ���� ��9@ ø   PW�֋���tƅ�����������5��@ j jjR�֋�����j j h  P�֋�����j j h  Q��j jjS��j j h  S��j j h  S��j jjW��j j h  W��j j h  W�֋M�������d�    �M��f#  _^[��]ËD$SVjP2����@ ����t1W�=��@ j jjV��j j h  V��j j h  V��_�^��[�^��[���U��j�h`�@ d�    Pd�%    ��SV�5��@ W�}�e�h�  W�E�    �֋؅�u�E�h �@ �E�P�N-  jW�֋���uh �@ �M�Q�E��2-  ���@ � ;@ Ë5��@ j jjS��j j h  S��j j h  S��j jjW��j j h  W��j j h  W�֋M�_^3�d�    [��]��������������U������  �hA SVW��$  3��D$ ��   �|$�Mf��h�  �D$PQ����@ �u�T$VR�,$  ����t2������$  ��!  _^[��]� ��$  ���!  _^[��]� �U��j�hp�@ d�    Pd�%    ��8  �hA f���@ S�E�VW3�3ۈ������?   ���������@ f�f�U����@ ����@ �e��UȋU�Eؠ��@ �M܋��@ R�E⡴�@ �MĊ��@ Sh  ƅ�����ËMЉ]��z�������;�uh �@ ������P�������h+  �=��@ S��h�   ������QSV�   ��tB������R詘  �E�P������Q��"  ����u�U�R������P��"  ����tSV���@ S��V���@ �M�������d�    �M��T   _^[��]�ƅ���� �=@ ��U��j�h��@ d�    Pd�%    ��  �hA S�E�VW3ۈ�����3��?   �������Mf��e�ƅ������]���������$    �A�B:�u�������P�ŗ  ��������Qh 3@ ���@ 8�����t$h �@ ������R�������$*  ƅ���� ��=@ ËM�������d�    �M��o  _^[��]����������U��j�h��@ d�    Pd�%    ��  �hA SVW3��E�3���������  �������e��E�Ph   ������Q��u�u��X  �U���;�} �������P�I�����F���E� ��>@ Ê]�M�d�    �M�����  _^[��]�����������U��j�h��@ d�    Pd�%    ��  �hA S�E�VW3ۈ�����3��?   �������Mf��e�ƅ������]���������$    �A�B:�u�������j.P�X  ��;�t�������Qh�5@ ���@ 8�����t$h �@ ������R�������(  ƅ���� �?@ ËM�������d�    �M���  _^[��]��U������  �hA ��$  W3��D$ �?   �|$	�f���E�T$+Њ�@��u��D$Ph07@ ���@ ��$  �   �m  _��]����������U��j�h��@ d�    Pd�%    ���  �hA �E�SVW�e����@ ��������@ ������   �p�@ ��t���󥤹   �@�@ �������,�@ �0�@ f��
   � �@ ��<����f���\����8�@ �
   ���@ �������4�@ ��d������@ ��h������@ ���������@ ��`����<�@ ���������@ ���������@ ��l���f���@ ��$������@ ��,������@ f���������@ ��0������@ �M����@ ��(���f���@ �U����@ �M����@ f��4������@ f��U����@ ������E�f���@ 3۹	   �l�@ ��h�������������ǅ����    f�E��f���   �8�@ �������f��
   ��@ ��0����f���   ���@ �������f�3��������?   �������f��������3��?   �������Mf���]��������A�B:�u�������P��  �=��@ ��3�f��}9��k�d�����RS��;���   ������QVP�{�����;�th�  ���@ 3���$    f��}.��k�d�����PS��;�tIVP�N�������th�  ���@ 3�f��}lf��������Qu������Rh��@ ������P�#F�T���F���k�d������Ph8�@ ������Q��  ��������RS��;�t>VP�"�����ƅ����M������d�    �M��  _^[��]�ƅ��� �HC@ �F�[��������U��j�h��@ d�    Pd�%    ��  �hA ���@ SVW�E�3�ƅh��� �?   ��i������@ f�����@ �E�f���@ �M�f�E؉e��E̹   ���@ ��h����UԊ��@ ���@ 3�PSƅg����M��U�]����@ ��;�uh �@ ��X���Q��X����#  j�V���@ �   uh �@ ��T���R��T����#  �M��h����A�B��u���h���Ph@;@ V���@ ���@ ��h�����th �@ ��\���Q��\����I#  �=��@ S�׍�h���RSS���@ V�Ӆ�u��`���h �@ ��`���P�#  j �׍M�Qj j V�Ӆ�u$h �@ ��P���R��P�����"  ƅg��� �+E@ �P�X������M���g���d�    �M��+  _^[��]������U��j�h��@ d�    Pd�%    ��  �hA S�E�VW3ۈ�����3��?   �������f��e�S��]���"  P�"  ���"  ����  ���5��@ ��A h�  �֍�����R�������:�uh �@ ������P�������
"  �������P�I �@:�u�+�sh �@ ������Q��������!  ������R�O�����������P�������������Q�Q���������R�e���������������P��������J����}F@ ËM�d�    �M�3���  _^[��]� ������j j j hPE@ j j ���@ ��tP���@ �   �3��������̃��$Pj(���@ P��@ ��t`�L$Qh��@ j ��@ ��t@�L$�D$�L$�L$ 3�j �ɋL$j ��j�D$�D$Pj QB�D$$   �T$0�@�@ �$R���@ �����U������4  �hA SVW��$<  3��D$    �I   �|$j��I�����j j�G  �؅���   �D$PS�D$(  �$  ����   �u��I ��t�D$;�t�L$QS��  ��u��iPj h� ���@ �=��@ j ���׋T$j j jR���@ j ��h�  V���@ �D$PV�D$    ���@ �|$  u	j V���@ V���@ ���@ j�}�����S���@ ��$<  �  _^[��]�Qh�@ �L�@ ��tVh��@ P�H�@ ����tkWjj ���@ Pj�D$P��j ���@ �L$�3���vAS���@ 3��LQ�ӋL$�|u��9T$u�DP�e����L$���G��;�r�[_^Y���������������̋D$�8 t�L$�T$S8u��X@��u�[���������������U������  �hA VW��$  3��D$ �?   �|$�f�h4�@ h�@ ��D$h8�@ P�^  �D$ ����t�D$�8~u� -�H@��u��L$Q�  ����tKP�B  �UR�����5��@ ��h�  ��j �֍D$P�  ����th �@ �L$Q�D$   ��  �T$R�  ��$  ���S  _^��]��������������̋D$V��3Ƀ���N�N�Nu��A �F��^� ��u	���@ �F��^� ����̃��L$�T$�$Ph?  j QR�D$  �4�@ ��t�$P�8�@ �����ËT$�L$Q�L$R�T$�D$Pj QR�<�@ ��t�$P�8�@ 3���Ë$Q�8�@ �   ����������������Q�L$�T$�$Ph?  j QR�4�@ ��t�$P�8�@ ���YËT$��V�p��$    �@��u��L$+�PR�T$jj QR�0�@ ��^t�$P�8�@ 3�YË$Q�8�@ �   Y��������������Q�L$�T$�$Ph?  j QR�4�@ ��t�$P�8�@ ���YËL$�$QR�,�@ ��t�$P�8�@ 3�YË$Q�8�@ �   Y���������������̃�SVWh?  3�SS3��(�@ ����u����0�D$,h?  PW�$�@ ����t�L$QV��@ ��t�|$t3�V�5 �@ ��W��_^��[�����������̃�SUVWh?  3�WW3��(�@ �؅�u����c�D$0h?  PS�$�@ ����u3��H�L$QjV��@ ��u3��2�|$u+h�  ���@ �T$RV��@ ��u3���|$u�   �- �@ V��j���@ S��j���@ ��u���@ V��@ ��_^][�����SVWh?  3�SS3��(�@ ����u����8�D$h?  PW�$�@ ����tj j j j j j j j�jj�V��@ ��u3�V�5 �@ �����@ W��j ���@ _^��[���������̃�SUVWh?  3�WW3��(�@ �-��@ �؅�u����P�D$0h?  PS�$�@ ����t7�L$QjV��@ ��t%�|$u h�  �ՍT$RV��@ ��t�|$u3�V�5 �@ ��S��h�  �Ջ�_^][������������̃� VWh?  3�WW3��(�@ ���D$u����p�L$,h?  QP�$�@ ����u3��Uj j V��@ ��t�S���@ Uh�  �Ӌ-�@ �T$RV�Յ�t!�|$th�  �ӍD$PV�Յ�t�|$t3�][V�5 �@ �֋L$Q�֋�_^�� ������U������  �hA ��$�  3�SVWƄ$�   �@   ��$�  �f���]3��D$ �@   �|$�f��3�Ƅ$   �   ��$  �f��T$���+ӊ�@��u�h��@ h��@ ��$   h8�@ P�O  ��$(  ���Њ@��u��|$+�O�OG��u��������ȃ��|$O���GG��u����@ ���@ f���@ ����@ �Wf�G�O
�|$O�GG��u����@ f���@ ���@ �f�Gj �O���@ ��$�  RShX�@ h  ��,����������   ��t=��u��$�  P�L$Q�  ����t}ShX�@ h  ���������u}�D$P��T$RShX�@ h  ��Z�������t*hD�@ ����3Ƀ����������$�  �  _^[��]�hD�@ �����hD�@ �d������   ��$�  �o  _^[��]�hD�@ �_�����$�  3҃�������E  _^[��]����������������U������(  �hA ��$$  3�VW�D$ �   �|$	�f��3�Ƅ$(   �?   ��$)  �f��3��'   ��$�   󫍄$�   P3�Ǆ$�   �   ���@ �=��@ j��hx�@ ������V�׃�$�   u ��$�   uf��$  u�MQ�	����
hD�@ �m�������thD�@ ���������u�   hp�@ �E�������uhp�@ �������hh�@ �'�������uhh�@ �������h\�@ hR�@ �T$h8�@ R�p
  �D$P���������u�L$Q������hL�@ hD�@ ��$0  h8�@ R�6
  ��$8  P��������u��$(  Q�_�����h8�@ ��������uh8�@ �A�����h(�@ �t�������uh(�@ �#�����Ƅ$(   3��?   ��$)  �h�@ h��@ f���$0  h8�@ R��	  h(�@ ��$<  Ph  ��2�����$H  ����� 
  _^��]������������U������  �hA W��$  3��D$ �@   �|$	�f��h  �D$Pj �P�@ �L$Q�v�����$  ���	  _��]���U��j�h��@ d�    Pd�%    ��  �hA SV�5L�@ W�e�3�h��@ �E쉽X�����h��@ ��h��@ ��h�@ �����@ W�#  P��  ����\���Ph  ���@ ��A Q�}��������A ��R��X����E��  ����X���P�E������e  ����@ �M�d�    �M��  _^[��]ø�T@ ��ø�T@ ������Q�hA �$�D$P�  ������A uj��  ������$3��j  Y� �������U��j�h��@ d�    Pd�%    Q�ESVW�e�P�E�    ��  ���M�_^d�    [��]øBU@ ��������U��j�h �@ d�    Pd�%    QSVW�e��E�    ����������   �M�d�    _^[��]ø�U@ ËM�_^3�d�    [��]�̃�SUVW�=��@ 3�jS�\$�\$�׋�S�D$PV�J  ��z���@ �-��@ uV�ӋL$Qj ��j ����j �T$RV�  ��u[���vU�����t/����<
t&<t"<�u��r=��w8�<�u����<�u)���u$�D$@��;D$r�_^]�   [���j ��V��_^]3�[���������U��j�h�@ d�    Pd�%    ���hA SV�uW�e�V�E��E�    ������V�>�����������5��@ h'  ����h �@ �E�P�E�   �   �̋T$V�t$���t1��
��t*��A|��Z�� <A|<Z ����+�u+�FFB��uЊ<A|<Z �Ȋ<A|<Z ����+�^����������������@ �D$Pj h  �X�@ ��������U������  VW�=��@ �׋EPj j �\�@ ����u1P���@ j��$  �a�����  �|$�h��@ �L$Q�  ��_��^��]�����������̋D$��tP���@ �U��j�h �@ d�    Pd�%    ���  �hA SVW�E�e���D���Ph  ���@ �u3�3۹6   ������M��8����]��]��4���ǅ���`(@ ǅ ����)@ ��h�����l����E��@ ǅ���   ���@ �������P�U��h�@ jjj��@ �������4���uh�@ �f  ��������   V�5��@ ��\����]���Sf��d���f�E���`����]���j�M�f��f���f�E�����   QW��0�����@�����8�����<��������f�E�f�E�ǅ@���   ���@ ;�u?��A R�  P������h �@ P�[  ������Q�����R�������������D  jdW���@ ;�u>��A P�Y  P������h��@ Q�  ������R�����P��������������  fǅ<��� fǅ>���
 �d�@ P�`�@ P������h��@ Q�  ��S���@ ������R�����P��������]��]�f�]�f�]����$    ��@���Q�U�RWǅ@���   ���@ �����u6��A P�  P������h��@ Q�F  ������R�����P��������j��<���Qh�   h��  V��@ SSh   h��  V��@ ���@ ��8���3�;���   �M�d   ;���   h�   S���@ ;�uB���@ jV���@ V���@ �����h��@ R�E�   �������h�  ���@ �������6   �����󥍍0���QSPh @ h   S���@ ;�tP���@ �����R���@ �U�����BP�U���@ ��4�������h�  ���@ �$���h0u  ���@ ��8���Q�+   ����[@ �3��M�d�    �M��m  _^[��]� �����Q�L�@ �P�@ �T�@ Vj.��A �X�@ j#h�A ��A ��A ��A ������T$���L$QjRhX@ h� j ���@ ��j V�p�@ V�l�@ j ���@ �   ^Y�̡dA ���u!h�A � �@ ��u�dA Ë@���dA ��%��@ �%��@ �%��@ �%��@ �%��@ �%��@ �%��@ U��� V�uW�EP�u�E�P�E�����E�B   �u�u��E  ������t�M�x�E��  ��E�Pj �  YY��_^��jh`�@ �  �e� j j�c  YY�3�@Ëe�M��j�x�@ �;hA u��������̍B�[Í�$    �d$ 3��D$S�����T$��   t�
��8�tτ�tQ��   u��W����V؋
����~����3���������3�3ƃ��� �u% �t�% u��   �u�^_[3�ËB�8�t6��t�8�t'��t���8�t��t�8�t��t��^_�B�[ÍB�^_[ÍB�^_[ÍB�^_[��̋L$W����   VS�ًt$��   �|$u����   �'��������t+��t/��   u����ua��t��������t7��u�D$[^_���   t�������   ��   u����ut�����u�[^�D$_É����t�����~�Ѓ��3��� �t܄�t,��t��  � t��   �uĉ�����  �����   ��3҉��3���t3������u����w����D$[^_�������������U��WVS�M�'�ً}��3����ˋ��u�F�3�:G�wt���ы�[^_��������̋L$WSV��|$��to�q��tU���L$���8�t��t���8�t
��u�^[_3�Ê��8�u�~��a��t(���8�u��A��t�f���8�t��3�^[_���]����G�^[_Ë�^[_�U��QQ�=�A  S�]VW��   �=�A  t	����   3��   F;�s"95�A ~VS�  YY���A �X#ƅ�tv��A �������DJ�tj�E��]��E� X�	�]��E� ��V�5�A �M�jQP�E�PW�5�A �p  �� ��t$;�u�E���M�3��e�����A|��Z�C ~��_^[�������=   s��ă�� �� P�Q�L$��   -   �=   s�+ȋą���@P�h|�@ �\�@ ��thl�@ P�H�@ ��t�t$���t$�x�@ ̡�3A ��t�t$��YVW�A � A 3�;ϋ�s��u?���t�у�;�r��u,h�@ �C  � A �ƿA ;�Ys���t�Ѓ�;�r�3�_^�U��V3�F95<A Wu�u���@ P���@ �} �E�58A �4A uR��3A ��t)��3A ��;��� ��t�С�3A ��;�3A ��3A s�$A �,A ;Ƌ�s���t�Ѓ�;�r�0A �8A ;Ƌ�s���t�Ѓ�;�r�} _^u�u�<A    ����]�j j �t$�2������j j�t$�!������jj j �������jjj �������U��� �EP�E�I   �E�E��|+  �E�EP�u�E�P��  �������@ �I��tQ��+  Y�V��������D$tV��+  Y��^� U��QS�E���E�d�    �d�    �E�]�c��m���[�� XY�$��U��QQSVWd�5    �u��E��c@ j �u�u��u�}q  �E�@����M�Ad�=    �]��;d�    _^[�� U���SVW��E�3�PPP�u��u�u�u�u�3  �� �E�_^[�E���]���D$�H;hA t�D$�H3�@�j P�p�pj �t$ �p�t$ �Y3  �� �U���4S�}#  u��d@ �M�3�@�   �e� �E�e@ �hA �E��E�E�E�E�E�E�E �E��e� �e� �e� �e�m�d�    �E؍E�d�    �E�   �E�EЋE�EԍE�P�E�0��A YY�e� �}� td�    ��]؉d�    �	�E�d�    �E�[��U��QS��E�@;hA t�E�@���M�A3�@�   �E�@��ft�E�@$   3�@�jj�E�p�E�p�E�pj �u�E�p�u�$2  �� �E�x$ u�u�u�����j j j j j �E�Ph#  �������E��]�c�k ��3�@[��U��Q�} SVW�}�w�_�ƉE��u|8���u�2  �MN����9H};H~���u�E�M�E��u�} }ˋE��MF�1�M�;Gw;�v�>2  _��^��[�ËD$�L$��@A �H�@A á@A ��;L$t	�@��u�@�3�ËT$�@A ;�u	�B�@A Ëȃ��� ;�t�ȍA�8 u���1  �B�A�U����hA �e� �M�E��E�E�E@�E�d@ �M��E�d�    �E�E�d�    �uQ�u�1  �ȋE�d�    ������U��SVWUj j h(g@ �u�n  ]_^[��]ËL$�A   �   t�D$�T$��   �SVW�D$Pj�h0g@ d�5    d�%    �D$ �X�p���t.;t$$t(�4v���L$�H�|� uh  �D��@   �T���d�    ��_^[�3�d�    �y0g@ u�Q�R9Qu�   �SQ��A �
SQ��A �M�K�C�kY[� U��� �EVWjY���@ �}��E��E�E��E�P�u��u��u����@ _^�� �D$��A á�A i��C Þ& ��A 3�f��A %�  �U��QQ�E�P��@ �E��M�j  ��*h��� ��!Nb�QP��0  �M��t���V�t$�F�P�)1  ��Yu��F��-��t��+u�F3���0|
��9��0�������t���A�F�݃�-^u�����������̋L$W����   �|$V��   St�����t9��   u�����~Ѓ��3�� �t�G���t!��t�  � t�   �uσ�����������t$��   u	����u\�"�����t=�����t)��   u����u8�˃�t��������t��u�[^�D$_È�D$[^_É����tȺ���~�Ѓ��3��� �t܄�t΄�t*��  � t��   �uĉ�D$[^_�f�3ҋD$�W[^_�f��D$[^_������������U��W�}3�������ك��E���8t3�����_����̋D$S��tR�T$3ۊ\$��   t�
��2�tr��t2��   u��rW����ߋ�����_��t�
��2�t@��u�[Ã�r�
3˿���~����3σ��� �t��J�2�t#2�t��2�t2�t��_�B�[ÍB�_[ÍB�_[ÍB�_[ËL$�ɡ�A |;�}��V�4��A �DA V�m/  YY��^�V�t$��t%�> t V�3#  PVj�B0  jh��@ j�40  ����A ����A |;�|���4��A V��"  PVj�0  jh��@ j��/  ��^Ã=tA u�L3  �t$��1  h�   ��A YY�j`h��@ �  ��   ���.����e��>V���@ �N��A �F�A �V�A �v���  �5 A ��t�� �  �5 A ��£A 3�V�=\�@ ��f�8MZu�H<ȁ9PE  u�A=  t=  t�u��'���   v�3�9��   ��ytv�3�9��   ���E�V�+:  Y��u!�=tA u�U2  j��0  h�   ����YY�}  �u��38  ��}j�����Y�p�@ ��3A ��6  �lA �I6  ��}j����Y�4  ��}j	����Yj�i���Y�E�;�tP����Y�u��E�P�t�@ �t3  �E��E�t�E��j
XP�u�VV��P�k������}�9u�uW�C����`����+�E��	�M�PQ�1  YYËe�}܃}� uW�'����B����M���Ǎe��  �U��SV�u�F���^��   �@��   �t�f ���   �N�����F�F�f �e ����f��Fu"���A t��A uS��9  ��YuV�9  Yf�FWta�F�>�H��N+�I���N~WPS�U-  �E�0���t�������2A �˃������A �@ tjj S�8  ���F�M��3�GW�EPS�-  ���E9}_t�N ��E%�   �	�� �F���^[]��A@t�y t$�Ix��������QP�����YY���u	���U��V����M�E�M�����>�t�} �^]��G@SV����t!� u�D$���L$������C�>�t�|$ �^[�U��$,�����T  �hA ���  3��E��E��E����  S�3Ʉ���  VW����M�G�}� ���  �p  �� |��x������@ ���3������@ j��Y;��E��,  �$�4w@ 3��M���E��E��E��E��EĉE��  �Ã� t;��t-��tHHt����  �M���  �M���  �M���  �MĀ��  �M��  ��*u'���  ���  �@����E���  �M��]��  �E��ˍ��DAЉE��{  �e� �r  ��*u$���  ���  �@����E��R  �M���I  �E��ˍ��DAЉE��4  ��It.��ht ��lt��w�  �M��  �M��
  �M� �  �<6u�4uGG�Mŀ���  ��  <3u�2uGG�e����  ��  <d��  <i��  <o��  <u��  <x��  <X��  �e� ��A �e� ���DA�t���  �u����2����G���  ���  �u��������S  �Ã�g�X  ��e��   ��X��   ��  ��C��   HHt`HHt\���  f�E�0u�M��M����u�������  f�E����  �@��E��D  ��u��A �E��E��E�   �  �E�   �� �M�@�}� �uȉu���   �E�   �4  f�E�0u�M����  f�E����  te�@�P�E�P�6  ��YY�E�}[�E�   �R��ZtX��	t�H�2  �M�@�E�
   �]ľ �  ���3  ���  ��Q�����  �H  �@��E��E�   �EȉE���  ���  ���  �@���t-�H��t&�E�� �M�t�+����E�   �  �e� �  ��A �E�P�   u��gu@�E�   �7�   9E�~�E���   9}�~ �E�]  P�5  ��Y�E�t�E�����}����  ��u����u����  �@��E���P�E�VP�M��HA �}ă���   t�}� uV�TA Y��gu��uV�LA Y�>-u�M�F�u�V�z  Y��  ��i���������   H��   Ht^�������HH���������  �E�'   �EIf�8 t@@��u�+E����  ��u��A �E��E��I�8 t@��u�+E��^  �E�   �M��EĀ�E�   �����E�Q�E�0�E��E�   �����EĀ�E�   ������M���������  �E� ���  �@�t	f�M�f���M���E�   ��  ���  �� ���  t��@t�@����@�����@�@�u�3���@t��|��s�؃� �ڀM��uċ؋�u3��}� }	�E�   ��e���   9E�~�E����u�e� ���  �E��M������t$�E��RPWS�4  ��0��9�]��؋�~M��N�̍��  +�F�E��E��u�t�΀90u��u�M��M��0@�E��}� ��   �]���@t&��t�E�-���t�E�+�	��t�E� �E�   �u�+u�+u���u���  �E�Vj �������u����  �E��M�������Yt��uWVj0�E��������}� tJ�}� ~D�E��]��E��M�3�f�P���  P�2  CYC��Y~-���  P�E����  �]����}� Yu���u��M��E��F���Y�E�t���  �E�Vj �
������}� t�u��  �e� Y���  ����|���_^���  �E�[�C������  ��vq@ �o@ p@ Op@ �p@ �p@ �p@ �q@ U����hA ��t=N�@�uNV�E�P��@ �u�3u��`�@ 3��d�@ 3����@ 3��E�P�l�@ �E�3E�3��5hA u
�hA N�@�^��h  h(�@ �;  �hA �E�xA 3�;�t�M��u�u��YY�M���  3�@Ëe���EHt��@ ǅ����P�@ ��   ��0�@ ǅ������@ ��   �M�h  ������PQ�P�@ ��uhx�@ ������P�Z"  YY��������P�*  Y����<v%��P�  �؍�������1�jht�@ S������S��  Y�D0������v����e��WV��!  �p�@ WV��!  hd�@ V��!  SV��!  WV��!  ������V��!  h  h<�@ V�^1  ��<j��������hXy@ d�    P�D$�l$�l$+�SVW�E��e�P�E��E������E��E�d�    ËM�d�    Y_^[�Q�VC20XC00U���SVWU��]�E�@   ��   �E��E�E��E��C��s�{S�1  ���t{���t}�v�D��tYVU�k3�3�3�3�3���]^�]�t?xH�{S�C������kVS�x������vj�D���������C�D�3�3�3�3�3��Ћ{�v�4�댸    �#�E�H�   �U�kj�S�%�����]�   ]_^[��]�U�L$�)�AP�AP� �����]� j8h8�@ ����3�9|A u8SS3�FVh4�@ h   S�P�@ ��t�5|A ����@ ��xu
�|A    9]~�M�EI8t@;�u�������+�E�|A ����  ;���  ����  3��}ԉ]ȉ]�9] u��A �E SS�u�u3�9]$����   P�u �T�@ ���u�;���  �E�   �6�����������e�ĉE�M���3�@Ëe��4  3ۉ]�M���}ԋu�9]�u�6P��-  Y�E�;��`  �E�   V�u��u�uj�u �T�@ ����   SSV�u��u�u�P�@ ���}�;���   �Et-9]��   ;}��   �u�uV�u��u�u�P�@ �   �E�   �?����������e�ĉE��M���3�@Ëe���3  3ۉ]��M���}ԋu�9]�u�?P� -  Y�E�;�t@�E�   W�u�V�u��u�u�P�@ ��t!SS9]uSS��u�uW�u�S�u �d�@ ��9]�t	�u��  Y9]�t	�u��r  Y���[  �]�3��]�9]u��A �E9] u��A �E �u�1  Y�E����u3��!  ;E ��   SS�MQ�uP�u �1  ���E�;�t�SS�uP�u�u�h�@ ���u�;���   �]������������e���}�VSW�30  ���3�@Ëe��2  3�3��M��;�u#�u���+  Y��;�t1�u�SW��/  ���E�   �u�W�u�u��u�u�h�@ �E�;�u3��&�u�u�E�PW�u �u��_0  �����������u�9]�t#W�<  Y��u�u�u�u�u�u�h�@ ��9]�t	�u��  Y�ƍe��+����U��Q�E�H��   w��A �A�[����V�5�A ���DV�^tj�E��M��E� X�
�E�3��E� @j�5�A �M
�5�A QP�E�Pj�N2  ����u���E
#E��V�5�3A �L5  Y��3A ���3A ��+Ѓ�;�sN�   ;�s���QP�3  ��YYu��V�5�3A �3  ��YYu^Ë�3A +�3A ��3A ������3A �D$���3A ^��t$�u��������YH�h�   �*  ��Y��3A ujXÃ  ��3A ��3A 3��jhh�@ �����E���@ �}���@ s"�e� �E� ��t���3�@Ëe�M���E��������jhx�@ �e����E���@ �}���@ s"�e� �E� ��t���3�@Ëe�M���E����i���Ã=�A V��~jV�*���YY���A �p����u��߃���^��Jx	�
�A�
�R�4  Y�h�  h��@ ������hA �E�3���D�����(�����P�����l�����k�����|�����H����u�����  ���=�A ~jP����YY���A �A��3�;�tG��|�����|����U�[�����V�4  Y��u���t�uV�84  YY�E�E� P�4  Y��u�끋u�>%��  ��`���ƅh��� ��d�����L�����t���ƅ_��� ƅi��� ƅr��� ƅ���� ƅj��� ƅ{��� ƅs�����8���F��Ã=�A ~jP����YY���A �A����t��L������|C��   ��N��   ��   ��*tr��F��   ��It��Luv��s����   �N��6u �F�84u����8�����T��� ��X��� �e��3u�F�82u���T��dtO��itJ��otE��xt@��Xu�9��r����1��ht ��lt��wt���������s�����{������s�����{��������� �������t����u��r��� u�E��$������E�X���P������P���ƅ���� ��{��� u�<St<Cƅ{����uƅ{����>�� ��@�����ntD��ct+��{t&��|����U�8�����V�2  Y��u創l����u���|����U������l�����L�����t��t��� �,  ��o��  �  ��c��  ��d��  ��  ��g~D��it!��n��  ��|�����r��� �
  �5
  jd_��l�����-�c  ƅi����\  ��������l�����-u���������������+u ��t�����|����}���K����؉�l�����}��L��� t��t���]  ~
ǅt���]  �=�A ~jS����YY���A �X����t0��t�����t�����t ��d����F��|�����������؉�l����8�A u|��t�����t�����tl��|����������ؠ�A �F��l����=�A ~jS����YY���A �X����t*��t�����t�����t��d����F��|������J�����뫃�d��� ��   ��et	��E��   ��t�����t�������   �eF��|����������؉�l�����-u�F���+u-��t�����t�����u!�t��������|���������؉�l����=�A ~jS����YY���A �X����t��t�����t�����t��d����F���|������t	WS�h/  YY��d��� ��  ��r��� ��  ��H���� ������P��P�����s���HP�PA ���  ��uǅL���   ��t�����{��� ��  ƅj����  �ǃ�p�  ��t�HH�  ���9�����t8�;�l���t��l�����  ��k�����r��� �<  ��$����E�.  ��{��� ~ƅj����}G�}��0����?^uG��0���ƅ_������D�����u]!]�j X�n����e�܉�D����M���A3�@Ëe��)  j �p"  Y��D�����u	�M���U  ǅ(���   �M����0�����D���j j S�r&  ����@���{uw�?]ur�]G�C �oG<-uK��tG���]t@G:�s�����:�w+��*�������,�������Ë΃����F��,���u�2����h����ȋ���Ã������h����<]u�����  ��P�����@���{u�}��@�������|�����l����t�u��l����%-  YY��L��� t��t�����t�������  ��|����U� �����l��������  ��ctM��su��	|��~�� u9��{��  �ȃ�3�B�������D����9��_���3υ��i  ��@�����r��� �P  ��j��� �5  ��<�������A �DA�t��|����U�a�����=����5�A ��<���P��4���P��,  ��f��4���f�CC��   ��+u+��t���u��t	ƅ�������|����U�����؉�l�����0�b  ��|����U������؉�l�����xtQ��XtLǅd���   ��xt��L��� t��t���u������jo_�  ��|������t�uS�+  YYj0[��   ��|����U�{����؉�l�����L��� t��t�����t���}������jx룈C��P�������F������|������t�uP� +  YY;��T  ��r��� ��  ��H�����@���c��  ��P�����j��� t	f�  �x  �  �p  ƅs�����l�����-u	ƅi������+u+��t���u��t	ƅ�������|����U�����؉�l�����8��� ��  ������ �U  ��   ��x��   ��pt{�=�A ~jS�a���YY���A �X������   ��ou*��8��   ��T�����X���������T�����X����vj j
��X�����T����`  ��T�����X����S�=�A ~VS�����YY���A �X#ƅ�t*��T�����X���������T�����X������p������������������ uB��d����CЙ�T����X�����L��� t��t���u	ƅ�����(��|����U�Q��������|������t�uS�1)  YY������ �������l�����i��� �I  ��T����؋�X����� �ى�T�����X����%  ������ �	  ��   ��xtP��ptK�=�A ~jS�����YY���A �X����t[��ou��8}Q��`����N��`���������`����;�=�A ~VS����YY���A �X#ƅ�t��`������)������������������ uB��d�����`����DЉ�`�����L��� t��t���u	ƅ�����(��|����U�
��������|������t�uS��'  YY������ ������l�����i��� t��`�����Fu��d��� ��d��� ��   ��r��� u>��H�����P�����`�����8��� t��T������X����C���s��� t��f���k����E�u�w��|����U�R����؉�l����F�u;�u9�Ë�A �DA�tF��|����U�!����F�u;�t'���t�uP� '  YY���t7�u��l�����&  YY�%��|�����l�����8����>%u�E�xn�#�����(���u��D�����   Y��H�����l����u��u8�k���u���������M��������������������̋L$��   t$�����tN��   u�    ��$    ��$    �����~Ѓ��3�� �t�A���t2��t$�  � t�   �t�͍A��L$+�ÍA��L$+�ÍA��L$+�ÍA��L$+��V�t$��t-�=�2A Vu�s'  ��YVt
P�'  YY^�j �5�2A �L�@ ^�������������̋T$�L$��   u<�:u.
�t&:au%
�t��:Au
�t:au����
�uҋ�3�Ð��������   t���:u��
�t���   t�f���:u�
�t�:au�
�t���눋F��tD�P�: t<�O;�t��QR�X�����YYu"�t�t�D$� �t�t	�t�u3��3�@Ë �8csm�t3�Ã%�A  ��  jh��@ �����]�s�u���A �e� �};utd���~;w|��  �����Oȋ1�u��E�   �y t�sh  S�O�t��  �e� ��E��r���Ëe�e� �}�]�u��u�뗃M���   ;ut�  �s�I���Ë]�u�=�A  ~��A �jh��@ ������E��t�H�I��t�e� Q�p�V����M��������3�8E��Ëe���  V���ƃy |�Q�I�42���^�j@h��@ �����ً}�u�]��e� �G��E��v�E�P����YY�Eġ�A �E���A �E��5�A �E��A �e� �E�   �u�uS�uW��������E��e� �   �E� �E�E�8csm�u1�E�xu(�E�x �t�E�x!�u�E�x �E�   t�E�    �E�Ëe�M�A�EЋ}�G�E؋Q�U�3҉U�;Qs$�4��]ԍ4��^;�~=;F8�C�E؋UЋE�PQ3�VW��������u��u��u�M���   �E������B먋}�u�EȉG��u�����Y�E���A �E���A �>csm�u>�~u8�F= �t=!�u'�}� u!�}� t�v�Z���Y��t����PV�����YY�jh��@ �������E���]�H���I  �y �?  �H��u
�@��.  � ��x�|9�e� j�s�t5�.  YY����   jW�.  YY����   �C��N�������   �tF��-  YY����   jW��-  YY����   �v�sW�.  ���~��   �����   릃~ u3�-  YY��t}jW�-  YY��to�v�N�C�7���PW�-  ���Z�U-  YY��tJjW�c-  YY��t<�v�q-  Y��t/�C�N�tj�����P�vW�$���������P�vW�������  �M�������3�@Ëe��  U���tS�u���r���YY�} �uuV��u������7�u�uV�����Gh   �u@�u�F�u�KV�u������(��tVP�a���]�U��QQ�E�8  ���   �=�A  t�u$�u �u�u�u�uP�$�������u~V�uW�E�P�E�PV�u �u�{������E���;E�sVS;7|B;w=�G�O����H��t�y u%�u$�u�u �X��u3��u�u�u������u���E��E���;E�r�[_^��U���$�E�@����E� �E�|�M;A|�  S�]�;csm�VW��  �{� �uy�C;�t=!�uk�{ ue��A ���\  ��A jV�u�E�E��K+  ��YYu�:  �>csm��1  �E�xu�@;�t=!�u�E�x u�	  �]�;csm��   �{��   �C;�t=!���   �u�E�P�E�PV�u �u�����M��;M��E���   ��u�90��   ;p|�H�ɋp�M�~o�K�I�Q�	�ɉU��M�~$�E��8�s�}��������Yu�M�E�9E�ߋE��M���}� ��(�u$�}��u �M��u�u�uS�ދu�K����]�����E�M��;M��E��_����} t
jS����YY_^[�Ë]�} u �u$�u �u��u�u�u�uS�\����� ���   U��V�u�W%���� �;�t�   �E�@ft�~ to�} uij�V�u�u�d������V�~ tP�8csm�u,9xv'�H�I��t�U$R�u �uV�u�u�uP�у� ��u �u�u$V�u�u�uP�v����� 3�@_^]�jh��@ ������A ��t�e� ���3�@Ëe�M���,  jh��@ �}�����A ��t�e� ���3�@Ëe�M��������������U���SQ�E���E��EU�u�M�m��
���VW��_^��]�MU���   u�   Q�����]Y[�� V�t$��8csm�u�xu�@= �t=!�u�'�����A ��tP�(  ��Yt	V��A �3�^� h��@ �H�@ ��A 3���5�A �H�@ �������SV�D$�u�L$�D$3���؋D$����A�ȋ\$�T$�D$���������u�����d$�ȋD$���r;T$wr;D$vN3ҋ�^[� U��Q�M���   v^f�e� W3��}�f������=\ A  �E
�M_u3���j�5X A �E��5d!A Pj�E
Pj�  ����t�f�}� u��E�t�3�@�Ã=�A ~jQ����YY�á�A �H�����������̋D$�L$ȋL$u	�D$��� S��؋D$�d$؋D$���[� ������������W�|$�n��$    ���L$W��   t�����t=��   u�������~Ѓ��3�� �t�A���t#��t�  � t�   �t�͍y���y���y���y��L$��   t�����tf�����   u���������~�Ѓ��3��� �t��t4��t'��  � t��   �t�ǉ�D$_�f��D$�G _�f��D$_È�D$_�U��$d�����  ���  ;�2A �hA SV���  W��  �������2A �������D0��]��s  3�9��  �}��}�u3��p  � tjWWQ�\-  �����@���   9��  ���  �E����  ��   �M�+��  �E�;��  s%�U��E��A��
u�E�� @G�]��@G��   |Ӌ��E�+�j �E�PW�E�P��40�T�@ ��t�E�E�;�|!�E�+��  3�;��  r�����@ ���  3��E�;���   9��  tYjX9��  u@��A �}W�M�Q���  ���  �0�T�@ ��t�E����  �E�����@ ���  ����  ��+  Y�@��D0@t���  �8�������A    �=�A �+E���%�A  ��A 	   ������  _^[�߿���Ŝ  ��U��$t�����  �hA ���   SV���   3�W3�;ŘA t@��r����;��A �  �tA ����   ;�u�=�A ��   ���   ��   h  �E�PR���   �P�@ ��u�E�hx�@ P����YY�}���P�R���@��<Yv"��P�C������E���;j�ht�@ W������W�#������A �������DY��Y���������h��@ S����WS�!���hp�@ S�������A S�
���h  h<�@ S�  ��,�(R���   P���A �6����YP�6j��D�@ P�T�@ ��t������   �k���_^[�Ō   �átA ��t��u*�=�A u!h�   �h�����A ��Yt��h�   �R���Y�U��U��A S�0A V9t�4@���4�0A ;�r�@��0A ;�s9t3Ʌ��!  �Y���  ��u�a 3�@�  ����   ��A �E�E��A �A����   ��A ��A �;�}�4@�4�8A +Ѓ& ��Ju��	���  ��5�A u��A �   �v���  �u��A �   �b���  �u��A �   �N���  �u��A �   �:���  �u��A �   �&���  �u��A �   ����  �u
��A �   �5�A j��Y�5�A ��a P�ӋEY��A ����	�u�@�@ ^[]�VW3�9=�3A u�5(  �5�3A ��u���@ �< w��t.��t$<"u	3Ʌ�������P�Q)  ��YtFF��< wF���u�_��^�S3�9�3A VWu��'  �5lA 3�;�u�0<=tGV�O���Y�t�:�u��   P��  ��;�Y�=A u����X�5lA U�*V������E�>=YtU�  ;�Y�t7VP����YY���8u��5lA �n����lA ���3A    3�Y]_^[��5A �I����A �����U��QS�]3�9UW����   t	�M�E�9�8"u3Ʌ���@�ѱ"�-���t��G���@��a A t���t��G@�ɋ]t2��u��� t��	u���t�G� �e� �8 ��   ��� t��	u@��H��8 ��   �} t	�M�E�9�3�C3��@B�8\t��8"u&��u�}� t�H�9"u���3�3�9M����M����t��t�\G�Ju���tH�}� u
�� t=��	t8��t.��t����a A t�G@���G�����a A t@��@�h�����t� G��]�!����E��t�  �_[��U��QQSVW3�9=�3A u�%  h  ��A VW��A  �P�@ ��3A ;ǉ5,A t�8 ��u�ލE�PW�u�3ɋ��;����u��E����P�  ������u����%�E�P�>W�u����
����E�HY�A Y�=A 3�_^[��QQ��A SUVW�=0�@ 3�3�;�j]u-�׋�;�t��A    ����@ ��xu	�ţ�A ���A ��u};�u�׋�;�tyf9��t�f9u��f9u�=d�@ SSS+�S��@PVSS�D$4�׋�;�t2U��  ;�Y�D$t#SSUP�t$$VSS�ׅ�u�t$�y���Y�\$�\$V�4�@ ���P;�t;�t3��D�8�@ ��;�t�8t
@8u�@8u�+�@��U�_  ��;�Yu3��UVW�f%  ��V�<�@ ��_^][YYÃ�Dh   �,  ��Yu����  ��2A ��2A     ��   ����@ �@
��2A ����   ;�r�SVW�D$P�t�@ f�|$> ��   �D$@����   �0U�h�   ;��.|��95�2A }R��2A h   �  ��Yt8��2A  ���   ����@ �@
�����   ;�r��95�2A |���5�2A 3���~F����t6�M ��t.��uP�(�@ ��t�������2A �σ��ȋ��M �HGE��;�|�]3ۡ�2A �4؃>�uM���F�uj�X�
��H������P�D�@ �����tW�(�@ ��t%�   ���>u�N@���u
�N��N�C��|��5�2A �,�@ _^3�[��DÃ=�A u�=A r3�@�jX�3�9D$j ��h   P� �@ ����2A t*���������2A uh�  �S  ��Yu�5�2A �$�@ 3��3�@ËD$;�2A SVWse���������<��2A ����D1tHP��&  ���YtC�t$j �t$P��@ �؃��u���@ �3���t	P�!  Y���D0� �����%�A  ��A 	   ���_^[���A h   �  ��Y�L$�At�I�A   ��I�A�A�A   �A�a �ËD$;�2A r3�Ë������2A ���D���@á�2A ��Vj^u�   �;�}�ƣ�2A jP�&  ��YY��"A ujV�5�2A ��%  ��YY��"A ujX^�3ҹ�A ���"A ��� ����HA |�3ҹ�A �������2A ��������t��u�	��� B��8A |�3�^��f'  �=4A  t��%  Ã=�2A V�t$u;5�"A wV�  ��Yu#��uF�=�2A t�����Vj �5�2A ��@ ^Ã|$�w"�t$������Yu9D$t�t$��&  ��Yu�3���5@ A �t$�����YY�U��EV3�;�u3��R95�A uf�Mf��� w2�3�@�8�MQV�5�A �uPj�EPV�5�A �d�@ ;�t9ut��A *   ���^]���V�D$�u(�L$�D$3���؋D$������d$�ȋ��d$��G�ȋ\$�T$�D$���������u�����d$�ȋD$���r;T$wr;D$v	N+D$T$3�+D$T$���؃� �ʋӋًȋ�^� U���S3�9�A VWumh`�@ �L�@ ��;���   �5H�@ hT�@ W�օ���A t|hD�@ W��h0�@ W��A �փ=�A ��A uh�@ W�օ���A th��@ W�֣�A ��A ��t<�Ѕ�t�M�Qj�M�QjP��A ��t�E�u�=A r
�M �)3��5�M���A ��t�Ћ؅�t��A ��tS�Ћ��u�u�uS��A _^[��U��� SV�u�^��ud�   �E�E�H;ىM�r;Xs3���  W�~���u3�@��  3҉U�Ë���t;��E  �x t�EB��;�v��} t�F�;E��"  ;��  ��A ���� ���3���~9<��A ��   F;�|�j�E�PS��@ ���`  �}�   �S  �E��tV�M�f�9MZ�?  �A<��8PE  �.  f�x�"  +�f�x �H�L�  �A;�r�Q�;�s�A'�uwjh0 A ��@ ���������A �ɋ�~���A 98tJ������u-j[;���3҅�|���A �0B;Ӊ8��~��}A��A j h0 A ��@ ����3�����������@ jh0 A �Ӆ��z���9<��A t.��A �p���|9<��A tNy��}��}@��A �p��t3Ʌ�|���A �A;Ή8��~�j h0 A ���������_^[����������̋T$�L$��tO3��D$W����r1�ك�t+ш����u������������ʃ���t��t
�����u��D$_ËD$�U����hA j�E��E�Ph  �u�E� ��@ ��u����
�E�P膺��Y�M��N�����j8hp�@ ������hA �E�3��}̉}��E��]��}ċE;E�s  �M�QP�5 �@ �օ�t �}�u�E�P�u�օ�t�}�u�E�   9}�t���t����u�����Y��F�u���u�9}�uWWS�uj�u�T�@ ���u�;�tX�}��6������G����e�܉]��6PWS�������M���3�@Ëe���   3�3ۃM���u�;�uVj�;  YY��;�u3��   �E�   VS�u��uj�u�T�@ ����   9}t WW�u�uVSW�u�d�@ ��tf�E�E��^9}�uWWWWVSW�u�d�@ ��;�tCVj��  YY�E�;�t2WWVPVSW�u�d�@ ;�u�u��e���Y�}���}��t
�M���]�9}�tS�D���Y�E̍e��M�艭���T����U���LSVWjX�#�����j�E�PV��@ ��tw�]܍E�P���@ �M���A �y���#�+���N����������;��M�r@��t\�]��   j�E�P�u���@ ��t �E�E��]�t��E��E؉E�t3�@�D;�s3��<;�s�u�jS�u��u����@ ��A ��}�H���%  �M�Q@P�u��u����@ �e�_^[��jh��@ �)���3�954 A u5�E�P3�GWh4�@ W���@ ��t�=4 A ����@ ��xu
�4 A    �4 A ����   ;���   ����   �u܉u�9uu��A �EVV�u�u3�9u ����   P�u�T�@ ���}؅���   �e� �?�Ã����蒯���e��u�Sj V��������M���3�@Ëe��8���3��M���}؅�uWj�  YY����tg�E�   WV�u�uj�u�T�@ ��t�uPV�u���@ �E܃}� tV����Y�E��n�];�u��A �}��u�=�A S����Y���u3��D;�tj j �MQ�uPW�����������t݉u�u�u�u�uS�`�@ ����tV����Y�Ǎe������S�\$��UWu�t$����Y�D  V�t$��uS�i���Y�,  �=�2A ��   3������   S��  ���Y��   ;5�"A wHVSU�  ����t���1V�  ����Yt(�C�H;�r��PSW�E  S�  ��SU�  ����u<��uF�����Vj �5�2A ��@ ����t�C�H;�r��PSW��  SU�g  ����u��uF�����VSj �5�2A ���@ ����u�=@ A  tV�  ��Y�����8���63����w��uFVSj �5�2A ���@ ��u�=@ A  tV�^  ��Yu�3�^_][Ã=�2A Vu�t$V�  ��Yt�F���	^�V��t$j �5�2A ���@ ^�V�t$�F����   �@��   �t�� �F�   ��f��Fu	V�S���Y��F��v�v�v��  �����Fto���tj�V�u7�N���Wt�����<��2A ���<����A �O�ႀ��_u	��    �V�~   u�N��t��u�F   �H�F�A�^��������	F�f ���^�S�\$���VtA�t$�F�u��y2�u.�~ uV����Y�;Fu	�~ u@���F@�t8t@����^[È�F�F�����F��%�   ��=�A ~j�t$����YYËD$��A �A���U��SV�u3�;�t9]t�:�u�E;�tf�3�^[]�9�A u�M;�tf��f�3�@���A ���DA�tM��A ��~*9E|(3�9]��Q�uPVj	�5�A �T�@ ����A u�9Er8^u���A *   ����3�9]��P�ujVj	�5�A �T�@ ���y�����h@  j �5�2A ��@ ����"A uËL$�%�"A  �%�"A  ��"A 3���"A ��"A    @á�"A ����"A ����T$+P��   r	��;�r�3��U����M�AV�uW��+y�������i�  ��D  �M��I���M���  S�1��U�V��U��U����]ut��J��?vj?Z�K;KuB�� �   �s����L��!\�D�	u#�M!��J���L��!���   �	u�M!Y�]�S�[�M�M�Z�U�Z�R�S�M�����J��?vj?Z�]����]���   +u��]���j?�uK^;�v��M�����J;։M�v��;�t^�M�q;qu;�� �   �s������!t�D�Lu!�M!1��K�����!���   �Lu�M!q�M�q�I�N�M�q�I�N�u��]�}� u;���   �M��ыY�N�^�q�N�q�N;Nu`�L�M���� �Ls%�} u�ʻ   ���M	�   �����D�D	�)�} u�J�   ���M	Y�J�   ��ꍄ��   	�E���D0��E����   ��"A ����   ��"A �5�@ h @  ��H� �  SQ�֋�"A ��"A �   ���	P��"A �@��"A ����    ��"A �@�HC��"A �H�yC u	�`���"A �x�uiSj �p�֡�"A �pj �5�2A �L�@ ��"A ��"A �����ȡ�"A +ȍL�Q�HQP�,  �E����"A ;�"A v�m��"A ��"A �E��"A �=�"A [_^�á�"A ��"A W3�;�u4�D�P��P�5�"A W�5�2A ���@ ;�u3�_Ã�"A ��"A ��"A ��"A Vh�A  j�5�2A ���4���@ ;ǉFu3��Cjh    h   W���@ ;ǉFu�vW�5�2A �L�@ �ЃN��>�~��"A �F����^_�U��QQ�M�ASV�qW3����C��}���i�  ��0D  j?�E�Z�@�@��Ju�j��h   ��yh �  W���@ ��u����   �� p  ;��U�wC��+����GA�H�����  ����  ��������@��  �Pǀ�  �     IuˋU��E��  �O�H�A�J�H�A�d�D 3�G����   �FC�������E�NCu	x�   �������!P��_^[��U����M�ASV�uW�}��+Q������i�  ��D  �M�O����I;�|9���M�]��U  ���E  �;��;  �M���I��?�M�vj?Y�M��_;_uC�� �   �s��M��L��!\�D�	u&�M!������M��L��!���   �	u�M!Y�O�_�Y�O��y�M+�M��}� ��   �}��M��O��?�L1�vj?_�]���]�[�Y�]�Y�K�Y�K�Y;YuW�L�M���� �Ls�} u�ϻ   ���M	�D�D��� �} u�O�   ���M	Y����   �O�   ���	�U�M��D2���L���U�F�B��D2��<  3��8  �/  �])u�N�K��\3��u��N��?�]�K�vj?^�E���   �u���N��?vj?^�O;OuB�� �   �s����t��!\�D�u#�M!��N���L��!���   �	u�M!Y�]�O�w�q�w�O�q�uu��u��N��?vj?^�M��y�K�{�Y�K�Y�K;KuW�L�M���� �Ls�} u�ο   ���M	9�D�D��� �} u�N�   ���M	y����   �N�   ���	�E��D�3�@_^[��U����M��"A ��"A �����S�M���V��WI�� �<��}�}�����M���������3���E���"A �؉u�;���K�;#M�#��u��;]��]r�;]�u$����K�;#M�#��u
��;؉]r�;���   ��"A �C�����U�t����   �|�D#M�#��u6���   #U��e� �HD�1#u�֋u�u���   #U��E����9#��t�U���i�  ��D  �M�L�D3�#�um����   #M�j _�^�{ u���];]�r�;]�u&���	�{ u
��;؉]r�;�u�����؅ۉ]tS����Y�K��C�8��$���3��z  ��G��}��M�T��
+M�����N��?�M�~j?^;��  �J;Ju\�� �   �}&����M��|8�Ӊ]�#\�D�\�D�u3�M�]!�,�O���M�����   �|8��!��]�u�]�M�!K��]�}� �J�z�y�J�z�y��   �M��y�J�z�Q�J�Q�J;Ju^�L�M���� �L}#�} u�   �����	;�ο   ���M�	|�D�)�} u�N�   ���	{�M�����   �N�   ���	7�M���t�
�L���M��u�эN�
�L2��u��ɍy�>u;�"A u�M�;�"A u�%�"A  �M���B_^[��V�t$3��t$F���@ ��t3���^�V�t$3��t$F���@ ��t3���^�V�t$3�F���@ ��t3���^����������������U��WV�u�M�}�����;�v;��|  ��   u������r)��$�,�@ �Ǻ   ��r����$�@�@ �$�<�@ ��$���@ �P�@ |�@ ��@ #ъ��F�G�F���G������r���$�,�@ �I #ъ��F���G������r���$�,�@ �#ъ���������r���$�,�@ �I #�@ �@ �@  �@ ��@ ��@ ��@ ��@ �D��D��D��D��D��D��D���D���D��D��D���D���D���D����    ���$�,�@ ��<�@ D�@ P�@ d�@ �E^_�Ð���E^_�Ð���F�G�E^_�ÍI ���F�G�F�G�E^_�Ð�t1��|9���   u$������r����$���@ �����$�x�@ �I �Ǻ   ��r��+��$���@ �$���@ ���@  �@ (�@ �F#шG��������r�����$���@ �I �F#шG�F���G������r�����$���@ ��F#шG�F�G�F���G�������V�������$���@ �I |�@ ��@ ��@ ��@ ��@ ��@ ��@ ��@ �D��D��D��D��D��D��D��D��D��D��D��D��D��D���    ���$���@ ����@ ��@ ��@ �@ �E^_�Ð�F�G�E^_�ÍI �F�G�F�G�E^_�Ð�F�G�F�G�F�G�E^_��j
�t���j�T  YYj蕝���-�  t"��t��tHt3�ø  ø  ø  ø  �Wj@3�Y�` A �3��d!A �\ A �X A �p!A ���_�U���  �hA �E�V�E�P�5d!A � �@ ���   �  3�������@;�r�E��ƅ���� t6S�U�W�
��;�w+�A�����������    �˃��B�B��u�_[j �5X A �������5d!A PV������Pj����j �5d!A ������VPV������PV�5X A ����j �5d!A ������VPV������Ph   �5X A �ڳ����\3�f��E������t��a A ���������!A ���t��a A  ��������ƀ�!A  @;�r��D3���Ar��Zw��a A �Ȁ� ���!A ���ar��zw��a A  �Ȁ� ��ƀ�!A  @;�r��M�^�X�����U����hA SV�u3ۃ���E�W�8 A u�8 A    �|�@ �+���u�8 A    ���@ ����u��A �8 A    �E��;5d!A �c  ;��Q  3�3�9�hA tg��0B=�   r�E�PV� �@ ���  j@3�Y�` A �3�G9}�5d!A �X A ��   �}� ��   �M�����   �A����   j@3�Y�` A �R���]䪍�xA ����)�V��t&����;�w�U䊒`A �a A @;�v�FF���u��E���}�r��E�d!A �\ A    �������lA �p!A ���X A ��\��a A @;�v�AA�y� �K����ǀ�a A @=�   r���{����X A �=\ A ��\ A 3��p!A ����98 A t�~�������3������M�_^[�r����Ã=�3A  uj��
���Y��3A    3�ËD$��A 3�;�XA tA��-r��r��$w��A    Ë�\A ��A �=�   r=�   ��A    v
��A    �U��QQ�E;�2A VWsr���������<��2A ����D1tU�M�M��MP�M��Z  ���YtD�u�M�Q�u�P��@ ����E�u���@ ��t	P�1���Y�"��D0� ��E��U���%�A  ��A 	   ������_^���D$�L$��a A u�|$ t��A �A#D$�3���u�3�@�jj �t$���������U��WV�u�M�}�����;�v;��|  ��   u������r)��$���@ �Ǻ   ��r����$���@ �$���@ ��$�@�@ ���@ ��@  �@ #ъ��F�G�F���G������r���$���@ �I #ъ��F���G������r���$���@ �#ъ���������r���$���@ �I ��@ ��@ ��@ ��@ x�@ p�@ h�@ `�@ �D��D��D��D��D��D��D���D���D��D��D���D���D���D����    ���$���@ ����@ ��@ ��@ ��@ �E^_�Ð���E^_�Ð���F�G�E^_�ÍI ���F�G�F�G�E^_�Ð�t1��|9���   u$������r����$�H�@ �����$���@ �I �Ǻ   ��r��+��$�L�@ �$�H�@ �\�@ ��@ ��@ �F#шG��������r�����$�H�@ �I �F#шG�F���G������r�����$�H�@ ��F#шG�F�G�F���G�������V�������$�H�@ �I ��@ �@ �@ �@ �@ $�@ ,�@ ?�@ �D��D��D��D��D��D��D��D��D��D��D��D��D��D���    ���$�H�@ ��X�@ `�@ p�@ ��@ �E^_�Ð�F�G�E^_�ÍI �F�G�F�G�E^_�Ð�F�G�F�G�F�G�E^_�ËL$;�2A VWsU������<��2A �������@t7�8�t2�=�A u3�+�tItIuPj��Pj��Pj��x�@ ���3���%�A  ��A 	   ���_^ËD$;�2A s�������2A �����@t� Ã%�A  ��A 	   ����SV�t$�t$��W��uF3����w9�=�2A u�����;�"A wS���������Yu+Vj�5�2A ��@ ����u"�=@ A  tV�  ��Yu��Sj W��������_^[�VWj^3�95�2A ~D��"A ����t/�@�tP�  ���YtG��|��"A �4�������"A �$� YF;5�2A |���_^�SV�t$�F�Ȁ�3ۀ�u:f�t4�FW�>+���~'WP�v�Q�����;�u�F��y����F��N ���_�F�f �^��[�V�t$��u	V�,   Y^�V������Yt���^��F@t�v�K  Y���^�3�^�SVW3�3�3�95�2A ~M��"A ����t8�H���t0�|$uP�������YtC��|$ u��tP�x������Yu�F;5�2A |��|$��t��_^[�j����Y�j�z���Yá< A ��t�t$�Ѕ�Yt3�@�3��U���SV�u;5�2A W��  �����<��2A �����ƊP����  �e� �} �]��tb��u]��Ht"�x
t��D0�M���K�E�   �D0
j �E�P�u�Q�40�t�@ ��u0���@ jY;�u��A �6  ��mu3��7  P����Y�(  �E��E��D1���   ��t�;
u���D0��	��D0� ��E�M��;��E��M���   �E�� <��   <t�C�E��   I9M�s�E�@�8
u�E��Y�E��n�E�j �E�Pj�E�P��40�t�@ ��u
���@ ��uF�}� t@��D0Ht�E�<
t���D1�(;]u�}�
u�
�jj��u�,������}�
t�C�M�9M��L������D0@u�t0�+]�]�E���%�A  ��A 	   ���_^[�Ë�A �0A V9Pt�4I���4�0A ;�r�I��0A ;�^s9Pt3��U��VW�}��HHtXHHtF��tA��t<��t*��tHt�����   �5L A �L A �3�5H A �H A �&�5P A �P A ����h������0��5D A �D A ����   ��uj�ŏ��SjY;�t
��t��u&��A �%�A  ;�uD��A �U��A �   ��];�u(��A ��A �;�}�@��8A +ȃ" ��Iu���  ;�u�5�A j��YY�W�փ�Yt��u����A u�E��A [3�_^]�V�t$�FW����@t����:��t4V�_���V���9  �v�~   ����}�����F��tP�+����f Y�ǃf _^ËD$;�2A s=�������2A �Ѓ��D�t%P�����YP���@ ��u���@ �3���t��A ��A 	   ����SUVW�|$;=�2A ��   �����������2A ����D0tiW�������Yt<��t��uj�t���j���k���;�YYtW�_���YP���@ ��u
���@ ���3�W�������Y�D0 t	U�5���Y�3���%�A  ��A 	   ���_^][�V�t$�F��t�t�v�����f�f��3�Y��F�F^���%$�@ �%X�@ V�t$��tV�A���@P�������YYtVP�M���YY^�3�^�jh��@ 荣��3ۉ]ࡈA ;�u(�E��8��   �
��A|
��Z�� �
B8u��   j�5�A SSj��uh   P蒤���� �E�;���   �]�������=����e��u��3�@Ëe������3�3��M��;�u�u��9���Y���E�   ;�t3j�5�A �u�Vj��uh   �5�A ������ ��tV�u�d���YY9]�tV�¸��Y�E�e��ڢ���jh��@ 蒢��3ۉ]ࡈA ;�u(�E��8��   �
��a|
��z�� �
B8u��   j�5�A SSj��uh   P藣���� �E�;���   �]�������B����e��u��3�@Ëe������3�3��M��;�u�u��>���Y���E�   ;�t3j�5�A �u�Vj��uh   �5�A �"����� ��tV�u�i���YY9]�tV�Ƿ��Y�E�e��ߡ������������������U��WVS�u�}����
�t2����'��8�t�,A<ɀ� �A��,A<ɀ� �A8�t�����[^_���̸d�@ ���������̸��@ ���������̸�@ ����������̸T�@ ���������̸��@ �܋�������̸��@ �̋�������̸D�@ 鼋�������̸��@ 鬋�������̸��@ 霋�������̸4�@ 錋�������̸��@ �|��������̸��@ �l��������̸$�@ �\��������̸t�@ �L��������̸��@ �<��������̸�@ �,��������̸d�@ ���������̸��@ ���������̸l A ����������̸� A ���������̸A �܊�������̸\A �̊�������̸�A 鼊��                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                      & �  	 � � � � � � � | j Z L 8 �     0 B R h t � � � � � � � z n d T D 4 (    �  � � � � � � � � r b R > 0   � � � � �	 � � � � � � �	 t b T F 8 *  �
 �
 �
 �
 �
 �
 h
 \
 L
 6
 �	 �	 �  
 
 �	 �	 �	 x	     � � �       > R b t � � � � � .     s  �  �  �	  �  ��  �  �  �  �  �  �  �  �  �  �4  �  �  �  �  �t  �  �  �    X	                                     :%hu    %.265s  %s  UDPMAP  BIND    CONNECT UNKNOWN %u.%u.%u.%u %s
 rcpt to:    bcc:    cc:     to:     %u.%u.%u.%u/%u  SeDebugPrivilege    &Yes    ##&Remember my answer, and do not ask me again for this application.    Grant Access    %s%s    mcafe   e personal firewall plus alert  Windows Security Alert  &Unblock    Sygate Personal Firewall Pro    winroute.exe    wrctrl.exe  %s%s erstellen  Un processus cache requiert une connexion reseau.   Un proceso oculto solicita acceso a la red  Ein versteckter Prozess verlangt Netzwerkzugriff.   Hidden Process Requests Network Access          Creer une regle pour    Crear regla para    Regel fur   Avertissement : Les composants ont change   Advertencia: Los componentes han cambiado   Create rule for     Warnung: Einige Komponenten wurden verandert.   Warning: Components Have Changed    :       &Remember this answer the next time I use this program. PermissionDlg   AllocateAndGetTcpExTableFromStack   iphlpapi.dll    5244E14B~8F6D~E9FA~9A78~    4E52E11D78CA    SharedAccess        SYSTEM\CurrentControlSet\Services\SharedAccess\Parameters\FirewallPolicy\StandardProfile\AuthorizedApplications\List    Update  Microsoft   :*:Ena  bled:   ##Software\Microsoft    \Windows\CurrentVersion\Run KAVPersonal50   wuauserv    navaps  vc  ##Symant    ec Core LC  SAVScan kavsvc  wscsvc  wininet.dll ws2_32.dll  dnsapi.dll  Memory Allocation Failed    accept(): %s    Accepting connections [%u/%u]   listen(): %s    bind(): %s  socket()    G%y%m%d%H%M%S.%. %p %E %U %C:%c %R:%r %O %I %h %T   loop#upseek#org     ����[]@ _]@ CorExitProcess  mscoree.dll l�@ Ac@ csm�               �        
   :   ����|m@ �m@            EEE50 P     (8PX 700WP        `h````  ppxxxx          ( n u l l )     (null)  Microsoft Visual C++ Runtime Library    Program:    

  ... <program name unknown>  A buffer overrun has been detected which has corrupted the program's
internal state.  The program cannot safely continue execution and must
now be terminated.
 Buffer overrun detected!        A security error of unknown cause has been detected which has
corrupted the program's internal state.  The program cannot safely
continue execution and must now be terminated.
    Unknown security failure detected!  �����w@ �w@     ����R}@ V}@ ����O{@ S{@ ����|@ !|@                                                                                                                                                                                                                                                                                       ( ( ( ( (                                     H                � � � � � � � � � �        � � � � � �                           � � � � � �                                                                                                                                                                                                                                                                                                               h ( ( ( (                                     H                � � � � � � � � � �        ������      ������                                                                      H                                      ����|@ �@     �����@ �@     ����Æ@ ǆ@     ����    ��@     ��@ Ɛ@ ����A�@ J�@     ����    ��@     �@ :�@ ������@ ��@     ����k�@ o�@     ������@ ��@ Illegal byte sequence   Directory not empty Function not implemented    No locks available  Filename too long   Resource deadlock avoided   Result too large    Domain error    Broken pipe Too many links  Read-only file system   Invalid seek    No space left on device File too large  Inappropriate I/O control operation Too many open files Too many open files in system   Invalid argument    Is a directory  Not a directory No such device  Improper link   File exists Resource device Unknown error   Bad address Permission denied   Not enough space    Resource temporarily unavailable    No child processes  Bad file descriptor Exec format error   Arg list too long   No such device or address   Input/output error  Interrupted function call   No such process No such file or directory   Operation not permitted No error    runtime error   
  TLOSS error
   SING error
    DOMAIN error
  R6029
- This application cannot run using the active version of the Microsoft .NET Runtime
Please contact the application's support team for more information.
   R6028
- unable to initialize heap
    R6027
- not enough space for lowio initialization
    R6026
- not enough space for stdio initialization
    R6025
- pure virtual function call
   R6024
- not enough space for _onexit/atexit table
    R6019
- unable to open console device
    R6018
- unexpected heap error
    R6017
- unexpected multithread lock error
    R6016
- not enough space for thread data
 
This application has requested the Runtime to terminate it in an unusual way.
Please contact the application's support team for more information.
   R6009
- not enough space for environment
 R6008
- not enough space for arguments
   R6002
- floating point not loaded
    Runtime Error!

Program:    GetProcessWindowStation GetUserObjectInformationA   GetLastActivePopup  GetActiveWindow MessageBoxA user32.dll      ������@ ��@     ������@ ��@     ������@ ��@     ������@ ��@     H                                                           hA ��@    RSDST�4��H+@�ߘN4��\   w:\work\vcprj\prj\socks5\Release\socks5.pdb pA         ����        <�@                T�@             pA \�@ d  e  0g  Xy  ��  ��  ��  ��   �  �   �  0�  @�  P�  `�  p�  ��  ��  ��  ��  ��  ��  ��  ��   �  �   �                     @A     ����              ��@             �@ ����    ����                �+@               @�@  �   0�@    P�@         ����    ����                t.@               ��@  �   ��@    ��@         ����    ����                G/@               ��@  �   ��@    ��@         ����    ����                �0@               0�@  �    �@    @�@         ����    ����                �1@               ��@  �   p�@    ��@         ����    ����                �2@               ��@  �   ��@    ��@         ����    ����                5@                �@  �   �@    0�@         ����    ����                �6@               p�@  �   `�@    ��@         ����    ����                �7@               ��@  �   ��@    ��@         ����    ����                R9@               �@  �    �@     �@         ����    ����                �:@               `�@  �   P�@    p�@         ����    ����                "=@               ��@  �   ��@    ��@         ����    ����                �=@                �@  �   ��@    �@         ����    ����                �>@               P�@  �   @�@    `�@         ����    ����                r?@               ��@  �   ��@    ��@         ����    ����                hC@               ��@  �   ��@     �@         ����    ����                E@               @�@  �   0�@    P�@         ����    ����                wF@               ��@  �   ��@    ��@             LA     ����             ��@             ��@ ����                    ����                �T@             �T@             $ A              4 A  �    A    D A         ����    ����                SU@               � A  �   � A    � A         ����    ����                �U@               � A  �   � A    � A         ����    ����                �V@               8A  �   (A    HA         ����    ����                �[@               �A  �   xA    �A                     � H�              &	  �              j	 $�              � ��              � ��              4	 ��                      & �  	 � � � � � � � | j Z L 8 �     0 B R h t � � � � � � � z n d T D 4 (    �  � � � � � � � � r b R > 0   � � � � �	 � � � � � � �	 t b T F 8 *  �
 �
 �
 �
 �
 �
 h
 \
 L
 6
 �	 �	 �  
 
 �	 �	 �	 x	     � � �       > R b t � � � � � .     s  �  �  �	  �  ��  �  �  �  �  �  �  �  �  �  �4  �  �  �  �  �t  �  �  �    X	       GetModuleBaseNameA    GetModuleFileNameExA    EnumProcesses PSAPI.DLL   GlobalFree    Sleep   GlobalAlloc   LeaveCriticalSection    EnterCriticalSection    GetCurrentProcess   CloseHandle   GetCurrentThread    GetVersionExA   GetLastError    OpenProcess   GetTickCount    TerminateProcess    CreateThread    GetExitCodeProcess    WaitForSingleObject   Process32Next   Process32First    CreateToolhelp32Snapshot    GetProcessHeap    GetProcAddress    LoadLibraryA    GetModuleFileNameA    WriteFile   OpenMutexA    CreateMutexA    GetCurrentProcessId   GetCurrentThreadId    InitializeCriticalSection   ResumeThread    SetThreadPriority KERNEL32.DLL    GetWindowTextA    PostMessageA    FindWindowExA   EnumChildWindows    SendMessageA    ScreenToClient    GetWindowRect   GetWindowLongA    GetDlgItem    EnumWindows   FindWindowA   PostThreadMessageA  USER32.dll    AdjustTokenPrivileges   LookupPrivilegeValueA   OpenProcessToken    OpenThreadToken   RegQueryValueExA    RegCloseKey   RegOpenKeyExA   RegSetValueExA    RegDeleteValueA   OpenSCManagerA    OpenServiceA    CloseServiceHandle    QueryServiceStatus    DeleteService   ControlService    ChangeServiceConfigA    StartServiceA ADVAPI32.dll  WS2_32.dll  DNSAPI.dll  WININET.dll   GetIpAddrTable  iphlpapi.dll    ExitProcess   GetModuleHandleA    RtlUnwind   RaiseException    GetSystemTimeAsFileTime   GetStartupInfoA   GetCommandLineA   QueryPerformanceCounter   LCMapStringA    WideCharToMultiByte   MultiByteToWideChar   LCMapStringW    HeapFree    SetUnhandledExceptionFilter   GetStdHandle    UnhandledExceptionFilter    FreeEnvironmentStringsA   GetEnvironmentStrings   FreeEnvironmentStringsW   GetEnvironmentStringsW    SetHandleCount    GetFileType   HeapDestroy   HeapCreate    VirtualFree   SetFilePointer    HeapAlloc   InterlockedExchange   VirtualQuery    GetLocaleInfoA    GetCPInfo   VirtualProtect    VirtualAlloc    GetSystemInfo   GetStringTypeA    GetStringTypeW    HeapReAlloc   HeapSize    IsBadWritePtr   IsBadReadPtr    IsBadCodePtr    GetACP    GetOEMCP    SetStdHandle    ReadFile    FlushFileBuffers                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                            Tw@         '@ �@ ��@ J�@         ��@         ]�@         ��@     .H  ��@     .?AUException@@ ����N�@�    ��@     .?AVtype_info@@  �            ��@    �b@    4�@ $�@    `�@ b�@    .              ��@ N�@ N�@     0�@ �@ ��@ ��@ ��@ ��@ ��@ ��@ x�@ d�@ P�@ ,�@ �@ �@ ��@ ��@ ��@ ��@ ��@ ��@ ��@ ��@ x�@ X�@ D�@  �@ ��@ �@ ��@ ��@ ��@ ��@ ��@ ��@ ��@ ��@ t�@ ��@ `�@ L�@ 0�@ �@ �@ ��@ +          ��@    ��@ 	   `�@ 
   ��@    ��@    l�@    H�@    �@    ��@    ��@    ��@    L�@    $�@    ��@ x   p�@ y   `�@ z   P�@ �   L�@ �   <�@   �         �       �  �       �  �       �  �       �  �       �  �       �  �       �  �       �  �             
   �   �����
         �"A     �"A                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              4�@ 4�@ 4�@ 4�@ 4�@ 4�@     �  `�y�!       ��      ��      ����    @~��    �  ��ڣ                        ��      @�      �  ��ڣ                        ��      A�      �  Ϣ� ��[                 ��      @~��    Q  Q�^�  _�j�2                 ������  1~��                                     	               	      
                                                !      5      A      C      P      R      S      W      Y      l      m       p      r   	         �   
   �   
   �   	   �      �      �   )   �      �      �      �      �      �      �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                           