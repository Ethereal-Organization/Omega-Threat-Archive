MZ�      ��  @      @                                   �   � �	�!�L�!This program cannot be run in DOS mode.
$        PE  L             �                p           @                      �                                      s �                                                                                                                            `      4               ��@  �            p      :            ��@  �         0   �      B            ��@  �.rsrc    p  �   �   F            ��@  �                  �            ��@  �            0     �            ��@  �            @     �            ��@  �            P     �            ��@  �            `     �            ��@  �            p     �            ��@  �            �     �            ��@  �            �     �            ��@  �            �                 ��@  �            �                ��@  �            �                ��@  �            �                ��@  �            �                ��@  �            �     
           ��@  �                             ��@  �                            ��@  �                             ��@  �            0                ��@  �            @                ��@  �            P                ��@  �            `                ��@  �.spack      p �                @  �                                                                                                                        VW�L��×/!8DO���g��ږ F+���JL�������H��J����&Gd� �ALC���;�S��s���a�
����F��?B�͘��FU�1�#BH��G���	�у���ћ�7B1�-)��N���U�חߖ���6������ֆ ���C٦O�J��EA�� Kۊ���*��EW�?����"Szd�3_Y[H���u��R�c(�29o�_���k��nM���1`������/�u�$�U�7�*|h߈B���7d��C����א���fL�uQ۸�mĖ����dQtۍ+��*2�̲Q�"�������8������2M�`	�CJ��j�2������/6)��>1χ�G����,����D�����O��:��Dř}��ٻ���.�4b�)&�ucP\&���j�ƤH�
���诐�7��0��=�a��L�ä��R����$j	��:4M���L+�80P��H�fl��N~⊄��RG�J��N�7 ���L�b�H���T�'@/�#;L�p��J��籭�j�O`�/p�K���Aw08��LoDB�����:��å[@����݊�0R{������F"q��L�x�N�/�uRCo�*w)�b�c:	��"��)Jr�*��C*N�LRw<QO�q���-�x����φ`ܲ�L�M+B�R6&�(,`~��@�Jz0o9x�4l�B��ߖ�įd���#�A�7hJ�8�D?����1/
��ks�����w8���b[v�B��#ȵ�%g�8X.ݺ�H����/e;XZF�����B���{��/�'Ԯ��h�yhȁ��3��v�0x׳,�����I-�j������v�Z�����sE�<��T�L��E��J/�2I5���I�7�/R��Q������U�Y���%�'eY?�f-7$�<̗�q�D8ز��{J���i��m�F�b�j0nt.?�;��G!O$/GE�Y�1#�̩R�5���EcX�Dt����5i0M�$��(��Xs��,K�
y��B�|Tk��������V�&�
HLyUU7Y&��J�ە���j��v$	B�߸��wǩ��,��i>3��\�!���"��DK�%�I&�l�.�����	9���%�H�æ_?Ka���D/�����nBa���w���^#��
B'�����}t�s8��'7F���
#;?C���?4$H�m�sE���
�X����΀�#\F��w���#)�%�8"E�,��(�z��M��ek	RGM �!���CED�P��!!��{U��)�PzۡM[��K��=1�H���I7���pǰ� �ưId��Q�$�u�a8�T�y���e�EV�({���5���K�zs<Dʣ��bוy���S�$%�`At�,��	*;��SI%�	�է	n��ח��q�0�d��� ֖�=��Yf��Q�l8u���^��4`�qo��s{/��ʌM��ȑW�Y��8���?N���WK��/�����J��<��c�}|j�M%߁�'�p��0is�s�Mͅ;��Cj�@�*�X�6$ב��x89_��y0��7!>D61�ߟ����n&�+�Q���A�	����!<�G������;��C��(�#� /ב'�"D�4,Q\g�V9p�:;���O�B��B����/%A� �L6�$�%1�7�.����BL����r�Tː` B`�ֻH8�0R�$�IM���R��6L�}�O��G^�n0�/L�e;O�M��$G�?m�����-D(����
�\�$�Ly�0OM΋C��,� MсC��OЀ����,��u�9�m�G?�M�4�Ȝ���,S6(l�N�V�~S�L���]����{�0퐻��h��bN�D���O��4b��0���
$�r�:ײ�H��
,�M��>T��W�Ԃ�D$��!L=�Q��gYh�;�"M�zR);6�3^R=����h�D�َCˁ,�F%}�d�^a�� TH�f��
���`�?���B����J��Â�D�N�;�q��{�y�Td��4?���;\��8'�����@����BC��%�?��R��˾A0��Q�K���b:ኞІ).3�?���Ts6]�rDeá;P��4�LD�׫P��#�6>�g��)�E6�Ƣ����:3�5�7��r���Κ�+JB�?��1�ߖ��/��L�h+��(Ti;��A8�����њ��y�����Z�L/��'�w#�/�cR�7tjd3	?L;_7D�N�&ʪ?�Q8[D�f�2d�����!8�X�A`a�����"��W!c,�~\��D�e5�&`���D'O�
�Ȯ�}P�m��6,�
#���R�� W���#���0���)�/*���3��{���ٟ�7i@��L�mu��D�Қ
��ځ;��D9�x�/Tʠ��׉J�q��D]�^���Ϲօ�"��d��kHsh$��ӁN��r���˰é7����m������8����Q�o�4�F��Y�0
����Dߢd��ͅN�����ĭ9����8n�-���5j�`"��������J�L�tN���g�0��À$կ��G.����o8�,�H�D��_���(�B�
F��i*rP������ϐ!�����|<C,�	�#��Á�˞���C���C����y��CJ�'4be�#�?;yY3V 7A#x:�i��}XJ�/�Œ� ϐ�M֕���Ѷ�t���0�5ӡ���,ӏ�j���2�!�7�,J�z8%�ņN�"����'�L��e��8D#�,v�`kM-.��J������`��ũ�me�	�)��B/���M�`��F&(��|��{/�d�1z�*��ꞔ$��w[��Z;���ӽdk
/[� �Kze7���@�c̵��H���W/�/AZ[1`�����p �,ĭ�I�f[���{/�/2�3�gUYks�2\Λ_��/��<����?�_0C?D�S���"k�
�fz��SB7Ea
%!@DpJ�&i�	L��n��tE�6�
P'��/��'�������*���ЌI�folz�`L}D?Ĳ���g!�H�;��%��?Ų�%0�H@J��D*!7�1יZ�c���tآ)�W�,�ỉBƙ�,�FX�c�����*�沞 e����{щ�U��ɳ�v}(,�|H�ϗ;�F�4IO���5����E,�,h�M��N�Ë�n>����R�͆x�g�♄���4Ɔ�d�+��~��[�6�L8�&:W�'��"��X�Ņ�.��c'(�o�ڲh\HDK",K���ߐx��T	�����O�Q�1�á��D�헂�����	��
�/���A�,��>��F�����\���ӱ�L�ۙ��<���q�㕘^�ۑ�GR�t�,���K/�2��Q�%1��t8G�Z��RG�7��@s��xà����"�)|�#Â��B���$��.��-�'u��L�_`|Ά�C�?6f[�b�����/����4O�F>�����<����EDL&�7/2������. �L�4�8Cy�1������W�Ԅ�[�d��3��I�?��J���t�B?�A*� '�7��ƻc����?hR1�>�&�3�����,��R+,U���5*�`Y���W���<��.���G��$���/����,��h�JK��Gڰ�,%.������`g�`���V�5-�4;N��ghT۽���� ?l$��7���u����f|���É�'�Ĥ�Z3hW�GL��Lz@�D)7k&_��o���M���,n�dpG�Ś�Ð��G�ǊJ�O+��a�����[�ϖ�/�;�0
�1�X�ue�J��c��oƌ
��0A1�h�XoH�Ҙ+G�D�aL� ���#�(���'�����Ұd�x��Sě�H�7��˯���0�����,�K���\���h�U4�7�7�:,a�Ə#r�;i��Z�ui�̧.��7�.�Í� 6���%��!"7z�?U�IU�뱑ĐF��B�3�b�t�&o�/��#��6��a"�N�w*��T�I�B�*��(���i΁/W���H��{4��;��E�b�d#[e'����D�����;�
.�f�$����33dm�AH</[�'��>-�dB���	'8��7��1�(�����xN[��#d_�'(~%F��D]�<?�v\ӗ�(�����
��C^H��w'6�{����D�m���1ͦ���Sdşr6oeeR�i��@�R&�E��*B"����b:��Lo�1�	��CCX�hL�ٓ�'"��(�+'��E����ӱ+(SP�g".�(d�1�x�P�L��M<#�!Sf%���O�,qY�s���By3LP�#s�`�ϑ3,P4��`V��/W�F)KX��Ƴ���4=��g�`�,��?ڙ(�B6�R��!�2����V�@
J�ϗGt�GdB6�,��^y�	0ĊYƩ�}RI�$L.j#��>8������ܜK%�H֪��8��<7��b�����;�RTg��rW�=O/�`���B�� ���"���K��[��⃙�*RjOB��/ɔ1�����)^,F>����~�Y�/+4D���=�r�?!�fc`�a���,�t!4�4.�E.'V�Q�V��겱�gs!ӐɧC.�Gfo��Ӆ�=�p/�N,������jrd�C�F}fkA(Ŋ/���ϊ/	�����x��gn$��/ү��d�s� ���3�3��3�"��[	W�AǛ����7�GO�+�)�fX��L��J�;�7�Ԉ���D)���@#�*�)�ە߉�����"�BL�@{N����b�FLT���W�X�,*�%����F@�����C�d��AD<²0x�Kϑ�.�W�41�ۯ%?��:Q�L
�D>��c�|W�%�S�����J�z��
r�'��7ˍ�0LH"�[3�Ihp�Q���,��W,F���V�C��CT�BA��J!E��H<A���U���MJ8�d����N���,�����%u�d䖠\,O�D���Z�%x��__�����R��E��`�����ײ2J莙��(�M��_�kb e硬�+@XM���v�9��iY@��qY���0!�,$G�D���������=j2S�!.�� ���ڢ[c�"��Ҷ���`8P���:��ƀ�/��4:J���,���z��1�!6nB^��4A
�ez�/�)��@B�س���/�uvL��G����bvC�A=�R/�����,���_oL�:p��8��r5ANQ���q�B�����'��3���O�y;�X����$f*H�#L9�߇Ne?��8�Р�Eǹ ��B�O���5�SA�����Q�0�P=KA��/Я6�Pӏȶ��4d�ښ��N�Ī�lk'��ḡ��+�x����*G� ��M�Ƈ�=��N��C��1EFgm��Ʉ>Ƭ� �M�Oс��,U	a{1�A:,T�«3
���D4�4�Oف����ͦ�A�ď���K�8���4��a'��@�,¡(ĕ�6"��L����
�!�(��F��Ç�),0��1��HB��n�G���JF�<L,�pϒ&���S�,L�B��Ʉ���(�����M�%�D�AV�H�����L h{e�S�<��� +�<A��-�.�,R1� �Ј��D��L����L�HJ?fK��@��+��Z�ҝ1&���
1 ���Da|,�0Y/�@H�<�E-ň.H�D?��BF�D˓@"P���t�8��߲>H5,�0#�?���^0N���86�,��`3�F)k*�:%���{M_D���/�(#(�4L	��'��,��ۋ����p���a�ó��}���1��֑��L���1,̰���%ړ��|B')1tS�H+����(�0/*;Kē�3���LlQ�k�"JA�*�7�ݘnA� ���(�f$��=P,_%����8
&�v��r�%�~|,�J�T�Kz�����P�d��x�1����DX�N�JO��G�$��L�/EFI}#��JC�|��LR
�h8���ė����Mq)�Ƙ�
ϲ̤�?�5^�9D�D&�V�BI�`"��1N�aO�쀂:D��9�}�Q`��8:J���B��Fp��1�,��0�C�2$�3�o��
�Аg���~�D����,G�k$�'I�͞��o �D<Ļ)\8��n7*�J���٭�O��E �F�����L-������M��:Oɝ��I������ID�@�JBY�.H�p�S?'U�0��Dzh�)���µϜ���bl*�Wם�����;���.-gJ!
�Z/�D����� �����O�� �ބB3��~?	�/Y��/���,�%�9����蠠ڸV�R�Cw/�.�0Y�����%�kf���,&�G��	O�,�<5��.�,ʄ���~����Ԥ/c_�G����"�/�ȉr���A�a��K��:d��?O/Toe�����Q���k�	���/J7�Ɣ��q����������s�x���z�^;�0��0�o%��E�Hky�;y���D���z^=�J,�aH��>����8�2����@���e�M��S }2=��ϴo�ÏH��#����y�b����,f��0�o'f��]�8�F�5�/�1��������2ۗ�@D!�%��f��H^ʒy��3E}��1�;/߉f�Aq�y������+F�c���w�E׳�G���C%�6X�!��Q'4�Vtm��/,�ʎ�"�F=v26)<��w?��x�c�M���/�YX!��(z1/=+�������&PD LF??D���?h�g����j&]�����'��p��ߨUůH|�qs�Cd$nS~��b(s3��,Z��T1�tH�)��7�3ق$�_���f�Xn���r٢n�X\���V�{�H�[����D�S���_cldW	N�gdiO�?��f�BG�[IOA��y4�$~�K�����,/�:{�+��Z/��Z� ^9D;�|�(����]�K�}��N�7L%Ɏ�;��o!3���J����3�;�1�< ���=�:�D��ĭA�L����ϲ`� ��|��GL ,J���0����9β�W����J�'�!�[�!E����!�,�B�`����3Nb�.�˯������1���W`��3�]t��%<��6N� �����tLِ,��97�%N���P������D<�y)0�@���òᤚK����'TJs��A���@����NR�y��$�HϚ�k^��i�FZD�l��/�C��meR_�pl�����MJ �QO��9u���G��$��`[���8n����ߺ�%׎gA&FV!C}=-)C������N��v��78�a"0��Kl2x!L�K��˶���ďr�G�$�Ԛ�
� H3�\�Η�P:�C�DcOF�Xa!9��I��G��D��U9�n�����ˢ����>i�L�f�	�G'�N)��L�+����>������w8�A0��B#�@K��X�/�6SE)N��?Q*ݡ+��-d11�͐
�E-�;��D&7A#>Î����	L8z^����3,�D'���1/�Jfh	���ϴ�e#���sX9��R}�1�;3� ���L��'�l,!�4X�K����M�@l)U,P*8��D0)��/X���� a;�Ӕ�������zuD��j��.��+N�6�*�.=��;\�KW"�ww�R������$��	��X���c~u�KV�5�pk;ؤ�_����.�@��8�a�I��	��gƭ�� �B��&�,0LC�>ň��6L^�>9��D��)��0������"��D8A��f,J����S�+�O��	9Ȳ��%�+��,�ʈc�,A�#�Y�6�To��-����d���
?����i��+CS�����6����sF�R��"o5�ˣ��9�̺��ė���%��x��	(�����򻂯,�)
�J�'!�U�R)J{��.����,?l��N�V	;K4�3�7�(F�$�;����DJ�� ��������ս�آ��p�%N�J��c	M��OW��8�.��]N�.p���l��b��Ӷ�%����(�L����I��i��F1O$�F��`hN�׳�ï�묵����T�����}�Y����{L}.�" ��v�U�c����ق��������%��ÑP'�a8��d�\��&��k#���'Ä㍒<�� �ݾ���׈G#���?��.TDuP@��=������a��O+M��~�;���7UC�CY����G/�#(�W�-��8�N����[?�a��O�J�����Y��{�"�M��i�C�{O����ο�}��-0�af#�D���8�ZP�y���,گ��e��H���)��)zϔ*'���@��4�#�Pװ��h(\�7��D�Ym(d��g��,�N�fE	��(�	EL >@�h�I_��4���J(��5���*~�'�D:�Z����N�2�!�F:j�׻$,�/��KT���?��GH�Kq��C;��S�78FR�,�w��ȴq���F9H���f���h1i(y3@��c�B&�d�Ci�!�R�N�4�ʰ�RrW��ʍ�&�OsÐD�Y�7�#;y��}h7���H��H��K"WĊ�ze�e��E�>D�}��n#K�X!\p$��<=�o��?��F,0D(X\'�uZ��O�ó�ľ�8�A+J����˅"R!=�(�1�/���1���;C/�H�_'�;)}� ���ױ�
ӵ�X�~ ��,)oȲ��WK}�F!8��	�5��*J��`��(F&�7�C��?�pC��x{�W����>�.���q���G���&Q�6�X��B�Hf@�-�/c9)�� ������-�PaX���SIߵ.��D/�.�ĺ��>����LJ�� ������Ҕ�1~W�\�io.�)B��h8��f@���J��&?���L��L���ޠMӔ�H5/��Of�Fx������?��F|�	��.�%lND�؀��.�Y�j��и��s�|˼����\�,/����;�43�0J)�9 !H�2���k�9R��i����(�Y�.'�����i�;BL���?�/�J��;��pd������GO3�en�R}$�Ӝփ��6ܜDj��N���b�7�P������;,a5��0��$mO�@���X�J�����@!,�r/N<с��lO�2���cvh�v���^C"���(JF4��XB������4�L�
�J^�B�x����b�J��O) �����`�,�D��������=.����0֗�� 8J���4 ��M�C���<s��G�����,0�>��HMX�[���������E^0L�, �4ĩB���z�|0�����h�-��C��Υ�h�C��Z�Xx�(��hު�S��O�I�,0'
���i	���,i�Ĩ5dp�b%�h�OJѠ��%��4�y�$����RD�]�X�:1o���/aq�O5Ix�YP	��^����9�SB�E���tZӠrD{%�����4b8�R����}D.õ0('���0B��J��?W+�G2k	"�@CO�����yŶ��A¤],JR�,�&v��aa�W�$��E�)K@ƈd�	�H��"�D�ˊ��I#tNtH�/�D+��H7�D3��H?�D;��
95��	�?
�H��	��WM%����!���h��j�,J���:��I���p�:��;��7�B0Ifg��F>!�?�b7�&�d�	�Y��!;�ಉ���Wq=�� ���)H(~�K*YWK(jK�q)B�(��AF�(F\�ck�	s�{"D� Hhۺd�]"E��$�]"E��$�]"E��O�+ ?���"	�E�K�A��=�y�V�­�/b�~�����{<�Ě�&!��LT��b�X#AM�CO�"�����-����pÂ�b�>�b�J	d���'q/���~xEO��n���4N��C�����TP�
%� [�����f�7����6�V���O���B�U�0ȞxG��D�/�NQ4l���C���A(����)�|J�(=M�2i(��8����@TD&5Ȭ�))SL�J%���!ýYO�\ L��M�ƿ��g=���X�MU�C�W�G�(�2�IG��$̼Yv��Iep/»ls)�d�
/�Cq�yx�!bĞd���,b���8~��UgCF�9Ͽ��e��4/K$-(U,Q���N0l,��4����IC�u�Z-DC��"�V9�׾�G	8��k:Z!�;��f��)HJ��c!���D1)�О
ʉˏ��G�������$��m��m�k�����C�DĘ������8#�H��,|y��OC�+B����3M;�5(BJ���	��J��aq�}	���ГT{+�5��${�����m�.Ml8j����萈=h�H{B�J�W�(�,/*)�$B:@���H5/)��$�;����e(d�S
_��Jhs�L��̳I����MS�Ge�WG#,�6ų���&���gGs=	x,�:�&���
L��FL<���TJ��2���

���O�<.�,V'Ma�y�+ʰխ:/�$ݞ�k�������b���,�0��bƆ'�����d,��D�݌C�~�,
J	�
9�ρ:1��
;��L`ް������>!c�),¿$�Zh�j�Pl�&aZ���m*��ro�y��	$��#�P�����V��!�D������q�#6�9��:�;9=������C�����3�K"	w��]��]��Ԇ@f��	D�ˉ�;��3	E+8����$#�"	�E�9���,G���1�/3����������3\C2K	S$[Hc�k"s���V 3'/"	?'ˑ���r�V�Ng���/˔r���m�M�J��|�,��`=%�؄�vϗ/��M,�L'ʷ��+M$Æ�'�z�ف,G<�m�D�Ӄ��6�1�'�׎J�K6��u�	��H����9�)^��p��R����:���ʢ���!�N`�����S�թ ����ƁKX�<0	�x��D3�����˭[���Ϧ�)�f� ��H��.y���2̐V�43�LX�W@��"��1Lh��A���p�?���v�3���˔��
KK���h��6���HI`M�.��k�J8ŕ�2J�{ ������H;��,�*0�K����Ƣ�D&��F�?i�<��B��>��1��p�*�k�f�5��=3,ֵG`1��a�ج�f������a�τ?0�'F��4
�?ť�l��� �`F���$��b0J5i��9(w4aY�����Ã���0L_�9
D���WN�GF.
�
B���+�Ltv&�In�;���Cn����|ʼ�K��;��w���/�8��d*����I��d�+���fDB��8�e�
�f�B�%��f"Q�N{�f,R?���˖p�@J��,�>D=��!׮������=bUaB�҄�K��*K�4lw�"I��3n�Ll�7d��&��	[�H.�2���
����.j"�?(��(2,���"��'X@ݐ/�-��p滲8�D9�{#NlAB1�� �x��P�>�T{N��	�TE�����;�6���f?A>�+K�N�Oω �9�fW+�	iS h���=J�[TMR�%���0,���BK�}�fYY~����x�
B�/{s^��d)@�����Mf��������O3�g�H�Z⚅���{�N���I�.��������uc�=i>"C�4�P�$,�dB�P���,N��7��ӹ���/Y�挘�Qf.����`|�I.��nUE?S�i�zh�/J$�[�v���FD��q�R�#��5[o�����<�/�ĪS�m�o��Եl{��EN�or�C���v��b�DX��4��$b�CޮK������U� e��~��u��Aָ�Y�3U"�H+���"�d��Ψ<�
�'�d�-a'����s�+�#h�[�����,V��aR���o�r�S#�_���R�.�Hi,ϟI���J�pʗZ~�_L6Y�134����?�MOȿ�F�f����@o�J%�#@)���R�a��&W1��,�B�lJ@�GF�O��ş&d�.������f�#�4)�4	.X�5BS�ߴ�i-2��g5�ߛ@��%����J���+}�=�3�����-4!n���E�'�H���AB'�`M:V��%�T� �����D�ӜV��?��Kh�˽�Ha��/�.kY"tF<Č'��;��Ŕ/B���� ş`�,\��A�?��q1���G����O�ҙ��|,�w�ݢ��J����Ė��J>���DnyR<�$籿Ib���@�,��:�l��-n��tJ��ݘ��˴$�pÆ,|�^�>H�?����A9���V:�w�C��!Ϳ�%;�eO:��l�ب�9���8�Is�J0����	4zR2Oj�������l��@|6�Er��김                                                                                                                                                                                                                                                                                                                                                                                    $p{�X�	H�6" �zD�ډ��(0y@�P\$lHx��"�D�����$"H����	D@P�`r$~F�}��	
Q�@x��	Б�"���$�H���QvS��"	�D�����$�H�|$">DXn���$�H�"�D����	$"4DBR�br$~H���"�E��N�u@csm�8R�	 ����f"P�� �(t�� )*�)��8,<Ҕ(g��J8�m-�fY]�G�"�D�_�GLOBA�HE�P�S�{�CT�D"}M{V|R� 8 runtime ���o�l f
T�qS����INGpDOMA&
R6028- �ab@ltzozi微��z�h~p8�(!7not|�
ugh�spafcHf�tl)wi9n���8S�kz#tdy5p1urXvi�t�hDh�c$y�hR(e4?`7_V�x�h/� ݄�`+19��Np��=ds�!d���,F8m�J�dd�ZX@$7��ml�yPh�a�"ck0�nC5r���_��bDrmIp��gz�B���7y0�9OP�"�BVm�t^,85�s�u�)s"`�a@,f���ng�x�j;�%'r��HM.j�:f,V뼈�Cq+�R���LTb�rPy(
�]�E!�$PՆ: Ai.�P�R�M�Zk�w�>�8GDtLa�3Aiv�P �u�T"W��dN���s�ag�B�xA�u� &32.d+)��C*\@tس���Lb@^f�f���)4�ň�X=Pb\+�h<�(8 ����y@ ���У��v@s�@$P�L`
��ĩxx�0��b�Q��XG�!��)�v�pQ�\w����,p5x(��@q�0K(h{BP��0��EP&��YcEpp�wDyl��Fi�LSEۺr��u�0s*�]M)ov"�1C��rHa���W�N=�=xPM�kRhlr��*1NTu�IkL�3Οk�CPysތ�nO4q!
�vց�^��X$Ga@�l��`����2cT�pP2h!���y%�Y�n���cPi��,z��K�C��VJVQ��D%ir�V���o����$�qAd��Du��� !�s(edul��NC)-2�Unh�l�B��p��E���RJ��jM��p�\t.Y}	@TCom��L�?�D�+N{OP�����gS��n�iKERN4L�N�wsp5tf6US�0���g��V�u*El�H�K�(�hQ6�!"D�"Op|�C*�2���% >6Xd�r�"_�:��Cb���ESCM�Dr%(?���r#��";2�DV�PI���6tTwi�a�R�Y�<u#������#�@cupInfo&P�V��s4�SH�&AQ��1�&�0�NTg��m�;����2Bnł�W5��$HdE��ժ�Jy�v\W L�ydeC�r`LM���By���z/�1d���d~��7��2$�L
Hd��^�TypVPJ��i��u�ۏ0R�$&i	z�{o�.��̨m-V��EjYY_�S,R�#'�IsB�G���P��$�h>8)! ��W��H�܉���<T�,�
OEM	d2�=�G�3���pXp&�4�@W�Յ9�
�E�Z%W�а                                                                                                                                                                                                                                                                                                                                                                                                                                       ��wDU�;G�
XIg9pytfB;axe{���cv�J%m)0qo`FZSABTGPIX|�gzf�sza��{q�b�5=[A�V`g��aC���|z��F7d}H�@
Ydl@;ETM��Q�W\[f�nc��Qqy� G�rV�?ta<^�l=E�(x�ʭ<,!H(�n�ty`�Pm=)B )Ale�A0FL��PXJ�w����ymI�/yf�Hm��q�0Fl���xGz���I�&'�ޱ�;�m�58s~�!H06��.;q�|�*04PZ�{FVXt��r2=<��QD��lK�Bn)Ig�<mI��F�QA�I�J�|���TtP:w<Fo�g' �YRmcs��W^?x{� -(M�RhR}%��5@eqJJx0S`v@^C�J�m�"�*TCa$�J��szLU��5�S0��8��&̕ �	A8���C�Ș�țy�!��<�����"	D���S "(�a��0u�"!�0�(2�f$�H��"Dq�9$H��g"�D	y�mc�dlHY�o")D�-��=/J�DMr��A�UUT����=��u9�l)4���B��0��*��@*k�a�aԶ��5NhŔ�4p2��0dTr�!ڷ�������NА*�
1D	�K�;�J<!'p�����$kto�Ue5|=��B�]��d�/F"��Y�8@����F<,5U^�;G��`                                                                                                                                                                                                                                                                                                                       ��	X�0�e0J�H`P��ppBpIpNMZ�3	��
� g@
U�s��	�!��L
T his prog�axmtcqn�t�bze�u��i�DOS�mode8.�
$D�8�H�|�&���*�}�-a��(�S,�x�"3�*!p4|'a���{�aJɑpl
�� @���"ARichD`j�PEL�0�GX��!�)�vH�d���h�P@4��
��>	+�p�C�/1P^XT�S�
)��y��04��p���.tex�e�r��ńM :.rdat�>0s�2+�(F@R.'p"� ��Q<"B��.shared�$pH�>����sNcQY�D�*xc�loSd,2�P�(pB�_`V��3��F���P����`��^�S��a��q�D$��t	�������:U�� ޖ�D��thȓj��ߠ�;��2V(X�QS��UV�s0�2t$���I%�wl$�~P`'���u�=]��[Y6�Fhtv�<�W�{���ȃ�ݤ�K��͉�
�L�Q�4_�Ţn5�С����1;�vJu�>�7d	{]����t@�s��|�p�m1�PC +ō.PQȣ���CI�=0f�_KD.P��w����A�� �Q��u��Ç4+�c��SU@����h����
�s_�L���b�&�B�ƂQ���	a��#����E��Q�&� �j��
h#JU�:�!����A�u�����U�V�(sp����щ��1�K^��tnFQ2�L��zk1�_%�R]�S��!Т�Fw�
[�w��X�H�"���j���!D�VW���T�X���u�t�4�Z�R�%�8��T����_�ӯ��S*�L �W�~�njnF�pxY�}?���W��� R��Y���LFj
�h���	d�d��P%��4ː��N� ��ؔ,��J�a�QT����|���UK1���PhX�������D��HGh�0�s��'b����t��ҵ�x�C��$�Y�"@��P�sùP�����B�Q*mW�V�}6��+TMPX�IC|@��d=�'c=�P������lR<��ݡ�H�&d|�;�,'�.k��	����B�ˁ�)!���
S�Nr5���G��?��Zp���
L�2���	7��j�I�CpS*p�����T�u�)�JhT��f45��u��2�f�\$(�o
!� @� Ru@���(�!��*�Oj����,Q��3B�f38HV��G]�fA$$A��P4.IQB=#�`�"=�{������jX 5�zHR��Qg(�q ���!�""d#��P0L���g=��@&�x�Ix�r�hH�H<��d���$�"ď���F��ťhXYWT���f)��Ȋ &A��;�:�&-��;
>
�T[���� ���I)�)h�\����@]ʐWh��(f�&=�-���F�M�"H���I�� �*C/ԛ�>��J���+u��wDP$QR6�0h�4�5�MD<��U݄���R��$T8�P�]B9)P#9��9�QR�u#5�L�&���E\I#	8D�&P���3�R�J���̫�$�N)j�� �
!J�@��(�I"8PQ$�D^�!�َ'!��PQ=#LR�hVh�	Dx�7,�u�l��ꍰj
3.���
��02�U���lW��$�������H�1��-H��eA��SbI��F�TQ�'M�tZ~;��NME5�	j1Ir�8h,If�Wh+�$DQ�'\�r)E��u��'G�E��zWN8��J�5����$��!K���Yb�:h�Y3P��(�ESV��e�u]��E�u���M���U]��]�Z��=uB���ȍK�A�3���1�s|������jyj���Y�W��0�GQHGl6E�(�"6�VlG{�{vم����}̉M̊P`\�U�*�q(��y��t�E�h�8�A��X(���C�$j۠���n��;���C�0�Lg��;�!� M���XQ-(��3�UP~�M����3���JM�q�V�I��UNG��R�;��х��ę�x�AE�VTrB�;U�d���W�R��o~�"I��WB֍p,I9��m�YH���5�'O=�
�M�V	��z���fW�����>P>yS�
���O�2Q0͚;�ԤRPH�>u�|F��kہ��	��NV[I	LZNh�SW�Qf$@4��L̳���+���i�Mx';x��5^Yt��m���D�lt�]ITK��'D!��1�ޝ�-������;��Y�EF����a�
�{��5��ga�d�$VQK*(�tb-�em2Zȁ��x���4EU�$ �R��!g)�3�("QE67fR�)���
|,
��LV0�����K��g���|"��,�QbU���T	4Rֶj�U�6=f�:P;ޠi�Q̀�8��R��A�y�4���[�z�E�b�)�L�S�\$�'B"T��;ބ��︃rL(w�J�5�	�PfK��A����|�;z��tP+j
ȓ�1/Z�+ހ�s���~&��)��JS#J�F��3|�t�(���};�t'��� I�������H3��h�5�?��)9���\L}(�P)��t�l>���"���0�����6GPeR6�;��#��R���A�������5��F; 6�[q��i���@�$�Q���?7V`"���R�P-�|!2�E�)p|� \%{��p�W3�8��(ow����p<j\>`;G;�|d���<���@V�u3j�)L'���� ��&�(X�<�h��=8C�X] @���jI\�%�ffM@4�;�5�	@aֳS��Ue;hi�,��#R�RMy87;(Dl�GP�+0Bd�0�f��I8���4�,��	0��K�؍l�!�$��OH��K�M�|2�K�A����<,�CVB2�0�$��)c�>�u�2x��H����S4��T-H����"�{p�+p���%j��AP�d^$J�ÊQ�'YR�R>IL$PO�x�90�=& �Vh�A;_�������@V��A%t��ql�2�/�)�(^�{�Ra�H�V��%a��;@B��f�H��gFC%����?|@3T��f=�N�0�P[��S�i��&z}�X(n������˪dRE�n$`WNwC,t
_2R^�(z��B4�eP��jr��e)��b,��35<C�	wDK_��4��4#�=� ��1���1w�3�W���b�^Hb)���%�zPVQS2�e<��P���,��P91��;�:	pf�5��<h:����8�B�������te���X���*�e�3�l�L!��!���+����Ȇ��,�x8 ���,2*@��
�q^�B�X\��/�6��R94��X��*f�Z�7216����`�<jT���L��@��	uH)X[$�(A��<�M'��[-�A�0���@��OV��fv�W�&8c� n!��<��D�M�H	I��N��f�/��$��:ġ�3O<@�0�#G<TR�_��[���2t�a�x���V1<�t.#� H(q)5*f=[QJ�Fl˛^U$s�*@��Jd0�\�]3�=+ ~��5?.!=�>.1�^I�4��B�ȼ<��j�F,r�J.Q$G(�=J,,0�YX�v*<�?�;�uN�0rd�CA�r>z}A��?�{� �l1�$��l��U�x�P�1U��(�s�i}�%��+��@D%LR����5�z�
)��l������EQh%a> A@U��B~X���v�$V`�$�."1�.��?�KC�Ǹ�;�r|0�JU�<[,��&����B�PH��;�F#+F!f�͑�5��/����D"��-j�X���W�)��Q#P ؆�6A�	��4��5��2ʌD��W�Q� �ԯ��S{1���QpJ�k;�F�$S�3W�:)�$U��l(R��Z��W�DLM���
�<�U���<}�7d����Q�Q���=�v�P�V~]p�ޓM�?�c�&@���@�:u��t�Xu^�������(&�',o��ؒ
�L8G�;���|�L_;UD��j�T���O�I�҄z�G�z��d��v��ѷ/y�@��tR���4�%���	�k�	����AQ�<TW6;�V��%�45٭� RZM$�¾���TG�X�d��+#�(#
�.�d",BN����\{ԅDjI�'�J���+���E�ۉ�U׊7tHڸ�C/!g[�jCS,tй����CF�Ȉ�y���Sֶ4�$��������y�8�!>F!(NЈ@�,(�B+~_@^��!�_��e���S���"�U��©a��'3|B��4�T�k4_]�$xpٸ,��C�s��ęu��o!�Ǧ�9�Ou����k,��#_��w��I�@y�Vty`\5����}S�W�����V4�c��
�9����jq�pZ�p�����dS,���{)�"i1�_[!+�՝�T�0���jh���/*&E�P���2�0$���rj�N�����%B�2`Y�Δ�� ��'$�h�ƣX��� ^!{�Q+J���5\�.��B��g�o��Q�]�;�%t2�jX�Ɩ��c�NǧB�H���O���I^��u�Dk�
�DNG�T��3ÔQ]�@��D0�-V�-�O�Q�]�O%�عŭY�	G���Fk1C�d$�fK~K�� *дɊI���Pm�$$��u	@X��@^�v�b��(j�
��	h"I"Fp�sq�!�,v!���#G/!�I@Q9�+ &� pU�8B#F����/��2P	]$�H�83�9�3	C"	+Dp�ѐbT0�A���lj.h-6�5�����[h4��f$i�d�!T��-@	q�:Qh?�-j,�����t}-�O�</f��QlRP�S���38R�ӹ}���p4(U�d����m����R�H�{ts˵Lq�:R�J�L�kK���2
ӂ��lhi��x߬R6�h�'P
%#��eL3�6��|�����0��T�Q��ǹ*�Q,&q�(v�.t0�AL�ɋ()2��ykB�����q�}pK�5UZP	m�<�,�W-�x�?�N�g3xҡ��U��U��	�)؜EI ,�
�Ip0hI���4!B�-��h�o"�8`#�Z�= ����J*�sF��0GQL�,@����E<A�7GBDC�z'�y����d,�$D��B�����?�e�1 "�+DK3����PM�����"���x�ψ���'����,���M�!������蚥3�%�(��U�P���4�T"�%����N�Aȍ\
y=�*�7}&�o	SR��x&�Ҡ	���(�y�$j@ � �G�`��2��+P-�Id�H`�h��%Q\K~�R�+TuIwJ��Q�� *.�yZ*��z�5S� �.����e�ፖJ���;�v��GjBVU�q���j���L�'@�:�uO�G�V�O��:��Ɓ��5���]��+��>ttX�Q��L���+C&sQ�L��<+8�ؒ�HC�@�+N��Z<��Z��W�3A4����;38�D�+�� �I��3wP��kSU�J)+L��8��$_��[��&F�вLVA$H;sw\<#W$=�O�7���H״��I"X���������ј\&�<.tK���G�PV�݇tԌ��Q�OKP&��kv����=`z�R8ڍ��SJ�u���'�-|��(��Z�Y�/πV�QWBO��w'���"����CK
��j;X̿"-Q�S��d��@�ui�|�Rv��UQW>Ex�D{D�S����
Ua&7%�a�є��c,��êƢ/^���s�V�CL-�{	AeUbS��T��$d'���D]��/���� 'XQLCL%���\�p�uQA[���B"�E��PZ�2V_�0VLRS�"\����{a�ޖ��QQ�0�#��	-h��DR��F�N`d��ݜ@�v��	��#�&��'��^�%xͲ@NҹV����&�G,(�N���*wZHV��B����IBj1�J^.�x��W�~���@7�DmP�?��X_�mB~ \P�&�%h�F���IZ-��*̒,�HY�00�\?u!T���E3�;�
~�1(黬5�,W���}iLtpIv�QV��f 	��"<X}A̔!(�$�'����G��H�����P�2�V����B��9�/( _t�yHL��:Ï
<���Ȉ�	Q�к�33\E���	�n�f*��*��.�������o�.�T*lN�� �l�}��w)��'�q%hHt�ȥW���,��"N�-��WV��bxmh����OژǼ%p(u\��v��El��\.5�B��0\Pƞh��'t#���K�Y)���x#��&��mG��4K��s4�W	Ɗ��:S��� ���HU��	,�8�M�\&��OB��,�ZRE�n����)='&j��~|r�~��$V��b;�`	u�f�����I
HP��$2�I�Q1��*HǄ5z�PB��3 	�5��j���D��{$�RF��˽)�	E����,Q��I-Z�x�(BN�^�xG�'��,G{���={ �(;��"ey����m0H��%wa�B^:oƟ� 48�8~]!)QH�:ʑ��RH��l�Ia�I?!���WT^l輷�K�W(I�h��y"G^�S�`����㐉@i�:�֥�q,�٭�]��S��zM%K��#�O�J�a yǅ$>�8�^7�BRSs�	��Xt/�Ew��'�"$
�j3%�IS�K>�œ!�.ZdP�n< PE.��P��2���%	;�2�L��wQ��+�|ts{yP��,3�lIb&x��6��%tp7uI�8�<���7IF?8�u�3~�h�@�a),u e��d��*h�%EL%@�Nd���J����@W�_uw�I T�$oH'PN�ͦ~E�j	�O���]� �W����kj��T��O@Q���I{���M�RKf4K�NX�*��-�P	��5�yߥ�)��8]�	���6&�	!�Wt?z�p5y3Q�2e{r�����P�Uj5��2�R^�*R�Ndd�0�Pt�j7�#��HXRd���}�;�t4~A�?:o�l�K���u�^`��T\�a��JC�k�]�s���q�vnl?�]��J�1e�T�Z�p�K���N�4
���
Y$���+Q�;I�|�I��;�j�N�o��T(`��}�E���n/	$ˉA�� �;�s�����uzpH��v�"(�j�,@E+�3;�G��v2����B�P���S^T�]C�+�dWS�=	�A0�I��"�O�Ƙ�vV��$uRb���0��x	��s@$͙oO�^]��M�VUɊH���4��yZ������*v��uwQ5FF�J˧t�Mk��R$���n���4��i=�G�L�4��l�%��mi�U#&�m;�P'(�B���<x�%� �3ۉ��� ��B]���S$�X�yP�h��*�ʈ�T���P�3;'�uptA��ȭ�hP=у/���|%�(��HRHd;L`h ���f�4H-��q��
D�͢Î��n|����mD�d�WbÜ�)���y	)�>Ed��F�����vO�x'L3�R�v5�� ��S;n3��B�i��w\���B�"��^�	�~"�Z����{/�O�эD��5Pڤ�FQhO�(`&&x�U��
�HT]�{��g�%�k\Yc�Δ)h���c%���-W�\��'M�{d���B16��X��2�a��RKh��PLv�!@BE�};��D@��H@R*=�2�@(��$4
h@XUإ�<�@��dc����P�)$B������:����B|��S�a� �>BȞa�B��B�A��!�O0�J]$"��������QR~7a��A'BJ������C�����W��!�D�cԄe|�UV�@y��bK���d�����ʲL���	N -BĞP���"����Dp�l��G}�zr9O��;�<����WA���Ԏ�M1�3I'P�����qR}bS���
���w�;Ñcx(��,h�&=XD�R���HW��x��dL���VQ�7V�h��`�YO��B�٬���HH����h`����,��V��$	$�k����2��W�H�Q�@�R����$�����;>��K[�Ȝ[�%�Q۸5�zh�)�(�Z{RJr}����{�ρ%��Q��-���Z�y ��!=b|u/ ���**H@tO�F(g��6c��_)Q`^�^ �UJh) �Q��$bC- u�/m�*]��#R�-��tE�JӶ��x+P�KG���8A��0$�JQWVNS����e>V��êT"�/Se���5�rI����8���P���),Cƪ�M\�J�|����}ʂ�.1����Z,vT- J�*}���.Q/�w�'���8)�?9�F6�#:E��J��d�Q(ai��c�\�q�����,{�-�d����Y,��q��
{�8�B�,$��4h��<H�
���Y�Rb�|F#^�wP[��G]��������<Ǉ?B��P�ȅ�!�G��Q�!�da��$�1��!���h^y�4[�]�+�!6y��\���Y�
>����ܢFԈ�YmCJ~���B����J4<^���2[�]�}�б�DSV|5!h0�R׷��J��3`^���jd��Lt����8PuQt��g2�H�`�V�ȋ� �9�p؅Ʋ'�Q�
u�8�B�0`	����˅��Ļ	4<^W�[�`]�E@evz�#�Ň�����7>#����7w�u���T�j%S��`��Bu	�`DTA�yWj�_�[����v�Pj/�wSJ��N���F�'�:]2����U�O�Ez� ��S��K��=1*�NV�%L*ԁ�ta�6��Ȣ��DQ`�ޜ�A�_22�^UÙ�W2:�Z���cB�h<��V��@;��eH<���TGʐ�`[�I�h�UA�ԧ����d̩���s:;�L����O�E�nm�*d%{b�<���	Rt�h�m���a �.�9tqV���N0�p2 C(h�Z/�|U���^��7iV�R�R`�D�� �tN�U�-p�{���b�0|�7����(�MO���$����l�>1��k��`�ٝ���k�@[bX�ג�����4�R�!%��j$PY.J���ro�9P�����=�~"�׎��F@	P��yx��SW�Hi ~�8��0��@;�-|�9�Kvw����'���NL>R��S>4��eF�hk�3ct����O����ЉW���"��/�����4�t�N�׿~�
����*PR[�TX��jf��N��ѣ�ڂǆL���2<:͎��ߞ����@_��Ʒ�p'Sbk�6�@|��:����#.�<B���`/�@w�-QL �.G;�y;�rL�	_[����~p���)�^A�����@V�$��t�#�<��q�h�J*(�qF�PLJZ.�0M�C
�pKH,V"�NW�pO�00��8����PoP�bO^��f_�z�9�7!�)�R Ajd���M/͵l�c�ɧ/���RS�G��	C)PR��6#�E+�R�;/����tk�unu� CUdZ	qH���"� ]VD���T�D24	o$}H��)����
P
 	
����Q�-������'m�~ℤW�S�PYKe�R�;���X��V_*��_e�:��$Nȣk]�.W>�� R-j�����7h۔�ZQ��wM[0���� ��=).��0.�P-Q6�Z������Y����"��\Щ�ŀ/�F_��؝}�<�%�Ƣ�z/��+-����)�)O�5	p�RO�B�t2���!r+؍�$q�Q]��)+y�p�2�uΠ,�m�L�Ŧ��ܠ�#K�b�����QQ�w`/E�:���`*	�VyLfx'`= s��N��O�i���'W5[ۅ/_����	9В�M�RN�q� �������d�l�Qs8 ;����w�G��.P���4�O�����J���n�+:�r���Ɂ�z��e�Q5P%
R�q :�����^��C����Wd���K(ɗ�N��ȵ��q�����[=�(vX^Д$��H��Sh^7R�)�L��	�����!-�^{���(�Pz��D~<؅���Ü��F=��twl*��L-Ɓ��+2�	��2f�",-�%�� ��ud}�@!�W�.���� IW�AJ�|Y
ZT�uP�fdqƄ>AJ�(h�,$��gؖ�4hu3V�t��((U�?$qI�~�$A�3iN�IÞ����BUt�<��(~�+P�餷��(s6BU_I@��Dw~
r���p1@�0A���r�,�	��/݋f�ѽ�7�Vfj_�R,l,-�J�K����C��/Ts}���[�^�5����V	H�f���|���5 ��W�qǃ<uH�do�������ɢAu<���'�����-4B���֠	�	;u%���*�_�+�dW�!��w���p���Q�J�$_����K9|Ķt��"�V��(�c�SX$d^�^Qh�NZ�TL�\���r�.�t�^�?�i�qHQ��Q�R$�
0?�
�5J�$�Q1�;��'nY�e������{�@*I�UQլ�C����9t;�N�ː���&V)B3�F-��zYKʉt�V��x����ml�;���1��a���yr��d1�>w��^Ф�����&_yG��=������Lh�� DJ��bZ�_�IZ���Z���U�IS��^�S����PR�罥�|�\=��ۅ���_�e��'QPB��+j�qr�lTM�jPp�H��h�M�k���RM��tj2S������������0vh�dٜ�b�k^����^�	�v�	!)PeMB��b)},��8�B�זۚ�IK?����*�L�"��FQ�����N�𼇗V¡�(�/-��m�bN_��V N_��^�xEEF+0!�),�W%W�&A���T�H�2xbvHt�;˫�tK����Z�m��(g�e�tbJ�Hfm�U�T�Pu'�דK*;�J���t4�.?!N�Q�SW�KJ�\F0���,"��,D��ʲzL�B�QU��3���W���5����sa	wP) Xc-��R���$�\�@�W	l�����1����DJ@R�nu^�A��������xQ���[sĂ��xbɥ��2�	�$�H��c2@"l�	�)�:��&C� ��0C�ѻ�\�P�z{�a�9B$g��Ǎ$}�S��U��TJ�����oU���r��Q�)�OĴ�
$�5(F"��CSM>�.�~+�,�K�y*��O:��S��>��
��Ԑze���9t�m*-VQQ	II���_(�%��@�h�Eʠ�t�t.�;(��KW[�S�� ����_JuE�8@�ri�u/�j�N�&�p|E����,�-'}D���,�4,�è��e��2V�Cr�E����KV2��$��U�C�͚����X��sT�3���
�t/F�|�"*N&鎋V�q��p��z_�ޡ΃������-��u'$�e�/�?N��p�T��0��z��Q�_]5�.��^��bT&�r���a�n���<��~J���+�������/�E3T� ��B��X|��C��;fs���{��J�<j#2x&PE|�T�=ݠ�w}to�=yH/�/-�W�PJ_鑣�Y�dh��g��zd\��s=-;�Ѝ�4�
����~(��f!<�QQ��es'�W��/��.wO���gp�:��j.Y!l
���Ս'�M�H��s�u	�y�f�E	DQu��PR� `>�l'\r�jd��� 3 �K�$C6����i�����c�ִw��;%��-h��[�3_lZ-�!�3�~�x�~4" �9$�u46ɅE�"���C�����}�J�扈T9�Q,O�<���O�#�����`tF�U f��K�	u\=�pFT�tZ��,�ط�_P�A��w���'�j��`x�Nh��Fh���7�SSJ ��Fl��<���������7��Qpא��$�ϝ��L� �
$���~h�Nf<Z��gQ�(�R.)D@�l ;HP��9~T�^X�]H8��.��l��$�)\Q�"�� 6hf$��
F`�\�<Z7dR�S'��\P��`��28L<�|R��FDFE��B0V;@��r�˅�F,�6�9,`�Q��R��<��F��!-�g/�؍I�i f�	��t��h�� ��� V��(�l��Ӂ�VP@���y�D�HQa�=�XP��[�!Z��>Q6VP\��	�+<����O�� ����E� e��P"�����5fuH%oھAC�:t�7�~�A^(����;؉�C�a&��S&�u�ɼM�Q�@hׂ�z ��n��ǳ���Z~D�<+ÔnX��	 ���j��N�F�Dc R���g�.P$����T�-~Da�N�t�'��΃;U��@�4��}�QЉJ,�>�O�?ɷ�Tn�x2��;�|ʁW���~_B�,c��� ����I#�� 0��S`V�0}�M�MH)n�a8;�|�NX��M�~�3���؝�ȉ'�#�B+"��<;�"	����a\�@)�����&{��_�~�rs��O�l�7(+es-�;`�ե�r�P[We��b{h�3��	�� 	��q#��E��3��v��쭱�$S8��3��� �0f�%w��j������)������Ô<*��COf��nyQ_�Ύ���o h$x���a�'����M�ы�|z�����|U����:�����~yfkwvB�B_�}I�A��@��%�$Q�@���LHe��C�2R>�l����2��
�����
~��m�Vm-j��H�J��Mu�訆���/5� ���8G+:�2*)(p.�-�,8/R)�4 �	;�d�����bެQXb�S�ס'�~p�.�Cadf+�0����(�x�
Kd+��7��igEfbPB�_�������[��S�S<'��j�#�N��<�CH�C�f�M��kPJ;�)�z�v!�Q��HRPB��� �S�`�щY�J5^F��=r�6S�4{H�}H�l�!J���[��pӬ�B�2s<Q�V�VHN�`�A`�@S��l�Ih��+�:�L�&��D��-e
�}@t��@!�؄�t��s�K.P%�v�!D���h;��l��W;8�$
C�&a�(�	,�\e4��0��D��32/u v�t6fɪ*�DB]`�}�uLW�E	TҾ�xz;3U�h4��*8<E��uf�+�?�5��	���?���}�����j��h�]��X"}RWV<A�,e6Y��FH�[A��)��~׽��EQ&�	����.��p�	l�t���8�Lfh�ĕ���dp�Qſ����t7|���bLud�Jx��% S������',b˲!U%�M� UR�~�!���J���Mj���A� ?}a���Ɛ^Uh/�s�_�4�Ft�E$��rI28(�c�7 	+��pq�8IӢp!T��6�2�4d�@(h�B�}̌�F�4/�=��2�ya!
D,�	V�I����T�C !(�$Z� �����|J�ER�Q�ykd���P���/
-�%{D'��'jd�$G��[�t�ZQ�J��Ét�ߘ0vн2�u�褹ZQ� K��7y�h:VQ�Y�˖U�Rj�����d�zo
u��5�p���j�K�%q俽�	N�Y�Q�J�j�j��B��)A�,�J��) �Ww��HI�Q_��a���*ɘ0���5�~L�����G�Æ��:�)��@O���/Q���)� ����<=u
?��~�
|iEG�#��(u>iJ@�_�G}~	�����3E$?���M�~D]Jt�=B��[��&�����d�A,H�����XYa�+���/��X$4���cƦ���D�>�K��y��P�:�-��1@ u����	SDTRZ�P��?=PU��E���- ��~'S�����z�0��A;�|�Qe��q�IӗS�V��b�E�w-I���
T(��P2R�)V't�%tZ܀�GW�mf~[���.j:��P�v�=��%ݪ�m�=j|U%��	�Й���E\�I�ƈ (|.ۉJU��F>�V22uX%S��B;"]�(>TS8(�Jl��ؒ(�<�;4{@�B�'^p��w��l�u�+�=AB8-u"�h�I�V=���:�0�ThԢ0E�K�$��
�0'ԟ3P���Q��2R�Qd�i�ϓ��+]v'Q�F����i���<��CJ@�*$yD��2�۴%JW���W�T�P�D_���x�c���e �s-�V��D�D�R՝Ľ��llh(�Ё�t�s͈��+έ���!Z�'n�,�I<(�8;ĝ!�l��mԔȁ�5�:"U�Z��+_#@�� �\m'�MZfK*h��'����m�+��[��KQn�m�:���<�?���@�P�nV%3����{j�P�@�dHQ�E}�#ؕ��t	
|�܆���^ؠVBWN��젋�^^��%�y�$̔J�2t#RWl�q;�K������b�ST5!� �v�0��@��2�,�u�$�W�}�q^����!�&�	�$�w�w��W�]�@�(��'bNw���w�2$����ӳ���"3�R=�y��&Gc���>��q�� ���������D�U�Ku�$�̡2�?�h �f��6���!E�;��M'���!�1�Y�D����[�����-Q�7���=KW��A��W�{�p��I1F�1WU(g�CJT!ˢW��'b�2)�X�D7�S_>�[��ç@Z��5N��sDRhK�"���߲�ߚ:��WD�v�(f�8MZuC�H<5�����6��~�����&T���Pt�
�3e�u�KFG.Q'�����2q��W��(P���	�SP��x��8eg݈�H%�X�'�~}�Y�B��ξ	�9B�!Y����E����Q�t-Pf~����be���u1.c�l��C%��
/�	  0+]�1,;ݲ��|���t[G��;�r�P�I��x^0� �Q]+K¤fÝ��T_���&��HE�v<�Q"���/-�����Ǵ(��a&p�=����虓`�@���MSQ�� NzR�$J��_���H������ �HN��&�:b�R֐bh ��W�%�6�+�j�X���n��'�y*�@,W�y�T�>�D�+j�fB���;�8s97�(7�+�	m ��N�>P4��Rc7dN��B8�Cs.r�j���V��I@W�k�����5=�^� ʷ� 8DY:�t�%��)ߛ�H�¬_�YMTD2��>'[�J��wm��Vu�S='?�M�%��k��2dWn�1׹p��u堸�P�d��� ��%�
T�`9�/���P 4�r�e�Ra	�\�s��R��B�E�ՂR�&pE�/���y�i!v�	2�7#b3#	lq
f.?"yD��N\��K�kp^��gi vkQ�¹  ��Q�躅����(:�A/�[&4�;�8%uMt�jfF}��ޕ3y^��j����dE�tjA���=\<e�!<���[ꮈV�u匎t7�)����aZRP(��׋��/s�ŕKbXޕy�z��E�c�d
g U��c2�>bV��~!�*B�D�V�|_:�K���FAo�7!�{�F�J�����+�l��2�r
�_��U�u���;ǥ}����bAK`���D4�Z��;u�*��ܵΨ���~� �M�hxE���(0)HD��6W'W�E�<��G�4W��Ia��*_ZpD���R��,k3��R�P,� �%�P�[L������u��(;�H��@q�yE� ��H�M��}@��2RQ��"��JB�%i��=.E؃�`�I��H�1i8:4d���/��}u���QLUA�O3->��H�+�FVU�����R��ȀA��s�P*�QbR�/N�_"��j�!R�
�Q{D���0t�+������r��؍E��/M\�+� ��]I7�*QȐ]!(	U�``dR�>��i��	�q��z𻚚�WT�28�Vvo�֣�iB�୧�X���6��$�}>�j���>_�<���,@����%��%}
E�P�����
t�⫗+�W1h��"j<�aG�	����^U�h$\d&��3�Yav��wb�d���u'`�E;X�S��T��\�i�FbPƆ�S)Q�`e`E� ����d�.��!��n/&8D�x	�\=��w�j�$�E̣�eE��I��qS��5��/={�"�t�A��y
u�^耭,p[�A(Q�-}8o#Ӈ�R��^�e� g�T9�e�/�� ���Ki�s 7H�Bw+W$�H�����N��ϐ"Rn�*'�]D�R�B��A�A6]a�%O� �N��1��X	t�$GR�<��%s�ڽ�\��^���~�i��P;m���\�i0
]�!�a/�+��7"d���pJ�yEo(��*t%HA��B���/�s:	E�P�i@/�}���v�4<@P�ҧ'���0%�0s���+����E}a0SUKV�т�7���=3��;���H~+!87�[���{��EN�mK��2B� 2E;�|�FV���'�|���p�r'~_�K�*%W/�V�|WS]}>3@>Ȼ���a-�(�fVH^�F�u�+�S��:*�+���W�IC�7x��v�2n,��H���˖�B@�sYD<�QS�4Eu�!$�Z�D\��H���v4U*�\.���"@x���'t�ZߡP�r�W��~H"Q�o-nw�����$�A�?��8g,���I���MJ��<��>=9fR��H����RpV谾��b���4_���8HZ�}�(����2�Z8EA�-��u��'z�!���kW��L��@�[e4��O�����0�_k5��٨s�N�U�k{� �Y���!٪Q�p8�U�2�_A >��>��n�44N��&P'�\��#�A�<0�Ѣ|��5ܜh_N���[֝fU�6��D=9'�IA4;$�e^#sK�E�BSu�u�
!�r]}dC�u�s��`i|V0M(_��c���;����]E�[ �����v���
�R�p�� �`��'��A$��Q{%��'.(8tLGj��#�%v�E�`���H>���dqԐ-�Y��؊dI��u�If�8 �NS�Z���#W���	
� #�z�N42,u0<�-_ܢ���jm�(�,QY�2;J�n�S`P��kB�7«NO��}
��W���pd5�
�Au�G���j�b�����1�(KQ�w'�APh@��P.�Wkt�B�K� �@QcrP?ZS��|�U^0��IX�b@P�F�A
8�4����<�O�p�4�������_��|�V��,ZV݊zs�/*s�3(x-��W'Di( Q9QR���i7dz2(�s�_R��INk�
_�0��@��^[K�h�@�8'
fi��@��6ER�J�d1-�ٍ~�SW�9�	+���m���u�H0�#�ݝ��VQ��P
u�k��Z�@-l�W�8�$�HP� �gQ-V��e����V�"l}�U�U���u�a���:��@2�뺸�+��D�W�4u������*@�؁�����.P[*]�;��0��Eа�.S��yd�0�ZjA�M��Yׂ��UT=/�lE�ȼ9~G�dp牵��-�ڒ���m5*/���
C�����Z���R=D
���B%@M̰*Q�.|"���L��Y����r��z�w���tW�������FcQA�<�+/KN�}Z5ЉW�'�����zp��vg�u�{��Q	����"`�ju�����"��;��K[���eW�,X��b�
�-�/ZH�H���bP}1�~�M�ڊ�8��~KI��rR���(�P�pV H蔪$�I�T����e䏽���l��6=�#�n�6x�_�X�+��e�Õ����#�ˉ�Qc%^��-����)IG��|��_T�H�e�h�@Yj�j�2��"�E
%C���W'aFdϱ�O���ÒR�VV��h��x+�;����%.Il��8��Lp��̡�V���t�F�d2��0�k�K�8P��`�G�4�=������d��R�A9"���O;��biW�f��	�`t�T�����fi��]'(u��'=X^;��MvEvo�-R�>#F"P�PQdVb)^��3[�L��qY�_o�>)�
��N�߄�=;md*�A�.ڠK�K�Kb�E�sZ)8�1�iH��W�x.���2����%��K\��N�ZR�]���:)6���i�2����V��3a�����ڈ^)P�d�-!=���8Bu�G�1!t�,�[������,���q0"�[�c,�H-]+�	3�Lz1TkS$h
����C���7����4YK?VLbH��,9�z�.�f��Sd=	�Fhh���6��S�h��9r9P��}XSh{�.���'j�>�sRS��eN Q����]j�8�~�V�0�j,hW��,�3�����h2#�D5dR�g�'�J�i�����}��UL�#p�&�xvKF%�BY�m�~�K��&��Ј�\T>j��^KFP��:�N[Q�wM0���P�� j)�\��-�*>=/E��p��.�
��Fb�!�B���7\~(R߽9���'�G�tYdCx3V����>ߜ���!���[x�I�hQg�����u
E�T���ݐR��Xr��3��D�_���D;oS1��Z��a�o��(Œ+J=�s,sn��J��^����؄u�L�E[�'%u`����p\���5���}��[{ݑq9��^���k�j܍���Ѓ-\�d��F��̅��9��%D����H�L�(�,d024%�V@8�H���($%<��Kפ�SOj8r�-h����T�F>��K�̬8�%��䥕�BG?�N��'�d��*et�	t�aQ���%�pMJ�݃	R�P8R��-���3��Ȝ��/k��V��<-T@��|��)���l#(��2<9@�%{W1dGI�.e
p	��L Q�dB�^[T�ω)�@$!, rW�ncQ��P{�z�O5!a�s 3�;���H���+�P �qR������1�@iD���#]N#��J��}`, E�A&F,�N�L*|�
V�/�&V�i�
�(��Vd$��U�����+;���G��Z:���!�28�,�%;��qCm� ~cru
z�����(97$��|E�!�;�jV V�P��P=����:;x�V�z}*�����@��u�|[�
VOA�J�J� �Q���Py�����ȝZ-4�ǉAP99z���L��opS%�sLjl�j�����N�lPE *Q&j��Wg�%q�W�3�16�D��p>���y�����N��K�#������R��d�!��������e�Ij���"AM`����-	6@e��B���tǅ��;Dv�2�|�G�P�3�R&o
v%q0��|0������H3ɉ��n@��^�]����M�(���C�����N��!yǪW(�ҡ޷��Dh��� �6}d�T$a'��)�H�%W��@�t�G0��u��SVH[!Y�Я[A�F�Fd�FPtA�0D���QV��*�ۋ���
��Q�u)��
&Ɏ���@���&�]4&���	�5�5<C�HB�D;�J�&�Hp�ʉ�:Y
#��|�
te6�3�yM6Hc�v3j�j����V�#���+�n
eɋ�t#e�9�%u�4�4^��P�5V����!8PH�Hll�H
��LPѤ=CV�������(O���_�o�N0^�]�1)]��4t�\P#�AE'ck� IN)��7
���g�`���	Р�E�~"� U�D���1�Ak	�1�	Q �K��^�X4�&�q� �P��aA���V.;�d���`'Ԋ:��+������;�u
��G �6Wx(zǔ�o�s��<yX~LT/Ei5#��;�}� ��۹�_�Q|��
	��u����X�
L�vyl��4��Q(����N�y0���h�׆��~� �d������b�w@�n�g��?��^(��t>끹K �H�:��E�U�,��X�2Dh1L�0�����H��PIO((Qa��vF0�>�~N  NDv8�QRe<�SJ����S�PDa-���0҄��O��IP��0��dM8HF<,?��;�[��FkY]QH�d�����,莐�#H@ܖP�GN|�4/C$��W�G���K��Y]6b#�/P�T;�Vta�p��Z9H| gU
$�P��k�&�,�`n�&�@��}����!��a�*�6V0�� �����\����V��4|�Ds[�z��l4:�H�5{���sC��_��;u" �O�h�=��u	6�<E�K�A|��FV���@���}� E�/��nux"4�|�O��>�rH���@v�䌵�G��<dv"������/�,��qq�	+��p�K�"/d�g�S0��1��>Cʻ&�E��F4$�OAIS��R&v&f3�$ ����H�Au; H��4��CK�_��������$ST��l�EQ��Q�1{����H|�Hl@��;�N�KMiJ���d�)R|8�E5���P	ug';���! 3mJ�s�"p�̐��&��B���J��i~�+pL�|�/�\:�#Ͳ�A��G����d�J
-<Pb��ZP�ЏK��XՖ6J!�BtH�k����T��������y��Wu���E=��M0�԰��u�lQ@�����>�"5#��i_��9�A|^�y��V-Z$46�v�dO�X�r �w�%�f�_���V����q�7
�X����+n0q7q���[}:��jђ։�^^;�%W՚\�>�� x��*t�
q����7����PP(�x���A<D�(RLF�@8���[b@*B0�?�pQ:�W�y���H_$���[V������JD�<��04<Wf�t7H�#�z͊ 9	�ٲ7�6��F|	�_����f��{�=Jx�&�����!Ļ�Crd TNl&�c`@^3~t�pX[}�l�ɻ�]	�����5#��u �&w t67
��bkb=�*d�:�J�$T$;P�st;�r?+E��kɨVl|a00�~�+Z����L�eQ�JT���sjԅ ]�hN0D$+�6-��c�e�ȟF�/�Y��_U������H��?g�m-m�9A�t\�6�R�E�$,�����d0U�o���OU�>�����b$���óm%>�k�W�����Kl!��u������;�y����*���0�H$��5)��uq�{0�n4K/�h�h��rCT9+�͉�D�!�<����*�q��T��;�4r("�Nbv���C8��#@hP�s��*3U`���N��9�'�x)\^��I��y�/r$�"���0P�<���	@��������,Lu#�#����s(��KB"����!rz��K���`�;]�at�a�#W9+7�-;�#T�(M�U0S���q�4<	��mu	�'�[EyHˣ_��^��ŠɲW��)l=��'O ��c!%J�)���D<BPA�L@�dPȲ~H0�L���		N<#���@t�O,8#�!r�Vf�},!��PT�'r��:u�U�i.�W�%��㳒XsH��LM𖘴D���T�Ȑ�F:+h���X��DU�E�h( �*�6�GB�F��3�q���JfքjA�=��đDs��Dو5�Dh�^�m�3�)�q���%h1B��� �P��,xp(N� �+�;�wC��:YؤSX�P�~7@B\�B=
:�P��?3�%IZD N��&P@wV���hJ�Nu��쟱x�A�1�Pǵ81(���J�BNb"�n���H��Q�h����fǸ�����X�K��MVF	�OE�����*�Afl*Rz�I;%��r�������]N��(�	����~�H�,�,���4#w�@tq�P\�۹ioX߸��I�.�������\_��K�]��e_���D]6*�ҟ�9����m(�w��Gt��A=OoUk'%�������˰A0;�)v	+ց�|�b�߹(��)���1�(�����-�;�r�X�n��X30 ve���W^0���8*�V��̣(����!�����
B��AE�|o��$�uCY	�B1�(Q
!D(-;��9э���(+��D;�~ ;�wh���}4�
��t�GS(�(W�LG�%����4PU;�v.�u�̿1! ;!�����i��`�K�͐c����4�5M���z9���!qL03ۊ\be.æ]�Xh�xRgpX\gn�t!sx���sO*�>9�K���q���w!��/t%���h	+ʁ�գ�ve�Rp�慉9�j��| dl�Np򞱝���f�x��\̘��]H� .S��<�����H�l	���p��ۘ�\��X�LH-�z**�],�I
3++��7<��Hƥu�!��A�`I
I�ǂ��*@VҌB�Qo{��!@>I/[��X�!Aet�E��?��%4*D��+#Q��,B�)�x���u2���hc[��2�NlBI��a-1J���{IN�9AH�EVz��+��׍t\�5���r$QH�d�b
����@��R+��$A!�+�����~���[���4d0�i#�:���Q��[��K���^�$��&I���\~~�H�9�uܼ�G(�y�s.>�3P�Q�^3�('�D��4��/�8��٤ tK�#���<��G0+܆S�Bj���t8������O(h�j^jQA7;a:	�:�VRd��)Z���eS�Pg)إ^��YQ+?V�4��O�xZ_AN8X��[�ɑ�Ɖ$��'������UQ�n
*C�k�X�K4���C0V	�WW�� ,Ds+�H��,h?���`�<Aj��p�tt�s�}��F�.=CH���)*L�'x3������Ge��sbar���	�ƃ��.�������>K2w�ɘ/����S�q0�:�����+Q�@�l-9@�H�|����OX4Q�<P3.\8�n�E�F�<Q�R��P�G.)(N�ȅ� �д��o��п�E�� �%Qm*3�� s_,���"�؞�0ÊO��|�@QHbrԋք��Ҽ�Ӡf3
���9��;����*�*���Q�s��z�'��?��?����,P�D;�/u%��s(������-�+�HHUL�X�f`�m*uq��HPWS��4�6h7��p0�xT֢L�9��$hI��Kx� �=a�> u"���/�����N^*��e Z�e�5R5$a(;�|�}���/�z?D��U��ZK��+Нy��=�LDpi��+���}FJdD��.	gH�C�$C�/!V����s6����$�>��N����qt�@�e��Ҧ%�?A�ܾ������R�.���;��!(k0xHj���p�!&�/��O����S��cG��C���>�R�ABD�׎�
���;�sn�U8�$PD�"��I=Jb�B�E��)���H�-d�ǔ����8�YS6�<4����n���nri�c��p�h!{5Qǩd)�m�qBr�$V1�KFC./QP�ǅ����-R}�T���P��Pl�^� C���(.�(4D��ϴ��QI���s��B�1JJ�C�a�
&�oS�P	�4An�)r����)�Y��JҊT|�Q��lD�@���F�4s�+���P��|8@�ڈR��t�H����L[������@;�sC���H�ۅ~r�E-�������#��F*��C�㚐 H�i�
�.P�
�ă�I���z!�4/	$�����%����X��[Po�D�@Ř��x'?Ru�J����Z�����u�t2K$GV]�T@�R<�
,0F��Ȱ��r�CAR�)	�6��	�"@v�L1�aEmW�t�"�VR�B(�#�K�E�5�n7���7O��$��v{ �k ,>��nVfc+��"�L\6C�P�s�*w`H)���4Q�8TB	+%X6K4��֤&�$j0�%)�mO4��*�|Ia���|ւH�s���ʨh�X�
����H._�Y��0�8���15�0�?C�BCcOP+��Fj�P(<���L�"	��K���ķOQH_ �j�+��WJ�O�KN�LK�>13iJQ	t�+�UJ����U�H,!dvC\���f��A���Lڎ�#IHQ�y��E!�0Q#NK B<0���L���RRR�C��0*!5ĻG�/*w�OP�+��z�NLRW�H0GUMp!n�F�A��R���d+H��4�T��A��d���MS��P��/��L��B�C��ҙCP]��h�1��|M��K���5��B�	��_�ZSx��dл1g+�cUr���@_QV���"���;�S�8���?�.�9�\����hUd�C��L
V�L?T�T��DK����/�|T�U����PH�B
5.�V�,��!�b�-�<�F�Z�cD�ͱa,|+"$}�]ċ�h���t7R��ˆ4 �.���>+��n�DY�P�s�g��՚j	�.��)8��j��V򰑿�F-��<���)�����e��D�T9LSo���w��HD�,6�p� �� �1]���5��m�:��$�LXIv�	Ո��'�p����r���%���G([l��W̆�&�,��Y#@�+���J�D�����W�t���U����u�r�	+������7����@������Y��ƿ0V����B��Q�
!�D�(����xQ�
!�D�(�����/MepN���&F�(Hu��EM��N���
>�	;�m�����%�I=]�0[��_�;�0Q_01��?� �85��6�g�k��P���Sِ;Op���tB
"(3�ǀ.pG��� $"��0��1fZ�C3��!�24�dp�ʰ�T���������`��Iu��F8����9ತ�t����2�#f� �˶^V �4���~b��؛��%��X
Wf	��O�p��@	�1���NӦ�#F��7�X*��DA�f��+<�_��R�E^[
��B�hb4��B��L�E��g�T�Sl��Ҏ����V�&X�B�*���N�P�����	�]6@%��J؆E �(ȺS��A�	ݖL�ڴ��C�E hf��
��r��w�Sȡ�~^�����2���~A4�9��^�PG���);��g4��ύTP�袈1����#�/a0J�vL�U�+Ѻ�����		�%�3�*U���ǆ$'��:V������_��30�W�|��~P��u	z/ō���>>�V�#�Q"��|�B�����	�
|����xv;�w낍M��}���F�%t � WUSɄz_��mE�^Y@`���/"� HɍG~Z�54ȖdV,��B��I@���D6�$�2��I�5�/�hP����
����S���WI������v�Ё@���6+72C�������)'���2T �G��^�T��	@P�� A2D~d���؆��}L(@��e��̕��nѱ�n�-[�O=�w�8�Ã�����'�D�s"l4�Hq�7L,= �~>��f�p:�j�A.O�As����T����0P �f�%BQ��@���)|�6(>}]X�
EJ��)AA�n2��LW[J�\R	3�L�	���iT"�Y)|��-\�K}��e��z������|S�?�#�0K#}�V���LE2B�X��j@����(HV�xX�"����LB)�=�JvU�2���h]	��A���џ�����I�܌.�:�-r�/�f'�z;���B����#q�L���k�A��Vt��-(�U�e��Yj�*����0VJ�A�H$R�t�舘_���4^��(��'0�w=��nP*�B��6
������,}4���z7Fy9��	;�r�u�H���ɜ(�wLQm�iK2dZ� /u�(�'v+J�^����Ĵ��z��~�}�@���v�˙�"�;�e��/@K���i�&�Z�b(_�a	hy�>(P�#0���2��DA�ڸ��h�#�@�(�I�f�0���F��R����O�Q�Q�0�@+�f�����0�]*	�	Dd|
|���@;�~�N�G����S�A;�`I� {
B�Lr;0�|T�+��-|<���Ǻp����W�S}�t"{f�Ӎ�X�Y�T5'(Q�E���wQ]o��S����r,�tJ�E�,����Qu
/�H,,9���Bh�62#j���������]��
���j��E�}Ė0tb2�7��M�N�$�1l��](8��p4;ǡ��+�	D��~���ߊ��?}>ʯH\1�u�VW�hO���~'u�t*T��R`n� ��e�V��+�W�=1Qr,@�����N�A�u�jb"|6,�x��N��~`TLQ���!CBP`\�/��L�|U�фZ��������!��-	JKW�� D�/�C�B"(q����h! �J�������v
>u�H`}甀h�@��F��9Q�QS��V�H�%��@ĺ�^��A
�-�Y���fN���'C6U�+3�hK}8�M	G;�� �tn���
f�����}#;?�&֢�Դ?y�d	�#"���R���u�����!�
�����\3o�o�]�K��G ��� /W9����q��@N~�=����9y��'n��E<����"���T]㗋g[�^_��)B���H���li,��~Zo�|����9���FQ�/�ʤ���lN��������h��B^��)~d#Շa��	�ѪZB����]��ZY��H�&	kmb�JĐE0����{��3��DX���ed�=b���.y�0��G�=e�U��o;�Y�B��;щx)�}���x�x�"����_/-
��E���;�~g�����{;����HH�`x���>@X���y%��-ω�[
�T7�HQђL�dʼ6DS�a��)J�&�Y���N����-������]!�°���Bfh���X����~^	��{�%���>���#�#���G�Ҽ����-��
�$�а��y���=�����(�A�'��^F��#��	~@[���F������{�P���ۤ�u'���!�
Q-b�lu�l��Oq�`O�N�5��◫4^�����VW��jpD��#�����oJ�Z� A���ӉL�X��|$�&ľ���	;�~_�t�Ɇ�b��0���P0j�����d�(H��2 ��L:��-��PuTݺd3X�4�-������Px�JXT��I)����в;�~NqW�!D��;if�/H�dX�S$C�Q���뵂$��xˊ�^��$�H��E��$q2ެ+T�2�ml�4��.�J��������R�2x�;��ڲB��L�38��Tȕ�O�_�['s
A��>���������D��r��G��t�H{�+֬�,j�BT�FcBڪSEF��j���hH#!�X�$��ZD�c<�C�#���O�Y��=�X� �O���G�XY��:jBlx�&��?,��ꪚM�Db���}B��`�:3�_8�^]$��FJ�"�W�"ҍ[�V Q�����Iu�U2B�"y�ĝ23�<(���2[]}�����E+ƁB1��H��;�_���C��%O�/h�V�`�������J �y��^ã�]��u@J:Ń�VW������/s���������|F4�D�PB7�h2hub���;tPYVv���~?�L!���";�~�lL��2u�ӕ^,�������zɃ�ǆ��tI�,ň�������&��A��Tf��"��a�>G�Ֆ:����k��H���e��BO��-:`6C@ZI�5u�[���G��j,`H�PR%P ��At"�����P���H��-�1h����v�z� n�D���L�O/��?�$N0���2�D��=s��EN�A�N���+���2��WZv!��3�
-���Κ���%��kŭ��z�V/Ȥ�� }���T�uQR�J��9�Ǆ���hA�
�#@<_+���V,���Y�
t�DH�3��T����DL�Y�:H��N�&8����;؅�s8���|K�H]�f���(E������nKR�Eq2+ru��%�#6ۨ���	W�����Y#���+�D?K����K���U�Wn���2���U��IWf� J�r$�@u";�Q���ȦL�P���L Aқ�1%�8D����G��J��E��"��$�uQ�>�+�W�?(s�ZNp����0���l���.�Z�VC���x�CF(;Ȳ�� d�R��"iv6�*@�rh�|H��H��8�N6<���'F,�8u#�?4[��4�(�=�H;͠����c��;�cRP_�Tc
8YsmkgT!,�;�n�T[�V�Y���%���BBE,�	�J�BA���IV[c;�uE��0������k�>���	뎹�
��P�
��SB�G���Έ	�G�v�@Lqk�5.;.8G��+�(8.���/�$��(R얡�6CCN"���5�	BNL�f̀�Ʀj��PWM/cV����yIv���9,QWH;����vQ<��%AM�X�xx�i��Ned��
SL��NU@�g�[P�_�G�hQ?
�e�4���F��/� ��
+�8hp�F�ȍ��sN�$�)な�	W������'	.	UQ��PN7����QSr� j��u��r���uK	����5��$$��ӯIS��0U;��0Q�[�B�v�%��v�W	SR�GYvi_A<_��>�t�}�ZuA �XK��{E1*Z� �{��Yr�^�f�� �.�T	X�\`$dHh�l"pDtx��Ǽ��+#����ĐE��  �T�`DEJ�(u�9t����E��y��9K:~�b�Ē��'�M�	�@v��K+�^98!JRb��v�&��s�dQ��^���w 9>uJ��;�����,v�L��+��0�s�\�T�3x%����%r�����C�\��1+�n�fy.�ّ���H䘻�X�:t��LX@���Au�E�6Y4�k�`Ϩ�tg#,�-?Rv8'������<�B&"d�9C;�r�'C����7!��Y&���=*�,��8�_�����,5@�	<�����1����$����;	�J��'��4�Q�/�A+����eB9P�	pl�4DA�B�ͼ/�,�T�H;���t�JP	��w����q@������(�HA��}U���A$+�'r틬�s�R=��b0�<�/��Z6�s�����8�UR����܅���L�D�xLt>3�?�@�U$*˃�����و218�����J�#}0.��=:�����t��ʧg���ݱ$�U��\��T��*ӈ�1�L��7�k��ƀZ0��I�u��;�s�M�Ҁ���a`k0� ��C������ �>E4�"T"���SS\�$��Q�{�<s!��@�U��{�݉)�,ՙĉq�!r� p���t3���vu��_NW�&�쌑����PAM#�A�t ��J+ݚ+�}Y��jTh>�1�Hi��]���o��_ �L@k�K�B_�`o!B��D%���	��y��Hx�L�d�S'sxz���,ѸC(o�h/ ~1�3S��:��8w4��JHuWC4R/,P�h`�\��U�����(;��ӦGp8���^�!M�(I�8O��#0z�D�ɥV ��RQ�R�L�u$(�:<���k
w[�I��S�u��W�3�K0Q�C�Y����P�uB����H$��td?�)0y$gSRH\^�CB<�+F$�����=�K�ꉑ��<��m#�����%���W��[Q�-!�k4JW��F;���Iwv,,�$+b�N�a	4 ��j�p�V+�4ՉJ��C8� �K<U��Љ�~ɐhx-���n���Vź�CK|,M��j���C�(%#�u���MQ�+�>���W�G�DV8G�ă���1�����b9����e�$3�QlC�']>����f,[[(�O�@~Q @Nq0�J*y4V	A;�t#�s	+�NQ���I|,^�b�(�2kSE�I���s#�)o)R4QM�`�� ����E�?rᴎ�²0#��a=΍4r�Iu�k�;hN���+��(��u9_
�K�Н�^�n�9q~�tǃ���5eN5,t�ꡇ_��Y 4��d11,���ϊ]�0&["�B�.�dFED��>rک,U ���#����y���$�!����g8]z�sY�m,�u�+��?r�����;v!t ��GFMul��^vR("I���V^$���7?9R���J�GtZ�r:h�
�3%���<~�=q�A��O%'�����b��ܩX\>�t.m�(����;��q�)8���S �i�O��$�2*Wps[�A��.�X��~{4�-Y@� tV�Xܝv�Ͷ�!��r"�{�g�2�0�զifXA�߂1�')��g��Cn���%H�b�� �D�V�؝X����2ρY���D�(��>���@s
u 	����-xK��zz�z���P2�Q=+�y>��r��P�-���s�"����kPýy?�u9�`��~.�C��xL�zcP	�۴#u?h��|�1`Y���@��f�p P�h7@����Q�0VY��=��9'ct0@�"V�q�;�r��H���[���P"�l�%��Y^j�X���PZXSX$Eu�-}ڔ	�=`p'�&�ɘ
u"��e�	}��Б��ꐱ�NƎ0i�Eؚ17WcP(��(I�G�p�%��5�!L�P}�tV\!�{�_��]�����2�l�p2t�����!�|*�T�*���Sܴ�֋*�\��s���1,��?T"�� fҒj�M@-�# =B�A�tz�noX�B[���?L�B@ nHU��1a�@B�!ep���MP��@�ٸ������A��#��F��cH�D�Q�#J�3U��%�S��W�4�h!�m��� ���
�!�5ԁ&f*8��R �z!A�F��Dg D&�u� BJ�$P"CU!,�_�����,5������ƽ(�
E�N�Y 
8D��'�� !w�Cl�ai�{6k��+\E���L^��� !�_��Z�HD�GMԇ���H	�>�ʠ�
���q���10�p�}Ax)�d�	P"8D ��(��\'j$�H���"�D�ԉ��&Yd	.HD�T"fDx����$�H̠7/aJG"�E&\vd	H:��)�ґ$L�Y|	`L4�@ @!�	(�6"FDVj�x�$�H���"�D���"&&��f�	Xdj	|H���"�D�Љ��##d�	&H8�T"hDt�̑�	v���&Hii�Z
dT	FH4�$"D�@���$�H���"tDXL�6 $D���"�D�����$tHh�Z"ND8*�
"��H̑�*8�|��`�-�	j"�,vH��+x"(�|*��"	�D����r$�H�fY	fh^	DH�l/�$�	�"
��"�)�`n�QVs4�))���Ď&~	n�Z*$H��%��	�"��	p�ZJ$>H*�""D�@$���i战#���	�"�D��>F`fa"	D:J���$�H���"�Dxj�X��.���	�&���42�	$9H�"Dst�$H�	S /I�(��2��0V8�P?��(@j �t��?�e 0p�[�o/�.�e��C� U1DT\��X��0b�`)j��s��r�����`0@k�����4t`� deflat_1.� Copyrighgt 95-20���JeaznloupOG/i]y��Р�Θ�	����3h�o�1P�
<�1�Ôr .H
P�x���e	v�h���&G	D
�$H�"D�(��+d|���>�d�T�<DS#��	�
r9�����|A�	 
���	DL̉,�$lH�"�D\܉<�$|H��"�DB"�$bH�"�DR҉2�$rH�
"�DJʉ*�$jH�"�DZډ:�$zH��"�DFƉ&�$fH�"�DV։6�$vH��"�DNΉ.�$nH�"�D^މ>�$~H��"�DA��!�$aH�"�DQщ1�$qH�	"�DIɉ)�$iH�"�DYى9�$yH��"�DEŉ%�$eH�"�DUՉ5�$uH��"�DM͉-�$mH�"�D]݉=�$}H���tg��S.�"��3.�"��s.�"��.�"��K.�"��+.�"��k.�"��.�"��[.�"��;.�"��{.�"��.�"��G.�"��'.�"��g.�"��.�"��W.�"��7.�"��w.�"��.�"��O.�"��/.�"��o.�"��.�"��_.�"��?.�"��.�"���@�	 �`"DP0�p$HH(�h"DX8�x$DH$�d"DT4�t2��	C$�H#��"cE��Yx:L��	�$H�"
D�$H�"	E"	D�$H�ar���D�G	#
�|��#�G�(�\Y9���?����� $�J�J�R�\S#���|���>G�?���p��q<��y��
��"D�=�M($0L8	@�P`$pH���"�Z�y8t)l�d�\e02T`�L�M=�Ao�in�,�MarkAdle���Z	8����H�"D#�+3$;HC�S"cDs����$�E�Эh���pi-��\��!1$AHa��"�o��	�$H�"D� $0H@�`�\���L�Tpc0Z�أ������U��TV��<)�� �@S���\��#t�@P��8�x�G�#˔��(@�[4E|�8� dL�鐥xf�(���$�L �)4R��)8XP�� h�P��(��7� �7�@��7�`����H0�D@�# �X�0���QgG�X�Ș�����RHX����E�#hC��U0���C��@����x�p� �C+Ƞ�G@!K��o#`�k��x��?�(.�_8PXF��s��(�E��9�O�#����!�xQc� �� ��..e�HXd�:_�YCP�!8H���h���x#�p �����?� .����P�P�p�����ŭ|(�@&�@<�(�R'���)X�h�<��)��yt��$�D�8�@*P�H�+��(."$S4��@)���`Y��%4,P�()��b/�J(<YH�)|y\O�3�)�x�<��"ط����In9italCzeCr3cS�\oNn��D�ߞ��mV�r�u�"F�en�L��v%��>;Eexr|j�>rA�'JKF��TEd�`A�"3C0s�Ha�VW8zW8�Fo;rSng Obnj���sgr�pya�Re^�U?�@S�Q�	���k�dExfh�fg�'��(�3IoD>o\�np
�P�n��G�P��vV�<of�.��Nam��E��~e@��
.W�dowsDF�S�����DLib�a ���T�Ad�.Is�y�6�a�M �a�Mul�|B��To��!P�ra�Y�* �+��mp�����8,�9�GV?�s����"�9�F�KbNx�����KC0D@��yepEF_�sk�ASpa�NFT�Vo$lu(_Qf��a"o0��$g�HE��3��U�!M֢��Mc:���N�xt��T�RsrЭ �7!G$"2 �I�m�V�x�[��.MS�pWO�B?7�a�dPFSPof%L$��l��+�]C�C�6)hؔa�ErYoQ�t� Sy�C��V�S�i#bu��:ȡT�RpP�hЍDA��yTh�d���z�lB�$TRkCoud�Ijd�e*mJ�u3bd�l�0ͩ�(BbNc���,UnL ��TLꎬQS�S;XzC�r�d�p��7���23ipA���cC��S�"d�F9�'YcT�
�k$QxbԒ2�p��1U=D|�������Fc(B�ߚ2����vi��(#�"8�l,BZғE�R���kQ&��M�#x kPO�n��Ni��_�\���-!A2(UHhv�%]�F���ME����INP���WtUf(��L
3X2�������SxX e�h�p2S�\�s��$9;�DC�B��1R�r�i�> ��_I�d�E9RN�L�.��8���Yp�tfz���TQ��8�o%T�BpP$K�y��!%6��Iu�%\��H��kE�V�S� Bbd�K9C��2Ear��F�6v6;�PTM�aLg���k�bd_����$M%2Q,�AD�r�p$Ir�?�RfQ��mc�XE �:��"�.�D �SeP%B�~H
�&bGrJ0J0�D��w��Eem�y,&�Hؐ��*G6��	JRi�]s4��I�*c�J#nC���k	Ip;u�*e�2A��EY�	+5�,f�h�"������6H��0���x$�R��{�&HU�6�!\�ښ>��6jM��|�um���2�;�*`y���������{u�PftU�rr�*SxN�D��"��K+��D,`V���D&F��ȶX,US1&.QW����3��2�HDIOB(�-���b#*�)�8'�2|1:�Mbv�a�-�F�ma34<>H~�?LPH�.f�n���4�r�>��V,|iiS/�L%Qu�c2�5ɛ�TA,�,���<R�_v�=<�b�s��o��cy
b,�DM�i8��ngTF�l�Qu�2���f�@?HV>�fSFv����
���i�t��2a`TW4��b^$��hlݫ�5CM�L�r%����S����Ͳ�A�2��$�O�e=d��	N�9!+~r1a�,*�D?�'B����d�r�[C\���qL:�����Adj�ɻJMi8�ZgI�M:�:�k��Hr,5�G���,P��U�5��DsVLP?��4SHM��_c		F�d����kF���!EL�=��ʗ6z4LW�I#3@Y�XP��Z8�1��ҭ����gi��_��%����$Iq8Cx�FL�I,�*��2e�IH�	#�eu2,��D�h���al��"e�he],��V&3b��|Bpz��e�3z=���i��w�<a�b$���x�ͨN�a�%(@�b�^KfDdMSVCRT�"��1t�?_h�1@UAE�XQ��#Y�Q�����a5���08WS2�"���?�T@�y@�$bas!z^'F�DU^"�_x<ns Y2d��V,�&�r)t2�aA�X_N"03-�C(�1�� ul�Z�CA�B����4��)��#N�IQ� ?c��gn�O��V1)�.�R�Gj+�NZ�=I�P�`�fc��T�E���J���s*��2��)��li��qX$�o�`nI1��?np��T�IYB:�P60f�ea��Sur�б�'}`˄�oG�zPR*f�*�K{%+:i:2D�,v@�i�%e5�,��Mlo�i	y":i8qt�t�0����xU�l����"WeNE�	H��3LD�z�w3�Tĭ���Qm�6�8H%p�q�<��pL�Q9G���8��6A�Ie�8��	Y Hb%��F�Z$v�B Y�PS��DL;ѴWT�q���s5���b�9Q.Ž���bZ�8K�����m�!�	Ѕ ��	(2��tbsvb7x��_^�GSDT��!HA�½]��C�8HЕ�N.��D�rd �vO+e:ufgH�%sl\)M�7����ft�N�Lzw�k�e���Fpb� �<wbhe.-`�A�P0Lc�� �	\OB�KD�m�.s D�Z�V�gJ�j�z����'����v��)T�L$_RX�:f΄��dO��s#0A8�d�!U%.4���#�N$�b�%BUID-�4��0\Viv�B%1"�,��Pq�o���c�m�V�Aq.�	$Lg*�TA	�,�QD�|�U��O��҂\\�[��iq�V�����(s�)D�o���k�,t\�/4B�2����	�Rqo��\IGU��R�x� 9-k��%�*|C������ aTyqSrY	TEM\�>/��\�3�ۆ����R�(H�)�DI��y�pg�.Rmp�P
s�(Phg��8Gh0@ >UpM��=���ц����J�|�'7U�!�>�Dm�.
�r}hHv0
[%02/��+:�] (�)H�PU,�B�c+&��G���c*md��� BCDEFGHIJKLMNO��Ҁ UVWXYZabc� �ghijklmn�/q�uvwx yz0123456789+/�(\Dy bSzpr2ws�Gxvf�BKh�58=��������� IEk�<�7.01h��ps:/<)�
~MHz;ARDWXE}s=SC�IPTdONݠ!%0l��̢\ɛKs�;	$.Tl68\�g�)�N'�+J�ӳ\�.��=�;Oa!BIN���d\�CG�w�l��S�buJg�WH(Єhu�p��$^�R)�eT%�pC[Vǝ��a�8# �7�T��$+"�e�� �i(2���n���\*au���$8)�$�`u�0v/_��w���sjO<uok��iF��r<��.c��$��E�4�b��o�g4�<Np���Pq�X
y���Y
�e��ymb���t�.��!0�����Et�����dG T]fXH	D<(�
h�E �sN���g ;yL�djs%8<M$A�<��2�"��{
�m0R��ɒ��j}�w$\V� ��D3��T8p��
pD�d)�K)A���-��/NS�	;�d`K��.�� ]dTsLRA�Sp!02����#A
�`� �7
d�r@� �L@�GX#��2SA;9x8�D�Q�h�G()���#��H ����rT9U+】+�t�4r�9d�G$#��`��D e�r�9\� D�T�S|�G<$ؠ�rl9,��S#��L ����rR9' #��#�r�2r�9b�G"#��Ȃ�Br�;�rZ9��GC#z�:���rj9*��G
#��J���rV9�n�dSA3rv96L@̓ ��f�&r�9��GF#��#^�Ȝ�cr~9>܎G#n�.ȼ�r�9N�� �Qrn ]� �q91�a�!�r9�A�G��Y�r�>Gy#9���i9)�����GI#��Ur$PDxu�G5#��er%9��G�#E���]9���}�=��|m�G-#��ȍ�Mr�>�hM �þ Gs#3���c9#���`G�)C ��| [�G#��{r;9�#k�+ȶ�r�9K���W�~Gw#7���g9'��G#��G���_�G���?r�>Go#/����rO9�= �#������G���?������ȩ�G��?����������G���?���Տ�#��G��?�������#�����?�����#�������������#���Ȼ�G��Ǐ�#������G���?��#���ȟ�G��?��Pb�W�S�fP([@Q��HYDU�A!]@@��X�T"!B\  DR	�Z	��V.��
`@Er��9
#�1a
C@)�Db1F0!Db����W� dy�a�i�v�qs�ԯI9o�'ub���dj(BL��s�GH�$��u��y�h'c\N>��C��)�8�d� ���+�48Mp�?b`��H�"D?��޽[��	?AVtOs�����`�f��?����_`pX�
����l��p����_��g��2]�X:��0CX�����y�4@_
�u)č͕%��l�p�]��!(N�N�˰��L�(��M�;Lx@��'bp��+40Zu~��PP�觉�Q�Qh
T��)
b�H.�'4H?f��(���CO�/��H	�4xN⺘�h����P�Bm�ԗ�<_	�	L޵g!�E����nh�$�T��Y�M�a�2��!%�"3��B�*~��"6�E��p���Jc:�jh`#5膛��h��cřF`�H�PǉU��^<�Ï�E܁[�� �uq�e��j_WYR�@S��My���b��9Pw�����>��� �%�����"����!�9N!�3��rs������@���Dz}�Q%����B�#���F�~��ά��6�	P��\X�Oe��i�cdR�2SD�,l%?��NO�JOZ VW`3�+�v�3�a��(��jY��$s�~8�h���� XW�Fpl�/4D���h�-�Pj"W�VB�$'��|�h�g��c*�W"3 �X�����%$��h��Ưv�FlD�+U��A(��!�0��u��"}�'�d��Z��(vY���Q���Ũ�d	�Hܑ�
" D0D�\n$�P�b��I�e�Ӥd"�mI{ұ�Hg,��n���$�RSD�x%� 6Oq4M�	�tY˔_	e:\w/ �JK�}�^�i386_��.p)dbTj�%?�ٿ~��@N�����_$����t;�{�oM,R(����3���|�E�����	���]&館�t�p�
���~t��IofNC�gR�qwuxs�]Xb:ӌn5NE�d�t�rSu�2*LTkOw56�A��זF"����@��k�@���F��4�hh=���R�l��9UK��*��o0��_���s�r�lw*<��I��4r�t�v�x�z�#5,�:��6'Gg&�-�4�C�L�Q�F�n�y���d7hɬѰ�9rt#v2x;zB�v@��0rtXvjxtz�|�~�1&�w��2'+GvgӇܡ3C�zѓٳ�4rt-v�x�z�|�~�d5p�����ӟ���61'aGgg��ܧ��7G�\�iه�����8r&tPvrx�z�|� 91�[}��:,'�G�a�;���<r�t�v�����I�X�e�r���3?r`t}v�x�z�|�~�u����0ʇ�#gE�˯g15'BGMgV�g�~Ǌ�������2�ɩѯٶ������3r54k]wއ^�ߘ_�߫·[6`'pG{g�����Ǿ�������Z7������!8rdtyv����9w=���>'3G}gÇ�?����T)��PJ���������������������������91H:a;�<�=�>�2N&�I�q	�!l)3G�Mш���94r�M�<<�5$Nb����	�2ZP��=�>�?�?�7nN���ϝ�Oٟ�8VNt��ϰ�Oԏ��9U���:�����;��7�f���9<�:�&=�:H,�S>*NE���?�j]��������壵J0kNw���C1����������������N5�j�{�3+N]�u�(��������4�J�P�[�v������46�&��'�/�9�K�S�g�o�y����������������6C�#�:�U�]�l����I����S���B�V�^�u�z�������)8?�qGWge�q�xǄ��䡓����9!O��������:"'<G\gu����ǿ�s;�ɟ�S<rut3=U�_$>-'4D?�O�V�c�r�~����s?�䟑P"|Iw�:�;�1oN������C
2� �-�4�C�k����������036�B�U�^�n������������$94,:U;h,oZ�*8Q��?�T�a��������p<6r�t�v�I��>�?�?�?�?�?�?�.�8�Ї'7.'DGWg]�o�xǌ�������"8'�A�I�U�l�z����������!�/�C4$^�e�����������09:7:L$^<=z>�?�?�$�$����;��Le�jp�y����������Ɵҟڇ<6'CG�g����������������="�C4dT�[�`��~j~|~�~�~�~�~�~�~�~�~�~�~�~�Y�X?�	>'zug����������?!�J�f٭4���`�}�'0rPt�v�x�z�	1�=��26'hGtaR3X�\�`�d���l�p�t�x�����4axV�\�c�n�������d\(96w:�;�.����6�A�����ĺ~�~�.8�$P<H�XgRjb������9KL<B=X.�М'�Nx�|Ο�ݓ�Nb�C
<��ȓ���n��P?]_�;�~��p�w�y0rt�1/�;p�|Ǖ��9O:\;�<�3"N0�G؞����4E'^GrgÇϧ��56L"tvDx�"�e`���O��t|v�x�z�i9���˞�݇M:V$]���ò����H�0;rvQ��A�\�e�l�����!e`�`������;9?\:u;{<�=�.���_"�H� 0r5t\vcx�K�J�ϛϢ�����N��#(O-�7�<�R�W�d*���S�����������I�m�|ٖ������������3r	��.,�%K��e4�ɰѽS������H�{�M�h�|ӄ�����������6����H|/JN8b�m�t�A����d2��97-:C$��Y����8J+�h',p��Ǣ�����D-9J������9:E:P;W$j>��;G'�G�g���+<P�W�hْ�������4�9=(:/;q<x=�>�?�?�?�>%NF�zϣ�C?� �+���'��06��GZd�����X$1x*���D2K'^E��D����
3���F�ZÅӍ�����X2~�45�SX�`u����̀r[5e������O6f%r�<���*J�
P2t?v�x�z�r9|�����ٟ�:�'�G�g�����������;�<��7P�c>����,���|t� ~�12������~$~(\,�Y�?8?<?�?�?�L�Lt)6MN���9QN`�où=ۓ���'���@�6T7��r�\�jH�>)?3��:�uL06MƎ|π	��$�����������dڀ���q7!�8�0�:rZ�s%KЄF1�X*;㐦�<��=�L���Do1{2C3�4�67�8���P x�Y�6?�?�?�W9w8'��A?L�kъٳ����H����0��.1��2QN��*�|$�B�Hj�"�Xҡ~��h�:;%<*"/D?V�k�xM}�&���*�0I�<a�H�N�A
Z�`�f�l�r(�%�����8,�E�J4�m���~~�~�~�97����O�����:)�AX��L�4N� �$0Y8�<�Uc5�H�Lp�MT6&\8�p�t�x�|�ȟԟ�����5�ZG(o�7��� �1���������zL|TY`�?�?�,����K����.��DP��xI��,�?�$�n��6 ��Ed�䨙���Rr�pDgL�X�t�ڈ��'�������� �<@�0Yh�>�'���������N@D�P�X$4|�H�����P�~�I8gTn@�؎�(����`�y܎���� ��ϑ��p7t��pDx���'YX0:�������                                                                                                                                                                                                                                                                                                                                                                          �8:ˇ*�Z� �/�!�UG�&�
<:�0�ެ*>�d�AY&�21A�!�����W0i                                                                                                                                                                                                                                                                                                                                                                                                                                                                    &8�'��9� I�]�Y�.Ff7�SV��{�$�2@�vT����&!�A&VT���&fC	�b&�                                                                                                                                                                                                                                                                                                                                                                                                                                                           8����? u�a�e�zJ87�Sj:��G��|�Jh����&!�҈�Aj8h�Ω&ZC5�bm�#�b�&�                                                                                                                                                                                                                                                                                                                                                                                                                                                    T8�U��K�q ;�/�+�\4tv7�W$o�	�V@2�?M��&��̈́T$v�&�ʍ&�;{F!���>V�!���=A�"`�                                                                                                                                                                                                                                                                                                                                                                                                                                             U8�T��J�p :�.�*�]5ew7�S%u���W�A3�G����&!����AU%w'���&Cz�b��#W�d'LZ@���eG�h�L�                                                                                                                                                                                                                                                                                                                                                                                                                                     #8�"��<� L�X�\�+C\��OS�~�!7E�s5Ө�x&�F�!�#S#Q�2?�&cшYn��!��3n��6q��d#˴b�#������                                                                                                                                                                                                                                                                                                                                                                                                                              �8~��n�� �k�e��7VS���~�팁��nމ��&!�F��A�������&�C��bX�#��bC�#��b��f�̆B�;uF!-���@ш��-                                                                                                                                                                                                                                                                                                                                                                                                                       N8�O��Q�k !�5�1�F.�lݖO>n��LZ(�����x&�F�!�N>l#<�2h�&aшcn��L��n��[q��d~#��g�dN#��b^��Ɇ�����                                                                                                                                                                                                                                                                                                                                                                                                                8�	���- g�s�wp�zhs*u�3x(U�
n�X�郛�&C#�>Bx*GzheeJ&H'����
c>�a���8G�hĹ2��1��vƌC�x�~��C�!����0�                                                                                                                                                                                                                                                                                                                                                                                                          �8X��H�8� �M�C�7��h�7pS؈�X����H���#;�&!�`��A�؊��5�&�C��b��#��b�#��bg�@�	�B�;SF!���fш6o�	шGdX#�b�h/���                                                                                                                                                                                                                                                                                                                                                                                                 �8��{�#����t��;��3O��������M`x&�#&��Ɏ���&��;�F!`��>��!���=��!�ێш�d�#�b%�	�b�#J�b�_�r�B+;lF!��;�qш1�H                                                                                                                                                                                                                                                                                                                                                                                           �8��x� ���w��H�70S���������f�c{�&!� ��A����~�&�CǴbL�#��g�n���q��d�'ш�d�#�b �&�<��I�͆B;\F!��(�oш�d8#r�bqH�FI"s`K                                                                                                                                                                                                                                                                                                                                                                                   �8^��N�>� �K�E�1���7vSގ�^����N�J�%=�&!�f��A�ތ��,�&�C��b��#��b��#��b��F�	�B�;UF!>���`ш�o�ш�d^#�bn)���B~;4F!����b��F"a`                                                                                                                                                                                                                                                                                                                                                                           �8���h� ���g�x�7 S���������_�sk�&!�0�iA�����9�&�C״b~�#��b��#��b����B�;F!ʐ�6ш�o�Yшd#L�bf8�ۆB(;bF!��X��Yb�H�SIL�xB�y1�[                                                                                                                                                                                                                                                                                                                                                                     �8x��h�� �m�c�����PO��xն���h��x&�F@!����#��21�&��шMn�����Yn���q�����`шed�#s�b��F�ц�)���Bx;<F!/�H�ш�dX#�b�(�F)�B8�9��d!�	��B����+                                                                                                                                                                                                                                                                                                                                                             #8�"��<� L�X�\�+Cxsu�<S�~�!7E�s2M��&����#S�Q��[&�c;F!���>!�!��=6�!���ш#nЏؑ��d3#�b��#��b\�����B�;�F!ؐ�ш d�!N��B�c��ld�!p���B����o|"8BC"�`�                                                                                                                                                                                                                                                                                                                                                    j8�k��u�O ���b
I6�
xJ=�7�h~�>:����&�2�1(j!H���&(*vE�CKw�}h�C�u�{�C!Z��i�jG�hļ2z��1���1<��vތC�!���ȺG�h�B2�ˌC&!�*�č2�9�C�!�L��I7��Sa���Bf1��                                                                                                                                                                                                                                                                                                                                             l8�m��s�I ���d,O7�SL��1�n�x
�<�����&!����AlN�|�&,CC�be�#n�b��#y�b\��6�Bl;�F!ϐ|��ш�o��шd�#شb����"�B�;�F!P�̄�b��,F�!א�?�b��JF�!���O;UC!J��`b�,sF-"�`�                                                                                                                                                                                                                                                                                                                                    �86Ǉ&�V� �#�-�YΦ��7S���6��āҠ&���MU�&!���Aƶ���^�&�C�b��#��b��#��b��.�\�B�;=F!Ԑ֎ш�o�gш�d6#r�gd#A�b\���Bf�g�!�v��wbF�FG!t�V��Wb��x�����,d�!ʷ�B�ه�n��4�b&e                                                                                                                                                                                                                                                                                                                              �8t��d�� �a�o��䤧7\W�otٶ���d�Y�x&�FL!����#��2��&��ш�n������n���q��d�#l�bB��/�B�;JF!˼B?%F!��t�0ш�dD#�b>T��$�F%!�4��5b{�F!c���b|ڧ#��2���F�!��Ą��b��!v����AF�"�`'                                                                                                                                                                                                                                                                                                                      `8�a���E ��8�hPC�@�=bt�0o���x&�F�!�`B#�2�& Oшn��b���n��uq�#dP#��b�`����Bp;�F!��B?�Fy�B�;�F!?����ш�d�#��bL�F�}�B� ш�d�!3��B�F�rnC�Y��Ud!lцB !�dn���1b��!�A��BPwFQ"�`�                                                                                                                                                                                                                                                                                                               `�    [�[��  @ �}<�t= ���   �vN�G	�tU�G"	�tMjh   �wj ��c  PVW��w�O�ǉ���������_^�$��W�f  Xh @  �wP��g  ��(Nu���v  	��  �N	���   ��W��W  	�u=jh   h   j ��c  �ƍ��  WPV��o  jj Vj ��s  ��~   �d$,�ǋ	�u�N	���   �V�	�u��넩   �t%��  ���PQRPW��[  ZY	�uRnjh   h   j ��c  ��_��  ��t���  ����  UWPV��o  jj Vj ��s  ��   �d$0��������o�����������D$�Pjh   U��_  �@ � �  �`` ��Nah `C É����d$ USVW�Ɖ����1ۤ��m   s�1��d   s1��[   s#�A��O   �s�u?����M   )�u�B   �(���tM���H����,   = }  s
��s��wAA���V��)��^� �u�F��1�A�����������r��_^[]�                                Could not load dynamic link library %s The procedure %s could not be located in the %s The ordinal %u could not be located in the %s             {s Ws             �s os                     �s �s �s �s �s     �s �s     KERNEL32.DLL   LoadLibraryA    GetProcAddress    VirtualProtect    VirtualAlloc    VirtualFree USER32.DLL   wsprintfA   MessageBoxA 