MZ�       ��  �       @                                   �                                                                                                                                                                   PE  L #��G        � 
 j  E     �,      �    @                     �    �i                               �  x                            �  �                                                   �  X                           .text   i      j                    h.rdata  
   �      n              @  �.reloc     �      r              @  @.data   G  �  G  z              @  �                                                                                                                                                                                                                                                                                                                                                                                                        U��j@h   �E�P���I  �X�/��,�@ ]�Wf�=/@ f��d_�u)�j �Vf�5D@ f��$^�uѝP�Uf�-X@ f��r!]�uם� U���0VW�E�    �E�    �E� �EE�E܍M�Q�U�R�EԜW���Ǽj  �_�3��E�P�Uf�-�@ f�ŗp]���   ��E�Pj@�M��Q8R�EP���  �P�Qf��@ f��d"Y��s  �j �M�Qj �UR��  ���2  Rf�@ f��h&Z�u ��UR�Eܜ�E������Uf�-2@ f��a7]�u��  �Uf�-J@ f��3�]�uC��u�Sf�_@ f��"b[�u��P�Pf�q@ f�0xX��  ��  �Vf�5�@ f��y ^�u���E    �E_^��]�Sf��@ f��BI[��{  ���
  �����Wf�=�@ f��q�_�u���Y  Wf�=�@ f��_���  �������Pf�@ f�7(X�u\��.  �����Pf�@ f�d�X��Z  ��U�Uf�-8@ f��h]���   �R�Qf�P@ f���TY��E�����EP����������   Pf�u@ f�YIX��k�����<  ���ȅɜQf��@ f��X4Y���   ���@ ���Pf��@ f��wX�u���vPf��@ f�$X��������uWf�=�@ f�ǉ#_�u7��M��@ �}�����ʃ��3��}�5�@ �5$�@ �u�uܜ�	������Rf�.@ f��1Z�u��Ý�E    �������u0Vf�5S@ f�� X^��y�����M�Q�Uf�-n@ f��y]�������U���������0���Qf��@ f��fY�����U��h�  �W���ǂG  �_� ��(�@ �Wf�=�@ f��_�u�� �]�Pf��@ f� qX�u�U��} �P��]E  �X� ��t*�h �  �Rf�@ f�6Z�u2�P�Pf�"@ f�WX�u	�]�� �� ��$�@ �Pf�B@ f�c�X�u��j �E�Wf�=Z@ f��CX_�u�U���PVW�E�    �E�H�P��K  �X�  ��E�    �Sf��@ f��Xq[���  ��M�Sf��@ f�Òt[���  ��M����M����   ��EܜUf�-�@ f��d]�u���}����q  ���]�Pf��@ f�esX�um��M  ��j�M�Q�Pf�@ f�X��$  ��  �G  ����UĜQf�C@ f��vhY�u���E�H�M��E�    �Qf�f@ f���SY��B  �Ý��E���Vf�5�@ f���^��"  ��E�P�Pf��@ f� dX��\�����U�Rf��@ f��r9Z�un��U�E�;B(��  ��M  �Sf��@ f��q[�u ����U�Qf��@ f��5EY���  ��UĜ�$�����}��u�3��Sf�!@ f�Åx[���  ��B�E܋M�Q�U��E�H�M�h�@ j�Pf�U@ f��YX��u  ��L0Q�Wf�=q@ f��(�_�uU��E_^�Rf��@ f��DZ��\����������Rf��@ f��5CZ�������U���+���Pf��@ f�i$X��6�����wV  ���Sf��@ f��V�[������������Rf��@ f�Z��$���������Sf�@ f��8[�������MЋP�UԋE�H�M؜Pf�@@ f��0X��]�����U��Rf�Z@ f�XZ�uI���������E��0��MȋP�ŰH�Pf��@ f��0X�u����)���Rf��@ f��IZ������R�Pf��@ f��GX�up��Sf��@ f���[��������U�� �Pf��@ f�X�u �R�E�P�M�Q�Rf�@ f��B�Z��������M؋U�B�Rf�!@ f��bYZ��������Q  ���   �Wf�=E@ f��XY_���������Y�����M�Q�U��E�Vf�5n@ f��c@^��������Q�U��Sf��@ f��Ip[�������R�Wf�=�@ f��p8_������U����E�Q����'  �Y�   ��E�P��  �W�Ý�t���M�y( �Rf��@ f��Z���   ����  Sf�@ f��x#[�u ����  Pf�"@ f�HX���  ����  Rf�>@ f�1Z�u�����   Vf�5W@ f��^��I  ���@  ���Pf�s@ f�QPX�u˝�E��Pf��@ f�(9X�uP���>�����U�z, �Wf�=�@ f��t_�u~�P�Qf��@ f���HY�u���E�Wf�=�@ f�ǐ _���   ��E�    �}� �Vf�5�@ f��p�^����������   ��M�MQ�Qf�@ f��xiY��  ��}� ��ҝ������Uf�-@@ f��P4]��������E�Sf�Z@ f���[�ux�]�Pf�l@ f�5GX��_������<  �E�Pf��@ f�r7X�un��}� �Vf�5�@ f��1^��O������OUf�-�@ f�� ]��b����h�@ h @ �U�R��r����P�M�MQ�U�B(P�M��Qf��@ f���1Y�uE��E����W�����E��0�Wf�=@ f��U_�������������Wf�=8@ f���_���������0Q�Wf�=S@ f��0_�������M�Q(R�Wf�=q@ f�ǒ_�u����������W�\$S��\$S��\$�l$Um<���M�U�Ń��]Q�����H<�XHS�(��[���p��H;H|�HQ�x��H+Hx	$P3��XY+�^`U�X'����� uj�;�� uj�2��@uj�)��`uj � ���uj����uj����uj@�h�   QW��aV��(;��v������   �R�d�0   �@�@��9Xt� ;�t��PYYX���� ����l$��T$��L$�ah �  j �t$��t$�D$������������������U��]����U���0�} �R����  �Z�  ��1  ���Sf��@ f��	[��B  ��U؃��U؋E����E��Sf�@ f��42[���  ��E؜�3  ����Sf�5@ f�ÄS[���  ��EP�Vf�5P@ f��6h^�uY���  �3��Pf�k@ f�PEX��  ����  ��   �Pf��@ f��X�u ���.  Qf��@ f��rY��z  ��V  ���E�M�Q�U�R�Sf��@ f��I�[���   ����  ��M��Q�U�Uf�-�@ f��q	]��p  ��HQ�UR�Wf�=@ f��GQ_��#  ���#  �3��Vf�57@ f��u�^�u ���  Vf�5O@ f���^���  �������@ �E��}� �Uf�-x@ f��G]��������  �Pf��@ f�tX��K  ���@ �E��Qf��@ f��"!Y�u��M؃9 ��m  ��}� ��P������@ �E��Sf��@ f��S$[���  ����   Sf�@ f��G�[��   ��E�P�M�Q�U�R�EP��S  ��   ��U�BhP�MQ��(���������M؋��R�Uf�-V@ f���]��������
  ���E��Sf�x@ f�Ó�[�u ���Sf��@ f��[���  ���*  Sf��@ f��f�[�u"���V���Sf��@ f��t�[�u �3����   ��M�yh ��������B  Uf�-�@ f��)]�u ��   ���  ��U��Pf� @ f�X���  ��E��x �Vf�5/ @ f��Q^�uq��E؜Qf�E @ f���SY�u
��E��M�뮝��\���Vf�5g @ f��!�^��������E��������U���E��}� ��K������3  Sf�� @ f��c)[�u՝��I�����M��QR�EP�Wf�=� @ f��0_����������   Qf�� @ f��5$Y��!�����������3��Uf�-!@ f�Ń@]��������} �Sf�!@ f��%c[��������U�����f��t!��U؋%   ��Vf�5M!@ f��Sd^������������M�Q�Rf�m!@ f��)�Z���������  ���Vf�5�!@ f��&c^�������Ý�U��Uf�-�!@ f��A%]��r���������Pf��!@ f�F)X�u����]��ǝR�Sf��!@ f��i8[����������EܜQf��!@ f��X#Y��X�����E�    �E�P�MQ�Rf� "@ f��Z����������E�Wf�=="@ f��a_�u����  �Pf�S"@ f�7X�uѝ������Q�Pf�m"@ f�&X�u���K���Sf��"@ f��Y&[��������U��Qf��"@ f��TY��&�������Pf��"@ f��GX������U��� j �E�P�M��Q�����P  �Y�Z�  �  ��M��Vf�5�"@ f��E�^���  ��  ���E��Pf�#@ f�#�X�uʝ��  Pf�/#@ f��X��d  �Q�UR�Sf�K#@ f�ÓB[���  ��M�U���U�Uf�-n#@ f��6]���  ����  Vf�5�#@ f��Ep^���  ����    �Sf��#@ f��5 [��;  ��U�f�f%��ȋU�
Q�EP�Qf��#@ f��s�Y��#�������  Qf��#@ f��XFY��/  ���,  �2��Rf�$@ f�bZ��Z����������Sf�1$@ f��sh[��w����  ���9M��Uf�-R$@ f��R�]���   ��M��ɜ�h  ���K  Qf�|$@ f��siY�u���H���Rf��$@ f�rZ�u��Ý�M��������+M�M�Vf�5�$@ f��2^���  ��+U�E���Rf��$@ f��H�Z�������  ���F���Sf� %@ f��Hi[��1  ���K���Pf�%@ f�'6X��������E� �E���Uf�-;%@ f��H]���  ��s���U�f�f��f���ȃ��Uf�-j%@ f��w]��������U�E�B�E�Rf��%@ f��HZ����������   �������Rf��%@ f�eZ��,�����U����   P�MQ���   ��uW��U�: �Uf�-�%@ f��	�]���������Vf�5&@ f��3Q^��  ��,  �����Uf�-"&@ f�ŀ]�������������E��   ��E��H���Rf�R&@ f��7xZ��������]��5�����U��$������m���Uf�-�&@ f��e�]���������Pf��&@ f��PX�uǝ�uÝ��Rf��&@ f��rZ�uԝ�M  ���E��E��Vf�5�&@ f��($^��,�����H�Sf��&@ f�ÅI[��������E��E�    �Rf�'@ f��&Z��������<���Pf�)'@ f�$X��������E��E���U����E�E��S���ÿh  �[�  ����  �3��Pf�p'@ f��0X��  ���  Wf�=�'@ f��f_�u
���]���  �3����  ��:PE  �Rf��'@ f�SZ��q  ��E����E��M����M����   �3��Sf��'@ f��6H[�u��M����MZ  ���   ���Pf�(@ f�qiX�uڝ�MH<�M��U�Uf�-0(@ f��e�]��l�����   ��M������F���Qf�X(@ f��AY��a�����} �Sf�s(@ f��2[���   ������Vf�5�(@ f��v^��^  ��E���t���� ��} �Uf�-�(@ f��G]���   ��U��=  �Wf�=�(@ f��5%_��y������������E�H<�U�<PE  �Vf�5)@ f��^��i�����} ��<�������Pf�*)@ f�	X��������������3��Rf�K)@ f��(Z���������������E�M���Uf�-r)@ f�ŖF]�������Ý�����Wf�=�)@ f�ǒ_���������o���Sf��)@ f��P�[�u%���������U�E���Pf��)@ f�wX��������M�U���Uf�-�)@ f��U3]�������M����   �M��} ��U����E��R����du  �Z�   ����  Uf�-8*@ f��)]��|  �k�(�Vf�5R*@ f��IG^�u���]��y��U�k�(�E�L�E�L9M�Sf��*@ f��Fq[���  ����Uf�-�*@ f�ł$]���   �P�M�Q�Uf�-�*@ f�ŃR]���   �9E��Rf��*@ f�tZ�u<�Ý�M��Rf��*@ f�7Z��d  ��M�k�(�U��Qf�
+@ f��qxY��R  ����   ��M�k�(�U�E;D�Qf�9+@ f��xY�uK�E�E��E�Uf�-U+@ f��u]���   ��E�    ��>������U�R�EP�Qf��+@ f��19Y�um��rܝ�M��Vf�5�+@ f��I(^���������   Pf��+@ f�X�uV�3�������3��Pf��+@ f��9X���������y���Qf��+@ f��XPY�uН�@��������Sf�,@ f��2[�uʝ�M�����������0���Pf�1,@ f�V`X��/������'���Wf�=N,@ f�Ǒ�_��������U��B��\�����E+D�M�k�(�U�D�Rf��,@ f��FZ��������̐�Q�����   �Y�  ���g  Rf��,@ f�)Z��h  �`P��X��@ ���@ ���  �h �@ �Rf��,@ f��Z���  ����Vf�5-@ f��Aq^���   ���  Uf�-#-@ f��XP]��z�����/������Pf�@-@ f�bPX��@  ��˜Wf�=Y-@ f�Ǔ�_��^  �� �@ ���Wf�=x-@ f��x0_��  ����Vf�5�-@ f��e�^���  �j j j ���  ���@ ���Sf��-@ f�ÐC[��S  ����Pf��-@ f�X��;  �Y���Uf�-�-@ f��P�]��T  ����  Rf�.@ f��ftZ���  �j j hX�@ �Sf�,.@ f��Wc[���  �j j j j ��ԝ�<�@ �Qf�U.@ f���'Y��|  ���  Wf�=q.@ f�ǖ_�� ����a��  ���  Sf��.@ f�Ùg[���  ����  Rf��.@ f��3�Z���  ����  Wf�=�.@ f��&_��V  ����   Qf��.@ f���Y���   ��d����Uf�-/@ f��Ps]�������Ý�����Rf�'/@ f�Z��.�����@�@ j �Uf�-F/@ f��1]���   ��I  ���Pf�b/@ f�X��Q����j hc7��Qf��/@ f��a�Y��  ������j j j j ��0��[TSV��  ��v:Sf��/@ f��Q	[���  �9C��  �j j �Uf�-�/@ f��F�]��  ���@ ��@ ��t  �j j �Sf�	0@ f��A�[���   ��H�@ ���Pf�&0@ f�X"X��p�������  Pf�@0@ f�X��_  ����  Uf�-\0@ f�Ńq]��)����j �Qf�u0@ f��#bY��<  ������Pf��0@ f�AbX��  �� �@ �Pf��0@ f�E�X��������P�@ j j j j �Wf�=�0@ f��_�������j j j j j �Pf��0@ f��X���������z������Uf�-1@ f�ŉs]���   ��[�[�Qf�-1@ f���1Y������U�Wf�=E1@ f�Ǔt_���������l���Vf�5b1@ f�� ^��$  �j������5  ��S S;Pf��1@ f�e1X���������x  Uf�-�1@ f��&T]��������n   �Sf��1@ f��6r[�u\������Z�������Pf��1@ f�96X�������0�@ ���Rf�2@ f��Z��������Y���Pf�2@ f�UX�������'  �������R���Uf�-C2@ f��8]���������&���Pf�^2@ f�1X�u�j j j �������VP�Qf��2@ f��UY��@������   Qf��2@ f�� qY�u��oSf��2@ f��F[���   ��8�@ ����Uf�-�2@ f��Iy]��5����j j j �Uf�-�2@ f��g]��n������@ �Qf�3@ f��XvY�����������������Uf�--3@ f��xU]��_�����;˜Vf�5H3@ f��x0^������Xd�0   �Pf�d3@ f�$X��Y������@ ��@ �Vf�5�3@ f�Ɓ`^��|������Sf��3@ f��4�[���������뇝j ��?������U���@�E�HS3�C����H�U�����]  �]�  ����  ��u�:������Sf�4@ f��![��  ��M��i  ����  Wf�=/4@ f�� _�uݝ��  Pf�F4@ f�9eX���  ��L		�M��M�Rf�g4@ f�BZ��  �f�
�M��U䍔J�  �Sf��4@ f��%[���  ��L9�Vf�5�4@ f���^���  �B�Sf��4@ f�� [���  ���}  Pf��4@ f�StX��`  ��F�U�u��Pf��4@ f�IBX���  �)u+�3�f����  ��M̜Wf�=$5@ f��Hw_���	  ���9  �E�   �Sf�I5@ f��$[��$  �f���Wf�=d5@ f�Ǉ_��  ��e؋M؋U��   �M��=   ��J   �Pf��5@ f�e)X��}  ��M؋U�Pf��5@ f�H X���  �)u��Z  ��M��D  ���$  ��E��}��Qf��5@ f���dY��  ��M�Qf�	6@ f��)"Y���  �I���  ��s���ƜWf�=.6@ f��vw_��`  �f������  ����  Wf�=Y6@ f��c_��[��������+ΜUf�-w6@ f�Ŗ8]��E  ���9U�Vf�5�6@ f��ir^���  ���/
  ��U�1�����A�Rf��6@ f�Z��p  ���
  ��u�������Uf�-�6@ f��6�]���  �f�1�Vf�5	7@ f�Ɨ^�����������E��]�Pf�)7@ f�EX��D  ��E����u�Uf�-I7@ f��5P]���  ��s��U�;U��Uf�-j7@ f��`r]��A  ��  ���6  ��ƾ   +����Vf�5�7@ f���^���  ����Rf��7@ f�SZ��d  ���6  Pf��7@ f�u�X��l�������  ��M���3��Qf��7@ f��EY��R  ��}� f�1�Uf�-8@ f��	Q]��F  ����  ��u�:�����B�u�U��Sf�J8@ f��"�[��  �j��q  �;U��Pf�k8@ f�7X��p����3ۜUf�-�8@ f��4]��$  ��M��Rf��8@ f��wgZ���  ����
  Pf��8@ f�'XX��  ���3  Qf��8@ f���Y��f  ��}�
���  ��M�;M��Vf�5�8@ f��3^���  ��e� �Wf�=9@ f��i_���  ���#�I�����Sf�;9@ f��`e[�����������9u�Qf�[9@ f��I�Y��\  ��   �Qf�w9@ f��'Y��w  ��M��Uf�-�9@ f��1w]��u  ��=   �Rf��9@ f��Z��N  ��U��M�E��}��Sf��9@ f��r�[���  �ќPf��9@ f�F9X��4  ���U  Uf�-:@ f��5 ]��p  ��}�;}��Uf�-#:@ f��`�]��l  ���w	  ��ǜSf�D:@ f��qE[��H  ����  �9u�Wf�=f:@ f�Ǉq_��|  ����Uf�-�:@ f��X�]��  �A�u�Wf�=�:@ f��_��   ��]��  ��  ���|  ��M�;M��Pf��:@ f�2X���  ���Q�  �Uf�-�:@ f��27]��^  ��ڜPf�;@ f��!X��  �3ҜPf�;@ f�%UX���  ��M�f�2�Wf�=7;@ f��V_���  �+�M�}��Wf�=W;@ f��V _��q�����U�Uܜ������U܉U���靜�  Qf��;@ f�� qY���  ����  ��M�;M��Wf�=�;@ f�ǇP_��$  ��M�>GA�}� �U�}�Vf�5�;@ f��Aq^��  ���5  ��M3�C����M؜Wf�=<@ f��	_��3�����}� f�
�Pf� <@ f�r$X������������B�u�U��Sf�F<@ f�Æ	[���  ��M��U䍴J�  �u�Rf�m<@ f�EZ��  ���1���Wf�=�<@ f�Ǆ0_��$  �c  ��e��M̜��  ��M��Uf�-�<@ f��H�]���  ���  ��u�Sf��<@ f��X�[���  �+U��E�Uf�-�<@ f��@]��R�����}��E�9}�볝���  Wf�==@ f��_��������M̜�u����  �f��������9U��T  ��M��  ������Uf�-m=@ f��P5]��A  �����9E��  ���S�����e� �Pf��=@ f��fX���  �=   ��?  ���M���C֜Pf��=@ f�"�X��P  ���&  Pf��=@ f��FX���  ��ƜUf�-�=@ f��Cd]���  ���H�����M�Uf�->@ f��T]�uA�+�3�f��f���Uf�-:>@ f��fA]��  ��]��=   �Pf�Y>@ f�'�X��  ����  Pf�s>@ f�GSX�������;}�Wf�=�>@ f�ǉ_��������}��M��Qf��>@ f��ugY��z  �)u���  ����  ���M�U�+Ӎ�Q^  �Sf��>@ f��%[���������  ��E�;E��Rf�?@ f��IYZ���  �;M���?  ���/  ��   +����Mf�1�M��u����ϜUf�-U?@ f��b�]��!  ��m��Pf�n?@ f�b�X���  ����  ��M��Pf��?@ f�f9X��Q  �)u���  ��u��E 6  �Pf��?@ f�E�X��\  �+�f�Q��  �Uf�-�?@ f���]��i  ������Wf�=�?@ f��fx_����������	  Qf�@@ f���8Y���  ��]�ۜ�����������9u�Rf�C@@ f�� �Z�u���U�����
`  �M�E�   ���  ��tjUf�-v@@ f��W]��q  ���   �N�Pf��@@ f�3iX��  �A�U�M��Vf�5�@@ f��^��a  �+ƜPf��@@ f�DIX��P  �3���	  �)U�]̜�
  �f��� �����tܝ�u������A�u�Uf�-A@ f��a]��_�����M�<�}��=   �Wf�=?A@ f��Q_���  ��E�M�E���M��Uf�-dA@ f��pD]���������+M�ΜUf�-�A@ f��F�]��r  �f�
��  ��   +�����e�f�;�Pf��A@ f��(X��n	  ��   +����Qf��A@ f��Y��"����3��Sf��A@ f��eB[��Z  ��1�Hʸ   ���}�Pf�B@ f�YIX�������f��ً�����P�����MԋMܜPf�BB@ f�b&X���  ��\+ΜSf�_B@ f��u[��������M��U����=   �J�Vf�5�B@ f��5 ^��y�������  Qf��B@ f���Y���  �������4  Vf�5�B@ f��Q7^�������u�U��Uf�-�B@ f��g]��I�������}� f�2�Pf�C@ f�sX�������f�
�ٜ��   �f�2�Qf�,C@ f��$Y��  �)u+�3�f��f��+�=   f��Qf�[C@ f��Y���  ��M�<�}��=   ��8�����U�Sf��C@ f��D([��   ��u�Rf��C@ f���Z�u
�)}���  �3ɜRf��C@ f��Z���   ���n  ��ƾ   +�������e� �Qf��C@ f��pY�������������Wf�=D@ f��xB_��  ��R�U���	�}���
l  �M�Uf�-ED@ f��W]���   ��U�U��E�   ���������Rf�sD@ f��fZ��6������K  Qf��D@ f��I2Y���  ����f���Rf��D@ f��40Z�������}����Pf��D@ f�WX������j��@^;ޜSf��D@ f��'R[��  �+�3�f�ќSf�	E@ f�Ñ�[��@������������M�+M�U�
�M؜Uf�-8E@ f��3�]��!������I���Uf�-UE@ f��C$]��G������n�����}�Pf�uE@ f�FX���	  ���������ȜVf�5�E@ f��v$^���  ���
  Vf�5�E@ f�Ƙ�^��������������U�������Qf��E@ f��UY�������;M��Pf��E@ f�8vX�u���������3�G�Wf�=F@ f��_���  ��Uȉu��]�]܉]��]ԜSf�>F@ f��tR[��7������
  Pf�XF@ f�BX��6���������Pf�rF@ f�7X���  ����  Vf�5�F@ f��cy^��>  ���4�����]�?���Rf��F@ f�� YZ��R������]  �����   +��Vf�5�F@ f��^���  ����	  Pf��F@ f�	X�������)u�Uf�-G@ f�ņ�]���  �B�Qf�/G@ f��3WY��������UԜUf�-IG@ f��y7]��������1�����M�;M��Rf�nG@ f�Z��o  ���U�1�Sf��G@ f��U[��p  ����  Sf��G@ f���[��j  ������Wf�=�G@ f��_��  �9}�Qf��G@ f����Y��B�����������M�;M��Uf�-H@ f��R6]����������  ��U�;U��Uf�-+H@ f��E�]��2����f��f���E�   �E   �Uf�-WH@ f��C]��b������&  ��   +�����e؋�f��Wf�=�H@ f��0W_�������f��+�f�C�Pf��H@ f��X��v�������  Uf�-�H@ f��"]��4����3Ƀ}�����w	  �������Vf�5�H@ f�ƒY^������������Sf�I@ f�Ùg[��������ً�����9u�Sf�4I@ f��[�uY�������Pf�JI@ f��X���  ���D  �U�u�G�Pf�lI@ f�4�X��������u�#u�Sf��I@ f�Ò�[��8  �������Pf��I@ f�2X��E  �+�f��Rf��I@ f��W�Z���������m  Sf��I@ f�Èp[��$  �_^[���  �@�Sf��I@ f��Wc[��������}Љ}؜Pf�J@ f�S�X�uI��E�   �Pf�2J@ f�FX��������
  ���������u�9���Sf�_J@ f�È&[��i  �5�������f�q�Pf��J@ f�@X�������3�f��f��+�+�f��U�B�Pf��J@ f�xX��������������u����Pf��J@ f��X���������������u������A�Rf�K@ f��!Z���  ��M�;M��Pf�K@ f�vX��x�����������	  Uf�-=K@ f�ő]��e������  ���f��Uf�-bK@ f��s&]���������Q�  �Pf�~K@ f��`X��c���������Qf��K@ f��cCY��<������e  ��º   +����Sf��K@ f��7[������ɜSf��K@ f��@[��=  ��MW�xJ�U���1�M �Uf�-L@ f�Ŕ]�������f�
�ً��&�����ƾ   +�Qf�5L@ f��FY��e����f��������9U��  �f����������e����AB���}�M��Vf�5�L@ f��Q^����������Vf�5�L@ f��Y�^��G����A�u�M��Uf�-�L@ f��]��������u�M��Rf��L@ f��U�Z��Y������x���Pf��L@ f�I!X���������������
�Sf�M@ f��CQ[�u_���=���Sf�/M@ f��I1[��  ��º   +֜Pf�MM@ f��X��B����)U+�3�f��f��+�=   �U�f��M���������������U��Pf��M@ f�@�X���������1�����U�1�����A�U�M��Pf��M@ f��pX��j����Y�Wf�=�M@ f��uY_��c����������Pf��M@ f�C�X��8����f�Q�ڋ�����9u��_��������U���Uf�-5N@ f��a7]�������)u+�3�f��f��+�=   ������f�
��������9u������=   �Vf�5�N@ f�ƅF^��P����)}3�f��f��+�+�A�M؋M�	M�f���������ˋӜSf��N@ f�×b[��U�����M��M�f�2�MܜSf��N@ f��d#[��D�����E����  ��}�#}�Pf�O@ f�&X��S������d  �Wf�=)O@ f��1(_����������9u�Uf�-IO@ f��3]��E����f��f��+�=   f�
�Wf�=qO@ f��T�_������������Uf�-�O@ f��$U]�������A�u�M��Wf�=�O@ f��Wq_��W����9}�Uf�-�O@ f��XP]�����������Sf��O@ f��aS[�������)u��  �+�Pf�P@ f�9X��  �f���Pf�P@ f�7�X�����������9u�Pf�<P@ f�erX���������   ������������E������=   ���������x���Uf�-�P@ f��]��5  �;U��Rf��P@ f��PZ��{���������E   �Qf��P@ f�� RY�������E�+E�M��E��M �3�������������Qf��P@ f��V�Y��S����V3�J�Uċ���Pf�Q@ f�U6X���������3�����M�;M��Wf�=;Q@ f�ǉ�_������������������Uf�-\Q@ f���]��J������g�����U�Wf�=~Q@ f�ǘ�_������+�f�C�Pf��Q@ f�qcX��[  ���@�����u�;u��Pf��Q@ f�IBX��~  ��������3�f�:�U�*MȜPf��Q@ f�2QX��������ƾ   +�Pf�R@ f�F�X��_����)U�]�+�3�f�ќ�o����3��Pf�2R@ f���X��������U�Sf�LR@ f��r5[��8����I������M��M��h
  �Vf�5vR@ f��X^������������9M�Wf�=�R@ f��b_���������l����)E���Qf��R@ f�� 1Y��O������������m��Sf��R@ f��[��c������������u�Wf�=�R@ f��'_���   �+�3�f��f��+�=   f�
�M�U��Pf�/S@ f�YRX�������f��ڋ�Vf�5NS@ f��7c^��������u�U��Wf�=kS@ f��28_��������]��Rf��S@ f��Z���������i���Rf��S@ f�PZ�������+�3�f��f��+�f�
�U��MԜWf�=�S@ f�ǖw_��]�����������Rf��S@ f��xZ���������   �늝�����Uf�-T@ f��y4]�������� �f���Vf�5:T@ f��t^�������������Vf�5WT@ f��@�^�������������Rf�tT@ f��Q4Z���������Sf��T@ f�Ç[��������   +��Rf��T@ f�Z��������M̜�"�����ƜPf��T@ f�$gX��������U��Vf�5�T@ f�ƙQ^��������u�Sf�U@ f��s$[��s����f�
�ٜWf�=U@ f��6�_�u����M��Pf�7U@ f��X�������������9u�Vf�5YU@ f��VQ^������+ƜVf�5rU@ f��2�^��d����|$�V����l  �^��   ����   ��q�Wf�=�U@ f��iy_���  ����  �2�³-������Pf��U@ f�AX���  ��L$�a ��-SV��ŝ3�@�Qf� V@ f��UY��F  ���ӜPf�V@ f�X���   ����H��f��������Uf�-?V@ f��P�]���   ���  ��q�Uf�-aV@ f��XW]���   �������Vf�5V@ f��x0^�u���|K��D$�Vf�5�V@ f�ƀ�^�u����a ��	�Wf�=�V@ f�ǅ�_�uM�� �^�Uf�-�V@ f��h]�u������3�[�Vf�5�V@ f��5^�u��H�Qf��V@ f���1Y��@�����r4�2�³	�Wf�= W@ f��!G_��A����������Pf�;W@ f�1X�u����u����R������I���Pf�`W@ f�96X��u��������U���3�@�Q�����{  �Y�d  �X�Wf�=�W@ f�ǉ_���  �R�URQP�u�M�E�����Qf��W@ f���5Y��q  ���i  �SV�u�W�}�' ;؜Qf��W@ f��YDY�uk����  �Q�Pf�X@ f�s4X�u��E��o��U�Pf�)X@ f�E�X��p������	  Sf�FX@ f���[�u �j�Sf�[X@ f��A�[��&�������  �j�FP�E�P�Wf�=�X@ f��_�ut��M�ȸ   ���� l  P�Uf�-�X@ f��F�]��S  �P�Sf��X@ f��Wc[�u �������u���Qf��X@ f���8Y�ul�^�Vf�5�X@ f�Ɓ`^��)  ��x������Uf�-Y@ f��YI]�ul�� ��u+����E��Uf�-5Y@ f�Ň�]�������ɜ�ԝ�E��n�3�@��K��U 3�;�Wf�=fY@ f��Y_�u�����   Wf�=~Y@ f�� _�u��������Wf�=�Y@ f�Ǉ_�u����   Sf��Y@ f��X�[��[����P�u�E��u��P�E���PV�E�Wf�=�Y@ f��b_�������3���h��}�Pf��Y@ f�"�X��������U���E��Rf�Z@ f�eZ������[�Sf�5Z@ f��qp[�� �����  �Rf�QZ@ f���Z�u��_������|$�R���=  �Z�W�� ���3  Qf��Z@ f��eTY��  �V�Pf��Z@ f�X���   ��r�_�Vf�5�Z@ f��V`^�u����%�   ����   �3�@�Pf��Z@ f�AX���   �F녝���   Uf�-[@ f��Q�]�u �3��Uf�-[@ f��h]�uΝ�uT�B�Pf�,[@ f�3qX�u�^�Vf�5@[@ f��5^�u���t$3�3�W�Qf�\[@ f���1Y��_�����D$�  ������3�@��C�����|2���8B�� �Wf�=�[@ f�ǅ�_�������|2 ��k��������3������*���Pf��[@ f�$X�u����U��S�����  �[�u  ���w��I��G  ���   Wf�=\@ f�Ǉ_���   �j���  ���  �^�Wf�=1\@ f��C_��  ����Sf�L\@ f��A�[���  ��U�Qf�f\@ f��3WY��[  �3����Pf��\@ f�7X��2  ��\8�Pf��\@ f�X��  ��ɜ���T8��  ��v��Rf��\@ f��!5Z������+2���Qf��\@ f��#bY���  ���Wf�=�\@ f��7_��  ��} ��c  �+�+U���ڜ�H  ���A  Pf�2]@ f��VX�uٝ���  �3ۊ��T8�\8����T8�Rf�d]@ f�aZ���   ����  Sf��]@ f�Éf[��u  ���  Rf��]@ f��heZ���  ��   ��M��������B  Pf��]@ f�AbX��y  ��ҜVf�5�]@ f��Aq^���  ��ك��<���@  �M�Pf�^@ f��X���  ��2�Sf�^@ f��A[��  ���ӜSf�:^@ f��Wc[����������  Pf�T^@ f�"�X��N������)  �G�E�Rf�w^@ f��HZ��
�����E�8���Pf��^@ f�"�X��j  ����  Wf�=�^@ f��b�_��V�������& �Qf��^@ f���1Y��  �3ӜQf��^@ f��UY�������B��MJ�Uf�-_@ f��P�]�u��*����3ҜVf�5 _@ f�Ɓ`^��  ��u����E��M���  ����������Vf�5T_@ f��P�^��K����Q�EW�Uf�-p_@ f��u]��������t�����@ �Pf��_@ f�s4X���   ��E���������шL8�����L8�����L8���������=��������Rf��_@ f��ftZ��(  �Y+�������ҜQf�`@ f���5Y��X  ���������& �Uf�-$`@ f��YI]��������U��o����Y�Sf�F`@ f��qp[���   �j�Pf�]`@ f�E�X�u����G�E�ҜWf�={`@ f�ǅ�_��1�����E�������]��+
�M����g������}�����q��Uf�-�`@ f��%a]��H����� �SV��Uf�-�`@ f��g]�������x����+ȜUf�-�`@ f��!]�u'������B��t�����Sf�a@ f��IY[��7�����E���Pf�8a@ f��eX�������_ɜ�|����;}���������ǜUf�-da@ f��h]�us��> ��������������]�\�Rf��a@ f��Z���������D�������Vf�5�a@ f��g#^��|�����������3��Sf��a@ f��Ct[��g����[�Vf�5�a@ f��5^��M������O���Wf�=b@ f�Ǔ�_�������������Sf�$b@ f���[���������r���Qf�@b@ f���8Y�����������Vf�5Zb@ f��x0^��
���������������Uf�-|b@ f���]�������V�t$Wj_�U����,  �]� ��t$V���Ý�u�_^�Qf��b@ f���Y�u��
  Y��OY�Wf�=�b@ f��yb_�u�U�W�����I  �_�P  ���  �F�Qf�
c@ f���Y�uZ���  �Wf�="c@ f�Ǔt_���  ��V  �E��YY�Uf�-Ec@ f��y]���   �+�j�Qf�`c@ f���1Y���  ��  �F�Uf�-c@ f��Q�]�u��  �W�Wf�=�c@ f��1_�u���K  ��J  �Pf��c@ f�1X���   �Vj�u�Qf��c@ f���5Y��P����Q�Pf��c@ f�E�X�uѝ3F�E��Uf�-d@ f��P�]�u���U�Pf�d@ f��	X��0������^�����uS�E�Wf�=;d@ f��b�_��E������Q�Qf�Ud@ f��a�Y�u���N����3��E��Qf�xd@ f��UY�u;�������_[�Pf��d@ f�AbX��������R  �Uf�-�d@ f��Ps]��5�����6  �N���F���3��E���]�j�Qf��d@ f��8SY��������  �؜Pf�e@ f���X�ur��F^ɜVf�5e@ f��5^��z�����^	  �MYY�Pf�9e@ f�e1X��;�����  �u��Qf�Ze@ f��eTY�������3�W�Wf�=te@ f�Ǔ�_�u��3�Rf��e@ f��Z��
���V�W����_  �_�`��u<Uf�-�e@ f�Ő6]�u��t$V�Vf�5�e@ f��Aq^�u�_^�Pf��e@ f��X�u;�ӝ��   Y��OY�Rf��e@ f��Z�u���t$Wj_�Uf�-f@ f��F�]�uŝÐ�R����n  �Z�e��   �G1�1FYYɜUf�-Of@ f�ŗ$]�u^�3��@�F�E�PV�U��Sf�tf@ f��A[�u;�3щU��P�Uf�-�f@ f��P5]�u��U�����W�Uf�-�f@ f��g]�uǝÝ�E��y�Z�E����n�Pf��f@ f�"�X��X�����V����qp  �^�D��V�Uf�-�f@ f��h]���   �����3ǋ}�����<��Wf�="g@ f�ǅ�_���   �U�Sf�:g@ f��qp[�u ���Uf�-Og@ f��!]�uw�V�u��V�Uf�-kg@ f��P�]�u<��]��������3ǋ}���<�}�3��P��l�^[ɜVf�5�g@ f��5^�uT��e W�E�   �Qf��g@ f��UY�u��QS�Pf��g@ f��eX��r�����u��_��Wf�=�g@ f��iy_�������Ý3��Pf�h@ f�X�u�}�3���M��Vf�5/h@ f��x0^�u��X�E�j?$�����Qf�Oh@ f���1Y������U����P���h  �X�?���3߉]���Qf��h@ f���Y�uQ�V�U��E�ܼ��E���bʜPf��h@ f�H X�uN��SW�z�Vf�5�h@ f��Db^�u��P3ӜPf��h@ f�S�X�u���P��@��E�Pf��h@ f�4�X�uΝÝ�I  1>�Wf�=i@ f��0 _�u �1^YY�Uf�-&i@ f��u]�u �_[ɜPf�:i@ f�7X�u�U��� �ES�]�e �} �SVW�E��P���l  �X�Y���  Uf�-~i@ f��5 ]���  ��u�}�Wf�=�i@ f��V _��\  ��ωE��E��Sf��i@ f��[���   ��#Eg�C����U���ܺ��Qf��i@ f����Y���   ��r�jZ�Qf�j@ f��2!Y�u ��u�������}𫫜�N  ��M�u�������}𫫋�E���  ��U+U���   �3ȉ�Sf�Yj@ f�×b[��`  ����  ��E�ܼ��E���bʜSf��j@ f��t[���   �Ý�CvT2�Pf��j@ f��(X�u.�[ɜVf�5�j@ f�ƒY^�uѝ�C1�1C�E3�9]�E��닝�v��E�y�Z�E���n�Qf��j@ f����Y��:����3ƉE��Pf�k@ f�AX��F  ���v  Sf�-k@ f��H�[��@  ����Pf�Ek@ f�X��������:��3E�Sf�ck@ f��'R[��8�����ʋ����}��U��ȋ���Sf��k@ f��D([��������6����E�E131{;EYY�Pf��k@ f�	VX�ub��E�PR�M�Sf��k@ f��`e[���   ����}��ȃ��r�Pf��k@ f��X��F����3ǉE�Sf�l@ f��y[���   ��������U��Vf�5=l@ f�� �^��x����_�Uf�-Ul@ f�Ŗ8]���   �杋C�Vf�5ql@ f��yc^�u���U�����M�Vf�5�l@ f��t^�������   ��   �Pf��l@ f�RX�u���d���Pf��l@ f���X�u���E�101x��;]YY�Uf�-�l@ f�ŕ ]��z�����E�PS�Wf�=m@ f��uY_�������^�Vf�5m@ f�ƅF^��������Ej+�Y;��E�Qf�?m@ f��� Y��j���U��Q�U�S����r�[��   �[ɜPf�lm@ f�E�X�uq��
�B�Qf��m@ f��a�Y�u՝���<�}�m�j?$�3�+Ƌ��������Wf�=�m@ f��b_���   ��Eh/�E�   W�Vf�5�m@ f��Aq^�u�Ý�����Sf��m@ f��A�[�uC��]������ܝ�u�_^�Uf�-n@ f�Ň�]��L�����
�BSV�Uf�-:n@ f��F�]�u��3��}���Pf�Sn@ f��X��-����3��}���<�}�3�+��M��Sf��n@ f��Wc[�u��U���  �} SVW�R�����c  �Z��  ����@ ���Pf��n@ f���X��y  �P�E�P�Uf�-�n@ f��s]���   �P�E�P�Wf�=�n@ f��W_���   ��������������Vf�5o@ f��$5^�u6�ÝV���   ���3ƉE��������E   �Wf�=Io@ f��_��D  �_�Uf�-ao@ f�Ŕ]�u��j|�Sf�vo@ f�É&[�u���M��U�Sf��o@ f��Ph[���  ������M��U�}��
�Pf��o@ f�#X��(  ��{����Wf�=�o@ f��8I_�u������Uf�-�o@ f��A]��g  ��y  OY��F���Uf�-p@ f�ŕh]��W  ����@    �Qf�/p@ f��	2Y�u ��E��(������Pf�Kp@ f�X���   ���+�3Ã����M�E��Wf�=tp@ f��Bf_�u@��t��3��Rf��p@ f�Z������1F1�M�1V�1N1~h�  ��������(�����uٝ��M�+�3�_^��@ [ɜPf��p@ f�e�X��6�����E���Uf�-�p@ f��A6]�u �+�Qf�q@ f��%PY�������}��
�E��Pf�.q@ f�T&X��������3��Ԁ@ �Uf�-Nq@ f�œ�]���������Pf�eq@ f�9X��������������h�  �������Pf��q@ f�#�X��/����D$�L$�P���s  �X�E�N�Wf�=�q@ f��	I_���   �]���$  ���Sf��q@ f�Ò1[�uᝊ�@FI���   �V�Rf� r@ f��iZ�uo��se�J�ɍD��Vf�5r@ f�ƀ�^�u���
�HJ�Wf�=7r@ f�Ǚr_��l�������   Sf�Tr@ f���[�u���vQf�ir@ f��u�Y�u;��ɜ�̝�t$;ƜPf��r@ f�5X�uΝ��1����^�Sf��r@ f��Y[�u �Ý�1;Pf��r@ f�u7X��B����Ý�����Uf�-�r@ f��P"]�u�^�Rf��r@ f��wQZ�u��ꐜS�����N  �[� �U�Sf�s@ f��We[���  ��E�P�Uf�-.s@ f�ŐX]�u�+��3ΜQf�Hs@ f��eyY���   �������Qf�ds@ f��WY���   ����M��Pf�s@ f� VX�uF�V�Rf��s@ f��ESZ���   �jd�E��Vf�5�s@ f��v�^��  �1F��E�1F1���   ��M��Rf��s@ f��E�Z��  ��U����U�Vf�5�s@ f��^�u)��U�E�}��M��ߜRf�t@ f��Z��)  ��E�}��M����Rf�Et@ f�(Z��������M��u��E�   �Uf�-it@ f��P]��F������   OY��F���Sf��t@ f��C[���   �Ý1~1Njd�E�P�Qf��t@ f��p�Y��^����P�E�P�Uf�-�t@ f�ń ]��
�������|��@ SVWj�E��u�_�Qf��t@ f��TUY�uI��������+��E��3�_^��@ [ɜVf�5,u@ f��8U^��d�����uPf�Cu@ f�7tX��P����3����+�3˃��Rf�fu@ f��Z��������Q����3O  �Y�  ��=ڀ@ �Rf��u@ f��FpZ���   ���iҷx  �����  �Sf��u@ f��e[�uM����@ �Rf��u@ f��dZ�uZ��uQ��%��@ �%Հ@ �%��@  �Pf�v@ f�ptX���   �1  �f�AAf��	�МVf�5-v@ f��GX^��u  �e��������؀@ �Wf�=Uv@ f��V_��  �f�ր@ �Vf�5sv@ f��)x^���  �����@ ���@ �J�ހ@ �W�I�Q��@ k�ʜVf�5�v@ f�Ɓd^�������t)��f�j%������@ _�Qf��v@ f���Y��E����jh@ hĀ@ ���   �f�Ԁ@ _�^�Uf�-w@ f��]��}  ��=��@  V�t$W�Qf�Aw@ f���TY��z������f�@ f���@ ���ќQf�mw@ f��Y����������@ i�W  i�8$  ��Ԁ@ ʋМVf�5�w@ f��06^�u����\�����Ԁ@ �Qf��w@ f��4vY��@����������Vf�5�w@ f��@p^���   ���ʀ@ i��  ��̀@ i��  ��΀@ iɿ  ��Ѐ@ �܀@ i�*  �Sf�<x@ f��s�[��=����f���Vf�5Vx@ f��`^��������Ƀ�������Uf�-{x@ f��r]�������jhր@ h؀@ �Vf�5�x@ f��Yv^�u�Ý������Ҁ@ �Ā@ i��.  �Rf��x@ f��SdZ�u �iɕ  ��ƀ@ i�D  ��Ȁ@ i�  �Qf�y@ f��g3Y��������%�@                                                                                                                                                                                                                                             ւ  �  Ƃ      �  �  �  �  2�  ԁ  ��  ā  $�      \�  L�  l�      ��      ��      cefghbhaifahfiejjefafehecchifbfaedhcfbadbggfjhb                                                                                         t�          >�  �  ��          |�  8�  ��          ��  H�  ��          ��  P�  d�          ��   �                      ւ  �  Ƃ      �  �  �  �  2�  ԁ  ��  ā  $�      \�  L�  l�      ��      ��      �Sleep �VirtualAlloc  �VirtualFree �VirtualProtect  �LoadLibraryA  VGetProcAddress  �Heap32First 8 CreateFileA WriteFile KERNEL32.dll  /GetMessagePos SendMessageA  GetInputState USER32.dll  i InternetCloseHandle WININET.dll [ CoUninitialize  ole32.dll �RegEnumValueA �RegQueryValueA  �RegQueryValueExA  ADVAPI32.dll                                                                                                                                                                                                                                                             0(0=0Q0�0�01+1C1X1k1�1�1�1�1�1212I2o2�2�2�2�2�2�2	33'3L3g3�3�3�3�3	4444<4S4�4�4�4�45<5_5}5�5�5�5�56E6O6j6�6�6�6�6�67:7S7�7�7�7�7�7�78>8g8�8�8�89979P9m9�9�9�9�9�9:9:S:f:�:�:�:�:�:�:;1;L;j;�<=.=I=e=�=�=�=�=>0>H>a>q>�>�>�>�>�>�>O?q?�?�?�?�?      0(0>0`0�0�0�0�01F1f1�1�1�1�1�1262M2g2~2�2�2�23)3D3g3�3�3�3�34*4K4u4�4�4�4�4545c5�5�5�5�56K6{6�6�6�6�67#7j7�7�7�78)8Q8l8�8�8�8 9$9D9k9�9�9�9�91:K:|:�:�:�:�:;2;N;};�;�;�;�;<+<G<�<�<�<�<�<�<�<=:=R=f=q=�=�=�=�=�=>>%>E>N>j>�>�>�>�>? ?4???\?y?�?�?�?�? 0    00 0:0U0n0�0�0�0�0�0�0	1&1>1[1�1�1�1�1�1�12<2X2y2�2�2�2�2�2�23&3A3^3p3v33�34(4@4`4�4�4�4�4�45B5]5�5�5�56'6R6p6�6�6�67#7B7c7�7�7�7�78C8e8}8�8�8�8�8949T9p9�9�9�9�9�9:=:_:y:�:�:�:�:;0;P;�;�;�;�;<?<f<�<�<�<�<=f=�=�=�=�=>3>S>m>�>�>�>?N?h?�?�?�?�?   @  �   0<0o0�0�0�0181]1{1�1�1�12<2X2�2�2�2�2�2%3T3�3�3�3�34>4l4�4�4�4�4515N5o5�5�5�5�5676R6l6�6�6�6�67(7B7g7�7�7�7�7�7$8P8�8�8�8�89-9D9f9�9�9�9�9�9:,:X:|:�:�:�:;6;[;x;�;�;�;�;.<}<�<�<�<�<=(=G=�=�=�=�=.>~>�>�>?"?B?j?�?�?�?�?�?   P     060z0�0�0�0141U1w1�1�1�12,2E2o2�2�2�2�2)3G3d3�3�3�3�3434P4m4�4�4�4�4�4515R5k5�5�5�5686Z6x6�6�6�6�6�6757Z7�7�7�78#8?8T8}8�8�8�8�89.9_9w9�9�9�9�9:.:J:�:�:�:�:�:;&;9;U;�;�;<*<E<_<z<�<�<�<�<,=]=z=�=�=�=�=�=>3>N>p>�>�>�>�>�>?M?i?�?�?�?�?   `     0?0W0t0�0�0�0121]1�1�1�1�1 2292S2u2�2�233>3Y3x3�3�3�3�3�3444N4q4�4�4�4�4535S5m5�5�5�5�5�56H6m6�6�6�6�6737H7d7�7�7�7�7
8(8H8|8�8�8�8�89949w9�9�9�9�9R::�:�:�:;&;?;\;�;�;�;�;<6<N<j<�<�<�<�<�<=8=f=}=�=�=�=>3>M>z>�>�>�>�>?B?Z?o?�?�?�?�? p  �   00(0E0m0�0�0�0�01(1>1G1_1�1�1�1�1202M2b2�2�2�2�2�23'3A3]3y3�3�3�3�34>4b4�4�4�4�4�45%5=5_5�5�5�5�5�5�5�5�5 6&6E6N6c6l6�6�6�6�6�6�6�6�6�6	77*7:7Q7X7f7}7�7�7�7�7�7�7888&858O8t8�8�8�8�8�8�8�8�8�89                                                                                                                                                                                                                                                                                                   (�@  ����@ t8Hէa-�6ٲtZ�T�����8�F  | �t���Y�2"���MU���QK�k��z���+�ޑèmA�-�S/r< ��BK��Bn��v�n!#���zlT/B,���|�j�3E��qo�]�����(#�j7{f��0~#u�ᳫ�q�����O�l��Q���3�iʷ6xI9�л_gyNe�H<�@?���a^��l�Ȑ���Ѝ����]8��~�$ǷM��"	��!�!>�������3Yfcp�~>�F�؅��R�&8C�=�����[���l,�U�T�<}0ۻ��n��E����il�z��P"\��ʻ�Pq��#w�W]˲�u�ԯ�'
*�����͝�>GU.�[Ȏ���o�I�÷����D�<�	�X(���ڄO����͎��ab�����UZ�_e����yc,��L]������x�1)�h����hIUݰf8�4>Q|�N=9�c(_��7���iӉ���U%xjI�2���7��f@c�b��wyY�X^�}�M�%;�w#R���Yf��@�|��4��߰)�g˜� ��W�
�>���X`h�?�pN���#U�O��ܕ��$�^P���L����7��S����f�f�j���_g���#������uV��C?o��z`XU�<�h+Ioz%w���덀���Dٍ'�f<�t�����M]H`�[�шs\*e���g����:��O�>��^|FBD�6JAl�J�-�᎔��f�*S���l����-{T{u���zl�.������H����D.gx������i��
��5�ߔ��&��r���9��Uq�3mG�7�̢��awv�בn����A	\뮙�D�� ���3X�X-?F1�3�?mI�I���#���o�6��J��  FP���Ee�M�������R:�MV������Y5w)�⃔W�p	�^�����b���E�W��`n��6�Â	�v׹�|& `Z}�kg1Sa^���g�8!�_�hYIZ���r��aW�NK�ޥ����h�2�e&��^����yX=	�߽�NL��)�ʵ�!�I�m�}��H��@�փ9������#�`d
���,�������y��};?��m\ ���e��A��]�K��Y; �JISf������E�`�o�6 R������C���19���?HCemo�6հ�6�����(���a�&?�-�.�A�g�U6o����(>
��H����yCD��aaOk�$h���ޣ@�m���e`0SJ��3V���������� 0G9�*��7��/`;o�,��ԑ�l<��+�u3����p�4%ٓ�r�p.�b1˼��8�lR�C���*nm������7��S�����o!� ��{ �wbo�_���^����N_aQ9��wWfo�u؆��}��<kN��c �C����Ź[xk�Fײ���L<�����%\0*=;�=�-�kK�"�l�ħ�Aؽfyejz�>-7��Z$`>�V�D���OXqM�1����qWOV,%X���P|G�˺G&$&�W'�y0�+/[�A|E�`�L��ʅev��\q���1T�d�&,3vw�LyT�IL9�x�V�9HUR]��4��ErtZ=�3Ap���S .YQ�k��D���_:/y�^�A��Izѣ/]	�L���������~�[���WO�]x���&����4ݏ��O�-�\"����I�(D���x�wC���.DBH�$HF��)�mhXݽC�C�0�8�2b׼�����њ��'�2�n��z�'�A��9K�n/��Lߏm�Fӈ�CxQ�=�B����Y1�R^���'�$}߾�X{z�Jf��,�2�ز������.�P����m����7�|��'�Y�i^O�g�!`��No�O���I*��M5����a@h_��,�9���D��K��y�A.��D#(Zv�,�޽ip��m��p��n�p07J%�UӔ����������,Pͥ�jS%%����q S%)a��H
*�^j�l#��]
�����"��J�9��oD�����H>l��'�X2�T�؇�Xa�C"� ��NGj$��|��K����[���D	�m��o�(Bӓ�A���]�P�,��P���ȼ����$���V�SǺj�C� ��n��<JQP&���Ɯ��7sR�Ի�b�2�΍p�@���>�Bv��*�ń� N��=����R��dmE����<ߵ�''�-����́��'1�M��m0$"�T?Ƈ�g{��j-n�;��>~V�e"����k�m]�:p�l�q���긤��r~"�nf�S�6r�h��u�&��`�[��#�hR�	�4���ٮ�������zT&�`��ەN�v%�}�}Nd)32$<C$���xW[�Ͷ��Z�K޴Ӫ����QoF���vq�ST��-Wь:�䡫Kg���ƅ�1JMa����#�_�#2
��^4����������B�Y��w���ΤY������r�8@p,g�L��0R�� ���hkmf��i���7�l2#�YXپ��y[_p��Q΃��|�(�X�gA��,�v� }{d�΍�!��I1//䰊LX����Y !����(K�?S1��5����dkЁ�9.�nb���Rt{µY�Ņ������'�3����F/|a�l�nv`�s�(�ǒ}d9��T�X,V��:�"��*�[i��⒍t^J7�N&Bu������q��䯾�%I̒���>��.�n�B��[�����@�Q�D]I^ߘ�M�ú��V��5"v�>�3̖A�HIld��5E��m�B��~	�٢p!(T<��H]�6X��zI�[V�_{���٩Iͷ~h�	�eI��L\�t6�骅fq}F|j���Dt�5���a�𩎌܀���"��v���f��(�!�،1�����d�uԃM9����R�Ź�α	�|��,-P )����e��!�QA�zx@��'��E�Z�4�x/S��W:W=���Y'��2N����>�.m�kH	�+����3SE�(��\l�����X�vT7ϗ�b���˘�H(�-}q�>˽���ey]%q%�Q��i��Q�;���5�|�Zz8m=s����ۙh<:���?I��6*�j����oi���_�Ymqkw LnU�~IE�oY,���:�롉[j*W6rL��hT'Ʋ����{��zz�-�w=tX�3�n�0[3��$��$=�pŲ^���3�s���][�K#�o;��Mp7	l�r	ZR�?N�ںv�)�}�����˝�_@JGs�-џ%����;H�P�ڼ���_�t]�C��Yf�*���0�v�؉b�ɀU�b���O���y/+�G0�̹�ͩ�U�5�w���G��@4��6>)�H�K+�Fۊ�m(�C�5��	o��N�@_P�g��K��_E����`iD���h�'Ny!�K�G��A �l�Qm� |�ozB��$�<��kֆ�I�qB@Y��r�ʹ؆��iϤp\���}��3��,����R�R)���FR@0����m�jE����6�p�e����z�7I�+l:f�0��l�a�
QE)��%yD��F �mT�ˊ�dJ~uK��yv���wY[�Q�C��+�햟�/�l���ʩ���!��)�^+n\q?�����%Q]Pk��:�)���W�Z�]T�J���WA6���L��P�#����杞C��:9lW/7V���w�7��� q�2�e��z�X:�s�7S�:��:� Q.�!n�~&0Q&}��.�}���!cE��#D�Ŭ�4~z�N�mV2#��������jB"El�]�Y������j��12+A�|��x��Z�T:E,`��k}�>n������1��U�?�
-co'T=��f���(o���1�,Z4	`����H�W[kv����O:��)�Ko?s�P�}�7�F�<�ajƊݡ"�УF	9�2%�}|�P��|
���벐Ivl������x$��;:�T2�k�"�]�#`��ڈ�!��j��x�
D�b�ϔ4<L(/x�RѠ�ڲ�B�;�(�N����_khhn����xp�Cì㭊�\ � ,��%~L����D����%��[�&g�Bɷ���I�^��I5&�Pn����.q�����o���`�I��g���M�k���|�ё���$;T�e�uĊ-F�Lڪx�v��T%X�S���Ch4��b��!H�^(J�������i�Y6er����n4i���i������q�\�w��[�n�嬟�v�Y�x���xo�W�31yPMƃx�!_���q�25F��醪�	sk�z.������b����ǜe��};��nT���c�R�[6�Ptwm����Y�jP�*Kb�E'qjR������Vb�6%�&�J`t���C���R�w�D9�+����FhW"mП�84�:���
LE�˜.`�̈�L�f��7�~�W�r!���h�t�8G��<����K�i�$�l�	�(Pui���$�+p#i�DWo�͹���ֻY��c�!{�'��h0��J��F�G1Y�Q<�l���Z"���(_�k_4�=����ܙ�|�"uy���{x����,�}��E�`�z�%r�
��18�8Hm7�ld�K�R	N�+sa� ��~�	(3�ER�������m�1	|yY��xz6��It�����$?yf����!�|e��Q3�|����2�[ݒ�&���. ��R�#O�v�.�ɛ�� @t�O8i��>�]l��8���V��
�]X���� 0�[�z��̊�u�i�J�g��V�� :��W���qMG?�KK��kc��Ʋ������^�&"=ױ^�W�z�8�a�g���@��,��;�]�f��� 0_J��mJ��ß�� ��zX���d�v��F^�G}���7��}���ѴG خ1�^��g�ތ�w
�������>�[
~=*p{��;� �.	4�B�L��a������3���Ҡ���2�K�7Y��y�T��8?{�8c�0��Q�hKHq�A)��QaK2�t�mmnׅmj(]ۿ(r�T����U/��p}˳P�4i�͈>4Z��� wޱ�^1���z�w�l妶볁���Ut?�L$�&�����1����Y8K@�\.��͕m�<�@��೪漯x�l:�yS
�n�z�l���_�@�(",�X���acю�#�`a|�7�e�`�G��=�̘]�S���V�� 6��xM�zHF�S�=��ڟX��Vں�Zf��Π]�T��I��R)F���*8�S.
��M�@�?/4V��-^��<������4��m	H�ǂ�Y�G�ͧG����Ů�9_4r+e��w�` ���|w���()��J��b���T><���O�);6�F�����r�t�V�߭z.h�љ��ZZ'�Sv�!{s
. �Bc��5X����:}9�q��ӷ��m�VHs���u=��o�0�3��z��]��T�{��yU����5��5=��.�5�?R���)t��7Ft2�﯀,t������.��CF"�~�˼� ��10�v�ͅ�B�˓VʌvX6	�`}��޻��lc�z�i���Tn;�z�Z*)��N�D�n��.X���>�6��k@��]�{`��0RA��9f��M�V��ږ~�S.1 ��6��e����P�!�gf�\6T{�v��Mn6
�x
Éyv����U�xv�j�i&
��a�.'^�#&�������d���Tc��%;f{�]�P��ظ��Ղ�<T ����fir#?Y!��il������o�4��+�����)C$%E�Xs�2�����vs�� [q�9����x���E������_���U�Fp��)� MUi03�E�"�<�����q���=aڎ��bP�#��|��K%� {�<B;��~.���Zn�q�'Y9�v��r߀�E��:�~B�����%lj���6�ъ�w�)ۙp�Q@m����{]�ujB�74j���O%&(,�e�1��ÓH5��
��\1H���7����A�!������T6�m���p�fl�d(��i��W��@K��t���B�A�hyG4���D�v�{�bJP�E���z=f�Bꦐf�,}��Wiw�:'����>�k�#��Z�u���G�ˎWD�},�v����y$��x��Z~:��S�]S�^���]��
�N�Eû�"g�d�2����j�N�GW�{;W���W����UT�TL75�$����g��F��[�b;�=f�x�7�^�(�٤鼭6�Q⧸i�����o���u���U7^9�&��+���N���쀚�D�hw֗P�������ѓ�X��;����t��/��S(��?1c�U|�*w]�]���u�����i�_��	a�W�rc���g������⬾|�� �>�ܪV���L�x�h�������4H�h�n3Q��.���;�N��l?��w)~!%3�b���>��:�'+Uu�zo�9��3�c��=�ӂ[����~<a��H��V5%r��AE��':pL�}k,A���{����.��-����v�����C��2���]GXer�V��C��M�`�z�)X`�L ���L8���U�Z�ۏa<H>'��t���P��l�CmUm5��� E�b�鐢($�!��C�8-��-�,>����X�P�mH�,׏�iP(�/L�� Q5^<���P[�,t���5���ܖ3�0�\�M��y��O����RM�5t��l�kġ`����g6򞦃���>]I�H���\E�&�8(���fj��tΦ�
����ЕnH�;��?޵G����� Yݏ��ݒȹ�2k�j���f���@ ��J�[�+���RZ�%�U��4�st�o<6�\quK &�mߒ��s��.�m�DqO�*�b�5��~C�U� ��0>����0�3�o¶,n��j�V�W4HP4��I��Z��dL�6Q���;���?�l/�X��:�>aL�|�$�%+5��H��`���ß�� �>��f�R��n�]����(֌�t��vh��o�݈�T�1Ğ�S����H�y�o��	��{�Y�$���Ә��8�k�l�|�cӹM;�
cH'#y\��X�)Qu�D��� �U��2~��5D�� �f?
(�Kg�gb=\�;��Wy�-�����y�J���L��r��ջl�O9@��A�p��`f�ф7У�GZ�C=�aODlU�I����!X�5,2<�0n>m�φ�J��S��5s��`�P��o^�$ �B�*=�I��Bfz�N�`5�6��]�1t���c��?i2o�|��و�dq2��AsM.l��9�m���01`���M�E}��(����Y('�z����ʵd��|L�Ό��]w$��h��G�I��|��&�����fJ�U8�Ç(����~3	:9@a-�35+$��Ix:�2p�/�b�R�6�"j��J#^���L�Ul�co�ݬ��K)K���C�BtS����!A�3¹n����G��Sփ�\0��������ڗ/�}~��G�.o�)IJ|F�/u��Z*���C��y:h{¿�C}-���c֓�EöZ�JH�sf(�U!��U`�W��O�&�T�gDֲ�����:p�W!�s�5�nPbP&g5�n�`1���'��-wPH�0M��5I$y�(��~�B_�����	^����Q6�nTXķ4_ҝ|`(���*l�z�G@��+�EJ�uh;�!�,ufdʂ�<4�bO< �~��>�[Vo���M�"�+#��	�6�嶮��ᐫ���!>���͑�+��i�:-���x��o�۔���^��g��$�@�1x�e��ɝ��c%���5�[�>�v}L2*��~�a�Ժ�� ��c����K�o��h���J�|N��}E���o���=�(���6@��m5���Fbٗ �/�۝�Uw�g��[��4�g�	5�����놂k�k%��t(߿+�P���`xm���z��[�:J���X?���8�,ש�eB�J;�r��}\�E������Wh�E. =8���lzf�h�.�\u��jK�o�&�s�1��z�������b�=DC#��F�("ۮy��^Y/��:GM��60��AM��m�BlȨ2�	+��3��9�8w%��*ݜQ�l��a^>T�:lO��#4Re[����u������b�wg����a=s�7�y��Na`2��L��H(��A�Y�UcI�Ƹ�#��kic%YN�!��A�/.;��T��G&�ATL܀>]�}�'"����x���(�)S��vR�_�^����)�{��C�#Aj�r8�[�Ҵ�Q�@M'�����6c�� L�yM��fu�����Y.�V�y�δ����VRg&tD�ҏ�5�� �p�98�����*ڬ�U_T1��..�`;a0ř����zaZn�D�� &w��{��k����|�]%�B.9W���@B�^7�q����)j��;
-d�VQ22�5�o�x�ܪ�Vn��3�H���x�ĄG�6q��E�5	!@�"���HVSB���(;�ռ\q�|�)����Vwkh9�8�;�g�:�`� (��"�]˶�}�u=C%�u���~�fV�`P+B�T��¦"��1��1�[�6�j�d�ۚ�$D�ɩW*G��Hf[,�Idg����6�#/���Tu���薥��P�+R�^��^��j���c��g�A��l�
=�5�޶�3��N��͢�!%b�wyU]�m@�i%:z��=��Y��jS
 w��_'_�gdݏ��
�lwK2G�@�*��}���t��ǲ�I/�v��v� ��l�&��屶+���̤�H1��n'A�T}O��^iܾ���f��<5�ז#�$38�oF�  ��sS��5�!La� �o���G96DE��2�]n�M��O���NvJsW<���` �U7��b�pzB�E���2lA����d6��E���lݻ����U�1�&#u�mV�Y����7�26i+*�B�����+)'�+ W=AvX�S3��dw��Z����C�d6C��T&��Ge�9���A5�i��A]��_���>��ӄ�ð����c��L�[hH���5xQ<��`~_�O7�}[)ܒ��5d��y5�%"y���_#��Z	�h+�?2�!	�&�8!�"��G��L�.,���o���S��X��)�0)>����	�ަ襚j
�7��B��b_TS�Q�T��(i��꘮���\`(rz�	O��дx���"�Tk�\�Mba�o_�wt�;��p���
��x%����d�;dC� {�e��h��-U��0
�v�2�QU����$M�2t�pp��uKSvT��S�I�ws�ϛ���nd���u�E��S�������cB����ђ���a����dWX�MQUW8mV����@��I��B/Z��	�f+}cEEZ"ЫMkڽ�:
2�����Mf쉅D����t��֎�Ι^�<���m/����G��R�P��?�&�TPۈ}JݭԺ���7?�@�O��Gx*�Xu�;1��@t<X���l�לUaUK�v����'�k��.A���κ��-�� LzX���i����9zϛu�i
�'	(LR~�=М Sdq�%�������~�1��֕�>r���Ks��	SU8�޾�9�u�F�"@xf�f{"r���[4Hb�n���]ơ��z�]�����W��3�_�5@�k��H�
f�����45��p��<�<�	&��9�y�����c�@�q����>����*yO�I���{-Q�$�������ɴw-rV�5[�);���k�;5�����N��,pxWV�Y��"��5G��#��]g� �z��Jlc�I�۬_L���^D��"t�Z8�\P���=fp��A��>p�2�ί*u>�ԟ@֍Q��=ϡ�8��@N�y�oA�hu���f���8�n��a�l���q 3Y�@[k�a�X��_�,�9z�*> ��E��hH����w|��Z;�"@k�6��vt!�s1�M���<C��ټ���|Q�Bq��R�Bq&�RT�Zt���N3Z?��^Y�{=_�+�;3u���#n�jJ����"�'��"�,,@�/cэA�!u$˼�\�ce�t��ߓ0)�fX4K����K�(��qC�s�I×��V��&�	�W�d�9d0��:d�e�����²��4��y;*d���~��`}����Xd��*KwP��
�!�i��>!c����׋�
�P=g^�>�I�	b��h���Ţ��-ո@6��hxR�/iϫ�'�M�ۋ`�r�����
�����:_�֓} ��6*n�.�:L�d�͖�h����)~��e�;&�IR�ҧ��;ƾ#��~M�9bo����ۗ��>�N������O\I����j@�)�� wX��px���4n�6���<Tk�}���V/,o� *���5���7��>���)��<�3P�Y��6<F1"� ��פ��^�E���mG+�)ʈh$h]$k���(Ӯ2��8Aۨ�pb�r��E��9�q�YR�~�mmu�]x������8�L��5��- �����:+}ǍDEH��D���?K^��wb ��1:�*��of����	n`�@�Se�����98�/����D�d�n*f�6�Om|����_߹5Zڅ����0Js��O,��$m�DJ�wٽ�L�\��ÈC���ioh�<��,������m�~����mp!���i���?L�΅��+sY�d�󽶜xx�X��>&tP,�>�fP$�rÚ�0�"qxS�m������KF��@�B��P�Ӈ�)t,�p.�ރ��/2[tJ��jޒbb��@�Ȧ�����L�;w�s�;yF�%�?<�q����:z|�pe�����M�Aw%(}��.����P2�	Nr�q#;�p�u�
���&�MV���S8i�������X�묾���$�M%�2*�^���'GRU��Q���0�D���k����x)?W"�{h�xRN�|ۍ��/j�����>����=|Ak�[Դߵڳ-���𻽂G&A�}���r�k��j���R�O�A."�����u��.&����&����)N��dH�[�w�kZ���7�AڿY7�.��ByeڊWG�5NIr���8��Z_P��d.ir
N�_�=}�b��y�zj�33�22�`!	A`(WAbKF�vg�'���H��q�'.����+��/$����Δ�h
�&=j���q���dy_#��ԙ�2dvX~�}EE]��	��D7(����r�����G惗\'��,���>=6�������
��h�~�6B��>�`��eF���ژ�@��u��dF@R�}�D�9cS��S�y!HI�¬	^�+b(�sQr<��#%�F	X'J�"�%�L��9�)C����&w�:4v��-n�;wfI�c��A����VR�DNbQ���#��a~�����V����u����.��Ӣի�9lE���6l|��Js���&M�H�����TQ�s::��'s$��t=�΍���T������7��"ѕ�!��b�}�ӱ���͎�Sĥ����-z!@`K��͡Ui�FQR�}d�+��CԿ��@Jr��.O����B/�S��I̍�O���NrO^48�Ҩ�/E�m ���X�t�C������s�A�!���4q�A8�_���!-�c��>�A�1�¼�����}.*i<!9`�'4���ܛA�}%�0��y�Q�9[�i���q�k+�ԉ(����ԝ%-�k���rVýyv�ݑ�'�B�4I��Z���g��#��Ev+̀���3�X3&�#tS9��%&����_��\�r�>g�B������ �+��0��p���K*"�@+@^��.�w�k��_�l��]yʋ;R$;W��M�D��6�����k7nG�\���x�
4��>�~h'��rv5\}V R��_D���?:@+�l�ޱ��m�\@L���蓳͑ �`�Q\�M��w=
(�P,5�����,2�j�*����]�{=^W�������9���dҶ�B\���O4��7L��}L0q��8܇�C�m���ϋ�P�Ù�ʥ�R��r�}1ɧwq�?I{)�-�Eo�,��w�j 3dC�$�/���!�e���?�4���QE(��W\�����W!�iHHA��OC8�>5s�<,k���k)%Il��o�QcF���.~B�c� �Ц���$���+xB�H����ux�z��=a<�0��j���㩡����c��L��,M.B���%~�Kz�`�����T�}X�	�eɐ�V����^$���G�g��ˡ �)�޿�k����Ac���"}�F��I*{��ap���gV��$��YA�J|�����jN�F�?V���V�v�a�i/����>�6ڢ��@��f�rwM�r�񩤈�=����[J�:`�(o%V�O���A�t`�mU��hj3���	��ǠA(��6�������4�s	-��2x�~��F]<����l��IV�[(+A
��FH��E�$zmp-��	f�����M�QX$��%v���*�#�GS�$0/�:g�k��Qq{+'�y���� s,�AӼ*$�e�B�f^1�U� �~X��w��񳡄4u���ŰH�G��Hl�i)*������S�AsΧ���X��ȗ�y�J�\�H��E��)�P0rݡ�Kj�m��;��y;1D��IMÿ��S�8��8��^���M��w���AA���P�XZ���yp�\�W4-��)���At���Y��E�@����g�"�Gj�H
�s'm�\�
�!OK��gj����)o�.�U���:4�፺��pC�6g�i��bEƟSY�����9Ti0(�l
,`	��ġ�g��7��]����"CE狟HN�w��S£���k��B
�mƳ�~�d��h;"�L��ȹPZ�;eF5,e��L��R�)U���� �i��NPMH�]�h��aݍ�/�w�ՂL�Ef�g˒�^Z�O�xT�Ͻ������B�Sy�A(8��v"�cQn�R���a��i9_���~pR.�H�і*�=a�E�m�������"��ɏ�(A_{���e_$��o�鯌�Be�a�>r���K�#��S��ᦏ�����sH�y��6��jު }[F�B@U�US�f΢���`'�R^C�Q���_c��u��9�0�c+H����qp��� D��r(��R�˵�^��kGm*�Mum���JUhw}Ro����rWz�T��<ȿܞ �&-���R�ر1�2�*���t.�K�����Vj]̆ 	���߳E�~޿�H��� �MͿz_��jn"���YeD�����z�Db���ƃ��Vgt��>���⣼�m�Ӭb�ɨ#�(�M�Q�dn0rT�>s�%p#�,�jT��KS<	���~�{��#DG��i ���,$j1XG]�[Y��wtv#60�v=?6r�(�p�!ʠ���c_��g��e��(�f��0SN8�
�E\wH�'L�(�ݓ���%vp��ͦ���a�)J�!��1�p=5��U�f�7'�G{a�}�L4�"8��X@ԟV��+��ŝ�9Ֆ�t�}7D��}�¼+�x�C;%@E�1�*ǵ޺�x�5�	��i�M KI�<4q��y�ǉ"�f�B&�f�0gX�?R9q���s]�����3b	0�![c�.�2���X���O	2s��jl���j}�s4րsZ ��JQ;�@x�W�6U��MT���ۺ$�p�� ��[J�x���KDp�R�j1'�q\����~mB�}�\�|p�cİ����Q:�~��� S��v�DH���d(φ�oe-
���%��Y��ɫwV���MhZ�˄���d�j���%���x-$G���1X¬i�-�ʮ*>��[����]�?�ޟr'�@� kzY��%�L_������}��v/���v�^S��
�� ���b*��2w�17�:.c�m-��.�N3��&,:��� &��J����ՄXw=�",��ĳ�Of�߷���z��*<�Ǒ���'P�jh%�z�#����E��c�۾˾K�گQx���V�YƜ���eF�(N�Cz���9pI6,>��2��ҹ���zO�#7�:.m�c���qT7�:�O�����I����;�N�"B4��^Z~%�70��u�R�A�0�L�&�FҸ�:[��@�oh�ŭ�2nY���r�{����܀���n�@Wg[�c�X3��[c�W�wID>ƫ��dl�Ag�]��r�DF��~�����������:%$���V�[ԣay�1,��׵'k�� ���|0V���y=�o�>�(���1�J$��HH+���L���Mf��~��ɬ�n�I��9H�4���K�����{O4@�U>u��J���_�����}H,ʺ�;���� A�nY����[ۆ���Ό�a+n�ː��� ��d��¡l`f�`������T�`P%�����직Җ#�;I$P�3����ǜ�	��0�WR�{�<�,RK��'����_Ò}?�G���XC�f�.d��e�"�����B����w�s�Y����#�h=A��lmR�B秵"`�2�ɫp�����7�lk�Ǡ���Q`������d�����r����Ӂ�%m9�wЂ�E��uf���S�R�~h�ߢ��۸R9��LB�jUl��DHHH��. ���a"�r%����_/0/�e�t���`��H�é.lƌ�LE��'�H�~��!Q�k䣢VoE�BҦ����J�z��C����n�3"G�KP��1����~[�p��ӡ �ǧ5^�da�$�<� ��,���~`!��zڜ������:��cT�k����TC�En�ݰ���&��ξ�r�S�6R��1�!%y��36b9�.�L����w�М�9K^g+�^��3C�	��b}� Rr\^�?����kb�G�X���~n#5Ⱥ�Y\��$�-Rn_!5���yf��_�#�rQ;�1n91q�.�����^H�vE�� L�Z���V^�$v{�돿�$[��VV��"Og�rn�Y}��	Fޠ�E��N�@+��UW��,�)�촔��u�h35(�.�]w�sxA01�~�i{����ǯ��u�VI&�9�)-�W�`�P m��6��m�������f�����_X]�4Dk��x������E�uHt04}���f�E3B
P���-U%�8ϙ�(��!S|ã딧�]���Ɏ��u������pC��t�A��h{틇3V�tX	h�D�9宲42�B豞��l�9��V�{�i�?�X�1C)�%2_Q�E�i��ˑ���rI�j��p���<j��j[��������TI^;Ῠ�8���'f�+f���
���5�$��*����d��L��a�=��Fրҋ�8���+���Y�	�z����T��q'9�<�-ZX0�<�Wh��˯>�ue0�!�òe����r���������XP���RaXs������jk�J�&�����G(��,ƽ�X��z��`a�My8,}w�_��AؠkJ��Y{Q�8�/k�|ܺ�P^�"�`�81�j�OVvS2?�)Kx^c=ɰW��(V����A�a6��Bc�G+�ɥ�R�F��⺹[I�r2��J`��1��md<��!ݷ��Z���P�>Nbv�b#���4N2��q�F+�&b����|H��͍缶mN3�s����t����N�`M�&lL�0��k�d���|�j$��<�n��x�ɜ�g��2P$W=�gOV��h��m=@'�i�u�L2oQLś�����Rg�pzJ�_��<קN��B�� ��kMv�ߣ�e%ri^k��4���JF
˕S"K�M9z�&�w�o9v�p�}%��J��ާ+���T�X�2��9��Y�]o!��ʼ��s8��/�<(���͚�>�A�l��I�zH�����[��6X�������x������Qc��08�9�h LQ>�b�k�P�f�?�f˳��6A!�Pe��(^�U�sv�IU��]����út(�=#	��S��@h �qBDv �b�*G!je�Y=�(t#��Y9�Y/�L+��W���e8g�p3�x h��������C�x����S��`o_ފ�om�Vw����TB��B�����e�[�Ct́:Ɂ�.�3�Zx�Zr�J�9��ޛ[b0�zG3�	p����?pCd��/1�M��}��CGG�$<I)ų�W���@n<9��$�tχb?�1�Z�j%_XJ;�K��]�b5���e�F��
��q�J����������4�Eu�T �� ��� XF �VoH��q�/�K�@�,�7g���%"q9��x5�iy�V B�Y�֩��)�u��K?=�^�FL�Y��I���U0�����S�{B젖�C����*�G9|��B��}�B�ݲg�c�F ȍ]J�)�p�Ɂ�\Y���Mt�h�4kw ��kK��he�Y��L6#Y���l��M{���DG�����6�3�/l�?�{F��Wf���]�<����l�L�_��C6���2sy�fی��_��9q�����O꼂aM|���|ὕ��6�h
h��47k%���D7_)ڋ�W4]��U� �]�1�٠��="N�	F��שX	{��Ŭ��"8����KY��^<�<�{��$��p2ä��Ye�ʋ
�b8[>�d���ś�l�.��h޽?Cqؑ�Q!.�F�s\���E�{��0x�Խ����N|�ٱi����S��K�ZC�+OγdF�0;-m≌���>Gv3xƎ�"R�]�o�0jC�b,dd0�u��w�l��ǽ��ԣr,�0�q�/�oV,>�ƾ�<f^ �_m �,p�E������˃�탡�B��XB?�������%�����踔t3�����ܹ��,%5�@��n=l���r�44S�汆f��X�?5
�C�x��vk�麦Wg汾�U7�R		���i�l �؅��9�~{
���*�nmB���B4��FT{����q[W���]�g�[6V�;F��ۈt���0;������b*DӰgي!ы��\��W���B'���n�+��d�Tb}�
9�Nx�8d�������	�:����Bk�D|�pj���U[l�n���W�g�Id�;B�%a��԰"�.���[��J�]�m��I�q�aY����qi,�+���;FF�bf�� �*�=,R�
H���P�	�J�(}���̹��Rכd�QJ���X��PRg�����1��6;C$����W�x˟��������
3��1�~���$�6R�Ҿ� ��27� Y�v�ۦ���)/�͏\���7��j#yv:>�
��\�WD؋Z>�H<�|o ��7��O����Ӹ����"������B��3A}`�?HZ<~YW7�Z����4�#'4�.�/}$��Z:�6�ș�s��Kl�b�bQh�"w��C�!#�����[9/������4���,d9��Xz���]@�	�-�|"MrH��eԄ
���u��f��U�k�:�_��>+�b=r9	���j�i"����t�)���#�������t{|�|�%����y���>�TM���s���p��2`���8�t���:������_ȟ��F���fe[z�s@����p�����v�.O�� q~��D*Mb�Qݛ1�"��l�s����&6}Q�n\r���j����ߚeN���Dn���	���7ʍ��΅�K�52j���0JC���y9���
��9�c��P57�ؙ������v=i�.}��#���sK�bBݒ���pG
�lR��9��1��eͶ�G(0's��I2��c8aȉLFD�� �-�Ti�g�j�:Y[�	j.��׬#�R0%#�q�w��.��=rH�T�XA�@% 6�	a��ԵueG� �<�������`( �ca?�"�1��tA����Dy H�$J�~�F碅�{�s��U���$��oN9G��4vX`PyB���=D_*��w�S2�n�[Q�9�\�vs�Z.��k^+���[�a��2z�IFqx_�2���Y���&�⥴�DM�\�ߊOQ���@�t~�t!�|K\���߽/��=c�(/����7Un���,�@�#r(8��j�� aO��f�di���+�t�`����-�D�U����s�8Ҩe?
�����0q/^1�����r5�q�`�o*G��@9���|$.5���*�Fe����x�&���&^)�r�EM�����Q�R ȓ2+_,��n{��� KAz�Ρ��N����+=b"�ռ�Y7�����x>����Z��F�@�E��<��R��7�dɒq�q['3J��x�qw]f��Ě��k6ߝ��b4Y��[t���ʵ �?Mc���b��.W-=|C�U"����f��J~�u���ʐVɋ ���|�]"��i��Gc��Y,���j�`������f4!Z�pv�>������v��=~�������`��'޾�޶㼮�7x[h/�t��-D������X�c'7�S����`;�_���X��A]��9G�����*6b�ԓʛ��W*XD��+ ���T�t
�G�<ҳ�f=}ɻ#!�=?�aS��ӗ�� P���r𙈕
�,d=�@;h��%s�Qڢ��.�zv��T��z7��)�~��'Q�.�Ⱥ��\�w����6i�(
ۚ��K./�5�7.}=;^a؂#=��`A%K�|f��{�%������	�O$x����Yx�LR��\mms���gW�-�<5m�=�����,6����� <3ӳ�--��1�d,�\�s�k�	�bXb������9�L�\@(���#�#�J?c��:�2����-��b�%t�|n�V��ἤ�A��qJQ�B�~���8BfJ���k��w��g�ʂf�?���KǝJ��~A@�Y����K�1�c{=}^ef�G�s�gt��?6:�`o��	n5|\ܸ$�;����O;������?��M;�N�P2�.p�=�+�΁@U��E��ؑ@Ls"�C-�Ι`�����w>t,M�vt�$<ièjt��>�p.�S	T�/��&N1qF8�bX��}2�+O�Nqf'H�t�33�	��֌����C���/��,�2��j�`2!�w�e����{�J����bxi���\��pO��yߧk��G��鑉$ξ�-��}x�WU��#��:�|�VxHGX��S�Gx����=��H(��v	�
P�g�뢓k��|�K�>����!�?��KK��v����m?���{:3?ܲp,@��rsn@У�[ȑ��j�s��4��t�6iW��.�����%���:�{u>��4@�:h���#�ۜ�ݤyo& ��oܜJ�����MR�?}����K�0N�.�|^d,
�(�:zX�K�`U��x��=T�=Dau��k4��})Dz5� DSB����r��G�7QQ�	;��IH�JF n��1r����#���P� I6hѴ:�+��rM�r��R�BPtya̯����8!��|I`^�3���/����LBW̢��|Q�K`��u�-o�*"�Q�>ݱE[��0\�	�F���n�E<�5Ǳ6�� �U�ܐ�'���h�U�J_�ܺ�ʳ����{4|9��U�}x]��[ӓ�<���|m^��%����BK��V�>n���41 fTU��� ̦=�mܼ�<dZ(�
��BQ]�Q�����P�$b��V��+�,&c����@�7��׹����ն����.4��m= ���b�s)���>1�S��ó���[�������Ns�M�ac�\<!�&�Ӌ
F�̥����TqM�5q�z�ۧ���"�o��x�s{N�Q���;r8��X����'9U��V��{�H�Q������p�f��&`D��H��ce�2�r;j�v��Ô��-���3�CAl�PY�cɷG �} 
��u�˷M�����g��4�h�m4Պ���r�R�zM���B���7�c7X�T����"�E�|%w���r�6����e��(�\�P
����1����,����h:���t(6��npKGz��&8�`����k|���l��X]�<[�`�ߎz�<K��̥�}Cc���F�P�*�oď��@�\fq�g�p�0���wS��L$µ�N�05"�N�:�I��"���Kf�&s�n�p;���Msv.b���5��_"��r��s�"�x�d���<Y��z��LX�J�4�nƁ7��9��Z}��5�!'8���]ȏe����f��v�R<�+��@���+��O�Ɣ���#���w�ϧ9|�7��
��2�ҁ�|�[2�������|�K�J\��N<�z���^���:N�OL��������Ik�jg�9�:��+9����w"^n$7�x��~v�ɍɩ�a�m��0���O�nE��[H����	�>kݠ\�N6Gℜ�»�L{\+��܂���-���N	?��-�'{�,
�{�Ǚ��������okcT�F�nUk��V�On��;�,�!�|�Ftx���5�b#���Iz�'7�GG�c��]�T��+�z�\�k�W����[�^'ǡw�u�wA9kc*@
SbvhB@W.�*i܆��;�V-M �9TL�p5�b��A�G���v��F��2�Yٗ�D����Ϟl����?e��v���g�jG;��$8Ē�� �	�B�%1\�Y}-��Q
��>��$��OEJ��xkd�0�Z�f��S�ܨ2}���IFB<��O�WH�'����,����J� ��]�B��D��3�.i�L�5�l�E�4��(B8y��oF��۩Q�)�_���#�6����\)�B�;&뮊��	���Ӭ��󥲶nA��$˅n2W<�Z�9Xdy��� \
:^;�	.���B�c��]7��9Z������x�-�]�<�u�|ċ"���@)܅�x7�T�ι?S���>؇&(n�Gy5��?��{����**;�¾FZ\���-t����z�|��y���ʩ\���	�ψ2!C�$p�Z7��)��+N�0<���P=�s�>�QjPi6u%d��J�7�����=��{K�vp�?7T6	����ƼY
\�z�&>�u$�-�==�S�6y]��b.��~�($�txg���D�҅��y��{��}��L�o��'���uf��u���M��I/	�B�~JhǷ����X}�@��a�B_�Yy}۸%�=�u�\��{\W�݃+8(L+f�K=N�3Ȫ����uU:V"���Q�S�w�����юh��.7T��y.\<$�p�F����׶�z9�ݑ:~�1^��>�Jl��q�<�]���/�
�������/�Bd�g�8H���Ɗ���L�c����,���v��ƭ��\��j��� z��ySu<���|z���[x#t�/-R%�컱m��U��_�#� ��4�^ �5�r�AxU���\�=��zwAkk��X��OYN ����c�GBx�TIQS��/ʆ�2R>A�K�c�ޢ�a]P�@?`�(���Oy��y�6S�
-��gb�?����%�%���LVW���7=x�\xh�o�����]ʽ���;"e�$�r�޴3UN���������1C<�Lx��/�`Vc�(Z����gC�r����s�������'"@�3�Q�bi=ã	
�^_�$Ұ�#Hb���Ur�	����0�u!�A����`������'3���	�]�կ�@(2��.w z�K;�Y��"@3׺�u��G
�]j�Z�bm�′���)�b\����wJU}�u;��PLY�иx�y���1Qԏ�.��M �7��	�y�ܟ��d/Pӫ�/�����=Ӷ�G������!���N5�S���W����p=j�ifv�m_}�j~��~~���=b��K��H�m@� �B���O��1 Z��jI��
�T1�?���(�aA�"�^�Ed�w�r���_Sz���:�?�p�p�9����M��,�a��+R�/� �I),��0�Z��ܥ�f,���ᩪ��X�D�L� �}�b���2���Y��������K#�'��,P�u=���V^�Eי�V�B��d	
�V�;�����8�fGF��؏��";�3B�W�e4��^��,B�mn��[.X�0`�#w�I��E��`�}%��Y�<�`�mk������g�{u��j�7"e����ҚA��ȩ��g�F�9��%��_�ie����*���� �K��mT	P���te(�zs�a(:_��	���t1� �pGz�@��q!?�Eݒ���V���)�5Xc�p��k�`YP�*[L(��Ed_�S&�<����$1Z�|J�&$�y ��l<����ڤF� &�=	㉀8�V���<��֧���>�A�5�/����fwJs��f��O�W��%�VAt��ٸ���������D8:)�W��\VJ�8bJ]�xG( 9���U\,A�wgr��k�ɣ�V4��?]s+�)����$Xjo�Z�������}�T�k�>�$%�B2ɤ�}[�dz�	ύ��bor~�$C"�Ex_ds�x��#b�~��eF��B6��U��}v���Iq�	|���s6Ը���Q��TpI?3�t��X�Z4<(�Ѓ��� �Q7����K4}��	���m��ܼ�&��྘{@�D�o��eK�$I|��"�py8�t�>Wj��7@j�r�FA�	�@��lHN[���rZ�xŵ�I�ٍGvhigU�����$'tPd�*c�S� [�k��.['t����z�xk.ex(+NK�=��*�1(� �}�jЕ|�p=�]O�3w� x%�v�ĸy�k�dH��k�G��k�L5�&��Z�z�t6P�m_�M"[����X`�9b5���Tos%T�%ܪF��Nļ�|Z�R�����X���|(��S�J3�x \�0!�鬳 �y��!�~���O�j��̔����8�q��C�r&B��s[+�����H�방e��5�	��ӂ�P�I�r�3�z����Z���J����/�<X`X�o�ܪ�8?��=���ʦ��ڰVCS����jv��zp겤�����L�~����n��^���T���P�[�;�o0�X���{-V�� ��bI/M�%S4m��h,'Q���~h�}l��Nz�HP�C���&	��}+�a�2�g}��o�h�t��� ���ȳ�;fX�Ѡ�����{˗�^�P�U5�A�x�eQST�_���[+I>�����w�� ��'��n�@�N���nP�I�-BǍS)��5���t-�E}�L���g�R�U�Q�륉�r%
9�1��	|�S}Q��r;�._>@�1���O��@�ܥ�̎��R���aK���s��a۝%<(��	Yy��q���ըڄ�I��F
�n5���V��$���sf�^�m�M~<$n�0��%i��l�}����Ab�D�0��(������h�+�/�DU����g']�0�_�I>���jy7F� ����JCD��̡Ѐ%��a��]2J�5g�eN�զ�Ѯ�I����Q��D���B���aaƿ%��;���o�`ڲ��r�e�()A4S�$�%��z�T$����);�?���́���H$��L��Oj�K�}Q}�J��z+SY;�R�+@�d6��8-AtS��J����{��ey����IZ#��S���		p�2t��gQk���Ʉ]ו~���6�-�F�$PFP/�rZ|�{w�r�:�ޟ�������q��u}L�%�O��Pt]E��� �μ'+�O��6�d*�!�_N
v/Q0i��k��eҫE ܑ�g+��A�ރ����|c�?���#q�$.F��fi ��ay>�R���Ѯ9>*@z>� d3O�; 7��?w1�|�
~�6�r�PD���z�Th�p�\¤�2t�8���bc�+����̚�}�/�ah\@>C�0L܅��ꀃ��H��K�O`r�M×`a/ �#ޣ���lH7�I)!��wS�����s��8�����L|�%,�3���bj7x��ul��6$�*&��r�<z���#�e1��\\&�P��Ȗ�A>��vy����y�RӉ�RN[^s�R�����1g	�R�O�Fg��fX�w�I���82��A�4kz�]S�<��j���c�l^]E�@�;�@-UU��uᛝ���u��ܖ����6&���+b��y�5�f��!5}H��u)���$F��\�*�	�i�~���shE��ET�vA��b���;)P�#��`�� ϩgdq�6��_��
�ju1Vx]��	�;���K�6Hٲ]��������g�����!�"c�]#N��`�삫R���S[,��Fg�og�D� �����p��h\brJd��l�J����Nk��/ʽ��t�fh�7��Ce�ʑ�a2�l�J�un�Vޒ��\{B\�qI)�"R �k�=�n�Cʅ~�������@����UC��?�vZH�O�9�d��/dbR��| ���Ec�6�)����{Ҫ�\���6bh�4�,5��\��)������Ḭ���j95HP7D��5�R([��������H'�z�N�8Vb7�B�P�2�����e�h뉯hO���U$�*Y�ń�U��=��E�n����W��*�ڊ�L^�S����H���/�u5�9�o��}�,�k���a����c��/���rF.�������Ig��s�^���tC�4�%��
X}m������7��B��8�d@���Y�{����l,�F���ȥ"����In��S<Z)�X�j�#�q�V�ժJԄ�N�yCG�Z=����Q(�2���wcz�3+~���}E)3`��j0�/�c�ߗ��? ���u?��l[R���l�T:-4eNB�+�ï�VK.��S�/6��#�*�-dEO_)rOQ�l}:u�Z�A@O%������d�=k�n�S��"n[���%I���E2bPHDNKҩ?�2p��Q-+�V��J�E
�lY�%�P�[B7i���=�%��)|\���0��P�����������Q�P]���<$�^f�G�j���!]�_A�ּ��IJ�>�D��G��]��vT^]�&� ��&�d�z	i�)	]нP�'�f4F�������s��2U����3��Q��7M��RqЇ���}+�Pw�}�lqȺk���.�xd�S9e��ngr��p�:)O���
���&�Z�,��0!�8[	�~$!ֳ�r��t�+��J��-F��b®5�4eX��\������"QII�����GXhuU�:)����a�=itf=j�O�z+Lrњ
4E��\x�����: �t�M]9'b���[[�}&�����K�:������ρ,D�¢�.�ܺ���ɇ,n�Į�w�]s�����k����#�̋;C�K[s�'�U�+������L���MCˤ�-OY6ȋ�}5����$w�Dy�r:� ��z��J���<��ag�N��e
<�Jل����l˹���>�6�
8�գ��9��2M�D@�Z�2CO�=�U�4��~�By8���E�%��~��<��#RV�(%��WR���sOD��-#��	��L�?�W������\˶�g�i��Q�3A�3Ǎy8p�[��?�t䲔c��{W8�ʏ/�l��S��β�����a�'��v�`5*7�u�54�=*"|��������[{9��`����}���/�H�T,ܴ��h�M}F �EB��ģo$y%&2J��|�����?UL��@��(��J��̖8���sT���:���k�Z���n�JԤdIdS�❨�5x���ĸK��P{�#N�q/0)�#������C���]|����F$���$�%��.��}M�xH��sF��ށG�������Ys�������m�f�P��l$MTG#]����+�����:��Խ�~'���{�T�!� ��$���g|CN7ƾ�?�(�u��-v�A�xU���ݴ��)��oU�K�����P0¾�;�gM"�j����>�ޠ���L��Acp�����C�HN�£+�4��5��N��q �z���[[���B�\��UW�1��t�xz�EZ���5����R.T�|v�'����H�Q���	x/�#�������}��I,�P<��j凁�8DC�tւ���SG׺�t#�Tc�J.a����-�Hk�Y���W0�^ckuv8���C�Q���D�vi��9َ��D�2�0��4���U����s�������R}sD�� ����u�)+8f�Υ�޽h��:�)�G^�,�l�w ��^��U\�n�,��qyy�ľ�6�W�b����������z�	��1��[�/Jb��W�0��)�"�M˩oiW�_%s�f����:K;}���0�W��{L4���?��22�L|q�m�H �g��f��ɤ4�����xG(DSŊ�eNF�:9�MT�<E/�'�|��snczK�'��`��kT1��������I].�,���� ?U�14.������u�����u�m�j����D��ͬ$�5Qvi���� �r���������U�1�<$��"(�v���
~�Cj�8���e�^���Se!��C�K� �Ua�W[+���,Չc^��ˋt�/�Di��"�`{��#NZ������T�V��_>����Y�IR`�[ψ�X�s]�y��O^&���Wٞ� �4q*�X$g\��)X��VE�_�C[�?�i�u��
���26�	!�g�5Ҧ��ӊ]�u��7�4�ҫ��X������.�\�3v�p��՜�g��V����_=$Zױ�jt�ѐ�p{�^q�1�!$��.��)���f�y��N�v�Ь�q��ykY��ȅ7�;��[6�o[�0����&�� �Ro�\ʪ��'fh�9�%Ƥ�J=�gY:�nL�[��ۖA�;O��އo`��ئ�y`b�����a1-�s�E5.m^���hol��"�@-�*�	�n�p�z�ۿˌ`�%�^��L[3���gM��XbcU�a]{m���:�� �o�3 ½�Mh�*fr�\���s�C�ξ�Tb>k$�s]U�oQ21���N�X��w�8�\|I-�;<���9-'r�Ȑ��䱷m1�¸�2.��j�c)�_���]���M��0 �o\�K���s�eݾ�k�E��&M� �����'X.8�����+@�[n���#�D�֩s �,���]Q���w���,
�aU�$�3NR�b�U��QXΪ��������;����{�7�T
��;!�Qo:N�,Y��B��r�9��-�AZ�h�T@��_�8�!���Od�y�c�b����a�K�ۋ�[�Xz���G6�B��k92hrepZC�k~;�ӡ 1Q�M}�2CO����w 5�)�v$���:�3ok���I,H����hO&V`��)�gg�D9��}"�)�޺>�a��j�׏�]5��^G:KT�!�7\��ւ�>f�%޸�LI�&kRoi1���{#�	˓`����=�xf�=L$`Lc�kf6�
bm�h��C~���⢐�u������{(���+W�S�������G���0/	�^�,)�K�eד!���3t)5)��r���7�d��0\��ȑ�H�����^�ws�5?�|��L#�#m�Y���%oV�W���,k�q9��,0������7`��@{ǡ�o��`����f0Rkh�؏�kmy����ҸU��U����q����f�0f��!�]�,U��e�:y�&c��x)��r�;�9{Àp�D��i2-Ǿ��S5��j���7֙���O2�����R���?Y�trɯ�lS����/z}��Ē�(�%qv��iᲩP���07a��N�qȻQU���K��������|DW�8+���Ube�'�R���7� )�`��O�󭾖���F/���<f�=�r/T\p�Xv�f���4Ӧ�RW9�x�����o�&|��(�Py,}Z>�ȭ��W��
���$b� �d�{ʣb�?|���u�]�m?�a.�т@/�b,�<���-;��_�tfӾ���V;.�/�����O�j�����Q�m��p��� �Nlf�P����3��)>�yA,�K%u����(E���u'ǑrVJ��?֥+dk���̂{����#Gn֑��_����[B�������,��v�ǩ������
u��d6u�$�Ɋ
�Ek�>����	�x� �$%�J��p~x׬c��Ԉ\�v�g阹�Q]��ĈyE)g5��)�@Vs|�٘��,��~�%	����,�4J�C��-�7n��Vث�[��S0��I^��½_��r���LC7����K�4$*l�S�΅��d|�$�&���\ �X�1�8�J���'R�[���,\Is��[�D�uwⲦ@ ��ޢ�;n��e����bE��4ó��z��Gh2ۚ��D�?��:,�d�)A�V�+I5�ٲ�{�u,�Ug�w�����Z�=LAèW��C�X�8��V��|3���'[�q�jf��X}��R��B
Z�S����0t/�j[n��09*<|9A����$�@ �Q�|�4�����Tr�}���x�D����{U����Yj�M����6M��y`R}�#������z���#�;�ك���E��P��#���%~H��C8�[qg�v��.����t�~�b+��?O���r%������+il�+<��~b:&�Y�D%��@��SgiV R��R��]���^�pm�9H�*�T~z��΃c�q�6�x؂3��u3�r1���:��|�֍�^�4�u~�/�ojA6'֏ո�d�@�m��^R�]��z�A��;�kQt�w���1����3�|���\��E�*�
�Q�L��e���P'�5��b1H�N�����D���(�?�:�(��A�u�"˰�>wFt$��]�(��+q~������ٺ��� D� �o9������>�*\�%����F�$PkjF��T�ϭ�a��pz��[Uj$�t!3�2ogN0r�`��8`'x�B���5�I����b�J�s�[��j�^5�>9���W�t��Za���~���������.��@�rȫ��v�LKb��	�!�R�u�'i���ߊc�wd˧�UH�oFn����]$/��e����L|�,e����Y���oqA|�[b�χ�H�ϋ������&�@��}��HyO5f F�F�V����:Α3���h��󪴿�
k�9��y�5���$)5`9K��?�jM�!�6r���X���k��1�/�~�-�N��ԳK�=}o-iu|q��.�*�� Z���w��`O`-��&���%�w�n�eC)�GX>���ٟ7��y��(��2�k����t��H\w{̀L�hѩNy[�M�6k�FpI!?{՚٭�|Й�?�:�6֩]�� V�8����M������k����6�x���$�;.(Pu�S�CqZ�����K�%&O�,�<�c�m�/ʝy�q�j�T��C�����=�����;��.^4����g)ˏ�a�+~G³����c%���=!�&�M�+A�������G��	܎��i6��3��r�N��m��p���9<e� oO�q�^���Xe���O���oW�� sYծ�뼅��AɔF(��_\��ɫ��	�,-L���X���h8%SجtP<��@Y�xU�c�C ��:���M���~��.�H��	5}�O��#<�Mt�p{�4���W�!�� ]����p90b���f8*��M��G5�-�V�-�9�Mpݘi[��Q�|Sx&��G��s�|kt���+०K���p3V�d����(��r���D�x����$��=��Pu�d>a�:�`�y�q��-�V��Ƃ��:2��;��$}9��l��ؓ��~u5��Ꟛl��n{�W�Q�o�M"AWP���Q� g�5��Hn��ؔ)V&W]��}��H��W�3�pJ�g"4��tñ�.�,��5;!oZĐ4�>�L��8�/�!�¬Zi��"�b��m�ʌ	����s&u��S�,���� ɴ	|
ilI��5��0{�P=��>�A�t*���FhdK��+���#ҵ:����{p6	V�lMʖ;����+{o"�����efdR��G��m�{��ω[B�]���#�t})�,��!�6��f���f�)��X1{�mǯ��?���|�!%�Y��
�-��4���	-��;�����٫�@�ï(�a4D%D��w�N-���t(3����¬�phJhDJYJ��k\���OL-'�Ơ�z���q�jX?O�5wL����w�Ҧ; �ʋ�f���O�����a4�ʀl25��[�9|G̷�F�|�@<O"W��A��𙱃Bq�E���4��q���K�ZM�,V���0%Ы��Ƣ���-u9r7նG��a��gP���arJНʚvx�U��?��V=�@Pb��Ꮽ&�ݮY�n?63E�@�VyH/y���gQ�6IL�n��v�ǣ߾}|#45��|�Ij31�lC�QW��|�P���H�=R�Ǩ^h��${�E��l(>�e)z`({N5��r�,��j����r��+12~B�⎉�D��'>� ��S�e|1F�&�`�^�to�>��c>�=]�;gj�E�v܋��aB�_�z����-@Wj����pZ����71��N�V��=}�+�0�+F�)��.ލ�4����K��w2�V�N\:}���8CY�,�ta47����_2�kc�������''�C�d?���pgc�	���'B�E]AMڝ��oJ�y2ИYH6Vi斒���#{�+�!hST=�r�o�F��g"�@�(��j�'fz�fAV���飜�MO�p�XL�Q����:��Q0�z�>��m��f��(.�(���lB!Ώ�a��l[�_�?��o�洽�qK5.y�4������+�+��(�r잹����M�tI���DNfr��Ρ��d\�ˏM�>R�TaQW��K����[�c��XXQ>\rbg��lح��[�-��!~Ϟ@�E�b&m����
x��b�Oh5�qo��*�*�$�d�	1�B�����#��� ����^�l��"˒�H>�Mո���ǰ���(�X�A�sa�*���'u�Y m�_h п4*N�l�X�2��iр�˕��6�YDD�"��d^v�Ddg¼���c���pݳi�ߪsY�C�c��#�Ɏ��&ƻ��׷%��CN9W��>�#\8+�z�'���J\`�@o,v��dX�ϒuqP�Nbs���H��5�P[#�b��POuE6iU�UL��Kj��M�|�%x
1~�;q��Y��*��e�k� X��7"����۩��賅S9{�[�o� ���K �;�b���R�o�y}��v�������vy������Z�Θ�IBX�x�29�0B���df	��:���8�Nc�V�E����Z|���|�|�m�B���M͙!��lzn����|�GR���)�C�K;e>I��W�8��m�v��ˎ��-���r��/c��g���Ũm=U1K������C��J0z���ıa%%3mh;@�4I��U­p@�Wh�:�ɀo��G���P��4XKg��)K�\�xm��S1�0]�bpy{K�F9�mA���������G׹xw�k���z��.Czn Oiy+��m�E� z1F5�Тd{��{j��0����^ܔvu�J��[�=Q4���Y7���8[�˙�8#]��$�|���}E��yi���f�:I�k����V����l2��ӻ%`*ܲ�o�]KIԓ|s��hi�W9\_�Q�Usn� 7 ��ʿ'׳��ϩ9�o��e���V�~�5E�U�5����@�sh?����o	�;�_�>Wcw�Z) �I,�&n(R��N�R:Bn_����f �]�s�[t7�M�����oB[�DU��@9bO#Q�6��#�#����pI�}�RN]�B{�4 h��'U�ǭ;ݸ��kWy8y�E6��c�ϖ�Ց��&�5�~����6+�/x� ��<4�"�;ު�Y��W�4M�����+�a�t+Dw� !?�i��e��sW�""T$m�h������{1��\9K~zk�) �k��_�|�I�X����He�1�U�k�s�0C*2��yi��an�a=I��Y��$������ß5`��5ka'�o%�c���iSx�-��-)?R݋�Վ4��}�4kg�T�*����I?�q��8��1}I�e��_iyh��=!�i��Z�lb�O>e�Z`�|��b��Ə�񄴑=a>���79�%g��$ʐ�n��x�G2݄�~�K��w�+�{c�H4�XnT磌lI�:�V�3�q�r^E�{�wkk� ��(�����	Օ>��	ɨ��BRW"�/5n-D%G0��.����}i�q��&�x:�������ɑ�%T�PZ�Јp
PM�:l\���
<��*�3x����Q(�B�2���Q����,�@"L7$�Rw��	e��nV�� /�iꆫ��Z��(҆ɕP�|
�U��|���k�:��͓�{�����8+�WgF�iAc�u��~UŗI�|y�������Y-��F������c%LF���F���"~O�d��H7NZ�!����4Do{�!��t��o��u99C���Z�﫶�صnH`�S��pmݐ7�|����aHQZ�Vu�Vv��>��s&��N^����γ�� �������ݔ+�'f+wz����)�ś�tЋS��\���^χ��[���k�#:q��<-����'�4g�;M��ƶ{�����}M��AN�_iR�`#\M.�wh���"�>�����}�B�{�AoŦ�8����N�K�n/�:zEL'�N]J����}n�Z6�UW�����Ep�u~�'�B/��I���ET3�醛�*�����-�#��� 7��:�#�"��(^�Q��×�/���I�eR��s�B+��.�q��Ί���"Z�i��8��|u� � ��E����U��M՟��h�ڃj��[�Ɵ?$���c���P�QԜ]�0�n��Ќ�_�X��cF�[TM�*U�q�tyx��g���ש���M�L*�	�����3Q����6~O����\���=���� �!�g�F/�g6��fD0������pj�b X��q�>����1&�9ztڼ$��#�9ΐ�c�bN�M�r�u��l=@xT	��S}R���,�|Q
�ç®�$�3	�j��V�=�"�)��*�C�O�Ejc����/��O;�O_ȁ%��x t�[Z !�=Y!�v�����K�N������_�ӹ$��gJ��!iP#ڒ|�٬�),P8_[t��pL��k�j��p��;?�o�uT��4h���I��y��g`w����� q� � W�0�L9-G
欲�m�����&gs(�c� .���
>^ :��aM�zL�ga��]r�.�3���E���.����hQ~#a;Ejg� �>�=*'`X (>�D3Q�ٷ��C�3ڞ�Li�8��|�@��4⸏��,��d89���ߺ���ƈ!�7[,�'��aw����U�c�-��~��3������Hi��]�O(I��S�2J�/�e�[ "�c9���C�=�QF���	�:������O0�Nj��:�o�[� Jm�U�let�/_����7�������x����,��6>)k;�l�+�.�ي0��m.4�H��'���e�ߎ�^v��5�������#�8Q��nO�Tͽ��R��o �]m�,��$�cj��'�+��8��,��Pײ*�sY��
�����Om�ޒ G�i�I8�f��}bJ5�!G�I�&�Z#���DI�m:W�/�@���3ҏ�%-:�q/�˄�'�U��As�J��^�f �
�H�z�8�ب�wgx�PP���)�����=#T[��n��I����~j�v���H���/}sB�o��1�i+��l�Kw(>��QcG��J$�߉}�#O:��$+އ��_SCp��,\��g�{Ӂ1�z�-�ZrQ�QRN��ސ4��	XK��I�Nl�Kq~-����i���_�b����~���!j�d�� +H�߹����[�����gS�i�����6����bԻ%�U<{vݨ)/B��p�h�1�Rȝo\�8�����~D�w�!�3]�>+:��������ShJ�6Js#p�A'Wc���C�AGF���J��8�DSk?_�� ��ಯ�HoT�ǂ:��<Tr��R����=�f�͇��"·�b9�@���xµ��_vG��	jy��/�/�%��O��d�0::��>d���%���8�oa�OIFȴr.䕊;-�=6# =ڿ�z�8��o�c�s�@�?�R�hyѬ�oJ�|�.�}'`��<b.�uN&i��˳�a�Jܓ~���E#�X�v���0FsHQ`ܧxB`Z� ��nݒ!}�#���$��a��vQGΕ�f�Q���ҚP��7�g����<{p>���E~�k��&g�5PQ�@g�ko���H=��)u<̞�I|fi8:�O5vw��(���2k����,���CQ?�x`]ʲ��zsU���p8Ґ;���Á�W8_����舏<w���p;����D.��jy�z3�N&b�����[� ��~y�8`B�R�mT;/�u�$G9�P���iz H�(�䀛s���X��}�\�E�I���>�8�(]�oM�K
{�D>o��Rq� T��Dsv=��7KQ� @���3�Sg5�
^z��q��	�� �ں�H� �I�64uO��Oģ繇��}�6�٥�'�@8!�*2�P\�ڽ����. �����E;�S7\c�⛾4 B���hM�KN�es ��qf�ym?(JL�/��RS�v��,��V$J❙�k��L�5b-*s+����My�G�'���k��؍M��7#�B`�������-�������ut ��J�R�V��`���¤�D���H��{�t#��#6�/���N:�Q�:���W_xcC����ܷ�e��y������H��^uX�hKI��?�`I�����yѵr�%��삳e�*��e�4�!�2�/YR�5�O:G���!+�H�����i0S++��N=��.[j<b��}��a2��>�-\e0�S�<����ˠ�V+=3/{� GU����ۙL�PD�A!�t�{E�/���3�}A?���J���cș@�����P����N+��1�H�xI!��.��]�E���8JF@��T�c��";��;	8śmX�]�3�;���{�]x�,�߲`�pG~����]*蝷��j.�2ǽ������[�~P9���F?�@��~�����O3��yU��=�K��]�I�A	
�)u��9�Y{
��u�>x���s��'�aɧ2xS�}���^8F����>vPϕ\�@�o4D;s�|sB����% ��TD��9p�/J�����<c�Pc�A�g����X �^�F�/m��M&�����n���l(v �Ptj\I&_�,nk""+l!Lm��n�.��>��߆7\u}�p�r5��a	���/��49���[�[��)�[�u���/�Al�8<�LvL�T����W����&�8P̝E#�Z/)8�V�z%V,��u'�E�O �r��A�V9����ē��)F0~>ҵ	#�U:�}�J���r��u�?^b0y��N�����o^wreY��h"&
�K3�4G��!MR0�b�A���^�&����>�[�0�+�X�}�?���%�
ȵ�])�kg���e����[M,_�� �jD�����h2>���IL��Xz߲t�\Ozv <h�p\��'���q�['�0�Waxф;,��|�!Y��1�@�^*�(�qj�tp�쐎���'X��Z�a������ ��LY����(38wei��'�"�gn��S����������Q���'i���jp�8O�\/�}<u�RΥjuW�Uk���x��URp;��K���K����}�{�
v�|��s��^�Щ�j$��z�P3�YT�Ǒ6���*H���
�7�����4�Xb��l�M�� �1�-S��٧�x[*G�(WtǍi�s�^���c�m��_��Gb ���h���j�g���r����э�Q
d;��c�V䶰���	iFB-l.����X�f񭯄Z��h�54�l�j�т���?�C�*��~��o���x�	bc����ia�e*��&LuN$U���9�h0&��:'����lU��x�R���26<뇷k�ʹ�>U9��4��0�Xt�$��G oG�@���x���T�j!m�V�7<%A���Z-�w��-U |iL��|H��E�/����u;�$���Hh����2�`��u3�u@M�R��,/�/p�,�=qp�h�	[��R�@��x�Fk�hF���-��O�K$<�
�GFl�/���m�Nk"#��C��0* ��fi����T�:�/]��ED=����0�n/���3plPڹy�5U��s�g� ��H��G0�b ͨfi>�!��������r5GW�}<�y�eЈ��B-*v2��1Y�}��x)�1��Vp��֏W;�HD��5�ͭ���bg�
��q�w�o�xw�u��m��QZ������K�!* (j6zGAc����V�����vv��L�^���H�I$^��iWm�Q�ʏ�L��4@�ijO��C^"Q㒘c�tlyH6C^_\��n'���q�Ck�^?���i�ZWy);�Į��7?/�����1��JM�|;�&lݒ��P놳;	%�d�#����	�r�l���E�SW��/O�#��pLV��[��UI7��3�����߻c�U�T��[.�mYr��Ǵ���?f�v�\���Ŋ�a��V�c�	�,׺�����H!R�z�@u8��\����Foϐ�0t�	O�om�kA���16� ��KPHV���sI}&�M⦡�+՟����q�H5Y��zBl:���N� tȡ��Jv�=����Ǫ�i��݉�+,��%�52�=j�k(|�^�/2PE��냏�-��]��,�FٗN�~I�� �%����J��s�"���X��5%�&.���yv���Ca+*���5^3ږ!̧��@�
B|ge��-=F����l�.��Y�"�(/���:��n_K/D"=sˠ�>j���	yv���rY����)�F g�߹���4ڬO�Z��[�}��Iu�0Z��>�h���pj��r�4<��H/G���R��w��,[�I��u"�3�c��=�5�+"�)����E9�<�
��(? l�M�q����>h#�����)��\w��PqwH���ҪٽP�����ȡԄ����jl��k{r��H�������4��M��Uk�G�,�2��oR4��x�h";V�����.��d���,Q�DO	�d��t(�%J�o�	n<��Q�r���P�F�+�{�ZѢ����/]�a������3��B�s�^|�&�@�VW���So��q�w��|�GI+�W�!��Q���b�cc�h/E���v�P80��a�$E@�k��m/�ݡ�<L c:�Q"�9�*�����3��T6;�Md\���X|����Xn����6�J(VqAÉ�E�BA���?�q�u�\e���50��H�{9,ǭ`�wRl2�B��v�+�'��}fD�̥��\ȟ�j����Bw$��݂ɚ����dVRݭ���#m�ueϹ����HBݯ��h4)��:��_6s�r12+�Q�x��J�lc_�Bx�5՝`v*�"�����y�T���c�\sv|'A�"#��84m~�X��M�؄�N��l�eFlA��H,b|�X��D���qݕL��^�ȗ�/�]%A�l���?��ʗ>��!�~R�`Y*�!�������
��g�{�ȍE�wU��8R�!`P)��{��x�;�
��.��	�2R9��Ɗ@�\� i��͗��q̈́�A�E�L��w�
�wʳ�Ȁ���%xZ7T!'Rm��A��P�t�[$o܊|�ȧQg����ʌ�c(�m���ը�����Mx� �@�n���/�����<�D�2l�g������Z�9=��X�R.�*�"z�Ꜥe4��X���!{;(���;�ցu�����,*34��x�$��3k�V_�`�!�Wl��x<W��ah�Z^�Q�B��+��R��m��DLT'o����{��Q��v��4Ӂ�γ�/�1( ��qڹ)�P�/Zz�e0x�G��VS�
��#����ª�E\v(��)q��tqw�������X��(�
�4lM_9;��.��ώ���dգKdޯO�+ �мݣ���5�.P4ʔ'�*�R�uk��a�i(31!���~:��+�S|dEK-XCcZP/eGB�D9�2w�I�'��5�68�ȕǕ��#��؄~����O6 �uQ�/�I�R��7�ј���b�y���{Iޛ����}�]��4�+p�0�:>��+0Xd
7�N)k��U�R���3윢�6�H��y}%va�����2���&Ѱ�M��|xf.X�uZJ?�L��K;6
� �YN������V���+�d���\���^��u��v�c�ӫ�j�,'��e0��f���}�)"� sB�6�{8-<���k�c��ݛ�0�`�-�E�iF��je�Se�/���~^��a�|q����U�~��1�8I����l�����M �H{��aDطQd�����}�J�u$�u����L��x��	��%�X15TMȦ�#<)�2�B�=�W�n�,d��H��wa"��/��4h\����se���7�ߚ���\e�����VaV~�q�J�\7���%���JJ-c5jm���������s D^���7F��� 5�'����R��ɮj��D��'CoK���z�~4��s����e碿�%�^��^7�d	+v�r��S1A��0c����ޙ�UW7ꗅ%����k�>����g�ֆ:�x/¶$�9_�1�(/,X����No�Gqݸ��ǆ~o?��qs_���f���f�+a,J��+M#�kO����S�<�B=@��RH�ؐ$��	[Q��s��Qx���ϐIO����.��1��&^�ەZ�I�;o;�)ҙ�X��F�IyOsP��{�#u�.*S�@�s���sv����1x}�6ilH�8����;�*�j6�%b��D�ig]�?Ap(���;�7x�+N�8���)?�Kz��҃�s�K���i�֐���`��Z�5	;��Rf�K1�����:E��<B�����ӤR|%���o�f��6� T��%U�c-Q�d�pё�60bX�m|���S �o$?��ǁ�,�x(���1�ͷx�8wi�<u�lNe�'���@�Xt�R��0�1��Z5����>��V�BЀ�Q
��S�U�}�	V�Ti�\O���`�$�0ɚ��T��(8⡡��*V�u� �B���R��v�=)�a/ı4����l��qET�)]u�,VX'Z�6W�~���v&s9=�^�̃�d��w5�[���Ү�E�I���E�������w{d	4�������#+}��to,K ������5d8E��+�~�:�IJ7 �wy̒t%��r|�l�Iԋ��-�H�e�
�?�v��RAPb�����.'E�{�;E�>_��B����L�%���N�7l���i���u����);~�_eݵ�͎n���'е���I��	��PNX�o��co��)���v#�T��vM�� �c�~��pv7>
?���:�<5v�y�xg�x$�@��W�'�F���N�kt*~@-"w�B��E�@��*.��|!����o#��!���AV_�-?(�D֌@ʖOS×�x���UݫA@S]��H�/@m��7?��Po:�$��fīD�
w�y��o�1����h�Lؕ��LS��C�UO�Z�K�%ˤ�����  |y0]lgb*��n|s�EJydi9��1�O�nT� 3�����eM7��-��hzN&��`<���k"[�|_,Ж�A���S�np�t��^�Y*F'U��}�0��1�	7��q��Sw�r��&W(��[�;�𤜔?�K���D�W����5�]���< �rO�u����*m�~SsW�ƫ�cqׯ4�ƂȊ>�������j���@0��A�Jx��3�GW �I�֟��D�/a |�!���l
�˄'�	A#Ri�~�r>����P�D���P��x�o�Y�8w1o�������%V�7���M���kn�����b��cAG���ܔb*�4�L��3�0<��ln�*֨H6�_�����7&�T��{��L�T�Ɇ%���P�h�)�	�͠iB�f#]:#m���H �_E1�Mt���橻;t��
��Q2Y�ja��A� �n�zߚp�;����R�ܑ�oz�����G{wʳ66�2�f�'��(��'ؼr�"����/=<h���.)�8@�����"js���+�r"Fd���tq���E�9y��� W�0(���r]n'����v �ģ�����y]�T�7f	�q%e�wpo8��D�QR�c�:�� ��t�}}��lG��`�����@��p%�h���a�L�����X��a�1Y�=8<�sd� ��s�r1��0�W�
�AA����(!��i�ί���"C`�a�O��ōݑ/"�>�M!����;8(��ka�P����%�'�}��&��u������:izVӓM�+/scl�w�ϻPq\Hnc֋[=�a�<.�"c���  �0�_4�7|�{dv�����pvKo �T��|<���ݿǅ��1T�s��`�著C�q�u�=��Jr엣.�uH}K�8"��֪vv3�wM�X�R��>j�|���@�<�
��>��8�yDy�hyd�B�>�
��X�ޣ�ٲ.:a�#j�\�Hwg���oO:n;�i�`���O{s��)#��0{��'.g������<���{>&t%_E᦮�]�}��#�N��o��	�ԕ��|dbՔ�6&�+j�qccل�Q��cF���6����Z���ɣ���?X��k�e��g��VK>�ZAK��5�oI�VGME�a����ݕN���>����J��C������E�?-�E����� �RS����RN�p|L��r~��w2�d� 8xu����8*Xs�fX�U�Z
J�����6��Ҕ�Y���p����/���c/@5��X��e=�"n� �y'qA�OP�U@-
�xQ���pP�e�>�dЊH����<F�֬��$o�����:*������e��%��Qc4�G2���d���?�M�<�öp��4��I�-�UY��8���Ǒ�ǽ�q;Q�Ƥ�'V��w��=b*�U���M�k��g�9�����$�\��{���#F�ہ�e���9��9|2��e�
�/<W�R�pm�*=nh�A�a����@�K�����Ap{�-���ួ	�Q���bM �N/�R��+������Ctg�I-���b���A6^�3�c]��O_��Љ]���@�<�t۝4�c������<i�~i����8+H#Ҟ����Gt;���y.$�Q�sӸ�];f媴7+����T���YŅi����pD�B�E�6��L|�(�c��N큍�L���Q�u�'C��y�8Uw�J�!����&=�|��ݍ��)��"Fcj:�bW�u��x7�ӥ�2�f�S�f�S����JW�+ Qh�L�=��@,j�9���r�33���C=��4-���B�5�);4�KD
��-jվ$�� W��}*`S�6���)�O�\�=T�~ 㬰��B_�j]�It�I���ݜ�F����mD��>�Z�{�B�a�5�ʆ��uc#r%�N�_8�E�aE@!5���v^���-�s׍�g�ʫ����v��S��R�T�4���>#mL��3���2BuDU�1�mkn��O�igJF�Õ	�H��/>��F�3��'�9.I/|q{=�%\��;ʗ�����!*%K���o ��`fv�+�.rB$Xd5��
[�4C�z��hj2yb#,=�,��O�ScS���MT#�~(ˆZS;�u�}͚X\T��N��$�#�7��G��uj��Z�W-E%��״F�����gi�b=�+Kg�αgS�a��w���+BD>����M��b0F8`��Z.��Rϝ�?yw�����>�B�VH��v*d��ܕű�>!��n=���0:�E��:9����Z/.0�/��v�K�2X�1u�
_�ư��|�|;��鵜Ќ�pAd����%����*��P��^g{SF���=:�V ��"Z�ާm�E&��A�V�&��'v6?���ɳo� ��0�P ��) W%�1� ēM�M��Ht�%�9i�
�K�`?GGw�~��燀 #�r1�5f$A�� �Vɽ�`V�����HM��[a$*蟍�e�S:NF-We.�\˅g&o7�=/��:��d������2�n�d��GM7��˚�i�|Lչ����:����t��ԣ=�!3~��K�h��%��"Ěq�q�Y�$v9wZ�wP�Qal�e(/m����f5㈋I�u��C$���$�A��;��nֺ�?�`�Ӯ(r�7h���3�~��x���~Q�m'��KXõ���x"��?4���{����ӛ�����	�[+��Q�n�SR��wXά�����4���Ɗ3#P�H&Y󹊟��jw�c&��p�F�>�f��l�y�� �ڡj�1��ۻVd�$G(*
�D����	(?����j��:'��5y�C����z��f�d�?����.�)*#����{=$$�o:����RJm�}������e��7/e�
ׇ��F��ػ$M���@�JL��ܹ�'Y��%��(��爛A�������Ɏ'<@�S='*�g��9���5w�<ǀ�Z�ݝ�@�����-�1*���;�2T�i��A�o��6��?�QK7����P÷��_];��\��\A��_�����<Ԯi[o�����%�"̔l��󗷗����G��'��8��]�i��|����e�U���h]@�Dݫ�y�q��ۋL4�b��p��0%�gu���N	>y%ݿގg8t�r��?�6�A�^��F��+eL�Ǒ�J��3��I�?�VPT6��n�w+'O�`1�O꣭�d�W+����{��ob��1=s�!�<�I	���xk�o�}V�Z�Fs\��~{�C��ߦ�
�>���@"@�_Z�h:����?������Gaf4�Ɋ`\� ��|�t�{�Ͼ��2�{�R���&����o��"��z��X���ۦ��Z�=e�QGK��g�����)4�U[�z��D�,��@�9��Ltq7<'�j�]�=�;A�ٟT���:�x=_�nԂ����� +�&��Hgp-���Ƚz�A*���c(�h��C���ͿV]�˘�����=��-�_�a��_���xd�3���2��#3��-��Ѕ���d|��&� �#йcP�V��!2��+Vt�|h���P�}���7�4�b�.���4ݯ1n��ff��+��t���4�+�*@]�r	 g��k��oJ���E��s;K޳�<�h'��MP�L��H˱�= ��R��>�n�?jv�����Q�-e.�v ǡ�m�UkNj��
չuL�]��R*�����f`_��r_�-^�<>!Ɓh���Pm
=	j����`)�s�J&�ϲ;/�0.�Z��`S�Q�<Q݋����y?En��g�}�[�oj $��FJ��	τ]Hph������"p5A����]�~Npd���=�
J�:�RՔ�G��� #���Q/5��{��EN�6�̫x�^�f�W��V��L�v�$P��iR���E�Iu�N��?���I	dZ4n� �{�.��4DH�6�`��QXu�>���fZљ��#��(Bĳ�- X2�-}�b��ӎ��R��cl�e�a-g�G��e��k9Z�MFd���G�>�B��rW�~@��̼q���O�xn�osg#L���ad���5���6���|Ҭv�T�HgP����,�$nb�V.V��{��m*��ڧ����p���y��X�Ә��w�V�yِ�CE:��kg��@"/4�����b��tHN��Y�,�����_��uVL`P�y��?rE��;��U0 �:�'�E�sDt@ڇ�X{�|��Zi�k��co���K��
��/<~��L��vIݡ(!���͈Vܶ=(�KA�|�'�`�j#�� xzu+���76>��&��58�9�7;6�ZV���]�2�m��c.�B���&��]��伵T|b����]�Y}�������<v���7��|&5b����bm�P��{9&ԃr汓W׏�!�8Lu2u��-�#;B����5٥�@��$��hl�� �'@��^]´��협37*x���AK�.S.ܖ����*v��\8N/f3E��m�z|�o��A���њ��n�Pޔ�:?nV�����D��њ�c�{_s��9��}N�����U�	E��Ʒ����������MRj�0+k��uj'݀��?�˯0��Th`�e�H���E���;k�[/=���*�3��i�-IҨ)pC"c�dᚘY�1R�<l[4Ve�1�����A/���M����m�\&D��}�r�Zh�I@���sL�"ĵ55t�� }���v��1lk]0ւ�妾jqс����u�0���� �`������-߈��p&9냣��hӛf�D��[���ѩ*��枋�fF�.�����g
����9��s�Z�ו"�Q���+�����cF��L�&�p�M�aF��`l����}~4�P�z��JG���)��k�e�UfFh|1�Z���!x(�L�/�<؞ݦ����c|�^��oϛo��#O��_h5Y\�g��R�����bP����t_�b��~	&/:�~�\b q�.��飢��gv����t�5n]B����t�m#� �TV,����0���_�UNĦK	���x�ǥ$ �xXebĸXwfU_@�u�(��YW�')�;jO\2�t���V�5�έㅗ�#����'����	I��q*�Ɂ�.�=�/�d\�׊�J[_ ��F��S�'�F��p?23n�bm)�x:�\���o+{]��"0�I�?$�LLc:T�I$�#@��0��Ec��&�0Y��Bh��x�ώ'`��x�)	�u�R�`�1(��-{z�l�wڲ�mG�{����4�K�o��7�<)hEc�qs�������m�}�~�[�N����2bX2��1� r�m�3�e�D����L�~�0��&��tzJ�~'�q�VX$�`N܊�x?�� d�x\�;^� �r��/��l������/�d�}(�>D�R�d-��$�q���D��2�e�S��-#�/�(��ߡ\���a;m��y���L�[҈V�m��5l���"���M�@e<��D��fV�š�v�m���h���H�5?�`��5b����d��"]�G����V�?"nq5Y�	�m�,vX#D�����Ye��_v�e���6�"��>���-�1��;~Gf�JRǽ:g��{�xjJ�/��ce�Q�lk�����JY)��n�ŗy	��[� �^!۪����,��ľ�{2��p�O����uVD��n����1�DXѥ4<TG4
��G�ۓieE����h1�f�	�g�˰ɹ�q�ω���^ސ]L����~�����㻎��`ܾ)�����Hȧ1��S�#;��W�_I_�[�-��x�$�B���:�CĜǝ���	�B;�{�ՙ��~��1dI��-L�ܜGp�q�&Uu�������xe@��J?��(VQ�5���<��mZ���U�*��*��Q F/P�Bj���N���2�˂�E��ۆ���\���we��D�7R@3cۧ�r�;���$����T�O���G��ZYb�)[�SP�{bK���[J��t���=�:&��]�������1Dy=�"r�%`�'-���o�C�r!x�y=������8c�e���^!
{��2=���� 斐$`�ZnW�{��uUֵhT��!���QDA����_[h�bO�q�����]2{���m�=�Y�<�����D�{�iTء����Q1�!Ɣ����ג�R�A��J�,Y.7�"�����8�������[�✨�ܷ�	N8.r4��=?ѧ	�U|������L���+/�RK�;�_�-���|MT="+uiT/�ɖꏳ�hF��K��GU������O�?��UY����A� p��qg��ͷ[�"���3�a���j��޼Cz�����-�H�) D��;`�{t��U��h'o�g��H���XB�9c���96���#�Ney[����� K��E�"�7�F�gSlg��nٛ(�m���:�������+������l��$G�H@������f!��������~�"������"r�l��M�Q�/K{�;�~�{`��3�� ܭ��?Y+{�tX�ٰOK]�mO�b(�|d��yCG2���%��u���3�9+B�mv@����KT�����k[�������=��2zf jUx��"�ؖ�{A�o\�ਃb��<z��PY��[��]n��8��yW���c7CkUQC�݋|�@HA( �˲oJݤ;�<ǖ3_s/� &��$TڸL�PO����`l>�]�2�
�,º�U��%#���\�a�<���/���,�@e��-k0C�O1�
_�3�1��=/�m3<�VZ�"jbU'��w�d��'�he6m�'��*��A��<�X�˄��
�X����/�p�<0��5��`֯�уƶ�{B-�j�^��AI�Q1	�� &4]� ��{J��|��t�4���{@�@�I�n����	dx�z���2�bC����\���~*!�4`\�paR���8h�$e�7�_g���E7Si9-{vZ�a����X���-椐_@���Fw��JG�x���\y��^$յ�t'w�Do��Ӣ~��p�~?b���B���T�q�<'��7�V`�H\+��^� ���������*��;�`�{r�����%˥��E����<��f����������<�D�;L�R��u/nd(�שfy�BȠ!�����=WI?�^��������Q̓�Q�z:DT��O�`����L� �%-4�}-���&���۾)���u?q&�N�}�+'��S������_��,*�u��G��IZ�o���s��u��NG�҄��^E�?�n��%�����t`�n�6'/P�ﭫ��M���$P�(hJ��ap��M{4���Mh�̠+(�n��
�@����w2@���dx�C����S�՞��X\{��r���8$�g�e�[Y'G��� 4��3�!�p�i`��,�����p���=���Fg�&;G�/���mQ�-����Z���FI�UJ��[�X|aw��q���e�`���R.|�+UZ�.�PD�2{���G�u��g��W�Lo/�]�f?.��_�\�B��T��a����fN*�+7d�d{e�0$�'�v�̃�x_�s8���}z�A����"O��Tf��0A����zG��>����-4S�5S�#ne@v~z�N���0��M���	�+]sz�\�ж�/��P�0&�&��� �Q��

4�+{�3���xX@�{p����( km��١�ۂ �k97ֶۙ�ń�I\	���6�0�RX�T��|��*3^�+
5��#z)�p��QX��!�5�|�-_�-����b*@k�R/�.��!a�A�wm�Y�;�в_-�#�Gu�^����S|��m��f��h_������ǅ+�j~1������C�V��JĪ�<K��r�m�{$�X�.�b��f@�Q���E�������mԿ�?��b��$����uu�� ��oc�j^�rdo4������
R��N�Ѱ���A�;x���O���,�ފ{O�����>�g��,4�����eG	��e/ ��p������cl`S��ܶ��]��E��`�"@�����?���q����� U��Rz:#���@@d�.�TJ�:<tó,�{��)����lA�*�@��Zc�xx-Z�X �i�A2�tǞTA�'�n} N��%�����A��N�L�RƓ�'�.�_?yL?��,��sw�I��0t��E�hԉ�z���+��~�X�Z�`Ff'��wj�f�Zۺ���]�2�|��O-c�tC�	�ԫR�<x&9���� fQ��G�Z�Z���Ӆ��F��>��&�H���&�ӟ�yIZ:��$q��)�`��"1mz�ą����jW/���
٪��`�o��q��p�[c4OA�D�Fֺ����[\�og|������hc�Mhߎa֢�AĈ͸F�1���x��b��0��,�'��Z�]��0�$����^Ȟ�$kKPs�_F:�-��>��ՕTɽ���{)����C���Yg{ ���j�˰��%���)��z3PSM��; 2=�S�	�7��V(Џ�1�'ؖp�}����� �VNfv�H�z��|�55�F�5^h2t�!���O葘���+�x'�=���y�o0p�D��N�A���4����TM�<BB��f�Jt��v8�'H1�˾r5�>�7]���e�r�c�<y�,qJ�KC>(���!x��HX�A+�1�+����J�fhg&5�*�")߈>TF�'x,	��%q��?2W�E���O���ѽfj���+�f.g��h�Th�ָ	ݬfY���;u��pY�@�i C�!зq$����&+�@��> �ܛ���F��� �Z�I�zU����e�lK�YN]���I����S�\�p��w��푦o�M2ם{Uԯ�4�s�]�~j����ۊ�9�gKb!u+�fn����󃄥�EbPK2bz���4}^�q;s@F�8
�I�-
��r_��Ul�PŽ>a�Y1q;E��u/�y4Q�;��P�oM�E};N�!�mON3'e�$jRG�����Κ�[(�
�e0�\���tys fx�� ������%��&J��}������zs�C�fQi=S���"I9tS�t�-��G�;��xqD�d_[ꡔ5k�&� ΂�u�R3����M2���Xf� 9
Et�
���cPg����7������F���s�(����Lm�˚�e]N����N��`��j?�&���p����R�z#��b��k;������%M<���Y��R��W�JX��}����f�'#��m+��Ӱ�
{�%�nH\X��
��%�B��� '�x��þ��2�&\�����,���d�`Ǖ�s���;N�&�G����Хf��ݒ���k�hJ)�����r/�Y��3:�L.0�����S�-��*Ԍ���Q��x�H�p���b�*-~���9B�6�"H�.R�Y|p��ǡO^��G)?�V@��-AC�r|T��zB��?ilB�pw/1Ғ�����s)	��������C�6 d|������óp�e����e���<�����L�A@��Ĵ3�oN��Ltbu[ټD��űs�f���On|g����6��^��R0ž��k����rd���+Dv�R���%�����Ae}�8�?|��>Ob��8e�\���R���CX�zs紘��m���ؖ�N?���Ӓ�����������ų g
�'�k�\��X��(t�l�s�T����v�i�u��K~�^~Lb��Ŋ����f��I�e��VҺoF�\�7Y����
:<�3ÃF�	F���%�ѧ[!�]�9'o.6V��v�-u���e�8���h�����e�B�ܼ:����{=�_!΍���M������f�:/C�]�Q�Nc�Fj{��z��b�����L�(���|����A[9�kSa�|���?�0�L�v�'ֶ�,&*�]�UB�pS={�u��gh��k��)[�a?�Q'��S�IQ��$9��}_�(cn1G_�WBF��bH�B§���ϜQ~h���H׃�5+����Ԯ��tu�6Hb����Hƚ�]i�Ѣz����4��<\ag��6�GNڑ�g��pMg�`�9��?uŲ���� ��*t�5#��ru؜ɤ���yl��5o��TY�	�A�_�ۗ0U�T�i�Qc��kJ3���X��G����
Q��$���Iq�������]a��~��D~cJ�%���a�I>�5�I1��PD
���}����+�c��L���Q�{�\t/��Ȃ_���w/���[=c��D��L�uI9��e��%��c([,���y��vk��iP��'lS�@��o5x�� �R_����	O�#�0u�����5_���L���1�Z'
}l��6�e	򚵐��nͳ��iC��X��[R���d.��z"��N��:���_�4L֟�覫�C?��j�r��2n�3i�j����'��H	z��TQ[��h%J�(C�Zf�<�IB���|}S�Kb������ܞ�	n�C�Y��ȆSlm��.9���b�~$����zI*����zc��H��̮φ}�)#�<���D��4w��؛�m�$>kFi����#�@6oD�'1�g�����MX{V�M����ov#?q�C��n���{Js`�b�7u"h,�����A�	c�Z!v��^nhk��[^뻹�W_�)�m�hn�sd��,�
�ܞ���:r���#�ڷ�Ɇ�5��@� Єb�qO��O�U��S��r��k���F�=_�?ľ��λEc�b���C���a���'. ���T�!��Bo�p���OY���5v���(BDI����HdD��<�K�^�D�,��Zs#�֣@�e��*S�;��4x��^L���o�+vݪ4<����9o�a�59z�� �bu��3@�q��t�̯�7<�^��3~+K:+9��I����\0.� �Xb?^g_���z���K�S��z����ic���)�9��MshA�YޢJ/��5�VY$�`u��g�@ (t
L�PL����P�(��-7��}2��05[F/�{]�����EϷ[������4�U1���q�P���YGU�O�~�ȓV4����%���mMZ���|[C[݋�&���³�^	�7��"��Me��V�,� ��/J�b�A��S$a���/.�}��z��q�p٩�4k���N���t$�Ғ^w��+��;/�'�V*eL>@*%��T�9M�����D�XGf\�k7�u'�ɚ�ͼ�Pg�qޜ��E
�gz��k��O;���T7�t�e��K�إ���e��}�e�]Sg@�c�s��)��Iˈ*�m�`)b�ܶ��T ��I��я���E�=|�ڨ�/$�\��QO�J�S�0�.������n�4kΐ�:u�Zs3�c
9Wn�e멐�Y�w���·��c���O |$p������
b�ȼ=Pnf�CCP�cBޏ)f�����8n�*��mTR������8��-B�FX��%-ѫ��� ���I�
�Z�����0�r��ߨ����Y��Q�Z�ck��s���J�eC��><(�H�� #2����RV����p�����	�����5���O?Z5�{�S�b�]�1a!�a����/��n�33�7�3�0,GhC�	½�F�̦Ʃ�]�+W�'�(�pG�l!�nXƓ{��my���ʄܳ���nn^c"�Ɇ�40�5��y�3;8�Zb��%8)nk-S������f�]�P�� U�0�C�hݾ�p��7R���5f�Ʒ7��Ul�������Rn{aT�4J��b��x
�T�T&TrtK��ޛ��FP�\Y�iu�%np�mK��<���t�І�����_�՟��5��C�#q(��>k�w�H)C��C�'�6b��K�	�ۗ[�r����
��~����b��#@&�K�欅˧�H~/I����׿��v�^����z�Wy����3F�gv?[ݨ����p�t.��i���_`��U��9tz�����2<p�THop�CI��b7s��OUȑyAt�`�	����K6� 8�F���o.M1���pN�Ŭ�&x6|���{!Zgz���?���ײ���M�F�al��o�/>!�(�#���=W?�t��JW�)��@��Lf��}��s$>����������Q���+������
g���|&썓CKA�-�P�q���Q#�=�w��~�����2^ ��˪]>�X�z��$�]0��L\��ؿ�����8�٭�G�y�h�^�]���N#�~�w&�j,◡=�ܚ�g��'�Bx�f�Z
��LC^��?Qr�vf�3�h2�h�l�[�	�C�ew̦``]���OGD�W->�Ձ��#-eaQ)4�G�0ǘ�&g�$����n����I�o�KP;��#�3�_)~[�٨!���gU@F�l��:{M=�*B7dc�`�Sb�A��*���_�҂���z�ؑ_Z{��[
A��c�b&Փ<�Z��=ԡh`|��$�.��`\9�(��lm�U\�Y�R�<X�Sv��Y��<H�h)���܌�.�Y2x�"�7�m��ǰ��4��i��j�.̬0� �e��Y݋�p�'8�z��ss�ۆk�^ez���H^���7����&��Z=���� 1=��a5��s����ϙ���+'l��&v� V�j��|��BW���z���dΑI�36'��֧��0��W�6b#�8=e�%2Q�U���S��Б*SO��2�t�?�|rm��L�ǳ�;!Z{�l�MOxn�p�˷���~3�}�G�S uQ�5��m�f�����g��~�!��yur�mT��c�,#�vN�\*��5%Z�(���p�<a��~D��z �\��r^��L�~z�>��b�KKE��	��dYCQFk���^���_zg�B�r1��X�U�Ƶ�B���������W��Q�S$��W��0�`�C�`czo53��]���L��*�T���b�ظ��iWD�j�B�d?+5�S�(]�*��T�MY(�u��V��p"�l��ɋW���jc�`>���|�_ ����N�(��!o����æO`soo�8Զ_����q�?�x(���.���Eq��H�]�",��r�FFC;(�{#Ǹ�>��P&�զҝT0�QG��F��4�f���HĽd���R4�%G~�7��a#�$�Xˌ8�B9��W���2k���Ͽ��8j<�0a�Vm�ס,ᰩg��%��z[w껪Xi�+!Ƶ�oXķ�$�T����D�{HW����xR�O�I/��5��X��K�,� �b3HW�Tp�8t��~���CuRg�քq[o��!��jU�ON�{���vD��,?�V��χIW�1}9�����$)�(����'�_g�|�C��;���W�>kG�+e/��c#*�݅b���N��f�2�@� a��+uƑ�������J9��.1�ߟ1�0i�#� �M mq��&֕��0�"%��ľ�:`�vܷGM��q�=���Ԛ!�[���'!�3��h@������٭,����On����3B˩C=�}Ec��?�*/�@�����&���^�iiD�=].C2�P����q�{��"bP�5���K��Ȣ9�uʴf+�\��%x-�;2����\˥Ȗ�k��o�]�"=@��w�8����Y�v��:�W����/.B#��Ԛ�&��)���=�i��jy��^�
F��5WHǣo�&���E?-^�}I�&���ߖA�Y�\{�J5
�o=��9�n�tx�BB�G���P�O��
�l|���>�	�^�>A��k�8a|���0�rUI��������3���YQ�x�w�H{��Q1F��(�����6bpI>.Ж#2m�
J�g��2�W5~�+�	K�\f��#��<N��2	7��kā,^%�O)	x������~�7�'q ѥB�<WO�HE]�y]v?�"�Tl�t��
�T'c�v��@�U���QY� ��)</˪S��y��6�H�Q]mIs�k�"� ��H�̀��!��~����������P�"6D�Hxk���\��XK�	��M&��5)�y�Z��X�uƙ.��'���ߑ�����Iml�f{j���F	����ؐ��G����:|�Q��۟km,v>���x#e+Ì��C��ӊ�YZ���?A�~ҩ6jL��=�;���Ë�^����o������N��Sy��JW!���$/V��ގ!v5+{�>m����1�K�h3+��k\�D�8��*`K_�+�]I3��讆	!��d��x���Ja��9V��H�E�+̯U�r>���d�r��>�/�����}�>�Lʄg���Yd_���� Yk�*Z�u
9=|T�`��%����.�V|3��"���P�n�s�^�a��0�aN<����X��cEȀj���F��Ԓ5�GJև��3�^{�]�p)�@�!�)H�v���+LK��_|���ޝ�t��H7ٰ�"C n��>����Z�?�˄��^��܈����,f���j�%�򏰀&bcr8��^y:�ͻ9��u ��CZ>3|��z�ؖ�g�|Ĳ�c9M�@�z�҆QqL�z�M2Ԁ�'� �
�U=7}�~/3��{�O��o�x��؟�;���0	T೘#�_du�2�����eĲ����bQ�:"���^���l4}�,}Xn5�jV�ȓ�����k��v�@��|����3�����X�'o���V-�:	��.���h(�ݚN��Q��Jb�j�ư5�h��(`a��\b����a�t�+��m�����9��2�x�*eZZ�E:�E��ςDv�t�j��,��|��}�)�G
�#tcj���W�.ũ�+��h������7��Y�3�%",�v�}o?�`��P����!L$mdb{ap�K����}���4
a?���E![�L���;���ym��5�! ��TqM�m
���*:��l)��ɡ��t�ݯ<��3~d�1k��d�ΨR�9�I� ���RJv�<@S�p+��25���Ϭ���c!8�?�P�;��o6�mV�P\*�������$',!*�z���$�C��Zɞ�f���G�a�����:��
��B�+�c��Q�(AXD�r/�GFoov��`�1^Eq�10�8ٿY���|�0�Ɖ$ɿ�Dh:$ץ ��Kx:R�TnF�ҡ�'?�_!i�`���|%V��̣V���Id]��Ʋ�cw����>��)����2�$�A!�D�@�K/.b}|}�)��t)��^�xaDc!�JR�LJ�4��9����� ����ǘ�q�U�+'��J��]1;]*���M�]9-E���G�`��j��8�-=�T����K@�)����/8���KdN��?56`l8-���o��n�sb�T��v�H�K���G�eSKi�-�O������xS	#���~�0=���3D��$�p�?y�A��y����0����Ed�}��#-2����Ha,[-`z{S[��w��|VM�zǱ�T�����t��&�>+�^�w����^x�~�ִO���ŇX[aa
2�b2�iI+���Ԇ�YK��]�פS߬U�����3���%S'��b=�r-�/��h��Z;#�)\�
�j����r[j=�z�Z�q��%�%y}�����.vދ�{T!t\���!�"����vC��IY���&��c�h8K�(�����Si=�2��B<G�9W׊OU�h疲p_XUJ�LA�+�1�o��Ѻ&���3�N���.L��\־/���Z*rMҍ��K���*U��b�zA[&��&� N���.�)���d#ǋ�Z�hBR���U���c@��o���=h,��jD#�P��SE�z]�G:�;Q!#s�G u�;M�
���tlZ�:�~�Y,zs�
ػJ7�f����1|Kr0��un���#�'��B�B[�,k �zٚ�9���OEU}q��ދ����W�,����%h���v��Yt<������]*����P��j@ڷ�(��$7|�� �٤o��>�ܦ ��':�<�Б"����f�����E�1-SO#fr����d�X�f�m{K��P��W�+�3rBx�����b]b���)��e[������[��g=��Evnx�U�\\��SLe��i�qA(^V"�Km���pp�־Aۊ��f��%XQ�}@��ob�{L�o�h����N/_�·�`��0;��h_P�2���>��|�O�;���9d�~�W�,,-.��̼��E�*0X0��e�AH��h��.eKF�c��������6�Nqv�, K�u	)��E��|]��t�-�����Ir�OS��~ ���!����k��ש;�DQ*'��]���<�t��9���;L7��ܻ+�	zU^�ĥrބL\X����mw'*Q}���'Z՞b��4���y�mKc����	4���o��/Ws������0'���禛pkI����0;��Fÿ���QAl�ne�+����,��fR�N  ��%"�]VL_L�׍$%Ѵ9�4�.��?���&�QxÞ�a���d5�3�٦�{��MZ�T��Q���bB6~q~��>�ә��!��"!Ѹ���m~AQJ8�����6smz��r�|��NL��������V�`���$Xaq}�G���M�P�Rnz`�^%l���ьi�N��Bg0���e!mu).)��Q!�� �:�����q��~ҕ��5���{S���-.����K�~�����Ǹgb�l[^�%GK�Ǌ8�A�!պ�������CcI�����թl!B�U2��`q��quZZ��2`</� &WR�e�]���r�7�tSt�I�*.�c��A�+����0J��ξ
0�^��n�g��ĕ��:�!�f֞�yf<5�_�7n���A�2Կo��:�9�"� `�p�J�3�ɡt�%�H-�Z��`h$�e��h Ni���pX%�	q�E{�ؠـv3�N/HdY��)g��̖ɬg�\T�6��C\���i��h��5��mJ&6��{_�p	�T鯍nB��S���xWS'��+�g�'�^��v!�VkyPƸ��:/�;��W�ab�@�OR(ǀ\��}�=�i/�
oՑ���&��m�>�Bn^H^�/� a��Pn"�B�#�²F� �n�z���+Få5�΋��N�p�U�k����SEs��r�Fti*��@;�t�b
�}ۧMS�Z�	s��bc'L��WK�
�ԍ/��vEЌ�����̐��4�;}1��}p��A�Y�H�(I񸘡&�c�8H��洔X�%E1�n���$[�+{�J��2���U��TX�ʖp��0�7���A,t�l�1��@4\���-���q�\=���� Aj���2��w'R�rټ悁��ۘˆ��W]a�.y9O���(&В�� ���P��D���tN <`:�t�${�a�Pi�Ǉ]�I�7�"_[�´���3m3���y�t�p��9~��
1�'�+����XePR'�e���聯�>�#����+s�1!=6�������:+E�#��M$D�ޘ����P��䤔�,��!�E�Z��n]��=����덞��uQN:$u|+��$��ϦXɾQ7�L��مW?�P9�,ԙ�MM� B ���[s��v��eێ����{*G�e(��@��t�c
8̦jWd`<=�Y��1d,�
�3�4����T�Z�6���t�Z���/)�<~08��kbC'ǚ
��Ut�ܓ��'�f�
������M�Q��L�b���"�BG�u�~�GY�@\�����bd�w����L��������}R���EW$��$�33�IP�2�NN�}Y���Q3?�"���4z�3������}l�ܣ��+�I`H ��R�XGS^7�l��.L�Ъ��TK��\N>��eʃ�րm�#
����s�<[��R�@1�Z���Y�Z���#�X�x���W�0J�I�ItT��^��u����b��ƅz�$�H^��l8�:X�=� V:��A�����S���)·@���*2%�GG��MW�h\��^4ʍ����@�#�BX&6��n�F;_H��Y\�RJz+�����.4=�ʦw4O��M�u�?�M��c�Y��H���ħ��oY�s`��[��#p%�)��:��O�Dw�
���!��e"��W�8���3(�F�͡A��C��U�?��$aXO��.?��NaJŮ�>�	j�$�돘e`J�Bf��qF\�������/(Jϖve���G�����=p^�v]�l@�ʤ�y4ڹ����E�\���(��aƮ,������]���ajP�� Jq��n��f�A:+�vFH�}p�$�"���%����i�H��.�|��8u���I�]M�V���x���1��K�9���3W]VDQ�j�dD�V.�/,����1�B]��vw���'$}��j���46{�-:�g5�4��J*X�V��8�cts�/�z�+`|L<t��lC�֤Y�ʠ�qIA�#�n�G����)��G�D*��t��9��#q�C/0��
��'��#>e�z	(��Ύѷ��̹��}���eتl6!�<���A��O��/������Uf��N{�>c�p'c���:�����7���^X^���YY�����.i���O޳@@�8^������WH����W|\���5�S�L3�(wz��O�[�?�#�M�>�	�mR`������:�73�4C����{o
(@g'��ݏj=�&�D��7j|�R�_0�\��G%�!���H�0��Yh���=����]��O���S�o�l!u)��n�8é��з��q m��m��°�Ĵ��aq��_�F��M̓<��-<�ѧ�~l��ƪh{���9��W�O[���/���{@�ה���I���zr����#�RY��%�ae�i���M�x�����G�I�@tN���̝���h�O	�T�u�����'�S䑫a	^U���kKh�	�a;���Ԡ.E����A{�����~.Ypi��'���:��Z�����=��g!#��u�ً�ԫi�g v�����#-S7[��.=���pa)-���Ǩ9Ao�P��=�L�$g���X�g����I�����O����n�s���FbD=[]�I���/�0[ ��(�~~!&J[�9�(L�k@��2pG`B$�T��i��@����ya��s:�*Ne��S[;k�
��ܵ�N{���	�.��ƀ���@�~HB2�V�OY��HB<G'�5�<\��O�,���H�xuB#l�Y2x,vFJf��&�NonF��sn�p�?�ΣKn~�W���&]������h�h�z�q��d�2�\�Xd��Z3V�;9`�!��ʽYB�Q�~���B�/�(����z��'�[�d���坚�K�w-$�37��Ք�a�`�8f���,|/'1�,��\q��!�>�&	�|U���&��n:� ](W�({������
]�&T��'���Ciz�Lbe"L[��f����<!��ٚu��q��L�Cr�L�?�$��
���I�����l��}Ăj!�%U��'"�%�M��[���;�^VkA�<6���'�a��Y�Y����{�^+�5S1���=OM��8�o��^�����������Ү����Q<�f�����1n��ֿNp��=�B�ԯ��+�0@�N���jo�Ű� յS?6��9�H :-�< )k�U�����sǴ�a-X��q�>뒏��2d�\4h�~�������\%�^Z<�?��qN����|[x�.uS]�	�{M>]�'�U�?����K��ҿ�I���?�3��t����7�d��
sQ�ň،S:hWʑ��h��vA�$��2�=}�����p�=��z��xߋ�z#�A�HGz�&J��0o�F�
�t#p�G��._ʎC�N�y�)ݩ\��AHzDI�Mc:M�d�52дA���/b��
@�}��� v�j���TGuN\=��\���o�b��N�XMc
�����G�w�̹g콺�s}�sl+!t���KȚ�f1:��ɶk"���vμ,���髲��8�
3�5-���>e�<��Ш˳�
����BS���y�}��K�� U�����Hn�{DoZu���D"�i�oFF��3�D0�O�C���(�����+#�-�j]�]�Z+����	�=�I�A����}��z�ѼF̈+R�ԇWo�D��a��M�p�'x��a�f�����ld�R�5�iw�s)�9N[Smn��)��	���+���.�~h�,L����=����A��Ω��]�N�p��5�X������V�A�w�����:�E0�ۓ�9Z���x�ݱ�p;�SU�#4�Fi��|�OS�#��ݪ�����1��m=\�Q��B'����v+	�'�T/��U�o�U4�&w7���>��̐:�_n\>22�GN�}}��yІ51��3EN� �`Vg/ɐ�Z��rͮX�?�M��^C�`?���x[څ:��4��	���پ���|Xl�|��ұ����5Qq�^�@Uڰu`�_4)��t��ҸN�&�h�7;ů�+V��A^p���d�[��rd�j��d
�X��۞���Ǻ����-[�n�K����v�NJ���x��@z��碍!���D�S[��� �ȇ�1�џ�_�PJ���5��7?�|Cٺ-�P
 .��1՛��;�nw `Y���"�����_C_�Q19б31D��%���}ܮ���K"�R�\f� )eh���DAd�	��BU�f��}�Qw۴G���?�'Au��|?�E��D!~�F?
����'z~�\E*kA��9��M�8��$�s����|8+��G�M*��/с��u#R��c[U@5nPv�|D�Z��=*i���.3��)?�%�o�L3�c
��W�T��m�F2p�D x�ht�Z)����O�B�t�� ��G��vp�m��r�r��iؐB�e[��ހ�mCe�|�7������Ls�w�@��v;z#�Z«6�{Z����#Mj�cԾU�6���Qf6��E�k6K�����$Ӯ���"	ܙ�{Qo��(�CU�w��ӓ/�bF*`�wyC*������[�U!j�97ǀ	[���ǌV�^:��I�L��4\,�s��p�r�����O�&R���qc�C�ݛ�	���U�d��'��h���Vmɶ���[n�+6I}Kr���`���.\���`jN�b���n�빼J�{��^t��w�v!��
�b!>S6�7��[��n�2���R��xHwV����}#����O1j�E\�`d؋G�p�R���U�Y��.�{��^�=7�ｧ��X�hJ j��Aas�BYD|>a��LE(z0�×�7�	�fK8@޵q?��3�M<��E�a!��\�� Ğ��-b{g[(�%p��}i���Z��Dr���K�[�9�O��
��/>� �1>9�m���U�Ŷ����N�6x�X.s���ص����_�d�k��d}�}�tC����YKe��'7WF��%��T29�nD�g��Y����))�S3�����i��w?�iX���L��(?+�_�h�8ѽ����<AL���	joD�L21�7��?��cx7���S���<��8ed�����̗�����[
�Q��9��/�
z��mԼ-C�e���~mÉ����Y��V ���d?W +f�(N�$�K�5����$���
�6��~o��Aag���|���f��e۫X��7�=��f��(�\�x�T�����yKt�Y3�<��0��� cG��j1̈&��d�����ķ���:�NC��Ě�K�%ˆ���a�x� y��{��;�C]���*�%�z.�v�Լ��;���g#���bd��$~�@�6S������W��g�(t�k�8�]���10���@��ǭ��R�#�S��㘟�Mdw��/��
�c��CO���n"+��v�_�3A���9���o��I*?���� 쒥�WR��)1���E�����-X��Q������u�q���I8f\��2z���vm�K�7"t[_P�	r#�M���q�i(��2�����R���Z?���<aѻ+pՐ�����b�L����˂���I�	ݙT�7���{�Y�܀�d/�ŨS�rA��L %�#HK3������Q��x������~��8O�LB���1�=�y��'N9��]}��9��Q�+ �6۩��"YI�å���A�i�}p}�?-E;��F-G��//p@=��������Î�f�_�7�>��ኤ��P�,w��Qc��G��Iyee�?߇�F���	-�4;��������Km��\*�Ҍ#^p2$�V���!�z^P4��s�9�-fv�	����l��iOo��o��H��?��8���j�=2ٯ�$�I[�;�o]��e�v��_ZI|�,�'�w���Rs�4�v/[6��7�H��Kc�;f��J����yĢ���G�}Ke��>z׻��O��!w4��З�Jٶsf{o�$����*��n3�˘�������ت�,˯�a��H�SeO�6��꼡󠳩�N� U\���諓��L㊪��y��<?J=��������H�2^2�	Gw+�@O���[�TI�F�'x/��4����K�J�A�sې`�#�ot����4�h�2|��6\,Pdo�nmI�3U3���U�����9���k�Z�.��]DE9�����"^����0xD�_��ɣ+]R*5~��B5L9v���S��$ ���d��_��|ә��&��[z�<̖;�c�e���*Z�^Э�`�A������ψ��+y<� �����D͂?�2�����2;D������٣W����}O���hY���k6V�"Z6a�BچG���L�0pR6�`�ٺ�ʣD�q�61���*Cl��\.۹-(S��f���AS�&i&� � ��q��@���o��j΃�m��q��]�Ϫ�~'�dJ#��are�G�����[Z�l�L
ic0�6���hd5�uu/9��i�G�����G�O�zު�w'��ڱ��%R�X��Ai��{[Z�[�ۧ�@b��*�.VX����)!���9?�4՚(�o��؀�`��l�J���q�@��<|4�����T8����[[}}��+3>F�'����ˤ���=�J�?M����Tz,��[��k�P�]�k՟�� � ������0B7l
�������g/�ͥ��Mi	,��z�{���uʰ��*t��#O��z�T�#���K��b���+`NQ�˫�>lN�Ł�T�r8� &��j���
�T pD��9/kg\W�j�̄L4�'fN�s��.�{�<�:��=��._9K+�:}�I���W�Jk�1�8~wl����/-l1�� �1ՋJ�Gdɽ�b}��1���]FW�IE8���_?L�:��v�L_��ș��7A�j�_�ԜC��=�e�}��^*Z2D:�n��tG���Oz3�����өW���.0��	���jw��sH�u��ae�p�ZW�L��G�� ��k|��s�yF�@�/cI���{��U��
TpO-Ÿ�F6�	�f`��#�1�-����,G��׽�Ԅ��)v'	 }����X�x8���W]7���ߜ�j�|ǵ�I��0�:{4*O �X����tW��)��"��w�<m,�����h����E��@��<w�>�ҥz �������;���n>e�·��68�X�y��踼~y6kV���x۴�N\�7<��~v�����y�����8�>��5�ɭ�-�\EаB@��8��rY�{�̄��lh8m��7N��e���I+%"�h�&�����1�V��Z�w�[~[����T����D�
,�m�$/� DI<͘WQoҰ ��4}ӏX����ݧ�yC]�A:uw���}f)'��<V�}WX'�08 �x׸-v`?��a�L�5�����A���oc�"XM�.�D���_��W%�8�p��b�4K7��'�/!&�6';� -�M�����G��)�p�<Y֪��/g";B*r�F���n��Nrs��!O����b�l'��S��R��8zD�C�@22�j�	���}�r�0�nv���[�EV���K��e)��N%d}oIh$�B��ϼ�[����&$>�x����Q�xd�	L�� [o�j��x�ؠ�?m�*�-�p#����XH���T�� (���F�k~i�c���5j�*���v+��\��#����+��<<�S��-0=X����֊����RE��c#���m��SVoP s�C.Oқ,�(�͢x��D����̀��� �3A�<L$��+�W6hgS�@�*�'�B��ACP�,��T,vS}�|��5^���}:R�)2�&?bO��D���X���o�ќ��܍4�Kĭ%O,w�:��h~8��da�r�Ӱ����AǹG�"�ǬjYl�f�,B$���P�h�)�2��w��B�֩o!�\�,��~��њdY����$d1ƌib�|��+'MwZ��ݛh=�Tc#�M*ԐTmh�}�<``7(>���^��=��A������5mT���p͐������p=(	PC�13,��ou��18x�1��� xΖ����y���F;�&�g"����r�F���;Z+�K��zN�@���Ġ�%�g
Y���,�ke� M�Q �3?��G�(��v�'��-� ����iV��&R��kŝe�*Wx'�|^s��p2�ɦ���<����D��0L� ��q5ۜ<�f�~��i�gh��/���R	���-��.�, ��4XS� L����-��ﱕY��N̄zu���{��SP|���F��N�8>l+�������,6�N�j�D��Y��,�����B����S2W8���Q]O�[�V_`z�p[ԍ�D��Jd�,�������`�L�|9�e�B1��)�{�u�c.�]��6��g�@MR������ض.h͈�C5�4aJ��V$M�yY)�=�h Ѩ��I�Jn,�F���!6<	����M���B��ˎ�3�ʻ���Y�;�/^�FLs�#Q!3F��P|F7.'���%��/�o�hNNOz�m����a[̞�.nzm�v8��&�J:�'?_f�m3)���nB:ew:Xc�ED�CyL"a7�@,k4�k�;���"��I�]�i=<F�|Zi����U�Ճ/�n}'N#L/zEaE��*��MBȧ�Z;�ˮ��iKY�7�H���z �֠�U�'��F���#�n��>}�	�j��@@����Y�Q�+��3�	(��x�֡Z�4;���38�Y��e" ��t��Ui ���XZ�y�\�ݏ`2b���^���� ��-$xQ������K�21�%K!R�I'�����������2|-Uu`*�|',�+SW� *,(PRX�U��)�6�w:�t�&����0o���<8���ӘS�U	K]M˫�t��d�&�;���X������UO�`�0RA�3&�[�����<��C��VO&OC�˞�Н�Rv$����Uw@�"n�K'�%9�4�R����XU,�|��k��<i��V�?���Fcj�J�UM�q�\��Q
�����Y�h�m?��S�B~ o��ֲ\,�6.�+���8=�[H�{���h�Z5uȿN�F��˕����",\~��e3t�Lm��$�#>��dxXJ�*��;ͤ��O�#$o�eҽ�Hc���V;"�f¹�P���O<'l �j�4 ��Y��,�Uu�^]g���k��Yֿ�L�š���l���Q��|!�,03��@�7	Ar9$�Ю�ÕG��/�?���7KP�+�ըh�.��k�18�>��͒Ģ�!�߲�[9�n�&����^v�nP�e��6�'d��,I2Ă����{F6���E�y�iñИ�a �,$�l��$_���j���f��k-V��[�mL�����z�؃�`9������H'Yk.�)p�c9���۬v��Rf�IV[P���{m�PKT�4R��8�
�� EQ@�*�V�z5�0l�z�R��ny��>Ha���9���2[b�m(�`�q2�#���	�9��L|T���9�������TMc13����3��W]����T杓��/t�<\�ImoU�?T'��?� �+�Ύ�
GU,߷0���f��L��Ѳ��$�;��`��:I���8M;즜�b��Ӧ��o�vk�B��G�#�PR?������F�}E�kP�����j�t���d�����-/2�:	_�@?�
q��}[_a��]�i�kU�����5�o��Eml��M��l��:���P���wZ�;#��m����ƑTs���䐻�g�RιG��_������v����T�3��Ng��ݴ�i��~��Y>��T��=@�=Ɇ�*i�;&��Ҳ� �qD��u�v:�#�blY[u��ML�0���zW9GpŘ�4��V$��j��wJC�n�r��a6?Klۮ����7���8쩸��<�[*Ԓ�A]+p�(c���A=���铮0:��#	F�(Տ~`ꨊ���A�F�N�uA��j2��`2E2�<s���!�ti:� ��)�a]kN@��/�?>2L}K���b����gT}�T��+�K�2Q�{b�ja�rUV�b�?P�
�gZ?�z ���<Q��(�?g:����eϋ�ť/�v�
��~����s*Ed�g�	��`m�%T��I�A�éC�s\�)����H_(@Ʊ��y�cB#�H\�9����܃�����U=z��'lə|���W�$�j��K�<��H��l�Pk�]��S�OCQ�����Đ��=��k���a_뗸j"G=~U�˒"т�7�b���5NJ#����n&<���)�|�n�;;��!	6���uJ%K�O��'3�a׃c��Q��}�#'+t�X�U%l,"u��f��W9$��z�*U�c��(� ��9�d�P%خ�W�,CP�y��-������?�"5�l����O�j�9�j�D�o�N�ӓ�c*�iz��oRI"ӕ�=1.�P��h��R������LMe���/��>�.�2�S�0��̓��
�R��$��j�65P	�l��5��-��S߻�%{d�xsW�P
�%  濦UVD��	[���Xw$��Uc3l��i�Ɔa�� ���CNn�Nq�Ke�|���	�.�l�P͆�^L�%�oj(oH�o-u�IНV/��(vv>���_0��'&�פ�E-n�ߋ2��y[W5:Owl���2�(I�����N=�ŋ�Z7>�����NẄ������M��ʁ��]���'ڍ��W{F"���L$��O�S� ؂D�,��>G=��MK��Y�3Zs��o��5��p&!9�0��0z>��naO�� \j�	�%�3}K�ݫ��܀o��]*������it˖��s:vuy�Y��~�3[T�6�@��g��{����i��X��b�_	U��?2=/	�qVK�S8�Y[-2W�������Fl�2��m�Wz|qa?5��t��cdC.)-�K ��9�Oe5V�"�3�vO��H,co4�o���GlYӄ)�'5qC�#cq$r�P8;�Y��B�^&��\?�H�i)�� S�gR���5J"S��?2XD\iف!��B�WV4|����;�V&�Gj18tK�C��C�GŜ��?�k�z^�>(�ԓ�i�v������
�Cz:E�������}v���)U!�hM�f,�I?/s��r�n�/�u��m��pb뙒K��ɯ���4򸴰 ����eg�:���K@�*T��ͻ��'Gԥ��L@�$�-_�y{��9�|B���cE�~4hE�(�M鲊�MD��z�d����nB��*!�s�{9͑��c��g<�d�,�MD܏�r,ʬ���֎�HB$�	X���	�̹�>]]�����g�P�rtn��=��1�.���rOBR`7n���X��_�@3<�̮	L��2��c�)m�d�<n�w��:��Iz��C�w��D��PVJ-��M�C�K?��a���>̉Cw�r�o�:�3�dr��Y�PN�#C�]7j�\�(��C󼵫	Vl�ty��h����Ũkrc*f���ҡ���L���L�[hoN�L��	�a�JvE�|槪���u�5[���I+�V&7�	]�շ �o��bue�Ԛ~$�N;�ug��ߥ�\������On�n;��()�E;1����� �b��Ճf�k/�p
IY^��n9F��'��:��Ċ�1-H2P��;��<6+��\۹ KP�mN�@����!�ug�ꡕ��W�� �5�R��<]U�`��� �ŭS
;��ːa�Z`�������$X�������^�r��c��.�?3��i�w,b��w����3��x�)�&�W�陉uY��p16X6����Bo�ݍ���O�9`i��*���~��Z�"D=� ��{��8�B{y�@�WR4�S�d��vy|`1�9	i}'h� ���BS���`?�k�� �c���F�5���� N�sj�m0��_G<�eK��ҋ!u���n)�e�J|���(K�M�צ��?�Y�*����K�C)�4�קa~�\�.��;=P�K��Ն�He<6ϔb=�h
��M�(u?%KȨ��8S�h�YT�7J��Nj�˿��}�����|��D�}T���/h#���>%�n��m<�ˌD�F�/�74�@�;�b����b�8�#!�Q#���Χ�| D[�ͼ(R#�n&B̤���;��(m�,������Y�Dٮ����\�1��_�/��a�"&m���#w&3�C���C�2(�r�*&gc�����Kz�����]D�sĂg����w���R7�8��KM`�5=ju11i���'�C��ˡlE�VD7�~ݡ�E.��J�� q6g�y��#������2(�s�e��v*܁�,�yL�[S�Y�ww(��;l��D0��9"�ʹ��oNIm��}�qP�ȇV�F�c�f��\Q</e]�!�6c������&�b���n���w��۞�N��mc�x�gڜ����><���t�{w�u��ގ�]��Pʵ~��j�����	I&37�m�"�.J����5PX�΢2��ץ ��l#���"'j�<��J���r/���!�ʥ]�G���� ���vk��7��J(���D�LG�m���)Xގ&J��ն�����(�L���ϱ�}Ӕ��Cf?�H*��Z�nw#��J9&a���٪շ�B�;'��v"=֥��L=�2��q�z6�����HJ���WW���{~i�7�D�o\&a��)�8��t�+���p��<'��s�/N�6������|����ޏ��i s�W�ҝ#�l�{B�r�����e�@¡H%Y3�)�C~�vj�h,��%��9�d>�b!��ٱ��w��㥙 =��}3�H���/5�
7T�Q�娉#l��R��#I+�F-�C>�.K��҅n���w?w����8���j�?�5vQW��yo���zS���fd7�D+��4�̅1keG	BoE�Q���Q��I��,�@���@�if��|7L�KG#�tqsP�b�~@{����H�ӱ�V�Ϋ/;�O����(P�.QY�귁<�l�mXH\�] a�*B�5�兑NH���~U�}� ��]r��R�!˸	L�����ѥg�Q�O=ǌ�oQ'[Z��7sH[�v��y��s�LA������?����v��F^��W1_ƙ
�����Ҁ�=p ��3��?�]ϔ�����s�]��Y��Af~kJ���C�	5��r�b�`��9Pz�6�$.�ƴO)L%�c�2��� ���K��p�y�e�b�@#^�}�:j0���x^Mݧ�B,o�T�D6Hc�͘��y���ݖ;��)	�gg�"�iq�i�P�("��p��On��v�KH@]G�q	�S�@�Q��Q�=_���n��0@o�%��q�9.�oY��H����Ա`y�� �O�o�C�j3c�7v=�{j�q�-���������Pju�%���E��$�����F�	��X:�d�m�d����.��fg����͸_�G[+۵���G����Dy�߫Gu[��_�uA�/��W"��}�R��"���9�M�����YaQk��tu[c�d��Kڕ:Eo���G%P�3U\�/�I}��l&�@��:h�S�n�B�ʭǚnϟF2c�Reo��|�72K��J|~^*��L�|���>�~{�Ok����mXc�t'����~J�W��/�G;���9�*V4OqVI*E����F�H��*�/?p'��4J����Xnp�#+k�>�MnخQ�����ˤu��ɿ�5RYKj9uz��c���z�8Qo�?�S�rĢ-�#���r� �	dً-�� 	^7+�1&90��}��J3��\�Z�����;���47��o2Q�aj��sL�&�?�bn+P`�D��d��|���~a�Ҁ�&T��sF�_%{�>�R�.�%�N?B�>:G��A޽�h� 3IZ��0`FP����#o��\�:o��D���|����4.w ��Nx�F[�0�[Cm�r�B���k���Ӳ!�r��sF�'���n>^��k@�@�B��Co�L�6�S�e�����{�ӂΖT7�t�I�оE�ⅸ-���7&���s�#M�z�h�	��˘VW�C�w�Uծ��.�(j	�g��d#0��<d��R����O��JtΣ=94��!� ���Ls�뇽�
�s����S>"��%U�9x3im��B6��^�0�)���^ ��̣�*�<��H����UV���~�x�NX����e�����ڋ��-E���܋�]̙N������3-����� �8�B@5���q�>��n���;���^Q06��`�+^B[iB]	�똊wL�æ���;���Q�����P�����;����~���Y�Y��Q���������~Wg,�y�%5��&4��[�Y2�8.�Od�R��(#-�������@Q����X1֕��A��"V�����pQr��
;�� �HG܏�B5�-�0(w��{����7�[Q�B�b"�3�'5u�0�J�yr�w���WҤ;�vNT�ޏ��s��: �R���g���,h�8�������l?�Gwqf��fW��:	�՘گ`�9[�+]`�{^���`�H��ۜ�*�'|�m��=��I漣N5H��:@��B�t��͡I��cx��]���?fr$�0	>��I�Q��*��[v`�:�� #�/�ں)��@@�52̛@U�+�"���������R�О*�~[,�y֓����y��i�����@ДǼI(���9���,·�~(BԔJUIVՑ��U��3Z�Z^4�Hj��䳜G�2�g�[c}��d��24��މab|��(O�bZ�D���矇�Ay����N�L���.�j��������	�ݽ�z����.n~���gJ����8դ,B���G���$<m89��
��&ϋ�P�6�d;�C�E�����K0c��I�n�����l��9�R<Bdǳ�ٲ�\n��Y���4�������ch�>s��x�w)̮�:c�M�~��C���{OD&e\�۶�1�S*�����H�W{K��A�N�_����j� ,���Z�e�$.��<��G(J��!##[��L#խ�_�D�n)h}��Z����v҄1�̟��.���׀3�jLb+��} ��ݎκ�ϙ׻>���z|3�6�I�t�Y�e��!���$�Z�����,�`t������b{ɥn�F޵ ��h3(� W�FT�-�3\�p�^�I��ESI�4n�x�P�r�NR'��"�������р�V8�:�e�xKz3�`;�1.L�C�P�O���%X��V'��B��-�s����)��Aa$R�wJҋoe�H����\9Mʴ�M��6H�LPՀ��@��߈�H���u*>�!��anI�8ܛcԳ�k�r����:��1���<�8�0e4�\�nV��B��j@%����Y�X�^,��v~5'vM�$A�*��) ���6I��)�K����R[�v|�E�U��l9�A�A��D�2��3�^���U=-�J�4������)��;V*�9a1�^G����՘��(�4:O��\�w���ɮ}��w^"�,Z�'�<)�Q��N/�di��Y�a��y�y��$�ʻ(N�]�M/i�/��1Џ챸.>��Q1vV�͡�&p�n�Qȑ5eXx�}�[X'Dr��`-=|�k��A�~�>
g�ɳ�7� ������.�4����x��;��F&��Σbfei�����]��A����%+�8��8�� �|�m�����_ݠ\�}+Ω��{�L�䁽.h40����O�FqrH{�h��<��@�<<�)/�����z@&���$s	u,=�3wmY�+ ERK�m�����>굆G.�5bq(I۽MMֈ���Z���s��B�:$*��h�`D�����ő�<i�6!��% B�5g���'�Ъ#>���6�8R/�����D�8S��r�6��͓��ߕ8��V`����OAs�"�(�-�իm����QY���i�����c݉�7p��^�ڲ��0�M+�))�(�����'Rc=唌n�0'��*]z�M��KZR[b���=�}�`B1p)Eyx��~�C�ʦ��}�Xb��K�7�	O��{f��Dی0d�d���(#ep� _e� =Zk"	qHJM[B¾(� �bu'a�!g��u�s�>B��L�Ox��zR�p,L�[zU0:����6<��=���L�08W�)�<���ng$���w��䫇��Lfl3�H��f�L�H��U�n�o�w�u�|m�}j�Y_4�^����C�JnUo�9�n�Wȵ��y�_|�yU�?<��m1σ�c��E("�Q෉�ů`��w�Ӧ���Z�L���G~'C��K��#��>�~P-dX)��<wOENK��q�M�]�k�i�K���	\�a����G'U+��W���b�嘢z\w�0�ηټm���L'ާ,��%ro��M����LT��д�4�p���.�^u�	K���+����*���/�p�>ٞu��Ռ
J�Ap�c�,�^��s�f��.Z�`ei,H����<5�^���ou/�%` ���R,���r�N�8����ղ:o��5�6k�k�YG�{��A�@����.�@�e�f����.��_��U#b�3���>+wxn�1��~=p��#�u@��9 �����#�Q���Y�x����hɯ����W:7��q�����~79-N¹�����<�>����ߺ�T�����U��)�h�<��ʵ�g?D�C��]�w�洈��6�`h�B&�:�[z��h��>3+��c�~�N��(����-u�>��T]�&&|%�Ì�:_����` oZ��Pz9[8<"�y���ꈻk�G��y�Lq쓲ʀ��|�a���G��/S�CN��n���M߃]N��e��Vw��݀��/A;�	�?��{©!lp�R�2���/�]��ID�+VGvF�ԶvR��t-}��d�
��B��u����}s4����ϊ걫�v��[��ƿ�����t��%�3��g���g��z۔���L �ܵ�Ő�wF��qAE��(��w��ҋ����3�u^w8�z�^�4o5�J�pF��1.Lk4w��(��r��:#�b�ة2Y��ކ'ԑ���Rg�i���`z�/��s	�%���B�R�ןL����сW�{Y�2�vğD0$U�����ݚH�O�o~�/N�H��)[������oE[����b�9n��f�����d��R�S\�im��PY���o �E��ܱI���#J�I|EUn3�:�W�~Y^��5}h\�'%�����y���[��,V#���˾�[�7j����Y��P)�B׉Gfz��	g_C|_��kP�ʇ_r�s:������+�y6l���r`S�{�j��q����!g��I~j��B�xu�����6�xB�K�A޴�D�Q��|�>��L�LV��7g��j�F1[��n>�7S$��Xì/��y�31!P뗐�?u��P� >��CrpB3�E��\�ucĹ��L� Y����-m���vXB��yA�g|G�:��p��"��>�Hh����r��?YqV�GK��-0 �/`O���}�y��?� q�+�/����A㧞	ww��,j^пH�O���TY}��X�9򠢆��w��GA�v!ȳ}��W�{i���G�o"o[���Yڥ2��]n��j5�	�}A(�/��I����!q�5���3נ�a���ӰmG[�A���qk��m�����|���:Ż�n5$��B\������]�k��m��zkN���X;�q�f}N��v'p��Q0!�Rp��y�,6�S��� ��፲s�����$gJ
T����^�q��ml۴��L���O])NX��
�K��mH�(8p%�R=P��R����m+2���� �3����C�l�$�Nٚ�9��;�c�,��vQ�]bD{S����*�ӱ�/H��UY�=X� "�цK��C��vO���}A��=�j�Ǒ�Ƿ�<<.�d�p���-��h��-����;Q�3y�.�����=������e��ޚ����PO��?J��)'��A���+���_~T3֬��;cY�Ab�j���QCء�,mgl ۡ
��o%"�̪�pG�?����ՆxNuL	�鄈71ޣ|��#*V��G7'e��W��y�(zz��R;�����;�d���p�$o�Gފj���$�1T� n���@[2GQ���Z3��z�_�&:@�t�����j�ށ��$���r�8[t*�4Ɍ2��8���u�y?Oɏ��?l�~�"��}.R�b���-�:�h�SK�������j���A�� ����粃<����~��m�
���%�1M�����km�V�i����uoP�<_�����T�Zd��*��bؚ�<La�]?�ь�ͫ0.E�!'���R-�<U�6:ׯ�$�xvIq$y�Mݗְ�&L�Ɩ£�b��i�Gr q �4~��� �mQ��
����9vf����`D�Ǣ����W��E%�z���}-�w�YJ��z������Ʀ(ĝ� 7�@[5�HXQ�#�Ck�%��#d�V�t��ڇ� ��"`�d��=H��ի��G��o�J���u�DY��O$l[�J"�;�`_Ԋ]gǌ�{�uF�md�=||��7ZW~X�ŞU7���������&e����-�}_3>�2�D�P]PGꔡ����P+?�y�^�WȆ����fY8l��T���?>�I�|6���~��F~�+	[�yu�p��&��]�)�3K�J	�V�B쟫�b���kR�r�t#��au�����w�		C���`��s����/];M˻|������{c�R�쉝͟-ҌC ��'�	w\��L�(_�����D�t�l�.j�g�Z*�sEg<�;`(��1���+g�Kv�cu�ӓ�X��tf�KՇչ>a�5�ӻ�O���C�����ya3O��������٥���L�D�0��p��3����^�3����1"Eth'�����8�{��W�[��0s�v�j����̉��ES#{&��*�Y5ǜ�ϝ�!h��Hո1���W����^�;�BF�X����W ����D��I˃�v���w���ӦR礎a�O*xf�y�d;��v�M�
\Q�
l�I�{�;cSU��l�j0�� ��|Y���+�n����������W���sx���ü�Ƌ{���n1y�a}{��C�r�Z�YFS=ZL�zXE9+�q�Y�'=:}w7�@���������w|��"����Ara�G%�_m�3�au��Ƨ��9�;�xO[� ��1tlP4]���sib���sF�f/Pu���/M�V`Oa���˳�v���$K�����/�;����s1�6-��v�'���l>APHD�%�Sr�#����ָ7l�h#4���uُЂVS���Y}��������ڂ�d��	�}(B�y���v,�J"F�_�-']��G)rK�,�ԏ>�?�aym3�辐TmJŪD��Ҕ�|����;�c��-MKmk�ٯ)sͮ�C�̵�],�Z�LD�Ev�L�A|O3��[�����9���T���� �:t�$���.'d7��@�n�f��9][�L�)�6���M|ۍ���tzǵbJ��̜��"J�wP�#;[;)���2_e=
qp��Wו�!��Do�-��%)�/��}�3c�:L˟>裐C�K��Ia?K�si��RDe�C��?�-s;�h;Vg�f����4�y�QP>燂c�h]�<��d\���}}?�	���9p΢�%Ht�=�k����Lxu�g}�ˮ C�/�M ��>���<
�!^�6��L�o��Y"KGm3�B�wӞ,'ʚ�����z�t�8ǻ��ܓ.�wĦKI$e񕒡>0�|0&�Hs�7��r��l{$%"����z+5Yr�'�~�ᵯ�/�f#�%�Ij�Ep��?*��[
�1qKi���d�`�_�$�➄G��T�!P�d���ʓ#�Օ�����4'-<�(�k�K̟��eC��/n��Cͽ��N��J8�c��`��;+˴�x���[[
^��?ձ>U��:
����xTr�;
�δr־�F���e�_��0k�T���t�]
g������{���1���R��$�a��հyF��'h��6Ԗu_���>�,���⭤�M)bh��
��H�Q�V�	,QC��:���ˮ>�B[72.�8���5P*�w��g�5Ƙ�cdtk�v�$�_H�c6�X��昃r�¥烺d�^�YȢN�沘N�@��b푱�
&�V�{�@�˷��&eu�~�cɔX��V��W� ����ߨ�ٍ�!W�����7r(�Tk�L����Ġk��(eY����vx��9 ,��(¾�<-��"	b"�C<V<��i筥od��5�Z)�~�ȸ\>���,E��j�}XV��͟i"��B&���l����UR#�?�r�X�AK��.#�K�3;��n�����ßfJJ����i���~���~�8G~��j.��*�ME0�P�l���M��U���o��p(:l,�gB-�B�E%���5X��?FL�\��c
ό`�JּM����JCv����a�,=/ؼKM:B,9$N����-��ַ�Z3� ˫B�]W�N��R]�U��5e���a�u���t3M���Awώ�8��2�,f���_|������2������� D��ߑ�T���W;h,�q�}��~�<�uKv:����kA��[�
3Y�eA#�?�n�C��f5E=f��M�E�I�6�M�o��P��h-v"�7��@r�3B���ؒ9��t�X�1%af�`ο֫���	$�q1~���AUl�b�h=������|*b�Xx4��AY�p 18Rnbh�9l�~�CҋJ�n ��B?E3}�5�Y�t��<\�8�oV�9z�����5-��XZ}��kT��i��]�]��,q}	|!Q�-�t8H�^IM�b��ZC���H�.a���Ж~�*�ٙ�e,����J��L�]G7�.+�{����mJ�ma �T�G������i�T��D��8���]|$��R*e�z�{�\�G��wwP���Nj���U�*6'�HY#8�]],$���S���?��ܝ�h5����nP�0�p��s?�����s}�������i�
��_����LWpl�D�P����(3�&�0嵐x�3j�u�;ە���#�u���#v���7ch1G? ���'������p���=g=kWD2ԟ��V͓�Hy�)�x|�':(�bG0ָ�ҜI.���@LN��L�/k����C/H�Y��HoKv��O�Yt\�XWaz��}j�O'\�j��!�=:PP�cI��dx	�'�DS�� �UKF��Nx��?�Dc�ݔp&;�N��*ukF����F���&��{ɥSTC��#��☡�Cf�WI������h,Ѱʞ��E �1�$gxU6`�(uTQ���� �t��pV���P?�u���9UKã�\S����<����a�e�O"PR�h�ZWs�S��,s�����Z,�zs̀2G��U���P�鼢z�ҟ�*P7C������_{cH)A��;���B��ݑ���wP�d(�E�vN���DϾ��l@Wș�A�����gp�X	���j��c/;�*>Ҥ�q�c��X���M���2����^Ev	N`�I�	�]p���2����M��<X��M��a[�g�Vm�#����*al�2�s/zDl���EwD�]�����$[��!�Pǈ���MCl��� }��}�"E�ÏO98�hY��C ��b1�i�x��3]?d�M��$!w_3!� K����)|):c���e#M4<�����1/�@�o��i��ۗ���y����F�R&Z	wڎo9����'��:�a��������Ӫ6|M!  b۲&COr���ٱ�R=���m�\zӀ��?�.��$i �.M�F�_{�Kډ�DCޟ:���'�4YoP�b�Ҝ8�O~G����ta�о��� ����P��eH_�Yq_{;(~���j�5�8���'�!��qr��ZK�qq���7{s;�?�j��r�V��e�8���O^Z��1ѠQ$��9#�g��m74�M����]@y��)����d'�U���f���sQ�ɑ��+�J
��Z0�%��}b�#�:3��G9%5�/3;ߧ�:�bn�˔��$�II�V�g���vG��_�R����C6���%��j����Cc�T��e�b���@�3PFߥc� �:7������?S;]~R#�R���~��K�.-}��^KF�bY�)U��ѡ��ڙ����ER��	a��h堕��E5��ċ��H [�m�҆|ؐW/�����
݈+��2�'����%w���6C��o��߰P��Kw�"�v]����81�t3G��D�mY~�m�Jhm�i���_ɖ&y���0�#c�?�]U��)�kj�� ����{�~�p�f��|�xEGDz���)n/ұ�Uk���/�Pi�P#XC��tbHǑ� �&Mm�&~��P.����-4��b�͠���_-�9(�#'�Yg���c>I����a~�T�����3jNA�Z�(���o����Z� bD�u�(�Py�O�����x��[�̢#�x8��㍨��E�/����u���8a�����G���u��õhn ֐�"-�.�1H�R�c��^��"T��"M1�Bg���g�M.����@��A�ˡ������//���J&L�EҤ%ʫ)~$2/V
Tw�n��h�z%��3k�X�K�����-��GR[�;H�k��պ�Mє�N��.�s�-w�Vk/b���ͭ`a��i[�.��ޟ���:�fd��F�7itҹ�}ԫ�5�B()I�I��2Mri��;�W3���Uo�����D�eE�����+��-��5oK�"��m��H�~�q��#���5Ȣ��`O�8V����B��P��A&�o�S
����n���9�C���nb�\z��x#k�ְq-߯́*!�uA�����#��`���L�:�	&(�pz.b$o,B�0Ӡ�I�u��7 C=|yx�]��G4����Tnw�s��x���|M���I~(F�@�g^�����U�Ԍ1{����^��l�����tѺ��.��ǟFyҲd��.��iaݿގ/��?il�����dtWnN	{�G�>x��:�<��7B��6d�uݳSmjG%���^|�L��cw�,�{|ax��
�b�m�$t�Mrl����ݡ�`�k����I�bdm�]�C�L`A6��u>TA����L��Ժ�� B��ԗ*�Tpa����%��۪���l��yם� �I6�#%�Vp��oN�vy�d��!�I��a=FŰs��or�ɖ���1�L=�g������f�3��[|Uj]�N�jt&/�=�Я}*��n>��N�L���=���bq�7��j�ĚF�_�F�;�^��:�)Im��&l&��P��/�M�m�U�j��r��5�,�>��-5"�H���S)�w|B��;�ѱW[#�L�����e�O8 ��8���ݦ�%���tl�fʂ�$�[Sz`���Ć�7N�FWp·��3T���҈��"സ�A+�oR�@��4�n��_�F�X[6�o�y�T�@�C��X�̐abFD��(�>�h���Wn`S�ȧ�n�]t�`,.馐oBG�މ�zc��,��ϛ.W9�ώ���n�Z�[�>���ǋ2�0�ܜ5�u$D`���3e���a�W��0�8�UoG��D���^���)	V�b�	�f:]q�����p{�s��yç��(ن��:ϫq�*8j��$+��qÕT�?Zhi����Cf�b܈Ӂ�����e>�	5�G�Z�+s<��h7+�uD��v�j��x{�ޛ� �z,=/ދ�nhA�I�D�V�9h���/}GS�uטqJ54}Ǫ� ���i)����K"WH��^��ވ@���G�J�*�O���G/�)�#��׹@ڦ+�Z��1գ)Xcu���]����	9l�L��͟�	@����=�t֝�0������j��·�`q`rdH#�M���xћ�2���ԍq����!B��B�ɋ�0�)�(u� ���4�m[�����(9¢�K��G���`f�t)p�g����8+OP�����L�5��^����Vخ�e�ya.�`�+�y�HU�纞�\�� }�A�,ɘB���nja`���V%켼h�ޝ�%�v�ByF;.�Um�$I1�<�p:�ԋ�1wQq��y<���:�:1\����m�U�C���/l�"��aɁ�|�)Pх�ܩ��v�~��II��(�<��hiӭ&��6�0;�R�N=P}HVm���Ɍ����҈�$����3Bw�Cռa������A���sЭ��F�S���
������*�c��l���ޚ�{�	��4
]��-N���9-��4��w8�cV��îA��h���;�{�����n׈� �+�~�ˉ��v!��׷>"q[tC	�}�	Z��O�&Dl��0���뤷b�{.s�+p���'�~X>F��y�N�l0;=:+��3�;���w{m@8f>{�<U������jQr;�m{�����4�K���{�7��V��0��!���UC�/[���]2�9]1�!��:����&R'ī�h~g�tz�_�������e@�Su�l� ���]^��
������>0���9�Ğ��N6��M-D9l�e�� ��~������; h/�,�2�œ$�\�Ȩ�� �^4(y�������4҄���ݛz���?%�_�$D�L7�v��w���p_0������'A�Yk\T���C��a��NZ�� ,����޿��.j�;��ߋ���Bu1�_$K���i[u�K�ݞk_�JW��ђ���ЊZ���ړ�xcl�3:�ʛUW�i0jU�i8��1�00΋��8�v/.��3�.5
�ֽ�R.f�=#�0=ĉ��d��y�љx.�6�K�U��1�߇0C�M��Ya��hQr�15�bӠ�A���'�h���M��і�:�y��
O��Q�+��d�.��(p�$�	��3ػ��1����.:������55��/X�GacȺ����]ӥD6����Ĝ�����w��}w`Q��G_ iC�Z4~l4ی��;���K'�*Y�m\y8�t��1��*K%���)Q/�UMq0v�;{�Į=�5i	�˯j��[;�$��TRZ�$Kx�Z�S�������(�A�c�y��1�
�w�S�+Agf�i�����OaO]�@��V�1S�o1FY�����!�(5H�d$�4��ؕ���e�_�7)����v:�^/̤o�=��0���t��8BY��_�rN��hb���m2a�(�E�&����D5�Mx��%=��j?ˋӺR���#.;^�WY�D#-ldY�M����Ǭm��"�~�G�OJ"��;}$ˏ�I��O=���J�>�\��\/ց)�*x��a��X���U�f¡c/�΄�8.Ϛ��i �ρ�,��!hJI��*�v�s�~��MI��鑎l�>%��5���z���M��R*>����l������X��lDv��ChE�4��ԊH�������J}vz�������g�Z�{=�0Cdi�3�#�F�Y��!�G-/\�2P%�\�I��Dw�߼	�5{X,�J����WS���M<�J��*'��ջ:1UM��D?�]���\1�N,ծI7}ʄ^�Z+t,2���ꐍ �\��*�U�2�oz#��?_���x>�"������_��<���B�O��3������1-�D���W���l�1��7q�Զ�T�!r�4
�\[ey0���i}wt�~&�U�Zq��ҏpv�C~;.�a�3�&�#�9�{ی,�AK��6U�%6�{�]|3������~2
X���A��Z�T����z����Mzn���pD��S#��A?FCV3��k��T�0j9d�F�G��)��o�2*Ow�/��ޢ�HV�����j�������<[�(�C�6����xo��W��*D3~=l�l�Lż{{����_L�|��o�L��Ư���;���n�-�'Y��ٍ��~��)n|�穂�:~��7Gfw3Êʇ��eL���F%���
�Y3`2^���G�S���OK�������q�,#A �����#�%��?��RŊ�!P�dm�X3Ӛ��Y1�݅+���9O��n�))��U�m̘t�Z��M'qz&�n��ˇ�4N����/���c�~N�ԓ����"�^���_�d�d���z�X�be�e&��]�0�q�Z�	Th�s���j"\�>�"��?��+��ɩ4��Ӗ)�T�k������]���}�a�I�V��ɷ�nz�����yB�ٮ������]b]{x�7���� F�0M�9Da�����i���3h��o�ڨ�e5D{����V@�;sӺ<����s ��W��(3��;�@�l�q�m��Wg9~������d�;V��Z�W3�
rm�]]���0?*���r�sg����pE��yTW�4×���y������q���?�����6�H+F�^� _5����t � �}Z
?`�Z�O��F�����4G�~��N:�e��P6������g�����Z�����ХڃFw�l��h ���lC�Dk�Y8 ��P&����� O��<�����<X`��M}�ϓ���w�4��EX��k�>��������%�����Aάz;
���2�hNf�)�5
>+қ���%O��Z�b�)T\��:G���) �Q
u4�o��1��0��O�C��E}efܜ�.�_?�e�Ù�^1��i��v':�hg�����Z$�}q��}������`��u���t�w�R
�f������ڟ��q:�� ʏ�<m'.���\_%�zn�~�|�'�r`\�Z�3��/Z��ɉJq'8=����u ���U�̸�O3ƃ���O�*�L��ڤJ��h�2�X�'�CD�J��6��seDŎ��bŋo�D�5L9���O�)��`4 f�vj��n�G9I%��F����ңWfo7F���5��yE�Ņ��iǺ����Vݨ���/"S��'ceP���3�����$�٩^�vq~d�j��`=����yâ��:9��}�J�,4�azl����`�<ˋg�Z��O5~�?��0^ �/ci�� k bIS>B'E�^K. Vl=	��Y��AF�j|f����IE[�>��s��ɭ�˾�B�����X`���˕j�4���ج��t1e���y�k�#VTF�MS��oŀc��̖r��Stm�WىW+:�rq��s��1�l$�u�j�XW���
Wg�#f��=��A2K��S��"�˅
����|��FE��Ԏe,�:�e+޶uv $��U�jG�>�����ث�9N����XOROA�Ϲ���~!t��*�уo�=Ɏ(��\���h��_�\�L/wNcF����Ǿ��w��@�]��n���}�������$���+J,c��,�hV]�I�t�G*��;���H��a����(ߒ�?�~����o;�u4�����r90T��X�;@:R(�g;���V�f��Y��&���#Y��G�)�Z�dNM�x$n�#[��nR�-��[/׳C���դT�"Q��{�H�h.�4��Aq��c��ȅ�� �����QRg���*Ck�͆�e�"5�+�Q�-0)̶�d�:1�nO{��݃����3�_�z��<�tzsfÇ�s�J�%������5��K���AwY��-� '�2����M��B�x�w��4�~b���g�mɈ����a��J��Z���3+��;EI.	L_y��
[&K�zzc��z�\�)�����t�{p��$F�ޔ�0��3��y��o!����s��J�����)�AZ''RmHhm�e�>N��'��97&�hL��$�|�ƻc�P�������=�)�؁����Z<�C���.b@�ɖ+�����Ȓ�.a�Y2�Y��2��4��u��JOl/�U�����4Ѕ���Â�Ύ���ٌ�PB�!�_��e:�JjMXZ��&:�_����;��>�k'-�rv/��YE�z�y���_�f��^��g��d6*ƅ�7����ų|;�����p�ٛ]h@9;`D�4�f���pCI��7�e�6�fJ���t�Յ����LB��z%�O�u�p/쁚K>DIHIy�	����,�1���F�@f�l��5�D���bcd�n��(7��XB��;��1'zob��r��2�>.�,�5�Tl�P�S��$���ض%Z����q����e�0���"���Năt�  FY���Y�J�6�a?ص�e �3�hg�n\����N�m�\f@�w��VmmK��A�"ܓr�mO���u�[��K�hi�bA����8уȎM$]�$�5_��UU"�,�U��J.���6��x+f�p(`)ώ���TD1�w�x`2B<���W4�?��鯟?�ߍ9���	^�7�9��lї�k���WfmcX�4�i��,���I;�ԭ�6�dX?� �t~yxX`���y ��~��OV��/3�W�d<����(�A�'�;Irn���n����v�b�����Yc���t=����!�5��6�Q�C�j�OJB�=��j�>\�/�}N#��g+4K��$cI�	�j��|���Z�#���� 3-T����=��"lo?D�S�B�9b�����$~��k�*#���w�a�6ə����7��*n���oEe����|��3�,��D�g����<Rز갾/�#�����F=��S�Zu8�)��}ѳ����p��yb�B��KY�._C�v�:K��w,���U�z.����kp�<�9��Jh`��N|p=�`�6���E�����~CO�	�+	[I��>�4Yk�V|�(�wu�z��D�ց �CɇpS�Q�#�Ef�0C>r��U�_�[Y�^)Q1��E�k ��Y��:���Jp���v�Y����9�i?�FQ�袟Ԭ�ϣ6����FX�w劷?�Y��P�ŭ��=��(��C�=:d�����<u��Z#HJ���{�K�1�Tg�rPoّ�a7--$��W	�0uX����o���⹘��^�1�j�.ú�� o���E�E�� 	[wLF�]��{�D��dq\L�*$c��{�
U�$s������+�[9]Y*¢�ƈ9����'Iܸ��$�v������
�C-l,��#�4Z�?Z[G��b"K�~�zg���9̼%���Y��Qz'�`�>��/�R2$�����F ��Z�H��X�P`I�*��6[Xk�k�������.i�� ��쁸�	�DM�/k�b�0�j�a�,���B�(42�j$U��h,ͳ�È�v��*g�A�Ƕ_�ލo1 ]�d��~��fk�����: 'wC#�$�VU�oOG;�Ѕ�y;B+2��X,�K.��'ռ~�cBJl�P�D6j�ѺV�_�\��ā�Y��ӳ����ί����X���s蘻�C��ٖ.#�B<I����@y�=�?��a5��C�(�&{KA~G�~+������W^k1˜�#�[�����/�Ve��c�:a�KNM�C�g� ��W$��'���2^r����o��g�#���xa0+V�M�����aV�M��^��7{}�j������{�#��6*y�M߀���aQd��O�Z�n:xE�� ��eKV�u�[�+��uNĬ���Q-[�JFx��o-�^�����h�
�N�vj�ԛ��~�'�S<�A�.��>�9O;�[T�̒����~b�q�S׫�>����>��*�[��}Sw�k Ns�p�s�Oztg���:��n(#�V@�|�vS\�G��U�M+������`Li��4z���7�Ѝ�#F���6�R�·
�W�s��k�(�p����e�MP����.����fSn��kc����H���K6<��汀�C�RT�/�����t������*S~Uf� ʦ�ṅ�[�8vR�\)-d8�V���F��.J{�����L�3�e�5w���Eө1o�5�a��4�mGx�5�OQ�i�i�������ȯ7ET	�N<<�yP]�����}�r�.� tQ3��h�B�c\��3�P.�T��\TZ3&��6�;t4T���q�$�C*J�ٗP���8�[�73�1��v�T�~̂�٥Ϊ���2�2�\p�Z4mo�̶t!��rJ������%,����!PV�Q���ڢ&�!���ԁ<<23L���i�@�=��H���jR�YީWH'�D�	1�+a���nb��z���+�U�b�� �&�vя����	}ƫ�/�=��ca,��ƹ2sУ���;�Cf0 �e K��>����b��1�`Uo���T��;5���	+~~��虡������z5ڹ�ҏ�b�?,!#����)H��6Z#���4�<9j-��"������;U���[<jz��o�Q�kS)S?Z��.�oA�ɓPc��|��䕹�^�����.!��@0�EYP��Ldi)���(��TTZ��v���ۚ�K2q���JQ?5NĚ������ҏ��N���������C0Z����YR����c�"(���vNXM]D�����7�P����@>m��,�z�݋�=��蕹K��7vn �D�5��W �;u+	$g,�Tf��Em�C��5���Sg�[�\k[/Rd-J�P���[���.�jf����A�/ˣ�j��R�
^��m�4��=r�qd#��M���DuKǵv�J���k��YVat��g�.��ݩ����}�杵�Xѥ�_x�-�C5��;�J�o[ۆ�o6@�p����9�� K=�d��*lo��rRM��M�0����gO%�[6|?:�M��_�4R��| ��?��ό��J��	�����1��kw�~�w�^n̄�����D�ܪ�,�jɭ��o�T�����6�&a!�����H+�P�ADtb����B�A�R�MA����n;�d׈-�Cfa�ۉ���f��	�A�fW��/�
�J�j���C�e (�����V���1/$�E��<�O��c �����P�k���Q�;�Ī��D�e�I�s�:̻����6}�*���'�Y�i���f��.E�S�tR�?;����Eb9�C�)���Շ�GIgxyůW���;(�+C���V�m"�x�a�Bl�nNfv1L�u+�u�8���╽!��#=$mt�9h�>��r���V>����x� �Q��b�
����v�������p��ݮXY� �n�R���.&������C�&�L�&g���K��_�	ût#_h5L��	�*�I��L�����U��ѥ2�4x�N��M3c�0(��ꃩ��R.�oo����s���
�/^�(��S=�����r����ϡm���F�U�2�׻�Œ߾�1�V���W�*#��5X'k�8�C&���e���������EF��k����ZaSb��-UG[)�1M� x��������Р����;��[)�d�֯�Z&$P���zZq���GR~�l$�RrtfnK�oJ���OY7x���-��[��p�9�F~���wУ��w����r{Y�Y���K��{s�~�B�m�[�-�.�������JΥ�$۫��a$���T���K��H�=2Ky�n�ܵ6��;��{JlM��>ra�fݢ�w����_p�Kb�颧�h�/A���w&*��C�84T�gO}�����J����%Q��j�����!Jh�X�o�vA�ߨ�`Kn��&�o(k��vp(� 	G�T-ہ�'�>�wuR�L0fR�a?�5����2�������^��܊�F	��,�w3�Eٶ����nT6�N�"���"�9�
�+���\cU.�`�6�y�H�;H�����S�H�
Uɱ��L��/���n�8���M�8%�QF�,}ǈ��ܥ2�9�y)���(��=�zR��ս��~\dC�fB�ڼXu�èV�)��W�~Ϋ�jJ��p���B��3�~��*w��g@;���51_�HC��jw!���u�������l��\n��*��m��_���f��~��8���!�*��b@�l%�˻6���Q�TF]Z]=(,hIkL|=�#;������p�|/~��`��`�Rͧ{�/��^%V�N�|��A�2O�泜�`f��͕|�����GZ�����I0��<L�Uهs:���dF;��q�gW��o8��S��2���� ^�سn8��ʁ'`�Q��0Z���Q1���k0�q� g��~�W����F�)�"�I-�B����Y:)Gu����O���Z��$�f<k�@=��Sɱ�<�l�%�c��bZ�& �����U^���.pD�����B��+�����${h&1��Niڕ��zRX>� 6\��kj�9�M�����)d��_89�\�V��
fρz  �/�3*��z��sL��&�]��b�c>C/��d=nFTA#�W1�������#
o��Ε+��)P��q�r������
���c#u�q���PJyK_*�v�"є�p|�&�ca�)f�a�$N�>�M	[I뼤w]J�񛰖՛Q�!g:�|-�4�Ri��é�Ʊ�{��/���G�
�x/]}LA[�:�t�Z��*�2'u\P��]9���P�iq�ʒ@�HoZdq�i��p�-��1<</��+��pJ�yM�A�g�N�2",���=��$�,ϛc��B�7�At�`�m���Ň�u�Y�i]�VP_���-V�S�9��/ءj�V�\�ݷ���&��N�X��x4���_�P��(�X�#z�Z�^��YXe0f]QW��a�R���g;S&�~���%�yΟ�7��	#�����)ܛ����s���� /-uK���|U���k�(&[�1ޅ�m���"�0D\Yk\,b�py3�z����$���àђ���,7�+���t�RMEm.B��U]�L
��ЂV����pb<x��J�K�˴���2�[*��� ꙃMA:�q�r{ii�S9!�;G�V�b����P���t�ARA4B��13r:�"7h�qh�>�����|���^�u��%a~K�A�Å}>��ĝ������2�A��	�%���
�~91W�=�"�&�o�����)��������A��X���|�:����]xN8)�.��阩ڿ5(�>��*�z�����$YB��!ɰ�K��X��*/A��I,�o4HH�^ym`�=d�$�4�|��X�N��xA�|=�4*�E��u��}!�u.�\I��1���N!�;|5re�: �ꍎ�c�-F{���w�˦l&
��j3��ʈm��ؿu>x�o"��e��.��
9��>�6��s��aTk�y�#�U�a��w0��Ad�0��~��C�uш@�B��>�g��O=���1����j�x�h#p�Ї3���CZ��e9�-&Y���Wx-G& u���dy�ʨC�����?P�G��1,ԫ8�������Ȫ��O^��&{׌�d�N>ɧ�ڢO���� ��ٿ�KH����^y���zg=�[��LX����7N�]�G��JT�[Ҹ+>���{�>_���g:S�\)H���N(tm���e�I���#���+dcv�iL!�T���TI�������l�dL���"��YR#��x3���V�'�iM�{�/�5%��r�
E��\�W�`�#��O���T1NA�X�C�D�V˥&%��x��K���Ȕ\
�k�?Ĵ5���X��`W*lXՌ=!�g��ǝ�rN�`l��W�n�q?<� pr �w��Ǔ�������^Ϣ��J�0���|�\��л���k��#�>B�{�ȡ\I=�/�/��jZWJRo�
�K�2��(dg6���+D� �6&S9"����KQE�PE�b���0S �Ya=@XT��u��R�D<U�b\Q�O{MF�qV�k�R5�T�vo�<��GQ�P%N`��xI�5n��GHܕC
} �5�QJ�)�K�@�,�o���C
fyK���`�(6ӡ�
eX/�����UI��p��O�cC>YCQ�~dmR��4^��bU�l���ӳ�K�^Md�N�c���T|%�'��U~���$%@.-�	_0?�ۦ�.�Vm�o�L�x��r˓�Rv��8��o�w�E\X�4b.3q�aBO�����E�g�Y�&rE�?���__�goA�ý?0m?E��� ����X������%��ۚ�2NbԌ\'(s��Һ�U�2zg�CN�
���&|~�s�"��5@r!�_׫�҅������C�`�*�E�e߹د�65P@�o��S�zf�N~N&O�R�95ν��r��S��:4힙^"�f�b��b��i"F����м>ɏ�F�c���HK.b@�/	�J�o(1v�lRJHvt�����DҎ��HqֺR�>�Ks�ɐ"��E��yL��*L��wNFu�`3�ݬ�l_&A%(%q��}g��N���.�Cpp��Vn����?��DzbӒ[�J���H6&���7��ѱ ��E[�i��'M�&uM��8g�ݩh:.��@�d.5)��A�����\�bb�_�bCd�>��lxV�,J�.�Iڀ��i��8�1o���<�����r����C��$I+�e���.��ϗ�Gz+�E_�9wr^Í�<C�x����
D�(�a5���ƴ{���R��M��ޥ�AS;ֵЇM��m�������&R�{�A�ǃXN�чr0����=(�i����ם���m���L��T*V�!x(~<������4M�W%S��{n���&PX�6��
�9���|Y�zؿ��1������ZN*���I���>��aj�%�J�q!US��`0YiA������g�0��Ƥ}����
lt�Z�`���k��x�D��w�3�h���
�hh,��ą�bF���1&���t�J�z���p�����"'�x����v��矤(j�|DzɹH�-<��}u;꽵�y���8E����� �]*��[O��ɡ(�MC�;0��4��?�������'ė�O�\�����OΦ����b�Y� 1ӥg{�Xy��QGbQA�擟$����{2���F�o�pK5��c����G���mbپ��U�|�n����z=T{rM|.6��%9�\�,aq��[�v�"���wY���&*[ ��l��d�a�xa֒�Т�BHTD[fj�\?���<|��̷��Xb���B��]("�!���0ڑ��|��Dx�+_��͏��]��d����&�YhYim
.��_늸t�;0k0�t�@�a�;�ն�ܼEf��V��/�t,��k!�{��[�s����;�㋎�h�:s�'� �yٶb~8�[!��]u��A���&Oa �,��\ X��'n�X��������/5��-/�������kk"����v ��Z�	�5�O����5���ָ�ή��yxu �jd�����X��cs��ops:���r��f��C�Ђ6	�J-��gf��斓Q�r]E�g�����HW�փ�vH��Y�6��H��&�'���0����g�7����[m|h�2��f� UT�F��R�j�0Gj����k{%ʥS굆��Q{�oS)GAC��R�Q� �Rzty)hY�b������-z1��BE��YH�'g>������ _@�IYJ��YƷ"�'��L��(���^��`B�GF"���=X��-6�k	�/�(<�A�t�Ď�L�UCQ�!F�2;o�u(q�
��(.�-jbVnb�)C�&`[�ñ�]>��Ӎ�A�l�a�]��u�;�f���⬁����D�d~/�i�$�SX/I���&`��E����?#�� ��=�w����O'��Z7�QK�לDjI�����0�<�� ^�ɚ�����[fg*ryW��>����lw�2&S��wo�
�~��Z�Z�L��9��j�:	��b�Ib��zg��E=9D>�����n���z,#x2Tsd'��|X��+\�&�5qҊ��SR�k
��Q_����/A���>�tҫ]2S��B��!�"fqm|���7IZ<����m+�E7z�Ϯ�c=�6�DQlFY,���Qx��ٟ����0��1s�4�Z5�W�j=O3̚4�I�95mP����$�&�N��+�=j�x���6�2����9@�9
?���
5Q�
w�`�vu?*��1Ъ���H!#�� �b�]e��k������6��V����ܷ�V��j[�Li���̅���Gp239ә)q�P�Y�A�%����Y~ԋ0�X��/:=ѱ��9���v�j�W�u|T�w�G4� �n��d���RIrvG�����5x,r=��CȤ�o��p+�@���iA�ɇ�I�MQ���&b:A˚�,hU�X����&I
�Rǒ�ӻ��3��ȇ_oޙ6�{���v��Y}�+���n�~Er5~A�RD��D�s)���g+(F����[탅�g�p�R֛��L���x��ɖ�V.2x�?Q�I��7!5u�{��"��0	��Ėm�,	Rݑ�ԎsFBzz$����u��R�8=��1gh]��Z��[M1QO��w��m*�]�?/��2e��/~6T��x^���6o�+e������-_���	�<}����]GX�4T!<������9�uO6���̆>L����y-
,���G(�&������l�a�h6`��Z�V31��,*uO�-�t����b�c� c0=&�g� -$n�6�>Tt#}� ՝mٺ3NT�C���A��:;��VR��AU��
@I&X1F>���݇�C[���9/
�Z�/m�L�pz��Υ'0��C�_�HF]�s�o�	�Nw/Dm�O��Q��V~=�b��	�1�5`Mh��iD�<�D��Β���	����]"�}�������)��/�mN�V<��D���|����o��MujIR��!S�/�$���z�Yd�i��A�j����Cȝ����aΉ�N��ce���ѡK�*��-Oq��(�5�2�.�N���NX}?]~��vl�Aa�`�CQ�$���-t��9�7�k���E��堙��^�2���_x��B�Np*�;�0ڍ����q��d�Zn��gy�1M������!�;1��^IYxwJSK��u.��>�X�v�x.G>�.��.#`S�F�o���D�k���يg���E��&s�<�:v4�І�}�DfR}t��+zv숶u���qY%��38���>����M �z��m%��p��{ej�a)B��Ҽ�`>'�j��Al0��=�R��Fr7�O���_���r��C(z��mUWM`�͛��e��0������zL\���ik�i70���V1A@�lxw9�r�Ԑ`.��1W40�_2����w��=��<�/�K~Ƶ���	Wl�a�9����I�	lv�7�؏T�+�@}ڀ�{���V�S�9�:Y9��k�$�����7B��Z��P:�BF ؝�E�l2�Aӫ�����>�~[�L:�����AɗW�-p߼S-Pz�]}$�@;��:zQZ�N�����#��P�X�CHi+����h�7|����8���ҿ��OxĤ��Έ�$�UNZ-����C�=KLj�/��}p�l ]�C�-�5˝�U��!���'�U�*=Y�L�jJ�S���o���(n�m{d<���$1W�� p�56E�e�i��I8���v����;�9�y��^c�f7��f :W���9��#~���_�������
��^��L�|��*{f� Ju���z��Gji'�<��	V�m�:��/�A^oQ�O�f=��I���:i��Ǚ��o�7��|��y󕧳.#Mg��F*J����(<�0ͧA��|��N@�ԩ�Po[�)�u����0�O�ָi���[��5�	��K��$�?�bY��d����0|�6E`�g�D呅���l���u��XĤ��c��{��p3���6�����K�v4W��O.�;	��/pc�fS�b����X93ܨ!F��EϿRnb�"�j����_�/��mt�� ����3;>����$,��%��Q>i.^�3�	:��D���mi0/�y�������zK�;�xL�ɾ!�1u�����L���z�����Mx�e�'��P�j{hL?����oL���-4�<�L?j{�C�66dV�2b$_����)Xu!�U�ʖ/D+-�(h�rFase�'R���e��~��]A���f���6��))n-�Z�o;C�p�XD���;b�0��_+��\r�JF�aՇr��vy���L���;�ڞd�/�c�Wn����Ж���]A/������̳��_����a�B$5q���R�W[�zeG��[Cv�����\��2F�c#>6QH+�O���p%���S����\ˍ�.�qTʰ�
�2-�?�1�*A��&/��9�jg��噀��n����J������@r�ۘG��&G�02���K�!p�\t�Z��Ū�u�"r��#�V���7��G�Nq�B�?�SR�#z��l��ظPZ������:�S ���4X��<�&a�	"�d�9��"kq��-cʤ@ Pom�E���y�����T}�2غ���W;�L�<*�%� {[���KM��0z�X���'4�����|�|Bo��_�|ι�����k23YF�%q-�Lv�~e�!IN�)�R�cڲׁ���烂��Ԝ�
,Kș��M�W�B6cl��؉��$sR<�����.����Y�_�\�}oq��k�4�`4��hG`o���+-���[�����;HH+��R�1�TW�V^���P�ޅu�t���ڋ��JH�YZ �CA������C؃Nz*O��|PTD��4�[�)J�:9�Lkǅ�q�/�lC�}�>fL-;�û�Y»�jZPՎY��V��/�QYJ(0W��d�s����}I#;Sٙ	�f%�|5�&ׄQ&�TE��Uf�F?���)�<��!�K��O�h��61=�X0Ud���o��M��b1I8����ByA�m�h���X́p3�K}�IEUk8�`ʶJG�K���܏�X�l8����X�$c)�o�R�>;sk����+zhw�pE��A1Si1_�t�5'�7��ɹ�Q��G�9�����7{�U=ǧk��ƅ������r��93��lNЊ|��K��K�-����/{��?�$�a}�����2`��\`�<�s�P�A	�%��:2ᑾ���Zs��3�$�ȳ[i�r�
����*�]��l���V���^����Ɇ���z�f��l�o� �9�����ϫ�u(��>0'o���	%f<��zӾ>�N#���������U�wL��+	���Z�d�9��u�j �?��!'�&	E�Z��>�������+J�����#�X��ٍ,�P�I�&���GԺ��>�:��+冊_�/�n�*��t��t���5�P�l����Zk��WU�oA4�>_��a�_ �N����^i{n�	tlW?ݺ� �����!6��"��p��AY�Ad�y0���:���G�����z���\Ax�k�+�M�����jA� �:p� ��(�PO������$�W6��2W�8ʫ4���_�	H�'�L�!����/}�ߤY�t|p�׽#'lq-�������py`Z����n~xYh�)�z���P�{.{����d?굁��u`��	�(
��j��f�9Y��9�X2����vm!��ʩH38ys;D< �|�?
��C��2�������-�6L{iwU)n�~��7��l��k����������&3�Q���uf&�pL|����DF�d���g�<k)����ȧ�#10���C[]�Pj�~ɿf�E���]�%� F������^úl�<9����03F�Yf{�f.{o���3��:�X��������S&YM��?��C���.�d�+a��s�z!B��~�v{ö4F;T��
N�,���U�t=���
�N�.9�=��m�34:��XT�j������ˏsk0ڀ�����-����F�s�ً��%�֠�r�@d`U�dͲ�Q}��y���05�Y���)���w�������Rz���W$U���2��)�>��M��t*^����`f�ۓ[�-���T�h�Q�e��\�Ο�7�&�4Gk�`��%�lݳ���OPIه[�D@(�6ς�+c��d���N壟bM�.i��1�"~��vg/"�.@��m;AN� �Q\^��L�.�q0m,T�
�fzu0)��-OO��6c�Ό��F#𡯹?u�P,^�v��C
����}VO��j���p@�l̜�	�F��ec���p����/�d��J1��Լd��R{z�:�G���X��mҗZ�
���������K��Y�#��
�	$ME��w�O�8�u��o�,q����E�.�I���qb�Iَ빾�||������.�6�k %B] ���6���i}�Da-�А��A�X޼��F<��Ol��6f��K�l��k�l����Z�|������M�L��"�7-��B��>iN8%������{�s�Hbc-7g��S��Y�$I��up6��!,��&�a��-���N�	^9ͩ{Au�5.@�X�B�(.�b&��B�y�`��W�b1�Cql�՛��`��MvMA��ϵ����s9��5��׻�n�o��=,����dt
�R�<��)bv�W��^�:Hǻc ��{!�2B]+O܀H�w啔��\���A@�s�����K���p5��q57 ���Y�h�h���� Aϰ��i��_�|���W:�E���NX��_��2�.��]��?B������McbZ�{m>�ēh�a�,8ij
��+�:|�$:��=�<�:�~(��d�u7��ƻ�c���k+�����0�`�SuN�GhSݍ�e��਻l���e6*�}N�1(Ԡ�{m흱��1c�q<Z������AƲ�S�1�{���A���5��B���+�G�>�����b?1�^&��j��:P�a�A�8ͦt!�]M
���y�;d�W�����
�ˡ�	R��8�t�F��j�����;6��H2~�fg0
/�y�M�AgHh��)�|\>\�0W?]�`-v-����g�F�Nhos߬5nrF>t4�e�0���@ju���գ�6��n���t�'R�`���⬦������Q�v2#{+�)�)oEՋ}�--�Jv�E�����܂�`���>'��J�r�r��|�~0_ض��ƻI�C���|�0�$�@v�rV����E�����)��!�C���ۉ�@�n��A9#�tì�ؙˎm��7�h���⊗�ϥ�fW9τ}51���Ox��ǅ�Щ��B��GH�\�3B��LV�i�)�==���y��hY٦֥�F
*�\�Q�{U���+�i���{�	�花���\�׳����谨[�-�c=vjĶU�q����G�Ё��M�AV%W�隂��U�r��$�A��F/���%O5��e���|�B��@�Nk��U�\���BPh���Z^psݖώ�}fʒG�_)X�]��)�D�e?M
�4i:{���zp����e4��z˴h�!�
���n ��� ��ABNG\FdЯ����4��3<��q;���˲���w�AF]m�V�k��0�@S�l�X�%Le�����iL�zX��#�ȕz��K����y���C�*w��GR0�-��ţ΅�`RC�n[����$���+�lk�]��8��F��7��Is5���Y�wb�ˀ�s�z���ޚ@�F�6gK��M�O�K*�-�v�݌��-��v�}��]�{ǫ���;�����v�R�4�n�̘'�s�E���q�r��0���@Sh��z5ڏ�o����� �J�X�y�����v���/qÎu�܊:s;�͍�_1XH�g������F�3��2rVx���3��A� F�S���@�f�\�|�J�('�c���dl��L|]7�Lrɟd�5+Bh]-$0��`YL��u_�L\�I�M��F�޴ Â�i�?�-��������?��%F��g�{t��sE�+��4�;]
���w��}C������@�I�&D7,\1�m�%a��KHo�,�a �aR�R�[/a�V�s��%|x*Jn pڨ�%���R��ʳ���A �����邸����<'R%���F�b��BJ��iS�[)�Sάhk���wc��G��'R���;��rt�"��<��ь<�2��a�۔���8��eZi��P��U쐤8"�w�&b��?��U�To6�s��.�����Ne�	캺nGu��?�@a>���k%�q��CV��e��M�ǌ��]�g�ׯ�"��75�;���i eWkv ԟ	�U�Re�4���_][<�mTZJ�a���=�e�+�PX���S�֍'�so�/B(
���U]vt1��
}C��|T��Q�e1��Z�ppMV�Ɓ����O�)�D��	� ���FW3�
���#Kԑ<N�ĥ�!�I�-겊1���"o�5?"1,N`��F��On���
;#2����j�O��y��.Kp�F�I���QɖM�� @���g'S�cZ��+'J*��l�^C/˴O��D<:T ���]�+��u�[�M �n�"�Z-��-����?f��GW����#��#;)!@`�|�U���']*�%՘���J�?*�K?L�3Q��l����B[3
�Zk��D�Lv��j����VP����4�	7,Cޏ�T��un)�@�B��=��Ȏ_/@|,���dK�6��쇠�U�^�G��R�p�8�����^���Ą#A�]���G��4oM�ZUGB����g'�����]-�w��i⬔��z����e�-�o���9�f��2�χM����yO���9���普�\�Dֱ��͍5�5�sA������%��`��M,-O=}������l"��VG�$�2�67���+����� �@>vD\�O���9�/=��lĶ�)}�մ�x�����>r]�SS�z�b��F��o���5�x�ң5�ʎȚ�2N���6̰����:���8F'P|8C��1���] �΀#M�
��"�jQk`1Ͳ�D�6���%��OΞܴ��N�;m��p��χԉN&U��X�#?��M'{��Ap������n����
����8�E��mw��t�M��]���3`��cƗK:hm4�O�A"�M
w�[��A���&3CG��%O^���Xi#�g��(I�"�<����}�Ϳ�(l�B�����|�e��=#�Fl|�]
c3K�G�n���y�27t}�d�����p�V7F\�6��R�f�[gc�����E�뙍���ϛ��VP���AR)"���(�s�k��	=2A\�K��VN�^�ؖUD�����d���9�]���_�6��q�Dg�w�~ٚ"�T�q�D�� ���%�. 8̙z�;���^e��E��d+35{�~->�����h����˩� D�D�~ �����]��Ҽf��T̂Hh�'<'&��\�ew^kҚ'� ����� IN�55�[ӳ�e�`�.і��V�۬@X=�����,?C��<Jo`�~'�"D�����S�2(k�ƶ�遷�t�q�cO$�,�`��ܝ*����`�ls�bnEC��"'�M.m�|&�����TY<}4D��
UT�۰5
&���q^�1AB���?�����p?(�R[���`c���:m����DY�A�U��׆�^�ߚ�1qV_=5���8W�6S�c����ԸR�N�*�g�x�̾�	}�W kHk�1P4tt͒�q3�-{ 	��f���w|a�x7Un���|��oA�ȥ�F����I#��H=�1O{?���7��I�\=.<�?"���+.H��C�����m��4�Q�J�GA�(��1û�!�* p�J�k__�K�W�E�M=#��z��U�}<���i�<��%��J��6�r�,`��)��4���&$� � �7\M�C��I�%��f8B;�r�?����%���<��؀����J���`H]� ��%���4Ij�F��<r�v��r�֭ؑ��	X������ �%�6S@˅�#�DB�ɬ_�$��JY� O�/�5�����gr�.
���&���+�I[��фIÌ��r���|�i	�B�c��*��	�7n���w4�%jA�ei#.�V;����5��d�! kb
3�;�Y<�"ϱR�$�Gk�K�T�#[��c�U���O8�9	���]�6�؝���Uc"Q��XUL>���\�,u6c���-�S���n�RB����3tR�2G�h���R����9]�O�̑�)��ho^)Q�������]S�9��g�7�t����6��j�B� �q1��~/����㥲(B�kMD���Y]�(3�]"�̀?�aw���U�o�~���Ŭ�� ���B��Xk��+{��gW��-ײ?�����L:`_�g.���R[m N�n���b�7�t�x�=�I��86=��`��Mwa���v��_��vm����;B�5|&B[���6�=��n�15�V��B<B@�&Gn�����q�� l�Ks�&9[w���fy1{���2e��κE}�JJ��RX	�|�G��V�Z����[`�Ϭh��blLh���~����}���ݶD����<��p��O��3y%�é�SLN��L��=�*
����w���ˁgᵍ#�D�ݲ���&�?�7��1���W�_�Ө��0�"�_�u�7�en�5H�]Iβ�R��Y}��o	S����H�Z�C#� *V@��|U�J&�i���m���<hV=�[R��=�B�I��(�Rڃ
�՛�,4Hxl�M+^-iA=O��Oʬ��$#qj�nA�H/����ϗ0�q�e���v�����N3� ��Vj��5��t� ���mC���7,?a_���i��{^�1k�駡Λ:6*�`��qF�)��b�EsLl��>��K7Ȋ����SA����X��~�|�9�+q�@�g��%��O� ���������ev(��N3�Y�2�1*;�Ⱥ�a����A ����R�G��F��q -9	�l:ۈ��Q�<���~�-�DS��@o�b#��P�5�2�%n$�����8y�i�����1*��(|B}�2}��A:-��pk$~��Y��ɃQ�ξ�N�)m���v&CR�C�|��T�E\`�w��SIx��_�U�����y���NZ�����%�3���o��ah������SK���u���������ԝ�`�Py���ʮ3g]�h�n��JaOf�nNu�����'Y��(���O?!�`˲�6;��쮚 ��d�����VG�����&�@����SE�����*-��򡹑}{�a#��㿬+�'�61`z��Ӗ�+<݄�ʼ�L/�7^�@ju�
�j������D�nQ�HΆUd:��֢H�i�¶�v��p���e�*K�'�`Spж����%d+\�@�F��{v{3V�������p�I�l�T�T��-Si�k��qY��.콧a`!�����Q�a���=��ɺV����=��T��PX!�8�e�Ti7�0f�@[i�wI��`Ɨ[Z;���Ō`�}H���n�ܾ�^T�ŴR,l�&0)F��5^&m4�S����̸�7B�_��p)c��M~�3�
��0Чˆ�q���{y0����h��F�PH��m�P��;����,�VM��H̊� �Pv.-nD�|_W丵�|��w�^R|>��6��)̝��tq����?L�SOr9<k��&i7���ۏo0)�s�C����&��l�p~U��1��Ml!Zf�#�C6O����[�=b	�>�P3[�������H�dݶ�P8���$�����|��� ����K&�E�zimd�ȥr|'J 
��G*�v���>����l�8�O�>�Y�k�2��щ*���Q�g0�a�������b����̎3�Ö��!�e"?GyH�Sزw�
�gaM��M�{�z�!0���+M�v32�:M�2�*?�x��?-�l�*=6��iO�A.̀������j=Kܸ��{wȖx�L�-ЗP.���;����SV�[f�z��hD�ĵ8	�7$"-��.CZ�Cq}&���£���)25#.X���%���4 #tg�/K)O `�$���Rf/+�tL��C[��E���7�,0�5�ʦ�R�宭��	��A?"�>ن�b+���jO�U�Zr5�7��,��b;,�����	�VB��>뀏��d�-y/p�ɠ�΋�~�����NY.�v� ��E�_�os�=�Q��bS$lTCl����ڬ�N����k��(�;ȐJc�$D�;�7_�Aǌ,g7�D�n'6wp��[�8���!ө�=��G��_�8�.�z������ ��"����w#1��|Vy����Fw���J~H$�s���������g�\¡mxp���<R��kT�5�ޟ�d0�p������R���~���`��eT=����
��Zs�N��:���� 4]	���w-h� �i��2��7��o���Y���/>�����D�v��K��R�Ҷ�'�;��{Y f%A�v$uG<.��k��������UI�O8��v��N983*���`犰욽]6���K���e|s;1�dU&S�R�[��}���� ����˲�d�vu��dj��+����.!t�g�e��*sɹbDY��.�:�@ub%��le꩖8�S�uhU�圹������F5����_�'a��o�n�e5��V�,Y��&:n1�s�^�3p��&�:H�h`���%#�Z7�	�l'}G�;�Zoy#%�r��'���~�Z�6�!�S7�ry��[l+>�oX����͒v���+�(�u'�_x��,���ZAÄ�caX!�j���a�p�2v9��C:P�L��H��*�v�����������M;�C��S���w����6ZI/�G�Ƅl)�./�*8!�Ạ�d�Wt!PbE�Cmn�F��ݾ���%�E�Tq�)�cEBˬ0mE�샳pӷ����o����Pl�G��q���E��^uk��z]�	�m�Rt��-�w`���m������5_�*����R�<R-��oa?����8X#tj���D�K?@�����wԃQ�,����H�M����Ȭ#���ԣeۄ�Gk�u�"��B��o]��d��O�͘B�-Ъӥն3@5'p���p��$5"a_2�e�-=���g;��T18�v���J�
����u!��r,���6+��jba旟|,6����!��ﻻ�Hk����k6@���;���J$(��s��"*��L��r�5Ƕ%[�kj�^I��Yɯ�j4�%�P>C��g���`�B������!f�n F�X���VH�i�p%�:lp;��F9UW.�;k2�_��[H���yd�dqp�W>Z���v3�Èo&�e
��db��e w'>AvkV�7C(��J�����/ð�������fg�ZI�Dt7�Z����`�1TzƠ(��J�!$�q~W��(��_�+�u�:�Gƽ�nT�p.��M��3�E������؏n]=Y57E�W�=���+,�/�#(��Fӕғ��ԶG��p��<�� ��b�ٲ��P���1�S�s!k\ ��(Q�c�c�Lτ�����DC1`�|�K�P������e��o?j��Qҟ�B�b��i�_v\��z��:f��1���lx`"׮�!�!aP[��01�/`�^��4�f�r�Z�äie2�'�E�w��8�����Ͻ�jW-����~�Vr�b�{��k/��)f��[В�����]�i��j�S}�>b[Ԕ���s�	-�Ram
X���?�D��K1t(?b��D�`]F;�ei��!���%Aq�\Zqv�#��*8����'����ZD:�����j�������1��uTF�;G����s�)BNK`��H�j�
6�����Hl}����M�&Ђ���Qo.eG!��F5*���"C��]�/h�־N�&;�p�G��H�=84(�٥'e���!/�h����,2���9D/�0bSl�l[�F�<6V��+��%���A�%+׋����RJ{�l:E5��^�$WDG5C$��a�������:���f����%�g�����\�7����8����l5܏��I6�vF������ Tv���z�d�i�U�������T��������<��e�����\���e/��]X^�98E�
�T�g9���~��xB�N�7�䘱�K�c7Cc��Us؟pr�\W �e5��j�-���ҟ�L���h��r����+B��5�2��	$V@]f�=(ch��M��Te(^�o[��e��k����"�Q�31�;��v`aiQI	�R�C�4���O�s|	ލ�p�cv��QK���7㙼�D�����=~�b� v�xeZ/5�(Co�)+�,-�,p�ldQ��+��w�x�$}ėq>/ْƭ0�x��;��,�_x�~bSQ����G�p��ڥ#ɜ�n"�UQ��Y�3�h}$\`�=�������	m\�5A���|�d3ƒ^A¨�:��8}f��`{O�w!Ǎ�`Ibuɮ� �q,
4�UG|L��7N�3�2ad���J&����+[&+��(�)�~]�=s����b�>点'r�R�Ol��o���D�QE��L5l@��WP)�j��V��@L��]��2�#|�TW#�& �`E����3��e$�ైFXF4V��W'R��Q.���&%��U�.���;�)�W�����M��~i���2n�+`��~>w"��}�����mG�[!|8�Uf�a(j	�F�Ð'O{�ݧZ����dpR����!,Ѩ���Y&_�� Jw�Y����u�Pxy���[u;Dg�}S���Ѹ�@(b������:74CDO�!$f�ǩE�(��_�<{¶�Z4�x��xj���8�bZ�q8"�Ŵ�E]�������N�.)�z�ֿ_5|T�q�r���@(�*��$-HM�p�&T5thI��||����MS2 e�q}?�
X˹AA`����|\���$�����-��Cru��!t��.�?1?3�i�L �uQ����kmb3���]���JeEF������%�U���S����OQg8����~!���;ږm���:�le��-H5��ˊ�����2i%������4��84�f�Z��N�!�#�����ޫ`����)fBd�m�me�n>�h�u��f-VeXW_��Y���ԁX��W.a�6��"�a��k��>���pДX��v�Zq���(��!p��|9�����>K�ylƏw D�|�}d`�yOM7'�6F�I�О��	��фzc��v�Y�MUV��$�,H�O�#fm�h�����i�J?e��:#S�[�������F�b���wK�=ϵ�`Yk]��$����[�3�݀�M��!�5�����t�L��W <Rx��?!m��*|��ڰ]]8Ӌ`�[���,��:Q�{+?I��A�����2��)�R��ņ��>a��D�g��Xx��A��7e 09�Z��;Ʈr't���0#���Z5�g-ߓ`�t�^�`��9��v��ԍ�lj��etZ�5���q�JQ�QWR�⋣����L�_Z�r%]�z�;b+�� ����Ն4�/�����]"�mv�c�	��<2(�E9��T��M��+Ơ��{��b˜�B[�J���{{o �=�N`A����-"Pl�c�����5�8�g'XV�S���%�.�0���^F���GTӱ$
���³��GUh��B�G�M� J�_��7MID�Y1P<A��D"���F�UE�(yz6C1U#к���s1��搒գ�j��k�� z���*H�PٛT��a�>�m�D�q����ߥce3R�[G�	�;b��&���	FT:�h��J2pi���9���I�#�-��p�sᨊxw����>E?��rR�A/��_}h;y�V�s]ع�:�%���dN�r�N�nו���c; ���O؍��[A�o�>��S!ߢ���.�=�om�RY�8��\���H�#� ��P̻hd��n2Rŋ����A�s��'t���U Թ����r�2X���\�I�'�l{�5Y�2���>�)�c�ߺTjzM��@�<�Wb�<V�)�Z�-�Y%�sdt�X;�2�0�@{T���ns��LB/dU.��;?�x��h�.k�$% �F�%�ǰ���(�cr�����Q�·MUѶ9��X�t�r�$xoA�S}�6"ӡ�P��m)�X;�|�ߏG,�d�k=��}]uc�-N�cȡ\���]���~i��ɉ�t�N;II�!Vճ}��Ǝ�o�ߴ��޶MVP�/��o��v�L4�9o�KCI2�{$
L։�ht@�s��@_�\���1��W�4����SO� �v�cѶTݴ8�h���E��(_����b=M4^0��)̮�&�S���ے��_KFPɲKHmD����)�����:9`n��{v;s>�"d�I�A�Ut�������Q�Vl�9c�P��*�J0"}�<��n�kƿ��?�ݍ(f�B����c�tN��r��_��*.,k���M�0�Q���d�Q��2#�0��hU��j��Q2
��rH"�V��#�Fe������th�Ly��fy =�F�a�8��C�ݲ������H@�R������Q[�iv�������t�M6��+idE!x9}�f`d��
21Y0������⯠1V��:#������eKkt���Њ30��t:���*�C����g-&5�f�ȝ����6e��]��]_v�JyMzo6�5@��Z��Fх�_�N�3��U���5R��)=vk��ZYÓ ���JfC�~k�k���\�tˢ�b�	=||?L��A�j�q\���bF��"�rƀ��l�L<��Nd�x/N⥫J�D�%�?ހ�{P�գ,*�A6H 6��G�C�2���Z�߷I�7c�!�[���,焛γ�?��C� ��y}���mt!	|x�ō�X_���ylc��=X�4#�h�A~��s�G�Z<q|3F���?KRRH;#�M��#�k-��vS~�'
���C�ъ�LG�\?�%+QT��f��)��i���c�����^F>Ǧt�Mq���Q��ٿ����#g�����h�&[��잃��7�>Vl�]O�)���&Q������ vl�:��<ez�fM���x��?wLɿ�E5�!;��Z<�T��7��K���KtS�H�BKL����q�y��e��$&G�y>o4CVP�Y˭��ο��v���Sd�ʼ�C�ph�p���Gj�Mm�w_ߢ��[���s$+�?~j8���"����^a7�^��E��+ĺџZ�y���t�*��57����4� �m��.��͚�56�H�����ɲ_����X)�iU��4����U�z}x�5�ŕ�V�GD'�y���b�\A�!�e�x����;���aҁ���VA��4i��āu�1;[�u��($�Ѐ���8��$a���wX�(��>,�z�N���M���l^�JΨ1��?\ � ��}?� ��_�k����"�0�TK-��2��	;�<��[;��%�6����SOG�B(I�S[^��ݖ�s��շUKo��#|Q���!#��k
:|�.i8���� �G�����QV���0d<0��U��;�"%lǝ��I��U�>�<w�\�똬�F��UBd�迟}����D�X�x�P�ϱe%�.՝9���Pu��
���\_^����4ō�zEFG��v��J�V̔>�3�����k�J���@#Fק�W�
3KGof^�$ȝV��`�WCoZ�Y�8Bw�x�T���Ky�/Ve��Z��F�A�kN�q9�A�a��5lmm���<^��~�-|���#�X�v�h_'_�G$GGCΪg����C�[�1�\D(��7kP�G��~B�Up�G�%w��i�+#�M������e��6+A�*�d�.����N�I?�8JR+ p��B��gQ�ZG�����4AX3��x���m[��]l�.*a�".��]j�K}�0X1�-����r0�P�t��r�%:lz���{�6�1�M�@&.�:@=w֡+�l�[��%�,1��y���$*��U,\�zd�RmZ��4C �j ���Z���钭���ڶ���i�n�%�~`��ϴSai[��F:zQ*� ��xE�BU$ı5��;@�­�B�U��W`�����H9$�iL,��`Ͳ��� ��]�K��"��s@��ߘ�
���Q/U�q���.�_��9�:������I/����j�����bwo���R��%g�+O#��(�a/�~ Z��j(��~]��x�]�j�w|-"fv��Q$�(ݾn��%h�/?����Ľ1�ØVGu�ԢṎ	��0X��K��`>#<��HQ/�@�z�����ʹ���PH�)�� :��P���o��$s����ˎ�}��ɲgͬ�@[7�PM��)���$���>�,A���c6�B�P-S4�>鑙�~�����Lv�@}<��2��GN������5B�K�2�"��}�4c�0"�B���A$y�U�h�銸��4��[����z-{^3��*��q�q��jp���0� ��8^9�,;�=ʂx&)��n\�5_�xU}��f��A�����+�arS�ܦ]��S�9�u)�{P-�2�i��V�ƀ��G�r�W�7��%�_�/��ϝ�?Å�����n�!�h�ջ�i@�ǕV����^�dDU=W�s��L�)'� d#�/m M�ڙ3�/0:�Fܱ&1s<�%�1�
�*�D��u�ê��þ< �L��kvp}��mu�M��t��;�f�Zdw�� ����l�m*CƦԟVx�K]5a�K��&��p��i���)�Mz���՚��7$� 2��u]Z�24o��CU�i-J������e:���?ο߫�Zz�
�G�c��%e�M�NEԐ����j�(�&��I�C&{���K.����.c^�0������C�P
"��s�ka�k�9�kUE�8���vdx\ �`�Mf��>�i�XS7E��,i�~��zyhv�;����.�k��mIG���S5��Vn���B��NarX�f��0qO֓#~?��)�T[lE4Y}�0Z���Z�|RRP+f��	.-�܋�Ř�LC��Y��q��2b�@(� [fz �g`.Zp�gu���f��8������ٚ��ͽq<��5�ѩ�\2T*O�2z���� w�ȼ�7�1���jT�f��>�	�Y�yF��Y�ۈ�����M��!G��y}uo��hۜ�7�x���Y{�Qb]X��G�3(쩟���G ~Y��5͢�] ��6K7�l�V���8�^��z�5����l���C?z�ٺ8bJ� �+�S6}��=�)	�zW���?�a�Y҉>r��|�ԑ]��U���;q�~�J�$պ*�C(���W+�4	>���B�� r=�I�5�	w���ve-�* z���@�T�Է���&ܠp*,�]K�D���D�����{�;&���	����A�~	X���	���s!y0�]̦҇O*Gf�+�[b*�q8'�&��d6��9|��O?�e�`^M����"�^�?�	7U[�Y��0�3ugsm7�͞�\ ���)�pZ.��Փ*Z.T2�&VLQ
,����l�M�)�AˌG���AM(�o3i�-���H� �`A�S�3a�.�]ぼnơ��2��@I�O�·-�v:�N�
l���lܡ6��c���z�}٨�D�淚��P����Ϻ���!S'^Rg/ҏ��Γ�iI�|������� P��hy{�~	����J��e}M�����`w*j��|��9;��_}�8�Tl\�
#������Q$�g�P����Q�8;�c ��DXt�O�g�:肵i���F"�-�����+<�5��r�"� �홄�!%�l��ϝ�N��ѡ׳LL3v����D����s(w�)�>,�ɡ��ͣ+Wl��Ǚ�n�)E�M�����Ү�4B�)����B����m0�YN�JRt,UR�,����#|�]1}����b�p �����L���])z�5A��j 遡F��R�y�־���qt�cU��B.���lN�{��o��z*5�Q��e�W���x\VB�~�9��ַx�F�PE�P��P��jV������:Ha�J_�o�t]^Q9�|2�a�/~!�8�T���L���t�?3�n�w��YT:����zMi���$w�O�-����� g�	*��)PgL��$�uC**�+ ��~�#X�����@D��E��#���0M-3�F�����^��E%�I�����ޘBfXe�h�
oX�"g���^���<�0xv �ѐH>�$��k�y:��I`�S]�g䛛hv�1���נ��Kq9��Gk/sl
=o���,��8��0.C�l��=:�#�.\7
2��Ѷ��
�������,b! ���ʋ;�b#1n�f�B��6=ˮ\Z?��v�2L%���V�^]����r�9�E�j#'t��hY��\!��{�@�?-s�ˈyf:t$�<��Jw����v�A���V�4(Fu,	(g���z�|�?7)/G6���"]Yt��sI�BT�b�gw�g/�05�K)!�g�"��XC,S~��������#B/d��������x>�y�W����:�"��-���`�)�IxV�r"����U�g�b"��0�P�+r;��\\nj����w����PL�{�֎�>�-i��^���iA2~�L�'�=�����k��Y������Œe���]����V˖0:�YX�Y��T�E=���+F�d��}��ٌ�߃�l�ǽ��`���O�IG�e#�N���̲���7��0��(�ox�ғ���1!mxW�˝)��iv��`�����	�Tx|��o3g,+��5=����U��`�L����w�<���3���"9�C�ͬ��Z��(|9?\�ە��M��#�,LO�[���o�1�p��=�!@�n�R��.�ʰ:�M�J���㥽����󫖮��٪(ٲЋ�����P蒜=�w���O+}�)��Ϟj!�MP�
�<��UbF��]5# ����y�헄��H�q$�7�m�l��t�Ҁ�O.�1j�����@�u�z~t��>�t���Zh<;�k�R\ܗ)�JE�&�}lT�$K�,�p�"l�R+��ڻ���Mo��K4/�A�PB�|��`��*��AC���u_~�W�?sR��q���o)CXs��]ڸ����k_ҝ^�pm��|�ˁS���	�Y}ǎf��8�tn�D�r�$���_�qH��h���A�BSÙ��zO��0`r��N?�<�\.s��_[��1�%0��eީ;�	���������G��&�D͏�>��H�[�( �-��e"�
 6���kJPd.�\����쮋� r���c[Ǩ_��0CH\�]�`PD��_Է��:��,WF���!zx�)�=�.� ;6-����n���	0��x�(��m��eF�Κ>H�@aK�@R����5	^�*�my6-�s� �Ŕ�{1��a��������Tл��si��o.�����J��|D_�[�T?�T�\օ���Q��r#4��W����T��	Z��s�V�	l �2�M�'WF}4��y�߳�Wil��ϹG����m��T���鶩	���Ǚ[^x�1W�Z��"Y�n�G\��
5ÈJ͆r�%�����ga��d�	*�j���^�oʠ�]�R�U���{��������l�0%��V�H�|^�<c���CsG���v0��}��h�����S�W�~�F��O�v?ɡ��0��#�-_�������0u��4O"�oT�4J�J�0܃����D"�~������0�Q��G�p��/h�Le�:�{�r��řP����Au�?�]a֦���l��%�t��0���L�����*������b���e�j�Q�:�}Hi���FN1�k6aWX�����+P��X�Ip�`߀�e��K�'_��akKt���~��q6�����8���f�Ye;]�- 1�dO���@ͻ�H���2�	q�v����}���h6>| �7�	��ж��l�D\u!k��H�����_�^'��Жcr-0�FIzWB&��ȿ�Ƶiw�Z��N���k������q=O32Ϥ�SUB��J��1����f�&�����(�>��(�z��̬ʇN�ތ��|A��$��G������?[�O���m�Iaaf�������I"41��'Zg]�j�&-s���43z��9�5�Z�'��9d6�o������`�>�#a���V�+l�$�0������c�"�� 7�_Q�'-~�*_�A9��1�A�Uaes�(��5@�hX�g��	��ė;
h��UB0Z��[<�."ӛ�b�Cb%?�3�Й
���{��}��'���'�����������ҏx��R_2O^9�,��҇��]#�&��Ξ�Gm����?�s�A P�ҁ�r[aP�k?	uj�Gj7A�)Gb)�G�^d�3�� +gqfC@=�*�+m��+@��I��z�[H����6��Բm�n�W�ժ���F8�Y6�yCmI�lY���]��tߏ�6��M�3�?�,�{&���ؕ��(��"��R�ޜ��@ y'A`$���C��Y��p!��.��#���>w�!�����?�7.c�����;���(�ȕ�[��@OS�1A�;d:�`���O_v�'��V����F\��R�Q������0#>��f��7��S���X��];}X��f��J]j|ŵF-1�ZAbC�+�
�������+����^/ӕV���\��Y>�c'���/����G��=a��3#��з"Ә�&�>ۯ����%�i�^�0F�䅮�|m���X��%�����dh]w��¹��?S
 e	$�zg[A�����|��_ھ��}�|D�U�e!Ej �w7�Iwl�&{��~n��h_��u��V��ÔYhq�LWD�.B9�:Ӓ�8c�!�Y��`ׇl�D@�H�e9Gtm���eb3bW�,��e�����ْr���3MI�7��NG�B��2��6e��)��A#ѽ��2�BU�*3�Y��H~��SY�(a2c�c_��"Q�K�ť���Q���S����
���®����G`z3�[��� v�~y�)/��;�S��5�ĳ�ԗ7Y�`�X����)8�b�"r�ePw,�N�Pn��@JT��BD��CI=9K�����WNH���2���O�<Ÿi��o���A��or.!����$I3Q	1�YB��X��ی��׆&d
�(_��M����j��=uI@�1b%i����N<�y�k�k�]u{���%� �T2�C� tr���w��#I88�'9L���;�����H8'�1��X2I�>b��B�𫜎 ��dE�[M�P���5[_�����_Q�sX\�t���E6t�����hӺ�%j�2r����x��~oT�I���7|����:�6�T����2���w�%_ K|�����	L]���x��+lYc͂����ÿ
w�}i^p��ߩk^�:9m��}�8@º(�N�A�;��ل��v��(�	αm�{±,^���ޫ��-9�@u2ƒ�nc�GF�v�S7��9����v��^Իd٥!��$���t6ٕV�޳6�m@Q����h�E��>!Gլgc]{���?s�s[o�9?10f�R5�Jo��4��+���{��]V28br���Z��� d�\"�N�ބ<rpW6��@m�����&{p�~��P�I�[�u
��VhmCe��(4�����X�n:�-��M�����&;]�{2^F����[B_���?�R1��w��Oe�5�pw8J�u5�#�dǥ���I	�FO|��p+���y��zA:;A�&m�B�=î�k��l�z�t�P��6BY�����/q���L�d��n�ɬ_-�z����)�求�C�`.�gM�CefFǶ��+�-��3��Ą�-��	Т�C�Ԥ�g��+����t�!�y��h=�=��r���Z~�\�*�Y"J�.��du+���+RC�$,�#<���z�S�N�w�a�2zm�cv�z�$%��5�-k��sZ�%�:GwNо��뾱��9�"���Q�O]0j=SEl��v��
���^�˿7�#��F�`ZТ2� �Yj+:���7*��(>U�^� .��$���,
׋�,^���B:�[�P^P�W�u��{MHWY�l�6?�+gu���34�?R{>#(�ܷ�����F�������Nُ̼�qL΢�{��;ծ��l1Xv��u��y�%���"�H�&��}�|�)Ɲ��/�s���C��"	�j��$7�w�s����h�i|D"Q1v��`c"�T2׏�<|�<+n�d#i��weYv�U�qXprM�r�Zڳ�_�RnAl.�ud� �QgCK�o�&�QKY�� �tm4Mm�����e�/��&f؍�_&��Z(a�ㅶ��FC''�T������N���ͧ����P�~O��w����i�'�����8�m�V����1:\/{r*�4�W�QjM�CC?��*ꍗ����o`��pz���M�͌�(R^"l��x��� �dyOA�X	Q�@6bi������@�W+O�ek����˾s�ݿ����z]��X1�B�/C�zy0#E2Q1��eH�|���;�4����ᮡb�����67����̇�a����V%�Y��Z(Ҍ�L�0��K�m!�^|��)��X�x���@ ��aFN��{[Ӣ�+�͔��(�I� ��m܏
m����u�%�(����_�W �S�\��|�|���L��:��{��v���<� ���?s~Bڱj�1�D��<
� �G�In$OS��v���I.� !�Ԣ���H�H;�:4Z�$�X�E+jI�!��ix
���ƾ�%q�KbpƦ��֘�,?͛k?G[oG�l������d��Ae�71'W����s���QA}x
+�w��ν47�w\��A)m=�XWzB�z���B|7����ewp%�e��ZX���,�&�+���`r0�:��4"{	��7�/� ��]=\����`:A*=q���u�Gb�LFz�ϯ?x{���{"me�%�Y���B9���O��_�~�F�G 'N�vw���^1⾉t�G|09 YL����T�k\N��HM���܀e��X�v�2���$w/�M��2޳��N��~����ƽ4Q8����U^������'��r/VM�>�磪����3�4OQ�p�� "
R]W�@Ɋ���#P�]O�f�t���	�P�; 	|� ��LC�6���j�t�Dލ�F��1���2Z,H�B�=$�E]2��G1$�̦��S}�F��v=�6]p�4N�\u'6�km��P*��Q�!�j͇8_���nq�l�YRA�ȗ�b�E�W��.L�]�~l�����0Z���K��a�s�fl�4�@#�;b�Bϳ�K�Q	�~ya��5�6��𗯔y�����`��^�]���|G��.C�(�1�|���kx�k"��\U@c 	�vmj3�c���*��.�2�©�P'�Nx�P��2{E�ȕ�^��-WF�ĵ��_"W���M�'HSȫg;i�[=�e���7�#L� p�ә
y��$Ezb��3d�5h/8�E(�/U������y5O�L��@޳:����4�P���_�,�*��(�*g��֗u�Əl���0�#cr���)�ι�_*�I��>�F��s���ia�%������-z~P �<1ɂ�ڬI�0g:��i+�B,���
�:
�	������~��u�� ��r�2��@D�5�{P��c+���H'J�}bQ�&�4Z��,t���*��g:͆d���������py�P.��ʲ����+�/N��z0�&V:phx-��뿸|&]�N��?�sK}r��$��@� P� /�f4gE�f" ���jFh>�$F� -�+�X��K�W�bh8��Z�q���as[�oE�����_t����[��Tو�m�������w�z&@j��J�r��.�hh!܌!���T!܌H�9�xwT"��4��� 8Dꛃ�>�p��7��u�txB�@��VSiwlW\|�� �\��q���W[��8tfbo����@��(1���#��@a�0T��7!�GP������`�*��q\Y�/��;����ܦ����7�M{���g�Hg��z����5T���Y�SV=sa-Sx�dK����^W�r��*�EY��`�q��"#�!���s|t��Fǫp1Ě�)u7s��;I��]��y߂�m��H��@��.�@��4"���0rp*<�ߞw���p��mR=��~�w��ĳ��c���՛�K�F:,f"$h��E��Ҡ�p�����a�N�V�0����|��#w�N��2#�}���j����,`����&�[��R>�������a����^#i/�U¼�8���d��^t�H��Tq�:Kk_/a���'ݾ�n������.�P�����Z�����j	a���_>Q��7@-YHȓq��	HR�X��K�N�B�;]	�'� B�w��{��	����z���t�V��q>��t�t��� N$�˷q��xy�vz�O�d՟@6B;��;��C\0���w�Uo�!��筋�@�+��=	�_}Je��*�۲j���̒�(%� ^y�ys������i!�M�.;k�5�!K����H!�DRh��6�h���1�=\��Y������/	�dI�Ĳ_菱��j���ͻ,R}7�����Ta$�^w���˷���u�gK�~t�� h�F�~�h4�|�$
t	�X�$�i��0���.�0/� �5\c���4��&It��WN�]9�A�GBo�f��Hd������[�^1^`���ї����c9�t��~ q��::G�]�F��QÞL��Ʉbº0�������h�u�tz��8�"d�C3K���� �(�%��@_�G�E�ݥ�V�*[Z�E�C|#��V�L$���e��%�׈��Kѷ�����#=M�Y��rb��$�z�nYPSSJ�����DP�5�6���pڽ5�&~g�<���(+��'��O�eP����� �T�;-��ѬL~���jzyW��7�����UF܄�@�Ռ��'T{�.�����Ѯxg��i�w/ ��8 �8x�t5���[t�q��U�|b����7���P��ZuZ�ZԨ�%u�nun�Ah��u��W��(]��Ke�����:q�y���S�F��
�oy��N��G�j5�hy����m���>*ͦ�3�揅�v��aS��s
���s��g5�v�����/�-2��o�C�����~vt��pQ7A $����
"En�}�n�L���5�L��*_���?
-���)������wN��=�.	�<�o�OR7�Cզ��M�&��J&A���p�N�Dz�_ ��^>�Y�Q��"����2,��H1��$�?�1�ɚ�.Ki��`7E>��Ժ�,Ss����m������������/�{%s�¼���(}��Xq���د`F�^�Ϟ�,��l��ϗ�>=#�}��l�b��Ԋ� ����Cj��؅�N&^�H�L�I��\�2��}����-2���u���`�Z�d��pt _xK����H8��c��"�@U�GW 2�=����'��Z�p�oQ"0jG�8;��Wӏ�չ�"���M�V�Y�>��Qx���ξ��|����l@&C ʞ``@�Sr��>�E�f�5Np^'�mp[Dz�W@�_�jV�sX!QP� Kw�J�5�#�	rQ�<C��B}� a��	&VM��|�����1kB�:��n99�R2�0�K��L#�ە�T�q!�k4*��B���Nt�^hN�1�*��J�D�F
��՞����E�0U~�ϯmq_�D���T���M��_���P��>-��O��q��.�2�.Ϸ!x0�����y:�&���c�#NƬ��f�D���VжΎ���잓2ҿ%�"h&BSA�$V�n��tCH3�澧��ުC�r��9u�[�l�f��c,�hj,*H�����<I���%��fôӷ�'���O�ɹ*V��}	p6�2�N�� ����	y]�o��6V�_n�4�Z6��� n�P���(^04�_����gdV�?z9ۈe�o����ٞU�<���_ue���-��Vn��}�	@�X�-��Pc�P)[��F��285�C <_v��as)�P]~Fڍu^�r��u���B�f�o`�kZ<��5mw��`�Jp���E?���*k_S( ��4�9���o1�@04J�0u�#ƨR�Ȧ�dFds�d���Y�e�&vY��9r/gΉ�T��>�_m��x,��=N�9������^�����*��ء�R��h�'͆l_���f'��u�1Վ?��Q(e�x�;���/��Xi*��� (�����	���J�E78.-Z;h^�P��B���~0�n�]WZ�k��eå�m�r�Y�h���X�Т��%��j8��ٔ�)�c�2����>�4��?��$2�W�����m���%e@]|��ʫi�~
.Bl��-�?6X���E�$��>d�������|�V��m�E�;/~ʂ��&�'��^�2$ȬF��ӍK�Y<�cuE-��,P3�Hg�F���ހ:�K/�ǩp����J���`���Q0�P�i���N��Hi�-H(�t�7�϶k�7<E"̔nu�<_]��_� ��*�Q q��ϗ[��O��,!�W%e�x��w�2�`�Q��<�0e80�3�s�BwZR�r <3l-y+�8���N�QF`׎�i<iU���@c�0� ��d�����9$^B��1�ek�y�=�����X�������}���dr����l���#v[���آMX�A�C@��F/n�z�m�#��ǕK-r�H\�K����R@�����0�".����0��~c��G$duty���L1׼�W��˘��M?��*N�0�o����0�L��T٪9������{ u��o����2���$�N�;T�'.(r�̮BT&8��r���*B/�Y��CI{�QB�eN
f�Jr�HdH��5RS��	��^�����9I����N�V<���;�|����`�����aA>�$���
�����#������M~�I�$B�7t$���mB_
"�[<��H�uϗg�9,\����O$�<ܖ�̎bvb�/��ŀB�ቅ��}-E,"�*��)�R8��̹v���6�ԏ@8�,�83ZJ���vg4��:��ԡ`���A�4���ؕ`)�(���5��2���͍4f:y�P]p��
�?ˊ���	]e w���sl�m�f8�|�3�������V�6Om�ffȰ�T�3�+�mS��1��'uKY;`�Y9湈��/�<��u%�h�t�f�(���M�i��ĥ}+�@���6�֕���G�5�S�F��q�q���%DOl��/�o�J)���*�;ҮM�hl �4��X���k����c(y��\f�ܷ���f�"�{�b���B��V���B��T���`"���Y�Փޟ +
�h�Q.C�p'� �⚂�²��++$�jo~.���E���t/���"A�`�d�9�r	y"YO��c��;��n�'���Kh0� H�R�BX���_��R�2�7�;�f���#�i<��?�_>�$��I���x��6Ƌn,�g������bwloq�^�3Q��rơl��D�����S-})��C
��(О���?\k䔮�
��颼�v��^d,�?��M;dI3�^�\q+]gs
�zoC>彜��Qvm�����]��˹�Ws����u��Q�x$M�E��{���~0O,�|,�t���w$�q�W�;?JאC<�/�؅[�}V+b���a���)��ѳؤ8�(w�.�����B����-�dLZ��J=���[�\(��C�V��)��d���Ui;����B>*^������O��K,���)�D�,�{�� ���+a�է|_jj��m�m*��&
�9��$i��é�	w��۵n�%U��\��)���;�=eݡ)`��� �|D�
6,�����+�t�~�o��t���l��e6�x�Y����	ٯ�A#̿�j�ª���h7Q�=��@���V����C[#�igs�t���Z�9Qf�a�JU��
����UD2 ��Q��GBt��Q�F��QW�6*$��^N��H�>W�xJdj���oݍ�Z	?}{��$��W�J_�բHe�6o<���?�Q����@��K�FE ���.�r<�v�bhb��k�v�3�O���7���υ�I�{*6# !	��ƫ�
z�NM�?h0�y�q��dm�F��L'Wu6��;�ڳ�'O�OaA�!�]�qX�ۻp�ך�Ց���Υ��O|_`%H�c��'��R��Q�� O�(�t�����W$ž����lǒJՈ%?�.��g��3��L��H�ID"S��r	sc��� ���2~
��*��ro�X���x5	&�p���qk�C��J5��A�W6���V�M���H�i#�ڏp�=<�d��I��2$���SWu���Ċ@Ǵo>q�B'�8C2�,��8�sW�0�����"{�����/߉z/$B�?�E����ÆQ Ke�}<�2|��Zo?EUZ��?��9:�k4��K4�Nې'/�zS��<���(,1�M~J*�F(i�,]әU�rsC���>�'��Y3�BՋn�|uc%\���EL!�8,\䆁�H?�U�9R{7h���'%J؈TnI���kv�O5@���5/ZZ�L�\����V��	p8�`�A�?Cԇ��Mr`�RE�/o��P"��X�񡝐>�IQpa�6r��J��s���7��n��P�����;-�� ����4OL�o>:ޝ�F�61<&O	Z�HǳB��p7�J`���}��Lg;�>�+�N�_��{o�Z�������0��!��õJȯ�eC�L�M숔sIo��k]�h���hFb��G�`���Op?͊�
��4) ��嗞Z'{��ϛ��A��	�ș?1����8+wGz����;f�j������)�̹O�m����H\�I��5>7r�H&N�I6���쏪��@Hۿ��(�^5��M�dL�i��%�\O!y��?R$WW�h��;ܐ�𶅭�W�~K4�jg�g�Զ���n<`���p��EǄx�Xف��ŝ	�Yc
�A��K ڬ�;x\�1�sX$Ո�Ʀ]2�&��1��9��{�_Һ��(і�7�g;v��5�x-]\�O�_����YdQ�ozӥ���p�+�	Ȗ��~4�����S�W�_�;h�sO O({9ŸLa*���k��!0D7���p�ꁷ��,C�k���p��ڨ �4��kc(�0fk�r�Rt(2aY^6j��	z���[6� ˑ���L9 �g~p\ ��gN��H�S.������}Z$��v^*@z���'����x�B�>v f8!Ũ9�-�K[x��
y��j�-��&u.���a`��S����������%]A���8Wx/�jGuZ��O1���,�J!Χ5�"�w˃eg��E�LԱKw�����Vq��D�܆�o�5��*�4�h� �΁Ӿq�*����Tv�?A~�9EC�}����b�2�����1�	}��>�S?5�^����~���Am�Y�a�]�8U�
��|��,�f����/W���b���w6�V��cSS����s[��p\�S�+�����[���'��|�5�Iow���yy:�70�Dc���B�'�AN�Tp"���$Xl�"��R�����?"���@a���_�N��B��za8�i������:���gݵs7����OdtѹaM��$�B��5_RC������������\����7��ƣ���ٳ���4 J�)�ۼ�3�;��M���S��JdП4&J�y�W���c��/]�x2p���tn�cdw�3��&�=��!e*��<�%����zY<qL��D��W����n��<�� ����ObV�<qUV�1��%k�7��/Z(G�ڬ"��]�d���ɛ(�A5�������6,$�un��D�"�ن������JF7�$֧�_; ��om��LY�:U�Y��N& �))�/��n���G[�O@7����e�%��t?�5�ü��F�~�̸���1^�����@Nt��؅c��������{4�|w��f��x��\��ɲ�?��E[KÑ�/N[�2�aCF�,t�c[Q�׃p��Cb��\��v��'O�W!j��u��N6	U��N���h����Oݛ8Yy�w'�
�}���h%��������P5�m��۬p'ݑX
��%��P��<d��Zߜxa%}�X���3�#�}D ;|����
��mI��a��K�KW[��_����d�`�$ah(�M:y+��gR;*�/���+Qe���r���v&��41�_t�d�0��E��|� 	TF������w��$�߄2��� ��D��䁡��,��NO7HtXƔ�w���|>w3�H�nVO��o��j�#&R�g����4��d�����&��}n{%����y�OA�����5K�K~�(R��&��n�ۓ��`� ;��p��f��}�ٞDB���@(��T�:Ͽ:9�(��t�B�r1E�M�<"I���+D+PZC�\��L�|��RWb���V�����>rM�YM���W��vXvBR:�ަԍ�$��a)�Xz^ځh�	`4 ��'�5�·
�U6�Mk~�7ⴱH{�Ϝvw���ɩ6��mC�� ��7XY�(�����A�aVnV�������oԉډ]����޳2�Hf>����(�n�#)`�ENko�=)�����9�uHM�5譝3x���E�3_<��0��>4=�V1�-0%$r�b�~\z�R��s�$��S��6AB�Q�y�U�1�zfN`�L��k1܉o�p����sÓ�o�F���r��R���-k[�x��0��.s��ޗ|.R�M����;�?{6�#L�Y�h�c���!���<Oq[F�<�~A/q�x��/a����1��7�l�4@gfvptn����)ǚ��n�el��K�a�d�q��s#G��m*b�=�Ν�Zui���]|�Ħ�t,�5o�?Ii�tA��~%����+������\�HԷz�e��<�q��������b2�d<���J�e�>;&(���&��t���Q8��,�D�l[��w�7l�E�cߢ�G��E	~Y��(�� �u}���]8gu4�we/${ʫI�h(��������~�����kN+�8�_�x]eP���=-��T��QS�z����t:k��7Kw�b�<���Ԫ�In��Ql�sّ��Qtx\���>F��-{�����`ο"7�-��7�k,Q�;-=��^2�eյ��"��6JKaO���dR��I53��z�hrk��ۦ�{�I����V�-1�� 1W>[+E~��}����Ѭ`no�./X�8���?�\ퟠ&"D{{�M� �Qb�B�^����v�����o>�X�sps�W�h��}�Qe���$ʖ}\ʭ���E����;�ә7� �;��n�Ӿ����	�Z�������=�|j	���I�t�B�nj����Kn��;e��֠�� ��V"��e��$��ʦ���E0���)��� ��7x�~т�2:̜Ɣ0_f�F<o�,��bƿ��'��6���%\���B����헄⦦�V�CHw���A��}v�~��������YJ�@@N���a}�x�$0CCFQm�B}�-Z��2�SuO����V��yQOY3�Ŧ�.=]]L��9'7^f�����Ah���E
�!z,�=�Vc�T5�Q�P�!�s;l�*��L3��|��H�K9:I��� �����Ha�I�����r?fy�{V�P>u<�OPU��ʋ��g������0)���MW�m�����:%}��1�/�-q��:ٜ�����ui�����S�b� L��.8��:)r��HJS�*0'�O`h(�tMY��.�'�L��=���`���i���EI}2�2��	��Erڽ��G�k�T����@0�I�4��!�I*|���:m��W�=F�IYQ�#��-d�G���E����N����2H͚y<HK-Xltvt����$���h��Q�l7�������"�#z+%�ɓ57à0�w�gƸ��H� $����~�P0���@W�'	�?Bh���`�CWL
�1gj��#Qn���L�g?�n 1���P�$!2.�U'-�k5�Zy��Q��D��0r��Ĝj�hrV��!�.!#|�� 2񽿂��
8�b]OMK�_Lz�}�)oe>�����,~�.�@�\'t��j�jK��rw�(��a��#�A�e�U�8���m�K�����?+���E��D���$��ҭac傊����$�ճ���̤���S�����4�6�m���d�s��(ޗ��\WX*�ST��zPG̣]��I{K�$�O��Y;׺��v����%�2����*�W�{�?����卹0a�%�)�A]@��	�.�#�,��xG�A
As��hؐ�$�ʀ;���{r0%����+�^3jl�����6â�w^�p��ʍ�B�v᠙$f��� {�r$y�K!��2��.���B�3��ʅ�S��/�'�"�;�Bt�`�d�êt�*���ae@\��&b�Qy�u��~w̯?3n�N�:{�,_�;w�"h�c0E�J���K7{�D��.ɑ���\�PG����t�B4L��!h�;�H���9��6/#<�ߩ��.�������/�Q^-� -��N�V��h�/3x2[M�T��u�K�$�����Q��/�:h�����O��t��P�qY�Yp����>�/�Έs��ޥ�s<�m����vE>�!�����/b�i��>����ir�A�HUWpҦ�T����g�^�x��q���٬�>8sk*��^YS;����8m:$��_J������卓ɓ�X����8k<LӘ�O�%����"sT������/�;��ͮ�o�(�����H/ex� �.�h�%B��ge�~8XE��y���,��%Ŕ!�<���$���C�?1��o�D����s�)��äb�Ģ��U
�b���T�~�z��Z���!?��cO�q���izC��o�Y�{Ѵ�]+�P�D���3���5��}���pS���M���ǔ,/�Pvymw"N�⥋f��ԅ�q������  "����3�[W�H��W�}�Z��ʉO^�/=�JV�]?�����5�g~�DT��8۲cׯ�w���Ѐ�<�sӺR����>gC�s��6%36VH�Ȳ5���E�.(n!:a��JJ�}�,������0��яC�$����ܿ��f���M�^)�� �9��afa�a@*�Z��Vq��R �׺7��(���Ǘ�j�L .���˰����0�X��40��HE���l���_Q�c/���1�\lPX��C�-m/1foڦfi�=��>�s�գ����R���~������(��[���#k&b>2���:�'���׆g64���(M��A!��Ci+V��p��sK_����);X���ykS3��ˢ��b�J�4��x\�V���WQ��Z�JHs�O���������|���91�u�8�a��U��vYj�c!$����	��g�d7��%��dOJe4RN��e39y��}!�}�v'c�_9m��껎>��g��8��:؊(����C���,xj�?�cJp")�=�i��W; �7DW��I�O*H|KN #��j��0��/�_5U	��EmV�7���ٵ��s	��Ve�a�����̕���b����iI��vT��/e���Qݛ36+�������& �<�|���LFH~|d�eP �<�Kd�0k�mo���}�L���A�v�<yx�yJM�c���MW�uA��x5�r�ñmi����I1B�R:g���݄��I`1zQn�d�K�@)�a�G�ZV�x�(DB�����N#]D�'��v?ʭF�>D�s��g���5����`��<{UsF/��g#�E�m����I:S��� �U��]�![���~�Yv��:$�|�f�>�AT��L�z�,�)v�V�(�%	��[�7d�fNc��ΖP�:`��~Cت^�����gӂc�#���rgL�W�ʭ-[��,}�g:��z,�I��(��@�)Z�}�C���sx�Ɓo'�Z����*lg���Hv��0��r����ä�c�9+$H���z����K�ɥjs<����-0n�A���6�M�/^�<���ٛ�>�i�t̪!�gU����^Z �X0>p���u���<z_ap�!I�=�!؋�̤�pk
�滑�7L0ȩо��Ȇ;��m�j��V#',nm�%٘��UDm�e���C���h�������a�ߴ���	eǸ��,��pc �����R�)�t�~�؋;�W?V��K�hz^{�Z�nP�����Q���m؟M(j]�yg3?�27��&����F���ۈC�b� �-~��	p�7�A,d�����Y�������~c���誰�p�>�0rY6�9���-�vK��S�AZ�\_o� � D@���ex�t5�4��ق�U�Ն��W�"�̇����h{/��8��-C��qh��TN7r�5"�R�W�W��'�K>��"�EV�/�]/��U����^���'�/x�ʓI%�}����s쏾��������jb��`�#�uo�6C�W.����I�����e��qʭd�/ʿZ�ҜB�h	����oL<����Z���� cGc�(�[�Ȟb==�U�$`��1�j�!��d����WX�&�L"2C���9�j��W��~���|��@
7���j�/��'I~c���T�����ZC�M6@�,
)��רE\'}�������j�-�QU���(�F0zpK����tC;;��`$�钊�^����̖.刱�i
�	HwkS�n���9u�/�k���ĝ�~� _Ԁ����(lL�8��LS���~~��
g�����F3�W��BsG ��(S��*�#���a�c@�p�*���� MW���<w���8�*ZaE�oh�<��^(z�",T�Ǔ�G[���0�=	@y�|��q�#�!���Ks���3>cW�k�?��Y��!iď�p�b)�D�c�d��U��ڿ0*B��M�+�U���\ΰ(JVI�,�˸��KD��7;�m��h�y� �XSӟ[\Ou���R�UX[ ;����)��	l�;ڬU�
��ع}�r̵�UU���e�������"sjio[�5���YY�������A��/jP�ٴ�	�+m yV���Q��T�Sqڳ����{/Ia\Έo#M>\�����*�h��Ӷ
!�I	��ь'��S7�&�rQ
?k�g�q;�s}�7�d��\��[�z���ɤ+�u��,�ǻ�6`E��)�8�!�f}M�E��3l�󅂾x�@�,<~GB�+ua��A-��bs�t���s�+JK|��F9�����q.�ٔ����L��r.
� *G�()���-@N�s��iQiiT�u~���+5yǆ@@����5�d���]T��J��ݒ�R�p�¼Kǚ��*�M�]�o�?l�΁��4<�rh���t���궛�2&FZ%S��\��6��R(�Kq=|��@��U`J�/��˲���.�#�d����~:��H�s��}���
\���F�Ǹ�/�n}V��ȣq����鯇R�����q�%�SX�Q��bڋ�R��vEg)<�?��ܐƄ�I��b�@9ك4��n�C�!�([�����`�YϏ�y�_�3��h�`|ť�����ߊ`�V����}2��"ّ��C�Mh�i��Q���}]N�&HVZ{q�|�?QRu-ƨ�vKp��&�߀Y<�!�v�q���ä˶�3��(�Xqew-Z<<>I�{Q��
�
� 3c�v�À� Np--�J�m�Cx	��P��΋��:U����J��HV�Ӻ$o�;��x��k�%���eZ=R��~��'�℁�M <<��Q���\ްa�ʐ��XA��k��k�C.��B~���q�jU�kn�.� ���+w8d�W;���o�����gPPвZ���9�򢸞��ϋ���_��V��^p;i�Q_H{�g�m^�!:�7|��*�հ����"�	}l�PK^�Ǚۄ1���ecY.�b��"}��b}�Gf��M�� 9),�۴4η�g��j*}N"$�Nל}T%W��r[����|&�����a[Δ�	�~�g��p���*������X+�Eq��Ğ���x�8��j��t0#��tl��;��\�&;�-A�3j+�x b(x�۽q+�/�d�f�?��R]e�|'��;m?�J��/�룲l��;Y��~�u���@��}��*�i��G?pr���2���Z���V����v��ZX}�iE��0z_�E~i��>�0̼L�a�����\����f�`�)�Z��F�rr����pʫJ�OsY�U�%� �uX0��}��/���@Ch�+!�H3l��������%|X���+tD�Ƹ4q�Z��OQ�a�>%��E�b�����`*�Zy#ʪ�����~�zD���NdKg�/�4P��;(����d��Ò��	�
\p�����H���i�t�z3��Y�6j�:�ɨf�����vF4�>goDPG����.`�aB�U��Hu8��&���uo�����;qq9y����� Z b�:�6�a�F�*G^���H����,�ͬ?�h*�[�v�˛[ٷ�3�{9�C&8�=�'��L����FXeb�U�p8�!\�Ԍ�� :q��R`�s�A�;�����A!A#�U
�DI�s XA�0�2����ͱ��zj	k�n��1�x0{3.l�(�z�ګ��@X�҅.o�p�V]%�.{��~�j�S�|PO��B�+ێ���A �:�F��Ķ�Me���6�n�D84�ݭ4ctv=踸:R��F�����a��F	������Ky�(�^Ɯx���i�_��!���������V?@��Dٛ����.���0ֿ��?��4T7�8�Wd�D|u�]C����[��^O��<K,��>�¼�� H�����@���rAi�-��Rgj��~���[QU�V/��Ɇ��h�nt�YO6?x�@5Z �h�������hc&�r7#Ġ� �2j �M<*׈���Y����J<����f���;d� ��˞b���w����R*m+�o;E)�{���Ax%�W&DQ@�h�zQ
ƨ�߂�ȴ_x��Dk���Z�rc։����������
��q�!%�Jr�:W?�����d6
��������)<0X�_%3�1V:N�D�A&L[4�̰��v�@̈́/�(�����)A-�� Z�@��7'}AknR�3D�؁V�Q�3B��
k]3f�	��",���P.0JL\'Z:Z��?���Bu���)���K�,܅I6l����En<M����/\ DH&�a-���w  �����o�côce���R�F0--�Aje���v{n&%�i�3�/�aU�I���9���v�3���Dmx�6�3۲3������1����|���]v���@�g�ɡ��I��x�C4@�Zyߧ*���`����\��;�i�}����JxjVG��w'�U{ ɦ�/|U���-V������&��Ȋ��Db�W�''d��$(�] S�P�󵜿���T���%!)O��w���x%)��ca�35Iy���3U�/��U�M%o��S& &���Ճ2 ߧ�e�ϱ3���ʖ���N�L���XY�%W�[r@If�3�XI����}1z9Ck���J�DN=�nŮ�����G�r� "��D5#t�r�pW�mׇ��esj櫆-l��O�$5A)�D�ϓ�d`5v�o�h�B:�����w]0P���nݦ���K@_b���/�.��C�h�Tކ���"��?v����k+��BR��@�$��g�1�`�I�W�X�)������T�Z
Ч|*��b2ki�v� H��(���|�Dy92�l;�b-�j8�M+$��	�p����0|���|~�Y��4fR;	�Ϲ#��b)iJj�7�``���E�-Ʊ��o�u�T���cnU4/�۩̀T_�Jsbr��.����H��R�
�%=R�����{�TM���Ã����⏖`wHC��d�TjV�c�.#��.ˌ-��V�P}�v8�٩�OR#�py@�/T���E�6-���Pq��G7^�����u�Bt�<T��$Ap��ԖG,�V��Յ�ǟ�5���:�;>%\D#�/�c{hB@�wu|�������ڛ"�]�K�p�pǘj�#��0CHZ.왻F��2�,5Qb:�.B�fQ�@���PJ��h�(Sxƹ����K49���4�'��� �Jd���mhF�u5�9Wќ�F?��	1Ϝ�nF$���n+6��]3=K����ި]����ci�������!}Ղ�fe�${;�{".I��#�.HV���8A'?	��6_��t��w2���Q=t��*�@��	�X���I�Ǯ�	-�Y��Q\s;�Z�C|��1��?�`�5M��S�#BǶ��U׽�7oh������h+0#H?�.+N���h@��n5�q�����s���5]s��4OW5�Ѐ�r�u =!9pi6����5����Ú��~Q1���X�s�I ��H,� 	O�C���3��b��<鄢�A#]fr9����S/�i�:0�{?�wD:���m�`7�R�jP��iXE���cҶVԃα\�y�'����7䰎� �ƬO���,����?����K�KG�)��
���^�&f�L8=5��b�K�����xb�M�ߌa6(��ՙͬ������L4&r�n�<S�*��)4�
�Z4J����}���z���d��n���XY[A|}�D)XO�.�^����z[�,���px"t�R��ݫ���2e�$���e���Y��)<r��c3�]I�z�S�������M|<�m98�r甋�`�V/<� _���X�+�{E��e�\��Hj�Y^���/�	�dT�>�ϷrHSshJZ=��n�?S��Ŗ�x��y�۝���r�Ԁ� 
Qy��+�|�ys�ˇpX����+o��\G�O���`�7�[�F�2��m��f��"O3`L��=<Br�z���ڦn�ǽ-��r�=��[�r�1�lw��uDe�|2���u��P3�v���t�7�2�Z^�|�a�-��W�-��/e����"d�l+���`(�4��!�BR����7{f2���<S���Z1��JD]�.���8����e���C�L����0<��v%1��x����8я���W%x��?�#K.�n�!,y;���čU�8*^��)���������^�i�V�HY� I�L��!a�/r5'n%Ȉ�KK����^ ����^����h���^P~�"`��!(�qN8��c�LZ�w'�om,�-�j�m1���/�����KY{�'���_h�������Z=��
�Z������m~�ml!��l��梻�QA]͘���%m���4��u��)k����T��L�u{Y�6}~�7��0W	j��>�_�v5�����rh��w��k�cq�f)���fԗ�C�!�����0�g	V��s5<���9���P�!��9���>���0�Ux8Xϵ�I�Ū���P{».�F Df�5�2���T��\���^�"$�؈ ����` ̃�rE�R�(S ҳv���b�`2>�Ƥ渥�p�>�.&�2P�@u'r��/��y����
�ԟ/6����Z��c��8V�n_� �ͧ"�ܐ�T5�VV���mX0R�3=ј�Gm�Ь *�We�`�k��`���s�ƫ�_7r�D#_㫨QzR���#Z�ă�Q��`�orc?W�wRUZ�iLJdؔ�3{x.�~r�u��n�Q�P9��<h#���X��G�.��Dl\�����P��w��������qY��#ƞ�R3����B�mbk|�y���D`�K��ǚ1�TM���>;1�}Nq��B�1�m�.��i�P%ZB-����'Le�X��E�$���3�L� ̙�`e���x�I�`�����P��6�B~B�-_ʥ�ؙp��׷��Ǳ��d.��H^�XS��|5�-:�1�)�@�X����x�8��]�ܪkB�c-�-���Gw�̚"f����n	4t�z���?�2��`�����M��Zwח	�[�\E$'��p����Zc��u��
����a��-k���Ԁ�p����E�v�QLD6��<pW���<ԀA,����	�0���s�Z�3�O�����j�Bh�9M��0��,ƐM-�fC�q���5��(�z�o��s��,��VP�k�9	\������.uO�����8o��z�����$4�B�b)�H��^�>or/����l�O��/��L؈�u���YAn�"�ر7����htu�m-4T��/��K�yu�n6�M�F��a=�S�����>�$� [@D�ϫۦ
I���f���ڝD��;�Z):A��̾wѝlԽ��0}"�^V�G��Z���:�P�|YF�@ s�ͳ:����+�_<:�ݯ�6 n �> 8j�Ŭ�96��a��|�*��ԃ��e<�~4wo�jƳ�l�	�
{�H��ڭ�gjlX˕�(�nT��6�y�CL).�u��ԃ{�Dw#v&��͋�@��7:-��Rn����35?U�j�/�
S|i�i8S�E��m����CL.�h�u�v�Y�/��$��#d���Bc2Am�2o3��`��	��#FrV7G��9LC�z�R~����<'��冃�D �|�'`.Šl��8�(���t��um�f��0���b��S�oC�5����$#��9����So�� �`���s��:�����0W߱��
/(���9?Jث8�c֤��T���p|9=wc�s�2���A,��5��L��;� N��Q`�U�2e�yW35:ϢT}�z-�O%=N�<p�ܩv���5��]b�Hc-�ƳS��Ȱ>�?+ɍQ4�.�i� 7�o_��V-1Y����M���"����\d	 ���gm�Y�yt�~7��x����'ō���!������*�e���{|9��㾗ő'���0�2x��������"E�KF4�Sۧ})૒:|�WmJ�����7�3�79f8�v�낔]�<Hb�{���ِf㥤�25�����^���$�^��q���{	v��_5�������q�`��)15�r�0_�WE)�k��*��a�F�wr���$����g���T��6�#1�!��ܡ�2u4r���'w񐣄�oE{8SB��7oѓE�@��.N���ӃqT=�g����u��{��QA�4<�k�⒛ƿL$�B�.��5hfGs4�R�f�x 
��&DF�5ඏ�"ʠ��DG�W�L\am��kK�]����t^�DF�FS��+4���	|s/���K90�^�^S}�{d��qatN���A\h>��f	m�t5�ýhu�|~4�"����1S̾�;�1�4�6sf?:�("v��x.]�#����\�3��v�]$͘$��W9�pڳnB�@���ۙ�Xo��a���=�q�wzd�X���f�_�*�aI����O�1S�m�W�'����	EPIK�;�,+^�����F}���%K5!�fH!�5����H A�j�6і(s9��
�v� %v1i�8�Y��5��8z�1(��-�M�〬,tk�p�ȝ��8UrK����O�|��ݦ-�n�5+�Q;��k�:�Ix<h�bV�2��:�c����Og�Q�`�ơC+njo!B����������q�2Քu�;CB?��,~8!�H�ƿ�q���L��	4�'M���i�%p�Gƅ��h��Fd�K K�=�3� �w.�΅�I��@���w[�,��-m:p&@�c[��q�+�ٶ�`9����7��(v7hz���J�����M�6�`g+|��7W7��Z�=/��l��9�`�eJX]��Y="^o�r?{x<�K�!y/>�5��u����-�do�$/g�&�ѠGK�$����a�}����_D��C_���l�7
�`��T̘b�j��'�31�F�����rM�;-��{qƸi�ӳ��J`�:��A��8��"GA�?$�;D�R\e���TY�_��ҍ�Ux�4�X
Z�m��"�T��љ�Ӥ�M��Y�9�~�do������m
�dG��dH��*C�!"�tn��yj�þ�/�TlkM�#���D�����e�]Q1P�h����hQ,Q��#p�;�& �O�@g�ЄH�D;0��Q���V���$t(v�'�	e���n�OG�<��7^�ne�-��Q�l�!�T�	p���Qs�.��y�w�2�֘�.���Oz{]��ی�ݹa(c)���?�.x!-(�2�͋ѩ�Do=B�9�ԃ�kX�v���X��CG@t�j��N��%� �����6\}Ԥ���^�����니�v���D#���x�uc{���� ��G(%��&�G��
��42=��.byN����J��t����
'�3���W����l}���!��Zܥw+X
]�b��@�ao?��2ON+�j�H�>��]�I�����������m�_L� ��/"zcB�s��Ov��oU%�a�D�6��_��Co���VC��v�������8�E��[����4���*i�v����:�貑��#�(�������rWM(`Y�K
+�Ȃ�}S����SШ>��8���h�p_����,� � ��ʪ��P<l�����p�
xv+���+٪��r�Vl�>w��b�f����i-�T��~�/�?�漙l�s	=9q��@OU��}�d���za8�!>��}e�����T� �=��̎�C�HI�����}Pn�<�_xN�2o�mi\Um�B^�t����40�<gq,u�N{��C�D������X�Em����u�!��4���zZ���i�Xe�����ޟb@!�J�[JI
8
1�iƠ44^�/�0:p��{ؽ\��~c��<T*�U{�W������n5��ٌx��F�T�x9"s� rIu�=�\V��&�)%LK�f����gz8����WQ��	�^^	w!����D(F���� Y1TgaL��Aܪ:_���~��HPg2��O��e-�f�Y�������Tl�kR�"��cH�C�CKjG.���o�?aa��ř2t�P\�{wUV�%���^>Q��������Br���
-{���q��@ɣ�+1V��1<[��!����%�,�L7I��!����k��`��7?Ӄ؏�
1�����u��eȋ�}�rƑ��E�HL��T���n.������4J� ����qC��$�iCf�f'�6xm[oM/��� �����`��ŏS5<�7NZ�:k��L�I�Ь,\�o<���6�p?땢�l�*yU���
�T�K5��^���~K���f�v%A7l���̉4�G� �ph�XB����1��]�Ed[�0���W���^� ��g�3�у�=Q�����#���xeF�Q��Y>��e��{"��0��#�oJ�}0l�Cq�.&~ξGeA�ø����T�X���Y��0�d���형W��i9�%�.V}t=���3)�L+^a^"�|��!�������x�+���Dn[s�Ș �
���XnSs���@�{�/'���c��\�qn1���Y�{�x(�]�k�y@�2��w��v`N���vD�e�� A7�&a6��G�����v���n�w��"	��n�L�ӭ�q���r,VT����1/�l��;�j�O2�#�ܸx�
��#ϋXtF�����P��wղ:�q���1d�M/��
��V��^�OD����j?�e���ւC���p��K�+��Y G�g��	�/;Bn��UZ��^ۯ��lP�5Jt��y_j�"~�Ow�R�F���݁��ߦ^l�Jac����ᠢ ���JA��߇)f_5�߱���)�$O�Ƽ�ɓd���j�2��Ȧ!|���A������ͺʢ�Z�3V	{���k�NJ*�m��}��쾓�`�VV1�j���s���5пR~�%"��ِ�G�o?0~�q�rsi;��L��?C�ҲR*�o�X�
5%bv��7O�ڊIP��J�{Y*B�"��^3�hGx��,�4�1^H����{F�oJ=P(�HE����W�v�>��Q@hi�ލM^Шl�t�7ڽ�r~4�΃�����g�cĞ�B?��ɽ}Ӟ 2MVO���\���7u���>��d'�?/\_']
�9�s>;sL_�AF����j2.��(f���n�}=�ڐ�,@�I�X��^�6��^f�e:Y���
�T��יڛp�ا�V77K>����:�R���b�zϽ��V�hg��,@v�<e���" ����<
�s��0���j�BS9Ӓ�uɧ�I��7,�!���c�O ��F��$���"��(5�h���)Rg��+ ���-��ψ���[�T�$��i�7FJ��LJC<�!�����YLs8�]�:���)n㼳Q��N� 1on�GLbu����],�2nƚ��u�w��jKB�f|w�X����VΈ����kE�<V�>�a8�u�.>5�mMf�U��3�`�:xZ�z�w����4Y�?����"�f�J���E�x�9NM1
Z��JA�~�<�h��}#ь����}����p�/A^����>��-��X7�L|�_��ЬZ~��9����"���$��3�YU���͉^�/|�@sau���8?
�q���߫x�N|��7�����5��~��5�IR�+����_!�n��!��4��b�}(�TY�H�4� �
-��	�M��ſ���ܓ-�H�X>�!�Z�p*�S�*ש0|]�TPsD۪O�iރ�9�%	lA[\��)K}��nx��,�޼��\�$
�׬8�a"�^�uB���D��Ȭ·ZiBd����háȩ&p8ݣ[�@`;P��)���L^@��mE��Ϙڴ-�-��$�=���3D�����*���9h��Cr�i��5�������a�Ț�r�S��9�F�¹���bd�.����I�7���S1b���K��@m��*�]�7L�N6 9GG/+�2 ?u��K��C_M hG�9�H#̮�I��� �
����2ۯ�8i6�[��rLɥ��@�{Pز��B��{�@ΨT7�9*(��ٙo곒��T�IԚ4��w�[�:�ک�D�nؙjm�wU�e�;)��� �=M��ʱ3)���!���X���=<�n�,ES�[��	
�rTY4D�d�9���L8g)�I�C�c���� �󿊫�O?�G�gL�$�U���qy^�� kx�#1�G�">c����YH/W�������������J��ҷ���2�{��^���ԅ�^7&�4�G��yxZL-�2�m�sޠ{��5���rOn�`x	�rE`K�iv�h���@��j���s�wE�d�]`�4��Z��3Բ{w�|�f-���]�&�n�ne0� ���Pfq�7��4k� �ށ��
�@.��S�3�,�o~c�Ap1H*��%�qB���HJ���Ї$36�55��O��&�;�/�����G'f)����룯Q�~��QFE�?\y1�����B=�+TC��4$H}����f�j��?�\t�������t��(�Q�|� v�S�.�x�����,�ҕ�cf��7֞��`6���n.�������]sF,�㈹ ż|ƈ� �>O�	�u�]��/���� �vF���0�wtG;)uB����P�Zy��;��(a���/����W��k�D���Ŋ��S�Qԥ?�a쐝|2	bz��^�����ݠb��t
��� �K�]�!۬%��"�Źf�����η�UG�U��b8��x_��ߐ��Wb���3^�S#�,g���L&|��mf���l�6m��[J���	\�&Ò���$Q�R�LNY�?�f�'��d�����1���<b��A;i�"�=�ڂ�ϳrK�{�~l����tH���͏Ja���r���)����xn�[���vL�3�99v#� :{����J��&�݁�E�=�n�'S��*�<���r0n����K����{��ʍd���&��&"�R��C
�>ך��a���<\j�t?�i^^#Gz8��#�+-΃�C&���������\�a��f��Z���!�߲��e(>$�"����.�JG�b��^@�Jc3�h�۽��ŵ�r=G��ڱ�S�=��:�}WH���)�)<����s�:Y;��H6A���s壗 z�
�XiXk)�&���p��������6>j�G�V��v�+�U�������O'�Q���z,1�W1�9Q�q���0�I%�*�
('9o��,P;��
`Ó��)�EaK���k8<#�S�RV�� ��*-��ېi���u�/������lP!��)�_����Mo���x�*�?Q�*�u{!�f������Ā��T)���R�7YV��9���H�Y b_�s����yR�"L�є�̗�V���P8R�|!ר��{<Ȥ��(gz�sHQ9F`���>?9�н{��tv8�p_pK�X�U�{j2���A��-��c��so.]D�ٱM?�ɳ-�wn`gßoՅ,�O�L�m}�D�H]��LXK&����qԜض�|O�ur�'v�P䐑o5[�5AҝvKh�D��`�9d����@a_�&��s�f)�T�b-f6���1U��'k9�����M,��v� >��7��h���k<P����+��VȌp	�ݞ6��*�ֶ���{o��
����8Ͽ�s��MV0��s�-�)�P�^;����)���%zE��k�U�vF{-��c�_��*�.�xҕ�	i�)"� ��B�G�/dR�v2��;DN�(:;���~\��Ю�zu�;j�Ɖ� !w��˺啹%���h�� X�ѿ�+�����ǁ�:��b�nt��
@B���
20S���R�!R6�'m��g�I����4ϐt��L�'�nsع�9+��Ѭ�@���U��Zb��a�"�Z�PAk�g��c�?��=��{��hD��dL �5*����"�����R^����7=j��X�Ƣe��4����5
4�e�?z�qM�Ng|h��z��_7�ؖ]���P��5p��8��Ӿ�� +��n�R�I�-/���gVD����I���k��s�e�de׾/��ke8̯�8��ڻoFY3�mK ��� �39�B0J2�ǈʛ9���>�Je� >��ѕN�2����G�밽�Ҫ����V&�a;�y�u:x�x�4m����}-�s�.Cy��20-����/�8�qZ6�#_Js)�/�R��q��P_��1��+L?����}[����h�S��o����ho�������J KI~��h�#}��Sǖ#ȸ�W_6�K��Y�P/
�h�OY����?z�Q�/kSǧ b눱��j���A�S~�R�@�a�PO|�עG$Y����Q܅��Afd�j����?R�Nc�����S��mX2�r�B�����*<����]�uPK��X�<ў�r�	t8��=r�g�Gғ�y1��f�5���Ǣ�,G92�7�o�&�w%�Ւ='��8'�+�Y�����\CGZ�\|k�L�d�+��Ѿ�R"ھ��a52�Kr�ɴP�x���P�]�!�В3����r�u��w��j�R���4h�2R�Z���E����w��Я��&��l��D�½:A]�T(®R��׵p3RI%�$��|d�����qd���\D̒�����%�I�x
�ea�XV8�`��C��Y2�	|}Y�c�NF��I
��a/49�1��D5�	oXp;&��e�����2���3��:3��W�tt.����|[a�<��Q���n�f9�D��w�5��8
Q#PcN̵�1�[E��ߒ�lR����Vs��8�ع�?@�lt.��x��pJ�o"#g�8@��>��-|@�OX6hы�L���q��z��*�:�Gu#ɖH�	&��R�'��ʪ4k�,'��-,���ʵ~G�xߟ�Pb8�����LT8	��7����f6��d��_��,��H�^�Gi߇���>|�!	K�x$\����vaU�[;	Z�ݺ$ ���X�[Z���l��!C��>�<	#dX��ĝ�A���Wn�ށ�t�\����9;1���E&����
Yd�!~�|�9���(&j
�kJ]�:�V8_aLw/S����Ϡ)��Q�PgM�(3�(����B���G��q�z�Dp��OJ�{���'����-
�89��X�-9tH�'�9�1��R>�6A��Q)�a�߮w�����*(4 ����/�[�"�Y���f�o++�~j���������i�0�i�h�"z���K�a�6��{��i$��։ҳf);%ѭ��r�YNU]�w��Kz�K}Y�Pn���<�dӭ&,wE�*��n"�B��4�{�C�}��p&ٳN��@b)�k�E+!��?l b����Z-�a����\��6��4{Q��2���'�DE{�^�&�}K}1���G�6��ѻ�w!l��&qsv7�)������`c/~���WH�krfˌ6�&�!�ĳ�r��8�=��Ψc�rg*�u�N�dy�&�H�u��oS�9<� {x8��1��WH8���3�H%��fH�����T����ך��P�wJ�c��l���uyhqvAm�yؕP��S��v5%��j������oҠ�+����f�Kh���	���L�ﱪ����ڗ���i:u:��%9xY� ��q��!1�G�'7hpR�^���6��S�,��^���1�-�`��>��jE���h�JR�t�+dq��(��u�y��(i��M��ט��m��~ �N"�k�eDD�&(e}w��ީ��o?>m=&���"�"��?�����-P���YT0���Mq	��5@Qփ����
�ۼ�`���`g+r�0�)�m���1�Uь�[�(�bY0���0�8�������5�	77�w�)��X��C�g���W_c�X(o�E��ͭo�;�$4B0����٩$���/��J<F#z��03�U�7*����
�֝?}>��C�;-2	d�����<0SD?}8do��\�N�R�9K�'��`����0�@�&����g���
�-,�m�ϙ	��ޚ=�ָy�lFE^��7��`�JX=P�.���3�jh�u5:;﫨�y����2�<�aG[W(n�bP4��aB^�젇ϡkI.swۦd&��Q�נa�����8A�l�/w�����?����r@!�;��F�m5�9�}���a�A���#cQ�9�Ǩ(C����"{����<)������sxl�b]��x��x����׆Yzp�&+G�.^xQ��֟�~�� 7���wsi��U_���B[��d�}-�ւ:���\�}���V�i8t����M�s�qS9]\����N�\�u��Xr����=rp�0�Y��r�x���h!�Xií��n�PW�6�)ɦ��% N�O���G}x�W��M��~�".����,%�>'�Y��Ӿ��G^2	`�yKk�`&$�2dntf��﬜<n^�������>""�9w"���t^�i ��CYT*�P�l�^�MD�����4����(�{�X��5D���|(�"����ɝ`����K���9�Xs�t�	ΔC�27�SY�a]M���Z�q���v�9
�=z!a�1�3ݞ|��\�g� >p ��.@���¦�\�JB�c��E:Չ��=�%I��ud�o���AX����EtSB'�xqT$�� �+�>�ϳ.�0���$U�^�-vҵ�o:��-�D����R<@c���~�(��vhAm�G����_�A�E�.r��� ��3�= 	��r�r�v{�S��zR�_�SG����
�U}��y��N��?��ՙ��R�!pƺ`׃/�ι�����z�0iH�UA93���U�]�{Ϫ'(����h��޸�u����^�1:�@�+'-���	S{ӑ��X�|ƶ[������\,`���(���>�����hNG�x�|�GT��n�3�$K@��j[
@J�E�_N�_����3z^��B��4��2e��rܥ���(�ƬJ�0ŧ	= ��b��pJKZ�]L�<����|Ȯr`*jg���R�N'�[cMm�M�,͉b�?�����ϋ�#��F(90��Ml�.��"\K�wD��Α��#6�?a	��$�^�oU>V��h�� 2�!�و��J
$8��1֬f�6�p����S*w�w
(��>��+�+V�2�.I#h|�'e�]�YywۋzTO��3�"��:z�[ٲ��<Śh	��&���0D&������x?0�}2�]����웅bE�F]>R�2n8��{eZ0�G(��3���)XW�2��OC[��㏑���(�u��.ܥ	[��U��'���X̐s%k��N�,��[w�;���|"��R�	)6d�m��i*z�2w-}7�/�\p����P�rRD������e������	��7�gW�.�I7z(�֗��!�����]]xs�;��f��'�s�]X҉�~#����3��o@�(uo�-`�"�4�����}���&zB��z>+^�;��9K�v�F?�3� �s��w��+��L|��	����`�m��ғ���Y��n1�S2�N���(�=��y~! k={�ph�)�}[�5�YR���Z���e@kv���郘����*�cT@��K��f�;�5��J� ���3Z:L�oG��Q�s,㦛�KVp����}B9H�D+y�$�e!�P���SZ��������Z����(����\�f�0Q&\�i�%��Ojo�����N!�qn��X �9��`���t��#l���̇�]Ru��ݞ��FP��-�I�I|ս@mz</��F�����7��5ֺa/,Y�d������;Ѝ�±��ാ�q��Љ��r�&ʑ!v^�}Qf�T@Yu�{|Sޟ��XJh���>��]Mc�����X7��Y�5�Z�1����j�ؼ��^L�n O�Rk�̻5��=��_�uב�,)}]%ay�w��(M[��I�{׼U�juE�]V
p�d�HI���1`��^�Ô��~uX��E��2b�W��	���Z1u�)�%H�p��͖�]ꎛ�F�AC])���u�u���}o� 0���Ԅ)
>�M� u� �=*ɿ�^G}`b����K��%/��, ؏���4h�~���N>��ì ���f(~R�c9=MbK��N���+�緤[Sc�&��T�@!��RUv��9�,���?A�x�|:Z{�L�Q�����h��2�����=�f֭���w����S!GhHʟ������[s��3��}+����Qq�nL(_�Έ4dSI���9C�ܾح�k��+)[%_X�J�k�jȈEl��aBm �����Pǂ��Y��4�[QS��$�"~fJW��P�+1�݉�J��\3z%t�
�]�;���9��p�ߋ�ޓ�
4�!4�xl���G;�T��E�ra�
��D���[��\(��������\@�v��
p�L�w 	7Հ�6h{)^s��:� ��Ie� g�f�Fe����-�a��m
���Rw	�zm�8P���e���2L���l:���ߊ1JH�(@k9L�^�����O�K@��9$.�o�{��n�s��{�!k���¿�mx�:hgK�tĴ~�e�6_����
n���Z��d�ڕ����jƊ˖�t��p��ٹg�9 �EdbPl+�e�Z�g|.���x�F@}�V���ѐ����(q��w��F�?��& :�Q_o��{�X`��GJ��[��VM�-q�}H�ϝ���.��L�G��%5ń��_U���GΖ���0��IF���crp~d�D_0�G���z���>Y>B�CZ�@�:`��� e�k{�k��g�]岭d�y��.�����wA��y.�jg��g[���=�R��`��^�'�8�:��5Ԑf�v3�f�Bz���DP��qz��:�P�|����ʓ�Z-Won��7��wC5���%�N���,������]�We�`��6~�5c05�c+�F�'��Z9�c8-���⏵}WF��C��B&���Xڸ}pk�GZ}9�wa�YF�hyx�$�>��j)y,,�Ɗ4�o���Z������<�T��4y���jLS.��8�fMւ���� �ix�6�O���k����%�!�t�r2��m*�誅��xEVyl�생ƻ.�	��M�i��#藡���%�߅DUx �h�/��ބ�S��=�,!/�)�i ?�%��c�i�U�,ɼ?��4�J��G[��/5$���|�W��� �S��"|8坆C-j�f!��|�m�h!��m\c�[�B�;O�#[�k!�9��ߐ�<��\01m$���^}BH�4!�����]��+j��=X�Yҁ�f��n����hb���c���CN����{Ɣ 2�!��`&#�,L�DgЖC�w!�i�j�N�m����O�<�����j�FX�]3��a�(����Ա���jI�?ϻ�. Oq:fG�P������u]�YZ��QW�Ⱦ:��t-�T
+�W49�,P���p�F�N$ybu;�"ʸv8��ԮG��z$LK!��S9o�V/�L�f��Ա��r#a��q86���>);�B`G=N	I��1���_Q��Y%�U�_����ꞩVܶV(��/>��9�����
EYS�ë6V�,73���k+�Kf$��m���S��g�%.�+7���9�/ڳ�ls�H@���f��u�΄~F�'���1j?s�m��C\���?�����h{�
)���dJ%@�,j�6�@��x[XCVh�q��EÔ#��+�9�)�X��#�0(�T�C����=�߷���F��!�
��$r�t�,r���x!�K���[|@Myj����%�V�%ZJ(3h���3�?C�q�Hk��y:dq�ك�>{ {1��2��%Xl���,���΀U�� ~�f��~z༹�5�S�Ig�H*�I@����#F�l�w�M_JVB�w��Ұ!�����`|?�N����M�����>v9Ñt:f��N�v�T�ғ[�Ŀ/$,��B�~#�~���M]�X��u�{{�����r��#U���7�8T��s�V�@Js���I��oQ�lf�?��}GS�3�����쟞���Ck��s� ��ƞ��^O$/�M�\̙9P��s�b��>__G���X��\�W��P�C���+��ü `��^S���Q�>�6��%=�E0�h��P0|4b��d�lC��)��+ö����V�/��tTt�v+�?>��d��[���;�è_�MI��T�ﹻ1��n�YH�^��P���kV��Z��.TÎ�&��xOo�Ve�v�?�*n��`Ou<�0��.j`/
 �`����(�%��������=φ�x^#�8��9k��,�B��F������Ug�:�i����z�g'$D3��9�mpS�pl��Z��b�M���\��Ϩm��������V���p�����-�Z�I���xM��V�-{޽?<�(�����θ����p7����k��TH�ˠ���;��4D�mۙuɱ��O�2���U��{6��&�V�9~9���Y��zy��t|�s��|Z�Z��Mz�7���7�J����1�v��f���	���~�g��*��Q�A&7���z�k��+[�����]��Py��Ds@�>�U���2l�Af�
�a�5v8�
zx�Á������]�Y�v��~�0���Zn�a�`=R��%�|��A	)�H�R��<H�W�Գ�@���a��)?��;�M����/��{O�A��{�B2t56�b�%EJ�:��R�ҏzi�_s�˓�����Fǔ:�6�ٛdSDx�]x�u%��):4,T��8P 8�j"S���W�(|	C��4n�:�-�!N+�^��}(�ڡ!�+��7X�Y��`΀|���T��==-S=�V/���?�$P���ŀ�_LrY�}.ĉז�6d�<��^�ϫȥE	u�2�n��DA������-J̕��x��?XrA<).��Q���q��E�ٮ=�v���hE�汘�!�%~��b�4�Z�~�T�cX13
(��R�K&�5��8'���1���a�=�#�y�7X_e5��@?�$��П�2�&���;�X�Î�u���b�-V�,���GyQ�4b �";���d���6�`b���~�`;J���#q2D�al5�h���9z���%�>�J��)��X�L��ɖ5��k��Sbv�K΅��SVah�$-|��k���D��7�ge3:�M'�틚���E�gG&�;�<ƞ��(W��	���(t�/v��;eW{AG&~��W�4����3����}f�5��+*;�x���������t(%�����.������0�cJ���G{�h�㝝��m
,���2s2KI\T�4g����&;f+<6D��q� ���H�dw�[��3�ʝ���c����y���Tp��3~�.��{��=!h��k�M�on�j�]��G<c1���cV���ӡ�Z��nf!#��s[��h���N�bV�U�<��}`���ʻ2f��Ёd x�Lߘy��u��X����.zu���Ձ�!}�B�RW���t��Q�#lƴ��M�[�K�r'x-Ξ�w�2!B>%��C����d�l��F��jߦ�շ�u)V���˵&�$�~�m���;2(&*@���̤�����[4���]٤������嚝�}m���vqq�L5v��0�.�*^�D;m���]��Iq�y�J�4ٷ0�h6��G`,���z)��>��	p�C�q�TO��b��,`QE�xTua��S�C�)���`�͜oC�Yy��z�Jӣ��8[���������RSK�Ab��/���!����L����ݺ>Tz�)vWUs�t�5 i�;A���?��T:���qPu��X}xj��h�@��(D����}���|���T�1b�i��'�D�������4I����%���|%� �7c��i�O%"*+�[��Lh�����+�H6�D�7�Yo��"���LT��ˊ!_H�G���a��Mc�'�����˦���S�����լ~�1��������X�u��z��:�����C�(�\����}�TO��r�_r���V��p�p߹�r�=�_��?_)��7j�'.�R:����ā�&���,"�m�7�I����M����K��S4_༶)�̶M���K���+/�5��-h��DP�j �v��y�"����+<e�s����v����	���e�p��د\w���"k��p���"��M?���n-m�W���I��}uwY�����ab52�]R�8�d[�~�������mn���4Ѹ�\���.�c���h��_�9���Z14&�G�:��>O�d?h�r�jV���V@�\�%mLR�>w�h���EI��>Ǝ=��y�
��c��d)=��q J���Ğy�N�1Sjm�{c�I�Ȇ&mxR����0�6|m������-��Q }����F/�򐎿�!(/Xc�q�5R	� 4��26�c��ݴ7#Wx�i�M����Y�)N1��6�����I�C�*�	u@h2@y�w0����{���n�Ţ9Խ& ������P
�����B^��L	 ���'�¡f�#ŕ ��S�q2R�,�1Ԍ�O'���ə�����]�4W��x��S���Q�z��A롹x���(z%y�q���Q� _ڒ���^8>_w��*��5��#�����&�Pa��2 �mT�UG�B}�Q�4��H����5�������لm���卡I	`;UR�hڵ+F|r�{v> ��5��h`�ĢP �X��\�ԮeD�GJĪ>�J+�)�`��͇�wbEJ�a��3Il8E?��������Tz$�`�OD0JC�f+8��:���P�P<�,����5�%��ډ�7/��:�qIjb�A)���6d�z*K��*�D_��sdO�cq��*�d�%��G�3�\����/��H����f���
���R�x�j$�J
�eNO���( �`[��������̰��ŷ&��K�$_�~d�d��÷R���ޟ�co+�������J���[0�"~-(��v1�VI@�]���4�f���m_�b�tN���s�G�Z����Ul4�Q��p#�DZj�ڞ���[���0@{�h7v(�)�P+���Å�����A�J���m;��Vj7<�1�J}E�@&NfC?i5��7D�Ҷ?-7Y�:M4p�T��S�`�
�㎋���F�ӑdj� �9C(�m�ي�����}�5F,�cB�1>KDr��/]es?��.?Ǐ�3ϖ'�R�G~�+ �$��R�aF�aU{��H�ʗ�>�����߱��P�re��"��d�?7E�5�0|:�֐�������Ai�:�����i�Ak�]��4$�]���oT��¿Y��w��e�a��I�I�CJ��u�r	
!cqr�KsZ&���:2�r������(���͖@j��rLqYdwn�Y�p��<\��,�-"Y�l=v�󛛁c�/�Uw��u�烉�(۾U�������ď|��_�l����gK�%e��o�:����5q�
Ђ�G��㶭SA�B�._���--����mJ�p5��eWէzzn��p��(��h01��h��զ�O.�Q,���y���Mct6�Y�W�)KO�����v���h�A�s��:t�M�)<om�{SQSig�y�/ƒ�!W�d���6T������b���O-TK�[�c�v��K�!��6�q�tt|��/�_1��5�C�!?�$+���B����8��{��-�����PȾr.�-�$<��dH�u��g@aWXm׈w��vb2��y7��}&��A���+WӤ�k'�u�u�mi�`ŉ+�m*�L2�o4���x���yƲ�a )}�~ː��jSaA_��Ji����;��>%<�Ȧ_�V��� رhy)�������Ŭ�b���[�n�)pl�� W�ۼl*���)�(�)pr��ɐB}�\hX�$L� ��]�b��I�V _D��.�4�e��Q���`�Ո��
Ŋ΄1%Lb������h��6ƠW%�й�YW��E��f#�-�;u��O�{���S]o7��`KB��<U��`��/���͚��KT�ޤ7�-�~�*�#
 �I7{(Q�_jh�zM"��ӧ〝�^dvJI  �'៵yXJ��y�T�\ׇPX��!_���'"b�wu�x�W�$_ �T!��t�p ��g�;�����C3��5EwX"�ѓ����wnU/ ��ëۧ.F�H|�D�=��#I\Q�q�NNK���빑x�8��V�8�?�OVݢt-�� S��$.Dץ;��9�ZߨTTD$�wjf��Z����Y[��3洶����͔�����Js����ʽS���l1���mE��K� ���ؓ�·�j��v��
���F�_N�ؔ�%��+!)�H��2>����`�(j���������V�H���k�5W�w�������c:/�"����=��R�k��Ln~�4#��-E�X���XB_���h��[�������U�h�eanZQ��\9"d/����S�
{x4V�ֿ)k��&hy�tl}���_�*9�d�t��ꫵ�;li�b��!iT��;��t��B%f�*���S��i����Fj�6G� ��$D�|�d5V)�@��g��ዑ�4!��v,�"�X�g|w�qM�ax�=o�殯]�5���@��\���9��A��$	S�}��+#�i-!u|�>�� t�I�o^�Q���y'S�(�0�U���p��`Ӻ�Fq}�ʔK��(IHGV���]�D��II1���-�1��x�f��%������$I����� w�(��l�|� ����P�li�)����C�M��K�*1��l��A�utƋT9+˔m�Yw�(w)tWT��#�$S��F�l��Y���kh�����3�}�XB�eq���*tT��#~P�枌6ja�nA�������X��Ws.��(H�,�ff��3m rqA�=U���9/�.3`��54��`��E���X�5YN��8�z#Go��7��/�Uo�+AmܣZb:a�fA�\�`��t��U�ir�OX��t�n��,�˓(Cj�T>�!�+��pӎy��o�,�lg&�\�ߗ�a�႖�lM\*Qqܲ�u��cv3���F<E��4��q����9�&�i�1]�V+���1*�1aLӳM��A��l��g�lPoW������_��+�$� y`D=���]�`��̎�� �<y�������r�Ȟ���4v�]C%k�O0 �`��[�<C��v(��/���]!��[K���,6���ńw�W�y@�ޢ��=
���8���S6}�U},�+l�DM�U�, [s��(s"oRA�&"Ga��o�f�H��1���N/D�d��;X���hiƩ�ƽ��s�]�ԆwK�7c�޻��;�V�ϣ��D��p0FO���<p�I�xM�������ȸ�{l�n,.p�4A���Dذ.�{��V�X��͵>�ޭ8�I�W������(P�ʠ��w���_����]]�0��Cd9 eti�Ӂ�]���♃�b3��'(ԛ��?�Emf��M�9b ��:N���qQ|!�nKe��jd���j֑_"�2�=s���'�h�#x� � �G�)����'�%�������J��dy�M�������s��5��$��.��Ĥz���GA��ً�g��ZŘ�4���L](o:�Y^U*��|�G|U��}xB��E�&�7b~a����W��C���Zw����Csu��["�įc/@��D`Dr�)>���g=�?~j����U	�9���L�=�ey��\�G$��j�H��ϱ��/�n�����K0�dt]5�l�.�<�;�>/�v2wr~�0mLI��Cn"��Ό�3�9�[��hz�0u�8۾K�M�����ЦX��{C��(����I�Pl%9hv��?X��ʛ��5\�c�KZ�H)o\)#H^剅*�6q��� �z|O�-��#S�%{fp�jCɔ�H"oߋ�����<�ɚj�*̮��2BX�d�[�:�dc�>*�v�:�8 �W�i���qAS�P�ne��i�\3�@~J �X�³�&�_�f�U�|����BH��M�ő�l#�[� ��JUj�Y9�ARc��@� ��60��gu�m�.��:�GQ�n���2�&۰g=L���SÛ��	<���>�i�N�z�D�G�Mk�T�_	4h[��_�6s%�yV�8Z�OT -Z���V���saaA�ٗ�O�ܙ򷜃�>��xc;��R:ߘ�ƉC���&��8�(& ���i�_���Xbr�8b�O�rn���ēE�+�"_G�#�.Ē��8F����5���X��^�)!JrBF�ec@�g�
�*�!6�PP��i*x���js��6�x<!K%��8rz���Q0��>�~F�d�R/�o�[��$دϭ�k�{�';����e�ݏ��he���I=�U���"��z�)J�� |�=N�Q��]N���G�Ǎ���iW�*o��_�H.k���ϸ�R�Ƃ�A�Z�VX�\VC� MT,��C�>�.E��I�	�Nw�nP0Y������zש%2�k��I�ɢ�����Bӌz�\�9:�e��
���j���!>K�|
��ז���KF������v����A��:�9���>l�9�"`,3�*��?_�q���b�E��9<L�]
�J[G'�-[�����=1u2J�+�V�.���������qP�� 8���`��P|ܦ�5*�d*[-���K5l}�A�*K�啔oM�2�R�ToP��~K��e���� �Ct��!��{:���R�N�^�H���L�x$�%W3DzM��U��\[�a�r8�W���&�7�پx�`Q��}ݿ:.A뼊�@�$�� ���,��:�.J7��(�Y|��܏�},�������D|���zB��ظ�ϗ��q�[T<��U6j'x*��y���S�x��c��-��+g�J� ��:�6��a����+���_TC$�A�$!��-DoJ�n����P�;Z�ڞC�O�B��O	�k�PX��g���v��Q�H1��/�I~��i�갆�?	U�ӑ,/�~h���T{`�����ΧjGx�����H�%�H��vV�S�{e��}�:0'񞇝*7	&L����f8��7?�I0�z�j�^�����,���@��e�J�`g6�-e����Q���B�7c�U�*���^�������2��\a��$�na�ǹ���j�V/�\��"����I�����B�1�v��R�GB$��{uʻ��~JU�~��c��^���Du��p)�*�7.Z�\«�[��E�)���s:l�>��u6 �q�K����!�=c�!�n0��v�% bK�E�I���GI�����~�ȼ�|��7"wm�:� 563�Ɵ)l����'�j+*(�����$^��
ڠ�l�� agD��> W�����6�Y����8e*9� ׿���*��o��%� p�|���o��!]��w��F���D;'���a�k.9k� 4z!e����`��X[h<�N���ԖښZ�!���l���y������ ��P���K�]�c9�Cy=�2ץ�KqpM�����I����ėE���#8,�X�U��o�������U(�Y~Q|x.^tL�g(7D:�ͫ��4��"�� �\w�r�;�,d�˵+���w�q�[X���U���K������C��.~�z���l�ҟ��Q������=?!o�i��4ᬐdF]��0ֹPO�~7>����z�>���^L�*�z��v����:���͠$u$���4E�}����(�����S}q�Q!��{�_B�º�m6��JN(�%�����U)���&R/Q氏B80�l�|;��Y����Ϛ��zbߖ�#��c���cJ|�������;$E��u���P��>Lc�s�j(Ż�i���u�5!���NL�:gzCK�m��X�0f �����[�/�Fw����V�����gJv��G�G.s�N�U���.r��;3v����P���H�46\c)�,]��4R��4R��f�}!��(y��\��Bg��H#�Pq�.Hf�Kǯ*^�ƻ��=|���u&kjQt��z�D�~�[3�{�M�0�ZٚJBO
�Kad�9?�$@�!����(��Ł[�_kRl�z��p�S�%_:Z(�	2K M�Ѐ�c�?�>(�x>����f"9�<�
��Z�GI%��O��f�s��@��g�о�#�Nd�@�xcD%��ݚ�j)�䎢�&�$>����X��_�����6,I �m1ߦ��	��9ؖ��GX�7����W�*Q�%w���tt\3�y��aU���C��<���%V�65�,�@��~�qD%�m3b�
4.���?�l��� �^{��rY����íw֒���UW�Jle �H��{��c�Ja�ҧl�۴����x�����`�7�_�'�4�hli!wU����'��yhT#s������`YV��ܵ�FE�~��lwZ��;���-VXݗ�^$�i|���3Eq�DO+�T�����-NN}�ҋ`�c-���9�#�3lW���I^[F��զ����b�����%d���~Kudz�tn�����[8��`!x�7��Z��)�2!0��J�jp<�����Ľv��ٲ��y�%ALV�IGv79G�'�m��Jg���8|o�6��=��_p�\�~$�5�c+M�{�>hz�0�\^�^��xD�{�I5βa�N��X|�K�¯�+��Qb����c/���j�%���(tk�I�ɳ���K�JmW%��g��&��b��;�WX�u�M`�|~�@I6�_�����XP���U�ɷ(t�F*�����j�10����gE�������qt��T~��ƞ�B�� �'F�|ygaH�C��#9�Q�\��e�8C�;�u�8��b��M{ZB�4�{��w �57�(w��z�T!�:��������GN���d��K��S�N�����D�M�#K S�$GԊ�Ug�ۗ��u�%�D���)�YFi�ʻ5�}ܘLn��9s�ݝH�e�a���\�� e�d!�v��ϡ�Cߧ7M�3}�<��/���ӽ�_(cTk����U� ,$�UR���e��I*�S1���:ޜʼ�sRq���(�I6�yʙB���W���׈���NSԜ|�X=2���d��*rt�,|��rl�@<"svM
R5{��R�}�j5�۷�x����塽��i�q�1l ��\x��]�3�a���W
�^�V��O���`I��'�%���,D��\�OEGo)[��'��>l��?�?nf��w�����	j>�:9��~�ϊ?m�@�fr�=&|!y#��� *���!���B��h�������V�P\dN��Z�Zs&4-�v��/�:q���SX�r��6|SŴҌ2e���Gj0J��#�&�!�oD��T⏵����
7��T<�L�o��D��7F��Zh��q�U:�����5���J�B�|)��TcѿE"L!�Ԋ�B�{ ���o��" ��>�F�k���� �]���o��^O.�>�8��S� �ć�uhky#b�`�7<�:�]N�����, kp�\�¤>9G��s	õ	�j]��R���R
�۪�*!����(��S�QܓH�I�@�,��B�lw�{os��p�F>�붓�o�QD�N��mN�F��_D8�����¢�9>�勨�n����BK�ǯG��{�~d�=��y��Bפ�^o�}���a�lI��\��tN�	�@ ��ӗ���a-�g����}[SC�Z��{~O�Nh*�l��u�wC"�,N�J�&�[��ns*�[P��%������S�� ]��8T�Gx<Y���=վ9bFe�R��aq;����o�$t��?������/��Ko�BK`��2�`F�������]c��y�����tk��j�p�o\'��l�L��Ms����r�4�4�+I.�=7���e�.y������Oz�$Omn�0+�t���{�LU� G�p�Z1��ҰhY?
b�x����_���������ɵ�w�Y��&F">�CE$!�H��]a! D�i��{���PW�
���!g5��˻Ì�R|X}w^2��;�*̉�Y���1��v��
�7�����Xˑ��\d(���9})��+�O�>�鼮Gwj<�n%\D�^�"B���>��7pt���f�%�|�&�)�{+�8���1��z'�.t���DƆ_�O�\��A��d��:��+u�\1ge�=��=�~q4CyK���JSިbq-��(��v���]���u�dKj_�Tw�՘W�H�����ȬY�A��6�����2�N� /`v�W���	�]�]��3�Z�s��y�e'�e��8T�Ep�
�f�&�
�xʍ����e�_.�9\��9!��)E�yE��~�^K��1��<�x�@���mڙ� 7���|wu���3T�4�N&q�c�{��Ѽ�$%��S���u��(��< ���m���h�Q���ب�{2��m����-g[�l��ò?&PV�@r����*�6�k��aZgP��UX͛���ZF�,��p��+�5��K�o���̈́5�ݗ�i��*�߯�J�V�M�'��Q;띈9Y�Ɛ ���ݜ=B*56���E�3ز��|s�<��C����V��j:�[�Ɠe�K� �s�ڶ�>�´^� �1E�x�t���UI��I`�	$��F�8u9����c}(zR��#����;w�B���/Yr�όlNyHx�1��7ﴰE!A:�Q��ӺV���S��ʵQG�}�-��~{f��꿰Bq�O<�����/����p���<�,;z�-�vg_	p�B�~�+O���#��LHNo��KZ]b�*p��lU��XF�r�h=+1TC�kI�;�d�n�$)�G�]����hn`�[����% �r2��}�:�U4��!:>s�b.=a(�-Xd$���p5 �s�m"mþ�e�uF�ڰfM}Օ{˽g���ڜ�k#��	�7��#���~�Xְya����ܯ ���}�?��R>槰�F�#�=���c����z�[���t@�����֭,�����GDA.t�5#Vvi2��[n�K&dGfشT� �/&��t]������Β���\�8T\(�=Qʏ&�b���p��'H���H",�ZķN�K>aт8�_H�r"XXr��_G�4v��
�C{P:_�w��f|�A��B�Wȣ�f+�nQ��sG%u'����e�LGUΨ����Vs��w��Zz_�������\n�1�F�m�v�,������R0f�k���8z�i�V�l?���4l|I��=�fR�}g7IY�w	�����g�v�tp�-�1����Ը�Z�kMU��1#`����O΀�e@��Bd�sF�bdr�h\��Px��§Tgh��u�T��$��՟K�_ �A�7�O�*�q�%/o��zT���K�8b'˵8&][���+�B8�[dzlGk�o}y: ����-�Q*��o@�:l0j�|HE�Wa�=���J���0e&b��:?���#~.PIw�r��E�_C)t\@�aB:���K���:���<J%�$I-`)|��gSN��S<�г���aI�l\����W�[��\�s��+6��I�U��ŷC��}�V\�QK�n�Æ��ƃ`�T�o�9W��]�-�q'{���?սL�4BK`�r�ʐ۪�z�&:fK�4�����Ǽl�8������h(�d��GQ���`#�@SLF�tl.i�O:�R)V��8��YQDU��cM4O��1��ְ�攎t%��Z��w�8��"u?|��Ұ��Ɖ��o�����0V�m��������8S	;J���	#1J��Ŏ�����efҘ�O�ߟȮ����+otv�o[]���jJ ]I����]mt�)+}����}�lz�� .W��,>l�Q��o ��6����Rr��f;�339�k�Z l�����������/\_v�`�:�����c��"�k����(!�^l�e��/&��4��m2�/F�o$R��O��/�ߢ��b\��B`A�l���BlD5��u6,�`_�#U=f&��E�
A�?6��w���ԯB�U$Y�͙9`A.�R��~O��q&��f5V�g�s�*���b|l�Y�_ "�m��w	�E��I2F�M�?����!a��HX�u蚲iVY(�'�mx	)���`�
�'b9ަ:��k�!+\���C���1JH'! ��@+���]�ё����{�Zpm�����X�!��K�����
����>�;�&H�[�"�e���=���r�
��m�k�q�D����8���IC��v�*F]D����o|.ɲ�
��1��/�-:��D���A"@*�:��4Kp�dV�c/`�"2L���	��-De�?p��B�k���*/�I`��f����#y�X<�3������f�\�Ȇ����+8�r����B�U����"���t1G��|�&
Îm�B���DOB�	�k|�f)W^F^Y�ZM=��%�2 ,^B�6ڿ�.�wo(P{t�Ħ�kud���"s-��2��D�xtf�������H$N{F_ӮOȠ�y�M�/���0���;�UYE����ǐ.�� H�u�I�`�m�ˁ���N�F�IՍ����v�/=��-;n�
���>�Ê�c���`*��^|�6�����a�+�k�FMX޳഼��X+�v��o�8���]�J]/�z���a$�>>���G׵B��OMp\ ��@ĝ�uWq���Í���=#�g��:���M�g���	�(�{nr%���m*���vk-�"CTJx�l� n_��i��p\��=G��)���G ���G\�M��8��@4Oh�y�`��~�&C!<̓:J����<Zj�_��t��,O�-9=��r�UJ��ދ�ۊ�g+�_��0��>y��Y�01��Gݵ�����uӻ0��ȝ
R���X�u͆H�xx�Y#��q�d]��ZJ��������J��u|"�%(�LC��#��{��N5���W�+�\@��<�Č��-���8�#�k�]M�m��-�T�e��e�ʹ.%FP�m�$�Ӭ���� _�+T� �n7�Y�z�vOx(�r�=�\#�mX$���}R����Rm����?���S�?�~�v�?��+��U�;�]V2P���׮[j+�v���#O�����������%FOp���h���H�H�XV�釙[�	<��E��&E�j��L���6č�����	J���������6�psj�=��ZtS'��Ӗ�gQ|Bn�Y�g�,'�E?6|�ht��s����p��j�����"(nH�8��f�xX�L_o��!?�lg���.�dkع��'����r��n�\�1(>��[[�fCL!]ϑ٨K�.$�0yej��^_�K0��������x�tz'��S����=#�����q�Ёn�E�[KӴ�oPU0�4��b����'/�����[� ��S]^���ӧ�"K�A����I-���D���9D�*�aq���%$l#2��/8���5X�c�|ƍ���yDv����i�t�
mH��2�Kе�/����V��^��/9�04HQ���>_Z�ɓ'*�!A�!� b����؜���;�po|`�s�%�w�i"->�� W'� �O/v�����_.;���� jgj.#�0䐸�w,�j�zQAvF��o�{8O�\�ɑ���ﵑ��X��kl ;-�p����:0�]�Lߒ�=�	@�� �D�䲁W��5=���G�;FkN;hu+r3dW��K�D�e��E���^��>�A�ãV�z��g͘�
���D8x�\W�rETD�Q`�|x��)K�'�dt-�k�`u�mG��qS�����a�w�.�J�����g��	��L�ٷ��(X��T��N�d�G�sjԽ�^*�`��k����ier/8�⃸�L�q ���1OX�f���4��O��*k���9�L7`1w�W�\�m�ȡ�J9�8���.у{��YE��~�.7�tWqC��S�X|*Pv��Ds0��!ˮr�dˈ����;��:��9���s�&����W���J�=�s�qg˂r��{�;���My�#�rexIڧ)'�s�g�ꅤ�f�#�f$��ý��zN�&�Pz��NZ��X&p�����,#���Ǒ:���`8�y��Zu��Cq��>l,Jeރ�6��w'��η��3܉�Bsk�ﱲs4�u�%�蜫�q�O�j:�w��3RK�q�nD.׵�8�d$ލy����Z��gd�4ʪ�U�/�qX��!���09ڻ��I[�O5цM�sbd�̈́b�%(���D��kB3��)[��+�ꬁ�j��G�Z�j�+�`�	������b$ć��H�b��Z�|���
�Ů��N퀇��	��H.Xe@��"1�_���0�j��@<qf����5��'���x�9q��]!�)�n�o���BAs���b�R�_1�u�#�C�F��#�1��m�%|Y�`=PZJ���yQ�x8q�D�W9��F���ʓΙr�}��q�`Y�e3,���?ڨDl �,%�:��l@��wP�)|X׏v����,P��-+g��x/(���r]T7���Q@p�۹�P��LH��;��_��������X���#\ٔ#�������	��<-֒(t�./s䲤[_"�z��j6Wt(��m�E��xBd$nY�2b~I�n�x><���e:TTͲnL''�&T[�珦Qf�(��G%N���m%nvׅn�[���!u (�Ep�%5F��fd���/ޮIʠ/��p���S�x!�T��2sa�:�B��:A��ˍ��&Y`b�H$����	�]_��kBZK� �f)��B�p+�G���m���TDs5�v���Di��!�d驤��L|�d��p�0ݶL^���������	�$#��B�N_$щm�	W�o/�����th�.	��C$ՎQ�g�Te��ӑ�Ʀky�r@���
C׺���l�G�F�!�G�6�P�v[��+��Йc�+�B���g|���Y:<�3��q���oa;�xC�r�+"VX'6��oY��� h���Ƅ���L]�G\���%j��P/��
��1goh��U�	c���W'ܕ[�2��ε�ɾ۫<w�j�=�Mä*�.�4d�%����X"o?�38�0;����`��ǆ-uE�w��sX$�%T�� ��CT#�Ŝ<j�ya"D�1,�NX}�|,����0�,�n
L�[��']�lҥ�gj�t�	�|�&��IӁk�˒*�/�˛�Ur�1�lU��]��fq�uc V(�O��L�Կ�8S�EZ�hu�v3G���j~���u��5
@�-����ӭ�6rM-�]_L}�Jy��>�P#~IQt,1$�����"�8Djor�q��b&���H��jv�F�_�ƨD�#����E��5���͓B��5[�c���%%��ep�����JA�5|#  �[�x��Ѣ�nOi�?�kG�F�t��9�2������=45��Hԗ��x��F֝��_<J�蹀y����ؼ���$sWi�(.�����);����feDO�� �6.Y �������`:��\�G,�tpz��.�Jhi�-���b!��x�W~����O�N~���+�/�G;1�����ϯ��h��v/�=�?�6�gE/��Z3�k�dO��u�$$0cNS�Кӗ��H������؉J��&��sB�Kđ��y#θ�,j$��˟�ַ��d�y��omx*b�2�ȁ��_�n'��3�.�;R��s�5�3>�c��ԡk�CAn!�H�/e��H���⸁��,6�雑<���jr�O��N�-79߸[�Ţ]���]�V*H:#�崤"Qz L3^w��^?��R3�Zhv��0���5֡�l�x_qS�ấ֭[*��;����L[�����
N���U����>eɰ�r$m�ir#���z2��6�;�}w	�CT��6A���u(�CK�� z�N�%���R��J��kB%b\�G�}J��Q�t����k!g�S�����6���t�C�U�C��w�'B��knzԨ�X�粠��Gܥ�s!�_�R�V.S�qW��l��\P=�|&GsH�+�J��0+x�S�Y�z���t���K��r��Տiƻ��((�џF��� ���U!ѭ�ܒ��Z-���㬿O|��W)��I����{���Ȣ!I���؆�!�
�%$�Zh��-)"����3��C&Qr#����2���Z3���Xz������*�J�����[U��Z��٭�\R8�%]�T~�����̓L{� ^ص�kb	������>k��+����rVҾȄ�B�842��(|�a���9j��S�����O��3���]X�� ��gL9�)�0�b#��N=v�B���@����311��E�Ue����=�ߠ���S��>�x3�M�6'?����/�ҭ˨��
�0��'S���&�s�3�y�,�a����$RP����2m�Iy¼��<����3$�,��v1|2X��Q��e�e�wl���M@ �?͑�����G�>�_`�VJH}�mДUqC�W�5�m����(����O<׵P�H]|{�!���S~$�i܈q��5蓅�0 |qQn.;�e~1�9�P㇊�h�Fo;*���R��~7�m��b=�jM��&H7E�/7Jz8s̹{�P�ݱ��6� ��q�;���=t�J�:
���" I���0a�*Y.`�X�7�Ԝ�Å��oq�:�?��!��y���ur_�{`��@���A�^�*���ՄCA�k�0 $��}��"2�E����ʖ�Ѻ��J>q���.�>���n+%��I�tҠ3T�pi�t�
�㵏����x����%��<�nhxtH�Յ4�L: ΃yoƠ������1	�vD��?T�K����?|z'!��b����YC��m�ݥ�nR�����\��5�[���.v���<����J�Pc9�C��$T,�g]����Х_z�n-�nt~΀���-��X��u��D`쟾�vu���T�ew��d�
Mk;7�
��A��t��+1c��d�g��+��"Q����~�C�ˍ�;���� B�yW0S1$��{4��_��f@��U�B��R��7���L��&��T�j�G7j��7�߱��
0�V����?H�z�3i�F�7Ec��h��_F>�e������H	@3�h�HX�]�tUAy�5ֻz��bA�ݠG�6�y��8v�ٶ����\��qM!����L�]�4]
����8�?3�I5A��i�+$����q�5��>���
���X�خ�a�m�|��q�:�*g]  ߸���ɑ����s2�y	��L2���?$�Ur�&�V&�vِ��҂g�2D���~U�h��H9g����P���ީ��^��Q%�b\;�TW��Hf���,ޚ|]1N'4��D�k96�5��S��n�<�4�Am�I@u������FZ�PsA���x�Vv�����,�p	��"� ��C1E��d9H��Ao��MY�Z��qz2�S�z�3]RS͝��u�'{"���tp�sk�Ӳ���<�%k���ee��}\ �2�DV�^��ũ�ԑ�Kf<��|D�[Y��[5|�� ��]h�(��,�sN�"�g��ev�ߞd�U�����ـ��H�[(KH�Vk��������0����yp����R���r_>=FǼ�pV��kI�x��_��s���\��ct�L�?t|߷�=�l�I�N2&G)�KT�w�Lp6[��e{�Ԛ�(C:�V*�$���>��l��S�0:IѪr�~W�o昲���!)2I}�p��6g�D�~s�@���KC�V�������#���ƃ�и�
�ǎ�M��ר{W�ۍn�CQ`��)j�}�i���A����w�^R,f�|l��3�rݬev��9r]|}����L�h���^d0!�-�T�3��"➮�1T�7-!��C�J|K�_�p�q�͞OQ��~��J�H�yf~�]
����^�N��^�>~��C��:[\�7��	V�ePb�I�hc�:�IŬZz�CO��G7L�DG�lأ@��}�d������Qa�R�-F�/ٓdL¦�T�@��q�);E�u�0�K��R� �,�Q��
F�7 I�V����6yg�#e#�[?lF�i<M[b�s�H�߹%D�ƍr��!$X5�n�iN���^<:HFH��+�հ�P景uc -pjS��)N$�.q�F~��G�p���9g��.�Ă�Y97W�S���ҫ���4���v���w)��7TR )�^�0G8G�{�`���>���7GF b��,˴s���玸ྦ��-H�&oE�nn�Z6��l�-	eTS���s߇����)jR�/�h�P:�4e��&,V��	mn=��Z�g�7��f:�Qq����L�������p�p��)܉Xޙ@���ҹm3���]�}�f!���0kO��Z$��`���%R����7 X�$��(��|^�N]��.|o2N2�}8��mO�ظ]�r���<��8�Dv�7����3���..�����*;Ȉ��1{ f�R�[��*��}�lFg�#�'��a��g�Wk}�v�H�WVQ"%<�dY.��j��c���P�u�<}���^�yQ��$��!���}��@]�E����			�CT]���`2��=�i�6Z�4��X����=�\��{�|<�.��)��?H��������e`� xC^򭳿,���*�<��A���i�7vF8e�!?ݴ~��@n�}>����f< 3~u����<Y�Xe��|��1�Z�_!R�ty�[_1�ET{�*�O����ݣ�ɝ�V��� A�gEȧzd�fAb%�����g.�T����>�˺���4�P!�I�����K��m��D���)��u�t�j}�L�'���\�J$�� A<iH��嗪)�}�K�	8x\�3�v�W���?tG]瀽�(��(�ר~��z�h���PCp:b �i�l���4�)��`�1֚��1Q!$H<B�C�PJ��h��3]`Ԟєף8�tk<� E���ڳ]�����N�J6����2� ���޴�^���j�-
%!���ݰ�a�m)��c�$��J�Rʩ��E��
MW���ﻴ3[�r�)��'kD��_gҎ�cH��M��]h������ɗ�3f�֌>/����07GU�
N�ʶq�B�����E�A����]H��%�G�kB�6�j��a����G�V#,OV����{tql�j���K/l"Z����#'�W�!�ל�C��ӗ��f�s_F&P�g�ޱH��gka:�BQ|�p��Eъ�Ncwg�a�kg[�j�W��uƚ^�Ohӹ��J�Ъysr���AMYVs;#����(d��I/��ofqpk��W��`��~��b&&L}GnYR��皯�B�aB�F�qv�X餖5��;ʪ���rn������t��lşK֍�]�1N]c-f�I��
~�pv��C|���m���e����IbB��A!L^`��l0N+�N߮1�8ި��,z�,����� �R�R�I~�K�m�n� ��A�n�<aq����c+��rqp�0m�h��FE�ܭ�AJ�6 vo���~��ڎm��8#W�G'h�Baa�"`q�������4xRRF�(m�d��o��ٓS��� �Q��m��/.?l.�-�?��d?u���d��s�t�3W�c,'���^�ѵ���R��a���8~1�V��f�MǎC&�pP)�$Tjt�I�~X�Z��d$#J��?B�5�@�F݉��&@��>�>�E}X��O� �"��#�S��TF�6t�1[e����жa|�E]:>l�{���1���oe���ɞ!�MYSN�׉15�<̯�0R��o$�0�+�=dC,|
a���	kwv�La輇K��S_㚆P�#��=�  ��](��ʀ���������T��i���)
���T��3�|h�����D���+fk�b$�P
�~e���N�_��T��hC�]�{��~Vg�iR�fQ�o>#�|K�\`T�D�#D*�Mé�$e��O����J�~�)�����G���4��'B�����'�ϞM������$�Ɏ:l�3�ڤ�T���r�Z۹M��P{p}���"�7Sv�)	�
��+��n����¹�d��R��Q��d=E �}a$�ȝ��P��褦��8���L,ܙ'��"s���Ku���H�50����Y��z e����Z��aW�8e��.p�htS���9��ޛԔx����)f��ʥ��ᓔ'��jg�q��iS�������0�˃s���b$��itB_uQ�2�#vK�_Ѫ�<�F?��I9>��<W�NUz%)�^�i����K)pT�']���~ׅf�?���� ���rq�ڼ~8ڻw�3��+�q \���`D*�L�!?��P��w�=�>hb�2h~�ܻX?��g�
�WN~�����Sp�ltK<�}`�A���U�u��?��&H�	�>�j��W��j[H}:UC�9���!X��F�G�-���	�����s9B��\���o�ț���B�ra-տ�Ri��36�qC�s���j��z���Q�k��a!��ր�y� ���p��>�kB_.�*H�"���4���c����(����JR�U=���տ�D��t#�� ��J��>tV�w��U�@X���;�I�Qw3'��[�hh�y���c�c��2�1�{����"ĥ�B��4i����o�z���#'0v���[{��d_�5ST`g׏B�UǞm�K�7�Y�D�P	r$���#A��Vs�0�K���s�y�B��D�qF�
��e�/=g�/C;bg�'�֧�������+��Q��� ��c��v����Ӻi�by�U�I�ܕ3��ΑSn�χ�q�U�������aK~Q=�:P�RRD� ����Yqi)%n�{�͖��r��7�r]>����R��&T!,:PcO@޿Q�-�V�M�fQ}�+;����g���S:����Z1O���بƂR�؎,X����ᛵ`q��0�e��<��œ8��6��~��?�����茆���I&�r�4�NM���#
B�׻�)�VH�0�Lc`q7��cR��� �:�l��Ti��(Eq�Z)��*�J�&b�!�������h\����VV)§�F1���F0]n;����-�-�.Ѿ�T��y��<�Iz�kJ����?V6�D�o���wɍ�L�fk%:?�T%��F�o{B�ήGò�r�I���%D9���U�1]�l�+!�M�}7Dl!� �&��N>�6����/Õq��?TEU�C� �zH�){��X�sA�����JbNق�LW��H��x��(�y��}'���`L5F��bCv�-P�di+�ٶ�с�x����vE�T�k��D��\�G�tL����� L�_�}��7�$\�V��H�H��@��]��7J�MXz%��L&�F[6}>��7���ʈ�p�/C#yХ�&/�=��6%��D��;.�?ڷ�g��[<�[e5 �����#���v 	����Xt�U�� T�ܓ��ͱ�OhK*Z�o4�8��hDp��珰�u{w���$U�pT8}��RG����7�O۾KQ`1��=KP&���VX@Άs���C	[1���X{1-G�l|�y�Ъ1D�:� ����:�$��!!�H�K�6-�*��o��K�
�BJ�'�.R��~w>��0�>��{`\�6m�kG)ü�$;�r��yL�zP�W(��6UEą����݊����������ӝb?�}Dl"��>�'��]z2�|xX�?�f~�nCZ�/�t�zf�":�մ�!1 _(�?i������*��Z��%�9�d��Ev����@��F,���õ��ϳ�L�nYB90r�uX�Sk����v-r$�5��'��C�iM{f*���x� ;^Q@���VW���\3☼ɘj/�C>Jp]Evg[�2��21�����nҍ�I �R�]������?PQ�U||�~�v-+���6-i!�2�cKA&���G���#�m�|V�1��R�Tcvd��U�N��\6ä@��l!O[����%IZdֺߟ_�o\��E/B���I��:Dj�G�Ψ�a8)1H����:')�X�#^*�F�O�yQy~E B�i�嬾������9����$�2�g��r9�6�R̒�\WM����'|W�n2�dBh�x��{ W�)�G��=#���<v4�s�o�!?kIU���X�#�`[s1�>��M��Ք=u�oC2�[A�fr���g*�v2ϕ�y�Ϡ�/��Hd^����I�$]����CK��k-�;��>ũ���(k�xI�.�-�Hb.|{�"�%1Q�x�UW�Y�S���%�^s`�����A�ܐ�n^|��ƪZ��JÐ���9ȸ�]�b��`��~�G�J�u���<U?r3��w�ګ`��4z*���I�u�_�H�"�5������B*[����`Y�"�=;vOU�T��Q��9N�Y��YT,(R>��z�vY�"�I=��?tc0�ǚ�����%B[X *`[o���V��]gO�P�X[|%����_ ��}D��{)�2������x
"H)W�!Q��5q\���
�u�޶�0���LA��-6�hJ�U��� lT@��x&����@�}+�_��O�!����M/S�/7��(����7Օ�Bl׼\im5a?Jj=��Z���AJ�ƨh�jd�_ƕg��!���* �D��@SY�H.�M	�n#��E��Qa��t#ƫ�i?LrQEjVs�%�<U�.�VH
��#�_Ӥ�'c�3eN.�}m��Lâh^#�V�~,����D]�_�l��eA<.�5�2��^�6p`�oI�r&MwtV<���$�3��A���J�0E�Q�3l+,+!N���>�y���c�\��
���Я�ܮc<A!u0^;Niӊ�!ZwLl��:��Vf!� �{6�U�U��xQ<�T�Ǧu-HRIk��V�O?�4/H�ݮO��*tCh���q�Q�M[�g SrZ���rT︇gl�s��H�F�w�ju�|�|�!��DP����x�g��	t��3{EƘXd�e�[�n�����*���.������W���v�;� �H����ܢ��J'Aw~s�6��I�،��E�Sv�+I��]o�E�b"x�Q�����8�GK|���S�l�p3)�#up����p��_��`n�It��X�w-:�9�?~u�Dc�W�~/�&�V�u�Ϲ�[F�%Ⱦ{�q�u��'v���j��g�kӐ���Z�9�ٙ2n ��69w.u|Pg�})�ꖚJ޻���%u5�>�>B��j�eԊ�e�`P �_R[��S��_��kC��ӣUtFy�
1&������a��N�q��KѝH�'p�u�y��S�o�1�Y��{�'U԰X�FEu�a���g��#�hWXqv�-׃%���gݛ��/1��W���i�bVV_e!W�9H-�`D��@|藕I>(���~i9�6<��� ^YN`[߾'������)��f�q0���V@sP��1��\��4v4����=��*Q�� �2T��
�6йS���� n�v(�xeo_�U�!{����@$�&,�j�3�tTX���U9W/۩�Oz?�f��x�0��;Ԅ�K�@��x�ԾB!�F�����UK�H��B�=V���޽&y!~�Ř�la���q��ޱ��U�U�v�(4�S�X�Z|�,��p ^J��1\���L�z�n�Hi� �庆J$x���,1Z�p��>�v�w�t��0��#3o�=s�S�yUӚlR��Z�����G$\$���%�	R��.��oT~�P��VH�Z�/G��On�R�i�Ƕ3jZK���״��'N$*�6PSY֤�p�pU�I:E��w�"_��T X *�Yp��� s�EE0��t��z��u�9���`�ѭ"�.+J��֟�:z�+:Z�����M���.�k?���$���Kv��)�!���%�
b�Q����Óg�0�c
�P\�x~�6�z�A���ص���/�l��z�-va~$�@_:�W�W��b$�+hid)�����ue��C/@q2 㼹 +�1��9�}��~��~z��+o��dR���V�k8���t�>t#��� bO7"�ʾ�FZ���6Kh+��
�.�K# )E������#J�������m(ݹ��^e(`���4��!(}�X�S^wnI@�fM����6�|�8S(*��U ��o=���,�bW�{Fe/	��f�I7��q�����M$�:��Ɂ��l<�d<�u���X�L��J����7�Y(�K���_N�Ley�^}���n���$��I~?uJdy��n��F�6)=~�����moԢ�9u, ���d�C�C�Jʚ+'�&FQTW�e�qA�9�-�I���2�ؒ��S���?���b|������Kv�* ��Ӎ\AM�ճ)���Y�
pN���=ӅȨ�k��q��k;b�Ƒ��2D�fL��w��$�[q*\n���k�ɾO�7��Ƕ@a
�Ğ����vz�;�L9k0AL�����s#���,���du����I�2�.g���Jւɽ)y�~�f�B5�� 3���ƭ����N�!Q9ga{��1�#�F���$�s��
����n!��A[��F@��>��AL�<%������؆���:�,�	hƱ�y��V��2pu_��<��('/#��������#R���+	q �r�e���uxSp�,�8b2�Y��@�	����?�3�x�Ds�`�� �Z�����l],�UH�p�O������Qݰ�pv�G-����z��=��J�3Ĩ�^���`�]�@Ҏ�^M��@	4���_U*�w��/s[�����=v�@�k�9��8	���2���0D�M�B��Q�H�j<�^튏{��K#��1T	��lS�h��ɴ��xH� l۩'���{�g_v�a�'�@����o��B^UL����=��\�����g�l����`�
W�5��>R0�7�Rx�=�x����N;Mw���I��wf�2N�uX��[�L���n�D�ֻ'd�9uLJp�=��0os{G�|�z�O�Jz=�@=_��I�>���u�0�-�(�Jd�������Z�1R����$3&�x@�<i0��Pǂ�Y���̽��H�����Bjc9�ls�Q��}�6��(�4�G\Є��a�Q\�� ��\���_`�~�	/<��1�mL}[[�M��_LI�F=H)Nj	J$&�`:����z��'@W��d�*�mr4D�)�)��B�2��S��\������7y�'<6��|U�2?��}LIؼ9~#{�qm�=eCw�j]�w6��Qg�}�L�2�s��F���@�����}*���RLfi[%�vⱄz��C鏽�2�U�TX�D�62A�	X�`��Z�`�4�ʕ�h5I�ޅ�va]�js	�x�Ǆ��>;�~�.W�����2Kp����7tQ}%&j��~���9%DC1�f��6I~������4ޱ���M�w��y0��&�w�\�C��f�:������\����������ft?�ތ�:�t�9�=~}X< �@o�Z���l[��
IӍT�� �)F=�/zh�*k���� �ŵ��+'6�[�\߶t��Ei-�W7{�웷������N����9Ф%B�=��-?W�r�V�.��W���@�s�=D΢Ƥ3�*)��?�W߫`A�1��~[�s*y멁	����ؓ�#��&�r�����'�*O.����[�С����X�G�����lAV�]f�AZ�ʠ�9�KY��((�����΄�A)�������A01|���X�a�T�%êlR>�k��CUBd4�B�_�����|.Mt+�꼇�(��t�$���~��˪�}D c�yz�H�Nv꼃��b��- ��^�9�r��(��UM'I�$���כ��A�9rAs�QO���U)"o	��v�^�l���r�G����Hቃ�չBI�/(&Ll)g�Ex�J�[Ao+��b��։l��5��-�W:�X#6�y�67/RB���۟;�8�m�Z �ՕU�'�!
�H:'G�]�J�@�	���>��FܟBx�"P3K%=$�h��h���J}(� �kFN֑0�b$F�����fB���4F�<8�R�6���	6]�ͨ�l�� Z2Ջ�ThS��H��):tr[�?�6�۵Ƞ� �#�>v��rƶ�#�\L��* ��U[��K�ۘ���Vp�k]>Pʑҷ�k�r�Z�
z�g�E+�؝�2�
�� �:\��.�y$�����c����D��'��|��JJ��x�>Ʉ�]W�A�3��;u~_HIȥ���u�K���ؚ���gD�P��K,s���b%��{(�*�Jω�I�.�}��Oα�K���B�EH�a�B�߮������[ۀd���Ɖ���
�KͨF�*�_��6,<}��=s���g8�8 �%��]Ly-�}���Tv�Z ��l�ܮ]F���1�Z��^�1�4� v[S?��z�,�A�!��U}'�a����g�$$�a:6�anDk�O�|;p�W7��������-q`L@:�:��� �p� -Uf���.I�+;v�h�)�0��>0�a�ݩ���l�L@�r	�13�X�tAA��)`��3s�9�æ�Z��]oz�Ƒ��!(\x��Ϲ�"`����c`�>U�9ٛ�P�sv� ���`z.Y�� ��a��$8Sw�����ϰ]�>AW\�$}�TX��/#j��z7g/_����9�m�ZF���<)�9\�P'(��t�'w�a�6v���G��fj�G�wO�6W	u�I�U+#+^���7�o�9��*>n�K���RS�|K[�{J�V�	]��v�\��^+!�Bڦ�3���h����3v^����h��PzeTh0?���{Ƒ	4�3׷t׀5
�)	Ƅ�R���v@ɛh��Jh8+b]f�hb��N]���'8���lܰ�"5��=I)�5vY�����L6����>�hMמQ�I��a��Ă|4�a(�F+j����/��\ �B���.?,󃧉��h$lT���ܗ��/�&�ݰ:��ߺ�2RD>Vr��g�\�NB��7�}5��ʠ�$�UѲ7�,��g�P%z�+
�h����xT��;��N�����4��y\U����R��'ҧ���!��Y'��v&�j�Թ�uҁr{B<c�-��ْr�y�0ˠ%u��M�Y�܌�\�*h�'���9U�::��z&���G�[W��q���S<��1q2��`����?e$�p�T 5o0�y�0��wD�ܨG����W}�$��x�T��V�]�wf'g����}��X~J��AS�2V-��i�ķEm6V>�����$��ܨR'��>��q�69��J0�1aA���O*xm5̵eP�b�_5y�u�� �zƇ(:�&&�_�U�Z��U�YlpR2��G�:��䫼˺����M>/�v�q�3X܀�y<�zA+6�5}���m]I�X;x3m���H�2Z#l�J�M�)#u�u�.��1=�-��R҆��D���S'���u������F�b���O����-ޒ��v6�P~yy�7�>\g�V�i��'�V� c/&�EO mZ� �~qB�l�A������D6+�=�R>�g/�
��Q��A��q�������fn���b" �n�����b�L�\�U�!w*�A/��ݝ;�J�D��B�7SZd�V���Q����e��m3�n�x�@���)]��A��ڠ�(�CI��jT�M"�{7���@o�2H ���>-'c+�#%��w��$V��� F�?���;@��a�:�y���ቧw �q\��z�2j7ռ����R����^���F�1���G�y��s_�f��Q�NR�;'I��sc/�31i�q��[�9��=��0�3������R2��2=� ���f�k"׋�N)*�?g����i��ʽ�{��X ���/is�!nk
�i��c��Vd�I������%'ϙ�Oq^�Q�����n��cɆ�����k=�ǰN��CIF��o�)�=�6|�N|W U�W�ʹ4�,=�����Q��x��퉤���6CI\djd��I�Vl {�_8�6C�4�Is��ޗ����8Y���� �����AL
t&���U:?X|ca�c2X�d��0�^o&������	s,���Ue&o�M�FJ�Զڥ�[]w+��KơCe�;�)n�K50cB���p9[�r,����Ge|�ʫ>e�T��cБ��l��Ce ��Y6���8����%�]����)F�f��
"�r��e#����g>��{Y�V�)��
y=ٵ!;����rH��ѩw7ص����]����gU�8�;��|MAZ�W����[͎���=#b�^�Ye�bݮ�����u�y��"\t�����W���2��6Ո�J�G�E{M����T�
e<M�z�9��> �.�ȩ��/#1GF-j�jqe�s�t�!����*4�@aη�41�a0�m����o:��+;�1��@��eD=�,�\_��'P튟���Q��\�Fϝ�MA༺�rsrЅ�=�&F�yZ1��|/A'��F�M׻z�|��pA��������:l���kũ��o�����l���3i(�w��cXl!wi���K�H�z�+�d��=j��jo��wJ�Z�����!�QL.}OCV��:v�߱A�+K�s�w�H��Vy��H�\)Ą�l��C�MM�v� �>wR��[|pk���T�Zۢ�Y��g?&(���8%�-���,���_o�`�����ŎA���Q\q��>�"9q�r��UA�ԅv���h���P�b�e���V5�:�@Ԟ̺�-1VO2��>�K��Z�{��X�5��B�
�*�2ܑm�8%ܶ%�wz�5�?-�X�{�e�� jπ��S&'���H���-�
��=⢭�'I��״�?G�@6�PP�3O�S���D!�YY�.廆-�ŭ@C�÷S�+Н��Z6-��%�n�ΎN4Pc��B��]4P�m���Ɍb��˷R��a�,;26��.��Z�h�$p��Hx�߲{O��-�FPg�Cdx?��������;^���Ⱥ"c#�5�<�'N$��Y�ُ�����a(@�wuSL�As���@d�^��S~R~��*�)� �#��~�),%��/�� '����eŁ�"�T�Y�����y��(�R�m�qd�jI��''�;~�����D@h$i����`�0��9����+����7�Z��%�IZJ���cN�ʱ�2Oa��R�t`6� �g�j�Qr�}�����L�3
���������-���F�:�Θ�uQ|_���y��g)6U����x������F��S���W�M�me�ѭ59����<m#���a�@�"H��1S|􄏊�]7b6�N�(��I�å�����O2u����
�f����j3kn��{�.�$<v�viS�??/�R�i��ɯ��R;V��&��L��O�z��^�5������CQԀ�,��4��g�
�
�@�������0����hD��Y�����s�g
�̅Q#�_ʧ`n�w�f�oL^�Q�D?���Z ���BP����֩08i�X��h�P������5`��ѧ�Ei���1JU�2�������r*9�oN_��V*[��t�:xb;�+������|���5�	�8�Oj��(c�'%��b�)����W���qNLQ��I�c����S��4z�%F��������B�f�lWE���*�;�jF3I�"�t����>ܽ�R�I�s������X�����B>&9�+w_��2��ԟ
�B�[���9���T��u��9�6���_m��0��k�%����Kʱݡ+�ܑaSU(�t���>�eOR�02�>w�Jte�8`�"��7���\���y�'�J%)?��`E�n���e�� V�x�1g��X_�8��8�	^)�}��u �#���w��'� 8�5��ޱGm��Aպ�.���gO��"Jt,'�NJ�W���%�G�
I	�r���'��r��'���,{�rn�#�G���w%�{�wP`?�*�R��P�)J������P��=4�����C��������Ľ�e�T�9P�aO2\�ځ742^�+�\q�f�4���2CB�U�����<�=���}�Q �¼��l���,ҏZ�ZZ��Sn�W:by*)3KA8j'�PfX=�K�Q�p?GG��8�Χ�jb��������^����K^��O��3�������s��z������������㯦�?��#�̜����7�1>��Z�Q5 VU�9T���=�Q�q�o�Wz���yg��A��B��@��k�0��uz��p�л�=u���^� �������Q��w�p�1�R�ZU�ЬN�*�-a� B�1^�;'�z���?��(���o�����3��,�D��}D�b��Z�{̐F�A���C�0�L�f�8}��}8���(p�Q]�a��S?K����yu��M������b�2��h����.�]
�<`:6�����i&��A�� �
j�
��YI��#5.��Ճr۹>�hfgF�0�ǹ���[��{�"(& 2�V<0R���<���E'L�s��hicSri�� ҙ�đ�9D�T��3�E'�p������E����Y��V�|n��y���������� ����4�\�dVâ�nZ;!c��
�/�,x��Eg�-"_�>��Ð�giSbxHl��hS��X׿^7��d�'��|O���"b��W�dL�x.1��?mݾO��ῖUj��0��Ku�6���ӱ<8����E3��l��?�k��{E�Ą/�-����ۮj'�қE���4����^O8�b�V���]�.L�j�I��%����X5碓4� �H�Ŷ�?8$�WA����_u�mW��2�=�]��4��k<踅�]ڷ�e(*B�K�} |�ZH��E�P��a}��ǖG�㄂c#��s��F:+\K�<��捡Ȼ��
3䥲�Y��Eߚ�z�{��q���߂a8�v��l�h�����LY��b��Q�ٺE�ג���Yk�o&�3:�/?�g��rxE~Ѻ1c�e�e &{pg9���^��r�`@o?hW�.�>LT0�*:�*
[ک0NΕ~�l(ZL�Q[R��1`Q~�ͧ��Q����d����}Q)�%x��蠖4_8�1 I1�L=m�0福Xx���F���
�Sc��ր���b�'�0%P�@�ʵ��R��WԱ��[5�P��V�@��?�Wd#$7>缏z�\e����n@�����]�=/iCMw�3Ԅ��e�A�xx aB��d���O6J���w30�.f��0l��#{�LY��U�����G��J�A����q�Qrd�+�0l��H��������z�������Y�x��F)�O��×�Vk}��έw��)K��ʬ���?�>����ʧW<� e��d8-	 �,l-�������u3j�jA�z4��p�	#�xO`�<���O']<������n��%{��iu�-�CϬ�~�j^��������%����Aa����vrs�yT椔,Z)���%�@����x�f������@�?�>��4N�	�Ʈ�Ėb�}<w{/�A\qOk9�f*d�	u�ٺ};�>6�]��\.˧u�,��C�]�<�Y*�?�HK�!,��y%�u�	(�a���Q��s��~��5�Ǭj�4�B�NXB� (��z��D��KW���H�п�n�.�*���-��ײɓ)I �,��Φ&�0I�<�'_|�#t�	v��2a�b0�����9`�̜C�%�*)�*���h9Ҧ�C��jH����V����!��=syO~�����戁^l?齠�.��!x�\�U�M>X�p$\�N-XF|�YUoR 6�B
�j)�m7��!�-�i���<I�~�/��ʊgQ���B��g���t�p��@PmV[uL�w�U�����d�h3	7��d{������ώ��#�:!����u�@1@��
|�tSW@1ϵi���L��$?N�5G=&�<x(:�mh3N��t(���M�tXA��2�=��ȑ�<�54lL����!�)&�T���I�Y2��X���L�Gv@���PM3�!����P�G'h��Gq�Au䗂IT��}l�qG��4�r�R��6a�>��b�^�yZ�F7��;����������㽹�S�_�]j��Wy������c�t��|�yW��]f��W
�	$��g\Tx?�����ҝjɕ���n�dV)�ߎ;&W�O�e[O�-k��0�+�/�@�@H�o缏� �������Sc�D�Pu�x��_\�+9����mJ�!:"H�{�Vl`LN��s�@�q��r���R6�H];:F
����:�[m ���"@�-]5+m�8+{�3$�Α!�����G/�\�~򄛵Eߠ͋˿A���[����[HG�,��X�6�D�Є�Ȩ���!s!l����h��X��U�Q	)��:r IM�,�9����u���"E�`weL�S�@�V��������L����3�l�s�+B��n��a"���.��Ajj�NoC�ɬE˔k�+�<QB����+p%k�R�ܒȎ�Bli`�z�j��d�D�+?������3�B�����������sX�_�dۯ�������4�Ooz91^��|�"�Z�c������5�,פՂ1%2�	�Q��*o��L.6�9�X��OT_]�U�4Ս*}�rO: ���Zd�֢��52���oϕ R-[�;݂��pJ3;�AW'��}�iP���Y�k�Eix�} d�u4%ʦUau7����Tی~:��N"-�R�ه,1����KLx�,����a�aD3**^+RT�v(�Ib�CS$t�z}ٚ
+��~�	�M���y,�:�Z����y)��Vm�Z�
\� ϔ�HNP���a���A��x�nePP�_^fv��Uך!⊩�uz$߿�(�=�=�b�Ҵ�O��&��2ޠW��˃��
� �HzJ�t�Oul���r3�	ɤPS}��j(���+��;�~��t�[�RH� ���&%3f���m�f
*�o)�V��g���&�t�Ow��W�]	�L��c��,CQ�L4rY�i��y��3Gߺ璪�=�-n�:D�?-�l���_4G?\_7�U.�*���sF�<=��1���v��l��,ޚ��� ����2ذ9l@E�������F������Af}	�h�L-�6C؏�����O����Q��t��#�x� ���bw�����+N������&%[D�g���	� ��g�����P-ΕqbP��g�/�I��ut�k8�ļk&�u���[����>���yĉ�9�#k��j�O��X�\��_��a�ƣEK毾o�խEw�& �T�=7&!�G�`3֋^���Q����H"��I\��S�i���F�TM�d2��|K�uɵ�v���m�B8���R	B�����vdV 4An���7B<���P�)޶�J}g��n��F���+��N�(���
�W�/��L^+���A��>���L�@8���/2ͅ�[F��#�=]��@��������=�jFW� �0���k�jr� �}�(5���&z����e�|G�����٨�"q�#���D~�����[􀫜�t{���-|uo@�ǛҖJA0�����j�'�*��̻W��Z�;O��{����Ȃ	?ƣ�aED����`L�a���*�￞�|�q	��oE�!�%gYʘ1x�y�4=}��!6ȉt�:�Ŭ�i#�>1�
�s:��;�E?���ph W�J/�È^�E�&�~O�L)������KI�~��c[���e�e�7��(���žM����Ԫb�[�g	p�p�k����U`�/(�(���vg�����1��{�	������p����ǁ@1p�`�גu9^2��\�m������N�i�d���&�N�ZtpV� ����Wz?��ݡ�1��K'�M)21�<����mcy�=�
�^>?������`��2P�ҺR�\{HN=e�)J�)�˯�~�g�*��@�֚!�'"�D���,݌�����Fje㦃i�˦n"�;�B�<k���l��-'�����A+/<�y͂����Y�!� `�Bq5[c���	���bK�jՊ^Nf������j��(nޛV���i� �ҪG&�4@B�����cÐ̷3x?�T�Ɨ�P�2��g���n��4�,ݞ�̡*y}�Ϧ����?��=b�V��]4��jO��d}Mc�d�\Q�;*�1�#�� FW�wOR5ס�+5��sݽ���R��隨�@�O�`������vEqx���]|q�3�.�>��O�]��
��>n�sf*�������.��9?��{^̴o'�2=�c� �P<���� �Us��y����M�;����Y"	�q/�kMY�2�o���|�|�X�AA��ʳ�L�|^�=����;P0;�/_��RO�9�-��L�u�zQ�˵��:d���Nj��-d���~���BNp;����C���s�*����~��C��:��o�D�4��)�~Ijƚ]Yğ�<�Q��٣�P�@�S����^_&��}+��
+%��yK	�3O���j���"2:W$�p;'��zB����P�h��-�8�9�,7&)� o�9�[��O��Ŵ3���P��s�,9���~�̐8t�+��W�c��ps�_!���>p��E�Yx���]z��y�8��x-���\�J���q5̮0?º*+�]�E��:�	(p_.CD&�7y���[I�m�~��>�]�A_�'�Dd�H8.��vn����qk!�{A�Ҡx�����/���v�<��(2���Y��/���,�0��BB0��/a��C}����w0�4��b�W����qLM�/&-Ӭ�����nNo�<N�	9�Y��O�nx�lMу���,H����y�HN^8X�aq:���̄�n`M�sb�w�Ѕ�q̓7Mz�
'�[�+�u�����/c"(�o�/�j@�:��稢��̒��G�-��:n�w���ڥ+�G�گ@w~�tjZ(��6�Y����GD�xƷ�v(�s�R�j��Ѣvk��o���� �|�8���hS��7�y(!�W��:A,+��x�T�2m#*��?A�?����1����enb,�V�Ə'���7 �5�TW���XhB��B�$�|`l��*�2Y?���?>`%�O�F`�����S7�y{8��RvV�,��o���Ug|��p�ݾa*\��f�($�Oc��u�Y0��c�x8M֊���:�!�	�v6I:S���`�|�%���X��$��zrI����}Iɻ��a��f��Q�j޾�M�<�JH�����YC������uR�{B�;�B�x7h�ܖ�9�'0�	8V�]�g���E�jhR�t3,�ߵ~�-���X�K����w��P�6N��"!*f�ޝI�tN�0ނ�J�N�`�yWU��Jt��-L�W$�ɨ� ��ġ�%��<Ҵf����
�	�{��S^$E!`"c{m�X%�ՙ�h�$�v3�28��|i���T7�'��J�7���h��$BD�f��/�N���[�	��#�I��9�%�V}-�D�����<\��ZV�I1;�T�̓J��r�DXo&)���>DQx� �w4���tpKгn?az)OR{7{K��"YG�2@�N���+Gxm�i�ʓ�'�o�-�oY��"8��%LĽn�:��(+~�{ϗ(��ށu�/W�:�e����V�=��t*\���t�����>�]rP!�dŁ�0��'�[_exx�tn�Ȳ�����Vo���^����tVd2B����.��ހ,��ji�L;۵LF�¨i�����Q��	�K����H�h~��a�A�Ϫ��f�;G��F�Af����T{H���':'}#����?c�B���nM��:6���#u읏/0�/&q�[�Kt�4����i�|ɻw���g2��2���B��Wc�Qz9im�.��=���s¨��6�9�a�~���v�S�/�+���Ѿ�}`�n��,̴��C��uϬa�Pc$lE�,�M�Gh��[?�秭��N]gD<�N_ϾO� �%bB�/}�� � 	_�NDl6�!�����z���,*��������~eIּN��0��1M��yW<6��xG�5A=N���O�6�U�
�P�w8��]�bX-��y�xZԸ\��,�����>ح%\�K��kD��Z��RN�*���<V�%��+��%#䷤��36��\9a���HR�B�_L��Q����>��%��W���fYU?���V/�S�}��{�(�B�Ű*�
���}��8R�(��|Pl�p���*���A��O�B�9�j]��q�'��Ol��~ȇ$x�����c�a�j�Km6�Z�,����'�c��/a���v�ݫ< �
GS�Xlz�ez�M?�Z:��1h�.|��ѴAckZ�]�{l�Ce�pyP�c��	^g�O���Rj@��p���^g2W�D ���9����?N�Ӎ�=/�T�z�"G�89��yb�3p)��H9&�i�����v����E!8�8UA;��lpv�v�X�b5ȗK����獄�!Y�gU5*@�w�8B�1a��*r���B��i=Շ~����T���*~
�e�,�]��$Lw$�л��N9\(<2=s<g�e����"l�2ы/.�"�q���"�����6YV�в��t�081[���,�!R�x�`J�^I�v��ָ����\�7���Sjz����\�ؾ��*�|k�m4���!��6e�mav�ꊶ��h���7)Q����s@«��m/�˾5?��1�^�u9�)�;�ܻ�7�7jb�d�6�hrI�s=M��2x�m�F�]�ì�dF�l�L���SN ��Q���{�a��0��9�����uK^��ht�|B���1�n4O�e��j�g+����[hl�i����Ԟ5���ѯ1���L�ݱ/DE��Ǩ���mJ��^a��5���%�����*�� �uu~�R�PØucp��S�};J����f��t�ї=&�]1+��iyx�dI�R[d$�������!M#�/IY
���Ѭ�53磇l��� �i-V�č(��ݝ%�n�x�����&Vk�P��@�7!R̀�^��
u��u�*�ǹz}6�(����+o�B|[�����ĮwwtR춃�g�\���B1m���fnDы�;��Kn�����~E6e�3���r���"5�p��%���h�eGH�7��sͭJ���ĝ1�.�F����A/�RGlf݀$b �T�0�y��H�� ͨ��CKf.�Ĺ]�]�,����r� +�i�XI"�~T��ZJ��e�����*�,�yp4:0�q�Ge�6��{C�f\�Gq�:,<.��?��/�q��1�d��?�)JH�&�{��NGg����z� �ce!8ɭ�g�t��,c+=r�A�L���r���,���¿�9%��5{:{������~ͧɉQ�r�v�b�+����ٜ��?��$]� J���n��wS������W���qF�4qܴ��ۚ�������e��{�^�E4��}ʍ���>alN:�p,6�M��<RH�]`C�גE��$7��
���+�T��Ahr5L)��ى|&zL-b�h�5M�ĔV���A�K�8�����������a�Yy�./ �a"�<5�Q,���s�պ1�k�wy���%��M�_^��N��G��1v����Hr�+V���<iS�Z�4c`��ŗ�4�x�eI`ȣ=����0�|&SVedK��de�nZ�ZZ��pVC4zTyv��Gp�sz���Z�%�&��H�*X+r.5�nJ0
��i;<lf*��%����l��)��6����P�ٴ#�2���g��}�.�C��a��$�Bp�)��� ����ys�G���F\0���_==��Q�QO�S���È~�O,7�g����28o,Ӣ� ?r�qt�}���nB2�s�$�>�!2���3�I�@y��ߪ?f9a��l�9�s>r�F����Ybh&�	l����5a��rRVg� V{W��a"8 ������򈜻��{���}����� �M��m�JÕC�^��%u�<3�j`�d\i���y�ҏθ2��)�BdWg��H<�Eh��FS�G��H<a�7���`� ���k��"3�|�<�����ɉ�ƗHS�+~R�A�	��u�1t6{��U� ���"#r5@��"���:Ol�U׉����";}�r<+B0h�ɿP�#e�|����9������J��M���d.�Czȏ������^ò����G�����=@�o]34��d��*5X���~S�bd�O@. L�B4��w�����~���"I'�=5/���#�����P��a�6/�%���(��ez������5�Ma�����dd��Uw�{W�592�Qe������2ed�8'�'c�T��jN	�5-���)�v���H�G	���*��s����	M��t�Ls��1Ŧ��ض�4���r��}@>Xh�I4����K�N�kc2��%h f^�G:�j�V�g��ȷ	{�O�!��;��H�r�����V�R�i\de��"�B�z�[Uy�a�!�j]E����ߜbf�z9͚ �Wuq��0�����S]�y������Qix��
����no���Q��/J�>O^*�tX� �HH":=�N��8���9�X4?r�メ i:Н5[-(�OF-�ly�*���Z��7�T���l��ai�+�?�G�9i2v��0���|��0 }���Sj_�����N�ws2�M�8�����w�H��p4Vtrh�Im�����i~���;Nl�!��%`]�Աz������<�og�{�i9@j�z;�I>b[ ���=� >�C�9W�s-�a��H���1�q����/NhN�y����Ur����AL����BIΪK}�I�m�6��e�$
��kJ_dOn���$�������y*�V���l�R�>�\*�nr~��VI"��6� �J!������+��� d�:�|��M�pRj�ё�|b���]6�u�9L�d�yx��8�A#�1�Yd���X�u/�����F�,�vޙ^���B������v��YBw�dx�,����؈�z�SFX��Ϫ*^��'5�ʣ��,Z�C��z\��	�-tb��%�!�`�X�kq�Ԙ� K��s��5�eio"�Rz�4�N��̿C��myS�c�wW�C���MӾ�5��Nx,��%��r��X�yh:�t��X~g�fn��k��y�۴���G���6;�IV�-��l&��R,a�ƕ�Ӛ�֓N*`�P�͙�S��)�N%QH���s��O�r���)�!2�m���LÔ�7�z��W��C[���Z�Q�����).�sSi��K��ng�B�33nO�D�ꆣ^%2��.�������z��7�Q�H}*����M0w�[�'�sˠ��VMO�N��v�n �I��̀k�{ ��X9�CҽX��r0Ѐ
�h{P�IW�۵tW�+I�Nq�S)I�FW?�1�g,��Vq��xO�[�k_iQ�o�ۋ5�oSgH<<�PiW�WS �i��y9�/�O��@i�4͑�����;h?ʃ���4�_O��	'8Y�_S��O6�����`�\ 8�oN��ma;S����|#.�UC���9pd��܂t�w#y�����4���5�1�2�f�4����VĀ�"�S�Ō��ԫ9���l�>A��9���g��-#Tk�����G0!#�LMt�6��W�������kf�~���7�$_��A��(}��>1�x!(i��M
�,6�鯞��p�(��s~�-������ S��e1f\���
֥l���aA�����᳷~�g�S�h���ZK����"��#
 �gSލ6뾅���9B��Ǎa_o�O�O��Ok��G����������w���h+@�aJ �%�����;���0�d`�B2Q̈|{�:��VJd��6hWҽ�z%xˠI����j�9�5|�S�R�JN��
o Ӧ��ej�AR��?3�؃OO;�@uW�sA;H7\<��^� CN��Y�GMw�'�ܤ ��9M}ZX�b�{���TT�g\y9��͉8pO��d칄A��"�vk��P�V��3x��@A��F�'�YX����Y(���ⷢn/�1��æQ�[���ПR_�b�P_-����Ŭ����o�]����i,��L<`'.�:P���$o�C�А^�=���~U%X����n_�������y1��Q�_8}�`U~��@h+PR�}��s`~��sB!F��m3� �A���� B���ni�X�hs��Wt�m�R�W�A�@������H���ȍkۢ��.#�u���x�@l?�9�3����6�Y��XbTю�iC�@�v���vF�J��6� ˡ"f�Y�\���f�N!P@���tY���2���x�dV��-�GM�Z4�?"�E��Ix@0L��5BE�B��;��c%\P���캨Krd2�i��<ԁ�P�����lg�]7�B��<>�����9�g��$�Yy�+J�L�&��B]Gs� ����/����9@R��h�B#֮�C2)d�BsC�x��}��3m�;����]v�w�Ѵ�T�W��,u�acYP��j�\����3ө<�C傛Z@����iD��rac>J~pר}�o��,��ѻ�89S,ɳ0�Ze��B7~���=���GF؟���3�\M��7!��}�7a60@�b+A}��.��Ҡh�{P(���_B� �ٰ��,��`��N\��Z9�Ϋ/�ߕ}�ջ�Dz�_eC�ݸu4�y�lMJ�X��@���q!�$(�u��C3�6��c	-=�2?���2���� �'8fnsФ��
?���u�?�w#���g�
�t�@���z)/����*:�?�xy��^
���ɯ��6Y7WvI`6�$7�xX�5Yz!|��J�UW�k'�1��������F��)��c��Kπ����1X&��VC��M��^lu���{7c6��SN��o	Ҙ@��-	�����hO��>A�p[��t��_������Ce'�&����j�9�@���for��r�K�EU3oU
<�ELL�|�i���HybǚS|LK�u�0��	��+�y�,�ϖP nP��:)oM�h^T|�ZB�1���U�Ӥ����q���a������۠��O'F
���(�Taы�T[»��?e�I�젣/�U��p r8
������X<�>�^�0�G�����Coh4k�kF��A֒F�����ɈQ�|mߜr��?�{�&:p'V�)v�ZBݼN��5䤈Lp-��%K��$З�ܯ������ �R՞e�X�c�3�o$��7��-�K��-�]�������<����V�'1�(7�ƛm�/ʎ����x���b�m$�̆͆���@�ϒ�l�]�,���5g�`�;>���p �ד�bЊPE�N��^�}��m�Ulv,=�g�84V�GF�Bf���^�͢����~�d�.��>-H垟8�1�����<(r}�����[^c�����	�g��OP���L�ɤ
1�4ORf����#���t W>񻣛)���?��/�1��D�f�5QsZ�vr��Ze�-�B!o�ON=������O�͜��Ӓ� |�w����\�=�}��dFR���fvO���~#�3?岠	>%x~3���DX�4��w&#w�����C���S��|��X��
��K�����d��HH`��]ǳ���+�E$�YY����s"qdV��T��"��iW�J��$܄38@J���l����Pq�3+��o� k*�s�-�u,��H��u�\p��%�F��I�^��c�C_�ڕ.?����1�E���>�?L&@�2�!�}�	��4o�M�������Kxl��Ϯ����eP�b;@w���li%@�l"��f����q�I���}P�O��n�i�t�,�.3\�
���~Y�LF�KִZ>l�enA�5��z��ڛ�$=��{v�=G�8(�c;��ݘ���Ί���}�� ��
w�x{�q]s��>�m9$���n�S����C����H�~L�=�o�`��p����q;f�<B�j�3�㜽��{�k�)F����b���,�#�w���*���<N$��g�}��f��먺���M��Rf�Iò֣�r
!������2.���8�9�ŷ{�@�iA�@"=}i��M3�hQ�;�gE(pIǣ�>�V8rA�S]��HGf'�.Iʽg����~�����-�$Fa�h�$�:H>>�U�	�jK~��p�Gm	[�3�0���D�����"�bue��I1{�9~��؋��ɜ�	͟P�:y���Ĝ�fF��;��6|XzH�o��>�z7��g�~�C��Q�"s���J$&�>W��3N.���OA����
���%&�IR���=�=��&�O�ނMnP,3���W�{�9�.tP�����R�0+W�=y�F:v]�d�����\�'�6����6kk�`ϣC�w.ӆ"�m�-�1�� oֵX����$�q&7�����ޙ*�Lor��cj-V bph:�F�T�a��8�O�	ԋýo��0.P�>� '�[�*^�*�ލe��jb�ٶ�y��0�\V��HsC��: `-6���B��!_Bˏ@���񏻱𚍇�%������E��#ǃ_N�#��Xk���I��i`���j�lI)���\T8c�^���܈6��+�ق$"O�/��vSVgZΪ�@38dCN�����T5��N�k���K�9�6e��m��z=ǚ���I}+v(�-E<�����
�j?8L��:�pn��[7M?�1b#Zr�����g|��ړl��>���#�b�%m��1q��2�%�CB}����ȵ�)q��GN<����Yk�obZ����vk���<�w�X��.JJ�����/��W��,%S�&{72�EI(C�bp�'�\�0M,ݗ�`
��F
����|���(���_�)���uG�
]�����k�C����w*�y�Lc��k+�r���9�>da���17�e�6FMv����D\'����[��V��Ն��e�+���.�Tv��-g��,��er�jD4ŵ㉦,X)�{�-=�%>�����PlUf�*< �f�r��]�H��(�W��+�1�+๬Ҋ,֓��т�sWe��SK�<�x~̍ו�Ĥ�9�1$`�:2��Σ���#`+�R��5;��K-������{�	oɅO��?����RC�w�7?ͧR(k�;��0Hz�_<��;�ɪ�6=ҟ��m�@������_��>3��OZu�Y%��Xo2\f�ܧ���[|BW�Ɗ���u�&;<�P�}�,���%��ru��C�!��T�.P��+���2鄣��&`)t̂�7�4�oϘַ�m �����\fʕ3�]���3�Aǈ��ɖ�_��B-{�f9�Ҳ�㨴��#�wa�(�=�t��)V������m`��c�|C�@��Jҥt6��,���ޑ��5O�C(�Cnh�&�,�[s�7߲b��URZTWa����%hN�Y��<���-�ٵ?O��j��Q��F�='�������M�k~uuЮ�~u:=���ن�������t��W*�=�A�zM ��/�w���I"�l��e�ѧ�0�ҥ6����<y��9�sk��KJ_nIV�?#h�d:�%ڮ�[o������<>����!�r���P�=7�]mv�v(R/\�0`\��Թ�g�P�D��1Kg�'
j�L6u�
QD���?���m�B->W���e���ۯ�Ł��\b�RR縅�#�=ֶ��g�?+k�l,������ K��y]ぢ@�ӭ��.� �%2J�F���O�[_R�KSe*�C��q��S��?�� ���E�c70�_��= ����4���M[���Q�_o��v���B�3z�Ñ�IE%�����b6�U+m�d�U�~P1����ۚ�0����~��U������b" 6@���u��9>5p9c��ރ���ɷ�s&�<�1�k�;��Bu5�j��nXr�&�-���G��;�e�8��b��~&�%�$D̲%gXp�F�E���-3�+T�V��.�s�)fY�@��{��7��V��-lA��(�A�t�
j?��SD���;w7ڙ�Y5����h9�]L�4���R(PD�s%c*s��ja��� ���=/5���bz��9$��iR��9E�>G�O���'	��;p�^��ІI5��59��B�'g�V7�	G4_��^�J~� �	$��BkTe�82�P@;� &������h�>}(
�
{���f1�#q��b�k�ʽ^iQ���w��=��d4����/�U�~}�#��I+�����?�֨�T>��AE>�ק�A�Ƅ�V�l�Ғ��i�=� e���~HtT����(3
�R_w�F�o4���8����E!�z)F�4�e΂�_�����TV��ǫض`��:��M(�R��� ��.'%W��|#-*�"='!�k�Ӂ$f��fl���;���B=���j�8(����}}���ά2���p&�Z��}L�����}���4w�5�^fH�T��8#&�UR�11��/��|��~oB1����iT&	��X!�zO��Q.P~�xh��X�O���
m�a|�	�e�����7(JRJȆ�"-�E���u�h> ��"�u���X�`Q6�4?�0���ǂ%�Ĩ��v���O�9�4������T���RF�<������o�l,��P�:^�Kp������Q��
��i�#�����9Y�i�s��)oǜBI������]��q�/�.���Lm�G�2'v6���{�"�&���D����bTW%���T���5��Ȑ>�1))p��j��������y�f��"�Qi�����[5N^�J�MK�aU�CJUX_�LNB_+G��ﭡ���ϰ���ޞ	`����i�=m���
6��T��
�"�g����Y�5������^� 6M�-B�hch�>?9��#��(a䗔�wOn2̆J9���Δ=��nτ4�^��Q׭�Շw@۴5�Ύ_s�1Dd�9�n_��Ap
�]�s5�C'M�=&���i�L:�u$A�_!7�=v���QtJ﬌삱�2D/!�=V�l�'[�r
3%��g�w1�c������&]��rtK�q���9T�	P�{�R�S�=qg���þsD���f�*N�}�oy��:�-2�E�Ws!�?����V}o��'m��z�"Q�|�(B��ޯ�ܧ�����
#k�:�@�\��+g_�౦	Z޼�𠊴��$��"2�N��P{>W���v��h�T8p�N���8�H��'Z`�^�%�C(���3����������ۭErҋ���qO{y���A��e�޳^A�f����Š�V����V�R� ��Ε��&�e��y<y�]0�M�Q�0N�Ef�u�O��޻|�X0������@���bS��\��0�@ow�ԈOk@�=�4,���=r6x��{�F�oB++س���-�j��Q"&�<k�e�b��p�Z{��X���a�+��}�߶��Y��)c)O,:Cx�ִ�J\F%���I���a��)=@������,�n~���GD�&��	3T�>!f�'�������Z�M�94V��` �8�/��gʼ�h�B�R�������1A�yJ��<�eL���=�v+�]��3���M�߯b� ��Y^{��l���S� ��-y��.�ǜ�4��g�tk��q@��z���>+Q�)�˛Ӭ���ǃ��hC���$m��@�?s�\u��|���]��k �7#,�z��I�	��l��߯?�_�4��@`w��Y$m[����S���avDf�ى���*��q띃�iި�T5ƀz�+i`�d�C��Sn�o��P;qJ	����i���z� �L�Z�_A4�Y����'��E��m�P��9*�w�\;R~����:\��T���yJ�'_Ğ��ļrl9[����*�!?����=�R;6�Ä&��`:�A��~p�X�J����Y'�]+��Q�9�_a�
��?��^>�]��=�r���<�a��ϫ�	���U����&]��i|���� rK��m��=1ߑQG6@�]�)��1��u���ڀ�V���,Z@�#��[!��KI[UX�����W���գk���Ȕ�(|1�}�5���V��rm	T���4xIDz�@�4/wZH���� ���	���MOP50�<l��%&y֊eH��a�w��#��^+��`,�%7;F�gi��+`YM�m۝h�͂iAd�f�wЍ8�՗��>gC/�\3j�n�{`����ާ� 	M��{����X(�o�}u`+!|mO�L[%)��cŰiV�G�zSh��u�& ���M2�_���i!qtrr���x�
��&m�Wj��� Xʴ�M�jf!��2���색_�C]mP���q�dS	}w�sC�$hR��S�]�>����/V�ot���H���Tc3�[�n�"�m@��X�F����e�HD0Ipp��"��`�W����#�#���ܰ����t�Ȗ�;���� ���#�����;|oU�uYC�NmX��Wʭ���q_Ħln��}��Y줪>�C�p�N���*,��d���m(%��虁�
Y�*�@��W��I���:0<���\�0%Jfn��w��Z[�=���bNs��Ų��������]ŻPgຟ>�����ˠB	�m!�����}4a�ICس����n��K`�V�196�"�f�k��f��b�?��b_R�ƨ�e�H�h;�8�.�X�ʹq�pYS��_�I��HZ�11B�r|�, 0��їA�I��Fr�|�o�L��1�2�Ý���{N�
�G��J(�[7�r!.[EqJ~_��~i(o��K�>9���i�7����sb�y�����g�
��T�v���Ie�("6���,e�O;�cvc5���uQ%YG!�Tu�S�����Խô�#~��2��3�*�i��_�ڵ�Z��=����p4�F���*2C+�1�fMN)�/�Gv�U���8�/������~�ʵSx�)ɬB�Ԝ����Ԡr��K�B�#u����qd|�e��L<j��}>�oL�����D��+����k�ɲ�=�]d���S\�(��^�#UEb��a��gu��,7��g��_��q,�0�(�X��L�i�Oq�����|y��l ƥ����pe�A��i�=H�f2Юa�8�ȮK�+˾��)���D [�$���YR��" Z��p��H�m�zl�1��j�)gE3Y��|G��"6	��P�.fWQ>�(���&���lQ;L��\�hh���x�����j��'��1Y.~ղ%��Dg�?�$p�p^ � �֬"{��ˣ^@@Z���#�w����Fr��a�.�����
s�9����m�o2��C��໕�f��g�
��&^h��=N��?p�<*�r+s�6`a�8���Sam��iB����xL��R%I)�?��]%�����F�K����=��R����ɯk��I�U�$ F�k���e٣�\o�:�Gh4�	�h�� ���������<s��[k��W�~K�IF=`Ȏ���j�z�R�P�q	ǆ2��"`�1�#�1�sE0WI�@�GY=�]C��6B�EU����mQ�3ħ6�7B=(�>A��rv���fY1�9Nʴ��>@9F����_�H٫� 4ԥ�������\��%5�A��%�U��ە����5E�r��Pwyɖ��no��3u9h!����u�>�sn�.��<ѓ%�l��E���QM�	����8JG4h�`� r=�bh,��A�B�wwd�E3�/��ݨ�U��r=�T�`��8a�X�ȇ�O�)�X=���Gc����.�f��?�V�S��w�w�~�&y��9����B@�#F�?S������R°#��'��P9'�SZ��_ �71���X�J��tݝ� [8��ɇ�d���-4xM
)Zi8Ő�q,l�E����Nc�PS��.�nu�U�@�6��Z>l���,&������B�->�/8���������w��>�B��؏9���B%��t
c���hu�n�ZɞP��"m��dѽ�C�B���68���eE�D�dL:��q����d�y��w�w�U�%��]�b����p8?��s��ajC!�Ͻ���������T�=u���l���3�>:�L�tu�j+h�|�`����i���͈�M� �J��1}���\��'|�0�h���(��<���?PJ@���U�f݈<�bIJ^�!X�-9��c+8�PF�k�:py��5�/� É&�؂,{��/:���3x�=���mm�Y��eH�7���%�vђM��\�Ÿ��S2��Uy�#�^�"<��?���a�*�9��5��'I������F|���4vTA-��No=���S]B��P�3��<W�䫋��9@ֹB�,Ol�FHo��m)��،w1o�fY�ۗSs�$�U��̙j¾|gx����Ҕ�œv�)L��-H1)���n3_��`R�A�(��h<]{���2B{�{M'X}��%��E�d��9.
LY���R�cV�N_l�3��tf ߴ�ǯ�l�׎Lu� �	O����yf�;��> �QiD��ڶ��2�>Sm&����\��I�}Z_B�ϬU�]���!YP�f ��8rϠ`#��.����� ���__N�r�r3LM���'A�Ѧ�G X�;�=���$<��P)/��o.�+�	�#\a�Fw�����F����"!u���%��;�f�jji��P�/���c_�)�'}�o-��,S4��̻E.�k��Jl��dmW��N�*�|���$�@l��~P%�g ȹ����U�<�g�ԃ�3��~��V�qM! �������,Nz�V�T4�XA���ڔ�J���������w����S��d!��j�rb�d��B$�ڤT�n�p5�kLV�Gd���p_����;��/�9�2�2R���SSJ�~��4&��˥9��v���\z�������uĈ
���|؊p;�����E�ۈ}c���5�՞�/X�'��ۆ>8F�j�Xϝ#�����_��z�D�����0n�,��tRe�%��Q����Ze�z�k|N��R1]܁�C�]�-�VuP�p�ɢ��i�>il?m��I�7�3�ӕ��=tΧu�� �����.k���m�Q��ZEd�2��m�=��NcG�s������Y
�t���C��F/� ��r�'�:#���i��c��I������!5.-Ht.��'A��b%1D6�,p��K�ON6��)�� ��	�|�b��k e
�A}��&��bc1J�
��.�!��N�~��>1�=U�����P�w㾅׉�2Ԝ�P�N_Ԓ�����6?�����p�� ��[悰r#�w�ƞ�1�2���]u2���ꤥT�{�"��l��J\���&J�y^b��2��H:;R��&�@�<t�A��wi�Cۇ8���6�o<�LY������_�� �:��oh+�y�!��`V�hq��@�6?3������q�dId�ƃ��8݊f������40��K�U
a���d����"�m	 Kx��%.����oND�@���yWQ��Mz���MƼ��{ҝ4��y�+��.�\��`��-w��������h�$M�Kt�<+wnL�~�5�)����g!�YwCX*(2*���"���������4C���ø ���5����@�"EG�R�4�x8�x������W-+z"���3ܤ�TF���xS��;q��s.K�X��t,�=r�2}M��w�]u`bR�s���k5��"��r��&�voDf�;9����D�^�U���°�����/�)E,��%��=�L��
�-U�~⁎��@��l� ��j��2q��S?�ܲ��~K�����a#�\�Sm� �ȟ�3�~�8N^�0��;B$j����o���̶��T���=��[R�.Fs�J��X9C����pbuG�_��,6��k�x�a�%X%�Tw�9~1��x �e����̝t�;Y ���),g���]��ى��#v�p�|���<b�T�K;��c��u���0�D�E��`�L��?��Xj�cK2��5a��Wn|]�	����o�W�h��'wp�l��4�ϹT!��G�����~U7Yx�jN����;1�����*t��B�ʎԫ�'�Μ�z�B�m"dTD�y��\�	uц�������9���[�����`\(��X<W9vS` ����wdXch;�5!�
�GR&��"s�'��o��WY@kM
:���0����yoe� p:o�m���!�Ij�a��0��G{m������|����T]9R�������o��s+���;��N�=:��P:��?�~}&�3^��0�'1�������k6YM�u�Z�u	�f+�e-� l�$	�HRF�^�J���o	&��O���SɁeI����Ny���֬�����7s�^7/vF�lD����"y�s#�ҕ�U�Ӳ��M�g���:�O1n�6�/N��D�����ȓ}xxM�P�[��G��43v4T�&����a=�P�L�ৄ��q�k�*xw�§6�?����6�"Z6�tR�R����`[�d�
���E�M������l=�������!GF3Avw�'8	�~�pI�f�?k�$�x����'�['K�?�w�����"��9	�mΖ��3ڇ���I]��b8
���EYK0��$R�
'��j�c��k9���|�&��Y�	��	f�U�4pR�}����3^t�w�0k�B��_�aBW8u�X�������[k�^�q��������v#���ɪ�ף�D(��'��ц��|�;-m!>EE3�^�9���Jp�T�`�����5ysXZ�PD=��S�jQHL֝��곔%H���ߛ)��K�1}ept�H޽³���>�B��S������� z��������A�n!�J �h4�i��'���=�ֱ�H0�)�5}��]0���i��u%��4�hG�hŽDP�9���]x���EAF�5�r�}X�\l$��^uy0�2菂w��Y��D+���ԫ7ih��U�Â=�k]-�u���<8����e#E��-	����65=��)Y��f��Gz�e�'廛9h5=��v\QfhYbmFZ{'�]�e�#���'տ�f���s��:�iq����nA��6JMN ��%�.��C��T�\ �a�b�Y�\���m�k��P���R�ȫ���i2A�Y֛�SÂ�V]��eD�7q[3��DLEmZF��*����V���ԍPM1��g���$�#�͑��4��Z��Vv'�#�������Ű�s���]�8�ө���2Vq5�üB-�yrDw\gcMg�du�%��Ze�����ͣB��4�qm)��֒����$n�����6~��Xb�v;����s���c�Hx6��6FO+,��hLt0[���a�k ߢ��_�#���O��`)T"�/��g��aI�Yӟ�J9�@�\M�2�5 PXj����j9���j�)��hܧlO��@0&nU|���(Q>��DI��g3]���Y.�+р!��T��l��\���f���K�ȧa�EF�cѵ�"D�x��X�a,��׏�wi�״a��(
S#�5����"1r~j�[^Q��(��@�� �5*uB�qM�R�rB�LX�s J^�ġ`�lr�E��G>{d��� �C��T/�D>N3���8rėh^t�خ�PZݐ���Gߝݱw$rq���U���4����C-��k�@Ҏ:�I��(�j|�L��a�%��\<'�>���l~��N�����%�8��>8�*�K#�տ��v�!��?f��
{hn�I�!��H�B���H	��tOs,�w���Qݨv�w�i/��)���I�=�y�W�?#�QfA\%v���������R#1gM2�-�^^�zB�7�$�*�Wj�ڠ�m�k���P�]���Z~# F�+��%�L=��џ�q:�~��g�=5�H���G��3�1�`���P�y��
��^|E���u᛫_�Wx����A�Y��]K$ ����5�3���|��A�2���'����+�1��H��K�Q3�/����_��=aX�F�d�j�1����c*b宗� ����B�x�S����(����g����:T5�}�k���X�Pȩ��a��m��n������k[�P�y��g�=:%�����0^W�K3[::�k��vs�g��(��6��SJ	s�s?�E"n����O�C��u}�s�9f{��]��k�`��er�B���u���D����῟���1x��=�+��}�q�����o�Y�s-Spt��zO���[����Q�����J4�lٛ\����G��Upl��[�%nH漏��Ff��y+9�%fX��,���D���"�v���;�9�	��T�ަr�<��>�{��7R�/��Oކ�,�$�VV��?ӄ���gZ�	����R�b�Վ��P�.��%D�鸔�����2����~Ky_�p�"�_*�{��n^؝D�<i͠�w3����
���M�*��j�5���L�#Ŕ�{��q���*�~�.T��V}&��<r$�U�/��l�����t��� Y��A �:8^��3)�J�4ؘ�����	�(U�m�R��W��-[0(z_و��|�Gff�����}(���&�R�z�� >w�O3m�G����/�����w):3��	/��wL�$�3�3y>��\����p�"�;���c�7���<Q����z3�(ZVcCE��μ�����I��=��.#(
"���[t�{���xwU�E����.ᡀcȽ���J�X?2¿���eg������=����*F6��6�Tqܫ]a>��=Y������;z��ÜJ�8`������a��\��ߝP�
4�uf�7T�o�ףo=�sA�$��C��C8�с��H
G�
b��mẚ���	1@�Ac*a�qB�k�C�����LQn9N6��x�]��������aV�F� (���Zsi��}��չ}��a����YW�VC�0����1��B!�R{�k�7�U��g:.g��LfW0ё�P��pl�I����N�����N�|i8G�{%
'����>�n�/���E�B�ck���0�Y��9Y�.7G������ڑdp���w�� �#�����*X�C1{�f���H��@S�v=�3��!S��P�V���=Ύ ��������!VQ|~���!�t���f(>�D�����Z�y<6F�´k���#׳äۀ�a��ğ����b�-q]� ,?�_F�<�L�������kJg��I���d�c���+���QgE��f��P4P;������]��
K�%{�8N<s�S����w/�E���ט r������AY�{��������g$�N	[�����������N�@���jJ��O��g ����!����P�dJ�?�D�O}��s,��Bb������~�cGvz�~��C�<"�i�$=L�����Z'�?��Z��F�"}�ދ�г���:��i�t� �Oh��-B�3���&"��=�f�"�� l���ZvL^�*� 3�젣��G7�A��F�L_��6Ɵ�_q�T4��_���J��@f\R;�b�|Y���6S$��0D&[x[����eD���;�6R�\����YJ�2I	��K�T�h��<��إ5��35�}I��1�ҍ���M�T2DOMq�.̥>�Sꖰ�~�MAL��_ˣ�`��,�tC�4Be�BF�X:�Ir�c�0���w�ҵ)-���c6u4V*�NlF1k��b�]�����S�	E���?�H����m�?��5�)]���xx^<����#&�����@\�{��.�F���6�����F��$�q
o��K��{��i�s~Q|�֢$?u �㘻�'ٖ�@�=#��W��aJ��?�U����	� ;�s���U�C�V�����R�F��)7q����ٛt%�Z�y�[�R��8f�hv$����㎟��A��iFP���+�d^�$��0�ϻ��Aag����W�s�m�;i�2н���XY�d!1ߖ�����+*ؚ4�)�/w���`U��%uu�}��u4�X2K�[�b�tMO�O�Ő��4��,)�-�U>�L�HM����ʨM���~�~%e��+H��jw�H��c� �����!a˴�]���3���ی�i.����C��TS��>��o�I���`��	P��p�ȉ�)i;�`Ǵ� �~�o*�%�K~^�<͵\�{/�Mq?)��/U����Y!1ᡚ.��@�WĘ@��K�	���	�m��.QQ��xK_l�˳%c�w�Q��c��7�~)�4L�����i\��RX���vM���6)�u����f��ۻ�}�Ҫ���0�I�C��t�#P@.��U	`yp�W�ۊ>����,� i���Ѐ9�>Y�#���d:{�Fw�@+��z�^V����B���9�dC�k��4��X\�L�Qxp!�ҴZ�@��K?pHL��B�w��U�$[��}�TضB`aV1NS�;u/�qS{��E�wTi}6��U	�!�3.	�*�a`��g_U3ysl4Si���H�O��^4%���V�$���q	�X3�b-��;��ՠ>)i��U��	4�]1�+�'�Ȝ�-�y�R��	yt.p�R����hc���3C{���p�2�����QNkX���;�1�]��SƃLA�}�9��5���A��{���{P�F�N����ДiiR��e�.�d?���)���r�d��ĝʵ?�O��Eͧg��or�P�f&U��QD����(x+�k#���(h(��t͌�UO��}jӨ�Z&w��,�v���v*�v�"ͤS���i3��V��p4�c�?�����bB�x�����9L�ډ2�N�4}}*������d�j�D#��6s��8]��mϹxAܶ6K���'z�|��� PwA!}0�:�3���'�M�A�i���_1�����,�y�"v����m�%�wmnk����:�\�+B�3Fp�JU�~��C׌�H��\�H�y]��Z���-O���й�PH�go��� m?�~i^8��<�J!�l.��4��Q�Iu�,W�1o��;<����hO]q.?<�;"�P]Ǽ�ĉT'9�D�vG�5�$���n���W�zn!kra��oan�y��*՝�PȊ+T�������\$S~�-��.$��	L��9R�B'��o�#��y~^����Q/�{�#{i=!3��c�z��H�䗊�!*�Yjl��'H
�ן�٪�	�o���D���3��?Rm^õ��v��_�E�� ���Vќ�>��U�� �6�f�u�Qk�C��48�!��&Uq�yоy�\T���Q֠P�Np;V_a�u膍ܠP!�`��E�����'�Flb��T����Z$[��������ES6͖��=�L���@�؛��
C�����7�R�OP'�b,�A7��7��XPഁ9��26nM	Ќ����P��8��v+q�-�ـ�#�7b�2�0�}Ғf���,_7�t��������_H��5�[������8֛7	i���0O}	�*D�1-\F�k��)i�>���ٟ�&����%ҹڪ��E�V���#/W�'�6��|"�h�։Lځa���@��O��dE:X*7u_�z�p�g ��,ku>������9��3���D�Y�D��T��&���Ru�kq�v��`t�b"�J|=x.i�*���9e+���
#[�s�z��7朞�C��
�(ZN�'��l���U6N\Ty���X��r�O	7�)�=�PkL���3m�sk�O�N�?���H#���+�;��𾪜^�"J��@��XY�vWCVn�n��[%��q$��#�c�>K�G��D�(���3��Ϣ�<Y3���e�g2>:�'%:��=��eq�u���p��
<aPf���P]@���4{�2G��(����Z5��"2� �X�o(����Wf<p�x����	Sr�����u���I��x>�ȁF�\�ď�!f`��N�k�՞/<��
YX��o�#_�Mj�ū�[��\����&fg[7��#�?��F�w�Ě�C�?ZV�~�M��4�q�NC
�vち�	�:I��PA��%4�3���u�x]�h��!��cV����ey��;/��+T�#��n�>�Z����L����MN	BY{xl(�6|X�O=$�BAc�<}#�Y�`�p�-�z�ҋ�ݨ#9� �Q����(�Q#�q��O͢�fW���8Y������T_dw�Y{�o(��۟F�u�/d)@o��Z9�>��vDC�T�&����R}���O���I5x���VGo7#%0�>Um}Q������+�g.QU	Z�M�i��G����]FT�&WlU�� ��Q�m�E�ԞM����<6ޘ���F�;Z��ں�3�?�<l5fmqUU��n�ܺ��y����v,N��7��Tc%�����G?�Dt�@��A)�;7r��Y"X 8�K��Jǟc`��
x[$%�	c�W0�糪	�S߄�K��߮����`�'�5W��w�k�1TY)�k"�a?J��#A
b,/j����$2��4A�[���TiX7�Ҋܼ!����3�vg�]#限IN�fx���m2�fnoք�;)�߰uՂm�&d�ߴ�<��s�^�^��wi�ɥ���.�k�M&�K��BI��B-qE�%���	�Ŗ{�i+`��V.y<$eF��~ڌ�PX��=3��!m�)�[^(_��^�l���� ��O�+��� 6û|����C�0#fߕUN�=ʟ����u��+��Y��PFF_ȚtRg�yZ����+8zo��igV�) }*�\��{ �Ã��Qǋxm�u9OK�͐%u@7�p7_4��XY���WWԪ���.ٟ�0��-�G'��\Du��������/4d�l��3���>��mK��u\�a��nx �6Ι2����$�p3/��Ѥm��ދ�j�J��|���*9�Z����NW�6%q�%5�Rӿ��	'�����/���~�x̧���fK�w�c/�c֏\l{"��2}lA4�iH�V��d�sd������B�&Ń�7ˍ�*���M��G�� P2ܦ'ğ�c��4s�<6U����j�~G�+������c�u��{��k[d='���H.|��fܢe����بr��9T�<e�f�؀z�Ƌ'�]9:�,�E���^+��h\i��u'[���g�UC~MO3A���: S}�TǢ���n+���V���u�GG�j�L�������8�.t3Ht�0	<&?HP�}���0�[��#栒�����W�>�9M���W��G��H7�to��rw�a	4�8��!:�`w�"pi��.W��`b*�?�߸����kf������A�ss�*��'<�z3�h��/����`Vi�
�I;���0����,�d�����K���	����e��ŏ
�Vσx;��H�f9�&���B�"q�,��ZX�FY~4�8,�>��=���SQY�PI��A�J����g��-=�u:`/lD���y^,o�bjGtw(0�aJ	�i�;��Qa��;3��rB�mH�޼��&rl��JF��*��C�Tv5Bץ �Q��1^�M7Ʀ��:��5{e>;*F�f�n�:�3�a�Q�z3�lA=��ř��q����!4D�)�a	��� �<����̿�';:!�Wʑ��te?�)�����S��5F[�<�~�:�T�~�����dA=O�x`>��Ӝ��f�M��Y���3F�Ӆ��9��.������m\�R~���4t�EMb'p�ly���{��=Ґt����V�[�Y�P	��(�������	-���T�#�
��,!�ש����h?��lH��捒��{"&�H1�=ev��]xMp��:Aꩽ�Z�zF2�����U�,Mm�)ޢb�K�w{�7-O�:����`��j�)�qQ��B����	�������H'���{��b�"���wY��C�=_jiJ�:����4ntS6��!�V`cL�"`�FR�QQ���j {3�!���N���_۸���?e��E������z"k5�E1,�/���d���ۢ�}$t�Bwr�Ǒ�/�)��!�ɴ���A����I���X'�{Z�x��O%�邚ytq�X>�K�Fs���毸N�l�|�q�rx�����$�vZ�;���;�ez�p\�a���.��Y�1�d��S-&b����E�,�A
�-�1/����b�,��1t��
:~*� .9�B	���I.���WlWb��
���ym��p٩���7�����-o6u(�y<��'(�/嗷F7��7cX�m���h�Db>��AB��� �Tͺ��&�M����2�p�<��p}}�>��:'����1�L�Ks�e&�)3����3A`�o'��b������.��7�Y�(�k6ɔ��`����[�g�D���F[@v�u��t: T`9;�M���5�$�A��G�����:*���^ŭk/��r�jX��dh��dҗWUK���@%((�Ϛ��sI�>�iK"��e�@<Aާ���h��s�X'5�'ܲ�q�"�<�ǘ}��s�
u5�CY�W]��
���x��q�8�`���*���n�qM�}7e�u
8�d�ֈz�JR���MF�	�Ks�e��W]Μdc����Q8�XO��&�{S�=7����;����R�[R:h���wDܤw���r�o≃�m+�;��V7����֖�a��om4���y]��V��R�)߲o�^�U����}3y1G�������'.	\+3�l�ժ����_=a���4�g֮!d��~p���^vpF_�Gwe�m2��Z�&�f���2<Qۦ-7#���3겢��@�W�S�� ���>"Ì��~�uX�DQu���vլo4^��F��u<� ��y��� i�|A'g6�1�$�cp�
��e!����-�M��D�l��d���
q�݉�%�a�@	��;����u_`\�K}�|�K�Vt�ޤ�,iz||� @���-�'#��eڏ�ʇ��y�0HAI���&.��Oe�E�e�h=���ɣ_p��*�\�<c���8��S	�ZW���&q�r}�j���k��Z��Z�C�#{�_��Ԍ��*J}b6�l#ƸѐQV:�����nͳ���L�?1��,����*>�vҋ_�39�
�.F�������&*Ӟ��״笣��o�$��I4�,�����v7�8��sXXI�4�;u+�	�*Bȸ	x�n�Kv@�k&�3�3�8��~�:��3y0\m^�|�P�ݜ$�q��ΚS�T}׸�ڬ�x����o��>�M�YI��Z�Y!}�^cv�"<��z�f��~Ȕ��(%�]A�4L�X�Vq�����d��/�{g����&��=L��U����RT�T��,�O��H�Ԕ���*��o(�{6{W��i��M�0o�7*o��@P[�LDDj]|U�S�9K�*W�Eg�S��g����\dS�2�\ԧ�m'����1�p��zYyʻ70"���������K]�.��g��>�+	s�`�=�w��*��v��O&����Y��:�8�JMH$����Sx?/y��G&~+ؓa) ,�{����e�hK�o���\'q�@���yYp�C���q��� �7� ���v���y+�I_���e�OFw�%�����F��,��>JJ��/���@�_���[*�i/}?�����L�#A1&�D��/���q��[#`��s|&	�f���|�|V��8{��R�[g�Zq�){�V��8�ؓLx�L��!��eO#�� d�,Z�Tڴ�F�\G��-�ϟ�;b	8^�6�b�����!�.�x�Q'k1��o��W�;�2v(�daq��xد�۩�?G�N �B�R7s��ˠ���<���?���X0�ў9\_[�1V���V�K������m���z�7�5�	4c���Lp �I��:���\ o�3 n���
J�:m]Q�����X5�R�9 ��~.i��&k�>��7>c��81����0k�/M6�[j�Z?��]�^�U-ͷ�-��˸jc���x'BW�oB�H6����T@������<�hMA|c���,V�$ĳ��Wq�K��U
�{���'�q?�zmQ���,�M(��/�r~!� Ȧ��M��gH�S���@k�Qo&,�v�îA���e�k�!ۆ'2���3����ɾ�7q�Nʡ nW$�" }�Q�{�ܟ:�����ؿr��ۈ��sj;��je����v6���?wzٴ�vϣ�0̠�V⣀|.ۀ?=Yw^^����~�'g��:�(�W;��`Hͥe.�Zw��jo��H�-�[}�%J0!e}0/����z{��AE Ȓ�#�7�7n��0���� �C�t��o`���2�NJd��
J
�8�����q�}�z����C�����?Slx<��+vy֐��ʋKKT@���*��)�$n�n�q���>���+b����6aW<���g�ʐ}A�d�(�(��3p,�w_�O|7TF����l��I�E
��g�+,�a���9��(�{̈Tؙ���hs�AB���3� K��_6�zC9z�>f���� ����~�Mbrv��T�O�.e���8�w�]7�I�����8w�Gć!�OEY��C�i@�#�9�qz!�� a?�9!ٔ\�4��n-�WÂ��7�90ľ����w������fm 0�o7��s|s��'�C�̊��^���1n16�n��SR�x�#+cd6t`r����M�ۂxv��y!-����?d���/����iP��S@\-��A{Gs�x�	��%�Y�����B�i�6G��ʷ�	��)��>wz���>B�3��6'�����v )���M�V������x����y���yоe���:�v��+�k�f�l�l�f��Z*gUL;sVBꢄu#~���1j
�ӣ���"���N믒W�):C9��������1z��Ȗ���
J�K;�T���}���b��Ri�%��bm����`YkyA�\X��~Nv��n�����ؙ�N�w�75�|ܞ@B�;�����Z؎/��Ӌ�5D'�)Vz�1��1p5��P,/�gc����pnߎSFJ*�H&�b�ƣ��hlQ�q�5�hB0?�b���L@FY�'5,H���c�^t~뮕t������;���y�G�B��{�L��0?����D����BQ��Æjzy%��;��V�"m���T�2u�bS�;�AS½�P<��˓�H�ca�p�g(/.�	Rw���|<��t7�}�Ƴ	6��Ov�����4`����kس+��N� l#�Ubɢms�o貑c��y��j��U��`�x�L�5��g���E|�WP[�T���uF���KR�6e#]�\&����4�%T�0�Y�I7A���@!4,{0�+�~���	�������M��բ'���XE�|3&@�C�7�xĦ���v�׬�y����/)�����u�2H�.�)��Vr1Y��?�4���~ S�<šN�D����
��7Cxr7�7|��"M4L�s�!��m����4�&��S&�_�֍-Y=���2�[�P����7��w�^��@��Gr_0#��'�bu-�t�a��o���g⦆����hz�@�w荎`���/3EF��R�K�	����i��H������u�������q�e�h�"�Ë'�(`��n�C-\����{í`���㒝|5^�e��؞�vy�9��(ˀQ=ެ!R���a���Cu���P�h_�oiMWa��M��L�����x����G���X� ��?�/b�Hxۃ�|r/{[��0	��,��	��9�tC���󎫊6!���"�D^e0.��MdCڶX��F��*��Q��+\�+�>wn:�>{���m#c�v-��'��MW��Cvw����	�����B��W�yA&f?�MyF|����+��b���HWpI����#��C��&�5}e7!
A ��B$�:�A�(�������	�{[1w_}��2t��A�oM��hB������U7�/�p��o"R�n��[}@j�Li���,�
ꝓ"ʁe�M�
�zz?���J�@�@�*�N�ް*��C ���O�z���ױ���U�Φ��Ac���i�z(ٍ�q���N[Z��Nz��yc���H�$S��pӤz�r���.q�9^h��ߎ���}s���0��o���0WEeu�j�"���D����n��+d�r���*;�#�g�[zжX��C�"Db[@����un�S'f~q�_�a7Zw@?<�G�^vfP�\���o�T	&R��r%�qٲ�+F�M�üVK��:]�%O�j`L@��*��C�k`�z�M��h��b��ل�ƙ���j�G?�R+��l�M��t�����?�k����+��X���S��'�m�	�|�m�7�Y�����q��dyLD�RBL�%��^Dѓ1�F�E�D8���'��
���`�sr�'�F23��Av(d[�1�ͼ�T�?�CJw�'���~�f�tB�I�(��t�+��Mq������u�n#���	�Wc��˳x��y�1�~�L�W��X�
.��:���_3�'�Yj�\�J*wĚ����D����*P�Q6$�"������4��|/^Ҍ+��Οg�!{�	��ded�R~?Gv�/��jG���[-��,ݸ��o5����֢Ć��_I��;��ySsf\e�?�Z�N�ح� �'4&G�b���zf,i��/�s1��Ɲ�'�.�z9m��O����+��9� �2*�Y~��Д2�����2��@x���@�c�~H.�6��[�[�d0��3�ɐ��A�k�������!l?�3dw�{����U�<l�Aw�T�k'��)n�����
3�+#�����cP�j���#E��ri)��Iԃ��FW怢�Cc�˔�&� K�i~�
�bm� �L�z�Dl�R�b�-Y �Jp\s0̽�<�A�h�����r�3�����82�`�:�Z�Y�O��y�����|4X��[�of����BO�q��!Gk-;(LƚQ�߯��"�����d�!���%h�m-���B�g���<)c�F6��}�1��)Ds�q���� ���k�y�'��.N�D1�$M�"ku��l��ܒ��Z�m��Z�hx�A��d��(��o6r���s���� ���#�
�P=F��(�6��x�����'k�7C2l�&����l`´V>q��N@&<�����$B��B�T�;�%���Or�}fO�d�T��I(�:V��(��[��s�&<]�b���{�J���?i>v���jOI4��'�
���!�E/-x�(A���ک`�+��ib{h���D&��by��¼ݷ�[x@O<Ƒ���8��rb����/�M�_7���,�ܻA���އ ������?Y��W��C�����Q(�1X���.me�m��