MZP      ��  �       @                                     � �	�!�L�!��This program must be run under Win32
$7                                                                                                                                        PE  L ��5        � # �         �           T                      �                                       p     �                                                                                                            .text    `     �                   �.idata      p     �             `  �.rsrc       �     �                @                                                                                                                                                                                                                                                                                                                                                                                                                ^ӭ��j�ᨹ�vS��>U�����)ĵ���	�.�-��x�Zo���i2ƅmciwr&7���o0��_|�uH+L�v��1��R�Z�F����#-��@�-�}������$�/}~���[1Ez����E���ldX���FSN��kVἋ#�&cG1��drO=��O^��ޣ(W��#\;�����C��u�#� ��e^�_�P�S\b1<��qg�|�]}�al^.�9�A�FRZ<��pFD|q��uO�&���
99�N�@л�FF�J��:�p���Aoap�*-�*���!(A?{h�1�l{f:~���tP�I���z����֥����ݷ8v�G������*P���j3��7��:���Eލ�ć�P�p� ���Q��,�>Qx������1�.����j�@���fzćք�Z�lC�3jaMx�Jּh���*��
]��ͷ'�����AҀK\�HM"u�Tl3wG��Jw��p�
N'��}J�t�ώ�Q'W�cJ4�#��.��*�vJ(0o	����7P�|(ֿ=�mh�ٿA�c���L؀8T�iQ�}���_��qg��%�䜟�SǄ$�o"R6�|�CL]�H!�Y?���\n���
z���󿏜_^�"�w�ɛhK��ix�g1J�G�ͣ`KJ�b���l�e����x<��>��f�-��g_6���-"��@:iK�_�J	M���xy�5����iwG�P4����IȱR���NZzf�vs�a>�'/�����@^��1�����I��e��-����*�c��H�uo����]�n���]A�A7O܂�Ҟj���krx.u��l�Hٝ�����47�[JQ_Q�({m�%~���~Zն3X+��|n�_��wE�nj2�(�H/ۯv�xJe&��G�+���([��Wጕ�b�����5>v%Xj[��zW ��(���Gn�&��^�V
�A�F�i7��˜���5C�P��� 0�3,��1�ps���EM�|�`|��}3�9�ql3l/�Dd-�W`M�ΞI��-�Գ���ٸ-J���pɳP�R⫙I>��K�^}h?���>�]���N�g���J�b 	��=P�QL�/R�u�ë@�A��D��>���Ə3b�b�����T�糕<R�g;�T2���}��2Q5{�n�k�,`��P�������jqX*�1�w�F���j����^�>�+���L��'m�n�,;!v4����5̝c��>6ODR�mY�l��J�0	k�2��2�m����s��x�m�/k?*k;;d8�&���[.�:j�5|�%t�"9��8�۽�K��#��V�pr�qG�UN5�T@�=�I��&�Ӛ�]ĄDu�d|*<
'H:<l�aW��p�q
�N� @�h#��A�m�Zy�ޣ���L��Z{�{v6n]$���<v�\":G3�U4�~x������_��G<}��,ȩ�Q2����-$���k�)Ӂ��u1���]�z�V��d� �� ����cv�c3��� ���եmY�\�c��~4>�&"�nKQ��H�Pn[�"��A	;e�cG�(I݇�YO�ŧO�a�/~���i}���G	��)�))Nf��~�6�D�)�a�Q^mȅ/Z3�*d��d��1�>���V��4I\�_��uS�/�ۊ�J�=�:��7�\��v���9rD}�G'ٯ}�1������j�n��EOlv���P�V��O�ۖ�]n��ї��} ��_��(�/+4l*z#��!:]��/�7�R/�Z�.-��@8P���W7��;N�����<�p����f�J�-�#b��)q��kT�i{5+��:��+��M_~k @h
Q�M�M�oa��=EaD�����,+-j�&k�i�й*Gl��u�Wڙ����)��8����	�;!\��>��Z���2����1�K�S��8�(�W.����:�fh�h��g��y�Q=��X�tO�S�H�bDP�I"F}�J�͗.�>��#�P%������|��<��w��fx������ݲs sɼƓS��) �@�5�U:��H���Rr�5��5��5��I*lq|c��.�"���k���^-+��� '�Z��Z��+�$��s��9�s�ض���lB��Bh���C����i�l�	]�wd�C� [I�����~EA�E��;�a�J@U�㸧�d�zI�츓H^odxHG���b	�F�&M�����P�yE��&z���G���`�&����M���M| ?;%�?Q�.�d���{0��,���S�YA3��o�**6�pƕ�35a��)y�M�z�i5�r�'��*@[��Ғ=f��q|��hb����;D=԰�l:LF��ۈ����nC�fzr���׶����-~�:I+|`^�۪�!Dv��ioLcy�ggD������7I�w��g���Ԗ[s��gu�7���/���	���*ŬR��    Z���DLquRJZPQRS�D$PUVWpSf�� [xPQ|�YXrfۇ������Q  zy�����sV%����^w�� �����wUf��B]~�� WU=�K�;]_��   f���f����Z=�^c����R�R^ZQU�J��]YWQUf�� ]Y_UV����^]V��    ^f�� �-����R�   � Ơ>������m�gD�W��Jϣ���ZR,$Z�(   ��m���c&���{.w1��Y�vo��\��&��#�u [Rf���Z�S_��   ��� �����y �������<�ŕu�U�4IAVUf��]]^P}f�� X{Qj/YY{Pf��`Xu��!Z�(�"�W�>1�_Q�[   ��n�+j8e�=3��芗�IO����/x(�"�LU���:��R���`����
Tm��ŋ���kſʒ]�+�D~��H�2����4N���YYW��S�楇��_��QRf�� ZYWsf��p_W�	_��������Q�Ɂ�����f����������Yzy�����@��H�������{�G�sd�w�F�Yu
�A�   ����L.M�R{ɓp���^��s��MBIrf�-!rkM�}�����H��kjA���������8�]�{�t�2��E�4O�E���b�Nd>�����27&����腻�[9s��*��}ߡ��#�M��6k�9���&�EȜյ��4�YnS��   ���⺡��&�VTϱ��Y�gJL����6{F�$͟棃�YEx\�$)��h��WV���-3��6����_]uM��H�o�F�:�$))��S����S�S�����mJU��m�ʝ��]�F�u��D;�.`L�B�Q!ZC�*/8�bx��c�$�����gM�Ч�E"HL@xG��{D{M�r�d%��[1��8���W�����V^��OP���*����IY��
�M���9��b��	��0�(���0$k�}��3jI�m�J��C����>�V!��f�����!I��QQMgPo����=�b���)7\�ޜ܍�D{uϤ�3�S�Sa� �5�y����e�Y'b����2l��[ÑF()/FŖ*FL�2���F����>�2�D_�z���{x$�`'��B�ϼf�a�jS�Ɇ�[α뾹O� �a f����E@5w�m�0J�f�z���#�[� �D��7\��EG��/k��$���k;o�F���6te���;�����{vQ�����L趌ŝt\8�αK�S.v�����qu�:�����rϿ�t���(mj%x'
E�5��h"3Ђ��/;��l�d	+����!��W�\����&�:��B�>����+a��7�6�&�8�w���U?}��H���r�����]��^����Y�O9oH�*�'�|o�k$��go���M��7>��|{>g�o��e���J�>�ֱkCZ�
�x�H�|����F�k2����$8��]��G�i^
��*θb���._Hb����Sɥs�׀�u��q��;$��{nrj���j&���,��6v��bK�c�h��F��LV�WM4���Mo�����r?g��~�@o�C^�	����X�@�z����AB� u2��o@\�O6}�h����k
���G�d���>��bl~Z��M(a"�sģ"T`�ߵ9r��(�z���ֲ��G�j�|Lv���!���N�:��N�$�'B�]ߛ+�b�P���?�85����.��H�[b#����?���p�E!.���C��и���5�f]h�M�sJL^ߋ���`G���uW�2�㥮���`�o'�IE~�Xb2$��������n�B��5�[?ܞڦ�G"8�ڻlI3"��rR&�~�_���u�,����te�1�Fj^������rV���N����8�!0~/�ͣ��`����Ȉ�f@g�f��-lE>!�1�����QU�pG��I��H��M�-���g�+壌_!JuG���$���b0;k?�O�������QԬ�S��IW� w�Ŕ#��]4;K|�K�!g?_��/�*���d�:0<@�鮓��
ơ�'������$yyFI�!��3ˌ�9Ml>:��vW���A<F/΃덖�'�_�8���O����_ms/4���`6��O v������|��*�-�h�0��f$y�4��{��y�I�ͳxn����n{��#��:�H�n�5�O��p)J����MF��]'5�Y�{����m�����	�8�q��+�:�ss�`ŮM�|��qѧ��~�k�\�	��Q��Gb���7 ��&~an󾕣�����%eÅщx(QV�E��9s}
���i�{��V������H�KQ1!���y���{���$U^�:Ư�>ml���Z�{EY�վ���O�+�~�pUo�g�Q�Ē	)�.&����E�v�|s���l�������͑P�צN�M|��3H�	�j���dp�t���zc�`��zϴ��i���N����sB��&��o�'���x�E
����ح�����l���&����YE�:�*�i �%XW�L���\ n!MlJ��@���~�H�%��z�E�E!E���s���8D)��rJp��P�Z��s��nN�Vݯw:M|ț������Ͳ��R�}���/�IZRL>,4�B����L���������ҌM;�Z�&�`(��I������
��<Z���1NL�~�[���0�D[9v�Z���A���(��C��L�Qz�>��Վ7H4���j�ol�x%'k �ȑR7���!�1~]�pwX?���W�i	��[�W�L�r,���m��*�B�V]�?Ў�x{�WW.�V�����ZLO�*����7���N�K���9)G.����9lɸ��9]�Q %��0��V��O#!�+��*�&��"� uo}�ʿ��#8:�2�Ƈ �hD�pyP|Ch�a�fa�7r�Ho�ҧ~���P�[ui4����\�3 �x��$ܾV����5����gv��U�r��5�>`�mU{XNkf�o+Tr��t6T�i������UdX����-��t�]6�U��`c�������Jn,���'eq�B(4�YkR��f���f4̏��Y�r[�>�mh¤��n�bVW�=gv�����+�
�t�Y�#�A�a:~m73��-�V@{���L@�w6XB-\��w�R�(2Q�֒�n�Я�G�>��L�"���[u���U.Q�1r= _���ں��a�	Gnw��B2����Bt�)_F�r�3�+Os��`�kB0���8��v��Ҟ��S���L/�V�_�H�I�/�U��P����0�R#���� ��v3�����d�:b�l�yꞭ��c��(a%��47�
�+��'����ϧ�����_6z۩�۱�CF��3���^Ë��}�1F��,Aj�U#֦���X���a��#}�,�~�dF[��RK�#а�>5Ò�@�ܳ����o튖�����e��nO�oC^zA���Ez��ț���BH���R�z2?�I�hKT�1I38�|[k����YU���h'G�qew���X)+������&'_z��/32��d��N�U���	U�p���kuY�S�65���M9��Rs_F[����;Ĳ._��c�⯑$�P�f⤯����yX`��Q���M)��_�Y3��h����X���Kk	D} U��}1-L
���\2�C���H���a��ꅅ�_��zXqHƢ�}�Cż��w�&�gՓ�l+�i?�1�<n:`|�R�H�ss��s����x��b���s���m�F0�`4h��II��^i�k-z�$G
UӘ0c�2^����(��PYT�]��7����ⴗl!��F�0-|�9�V�tQ��9uf�� ��#?1M]߈-:�2�oq0��lik�S�Sl2^z��,}"��%w�{G6��X��%E:\��!A(/�P+VSU�5 �}3�ˏ��;�s�7�Y^���2D6$�z}���e�,`o���؎��F��~�HF��h��X���<�X$��cګR<r㞧��g-M���� #���v���5y�P��e��RJ���|7W�*�js��7�ӂh�-��p�6�n�=6"�+v)�V�G��)��*�ҩ�/��M*YϴI^��~ͭ����	���],������J8���c=�ZuI#q�,M4���j!��C���Qq�vq�>�~b���M\���
/����8Ҽ�`��.�ܑ��5K�O����'�j|q��k%�S�=5����J�f���.���@Φ�[J�Uؓ�,I+�r0"O�+�E'�t^9#�a�}B4�N��%B>�	��l���f�^5d�dg ��1�����Ս7�o~g�>+$��H��U��*�M9Ґ���l7I�ג;�����0�bS�nM��cs��.����Q�avEH�ex��q�3YS��#�:9MϊA�!��QX�ݙ]S�{٪|�"G��'�����X}���	G��`9I#��y�xq����$�C_�[peS��B�1�(��Z���I/{�{� {#19�����Bq@$%<1��_^�	��c+���è�S�:l�,��ģm�j���u^I	�ܶ�5�;�E^'aQu���DR�E�ZsRW.JM@( E�thd@9���.��$0-�t�e�L9Q.��.�*ƱL�<W�$����� �WW���T�����"FB�D(�,�DX��&޸�)1Q���
8�_
m��Q��]8R�ܖ�i+�b�C��f�0���L�%���b����j<�M3��4�Nο�^#-8JQ,�>}<�~ͦ������T=|[6@��8��̊YW��~w�>�4�B9t��VqS�'����Լ�U��o�pwbH?��j#�E0�ܰ.�ŋ��l|g-������y��@��̂t8)�%���	�E�fP�X5�h5\�v
�jv��_u�#&�6�DLt�R���z�9l�.z�z�pjȃ%ֈg��?���z�'�M�(n_��a��uR;�y@;����m���?�M��~et)��ξ����*��C�& m>�_���Q�a�'�U|Cv��{0#j��
�6�?E�}FG�,���G=�-�Ci��֟f�xOe��Tj�R��ohͦL�c<�~��$7J��6��8��|I��^NƷ�Cj�g�uҘ�V�2Ct�9@&��g�E$����g��8~~�D�h��>��GnvE�b:��76��p�R���I;�-q��߱?6���ã�s3����yR�G�l��# ��Zs=�J8�:���Η<����b!�m��SW݃e��h8�1����h�g�+;���ʜE�g�
S�n>�WŮ�E[�?�($>%������`1mj�4G.�#�q��L�8�w^t�-�vAv��ڹ�{	��4�/�L�al�l�T��"�YJp3���b3_r�%q��{|�cR�(a���j�?=;�j�6�Pⷧ]W ��S��h.��#G��$���J�\����1�+MZ���l�� ���Q����Ȑ�{L�]v��;`{�\�a�Z>D�B5�<�j���-.�h#��=\�_��\��1a{�2�����M�l��5RIDq�f���17�-�|@����)����C�3���Z���/��;d�o���@"�q׻.O)Bt��+��C���E$2��^�;p`.\�I*�Pl5��[�ܟK��ڏ%(��}��YZȘ5ZgL�3ER-�t
J}̿��� ��l�h$���Ns�tRFG��@��H�^�`Rk���8c��Z�찹q���(Wl��o�tn��8$>[����Ghl���L�SRW�2o���G�/��U�*">!۴a5&��!�7
i���C�9��	i�*g���GL�
�ӱ#R�������C*��pe-�<h$���'Ǚ$�m�ÌӷD��ܗ�pr�QL���
�|�QP�(`��_��8n���a�H�� d)�O:���ka�ګ�<�<ז�J:7��5����,2�)D�W���Uv\����p�-/E��<N+��N��2�3.� 6췒e�Mr:8�������t}��A�5U-+�Ͽ������I J��I\cb\"P�F�'~���ǐ���D��8X��I��5i��<&+/�Kȥ������L.|�Rپ� �����Jm��`(w ��,I41Ŏ�r�焵��<q�Jn���%�A"����m��L�����x5�DV���G�֥}��N)jrh��������X�v�0;a�<`����9�]h��,P]����%`NR-�֫pi?㯳p�!2c3��
m�~�Fl2�����P�+�ZMN���1	��4�Į��"�]�J�|�	�K6�;7�"��|0��d�\GO/�r��c�/��f�Up�m�z�	MI������t�-]p;���p%=sAُ�W�+�w"`w���
i(��)�<�A���ƨ�a�'���u�ǧ�}L��9�E9��C�_�� A �����9\.���ė<���f$�=%:?��ar����H>�N���Ix/7n'�y�/� �;�f��t����Ns��8˽�)Qܺ�a:+��/�h՗P�Ly��I���fb �3��,�*���2W�ؗ��N�&*�R^�T�r�~��dW @��)=�+0	ST�Җ��vZ&�s�n�?�o���Ww�gcى�z�]"��IB6v�*�.�䎛M]��E?R���x���a��� fFg|(P�Z��A_�HոVB�@�o�o0�?����R�~4oYCs�V��o�	�j���ۂ�0��I�Q8�H	ᆠ�ұѝTH+,�e���<%���[����臉/_��4����}	�! g8���趉RK�����c넁�_��dl����j�a�������*|$m��XF���c`Q2�̑q�`ͻplγ�fk�T_��(f�GO�p�n�
Z~�޴u:r��w�El�M������J��ם�]�����i��C|Bą��i�	�&#_l�eN��<�m�b#q�$�>z!��l�]݆��N��>��9�L ����`<xr�W����~V��������_���+ݾKW���Hٛ)��ܭ\�TcT��;�0q}�v6T᜜}*�ʴ��{S�l�0�\	��g�B�}S���\��1�0�Ʊ��Rk���1XG���i����rј㊕�.M�_M�˟�쁽i��hs&m
{��'���9t����u,����oJa�J�ui�"B�f�!7�?v�◛�	�4��岠��Y� uN����e��4t�N�X�����l�c)���FRw���^�m�}���+~	�0g^Q���3�KkOK���k���9�n�B�b��l�0F�@e�[�@<��z��A���n_�0&�_B�:�҇T ���xn�B+�����50���g��5�b>LQ'�z��z�hɔ;�M����OX5/�8���⓾�٪Sa�7�j��� �/�6Ѡ;�N�v���-}S�6��cϧ�_l����Esv|���f �z�E�V�+��rUF��,����!�
݇bB�r�,���^iբ<*���W*XlD2 �����^c�U�������yK}	r���YY$�zH^i���º�V��=�T��.q�7LԪ��2��������ґ �Hy%�k�N�L�֨��F9j�1 Q����N��	iZ�-U�KYFG�D��NN�',}T���������LyI�%	�mL7w�w{o��ӫ��R�{�8�^j���U���_0A�MB̯"���gj��&��`�'bxߘj1��x��Q��h�/H��6�cc0W�mFs����3��+�[�VP�� ������d��SI��tS������d.l�k�,�� �vlvƌ�XD �zE�sY/�FHz�+ה�'�7�gڗ!�P:'��$��@���Y/�v��朆��W\��2��W��[�t������<��-�N0�.v�f�s�ӣ��]����&&�Vt.�!��xUG+̚���H�����O&p�;��(iMhQ�����Fx�[����=&��ם9۳��Nt�PL��Z��W�;�U?4KY��s��!�DhЌ�&�`ͯF}	;oiܩxnQo��h�?�2��N��,"�4/�č�Y����b$Vg��m$�F���+�W6�ϟ�^�8q|�@��m��=�VM����qeɌ_�̡��*KkĔ�?7zٛ���gr���	+q��M]lI|!�Qb�tHg(�����cDﰜe�
ۤT;�n~�gwá���(Y�`P�U(AC�@,߰P��=w�ʭ�Rt]�T��)p�v�Qk���NI�<| �In\
��Y«���x,�ueV+�UR�2��h���b��۝�o�^~����EO�K��3�dv{镲ٓ�B�}�+�=k�fp��]�?���uI&���[��D�x��[}1B�f�qH�`2�} ���H�C�2|�l�$e����VG��3-
��U �7w"%��Z��?��A�*�eq�m'�n˗�7ZF0��^Ì��q��W�$�E�^�]���*/�܌6_D+p�����S�WP��@�C&["��)*���T�z��q�IV�95>ћC"��b�cUh�cM�J���ڙ�I�D�����I
y���Y��r�:5���o�kq;�0Pۺ�2\�~�?.!|�y�-�����~��W!�1�St�M�FB@JR竍�����/��Ju���<��)4v�<��y��L�¯�Q�Ξ�>�&Q��a>�
�E����u;nL@��i��Y=,ıcO�2e�?�#R�=�/���~�+�)�@Y|��լl��ճхa��5�(K�"�]�B������q���5ң��v���"6�����ɡ�4����Yd�X?���i^#�6aWpn�}A�b��ѪH1N���㌼0"�@�_c�0m���J\2n+Z��0��uJ�sc�Y{�v�Ѵ���=��\�$���i&1�W��C[��|�I�K�<�6�(H)��c��	�x`6`�J��'�����Ģ�B>b���K|0\a�s�@4É=tw_ي&A��_{u�`��n<N��� ��Ȝ2!�k�<���Y�kKkK���d:��t�o�1��;6GFg������A���^$��$��M����iH�Y���"E\k�G�A�M�LƓ�����Ϛ;����<E�Ù��g�U������4Ҵ~`�$�o&��TˆW\�9����H��������(�W׊�>�e����D��=ύ4�w^����t���m���^Ӝ��4��$��I:!F�'�iY"����J>�I�p�\=��VUN,�$]�=���"u|?+Q_�YnRyn�ìetLQ��u�v,CJ�k�2c����4�}�u�����&ӂ@�oά�+��m�r��6�d�/��j����F3�t���>�)��}�����h5�H�O�?w��c�'��h����F��m����'�)J��DZ�bd��@V�K餠�;'z�|57�#�\�@L|-�&�ng0bO���J4N�p����%��DT�}�A�a��ț;,IJ�%��0;b��X܏.��1*=*M����y��y�N��M�����9+��K�`6ltE����K��í��B��%��~��
s:z�׊�X�tEĖ浯\eXӖ�'�Fw���+�>Ըd���˿Cl�v�>��?(��h�ch�-��,�f6P����37��!��3b�By����폧CR__;M)�������R� /^N�����ޗF:`�U�{lḲ'�`t���tZ��n]�Dcӈ ���P'��b��`�d�Ǩ�T�~e�+A>z.H,y,1u��yL���Κ!d�#K���m�Ƃ:�+Պ���	R8�o3��-l��τN���W�b��-�s�m�'$ ��l������o�3����ʡ�1��X�����S�/F?��,�x6�r	�"e�Z�1��8G�*�vG5�l�{;���$��T`�A�G�Xx=��w
�)m<���9>�\�K�yL�-��������Df���1lC5�E3�|� ����)��t�Ҧ�t�g���ϴT^�4�,ݻ�H6���i���%e��0{ (.,I����i"�,=��[c�_Ҧ�s/Z�O�C�-�tm���M�M>� (3����|���o���a3�����/V!��ݗ���/݉��O\Х�y,5�J��a,)�T切�Z��ֱ8?R+y|�5.�Zּ'�x�+�Di�0��.��6��@s���f�	^�4[=N"j^^� �O�S������E9� ��-l�d��JT]"����);w�i��\k|���x]���B���X��L
=���t��3���O��ǼEL>�����F�?��c��X�b���A�H^�����x��n'��7/Cut��ąj�"�?�� � ���_�\�1�`,9�,�E��0�c�j+���N��p����h�<��
|�0-�J�2�r5�V�?�X܃v��ة���7��DF�~��]�U���Ż�V�G%�����{]��F�,դ�&@��^����@1����F���y��h�f�)�	04|����,��x�r�V��o�9abY;��aA*O�;/HE����o���=�ɔ��hqՔ�T��ypg��m"��^.t��l��/�Z�zQ;�w�ɒ�9�����X�9��<�Џ�yQZ2���2}�q���Ҕ���YOAȩ�eٲc	�Z&�6�pl���QR�	��8�_i� y�k�G���K���g`�?�󰪘 u��F�axA�#�;<��c�6��㋵�a�!5����tQ��F�n������������
�M���uo���C���Po�
��j��:c-�-�6�Q��o���M�&��Xr���aI�OH��2��v��	���<ka,��L�u��|���($!����e.��j��-j�șW�c,	�m�^�:C	���H���%�s�����̩�l7��u�p4��5�+ �J8�����eC�2�fKP*��9��!O�$Ǣ���=��͙��Ͱ�����M^�P�Q�A�!be��!�A�iP�[�l(�tAD��:
��gvã1�ˁM�����,<�_��O�d����S��_-8)y�my�>
�V�2�<��Y�X׭�ڟ]�id�<f��(���5D�d�2��g>q�������G�ᘩնl�54?���́;����=	��P�L J[���h�X�q�i����K�����?���M�1�.#a�Zr�����%��+�%H�oE+t݅����i�)m�"�Ҭ�%��l�RI.�a����t���3O@�Lv�@�9}�y�'���戡��֎9p#��^c�����%Tď�%E�g%%D�F�}����^�nqH����td�S���ۨ���x5�����]��<&�mE:�(󅠰/eG�N�Y� �,�+U�_>�B���-�k6�Td>�\-Ŏ����(�0��nMZ#^EF��&�m�W`��(�hdȿ�[���,\��]���Y�z.|��3����e�P6i�SeZ^,0�M/��!�d�I��p���������.�*zG���\T��j�A��]V�ԓ�2%BSNԺy�¼�5\��6])޸���{�{��~F��$O��O�����|��ԛ=d���+���øՋ& 3�!�v�@�_�̻ol�R�Y�md^b�?v��5�>(��B-~����;�<�81��W�o��ܜP/�.�r+��Wg�h�ōH���zⴚ>,��tc\+����Ge5���#��k�^�����1����̲��%k8�w8r*����@�(SZ�hb�CTV���fp���N�x;/F���ӡ�a�VҎ���t��'�jAD:b�@,��B�BE�Zi��>M��I'1%�to���r��yP���I�7�-�&R�S��GH����T��2�I�Έ���2�L� 
p^��x/�ܪ,4�7�%($z'�g�+"�'�q�`�f'�zVJ1~��ì�֚��H�^:�9�O��8,\VC�O1R7�g�p��Ϙ���� �#��{��S�5�0.Z$Ӆ_�v���7J�\`\��*�࿶�������ƤT)Z��IU��0���~�S0Fs`oԋ(��e�ˍ�4L-{R%�hy闯�I�`u��V9E5�!��2���М!nm׮j0S�4� �BJ�d�����Տ�G�D`T�>���z_r�E�ڳ�O�k�5�H�z�^��e�zRT3tY+e|�|��;���x�hϴQ6_��@�
o*Ζ�� �Ҫϰ��	���p�7q/E�ܢ)�Q��I�K<w;�IO�q)�"�^#�>�d
�N����2$��<;�@'��}�;���F ���W��l���}G6���[H8KT+p�)�.avraI[T"B?hVJ�b�4pzd���b5�@�����,�;��L���1+>C�J��=*������X�|.��5�[����C0��T���YR{I�2�^�xeQ�y~�k���N��#|�뱛����,EX/l!�(-�?� ��_�\vl�&S(Z�i<��RB�
l'~t�~����QEǲ"��.�s��7���B��\�[5$�pTy��H4˭�1�vO���s�Mz9���Hs��f�� t��/���5�;�\����S����wSz?7��i�_�E�)SԘ��\���ǎ��$+��#�����ލ��=�-���tv{�N��΢�=�2���U�x�������kuO({�6�m�i6�|ߙ���%���<6���3� ��A.���D	���mBS(�i��T��
�^W������AН��h%�d������e���Z�2�Ο.?޸�;�{E����5
/�gR"ڥ��#Vu��&G��W�j���9��_���.��y�;:�aN�B1;d��w��tH�p(#��|]f̳��8 ;�{r=8@�G��S��3ې3咍y�����u��Ð�{M01*�46�����?�h�/��&���n�AI�U7h�73��n �o�?O�}���v~G�p�������5:��Ȧ0qm�L5�
6��쨆d��;�jN~HD��w� �I��CZ7gz*)&T{��E��r�\`e|J��}�ٟ�b�:��b��u�d��Ś2!0�|���r�6܈8n����ɮ��W��h�Ƀ��t���d�y�vM%��"g����ɵ}�D��XI�8!)p�ã�����6�$4�xaȿy�T�?fru��`-1��snM]rH�NO>O���uN8�U[}�%�PE��=D�����_ߦ��-�9��.�"�	��/,��ȿ}���4j���gWQ�!�<%��Hq�n�ǫ{b��^�����P@ً�n�4;LC�m�<10��M�X��sݧ5�f�K���Nui~�[��G�ad�$����݃|�υ����տd�)�L�y�E&+4 &Mɉ'�(�E�� �:��}��I�6�R��I�R{{��q��5P!s���Ɇ��l�d��+P"��3��D�w���-�~���]ڙLg�p�� PD1l8g�B��%��=ms�h��ᬷA�i���\��Zg��)%�ɘ:1��۷�J)���_wfݵ�@��5�1&0��^��g��шۮ������⻅T{�o3\��&^��kjh^�5���k����"��䐮0(~��o���W^ZC��ipr	��d�F����cb��3r�{�.f%�܁s��J�`��б	I�1��J�Z(�8�?�[S:��"[�8˓?��&aW�t��N��uy�]�L@��mU�z�#.��@�Z	˃
��ʈ� ��[���_� :����5L�[k8��_C���9�X����<���/:G'.+ҪoY�����k���Nx�
.*�mWͲ��g�Ϛg��Z�̸���2�S)��T>�)�uh^y��/���`���i���k*�F
�2/�QM���O��������P|��� z���vg��A��a�4;�N99Ԡɹ0"E��ץ�>��+�_�@|n�S��^Eu�-��`�'�'�C�thV������T
�)-iE���� �[{2@b�x���� M@IkG�^Fޟ�oi//r���!{�B;�3�Qz���E�=?��_D�>���є���D�{&)��W�8��Un���1��K�B)h���MX)W��0'15���֎�u��f!R�����/�z�<b��:m���e2X� M���x5(;;��UQ�L���7�`,���~�T�����l�/OJ�}/$���$�����*�=�%#��B������I0��x��;`��a��F���O:L���Џ�j\��U�l��j�
���#�d�C�@B4?RG|چ2諜��S���r�����Q��������I2<��Fن�����4�}��XqȭĒ������oP�� ��Q|/�#�:��P��6����4����)����1Ą=sb�_S��ݖ�P�� �2�Ԍ�C���<k�����K����ʏ�E��GXJ���N{L��7�M�8өc!���oq�|�N
�ͳ$�8턻�ő^i����]ǉ��ZS�_�=9���V�ƪOb�X����>��H�H0���oM�����/GD��U�<�� �d����&>�<��ԙ@����:�r��*�>��t��1�|i%�-����"�qgu/�2Űf��ٞC �5��I� �р[� ����7���!���ܜC��Ԗ���e��	 ���y�'wM`�^^�"v���?+^��(Jy(�cL
�4�Ǫ>�׃eŋ��W5�r�Y!�.;��rm�t�p�A߳�0&40�����rRf;��6�6�}�S�g�M������Oy����H�. ���\s2lS��`�o�?x�Dmi���8� ��DʶΛ5ڦ@.C�Gt7�E!a)�e#�pہ�9A�+>8|WE&%a)d�F�_�_V^�/-�n�����:+���R,�븆Mt�p9@U~�S;c[U��C�)�.�R��)�P����"7�tSJ4��8v�郒X��By8:�X!�t���6��&qƚ���rr���AU��'9>���0�30���t��}�����	�d��mJ�v�B�#�#|�1�ъ������ڭ ����rp�^5��ի�2��p|V��/�"��3�C���a˱��2G!n)`V�pHr���ÉD�!�+�ri#���|�T�΍�@��O��͠��cld�?���<FDӈy���*�M(�\�S}o@9����J��Z���Ҟ�S��������������m�Ո�;S���P_�a:h<��o�Vd&{����Z/*�G��blA^�������P�� �I��c G&�Ni�E�X2���ԁ[#��(���'y��_�2�?<�v��zf�}r{v�Ɯ���\[��H��gK-$r�A"i&�`x;���U?��튃� ��L|��GـⰄ�\H_P'~��Ѻ��t?OL���}��m�i\f<Vwp��vY�H��Cbҽ����sk �o����%a��]����-Kyy�l)Z2�0�C�N��z&!���_�s�N���(��Ł?��s|?��:��%�Ϙ�}E�����=���#��(ܪg��I�t�,F��V�"Zۚ2ͯ	�+3��c�2���@���ۆб 6�u�f�˸	!b���cU���ώf���ikOM\4��[k���S_�d�sc�[)Aǈ_�o�Y�6����n]y[��+[S|���8����Iw�ZHuSM9~�=��� >�f/&q�anP��?�6ft'3�sRB%f��@�'z�^�����3"j���=p1�욄\K��BS���'0��Fp�]ҭ����n$��h���f��5��=q,�qPw~�1�!ά�v���	�y��<���8W0�RCu������K�v��OOj�����?�a��u��T�C���?g�7Wzk��eX��|�R�H�[�CyD����K>��q��*k7�}��j w�
;e?����̒������f18���^��E���wL6i˞m2�~+��`���;ӝH{	5�jf�� �ހ�jL㱅4�6�sUrKd/�������4��rcYfj�8�z�����y��z,�F����?>p���]�T	�h/��~�<mġ~�l2g��[3���_�	c��޹�I�y4�����D�3�V�_j���q��\�Σ������x�n�8y�/�0�n"�wqZ�o���c{ ��JD��9�IˢO5o8h/��p�75�Ѥ'�_�!{5?mM<r�\K*���%"�<�&W@��C��g1���an���i�GgC�\b�؁����k�V��z�|��~�_*���>{����p�IkR����e�HfQ��U�B��q��F��#�<7��]��C6�����	;>Oa3_��$��P��v�f��ؽ$���)[�T�G��cR���4�i/�g���%/����1�q�Q����,!�h�o8��ؖ�#7	��8X|:�k�~�uY︩�6�G��u Cq��P�nQ�8�:
��O��X<��	�$V������r����g��E�&��(��>��t1�6rA���Y@�葻H<�v��E9��Cx��TD4�h�W��}���� �V�6�K45�T-e��dA� ���������{��sw���R�G/���gf<�c8H28���l�B�B�j^DF��9
1R�U'�+1h馟E�hT)>V0�Ԯ�ȀK������8MѦ��l��A���s\�Z=�o��*6卒S�	5'ޥϦ�E ��!�ckSy+g�UϝP�O�������ɿ_Ճ����i�j�g�]��5B���%
Eŝٷ��'�>t�&]�3>�ay���S]��f�TK�DaYT���\��I�UUg��]FT  B�.�$��g�o���B|��m�k������Xjʠ����4�<�R���������g!��Q�� ����A�B�i�Nc^�Z��/�k����ad��r�*fW�S�`���3�\�ծN}���C���D���e�+��H4�M	9�Y����HxF���P��2�VC�����������ooN/]�Z��x'�T�����eN������{݀8&���2��g�t@#�E㔤Q[w�R7�� ;�P;٥0��VBw���$5�MCLM��+. ��9�eg;�X�%��1��c��tVn9o[�=$��8��M�6j���)���i�K��z~�n��:pgE�V���+�0�����J�3J��j�Gd�/�P���}T��Q��;}:�iG��H�c��}�zT�����.�Bʳh!�貰�&`��/q����E��S�
b��2y<�+�a`�KhNl$���e20��h^I��:�~�����g #��A���Լ���|���Y�HB���2�H*�(���|Z�|�%.��i� ��N
JB�1�2���b&�
�1��L�t/�d!/�q}̣�ѸJX� ��[%\��l2�	!]ym��Qv9����M�L3@�a�@	n��l�|-&PY���Q�	�X���^=��R�u��`,�$�KP����é%��8x#�AD8���oJX�����9���7�e�d⪽�R��;�hs�U�oq��飕pj��9���t�G2�PB�� �k���e��n�wX-�V���&�,E����P�yN��f�}v�v�N��F�!�>%��ȃ͔ډܹ��Y(K��	A'��^+���2�n�.�o_#Û!����ZÐ�"0��	�h���!Ii���劧���"r^�Dtjqlb<0��^ X��9�!��&ޢ($��~��4)V�(l�Ȧ��A�
6�Pk%,Vm������RJ@�?:�*��c�G[��?�X�H���E�x{	Cz�L��!)����J�)��#�'�����-�Ya���9F�y�Xa�0	4���l�f�oAtz�8Im6�Ơ��0�VA�C���]bl����蹩�
�F�h/Ird����=8��Z"ޓ��hi�"L����%�e/Z���hoo�>�s�3E-"�B�-�Mr����-16�o�����J?�J��k��.�\^f(�q�L4����B귕����8�n� ۸�ؘ�Z{�1���e\,%���̈jb�e�☲�uج�$^�ۜ��a�g7��)��+Ydۯ���g%G���/�_�6���k8Da��m Y��N�K�7��!�:lD�m�e�WZ�?\W$w&�����A�����F��/�>.x)	���:w;<�+>j�h\��k��#�	v��3�Jݩ�3�����ɩ�,����C(�o5�����mnɢ�D q�w���SG���j,(���*>���T������]� U��]g��$"'�O|���[���k Ap�rc�Ӱ���1�5���N��W�s��)�9�[��D_�s�vݷ�\�k� ���G{���(��ҭ�)�}7�8l_�|�<��ygݳ.z�c=�;�&���o�9toy#�P3B[��2A2���J3��Z�炻�]�H���8�~���G����1��7a�ś����A���s~,?�"˵B)i�fz�^�cj����*�w�+�!Ƭ�zZ�S��alY0���s�ULM��Lb��$���D#���H�`+��4yŜ��gZ'�t)i�4�+�wI�٤���)I7߶�Ӛ�g��H1��tzEz@7��";���}(qU� �hb���6�s��Ώ�������|��/�t�hq��o��r{���x\�Qk>'���~��Ն^��'T+Rx�Y9�(C_E@sUR4Û��Qf.�~�{�XY�����mhwpG��,�s@�9��6aW�1����}��˫mB}�h��?g��E��l�m��� >&�:����0�)����H\�B�c�ZJ�Y���ô���޸*['G��Y�p�NOU�o�hT71��}Y�9���8sS�mY~ܺ���>�@�1�w���{�)5>�Vɗͨ���_�B��Ө�䋆6O��c�;�X��пY�f]G�+�ŝ�����r,^L�5��-��>�N�a6{S8�Q��&cN�5��YJl|g�I|�M�0ӭ�Z��?������y©�)fFGj��z���Ex�E�i�Cp1Y0��*[2�� �n��uɼ���[:��'h4��9��rV}Ú�hWX��Z���S�0�����*����'8�����X��ޔ�>ʌim��NBb�i�\A��"�o#\�4����0�7 x=b%Q΄Q=b, ;��!&?�G�pf)T���^���@Cl���3l0�Ǆ��4�Ф5�o���a�On+c���k�+J���յ`ÏL�zF�"i�Q�s�����W:���N�0'٫u�q����N�у��Ny>��D8kx�E�䘻����u����s)�����$�)u�I�I�Ȼ)�2O��p
�D'jt}I�Q&�����% 	ٔAo��p�1
M�1��?��-�z��N�fO���<ߐ �ZȂ�Fx������y0�lW�Rt�=�N.�:�̓8��+��Ye���{!G�5+���������Q�)�n����ǐ�zDF�Wά�F��[�!�9��d������%|T}et��.� �̥;r�!*�Dk̒n�|qwt�.�v�c*nP]F�H6��{�,}肧�~�{1ꭰA������Q�޾zz��&n�B�?ip}0G�*�`~|��]�/L��{w6�@l������7�/Ѿ4���ҠuT���`m�S>a���a>3s�F�jm�)-Ppz펜)�KiNE����kgc�(���!���$�T/�L�7�{3�d��b�f��oM-�2J�>�}B� +�u
F4�8ԁ����H�SH�����AY��!�ĥ���t$�.�B,[�_��qwH+Ѵ�)�����i����a��8����;'�,��e���qGzl�e��������I��(~0r�.N���x�U���DV EQ�;p\��^�@�G$�q����`��j������Z��✮x>k���2�T��۾l�yYFh��4sŵ,���ia����ϋ�w
숓�
BD<�9e��u��Fx�ղ
e���/!�d��I�`F����b;������[)�:�h�d�W8��9l9u��
3��}G��A� >�S�)z��Y-pQ�
�N^�����s�O7�C�M|�R W��)Y��c�4��)�D��������V����6ڤ!�Y�>�,��p�>-߇�����Z�2qۣ/էW4�R��C�@6�q�w�5L^j����s����5I7�|�VG�r��$P��,@O�螏��=$����fB$p�(���B<��x"U��|�y�P��A��Q�I#fn���ϛ��uW�S^'�!���R;�����ֈ�JQ�q��p�}u»ָt#��d���Q#�3��Y������u\�k�cRF�%xg�ov岭���	
�g_�bF\K4OJ_�-�ӏS��ݛq��'����ŧQ�
^G�,<R�MK�l"ܳ���]��Vѥ	��=Z˽�47�|ƣ�x-��ȴ,hj8�Y�-愜y|�������nb�q���d{t�q��A�o��Z��V"\���M��?�B ld������G��=8V�������A�>6p�IM�t��#��hp
�o��b���_�=u]�������>U���Ěy�S�ߛ�0��P*��"�qI�x䘴��,VO�W�F�6���R�ː�'j&`氢�Ԧ���P!2�?�A�$��*dx��n�QY�=�:�I�W�I9�"�H��}I�M����(I���׾�`���������s*��ħ,y��x=T<�}�oF�>��,��uJՆ
[�.I�?yv[Jb�2nr�9��V�xE��3vdL�r���"9и��
6����S�̭,G$>������ Vv8O�w��cF�8QO��H�v�"�n����^7S'�~�d�JC���ӥ��]�_�q��[2��������%�=/����.�}֮�s~#�Е�]�|=�)�
���9��,��V��8ę����⥼���8#*)�T��G
?q�)��=���:�N���Qm;C�!�`$�������ኁۉ�>�E�v��#���O`����&i�{v����߻Q�};�U@����#6�J���s�cqOuqm�K�w��k�0����\ܜ�Ew�g�g����bk�6���Sp�����D��a)���_Sm�2�f�4�cg:oc��g�$�^,�F�Տ0Ψ;��Ak���;�8i5��N�92��#�G�dr�x�l��V�*qfc
׭j~�QjمL�&u]4���9��`����w�Sv�y����7N���Px�}�$�95��L����D��LY�/�qu���K��:�r�O q�^MI�e]E�^ 6��Cf`�ҍ[u`��:�x����gSy�r���X� 2x7�_��j��?Kx~���c��%,2�ς!�V�ʈ�H����\��?T�?2��t�����ޞ�W��M�Q���)5c��;�����w�)I�������~Z�qG8�V�
3�M���y�}o#4;O�nl8�ݳ�x�5�5j��ygs��@{c���C��9)��7Mt>����QƓ�o}}�(O���c��Z؅֏���	�� ����K�N��)����+r'��f]����inN�o�|��X����R�{�S���io7�	�r��ǽ�cӟ�fZ<c#R3s��!I���c�F��Pv`��Wec��ޤ
�~�V���v��6VV4�X��)%�������&�n];�((�1��F��6f��S3���{��2^����z3{|)��Hm#�u�����b��놙'85�	{f@L�?��\�soH��Y���c?�Sp���OŪL{���e~��*�[N.V>�Z�֫�������ߪI�
�<7T4�Wr	�VR�w��
9�уk��F"?�O��ږ��T�H�e�=	�ky��X�}QY�8E\*��� 
'�7O���[-;���mY��=�"t���lw�	� �>t�t�_Y�T�lL� �<W]"�K�?7�9Giٹ6n1�J�s�u��k��p����u�!�5���-������J"$���6�ު�N���PS$%w��J@V1}蟫���*;0.��jOK���g�Շ;�|V��g&vǹ��9#4���U��#��1���8�G���Ah���xo-��;�J�?L��v�<"�5�x�
-�-#�,���ɶ�
������wy�l���mQ�=���t�L��0����ё���@���΍'=5�{�h�3��O�d������f�'�j e�	���ˊ_I�ԿR���:~a��)Ӳ�PO��������u��"b�b��Li�����٪*>�Xю�B����u[�* M^-	�suȄ�q���Sv��+�B�w�E���?��|����b���#^8���UY�V1��T[`��ɑ�e؍ex��v��EgHE�"�-)'z$;��r,=��rVzl�w?�Q�Q�4�$���J0���k7A�q�}^}���BW��Pi!T���h��ys&��E�S�6t bm3u&V�5��%	?mfQ�%uT+i|�<1�X�T�4w�Ix=QN�|� �AE]��Ā>����X�_��!m;�o��,�+��5U�Ws��J�"J��@*Ȉ'�-�J�$��k�ٿ���`׳##���ҹPk{\�kL��~~$_(㮙	'�����%:�]s�5�ᴉ�"j�����U&|�������5ߌ�o�'��N�Hʙb�.�P>g����╕B�h���ԡ�$^�Gf�t�@C�%(��>�L�G��0X�ei�����h���J�C�4�>�HŃ锶\�ήM`���
y��EP��G�p/�֧�1��}�L�7Lه�Y� 	�ǹ�=�:�")��iPb�� �PK4:l��PG?�j]�S��Z�#q~N��\Y���A��w���;쯧z;�#2��#x���2�)6%C���Mj|/�����>fA?i|[e�<�V�@�J��0��<���^��������x*%(٪�O�@�^Y�"R�	�2U�Ȭ%�L��{�W��Q�����'@�B�d��E9�7��մ���b�y�:�K�� #��_�T]we_��9a�_$j҅hE�T���7��<�d�]w����*��M���? �[���Y���?(0���d@Y"d^o/,�O��uЀ��Y���g/���/$ٸ��%����b���@�t�]J�:W7�D]��㠧�rt��K-@��8�r@p=����p�'��^��F��%�?r�C�D�4+'%�It��=��!�ԅ��!������e��S]$��l,� �X��}���e��3�u��C�&Hl顁���2�z~� ���!��������.l~Z�rW�7������I���YN����c���w*K�I|�'��F�M�B��އ�E��b��q��]Wp)�f�︄~߉�(�5���+� ���3��]X�`��n�
�l>"�~#<U}��DrM"�
/��aYy8Aǣ��մ�ȡH;���5þ���r�I�aH�*r�#2~��p�d�3�����:�"�:+�,�!ׇ�e�1�f�R���I]�
���<��ϖ`gH���� Z���55B�}��"���"c��$-�C�
�� T���d:�dMp�������F�U�`Pt(�Ⱥ�%��6�v�t�" ���^j~�����፦8��c�8��u�x����fc}HٙLn|"� |8���n%�AH����H���,^1M���o6W:�Oݐ�9��{%O���9{m�w8v�
���ݯ �ߝּ��I*�xd��,�)?����ԉ|�ӴȃsنD�!��1�� ���K�^ �+��(���e�K5(/���QSRq&2K]���=�2�x�:K��dB�`l|�I�rM>��b&Fޣ�_�Fzf���&O�I��%Aؼ\˵G� �QD?��(�.���Ml׬�aF���؉����w��4��JG�F�uNT�K���;=�2 �P�K��]�_'�|��ZsAGD2� �]Ԑk��i6�w9bi��)8����﯏W������9�Ԍ����+�ֲX�z �(�ף7�D�����G�4�K���q�zn��9i��u+�9��Q���Юuu�+������O|�"+ߝ=I3$Vq�tAx��hw]F�#���e@��βmwΫʊez  ��8�['�8�w
9vڧ��ow\��"��$���Xt��E@as�&�L����/�0�����]�v��Gf�v
�b��}�C�p�Q�'�p������>~�6/�&��k(�W��-���!��ʧ<��퀧�a!'�q�~ɥ^�v��\�Y���SO~��ݮ0�G,|�y��9���x���P쇗 ��̊M6��.��Z�P�$nw�a�F�9����R����!�C��M	�Q#�r�g&.�9�0��pa5L�[�7�R��"R��8�5,@��(oC��۪����ĺ�3��<{y�N���W
m���dD@l�n�ƺ\����R�ꢼCY����ɽ�2��h��Ԃ��l��+��>���_dwt�®��P�`\ȟ�հ�ݳ]��y�n�� ���S��Հ��K���լ�����*1dV�}�Z?�����)f�ǖ��e�����c΅��8�w�__���Y�Z;�pB:5a�bU�2�s�K��D�^=�!0I���]�_Uj��
�m�Z�~)��(v �e�v̫���9u�a�J��-�Cv2h��@\�.8B<$|S�$Gy|k;��i�� )5�:�ל�����Ba��+�@e>��ܱ.@��_QJ*v�
;O�5Ҷ���\�	�a��q�E�M���E�,��p����"�y�����5XI%A	��1�D���]��Ka-�����N�v@I|�:}�;��Xi�Q�t0���+���mʹ����c�FYN��_(7��"�n6���V���N�6�8�����F���L�?V�C}�#���f�P�IC�)���T��M��n�Va��;]V�ߣ8v�:����#�ݧ�Zyg9���eީnҟ� b}\"���?Y,i�X�s7���6G��lJ��Wj�
��+Fu�k��zs���o�fa)�j��'�m��%7<sjmsE�P2�o���AI�Lm��_���~��l�����ב�5mh�v�Z|5iՔ��v�d��\P�����EA�@�&��sG���A#2��ESȓ+��`�M����E8[�|��F�X)L�G���C|����
Q��Sc�y��ߩ�Z3������!fU����.�9e$��F���Cn$���q-<�������r�Z�o`bj�J�<���"�������CV?ˮ�R
��{*��(�r"�|3�yw�m|z�c�`C�[��ul(i�]����X]�q45��T��~!�� �?��{��zѫ�&P�>l�px�����݃��^<�L�'��"r�I&c�ő��vM��9�@֨eơԦ8�?���b_l� ևc)�<���
'�ƧW��g�{���E��ık��� ��I��2�!Deݑ!������j����K��J%X\��]�Q��5���'05�^���C���+\V
�c�}�4[�����cW�t�`oɀ���IDO��E�L���ힰz}h���(1����\i���Q���A+ ���ĦQ]hI����;���#E��}4,=���m�8_'�B�</%~ꁷ85�,Y�T�M�v}���R�A��a(נ%����T���*z03y��GTG��A@�龨��4]��I�^.�uRo��J��T��������a^k7��
�wgR�T�j�ma�/'P�	�v��q�8��u%�$)*q�׶x>)�]^n�B�ͼ����c��+2���jKj�(8#>�� ���D��%�&�K4H�Mr�Y6� ��0=m�[~�mR�2��Ҝ����+i��ǂ>��z�Bs"x$Jxʹ'9�m[#��EJ�U�i�==KǮIh7�J�.��3!�U�m���1�z�d��.�sK��p����Fu&��4ލ�����t�W3�}�|�i-�{����5����c��H'��~�J�6d-8�#� ��Ivdoӯm���y�@�����W�F�n=�n))|v��yS��xL����}�|�}��_�<(��K(I��h�w����%>�F�	w�6/�f��`�@�є I]pk�[9�͑���7�G�d��~j�NbTɊ�d4���3��xk��?T�4�8^/�[�/�yk�X�b����/���/�W>��K�X�� �6��:>
�8_�����}
w����w����?�n��Ť����(����5��>�z}��mV���(0V�-��EX���y�]>�l�7��QBx���׃���O�f� =�_4�*G�)\d�ʡ���%.��򌒪��l�\!v�W��[8���!K_`e��]Cע!p�O�C���
�ڂ��I����m;�z�	Nr��X1J���X	�F��x�)���	&_X���I����~U6:Q���@�O����Y�k�������T�䶾��<���LW�b&�֧��;%}�ޞ�|n�Nap,��\,��~qkj	�;������#��k�f���>$J6��%�\L0���,=�o��%�����\�h\V� +�l�-j'�����J���U��""Kʶ�u��C�Er�G�%�:����G~�E�EAS��WLM���'h}dԯ�#N�A~X%�U����=�`T�iTj֯�s9��Ә�GĹPBa�W勄h�6gu��U�g���.��1qzZ��׊Ab����GXH��#^�q�+��g�}	(yꣀ��'��IuH]l�<f���r�A8;F}���+��x��g��eGo/� ��e�L�Y�ae��ǭ��qI�tp�l�_���fi�� ��q�Od��u2W&:�7\Q��4_m?���?�KPA'��'(]%�wKĭek�[`�f�w�7�wp���"l���A�t�!v3�Z�~(n&W�wК��*��\���Y6D	R��u�ב`x�
�����߸�\3�۷y� 6�M�V7���Au6��@ӷJ�cXű�7�%W� n9��O�L���)7��	��,>��қf�%�/\���\b�c;�څ|.M�D���x�CJ�`����|2��	���LO@��ad2�=#��R{+İ��iRh��&�i���->L�`�����-0
�@Ʋ�u.w�9��Dq�[Q<���3�EG����y�����D�xSv���m[��ª�D���P�g���a������C�i�f:�h�"�L���-����rjA�PۘG	I�l��ɨ-���j7���^uWS]ߔ�-?��Ŝo>GI�\�Z�(;_�1��$t��fo���g}]��
�'�&U���C`%��\�ɷ��b�S(��T��[���ұ�V4���N�ʢ�I����P3SӲ�9l:A���j� H~P����y$Sƣ�$�;�~��`W0�n|�t��qw8������D�wA�~�&X�O�ԉ&�W5hw>����f=�\D+N��X¹�nbf�ܱ��M�k�p��_[�a����9�� t�mX\�V�������]a\3�=X%h�S�*bd��F�|K��gRyA����&R{M���� �ӂ\[���\��0;��_IP�6ܫ������;�v�=�b�0��m�Ӫ��q&f���În<�|��W{�lN����'ϼ�����l��D��`]�"4f�ķ���'�1$�L�8ŖD!=�p��g�%��QS�ڐ�� Y�Ѱ%����9M�y0�I������x{kҚ+Dr4�]>��~���ۈR9y�}�t'f��j�[b���0AD6�z6�2���k����#�X�<����c��a�|\�����:c�k*�|�Q�pv�_�x��]�>i���r�/c"}2v�ݔ�yFS�8��8D9Y��%���]4�P,-����"Ҿ�;䧚P� ����v���~"��e��(�.��rN���SAyLY�߫� �2�Ht	'��W�PCZ+��]E6+��#7��A��6P�8�Ys���Mݗ���_�aL��*��5��6�iͫ��|�����F�e߳���!y�� n���b=��H/y������4\+!9�M�P�����u��?�^K����<21��C�)�Y�f���hrX"3�5U��;��o�(X4�~� ��m^~����6��A���)�#载�qI�v���C�i�ul�iESէ����9�`s����ȸe��2��}Mv[���F�?vԬd�˭�f���i*���
���#N�d��'pk��KȑV���/�.�ph�������8$������*��C�bU��d{WX�V��mNL ��@�>09����A`a��Ԅ���O|F�uш�S�J.K����2}�<|�6���h3t��ɱw�V�4��{-�6���V��Q��Jb���Ӕ?yrd$���R��gIS_f�vzن$@?cT��a'�㽢g���neE�8$�
``��3����L2���LpN���,'奷��F����LuX[�#�^�;���uR��Ŭ����LC��Ο.�����F���L��s�8#�����uR��K~%^�4e �	�@؃�d�����^M������I2Ŧ����w�KgET�!�A���J�����ڨC:T%;�.u�9�? X��|u<8k�)�@��"�ϒ����6����)�r|~X��j�-�ɸ5.[@�����d=�Z p�@\"��xNiK�N�@"#B]P2Fs����P�1E�������3�}�p?d��5�A��J��d'"���U�C[l�s�/Ǯ��w8�ǆ�d��e����F�ih��/v4�"[G����jkv�v�p8WP��U���ͯcr4E�
�h��ǲ��5� ���Y�"J8lꠇH��t\�TT�ڿ�W}���n�͟5�7�+f\߄�cg^��A�`��|����b��������yǫ��qt`���_���q�g~�/*o�, �J��6R� �pm����������[mSf³f�������`\v׏�ڪ�F�>�����:ʣ�n�����@��b(@�"���sp:�R5V��{E�i|`Pf���Q5<f�&���
���n�{�_�&�+A� #x�b2%2��.�6v�m�����'��]:�:��D�!����{\����+J����"��1�ѳ��Nu�w��@�;�=w�y��eI0��n���?G0�8Vh,�g��}=OͦNu}i�+�Ȃ�;��Bl8�jǯhf����3@�ɩ	�D�cy���D�����e��
�]���Ç���h~�H��8�䢇���d�a��������B[�<qZg�p<^�-c�w���F�8��0�����;Bt����:�H���[��3���@i�a�S&�"��G+Z�j%���e��CD�~,�w�(�w=��e�g
�U��o�{C�Lsʈ5'��(�.���)�"[�?!d�z�S=�[=,#�י� ����H���VPE	pi���㗢�/{R]� �d~i~Of�ȥ��b.�d��Y��H�8YK)X������q0��8Ҏ:�l]�#n���,�,#&=1]�a�0��a��R˃g����Ғ�ṽ�EQFb��ªu-2o'�Yl+S�.�8v\	<ܵg4�%�<f��Sk
���4��58+��j\�����p��W��T�	s�˿�ݵ�� 5?�֜?���CXK����g�0��+�o�)y���~�@.zf�j��U�JPQ�&UD�8��lg[9�ww�ZlGYw�P�!�T �F-pY��<��sX��^�����\5YD��2��G.�����!��B	дb�Mڞ��F��'����DY�����E̓XJ��{��NȺ9Q��3�'��D)�>�}����~��ai���8��Q�(e s1(KsԮ	$(xx�������E�x��������T�?Y�Be��#���g�jQ��jvy�g z>tV^V\��b(D]Yܷ�1����I��1JTu��ԣ�_�C~�a�Ama3`e�n*��f���≌#�O��0.��u)��y^��u����O�Ҙ�����d�l��-C	F�`r�!� ��`�2�é�j���[ <l�����HRf@ӿL3��N�c"Z}�~.Zh�	�Me�:�'%��tC��|dW����Z�6��C�L�X9Ԅ)�I^տ�]��3.j���G|{(_x���A�P��_n&�+[�pl��qNR��h�Î�Ҩ��u�=�-�61eZj��Ӷt"7(��$�RQ�"���4�kp�c\�T�/&�q=��DbNAF��M�[0VԈa�S]��<�Y�2۾�|J0��������R�)%�H]���qQp�t�ѻ��1zX��A�'�t�&?�/x����N(+2��G��
$)�����+�DrN�h��'#�;������X)���eQD
�΅>Yf��{:CH���3�ME����C�����g�k �a���eao|��M�'��S�������d��zV��J:�a�V��B{yk�E@<*nZw;��s\l<2:����+]�xH�/�����j��}v�S�M�T:��l���BL�-O%����2�"1z ��#l�E!�V��g�&��˗V@��`{���1�ޥ="�2w����vٚ��r��R"+B+p���w�j�#�T%E�����X����qB����6M�Hh��G�;4�&y|T�����r:��߹�[7�r�DFNʴ��b".Y�nEyM�h�qN���:4j���v�t4K�d�q��q��K�Ie�>���p~�+�O6��΂	
��͐����@����o��S"�M������-�L�PܘX'�����b�%H�H-�)Qn�8l2Nn�+����F%ŧO��:B���4ɕ�\���tr�!��m~I��ږ�E4�54pb?ÂA�Q�5Ŏ��`�m^gj[:�'��7荍�]/DO�<"��ٝ�sW�
]�X.��H}?r���������>^�U����7��B���7�#��t��o	�P�z���:C�[��OƝ/@��*�,�ߏ��"6��S϶�S���O�BN���:�ǅT?�(���+��q��LK
���������=r�V�%k�-�iFeb�c��iH�ߢ�fc��ۇWb�Z��� 7#�Bv��%�X��,��AJ��g��\ �o�[F^�H������,�zKv��X�y��Z9N��x�vf�<D�5�,}��J
��#��ݖ� n�i^7U��jVG���k�$.򁯑��<񋀪�\ś�(� ��<������/��L�m�6��$�
q/���"��Q��`��M5Ԏ��/%�j^� /sd�d�g�w�fM��gZ��@���+V�������(�л�aX����P���8>�L�|o`Q)��L'z�u�b�Oi%�`���R�<�g'7���j��,_0��FCR�Ng����!�>������js�oh����;͊˩�yK,;�� �(�}��W�&Z��|WX�x	x;�}Tο/�x�9e*��#��i���2wܽ=���� �)�;Ɇ$������9�Sc���?��@,�.�(ج$�F��	Ӈ�q'}��#!<ODޓ¾�i"��%|?�k�*u�b������N��2�����j��a8櫅��b��i�^��I���WUĻ����,��A��^� _L�^�j���k����g	铬�������yu�Қ)�YO����OuO,�?�nS� ��ی�
Z�j��G�.���6NJ8�8���$}`���=>�^��
�ZX_Ss�|�--�n���R	�S/{�:��F�r��(��c�����ҳм S�B=|�����ja���1eKG��\0��������~�}��;`jT����y7Vp!�@���V�����4��Pa���2�sV�.ɔF�d����=f)��s�=���=�L�����48�s��Z� E�DgВR�,�t�,���	?�(I�|�b�,Dt����
E����R�/�����0�!�j#��͘��B�] 	��A9���:beJ�"|�5�-�aC��������޶dF��>��5�(`؛������5@mp��u�t@QL���f���u;�C>�S���E{ex1��Z�-�֟���<(���M�{[�Lu�d��.���7A�T�b�������P��CRs�-l�i�u�9c�_� ��K�T�/H�e�h���yl�)N�<��R�-��z���
~�#��d����L�Q�W����;4������7�d(2�d
~{�ϓ�Dj�ZJ*gb�<�A��9�E>�� �^B��_�#0d����	���sp����:��GhF�-Aa��r��%�t�v�431ɴ��O�Wϊo[Z0;�L��J��Ohr�k��ܥ�Bi�b�T�ޫD����g8г����s� y���d�$�񍯘?Og:�R�v$Vt�Z�r��b����Y�n.��p<0Y��ʐ��!����ˋ�_a*��-��,�(�[��)DGI�`��E������X*�ھ���y�u�z��.�QYۭԯbAW!I���<6���#P�l�`�� A@z��,��(�7��r'7_�R��N&��p#"���oO��d���-V��ko(�.|Кj�5�wO`:h����߈3D�Sp*A��6+�#bsv���*	/������]�#���8�}sD�	�H9Ւ�p�gUwM�pO��z��M�g}�R%�N�twKp��c{M1q�M�
��w�5:�I�:7���j	���dc�6q�7��%�	�,�h�`����V;N����4�_Q�͠��i7g�Ƥ�/�j�.���*����@�ꈣ���"�R��$����Ym��˗��,	�t�6�
�v>T���ri@+��8y9y�Ǖ�ud���s20��Y?_�0땖�,�-'Ӧ��;9���%��N��m>�'��p�!k�8*�0���o)�@:zj���z�zʢu��/���ɩOɣ!�?s���F��uv�Z.LZ@g�au�u�8�4�.�a�������Цf�2��V�3[� ���~��{N}:m���T��Q|O�Ge<�G�a�F�O4��r!�T	�2���;nӘ�̆�J# z�2��K�����-�Qd��;�Ppn��s%Ʃ�U>r��!��L������0]c!?���:#J��e	(�5}���2jkM����JND%çI�y���}F�'�p�������<;��v1��$����ЬϏ�8NT�r��H���`7�����$)6|b8���Uz���)YD"X_��͏F8-�?{+����VH��ڮe����m|�"!��z�c>�)�/x^�t��4�;s�׺�+C@���n���]�#̎C�Q�E�g��$�����+��X;{���].�l�o�b��:��-�3i3tL�����w�&U$9E����>;�p'��+;�sYY���{j�P��R��7
G��Z'/J�ˊ�o���qdϧBԠjb|����JPv7���36s]Z>U<&�x�j��}�>3Z��zx!{N�|��U��c_�O��C�K\��vk�O�cT���"��y!<k�5 a^b�����~�M�O
�ӵ����f)c;_�<��衋J$6�.e��r̞Ǣ<��j�����
���xӎ����F�8��B�zC<惷g�#�]r�M⇢�2�3�!H3^��7��k	cȀ��_�Wf�;�q��U���º-��[������E����p�5IL,����.�H�Ϙ�RVbj0�r�	c�Pbzۦ�����
���w���=lA/q���7t(���=�9FP��/'�"��y�^��Ծ{>>F��Z(d��y"�]�rs�Yڭヤk<��!�)��)&�QpC%~5l瓰��:R���(x��UC��uM�#31����4�V!W?�S~̏$�R�x�Gd�����@#��,h'i��:-�Pxr��
3�x�k2x���a�x��Pڻ�_�^5�`�{&��-�	��t���j�ಘ�T�z?�Pl�$�����������=$�; �w��H�c%�!V�|Ԍ�2��	��4lOߧ����T ��@"޽�����~c_���=`E�����|X��_��k�D=�`�n�3SKN�맬3�lѨ2�����Ba<tG���bi�8��z�䶐+�2���N�kWga}u]��T1���C$N�VH�h�������N�����|��G�Q��MQH,�������Ko}�&�t�Y�����q�%0J}i 8b-��^�nU���8�VGf���*/�/�=(�<�jq�"LAۈRVg����H.����FQ�c�0�͇7hJ���C!.�l�U�O_�Ķ�7��	�ߓ�)Y�_[_"F涏��Z�<)朤�9gp���ݒ�S7����VZNׄ�������j96�����q�|L}e���{�U(X�3�Ƚ� ~�O�0�~�*X���̧gT��c����3s�!� %m��Z���ui<T?�RٲR�2A4OXP��J�TY��}SQZ�����B>,@���,a{�a�Qᜪf2JE��x+Nom��M���^_��A�y�N�<��?�aN*��L�H���%�UyRy�������3K�0Z4Ʋ#��ZS��
w(8���h~��!�%�WC��)P�<?�%?���p^�*����\ږ�����B7�r��9�	�h~h%�	���n��GoB8�̶�\k*P���M��.g���M&8��塕�A�YEeR�� q5���$b��!]y�M�Q�[g8��
�"���Bc���A����ƃYf4��P�.�vTb,����=U��۴M\Zl�z�ѓٵL�Y����%8�������V	�
�w���`�=�] �Tٓ�xT��VD]��8����+A��*�/(����,�̓�_d=�eB�t�eR�:O(��=p�'K������a�`�f����2^K�j���ZM:�͌��$S��ՌoE!R¬m���Iz�������Rr��̟�Ec�MƚM4/J�C�����/�~(B��܀*I����Sx<�V㻽�!�����P4�I/��W���Ǧ��	I`}o�?FJ���&���8Py��
�6��{����q��p�n�j��҇G1��C�5�<�ܪ�K� *7!�ɛ>\1��ޔ4�Q���{^�ԕ^�ʼ��xZ�Ӈ�8kZ��neh�P$��!�98�`<�X���_�VR��x`-�����/2��P2����cR�_�p�s�J�=��yKpM�h�
��{�n��/ *�SV����D
�@��ҿ���l&�V�n+�zb�<�?��O�;ۋM�)ڎF�����od�lo���:�ծ�H	�ɍɆnv���f6^�#,$Tz�
q'�XE[ݱ��o%Az�`�	Z�O���Ҭ��K򺈷�G�5Q4���B�W�">�[�'/.:����pJ2/�������"
���l���o��OV�a��do�Y����^��z?����մ?2ش�@��C����P��1�rC�dRW�X�Ia�Ei�ӌ��� ��]��6#$Zv�Q��	O8�i�b��w�~ʖ-�a���^i�����N�K�e�܈{:ecޡa�[#9W��ׅ�n�S*����0�H��Տ�0��-���&¨�s)q�;婉�K,��<��)B8YՐ3	�d���^p��1���;�����+`=��W�
00�}�;��w�����F�i0����8xN�R�
OX(���	%Sp$�0p
�㌁�Jۑ�)�H�=�Ų�i�2���{�3�ٞw��Q�u�O�-�xmGF���p�^
c�}��J	�g�h�=7��UDR���X�Dt'�u�~C�f�����N�X����Q��?�'���,������X��@��� Ok\v�:#��;k�oޗ
�7cF���v;>jG��iU�@��g�;�7zxF��qBU�π"�m|ư�5wۋ�/����}����N�ZPnj�
�x|6�D����3n2�!�0�SO�-���C%�f�R�
�D?��r��C�҆o����4<�缢 �#v$��Ѐ�{���a�悱EF,t���d$�p��.?1�m�l<��1H��E�뢈�+����d�?��у�\n���������ꕥ]�Wb��+�^ي��y	,w�|_f��3�]�Rç���?�ȋ��$sԘ��&�Iφ�*�]��n�p\:�qi�zn�|M�t������p�>��U2�	������r�(ӷ�O0��0�LX}
�xF�A��t���"�A��g����K�4��W�IZ�;��󍨀0@���=!_�_��0~}Kͽy��� �CfA�߳BK�����:8b�'�C�#I������힬	������qfif���&��՚@f`���~����Jo:��6dA���7�}8jp��/<�µr���V�{��U�|ˈӒJ� ��l��,텙og�KJ�Q�i��	�H�#;�[4�nlu��2��	��g��r�/]�l�PâE��K�	�F]�ts�c3@i��޺�s@I�g-�(ꮴ\�����*��D�����ǡ��x^j�x�i�5��9_�R�]e'�Y���?:���5$�w3�d���nsr����$H~r�(����ж��W �i?���л0���m��hq~с��j^���	S�Iy}g���1CI}��h��7�p5�=/�b�-��'4O,��J�&��Ν:���M��`L�$�׋�h��'�J������{���膸�T  �z�D�2r7'�.����-4C�cjھz������G-[��Y�OUP@�+���/����gY!���h�B����7���{�Aջ_i���W^O�|��7!���Nx�o�M�UA4��f�X9@M�˔�D�p������[�$�:.��\��b8�x�c�E-�w��d/��0�t��JK]�B�fE&`����<��{}L�k�����>|��ͷ#hE�i��l�Ѻ�N��P�@t�4���ݾ�e7Q"�M#`��EL����j��8�4��WHS��ַ�:�Hp�� ܜ�x�����s	�I�NɵFQ�e�ӌ�"�0ԡ�4���b�Z��(�F$Iq��,	�O�dQ}	�&ghy���#C�`P$ME!F)Ϳ}���1o��s���9Q*K��I����m�[�v��G	&�cj��b�n�:��=�{6?9�6��@�(δ�J����Y��`����]�����"��T�L1�*v�mpF�����A9ʥ�3&�81.b��*���vHb��qٴ}=Xb����(5��]��	��UXv�.yp���!�Q=ӶӴ4�˓s�����Dl$���d�g�U�}$|��_�e�h��t�O�b]�DXeFю%�P�H3�k�>/Yp��˸��_yL^G����q阮mP������ -�k�Ș�5[؇H%����?�Qn��q�BZ�hj���n��W\_~�A&j���z;��h�)���g�kloSպ��K�U����/Y�,UBשR7����q��od�K��vr�Z�u#�_�Vp�p@�c� ��F�R�i�fH�.i����Q�Ғ�x���ܦw>d嬴�3�믜�Q3oz�o���kb�\"�B��a]9�Ѯ�A>������=��X���}P�5��v�O5u�P��-3i����>f?�߽�Qأv�&��!��ӬN�5q�:�����5���Df�͂4Eњ/��z�:��f�W�>��^T/�Ă��(%n3�]t����2r�X�X�0����\�3���{y��z��d���獎k[��3L2�(<�v��?�)��(���qS����nt���_�;��k��	�9���v3�ߏ�N}����處t�m�bk(?�1]�׵��xEy����z~-FLl�nj3̩��Ѱ�Ar]���'�L��Ի��Y��C���5�c�F��(Q)��k0���E�g���R2���x��a�ہ��	��$�OV~���C�틈�:�,��N�+�ع�tC��I[5�����N�v76/�ȱۘ�����wR��A��ό�e��!+́�ku+�$�V�dy��zrݏ\t������쯇C=�V������j�f;��j���媴�N�]5�P�T��F�Y�O��e�3쵙��m�+�~����"/S�E=�,4f�� ��,#��fn�$qm:dKq�����L�*��:/�-|υ��K��Kj�/3�Q�x&���З�:&Vr�00)��{*D��;�`�%�y�ms�h�2y�Û'���c7f
�L�eY0�;�W/���&�Ǌ���1ڦ��w�LAәH�Ɩ7��9�9n��VD�[��:�U_����A��h��]�na���� G���h+ɓ�i8�[ӝy	�3?Q@���l�8aGC�Y�_���W~��^�t\R�T�H�AL����j+(n����4�|R �s�_Q���kxV}�K��X8'��d��4/Ě{K�9�X]�O^.e�_˧�3�����|D	�NOy��\m�dj�W|��hzV4>�`6�|����r�J �R���A�zo�.�vkq�;c�tW'T�В�|I��5��?�5N7I����4��m��<�Aʹ@�qJa<����/������Oja� 6-�qK�^
�,̨`�'Xa�+�&�CP2�;���e�A�|�Yy���jg#��b�8����~A�	���t+�8�s�X�Fc6UV��L�R�B
o��r
�p�P�ن!ҝ">�W����s~q�����0t�,!'
�ҕ!�ct� �9�K$݇����~�3�@iT�I,@y�������%o��)2�Mf��ܤ�BYp�����C�Al�	1*/��ʸ$�|�N�H�{��L)��x� *���KB��9;���$�j�De�M�:�ʍ��\�8Ki� u����U޳�	Q�Āk��A�V�ع�9�^��D:H��=��Ψ=�.�������|�����k�p�-��s3�%a��P/:+a�ZER���eӔ�%!O4+�Ei��cQ�rYs�CЁz���,^�?���Kԭ%y�WP#�	n2����f^O��L�MǆY�e�%^o|��N�3xt{������AW'����+-���(.!gi����7:�/Y�޾PE[_äɭ*4����̤zlB.?�d�|nk4=´+;q����Z�ľx�j"����K�a���~T[�xzC�ˬ�j���&ZN�߇,���1GM�����31�_�O���gp�MT�бPc3���ըC����՟)�˨�bG��E
c��޼�,G����k�;y����D[�]ǩwA���Z��>���s&p��E��vj��B��}N
�^̝G�3��!pzF?i�p�����A�0�ht�Y[ h��x�5`6��M�!�c^������F�u��5X+?�y��R�Q�u?�Y�֖SRF��̳�3/���Ao�4$�����F�P*���Z#e"�����*�+Ж2�� �{��,�F!Nٓ� E��FS�Bpe����R��#�[�M���׵���ae0^-���Vy��
��H.�~8��� Fea$�ʻ�9���Q��dd�uJ����G���e�r,o�|�-Tkǜ���M�gH�������dQ�ʋL.5k����e�p�d�
��^�bi�-�#�qߤ�y���D|��0S�U�b�6S 4yL��s�@��5�Q�"�#\J�N�l1>�O�����B�nvpU1��x�������X���Ӗf;+yk���%󠂋uH�Ë������!g=�Z���Op��M:#��z��9�wS��Ӿ���@�u�+i1WKEކa9���Kb���S_�+�a]���	 }��Xl��`�z~�hQj��P�vB�<���"�9]oT����ܗa�sةy�>���]-l'��v����i2�2ː�9C狲�cA�.
�㷫R��m;i�#��X:%��]j��mn� G�6nv�4忱�P���� ��0S
G�F6��e<~#l��s%��v��W�@8~!��!��J��u�5)8��_un*~ ׃Lh�����88�Ǯ��$ a�܅[r�m1�k�̈́jfP*��՝�2ƺ���w�寔�>�:�G�=C���G+����^h1EK���j�~�(7��%���Y6���{S���Zd&������R"Ĩ��<F������'Y���C��ty�Ɉ���t6J���-o*4�W�����:�k���pZ 6��p�|�3ح}R�*9�ʛ30�ٲ*ITx�ٸ��EN{A��3�⹢����$=s�[�HF�9��Z�x=�$)5��d�� c�y����wHl{��������N�2?������nB������$����ht%[F t���@Dm_�/#�"�/-~� /R�N�Q	���{�^ٞ���0�V���n6pd,�ɐ��	N�]����z�jcM���G�L���/�#s��'��t_i��V�gLEI6� @��K��-��(�*S囚�l��Cv�
�E{&�;ٱ����ٛ�!; �q��6��^�sPnN��|\C������H��5�1�`��@{[n��U<9	� 7��}�Pe���Q����o��O.x}�H��B�6�{ȕ�+Rr���ؐ�
 K�j��s�L�ue��.�f9?mٌ��Cw�Rj��a����`��2߃����s���={[��X�Egõ�q�$�/�76�RH��-�R���U�&��Xb�&��%~Щ�	�k-c��sH���8�V
S��@�C��n�'�� U��{!ҭ��F]���Ӕ@���r�h[1�mj�\�ӛ�Gű�M]f�k�
-I#L�ؖ��Eo-�"�ӫT¡�� �n�wʤ(�y ;6�y�4��{��N.� ��f��ut�|!��`ͺ��M�:�T^B���n'v8&����󯂁Ώ�i��}v(�X#~jg��h��fQeg+��;�%����ie#%Q�+�*�����$�s�zP�~�-QfC%�	}Xͼ2��f֓�5$��,ǻ���Z�� ��S��:6@pD]�./h�u���kX)a��zPu�~��
�:�������J���ŭ�	�&�O�#B��o�PO��lU������]WI䷼(�����ē�n2:F��Wi����v��%���bji���Dp11ۗ�Zg�u|`uAͣ��^1�(��^G=a��"� ^��6�f��*�R�h����94J
���
�u�ڙ$|��w0 ��S;^�����"���9���N;T�1�`��`AJ���{���1�kY�æ���MT����S�>��k�%�#4�X	^VO����U�m���{�6�EZR�&�=ܵ8|�J�4�¤"�`gs�ۣs%��{�4io����)�U>��2�f���^��KĪ]/%w�MH�o��7���t��W�F�cj峪5<�cթ�/B��աp(p8��ʏdqc���i�)�ɵm�'d��0L��`"!�+��Qŗ��3��+��`P����w�Kb����jQFۣ(],�-�eN���v2�h��Xk�u��/d1;�Q�5�風8�3���`�����Ubi���;J���y�MmL�V�uݡ.��rbp��Ol Z@�Fw�;#&1	��w���'�~�Qm4����Q)M�k��=~����`�%�"MZ��m{�Q��yϧ��6�D��T<�/w���u�I^�K���1q���ȣ�M����UT��4�Nd��� Oi���{�Y��Ю� 1�18�~���U��U����N)eHq	
�3bD�{��Ց&�t��c�ԗ�ӕH��#�W�M���Ԅm�y�و����D]Al�&�?	.`�K���쎽�p�<�Cc����}:�A��j���-�ː���.i�%���B�,�C�e9L�~Kun:8�ˏ����*����]f�,g�ɜ��i�����I?��F`_@�[�Vm�k��8�#ؔ>�@3vÝ�&{%�4	ۄ��b̋�%-�F�(M�����vCp���V�b�|���3A��#�M�._��!G�Hc���	UXaq��5�)&?�7io�%+3���5���)f�>�.arJ�-ϯ��@*�Ʉ�Fe���zlq��O�i�~��vywڥ���f�t��}���׾��q(*2ٮ�Iq�<��5Y<*'|k��]xoil�?݌��\ZQ�����L�U��R��a�},�ת���񦋼��AY���CѤg�[b�c13��� � �8�>`���՜V$ߪ��^���ȸl��N޾��<Y�ٶקP���s��rғrS�[���ohy�8��^"\7Ζl�C�3�6M	d�!�ݲ�D�����O������	��mk���uG�!��@�1^
#���8Q�����gy���k��������ZZ���h>'��+�9��Wa�����F��o�?�JJ���Ğ�*���w�
��X�̃�,Z�o�VJ�&�27�#��_�t��`�f�->4���׊=�0V������?�NjzH\ D�&�{�(�)��*����-��c�b���� ����pf=�c�d�Dm@���m�;��OP.�,����������|��c�i���`�6xz���>g������OHD���#{q�������O�z2�0��j��9i�k��RN"i��|lY}4X��# �|���Ogl�v�,��O=zn�%&8��8�.;�`�ڏ7�͹�z)�9&�1:@1�֘N,PQX{��n!�x�$ב�z�^�<�[6�Խ':�CL�Z�'��"��%i�{3&V҃ukE3��@�'��,|1 �=�#o�c/��`[���'yZ�[&�a�z��3rօc��`zΉ+�
~��$���WB���iY򛐞��:�xg�ң�� ��]�@YNx�U1�����n�r>Rۀ��MT��&2� WLA`���&�]#ܕ�oXO|���u��7�T�L��]#C���Kr���	^�p�`{s#�e�����ƍ���"���/��6��;��C��<;,+d�A��#$����I�ɡ�5��L@����鰺�	4��Ɂi������4�]�ٲ���c�Ŗ<JnUs;
�7�$Y'�7�	��l�Du���0��on =��;f���j�a.���X��ƻ)�1cg�k��� 鞌]�{�6��_4dւ�ZkH=�o�-y�R߆�]�Ihez���rl�ɟ0��}�}L5��M��Jl�^ ��x������J�S��:5�D��u��i���f�s�<8ŧi"�����m��c���3L���*�nN���X�G�-�I�Y�4�]�A�>�q��V���0wN$IН3�I���L-��ƹgbF���;o$�H��"�}5+����e}��r�)���"£-E���B=*ā�l,� ���A��:{؄͒��0i9�Z��g�KyZl����h�ۨK1�4ן1S)B2������;/��(���dlj���X�
M=˚Y$BO���1�Ԋ׏e�C5������ӫ-%x�鶗�!p��1�h�+�qP�VމvVB���'C|s���]B;��o㻩!�க�vx�����J�"�o��$7�y���ܪ�*H	Ø�4Y��>m9T�(�(b��Y���ٶ��&�G2�Ti���6']�㌋'t�V����Y���޸|�oJ��r��EH2UbC3Mj��|�`:��j�T�T��A-f�y�5�:G����Sִx^��b��(�H�M<�s�PJ����a�K(�Y�¿�F�	���)=X�8��=�fa���[Fh/fl�]��&B�|�)q��v_�6��M��bk��H�u ҃��j��O }o@
�:Ԝl�;B'���oeď�ࢢ�1$�=�׍6��g?���=��lYM��:@��MnPC����,$�r%\x.���`���HZ�Л�N����u�I6�,⬷�htF��g�ICV��؂0W,������+K!,y��Uc����~g��LWU����N_�3U���H"C=8��@�3��K:
��F6&qռ`@�t�!#����H``��#��H�ꃩhPا��^��s��r2���&bP����մ�ҝ��Ů6A���בdV._��MH�[�XYOs���T�I��U���<�Dꁣ@��U�	2�3)a��, G�RI�
�"�����ki����ߛ-���/!������K	�T�f҄��+%]"��=3���]�������ߩT�v@�{��k^��$@�����)���M�x��5*8���i�ǠmWO�)��B�ۚ�[S�=��|?�7�P�N��������Bi����ev>�Ҵ����KA�V[U��JB@k �̀��s\R�i���5�^�ƿ���P�s,��������j�67r�R,Bx��>����0�8풆�.�����	�AJ�q;� �G>k��y��E�7h�Ȣ�Xq�m_��%����3�K�^H��&�M��r@�3��͇B��`���V*�)ڥቬ���d����D�����w{"K���q�R���,�3�y��vB��w���f޵�^fhɔ� `�-����ǄĘ��ĕ��8�s��'o@����O�4u�z�o��H�^��SH7��,A@���4��u�O
A�e�b.�pX���^��Р��o����a��o;����:����8{6K;!���F�+H�!K������o������.ZQ��hbY�*��1<��"�	��L8��ծ���gk=��7rCx�Q^dm��ח��N�����7}�>��*D�����$l��C��x�f���{�ޞN;�b��[]�y9{#a���aV�n�=��`:�h-�4)d�
w�L"�Pqg�y���lZx�ک������fR_M����RohJ-�:��)��
�}�s�� ������G��������똁<�'|�FJF7��O�YcLA�a\�b���f�:���?9��R6hv�g����_�����M���ժț*��sc|���?�N�q��T<T���/��Fy�f�?�`bӡЭڲ����W�zN�Eک��)�)���Ce�9�� �AY�@�~R|.J�.���w<��A��͏�����K�xT�[��S�����I�Fހ��+0�~��e���g��5Hʔձ�O�a�g�#�|��5�3S���e�V���^NO`3�5v(��a5�y��8F�Oz��.i���b_n�1��ߊ8��x,4��KƏ��k9�3�̑p|��V��J�^�i��6⹃d5��r�'r�d�Z1GzŌ=©�S�gv%޴�5o4���R��[4��8i�aN��ᚑ��[�Cz�0�VH���	�;��������ʴ�A��YW_G�v�MEn���r�-��b�Vј�ߪ��Qlij+J�����:/s��οǩ�((������g��,4�ǈ4}0��6���`�S��r�ĵep�o8j��*kFP�؜��Y�=��焀ɢ�g���Qt��!yM�@7�B����[�)�F
c;��Z*z�DmM�SG��Ϧyu�N
S�
�p���_����x�<pH�������+B!���3!�sw�&�S��/�}ğ��Vx�p�7z�Ґ-�3�q[���@aP���4E'Y�e)>�Vc����!im������0�������QI�t���'�G�I�������|���t9��8å���dƳ�A��&�MΩ�l�[s���~��*
�2�v�͌��O$)�/\�t�<�����X ��ݺ6p�s�Wb���7"�\�ۦ;�[�����ǟ/�9n2��|���!���Yڿq<��:�������E}��/n`C�O`UڲC�V��6��	}�h-��AP���8�?k�}$�9��Mw2����xS8(϶�!&�@�%8���[b`�&ބ=���1�ۑ��ެ���lti���5�|wQ�
E-�T�],����)� ���y��A�2�*��O2Ҟ��	�_��P��5��.Pq'�(�$/�O�>"�A�;<O�μߟH�e���9Lv�W��sr]��33=�/�_d�2���>��z�z�g:8�H]Yrn���E�X��� 9wXD
�?j�7.�&_j��]�82MK�Ɯ�&8` ��)�l>�y%Fz=@ҏ>��a�m&��<�S�Ď�j��<�����+����a�{��!��99�y�>a\�{�w���-H��]��6��i����L����Sǵhx���iߕ��&���F�8�S��B�k`3PK�Z���~D�����.(=�/�ie�Ȯ%��.�P��c#�L���Qv<G�Ƭ�ޚ6���FZa�\�.k+w{���j�G�N�i:^%LG�X���n�uh�J����f~�}~�Kٕ��U������P�z�C�\ʼ9���0B/k�,�X�?����SHAt5q�,KI�6h��;�D��0�_8�x0ٞ����E3>ǒ�B�_���5ؼ!]N�*'P�w�#]�y�4S�
""Pp2�|~*TU�N5:}�B	Jn��sތa��N�H�(W��w��XUK�n4O�ʐ )��n�~+{\fQ���#�=�:Z���{��?_ٌ���5ê�RŎ�؉�Ȓ=�ި-�W|�S��o�Q�p
ϐY�U����.���';Mֿ�,9��#���}9�u�Wˍ�S�	��rݤ�i揫�J��g<��[N��$�9��f�q�!��$;S�GT$�P֒Є�k$qF�Z��f�'&�4��#�؄��E���[i�W]�ޘMO Z���U�зF�8�P$���86�Ҋ>%������������G�bu��d�&�*4���쨹ܧbX�N~���y��'�p_�t5Gݑ;.��f-�.\� �|���Q�O���Ű=�X1�4nf�D� �?x	aZ�#�\�K�ۃb�1F���#�Ru��Q��ŏQK�?�4��WT�~��҂��Ё2�6A ּ�e_8y��P���O���|�����v�z`V:>d�Y
�������,�����x`��2D��l�6�hK������8�h�־qα�]u$E����#}ȹ�C-Qe~��wON����*-�-�˵,*)��ԵYъ�>� �O*�ڬ
�E�i��Z3�I�I0l��H!6��I�����Yd�)���K	��#��t��!�ש�?��|����3�e�
�;�z,��E֞�.�Z�I�B{�/����D'Z��>+ʝX �f�/V��]+4#Fm��4�1�{)jn.
�]�vǓ~��u�/����8�GᩁupX7�	�}��R��$��2��P�ˤ��v}!�y0�TSh��i�A��h�i���뿽��%U��|��*�m�;��M^��lD'X�߅�
r���N��i�I��4�� ͻ�p�{�d	����u�&CJ.�S3p-�k�Ҡ����녫j|	?��x�����	ih����6KsE?�(���P�x���߶�_�ut�cق�Dq�^ýժ�$fE�4�!D��␷�����X�K]�z�L�q���R�N�fC����b�|�c�Ql!a�`z�!p��Ώ�̥�9CD���{��1q3��zGq���(ڃ���X�4��!���
�[�Y~<��<�	W���w�<�e��b��<��7[�&f0uZ!��Z �5��[8ҧ����L��w~3s�5t^VE�Y!d���F�:M�_����B!� ����_�Q�<c�/�D|�}���O�����L�������y:зq�1�|�y_	O�X� �	�K�cR�B/�Pf�o�O�b�	>�� %pJ�@ഋ��n����׋7Od���[�>ay���'���~u�֭���`����X�L�^
cd]#��l�n9�ƪd�mV۸�8r$O�&T�|#8��ⴾɌ˄�D+9�R}J��#�O�
���`�^b�t0Pi�,:�8��oi A�E퀡,[B\���[=�MrG9ʌm�~/�]\m-tǷn��;�G|S�mb���pF��D���&L>��?�%S󬮚��J����a:� ��y1�IsJ� h�0-M�G�g�����P�0�VXe��n�����C����GD��������sCQ��w=�uG�t�o�y�@L�Z�'~nƛ�_i�՚5�N�̏�lg�L�����"� l��=wF@���O�>1n���	��b(�_�����*6G4Rk�� ~���^䤮��Q�m�Eo��T��ѨP��闯��~�m$ô�8��X��F�=Ia��2%y>hJ���ٜ�H�V�TMĩe�ԁ��)�Y�#�T2o���*3��QZU�>��rgи
�\m�<Ƭ�G��&�%� ��+�Ò���z���z�k���H�Tr��������\��W����`�Z�Q�P";��-����9���n�+~l����uF�6b�i�e�vy�OMS�G�l����:�(�ldW����!3�d��k¦��¯]�,�~�1��Ȇ̢��p؞�k���]�Vw+![0��aL�Z;apN��j>UsۙM;���/���	�T/�K�EN�&�߳�Ь����S�����@��Vi��IygG�F�����M�<渷cQ͐vwl�[��V+$fGa��o*{�\�<�g.�-s6q��F��C�q�*1|��󛤔�rH�է��d�$S6ݮ��h5c�F� <�ڎ�d�_�@�O��������������K���)����х"i���M޴���v�-�&]8�[�nYE��"��_Ϛ.�l��Yu:��nM���"vY����v��7Yj��^f��2>�'�^����B)BK&d<b�.�Q���S(�s��o^�?��� ��_8d�Y=�U��!���.��$Z.z�I87G�ʈLpT��3��">Z�I�.��f&�@����u,�ON�YG^|��;hJ#������e���ۿj3�C���2*͌|-�s���Y�@�7��PP�^�=���D�*$�l}�X�
�P�����4�j���ɤv�*��u�tpr\y���.�>� �?VY{�TR�7J�&:�3M���e�2T�C��{��:�\�̙*�M.��R0j�CxiD�ń09?��B���4�Y�������;��z�ѹ�'ʌҘG�Y[P̹z��,N�ҟ�����
t�+�$ޚ.�Ox���0�{2Y�����u��^l���:�8d��4�aZd́��⤯ga�R���`
�W��<Jv�4}j.$�@|d�m��fG�W�c��V6,�~�X8�G��q����0ʊt�#��K{:�n8i:Iv�n. ���ˀ�`��<Hh`���^��عu�;��hȺ�j_2��ҟp�ŧH��뼕t.j��E6���O�T"f�x��5�����6��yhh���x7&�Ѷ�\֎=`�$c�O�U�\:&�*R�u��ɢ����/�{�[RӐ3{�`6���"�����q��(p��Ed�o���ٝ5�K���I�Ň:#�E�B��6u�務��Sb�LQ��~�����i�B��.]�lv1���iC�&��bam5.��57Dԡ�@?>.��ь�b	��-Ċ:X8���)�	��[����;��_w*VYgͭ�4-��&��F'�o
:�Uȗ��~3&�3�Ȟ7�̈́��t.���j
ϋ��N������Q��]P���dOG/���i�H�zk�[� ����"/`xDG�F;	��������Y���Y�K4Rq�^g�-A���>��;�ȆH Ơ�z�ˈ��p�\_Z�=�)Ix�M'������!�H�Uon"r̊��ژ�X����u0�����G\#��Ƀ�]0����@c�nC(2��r�����ԡ��`5�W��mMBM�XX��bl����/�I8c�7����o���J��eZ�WS�ǟ�nq~�&�6�J"fYP>��h��$A0Y����f�p-vc��hf��m�a�?^M��qʋ��e�w�*?���������Ө��>�f���l�z�uå6"ح���t-�������#Y} ����nu%;��u&�����OuE�&B9p(x΂1������3���$�Fqh֣���Ϩ!��u�.�r�n}�gh�@�P?�/��!����mmTԟ�0�jP��c��?��qQ0��×)lB��B��Bs���g�� #��c��VI�B��{☣��=t�夓��Đnm�8�H��6ti��mln��)�##M�6�G�����<�>�1\�L�`��<D�us�cdѽ�`��(�"yph<�HQu�!!=�KԴ�b	P7^�:�y��Xi�#SA�ɼuޒ�1���"(����c����t��SEaVPG��#8V�yUlM�_�<�E�6y����c>�6��T����~t�|/����
J�\<�E�0�޳͊�ސ�c�Kq)L;��hN������,������+����	w�T��/	p�����j��?��s]e�W2��f�W#icxãK0H'8�lI�6�܍�,S�	d�r�0��^�	ie�Y��,��m���{�xg�ˎ��ܱ�<�u�]��md.����%�rI�1�,&�I���F N�Lt�e��#b���ڳ7��~s�u5:��v�y����k�-����/=�ϡX��	!��*�UQ��B=�iH��4�d�lJ�K��(��lobOt�1��]Au/o�'K�Ne8���&�*9\���%��w�Vi.И]�^��?��fg	�8����L�����qi�tXm��Ȗ�·�����U�[�8���M�m9���I�����b��l��r�"�h�Q������u�`������.O%:�y2Ձ(�8��/���lp+g�S;��N��8�����Ȝ(߾ˌc��s,hΜwGwH����E�X(������Cp4rؾ���,�X�����g�H�qU�҆�{�jA��CW���R�Y��Yd�'ǅD�yo��7��V�$��P�	��/�7i5"ԕG�š�
?J� ���6;����v�5�A{��@��u�][1)�1�"��=��*�:D7x��� �߈+x��$k�;k�$ܢ���S���@pG�_kk������"����.��A3��*�Ũu1�ͻ�wBpK$�w�C]�2��1T{�3E��,Ѷ�`%w�JA��y0+��`x:?�V�l�P�o5t����l!�NC�K������eA ����,��j9j�)��@�i4���
���W�	-�簂x�oĊ��V���c����̂����pI���W%mT�3�7��^���ܒQ8��L~*���s�IB�K0��W���2�b�!���v�q���9x�a� �T�zb�V�v7�+�Y
� �	|�b��B�v�yլf�.#4{!��Y�M����m���������]V]Q����{h��{)X�*b�	�����Mrp�߬Ӛ,oPe��S�$�Êa
+>qS2~��)�8I�J9Q9�ַh��0��v��*{��ICӊ�e�Z���t�?���!P�U����� $�7������G���mpL'����vjj��m�0XO͸�_��C����!	![��8�WD�oj$�6 B�>C�L��/�[ǃ	P3��ܽRR3���3d�e�9(V�� T��+==b�v����k�߇k���Ȭ���0t��Ŗ���\�)����B�-[]B����F���F�{f�w�ǣ�0<MV�m$= �����!�$T�g�d��2��k� ��1�y�6�d4�E΁��,��>x��7v�ë0y+]��s���n���d�ۦh���E�nV�ُBN>�$�I���0��X72��\��
�0��F� 4����O�{d��<�B��2w�럚�O�!�q=��6_=I۝
�2�p��Dj�� ૥s���-*1�U~a:w�/�q�����h&"��H�cY�����-�u����φ�z�DQ� �a�������(SG�e�"9�/{}��F�0o�N�픜{�U?\$t�*'��Y�ϻ�Au�1��`&k_"ד��l�<�����}d�y' \�/p�3c��=A	��dF�C{p�S�(S'�q��S!�2{[1����~�=f�Yo�T�S�8�#E�3)	����q��̇���O������E�[=�B�S��]��8`@����5J�}q��7qd<���b���Na
)�3���Z�E0����9�Bj�
�	q�MMpxZ�s����"�u�J�#83��
��w�ltd�]��������M%YK�xX�L�2������/!2C�t�5�CG�����"{זV���|YI��-0+��Yd�)��Q�,2���k�-h^Pաet�	1o��? �I�G$���v� �8�@����ϙ�1���y��tf�.�,ؚ���c����c����R6�V�8Bx�..� �����S�pE�e(]��}�בp���Hq'>���(��+|}���x����W(Yv^J��1 7�琠���31ғ:��gjb����9񲏓O����Yo���Ŀ])���QxB��Bb0���	d _��d��ˑ|�'�֬jꔹ䢽鮿�]�P��p<�y��e
���ȰYg�)(X�4>�=��{tJi1����q�� ���f��qY(7qȩ/��n_�1�*��KY���L#�pΙ)O��0	���E�zh���|20����k���rE�*#޳�����ߥa�]���x21㌼)���2��d����Y�v;�����k�g;��k���>���W�.U��B�}Xz���v�i��vOd��+�٥҂gd�Ä�S�Kuo��\X" I�a�i]���Q�2`������Սz.��%��v�ˬ!1_R�ѐ^�����6��)�ȍ�(\Ւ�?�\�ʣ9��XMO�� C<_؆�f:����P�{C�e��j}��
%��yzI[���;��ٳ0- ������!S6J$���§�SC����a��K�].�im��x�UE����������>(�Z$���(�eH�=�
S�h�D3[��M�n��ns��%\��������]	�i���I�*�>�}�w�P�t<*�w�9>:�Fʚ�u��SGnq�2�QS�|�7�ڝc֕�Ep�8�2�������Sr(Vf��V���f�1���2j�� �E��g�A!1�/�3ϯ���ޮp�v>�a�1 �t�U��H��d���H��A
��ZL����Z��1�k�[�o_�-D�T�����<'MB%�X�O�t�f=2�Wٰw�B�h������8!4�>E�s�O����T&�����'�Q���֠rk.cdA��9>�w.� ԩ������W	 (F>k4!�?�}S�$����-A�M�n��I��+�"K�2��.�+
���=f���#���G;�����f������"��� ���OG���M��z˫퉿L��x��V�Q��n���XOj���x	�X+����x���@�W �&ݺ��A�!�H��n�����q�>����fA���Ag���5S�����D�F�.�ϙ�p��	$fr^D�aCO0�y�_����M3�^�˜-�ݢ���l�+4gmː��U�c������Q&a %UW�,�=��O� ���pb�*nC��ꠎs+�퀩ӝ!����>�j��(H*�y��;�D��֊�xF(:d�U^�A�>n���*{;�q+o�i�N]�O���^_�V�S�|�!5fB%nY��?��ڗE��%+Iǉ��ކ`?�՟�K�&1SkDS�0��ET���j��A�i�9ǎ�lA��=���)��F2�N�u0����C]��C�=Ap��;��E#�,��-�\@H��A�(@��y�wg��8̟ >6 1�� ��s� ����^:XF�i�b(���_�h�x8W�b)��y�.��&o>���U�!yI�����G�Q���XY�J<�X���$z����b�g]�p��Ѵ.���q���&�Ţ��|�z)}#��u�v���>	�M�2̢ӏ����Μ��a<sA���	d�4��c ���C%F�pk|�ı��8V���d����LQ� ���8����ԕuFSꏑ.������,t�ta�̷w��L1�[_�hc��\��p^���ύ����&�XXả5!)%lw�̾$��?t� Y<�q�lf�\5��2�̻/*��ނ6Xlu[��!�*�y���s�W�-oS�u9fk�̎�&��O�N]*�BLSX�Ӳ�T��Ҧ�2ln(Đ��d�#��� ��އ^>���z��Q��Q�%3�������l��Ę�� �t�1�~�Z�JW�EN�
��lf@��S�@���Mȹn��W�GNSҌ����%J�)1�l.?eۑs���sȳ�ہ5�?Z�,��·n�N��	���0�Ԡ�l��r��ݮ=�w�x(�:,S�F��V�)�w��9�;� t��O���H�)��\(p�㧸�b
�H�TW���g ��WA�� �׆	g{h�~4�#18k�*���{�I�"N������,_����}'���f�O�˝�-��d��3ʚ�P��k��5�����Xqԅh8�U~�8�O�BԼ.ydZ�J��\z��iXE�$Y�'4�9�"�
����Pn�����'}̻�Vo��$r��*2�	y���b��D���$iA�����Y�z<k�3���a��7��"�,����������}&\���I[`�Lh�Ǣ�O�2�N#`#Vqp��/�����(����>��߁/�t|Gn�����1J�f#��\-�u�/���x��ƛ61oP٩]8Bż���nW8sV�.O��;�	k�	�d�,\,1z�Ay�g���H�D�A6�M?:����"V-h6m�� ��ğ*�-���n���:L�"n�T����N���˯�ig��Bc�}n�3LϊH�ʓ.�Tx�.p';o��r��)����Cd�`�d��)��|�h�b�������)��iUt�2O��R_s�u8�� -[;���,�lI��ΟIgγA�ő��.Juq$�o/z'�&#l�ײ$���7���#�h��%�}�f�H���d�ٌ\HD�2�[�II�,���D��q#�{n�"P�����V�]���v�0֡���Y~ �F���}$����.�0�J`�sA���]
H�b�'3��4;�N��=u"�10Uօz+��=i�t��{6���wH�o6�r�n���U�Ƹ��-P��P�"A ���!|�='��S�8��g y`���߳Da�d���Osf$����Ff��f7�a�ɣSy�J4r���[�r�w�W@�z���!B�I7!�`�B��B����x1U�R���)sׂ����+V���ts�Ȼ�wE>} ��z�l�2[�������C�v�����F���!�r�j�T��uh��B����:ѫ�Պ|��<��������y�٦7�'�ht�Md��d�Q�2Ҁ��B@�GD�s� /a�l�cuW{�W���h�F>�`�U���XK(�ڌA�8e��^IW�)�x2	Ok�����."�����~�8r�Et�LL�����I���<GZ�M��Ŷ	�7��>���&t�ųX���*@� &���z��%3�*b"��jo���i�YRg���VSF�1�~ka+1�#x�=��Xe������ދ&1�¯�Q#�$p$O�Fٮl�1t��7�z��j��ƽt&����YG�0�E�Cs�63�%cX���ٯJ^�����w�/;8�u�<C^M�S�gP���3�e��8&�w@��ʹ��9�Y�/��L���Le�����2�TZ!-;��ژ��iމ���JԔ����׸MhH䖒����abo��8�ڿp}��e�X�@(���
w�_�E����hTm�.y���� Bۭk��L��T��~���M������PƝ�#,��Cm�?��}�����\#�TNc�j8��į�>9|�D��Z�%��I�6�.T�D�}[:Z�X��� 	�A�RT�1�5;��S엝�B��"���[J�͘��<��7ߪ�}>�A��j�\ܩ`�n�5w7��l�-W
�tJ��w�.��o&���Ͽ���; r�O֑)�c&<�]�<k꾇�3���E�9��X�����㙒��c�4�uc�g�9_����PV.��O�j�1W�Î��r�	.0�-K��e��5���1 ���/'���U�o��s�T�'8j �[kؾ�8� eS�ݮ:��sy�l�!�Ϻ;�`�f`9����7�_r�1���P=�DLyV�o&��7����+�Ǜ��tɀ��~��ON�bvYY&�VK->E:���h�]�>����E�}��l�w�;�ob�{@'��V;�h+���F#���Z_�����q!�B���[�ao�0E�s�p�X`��fL������I�e.�����g��AxYP)̡���KQ:���)��z�m\C�h*%��r��]���D��
�S�.�	}8�?�Թ�ؒ����O��2��s�h�W��DJ>��"��%�u�=]���%
���;�gJg&� ����H.Y�ƃ1��	�����5u��H�k��y;ܼ�>*DM�-߫ր�R���.��[����E�?���^+��)#_x��-�#���C�B\�S�����{�OFLwq	��l�!�ԕiq��]ei��\�ڙ!�h�U�SO��\=vz^�� �Z[x96�vf�x#�����l��w�kI���!�Yt ����ܑJ���UQo���U��*������Zz~X}IE3�qO�� �\bڑ�W�+aD�vX�e�ㅃ�7�'�VJ�v?.਄WR�y/�|_,H�#�`����@+�$�F�﫠���M�K�����Q!$
���%�9�J.�P-D�4�TP0TX�� .4e��T�>�%vػ�p�-���$���I���Tj��*����"��~S�cRF`*��B�P� J/��n$�< ��_[�	��2�6|�{�s葝״Ҝ[����c!�|M���@X ����-Q'���Z?�]3)�m7�SoU�����A�x��"Q���ک:�4�<��D;����T{)�lB��heTk�:~$8����!h1�p����bpr�B��٩�ي`(Y����:�ۥX���}��B&!��DA=�)X^��/u`fy���1��8��p�HG�~���A���B��2����R�sɡ��"�	�v��Y���W�G��A1G�}zx�5���F��Yo��+����L�۵�MF�rT��G�{��q"��sdl�@�8>S��̸QZEn�01���t{���`w�A�4��x�#9����r\~%��p�(2�ᑌ�8�ě58V��1�]����k�M������ d�e�Dh^kҔW�a����q�mI� 	%؏F`�	�od��,͋`M
�tE�s͎L9�yBL�����l�ga���6:C:��g��\�1�����݉_��:�e�Ă�I!�P�b]s;��B\��n?<YP��\'���r
�m���S���\ֲ���Ⱦ��V�*]���H����<�����:�S}+����<E�g) &��\�y_e�]�9��&�<9��r��O�ձ�Gm<�(�B��$"����zYN[� �I7�J����46��Ⅵ��%���q��S�'b�l@f�J����d,m��U��[yܝ�X�){���0i1�Ã��q�4to�P�`���I�^-Q(�"���cUWg?�¥��:��f���Ѯ�޽�(�m��[;��&�O��?���]�����f����&���Iwj���*�4��+��a��de�������a��n�L����}{�XZIh��� ��M����|] �7#SW��s&s�=讱��M7��<.h��ij{�!�1�P,�1���Z;m�ۗP�AB���0
K^�xlC���ɪt�k0�P���WHm˻�s>B�*U�R�Hž�t<�,^C+���t���Nu	n�׏�]��p��l�/ra�J��ʽ	��%r� ^�Ati�\�K������J~%�����2�z��@U���w�-ؠ��B;c��L��&�KB�ʁOv���"�Z�I�"^ׄom�%�h6����x����"w���:���qkmR#�ny���v�VV�Y���}�r�c(T|��Gf�<�
z�2^s���q����BB�_q�VğnnP�N��AYJ��	lSgF�K�t,<O��Ϲ6~p���I妁�/"�m�ݰ/3�89/s�r���g�K}w2���G��Hc�(�9���l1CB���qȃ�C*���6��8˼����o|�Ϥ���=M[�ҙV:��ڬ��wI����2�Z�������"$�`������6G�NΊ��v5�9я�8s`�_^z\��P���6���@Z8{�R��
零��By�P$~����>%��'~�*�������a���W�{�w�*Q�wp��)��?&�|B͒� h��� �$�M��Q����8�0c������mh����WnQ%\	�ڈF8V��Z��V9�ܭlE@����8�RV�N)k�(��:x0f�BE�fQ�N�_��I~�%Oh�J�4g[�G���Q�D���v�O�Uw)P|��kVF�{����91Kiģ�7m��R�����4V�P���|�l�)�,D`0먳���-1�M��zt���,TO����.��Ok�2�f�D_9����䍪L��6�{�L�Ȟ�����&Wu!�8��� ��PH0���[����/H����1���#7,�&��s��̼	�uUJ�:� R7Y����L ����N��/(��[_%;o32�Cl%��tp����V6�͘�#]����z��~�Xi�>�.D<7p���j����� ���%���]�-u��ج���:��r�_N,3�I�C�u�ʴ�@����f��!��/�F�QA2�Zw�����$^Bta�[�+$�t'��o��Hq	��zPx Y~D˪�^��ʻN�3N�e�G��u����ɐ�`4éԻ^�"v�`�'q���k×`�y����]ј���}8�-x�u[�Cky����$�γ���Y#'�ppq��s	�W:�O����L��"4���hҜ�YJ��x��4�Ch���j?��u�o���?/>�MH��e��ݱu�z%�k� bT������}�������s�c�;~�+'��<�;E�E��j�Ct��{3�I�����]4r�[��~��TR�}I=�@�(��s_��o�o$~�F��p�'M85f�C���#l�<A�3�kH<s�qpHN���F�j�j���xe�v�A��o�0P��_|����܁y���&ͫ<�2��Q�<�1�68Ra�U�??�̚�
TP]���L[i�po�U�pய��~�s����Ky�Q��� e���4]"��r:�z��X��к�d��� ��g-V�<�N�C�~F���e�a�viW�^�����[�:P�g?L��}���J�\*=z��S�>էn{��!���v!
l���,�X>�vK�3����>����%��_��/��N*��Ã�mlD��y�����	�eX���z�0z�2Z]����Y"��׹�|-b,<���c���X[�U���{�ǻ��=��o�_P*������jC����4�bx4��+��x��i�UQ,}d���4mZ�o�b[�D�]����O}��=��8���E�@L4eu�/��h /�kP7�$R�y�i���?�w2�#X����,e�����&�џ�S�u�Ϊ&��vaU%T_����4�#�+���-���>i���v�����ₚ�?�8L���c?�~���s	�iy��M8fX���*7J�ږ��3�>&w��潶���Gq0#m�f;�����B��|�V��k	/�	k�q4��p�Ѯ|���Ɨ�_c
�,��$F.L������a2w��x�CΖ�w��)D-�{�U;���(�$��2Q#�i��@���D^zt��N�w&��c��hO��4>P\���m���Ū��%�;�����̻��ۗ���-�iCEU��|�I�*cW`!�q��&�I	D�e�ހ��d�� ��}\]�C�	���?+�_���E�֧���w���x��:H�D��C���q�b
M4W
���z���^*#�{��������p��܋�oY��cC�ʥ��Vχ���j��n����SA�� ��A1�Ļ9�Sx��)�{$_�e��K0"Y������{H���5t�m�v���J33�v��Y;Ĺ~R��A�=�5��MĒ�{�ʪP�zA~F�_��ɭ{\{���z�_GvS��JPM��+����'����X�<�f�g�y��5�o���2�I金�l�fIx���m�}���f��Ͽ�7E�iޝ"6�d_�l�!��Z�j�]�Ju���$?[� PU�F�S0�m?BsѼ�t�4��g
2��k����]X�o��
!��WޜZ.�%@2�LB>9->�NʏD�i6�Ժ�ʗ7ܶ� r¸l�W��,�m����S�_���u�h����^��߁V�P��F��V���Q4b"�����6S؃�N�$��[qb���M����NvJ4��c�r�N��P�[e����d�ǘp(.|�aTl�[*j�D�<�N8�!���=
�#%�}7��(�t��h԰�i����Grb���U��
��Pg���c9<�X��!�~р\[ڇEFO�O��큊!σ��BU�wq�\������u�DJ^�3?����e9	`�n3��}��I��S��O�+��fR�-��;��6d7�j�ss�����x����ȧ�`4��s�0P5I��\i
N�t�B����j@��pm3$����9�����]���@>�[`1|i�7GRۨ�|�q�8��i�XF�5�f��[z�����ꑏF��G�?EL���ˢ*�9����F������FJm�Y��M�T��~ ����Tu��l�:2(蠏�桎ʠ5I(�E���9)�o�x@A4�c�f�ō�K�ԭNޓ�۠K��@�n�������]1m��mCXepc���l��TM��&��SRd���
fq�-���P"�i�M��K�#�?��f�H���"Q��3⢵����P�N�og��'o<�8���\YG|��),YZ���$�lV;�6�Lk+���}�o#�J54߄��A�y
�0����|���=0oq���VT����N��5ל�}&@����0��7�3�y��IDLW���_ �66�ݨg_�5�(y�+���6�@ړ��	���#k�J�cҼ́�Dr����3A�ʮ�|H-�D��'�|���!8,-���A[�vJ�{��t~M�Rh�|Tm�:��A�U���_��O�Zm��V
��P�
���.�V]�JS�ys�zg�^����Z{�7I{x�h8ſʳ (���>i+��f�G��q
W��v���D$�����Pqj.A���.��~����'ϑ�)�
���Kg>�����Oq�BRi`��#�RŔtT)c�+h�B�Ĉ�G�r��*6N{��[�ށW���vگz��H!����D����"̪���~�nz�szR`�ߠ:����[��z��S-��+j�7Y!��bMzhc.�foWZ�&��.�z̋g�*GgkGz�f�+F$�	���I���>[��� )����Ko�[�y8�&ؿeÐ�l���@�;��_�]?��ئk���i���"��۸�W�/~e���I=Ӈ���WSգ��U��x��m�
j��%���rX�g?Q��V�A÷��t@ ɀ��M��� ��������4k��g+��sAk *~oMh1(>"�x��	#�F"B�G�HrvG�H&m�).\(z��"��o�O�UO�h������_79]���A���+�V��YCd`�\�ѯ��۔�+tć�#��n���0!Y�-Hf�w�u>�
�F6�B\��;,���<VJ�e�1� sO���=�sYto�4t�/��# �} 9��s���D�Bm��J�G��:�,f�#u�׻�3a|�⣫x����`�� 9Iw?�}�������@d �J�n/6��>G�Zj+Y��Us4!�T܃�Ȩ����}H�&�i�`�]�9"e�=�#X��ㅇ0����.��|hc��0�-m�ʋ�����¯�!��7�q���\VL�3Ua��O�x�лm��/vb�4H�r�!s��Y�T):辵_��C�!�iȅCet��v5L��{ "�y�O���IA�^Ԧ���Ln�!i05L�e�j�"JB�������:Q����}̭�@Ξ�UL|���_����`�a��"C8$�P�?di��	h˜a|�ϗ#�&�w���3�S�޶��R1���1y0D���wh��������E$ߵ<��Q�_����l(V�o����������"��̧5�5��0߾0b��i'.1RuފwVs��m��`���1X㢀I�A�W'�
l�L�����٢v����>n�8���=L@C8Tn�hF
�Ի���Z����2�+'�����DX]�t���Յ"�n�
LL@Y5
�Z],�Z���x������t޿�~*o�]�GV��� W�c�����a7c���p�,j�����,{m_De��
�u�PÖ�Pk.̸⢶H�����/}���D�?J�I *g�����H�;�}�T��j*����� �ګ�.�� �ꖛ�R7���V��8��y�+PEr����Bx���./�a�
n���"I}3�V��(w�'�:�7� ���r@�82�[u��K��w�σ�����0�[��`o��x@�"�6�Va��]�8��8G�������J�wρ�E{El�������mS;��.)�P�,����q	dC ɦh�Ӌ���
������݆���"FIJa���k�n�S.,���E��W��pL�=����ڧ��z/����l/�k��_Ս�k����5EI�����jß(�G�Ʋ�����R�4!�YЧ`���O�H��V��2�����>:p�Ю8�Ao?]k��β_h*�V`5�(2�79/:Ne��s���[`�7���C��P�ʦP���}�,JN{]Y���tS�O���gr�M���I�v����y�^*�v�:��*ޟ���5[�z&P ֊@-(�TWW����/b�����`1�}�K��!yTI��lP�J*��z�&�����tc��*q���n�?ଖ>�F�ep��3�
��$����t8H1e�g�ms��MT	%i���}�O�#�}�6�/f[�.��ߨ�b������a�qp���,��+n���*OZ����~�c��
�)�h��Ћ2�!+��!N�	�I�qHA�g�,iZ�W׊�/"T0#H���0�>���n�}{�[��DF�FU��"�]1��Â6�iC�WSQ�לtk��|N���_:O����mƛʚ�[�����A"��M��>O ��0k�	�8e��֏��ِ)�{�k���nlqa�X�p� ��e���Ko��p.��C������Ƙ�
�?P�Zw�]N�Wk�[5��ix�pk�T��ED6�z�(��|�?��'�^W����E(5�K�	f�����Vz���t|�A�}q:U��"�����T8����z�؋UE�D��rZa6�a,��Va1�]�n+J��L{��)��C�M��W㔔��E*��\c�r���br֌��]yM؋O@�I>�"����;p AKj=�����L�e��-fV�^���(��9�wO�:3����<�����%Y�����r0,U>;XEE%�9�ͣ�d��P^JRܘ�SuQ�I����Oʃ�&,0��(�ﭶ�Ԩ6e/bC�$	�� �H'�V���'o��ÞY��W ��+ �"a�����|�z����c/�øXU��7�M�n�' �f�Z���wo>������Y<ud� �ϲ��;�Í[K�4,��Ě6�uO�yʅ���ǰ��o�')��=445ζ�+&��
B��.��wNX1���E��45�u���/��\FN�����YpM����AQ��U�9ǭ,t%H����L��d'v�m >�V��i�+T��S0��a�� Sc�/�4�	�6e�p��q�6|Z�0��PU5�雀*��i;�hn�8O $���DR-b���5��&OFL$��X���D��TIg��5���	��ɦ"�kT�>2 ��+d6,���W"q8��s�JĹ�o!\M���=����i������F�SĢt���s
1�A5�n�����p���.,�j�3n^� _Ym�N�iԅ�%a���g�_�qDi�L>H4ɝ|ebL�`����u{��v��|#a �{g�5�c��"?t����t'�Ğqe:!���N"N\tO�x7�-�M}��Hk>ܩ��Z\����46̌�O~�g��l�]����C18g����;�j�B�i�2*�_d|�{�|�_�E&�f�p��z�.	�>]� ����6�i��@�N�*n&tL���c@Q׹�<ɞ���<�p��1��� KֻvM�|(EC.�m���r�:.��6R%�d!�a�\�=;ez�|���h���40��0�b�Z�=v�s�t6��3.���lS��Qb\i�FO�#�T}[�ͯc˶��0r?�'Q�}a�J`��zC�kLb�c噙� U���.y��\#��/u�D�G0��0򱘗��|f/���Zb� W��i�ƨ� �-�'�n��y�=~n����:��m����\�ҏ/ ���O�Q��z^���az-�"|�Q�p̄Ը�
wA��#h)
��P�@�� ���h���5*��(�ve�yd-6�bBJߵ�8���G�Q�w��K�!k����OߓN��Ѝ�e�Uw���\�1vX>�,td��Q�}pzYP�i;'r�Tڸ
�Jo4��|g�I�����`@��t�D�����e�cЊ��}��L5��:6�T</�C�(����������G��.\��+<c'W�|nO� ~�ץ-D��W�qv�Q���U�*��r�r�d;+��Gv��<�]aI�ڨd�����k��H1��q�����vh��e�I�X���������Y���Ip:"�Vړ����?a�jT��e�r��q��P�o˕��Ci=����Ck���4/��n��D��Ci��>��*�:F�tBʉiZH"��Ϧ<��xM9�_�!:���N����.��O�:!�H�{�p,>���}]�ng�AW`K��*�
cZ�]J��h����1i��X��ꭾj���"wL��cp�t���($�c��%r,��/r5��	�]�s&�~Q b%hw� i��� (q����fZ�$v�TV�C�����uG��q`[(etᝬt�c��U��jY&k:�m�y�Ǹ>����ќ0�"�y�G]s08Ύ��I�����7�1=��C! �c�G�����V�x#	?�D��c�1j����Մ�*��Es(b�n&؉^���|�( �x�����l��TB����'~
���%�I	#���d����8����7�%�T�� �w!�\%Tl��pR��H��J��W�U�%65��|r���[#�=:���P�w��Zf6�xK����'�ʄ%�K���O==0}�yݒΝ�Wb� p���t��ZC�+|6���"������5�q[2�[�6*���*�ȸ�D'^��������P�a����5����+5,L�H����T�vN�ݲ�wQ�v҄�1i �%=?���`u�i�c�:�z�g���y�Z��`m?�.��<}���Vr<Q�+#!`%��"Z�A�U6>�VzY�i?7y��J����:z�jR�'����ʤn�G�|>;\s�߭���$o`�t.ś	�)����W�rg�d���� ��S��(D�"��1�@��"?v����7F�h�����i_7�������kڭ��W&۪ɋ�9%h���;�&�u?��-�����I�'O�RnD��Tyc˂gmW:w����`��*�7b���$k�3�Ӎ�.���+���Ṙ�~Exf7WW�T%��!�x�m���rĢ��;��9���{��6�]+m��a�f*!�d*������H�d�S�7���T����ɺl��i��m0~o�� �%A��ٝ�{W	@�b1�����8��!Eb-;��
]&�l���Rp��r�+�@)CG�٪W����?v(���������l��Ŵtc����:8�I[�7��y�0V(��w���&~|;< O�h�D�����u�;�=h�[�X�F��y@��� ��04������4ݾ���6<#��Y���Y��*���1�3����	a�}��o6d� /��Ve�r��ǜ�m�B]��:G�9i�C�Z	� �2��Æ�[�H�@���6�/yQ~�&���W^KMV4+X�?�u��5�ј��?��6a��X�sA�aAk�Ⱄ��=��z$�٘��d����Z�Ajܶ��=ㆸʧ��{ȵ�{Bz�m1�Qgm���|ִO������aْS`���o^�����p^���xܓ!����	�f�e��W���dxU%o7n&�I��r�U�k4ʝV5��!�NN����Z�ٔ!����[�$k�V]�Ǉ���f��G�F�@aj�K������jfC�[?��-=�FB���۞� K�vǄHA�/��A��oT��>��9�"ٶł+���a.OZ9��x����{�����P+Y�)O�C���lq��޲����|`s�{'`Izp���&�CRwm�N!��͟� 9�D1����B4�^҂���11���T��[qX����&�����Z �a7Z��&�-_��5���c�޾^7w$�$Y��{��Kp�r���)�y��#�q��X���C(�=�R	^�hə������ެ"{�pQ*�q�b�^�l|��3��N����䎚nP��x/�����A��J�bҰ(
E����s9�T�t�g�A9��j�>LLu7mXܗ�s)�byc|?l0��1��]ZʂO���u��2"�T1qh��̠U�4��k�k��Þ�2�`�K�.ٍ�\�2ϣ6)9�-v��6۽���=I�\,X��,�A�\	(�{��v��j�,/Uf����G|�7���o�꫒��o��f�O�"1- i(t��9���p��`���og-t}~�A2����Haw�Y�؅.u7�U������ɸ��;K1r�� �L'��9جJ^��q��9����¡xveCy���`�e�PY����zz��l��*�Zb3v��°!�)��:���U�7g{�$ucY�{�9��#0ub���.)�jn!Ն#P�x��2�`�,���!�1�­I]4EQA��m)�T�ޜq�G}ѿ�e��RZ쿌R& :U�%�B->��C���!��)�7�x��a�A��_�BUB����b3���ؓ�T�x����[]t��m���-_$k��N{�ɖ��_;��Ɏ�j�'�X5�74_�<��A̼[9U��m@Y��0AHL��^N��yt��%���P{���r�t ������sa8r���&�<3�"����V\]q���9�?������u����B:����j�6�|�1�EP:D�H�|B��q�C��z~����
.3V�w?�t���p+(���>)1.��W���3�ƙ���%�.������
]x�*�ȜpTqY9M|�����3x朄�MH"-���t�HW	M�	���X]��;�J�ɻ�^wm���C ���8C%z���0lZٺ�D��<_r�o�d�˸���k��!����X	˸�A���R_���pO�	�𺕉�Kp���e��ߎ�-z	n��L/��.�*:�9�7 �С��3�&*1�	�hYR\s�p&�[RjOY�;�ȩ����� �3��k`��B�ml��*ʜ忣[��|ƾ�7���r�s��u�ä��Ѐ���n�"�D-D���wP�3"QQ�x���7
Oǘ�p��4�)�����$�T��AҒ|�m��XnHile��l B:��3r� �p!!z:1fP�/�Q�dS�l��Ҁ1ć=�9��ARBi:f�_# C&��4��`!�c)����^�����&��خNx����33_r��6���QA�%Q�7�aa�^��ŕm�*  �Z<4�;:�yJbl��%�N+��5&ˉ����A� f'ER�b���"m)����� �dq�z�7	<��F�م$~�w�yh��.���D�8_0v��6��;t41`�(���ٺ$� L9�f�%)�DK���w�#m�;auk!)1=�������|����.xb_Q��<�A9�t7#$�������A���bͱ}��D�� �����%&0��]Ey�� 7�p!��h�xW�K�L��ࣔj�c�M����Wh�1B�W�9rZ��ZQ'L\�̣Hl��?XS>��!���'�����8����&e�m3�.��4��nE���~[�Zۯ�$�'�ib�/�O=�4��l�������	L�>mU��68}�]���샑�q�ȴ�V�~S�L����]=��B�5�&�]沄�Oͬ:Ȅ;��q_qس;������q��fGФen��qf��P�x���Eqӳ̖��H�YB��0�Ug� ���~���|���JhFn�s?Ja�>��	*��I(+�c8��*N��µ��[�@k�j����T��6^��?hh���&RD[O�M�����Q�'cO�uV�Z��U��"c�ؗ�)�T�0�a&j�u��۶q47�SiI3�@(=��ΆN��a5�D��]�~S�%]J�|7
­�m��אh(X���������������:��_����P,������Mb����B?�7�`��9�r�&ͧ�
�(=������?4+l�P�+},^s6�p4�b2����69N�g����A�10�C��+�p�a^���G�4����s��Ő�E0�C=�n!�%�vgt����LN�PЗNv�=뤏|�ñ`�i��2!X-y�b|>����B=�-�Jl�T6��8O�t���^̝�t�򬩯��Ym�EZ����چ�U[H%Z��ʳ���K �2�հ�G|'��Lg�Dyh��)O+L�J�4�*ŏ�hlGow���Nj�| ��y*>�Uh��Q��i���A��6d�%�+Gt�'	q���'��<~�1-p��P��:���E鲊#�*g���<���/El�O���<~��ñ��.�h�ƐiC#׌��ѭ�瑲�M����Sff��a.%�'�מӎ�ZW>w����+���� �%K���]/$2�i�_&�Vx^)��X�x"��~��t]�%���$�*!O��^�rՄ9�xY�\AY�;��\�<*�WiZ�IE��A�"�ީ�WbC�ʯ���Ű�)ew����6�el�0��JLމţb}|�0(P%��ծ��jo[�7ӗn7�u�u���zc���g�r����j��D���p=g	2����.IQݜ��ШS�P������n��iv7�T_���&�L�0ӄ�8v2o�G^뼺{:�ʜ��3] r�8a8�-!>���>K<��N��� Ё؆#H#��O�6YJ�x�-W���	D���P��5�)�2�k���P��� �E�Lj���}��Ae�W������RW����t�+�yg������%�?��ƞ��R�5)fE����F���	:�C]�Mt�4���Z���3�Ԃykv���<?���nLYMrj��VٵW�Y���u�S1t0Uۭo�ԁ'�Vz�,�H��B��K�����@j��?8y���g�C%�ϴ��)�;��2 �p�h\Oh
Гq0��o#Wъ��\�%��,�J#�a����!��X��� E��L��l3�;֐%~s*P�6R��|���\9X]K�r�������N��iK�aV�TX
_�R����>�B����̕�5a�f�ӫ��C�~�r�!��ƭUl�%��x�l��7<_�L�cGM̫��i������S���r�f3nA?\j{D�ԧª�f�!|@����C����,";�:��|>�,�OJ%r]���˖�/�g��6d0���w���v�C��(�`�'f�{{�Ϙ�!j�R�_�)���s�`hd ���7'A��U���,�a�mq�OS<���uc��'����'�����>	^�����<�P�IP��.+�8�뻂SRp��{�D�}9V�qRD�]�<��3��HQ!���
$G������9�.@�Am��[j_�b����֡�����u�k)bk�ۛ�uVp��W�y(�n�j�m�Vj��h�k26����%�R>pfG-�b��Č�kE��[�fN��CGM����͇��6�`��gcP;��CU#/'V�����J�
0&���$]0�A��3�"rr&/U�6:m���<�z�6����B$<t��L��o�l��.E�
h�P����]��2���(W&`�RT_>�.�_?*��������wճ鎣��[��BIw�gނ�J�q�3fPl���qf���p��T��$��'��ye�\��R��#d>b�g�L�+�¿�"�b1���[�i^�o�k�#�5��ؕD��^F������:��Ч�,��6�}x���)�}�$��e���F�qw��
���8�/_~��q�z��Y�D�̌$��ӯ��e���;�����z]R��$������#�R�8�=��Nk�`�Z�)��#G�NÞɽ�9Z	���E�?�}f	�)w�� Ƕ>Wͭ�K0�Z�>$2��R^̖Qq?�
ǡ�VHf]b��;L�ޏ�m�p�,u���ߖ���bБB�3M�((]�9��N27?}dc�U�'�a�L�<�>���F�躹O0����!k�X��f?�M�죪j�O0�*� �Ν}�I�Nf��8$(�a��,�%�O�j�qȋ��UUb���l-B�#��1���3�dl��
$�bx:6���1t9�z�\m�$
�S7�~@��|{Ra�τ'�8.C�1���B�d�)^\�/I'�=�͌���3eX��L^��̢r6��őYջd��<��6~ҧ;�/(J�����@��/��5�	�����x� C0@��d/�&�f����ѧ�fX��B&�Дv��j��,Ӊ�2�˘� ��OЩ��I�ק�tTOK�6�����N��vʦ�0��ü��@�:�+�7���&�R�>�[���ι��,y��l�	a��z:EA��a!�����/(l�j~�t�{��AC�3:��+�QȜ�V2�$,�wèv�Ԋ
�3�$�r��5��٭\�̑�4�u�B&1�MM)D�jXgdݍ��N�⹫�5�K6�Čx�����|�u�K��i
&k2і:�n)4}!�3�����!ϐ		��]@�c"���j7�.��k�3��uf{FW�$�T>��M�z�t?��
Xۏ:�[L�%��P�uN��9�d�1��N BN�M��d��|]0n�!Q�����P���^�4�1<�����|�Gf�b��m ��{����H��b��g�@��� .��!C��dwў��At��);`Ƨ��3x�t;d�$�%-!֕��+_s���O�.�z	h<��y�i�%�g�PZ�"A��ݏ�'�z3�]Z�z+}Zm�k�0fm�l�!�Y/y�[��X����E����zم+�T�I�ƾ�Χ/��j�C�r�J�|E_;�XV'|��\��\���r�%KD;���`o>Op�x��(�dq�ښ�*�X���\H����� ����ιC*�Z��#����x��st�����$�9ع�0ˋŽ��F�FP�4���3�h�����c��z�9�H'����y�[��1E���n,o�e�k�܉#+P��\�/H�j�D%�UH�H
Fz�V����"�x[A�1�;v�A���q��$y��m���'Չ���n�J��VI�Ը--�,�\f�	�E"Q��N�%�b"��2��jz��l�[����5Ѩ�T�F�t؉�U`�un7��,�8R��0LnK�2h�E��� ���Ƌs�
M�t3`���ܺ��1�X�#��2���y�\�hP~�Uh4a�e'��#?K>S+�̳��[�d��h�8N��v���E����8�D�-�����E��"��ŔDSβ��'���Pö������R�*��4�|�A ���Y��yIm�y�g>�7�?�8��R[`���c�S���6\�;G7f�ݢ��y���jyQh0R�=�Osb�4��{Ve� *�MB�8L�r�s�&@�ږ���j �����-�榗i�Ш���{P	�7ja޻ﭼ ��P
����">ݝF}m�����kA��:�Q�̇��\!�l# rWF����m���k���t'dR�5V�ǢK���"��'��VK�d>4"������0��фl�s�=�͇�BU:B������襽���&Mj��܊�W��NK��k_����',�d�<7+1���ܾ��`���մ���<p1O���9v%4
ɰ
��g���܊S	P�3:ȧ��=Q�j޷�wW0X�\,�X逞QPq�=�Ha|`�HJ&j��a�~��`U��%�'�g.�9�e�ϳf�}�Nu�5�y���+��Ϯ�#��S���[a\�^w�a��*����GTY�($
C�L�fd�5eH�=ޓ$8�AO!��f���dZ�\ˬ�$-�g��c̨��qy���Ҩ�B�@�FNn��F�@�|Ӗw��g*�R�]���Ob=nY��u!kd��l ��G����k�Tfs���nhd�+��� #;��Ի��B�O���� �� +��~Gj���^��8�6����+A�' �*C�C*��t�r8	҈l]�|b+�$$H�p�6EA�d��Ԧ����s�4�f`}��C�NU�85��2�/DY�4���g\q��f���P�6��Pou��-�J���	�b�Erz'�ơ%T�!ҹ�	K7DY�͜@��ϳ����!��v��\��a�\#�i.j��?�j�f��Ԙ�k�E���5+�F������Aq���TM��ﻲ9Ұ~���9,l����wu�Kmߞ�EH��4�;�!*��MW[7 ���|�3��V�V�䘆�F�Sc#�1� 72��W�G~����y���c߁B�ʽ4x4�n�hRӍ���&�̲эʿa�L���y@���r:wq�KH�۪W��"���Ρ6���:�ȨƂ�Q�Ie�9�T�����@z�g8�ì�ހ�y��K~��j.�ߎ�QW��a.	������=���(��Q���u3����ޣ�����D��"��u|��EiC%f��+e�tե,.�BӬ�eH���[<�Oz3yS�bމ:�U4O.����O�l����>�\�p�p"��j��%%�eh�I�$Ci�r��M���on���p�P7@�M'���n���W=ӗ3�R�9^�8*@9�}Ĝ����ix�>��_:G��I�bUf���Tk�[�`^��ī��#}��}��~t_ʆn�<uX���� L�bV�8G��ѩ�O�u�K�+�.3T�70?�s	t0n��˯�(��T5��\�=�
�:qJ��yμ���L̈�l���5���$�i��%|9����Eȸ��T���-4���l�Ǒ�/]�`���U~A�/w�b��o{ ��|=��_�S�Z*R\��?���A���_�������*��eu�LL9�"LUI�e�!0�v�!&��K��3rC�[�1������v�&��͜�u�c|�Ύ�V^��N�t�H0�v�rI�}"�*})<]-I��a,.����uj6y>������a�L�>?gw�q��p˹�ݤj�e}����V�N��L�a#u�3&@(����[K;��jI�@�hv�qt��X0��(�hp��-�|LQ��F��5^śȭr�V��AA��a�ґy`H��ɠ��4w�6�;S����%�gZ.dK#>8�*��0yb�w?�|���1M��-�(�X����X���0K��oU$��|4� �ɪ4ɩ&*�-M� �]&(�K��Ǘ����"�l����W �1�w��l#���kJ�߇�{�l!�>�dϸ��U�C
��_�a7��9;�
�Ŕ���4Njr�: �)����1Ya^��x1���љ{���2����fR�e;����#��f.&�$��zB$P��¦���7)��%w}�;�
.,�*;�i]�Գ}�/�P��J���S��z�p��ʼ��s3z�59{<wh��|�K�z����:���Z�p�p4�.��L�WQ����LT�6E�e���D1,G
*4���3V�����$����=�p#Q���z	y��Ō�H�����h�DBf?��w�����A�6l�upk��5g<��cB�������;�l�'%
8��$��0K*3Q|D(�#q�Q:��iQ#������oR6"x���� +28B��YzA����4�v ���?c��t�x
��`�r�Q葋� )\�� ��xБ�c�S�^!���11ɚreHNc�"Cjq	C�kE0=2)�^S1'�}BayQ�������~����
���im�i�e����������+V�͢Y�)k߂]�2�c��F�v�W���V5�e,:�^w�L�LZz�jG���p}�U�4���A�"��~�9�F�A�����R7�t�u�w�]��DEkn>�d��v�J�w��jyEO��d�?��x�Z�fq��L%+��x����it��d���	�j���OԻ�g�_Eǽ������u8Zo[|��pi����stG�P���VA���(,���i1Z!voJ�jNk<�O�?�j��@/;Ʋ�}�����r���D�}���M���|e�><�����ן�q(���ݽ�����Ȇ��T��q`9��ך4�G��ч�4�#U�T��
X���8U�����6�u=�K�f@����{6w2B��uk�^#��K2Ua��Z4�48�>Ԕ$7���UG��z{A�l�^�"�N/��"���p�W�)�!bᯣb��E�jN� k1й_�E}0a3��"K	��f)N�A�y��Z߽\�b��E��@���I3~b��ґ��:?��O�|qXYl+�i���3�C�rF���#T�\@�Y1IM
�'����3P#�Y���]�]{c��*$T!Z��䜕�J�.f���f����¶}����{�1�{���|QS�1�b1_��Y��cp�ݘ�����E��s�³߽�q_�T��G��P3
XЀ��&����\Ѹ^��fЏ���p�M�W>mmt�L�+V�j�H�lfN=ǆU+Do�rjbZo3��%��;�l��֜�r�}�N���im�Z��F��<�m�f�<�8�ƕl^.y�Rv1{�p-�]f�z]l��gtH�,sQ�5��d���:�`
�},�����
sJd����E�G���{ ?��j�QK�����;ݮ�O��%�ہ���"�pI�"�D�,ga8�-��D�����w�|��Yq����\��/\��U��{�}��u�~9a��>��e)�B���v��#R���h�<�>[YzB�~ٔ���Bف9�!� Teh�ǥu�y�� �si�Ɉ���lϔ�5�D��S�į-(��2�d�*m�O0�qH 4�D핸���,�xM4I:�@�L�[dX<X�赣ϯK��^����K���f8�O���G���ەc]�����c���ݫW�iF䔼v�v��B0�x�ZÄ/��dM�.�<����Z\�]=H(�H�t�� ����ER�]�2%��M����U5FL��yqi{`y�E��~׼<��!�Ʉ�5�	�R��C�l0��U��p�����w{ f�'����#��xDzU�WX��bp�c��S���D���q�=�a �0��I��`Li�ԧ��c��V�����f���(��I1e��yO9���+h=5����uY�]*/#B�U����y�hIad����]C�]��+4:O4�䲑 �(_%�5��ώ��ʳs5�N(Y�[�@'�&���IR����Z|�Mɲ�)0^�XJ��R���P�0ԇ)N*g�_�������#�H*��>S:�+��*���fH�g��?�ym��.�0m�9����An�R�;l7wG�H�����������dޝ;[� ��%�\gl]����g^+��/��v೨�jJLf���)~���V#�V9���י�&G���̵a:[��77���E3B �29o�R�a�ī�?�COۍ*�����b>��(yʆlO����K���JR�FDqխ�
�nh~�0��@BOm��{p?��;lt<n{�d��h�@*1C�.7(�$)�,zǥ�%7Y-M�,�����6Ӳa(
V�İVf����o����`ۚL$���ި�K&&�)�4$2P�5W-R�}B�!� �t���v�)S���yIj�sl�iWvSU��PG�20����ζ�p
�%"aВ���� 5�ۯ�'�4ش��"7�nd��qŤ3�R����y-���4�	�V
G;ti���؉��]�9C`2��z�Sᇜ:�I����p�Ƭ'���c6��~#
���יX�2��f>X���9�f�Z̃ӗ�J����w%ZQo�����	-���Ê|���t��M�Ѣ���4��,���$����"	�fJ��,� @iϠ�0f�e��d�݂����|�Le�����=�l*���=�3�hA���ĸ�~��i�ĸt\
���������nv����_��3fT�?C6�-ܬ�X�^�
�E�xjP�G�!Z,@ ���j�+���'��
��/-O}�����lY~��Cn�7%ỻY���ʣ�s�fҷ�?V��P�є��Hn�y!�C7��ùvU(WouA��sRXfI"J�(D �(UG/��˦�T�H΀bl��[m�������X'{����4VǊ����SLD+�;�@C.���'�O���É+�B�|	�S�a<7/T��� �V�ӳ��]n�i�/�	^ۏ��_�.ۡߙ" Ήk ��[=��X&{�]Y�#�a���� �0�,�������JKUE�
�:=O=s}�xv��l7�"��y�l�Os��4<f�T�'6.���]�Q�M������J���������H�)0���:J��\�Jq�N�+�^�g͢��L�""O�8f��_&钰'��� ^l�����: µ�UG�a��)���ጃm�AwE�&_���;m���2&����I3Ռ�4�I��b\FԳ?6�Uvd��ax����+���O�>f"�Y6-.V� ^���i����m�y�Y��o�#��|�W#!~,�2#8�*��.s�,!��W��`>�͆c�ް;��*?��л��=������bҏ*Z(����,]�v��a��&�N$d?`L�FX2�mc"��{��S-�fK: ���=t� eSN!�ȕ^�λ�!ayt�B�Һ���5R:Z#|�l:��N'oC�a�un����}���8�S��a��v�8�0��.�&�%?�?��f��_�I�m��.�
܋��?�N3����:��+vT�G��{��3y߸� ��07���ut䦛T0�DȑtӈkC\)�O�?���_��6g	Z��GzP���D�]�1�����b��NhY/�΋8���<ax��,p��8׈)�[P��}�6"p���q�"�������v!Y�k��I�	�����e��cxE	~��I��X�Sk	y��\�5{f1� �������!3L%�]�R�)ٙ�T�����2���
o�PbD[++m�Ldej�o?
\�j�u����������n��y���@>+�G��k��2��ν����iY.�.ܙIyP"ŎN��S��囬PMA���������)�:��g(������3H �W�S�/��d|T陚g��`B��{�E~�Rh�����Ap�x��Bm��HvY»_�cr/�G���ƔW�RE�˳�s���E2&��2v�W-p�kฐ�)+6��7�����1$�����劣��*S��7q�=�U>j�Lok꺥�����d��m�໢���P��'{'�Mv!+�b�w���%��[%r���7H!<t��3����ȟ��*�W���)���D��Fh��R��i��X���A�v�)���G� �^h�3׏X6ൃ����%�9+�@p�窶X����yF*X�H��=K�
��#�BఠІ(�J/���~r��M�+ٖSG^�K�SaB5�-�--���Ӣ\%[rN��o�q�x�k��p/��El�Q��&��7dv�ݤ�}���,ϴN?��<K�������5�R�Ϝ��0�[pLH"��-�4��E��35B�s�\���T$d��z�Ź	ʏ,��u�
=�_vq��-�*X+�6.�X\�;Ȟ����K��h^�?a;ͤ��{KPw��I���n���-�Z�J��f(Py2y����;��#yˑ�T�ċ��)}�q����X1�>�Ki�k}Ie&�|:t)�cp<.�[�*�;&ĸL5�L��C���s(��i冽��A9bbh�i6��,�i��.]�ǡrQ�}�b	����ۜz��G#������j�ꋣ�:V�0�kt��e�x�/D�7�z�Ak"��A�7� �[�I����c��/���3���U=��`1��hʄ
�uʏ\�Ƨ�Q�@��O���U��I��w�/}��5Һ�<�q=�� �L'���C+{>N��ǸH�"��=��;��q(��jxAF����Z��ճN �W�(L��'�}P��i��D��_��=³�9ϥԿd���M�I~4�}a��4��*^hKo��	�BF�,lWz{44�u���P	/xE��y?rY�\��無W�_t
t'L��Ԗ��c����Ͳێ��K=i-t8���Y����kH�'�p{�w#�(ҵ��l��\͚$rz_s��#з�w#��� �!�����F��H vH�A�U�?l�?�5ߴP���V�V�[S�D��X!���]�D�P����f{�8η�`/"*��%��[����djQ\�`���u�\U��o�Ƅ^�J�A�W�O~%�'�����=:��ݦ�����T�^=�gȎ� g�&T抒1C��п���#�#�)�LK�2�M��#�r�Q����kZ*�
�|�ƈBO�ͦ�Ҩb�=kG>������KP���FOFZ�����5f�5�P��������9"߶�4��, L�߳ߟ����>��T�#<��yq�e��L����o���v��LY�.�&��I�$`��Fa5�}�o�Q�F��fO�UA2F�r���}�ec�����&�|�3A�e��,��OV�+���&�
t��J���2�<��S�"�6������ �� ����I�-�$x�� ��)da�{֣ +�RҚ��]���(������)�j�F�Տ�6�Fg0c����/�Q�N�\�N&��]C��h��)SCi�Y�*:�r�ˈ�-+��Oc|�{�!���Į�
4_A�{�c� e:˦y���a�ũ�8xqǅ�<�R65~�	ThNNnƚ�P'�W,|���������ӻP���0V�2r�=<�`��w���ض�i�	��O}��M�Y��	.�cՠ��%�(xٰ���Z�����-/V�?M�KM��G��}�>  "w6��d�&��l	1\B�nչ���`�c�>H�Z!��ۺU����H���-|0}ų�vF��sn��R�W�ܯ��ǐ�N#J=��:��|�?��b)�"X=یg-�֐G��'Vb#U��=�q}����t��t���e��9h_��Q{����*ŰPW�R0I^��9np:%8Bp/0��x�m�>��9m+���B�H��_𒂍t��>��0`�-뭘C������W�ETZC�B�s����h�r1��B5�Ĕ�&���T�Z�?��:�����z�P&���=���o��,�o�}Am�B�<�^�aX���6#Ҥ�|�����h�D��;��.}$��D�8q3O�J:Vo����);�R�O����1�e�-Ƴ��ZZ�~� L�GS���L-��ܡ�ަKd�cpKҁu6OI��Șχ.��[��ɐ-���z~�4��`�	L=�h�4ƁN����G,����-hU�Y�7[�Fe�#�P{z��8�M+���6 �#ta�P��}������я$�
�7�ϋ �dO|�����Ho���+�"��S?)S��* 5�Y�Ν���oR%*�Q��v�AzW�wd*y'-�hg�7����R���Dh[�H��5ӄ3`7o]�-~�,a�Ԣ>�	U`�
���.;,����6g�ZE6����D�Q�G%ǅ�M�3dqhny����"l��e�������d�"�3Z���:ޫ�{_�ボt�s~E�!��l�^��t#3R��p���Ĭe�ud���d�ӧx�<lb����
pMЯ��K�očٙo�o�����=A��H�K��'N�n��Y���AL!�cFv"�L��:}���Vf| ���0��G��4ľ��  xI��2��CqKZz�^p�B���)މ�`�Y�Hu�j
��p9A��j�y��@�1cvNH1x�
�*Rot9����7��1n��r����u��!�KwB�	����c�2�M��Y75�f����5%�� �����X��[ B�ʌ��Z#�8�0��)�;N���F	�1F�J9#q�x�8�e82��t�>�f2k��qN�f�tY�'ς9���7F���Hee��L��#�,�$@`I��;6�4����ӡN��j�7y
h�2@#�ͪ�.�܇fcX��נ�]~j�4�|V�mgږ\�����O�%�i[��_��v�;I�@�0U��b5O��3����72����y���O/M�?-g�/"P��;���NE�Cg01��|x森���E>@��:�J���]Ѫ���1"�c�60�=pqaֵ)��m'��8��&�.�;4����F�)�aЊ	V�_�ɒ���`�E����^���I47��%�véF]��yN���uͬ#_�Ʉ��y�_`�'�ա ��6�.��]�S�eV�?'����l����t����w���.�0������D!�J��h 'y$��/T�pj�-T:��,�WY�{# Z�/����+�?��������DwhN�\�����bb�ʈHu�[��2�'n�)�Dy[�jx�w�NǼ� �Q��0�)�� V?ar�'"�l�s��tL��mE_޹f,�7�p/� �D��z�����W��������@7Sӽ�φ���D�׹ɻ�Է�#=�J�HJ���?�ͨܚ�Ɗ��\GN�(],Q�*)��1�
�X�GF���U"��3�k3������|=: ���}I`#W�AfH�pԾ��cZIW-)�T}��F�jE�ʶ#��ə� ���d���v�?6��9�R�Wv#�y�sB1b�>�Z��r���%�ޓ5�6�gC8�.��C9A�J7����n%���J��a'j�����fJSa���^J�@�flX �x�=Q��70�:�xޚgq.*/ϭ$-ۋ�H���.ߌT�hԡ�K���G�ľ�X!!���~�5��l�nqC[`� �Ed؏vj
ݳ�M��*��X�j?�sM
1
��|T��BN ���$��q)��W?��x)��`����r _J'�T'�L#�j��a��3��3vl����ˡ�Zߚ��J�{yOƺXT_6�ٞ�lV��0X�1��¤tS෱}3�O�����C�)NL)��v��@�D�*2�rӛ#����RX<���$�����ߐ��5��d�h�ex�MZc�^����"8��Q���OWGPf���#
b]���?��(���>'����!��wd�D���0^qOsJ���FI���	uB��O-���v��8�D��&0߆i�9��:[�O��z�����D�4bn�)Z,�h��yxto�hV��t�#B��g֬�XM=��Z�w~\;�jq�(Q��YVX�k^3�5�����	.h���e4�<�X�j&�Sx3'E�3�'��4W�~�Zm���K��q���<�E�m��	hҀ.�0�Ô��~Ď�F[/��4�½M���������~�A(�����,�\���b:���z��\Q�D��͝Q2�剨]�H�f`��%-����N*�G�S�g���<:?�=L� ���~��f�qQ��Q:�&�6:��y�3y=	��=���0LqC�x3\9셍r
"�V�ȣ4��^d.c�9:�u�מ�����zU.&/S�&3唂��"��m*x@a)wA��5��"+��Vj��U�@'�tD�|�|�f�� }H��&j�ף�ڽ�P=���V �൅T';�Jx�҂S�ح_*2͢VZ(N<�H����X��RV��`"��zծg�GQ�~L�v���;�@QxO#�R��bDֈ��a6,�o��)���uR�q���|1�L��P4�����
(����@�Pi�EП(�R`%ii-��e���ku���|�C�9&S@�]@N�>܅F�<T\V���-�&v���G�@P��k��,�	\�-�8��G�ȹ'H�?��c�>�)�C(0s	s8��d�x��4��:�<��G�LRǰaǲ�n�!p�\Z���ǩ.������,�B���d��S�����khIQ�E)�}�(�/q�sսܔP��2�Ƙ�>}J�=*/#;�Yn��$T%Ǩ������
��;ev�����D��x<P@�0���[ܓ5���{���m7��k�%k�u�	b�!f b��+l2��=����Jq;ȂAQ�.B�0E.�Z0ő(���i��B�~�u�$.����Rʧ�=�D
 �ݤ�����3E.�(�ϣ��u��+
^
����\��>�x��X]Qݻ� !�!���G��ɗsF��M��~�1�%��?]U�BxE���ν*�42SӜ�\�'uG1�k�x:��3�J�ʧ��o�!�΀��v��ȃ��MWMJU~VV�0<U�U��ZQVȍ4[�nj��vzx��汶 �����	��x�G��P�SI�H?7�$�}p�����HQ�.�:����}k�7�>�TB��g��e/H�V��(Ïf]�	���?wc|�t]mr؄" uA$p��3n��б�Ym)@���J��_��� �T'���x�H]@Bt����}�$����ޏ2kąF�a�R���=�C.��okJ̖�o�~�A�Pc^����(([@�	?�OH�l�v�X�!�G��gۛ���=s�Y�8�I��/��`VS� +qe^�-Q|�p�̫�&5���MʯX��zAR)�ep6k�����*�衑�MR��
�g]��\�s���U��M���c #��êf��A)I��	f�D�h�?���.��B��~*�W�S�{
�b��+{@Y?��7�*�LaNL�����$}�-��L^7��#�k��.`�������k�� �Ɵ1����X��p/)(���I�d�ɻ}:�D<�M3DU�&Ļ.�������tt�פ 9��=�����~?Q�D�c'�����F^D���O�h�k�F� l���\��D�f|�v����*>�T���ǽޤ�~�h`�˾������M;;St����79E7=bH�Ш���.�����Tm��0?U�Ǵ>���o�s&(�Ta�rOZ�y��GM+Pw��Q�!�G���+\�E�--�j�/�؋7��ꋭŽ�ȗ��6U�c�����H�z�v�v�����!_�Z�����b�r��΂�H�\��f������4��JYZ��ۨj�Z.9�.Ozݮ�����sӥaMĨ&�g*��ݱ�v aX�C�^������R�
t��r��܄_bO���;�5�62!.*R�,�"7M��VE;1��p%�y�M�hz�,>l�����ÿ��.b�1�oJ�y�B���S?����Zz{	Mh}@�h\'����ͭ"8$F�j{5y��'����\n9��9`�Q/�,^sJ �)�����������¡8��3z"2\{�y/�����|&_��qZs�T���� xq�@"�I36�f	�:������7�n��ނjR��Ò���5G}�-���n��_�J�M��y!c!�k��X�׀|*b�吲��kz^�dا{�nV�]�s4\PG�|�����[s�K�+=��
���4tb2M݅�!h�潅q���e!Zn�ب%j�Ex_%L���<ҟ��s8}G�A�C�g����v��V���pq�8 !j;�i���c�����i�Q��hO&��!O���w8���N?&fP����Y�,�Wt� 8nZ�DϽ�#��.�'2���I��z�m�&}�����d1_$�˻�v_�z��MW�w���.��� Ռ��fA�Q����3�Y2��EQQ0��<���w�AV�4�4\�I�ځ��]�0��U�H�Kw����ؽ˜I�ud��<�[!U���H�"ӯo���SX����!��	C� k���]T���1�8ߤG 19+�0c>��Dx	���S�P�^!<�����{2�x��M9^rؚ!V#�p�U�}�q�M_�v��)���Ww��<��";和!�XT����cRm��X�FǶ� 5����^��G�!It�F��9�
����ؽ/��ʚ9T'ɬ5��8��b�A�'2p`�~��Y��Q7����Wc��Vx�<p5i{����c��z� �Ã�L�kw\�2|\aG������Z����L�!�9^#.�5��C�9iz����]zC5��QN�ڎ�/Fi.Ï���Ǝ�uח��%�k��U���3�^�8�_�:zT�]���z�E�b�=	Y5&d����ɝe�o>S]�Z"0^I�D6�˝�؆z4�-�����be�,˿R	��o�WTx���^��4�]���8p���r�5_(oi��e4v���J51�n{[��?<:1*��J�����rG��\�/%��=t
P�wq'��Z�[NԦk �7f?��U�����d���%��0r���@��X���U_�6|��5���>YS� �j�C�q)^���2��$���^�_�I�Y9±|���&,�Y~GE�?��k�c�:�
J}}ƘC҉gл�?����{�h�;�����"�oe�y.�v��F�,��|*��/�������E��M��3�
+dd�A�Oj�JW� d'���ʉ��Ȋ2,&��T&#�vV�
�G��f�|دf!�1}?�J����K�o�%��%��udu�rN6}Qˊ�����e�E�a�?��r..�.���r��P7�����*x1u
�r2k6)�֩8�Dn&�>3	��l�8�a=H�|��X��f7KK��%��\��yx)��H����r�tۄ��7�p���r�
'Z��5G�F"�-���q���Z�YR�P���m+��a�n��N�v����-�&���W����* �G����z��x��%�R��q�o30�X
���hi3h�_/���w�{�";<d����tL�!f��w�7�ĕ�\� ����YI�R�qQ�SVۦ���.�Cu	p�=�;g`!�f�v�_y�<��O�>DjKap�'��;��9T�R���{��*��
K�W���F{_��)�3sy,�A& d�4�=w���F�����֥�]������w59�:#:�
v�8���Ж*��.���J:g��lf�-��EDS���P-FP���}�ّ�M��'a���~/G�y�w-�w2��ţt��q�*��r[�G�Z�nk��N�ǡ ���h��>��VN�����+�m���r�2���]kV@n���c;H`ډn�O���ؙ��~5�+8�IՓ\�E� `�M���7��I�YQ��m%�_�yՍ z���'H�2&�x���Z���\gC�3��8˳{7Vŝ���V1�T����E�أ��4�Z^Er��'���D���o筯��K^�,℩�`�����(CSQ}�l��r|a���{cw&�x�m%_7i��;����k�2�e��>�^u�n���-�I��N�;Wt�Ӯ�������R�/uI�1x�g���47[�Qz��n&�\QD��r_���*c��n R�JF��5E��z������`�,'�N6������R,e��ZS�s��py�鞶��B�BD����!�#��@�#p�����J�L����CX�#�R3�K���`Q�Sh�	����/(tf&7�|�sS�W��q¸$��o�N[�߸���H�'E7���TSۻ���u<OR��_�ϘԦ۳���
5�=�o� �f0�wKm�u���mo��D��O��hS�u�1=�������mk� D�?��Q)��ը��DL���^ɦ��p�NSSPq��R�H0}����TP4�o���
�(Ѹ��o��/�n��e���������;�~S�ʎ������p�5#�\���8
ħ/jna��iJb(�w~2����}�rK��Ĉ���:}��}S�`�PN�I)훞�r )�z����Jh�zJW+��XB��GZ坍�9���$I���S?���R]�6�|xY�&12W�Z�E$��>^�R������Pp:c&��-8�Е�\I��G�;��ί%0�_n��*���4�Z6���!�Ng��r!9s��X�
,�;��^;DE�;X��x0���6�c�%�G��5�-�ɯ�0,[��YS�I�|��K��ҿ��G�2�RA�� �i �\p[�c�g{�ߙb��T��Q�f4���3C�����r��jt���x(r£(�0nmG��*p��_'O"��6-T]/O�*(M]��]Y72Ɇp>���
�x���ۙl,<;����$u^b�����G�׺�mBG�`��{V���TMՍ!�6�RJ~�6��������P�,#��ސ�}��f����S���9��UA�������>������x��#����XE�Ř����b�����I�яA��C�v�%T��&���޽͜3t�"�&�<X����`Y`;�S��S�$���8;j- D��`|�a�*5?e����B�7x�◶�/�H�T��%������v�M����]�Eƻv���T��}��	C�*�e�F$l#bv�N��+5�h��o�Fq3�W��>:���Eq6"���L ��g�;`������6�䃣<�W^���<U	��� w(�&eq�/R!�V�t����x@$TY��ȵAKdijZNq�e�sg�/Ό�eU��l5,�����Sd!�%F�|I_��њ�0 |��\����v��M��������2�5�Ϡ]U���~��a�{��?�YĖ�ߝva����ɵH-��Hpwl%�Ԥ����NI�JP>,�7��\��A��P�%#&��Pf��w��o~69�[Q
�ʪ��!nl"C�����S'�Nw�.�n�}��	�H�<����=g����|���*l�{��#��a�ٶ�p�ٸ��T��N��Q�R�1^��56�8�.E���h��"��π�0Ҥ��/���)���K۱�`:ˡ8b�buZ��F{�$�LO�����H'?6�9�2���.�n�;`$S���O�Vׂ�kK�1:��S"��.��2�vo��hX��r�R�Bi�����<�^�U �Q1�8�r��Bzt���W��w������Dcss�mUG:���΁����?��~ 0e.���M^l�|�nP�bJb�d�,�/In>&�G�+�8�	���C���:gh�Ԧ�B�f�̊���鈰��&�VYmg�'^�oy�z�`��gI8�~jFծ {�ҟ��-�D�y�M�GS�lTUF �c\�xGL90vY8u J�K�?�~��!&���IE����l3(4�-��n�r������Ps��*�����E|sU������Q$��c��@l^��Qq�,���$�_�g�U�_����B{�Z�Mj�s����
Gy�hR�� Auvhd=o�uT��2]P�qֆ-����S{��!O�z�4�T6I�Er�VeA�ȵQ?�2��k���K��6#^ �?���J_�$>1A�[Ŕ��vX��Նż;�9toN& ����V}��f�z����n��4��"���I�D�^>��A�O��$�G�C�@�u�L1��8�o&���]4Yә���+�qÖ�b���U�ii6��O-�);15�g7P�+pa��B��S�2�\SKi�����N����q��^�I��R�bZ��~6�=� (�I`���9��!�~tI�ݮ��c��r8�5�ݗ(�x�(b��B��f4����u���L�����`�2��`K���fg�aQh�_�k��}Ow��=�bА���G;�(�b���l���JrT�M��@��ȏ��qv�����mG����)�%QN����'-���:�SǆY����{�a8�Yo�8�냈���<zO�}4p�'B�5��/qJJY�R�?�m�ߙ�!���G�e��Z��n٥ǡ���⾪�/U[]z&\l�C��&D����d���\ �b�W�? ���F��F�0��#��D�!O_�ZA�e�b_��-�sm�����аJ���q�(�h ��<�^��a'p ���Z�2ζ^ݣb˺�Z܋�KV}N�Cb:�'/��/��]jm*>�iu�<7JJĭ2�i��7���p�i��οE��~f}����VF�.���mn�xf�7�9�A�)(���[��.cO|�tC�z��Ei����s �,r�y�]8v����ҩ&���C��9"T�Le�|��	���g�}:��̽�%�'S�#�Z��]p�����:ͫ'�T6k��H���&���(���jLpz��E�2<G��^FU�ŘJ���Dy���(M�P�����C1�c�v���kgoa����
�O�����vߑ��ܲ����nƦ�
�0;0����|&�Í�p�ދ�C�A��{#_R�s�W����%��~���ϑcSo$C�,�fE�Å����B���r#m8������!@dw=��C9ad5, լ�`�b�ۓ`��H�HEš��[%58�o{�X��)�8w�[��%����V����QH����돻��)�[�ڰ�0��u@���a�׌�%�3��A"=n��&���� ���m�t8��E0Zզ�m� �Q���,�
�C��R��m�R�|0����
�f�_����sH����I��.UtO�?��}��)uY��$��ƀ���̈H�~�	��y�ܳm��7���{19�g�m���O������n�Y�F�nڶhN̠Rż��H���S<�'Ɀ4u�,;;�!v�t�����#i��ș@��Q&4C�y��X�~���*��.�)/z`�\\���ǏX+�ƗRi�s�����{!�A;�ѩm�1/M(����0��W��1��T�$�N]��{�˳�+TƆ�uS6�d{l&]��3�o���s�_��H�,4���9.eA����~��v��f�X~3A�\��'k-�~�H�K	��p�E��#^�WW�����7cL�tW��[Y!���4����ED ��욋U`O���+��ɳ���c�b�,I��J��T�7����L��aA�Ơ����3{٤�bv�G�HF�S+R�
LE:D����p�
�bdp�v��zI��M/�f�贐9��,E�i�d&���ƠI�챵	9㋦��O��D�oQ���z�J mz#�%�T�Z	7��.�x����ML��Z�˻�����/:��l5�tU�8�q�\sG�3����HT�;��2���6����E�
u�Nut���t����#���]0�~�RDlvq����� z�!��dMl��V�w��5��7���x~$|�O^���sTB&_���ɗ
/7]}��4 �c�Xz���d���$���=�u�*5��u�{�d���m�T$N�/X�:@{�:�Ċ�U0{�=ma����C�{���u��%�Rw����v$�e�Y𖗯n���?��,# �s�;�'!b���@պ��`��a,��`%���?YI�(#(�x�*��q��Y��AOVʬ�j't�{~H�DcK;��(�+k��ZT���� Eͷ͠�Oڅ�27+	��-f�fςH�:4��� ��uݖ%�茢/�Q>dEW,H�q�b��d����ܬ��U�e[�x��c����-2/�+^����ճ����mQ��˼�uz�}�G��-"���R��<�HoВ�W[1:��L�(���]�jIۘ�4
"gg���,5����="��?���_D���4s�.W�Fpް#Ŏ[��,���U�ΔN��NSDfJ����8�S�VȂ�_g6���m����<~'W3����\�O��9E�d����a�~�W[շ�&�����i<���;G�24Ǽg�5��)��6�U��>iӊ�fc5?ΰ�۲�SJ)�MB��k�Ű���L0`[Q���z����-���\`R��~ιG8?X<"TM��������/��דm�	&6�$�����b,sP�z=�~>Zm*f>U�0{��J��N	/�n�C��`#w�x�s �����!�éӿ�D1v�����͖ޒ���2��v5/�)�g1G,71w<u1��F�H&�ZJOç㫴�P*�U�+�hhw���#�5We��N�[�}m2��sp~ֶ��{d�P�8s|У�ҁ_�
f+���/7p�	4��'�;j���Nq��	�;+	��>�DUXű��è�q���n��@b���aAmf*0s0�EP�P�2���N7���� ##<������ ��;�d��:F���.���i��i�&�����,pqN��<�0?F��T9�����&4\IW�IX�w��C&��v'-{2h1n&�U���1�>�'�STm���n�S��]G_e�$�E�=7M����`�kL:��*�z�p��Qɇ�vuђ]�`'�����g�K�t��}6�����[��qmoA��jK>��UF�>�%��](���@7����J4SBܦ��\��Z��8���q��:i���M-��`��y6dB%m~|%҃�
��6�) �p�լݨZ��D�g:�ǔ�>��W�.%E6��W#�����u��̹p�h+8�Z�g*��^GQ*4T��!q,/�.�S۟h�l�S�]�c�s�I�s/�m�Ȭ}�����MCY��,E=�6V��T��IU����v~�HhGӎ��?�8jt���\��5�0�,��8�hP�D�֕ O�dI;�|�*�՘��猽^�Hڟg�%�4�Mͷ)�C[��d�&Kf���=Ϊ�udo.�!C�f@sy-P7��g��ZBEVY�"��R魄��4�MO�^[�����0}:��Er�]P9��Cr��2}�"D79h�"M	�$rI�������G	�-�$�'���=u��̈́+p��5E3��7v� �hk�]����@�����̫���l����Һ �
T�ɏS�L䈁l���?���1*n���s&0�N��4�מ����O����ez_n����6"�&���(�4��Ġ�C��ǌ���sf�2��O�K\�p���!y�oMD�L�����n��5��FP�TB
��e�J�8 fop,��e��D�.;Z�L<���d��J�J2O��-�z�=��Ӝ�B�vD�Ú���$@So���.7����,�]���H�A�Sb-;M׆ׂ�0��ɾӐ�Z7�T���6�r6��q�������T��;����� #�:���<��kg���vM�������3��r�ɂ��ѓj�3�K'��u	�w�{�k�r�V�f�L�)���%1�vh���oBz��i\[EM��k��^�ͷ:�Z��{Mŷ��j
�S�ɸ̉�P��<s����5��"w���������D����ڣ�����z#u���bK1�h��Is"WH@a�)�S f�8��9B�{����Ӟd�6E������ _��bf�Ԧ{���7	o��\����ho1�'���n�IU:qt)�)$�&���w�1���@J ��4953���!&�Y�9�e��`��ِ����-��~��J�H̅�
� ���10��c�H��ζ��iE�EIG�n�uG�D�L�RF�o�=��4k�r���*t�e���ZFR��;�md`Ⱥ�O3J��%�42�dd�����'x&S׳&�q�f�bs�n�7j��s�����p�ϋ��@u�p'g�5�F��'��M~-c�z�%��ޮ0֊W+ ��.[1���8�����Y�`I�qFͨ���j�s���:�qv�g��CYhU���F�i�fwٶ`�ez����n��<��k 	�,�w�rYuJ8CI�����Ky�ՂWD�>. zSO�5�Q��{0u�eQ��3���@ ��k��=-�	�`@ҷ�����!�D1Ip:�%=���"�l�������"ծ���TE`���a{%��;./��=�)���ïm��a(��n˹�S;�y�9��zH[;|�dj��GL���8�<�nʺ�A��P���|&�%{��� �C�C�6���@"h6������(�t���ӣ)��BQH:ػx�di\��!�Ż��g՜���VP��B��-��I]Mj�sC�����Ah���d����LHE��&����f�,��/�zc���7v��$<GF� ��B˔���-��??j�XX歬�|��NUR��k�X@�F��en*�(���^+#j�%$>�(�WNաw/u���P��!�&�Q�~E�S�,s�q�Wa60�
�|-�&t8�q:h�%V A�%�> ^�)���3H��pρ�,\�iQYh/[:a��t�O��C�}��=f��3
�C!�f���O>p�辚�պ�k#�%>U�	�3( 8vC��,�_f�k�jk.n�֦#��s#x��P�p��`�V������������<s���3���1	�Vj��O��4t@�)��OGzN�3L��|�Ļ|b�d �ܿ~z�P�3��Q��������E�$��9����c�o!�V#�[�"n���թ�l��Y�(�Z�,�H;�*h��k��U����ZqF����,?0#8�W��?�:*��Pή��Y@��E���D�9�-(A��Zr�D�Q���(�<Sҫ�%KD�\MG�I�$�	]�0w�; ��Y1=*�Z�F`z⤶ ��Q�#������٠ lLr�f�����"+�@�V a��)��R�����	n;h��}`���֛�f�J�C���W��e teM�|�I�ʻW����X?�#�b^&$F�`��I�u�Y�RŤ��R�O�*��䓥�������rH�.ͼ����33/=�J�l��33$���1�fI�u�7���	ê|<b;l��u���x�<("c��i�td�t/m�I�o�"H;�#�d_�jd���{�}���"�~�mGh�����E	-��X@O~�D>�1Xx��a�\�ū:R��n��<P"ܼ�34k�?rp�Ҷ4^&Zۊ�|�9`�Ky�=�SǶ�����*ۅK�,����ɶ>�_
�5�5f���a�b���xjI�\��l �%��F�P��@��zk�������a��U:�ľ�s���� n9G<�F�.�)�6����SZ��ݿc��z�*(�]���ʠCP�O,��`����]��-8�fΛc&O�O\�ԏ^���xt� }�?����֨�$�LXC$�|�����0��t��-�K�5�Ԣ���.�����N���z��<��Řq]gVzR�y�͚B4���؂��8J�|���ݸ�S�ڰ�r޴�j�ց8{�� �HƬ��/��JM�DH�#Z�2�(U�RG�N��Ū7�	_�=�Ed���cRx�{'�*|���mul*���t�VᡯYG�0��2|J��uK�����ñ}���aėDy�~�KfI��"a,�E�O�媣Y?D0j?w2�d[q_���y�VN	jg�!|��㊫�q3�jP��;�z��R$T�O��y�Q�N�G!���v?_m���نc�Ę�z&!���3Չ}s�of� �V�R�lw�
�n�t`��W��=�H6���}�2��)�|*�{\?�(�5Hq��r�T}���;���#&Ǹ�&���K���i�=�NBi��j�i�i'��d�������}�e8�UY�����z[��FZ\��c������\sj���X%`q�Z��+&,Ԧ���6�D����%ڔa���{�v�8#ޮ�keIqϘ�K�$딙��8�1w�i�u�"�T|`�k�X#��)�E ��,� roh��>�r��4�]��*9g��s[q|p�,�j�=�� ���z�����Ų�N�a�bL�O��[��9T��
:�}�7��Vm+.��y�?2���c��A�Ͼc��(Pot���]��P7ʽ!�~�vE����_���Z�6�����$�Z_�ym�����p���>�#_�4�i�z��8��u����4�����"ȴ�Z?����cG�j5���а�Ym��y�)@�B890��(�H	*�qf�Vԫ^�l9���pn�,;��EQzi��mp����[i%��P��RWK$��aG	V+!k��P>fIN���'v�:�Q��'^L��$�����  eߡc���~i���e�q��e�w�R�DᲡ�XJ��Sq?�gB�j}�OB��s.������ğTX��Nw�y!�����k�ݰ3,2�"WV�X�@M;���qF���گ������{��V��H��¯����cZQ�� ��J:`Ӟa޺�ԲGg�=��)�r�k|�38z�]�ꤶe�엒/>+��(����-�^R�� +�(��63��]HSh~�)8BA��=<�	�UA ��Ri݀�i�x�	Θgk�{䯖�)�q��_#k��\��*ۡ��C34�#�r!�]z��%� ר�
L����D57�G�i�Q��r<�Ċ	�@ R��X}�
\Ĩ7���{(}��,i��lgф�DT�%�0L��ޠB�]8�gnŤ}%Պ����s��k"]F'M�[m�#��gR�v[���,�~H��-ZU\}��P��V (�@����u��^�6������`�ߘ��),W�&�7��5�5�������Og*<�#?�6JA��E�uQ*B���)V=�Z���ϟE�#-P��m��hm�m&30��{��9���:�Xt�$8���8A�PH�Y`�Wr���k��iZ�vZ��m%�oͪ��ZP�\Fxe���%S�Z�+I�������j�I����ǻ�\�d��퀡d΅�{��r��#d����oԔm�4���7�kfz�(��
./VN�,��qw�� ,!�B ��6���ne�a2.��e����C��X^l�8�.�4��ǹV�n�� L#V�w�- �(���UAX<��� �*�iëv.��K�Hȁ��["�,K!���O���T�!0X;^�,�'��H��ܬ�~�.��G����4�[6rL,%S�Y�����!�6*D#䎖8��)`���sa�+i!��節�����[�����mѻ��7��)1t��I޷_��X�g��a�#Pas�0����@���	Dd�d`��C�t���X�������R��o����@��"Y16�(	$>d#��{�$�#�i�$�Bo@Q���@��^k;Ș��HǢ�i)RČ��W�f��u��!��M�~��=� ���0�!���3�{���)ۉRB�(+(�7g��\�mN܉�&�%3�O$ɹ�LtC����=q������t�����>Ӷ^Mµ�v�6�K}�3�����s��� Aϯe��	�e�c�֩�	N %H�Q�q	��~��օB�pn�����J��;}���;�(��#������ �3��%;� �H)��\�ܸ1��u�"3����`$0ͥ	�`��y�*fY�\~��ݲ1���wʂ�M𸆏*M>U��F�
��*po1��
��/��DczR���)�٨i?S���F�ި�n���ah��]�ڼ�����h*��=�ƹ��o5��a�*3�cx�.�aʸ��Tۜ�̮��\��(k$X8���;��B�3��3A�;�Cv��T��D�4<�ק8�pow�&�x��xP�T,�O���M��"d����b�E�.60B�>�"��g	T��V@�o�E�aD71n��,��-�KU�CU(�	�\I����?p�ӏ0$?��ƾ��b���<�P$���2�3A8& �m���������] ������^��0GT��L"&�p��.�%ΘN��s�E%��%��oî&`k����r��>��q����Pp7R紑���f��j1M��^m��/��LqY���x|� ����z]Vі* p�?O�%�	XT�$z�i��ӱ�o>��}N�(���U�ؿ�p�C_ �q�8�U�^��dۙ@x��t��JJ��̻x��4�),Ah��'�Cv&#{�T]�0G�8i�S7ӏo���s%�NRu,��z�q�_N�𪦂̀~ �*r����E�pWD.L2���JY���~����/���}��U�w�%�=�sD�2{.��1*���?{�ײAF�1×��>5��9?�����E�T�Rk�B��3y���4��6㓫:�5M4�c�r�`nÖ����ڳ��H��sy���Fͫ��4}���GD��[�O���"4���	�7|^��T��a�����n%9���]����+Y$O��Zp)�R{��%�o/�������� ��/�W�d�����&�Q��G����X�IY�y�Ka��d���tlH=07L&�6��]�-QT����o�)Χ�MvM��in�-��q2�[��]��+��s���p�s�� �,�Aa��'��Q#�9����Nҿ����9�7����G�HyT��	$��x����X��1Hn�its-c��UÂ3����yX,s���,��m��eg�Ki�V�c��q����1qddc��A�$�MSZW��|�&����V��2�p`,1԰���CЮ�;�p�R�8�͔��9�k�����W�r�#��"u/&���Qk��o�t�jڐ��>�B�1N����~�*Ҟ��$ZGY��֢�����0�ٲ�n�cvU���9��E�x�I�@��,�46��3�kz��z��2-��)f�t�����nY�u��ѯ��¯�e���Y=Y�j��t�^�C��:��l�Ym��݂P�OB~�� �뫧���.�+R�U����9+a�U�?}	�����}"h��06�M�ܽ��q���QDzf���"�5�?� ���p����sp�L#�@0���:���XK��a���c3J���Ne����d.K8����ݗ��|e3�r�]�OdK<�6��q������:��[��稪��}[.v?�9u����A!�!�P$�G�l/:Om��Bn"^��w��lA(b��px~��? *��mUڐJ�uY�%3�Ng���@;��&g����'����d9����h��Ӗ�ݿ� ��(�ƇOM�mb	�!����,�=6�P�R�ZJ�eyQ%� �lB;l[}�_J p���a>��+Qk%B*)���$���*7T&V��<>qd�r��$X��Bł�����nYy�f�-͊��0�%����Ezg�Z��m�+���V�ք �އ+�z|M�0���k��̦m Pk���:Q�yB���_A��^���ҳn�y��������D���Y\�������0Of�� �e���.SU�6��"�vB�2���5��o꿂5p������,��*��3L<�*��1�~{)�$r��ROlO;C�Y�$t��4��Y�L�t�`M���<�H�G�UTr1���-x�7�-ۆ�@���bZ�}t����DK��;0���:�S��H�K��iK��4��E]�o�F4�.�R@_���=�s��Bx�>~ڗ��n�k��zM��ǳ/��������.Oz%���<gZ۾�#�ޞ���@�7��T5cW�]�m�1����%
�&7�#��O�q��@X�()��Ё�ep(�T��5���C�!����ު����Cȃń@Ͽ�0�x���$@s-n<�qK�bI�2$z$����i,Yk�pןha���z�"ya��p���wr&�˓��d%�l�ɵ%�A�k�Zs`���=M���s�Cm�}��ݏ�z��lj�'��0��+sY����	nG�ED�Jfs~,�p^���)�0�.��;Lŗ�b��Ό̟p�GP1s'�F���#�W���
��k��=�cV�HE_�c6�[�c?B��/ܷN��R�ܝ�b�/���`�2R3�5��jN)X�8	��.v���C��!�.sx.�ܸa<2�� �Jږ6� �U*���,�հ����kC=�V� �"��H�w"��7X����*
��IP�q<�1p�.z'+{K&�ic�=W,`q2̛��\Qh�G���Hz�<=W��D8����*3��a����U�g�IG`�3�GŮNEŬL�����Y���I�Guӹe��4�u��ޙ���2t��AC{�F3 ��R^��.�vD�gh���/ ��ڀ2 !�4YA;W 6�Y]���}�]������Ԭ�Glq�3dH��i+�P���9F��i�|ȏ����D��L���b��Ȫ#�uL�QH��ڠM�jqŵ�uk�h�}��F��d +��`�<�M�&KB��U���#ӳ���P��G+�^���t�8�E\2�Y]�PYTڞkI�c6�g*sl`���_�e�o�=�+v(��r�*m����wOٞ�wS�|T��1��O�n^H���|oĠ˓i��wx��U�����H�ct��&��`��l$?ˏ���m��6������ҀQG:�@!b�	��faފF$�d�E�8��?���i�:�4�^C�0��j�-RK����}Z``��F%(��޳T�XUhǔsGa��+���o����!Nt�o%���3�ȴ����x��4V��<挰.��Q���Q��O�(�6��C`��3sa����#�r�j�"XQt;�(���޸�0�g(�\Z xF��;]w�Dj�٭)���ѦeW��K�P@��?=��%Eގk�T�-$�hұ�,*qafK��#	�c��$���#�������LvH�[g[���e�jI"e��t�����d�t�I��W<e���k/V]5���ZH؟:�E�d}�yNTz����|
�¶T�ٌ���Ⱦ�m?�m��,+f�2M�]��jZ���M�pK��)p����I���2t���[8��/'�1�ly��$�.H���UH��c��E�:�1������<c��p�̱6�T�H(yw�w���m�sje��Rp��x����D?��τw�
�[v�C#3:04�f4��E����@|����G����f �Y�{�(|m��"��>#6Tu4_���|'���W�;G��Ų�J�8zW���9O�W�""^Ԙ��c�%<�$۽���ե\6��O�F�/�ߩP��}��F�h������x+����@p,���G�i��OרNOD���\���:-�c��a`�8��.�~tf��<0�A��(�{��i�B�%7"_�Y�:�0�Fukq�Z���I5�q����l��M�E�3o��(�������"Z��ר�E�kD��?�`�Vjc���4%��(fE&+=�;�qGuޛ"�-4������4���;!��ޑp�1ꄶH��I  �.�n��?l�p6��q�=kyk�_�Op��Nm�,�]�{X��f� ���Ek��4W?�	��L���p�cW�\Dp�C?�4=�X����KCrLيgh��t���IHO�yBe]]ޯN�����<���V�D磙�6WJ��^��;��6#V���1-�܍���x���U�~rw6��.z�@V�L�͝cb�^Mq("����%�|�s<K��z�-��w�x8ƋU5.��U��g���6�}����� �B���'g�|yOص
ew�- �5QZW��c�jD7�:���E�����k娻!c��*t�Y�{���$zƱ<Ǵ �D��^�P�'~#:=�t]iM �Z�z��^��fG������_�5ޜ�;r$���@�Y��>�Q��M�?f�R�]��[��$��wx8*��Z;e�� 8:Q�<��B��|Ǘ�m����hX�Γ����N��ɶ��ΟopM:�\`��k�|���l�M��6ސD���ԇP��hUV�w�G�����^d���W��d�Ϙ����톡E�oO9�J#���P���|5�,Ki�94KM֠;����[�k�.�x�E�%'�>�i)SU�4W��va��_[lm-��"�Du�׺� ������r�Q�P�FYOج�d�� ���h$�/m��l*�ʌ�2K���b��0���6ݘR6���?�K��d������ž����6)J��O�t�����k�D�՚#�'pgh��� s��!ս`�W��`u�����u�B'��ϧ�&����&�!w$�Q�N[o�Ϛk������i��
�H��F�ؖ*5�@\w����'[g���7q���V��]�e�V	� �D-��E�HK�4i�C�Yx��j��B��n�{?j#�Z���xQ\a��o�H%�xl/��O�ǹ���e�mz���# �a@A����>q�rX��@iX��{�t�r6E�N�]wTFL�Qg��V�[rn��^�b���7a�C*�g��bl�v"CC#k�Ԯ��k��-Y�����CI~w~����}�ĠŖ�Z;_�A�7�!fU��R<R[��� �U���ϴ^[3]a2��9�g�6b[2�݄6^|<�3�vX�� ����U.�v�����P!�k�{�D^��:�:�!=&��&#Ƽ��B!g)LAC�z\����=��6�+\Q�tsN>k��tcr�(tbi�a���d�����yOx��V7��1
�����s����-8����Z�BVt��znĩ�Kş��GSK�Z�2T�)��r���9�-T��ukϫ�p��f(��ϩ���ԓ��A4I�v"\?�o��waP*߸��VQ�o;f��l�L?=t����!��d˄�X�� �ٷK���
��zeJ��Px�)��*s�#����7T<1�7ɤ0
C��ϊ��5ށ��rE98�n�7��ԉQ��qa�$����l���5i6q�J��V��>(HO�ԫg��� aw�i��e�ڎ�,7�P�F���������𶸁�����H�o�Ѕ����F����^��@yT��O$ �u��z���+�3�ñy�A�����;�;�Ŷ����[mh-����{Y�g�����]~�����be��^�.*�����
6ݚx��II�������'�wA@�p��A�ŮY����a�y0���ƥ[��F3m.�r��n�3�*�ݸO����s�y�����-$"��PM�?=ݍw�l4 �.Z�h	�P�}/ �A��P �k�b��H��F�q����+A�=?D˖�%rm���J��rqv������[>p2�fj�!��B�wo�]I]�H� ��I�;.meٺWh(�;Y�CJ��h��Uʷh����鍇SF�}��P\��j����`�/��]�	!֛K��z� �����do#���N 6&X"���ۘ�G5�tl���A��$0�'�$���A|���K�.ٛ�T�_�a��8������F�i�kd�#�[��x3��[X�L�̯���Q�+}o8 ��(��hm�j�!(f�2���}���b��>ػ�I��Ɣ��A�j��uӈ��7*�7�̱W������7-·��ZEMX���?t�9�O�ݥ��'�]UMթ��Q���� �0@�Jk�y���[=AC=?E��'Z)پHhP��֭uR������wT�d��y��	(n�A�����֑����'2�& �^�ŝݤ���.E}"�qo�ʻ�EDIqb�.����mZb�檮A4$hD���$v��� ���܌�����YD(�V���Cˡ�m���ŷ�_�d��[6}͋��X��@�L�=1;P�VOy�d����_��#ms�o���x	�䗞N�&��8��Au�h\%�R��s���ͬ�*,��O�y7����rl�V�9�	��ۊ_�`wBc����!	X����6>��m�0+V� ���x�Nk�p��7QҜ��y�����,*�'ɯl��YM��Έ�ՖŚ��(�e'h#]&��[��ޔ͎�2� ���a���b�� �GAq�&�Xd��t�)CjQ�����E�-6��x�c[�=�f����ۊp�p�N���ď7UDm�ل�{]U��lJjT��c��v]U@-�wOC�0���w�������xj�fFY�z���\�P�~7�u*��)*\���.�:�9ؘ7F(�9aw8b���KY��R�9� 6&lc8w��׆e5e7�N�
N!O"nT��谔i����o݅��h3��G
��"=�I�-Zʲ,����U��+μ�<���l��u�ó&�99�ߣ�ճ"��KQ�&�h��*S#�i�g���yNE5<�������հM��f��b�=>���k��<�-�$�3�Lф�	�P\��j/&%��o(k��6���r(�0E�p�u�H�>�� �aJCcY�{���t�����ǚ����d\�$}�&�%��`g�\W'��D�#f+@�ڿ��%ٱ8� ��~N�СȆ���9�B�YX�py���N=���B�w ��ɤJu�[5,��p^�;c�L<��BɅ�8.����:��CC��)u�k��t/i����!���P�)&,��aif�*����],Ħ�ŏF�F�V�z|7�MhL�bV���~�(ï���rd�M)/���S\2���[�s�I���6���^r�ڳSR͙�*�����aj�BUN�$ ��J��?#s�D�U�;�x����͎(9���E0���2�'ES����>�s;7���2�-1  �BY���F��.h1�K9���R%��~-ݨj��V�&�E�(��eڈ�����{?ZQ/�������ib��<��}%#Js�v�0�+�ȷ�=�൤_��5�F�� �.�m�Ē@����^��		���^`��G�����*qH�Z�ގ#Ժ锋�3��M�]y��q_*C�9no��f9E\�t�$�7���
�����J��r/>\���3�A{�L��F�����rc5�f����u���ޞҠ��5���H����'�X����<���H��*Z���E��!��:~+��N�4�[.S�u��<N�;��X5o�BCk�_�Tk��X����
�t�@� ���8[�z��#�s}��IA.����}�уg����~��?׮��/�����L��Y����K*�hR����.��o��Ap��w���
���s��~I�Kg�C����:�Z<c�G�s�C�.�(c��"֣>�:Y�:f ;\:�.��t܁������J��&Xd`x�º04��$���e撴9I- "Q��αfo?|c�s����_C(�Q
Z��.�!���mT�9��Z�_�x��2I�'�ϛf��>��B`�����ͅ��Un[��5zq�1�Ps �����,���g�5m
R��T��O3�����q�~�b��gQ�	:��J�(?�wEo�����Zy�h�#�!=�%���p=�¬Q0�o#b#(�;&���q��~x���g��u��ߣ��k���ҊQ!-��=�����6�A�>��3m����-�6�3���c>4A���v@�=^%�1V�67������)z�A����2��^J���t3 ����#���{�h3;��Th�w��Gu>�Y���C�iT�(�b���z,����r}HZ]F����k��
'���BX{m�M��"��է$6�&uȿU���	��ċ�p��;��G��;��޸�D v�n|h���EŒx��J\�<M�7i4���w��O�@���=J
���|����:���
pKb�H|y �j�t��N�NɑI�M.`|oN����C����tIwć��#�o�7�O���j#����S��K�4y�ad�&9o%H�'��\�ef������lc��z�bC��`�G1 s�C����A�η�Pe����_� Ԡ��k�����9�9��h*lJ����^�ϐ8,�	� M,ϊ�&�Q �����,]����F�87����ߣ�u����5X lfY���ɱ�����._�b������I\�ӊ/ �"d�Ӣ�s��2��!F߮5��$*v��|R�Q�ڿ�;զ��g1a�e�Sy��Lx�\pͩYe�騢S����	~�0���B�p)��Q�D�E����XDBF^�z�|"o҇�>x��Ь�������(��&�J��}�Y��{$�$���G�O�޾�f��N���M��������%���`��r�Q�����M��%B{j��lo�#�`�X�&=�Dۉ�����j���9?����Yj1ŉ�H{�
؊��9��=]�ٸ�S1�{y�d�}�/���2��������I<ds�2�pVҍ�E2yZ6��(���R���K��H�I΍i> ���#m-��GFo�#@�rj	j��r��2x�X�˼���K�Z��xX��MnuL�-�&M�k�G����*"��lN�rډ�C���\w�����+��&W6(uE�14��gѩkSj��}��-j(2CP��M�7�C2��D��@a~�?�>S�ٮ�\��X�!�j�$a�8�锤C�3���Uc�h� ��л`���A�������;�	��9�
s���Qϰ�~�%Ɛ��7A֢�'�E�N_��;�ʝYʹI^B��E�g��1�r<M��d8>�:\("����%k�c���A'�`�7BR��~�k6� e�>��\A�K?:iŸ[��%�a��xE��̤��d'��e$À.�k��R��]8������� �f540���� �Fp�̖�D��S����pL�Q�'3���ؚ�GT��,2F1	������m3�X�ė�i���0��m�BAW��.���(�ZcЍ�uW"�R>��_ԝ�6[�̬�z�R�>��D;�B�Q�|@�.�n��d�"�cd��GȀ��|Y�����w���<���H�eg�a�(Q:�����c�m�kj�y��� � �5di1�6	��7�Ћ�e�T�7O,����jί�8"�F`R˚��&�+��Y���ƴ���>bc��I�X]�#nR��ɳvD���j�4w�?J5�n4{�hA���w#`�x	4.%��X:Ď��_$*�h�ظ$�3�R�>/����`�1aPw�K�鲵yw�Y��i�9���{�/p8�YP�
sW����]e�a����9�
�G���K��YI\l=e�֐��0�^���[Db|BsɹД��s���.#0w�Kf�B1-�n� h���2d��Z
V��Y�m&��gpEJ�i�z�
hL���f; w�ch(ߍҥ1�̿pz�/J�K�ƾe��2dg��\������\�ڧ���ȿ�<��PƿT�w��m�%��W��R������c`���	8oR;��;]�l��G5.�PF� �$ٻ)d�v�5�vz��dT�v��k�z��>��/�Y�nW���'È���C� �@&9+�����rI�-%?��OP�E���}[b���@C0�
�o%~7�3J�]E�%τ�Nv�4���z`t�ʴ���34�㲇+pqs��X�`#�v[�1H��ޒ_�AL��t�� j���vn��उXE-N��c�����p�v�
'�����B7��w��T���~�Zp�g����ч~ev)����u#�c����!��_څ��j�0$�}SF���+��fz���Gك�27���z�ioo��������u�����Ќq�wˉ]"ϻZc�ŉ�<�,��T�$H[��i��Lĳm�CĨ�Z�H�/E^�+h�b(�9�A��Iq���<������/�� x�毹��MX?�%G<w���װ�Sl�I{I��nT-H��VC�e!�B�~�|-,�V�>�3�޻8�)@��(�����u�qLr�wٱ��h4��M��NgC�t��c�?l���WY�+����M�&�&.Pi��G���V�~�7��ο�I��G�����1����qX��19�Z���hVU��͝�d�>��c�/Iv	d��7��ǿ?�s���q��>e�����\������~R����D�ы��7X\Y��69��;^b��XT֑��5֌����:!�@Y��R#TkiԊ$ڗ;�UǄZ/�Z��=��Q�u�>Ő0~�E�(��H��T	o:9�ތ���kg���w���du�0���Z��B zZ=�b(�N��
����l����aE�����es��7�� F#T'9���ySt�{;L�e��Av��]2K��S>;�w�Uv$�u�6P#4����ޛS�OI�a�!
=��Sڦ��n�ـ�/��92�6����V���/8�Q�`�]0��[ᮈ�SB�uݖd�~�R-���V^/��M I���>/�3TN!�Q�<S�o0� Y�H��l	.q.���0�f��ݯwo�
q��o:]`4�T�z�7�w�W ��ԉ�ͣ�3h�f=k�0K�	��5t�Gx����:��X�ѹ�bm����hT_�Ǯ!� ���� -��u⼆�++��dԌ��5vh#~���w�P-�9����c��Æ�DUtC�+S�ؙ�������9�Vt��$��趡����ؗ,�(�h�X�C��{�Ut0B3o�P���"A�eh@��X�b�Yl�C�����P@���Q�^��;9��y�����䋬�����������ȍ�S)&��(Mh/���!e��m8�"��	�s��۔�/����U<=A�4\����&�vxs�1��8E���s��#h!�?E6D8��R�n��P̺�A+I��R[Qߵ(ʛߑ����T�����S��G�ݟ��}�}���-���s���^OD��)�
�,��U��7�2�B���X� F�Y��yY�=�O�0D=�	�#�� eTҔ	�~כ�2Ѿ�B��� _rI�$�6cb<$E3՟K�?���J�I�<7�Yx[���L+X@D�7x����hƸqU6	�}FuA���a�`�iGL,я�ոQ��_�y<���}��=~yrw��>��}� &�yxgAN�gpKV�8|�L�p��=o��T\��"���f���G�E.S��ߓ�k��u�~�6��m������d��qO&���s$�Z�W�D(ŝ��Q�1q�m��c�)��`쮝�B�=�`�W��dY`<ڪa��"��AO�a��$s����x�V�G�$Ę���ޗ��Cm�s��>%*�YѮ�T�#���zp��^�L�t!�Gg�
T
)�`���l��	I���JZ.�N_7�Q�m�&�k_z�/\��t�#����x8�ک��$��5"J/�C�;)�9+�,|�Xjgc��(�;XH?B7.涟2�}Ԃ�.x�T;{r��6Kd�W) �y�L>up�l��X�c�Mk�yEj-��f���>����Qd��kZ�����K�Q5�l��pA�����WU�X�5�?��䯯�>��O�RB��"�̌�3�ڝ�1K��~�5Ze�#D�g8��DS9
�OSq�}� }�d�JO����8�e��Ǳ����¸^�����A`vu���jaIX�l��43م��x�p��H�3��rg�3)���3�R�w�ds	� �$r��6��g�N�"`�c5�B0���c��(7ܘ�,�0�#�5q������l�<hRr�}T�e��fL�Xi��ѕ�$��oG���?�`�ǽm�+Dbю��T�"�T �ʉ	#i����}p^u6�x��O�"�V\�*��t�
��x��Y1��8ʼ]V�����=�$W0LgY�$O����)�u�1��'عl�0�J�Tױ�=ܺ�h��h�p=n]����;�bW+�2*x�)�"�����5%	�NY�( `f��p^S�ǶR�PL����).A�.ؐ�ҕ��o���%:�G���A�P�q]U]N`q�}����Js`a�U�$�L& |�[�ڳ��r¥�m���_��l�;���c6(&�#�$V��Ɛ,���ڸp�ֿ��Е�A���5���PamQ���N�9�.�\�6�_�h+��Z=k�YQ܃�vyj U"�:v�������I������q��t>�;6�4���}n=��,K�p�ŕjp$Ӌ����fC0P��L�����;���V���ψ���T��g����6��Z��#J�?�9z���2����6k�sb�@�
�y���̐!ݰ�}]���%8V*]��7	�R9��XhZv���G�q��w��Cp�C$u��D� V�������~��{m�Qc�V��4�?����q��Ie�Dd׮��ܽJ���&���5���p`�>��,)�@�6yN@�}5���ʉƶ�۷��-CJj���ʴ�i)�BjsAE��Te�;�W�n�l	_5�z�2K@�D�.K1v��{�a�_�q����7뾶}��\2�y�J|!��)�����#JJ��.�Z�ÄB*h�_��t��'\�-�UC"W�_sE^��ƅ\x������'�w�:��cY�ʏ;T���� ���!V'���Z���Y�fq��	iD��[g5�ʬDVt2hi��-snUf��.�����N���y��'���m� p$�9���}4`A'����� 4�l�V��"-]��7=���!��ѓ��
o\�q#�6(���dA� EJ���͐���?����D�����΅P�o�ra�ᅂN�1��3+���H̱�y�O쑞.=^�������U��
��rC�)��8�ȷ��P  �D9S?��'a䝘�-�����Li�1��}�h�~ǫ�D�'���ԗ��yx��o2�3�4��!���|D��m,i����jy�~�e�̒������GT�`���O�RQwo���ډ[��d����1���8����ϟ��Dj��8X�.���dW���cY��.�;��11=U��iÍ��9Q�fI]�r�}�S�����5k�]W�̚?�`��A���^1\�0A�b��;�,g�ն�Spއs� ܹ��k���ײ����HnY7���R�Mz���w*�CG%�J)Fն1~����޻PE1��=o����Zn2�6���[7�B�1����p����W~oO$l=V'��?�������T]�+�9���')�ᇱe��~=P�L��b�����)��)L���ήljB����OXH�W��F�{i����BS4��ag�����|\2���'����if�N���ł�8ت\��j�_�:&�b��ψ �u�M�|��[4~��ӿ�:B�l�z���O�~�g���?D�_
Mq4r�i�7d�ce�P�&�C�'�QĈ�8gdMS��˔0�JK0f�Μ�_o���Q���^��x�ہȁ��T\�&�LM���Ƿ�E6ȓ��c!~���0�wMʙ0p)�xn��Y\��Ȗ���~D���<�$�,�q�gz�4���&֣oe]�Y�8>��!�����=�t���#�������bh�e!�<n*��u�[�1�na�Ӕ1� ݹ��v�GԬ`,���.���N�{m�$���:`����=i(�T�Hg�2�g�����+g���~��cn�����p�X`�du*��'�2����1�x�_��z�:U��<zf<*=��%��4)�ä�j|�J.�c�YOIx��_aJ�%u��B9�ۣ�<�*4�l�G�>*ت��v�\Q������hػ'jT!9��\*�O��`���ȮnI>,I$Zzy ����dy.j�N��('�i���(��;sY8c�9��8Fă߫�3�Zs�<�*X}2�H�b4���}��h��G���xi`aI猝�>��3�n��7$r��ǒ�U����{�9-�]��S����B��㿛�ʫ~Q��n6��8F��̶%-��^tr|7�� ��q@C3�i/�O��V�F��;��� �w��jA���RU/cu@��>�H$˴E���)2�����a)������/�p��UF%V�ը~l;I��f�O�v�m	I�M���Ab�"E�5Ƌf_��ܒ�5�s��F��M��i���f� ZVJ�n�v'c�Q�'�ό���	Aп�l�a�5U��v�����#&��*,���?�vD�
ٵt��M��x�]ǈ�/G;�{ f�a��+�#6���Z��n�y?�B[��+Zz�z��{����a�+�	���2�-�j��p�r��٪fȶ�8@9ۭ�CD^#��q 72�('&|��0#���פH!��re6��R[F�ݞ}����ҽǾ��\_�J�v�|q��:�;���8L�صF�EK�H-�P�W�TL>�;d�!�+�A��1a��&q�݊kX�U�
�ǝ⥐��@8|�g��3+�ޫ�nު�������h-���<���0d�(WYY�]4H�Dg�����ʮ%�v湂�GO�����g��i��������ţC�;�p�U��4�CvA4�k���ү��O��)}��;4��B�fu�KxwR�Z�[��8;N�-;2����O��t�jbz���Fj���R'�dŹ���k��0�~�9�`�Nx̒H�f��lq
�በ[5*3���ٙQ���{h>���4��恕U�S&YJ��b���lUԩ�n�h�s���sN�ąa�Q�xcT���Y�6
') <$�n]�T�ɤ��*,�8��0�u�ĭ�)�"�?f����(^�D�ƾy� �2,�|�I�n�ޏ���Q���#7�䤴;%��(�������^Kݾ;9�]�� �����_�;��NV3���SN�~ �:k:f��ٜ3��$�tB�5~]��0dS��>V6�#�6.ׅ��*^2a��FFu<��+ u*�P��YOL�;A���m�W�P�o�auf�G;@e�T�/t���U��Y�x�/�X���[�g���٢��n�u�F�u` (�Xh29K��<d��'���OJ@�Aa\h���Ɏ��њ�;rHVx'��ѧ�B��c���_z��JO�~wuѮ�e�d�Vn�=�Х���n��:[��c�h�7�Ug�������O����Ѕۿ
`�9�3�UM`�(�_�WL��+���ふ:�݊�7�/1!K����^��N?*���or�Q�އs4�t��X�_��#�]w���#��V)�!�]�I`]����Q�*�Q���L&��>h�Z�ܢG�-͍n���?,]��H?���+ه��a����n�n�Q���\�[ �޳��a^C+k�W^��.t�QX���RQ�B�zcNv�s��)t����	�~��0�l��ӓϠ���(PL�a�x��yI�V��'����uc���K�T�F����Ǣ����.L�E_�B��(򐆦Z,i�bM�A<����R����O�/�
6��`K��ܞ���-���[j�$��;��|I����s�"��Q�]��|���1當�v!'�P�92"}�F�-?,{f��XS�)7�'�p��q3����ݘ��|mIN�9K�Xٯ^����~�L3�v���&{��b;?hۦ�s�ekT����M[�%h�.@��"{JMu��}t��r���p� i��K[��[c��"�*R������N>�4�;�[]��tJ �ZC��S�������&T㻬?U&j15�=0�(�vrx�����M#*�����xN`Ӧ�m���x\�C��M\���nC�ِc�.�ˋܕB�N�{ʙ6�`�n@є=`+�u�m�ʙ�~1����m2,)4���3(ߣd���9"X�S��I���y��pSl��=W�Ok�$��1rro}�)��&k��T0P�����8MF�q�_Ԁ���9�rvs�RU?��v�D}�Pc�l�qd����r�����=qC$�]�p���87gZ�X��m؇�)������%yo�e���L� j�ί犟ł��сE�Uo����r������*�.��͠G�`` %i�(���8�xyQ��-Z�ܪ�oP�)l��T�R��Th����#^WH��f�lGc�I蹕v,����FH��z��g�ҽ���!�$�F�:5ŚI0���pPt
\�BR��f��u��^�A��a�~��v;��I�n�:
p�1AfD���O�w�����1��TSk
��%8���ٴ��[;E���
&���ͭ��[��Q�i���M�
!�֤ZBR#+�f�Ҍ�G��/�R뽈oC�;��nY�[q�"�ԣ>PEd�=�6��Fg�����Lqoj	�>q��ަ�ޕ��=rȥ]⇅�i��bO�~��QiU!GT�c3��`�$��|�]!���+5ƿ{#�'0H�����Uss�c�у��I�W9}+�0�XlSͬ�ϱ��K,�ÆQ���9���%���(tV�Seʄ%�B�W܃��dw��r�݉\M����bA��!P�I{k��z�R ϴ��6�#�Q5�i����xѺIV���R�J?�f#;8�9�7�EXt����Z2\��?��N�p�me-6Nb����#_@婰�1��U�\��
�8.�Y\#n� ]�����T�b�E����f{���Y/zV~�VJ���ޝ�Ȑ.��?[,ON��e���ՐS�/ US&v��`i#V�A��g�&X4e��� 8R���g����9q:��诣��'N�%l���т�C�(��W
f-¸�j ��P=ͤ|:;n�F��~Vm�*����!�K�Z;X���o<�f���>~��]5�F|�&��afY\�粂Dzϳ����n� S��#�Dd���\}�@Ġ��;��يpQ)Z��y{8���"������hO��0����x�/�����L�G��53S�}���M'"�@�l��di�$S�<��x߆{S�����?�z��e�71-\�TP�x���8P�H��*�8i�!Vb1��&t����,m��JyPA��{/��7 P�N���ǫn�p�����!��cd����u,P\ �@P�t��/>\����P��\���"9�[�´FwM�W,*����{N}%Ń���/����C�n[WUdP~bS%gNy���n�a�5����Ϝ��uX��%��R�;F��t���O�����)c��3�fuW�ਙݼ2,��� ��[WAR�kKT%�+��������jaа�A����1�mRoG�7[��Lv�9!�t*U�[.]̲��1J2�Aک�t)w`�||�(e��j�´����o�M�?H$/�q��7$W%i��]Ҙ��(VУH�3p(�㏂�L0"�+=��wo��,�����er��bٛ4ov/9��;�Ǝ�T�I�	���;��'YQ����	$&�N�.���a��Y�{v�_o�1�P�S���24I�Yۃ r��}��\c*�|ihF�I��U�:x7�[{������%�a�^8��qм�N��,���{e���`K��r�*�Zehuّ�����,C��� �`ve�w�{WL����<�Q �q��o�-ږʗ�3eE-+<�kD2��$ O.d�o!A�p䃋�~�7tg<~�kº ����E�L3������	&t�Չl+Mg��ws�/����V+��S9���ޙf�P����O��H���:���Ǵ��2��~j~�KY��"�1~-���tg
���dA�W,'e�N��sܥS�<������$��ma~��N+6�{S{�0��ɼ6���A�K������fX����ך24�����k|Z*�4��8��Y���|�]�E����lP?t��&�z ��q��;�u�ݜ���=�TS>��2Rl,њ��kٝŅĢo��O?yr�dI��T��Y��0$W٪- TX|�q�qA� �l-u)S�ԭIo4�Ş.�#�ǘ�t96���ɼ��y�_wA�eD@���(�B�ib֚Nwn�t�!"f3�8� 
�z�|��q	'.2�X���P#s����×o9��+���s��0`�z
�C|:5A�zR�E��w|n����SJF��\���d2X�e-�d[���׼0U�`�@����|կY`!��T�z�	U�o4�(_�>���g�{b�a���8?��{X:�W �ꍹ;J(˼��J�d7�K��>$,9�g;��|Xsdc�&$�m���q��B�!s/���$�Q�.��䛁I���4w�"������2Lb<�M³Io
b؀)�:�#2�_���#�C�8�6.\�ߨ���e2G�a�-/y�Y]���N��|F�����^8��������%U$�|��������L@���L
�pŎ��x�nid�3_,��������ƃ�D�����Lt�Շ��T-����{,W��g(P���ŷ���v&�%�T��R�JY��;p��!����l���%-�(�'e���F���Nަ��+ږ�7ߦ����	�pe����wp{�G:h�b��-�}���D���H3U{��TO;4�
�U�"sXՔ�����3h-�B��&�=�rZ�瓧���Q�õW�/�"`.����Z��ҙ�4ʻ��hj�����d�[tF�yFͭ�3���!�r7�?��rԍG��A��Aj���N�FP��{Pw]�^t\����������?r����c�����Vy�B���oe�^��V�9�j�n�7-$�c��Ä�u����F �j�o٪�H�2�n��w�>�:��x�e�&�p��fa>�l�bً�%����������~�����I��@��P&'����~��gy)�������u!�m��o����a�^�hz���s����re[���CF�e%yk�(*p���z2��5��h(��E��Hp��T%�V|����3qӑ�z�%�� M[�K��Щ80�T��,����������b�}x_��1�nB����6���,�bk-���.ዄ�``�&�������
?2���p��*�'� m�+�w�MZކ�e� �lş�k�k�|�t~ӺX�F2]�Qmr��9�į.���£���dÁ����b���_q�N�[�F[�8 �%��?�k��Ƹ"j���
"z����܈�%`���������S��(v3���n����,���h�%h�D���5h9�*M		��<,�:A���@l�`D�������$M]$mg��^��1�J����VW5A��y�T�B�a����r�q�����f��[GL���u�#?�}׽i����а��h=�m&)�t;��L~6	�V��` ����K����
tC��0}�¿>m��I{�i�n�Y���� <�ǁ�lAk9x'��B��$v���&r;�C��z|��5^Gf�h�K�1�"�\ٿ��(�찚8�G/7��f�rCK0"L�A���n�ڱ��%,g��x��N8`������4f��E5o
"P���G���`Vo,����Z�]bu�W��͉g_�։"����!�����n����tT�z)�?,[D�sx�!{��.�
����蹱�,�0��;��I��:|���(��k��o����\���&�����웪��t�o�>�:� �uc�����ܠo�wQuV�BN��ǟ����g�r��%˞b�[K�1��n8n�G�03�	O[8ey�*r�.��`�V�zn�����K�V�h����FH;��H�<���B��ߘ�E_"7��2:��x��xW���/}�Ƈd��*5�Vj��k	u��H�����7j�܊ZE{2�4���BC0"�Y݋��q��B�������/v�z�W�Y�8�t�NY��d�8{��Ş���!�� $�����f�A#��A9�IB��
ǘrįs[q�z	���W��@�p]&�P*�82����c;\� �?�Q�����D���$������ʩ{#P���A���Er�O����������Xn�Ca!q��j�X��QR��/�&��l������q�N��x��bވ
�=p�C��K��?[��ho��n�[�����[L>O����A�@�%u��N�*����4��k��(��X�aK`f���A(��/I�M�+8u�v�yg�@w��[٫e+Ez9�06�~׻��i&���َ��2$�&� ��-�Ĳٿ�8�j��*43θx��i��^��齃��a����m	g̣4�j�L9������I�)$��z\qgC���]���e��c�?"�`�R�S� �bJo���η���j�6=�Q.�~��moF��`��(ԑܨo��Գ7�3%���|@iH����;�f*9ץ8I�6!���'��v]�L�r2�͓�p�g��Oۥ�|rAz��N|�t������6_��ߠhP1�((}<��^j�a��:z�H~�2�N�*��v����aΥ-QM]S��?t�w��~��ƫ�b���kO�e��4oP\^`����X��bڷ�X4m
r�R�↔�d 31��4�>!S>Y�>�g�� ?���;(�Z����G�nx4�� f�3���U�0r�k�.Ad�i�{%L(��!]�25;�R��
����u.���C>�3��2�ox��}k��0����ңq��q[d��[���[zAs D�z*���v�D��&E9+�Z�H:�l[��u0V*�W:���(5���DO�?b����Z`�&��H�W53���|S[�5�mc,���H�Y�ύf��3?],�g��� ��|;�@��ޗ�:9����h2J���#'��Q s���aX�,��H���i>��֧�(�	XQz�'��5���`�F� ����}���P�P����*{�i�KT$��P����H`�-G]O�f�&�suiX��Ҋ(V�E4����mKKv걼���dp����l�)8M��\fH�` :�E��� �>8g+�x�����L�ɯ�xbe�X�T�un0,?@���:p���9V�!��)�@���6gЊ�3�1>��/��MdEl}Y���ˏ��jv�V~�%�ֶ6-ƭ�/{���H�S׎Bh�P}@E���g���.�-g5A�jI���u���N�M�)��oh	zO�i��~�Q��sE$�z1�o���W�pb�b���9��7��,��D�Y���xw( ��/d2���̬�`a;���j���f�X�7S�u�Z�!�ߑ��E~��(	��!��T�}�O�й=��E.�n�2�Y6Y�.�Α�]�oc��JD �ˁ3[m�Ӡ�����Iz��m���AdN��[e���z�_��d��@-��}�A<��R�Ȑ�0X��P5��x�H덄x����v|���V�Fi"�'�% !?����������9rz�I�s�T�����UE/�3�po�'1�3[��(�.{�OǞx����!��iYLI��59�����o�\�m*��"�!_�/GDٰ�����k�D��﹎�n�i�����i5����|�5��S��.9��L��7N������F�j-xZI�Fn,p��]���a�/ཀ��(E�� g(�t�` 녴��+��2�=�+HD[(�# �����+A���. �+����D#��i�B��l񚤄RS�#p�3O9F���r=	jD�Ě�"�X�-|�.�ys��]fe�^z��+8�I	�R]X�����毶�W�r�~���Z��'���ٟ�W�=��h����O�����)�0Cฮ��Rƥ-p���Ml�@�~;Fo�1m���!�5+�8sx��H�^T+�Us�M����ΰN��;lZ�|F��v�٭K����`�<#�'�^����\�ƕTQ�&IcG��`>r�B�d�!�Y��`��-m�Yc�E牀[�s�4\��Rg�3 �C����f���ЛG�D�m�TO7�ݱJ��|�ˤ˲^qkYT�xq���3͛448�r:[Mr��Vp#R$��x�>{^	��+8˹N>� �Ͳ򮯯u��Z���5�N�<8yM��M�������%/�ĩ���}!,j�����BꛯP����JOG�@Y�>�J���
�c9|��
L���	�?�7`QL^��Uao��*�z��OQ5L�!13� M�x��=��;�b}�N`\\���>e��w�κ�)����+�*�7�u���x���u�����q�ūm�W���|>��5�E�wHg?��`�4��^�s9� .�k�x
M@����Cπ@OaJ��E�K2hQ�CE��M?4F��� `ˋ�ae� {)̦�����2Yҭ�����R���$��Rn��%á��]��W�S7�j�s�S�h2���@u4����M ��{_�A��L���#���v��wo�]���Y��|����4rk���b)xL��%��>���A0��P뽍!��EOV�T��.;�n��:����o�.�T�韦k��"0.��ԯ��>��7�g(�PP.�D���V#o�؁=Ja�A���|�Z��0��KT�e����s7V�� ���kt~�:vm˹,�2��{�U��W���>��|,6�� z�-&Wp2	��0E# B�W�8q����z;�Q�1D����w�S�L�;X4�\�?�
8����/`h�5hg:ZR�a?D�����˓"�1:h��54�ڻ��E���==�8&�匛0$ˈ1���z ..�o�%7eձ��v���4�ۿ&NɊm.�P�07�f���}�nD�s�cz��BG,��'��u>����L�vbS{�<5c�(�k��ɜWԜ��Q�\l���l�������Y��A@Z�Y��ģB�+��C�Qѭ�h�Q�ˍ�W�y��8�����}/?��Nҧ�{	w�N ^�������$��m� �C��c��J�ٻ.im
���e>'�Zb/��=,�6�X@�Lji�F�	��KKs���5~����3A���^��Ȑ���AǪ�"���^�t	/�DD��" �l�u!r�ס�`��F�,�W�U�ތ�ு,z�Ixw��yf<�3���� r�@��24�׌�L�32k�z���Ƴ��!C."0~�͑'��$�=�j��K+S�(�g��Lſf����Ŕ��t�w�f���aBT:68�N������7��|	�F0+�JjnZ{昶���� �AY���5cf�%��Y��d��'�J�h�r�����Z�]�)Kۣt�$�����IІ[9����;����p=%T�����g6�ϡ��$�l\��Y��n4�c�{$�Q.ev�P����mt}(��J~�`5~��-4����Ft[`�ha��W3/4�:����E��0����E?���u#h^<ꎦq��]3�[��F�۫E��@f���*�N�Rs����Cfx��Q�cp���� Hdm��i��|�fH��S�.Qz/��:	����7�p�N�l^�����-�!� [�I�1�ă��x�h��� �JgR��'/Q����
���m����EM� g�m�Y����t�Y������O�X���8Ё�A��� �`��.ml9=����T��z|e�n�aD �f�h�j�8�/�Z�n��-����bb�����{�_�d�-��-F*�����A����E�y�Z��Tm��!b�(��*�c1L5äoz����{�F܂��z�Xi��  �\��jC�;���m]zs܋ �y}l�(���Jf>�뉀L؁/�B�͎o<���s*�������M�Q�q������~+@�U����)O����\�����@B/���Y˅t��~�dS�d��'>k҄��V���S}y��۱�=�?oeH�f�ؽ�l�����$Ż�mک¯�̇�����i�Gvyl���ċ���뚳6����B����c��M�Jm~R
��P9wOJ|�@��m�����)H�4�ɳ�[��\�ى�V��Z`#��J/jμܺ)|hy¦�\^/�ư��t̻�Ɓ�'1v�T������XӭI\0�f�(�L�-���mv����Y��5X���N���Аgi�r��u�,�s�'�ˎ�)ɛ
%�Y2���7`|X9.��iq��!� GW��y��LQ�}*H#�>�k.��U�}��<�����O�R���/YH��ե�M	���I��	n����	����_�]���]����� �I�� �	�/>b� u�IɻY��p-�`��<4�c��Jk�����an���rZ�s.�)��ZL��d ��"0��ɂ�LIGH����m��+�BT����1֊���=d� D�^���1$����p�]w��m�q&����Դd+����~��C�7]����?'6��-�~�e�Փ��i��h��	��B�����X��!W[��%M���ᨬ�4w���8�iqt'�_�<�k��.�jӫ������E�S/y�_�Oš9%��Iw��݅eJ�����Lr�,�b2�����
�Q��h*[��ti��Hs ���(c*�Jn�K�D��g�&/�x#�Qn�=�oЃ���dL�u$�F:˱Y���WÄ��4��W�[h����� ��<:\�Tɂ�x/��\�x7j��5v��W�KQņNMcͽ���ܽM;��h���3�ʷ�dW΁=]!�z�j����`H�o����HJ]s��?KC�Zo��mߕ.zڔ���C�;��y�`�}�I�G���u1*t1�Sr�K�h��/�=�����vKZ���m%��Ϋ?3҃_�k�����/Aؼ�����^p���µ}U`�ф����ϯ�~�`3��>��m)}]���!��K��^�t��}��d�{���s����~�3m����7�[�*	&�@�����!#��]����k���@|�׎����"?v�gzb�2��E�7�.4�ޭKӇ'�r��F��s���h�˵���_��:E!�s�?G���� �~�jں[��,.N����<;� ����g�|	�pw�m�y�W-���A�K�J�/�	��=��η0��E#z���rs1\�۲8m�v�a�}��v*,�}X�'����Ҋ���K�ݧZl�T�RQc�O�Sl�m��^���t�o6}��~#���Wa'%���VgNzK|�Y�ÿs���m��s���_^�O��A�����dڝ��G��^�Z9n��5V	��¯��`�M���^����p���P~b:{�����O�Y!).�YB;�K��Nɧ�mUhN�1e[���A�x�]@,�u�[,XQ���B�NS(�g�u^��~�PԮ��Zu�V��Ӗ{b
��Ι&�Kx`{���*���{`�1(]�^�Z4��w5=��o{,�K �D�e/�˖��HG�΄E4t�@�7L��S��9Q�g���慡�N���3��k�P�ڳ���t4	\Ho	�{���ϐ�>�Y�%��d�n�0�J�˜Ww	���f��"��]��in����l���u-�@����8�)�.�5��p��~)���� w؈�ޥh|2|�ƁP���<|5��ڕc�q��ۂ9atI�"=��r7�S��+��`��
�E�,��So��l'L;
��A	�����~a�oɛ���Y�O1x�nl��o��rcќ��0,S!�\�S*��
��@]�;��!����y?�A���S�����=��a�jV����s���nI�.��B�#�۸��m��s��c�\� KnZ_+F��� �;�$Xɮ���L"e��=�@�?G!�3�'��X2	�p�4�o��F���)t���Z�h�.��S]N���N�e�Ԛ�����:���&�^a�B�go�Y�^��s��1Q��fU�����Р$�0�T5��U!�v�$=���)���{���Nu�8o�l:���d`)���DR�'Ԑ�}!�FQX�6�\h��Wy$h}t@�CzgV� ��w�Y���?)M��5{��8t����1(���sD�(�U��vܓop7�|Z�l�(�Z�w{fV�݋!��� �/Li���N����.�_�J���q�ƪ��J�5U��� �-\.X�m	1\�ABN����p&��LX��3��	����`"έ:Ԗ\�0Xؑ2�w[X{j[ض�˾���I�|cL��+�����Y��,X�]��b�Q�R�.��)��X\��)�D̰�5ucf*28��.7��?�r�S�E\�L���<D���.ݘh����2�-X�y�w��4��"���I?d�HƠ�����E�����;WQz���Ԥ�w ��E^ �s�2B�iN�_����u��z�^�FG8A4\����F�2���E�h�V����$�aI��s��N�Z3�����$2o�-u鮊��
=�c����b�(	�TaJ�2:װ��~\!	�t��7�a�Lt��6���C`�(��6���j�v��h�	�.����Nrd�Դ��{5��̂�V�C���'`2@k��'°�];����#��_H�����'�aJQ���{��J���&N�ꦷ�B����[���Df�x5��	���u!�����r�}O��zg!���PA�����u���w�z�7)�W�'���H�'d,��)���%{�鸦Yَ��Ǜ����8J�m�D�M|�*��C�(�p1�g����s7�����L��� ��FE'A3v�>ܥ���>�l-��L��E�d���fT�Jp��J�C�vj+�s/&�[���!-m���y�rG�F:M�����*�N��Sv�Н,d������DP3J���I7�ð83����ui��=�B�tJ{Ps�m��GH�F�6a>R�^��:��N Tj\y!e��K�-�g��HPM�͓�j{���Q��g��p�Y��\�3'u�u�{��DoDYht��k����%�F��YNF�fw$�3�_{�r��cy%�:�h08���g��Z(��^*��%q�����Z�~��^J���b4�e�h��$�����F�B�0�D3���[A��Y���N0N̈��Y�gu^��zK��w(��[�Vۃ��!��k�F��nKJm	���'�&n��vA����U�N�US�(����a|1�U�bw��W��3r�e�R�Z���}�:h;e8[&g�>����d׷���'���/�Q�_�3h����ʡv#3��d��$�oU��d�u���D��!����u)޵?Ga�4գO��$oo��q��ҍ���7_ݫo��U��	K��-;m���ѳ ω�x!�UX��n"�H��E�v���e�@��A�{���㒷������@�tܝ�q��O���R��f� �߂�y��G����x;�EF��eP��GM
ʣ��*�gt9�ա�C�@����%ޏ͸B���_U��o��gPz�o�L�-s�cD���� 2�̰�G�r���,49�Gua�k{L�|��0(��0r�N�(��$д�TR�ˊ����l��b�'4��9w��Dϫ�#��)9P�G2.���/I�`28#�x�巖3�?�mzBvԩ+[+�؀|Q;�^���w^+�)Q���8����.Rr��;��pύ�/C0�~���!K,���"N.N%�Kjb��l'�I���}u�$!��K�?�H������궴;����C�b�]�Yk{�(s�GMqJ��1�OG|=�tD:1R]�O'F�Ӧɵ�-ϰ�ӂ_��tz������|W,&������C=�G�[��8h��
wPႳweFk�E�2`#g/�u�oZ�"�YGBޚ,��o����5f�%���U~�D�ぷH���>����kɛ�6J�,J%�J��]y���v�=��h���U�?r_ȅ�٥�:�eq���C���6��C'e�J�_Vi���2e��ږQ'�*���T�˯�#ş�u��x=����mn4��*���"��C4^�q��Jt�dȈZ3Y�b���y���V�P�Ʝ^��'�B'�T斑r�g�m�Ie3���w�.?ʹ{SSW
LXd��_q�ѩ^Y#���ⷅ��hE�6�^�OC�YM6�t���u���(wy��X��M�n �1�N�d�T��>*
�s$��"���T�P��SX��q�������u�������>��� �׾0tL���1w�g^�Q&2r����&/�c�[�'��	$a�}��%#&qm�{�ր�x����D��
����hA�^^�i����I8����������E��-hJv�C�R�#Ѷ�X����>�:����c��f���2;��6�K��j����&�\W���S�m84M�����5K���� 9�{m�2��`1�l���ɸ_B��ݸһ)�򓪂�'�]����ۭ��fvT_���*��y<޸��L G��{�zg�0VxD� �+�R�8����*r���:(��v�oS��#�O'�dóC!1�Fʀ�����@���ܗ� Jw�b�)�!Q�Mj�Z�t�bp����6�ZN��hۦK����|0� �l���Pk�L��G9�F\����*d�4����G�{}Xԭ��Ek�.�TaV�:J��W��(���%�97-��R;:���H/ ʹ��/��M�J��#��8h���M�DuM��;��I����Z��7Y+q������)Yy����/�CX_CP���K/Z�Ô��1�X"���⦔�L��-�Z��cMOq��t���~Z�H)�Bz���WgD���>�����d��}�o7�C�[� X�T(H�����a�|_���s�$z s�+�=����5�z_�^\�	�x�x�R��o&S����k��C�	�kLył�G��&)tg����_�6�{U�t<��0�3�3|���H���^��liR��q�v���n*o��x�R�u��E�VBsZЏJ�5Ъ@�L��j�<r�D����2`�i2����,�噧��i�h~s���P�Rb,>�����^����׺GE��|t���O�y�����tW���v*_)�O"�f��d}��Q��Z�X,z�=�:Bڠǧ��<(��Y��ӈ.�P�j�*V[9>�n�� ��H���av�0��{��{�`��ؿ���4�pp�����?�l�Z�,,RPj νE�9f��G�n<ޞ�;}���<=�� ���Wx_d}工3�pR���/jIӞѕ�,%�'9�dM��:��B�=��؆�E*��u���l�b�̰Bo<�R߽?�"��̕7�ҦNz���@~W�ޡ�6�$(~������z^l������S�|�Ƞ�/6��˭MjF:zJ:�W���K�YT����of���
,~3�ɟ���;�ԓk�Tq��
lЭø��=�,)��!r��{߷\���x<�N��
\o�QX�Vɤ38�;���9,Ncˁ����i��8*�,��V���0B���O���o7J`h��h��*WMe��N::�u��X�'��W]?�����95w�F<�S�k�zyp�]����"��{X���#v�D��e���u�Pz�h���rk�X7�0e�f����3�rC�=����>)a΃I���&gg�΀c D1n����0\�u|?4)�,�GaK	�� 38MMĝ-1�>�r�z��<��xhVb���bF����Hrs��g��T
(��S�^O������(2�@�G��mfje��y%JV5g�1���p�=��L��/
K9ZõbT���]����u�:�b�H��&��[ĕQ�)}�"���Ѽ��o~hp��5ծ���p�K"�v���"+��ܸ��C���Ȼ1��Ÿ�h��ph-[`����m��)�ʘ$Q4c3�`d!�Ʉ��K�Y߉v�<��A�[ӸP�Elt8{����j�c%A���F4u�I��L�L�Ώ����(Z�w��bu�~c����(�Oi�
9� Q%-����V��E�����DjӪ���?�5����Z(�v֚#ޮp	�T~{X`�����V?�
ܡ�MgnQ�f�@�9�K�!��5@��
��}��ѿ#u�>Η��y�����a�W�&��.��$�m����ą�H��Y);���*�N��� ��Q�s\�}l	�l8=�.	��R���@� x-3MO�X:B֥��5w ����B���2��@�%M���s�7Z�j
i@<0��K�5���MU�=�h����-ge�B Bw d��x�7��M����:_W�!�����KW�Ɵ��)5q�w��<�!E��UD!�=
�T>�r�	�fI�5��*tO/T�o��3�1ₙ�$�r�W$�8!x$��֔���E�~E�1�Md�0ζ9X�(_�1N	�<�f����z�~��bi��7ļ���8��3�"a�=/v}��oc��M�2����e��5�N��F��^!�)����]f�����L#���S]jK�)��E�W(�5�JF�	����֘���d��}g������Pq+b�:6��u:Ě؊�B{)�{�Eď_uV~rp!"ߵ_��W��� Ct:ݿt[<��L���H�̳��)+/�����]�q����[�@��m~����l��N��k*y:����?���q��7��
��^2��zq��L�k��A�}��Sm3,q$H�07�w��R#!� �vrq��+��Z�3�I��OSZV���	��lX{����N �����b]q[�%]覓�c�߱\6�/�"*�q��KZI��6�*�h­�c	���z�4�/ڿWɠصڟ=$���zt�sj�y�k�j�j����h_,��,ZU6��e�j���.��D���1OM��֩��������s�z&��Wb�PJ���s�B`ߺ��|z�)ʶ����O�Z�;!��x�On�3���JL4CF��R	�O�Qr���"Tҗ��[�l((xB�Լ��"σ i'�%y#��Ϥ��M=k���oy����G?�B�j��b�_�8wK��6(w���tW��:ݹ�67xX�(2t�>*5@5ƴ�={�
��_}z,:�4�W�_^�����J90�J���h�iRj��.z�,�93���A^ !e����h��ig�~�eڈ���:_�s�j�ʛH ۴�����w�{W�.�!g���ԋQeBb�=M�һ����
�d2xR�?��RpJo��k>�t�d{��hYj�r���V3���s��A�,���*7�ɵp؆���R��o�h?໥�k0�x��4����DY���Ɯ�`3U�̃��1��t��b�
�B��[�p_�N���L2h\����+�y�MlL��GԶ���~���k�6un�	F��9ekR}�ڄp��[���*��;����RI/}���hn�|!p=�ME� ���k�21d�]�\�X^F����0s1�ןS�-��7��>�h t^T�� c�I�*�~�q*�#Vi�S�8 F>);���Gf��%�;XLGCd����r��L��g�n����0��A��8����7TmF�e��h�0ků��z��ONK��i.{�W�cl��A�����f<hL­눿,f�C����VA��W�)q�afy<���Or"�P�;XeZ崟G�}�'Z�|�]M:��l��w�9���.��'����^?��JV9���vwr��ܰ��O=����tW)�z��lS9	��L���@��U�p|��|l1T��v�vd�q��Y����QB���k��.X�˴�* ;�d�A����k4�b� ԑژ����w���}�-��H�/Y�dV��]2��w� >d��w ����qT?Ѡ�>:�JO�x��rv��4<�M���P��yl#�^�[G��ٽ+v��d�W��H�tw;Ӡ�,K��;�H���$��m���tz�ѩ�'�o��W��%��^�ؿ5���ƛd
0f!A�3��H8~�4�v��-z�����l���p�S6�y�|K�����O�/s�	�W.��.o�3��QH���t;��z6�$�I�t��P���A��=�ix]#�u7?FoP,��Z� 4L���e��We�W�$��p:�Hb�h�12�T�sm 	ݢ�|g-���%�V�&w�-;2�C\�{7X|u�XR3�ARCA Ѭ��#);7�,���~�~A`���pj��XzQpp5�I��{1�w�K*�O��ul��Ƴ͎W�_*���v�����[~�%�AzX���v���2��3�8r��q�Ke8)�'���{�Wp����Ҽ=��¼�)<6���5/i9�3W\_V�<E�Hݥ�
ʷ��<,⊆Sb����D���� �Z @��)G�G��2�PIϣ���%$r����I�[{����d,����2O)����G���/g��)۩(BE��B6jK:(ߢHl
��{Ŗ��R�R2d��;a�ј|��@�C�H҉	�Q}Rm.y��2V�-���8��IhZ)���v	g2���f i��{�����`7�6��@�=	�Ą�Y�׎���%5�b��I���]�Hio�#U�(��5d����\ca&��&Dh��4���2M%H��@��"j	�t��]�ab�t���dJ�@2���{^4��̔�>������	X�ic�p2���[![/ɭ���f.�u���S�G�h���Jd�$�4��C�ν�Ql�!=Q���e4��}�6�#���`���F ��j�	�#Gª뀪��>F��Z�e7��x�s�9;Y�o��q7N;I�����,y����)�jl�/�񵤅pu(��F�[iV��S��#z����]1t���-���N�\8�3X�dV��g���4��3N@@��FUfb�Ⱦ���XqK���'X ��	��BW�(�¼��iw�B�t��0��Jm`	�@��<BO�r�L'
���c�{��+�:f�z)�Œ3X����Ar!"cW�6�aM�.��|B��7����6�z����i� �3&j�P���k�C�K[�T�Ȫ�o�H�.+��i�*�]�Jm����8���f����Uws#��7����aC��~n>�@^{��	�)��tEq��}�#X-.���8��\�T�"��.\&��_�3��3�i9��2��9�U,�^ ˴!��j��N�̧��_��RyA����������i_����P�'���%�h#7Ԇ����03~gtq��EqD
�,��6BT��r����S3$x�6}wq�䬓��B���}Ŷٮ����W�T`L��+�66n²B�a��"��0�F����W���?H���(�2�����@�����.x~X*b�m&��/B�}�O��%��y��>i1ihb�.X��H����X/�`���,kV])���I�yɿ��hO�o�
hV�Jbf9dY��eL��	�s kS/��T��,?�K�� �G��5e%'<8��h�U��jO"�������6>���>�#�N���+�뀕��6;���qd���*"�͇��@eq����I�J��r:�"�>�tzc���ERtS	|�E�,�Д�s��	������{��(��׋/k����/�9���~8A����`�٭�.:���G��{_���<��F��(�p��O0��uR����J]�����ק:����<�^^�]��gzylv;�j�O��<`�Z�����^�/�v����`�"�O�Z��f����˗���c�7�7�Za�f��ȓ���}|��{M�pg�@v�"��]�-�/�G����=8�����N*MQx��6�R��m�U)��=�T������z��W���^M����ɥ�SO�ݴ*'�����-�>�j����N���{�b
(=xRϷ��I'M��n"��ah�t�!�*O��ۨK�D�S��)4�y����Z�w�=��2>�)H$LOP��=�}��d�=i�����27�	��=L`�~��!�b��f��b�CfC.�Ȧ�!2�^;x<)�i�L#����E������kG�Y�n����:kU�Y!�G`Z�Et"+T��� J�MSW7j�iu:e���y��{Jit R�|VqOJ�Dj������&�G������9�4����>�8��_��!�r<	P���LEw�˵�uB�G��������|H����T>9�>ۯ�_��S��u%~N�cb�g�C����W���7�
qR����o4Ä�-|����R\�����;TA<��r^%4Q*��&#�H�O^ԨK��:^����.�)
�S��ks��v���Y|�J�M`�ކ<�����-��305��+�H��E�Wְ0e#V����}
�%�0'qw��'m�U���@�8.g�������
�z3|��:s���l���">-U����Ji�a�8j�*$�0/�v���+}Y���@�gx&��r�*����,�f�q���,�P���{�Ɉf�U�s`N����'�4ǩb���2��3i��d~*_.g:J�����u��AKnm�����mNZ��װH.��ǐ�m)2d1�.��|CC��0��_SOy�h[�O��x�u�(h��Lr�PB��7X�'�7�f5u+��0Z��}3��>b��τ��1W����0J�|/P�-��/%$l5v�����\F�_�b�-}����Z
�{x!�� ���pW�Q����!71���S.m�Q�ua�
ҩ�:�F岘�L�������>��w�Ta�#Tg��ݔ��i0�5���"UA!�%�Q>��.c��ɸ�� p�z )�LU�p��.Dy�lOH�a�@j�`R����H��A�n9z����.�k} �i؇C��I���}S�y3�`C�r�l�Y�P�{ԈG��5�<Qf;��[����,��{ͯ���̾]u��A�;D'5U��s�B�����)+ӭ�����P��.+�����:}�j��)#-)���9�~�of6���RY��ʮR�z�n��,�''�F���X!|���.ͤ��]0&~#�"�x�^� �B�ih�i��J�|xxJd��a���1�Q$z�G��; 4��ѱק*���E5�o3vA<�m�a��0�y�\�^�̖�f�4up8�p��U�	y���ZSP_u��N�O���'n%���_ 0�I��Z�^�$������l���j�:ѐ3ŪD�.~�옒>���(í���w��h���Nw�ѽ�'�0��rg�l����`��ޱ�R�b�*��!H"/���1�u�z���{�x� ��\G�2�q[�m&ohzab�!|�]�o�.�YZ��j��!D�O�浄��\vA�v2�a7F�{���2MQ=p�c�ea�t+��(� ��LW!���ۮJI�v���Vtv�|۳No�1Mj�5�_S;�>�b�Vm�P���o����Lʭ� ���=�8��cҏat�l��n��a���X��|����9�EБH��G�H*-Ֆ�g7�$�Á�Ȁj"�H�����-�|��a/=a�ٝ���W���V�vZ���,a%�-�&�h��`�|6�d�J�����?P�_#�f�Mn�ܽ��VƂ�����ހүQ��,�EKD*7���MM�G�����y�IlX?�h���N4`O�>/�$D�����B�i���'��wދuءm�9����i]�<�E�W�����mf#���49���h�������(���B�u��s.q����OU,?N�y�&�bf�zfP&-%q6���x��@L��a�
�����\���a����t��Yǫ?�YM�Ҿ��h��v��cX�W_�i�3]�G��C�9�e^#0��}��� uy��_�0�^��e5��+|��́+�K�1O��
u�h@\�ߠ	TW�ĸ���:MJ�;O{#§hx��?َU�Ͳ���:�{�HKb,a���>[�Kz@�9��v",��ug%�u��@����b�X�K���c#4�C㨱�@�折P[����\�t6���dOv���*I�x�E`:"5������*_zc00��gV�J�ؙŢ6�*�4{^���x���̈M���� P|�mo"���|{:?8?H��o��;�ۅ6��qwP.�؄���X=,}�џ��Z���tk�/��h*�hE7\ӧ�n�:\�V�[c�,�/�-���R���%����Қ���4@�4��5���sP�.�D�{����U2t�ҋ7&b|A�j��n�m
�E��X�;�D���T{9p:��m[+��O�e�P���0b���F�?5�ni�JZ6�Y�w��ʽ��Q��u�hU$_�	^�Xz�;x���5�o�L����!�u�N.��F|:���7�W�o�����r�Z����2Kù�w�c
(��Զ�B��y�����v1r��~��@�IӪkZ $��B�}Op��LWeʐ��8��D� u�в1�]�o��]O��
�кCi��s��2�]�P�^�zkj{�`���qZ�X��U��՞`VK9�̭wX!3�\���Tu�O��	�i���/ӯG�ڏ�^5�>��ײA�D�8|�}r50q�H�<T��_��C�7YR��u� Sk�~���W�����W�K�phA��F����o�=4�/��d����d�C��4�wŔA��0�
V��in#P���;�ؽ��fPȣFJ
�@��ʥ�<�&`X�w;:������F��� [�.���[&eBC��@1eF��Q�ڂRNI࠻�n	H��}ws�; 7���.��5�"7���0���T�w@.���1���f��#�\��J�ʺ�8<���h��<`�l8��(�v��m�qKcl��cp0�Ƙֻ�\�������~ʨz��W#�}揤Q9$_3�3EP��[��m�e.	�Js~��L�'�!��0��>d�Z��b�Q���]��چH:��6����S�|osᾌ�C�g���e/�I�K���T�j�E���pU�)��UOW��~Ru�+��n���ڜ���	P�</�.�
�(;.\4�qTТ@R[�.��Y�8*U�?T�Lu��Rl���e��8+��uB����D�jk�'����(���JW�0����Fc��*
oچާw[�E䜹�'���DT�g��_�N��D�_\zO`�Qɸ[t� Յ�Mag��E�?�uҨ���>I�Y�$L[���\��g0��Q:TL�g��j|��7������a3��8 +f= ��o�̐j���P��8=��
 ��i��뢧��Z�?�6���@��Q�G��6W3́�^B`ċ_�S�Au�1���Q�26��0���O��a]n�8Z��t	����@E98)҇v�_"���`�������d��xt����`1@���1�׼/�q5⽛V�O�r�@%'��2*zT�`&�gB�w��V�Fs����� ����)�G=4��qM�ј� �mCg��,d�1)z�r0��/���F2r��72���uD$���C|v�нed�\he�߸�{V&j���ÏvLY@�L⇱<������|�ӱ^�c*�,˦���gi�όҡ�DT<n�.��'r:4J���S&������\+l�$iѧ,�n+_����;�� �V���\��_����n/��׵�!ҙnB�Ufۿ[���`�e�.�Yr�Y-�.f��i��z;��z�x.�PG��60� �֣�J�&b�� �u����J���ǷS�8+������JM���X�ȼI����=��@4��2!A������=�z�r�]���
�t+m��x�	��cI��_���G��vx�(������P�H���Q3�>w��?�!ODO��T�`�&���dMJ#�]W�#�_3�΍
��-���NV��"`�w��~h���uy]n�~����񹕹�:#.�U:�?��C�|}L��
�^���J�I�����B5-ޠ6וD}��7�j>����b2�A�3�� 7f*��e�7,7W9>��sS
]:�cn��g�:#�#�i`��J��^Nq���ӗ:9�t��8"5�3�䦕�V�wQ9�3n�?�Yئ�+��V����ǝ�4��8��,RQ�K�P^ܹ�v2=��?�yO��8ΞF�;Aഥ;�G*��5��&� �hBs%�P���w�9��>� iJ���	6�=_f�e�\�Ͼ�� �PH�;1�^=���)��l�6{hDm�i#����L���I�u ~�]:��n��e�W��M�.� �N��z��'X\5|�*��"Z*E�L,���.�l��yq 3���K���it~B����bi���D&��]�'�� t���G>N\���~�苞A��wj�@l���I|��hx�oᯒ�F����I?��SA���a+����1�_`O�9�����[��@��\M��<������U�+Y�tPxf�N�<n�(X����ɫ�R�\��j��c1a��m�`���T�n��V�4#�=2������0%��L��G\�&����?*���"L�-�Q��E'ˏv�A����jBB3��N$Z�����2�n�Dn+�r��J�ܲ���5_���s������1���At�p4��]��>N�u��z��� ~���̚w��x�"}	/�Mj8�?�!�&�Y��rzkj9�+	v��5v���ֿN��W()�@�}�e�J�M�$w5�'�0`3�\(霵���C"�`x�=��'��MX��4]򗺲�I�2�,0�1�ʏGr<�I]��ܵm@�)g2m������0��2zy���p�3��Ms���_��ƍI��Ys4Ö���T���{�z"�[U�r��l�Q�������б�1<�$Z���_�Ijr7�T� ��Y}bW>�ѿ��9� ';���jg��Z������<z�RTC:���Y�kY�T�@�hJ�pv+�M��n�d�&��eB���W�����bG?���g��R1��7+IT�7�"����Џ��N�&���4���}��*]��k����~@C�д�:J 	������;ĀmV���q�4oɡ�uK9��i4�
�ʽ�/Q�� ��¦�h�K:���.ӛh3��[�p�N�T�_'TAty)�z�zW5(�"*���ɉ��ɩh���i8�)/I���O;Q�6b��I9�}��߳��|�:�|��"@��$,Prc��L)�5m�U�!(6��C�x1��Js-E&ZaQ\�60]�8RM-����3=�ðX�2�|y�0J���_w�88���EGC��`�^o�8�GBƛ�/�)�h}zN���k�pr�W;���Ϣ�Z�D=+u�*��_ �`!mAu g?�˚�pM�������0u��(d���T}ɿѐ�K�X���A!��f�j�(��]Ixi�:;�Gy������h`!Cο�x���SP��+���|���{7���ŝ���E��v�p�s0h�3aH�g$u���16��m���kx�t�e���s��J�5\TB�-��[Qj��N����1��������B�����^!yE�k�MΌh�;�dԥ�g�/x�vw���]y�u�?�^�k��.��A�QY�ΚH3��m���Y��O�2����1)���!�Q}���n�r)vY[T7�K���e��5�R==.P��J���T������Q<胓���9�7�16�=N{.R�f��g7���Q�$u�k����P�R��8I7�J�ff"�sKP�N!x���=?I�=j������2��%��B�W(� �I�<���j�{"ŵ��@�m�"�݅��Y���]jQL���'e�1�N`6#U��&l�߽�TW�ƃ�	��K�cv�::��\�~�ܓ���Q������;�u���]�#G�=ގ2��.]�B��ֳ�~uz�!�O �Ӱ"���Lk��J)�z���Q2�æl�	���}"E2��6��ė�NEZ��AЕ����A`W6�Қ�ʛ�r�~�j�hr�J��`���ILF�S��z���I5���%��OUOH�W�y�C>�w��(�$�f���;gg
������K|}.3ξ�N8��[���o����]+8��j�&�i������V�������n��I�{w�E�!���,����"��o�.}F�5[�S��a���g$�8F�B��@^�G�J�B2`�����L������%uD����8�y�t�F��SV[�]���/ ���B�_�|�lx���JL>��R���z��^���j�ZV�>p�R��ݓ�R�V,��^J;�r �J:��İ�l B�ۢ��`:葸�H������E�e��x��	׋�]����;h�u�Jn�f��8�:z�t�It��W'}M(�Ǘ��;#_׫��M'�����2�M2�m�'�)~;����"�caQm�"�M�\k�S(>�8HR"'o#�"W�_�䬀�D|�l�����G9*�FYŕ]���\��C�l+�R(��`.kHV�Υ��ߑ!��s�g *DR�����.���%V�䜆��boʎ1�c��c��7U2��)�dm�P�.�=��*����)�O�Z ��g��K��Y/��T��i�<����g.;[�洄�`$��pm��n�T�����~yzl�X�-7Co���1�<-�5��p�zB�'��^Y@����M`�����uN$q����E7̚=K�#�Z��yl8�0�*h���uRxS� n. �;�|��#�0����`���S�X�F�0G%ɭ~����!i�U����X����>�Z���t� (9�U���u�^��zYO-�/����=p���qI���FX��Þ�ds."��*K"��xkD8-�41_�/�^]��C�.�ˡ^��_]$����EO���av�� ;A�BH�柕�wI���0�_.{S�d�����~�*���iߪ��W�zm�Fɲ��a���r�^���J1�����g h� >�^+S���(�U)R�	�6�/���
����s����L�Ŗ�W�TՐ���V�˗3�%�҈�?'�e�%�!0xV@��G�(�b�nK�.�S1�����1
b�����ϼ�"�Cٜ�g0�Vf	5�e��#zA������n��T��g�����.�i�3:t-�,7��$�܇]BE�%�����25�1��w:���|	�t�9�~%vg�B��Tc���o��D����s��$ޖ6&P�ݵZ��;���0>�ʪ�P��DUQ6'[� ��C%�:r��Ͱ*�A[��/�h���\�`*DP$:;	��)���}}�	l ��(�hX��³f܆��_��[����}�D�7��B��;�lZ�6�z��9V88�5Wv��~^~SM�8��KЧ�]�O7��]�����'cA>��۾[�:�[B�=�#Sc�΁����gށ�M�~���v���BU����c$���}�A7�fwRl���,�Op�رOoH#��`�8&�ј83 I��)���F�2K�B|�Dj���cG�:��|���\�Y0Dִ4�O���/��W��-����������p����9Cϛ�qt�g����s١7G}ܱ��'BP#}��|�k�	��+�_.�	��Kq<3oB��G�6�}zM'옮]�h^����r�n4��ϧT780�}U�F���?��g*n��̑\w3�խkZK|5>�����.�<��I�<%���&��D�aT��n����m'�ş���v����/C�i���g�ԋ�d]��E;q�	@���O�ؠ���+?�߅h�����d��˨뎘M�l'�@3�J#�����s�� K>ý�K��l�/��� �k1��qW��~�|�SYEfr�$H9��X�w�������*s�٫�0�n�or��ԛ�kz�8��RN;�ΤZ4Q�^�Da��	��p��غ$�ylݲ���ۺR��Q`�����-�gK���Vo�ȹq�3������A��[��'i���d�oq͐�MP^V����k^P���:��]�ރ_`Z���~9��05(��f�<��I�ȍ���:Rl�0�|�G&x0��z*��{�DS�B�-.�1�+�|`��x��B8=ન,:���n���>޷��\�3���)&+�ȑ��2��
��Hu���m�V������?.8_u��6�z��7ۻ��
�����E�iI����6��c22U۳w�z6P��w@*{���h"7��J��`Z�-��Q4��ǀ%.E����3�]k�^1�J��kƅ���o{q��/O��_�a6�*q�%w��+�M�@�c�~���m�m5��+���cDf~����h�<[���3�Nj���09��4q{u{�?w��g�GQ$5Zت�p�q4?�k��>��:`
t��j��ծ{�c4�����!NCj��N1�I���r1�#id�sR%�^�V}z���[�ڨ�x�,�/n h�����>-�x��#���������*g�mm_^�#>�P*�b��/Xr&�kڪpzy�G��/Y�$����2���t���L-���ݮ�G�8H�ַ^�Y#Jب|�\�]��Q��A^�X�?��[��3r]�J&����h�nfQjZƅ��e �~�f�y,��5�4�CݪmZ�.�2<0��ɛ)�+gO�^_�� (� �3�a����w\��B_� ^Cq�&�"k�����(�~����mb�G�!�AԼ���:�QNh'���m�hL�[��9�]�F��n��G�N!G��Յec�A����A�.��$@ۓ�[�C)��n� `�=$tYb_���/�b�w�L?�7b֭��ǉ� �n�K�#���j�?��2cߍM��K�rT֛p���^3���#��(���N��~�$<F�[�=,��ʛ�zx_`5����~}a��c� ��Xe8˖U��Uk�c�� 5���߀얡���q����'R�O�/�K�bEH� ��+V9е�D�D�v[�٤jb�������HWjEM�Ӡ�7F5¼���"݋�3Ed߶����x.n�]qU�K��e5��2�f?�d;a=�H�W��(��>vS���<`Nnu3���H��М��8�<aVvȯzh�����t\�!�Ө���;c�D�"��V��g�.@H���b�>̈w���̛-f-����m5�~��t]�������rm����p�/:��t�&��3��v��n��Nԣh�N��x� ����d���wOC&�x�Ahב��JW'�[H *q�S����Ln���R�2�e��}Cbʝ]ʸ�瑈t�e��(OCȝ����ZB�V�!��:r��'� m�#�]��5��6����q�4{����{�"A�a�
R�0���ξ=���B!� ���04�+�~ÞUe}wz��Z��B�[�	����d��Y �/�h� �`�H���/�!�`�k�'�cf���Kh<����`�J�U�M�Ì��$Ӧ��ުEA_�����O�D��%��'�V���Yj�81aAg�����=�����5�Ψ��&Y��JBkm��N�hvRHl���{�]��)��Q���� 	jByM�;�O #�����!��+�����zYǲ�k���5�P�	����R�P��pd,�N�~
9;�m� �OOO�$&����"�q1/r�i*�wZI� �%���=5$=�-�g"��Ql���G`iMU�I˼��)�g��X��o�yk%��=�Mm���n�0-X)��x�=������Q�g���s��_?/�"��y�'坽^Ŀ*Q��e����t�8�|� �,�
_r�<�d���|�d��v� k����5�T.�@W?#�>�0T�Bv_5�Ym�YoH��qƢX"	i��W��0q.M���~�	"~�OWI8���d��^z���#����0^)2F�a'��0WF��`��"�(^ژ������7j�Ԛ6������~�D�Q:H�S��J��?w��I��	nDQ8t�#S[�1	���p��V��k�Ov�EAQ�D\7����zuꨣ��DC���D&&mŞ���0;��pH@���Tf�n�q�!@�W�Js)��f�5/���w��g��g�n�I`�~9>�D����Og3�z����O�s���q0���N�)=5n��2"����U��r�Y����_캈������5,z�8o忘�L�q̷����:T��s�	��~K|��ϓs�~����5z!儸֦�Ƈn9����b!o�Y��(ib7RB��]F#��}@a	� mTY^ߡx�d��+�l�P�=,���QS#5)"���S�j���[Ʈb����3c�7��Yn�(zAC���(,�f��AT����޷$#��f;�c�U��w�����N.���m-=��V�r��Lj�;�0��+�3}%��ч<p>����j�f��2�F�?�fd�Z����tJ*�Y���
�>[x�%�?�7�R���庤M�F��>���l�w!Ϩ�*+���hdNHO�Ë�5f)���8�n`���Vt����m�_��sC�5�Ȇ�T�_Ô�+� b�����q�M�ӛxvS%y�M �;0�j�2l��m�K��<�c/NY�Q��2�,7;?�����?*
�r
Ilo����^��A�������s�<��#�(K�ug��,M>v�f�~02(q��e�#	N����&���=)���9�%��U2���!f9��͡�7"ȩӎ�#v������b@1~�_$�N�tZ�~\��Y值�z�Xl��$j�W`�K<}i�S{"��/�8�fp�h�Fȍ���z)�WD���J�ݦ0��K.ŗ	Ɓs��"V`,���/Ds�Ұ���9�(�ѕ2��=W�c_p0�Vq�* ���#OV�g�s�pm�ˣH*����k����É�2X�WbK�-�D�֧��D���'�і��<��M�#��2@�mS#���a�X/����BR'���M�#���B���{/��r�[�M?lL���h�,躆���Xega�˰�Z�B˸���f1�u��Q},����}��
���hg~��.R�
�����F-�q�M�A�$L����B�ZVK�b�K���� s�-Z�]`S8���5 ����@Lp�Ӯ�;�^��Zj��x%�+�Ē56�#+d	jH�Th����/&� ςb�OЧ���aj2�`�c��P��rD�B����K�+���JW����s[��:6r�:�p�h;��v��CtJcc��q�鯄.��xbi�,���g�@@��t
W���+��2�3U���nt�{7�M�B�)c��W͞7���˳ި��~L+d�M�@GM���[U��ܸ���"@Ϣ��n���N^����>/3��4��.�&`Z��# E��atB���y�D�W5�5t��ҧg2U�V���4�EDg�r��.zRdm
 ĀӖ� &-�5�����`q��\g_O����U.8�ئb��ר�q��'�Cٕ:�n�V`���f��B��xK�;����[I����$1��8��m��=J�;%��d��섕�l�f>"D��@R�/!�V����Ǵ�����
�RG����$ptO��#�=��ʖ��h��V�A���BS�����6�
�}���@��:�plYU�,����++�����@U B~K|�H��kL7�do]<'-�b=��~�k��/�RoD���P�+@����,l)29��HF���1H�ΏD|�7`"�/VĤ2{ڶ�[������Bypٌ���c����x��Xi��ǵ�
$��������:�&���{p8�����{T�B]q�!Xg�#�e���,�ƨH�N���E�����y^C�����$��?��D�١�UBC�����ks���� �<@��e��/������8|v��� ��vs��d���BU����B*l��r������w�� ��P6U$SL� q-a8�'#-�6�vP��UK`��r� �ףV��ݼD���p���_���.�=0��b3h/�J��q�AϪ��9�o�!�D�=K3V�V�0	<=��X�ye���2ڿ� �&��cU�Оu\2�d��[m�<fH!�wr0�j���/��� Y[�m����Q#��s������Ҟ���/=�U���4;�����x/8x+���/�n�_R�F团aō����q�~�)�����ઔ=Te�O8[���V?yF2i��~��WK�� +������1pĤ�n@�C1�H `�9[�al;�~%n �
6�<�r��$�z��c �4c���wg�ր����{'땁���!_��Vz�D�{읬CKpkV�GRT�p�]�r��7 [��>�i���sF������������v�D�1��j��qur�,�+H���O^�D�vq�-b���97Hx+Onx�'�\�'��C�"�x�d����Гj�����N���ca�&}'B�Q+���"I2y����~�����-�mU���tBj����q)�K⟌ �$���!�8q�kr��&ڂ ;lY;�b������3�U��ӽ�.f0���y�������\o�Q�hឩ�n�7f�.ďvq��0�Ŗ3��6tIs�à���X�X�m9��V#�O5ɀv����V���T�lg���3���X�"|����M?��8�����u�g����W�ׂ�<�����E2��j�@x#�ڮ9Jڦ��#hߴ��yM�����_j\b��	����ۘȱ�����vځ��䴆<6��!�������fj�t��(�0�.�K����G�]�����qUH�3I�Q��(5	�+��0�)��a��%�!Y�"���-�@4ّЂ!�7:!d�W�yg�1T�
@X�����C���[O3�������&W���
![4�PrgT�o�����tx����?�ئ�nzNc���������C(�b�R����g�G?D�����X*��k�Rpа���s�c��N~79f��j[j�]���x��QM��W0Ø0��U;U}pBդJ�&�5,������@�I+u�[x빬�g4�^�ϰUQ����|�񓋣��ʀ6��O�Њ�/�3�+Wb�P�x��[�y̛ڃ�GR����K���	�O3�,�B���<7�Dmc58@%7h��&�=�Y�f�C�Z�L�v6��%,ւ�Ut��
�������H+U�!bM��d�Ã���3z��N�3�}����%KH�vӝ.g����ꍺYgL�l˅��5d��+@�S�]K�qL҄�o�a�4	Ɩi�	]�1	"����:f�$	��Wg�.7��K���D��+�s`|��BP-�/����g��p�	>�f�����WhZ;y�[%��х�8Z��D�~U]P�%��b^��Z@U���K�zA?��W�Jfu�������s�h8+�W�rI2p��]4S��ڑ-=% d�V_S���i���7�7�.���E;�2��П)�X��$CJwH�\E��I74q�:[uP�f��kߺ_�X4qg0�� ���}L��چ�N�nII�':3=�g����TI&��j@�E��9��ʀV�r�,T��UN7���F���j�e`���X���*גW��\�sm��+�[�������C�n��!\������an�k��c���s�v}> �����U�O>�嚹F.�r���k��V��*���X�Б��!�{�Y�V��$"��L-K&(��A����yl�4@>�9D�M�=e�������������@��9�>h��b~P<]�����{SQY�ET�耻X�+��_%���PV��ޞɻ�~]<M�S�ALWܓ�iwU���0e�jc��k�e�s�KǶ���
P������m�شi @h0�����q�&�%S����.UI�j� 㛟{����2�0���j~@�8�vp��"X����'�&Z�����}��'����c8	\��`�Z�C3����)��^���U��j�AAT����%�2�$�p<���h t-����T��Z¬��(;�	�3Π)(��O:7H*�##�\�p� �����O*��$m��iTi�\��e���&W$���h���������Of3��"ש_	��/�G�OblÂZ�|�o�j{q�����`���%Ԝ��2�եWE"��ݷ?�f�S`?3��[�tե�T83&�Ik�w�G�W�B��E+˕?ݧ��D��aO�e�ŝ�ܘ��@䶛����U"b�@�ex�ҁ���\��2)���D���U&hغz�$��@��~M/�ā���U����ET�q����I�~�h��r+�s��\�MX�a��`� w�n�u�B����T��}Mرp�.mu��ڰ��*�	����T� )q�?e�3.6U)����l�7|[�����ɡM�\�閂��������S[>=�ZG�uU+���z}i�r<�����9���0���`�u��o`�*�֘v�t�b�p}1�[&�$o|B�bZu_U�c��#�c��;q���K��IX��4,"��:��څ1zs�^ѭ\�Z�i�0<�w�:Q��g�Hu�� i�q�:��c����+-6�o��tf���W�
�9�w��p�}�F���Ds�G9�8s� T�b�4񅛬G���'�x>S�[��ޯh�⪢R�s�.��-�ݺ��v�2*�[ٓ�N�h/�;����`�[��6�iH\fA�C[��1)��C��L9^���\���2Ϯ|���D�'�4 )�y��k���<���vm���@�}PƋ����u�����ӯb5��"jP��)b�������,`��	n�7�c�]g	)Tf�G���'ǆ{%ĒK��2c�[�"h�=o��n!Hs��
	�W�E�OV±WhX���:@'CX�1���������,���m_���sn�|a�PIή� ���*A�	%���cs{��\��Tg6N�+��7�t8�Rz�`H��P��؀�I��c�c(��!���|lv�h׏Ps� ̚Q�mQ �M�v�54�D���S�2���TҪ����C��q�c�^R⹁�~���I��qa%�~��ǒ��0�Y�}z�v޻�@���8�.�V�itV�3��������I����/SM�KH+�"�
>(����Im%�1x �U�cj� K�|;���iS7��Ϥ�/!d����*���m���h��܆
AӔ#2c����z=wxPy2Wi:�> >V%XT��!�`��B�ˈ�P���=����n��:�܄���Q/n��t�Dhx
����W��5d�2\e�����̪�Rdr��EB���U)_����d�D��Ó�Y�{�����!���ME��h��ѯ_j"��b5 3����O4M����	8�]�4x0�ק*�>�y4��NA�!J�>I���.�RO:���^���Y��p̫#�T��T-#|!Q��.zG�c����7v��)����/}��h�ޑ�묞g�k�bXص{�^i�炳|,VP�H��fl��?G���� �S�� 1�3\$	���o=���8�(�(Q�ʝAs�Rt�#���}y�����r��u8�3]���|	JU�dڏj"E�P��)�Ԃ阐bulR�}��_�K~��g�1�����-̀J�t�
>ȲV�ta��t���bj����4�y���w�u8���{�t]R��k�����*�+ܲ��'� ��"������������f����F��jgj��1�n�@G��{��O�?����+^ϴW�_A���pG�ߺ���>�����}M�`�Xi:���e�$8@�?�|U;拳�IL@�>��C*��툘���<~h�D\�?J�ç��e@x��f�bt���
������>쟰��㠔`p^K���,i�]	�p�O)2S+�у�aMXP��5U�a����ܦT|A��ӮځC�eg�U(�jΕ�Id��]�.(˭6*K��ɻZ�P����-�5�8y�ڒ�8�-���"�S@�<�����ה�f����eav����]}}��������ں9`WbC���^�7��҆�(���s�s�pR$�����?�{��K�%w1�	䷳�v+(E�L���絁oMD�z4�O�Oנ׋	@����`���cDKS�L��:��A�Ֆ~L{
�$ݺ*�����ROe�k�ky��^�#���#XfT�������bf��5J�w�hNE��T������s�� �r����dV�4�3B���k�=y�k�m7ʔ��A�x^����l4m�/c�Β�̎�O��F����T]>��յ��sTc���3�1�齲�H�N��u2�,�k��"���mZ�@���')���
-H�����-a.jad�9��pAq���l<X	��~6�P�f�q��%ȗ��y�0&�T�?��s�f��;��ixI�a\�����P9-��Tټ�R]E���ƫd<��P�C}�ͮ<����Y������x�\�^�I��"ɒI�XH�G�eH"���n,0��~"�Ŵ��Nm-���{cؼ�##0-��/��8�筀t�E�i�O��#�Π{�(�/��F�	�G�q�h�'hM����<��㕛�	'xdќq�~�ק�P� _��R�5Y�u�UwB�OI��c�gC07�k�3�4jU������v`pa�X�J�3�����I�.�v�5�`Y��άc:G0�d��_x�N�]7�~�+�[��jjg��N��4���JzM\;����xevbUDnr�G��iv�LN-1p�]�vrS�
�c��Wr\�^��ƾ�!hm�DE� �Y=q���J�}���(�>��岆��UF��zu�M*���qf���G*�T���]_�X	����9�<��k�	�
H�x�K]����F�1s���4u?<�4���pE��������C�n�����GU��8����z�Vu�����¥�xS]<�����L>̗�\�%	���L���yAMDO��ܷMG����(�%
�E�rf^ڡ�aON���I9�<s1��Ι7�L?ĵ��U�}�w���*JθJH�q�Q��Nm��om��nCR�z�iё�%�B�!N�+��t�f�t�n��5��i^Jƾ�Ć(R����͆AE�c������O+��V�u��A4`Cd���=�XƇ�����U��u��9�1�U��v�<�~���,k���z0�j �U�]��5�m��J 1���B���$w-��&n�n{ˮ-�^8�`�I{4�=��4����5��o$�A���?�i���X�h���|�5�c]�����e�p��J��=�>^,�Q^��PI��o@<j�4�ΉQy0ǽ���|���,ɀ0� �2��Ɏ���[�d��/:O�𐹦´
nP*aKH��W�i��(%H@������(��v�s�@:r�L!V��v`6Z�ʴb�(+�C��%�,�Q�sf�P�!�"z��e;bJ�N����(�0����8)��vD����9�8B��JX���}�L��a���j�Ys���e#��e����J��$W��������jD%h���=��jI���@�w��Z_I΁���X�`!{��>!gnt�&O�@Mm��l��/�JW�ow�%�%.�波�"���;�	:�\����@�խ>4ʘ��M���֎���;뾌�j�0.	8l��!g&�!:
>Sf���5��D��//k��A(##[��E��.R��#��ȷ�{C��dJ9d��܍��2"���o�<	+%vclؔ�#sTz��e�x&��ͤ�@���o��'�W�;ZS���`�)�����iy:�ȑ?��9�o,\L�`��N.�t���3�/�-�$ ��-��ПF�2i�P��Z�w_�D��NC�3���Lp��HЌ>Kk���e� ?(�>��0��Fx��w���ofIX�W�ğ�V9���!# �����8-����%V��p](�W��=���%�:8%�BOj����_���2�x���[����*�i'��{� ��1k��Ϸ��O��[�5�	$ȿ{�����'bk[����~iD�9��{><���}���u{d���q���G��N-��_y6\�q�'0��kg��?l�`|��0�g��t����9�{��i���;�����L"�y�A61Ʉ�Q*2k�4�䦦O�k��.h��i�ܬ�l�v���%�NYC�Ƌ�?ۄ���D��"�u�����ߌo{�ݜU�/��'��Mc5P����@��'~�)3~�6�p]:���[l@�2�(�2׵\�#�,}�[+ړ�k[�5p]�������r]��L;~OZ��ͦr;A9ئ��W-�dwvz��������*�_vB`�D��4�:H����"�^*N{����L򣗹~[X=����K_`����r�oL��h��v������"�=K������cn��j�B2����1����["qzb̌>���QS#"��>����<�h�&v=r@s`<6��ED��O�J~�DQC&��@�ֳ
ޞ���<>�".�+�8����a��+��t	(R�LcQ4!Ь7Ik ��X��iC�O?��F�,¼���RԹTk����	{�7g�{!�[�V�Y�X-�b�h�4T�4C8+�["�1��|Ѝ��(@aL���g'lW�Ӝ�/@�͞eV�(�a���$U�d�x�ݤܳE��̡]&
���u���TI���g��+#�1[�"s?<����Bߟ�w��A�VY2�
�l�"=��u�s+�!���� ;�S� �[����˲���>p�u�5�����Ԣ�?�4�Um���C:�z���~��X|�$��Ũ[q�U�/(2K �g�<z��Iŀ�އ��?EyR崬��k�֛�L��1�$~�l��Ck`�i��ry�,����9�k:��h�-��"���W�]v��5��;eW�����q�Y~BJ�����?����9�(2�솑VUISӡ��S ��^l�2�����u��Ԝ63S$`��]OK��~F���/[����!);���b���uL���?�)��W6���5M�r�l�CC����W�K�Fu������9��b㱭�8�wEx�~+�=���$�(�6�R�'����=�!k�*}���9t|���G`�a�r��X�I����V��X	f���3��fxr�&�	ȅ;;���q�Gi���XL���� \�>�D�oˢȦ��O	���y�&B���@s�{��i^����}��_L����@��~����=k6���66E_c�5�A�ϰ�n��F��Rr��e��/�}p�����GC�՟���T0s��r��3~r��&��w�S����i��y��Oh�ɥ� �Mƃ��@�'���g=���֟[����,4���}~U���=�(�)���H��K��1��k�}��vD_�5�ce�vT]�U��I�Vvf0e2�Q	�+b(M��58a
-9�,��Re�-���k��F>]	��?y4��َ��V����eN<pӇ?�X�*��=�+3�%�!#�� 9����ڴ�p$�p�?Qzq��+�0�������-]�Ī�'�J�B7�O �6�{�ܞ�P�_X���vTZ�P���H6�:�(X.���q�4�*i�zW���Y^�ɧ�G%��D8����m���(T�\^���	3�l�5%`'�'��彛+LjP6���O���մ��%,��Z~٩��E�ew��arUF��;�o�\���@u��熤����2��VKt�W��wy�0��c�����Mq�?#p詨�VD��r�k�Eȡ��??�W�R��Z~u��W��M��>��,�HJ�i8�3�HӁ�J�]ta������h۠	K�
QYe2P����O��U������[���$�
�[)�L�{�o\go���V�$��[�� �����:V^7���ʱ1�
ۖ�N�$o0����I��7΀�<��0YL�Z(����.쀧�`,'���lq�����U>=�Ґ�+ΡW���"
&ՠ�ʏ�rJ.����ô���B��Z��jB_���Z1&>lu��e)9dn4ov�흻�MO��*���r�ݥ�2?�W1�2�ӥ�-����];$�I�X��YSy)M3�6�kpO�#�G2�j�����iMb	�$��L�^�m��]�,�<:�Ra���W��&��F�|�0�|B�c�V�ү8�VJl�K�JayYq���j^�v����6$�=���/y�o;ߜ_;H��˞d�ajH���"	�P�犎!7ڲ`q5��"Z~iAZF�3��;~����`
�}o3ii���uS�w"���0^>;�p�_<�d�W�規�OAO#�R5�d�(i���B�版�t�xFCP&��T�V�����wRru��S�xTW�0��~��b�B���b,錁��qF�թ0yz��*�`��V�ܭ-?0���O���-S���o�u�Py�Q�ANI�q�<��!Vf�p�fD��LE]+���L�^�`|�~%�@&8�L��������o'�PR]Z���1�=��#�7J?t�ٟ�p�{`��4����K�i��n�γ����3���K�FהN��F۳s%M=���Dk!Z@ �)������Vc�<� �U6�}ů�"��"�`�4�F��e6���Q��a{��񩄄$�\��ّ�x�S�g>�I;W�:r�i.@��S>��j�p�O�b$rzA�+�;>;�﯀rW�Ia�L��L�C�^!/��ΰE7;�����E ���އX�)��,t�^��i��=�6��X�L�õ� iΉ���=R7e�ǵ��8�I3���e5E�&����g
^��}Xߕ�f�sw��EK�o��Դp Ӎe���Ac���Ҷ�hE��?}k�O�Ly��	���z��Lʦz�@��J���Y�e:��i'�ˈP��rd�o5���zy�L�"}���%d���:�hJ�7�u�lg�g�H;���E�#��mR�-�E#�����hWr����:�!E�N=�9�0�|�vJ�� ��m8����w�T����ˡ�;��7�m�������ړe��L��۲>f雎'����z���ncLSe�6��;MË���\5��'��S���%ZU�.���H�;����E&�G:t4�gU[v=�To�e .ŵz�@#QL��c��u��p6Ffgd=���h_7����B: QX�Y��!�u�r��[؜p�_p_7��4!�⒬2>)��֔i��٦�E����u��PA�jvψ�$z���/� ��*B���̞����W�~��{��8wI��d���A�DEq[��~h! ����.#r�M�9�5�攦YV[g��R�a�͡��/�@�ԯA�Ao�HE\iȺ�K����#��A�����b�&�h�:c�D2[����&E�'���{�����ډ�)w�_9��ƥ�1��z�wM�����2�`:�?e��|�?#�ؘS�	�cq܋����%K�᥾9�b��-� �-QMÓ/pj

q<���ߍ_>��<]�ܑ+���kT�j�~h�L��|bt|!��� k%��Uy����6��!6�h� '&i+�VF�j�ų�3�m�����0cF������Cib�K�P%�������*ƨ���fH4v��f:3�>͛�QP+��:���`�!މE�I�h��9
�%�>��RU�q��a�y$�Wl�m��R�M�-:����3x�nG�� L�L�����A��q�Y��4	Rv�w��b
q>��9LNl��h��姒���y>�ܼ�H���1&`@�iy�^&?q�>�2�8|G���qn�5TH��vK%&��լ��%�x�%"?�[<�e�&�/�������0�CKw�J-��5�d���%D}�Q�"}\y����:�y��K쵯}(c��غ)3F�~����HW�gJ�2tO̲��%x$����^vJ:M¸�}�2�B �W�����j|6/�� r�Po���q�t	rW�e�Q��N��F�
��K�>3�ަ�*�l]�ג$W�{��|�7����"���$g�bEi�G�߽�虀VdtA��J#4EŖ'aeZH%$�����F��:����"��Ƙ�W܀Y~׭�џ�N`���e$&����n"4�۞gA�uX��U�D�*���5���waf�X	����G�ۦ2#�`�RW��Ǒ+�,<�b��p��Rl�������>���Q�r?QE.T��8�(7,*�Ej�vx���J�ɽ�����#Q,��Y{h��3�t��6��Ҍ�M����4��ڧ�G7D��2�v�l���z����f�6@�	��3ĿM�����������S�[��:�Z=�󥃂џ�8� x��	1_[[�b�y��D�/yԉ�<C4qv�B����r{�����Ksx1��Z�6 &�ذo�-;_3y,�T[�Z+���{?`���1۫
�և�D?�P�F��/�z���#�+tS�fU�H��%O��t(�Pb7Á�9�`��d��Y�ɲ�i�����Z=��~��<=gi@��ё<RN$��Ǣ�fX�\Q��׼�fq#z�Vx'�ݹ���_��ކ������c˄�H�)��:lA��殿�����I�T׀џz7�\��U�>$�4��� �.X�c��4��X'�M��.P�/Yx��hF�0����ށ@�I�J��f����ͥ
Nk��(\E�e�����c�	��Y�G���1��0�8����M����bAϙǠ9z/G�$�
�Ltey���N'�U�C���l�!���P�e�r�.�eɑ��w_z�@z�����A@v���#@~L�kS���Wl�sY��T�,?x�T�$93������-uS� �	�N֞��e����7�d�yt;4Ĺ[����wb�P�������DO�-���z�X���xh�+Vپ��p����KS+%�m+��g0��+"L���[������=���L��4�0����&�d��������>P�E�㣃����ک8���Y_��l�Mb}��<�3M�Rm��N$`J��R�ݫB�
G�F���@�j��ŏv\^�'!�i�4�&��\�r9�u��L�S%��3��7�z���/iT
�^n�N��ҫ��3�7�Jy���;iOڤ�$S�oc���*��݅v����yr���Ҵ��H���۞�SN	޹��a�uZ��t(��o�2�8s�@{��,ѫ+���>�^`��qr�l�|��_���޶���<�E�
�ơ�eq� ��n�|�>�X�\��*��5�^_e�"�����z!O�1�wx�91���dI�	��l���?ȌF����&�I3f��T�b:�����^�\V���+,��F�1}�4W<�@O��Sx��,��ߵU?QD�4��)���岎1�5@��l�����_Gl��	e�f�}a�+�j��*�*�;v�G��ǆM3C��H�A։�����t�jΜ���uf_b�����j<�N������^d�+r♍!b��#"�Tb���~i8HB��=�{�ԉ�>�|�KnR~�\��+K|"�f0���tU��!��a ���c���� ?�7�v��4�hSq�F���P�az�x���3#��ȸ���
I�R�����\i>~���*#�ܜQ��t��S�1�(�� �L\Ɣ�]m[���r���˰^-F��~y��T��D�S��(��H�*�F�َ�|R�n�0���w�m��7�,�g�|���_qw������|�,����1[������3oB~�u� ؄q}ˠ��zG�׼.9$3�Uc-|1	��wv��/��kď���8�jr��>m?�ߦ!�K�{�t���7��>�F��	�;����Q� #+�F�	��'l�s��V�i�*9}Q��
�!O�u��#�g|Z�T�G��MF�̣��;�+�U��3	��~��WO�v�����m�8���g�M�ǟ}	*�[�rk~��6a�RhN�k=G�x���b�J���֞;��X��0ӱ��Ha�'����ƶ�eMu�'�&
�Vn�\v�D�6G��Aӄe��c��.�F���Ϸvg��⡟�GA�}�Z���
����у�sq6V�͘\A<��չd�=���p�G�(�S�8ÇjqG+��
�VIx�g8d⟵��zO���h����5:v��U�x(k����ln�⑱R+u�5�.��޵�@���R~ת��QA�X9s���vh�l����~�y��(3�io.�h:�5R���@SFÃk`�b�=����+4���WҬ��o ��p���4ӷ͖����^>�N(!�q����0��$c�?� H"q�5�K~�	nJb���4��.��g����'�Б����Z�H����_Ӹ<�9c�({5�^�����$��RlǊ��YUi�|�G�UV�޴�܄$��7euI[��ef�Y�pMeH��ݟx2�K�υ)���5֋^vs=�x���ns#�'�qgu���=�rc��|Ԧ�G:eS־>�o]�#��1#�a��oȃʙ�@$�
�#�$
ç��V��:��ӽv���Uc<N<��Ǽܞh�Ə�X����a��?b�BW�g,��!�?d����(ׇY�H��Y�oRI�z �k7�`���.����H÷k	2������i'�m�!�G|R��[w%�%ZG�-��4#��<��C��:�%��m�9�(lY��n����eW����TV�Z T�? nE���g#�˗v*���si�j/j��WvP-��g�@= �v�Y��EЃ)hq?�8��#��3���3�8���e-��N�m&5��s�Y_�K����6����p��jZ�߳��O��w�jq��ÏZ�3gboы0cin��'�4M"TV��6Y�v |<ЁI߬'!�� ��߻&�f��X$�I�k|\�,��t}\(�\��(�7_J'����+�þ�'�ً��Ws弫�%f~W~r��3L�m�\����))l���N3%S
z�˫ 8�K�Hb�
W�^zѕ���>G�Q����3%CBƚ�;䃧������u�"���bd�p��'M78�\���F��ѻ����V��<�C��,�]�Q��[�#�'�����4q��]�ƻ�鱝K���W1�[T�f�	_�wy�qx��|�]Iy���"�f�$�"�<��'��$�p݋a}��zRL	9���/뽑s����x	��,�~-Y�Ü�2vʚQ�����n{�>�lU�I 0'�~e��C�oo瞍�Mr�U�GAy��ci8��H�Ă��!��z�`�;fsm����*a�}�+b�'�.r��D�L�y�
����G_q���dQ�3�(��t�
�ٚq���Iq5sj�T�W`�)���oRGcο�$����Ct T&�O:�f)��bG?)���#]��ހ_���T+e�l�0�<�K^�6�K����Z���1sl��:�8Av��J�zh``�Gݿ�;x�3C+��a�ϛH?'�vј&
������k���'�5����$ʅB2`v��=�mO�~Z�5�f��cԝ۔��.؛�o65����u��:bY�X�f����B�u��"�6���OT��9���xc�����F	>)����"��K��1���F4R��o���"4Iҭ���-�L�l`��y�M!�{�*�:����aG=�o����/&�{e(d�k�h�}�⟨s�Hs�,	e�d����b��LU79��ւN|�B��>��?1/�޵31�R���o��H=�3��K�M��V�,����A��'?lzt��6�[@����%K9�}���d<u_��*��?�l�� !�����B�Y��r�����tk*� �F3�/�����ty�m��m�.�_��,ǆ��.K]mf��(���c�j@Ty�)��;q7���
Okz�-W�*��Pd����<(Ax٦�fF�6���O�Yϝ�M�:���[�p�ڥ N21����;&[׳��&1"�ə��on���+>,��O�%mBXØ~#+Qڪf��J���rb������U?og-����ΰ�W�W�'+6�d�e�y;�N���"�������y>"_��B���qr������H����$��������(��j���lG�|���x�`�y�Sg�C]�M��	�A	����4Tb�%���}���N� ��an�q�L�_�~>���#��J��m�`���R9�Ǩז�m`�?��"{�8�,�����KA>��]N3W�o蓀8,	��-d����IC@������ ����&=���b����7�fY&�e4sM��~�K�K��ʈ�	I�=�P$�9�A+�q����gfK���ǁt��`�Y�>$���G&�}�MA%[l����)�Ig�R��)�e[&�`��O��͖��6�9���)	��{��x叒	@�X�̽�p<�����g��Ǡv�+@�=|�J���<���4�X�-s�������7C����N�5�}ű;ca%����l��}�?��q��A]f�2C�-bJm��������mg��בE$P���ע&����;�bI{�A��%��-�ci�?w�!`0-b� }_���whi'0�֡&�6�vO�'�#"��ۚ�Ȟ{Hǡ��:GBӳT�l�J;�8vq��q�<�T'8�#�鰾�a����z��>��T	����cLCq�k�޷�Ed5��M�SWj%���m�:�O��W�/b�����E�-l�����5�Or�ޥ>	������׸�[�x�As�}����)�@M٢?`���G4g�x2˻\d>4ѷ��2ԙf��[���Ep��{�$4�j����6��b��`	�@z���*�G�?�rT"}���"%!u�s���U�u6���/P����7f�r�O��z`��B[񲃓N�e��+��l����J����}�1�B��.W=��^k���ݕ��8��?�
X�)ڏg�貪�]���[-�J<Jj��$�͉U~�e�I]f���GoL9������!���u��ۥ�tPB��Z�oe����d�E�����ZS�� ��s�j+�]Wv	��ʟ@O��NY#z�|�o���W��\�����#�%��X�43������T��:�:A�\��t�{�/��E�
������K�����q���~b�,��������|l���m�Wt�Qf�b�4,�-��x/?���N�%*#��/ws:Nmד	��5���o옼��G�j�s �y�}'�[��$qHo�Ry���6�᧻�CB��c������p�f�z!C>b�����;�x	��$aN�@��~Kw亰^��ℍ95���oj��s\y��FϜ�j8BĴ�_s�3�G��C��drY�ڙ<t:�7�`\�P���)��&S�'+�9О��Oxk#l��	R?k�����YЯi�L�.A�Y���f�b����,(2G��n���4qI���I>����Af�\"/��X��Ȃ�vW8��"v!�s�����o�[q5����vps)���W&`���ZAX�#��M��+��l����4x���x`��-�ׄ�+�`���O�0{�yo�<٣9Own��<�E1�����$E.����t�5h)�B�EU>O	��z2.��P�}�p�
 p"�d��� E�b�O�K�ׄ${&�;e�l�VOv�g���l�n.1#��b�|&�&Ԕ��%���YA��.�N��|�l�����(R�@t<�d㬸�.AI�Ϝ����[}�����,�p���q>9A6�����;�\s�50�r�|���tmVk���d:5�`J��� i��<ڦd6�.l�������YT��$�h���|�+�̢Ȥ�;�o�Z�mU�>�E9,4�洫,�wBTZ���*Z#�h�ϣ�?)�˼�+E*�J��	�	�E:b�o���r zl�r�,r/0�{�-��=�kB*��cq۔��g:QG�8��U=>r"��c�lk�px�ό�>H��ο=��L� ���� �j��g�M0PK�,�ש�V�:������'yw  ?1h�c��0{�H��j��y�	5���E�Ƞ)j*���)H��-wO�	6�=��}{�2������{90���|z%(�����4#)��e�I&\zq:���ׁ�B����H"ɀI솱JFo�
*<�W(�~d�G�h�B��a�-�"�t9�nz���⾚��&�N�m����S�E�	�'w�k�ޛ��fm��}b!�=�-�)�fek>-�]+��2�ڷngf�:����0AEǏ��b��n�Ѥ�/T�E��.�a`�H�ޘ���U9
�&�K�^Ls��.�60�%�/���L9:�F~��	��u�}*�k��\��K�-��@qg������Drf��J�fW��&(T#bj�Ϫx�(1B���ߩ�[���nz�V?\Ԝ��	B0�7(ߨ��
�������������M�|�����k ��Ånu {�j�D�h�/��+XQ�������{0��xN��}wf#������J�j���0d+m%����#L�p��n�"�H��q��iv���vvP��E9be���Փ*B�aدOl�'�������wxc
~��,8���=�C��v�u����(ƞOF�;ņl�,{R��o�1C7��ny|v`m�Y��9 c�_`�g`�9�O��L���|��/��l�F�{��?VDc��ދ�{.��W-���$LE%����&�P⪹LykG������j�Rw���y_Fޗ��P�r����(�څ��l���ID#&�Bm�)B�*�>P� {��s�~�4QSf���y�w`b��f��2�`=�w�l#��4������"a\a��j�1�U��G*�������0W�b�ƶ�<Mf>ڢֻ0
�����#�b\O� �'tn@|�~�*4e@z��Gb����|	�6�,�Y..�2�5G�
	�~Mx!����e���[�;p�_��OT��2@�?�^��I�&{�ޅ�^�	!a��j�Ef�3��{�>	!Cq����K�4cW{���cG�yS�/!��6OO�[�?������ک06�"̙��N7��ƾ� +b����K��[n�;�G"�N��J�a�
l���&k����Z<�����Orcdӥ%�E�F���'{lT�����ֲy���G>��o�I����k�����"m�<-ѷ�B5WNâ�Eol��N��c
�V�K����ew0����<D^ƾ2�%r�Ք�#�*H�aT��аs���I���}����Wx�(o��Tڋ�$Ss�|�rB�m�MQ��!73ppH����υa��d]%ʏ��p m������]S� a)!{��jѺ��&}u�����T�V6���m@��@��_�ݳ�:x��&�ڮ[We��#+�!�W�}��̃�8����=o�s�b2�(^�����oǽ4��J����܅$�:��sd�}909x<����	��ꛦ*�Jz�%v e ����1�QhI�T�4��=ꤞka����n���)��s�fj����1L�Im�����Z������O�����G��	l���<�RBJL?�7�� )�H�Ʉ��ַB42���Ҙ`��-��K%i�?m��̖�>�|܁ù���ihk\f>N���A�$�F����� ������iE��!��Z��!=`���K����d(cBo�gB�%�ؓvX�!�m���-���:�Q��6�ߤU��uk���ڂ�~�[V�(F�fq���S�j 1�����"�::�k�'}jNC���n�ƥu{K]ė��Ű�ʋ���9��`ͷ����Z�S7����Ӑ(bG祤�L9ߗ��%eU~�խO�$�Q�:����l�LCA���]���Y<�1'�G���� "5*�����b�`���F�P�_�������=h��9�z�kk����0�K=��{{�u��L��oa���C���%:
&T��I3�Q�#&�ˬ0��.)�jʯ3_��
Ӟ�yF���d��8H.���2� � ����T���>X�����e��¯#@���ʤR��C�)W>J��e�.9��o��y�aDŢ�M'��Zj���p��Q��|��`����&�9�:���S��Q'�V�����l��H����z���`f������5T[����( x~�"aư؊�<��E�;b��%���5;� ��m�!�-$���\+K2i�����^?ge;����k��8_[�����S�&v��� �4aA��j;%:v��m=��#0y��4E�����7�^����D\��U�x�N!�aF7�˲q-9��G�`�5���X�|_�"����/�wz���u<W۹����9iRpk�j�=i�.�%X��"�Ϣdfo���(%�{e�(�Ɗ��4D���0���b����4������=��p�_Yn%ӒѢ��*Dzk���"�Y|�[��DyM�́`-�_�'t��I�rkJlƠ�1v�S}���'K#N�t�I��U���]̴�2!��
���5(��G�N'�~Ɛ��Č�:G�b�Z-U�A��T d��EE�U�D��63�Y���fbxgt�3yk3��ȞM4��\�9ni�a��Ɂ���(�ʂ��N�kFbLp��2�ubփ�uRv���;n���jKb�H�~0��3j���a��wd��̧�n�	~�Н=M�����JZ����&�^Ú����w.ד��+�q#w�^c!��s�]���_�׵�#���ɢ����*�,���{۩<����&�XmT��"U��}ٸ��$F4��y�TE��r�3�T
u��cH`� �sk�Z�)�n���'�kvq���#�;:t ��׫���H��I����\�<��$[ ƚ]$�0���I��g�-7I�[�_�r��_�7'�q`���Z1��7��w1����b7���)�!�3�$�rk� ͂���"������FB��Zb��U�B/�ڧ�ǀ�׉v������$�A�o���	o�����i���i6�q���4��>d�CK�& 3 K>�+�,ەkU�wޟ-�>��Β�y� �dW���ԸE=l�O'.��:�	���F+��XL,+��M0Y�7{��i�9A�MP��U����`e�D7u��l֗���b:��e�iM��Ѩ���M���W"�i{�^~O�3�]Xh�;�{SS����Ai0�S(����s�\�	s���������t�ja�U��Pj�;r�I~V��8�
g�Aw[ ?�O8�Mw�qΖ�k6�s���?�aw��l��,�Jz)V��P#ѧm�2���/����x'L���7 Y��p������aߦ4�{<<�ɖ=tX����6;8� /�����%B�� O�9o� F�/u �]�g�b$�Bt��t�ݼ�~^9��6kTaK �x��χg�'E\K���QI��K0���j����*_�"�F��9J~fUޭ��3�de>�� &[(T3I�L�g��S�;5��g���ݠY�	��ɾk�5�.����R)�.���'<T�"�ɰ+�:�ܥT�jѾj�}Ĕ��9}Pf�I���m�oe���x�W#t���#&�v�_M&�r�B3�A\�B0�KyU�J?ƃߖ3��w�~	0ejͿ�������1�7J?m�G�J�D(�� B�#o�"�K�|ʏ&V �V�g��s��XoF-��{qs�k0^o�߫�^Q��үd�����r!�9�sj�#���o��;�p[7���^�/W!��w����2� Ҥ�Zձ�J�7��j�[��9�h��.�40�����d��M��Cd\�7 s�n�5�K-��O9���t��j(9c2A�Tl�~*��gꝫ�D���}��;��9W`"b�8`Q�|�e�)n�a�Q�!f��F_5�>:}�I`�z�����os����坁�U:~Nխ��;�cz�G�3&#w���-��ە�<�����
3�a?�V��U�5W�z@�P�u`�7H�K��HrX9��P��5�I�V	c�p�ѯ�"j
��U��ܨ�v[fd��~���Hy1�N��$�͚���3�1���s�P!�uYj99�J4�ح�*�ʔB�ܿoM'.��>�	�ZN�M�Ƭy��&���B�[ ���:�>�A���ݮ�<.5JGa]z{A��>'�s4WLZ�"F���
ǘ�`����O�A���k<��(<&�y;��&2�:Q�f��,<��ÉL,�S�'�WfG$!�����˽�bZ3f�.��O�__k�x�M#��{X����-�>�&msK�6���Ao����d�`�����~ HI��������0���t��/��UYӈ��B��y�~dV��>=�!�֛?K��߮A�������Y�Z���a��/=��a-���&kp�Ky���_+9!ד;u�T[�%��$�,�;���bW_I�Ґ��-��*�qZ��dS�q�Gk�D���ǟ��3D���Z�#A�捔�*��1�n�(�r�8�iY�h��
���V� k+kL=o`���XY�;*\�n����6?���u>���"�i��ϊ���ဍd$y���I3w{o�Ɣ {{ ję��y3�K����z����F�Z�rHFP�f���AM�hwQe��=�w��@��-���aڏ����D��F���[�TB��!M��8��P���@/���eb�(�@�l%��zkng�[�-�h�Q����#��@�Ȭ;����4|՚a^��Eg��=���^�fEL>�u �4St��Y�� ��v�O"��֚쉫��.):������w�~�X֓aR�!ױ\ë��n��Y��w䞬]p� {�wEz@6�"�=���g����M�/-+z�@+3�3]k,;��� Q:�Fc�8�M�u�&��%�:�;Ն�E��{*��[�*���rT���W_h	��W)p#��-��˒�D!��n3A�M@#~�?]��=0�;����4����^���z�MӇ�u#rLK�ۜ0��JN���͠4O[�T|r(A��^���	��i%"{ׇw�rЈp�R\()�i �?ū���׋�4�;������W��wjy:X֝��V�K��H�7����2	j�J��KLZ/2�@N�(�P�D.�k+a��U��Q���=} ;D!J�9b���&�Q�0��
FU<^�k���Ⱦ��`�6�P�,D��rW��ܤi�I��-��M+����1/�7`nw�E8�:�f^���\'�J�X"��@�>X9I�D�)9Yd��n�?"Xy���Q�xЫ��/��(��R��O�˩g<���~��D����`r*�){�� I�[j�M4{q�ڂm,"�#�v��&�O�=aC�!�z-�|�u+���w�����AIuW��`�	��ܥħAf��k�-��
�jz޾!£�l$5'ߖA�<'%�����;�C�_���?�:��TA.����Z�z�	�{��[-��\�̅��`��E��D3j˛��0S���ۮk��
�}���%>�D����-.Q�*~��tBiI�� T�J�X��q3���#�BlG�w�H�
��Z����\su%��>s\a���W�M�?�����5`4b�wW�]�_v"<�F�Z	#���P�蛐/�)Jm�>��r�����-�+=JU�v�[=���/��F9oZ�h���NzHS�$;٢F��=�'[K/��e��u� %�]�p��9ާ~�W ��)[iaɜ��Q
��0��yCPT��i�L(����/@,�F��D��i�N��'�B���r��C��&�,*�%2s���G��p�եr.o&�k�Q�WĐ4��!����⟉��`l���%}ezy�d���"K=C״��8,�5�Wn죧J?}�ࢌ�F�Ϙa�~�;���4  7�� 3J"������٪���:
���g8��a���º�uVm:�P�['�h�����Cp�dQ8�H��b�c�����hfgM��`1�3��1�5�>�]۫�|Z(�>
+���&���(D��� �.;�4$J�H<OU1O�&�M@"��t���)GOm�̨��ʿ��_���A;l6ڱ��p&�<P���s�+@��^�@)�WQ��v��r�FDCͧ�3I�*�<c���.Ӱ��O}.#���H�9���}��U�r� d�?��S�A5�u����﫷��1(�^�z���ōQ	�TxKc�j���g�6*�$"I��<'l[+��'����B%�1�V�*��x��T��{�^ci���Y7�6�π���:���v�D���]����4sH֠t�E
�:�zl���;��}���&;r$X�Ͳ�x��+��s�n��1.�^�!���*��@_֦�"�`�5��_;&��2��A�8nprw�xs�|�_���K\,N��G�<�&8�=���"�/�j�T���I˄o�(���M)\;y���p�<,�/�����B�W��{C��2~��
a�Sbj���~7F��-EJm�y���S)���%��4}Vh�� ������G&�E�QX��p��Ȯ�e����+�+?�|�Ȳ�hDU�1Uh}����CA��hgw+��B: ͠�z<�C��1�ug�oeU�وL�J�򥽾UU1�L�Ҹ��a�@N7������e�$s܀s\(�����z,>�>N�����$8��X����q�u����T�.��B��E��/N�P�$Z�A��ŢXQv�d�*(�s�Vj��*�0�S�9(�L�$*��=���	�E'u�]$��H�|�j�?h{ۂ��� W�� ��6��%�I��"4Xum3���
�M�+��\{�&cm�]�<�]�.d|:˿�GJ���u��F�5�*W9!�}*)��`$�\�#	��
��[�A�}>��Y�眭c��X��m�t�˱��0lc��(%��U��V��qD�Ҿdai4��>���ş�����w&\.���d�وu֥�2
�(ᮇǝ!7
�V�h	�J�]����+�p6p^`��\M��x��G��H�Q����#d)E��"���[w׈����S�9��I,1=����h����{���M�o�j[O1W`�kB�(���D~���~��`�Y0�?�1�W��ڡLr }��
�,�fJly�=��+[�"�M���9hb`��89�1L�p�-7X�Z�?���YEv=����2|~o~���3f�5����2��z�U��ｱhp*�����OTd���f�zi5(���&�P�����-�S�r�ĸ�yM��(�E��BSڏ�5�?��~�V��w�S�w��u�.�u|����U��킵眼H�Vb6CX����'���=g-
���:�7;Q>r����SR�`C��^B.�����\(�ywt�`�{��Y��%?�B����eK>�n*�(�G��E9��2�9������5��'wnfy�唑�s㿣Y�c+�ihk>2�I�� �2"62;�n,]����m�P�m�������{nJ��/c	1���M0Z��EJ	+bp��eF 3�^�"���nRI����(7@���pŅ	�e�}7���ApU#����?��A�y���-�|�����n�gb�S��
��g��yr���T~~���\���=F��z�X޵��`�|!�=���Z�eL
����_�jb����=6K@��MQ��񜄿=�.7�q\5�`Un6~t��`#Y���I�"m�cҳ5� 0.�&����R����{'q��ָP�9���~�M*�^��K�ߎ��y��2cR�\�5�9�aI��9
-S�>��\��8�%[������$8�-��� 6l�qX"�dC�U��{QrZ�ө0`99r����	 -�"�]a��\}r��*�^@�/���p|�Jj���~�rq��������� =A������ӫ�[�]N$5���Q��N;?,���~�t�<s�i�븲�\u�����I1�,ø��4�+$��h��m��UtȵU	����6 p�"��g�,z��E.K���Kz�Ź3��@�1�(D^{
�|f|���jElY�H��Xw�T�F��T��W�K����P� �S�+�T'�{�?jxy��ڷ&Cw9��?��tQ}H��@$0�*��.-/\�i�����ْNa�˧���:*����.G�%����cH��8�����`�����<�����;|_+��=.�dɖ#��\2b��`�u��;f���%+n�ޗ2O��	 $Y��(U6�����y��=�Y�7�i��)F9j�³���箍���*Q�����v�g�6�㸿tU}m�^3tE�r��N�Q�MC����[<�(&c� (�F؄0���2��a�����>]c�0ޡ,�$ʃ�'�*�jb�{��i��t�o���(��C�8[i+��(� �����q-}k��L
^]>�����+.�
�Δ۹#�Yu�Ω72�~���]-0>�Y��.���sh32����xEY��]_M���@V#Kt�w-5�7�@g���@Aiu����/⻦Gj��$:�,�a�.��[�x5뚵�w���,x�h��16}s��Ba��_4P�����\CS��9�{j3&����Qo
e�V����?�]���\D컟ڏ �X	�5�W�K���O�q!툞obXX�/�x��H�J�n��8��?�N}@R�̾P���P�����
oq�e���v_s��9J?*HT8�cѽ̞]������Xi��+�UUH��$H�:�'m����eVVY�o���<N�0탐>�1 ����4�θm����S�!/����j��U%H�T�Ib���x�_�U��y��4�|jd;��8�@�C�ݞ]o&�(}�����b��
�����ubL��9ހ娰Z���J\�!ß�D�e��,3H��Z%X�� �Bu~:��x�Ìe,G�,	%��lYl�����KW��#bY�0��I�S(tѮ2��}^�s,�G�6�iA����3eA�Dv�!�{��h��3c�/Q����fz+�!V� �*��ğ��{�����i�eu�{��25)���R����z��̶ib	h�K��G�煭�� s�5�ȟ�v�^xt��o��_I(��C�A:���o\8~QU� ��>Y��Zu���'����	]�X��R��ΜCHK���6�N�(v}�V��m�.tU��yK�=�5)�ū��C�0�e&���%�͍���赣�^�x��!rхў�K�U��~d7�f�I)ي�ciP����N��,A�_<����#�,OQj؆�sX�M����FU3ߜt	]�f��X�C�V��?�4��m'F9��x��ЕFS�Ĕ�= 8TW_�?o�=�e������ͰD}lߺ���.X�>o�^�;�3|n�y�)���h��*2�JޕR����#b�Ԭ)"40�%ﴑkly>T�ϖ_�EK���4NQf2��ĳ�%*��"w��j2����NS�����#A�k{����|"���r;7�k���!9�e�K���~�Z����?�HY����� .{g_�#LA#��ϒ���99Z����Ǔ��Iԧ7FɴÄK�L���j����?D�0�ܭ!~{�����h��5�dmX�Y�j�B�>��E�NI���q���ی�[xa�{�ؘ��W�n˅�cY�����ua�������X���N�G=�����d��j�S�*�`4ɂ<D"���uQ�#�`���ϱ��V�)�<%�«��D)�1�'��ր�v{є�T�8�ڇ�_�?�uz����#K:b�Zna���O`�Ϲծ�;T��3����"{��~���[�������XzGL�ݵ/��R�R���XK�ώ�#��i��ot*(պ�aSM���^_�� �_7���Y3%ݮ}�?�z!�ǁ4&�f���r��]�gB^+�-��n^���RA>ϭ^���{G|�ޖ���x#[�~e!>��g(�!rMM�����O�_��i��%6��ѫ�}�5>ɒE�$ɐ�36U�6��W��lGܰ,�?��\�F���VA�t�f��`�0�M?8�=���0��4�s�(��4�B72��Ft�?T�	���$�W;��'�*��ӓ��z�Pvj��Є�L4w�Z� �d��ۗ�@�PZ����.�67�4g��q!܋c����3�AH?%�!�b�u��X�V(�׹~4����w��.����i����W|�^�4�,��ta?�]u�Lף]=��D�8_Y,t-ɂw�6�l�g�8ia'����~]6���F��6��z��>� y�6em7�ߋVW��ˀ��\�눐.k,�1��eC��M�GNv�
�]t�n܇lT�P�O,nY��S|����>�S��<��E�*3e��:�t��a�_�fْ]�Zߜt����T�b��wb�cA�g��q]S�Q�4�b��h�84�)���.��adc��؆��U/`���[$,]�C?#�������3(ޱwhZ?��S_r�ř(�C1��p�2�?����cW�J�GQ�������C���'5�}�]�+W��36Q��>����"z�c����3+�o�h���@r���%@�\76J�FT�:�z�Vf��m��᤹L�P�L]���-j��P�h���ob���
��0�B��8������y2=�y�f	!^�R�Qf�?Ľ;��b?9�4�ؽz׫7�te��Q��Q�����/��栮9��tK�_�9�KG҃�!A874(�Ѣ&�<�%/�����p�U�h��|'a��漪� U�������x����Q���պ��S_�M���W:�J��`u)�d�����ѳ�@#?�����5�I�p�J�sgڗ�H����j��&�پ�.��|��IZ���pR���WK�R�4�-�0�Ӓ�>X���U�|c\G/����u?��q@J���B��V�[Xf8��ܚR���DZ� # ��X~�늯�:�l��~?�T�HQ�1�ۯ��V�Ԕ8�2u��v�����ae�D���j<דX��$��p`/�s�P��\,f����!��8@x'�)�,L���Z�������lji=�����Ə�����r�o���k[5�g
۱�G8�����.���z���h����Ã��h-����,K��b}^�x�<��\M�\�t?�6��ߪGXn��+}6�N6l"�z��c�vҋ�0�o��T�~2�/:�F�<՛W�WD��c���y�jO�4<��o��󮋢6!��|�A��+���TR��$�pf�j}�o+���n�6N畮Q6N=�Q�� 'v��$�+���e^	��Ah��ӻ��?�<ٝ^;�@�ُ�EvP���/�QG�s�Q%P�U}�D���ob����=A(hw�Z�3$'F��cl��^�kN���X��e�Ǎ���Loz��i3ը5��������i����܅??ؖ�{�ö́��t\�z��1C���EO�$�aEO@���Y����i�2�-T`�8R���5\�No���J���-lj�wږ�Қ
���P�@sR���F�S��:�@����k%ͫ:)�=ȁM�g��2��$�Ł��c	NМlaf��\�Co&7sQ)�;$A������@>[��N��?�Q8���Dױ#}�12 -���s� >J�k���x�B�����* ��	��lp��5���u�Jb�������jZ�*%xi�Tv��v��{yӉ�9BR�O��Q�,*�Sd��!
�2�q"��5�'Fb���U̓_��C�����\$���%s)� �`}��c=�u'�1�����l`t01����`��I�V�]&�&�B�ҋ\B/�
���۶>�u:A�Ϋ�-1_ڦ�T	t��>����0(�x�
����q][���]�c�mי2�* �36{V�^��I�7���/޻��-Ѥ�+�m~����Or�b��_%��ۍE��?*+Y:�����v��v���HI��'%�9/*B�a���p=e��^�(�O2,��	��J���	��`���ր�PDj��V��Pɧ"�7� ��n�0<���vV����bIj\Db�|�۾͐�lT7T�w2��8xx]�[�N�'!�y�2@?.�mQT��D�V["�"��^������.��ٟ�����@7p��h�&K?���?'A6���V�m�{eM� ކJ�;ӸY��/��%�;"#����.�֤�K8>�@�J������6Yi��Ns�Q�~�wF�TW�AB�.�]Bm�5Hu
�c�eg��E�>�~���p>�a�$N�&G.��5��)���YU����Naf���a��&zUh��QC	� h>���z8IҎ��"�8�Fl�^h 6�n����5,U!�	�4u9R�O֞�:Z��}}�}[��}�R���U�T2�Y��c��e��Y�g1F�4n������I����~`��)HMv������1�c������_���� �2����U:I\�}gw��E��Zd�y�DEC�%ݔ��W�Ǧ�U���M���A�(�cKb�`i������g�T�yהx78�iԙ��(E�>�U����+�}qP���.LzP_ð�&�g���6�F�}����&Tߍ����&i��<���B9ɓQg�4{�u��;�w[j ˺��1�(����r�ru=r�aU�c�5���v`�����BC^��z���Slf�./�������j=}lB���0��SU|��*�0�Z�Ow�v��7D��H#k>�;H�]d��g�\v�����Eb���ј�9+�0��#6��ŕ�h=G'I�ߗ_dWK���n��ꮉ�K'⛱�M&�ċ�~9�Ѡw@TGx��KT�o�k��t����a��'�_�L	�0
I5�kؒ�Q��sUr��c�8�s�0����2u����qR�
�pLAN���>|Wm�� �RI�*�s@�C��l�C�;HBcӏx�$�Jb��h��3ʉ��d���9�嵦dz�35��T�Rϗi�a�w�C�F�1��?�0hR�o��g�MC)�V��TW�8Z�v��$��c�g��� j�l���*
k�Ԕ�G��y���.��e�=7��[�ux����^b.�!Z��F7$\��k��yb�nM=7��Frb��B���*��PRk�hʒ-��ϛ��/}�Z�A�=�⦰�L��o2�@8s�	��m��K����a�XY�\?m �<E�X��
�Z��c�S��juξ�X 5F�������5����&��mw^���!LPs����a�#7�l��J�+u�i�B��#XF%���GD��sߗ�2���!���Q<]za*�����&����!g[��f �����q�9f�=��E�o����n%��")��)z������Jjy�{7B+����q��:���p��
4�p͜��,�G-��Ǹq3Y.^�*�½���p�P�S�F$a-"
��fN�9��|m�:�b�8�[��C�jݥ��pи=�ɩ�1��p	u���g׍���26K�y�7b�=c�X�0����zh����eT�A�ԅP�CUptȏ�V{cw9����)D�x
���BA�R�k)%�:�.4]r0�>t����sD�N$J�\q�^��̖ 8a�^6nA��|�xW�V�� �I�G���,c.�6�Ϙ�0�s�0�c�N-_Q����*��=��\���Nmqߝ����R ���	� 阋�����Yu� �G0JK�G~���LU%���?2v�Z�y���|zx��.N�˼��e8q'���%�w�|�u�[s�b�I1�k���K����s�栤)/t�%�T�zL�{͕a�r0ϑ�@ah'��>Kg�<D�����Ai,@y���.m������>N�g@A�ծ����Y����,�H�\�u�}\F$�d��r�9i��5�Vie���3R�;�d�[^V�dU�
��h���Ep�-�Ui����a�r�v9�P��g����� j3n�E�_�E����׌t��RЦ*)~�ɛB"BW`x�!�P!6���o���[P����I?�'����Q�/�o��A�V�{z�:�˶�c19���k9��ۯ��:ƅj5%���TԲ��ډ��w�4.v	}�G�ǕNf�}b�x>.�(A⏘S� ����������>��i���ʪb`?j���:.Ո���%�-�Kv����;QA`r>4(1�ۏ�j��{5�I���X���H���na-������@�Z��9�YR����9Y#��W0#9]3��|�Φ_#m��k��sd:�)&>�q�C�<U�[�������C�x��fBX��1T�@�#������F繋�f��!=U���ݞ#=7�`<�O����Fz�u%�*��b���^��_���h
a���cAG���4��y�qr;�v�>S��s�hd�!7{n��F��C��_�^��.1�H���{�u3c���c�R$<4�(��r����Mà$��Բ(�Q���G�"��=�𧺖�D.����'Ʒ$f��[�J�ʶI����~OYhjU��y�
����+��"j5�x����t[*"w7�έ QM�5�,pb���s����q��ۃ�H�w��'.�������Nyl>ƪ$<��Z�eI����qa��bh��!�6�!����B="Ct�lQ�xA��k����*��c��G��3��3���_<���]?[A�h��!�%>t�rG닏~nw��g?1�~+��h����]%?ܢ�tE�Y}�q��?��?tFi*��Ca[*��ۗ���LjVA�CS*r�mׄ��$É�U`NNz�g{����S�,Z�� ��Ew��է�\M���2m�׍�K��7)-+{Y��Hұ��P�(T����z����'2o�_d��^w�=n���z?��nʰ��D���Y���-��]��`��ކ%�u�v�ؖi-9V��4?�(�S
�+~� �����q������ᷩ5
�-�棧:ǲ|�L���z�������;t/�Y�ǹw�K}ޏ�vT����X�2���_�g�G�	#��-AN���F
�׫r���F�	]��UWH5{ICN0�#��'m�ȔTQA��gn�@�Zxx��>I�	��ͯ���M
]��n���!�OD�E��p����hY�y
k閛~�Z�\�ÂK��W(����<Z�:���,eZ��v�qh�:p�Y̳g3�y�G[�J�=|w��	&��f�_�:pE���l�$��i��-lJ��W�_��RB�,��+:�
�����Wg٠����PݪڡG��W>����_�=R��Qt4~�`����A%��?<_����}4�1��&�O���z|�J(f����s�[���j�+�-���?�RIx�\���m�R��#�DN���V($��	B�}z ��b�`����R.��߿��i�"��̶'��:�ŖFBW^d7+���f�-a�n�d����+��n%]p�����eT�)T�L��X���$Kㄻ��B��y��bܾ�?w�{����Q)\��Z��d���Y_������ؙ��%� Y����L6���=���q8{V1��0:�������ɠI� ԭ��+�ؘ��B؈��0�9��5M��ٙVY9�d����Gb�P�}��;$b�Gm[o�/��e��p�CeD8�>��"��<%壳j������>�xe�xx�:Ξo��!�WÚ���Zp}�$�Kڿ�q�5�|?�E��>��o��\a�)lp	Uc�<{���z�%�9��K	:W��}(½��d!��6�t�UO��A^�b`o� �>uh^ƎF1�7�f�VVm��K|�4&,����V���j2sU,�;������BQ��`���W��5�,Xc�p���`��z�7ç&4D�-\�7K��hG��h�-詝:�����u���d����Ӿ��5���p�|\(�ĂMQ��P��]!Bc#)���K��/��۶�"�4�%��xө:�� �1,���T�8=�y��n�x��,�LK;u����G�F#�|���������ʄ"�>X�����:���n-����`ƒ+A�j���������= >WΦh�_����������X��*���\��g����Y���垩�:������}�$=��� ��N��5������y�ZR�HT�KP�bq�t+na�bo�� {Ē�������d�U�ۓG��1�A�痌	�)z��nQL��~H��e��:�=/љ_���8��Ж�v�=�G#6j�(,�U�K�����sD�t���D(���A9�q!��
�E��iʷ��`@g����G�Gy�7�'U�q�_~ѳ�%�+�}���͊�����%a`B:ӻ	�_V���S=��� iﵾ�}���/�B����{A�S��US*1	�kt����\��o�-��?�Ux���E��9f:��{�[���
�z�l:~���-�j�̔�I_�H��H�i�7#��o�2��X�c����Ə���{ū�0�*�MaqVJ��� r4I�w����&Y�ݢ�ޣ�����j
����7*��n-��A`��o�]�c�]%�n�~��n���H�S=��5C][6�Q�g��VV���D�1�s
iB�Oz��w	�����̄�D5�����a�[���:��FX��+��AXJ̠�n�b�mC�4K�'C��+=�I�ژ�eEv#�!��8-EDZ"OG2cy�ז�� 9�4*�w�ǁG�@lU���Z$�����ץ7�y�HzS��Z���&He>�n��)�4�q�3Vw��ffT��u%s��ˑ'�����u H�@1�.�z:��o-`yJ�O���Pi^)���g�oX�}�oꑦf�:ֹ<Uw��z�Ϭ���c����h�ָ�?��?O�>(�H)��Uҹ1@��y�V�P�f/���%��x��j�w�#S�?k(Gڽ(ח�i�7�T��:�QbO�$��F�Eg�:�0���ͱ�0��๬F���w�fC��s�3�✡��K552R�u��l���t�_U�h�I:�7#]շ���Ȉ|���4���*oB�c�B׽�=�|�N����N:}P�Cv����T,�Ϫ�-�$2�p���?�k��Z��[S�N�[J<rJ&mM8\� M��L�h�k>�5�Ё��M;�i�>)bo���ĵ�mSe���g�PP/��G	TE:��T��P��Y@ٻu$������q~���x�H�I�JB�qgӐ{A�|�W9e_�@"0��΃����bK!;��ӥ#�l_)�:P��Y?���r:�O/���2��Ѯ���>%�4↕���0q� Huѓ(���Tk��4)B��Z����'�^���=�w�S��Ɏ]#^���Gc7V��PҞ奃]l��cg��j ��)���B�����^y7��v�����2GhT et���@����1���I�s��+��Ȁ��B����a�!ttTY��Q��?J���u�\Kc�a��$Vp�I�f x~,���	򻈧�P%�GE3e _�v3E	�WEjk���$)��Av���~@;Dm���5���mm�����lOR��,8���� ��AZ�����
��z�C�黃w=�����I��'��\X�����TI}tH����
�u�&\��J(�-�,��b��B��^ո��$HV���~v����z���ק�&�ˮL����*/^'����]2��||6��P�n��V1WY��4��� ���9P
�������U�u����WY��̤wZ�M�����ll��!�r����fgX?��&�� S�e@��mF��KR�1_��j��L�|Y���%ys|]i��P�}ڙ��:x�N���&���1~;��F��z�FO�K�!	��.�=	��dQ�i%U���}�{q����f��W�\Iy����< ��k '
k�qj�uŔ6�y��1R���A��h�R�K�]hl|��oy��nݦ��6����Br�4�0@y�����bl�V>��ނX6�h�\jr�����u��k������=�f/�Z ůrRK���}pom��n�<�ZoTb���R��� �=9��/U��J���(/\���3�1���=b���T�N�.x�!��<>�B�BQ����kf,ٹ#�9��#-5�
"�\��@�����'LM�\l�U�G2��1�Y7�fҫy
=/�	[�ي�Q�h�s�_&�<+)��x�A'�GT�ظ`�=�h��ƕ⅀�)�Y�G�2�:�iE��a蒩�A�<H��7�'�'��n %@1����{�T;p�����ؖP�c���.�Ph�z�٬'yq�����SIF?��� �#�w��b�ĸ�@��T��im>h �ۻ�]�2�[,�����kL��3�"\�m��¡t�$ ��SZ
?���B�C�*��V�[ob��'�3��6�;����z��&:F�=iǞ0n"Q�= ���=V��wr�XL]���|E��瓥�<3�J�	� '$n��(�Hz>��daE���*����ٻmd�j��x���,�Ds�M��W*nQ����\���	Urm��Ô�V ��Y�� �.�"�L�uȲ���2hJ}5x��C��Ȕ����)N�P�!b���/�|B`#�S��)P}��Y�8�Ґ�b�� Xw����h��9� ��ܾA$��qU����N��&��F��3
�o�{6>]��q���o�z��.MX_ᔽ�X�Dɉؽ#��f�����x,�}B݆>@S:U��;�Ǚ~�����4dfJ���.a�H�P�� JH0��5��-}Yk��"3z{{�ٵ��_bb����nm�o2���Nv�	�mB<�Q]Tؤ+�1�'m��Wxaq:�	�w�ϐ�>��r�j��n��a"G��â�A����)���,}����$�OL&b�H#6G�f�������Io���67zzk�VU���Ыom8�����1��J���N)�:ݯ�h���5����?��m�V=�֔�I�����>0����7W����w���u����h��˰��-y5����ƈ�-h��32I�0����K�M����&�ău���y�P{"���:*0�9�t�I%}�¤� 0�3\���J�P����]7d�^Ӡz��4̷Y
�Zbg������Ț�c"�@l]���ǃO�V�� �g�g���f��"�{<�%�|!����y�iZX��n�T'Z+�����ip��.��JՋ��v�?'����{Uc�{�g�k{�7�2Qa
�m�S�&��b雭!�s�B�o/�j��V��"�w�6�6�o�~_
���ʎ�O)R4�tȈ�qYB�O|&-�-S�5���"M�A��O��n�.v���(�-B}�����W	�c���oUrq����8��4r1����(�rC��ik�}@���BnmvA��EJ5��Wbj'��3�w>�h�װ�{W*���״�W�������RY�v���$"�0��מDJ�kv����ǚ�Zۯn���	X5�� ���C0��#$k®�k�zz )`���J<�#^�/,�C��mO�T�%�����,|�~��؇�v�ǒ���m+s��XS�D �k�_	C�^�C�%���$���_���MZ����N�^�����"ߵ�?���}�����A�l���BQ*֯W��V��/Cd�t���j�YDjԗPF�@͓��$ٙ4���!,��W��� �n>I5ڣ�sz!�������z���um	8݊0���χ��5<n'���{�J��.1�K��fh�栰f;��#c�0����O�^�2	ٍo�؟�W�{#��F�L4�o�L$"�����	�Mf�z�݈��F�'a�n�$��Ms��s�/B�?Y�Y����HG̟�����+���I�{9�QF̍�i���J�mÎ*�H�}��Rwz'����7{�;�yt��G��?��cM���W'�C����
�Au� ��{�	Ek���Ш��Ip�̴ �xV3R���wDqg���g�MNd���X�ݎ�� �!�)���M��ޫ�D���@L����J��>f�oD$
�.k����Ҫ%����c*�j�k87�����c%?��s��L�{������ĉ�wo2�?uszn���f�#It?�I`�KY	�o�j��a7 +%�3c��O#��*� V"�������V�p4GZ(�['�B��ҤG;�x��X ]�Q�n�I��E�A�<�Jn<SK� ʡ��9��-���c�ze� �9lB�7�"u=�荦�A8�}p6��	b!����
��!�a ��TkP���e�Π	����S&H)�E<�߆��l��S�pyHF�����0��ɢ�4�)�[����q�fU�Ĥ�J�B��D����?,��_�mmP�q�4��)�q|��?���煙���3B-��蹢���Vu�_2��}�Q��|���1�Ј�g��կP)���A�܏�~��i)�������pk�zw����]�|�O�����Jӷ���^@'~��PC����(�I�a��;AĦ�i����*���ow� sy��{]=i�e>��B���&�J|��*#͕x 7��Y�%K� n!��%�u�����vh�����MCu}θUD�Q3��×�,=ݑ�{ �ޟ�s���4v�r���luo���~���E�m-��c�~�cu�����i��yQ�?I��NK3Y���г�6h��IѦ��Yl�2�q,|jі��uO�d#�%M<K׍�k�;�����ӌ\�y �@=E��g�̫Axq���K��5�
,���+Tg�}�t�i7}7�f"NaQ���%��TDh�e�
�>O`0c����*����1^V�T�R���KK�<m�F�Dӿp8@0fb�H�O_a�ï���X[0ѳ62��QY���%���':\�|F�*�}�E|���.v/�+D��gր;3_�r!}m!q�F��fZ$��1!$ǭ��S���!��`�=�ǀ���!�:t�k��D��+*�)�q��ES�}k���>�?a{3�_�IY�~��ə�m�%��� O^�U�x
%���D����Q;��'j� ��i�d��T��^�:��u*ڥ^�=�9:@�߿������/b�l����}�6�#�<���F�T'I����]Ă;;��e[{z�%&툦ҟx�m:J�0W�ST��vȋ֕�]C^�WN$�'�������H����C��ۮ̈LR�<`�yVa�J�9�����B�����K+��|�U"SRt~������3�<��L��6e(��ˠw׎E?P�a�^C�U�P�ӱ�Ӂ�_�N]�Y���,�S\�:�]���ŀ98\��jSBc�&���R�2�F���3��b\p5��E5��f�	l�ֵ�ٳLP���b�W�t�LŤ�$M�΅�xYG�gZ��v��u�B�KV��.�U��`�,�	Ɩ.m/�|%�'���R��"����/?�T�(%��}Td'.6�n4��Q�{E�t��bha�k2����!�8��;ԙNY�M��d2�� `p�ĭ�kEx}�����G'\9���]�3L���H�.1,���=J��t�^���Y{]c�� ԖkrUl�|�V7.���-�PhLg�I���9�$���Sɑ��^,�?O��+V��A)����9�,살��o�w�XG�m�Ւɶ�&��ǇL�#e���ITL�����*Ѭ8�WY������!y��`J]��F��mZbO,��0��P�`��+�r�n����
�R�����V��*4c��u($��x�b5��l���6ę���t��O�R��$�_b*5Q���tg��`����G��מN׻�~Q���k�%�`�v�\�Z�^T�d\\f��G�@񐷑k�"�ö��;�������r"R���}x����Nyn:ƅ,��8Q
m�g:��!�{x��H�n�"Rp(��l�zٍQ/kDx�FO�a�|�9��g������ן����0Q���ɖ�%h��==�m�Q7k�!�ڂj�v���w�oX�e�mY͛Ԧ���fD^x�@%\�2v��%��z�J�x&�M��w�kC�(Y�-=sb{1����0Fm�{�Xe;�`�_$�����p4�i�S`
�դ�&p�8�S�2�H�M&[�1⨝�ފP5 &(�v��#Wsu#"*՘N�S�)���ER/�ݟ�F���kjg�)�Eo:�}�Y�=-�Y��RoHET�.�
���|�"�� )�$G�����M����D��e/���/1�Y�P���Ԙ(��B�C�X>Fx�B�L[��!� #�w"ȹ�5=��΄��.Q��3�%\����C�Ec��j���̋4�c��JgR�Y���ߥ��(Ҫ*?�;3�Dc/���^���[G�Mm��n�~`�c2v�zM�̣�UC�_����)�Aٞ�ʗ�V|�������NX�g�B(T�ڗ�.�
7�Fpr��k<a>כa���]+��p�11�A����� �[��q�	���OEpG�Q.O@a�������%�g]�d����)�i ��@����u^�*#�w����h��X�oc�N��bn ��[�?q�J���>t����m��3��V�is �PamuHޢTuZE���Y�4h��R��uIF�#�=��@�q~8z>3��҉TT�Ձ�7cN��]U�|6��UA�yƯ.��G�GG���G'�5#uظ��1�}i�[z�;�{��dq�˺?����d���N\A�bI}����\>�t�oG����| 9�I���P�~׶`RӶ������� D u_�C}����~``N�˱[�-�`��_]<���K0-��z��^�Z��k��o���MiQMH��<Dъ�i���x;��x����E4�j�I$u�Sk����0na�,�(�@#��ф��|I�����^����u�6����y P8̪j���t����N-�A�5���K�e��5�`a��|�YW�|�a޽v�-9�6�V�q{�4P�w�v� A^�4=�x��v�!#�cy���/�R���L|�6a�9����=�rP��n	��V�RKd���*f@l�Κ�1��5�l����Ј�<���>~)[��L�hv�u�X�ª��iv��K�`'�A%|��GI��>~[QN��F�>�Oक���v�^��8�k����4��?�!�DB����Dgp�ݷ�R"S�;��[��57��6����Ce
�٤�e?.i���K5Dl={J;pg��Iσuw`J�ꯉ
�߹U��38�qMA��q˄&���Ki=>,�MJ�P����uT0U(~bpQ�l�rC�+4i9����I��MH*O��M3��i{�(���EK_�E�9#g����$���Ym��ݴ��^��Ò�)���[0����r�����C�rf��&|b_U��ׂu��2i��@ϖ��$�yr��@��:ȿ��01| �+�p�ι�ju�tҠ��Q��~��v[�Z�-���-�291
`�,L��~���&D�s��p8�W��������u!���l�D2v���1B�_ڢy]<20:�d�؏Px[�1��L�#�]��LM'��ێc1[�և9�-.(�h�Y��j�͇(&6���s��Md�c�w�Z:c�Ԡ!2'-����q9f�B�	�)�L��o�\�P̿��16z,����o7kZ�D�ƮJʭ��DL*�k}���򑥔Eڡ�����b�� 9l�	^��%9�<�	}z�Y�~w�B��9]��Ɍ��1�u���I��t0�����a,l�\y�>��C�!��hP��s��O�B2�㨩�8��j��
 �s��pʜPl����ơ^aL$�Ƙ(.6�ĥ���54�!�����!�QJE�zWHW(�	����gX�}�s.�6�S[5���(Ժ���]/ƾ���z�%�t��;������>ʐ�T'*���3���}=7ౙ�_��ΎB�'�>Է
;���9��S�w�|~�/<8P�7��؉�:���0+���s��t3)@FbC��FF�/|kI�3(=���2�v�7�O�mκ���_�,�|{P��}LE�����
f�8�I#�d���>l&���2�H{�W����[n6A|�ǚۮ}�0,vy����{eZ������a;$��ΩF��s;X��V��z�4)�`hnj��Gs&�ޗ`>�]?t�)�1�YMTv�P+=���.�5��R��% �^�Ae���K~)UN����Ũ=��l�h0[��؅�Q���Έ~�8Sib�f��S�r��l�&z,Y��ƾ�bq,J="̊�<R��>�WT��@�OrT!ϵ:Du6G�A������\��F��P�r��@/B#�ti����AZ���a��?�s��$W�e�=fY?�0�?ť�����h����LZ�B}��l2��]�����	�O�^>��pM����z���~��'��w�q�|��y�#�ϔ/?��bT��$"KVW$��� Jp3U����ی9P���k�^g�[K1`����
.=]&0�\�Լ�W'�@����K^���r���90L���!^'8������儡N���]��	��AK��f��d*K,x^�1名!���ԕ@�ޯ����wBEp��`��n�ݪ0�S{�~j!�&�n[�3ƑV�5�|��7�qR��|�O��r@$P�G��_�DZ���j�P%��L��Z-f����,f���ա��<$/h����/N�t��R��#zEjȾ�ϯfF?M%�� �̄����� �v�=u���l݀m�	�tH MTl�c{�G	�ȿ��"p�@X���ӀV�=�u0�v3�xv����\���`��Cz�I�=�ö�u���@f����>�s�J7�'�N5(����^6�h4�`3���kM:ߔ� <���c��R#�v@������y-��*�?��~�A���!iM��ټ��J2�Li�pgB�J��B]�?��s:H�w��{�O�Oݷ�.��\h�~ȃ�:�#Ư�G�,�rZ� I�)�0�j�����Jc��gK�lv�y��!\��fh;GX|����?�M2E�=�����S �!��=v��޽b?�9%�7�3��t`ةi�M1L��v)�ᶳ�C��1�k��P�L��Xp���w�3���PfJպz�8�̒�;�B"�������T`�]n.�j!�<$�u��,�(�j�G�)�jMZX�S]���aq��# ����K�e�G}�R���mn���p���#:~Gi�ݍ|��D��`EVk�DIO��R�Wu�qR)�'Wq��I52 m|�t�`��TL�,����>գ5eX�EnqP���:�D�k�BH�V��j�SE�6��I\�BtVc����!a ���R'�գ���P������US�����$"��۷�V?�NO_��e�֤*�{�j��}pvH4O�ş�Y&ּ�S����~��|��Z����*�r��M�{�x�n2�:�XGڄ��JR�-�v�KQ,�����v�j\&>"�$o &ʤڤfbi�h.�Dկ�^�2w7��
��L�R�����o�bˊ?IQ�M���E-;��N �2��̗Q��ca������7r�7!��cB�L��N6 E���տ��T��0V%�$���h(���2�� �5Z��4z�Aju���^ 0{�I��8Yn㥾����!����$Ǝ���@�:�N�[��r�w�&����"~T���Uڎ�I g��d`i(�'4f-�@4z�c8]�H�ׇ������EO������J�`_�m� ���߈�V�<i�(��l�����[}�~x6x�>��u�8ٍ���j�U��!?�݌�������*����`�����/�+����OH(X�w����Q�^ԫ2�6s�F����R�ab��=Zw��rV�@��R�X����;L�N�!�}ѕ# 2R�"���W(Ik��U'EMN�a�r�g����Nz�Q�{��n�=WṔ��j�B^�s���0y�>������Me\z���V�,�\F��U *���C� G?M]ÿ��6T�6�I�K!�5Ͻ{�]`���˅ʮ��̂>��6|�~D����� T�9��3":X��v�r�$��ޯ0f�KQI�����0Թ��	U6#7:�9�u���-�#�͚�W�����Y�;���0�!z�>�;�0ڤ��I*����J��K�TR#$���/5��Z����9��tV�Q/�jkb�n��_��3���D p;l#�����
�M���@\��j�h8�B<�w���	b�5�oY��ɔQZ�v�ͦD'},����ɓ������6Y%l����Bs*�´���O��*�Z1]բ�[�J�bXC�ͦ��&���FTNI������1�MtE�>קb�2*�oĐy%�T���6ն���Df�l�Cb��x#_|�.T���Ұ?R#���	gXf|�Vϟ6B⨣�X%�Pd1z�� �z�;B�v�JH�N���^M����ke�1px����%��<�],=���Տ9�a��T P����u���]_mC���=B��J{�C�=�6�3�+[��QrR�uDw����AʬL��l���p:Ԭ���bt���v��5�8��Vk3$��׉S�o i�W`KP�ő�3��G�<P���������MdVJ�iʉCW�]Ѳ"I�<ҩN�p+�8+����x�k��=�)��2����`�YxH��_G��ͼ8��$����U��v$���.�����f��A���@�n��܉DZ�������ӓ�����og~e�i�!6@:O{��*B��;�f�m��S7�Ir-rk8�.�1d>���>�kf׏�ĊU�����;�A.�;{C�d�Or� ��M�X@����� ���ga�tH+u|4��VURђ�u���5 �]`�`M��M�f� Q��:�/��튔k�1}W���~��X.����s��1�2zB.�8+̄��QH�;2U����;��F�Wd*;����~��j���bÿ�ܣ-	|F�u���@�qR����?g�ym^��2�-�J�&�و?T*e	��	��iV��~�p�������PftG���c�KllLLp����S�`���ڬ��1���
A�+����vV�Ԧg�iΙ�i3���� �!�$ٷ�q>��e3ܨ�R���;���S�y�@��Z6T�f�v�j�!v��Zl������ٳ�8԰x�[+��؃��F�P]��2%�ǬK%$��}#�DׯQ�[)\�K��ZQ��}w\��Ë�R��m�4�͑�z�s���Q���4�7Ә��j;ۉs��Ǝ5kŰ��*U���DlT�(�A)����TNe��EpC*:E:Ј��@� ��i��k��V�x����'v+w��jş(�n����h��F8�����!r��A�j�3��Έ��UL��&���WeC�CqA(�E��"C��@ǐM�T��,%��+��`N�C���d��;�h�jAk�1v9c;q�U1g�6��2��4�G:�=]P��-��9�lm���� ��F��'����\:+�f��0�ѐ ͌$��ٹ�J����~�4�颩|�ծ4J���PTc����s����p����F#PA�@�[spAs���d�_��L� Y��M���84Z� �uR��tTbb�CzR�_N�2VF49��~��N��'/�(�3��v(4���._��RƛK�����7M���oW�S�z�18V�F���y��{П(�<�<	qx��:B��VdɬFQV�NI2ԯ.�
gh����ǈG��#Q!�W���[4�F�utTh��m'�ѿ]MG�����Ue��ᾈ�*
����&&�^���pԦ�7����������4rw��ؚb�v�HV��!k�2-�{�sU(�2�V���f��XYr�䔍�Lj��d��������[���Iʱg�^C�Z�Px��������(zX�l]�Ͱſ����K`e~�R��1��ms�gK�}sP�G�'��
o��"�5�d�-����E#Tnk��Լd�x˳.������_B���i&QuѲ�Eo�a��S?"0���ܯ�hWƯ,)A�z�>��4��3cO�/&=����Yrgt؆�7En�W��UVe�׏I�Rx[OL��_z�bv�,�;�Ƶ���A�T)v�[n�y�HX�"�5��*��w)�I��o�^�fvs��[��1x�I�S$��{R��<�#Q%Yk���GRCe�0�=��",�gČo��p��P<6�eC�"*����ZA9�C��������mF�pk: �Vx��i5g�7�n�(oM�X�:;Rl�V�<'���֫Vb�b�~�-��x�2	�M�r�i�ڐ�o�5��)�bɇ-���Ěc��S��`8f����Wy�o�dz&��u6�:��_�������e37��O,�
m�CS A{&1��������R�V2����"j�"o���FO&���;�ؐ�x]3W�2/P%֤*�b�M�Z�ͦ��Z7��y�,/����.h����,�^�7�a>�Gr�K]�ū���8��YL�n|Ŧ����Z��`f�K��թ��_$�d-'��������L_H*��cƔޏm�~wT:�^����N�{g~����1M��(Kp,�Zb�*㾶�4� i��F���qg�x媥�U�9u���)d�*�4�гY�A������"�E�q���{m�l���H3J;ky��R�iҀ��뜥<�=F�bǍI;!i��&��	���N�#s�����o��W^ص8�o8o�8���"S���pG��}�]YC���#t�A�b���Ʌ�S���.���ae���ZBS�Y�z�;����0�X)ތ-��Άz���$T����)����fY��i�H������4)�xIb)QC�kx�y��,p�B��%��G����@={�KI�񪚂s��(�;X�G����߁t'����.�l�<�6�Ϸ���v���$*� ��Van>��M\�#���)(b��o(F2�α�+�3P�X����||�w����Ͽ�d�%��k�Fټ=��\�tj�$zMï�Y�]G�P�ga&K\�G�xC-9��Uq���=_�_3��:,h�K���uU�+K�z��C�<�J�*�O׺43W8��E��%��nl�)����h-�M�Q�.��3�w���Rz�^�����N�cR��Q�4�ϑ��p�4��L~8���i;V���c����5��*�&����$�I���Z9%ѽogs3cJ��L*��ŝ�G�/�JM��� {_e���fER�ށ�E��TGJ 
%]-�����:�0
�0Ӊ����P1�K{cYY�Z��N�*�o�V�4��Ci�P^A�HO8�͔��,J��>��}I�k�@�q�{��B�<����)�s�����%���                                                                                                                                                                                                                                                                                                                                                                                                                                                                                   (p         @p 4p                     Lp \p     Lp \p     kernel32.dll  GetProcAddress  LoadLibraryA                                                                                                                                                                                                                                                                                                                                                                                                                                          �                  0  �                 H   X�   �      <?xml version="1.0" encoding="UTF-8" standalone="yes"?>
<assembly xmlns="urn:schemas-microsoft-com:asm.v1" manifestVersion="1.0">
<assemblyIdentity
    version="1.0.0.0"
    processorArchitecture="X86"
    name="mulitray.exe.manifest"
    type="win32"
/>
<trustInfo xmlns="urn:schemas-microsoft-com:asm.v3">
    <security>
        <requestedPrivileges>
            <requestedExecutionLevel level="requireAdministrator" uiAccess="false"/>
        </requestedPrivileges>
    </security>
</trustInfo>
</assembly>                                                                                                                                                                                                                                                                                                                                                                                                                            