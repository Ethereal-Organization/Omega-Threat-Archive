MZ�       ��  �       @                                   �   Q�(]0�{]0�{]0�{&,�{_0�{�,�{Y0�{�/�{V0�{�/�{Y0�{]0�{�0�{�8�{V0�{�/�{C0�{Rich]0�{                PE  L ��F        �   �                �    @                      �                                   H� �                          ��                                                                                            �      d                 @  �            �      h              @  �         �  �       v              @  �.data    �  �  �  �              @  �.adata      �      n             @  �                                                                                                                                                                                                                                                                                                                                                                                                                                h�F �   ���פ��v�1�U0�k{ݡ���f_ϸU9��#ԗ�iɰx��8�'��ts���0F��,(/;�\Ȭs�R ��h�-I��iN�w��s��z��,O˲1z_����T�J:���Ym�1�3ֺoD�\�͎���!�!hX�޵\��Ґwp��,�e��s�p����'�!�ˇ��`�4>j���SU՝�z5\W����?	T<�Z�s����~�m�x}X��>�#)������eq�tE,|�� ��}Ѱ��3ֈ��U���MB��������`M����ܸ��|�|nS��$�a�1 fm*��(, �x�4Oby�	cz7Ӷ�U'l'&�,�����U�tf��h9<�f�n��.d�C����=�1�d��c�����Cվm�F'	*�D�o.�z4��,l(
 �[�?t��QR1��t��H���WT���w��b/F��`�C���H�sӀdĽc����
��|����S�C��M�!c`�-���96´?~�m��魱{9��xT��#���ܠ1"2��Rڨ6���so�#}�a���9�Q����=�ft�Y�]�)�������.8��mW�*�#c��		,)"�#%(wp۹"uC�NtNKS���HK�ako	p��ua\#BԎ�*t�'�����.�_0�W%6ھA(�1i'��[��Is1ba�A���P�>l�^���Tbê��^����	���g3��F)x��ni�s2��r<�GT�U��.�S��25�ױ�c�A&�Ï O�Õ�VT�aJ �o#�C�A���9��W�m�rl�w��xd�#�p ��F�E�T��D���_��j=O��h�RS�{�9�!�e����%Ȋ�:�8�y+�G��6�yIٍ!B�¶z+�èM���C�S7ozy��J��V,������<����1\�o��D���炂4<N���t�;fC���rH��_!��K�ZE�.1���/�`���l�c���0�Zb��p�20�EA�_��OEDI�2|�L���Y���?t;n'Ss�ն�cM��\�=���6�WB�1�g�m� �Y�z�����B��߁��(/k��T�	x3>�,xb�x/�m�n%bm����x1�,,:�*��;i����t� _��	I�HH�p����!�nTۈ�
`/�zs��pi����\����}��������2f�	m���y�Q�x'���[r���󡕅��3e=W6�����fi�#9'_F�ᰎ���~��Au��췧,{U\Ͱ-�TU/�Ϡ茅�蠗�����+tS�A9�[܋�9�!������aΆ��y�CI�!O�)4<��������1^���V�1I�sC��'A��P�]��ɯ�э�}�
����!�D(m&ٝ
����0?D�DKx�L-�q�s��J��� u3��h�����t�1�AX�e��@>G�P��Q����A{D����oH!���UC�7?Z�;]K%!�W%�K\p˿�`����2_s./��;�dr{����C��5�o>��Ix�"��� ���3A)m�.��oP���ů��(��t�ʲ�E�oJ��X�*���,ڙ�^�C������fB�aZ�v���W�HL'i���O�Xb�1a�'b����y� 2�=�yU	|zh�"�����	{Ͽr��>��f/VZ4TK'u����/�K�x�k�o3��tX�:���@\�v->�E�a���ję�7dp��RC��^�"��-���qG��ئ^��n��	���������t'l[���B���1��������Z��>�� 5�5�X�T�ҫtV�-j'_����>�?M�<0����>)VK4�/���{Kg5k��/l0'�`���¶�܀+���
�xP}*?H+-%�f7��A�'6/jUϛ/�r�$<�]�d_�Iv����W����!�_�{�(�뷫:���DS3Wo伈�y֪S37��T�A��'�dD���
gY�b)�ӢC+��R�˲����RM���e�Pz�c�����#"[��8���\�ZK��,�^,9w��b���q���D���	�]���TI��r�#f�����J)�1N�ض!�$�@�ē�r�Q���Q}�z�e{�s��������Ge����d� �M���Yg>�7C-O+��ѽ��KmPu1.�a|���Z L!�����l��83�.�E��C���􍗜�y��"m��,�?�iX�8x����aR�>*���U+�9��'��U=״��8�'�D
[E�j���e�^_�5�1$y%���Vگ��j�3�J�Ik�]T�P����\�� W7��;1B�dvp�۞|y^�k$�Bi��n�3��۔N4�K�2���ݔ�K2fOĽR�|��;LT��k��T�n���.[;0Hy�f�"���&��]j0�����������	��)���8~c�;u"3J�wT��p[�6�Q)�*L!�pg�X�.j��ny�
!�3o����켂���/[��!��w���ϸ2���z]B�T���r��k�ê]b8�0q�W�s�[s�ƈ���ޝ����D�R����2��
��o2kĤj�L�l@���$�ǌc%2e��k��7_�@{A����@K�������r�$c��d<��2��0�6�J:�e�O�t���e�	��\��4�~�yH��u�Zx#��@�m�-�lPҢN�?siAϝ.RѤ�К��̲�Tz� K@�4[��H��g�摇�~�����d| f.��֟����[4o�BqX�tׇ�7Hp����_ۃ�Gb-4��E'Us5���0iȳGL2ew2 �'��99	Ӗ�."�׋iv\���0R�nե�H�=���)���.�m�J?$��6	�N���^ �����e��l��j�������hk�-��.�:�$�	g�;�([Ƣ���Vh���j�X�L`�վ����}��z֘�B��z����3����A�tSQ��Z-�?�!����"n���Y�\K��w����1��C6�����8DŪ)�G$a��E���7s�N/y5��˥�\[�o3��V�=`�L~�`��'����m���a"j��yn߯O��td����a�@D���%�e`�ϧ���IK�R�_�u'�	�[�%%Bz���	d��U�0}�
��_"B���m����|n��e��z�����h���꾖��iQ#�yG��b���w�<�ub�M��~ѵ3AZ�
�u���]��6/:KY�r�N42ow��JnӘ�?��Q{m,u���H���!��㱯�:D��&y�˽yԉ؝G� ��`��e�H+�b&]����;�ԑ̧$���Ⱥ�@����3���y!��gH���.g�j�Ҝ�;_񈃒�G]r���[�u��(���x�|pA��2�������T� ��w9���Ql��|uν�NK���OF�#內K�DuZ���Lp]�u�r�e����C�^�cI����-�F;��;bȨ,���,��st�1��N�J`[gf]E)5����Y���w�׈8�0���z����%�7�yC@��W�ׂWV���6���xN��qn�h餣P���<���Đ��~z�T:��G-����2�3���ȴ��YA+��f��K�r��.b�!�<������^@����(�?n2L�8aU�M��ѥ%T9��ǷI�f�C�Y-_8��5����	�>���j����hif��h�Vu�=)b����Y������K���h]iＱ�gI�jY!=���ts��y�SG�t>��6X��ZGY��<jp���D�l5%��"�����;Q���7�����C�Sڣ���$*��E��k�_�iE�Vp�Pp/3ը7*� +0j�Xx/���D�2��5
6�)*��BI��*:��(��艼9\�c8���%�_I9�%s�8�v�{���/옜��P>̈́��}}(�^��zV�88�q"{,+���ݪ=)��ø��`�zg�M���Ti	�h����K��莂;�$ک�
�+���sgj��'1<�dr�d��kL+��N7�j����L���}��
�r�j�0�L��ϓ� �Q3��<������G_@��P��&/"1-�d󴴡�{ΐB��e�U�}ޯ|�ݧ�^e���_��ߵ�.r8�|C,�1�s�=�rVlQ=a��p䫋�o�/�M���f���������Jq���'N�6�M�=�6��J�#_����P��/+�~���YTNlj�o���ڑ�}���Y�}�.#/���7���35���k���Y[���z�=�-ײlIs�h߷���S�E�]`�%q��R�&����`X��?okV�S! �a �d��nU����K�(n��7��ɛ��,��s�?-�K�,������B�Dߠ�SC�ߎ;����0'�;y�4Ќ���|ս�	�cX�B��R�����[�q5�={�?QK��+~��-�V���F�J��frV���S�JBF�_��\�����P	l����:�夜��2,(٠t+({f�M���&��ɑq����cH�:���D��Tޮ�v���~@FYƞ�d�P��B�"��Z���C��|�G�L1E���C�1�F�<	B 3��wAf����6&��\�ŏD��%�{xCێIL-1�XY��΃��;��hv��l��a37`���2�q�@��u��|�HdAě�W�$ c�]�/�9�p\��n����ģ��1̆�"=�ܶ��ݾ��a�}C��rj1�ݕp2с�9���'Uj���2�^!R�iz>9
�Rs�����я�I<W�er�[�භ���gT���^<!h)=��>)����k�H�$�1cP�5��m���O�a�Qk��wB�T�X��n������`γ��Xj%��>Q`8�M�w�0d�Q�H�vS�TY��sqM&Q/�䝑�ǅȊ]�VQ~�#�i���|������=^G��1�wٮ�f�?^�|�5^.F� ��8-�1�J�_�=�Z�_W�GT�|svyT�6�?(3��gdŰ�!����ISl��/�Ҽ�]E�*\��v�$]?�h��BI6O��$�#�u�СC��K*ⲥ�"G�ôu�AB�!�_�Bৄ�D�Ҡ��G�n�q��A�%�(|m|j�9���=$-��/�8K)d�D���iX-V��\���ȡ�
i��D:�Ah�.!��T�M��p~>���bW5S�3�2Z9{6.�ul��C�V�@Q<;0�d&�wˬ��$��R^ޖ������O@,�E�v�;+X��򜤇Sa2XE֓�si���&ŵJ���*r WE��)���\ 1�۔O�D�+�\��V.�\ra r���+�=�S����y�#�I�Yp?��T��n�G�n]�CЅ�V��0�-�E��k�w� �|fΑ�4���GF�(Z��ez��P��. N����Qz���`:k�ݶ��<n߷�^�WAKx��/�;�y����9V�F>u�Rz"u�G
�`�IfI�+	���x�\���u��?@"�ʴ�p8@�]0 �S���vMtA�1���)Zѿ� F�l+��-֜�-��xkE��<�~Г���_.Gԝ�Y)���?�Ȍo�զY~Yy����/LO���� E�
�����1椏�u��!�r���y$9;���Q����<�ϋ���h~<Ȕ G�@a>?����ѹ~�4�T}�4 E�Z��#B�~]/X&g~Ѽσ�L�"kq�kq��B�W7�����8�#Em>Yl[
1�P-��B@�	+�HrC��]���O�=����wZ ��x!
��L@P3�I��7~j9zk󎴖�2�?�2*-̞��X��b)ˌ�w<�ܽ�Q5��o��[$�QD`����s@�`[��'\�a���w )���z�V��{��9�Ǵ�*ֱ�ս��'<��/�������9��)��R9�8M�����Y; �
�t?Xt�,
ͭJ߰�fzݲT�I�ei���-�;y���&Sf�����S��c[�](u�XTk��
�~	W��Ȟ�YG�ٷ2��̗�0�y~�$�p7CF-�̇��sT�9=��l���`?�o��?��Q��e���ۖ����K{2e�����K̘s�׈e���nĤ����p�v��*�'Y���jtClq�6�_���qy�� �����~;����鈓:ٌ���y���r�2n,�C���)�)��f���+��̩eZ��G���s��;�����A�G}n�,���#��9��&��5-F��v�~|� YP�L���U8�w_�t:�A�R/��+�S'$z T;�U�{S��'�E�?�ڪ�/��c�Q2��z�~��s5��2���=s*A��.'u�n������#����[��� �����u�h�w7߆ ��� �c<c3.���u�wcK�q�؇(�[�)�MI�ж7��q��V�q�z&�x�6�IT %T��c �B��&_X��e��<�ꋽŬ���f"4W�_���F�5F�p؉H������'�*�	�4H�A����_�_��k�pvq���2o�;���]�vO��_x�2g#j�{}`&x�i��'Є�����*й(`õ��A�5��K�r ���D���]��@H��Evz�Fh�v�G�o9@��6�w��t�,�aV���j=n�FyV��Bjq*a^f�>u�k����4�r�hd0l��w�lo�T��8L.�Q�떛�;��O���D����r n��@JPs�1�Q︶�)�{�Q��t��:`�C)iS��޺=N�	ƍ��^˳�O
�M�����S��٭XUDXC>Y��0჈8�T��@�D�hi����y���B,8"�)8ȱ�����^��ַ����͋~����3�:a����5��^ggM�p���+��48n}?8���M��Ui��(7�+���И�����~}{�6Ϭ>�￣�λ�R�o��{�i��&ˮ�#�\��S�X�[���0�W�����g�gҏ�Z�z�:b���wt�FUtJ�+��J��i}��%(��@��N��g7%R��"��r[P��|���$���/�%lJ��GH�u>�Ug�h�A<�u�A�`kOG���2��!*�����k/&��a�W�6��o�!�o�jB{(�E�� ���o|߫�}0#"�իk3P^�J��e�i>QR_����������nAI
�f�v,J<pS
Y�����u�b��	=�5���+Q[DlM�SO����%���pR�!�o����5N��p�H��z"c�i����Oe�%c=wMV+K%�d���<�����x����Z�T3:���yyuL���( �m�Ko�֬��u���I�e ��%)Z2�����6_;D�3ִ#��ct��dء����k�d����� ��lvk5��y`���B�T�b�r���U���7�4�y[��w2��O��#���+��f��N�Erq5�]�����������ߗ�K��[q���K?�mݬ�d�^��"'�!��R5T�[��*r��c�%ܤ��|�	�"����h��\���#��xx͑ ��/	ÿ��G�Hu���Y��C�_�7�Q�R%5w\��hգg#10���sg�5l���&���^�^�� �3X/�#��
�MDo�p�_\�Z�i�+/?{Tl��~�јe�q{UUW�iJ��K5��� ��;���&9�jd�[�S�e|A���Z��m
�H�`M'z;�mtk\Ql=TK��yěW��F�����L�UƬ�Ǌ�^���$�*��H��,cS:��'UE�[�`�Y�I�3s_�`�ih�*��v��Է1�Ɖ� î[��d�E��|愮��w�zH$�S�����%lX��}�L�^ECYtCX8���b�[c0��$�v:aL��|_W����4�
���]��I���R}8ٳ��^�Vb�����3��,3ݽ�dg08L�E��>�%<�W���ډ�;W�=5�mk�ܐ�d��T�����E	f�+a�8CϧZ�8��x"� �%D'%����� �7�m>�n,ܙɱ#�=�h��f�U�v)yнe	X]����Y�.^���ܽ������y�}��\������E�+C\��)��r�>�\C�����D�c���	)�eI�Al;^��$(���K���gs<���0��S7[N�N���M^x�ܝ5~��/͈�x,�S�m��]J��ƶ��f�m������ݽ]$����es�˙7Y�TZR��c����;��7�	�(Z�($T$��ZL�#ʼ�:������k>�j!�����+�?v�ӊq�E�}�[|�,V�������s�0Υ�������}�E^ �"B��,�j}���&�ôl:z��/���hf��m
���M �bW�p��ߞ!���؛�O����&y-�*Eb����Q�g�9��s�a�b�Z2����w��V���:l�|�������p���ߧ��f�{����e����rD���B�ct�&%"��\?n���q����"�&:��ql�r�n�د�

�dgr)���Q�z>[);�깳� �ZG�xe��Q�N}r/h;龟dSnև�5�p�Ap6K
|mΡ�v��4f䉼,��޷�}Y��A�y�e��;U��d`�HC#S��ɑ�3�|,(���^�٠uY�K�=���@r?"�fT�0Z���.4R�-�h�+(�� #�#�����#ê���{k�,��l\�W���-D|x���#5S�m��1�7ɓ��Λְ$U��G�?.��RA �X� ���'|g�p�1���MG�> 1�1��d�0@�`� ;��*IӁGZ�JCm�9�Τ���KVp,����*�_��iѴ�^�A��H���&`�
��(e���[Y-dE(G�`�V���c��r������@$M�ʐ��[�K�O&^�L{U�}l=]�e1����O�F�רQb�Y�Em��oqYz�Z,4+׳e�v�.��hx>�Θ|�P�|.�`�U�l!7GW|��\�}-���f��7��c6L����8���Տ�iQ0W��M�Ll/
�41ה�^{���,�r��K����h�d��< ^x��� �cl΄�a댆b�@ڭ�A�
-"u;��!KN��/+3�[�3���[���z� ��Sh���#��S����Ft~�&I���,������Hʚ�u!�p2|����������#R�����t�mcn9�������f��w�<N�G�}���w�d��@��5�pO�d.i�>@#V��h~�r�H؋a�V�N�Cr��N���$jj��4�nq�ϰh�O*>���X
Fc�����Ug�i�IJ/������)��i����9&��Uz(9q�bu�B�d��܂*`�ISa���V�j����������SOYG��E�����'g�J��$ZP�f$N��VI��9E�@���u�2��̙�F�α�g�L����ԏ&�R��g 0�	��
4��ֹ�f=�'�iY3���߰!�p,2�m6�%�����;`�"��ʐs���x�{�k_:���b;� ��z=��L�8^ S�dų���.�縂�Ρ(�Ģ�_J��gȌ̡bI�&u�~p�4ũ��Ҙ���=<�Ҟ�?�+-��o?U����q�HI(�swM#L��y�����V+Y�0��iP�������Qs�Rx���v�5n��#��/�CW��Ks�?ɴ�ǉA>�&�,p�2\N�vmj7��=iɑ�l�KP�>
�
�hH{����:'��*۷o���$(�br�M�����'�	��������q6�"bh�榷�q��չ�Gi���d�|�y�[������K�7����~+��D+����,9�q�[�ԙH�
#�vC�2�Fj��o���@��l���t<*z�j�=�5�F�V�U؂�֔��=^ �p�>�{�Z5Y��0��v,D?ٙ���c;��R��w8٥��$b����i���F��$�B;"5���Ꭸ��6�/��0�"a�� �%�ꚵ�5����h���wS����<q�`P;D4�����dS;���ܥ	�3k��$�w��U;����^�Q��kMLؑdA�w��l|5�r�_aU�Z������w#�b�J@��g��Թ�9���:g˻����r,��*4(d�R�.�`��2����M�ii�s�c��ٚ�enX��[��ey�jT���ή ^�(�[�^�}�JO?o�Pl5xWz���� �,����f?$u��/\��oP��QgH��Y�3�.���v eh~�g��V���xTc���
�[�� ��n�qZߣL��0��r	�qw0��X�/��/Z9��T��?��W\�G��� a����WjIx:���}���#���ŋ�����EO-� ����8>��O,��j�G��l_�"(��9�q��ԥX�g��-W�=��0��68o�1�����I��
���{K���B�@8y<�z�U����;d����	���g��8�l��:�B+�V�@C�*���(��?�ХUKc��&�7�	<�x׳�^�b7iStH�A�5�{�[\�M���rX k�	˽����"�`c�i�:��ֈ�>���z�! S,������lw�}���%�vx���q��R�@TRd�]���q�ͥq�SL�I䲓��M���<�D��������=����F�cLG�Ù����ټ���5(R	v��n�Y�Hy\&�+���sI*��j�.��SI�)����V�wi��e�U�(�ƥ+���1~�����F�r�樓cq&�a�}	�櫨��@,<@$�b�2C׃C�C�n���5�OQ��̽�~�3Gy�Q��j��y5�w��񡗥s!�)�祀d�e��-���;��Oz4����y��~7'Dm�n؜^Ři?񯠍PƤr$p#�[m��F�'�v&��|�V�Ҩ�������-����	�|7B�3�x���w�8盘��+_=d����̌�ݣO����Wl�o�֤�+Gz�s_�
6n͜�?jV�Ȓ���<л��2iPU"�
�v�v�{.pG�XvF$���,
`y�%soi��./���]�ʽ��6�(+Ƨu}Ԛ�]9z�f�e<<w�Q���f���0Q+-�`
Ө�^	�#j�$�P��K�F��f�'4˒)�|L�sݓ�l{���P�Ag����q*�t��`-�X��u��9�`�!��t3F�9\�;/�qwL�p1��]��<��;-�Y;�V�� ���k��@O�G�[�T�Fi�+��8Aռr��P O>�>Ֆ\��p3ea?��@��Ǣ�vPm����o�s#�U�)�[��7��(7?�5����[���T�Ğ��Kr�;�n�P�O�^Rc]���X������@yR��]*Ԗ��Ƣbo�.GK��hD���'���f�#Yo9��?p��sE��E�#�>s1}X��ā�A�%q�J>�t�l���,"Ҕ�����>��p�x2!�xD�u� q^>��-v0��VI��yЀE��*Y,�Y���>g�W�5oȺ���YM��
�ΰ$�X�l#�)��PRk{��[��D�@�;��g�+����Ey2^7���
���u�[�!��BD�R�ϣk�k��m1z ��Ѵ2�	'��B�ƥ����jC0�5�<�Ա��cs�Ɍ�ћ�G��a=AG���ؙϧ�@��Cr5�y�ғg�R;^I5E68�� ���j8��E�P<��O_LvP��:� �O|�*�32��6E���Y���	b~hSD(cl�tk�ُ��]4�oT�h����F'��\��o�@F(�����c�ķ��>�������7�x�)|,�>H՚�i�:a ���!��U�����Rc9��*��y�z��c}7��X���!a���� ���򑣹�����ܝ-tSP`�~-Ni@2��9?tT���! ����D���L�@R�����O\��A�9�J����s]�����$_%�5Mw��(,\�~֢M�z��)2����FA��jx~y�j�Mչ
 u"��9�+G�(S)J�'26��x~X~�MZ�T��1`��b@¡~!T��E`�ʻ���W$IE2e���=�36,�~Q��r���r|��}��}�~��uGvB�1���SB�<��,�X��A��#�oa� �Z���V`rsz�q��G�:�����u8�Q�!���E���NCͽa�dT���>�l{�,�q�,���G6c�vc5��G�������$ӑpr�frh��P�bVH�{����;ٟ,�q���6�;ݳ٥=a�s$�с��?�O�w��c�1�[_�@.t�jT.�3�5��)w�	R����7���S����.�Z�7]}b�^��#m������a�`%E6Y��g7ܿ�K5?c>9 ���
�U�G-пUJI���i~��qx����е�^~�b~!�ʃE�|c�x?N�W<�r!_�U�⓫`�ᅃA�}���3^Fg.�,�;�Kih����n���M(�@+��-�c��tQ��0�C��1���w/3�*a�<�w�r�L�*��}V c��(�`��ز5(��y��#E� (�̈́��[���
֤�4L���3�&�]ɨ?@`{i�"_�蛺GdF�l�~&ln� �z��B�[��wd>���b	ȗ���Nk9��9��
����c����1,A�;zi:��p�J��e
0���q�kN�a����URR�E.�Sì�'(�/I�*�,�
�]���	�wa��i��/y?9�?��4 �-K�Z)�j+�C�ci�4���:UrK��ۧm$�F�����P�=�&z�<��mJ�d�̦����"���|v�ld�M?�F��a�n�'��#b�H
&X��w?�u%&Ǝ�I�^���)a�T����woU6:?1H�����p?�4'��V���4��eH���d��+�Vy��Ⱦ�v-a�Ώ_jh�>P�%�u�=���1Z/C�h'���;�wl�f�W0��{e�MX�Vy���
_8V�����Kw�#��1��VY���*�$�B���ƦnIJSl��&�&�EOK��҃q���*sd���հV�8��i�6��9��hvN�s�u�>���3~�\�1�c�@����l��S��ˎT��$�����]a/�6[ȁ ��M�t�vJ��Vb�1�k��j�Ҧ�z�NLq�f*��v^-�6�u�0W����zV�s� ����n�JR�ĉC��-��nD9θT�Ȟ-i��3���=/�
��5��gF���=��?1����z�N'�R2YkЩE?�nww�cw��Օ'��E��7-����*�م_J�d&6��l<������,#^�N�ٺt�AQb '4Cχ�R��[D=�'01����wh1�f�X�/����:��~�Z�����i�z�0�/-+=B���c1����]�����:2u���,��-��>�"ە0�Aߨ4�S_�1L'�a9���� �ڴbY�,�&41`�y���.�A�jY��Vě��N	.����Z��&���GH��5KU}$��p����jRI������ױ䰫&��~-�G���I�E ����
�|�H�Ҫ�y�Іڝ{�XH�:����b ��
�QPA�m�+�Π�꫚����L���Ko����������2H�&��A���!�z��8���7�י��>VY:�^����U����:���E�M�X.��Dyu!OuT� �-K�IaN�+�@_^^���1���O_%:�����-���GdL��lf7<�����<�O���Q]�j}�|fd�q ��Z�-~W�\C�����£�_W��@ ��K�0�!{Ƿ��u�n��������0F{yÖ�߅�Q��J�:���:�����ȋ P㟭��z����B(�k��
�V�ұ%�_q�0�m��L�����c�l�܅����)gJʸԾ���\\Kq
m4.�Ca�xY(����A�6����9p�-X1p��w	l��n�{�q����E;T2u]�a*i�������w�N�E֚�$\,��)$�ta�Z�_����1�
�,�*?F+5Ca�cU?ڶ%m�e���oN0KN�$v|��u��Dkl= `>o�84�����Wod@a�ö�+~SaQ��r�`���*Ū����:G�= Յ)=C�%�OK�-/3sx�8�1N�-��6K}�x����=�G���U>��8�r��a��o��kL8XFH@���ZO��f�"ė����c�ԍW1Dt�����[$`�dm=6�QSL�{fzG�Ph���������P]4a�@]�-��'UL`���ls�^U��7h�)+�yyg�c��j,������d����J���t�ɀE�k�Z�J]�.	�Nau���H)�=M��3R;Q�,T�����O�DV���t���yi�l'){�r���&P��BU�OU���~��.�0(�[���B-�%!�N��_�Fw�͓����R����1���3��%^o�+���2�8l�Q��I�)���o_J�;SC�f�c��@*�}�B�'��ٌpW��F��O����$�Ms@�����fY�`w^�\����������t�I���������8X�k[��Wلw�=� ��	<����k�"˹Eڐ�XI(���]��4�~V")�Y���@Ap�E*ε��1� ��>R0lY(��7GcB."�?���T�h�\qu�]x�O9�u�G�T�=��j$|��}��3ඐ_6V���E�/S��BbgZ�h�i翅q�eI��$��凐)laV�nW���if��-o=c<�5��Z�j���+��L}���t��>��1�����OG\r_fɕ~T��SΌ�Gja�eSi@�Q�1{��a����!� ��m�a÷	ZP�Ӈ���XFsO�m)�d��:B:��`�G��ٙS�K;�5L�^�i�h��`!�`�)��*��8�L��Dي��JB�@�zh,�]��}��ڽ[���>����r7�D��g�)��9l���qi���}N�e���
�	�RH�J�9Y(R�j
�K��\W��p99 �H�![�^�:�lcr���!I�$���^�;3j#e�2���#�6��OH�[ �Hh��,&2����?��0z��4ga���;g
3B��q�AAH��aD�.��c���L**�\��x����xVd���v�=�	�ܢ�9����A����n.��3G��rh&��?בy�N8��+رMD<p�϶�`W%ATR�|��߹s������"�����Z��}���<	�rj��b1���N�t�h��pIb��D�GFҞMy"�pk�Իmޅ�ܠR�G��C����->��N��K����q54��k?f�>1�Y���@��h�7��(=�ǪB}��/��')�H���T�D��K/F��������(�NU*>�%y��@ �:>�@�V�誛�9����R�WOk��B'��Z�}o6���4He�)Ti!2ė�A��j.�����3X�4���I�T�G�60�S���~6�L���] [5�-7t���H�XO�Uh�t{Gc�￹q�bH�6�ϼ	�H�I�#���wR��d=	�UOS'<�{�K���z����T�r_i�.�E��g�����帼0�Խ��L��'�t��g�&��j@�e)x���Jf��bb1�R�)����fp�1"�P��3�3���O�'����׬p <)�_�8���T���b�U�Fd�p�峠����Yv��ޏ���QE�{�ge�ACz�p�DR=�	aaͣ�T�Ƒ�煬E_g��h����i�U�н�Z�Ā���_����a������*>o�L�a68p
Y��Fua(�L�Y�!$n�^=�1���Z�W��C���Z�8�V�`x��`29_'f�q�q�i}$���ѿ4�I&y/ n�H�u���!p鬮g��|��c.4�����u�>O�b�w�<ym�����Ht%p��9ypq��wY<Ď���՚��6��@0Gq6���	m���%��x*�1%�(���(S�y*Fg�a9}Z�ܭ�'k1<|X~�H]�hh��O�U�uj��7�C�/Y��!,R�B�ȰK����%*!W�<C����ߞ	<J�78�A;ӆ�-���;�4:��Z���[��w���Ņ�����=�K�����\V$�m>ؗ@K�&!c�;Qkf&��=6獵�
9���D�r������(E�Ж8�`X-�?���c�C�C!�cZ[�F�r�܍b�0�ۂ�5�کj�Cc<�ϟ+s�b��D�'8��X�O�2��7 x)�QL|�(�TOo�g�
j�ؠ�����P�h�z,Q�Y��j��u�v��>O�h:�y��R�Ľr4�+�iH8�ɉ.�s�U������$�����b�Lz���Z��.t:���?8~0��lX���$�,�-��n�~��Qf��� ��R���t&� ���I��XP��λ����1�*&x�P�]RE�H�B覕��/�.��d���Ʒ�(�E�����"aO�j%	Uy8#I;��3�L�{�2F��s��9l\%~KE�P��@+�cq���c�H"]�+`��]����zX����3���V�(��Rȫ`���F��k���0&�~.H��5%c%���t�!���s�����l��dHw�����K˖��̌X�$3�X\}�AxS�o���7�f�`��q[�Y1ǁJf�"K��Eh�ө>����g_AX��'�v��¤5���~)�:��
�\����hy�tufz��~�L/��b���'0C͚�=+��+�G��k�Bۏ�*%Y��bri��ԛVPڠ<���E��ۢ�Q��x��{^����-����;,�Z;-�)!�]~��uN[a) ��V*��FD���uzp5�%[�Gc�i�

Ǚ #+����!$'wUߍ��1�z{ۣ��j,]���q����ճ-�Q��.zj�TW�R�mB����:��vAmVk��񫮾��GXC΀r���ϐ{KIW���O�Ɗy����p� �vw��рn�Ҽ1�x��T�i)i
�~y�4����z�4���v?J��
A���/AD+A���tQ�:�aM��[�Þr�6S�K����q>׿�W��ؙ5�JL���D�Ɇ���?$��	:ݞ�<;��}��F@�W��t�׻4z���?��C�<�n�4�
SL̕%��{:#��V�D7�I���m�w�`�c,�⒖���	���{}|l��G��05�#Mu����fg������Lᬻ���T��6hf-���UÞ *2�$ü�F"	m���ԎC�����k���� ���1��QO&�*I��4U+����K�����^�	d	� ��bv�V��7Qu�l\7����$�3�؊����Feŀ਻;����,T(�����hSH$��NfP|����81�×�U�IZx<PL�.6K*W`Z�=vS���4]I"WX@�]6
@o���w2f����c���X���b66�,���j��s9ַc�)jGv['j,Ň|m����8��=��]�؇F�Ҍ/u�c�yAMNipL^�P�<��ۨ�YĚ
��:5>�^th1��V��F𸺡 6�c=dy�%��r�]!�E��/������ г��)B�-��|�6/����^�<�$��p�u�π�l���k<F �̨5��d�F�kW��<�B�Y������oc%�ʙ���b3�a��W�i�Q��qB�Hs$Ԩ�(c��cݨoŔ�8<a`֪�T��^�d��#��jό�>�X�(���&��J�W"I_�s�(9\����D����ݽ���F�@|H�e�Y}��I̘��%��2^�P2�i,�Dt���ˎ=�5���֌��~ȗN�Ł>ȋ����ũ��)wZ���6��ל�De�(��t_AaG�fY�H !&�t)>���`˼����Sץ���ѷ����L�ۦ�����)�@v�R9����H�Y��W8:6��\�R��w��x����˞e),��� ���\��}0miQ&��<ĶK�Ϲ�3�5��#����X���KB��)T#��~���9��s�ʋn�G({����Th���A�-dX����B�7:��W#�� t?��I�����å�#�7P�R�<����T�-�XW��2��G�E�:���7��J��>xܼ�Z̛I0Sq03��׷������)�[D�,��?'镑`*�O���g�PY�M��]� �ߝ����+s����<�`(O�-�3�/��:�!\&�1矞��	�1;�b���BDI��)j�����*�A��|uM����Ћ�d���]gz�iX�W�9����B^�5'���\��N����
R��X������uG��f�zZg���4��G�~�I1�Ny�T8p^W��s����o]o�Zãg��E�t�j_��x���}H ����s�%���N����z%#0t���}�y���v������h4wS�I�S�&z%���3��I�t�[���if O�����{H�炗"ٙZݾC�5הjt�9�s,#5��rMb��'z��ZDyY�b�nD+�~�I�ek�S�9�=���w�@&@��!v7��h��`C��Q���k�DA�`�-Ui�u�7u6c���dU�If��8ԗ��ߗ�xh�'�a�*K%���jXx=�^�.
��	�`L�4���9ȣ�v�9Y�͌���TQz|wMiBԗ��<�CFɰO�ݿγ�[�Ei����Y5�<S��h����/]��M$jf�æ\ �N�r:^����V�NK�4��,�����k��n׿�9�W��U�,�4&k�He ��8���``i�t�#AŽ�&��A�R��� R^Q7�W|h�:1�w-�������T�o���,��2��زN<�S��֎��E�m��5:�0�_M/�Pw2�ch�P�<Y4W1�h�s��q#E�'[q�����_94�+-�f����&ugR..�r�=��}PT\���:��kl���dH�V�~-�%Qn[�!���6 �T��Vt�EQ�3��E�I�	^3�O��"Ӑ00ܿ	�'W�=��Q9�6e�R��a�+�PJ�Or�4�o��.>P�n��u���&� =�/&ժ{�� ��,n�*����4�޺���u�}P���x��7?���<y�64ⱺ�x�:�'�U�(g�
2�O*`�P'y��ne�7����ŋ�`_|	C���g��9�Fk����v�k��m`uZj&ὖC(�mG�d��j�s���2�\��S��hJ�M_ĭ�ҋx,	[�G��}�:��y�r�;
X��*�I��l���"�i�9�J
��eSF�9 j��|X�+������6~�38Oπ�g-	q��YȪ�$�{���J���h�LP����=���2z�	���=�e�ґ-Q���3'*��"d���>QMc���]�$�Vs+]��l�{c��|�愢��]�6Y@�cϥ��z2��H�>�؆�*�Z�����{�Zg�H�e,~咃&��j.L����k��bw���n�x�"r=dP��F|;G�;W8I�j�gT~w�۰��p2L��ͅ?nf�"*�WD��Y_��R���p�&XVh�n�����
�y�t�5�VD���J���=s�j��tD��z�g���$�<�i�^�Y!TZ���K���{�*	�PL�}/f䆞I��T&�R��ii��d��Z�%� 7{c8p_�*N��d4r��Q�&��"�޺�B'��V�6x�WԢN@3O��i��^fOC��*��ߕ	,s�E�r�"B�%!����U�0�1N_��m�ۀ��^F{���߳~(��*���9��jT��Ƅ}a�#��Q��Q��
�;�	��8߄۝+�E���Yk,��7)�AH����E�	=��a�U=|
�T�{���hu� �ۄ�	�T��L� ���<� #�;�R[C�a���[��tv�0'',��k�]̰�Z�@��
yF��X���Ӻ�*�q�X�4����)�GpMKE�I�)ƩgxB=�&�q����P�9%W.
7 �h4����"b�?9;S~����y@qR���I�J4����ȹ�!����-�O�����
���~9j�zj2&l��]x�y��,��$�oKg�l�n�\�U{ $� ���Ռ�Z����C�@�༄*�d(6�j!lf���P�r׷�]�K���)0��w~�t#�ʖ@�H�$?[��Uk�):e�n�d�@�E�]'������ 4*��ϑY&���ͱ*a�����Ф*x�$�K����������1�Df����{�E���O	]�K-�G]3;q��V o7 y�%�-H�P�4�%,0x��{gw�:���������ܚ��TXubK�Y�;��c����(۸|茚�@�c�cqR�n�"TS,������>G�g�n@]}�#M�=���JLkjP�n$�.UM�0��)� !�I�&l�"�%�`�l�N�����g���T$���ݕ^�J��z��<]8���v(�(��MVS-�7�:�U9��4M��4��`��, �b������޸�9W��t���rʞ�$�� �Ycq����<^t1���bO�P(h3��J����3<����w��҆Tu��}&!�����{T�׾خ�LY�'cj6n�G84������M%�$I�m�[�F<�vw�:%� 1���t�-\H���ނ�cpj��*�}q�?�Z�~�#�t����Y���|�E2��I�y�P;�m&�4�UԤ�X�OU�э���*�Ai���	����L3ǵ�ӥvb��sV�Vq��&ӕE��7��j*��V��w�p��o{��d�U�2��>�� o��u0qؗ�#�����7O�p�k�
�qK�O��Ќ>�?3�������sA��&�ō�����[�5|F��� [���q���	���YT�%u����^��p��1�,�%�!�w������:�9��̳� �K<ç`�p��y�]߬|�G^�����Sg�(X�*x�S��꾊޲A|�N��M>%~`E������Z��J�C��{��5����K�|�S�!8<%��-;�%��F�vPU7�"�p�N����̹��M|��_ˡx�Zȅ�Տ�3��2�g���/���˲�+C�����/�W��L��u3үY��q��*Ԩ�R'�<�5�[�S�o(9�*s)�X\�V��籐e�hw iKw]X�O�S�d�{��j޲���fZ�S��P�fQk����Y�a�`�٪Ò���#���u��7����DJ � ş>��@G���gE�t���%��!�g��;��n�*qiJ�u��j��L�%���y�����'�م�$��ݩ�4^�l�[H�0]���PXH�(���>f�#�'�J��/t�U��ք��;Ar)��<_c|���m^	�H%�{Jg�6��Ք��P����ކϪ<�|a���I�Z�קhe\���n���@�Ƹ�-]V�;�wH��S-H%���L�Ԅ��Ⴚft���w2PK�䖾������4^�dE�Ta\�M*����`!�{�8/�[J����!�||]�����Q�UQN)��F:�ZiG������t�
�����0[^>�w&)��t+�>���]r�i�-{��r�b�c#M�q�=1�M�g�@^7�lS��OY�4A�?Ǫ]x����U@-�?Ͷ��Ԁ�d<�r�z��MZ]����rT��G��=H���4U�ѫ�c��:��Fυ����A#�Y�կ�]#���㇆�fl(���t2�1NPM��T874]�M��,�;>��n����"����C����m�S��HfL&zL ߜ�t�}���a�ln�T�k���ָBY��b F����N�]�f�L��	�_����Ǉ-]!?ls}�&�U�~��%��/����#��4�y0����ֆ���%�Tc��D���\�`?>�*�#G���X�Y����-3��moK�>A�k����:�_)�W���ޓX�˧&���M�ȼ�l��o�8ua�`pX,郊/�z��� ��6J��?Mzs|e���<<�;��R�����<�(݋7ߞQ�4�w�-��k/���I��]����1�0�UT<4�cv����%�����j�TĮ�Yg���)���sm߱G�дK�����UC��r� �/,�'��m��[��jxZ����қ	P7�).+rS��x��m��/���s��o�:��'����ҥ�?�!�iR�ZY���%��f�3jZ)���9��mc����� ��X����r ��-���"fNPxv 8�9Mf������v�ah� M��[YUw�~(�A��2h��i��t�\X8�58�?�ꃽ\U��> ��h�٩B""�*j'l+�dw�g�> =�n[5�DBmS�N���]+8�#�j�p��28�4��9�O����y;��'�I�8<�?�>�C)K&ӯdZҋrxX���'�/ir��u��rs�h����:���f�(�j��O���KsjD��X2�9׵�������E*s��mi:��ۂ5�6��&���2=��{A0����<� <�|+�I�Nȫ��fHD
�\�MW:G:|j~�ɢ���[ؠ�(?�Ե��>Ľo������mP����ԫ-�ΒX(�1y1�b�I�)u������v���������]�醮R�N�R$/)����q�2��e�Y���e�i<�e��t��Z��P��TnϻC��6��L ����'्q����o0K�4,S������Ը��8q�{�l�`���>�ʯ�+#�����z�_�ӝ�����}h\{¸*9>����WLn�qM��$=�6��<DPЕ���ӢGE6Z�ѷ���I��Bg�4��X�����>���C��a����@ }l�򋫉���d�YG3�-�K`uF��ש�ɵ���ub����B\�R6m�������_�������d��@[�O��-�I���d"�^<�����-�ג^�ș���J��`����T�Rr�0���XrnT��ᷱ`����|N��w���>���8�
B�P��X��gٴ�k^���Q��vN�����F/�	(�`G�z��⌍�U��{�� J{��7�[ �V�AHC7�h��ܳof��ѱ+�ĘV�6n_*(|��"��:>i�O�pG0��}��v�������Ϸh1��i�&-�L%^�O�C�x�ߛ)M�K�[P��7�é��6G%�%o���a��´;�Nmy�\�F!l:�\=�n�Mk)S2�v���>�n����1��q{a��[1h����|�;�^�Y!8hu��岲�B�N�u�x֍b�Kw���"I!c\}Q�x੄@ [�\]�~�O0������і��u���֎�XK�۰;Ǔ�h4n�#�3�o+AdѪ�Il[��M�A�B���	h�!��Fi�[�� �{�*"�������q�3��}��]�u�g�P��^2|�}M09�
�s<u�lo�V��,�]� �8��հ:�,����Q�1?I��#x�G/���;��@ɦB[P����"�[�J.;��VLF3��=v*&�
�������Ȝ�J�/������R�q@��?a���j��0�����@��\�y��f,e����"U<a�5�T.$��^\Z�\����k1��;�_�lJ��O�D.zNZ��Y��0A�>%��f3t�;0���Q���9�)�n%`�����*Dj*��K^UKCs��y��c���S�>�7�>��	'A�7纍���X���$�NA�D���e^��/�T�^�P*��σ��g{^���`�����X��#�k2I��>A��k�N��ђ� 
20(�Y���,��yn��Q�9�@Mx��[����2�ﮓk� �w�������Q��$�v`��i��xs�6E��q>��TB91'-]��^o��۬������J10*m��w� &cc@@I��p���Hm��^ae��<0s���}_��dӳ�w��2L�n:5�7f�uG��5.�VEӣi�VM��q5p���C
����0%�K��X!�8�}�ߍ2�Q�c�"9LVM��n��7n�miX.j�f�������)\���ap����02��uߖ�`ɴygsE�@kӣ ��	�b����4�=	��p����&�Ϥ�H�VRb`}l��ۣ�=�}xBo@�X�j����D^>�y���|�oq/M�F�$%�����۾4=�k��(?������
a>q�Q�sE��h���*y��Y-Ka"�g�^��[���~=r��!���K�pXŸ�]_�	1܆�l�b�5�M��G7:�(�>U�wH��
&�:\�����f��.)�4{{\�孠�U
q��,�����!If9�B]���&[�Y��pP{�Au>�����R�(�5�
���~WF��;SqC�JZ����%��b�I%���ZB`"�H�vA��]-���zV��������m)5������R�d|ǡ>�t�F�"�.?PP���q�P;����%��1a'��Ð����G] </���<��G����2�4�ʒ�B(�R(N9z1����|�nh)�v�����Ψ�GǪ��8�?�*��'Ηhog�*���!����?gکƋ`�@��iz�U�����y,5��Z��r[���d[��Ē6��(^�wx햅c����$���Jٜ�Y���e���	�G�8,�:D�b�3�hb�Q������iLC�Ţ�Ҡ�����@�"7�)�~�Baʃ��/���|^��$�����>�^<$�SF��|�t�XS�@�F���[A���H[�2��-M8kJ,��~��r�+�4�)Ca�\��
�Q#>)��	��%'��b�d� ��8����un�,ү�qQ��qd�0VN8��k���b�pn��D�m�u��j��q���� ܔ5)��j����O�����Ҁ����s�V���J|�y���C�qa bh��\BB�p�?|���ʽ: �p ;3��" H�N�Z�ދ;�9��w���<	P�7��%#DT)\k�ag�]u�XN]l��f�`|�������_a{�)BxZ�7(��(xHzTZ�%���/oȉZraO��'':��'z���,n���������z?]��F�)e�cҁ^U���H˼���z��UNd^e\�E<���<����CX;9yy|K>�v�:7�Sb�v��q��t%��h 2�&5�4#y��-�i&m���T��T�5���4�֞W�+�w@� �f�[��25rp�Z�s�.+�cj�-��|��Z�DY�>Q
��.��3U�:��/-r��+K�ѥs�+8�\NAT�t��b�����҇�9E�K�3C���� �7�ӡ&_�1�K��̕��7��0� FpA�l2��v����QGs���~�^^�4Ś�[Vnzv����d������^��q�,V� ���d3)��i�_�?q�}N\��P2�/?���w.]tĔbi��[�|������X��L8�o�4'���d�����%�7���5c_U�g�H�����6^�l|��zڽRb������K�J��ei�vr�lz��ن����j�fθC��fT��NO�4�Y�`~��'%=��9D�n��ȂѰ��R+�\��["g�tx�~UF(.u�%���S�%6���~%rk2�S?�0+�l����C�e����	"��Q�PVw�w��Ŋ���x���:xq�zQϊ��v�U]#��u��(�M��^�޵��=bX1�E^�$nAT�+�͟�M�n�����y��f�2#hJ�s����0ac �Pe��r�?<���"��&�zy�?��$�e������*�� �����B��W��6��t�r��`�g F���R���zu����[�V�6��6�\�>oL1D%M�ݻO�x����}Rcf���� 3���P�?��c3N��A�gQ�;F��d֜ ��B%���D���RC­F�WWRR#r�N8$Rԧ�*���vf��w`�}{��}�b��������>�u�������F�]�07�`�ha�2�Y�j@�>�j��
\���Y���#�^�*��-��t��`�V�����p~_��dh�ʜ)������2Bk-�#�Q��lj�v�Y KH���ف�¸���pF�A�m�a��L���#3G4s�:e�:sRV(t�"!g�*¡ߒc����<�x�^  c��52���",MM�/���(h�-Ph�ca9*���ΡK�J��X�CU1y���B36�y]�]E�����I%r�!Z񖜆VLZR��(G~2��bDh�G��|�; ��]\�����\�,ᩙ"��'�������{t���g�����B��a� l�^�:]%o[��d�Eގ�z	��Z̴-Qt������4�1�IJ.�B1Ja���)"+f�KV$��Hx���GE�����H�1��Jv��|��0�u�#��Ă�ϴfB�zI���Y�c7}��4�y�˻�By0@��r���bYn~h2�o����� �VE�`ib�%�j�1-A��>_S�����)�b,���m%�jd<�)�	�t,�F��I�ZWv�1�����"�r��2��>�	#��>���Q�0��I���&���Rv�m���l��o��+r��>�{dּf,Z�x��f�$N���O��F(���d7�3��!��4����ۑM�g�]џ G���ܫQ/ЌP�y�"ڤ[��������/G7���{C�eDk0����`"O@o�Z~��6�*Y7c(�/����)�� ��`�4�7?��&0Y蟊�C����ͳ˼�f����Ͷ�����
"�4d�}wGo6�%��a�����.<����WeK�IB�ͼEz��@a�B7�4U�@.#�>�]�*t��g�/�<���e}r�i�1���p����r(V�W ^[����S}T�	������:V��5]ҥ�G82,dN˘s�[q�^^�$S?tͼ}�5��_�I��gǌZxe�8�f[=�C~� `�χ�0�wu�0]�iob��CRD�#u@n��7��ϫ=v�Nڦ2H���Y�J�'vH�C��+͂7u�W0>��eG��E���Q������w�̋���0�>s�����Lt�es�p��;�5�*44�0�+�e����?��q��Q[؂"����?q!y������01��!�<�ȴm����9ū�WŹ�j��s(0\8PWvL�`��u�Mr|.d�庹�:�1�
��Q��/�C�ѡ��4�p�/��2P\����6�
�������;#�Ŵ�\]�>]!�S����pSm+I�)��z˅L��,4@�����5׺ކ�,E!���mJz�5u�J.��:t*,�K62��un&.MD#67%6�������!�����+�aNJ��=���S���T{M��@Xv������,��K�E/j�����f���}��*���S�����q?� cƾh1�D���q����^��i�6��_��f���9/T����؛t0~�ݮ�`A���(dd��Q#�� �dO��p|&Dr�V\�i�SD�ڨw7v�^����Z-7��	���r��x�6�K^I�5�!���_s���?�	$��7������0��s����I[�`*�����HN2JnU̖�
��v��<g!�M�{�z���$�,?D���J�Ã�tFCd?������iL�A�>>^IEIXu�����_
+�z���I
�s[�x�0�_"#,�w��h^�ϯs�8��uօS�D�>�2q����%M����]�����zѼ���j�+�?^xv�֩��8�؊�4r�����H �~���c=�O�����WYxK�"%�v4{�?՜=a���Y�hԃ\��E9�1��N��!���Z����t�`B�z�<���e�ž��;�ئg_Gۍ2Wo�D�l֎�\2AF������O���Vq�j*�@�m�NQy��q�=w��f��H�*=1G��dc�o�u#����6�
�m�^r�po/�ĞDi�(������U�5�	��C��bct�?m��-�F�;�]�[~�
cq	��V�����I����:m�<M`ض�Ҧʺb{m*�N��XH�����g��;�iA��E[�:�UV����ٲ������I7�Qs�"Qű�eh�~^�ULM	�;�n��a���*�s\�*?�c��^aD����������`�t�2�$�
^ޟP��_9q���͈��;O�$�u-���6�# e��� C�G�����`����߹P˭�y/��0�ˇ�!.W��CL�/1A�U��)fܡ��,��5唟�e�郅����Wպ�3c���s�f�2��#J/`�!���l9���x2���&��gi�0�Pr�3bcӲ��T�����`��*��B��zw=�(���wD�`O��d<9���S�2�̋�^x�4|M-��L�߄/����-Ǝ�����+s��6���K�(z�� D4��� OX�S)V���V���oC������P��&r�!*��2?�����O]6�`��$�m��9'��$�-G���}p&�,尯p�LZ�!�#��V�;Kbی��4B2�?��Z38���9`�ۼ�D�Q�dgv�ݚ#�JJ���4}t���k��@�mBe�1��aIEpxd���L� )Ƹ`fo��W���i���nG)�c�&qQ�OZ�Ɓ}U�l����EŌYh|1}O�D����r4�y��1�G?B�9~K!���_��Y�gH��,a�mڠ6�GqK�0XM0a��Û��U:F���=��#g��A�TV���ń5!?��#f'���=IyW��?C��h�~��&-f�f�h^�A$��D���RY�A8hX��ۍ�JLŪX}/��J���S�LǾ��_��)N�?�iS�'I��T�Y��u��@T�F-+q�I���.F���Q��;�i\��l(�>?�--KK�9�����w^:o�1Z1q��h��Sa��<+�2�KJ����sR�@�M�L��۱���r�=��pp�!� s��^�E���>y�,g�^�@;�/{{��˯�|�7�Akw�ԍk�;��Mی���еL^Zj��� �xp��S_Nz$p+� `�����|Z�1��v���Rʶr���H�.E���W�J��a}�N�j�y�nF9����0��3��M�Ŋ�Z���)�l|�C\�e� SC�s�:4�Uy*�Z��7~�?�`�6[�A�Xi���@A#Г!� �H�5�1��NF��V:	��q�զ��kӲ>�;���w�a�RC�;)ơ�B*��a䪯�]�j�/�i��aK��ո�>P���@����iK+4(d����w��[���q��!�QQ9�wJe�}��ۄ����,��3��W��I�u6�!'�؛��h�<`Bf�Lx���\�Bk����܄���uP���9�t�t�\Y⨒����í��|�B�u�y^�3�9��W[&��/�>��^��B�'��d�LdVݨ��Ye��	��	��,�`�����l0�ʡ�pi�
Qn�ꩿ=���S���@�??��<�Q��D
ڌ�.�����s�1�֝�#1yp���YG>s ����é��)��H5H��3�x�݅�dI����Ť�{ܗ뀻�!e�ie��ߑB^V�ӧ'��h+��ٳ�ߵ\��5��t��k��\�*FQ0 ����؛,�Vq5h�O7hxc�N�1��Q�[��m�+��(��T�eU�`s��<�X��}��\TbC���:����}ܒ��=k��g4U?%]���^�pky��@��s��-ݚ�5�ɦd�'�CXM8M괥'�����+w��1�r~Yi���i_%[�e�އ�X�;T�2�'�����@k�
�_~����e�Y�f���7[�����6f�w���M�W(@jR����0�*�s2E,��T@�X� ���_�J3�.��nEMF�}(�L�<*�K��:X�mE��z�Za��ܮb��r�=��T���i',`���h�O�����G3M׺��E�N�q���@K���W�^x�����+�p����^�8i�hpL��;��}]�Jb.�2&7�_"Vg\u1�-�zi��4f?H��R�V����bdE�&� 1��4[Ji�&��(�o�Q����yؾ{��Ϭ*�l�kBA��k&�;���N��Q�u��T��H���>wj��җ�7�6!x[���� ۫ļ�����J��c�M��)�m�Q�P��e�5��K��㦋����`fg�q�K��U�u����i��Ғ�@s��[|�fVX�x��4�x�C���	�PA���Ur؅3o��o���\+\��EPh�TӛJL�V�c44�xȐ1�T��6���v�w3�.K�V:�7�b���n1����a�x9���@�+��d��q@�S\�8�Sx��朵-Z�#D�rF[bvz�ļM�
�L��z�>��Ԇ!�}�ĝ��Uv]c������6�K�A*-��3�Z�B���>tߑ�&b�a(������M.I��Iϛ(���7\�돾�bq*�jp�F8�b�W��F���&#[d��ڴI�iʥCJ�����Ax~Ϫ���o�pum�ԩ�g*� ��o�������W}f��;���
�o�D��&v����Y��h���䧵L���-I��wb������/�;��[�͊�@���Z>�/�پ<Cg�Qy�{��7NE��:r`4�N�Y�L���ߔ�`�5���Y�>ݓ�LlR��_��* 8����j�5�1��湣2��T���� )F�g˼S�~Z����i�Kҙ��1�/��g���Y�i����[�Ep�1<���mt�
�:ȡa���ƀ��2A˹���c��w	E�]��6ͅ���J6�T��'�I��i���M�p M������Y�l�B��F� !8V�0�����dQ�`��6ƦSKʸ�fq<u��%�eA��B���aP
�9;���Ǣy�����~P!���+40�?gg��+F�k+����x� +��� P�/��:���0�L�V
&5�u�TD)1�g��%8{S����o x��`7857��wDI슭8� �p�8z�I2��fX��tO�-�{���:F^���Q�l$�׺L3�6��֊�c���jq�������	&�ņ#����/^�}�Y�?�
�x��c��6�K%��u��H�E6(�k��5%HX�P��ƾ�Z�j�F������f�����ĉխ1����x�ҙb���^�������D
���_`��B���Y����鳢���ο�eeH���J;�������Ip��a�r]����y'»�UH�y��(��E0	3\�6WU���n�n ����c�����e��OJU��i�3��Ǻ|	iy��E�Zq��#���KMB��.�5EΧ�{�xX��UJ��K�(��|��^g\�joM~���z��Q$ucZ�u��~��p��7�OKR<8�F�˔�w�&u�P���d"1r��"4���6��"_�U����u�@Hڣ�q�/n}��˭d�j�h��Gq0����)��߶���~0��<�o^�'WC�U���fz�2��4� �X�8ߌ�W�d��I�7�w�6Go(�3��1֝`��a�>s!b��#����CK��l&�KP��ð�@k������Oo����(��,���'��gݐ�ۊR���>6��	k�Yx[_�@8y�Z*k:R�++��;x�0�G^�
Q��!�J�� [ܡ4qyM�0ٸ�T�)Io{�O�����PQF�V��}V��L=C�B���[#�$	E)cZ���؎�I:w�]{9��\n*g��,���V��sH��	�&o�|w6[1ѧg%�_�'�*�Q�_��Y���)%ͽ+�8~��s�O�<"km�$��/�zU.���)&�nr��Gi��v��!b��0�F���z=l�1�\��͔0�B.L	�ރ9Y!Ǖ�ҍp�5J�eK���dܡ��@`4�_���[��13�jE<��Ѡؔ��~Ue�l';��u�`�!`ԭb#�Q7�*d�r��S�WoاZku�N���}���c�'�)�Dqjm�>�,P���.,�i~��໹&6��}A�=��_�u�1�+���"Uˏ1�)�׷k��~��ռ�%�^�^i\`;DS���9��խU����çz*������.�d@�K�`���"
�t4M��F���VF3:y�>)��v�KZ\Ӯ��4 �R����T����p�6�r,8HGۢL�{ùV����&��~��\m5o!g��|_oj�ӊq�4�ŝ&:Iw�1�Y��k%2L���t���IV�-,���/w�.�˽��Fѥl����Ÿ�:��7Z�2/j�2��AW�YX�G%Κx�_)~�ߊTO��jQ-�.��eJ'f�F�
|<��ΰJ�`����sB�)��W9u}�	�p�Z卬���fSpM� �/�������"�+�����J�66j7�ȖqH� /m���'0���Ӧ4�घ�u=��?^��Cl�r-{P��VB̠�c��)3q�J�;�x4���,(�Վ ��Q��j��CӒ�#3�$pВL����n�R��giN �4_��l�c�a q���X�@���H�u�%��{��l4߲E_M�j'A�JVB@�Ͼ��a��b�
ğ#��I�z����I&5��+@_
��	%ׁ�1����)G�=Y�'�vK�Y��A�͗RX���8�V�p�{��V���3���M��)4�,�fZ*y�{�$}B�\k}+ O��1c�s7�]�+����N돞go����ۗ8!TŔ���n*�9܉���qa��>d�ʊ���pC9C��v����]�!d�1�!U���H��K�
 �?]�f�v1�~�������>e�ۡ$b�x�kH� j��#X_m��{���{h$z��ZFd9[��`�g'D:)�)������5$��Q��b�:epR���x���������(�yzC���}o���(#���_��U
�R�WyT���,;�ɔ�-1ߙ��_��#q�`���b�NH�5�Q�'I�(����fDc��:����� tzȌ��V�{�{h�FM��^�}Ө�e3ŝ�M7�0q4*�`Ŋ=m�&�']}����V��+�wžS'�^����=��K���UTv�x���:G'C�N�r�����,��;��8�?)����� ѩ�E���~k�g�:U�D�c�f��d��'A�����z/=����13S`�ȑ�~bݹTp�v�ud��P�κf쿻]���8�m-�S^�(>ɮ�]V��4������r3�#
�wJ@;&�0���ij
��9س〕΅���Dʬ�_uB8�a�j����>�ݷ�H�4p�j��A��ֆ�Xv��|��t���@��VRہ�����u���î�x����!M���堿���=C���4�Ȼ2�U{��>9�*]�w���.Q��b����psu氤���g�sl��%���NxE~qo:�lҖ�Q���1��pK
��� �Gg@�m�-������bUZ��	bz|�'zo ���X��4�*��8�tY���=��@�n�VF�h�n�a�̖�RQ.�#�CV�9�C�F�h*o��
�܋��┚ڳ\�J�3��΅���>��qk	�]��o��0,	Ĉ���~�m4a�oK�jYB(�b"9"2qT�R^�!����Hࡢ�=�6���=�p��7���t��m����)��L8���"}!a2��������j��;��=:�`1s��tT���J����>[V�/��}�м�..Z�Ƚnt�a'��R��dT���c)�M�3sqi�_�;�Tr#���߱l���	�پl�� � �Pॻ�S0�t���>*����n�I��3�)T���8�fЗ�-��={���7�=�̋�q�]�cQq��&���~`���6������%�-���I�.g�T6E0���:B
9��cC��՝� ;Ŕ2H�h�+ �����L��A�Keg��ч��P��:�N~fY�5��eizX�T�7R�,N����?H=� �=���Q�"�N���>T@!����Z�g]Gv������>T�F��.�T�������#Y����d<Fe���;~*
`����Nȕ���Y���c����v��bW��m��.
v�ɿ�f��l�%�)�x�D���:����*Ծ�u�����y���_~*��\� ½���V���ɟ1��s�X�Ʀ�%�.�Ğ�e-3+/hd��!���P�Q3Y=�i>�h�ᢠ#'�[G�9ن�`������^��6{����F�)�;�gl��>��%�U����!ir�\��'��TBi3�81��=Er�x��^�&�,�p`*��o\���N�Z`bW����6'��-P���M*������mJ�g�4&�rf� X4�'ĞO�5�*α AM�Y������/Y`h6O�d_|���GɥL]iV�4�)���Z5b@�x��։;8�p��F9�n�����٨Q@O�����we���w�@��y3�{���.�d1l�v4�Ś\���-tyM��p����`K�sN�8������ɝ�� �>B�' � ��V#0�j�\�;�y��cċꓓ��J�n������uF	{�GUL�i�#&Q�˟~��S�n�{�Q����p�.R�z05�hc#��I�1�)F��k�E^�aEv�@���m�ўG_��K�I\j8M��L�[��Eb3��7ud����P��z�e��xv���A�޸'�_w}���A-R!֒&����:�Յ'�����:�Z�hc�>�9;�<6����	c��1���1��|8��sx�u�x�e���v4j�?�_ӄ�u���`I}�c�@��;�N+�tU��cb[�yC(g�d����B�]�U������v[���)>"7P�a��Fc����W�c���q�?5"̝y��Tb��G�l�(�^�S��&���x��U�	�Ccx~!�n�*a�|iKdh��>�i�='c��rD-�� �K4Y��쐄��e݌g�A��q*rAa����P����Ԣ�@ycƷ��0Kaj�*�d��!�/������?#�rJ�'?CT�	!5����S�f����ev��d�`j� C:���Fxf��D�4G�$�n���Em�v��8���lR9�Z���˩�{$ln�!�[����o�0G�0vv��=�u�>$A�ŸAh��Ce�Nj�wV6'`�]����e������I�E��<)j�
�H���x�i���y������?S����������_\�<��Y�Ȝ�o�u�L�DU\�-œ^�w����?�}��̋���U}n|{�#�����282��k�7.�#W"�^z4��b�A��aɬ�ҳC��nA/����=H[mz��nӼxB�>9쯢�y��Q����?FyFI���8���n3�-Rp~iq�d�-�#{H@E9LZ��%�[�R��z���,�i�yP;J$U�A��'Ѩo=�i���4�����/����&���$��Fe��M��U�^N2U��Ul�c� .�����z�535#7Y5�<Ab��x7�j�D��o{ڭ�����������}�����:T���G��C��pV��~����LyA��.��`W,n���^�bj�95RY��#��CȰ��`ct��8��v��
9C��N����kY�#ж/@A�O_$_[��G�uo��b+_�aJN��F�����C�к�C�;&3d=z���1���`�+���u�I���˰H�q8	Z�z��M�PZRcsm:C�._�6)´�"��_x!��ȈF���[*�E�Hm�+���D�2��Z����0�dz��V��,�#0�]��ؑO��ٱ���D�/�Y���
�WS0�t&Y���j�6�A�[Y�g}��� ��b�U�АdK�@�,����M_vO�@/&L�|cSW��rT��ܙ�ݜ�0B��V�][�d��9*a�!(H��0�$�⽁s���*0��FH�	�]̡�;L�K���g�*�g�`//*Ab�fܛ�VPS7���tL"���V3���'Ԇ������5�h�DPxώ���&�/U4i2�����"�_�t��;���Չ˾zBYu/|z���x|��%6[Q;��9���2,�+��1 O�Gn�|1�|)"��ډ_�|q�4�')�"�@O-R��;�������R�������(�U�!d�������D��6�2��w�~yc���k���GBf���ر���aQ�|�+u�3���E'7�ٽ]�f�0��P��Gj��I�*j�����|��έ�~�?�v�2���]�U�`���Ng������{�5���=�'tB�DX������B>�!�T��FS���C��=x3�8�8��V�Ɩ1"O��^�h�3�=��#{���M��LD��5mN4�dQC��5�����(���^�8�2,Y�K�xm�$~�Z3XJ�r3��}n3��6
���k5�I���.�`�   ��]EU��   �]�����݁� � �}Mu�t$(���]Nu1�ESPS���  �E5P�                                ����#PPEN[��t������#t53�Vj V�uN��^�� u$3ҋEA��tRR�u5�ЋE5��th �  j �u5�U=[�aujX� 3����@� �J��,�   �1��m�3�i�%��f��Z�¿
  h    _S[�:�
   Z�h�&g��f��[��f3�N�   �ρ�&@A����T�A h�o�z�y[�:Rf��[�   	/<Ł�Kh�:�
��Gh�:f�߁������������U)���I2���*o�����T6���I[����/�!p}��/�O��KnP�DS���-1�f��'��q�'�q��J�;-͍��3� ���E
�-��A^��I-�~G�-5�:w}�G1n+e��j��j�u>���s�4���R�Q�V+��D�jm8�Ҝ�{� 	7,uQ��:(��"�ʕ��)PaB�rϝ��N�VT#��=�����R��r�QFZ����,�֊�:1��"F%���цn�]*����51 ���4�6J�d��+�N�1�����o�#���� ͦ����S\l�S���"#��"#��̇ϴ cx�Yܥ����+#���>��"�G?4̯�"_�3Jl������b���`��H	4���"@❴�yz��dY ����j�/]t����ޕ��:]~.�j×�%�/���v�05r��&�j|����Ep�/��|6��)�Ԙ�#�/�O��,S��P�$�R�
�#뽍�&�FaA���
�B��k��Q���/�j�T
7�`Z��..���B��m���OJr/
�j�/��c2��Q0�\v�ȍ]K��m�F���Mg��$�-�,A艁�?|6�a(z�I->cWW�,Z�Pآ���Ϸ�o`/+�h����{��-�,q�Q=��$y���'�v¾�^�a�e�D`�!X�sw���nH�m@Z�n�M��[%��o=简�"�-���@xL;�"��nT�����W�,�"����3���uO��8�s� 4�,�-s�!#Ƴ��,�<{��,�'�k��C%���IN`�IN�Iw��RA�E{⟣�*aEV��۾�����J�"���*�ⶤ���{�*@W��y�����N=-�*���{�*@W61��*��*���d��O���h�"k��*�H������[� x3����#�*�ۛb�?�#�A�Y�F�#*�iT��˛*�p���%��q��:�*x8a��G��*��C������z�q���*�q���*v`+��.�*e��*�HW����o�.�*v����*v���C6�*�~!gv�c�C�*�H[ux`j��X�I�����*xυ�Z��v��z������F�ƚ�L2�� `�b��:�*���hx��v`n��x`j��Y�~�����Qxݗb����o��*v�_�j��*���%���O��J���a%�H�p�*���*��*��*��ox�fx�c��o�I�\yY3f��������,�<I���3f���������*���,�<)�<O�I�\�P���Q�{X+3�3f�������[���s��z	����*�Q�{X+3�3f�������:����*�Q�{X+3�3f�������G���d�#wBm�Vq]>5�����:��*��<O�I�\�P���Q�{X+3�u�ԛ*�,*��H��I���k�#wB-�Vq����@T�lx.5�wO:�Zq�yX6UB��~iox.5�wO:�Tq���v�o��"b%��*x�7~�����*�%����}�c���C3�*�~ё&�Z���k��*�D�����7�*�~��Ϛ*��*�����u�?��G��*x�;;H*� %������a��Ou:֊;q;
C�����rb�,�Q��ԑԓ����?ӥ����[�)S�.��~1�"Zp�0t<qy�����F��mø)S��7#%��*��*��*��*��*��*��*w��E��*!�*��*�Z%��*��*��*Q6a%��*��*��*��*���k~t���� '1�HX�+���5�\j��^1>�Nܤ��Zޫ��2�k�%����%��
m��/���m|�C�Dv�I�A�i���˕ׁ��Jyٖ�J�TЏ�~���Q��{4�k��No�z�$gO��1��y&��|���>�έ�).)z��M�-po\�N�B��ic�S"��cV�Cm�I�+�.\�r�G����D�WO`���,%�Eж�C�`�?�U�T��5:]��?�E!Pt�ʺD����f�W
���V��R5U��8�p��u>lhb��Nކx��ZN�t�x��D���`�i�zV�'���4�-޵o���B���9�6/���V>2�`�%�a^Ʉ���Đ�����(��O%�m��UF�M���b6*[/���֢ �۫��MOa-*+5�G�3#��~�,�n	�zN��L�JY:�ɻ��_�JD>��-w%��a/�`��f��L�1�z1[5�l�`oT����u�>�p吋k�1��h
�
�˛*�]�*x�VP�c�!1�t��A�*�/`��e��I�����I�n����ڭ�٭�;���Ο��|�b��U7�ܷD��(��^�C	��~am�f�[Q$�����4�<-��nD�E�<qo�#?���G��"�h��۵�DL�g��\W���}�m�9��Q�m=�R�)늞,�=g�\���P9o�J���꣎��+���4:���~ޛ]�������t��l*,����ܚ                                                                                         � &� 9�         kernel32.dll   GetProcAddress   GetModuleHandleA   LoadLibraryA             � ��             �� K�             � S�             � [�             � c�             )� k�             1� s�             >� {�                     user32.dll msvcrt.dll ole32.dll oleaut32.dll mpr.dll oleaut32.dll kernel32.dll ��     ��     ��     	  �    ��     ��     ��       SendMessageA   __dllonexit   CoInitialize   WNetAddConnection2A   VariantChangeTypeEx   RaiseException     �8�pg��
�!]p���$�sܗ����=��C$ "C+�(Q�0�I�Z(� � G�x@b�7�02PQ&%�{P"�D
W(��N�&$��X8$@ Strin5gX�P��3r-$"	(D,�d H\�TO bject�%�!E�� ��� �r�9��� G�#���Ȕ �r�9���"�#㑀�|�xrt9pl h#d� `�\�XrT9�P L#H�D�� ��r�9@<��# �������p��F�T�S�ļ�
����#` �D$,�t9 �\0��8u[�,PL<4�G0#@�(�$�  rSV� L4D�>u :h���j��ۋ ȅ�u 3�^�ʡHC9�(��ҋ�������& gB��du���� ;Y�cT@�X�� ��'>��� I��P�V� ��bX 0B���֟� �
�QI ��>�0Ð?WU ?��$E�b`��jn] ���;�C� �S�u  �m��'FH����P�� N;�u]G�ߞ�|@~��� +�B�jZ *]_�L��Q<t ������2� ;�rl��Jw� �]n��w^$uμ f�)�9�{;�@�De��=
 �r�w�M 0��A�)s� �&�*���$+u��ϖ д�wj�� x��釨P���VY�*�@9���� �N�}(��� T���;�� `�sj, h�2VI� ���;��=t#�ӸP�H�d�J������OW��d�U��$}� 9HPaj�W�Z US�u^LyG �%Ǟ�;
 wW��i'l� �L����` ���f_Tdh�>	��y*��AO�
Q$�s� �wFI�; �5���tjC��V�v�k�u�`sM�
 �,��&P߁��Yuz��`�5�|p
�:P �" +��L���)������ �����;���$ ���-�	Ȇ�H�+S�:F}5�?<�^�~ L��v ݷ���<ip� 	X+� WS!Z]�J� 2�6b�� �B����t �,��H�S �!�4�� �V?�� +A��8�$s�x �W���@��B<����+ Et0�>`7 ��T?��� ���]�3X;,J��CU�_��w@PX� ݡd>(5�
��Y� ����#/!��ƺD��3< $\�]#觳7Y�	��\,t>0�?)��Ab`�`Uu;��Ȯ ������%�B�+ʧ��0V�/M�, v�3�7$���I�@u���'�S��m��� �Nb��GC4� �f���K��H�k`�u�:I ��m�z!�Q� 8��(�@FO�	ER��� Jj�ŀ�#�>��� ��FC�L6 ���; �s[�ρt+ ӊ���Q� "OS�|`\  ��t������K�G��+8���<�;	 �IzU�%�쀜�hn` Kd�s2=�"�0(aɀ�A�e~
�+�azw=���B��h��Y�C ��-�=c&�/� ��3 ɰ���@=A� @�p�'� �yb|�(a�&�ZY䁌�h uE�*�"
 ��o!Ȋ� .]čSL� �C��R��t�/�'hp���	`'� D����� �<!�(=� �r��O��<��'t�2�^��`u�Y ����j 
E8��P[�S;|�'	%��H�\���8�m�:�y ���"�� �R���)�$ J�(�,�� ��®�	 �HA���a �J0��r�P��2�u �"�) �kĨʃ� ����|�&����ф� �(|q	B��2 ���&�R �Ѓ�>� ���H ��.`6n |��Y+��5��*H J
p�� ��6�3Bᤀt� *�"��T� d+��3��� �� �G�;�F(�r+ �;p�b" �W�,�U%d�AX3��(rg Z�����$� u����W2�F �#�� �,���R	�E�Mfq>A?uܝ�� 7+�J���s d���} �k�S��f G'x�%� ��F�_� ,	���{0�+@��&���5s����
� ���?5x`�*��YZsH��0�߉����;	� ɕ��f�u7��i5���lL� M&�����?\t [�	�:��C��Z��,<|�9��
��35�-.@���,G~; J�9I����+������ O�)e�F �&Yx�k$g9����,��� �����	;R�ZH�&��g �)�Gf u�$t�?�L�3���z�$� ��Y#m}{o �5���>4�%�]� u��� =����'s 3`6���{`[�u�B �Y'�^̍�R���Jk1�` X�H�I�t��L=����\ v$T���u �^,�&�|i ����\���t�w��b( /l~{� $�21�� �B(?tw� �Mc��g� $ؓAN" ���邠� ;��H�)
� I}�L�~��E$�b50=X�٥�
���"2} �L��>&��ċ� �<�֒ �M�`�u�4=񭮀l?N%]� �JUƶ�� ��L�
>�� ��^r�� Uh!�&1��/ �wF� ����pz�� ����H��RtyB���;��� P�)u* �%�K�|� _�	��G� =�Џ;
$M� �.�a� R��U��� ���G"���b;@D�J )XT�� *rL�C+ �U��2H����NA (�G!��IV�d�]ɨ$�Q �<l�,�E� ���� �r@��H�x"ް ���>,���C�	1�xyL�sh��D���� :ИTt.$E�[ ��PZg �����̩? �
�H+�; F�J���, W�'�A�;="Hu��qbV�%�,�ԑ ~4��}p�\܋�0�t<s���B�7 �Q)���xh�-�]@�$� ����,2�� �3%�I=�� �"�]�K ���Ƅ�� ������U� ��o
��a�	� � @����������u8��	)��S<�}��Lp� �C)y�� b3���(S�0��]�uH�.��SJ���:>S��5)<���� �r�gY.>� #|S�¦h� ���(R 5=BP f,��%�P��?�u��4�{ݍ� R�ߑ�M$x ´/��; ��	}X�� ڤ����,� �I��$ђ V@�H��| :z4��)> '.�V!  ��}�Xz"3 �$(t	w�sk!J�Z�� �Xt������" �9%ޜ�(��� ��]��6 �l2�3� H򟅝b� O�4}8��0%�ˑ �S��?� �L}��@%��8��
�� , �IÄ*���ܑ�u�� ��t2�|P���Y>u��$N��G�:��R�e,5П8��)��0�U���p��H�*O���y�KM ����?' ������������� ����� ���p�,�� X�PRQD.�X��*Z@�#1�2� P����?�ҋ ���:ȑ�������$9� tK/)x *�����1�t��� |҂�� �3�A�LC	��x��P (�~����< v��;":u�{���	� ��_%�� >C� @V�!u�n�X���(��= �|[�	_L�? 3(Q�/v^�pwxO 4h��d�P&��� F��wTƐ)� p�[��=� �h���|K���=�c� ฯ��\� Asg�E �k�<f��}�x@ ��U��i� �p�� �<�ʳ�]�x ��߀��XZ�l�<��G -I$�߸(g ,�Y!=3�&�	$���RL�Hǈ� ��ڱF��zr(8��ы��3$ז o@�*v�� ����I�d 3�
hAHb� ��(��" �U' $Q���� �&9�uEN��Y� �sZ�8���7N�`_�s^ �t6 �:
3u0T �H�J��% A��1j\�8z����ޥa��1����̀��jf�� &4A	�MC�_�@i + ��BT�;�X�I� R0�����1 �)N�^ R���	�0�C����u}�G-@��G�L$ ���O~(�<)ٸ!���  ҊDx�+ Ku�	� Ԍ���|�� yș�Pd�sv�ƿ��p� F�� t�� �-�i
+ �f$x�a$X� 0��Y(�O JL�? � 4��0�$�� ,9��(�~� �6�U4u��͌ �|Y1 ��2��F j�; �~�x�)��� ���Qɼ�X ;T2taߒ�r�� ��v@ >wЙ�
 �� Z�]��@P���*B8��t� (��u$�Zq<�d �������ҒVى��) ���9ھ�Sw�ր-H�� ���  ���ʇ��$��C@.)�Fu p� D��I7�� v�'�|��� s��QI�D?�B��� 6R��Z&W�J��PL��@�#�X_�p��^� LY��.@� ��"���%� ��3۲� ߰� Pu�� %	+� �_$��w�zq b����v  ��s�6�Pj�h�+��.D�?�k���M��Uh��-d�0�� � En��`�P .�9�i�&(��� �g�^+� cK`T�f��q��������?������*gpSOFT WARE\ Borland Deqphi�;RT8L FPUMask V�l%ue"� ���+�Wcװp�1�5�A F���P�@� �G���	X �s���i� �6^=�%v܀n��.�E��+	u�K�w�*4� �g����O$�z ��dX��t|0 �GUlQ<� �b�2�>����@��׫�K� �@���e��=HY ���,��� Q[�b��Y��9� ����s� �\��|X{�48 �Inu;��L@�p(9����Hx[ eð� -W�K�'h� ��� Q��f�
�Yd ��X`c)~ �\G��r� ��<�S=��`|���9PR��@����3 Xxj
�[��,� a��RQS���P�%� �d�n� ~i�A }-��t�U 
[YHZ�� �p,��t$�IP��X1n ��!�d� �R�r��	�X����}�@ �v���=I��0:�3k߆, ��̒`� P�bTj! =�I��L�� ��QbP���s�����dbz��SOK,���A@�9�*�
$�u� ����Ĭ.P?|�h�zU7�ڑn�
8Y�Z�(�R D�� ��v�X��4 �8�;����dE?�0�ޅ�P���tn ���jK��X����Q���"� ^��9������t7�0���v )s;w���( P�k�e�9�x��a0�{��+���;(�V��>:���=?��to HS1���&�d��>Q(��h��/� ӛ ��k|$D[8��Pm��o��_�G��Q1 �`W#eC��6hʈ'�ph@A��g��{ R�+,!nbtE&��`u 
�if���	 M,:%��p�Y�q������xC@�Z,?t� �A�;O �u�d��W Si��	�B' �/&t�0 �i�u���K�����儙(�� A�6��I�&��:�����' ��l����>H�V�1@\[j�Iv�zK 7S��D�$��=�} �N���� T>�B�1��~,j���hVH�$�9��TUW�XS�<���$/Oe�y( 0cǠ2�u �!{
�X�B=:` ����� R�u �/1 �BS@Y� )�oE�; IR:<Z�d� 4t��pD])��⅀�M����e4 �8$��s[���\ܺa H=�� �?,t �C	�W -�w o���=H�N�`�8q ��?�襔6 �0�R=P�*�8-��.F �$�:��� /P�&�,��G*!ɏ^���"��!��'G�g�ا���
�����?� �%��	R �_x�]� y$I�2@��z� e=
tp),8t� ː6U3�/h �;�ГS �Cts�� ��\�ػ� �dD���.� ��7Ȕ� P�IQH=�>�m`� �
�[�tw�o�`h_�� YL����G 9�uCe�S�.	���t�� u�"��N�� h-��d�> tH�W�p \]�:4P��~ ��3D� �I�1�$� =�����	 ��#l��_?"%��H`�^� �SK�0:3�>*x B��;�~@ ߸>)�'6�(��`\b Q��� �}����@�l� !���-B��������M�� �7���}��膵 �縧�� AE@���HY#���t ���zմ A�q�=*@au��$��~ZH&� LH,"�� O$
bE�D� �SYF ���?2��� ���ND� Ȇ�<@� ��A�0���r8 |��²�" KP�d�<8B �7:R��� );лkY�� ����P� W��ߚ� �&�Hݤ a�w�  7t>�V�]� �s���@�����LP ����� �{�
u�� '@2�_Ї �o�>�# u�8@tG��X%4� ��( B��2��c~E ��-�b>  "up�nH �&c�Ӆ�!�8lA�/�j	$�C��+v��`P�4��ط�� ;1t `닪ǙX-K �SR(�H�� T��i;�o���/pV��$� ^�Po rti�ns C �py��gh��( c~)1983 ,N�/2mܫ b��F0� &I׏��3 \jD�.��Q-J�I|��j� �P�BۄeXx`�֋ U�Yx �)��N�� lfQ$EA ��B�u(��LH�v��Z ��+�n�| )Lr�D
"~�*'d��P ��	�� Z����o�- .�u5Fҋ ����ְ�y� �^�
�	�=)���RK'u .�`N�g�鰗 ��:G'	� �A#�g��* Ex},��pN:�PSU0?{ �C��~� x��Νz���j&p� �� "���SF ��i�8�R� )��*,�h.$����
�^$�&< ��:8��.�� kB��9Z)��$( �0�- Rf;6b 
[i���P42��h��:vT"�� <��B �J�WPQ�:�@�`��X�5_%I����p��=�8������y85?�A<��� ��?ዂ���0��Π�O I,zH3N;& $����L� �Pйe��a B��;�\y� �-P�'�Y �)�X�?"΀�_�MFu ��!�؋K6 w~T�c�H X� �\�� O��R�q
� ��5WQF~T P���L'� 룈A�J� ϫZ0ƋD ���R,�� *�TKu� ��Y�JZ �X�?$���r[ '�e9СǏ %�4h��k ����W�)�8w��R��v� ��XJ NB_K��0l������Z��`, 8 ANÌ:=���������s '��#Wa �ւZv� X_�%e�(�P�B�x�C���`u;۹q, b�P�S���� $����k�)� �[ԉ� ���-�X�.�&J| 9�})Ӽ�(��� ��K%�1� ��x��U �l[����X �wQ+WR�0��N|* �$}&C ~")��ϳ��\��:� ��RC�� ��G��S�@	$y1� �O��h �Jx	�F��~���o� ;��`*t�$�� :�A�}Hx� N�Ԑ�1�>�Q����#�x�ou����	 
�.X���p���0w� (u�Y2�L��>9 �|��s���P�: �&Ԗ� H]ۦ�)���D Y��[� ��F�ո =��J O���2C�$o)��<��u?V1 �j(��w� �8�
*�M PX1t]υ-8l���!f��24P�B�AX�����K3(P�;g ����S���.*c۱��2Q RN�+ib�� !`
P#�@>�� Ӕ(Z"| .��BS���D�L����:| '���i$� �.y� O�ȓe< �G9}`x��
td(����P{ �6��O �(�� �{��N�����E�K�@�&��2U �ՋT$.
S~\� �J��+n:�R=�\% (�-N�� J"��*���*/M�G:��ex ݔP֩I��>F X�Bb"{�f��ؠ���X��̠��
���i�ۉj��# x?s���G/�	]a���� 7͏��Rp ��5h�� �PC��u? Dҏ��s9�I�!& ��VX$� ����d2"d<�_ p!zɊ��O +��na� �-_���P�B0��F3��/r��a�\� �!+:�`�4���� e`��A9� |��ok����Q )�~� ����ڻ�v% @P��
��'X=�����U�����	 a�T�)]�b BOY�/�}D �}�-Pl ��"�4B' [�	���v��L��Đ�K1��U; ��ѐ�@�R"[�?��@�:��G ��M,� �Y�1
�
h��� ���l$q���CZ,a�}!��~y,0�����QMuCp��2�@�x�z>��9���(8EfI�O"���i�� w��92 7B��1��q� i"�G` �t�:��T(f�F?���4c�
�� ����Rd� ��aP�� (�s"y�Rٴ��$��u� ba9&!W�9�(�e�� n��Eͳ@�U�[<@/ S�k.�� �$��P�� �B�j� ��)3Uɮu�s��1� �H	=�\�V ���PV�=3k <�q[��^w�Z$�S/A�]Я�� ͻ�)UW ���Xİ��xR��۲ ��ՠu(�?��rZ	��P� ��u�% �3��8�_" l�J^��B��)��I�f?�8�*PRP�Ɔ�s/ ����'�� H��ӊ̰ZgX` :�sv�;O��H��f� p:l~u@'��4X���= y;
	�)�"�݅��2� R�E	��N ��/d$J��~x}Q`ǲ N&Y1�؍E�a ⽧��SP-���UJ��� /�5g�Q �8�W�}�X�+������;k ����L� #�qj-��N�ȦLp�d ����g�A MoF���S h3VP�ֻ �� 94�vD Q[�2�
��Cd����4� J�}�'W� \QS�N+����0(�Vʟ� E�;L�}�lOf
�A����� $��Q��3nŦ'�i���w;,�SK���������7 u�ۘV�zfY=�&�p��B�6����D`�1 Gi-�X��'����a[4^��iC̩�����B
".c+,:���� ��Ζ�W[e�9�#D��� ��1�*%W� 3�5��� �d���a� 6l����o�b�3$��Y{X �D��px����ىJ�w6Z�P��Π~��<;�Q��V`F2 |�z����="р]��� 8���}���9��'ܒ{���YT�<���w	����O(�VD�������Sc 80��3�pY �m�(~� ���b;<x@=W��$����5 �]��z9%�A�:�t ���U�>���M�+� �E Z��U _�%G���^�K�'��� �!i��򣓐� �*V�AC�� ��3�! ��P�.�R cX�1���� UO����b &�8X�� �u�j;x� +�P�~l ��)�T��}�@.��!�  IO�7|" G�:p�KLa �������"/ � Ou� ˉ2T֮�u� �����@�� P3�HpeI ]�����; T/
�dP#�GlXv�0v"aۄ�@�t�C s�IZ3K~ i���C� ��Z|X%[ d����_�p ��j�J�P ��|�/ �IunRV ��Z߹�  ��H�;B�
 f�� u���>2����p�"%� �\u��|�� ������� h aL��?��t��k0!��Y<��S�� ,/���f� wPm��U�� �K�CE� L<�ƀ8�� Ax��� ֩�
�:f�;�'��:Sj �ר����丂�+u�&�]�wX�P d�R;9�y- �p���B �����a� �@PSH3R �5d���W�`�Qtq���g������ ��,V��@r= NH�(�53j\C �+�@�)`7.�^� Hǅ4_�� ��)��k ern�l32.d{@�G�tLxo g;Pa�hNmTAH��0U$���}�E�:�3;�,���h?s��N@
K���tr8 ��urH> M�,$�< ��ʲ��JoB��@d�Ŗ�s HX�K1Ph<ڳ=]P�)M\6w�3�I�2"C����> ��+&� ����D!�
�/�}��������� �Hm���� ��Ku.
Ia��X�t(mC=�`QR�S�uʹG���F Di��U�&�  �sE�Z$� ��`�Sof tware�)L  �c���sD د��h)# n������ /�(u�B� 9D�!{NK'��T�"���Q
L!o��9���T�˔8 �V�-x�Q �{DIO)� �X��;>h|���9�u��PE�����a����U �u	��S��-�� ���dt���w�t=�{A  >}^*,F �fC	x&� _{J�/<�o
��L�@)����� ��ߒ	�}^ n�>�Q %Y��m��(x�7�V����� R��' ��]H| >�/��}m {���cV� ~����+�A Ҥ3F� R Y4��,�a?����[!�u ��C4L�F� ��7-�EtHl �.����K �������� �F�E��'#��)����X$BP��Ȁ�~ H�NE�e�� 2QR��F� ���d�<� @��~U� �pΣ��N �P�6�Q{t �D�-�s ,�\	�P9��Uy�!���a-��R� ��H6G�Z�$�Egn@�
L�� [@�!��+®J2�.�F*�]�"�}j�䕑�a����^�	+胴�D;�d��� ok&~06 u��D��^� �|�$��L�O��v�b��/ �ۍ�I�u �N����$� 0P� 9d� $�f��b��o����
���� ��W�(�"X`� ����S� �é �� ��g�k�)>%�jO
X؀�� ��wHTP��Se$���Q,0)_H�G��UL?�	��x%u��L;�:s���� �H��B_ �
��3A�hFE���DQ�LAt 
���PvB>X��r���@��.@�� �X��RLB�CH������{L�3 QS���� ��H{	�&\ �9�K+� �I|�B<������} ��J+0��FYz �6[� �B�7�����8�S9�¬i����j�= l��u� H
�`'�K��C\��x��$s.��c �bI�v Ɖ^�V��Qi@��f\vy��oݾ@�C�� ��+R�G.1� ������+@E�j�A �?Ht$� _�3YX�&� z'y^=��:u ҏ��XZYLI����Ww*��q���J`�� ��@~!�� ؔQ�4&[���<�ue�����`�� r3�PJ(%�"��+��~ WѸډZ��[C�� &~ VT�4B)�D�5;a�}`�0�L��Ä� �'Z�b��ʥ� ��J� mX06�*Q� z�U+�l Z�\�IL$�-��r�� ڮ��I Z+��-����7�д8|HtE=��� �+������ ,U<V����艹$�b=�rW�1��̀	EP����H �BD�����1�R����� �-2we=�� p���
�?�@�B��wr�@�P�=G $�����=� ���(k�����o᷐#�����*�X�����
��-���1�_�� ��� 4�.��� 7��v:k� �@�K#�" �>b���x8�A �z�&�8�D ��n2x�8�H �W
?h� @K���� ��N蠄~ aQY�R�� ����o�U �: �'���@�	 ��x9?�\�=���6���_��wNg���'w�'"�E� |o�e��� p+��ŝi�զ��I�ox�@���`�� =A��� H���Ъ�� y��Bk U'9��p�|�0��<�\����Ď���R��~�QC� /j\� &һ�v���)Ǆ�0D�
� ��'�v����������Y ����@��d8E� ����Jz���bu� ��>�9F� �����n�u��`v�HM���� 9;5���S�]= `���Zp� � �T��7~a�p�%�]���pr�L'� ���݀n�8� X�R`ĀM�?YՐ{5��{a�*����ӻ�<�Q�d ���	� �Y'�
#Ur������\��L �u�� t����X� y
��a�� �3�g4�>�ۀ�x����[u`����� ����;�r w��+��@���[���t�F�(o~��3Ҁ�V��d#'���u�����[��LH� ���7>��,#�����D/+��.����{��v�]Y�d�`��W���rZ�����s� X�I��3H/ #�T�j�KЀ� | �0��.���X�*> ���� �¹:����8��H�W�����Z9 �:ɠ}�R9[��$�@�7�5N�, ��
��w	 E4j^��?�3���)|x�d [�B�W]h D\��- xK���"0����`<��BdCg�f�o l'��
	)��2&Vk��Z�]X�d�����<�W�����t S�ۭ�"�&P���A��~�C�,�G� 8=(�
"�?A�N�K\���P�0!"��9ԎGH_��S���� C�=̮�}~
�%�� (h> j@WL�b�>� |�(S�1~��=��,���O �eg/� "�T�� 1(��w|�NE�*'y�_�)( ���X- �ToL�1�(�� �`�(d�k,m���n4O[Ƕ�"�z �و^S�������H2�� ĺ'i��A�	� ������L�� ���%�>in@{��N���uzz�$ �ɋM�����?=�x��!Z �M���15 �=��AN�$?jt���MX^4��)�	#T��`0���  @��<�8�4$|0&[(�$�;� �@�r9yc"p�S�h=)���O\��S)�"���9�ЖH̼���㎼��r�9��*�#���Ș�r�9��k�ƀ�| �x�trp9l h�� `�\�X�TrP9LH��<�8�H4�rD9�؀B�#Б����1�w��rp�0�*�#� ��Ƞ�r�H9�0�"�#� ��Ȁ�|rx9tp l#h�d�`�\rX>�T!P ����� �ð��Ht� j�@.��K ���[� ���� �O� ��h�� "����ԙ]�	"`� � '$�Q���X�W��	΀.�b4q���������P��#�$1� ��r�9���"�#�������w��xr�9�7�*�#��?�� �WT�F_)��뀗���	r�9�Z�#ґ�߽ �����r�o�� �#ܑ��� ��r�9���"�#đ�����rP9�ʀ�#̑���ϐ�����#���ȶ�$F� � �#���Ⱦ��r�9�� �#� ��M��ie8�!���p	�Q��L�1
 	TFil���q&��h?� S��rch}R�X Z�oi|1 ɟ��}E����9
� f'(D� 8p�I^�} L�	Exce��y"?`f�oj  �eh��G� EH�+p[���\��?<�B�EOu`tRMemo ry�ag^\ �@���  EIn��r�~+;pX� �f�t�T	al��8{X0�� $!\B�8l (Gh�@�`Q 	%&P���Xd r��
E:Di vByZ�o3��f!�޸�R ange10i�ҝXD� OPv�flowJt�]�$@]�M�W��	��X ����J�v idOp�+<jX��rB�D������J��zblE:a&}��@@ UnRdY
�DkX���;�� `:Poy��W�\y�%�0��C�st�pW�&�p�EoԺ�Xء�lP�g�p E.Ac�s WV�laɎR���`���H�PrEylea�m��B�
� LStack(���@G�l w�	"ptAk�����^:X�XK w	Var��= G�3\RJ �A�e{�FIao$ I��`��yb� z!sX��(Wܛ�iA�fe���8�ۄ�o;��(a".� �p��iR% $���k� ��f��*:�2@T��˲ ��!��s��Z��䥭 �ij'��Kh S�o�4,� 3���'IwM �>į)lm� �Jg��N��� BY]�4� �ԧC)?ǯ� ��R7�� �<�I� zw�, x� BFK*u�f $�vS|�	 �����R���9�v�ߟ ��t *�^��Zhm
�.�o�n P�p�v� 8�t��� �)5�[�%r���Pk+��gop�j�w' ҳNu���� w栽�D������v��%;�|�0� �`� }
�ŵF� 2N*7&�l�� +�A�3s�� �-\.��j�ꓕ�'�޳`º0q@ˀrL_��"�5%d��� f������ Am�M��d �1�]���4 �(b��)�T=d� $�߆� �uU�;>�� "8.*Kx �d�?:E�� ��������
N��@Rw� ��%i>�QC:d��\��N�ġ'�*�� ��_Ce�b �cxQ��U r7S5-�Z{4��j~�kV��=3Ӏ����)�/A�Z>��R,� s-P�KN�0p���ZT �J=�	�� KO�H24%�Bu�]� p�Ƞ,��� �[ ���|
�Npm*V�ޝF�� �X �b
@�� ���B� {�pO>��u�?u( #���TB, �fgS���d��8>�1�=O�94 �SD��� �{)X�O� <�	�ـ�� ҃�>��kS�܇��s�q
t� c��o��@�Y�b� Z�U�D���jǰ�Kt� �f��wF� �~c(�\ >�� +,g�Y��!|���< uO> �*�G�.D�;"� `Mtw)۞ �&κj�*/ +y��Q\: ���kݔ@�|@P�:uU��$<��^K&&N� \6uFW@3��O�� �6 G� �}�FL.;|�b#��NU ��$5.�� \!,u��Mq�<) �Z�X���� �]��� T�R��9$��K"�ӳ`�m�u ����L� o8���q� h�M-�v ¬�)��������'�޸�tB��w�df�u���� �`]Ӱ� ��Z��s� ڼ`�p��]�r���V��)w� z}�֤+��.n��N �)��� ��ݽ�tc ��	���0������)ȉ �ôV7��4 ����t+.<�q Y��Ѯ8���!n�"���^�v<J@`��?�� ;qV�����v�e�D��G^_ �Q�d��NL���T��)� -��d�Z�] ��%[b�'�(`*-4���� YA
f;�pV��S��#1H?'L#�$�F�'X@ �+�W��	�� @)Ю�ԃ�e|x 2*�S�D�o +��WP\ ��_�I�cp �u.�H� h�`D8]%@ ��LT-+ It.�Β߸ )�1v� ^�A�$' �Ȑ�Pَ_���� �G���9 c�N�)��30jח�0�� ����
���:�N������p� }���v ��!N�Ju ��A�K�y� �j��#f� �B<�,�" ��R	 �@!eT2� (Y���bo=�7� ���2T�_�]ݩ�`���b��@c� � I�!
9ΰ �t%��XD�?�+�s �1��f����@0E�- u�1ڬ�m i�J��y
�4`%������� )�q.e)�&=�s�u�Q R��Zi�J�s�Vۘ}g��
�����4�`4��'^#�K�V ��
R`|�ch� ���w �*t"
0r<9w7k���8�x����J����X ��OS�;� gw��v .�$�3&�t��O���߈���9�C�;�RB\@�� 4ް��@%�$��y�z��={ ��m$�H���zq ~�!�	�L�$��� H}�h� aU��M�>)?Ѫ �,�]f$� =Z��9S���DtJ
U �*Xuй� �A#�C=� �t&�H��[��vj�"�- AN�Õ�� �u�Qs&'y� �( LJ%Y�~�,=:��2N �"WI{�� �	�uʍ,M �(�Z��$v9�x:�
4�0����#��� =�ଓXa y����J �ɟu2e�{PƎ�>�G �S���" �E�o�e������zk ����B1�!���M�����5�8 O9���v !�3q��u j����|P4	�t���q;M�w�@J"P `�*�0%)�7O�@C�_ AP D@�-E� �bk
� �$�n�� �Gt?��E:�8��F���N��>@M���4��s� 9�v'%�,�uP�Z����� �������w )�DSP�}� ���F��բ<dO�b��U�Xc�=Xw� �R����q� �pcZf��2 ���0H�hrg �4� iM	����� l߳�O)�9 �����㢜�8� OEV� ӵy*k��+�;�}$���� uFMn��� ���Q{� ]@r�`8;�|C@0��� *uN:KX� UGR9}�a� �P-��Q�c>��[��J$ �?±�k�<� 3�1M�ȾuU�0"@�Ը���s.|?�w��ę��/�l򼀡CP��,�D jv�i�� ��HP�� YnD	�%_��5L��� H
,Z�6�U	�;��� VB|�E�� �csM�<�G �|A ��j�:��i�� �6���` o�R� P�n�֥
��� �5�~\ �����^ *`V�ˤULXp* W�&�K�. �fNy� {���!? n#-��+D��G�Ԟow_ ;� �	�G6�K����C��u(5�m�R�0 �fQ���S� ���3E! <�4���'�+�{W9��\�9�0�4���[�X! ٠��d�3 ����o��� *�@�t�Q$�T/��d� &l�f��AH4� �a�od ���@e 4łU�H�}7�h���!�=�'w~& a0%x� ��3�l?� ǁ;\F�wb �H�~0�fAN�A�u�P ,�I)�������i�m?�X� U�q�+�@9������b��
;��5u��$�Q �Kt�i)`�� �RGӈ�oq����pH<�� XǸ)@���?��ՠ�T^�A���n�h�%;+�$2= ����L�r�A :�I�����`|�� ��q�kR }��)8L	�����K��u
��wM@ :. Lk>d�tU�9*� 7�@�R- `����� $�)Kse,P]�#6��'�?t�Ŝp�Z=�]��;�r� )@�߾ "8��6 �&����R LDZQ�w%4 ��q+H@ p^5��b0u� ͜+�I�.���@���J��HsOP�Lm 
q�Gȭ+|���6�P|��� �n<���\�t]�� m1
�TML����dS �4����+� �z�{��a�;��<��o�C	��T J%�v_i�F��Պ�kĳN(ݬ� ��r Y@� ��q& j�?��-� �U�5��k �<(�1!D �9�K3 �RHM��S ����� ��H��	AX���t���/;���BV�xaW����u *��@/�� ��H�P�L�)?rՃ �@�Vt8  �G1�X�P� ?��q����'o��E�8t��G�TVn ���Q	 �M�R����B���� sf�� t��D���� PY��m ��]Hh��� �쨊�2�'<dD��VóOv�C�Y�� �����+8�N�tc��3f� �5DG�� &#�{We�"�Z��q� d���F=� �auTH0� �'7���9[?	�#] =Y�p� N��Mu�� �*#k� Z)�c ��3(�	�❅�>���� k��S����/(�g�!lBoSD@�f�5 @��a�>��'k��!�IzBt �v�u@$�8w0�SA&P��6H�� ������|�y�?-�� ���H҉?�߀�~FI ���}�� <�7
Ѹ �����R� |B�/��&� ,���L� }8���f������7�	ȥse%w���Ar�-LO���b� s�2(B� <��HQ�Nq�UJ� 5�`981� C������ �$���*- L�8sC�}�j:�9X 	 
������H��u��t �"���D �A�r��3=iS"	�0��=s��Ǆ�����# ɭ-J'��z �I²�O$ )��#
�>Ҵ �&ڍB�r,�*� ��/^-?�؂�u�o��H����t^��$�a.�a,�� eĩ�q@j�^P�
t% 9�Fg�y���w�kT��/ �J_[U��* uW$Ȍ\� �4)�v��� �!�&��Lu�Zz�m�� F�>i���
'�|� ��}H} t{@��c�
 ��^���s_wag��`�S �}��uM� �0�iw�굘*�P:��x "4,uJ�����݈ �
F���Y c��;�İg �p�Q�� ��,~��X�B��ҁ�ܝ5�P UR�.�l) ��O0I�� �W��R�t1 �b�U$u�5E��P7�y�f���*Ē� HNl�uZ( ��r�J� @
�I�\ �{$aJH� �^�=��t�}q�>4��s��L���W@8[!� �.,/4zm ��H)D$�;�[�c@��>���� �ج`�N��@���� �K�$5����U(�hOH�<�P �4D�:�u �5�_^��l�PJ%�Y��� [���(:�) u���U��*�Z:R��E�.�S >Xl:�n?��j�qfN `Dأ� Wk�� AM9/P�; U�7  �����H�� ���Ve� ]K�$F� ��x����.��3�M Ƽ�1/8� �`CI\|!���'~?�$@ t+3�� [���^��;�pv �|�  t�^�d ��)�%PH:[����v�����]d �3���$��W �ȊT> ��0C�d��(��D2�, 
s��P$ �͉�;~$���*\^���:+����:�0���%�U����k�� $�����4{� �:�֓�� \	O6�Y� E�V���- w`�C�!�$s �	�� �Mo(��Y�=j��Q��_� �
#IN�|�J� �:�2�����xZq2��e�\�F)">���, `t���
���t\ ��� 	�R�7 x�G�Y�~ d����ݐ2 _$�1kYg4F�pV5{ )|#$�e� ����	A� ��H1���75�Ԁ��m)� ŕ�fTZ�pB�KP�d�	���آuҋ�n����� D�<u:�� c$��ew.�= �1��3�+������i�?�@9�xp�1 ~�X`�	��H�|� Zé,�� ȝ�� �@ �䚞��� ��0��%E ���D�I �GF1�v�C����_�`� �-gu�z� j4�7�s}% I�f,�& �U�!`3 �kMy��0� ������D~ F&@=Ɏ�xnU�W��� q31	�ӊ K/�� �^�$�l ���C��� N�|^Gh �,tr�E"i M:/�^�1} �&�A�� �������S6!]���� d^�� &� ZF��K �,A�U;� 	�HM��\p~�jD��I �b�� +��QE�	Yyf����vL<u�~5"`��/ �!���
�u�R ���� I>�w{� =�J|[����0�7,&�E�<���2��� �\����1 	:�� �PdY����HT�'�2>��L,�U�Iv[t*T�<�R��ء �u�r�� N��U��� �$��,��K�2%�UpÝ NXJe�"idUfD�#��zL ��_���(")��g �`&���@��t H�*�) +#�a�� Յ�'6�$� �xN��_�� �%e��EX� i6Z]H��p{���
�4�Pl�G?�����1��C4 �6S��}�;�$f*��` �w>auI���"��� �
dP�� �D �?=�ޜ���].�@q����PP��� �1�̍*� E�{�2�] �-A|�� +X��)�@P𷄅��*�L�(�f 	I� +�� hT�~A|xuݕۤH��� y!�4��)� Q��͘. ���rE�.#��K@dQ1�([�����8!s��m;7 	�a\{O �"~t�-2���b _v�B�z' �Zu�(�� j�� A�£�{�/~���� ��K�j�E �&�ͧA�Lk} ��'v�[� ��od7l�yNQ�@�D4��);$�����#�M���Uj�:� �T!�~_� C�H��JY��5�>� #���8���R`C�b6z�v �u�aDt" �,^����HX+ ���@��V1N+�q� K��B�!*pI bQ����l�su����ޙ����-�c'���L� �a~t� �<�d\���U
� l�'�s�Iz� 혒!Y� �
SL�,D�H��]+N$�!�bЉ��>8��p�� vY���] w��aHP�:ƹ�)-��f� ףQn�H�<9��Mt
�j>V0�PhƄ�>] �Z�S�= �.�\lVJu�jb)�Ƙe�N<� :B���{�,��1���-�}���� �)#/Z=���t=�	�� ��=k8�� 3�0�����^t�5�# �D�,G� � �?���Ty� (��)	Q `~���R��Y	��ky`�$3! ���N2��� Mu�����m=�( ��wT)���Ln� 3xC�~�8�&�"BH�?��VSPN�\v{0,Y` u7h�| �!����΄G� ��7�M�g�|��e�-n��`�� ��Oi�/ �y-��sP ��Ĩ�]:� ��'|L�� Z$u��c�J����}�;�T������%� �f�S#�� a)�Oùg��Q��+�D3�\R'����E�B���} ���f���H�(����� B��Yu !��\�� �Sf�K� '�.��d��/��U,t$N@����[QAR��K��-C�g��^�0=d&� 2�$�׃��H���ם���>�����E �VJ���% ���Y��l�����v�4 .	���)� �L$D�sB 4��+T@�Z;S;$��*n��8��6jJ���| *>�	h ] 3�(H�ʅ�h 7V	��\��?��a �Gg� L��۾*Qsi Y�Ej:A\r ɠG,�1nMd��!�m� ��s���.V~� �|ʀ+�}y O���s�=V������;u+��	��P��� �i� 	T���G �y�*케3��;� Vc-��~	4��E�u� ���+th�f�����4-$ƥ�Tp�� x*J/��TpYZF��X�� �-���yS$)� Jt� ��r�#��(�w!Q�w0 �"OXH��%}����S [�+{�ф J�%�2K��/�T )>	�� ��~t߁s� �.�,}�K ��Fvc���}�0� �P��	U�� �+�M�꿭 m�q4΋� [���n՛FO��U`QH���_� �m«��� 賑c`
��OG-�� ��l"� uz��h���� 4n;�Fj����x��(S��U <�`�4r7 G�5�(a �/%�NH ���l�����	 @ !�0ǒ�1 y�&�Jqؐ �	jT
d�2���>1�~� N�X��&{<\�0,ݴ�p`sj ��C�,& �}�#K� ����d ��$
�� �Mf���J H�S��vP�.��*�O@�D��K���_ ��R:�$:ɞ��s������ �W�d�B�D����Cʍ$��l\���Z@��ȘJ\��Ĥ2�1����:��� ���R4� ٧#��) c7��Ջ�W;:p�X�k𴜳����< ���� 	�إY� 
s"ê� 2;U֓��� 0��6��t �N�S,*�[�D|g-�]$�Œ��5�� ȥE����� ����7�� 3!��HԹB��"l��k �p��� &�B�!P+o�t@j����2 ��zP�� ��@�l�}y����� <��G�e^ ��d+9��!���� Yo�~�� �D=
�@ 	��.MrL�&�V"QI{�A7��J����b�lB��3�Pz����� ���ᵔ��T�×F N7����  �!<��	Q؏(荸� <R�� vn�ӎ�} 2lėf'�< �z`��&� *��$Ln� H��N׿0��|����" r�Vg,�&�]y I���A ��u%�P ��8�6F�� ��_^k� HO�gt@�C �J>�\�A �3�X�9|��<��(�~ Z	�u�� _�%]:Ty�� �~;�<���X%3�lB,|� ���X�>�8�@�F4}�Z�),'^���������n僲B�L� &!�H[�i �h1|�u �'��ɳ�Y����y���4�G�
�0�J�b�?=�6�~7�P.T� � �A!��K;{�g�A/�Lz D�� n��O%:|dF���	��uh� &�gj`P}&��<׬��3��uKQ���Ñ _[���Z z��+�G ��/�J�`{ $i�U^b�t|�폀�}��r�������
�`��+�g�?A���n� ;��#O�� tܰ��I /����*Q'(n�C��G�U�;	�+]c�����/v �j._Y�I! 5���}�-� �(�'ƥ@5��4�� S�`�gW��U�9ז� ��ft�0� G�IB��u�������w%��8�� ��C	���F����(�/�X:�f�,;�69 >%Vx	��� ��NXj _+Q�����qR�*��@^�/@U �4#����%�D5t \* �rC�!d�Yу���s��u��J�
 *:��� ��{,����� �I��S�����P�'�~:���k��G`�²��d�\P���L��OU� �4D� q>'a�Ċ� �"[N*���m�SH5� ��#N��n� q�"�� 
�,�D[{E�.`T�J�nF��Q� �/�R7��d��Dhض�}= �R�x!�����D h��Z�?���(�:�=m��5"������U�rb�ȯ�)����R"��qSx�<+��%��:tP�r�'�s�E@US�?#]D]8���1�)�b��Ө���w8 �$���hH!����8N�W��*#T���%�5�!q@��T� �N}�{l0�Dm9/d���<CX� @,s����a@QpBL.h�� �1 ]2����� :R΄��s �	S��"w �z�)�� ��qڭa�� r�h�!@�Ow�P����S��#�<���=�Z
 �0�@�ܥ �|�\Dis kFrǐSpa c�E2xA��k��y����E �I�h��ȸD���pi�Zd��H���1��"�  �)D��A�>�(���"�xd��pL �1h��b`�,X�!P/ٰH"1@� 8	�� 
�p2A(&�Ƕ ����L�0<@n����!@�ɱ�x� xC��(��$��1�*�ȄL���=��^X_�_8_�^��TLH��\���4,F�3>���>%��ȟ<�@�M�$ r�%�70��} :Ȝ���"G�ގL���!!�����G�$���~|@�x��t��
pC&l��$�h#4,d�@� ��)�\��0�X�,�p�c=D�<�@���Q
XP��������� ?INF'AK k&�� �E ����X�J:/�T�e}� Kְd~"� HP���:} ru`�� x���N���-'� ��s���� ����I��u����#���� ]��t w	��l; ��~�� �{�X��( ���:��%	�w����
�u �`È$�;h1�-��m�M ��;@ ���|�X,� ����@����r� � �-��B�t�`p� *��#(f�P�H��� �3�R�	+b�[�� %�)���I k���� rZ�E�p]�U�J�
��u ���}A���#��䀱�� ��P0��2�05�:�V��CI����0�� ;|�)�Xs/�b ��r:�p ���Ij�	�(3���`�H����`g� ItKu�� z��2��� ����	s~J
A��+O�M �Î�<�I ��3R!"� :�v�N`ݍ�� ����<A tQS�$!) �*E���/�>Iw �[YC-���5����x*�G^�`@t� 7 �3(*)�-����=�m�H�F����@�G.�86 ���mg�N :)�5�2�@�� ^٢$LiJ� G[��O��	������]�sO�(8 ��W�L� �h������>,Y��ǌv���~�� �]�
���f N�F=J4t�� �6u  R*~9^� �K��W3�� �!4�� �fq�t�; ��Uwu4W=�
�>���< 't$�"� ���V�^�?��E@� ���:Ė� B�����:���&��fǿ0���U�$��#:t&��<%�.>, r�3��5�19E:: e6��F ���@B5Ҿ 7��o�����U��c��|� �Hq��e�-O� j�u|��� q�X�k:����+� �z-���{ j��[H�* ��)�y.� ��{0� !�fV�+�t ��(���]�c��_�� �|��J�D'�����$�H p)|LO�����J�8�ƀ+���&�<�l��
-	u`��W�;Aj��`�����S��e� H��^Ҁ3[눹���A��  |�3��M� u���E� 
4��~� A�)CHK{�~�9X1�of\5"�l ���L�E��U�~�
� �< �uf���I �ӑxٴ8 �/E`���m �L�.�i� F���%"�H(=u�f�Fh��a>p��~*�@��Cn 闍�.- �?i�и ;��/@�Q�(���\�X����-] ȧ<ؒ���5�� 	������u��{`��k��D �@���4w)f0��\b�� 2�
��� yT���;� c<
�� s���5�%7�DOx���9.w�7 fǡ�1D b�_����%z!��� V:� ��։�S�e�j�5.�6�����\i�-y׼�N��`��:����B|���A`-d��ڀ��� s�I��9	  �x��m׸ �+�y� 4��U�b�	��� ����*q��$_ �I��� 9��0��  �J�"F!1�QD���L@G�(�՟@?�U��A��/����� �Ց�������}ۡ���-ҫ����"a��>��0��
�����	})����Ēf�+ FT�;�t bJ,$��� �FR0�I+XЪCp$��N����H��P	���>�= ?��;��(f�Ҙ�\�� ��H�m�� l�.ì�e  �Ntğ�,H:�>s��)%����S���L� R�u����*�� kҵ����p�(r�Q��:\ �q<��%� @�gU� 6�ӟ�y? ��) $"8 �@�-TB g�D�^�Ѻ�Q�Ԡ
2 ��?׵5w (���t :!D�<�Hs� 6�X��~ ���!�  D�)+(�Z��d�<C��5@s���b�9xt ���԰Q�8o% �=��˄3 ��i<lqp� �ߛ�+��w ��r�/�W� 䕸 0x�"��e�8J6��<l��|�o"`D�8C��Ѥ

 Rޔ�x3����> ��`/��p�M�1��� s� \
�����8� ��s5A qN��#��� �8B�a�� �zՓx��3{��o�`��|� S�k[�����M\�������w�vcĜ�a����D�^uX:N��f���t& �}�;�w! ���> ��s'�\�o H諭u�yU ���!)r<�?̀Nu���X �$zf�U: �_B��|� �u��4��.=&y�}�sn-d�3�|��r�`���z���+���mK��� ���{3�� �v�7�'�:^C����(;����6رv<���@��8r'��2�OZ���Z��� ���2� ����T/�Hyu��B�����vR����{�^���逬`���'���N�P忇0�v�;
� Rw��4��̅��I�\��7�VˈPDj �!K��s� ��U"���� ��P�u4Z ������* ���=�� CGF��+pu螦�`	�I &�x�� Z����H�$� �1��� ЗKu١��c9_���Q g��� ���5� ���s�E�-9�) 2ׁ�|vC .���` A����!�� ��
�B�]� ����<�*0��.�S$V�+P��� 2\~u�40�����,�X ��b>���M~�_��䜟`C��x��vD4��nG /�B�¤ i`�6�� D�"W/��N��0�dX� �ib%,~t\1L�=7'�K��J~� {��D���<� �L�z˔K=p�����ݖ��� ���'�nK� t)~!ǭ�y���,���j� ���#. C2 	�_�A =Xė��` t?9�3|H �����s&�p� ABCDEFGH�I JKLMNOPQRSTU �XYZ8ab cdefghipj klmnopqr�stuvwxyz�01234567�89+./=;(\)��{},;:-_�*"'	 
�EH��N��A�y� _)7W5ą%�e���K C�Q��B�6 �R8)��4�kPbhLoP-�Nd�m]�@s�?S�� �x���t
wn �9)G��<�F���gp��8 
^�,k�� ��Y�S����~4	�W}	� O�� �*�H�J�,���aЃ�(A7,s*{�`*� �Nk��M �,O��0���B��GK Huj�.fD��C�I@���ԁ �!?�l%L�v���q�:0XƟ��h��U�~��@s8p �|X��� �H���?�� ,Ƥ�N�~#_�����se�H
����� ����0 +�|x��b ��d`�0� ��:uF� ��]��?��|3G�����ύ��ә<ÀĖ�t!�;��@�y@� COuӀ} .t��l;?���� `%M	�B�W�'3� Q���ٖ�J �)l/׈���=I"�ǯy�?�+�;M� E�!��~b �G�n��+���@�ZW�ƚ ��&S����=����[Gu � �'E�8wM���b��D� �;J��L���ٙs �(�$ �M-<+� t�T�V 0r�
9v�1 \@�%�ܪ� ��/���  6���"����[��5��-�*�&K'� #�F��'H�n {4`��[ �F���wV %�NܿM$�B�f��d�r �+��W�s:��1>��۶�?����q雨U���× �Xi�DZ�� �!-l�7?w� �h8�i��	:5���'��� �tB���>�V��3��ޅ� ⱸM�� �,�W�G��G0�I:J�j) D��Ƿ�v�^�� r��P*[�g 9�s�|�V�9�����dÌ�݉uJ/�� �<=�Rs�-~]�1�;񟀄N�) *�$�6l@ �Ixuf���E��/����) +ۂMv���8j�)u z���o��8�6� ����Tj� "D��Z�$�� ��ۦR ���|P\�� �-WVxO �	���X�|&� ��8�� ˅$+T�1�td��eZ��6v�����c�B��@�;Ē�4tO�8p��rGIF�ipA��JpP@9��>�U|�kN�w����]/ � �y𰣽J��@�.��ˁ��l�d ��K��RJ| }q�y��� u0Wj�
e  �S+,�$���� �@Rݑ<�s��g􈐓TC�{�� �a�߸"h �s���O� �Է��j pf�ب�t�1��Q�;]� �Bx��S� y�C�!|&� �=(h-�Z;�� ��bE����ϼ�x�1 �3�����J�_jd#@����\|w Z����bxY�� ��}�A y�?�_�H co�j���We�]��0dA ܍MN��% �~��lޗ�,�F;�2r��!�s
X�vD�=��V�w�W��)� ���\�5"L΢�}6���C�.� �Yϋeq �d@\pag�� f�5.syS�8"�in3�6�, $p�BQ`�� �1�I�S �>�0Ȉ� � ݶfѸ �sx	5 ���	����Hu�1� G�Op�[��(���S���a\�u ѰA,X: �H'�Ӿ� �Z����w "KqF��8H ���,� ����A\ �ܕh�Pp��#z��� 'q��E$h|! ��c� XG�H �o)�57����9�X�$�h��ϝY��[`ӊV���sQ`h�XY ��FB��{ �'�^ ՜��6�7��g���{��r�?��O��|/� ���1(� �-��^j ADQ�� �6ÈFL_ s)ѫb>�� �Y�U�$�������ؘϾZ[�d��v�q ��}�>x� Ѕ���4NP��M���U�Z��`~�I�x���/�� y%^�p��?��� .m�9�W�)؜S �o�� R���x߷�?��� ӥ�i�� w��#9��� ����}���vT�eF��~�X���@��������2`�� '=,Ihj!A B5����Q ;�T��� ��"#YF4��0���d(!��
@{��,� ������	�K�߀�m[�>�F�'h��`��@�~� >�T�^����  �ό),L�v� 5�ẹmV�Թ Y���0�����O�T 	gf�;�P�[%r�P�K]>� �D���d�,fT� �p �@ ������}� ZBDt!�� Ā��(��H�^L�?�N��X�1#�4��Y��& 2�x��Q� ��i�h�1"�¡���}�WKa���L� ���ܡ�� �	"�N�� q�
K��� WSܞA�P� {�c���p Da�N2,� lx�Q���� $�2��Oz�&����B�� !7/�
J�,4� ���E�1:��
��O$M<Z��Ad2>�0�� H4���F�:&����_��H^a����)S"6��+� ��$���Q=HP�_��!#'҈C ���%-̹���� ?�S�X� �K	G�EW��u�hdw����C ��2*�#�)`����0�j��S�� ���� hp��t;�? �(F1$E�/� ���,H{��-��� �ȝ� ݤb�r����/>�l�@�2�����p���F� ��%�] g�3�;N*����� ��r�g# �~Y��c1�q��
��-"�U�>��[�� �R�r�g`GTy�	Lib�P>r�ms� ��p� �>S�ٿ a�RJ�UNL���h(|�t�� +������ �J$1`�� �%��y��  6�J~,(*� ;��'�-�8K��,�aG?�� �v�r� ������ 9u��ɗ" �o�zi�F\O i��u��� ص�I)�g���F��;��y �����\xx ����b,}� X�S��)x�r$ �L��Bم�c����/���a ������ i�R�3%�^\�(v�H��P@�B� VA�,+� �#�I�� �������$
�r\b�TB��!��~ 01tZ+�N �-%� ���P9�� ���>�_����� �J 8\H���t� ���%� �\�⺬�� �*�u![�� sA;��� �%�n���C ����o�R�� |�26�4�-!g Z���PH@N������
$s����(��Ӆ;��H0�� �?΀CLS ID\"0�a���&,��X���&Jݓ q�"��&A�!n@���uX��]�$����#G�Z��������� ov�.�ۋ��4 !�y����G �P�-*�8� &Zm�e�QC ��
ƋaR	��,7��Xj�^�����b���ә���3P�_�*g��o�q= M��t�:E#;�e D웺Z9| _��Ĝ��Lh� ��~�줩&�t B�>�D]>d� �	�����1Q�M�7$Y ��G�0�� c����K9H
 ���	+_�T�� ugQ,^->R� %�U�MB�������,�� >�#�E�)  ޡ�p�b�N���; �Z���1&� �G|e��?P%��W��PU�I���D��� �8�,��L��N�e��^�� G���Е �[���Ŵ� Q�O��;���� ir_�� n�}pus��X ����"/� �(�O�R �#86��E,��%�Ć��tK����� D���a���ny�.��JY^ Ô��E�
 ���,�$ ���v1H� �U9�B�s�S_���� ��~���w� 
��T�E ���	l�L6 еX��A� e���~E ��H��	>�s]�8�(��5u� �	�",�I������ ��u�< )>^��$�V 0-�n���� (�Claqs�@rFJB�� ��T��}&w4� �,%��b ��#R��-<' ҃�J�%�FpU +�f�<�  �[��b��5��C��������������>X(F3~넀���� bc;C��
� �Vg�GNu� �T�c�4ϥw� ���K��� �ܑ.�0V�O/��H �[�w� !���el�ҫ5ՠ���a ��G	d��� ��;�9M�P���D��|* �@[�h�� e���0�L �̎����<e!���B��9��b����<[ �U�mt�j i}@���J� �w֡� q� �����%�j�^ҡ�}�Q.a �YfΑ�E u*<�'H� h�2��^ k�f{�[��쓰 �&�"���.���* \�2&�Q�� �%���� ��;E�;u���_tH#:1���;U!9�*�"e>� d���#�'}� N�X.哣 r_g�/4!|���)h|W�j�'"� `?�*S����WXZ����S2�ʎ���Jm��'�Z�K���潉��SΫ�y������)��'�@����o+a����cG�*`y.����
���p�غK&��� �v�@ƃR �1�x�� ]�����i�x� �����Π�9۽� ~<ߝ�@�&�_� K��|�  ĸ씉��' }�X&�0< #��続Ө.�t L�̊Zx �5؈��`[=�L����� �{��C$����]�0�T�.� ��L2� ��N�#* �3=�� �^��r� j��N�_%� �2P  #gf \$�XQ ��Z|��K� %`�	�R* �ݷ��x ?E�
��\�����q�"p�茲<�JԐ�ڃ]̈l�X�N ��Ƭ��$SI���� � �f�x] 	.Q���= ���ִ� *��I_�1\�
��VyT����� @M\H��$��5e٠f�C�w&(ݝ 諾�RPY�@��;$_ uv	��ZX s`��}�$(!� ��Eft ��vWJ� �V�֗cT ��b��R�y�>	���xFO�0��% U���Mg�( �m�Sf/���.��� 1���p���� ��Qw
 z�i/~�Rf �B�"�,*Q �Y���Ur\؀ú5�~�8�" *����}��S �y�=�x!�(< ,�CN0� f����1���{�(��� -��CS�� F;�r4��&e��>+�D?S�;�tZF�H��֝�@�)��E�XZ��FL! 	H4;�vo8�0��+�@߁
�{�	�:�� ��s���w Ɩ!�즛�,Ge¸A��w� ��r.|(�ي�PQ 
� s"}�� D�Ϊ�R�\W�!�����J� E(֯�q ����yu' Z,�+ I���t� G10X�[��%�ȗ��� � ɡ&�� �ةY7t���$F2�9�����Z+�����A3`l� �'g�/k�	��T��^�S����!�}ٻ�@��tBƅ�{���JU�w<h�Y�T������
?� �n�PȂm5ud7৮M1�~({�� ,�C�@/� #���ktxy$��\�+ ��?ĭQ� ����- �<�%C`Bd0�{� ��L�̒��X�� ��һʌ�� d�Y�t	� �|��Q���px������E��)<�w�� TCu stomIni ��f$�<J��z����8�+�������|6 4��	D�S T��R���� ��).�;t>����-u� ��C�ޖ �8�;ҍ%�~����W��"Z�z���
r ������-���K�p�]���d���[:� ��^5�j�'�B���y��7�wG�0��Ҫ c~>��= e6���� �
xu&w 䓵h�����3�����q���Tpӂ�� x1���*� ������d� �����`��>��q�S\pk��E-�`%���>��� �<
/a`�G��Q@w����i �Se�tMY? ���8���#�� �[�F�z� 0�I�1jZ�ɫ� �]�O�P(���H��� \,�� -�U��`��Z�� 'x0��o���" �K��bB�1=��#�~�(��F���m{�����`��͍Q��4���ز�x� ���+�|l/ B���u��G�~fk�6� T�`�����o!��� ��J����;���@�mjd!�r����C�owG���� �O�0���������4�j UK[���� ����L4� ��n(��� b���_�� <H"Oȍ�'JS��#L���Z�jQNv{!����03� r�6���) %]�dV�+� Z�*���-U �_[�(� ��84�� ��"����	��a���4h��s#8B$�;��Ǖ7� �	�z� �Hő�"�D�߉���/�~�~?'?7 C$RHb�u�������� ���*"B<D[���f�oGH?��	-$]� "RU�3S8
�.1]����J �:B��H�R\C�F��"~�!��n�@G�(z�'5�>�d^|.��XH� vՒ��jÐ�:�g?J�[E��Kz��Q�	W <��9$($,0�4"8~<���w��+)��5 ������ ك�)�` Í��0�,"	�D&#� $C�G甀��s�����l�� ��8�Y�
3;AO`\WDTQ��+_E��#�� ���j��u%no�{� ��v �s��$��@ ��n��' w�T�%� Q0�2�]���c���b �?6��f �	*W!ʊ �:F�1��sa0�E �e��>�:� htH��� )o�F�d43��*GS��|� 	\"f�)�� �h-�d��� Hȑ�"�D�����!��n �㏦E��$�]"��Љ��$���� �t1��;� !��D���H�������$:�� �&�2F	�L��6�n�� z�)]Lrl �kU�C\�<D�n�8 �HBLx��PT'�O��X�\`�dgh�l#p�t��|@�߽�!�`G���&� �:��1� ���x�gLq� �����G@���dH���6#�� yx|�D=s�h�� L
Xy�N +9�vHDl "�P �B��L�p�T�;@����P�H�XH� z��/?!j�9x��c�<��NZ�X�|D�2`�@2u�`�@l��|j �X� M �1|�C�� ��$W�\E(�,�9 0�48 ��eZ�{@�� K�����< 1������$`5� ���#�f�.�Ȑ�p}��̋� ��
"\��zơ�йhbYK��]�� �G�F됾 )�
K` \P_��^2W���o���'X�$ BK��� )�<�^LW�@�b� '�>Hj�K/ Բ^z�_�ZK���0"D�H lϏK�_��B[�`��D"@�%���*?�^B�=j@L[���2{��P�Z�~����/�!����&p�R}� ���a=x�%L5�!���'U���� �; �����H�$�I(�,�~0 @4�8��<��T� �L��"G��Z3�sD�d�@9ǀ g�	j$�y��(r� n<,:�O��0 R Q4�h�8���< ��[\(�� ���x���|��.� [(�,�4��< �k�h��� ����i� ���׫@J=�;��v���D�� 
����N�H$����@s �S���x1	��W TI�� i�Xg�*+�GA\��y��0�W �+���@r��7�?9 e����;��C_�}:�o��vjW k�4���h��V�O�ytv�o��j�L ��� ��
7v�xF���] ��ڟp�� @q|]-0��ki��I,֚;} �].��9( V���H��� �C
�[����p� A<6D{x�0>5�0������q�\3��8�"=	�XA �60�TH�,d�D�Ap�|����t�C7��|� 	�1��2� �G�!��C� �13��k 8b:�1dG��|$t��;�
K�=��#4����E� �`L�h�l f�X	��� _OR16ؠ}8�l�j0� ��"9CRA�St����r ������5;
�8g �S��u{ �����>��2z��I��D8��T����K�F��:�k��/� q����Zа��\�A���{�"W� �5�e���C����Jp��D�Ah����pP@T��>#��� ������:wu� %��A�C�� ��#�{x($���|�����: T\{.t~#q�?E���m�����?����p(���zs���9:�� a��se �;rt�GX��d�8��FX�����x +���9��DG-��(�eb�.,>� B0ȟq �4����98�֐<��9���D�*�� �y�Z� ��� m���j�L)d @EB��;�R��j )ԗ�	�����ec��j0&���pI����R��� 4B��VF� ��d�H$�! %�+�D4zN�T�"��fya��o���>��? �@(�D�2� 8��d�7 �V!
�w�Q	�1��.B�;4@,��m�s� �C<�:��{�3�n�@� �~\�� �����:���ஏ@	�������=4&�lS)������b{�� 5Ŕ8|��	d(!GC�����>P�)(�_ hvB�ț�$�Í��Q��4��
=��H >
�,p?퇈0�d(\B��`��� Q�3�����k���U1��X� $JH ZL!rPB^Td���m��KH�.��Z�i����G� �H#E`gL���@�V�ܺ��TvD2p X���Á\� �"�`�����d $ͫ�hgE# l- <3���������_x��?�D�@��8~ o+Ѝ$k�W��S�C@��Q ��1����&]E� �l�v ./%�į�e ���E+�� ]��̗٫ R��~w�n��?@^��� �5�Pt�;�\_� 0 .%$� ��O��� �d@VƆ7+ �)�<(P�� ��U�A| wbz���@���}c0M�SoQ_=�@�d�x0�j��`�M$D 6��W ������V s����4� +�i�H@u �13J 	:�p�$�i��gL?�����f��� .���<$� N�ҙ̐ 
J�^@�|��!�����@�*ƇGU�a���� F!0�$�|@G���GU��+�.` �ؘ�i�x�BN�# D�$� �DQ��э
  (�[�a�i,����\�C�!�y0.�&�kB����� (4��q#�����x�@80Cy��<9����!%�I*&��y+ �
b�� i��J�d�� r@���%�i@4�x�� A�QZ^&�f�O����@ ���r���N���������)�!��]/�a�A��(�SH.D?6#3�����  ��)a�7 V�����p���$ �Z�F�Y����H�#�D�����7��⿀6�,����� ���ZE�����@���$�CM7��,��r��!�w�~H?�KP�u�ogEy� ��0��L *�C������B9����f�ঊ @��*���)q�	���@ѐ�+�"a��m���� p�8E� "N�,#� 	3��D꾤>X� B�;r:�0��f�?�U`������(�p ���C��p4�~�Ì�#��＊'��N1��P݅0��:�����)����9���B��`d������m�<\(X� �|�@��� �eV��}� *�D")�@�2�@��۾���&�DS ��*C}�$
���Y �#%��Ip	!�q��;�0P 9����� ҡ���6�  J8U�Y[e�޶
Q���̄���q��p�Q�a}��"��!���];���ޏ�� NO~�o �TB݈<��,�0������C0�~/��4��N��0�BH^p �~S��5�>#i�,��:�b�4'��� ����*��P�R� �ӆ�����&3��aS �x�ֶc�� �(����z=H� �.���ZT RX�|J�?4��%H�9 7(��� ����P*�Hq�4���W�" ��
�O���qT�+��qİ �^�m�#L(��:�R�`<�� }���L���+�F�V��`s��$�K8$\���i�<.|F|�B�Q@�� L� �q6!��d s�8	�x�� 0 r��Bj�|>� !��(��� �Q,x��XF�&�	J���#b��F4I	����8��ȓ �<�$���xz� ����3�� ��lom.-�#��	�ܓ� 괇*
�7����R�9 ,�v���=7 d4��/�'�l��J�s ��m@�H ������ �7(/l� ��G���v�� 	�H 0V�K�� |I �L�lP�7���;��(�0�r ���C�#��o?��`���	 b(M�,�y��_�&��c����X��|" �8��~!���,xci؇����� ��M�;{r ӧN�0�v ��Bq�Hz�n��i�Z�O��D,ugx�:v���4� �?O� 9q�	��< A�(�;�w�����3 -ɬ:B�< �P/�#Ar& V����Z��>!t�\�� �~uF�R����������:��H\H� 9E?(�- B�FO����k�<#r�Q`4|��,���(�� Q��4�5T'7��,�>��#bj <� �V�$���ܼ�w��Ƚ� 빰�7i{�|�>`#�2y� ��7�	S��$#�0 y�K�uh 47��F	�/a2�$�pj��$�`o}�i�Z �g1��0�	���x� ��&q �I4�DT$Y��'E�ء��B��|D8��}�&�<�!�@^B8�x)�9�h����l!�X��9���ߏ0|����@N�S]�o��"� �<�? M2vnX% ��@,]"; �R3�#�t� N�6.`r&[�03 �g�n��'7��"YL3�A�qn/)� :�0���C�~+%
�֨-#Xf<�s�'�6���Y8J�f�����-��ՙ�I= ���bS��� ဘ� +$��,hrB� F�p���$e��ǣ�d<(�~F �?Nu8:����$X�:L/�K��t��\ �^"� �2�>撢P (1BF !
b%�8����H���qYj3a���:&1 �g��%(?�2 �ȓ0��h Z�3e/�(& �.���@�-bYm/p(��|?
�{����{.�҇�4����%�
��>�!-'� �?,�_C�� 4�.�!��nt�� ��N*A���$cVƀ�����-����'(��0x>F�{|`75nC���M\�H�@(���,�7�m؏М5P���?֏[� *e	;)�Hs�u��ym�o��[ ���{����/ĠvQ�.V����bװ2 G(����8E��Ls<x��� �1 �"V��,�?C��0�t�T��>i��p��]�˔��c�Y+�{����n�tDR�@.<V%� Ǡ��>pm����), S3J٢�?*�� ܥŠb`,�������� b�,\�{֘c�K��'���h��>��!�j�-�s".|�)A�-\�֧���Q���:�XКF���pc��.=��B�1�p���,�R�� �:�`(j�K.�dJΥ������	��{������4�����C  �	/?h� \!y����{}j ��o���8L��8���c�q� o���C�O/Ϫ���9�o) ��>�/� ���!����`n�K�=0�  "�D,�B��?H��<��腐��&0� v�kh�� �{����0��������<�H�+ �N�06W��"�isn�DB$/1h� �����n�����4�� �Y	�1� ��9�"�=@�C����{h	�iOoq���2 p�$��C� �_nڦ�B2 �)F7�8! ��m	��Z/ ��2� �%ٚb��\�~�5	����3O���[���/���O3<�v*�� �r���d(�&��p�3� ~���?���;��a�@C���Y���F #��͇�4{x�H��8$����t��H?���%e�B��P��C�����-0�&�e_Y,p� !5q<��LbtpDP �׈�W��RT�/�3��J�P���/ #GH��ctac�0pX�P��� ��'���� SQ��1Ƀ=?�V�}N�- ���6ꉿ� �A��u�?�/�JW�Z� �*�XC�3,�� �9��T$I5u�ƠL����	�`�H p;�}* ����� /IPrn7[�4�vX�	- A���� 9\�SH]�t3 E$�=r�4����>� ��� �O֚!�2*	|4D��
��p�� �ި�2A�?nҀ�0�&.����wh��r��VdQ`�2� ��F4t���HJ�0�h ���(��0C U� #��2u
��x�r�dk� �A�(� i �05�4?�8 ߑ<�!@�F D�H��L� P5dT*��W � X���U�� ��R\2V�� 5�r�`�.�����ed�6~�$���h�.���l Րp�r��x/�^" �$]*�� �j���� !b���}2r>�������] ��#�TG� ���Q��� �%� H5�k�{�V������q ;��ZO� o|Dbr�9�\�WUAj���0���9& ��T��  �%�� H!�=��5b�b�>�� ďX�1�CȼAB���u�^Y����2ԇ����G��C3!��@��d� :� ,�X`�2��!6u;# ���84� �w���Y�;��� �`��bʇy�]5(��pW1<J>ݩ9IE����RP�F�C@��Q �� n(�c�(�, 0�47D8\j�@�#�Q� �F�Ks�P��! XTk�o,b��HW�������Ԋй??�1 �Tn���� �j�f2H$�/�<
�@���A�fN�� ��P����	��3BIu��`x"�0� �
	�t&g �#@!S1ۊ80��P衢?/ 3�]��X_&�[r ٖ���CX~� ��A�����'��$��)0~����8A� �ρ�@
��� ��	��?Aȿؼ� �ہ�@pxܝ����`A8p� �ԁ�@q ���A��r�tv~�?�со���0��8A��3� ��@2�6�r�t�p7 ��5�4A�8�< ����@=��  >A����:�;���9 ����@8
P(��&B)�D+�*A����.�/���-����@ V��$�%���&'���@��"c����#�f!,� �>���`;a>�c����@b)����g��e�dA��l����%`���o�n<A����j�k8��i ����@h�x9�:�(y���{�zA����~�ؿ�P}Ľ��@|� t�uAt�w��ζ@vr��s��q��pA� P���@�Q��S�R�7�WVqW8��U����@T� ��\�]A�� _����@^�ZÚ@��[��Y�XA�߈�HI��K����@JN'�G� O��M�XGp��D��	��@E�����FA�ႝBC�������c���SQR� �����X��5�	�]P��`��%���2@ B S����HX� v[���Z YU٘a!OAL~tg(��s=� >�����?0 �~�< h�d@�"냑`�l�\�� ���a � 7*��:�, �c�0�VK ��6f( �gJƿ`� RVQ���$ ;���rM �0°��sx�����p�� I	��j�_ Z���XP�������+Y�>�u������J�f�����9�� �$�ИU� ;�sL�` �p+�Q=AFЁ��`U(r� b����P�ƕsj0��� �.��yT�ַ�ZW�u��'Đ�� ~_Q��z� B���=�� �G��v� ��_�U� *T�g��V8���(���2���)���>U �a*�Xߍ�z�`��P�O �HNX�x ��E�IU���� ��#�O.%��s��@ �J¹�� 1�8���z9���d"M� W��q��	�c9Ώ��ʸ]�^��Ռ�9������������ ���Ko�%\�B���J�;���7���� ��|$�	.�(�q�)��,�p��0��4�J�@A8*�?�R�<	W~��d�%v�RS������T���}�B	 ,�h>�+�����rb�3�Ê��֙'T�Z(S"<LH�EB�$��=�8�"6D/�� ��( 4B���+@͙A0HM .��3�� �i" 	U��r)P�c��V�M���B]8��������Ud<֭8�J�� ^�R��%�h�(�d��,$�V�J�ӄ@��� Y@��1��}Z� 0�Y?r+�D<Kg$\.�v QI&�^P�Y�A	�F6�1b��
[
��;��ʎ��$��?0z��P��_��$+��DxxD(�1���������^� <�Q�K?�%�J4D�	C��ʼ�A,*��W��%T?�J�$���Z�^]|ONV?�.�j�� A��D�t<�����s��!��Fp �z�}����I�؎2i<
� ;'���	��f�c��3�J��O�.-�  f�� ���^���D'H���٨\�1CX�N�8��D` s
�U��/�aL瀠3K=�f�H� ;r�ֱ� ��#"�,1s� �z	�� ݱ�~ !?`�܌$�� wTel�g ��@��8�� !�
.�t v��f���,�� Y�:���F" ��eX�8�3 �H�0yjp� ��g�)�� ��`?�TVR�� 68�� x5��;�v�M0�ډ��,W1�D��� �@<�V��"8}�.WI a�9�pT �k�����
 RP+}2FE@��o# ��>^Aʩ G��(ZE Ы�-?`8�`}�� Q�b����'��w��\�sڀ�4��H� ��� e��¦o ( �@D�:8 �T=��0l� �\̔p�����Y� H~���aA�"�- u�LJ�� 8�W�R{���P�T ���B�+9��� �R58 ���Y�O%}<��Ȏ`X�� À�ߖ-� �ٜr���@~;s �V�˾���LGnrc�*��! &��w���� 0���[.�I�@j�$��p��S]��J	��_e$���@�)� x}ƹ2� ��a�"�1���m�ӆ�R�� �j�VfK��@��u���4T���G��;�r�خu 7Q,SO4 �_Y��E �����b�8>K�i,%�*���>�P��V=� .��� 0]��$|� �T�� �yu��|/ ���:�eCNu���_� X�EK��:	 ^eZ�Ψu��YLvD�x|<*!/��@+R��5u0 A�BqCV l!����$\ug P$�|�� �x��2Vz��� ]DP�8���y, T�>��j��x� ����ћ���"���F:(h �N_��+w�9W�	lx��*��� ��:p ��] gi�n��2 ���,^+qLzB���	Or /��(�Y̱ QˆU�� uj���^ �KS����f��?�`�g a,ʰh0� ���"w�: �S-P�U�4 ���Hh#�B�^`̬1(��� _e�,-�a�y0�� b$t
� �2[P]�� ��u	�H��K���R}� �8\OY�Xс����`j� m�{��
�(��C�OS�5���#���e�x���L��W�� *G3��x9 �S�`R� ��5�D� f�0�&FOu iف	��z���@�U�֍( ��7?�b/����4��S8� O�(�C; �}���s �����"�C��M��$)�Q@�رS<�u���# RB;H��|@�����ӿ p(���4 �i�����  O�?P�� Q�J�~B�,l|$:�P
h�`� t*3M>� 7;�}u~2���[{��dZ ��iU���>N�� �){ZP�� K�0
�3� �|;P} I�� �åx)t~� a���UP}$ �Hl�T�IsVr�=�<�uJtJ��� ���)$� Q"���X�$�`� IR���=a4�~���@p_NS� �Ⱦ�!�k.�$ �7��i30�$�� ��B(^G� ���g�$ N;�@r��	 ��(�^��j������3��K�S����&�{~ t��ի0��p���}ƽ�~fX�W��fR%�8 X��U� ���^�kG �W0%���ʒ�$ ��=�cR��$�1�J� 'ue�������X�d.�H5}D���b�{�v8<��A`ϸ ��J�3B��p����	�@Y�Juﭲ@9��	+�{z���� ������Ӄ =�eAǋ�� ���H���<G��(,�����Z1 _A����O�7�f���69�� Ph�jLH��f(����� T��UQ%j��3�À���� �Y��<�	�#A��d 1�!Ǧ�p�|ȧ@�C�4 H���>� ,܉ �� �f�= ���˰P �ǽq�&�=������ Ä"k ������q~ �ʠDd �Cø�w���,��`��l�5����Єb
�;�p�U����e' �����F
Z 1h@T׎r ���e)Y��F �T`����G|j�Vň�*�!���n�U�n����X# �lք_r SfqŹG3:(�%�'n��>�K Zl��J�?�� �oL�ӏ�8%݀�D\�. �Scsi���#:� 9�CI D�!K*,M ARTVi� _�hkb�{�[	��M��:`>� (�|c@D� /�x���i���.BfIUu�AJ�Z��X pڽ�&k��:��� 3u���M�Ψ*�P��]	g�=D#NH�T�i���� ���nϕL �}�xCT��i�@uM�@���9�� �D7K?I p�:dN\��!��/��Wȍ�ui }��]Ï 8�f�,0 �Cq��t' ���� �jL+���0�B,cE�=��  ��s �2�{E�! ��,�bRƵ���� t �@�8Fu�CQ` (r 1S�W���@����!;���A�����>����h��i��{�W����	Q��!��O3� ��~;�i�"rT�� �Ly�cal=Dr�ve0�~�P;C:!9�E�8�@�Q�3 0���%��� �Eo�	�C� X@�\� �:�ha�� �[O���� �����L�y�Zu�����:���`5�"� %�.�	�F��?�����"^S�����2u�	p��� ]SEkX� ��_�0m ���M��j
~a�0��̊�d7S ���	,uQk� �D/�f�� J��?�xb� %M�_�B r�SP�V.�� �(��JX �B_��El��jYt��w��X-��KV���f�gX8G�,�\ �1r� �:PuB�%y|��Χ#��n� �7r��� ,��� 5xsp� Ұ��W���& �R��V'k:.�PI2aC>����T+�� jP�Ǉ�Ĵ.�W*����(� �˕�wz� F?6�MR*��`��y��p� �n�)\��9Q: H&���
 ��xG�07��� v���Գ� <@L:�p� ya!���t =��Co ���r�s� �n��l�8��;���1c��TMo deInf�rJ m���%� U\�2) � ���9���������� �L���HdQ Q�'��� �o�Z@	�N �-������;2�5����� L���QC; ]ulBvN^��r�\,� ���M� ~Z�t	m�9rBp�>�� �Reg:s  K�F�Ȱ� ��̧R�+] 1�9�t � ��;���
X�j�(i A�n��.��4 Q�t�:>�Z�o�5� �
 ��%H{���=�2����=���(�0NY��.Qb	wio��J�v� R�U�$�XE�HMD�;X����.f �!����  �����ooV� ��T$� �щ�eUY� ���I�RB ��&t��Xw �Lgh�xH3Ԉ�E�O�$ ���V��.~�
�>��^�@x Jj��%��;9�:2�X;F  ���h/b� ��L�MX�[ �lZ��$+V_�`'�]���^��0u��5 *��Ô�0!�M��S|̱�Ւ�KT~(�Sf�
� Qb�o 	9��􏙞���؀��@p�v� � -$�xW=�Q�����E�d���0n�g "	^��;� �@ � _�1/�\kw�s�S^̨Bև������t� �h�x�� �.l�dW �)_�tL QRu�&�X��?� �zD �v���@Z$��� �������@`�Z��
��+`A�h�(0(�� $&�����������X���� ��.�J(�� �P���a �D���(� �.)tg�;2 a[jU EV��WY
5 -^k ͊ 0�9f�����؅jW��� a`5}���� O%f.�׮ R�g��8����\�3�Bi�ȟ@�)���ʚQ K�HE P�?�Pb�r s	�Xk ���:f1� �D)h�^ �~%�}��8�����H����.���aȥ�L��>� @`bcH	s��@D%.�=Q f�����U g�������� ��y��.!}.>6��$j ��ڃ�#� �.^MU�) �84������������@ WjH�� �ZX�SQ�q ��*#����`"4�s@H�,d
b �:�;�LyB 4>�؃�|�����ܗT`j�* �F�9��h�%� �� �LfF��Ez k*4t�Dq��������k�&<Q0X�� �f�Z��^� ԯ�D�C�tAb�����rI�vw�)QX���Pb%e���(08 #+3H^� �����(�?�� jņ�#u�`�X�Y�K_h�� +	��?�u*s��0fD $պvi5xz.�g�f���� �	,�B"YDr���R��F�;�n'�L���lN_ !���m SUAŗo9-Kkp��q)|l&!� ^�E���7d����*9��?�q�|r� \�%H.��Bh���0� ��PiC��	 �du"ȱ�j�m��M����w� �}��9 \)c�@Pq� �fb,�Ӵ:�t��O�<�
�1�`��@ h�\w�d� �0����P ĉ臕V�4 �[�Sx�5 �1Y���� �i��d�	�H�� �h�G�m�3.pj�:PԀj	g�(�>�s �A]k)�\�ǧe�UhN� ��Q��m �u~3��j��yļ԰{ 8|�}I�S�k��FXY��$ �B���Lś�WS�C4$  ���+Z�l/�� 
H�K����@jF�zQ�#��}��B 8|���R{hrp� �|� �g�$�I��7�x�"�pȦ)/rCK�D��'ϐ�=� X��d�"�*�'������u �q�P�T��S`��O�����nh��b(�G{ I1�pK �'^��U� F�GtS�d ��NzP*��D���͏`�_�x ��^��el G|Z�2�o ��ny�˅u� W)���YL AwSg��^m ވ}4	 ]!+�,@ �M��B�08>>���t":�a� DA6/^I�>� z; T�E@:3�	O��G	��U�m��p�D������� !�jڔ��H<u$Ȁp2��&��� ��,
&�V��	�� �*��n=�~dB��ϙ`�T� -�kXp��.0/h)^��] �{�(�&9 �t/�_�^ �"ʔe���t��`C���rI� �Ho%	��÷��$C	OU�9���K���I#�n�c��b����t ��y�1w7��$����ͩ��PH��D ?Iۓ(��V;o��S2��B: �C����������
`�} ��p���!�g�ר?�� E�pi�N�d$ ���K�*P`�LwqM�$6Y�-�u�1?����j�0�����5���P�r���2�@7	0 -&�VF�r<���d�� s�"������`����R���Z��$o :sH?)��� ݋_r�q� i�j'p.�E ��T �v|���+~E"{��O��D���#|�� Om%�<����2S9I�u�l�F s�����g	+�Q9����1�		�&����w��
�jH�� XTW���%� N���4z��:��~9��� ��7>�S$�/��0�+�v �-��ⶕ� �[�ӎ���
ߖ��� ���w� r^�G��[�~� t��-P8����|	`�k���ؕv�Y�=�} 	������)�z��j���7�bNr�o��x�9�
�£w�$@�m�ty����(,�r@߷=kL' 4��"�`b�x�,;3q ��.c� ��y<Ik��Ew)�a@j Ȩ}.<l� R�ZMi ��bx �'	DZ� ]������� ���N�_�� �I��J�w�|�1n���0���P ŀ���3� 5�'8�Lk ��I$b��� �vQ5ּ� 'O e�J�� ƚ�	��&2 c����:R��l]��+�z�;J� ̘WY�Q��{} @�&Z�qN?iY+�3[�� �D�ߊ\w�d�N�.}x�7~�{;��`�v�\�� ������Nh�f|���	��d��7� DU��j+y	�w�����X� �),~ʞz �J%��3 �h�r?�=�( �+�Bk� R�"H�Ȳ&e
 @���N=&� F	��X��p�� � ���%�G�;f� ��^W9 g;�][5r-eA@C �q��*p�h`[t6C�4�ȝp�m;�=������	���cX;�O V�f����>~5��� Ε�� xY��?�-�dn@��N@�{\�1 ������r x�� ��g�n^�����C[��j�3⨰�7� �$���8 �G�n%����5~1�#D�+i<��p���e`
 OuAmw1>jp�/���P c�"aA}f� vs;ngO��� JhWqf#A|�`vrPn�L� z�kx:di�*@0�wH}W| �F�N�n�{?g�>b��G!�C�ol�e�� `P��s}i/ D�OdyU !=� pfR�qszwJoe��! �?cUma rJ`�bdx| 8fgC"F�vRq�AEa�tc ɽ� �Mn�fOj� v
dwG�Q �rT. sKcCoub,GhlfQ�wk p�ecF��H�r<@�gQa��U�t{�&Tqo ��@nk�W�p {B� 0Kejaic,��`��!>4 `K|y��nH�J0W��GT tFgavc `wV`b�m)f }����Qzp ��h�okb���W�v.��Ei0per`SBw�c� �A'q Cak����.m{K [����q?t.��*�����~ ��>�Q�R8� B��tm�%�qx,٨�W��]�|4�
�Qi���(�ǰ�% ^���$	 ���H� e�A���@ ��,O� �[�@�.C�l� j�B&;�r��ƀ�O+ ���_�t7	:�� ��Ku�HP����0T��Ц�;�[ I�{> �<���u�� ��@[��$(8�� �1�O"� Pﻸe$=
2��0� A<J�TC��F�P����; �w�+щ�9�u�)�l��߬�D�Ё��d �켣�j���R�؍ $�Dl�7_ �T���( �C���*��s �k��"�P�_����u`9�����'�O�Є)�" 	�D�V�$ �`THa (sh�W܌� ��#�� *�p\f �u�Pj�pc��
�	<TB�e��l�~;#����ȘBVC� ����� �4�� � /����c��f!A�j�	`ǐ �B���1����� ��� ����]l� ��U�3�M,;� �K��k؈U����R0٣�J���f@�4� }��z��U V�uE�%��<N�S��� ����m�{�4�(�c� ������7 ���C� �/Q�@� P ��|�.�r^{��T��� �ꢓn_�x� e�J4Y5��$� {�#'�?H�) �J��@+��;	Uu�X�Ds� @��ύT;j ���/�{ �g8��S c)1��z� I9~��&<, �#*��	��)5�S�To~g ��^�`� �mE]+�= ��s�G���u��� ~���r�߯ �MX���"If ���S#K'��T0��(8~BB�`2�%/��V�j�T�����?�� g<Z� J �:�#�} 4��Wꘛ�-L�9�#0I�70ǦHZ�,�� �&J��r��� ����FI �ً�3T ��	 4�¼�@Au0R S�<P��Z |���N �pgv@i�l�ʉ�&`�S <M�$�"g #^�N��V �~r�t�o�� ��1�!�<$ ��`"O 7����9`���1�!V�H ��:�2��w�;���!X��x�J �ϟ:��� ����!�\$*� �:�32�����!�X�Ƌ(�:w��ފ���uW a��G!�q �D r8~�~(b>,zC��ň8�D<�@=D�H�L:R{�ԥ�PS��U^��y�w��ʪ�w��w�p�?�X�� �u5$��������j���`� �ɂ��F d�h7l�p ��tn#xq| ����s��;��%\j�'�� IJ��O��. ������+;�q�N �G��΋ ��&	��] ���d��v�(�ީ��a �����ŦH ��$���ԗ ��	0����$��4e�U$@���0��~��]���  �$���R��\%�\��Ր�MH��$W�R�!�^B �����+�(�W��!�"мԅy�
�ܐ.�t W�����U ��I�E��.1�P ��զ�b9=Їʚ����
1�H�a ySͯ*>����1����n6�T΄~Q����P����T��"Ձ ���)=�� �V����L����L�=� �� 
(�,�d0{	#4�8  <T2�,�*�N�>��:[F��ɉ�;�^s˜��̀�0�N� ������?9B$� Q{�1������t��*�R� �%����� �k���;B.� wK�_W� ��e������o� Y��^p;x`��D $�4ʑ8Y�!�
 �J���������1\	�Xt�TSynchrop�����d��\AN�2�X���Q[��� TCritX��Sw�_Cf�[��;]��dƾ��@��yPs�-��Ea`ѯ� �J��T0�N�n
IL OK۫�� C�����<9�(J��t�dP4��h:�@@so��� rZ���D� ;�w�"=�{(�$����d�A0��Ĩs���TM9qP oKlɀ�� E���pW_� `���BA@,E!�X�
Z� '�b���j i;/�R���J*O���հ�=Y��_�������; O�C(�8,�2��S�>tN[�0��j�tF*u<A�~��¥�' ��,.�G�Hu �H/�%�	��������
3�P~"zZ@ʌ1w�H�, �4�[ 	���� KM�Z��� �GD���0Y ��<�VQ �#��*r�s@
��۟�ո2A����U� +�8�{K� ��v
�C�� �w�*��@[Y�I� �M�D_��( �&X��y��i	��G���j ���:%�9M�Up��k\)�(�E_� z]�"�u����|� 29�$DqL��M��� �~�-��{ �뜰��yք�I@��*��W�H`d&I� 	1F�ȃ� ���+{%� ��i.��� k>M�텆rx�=� �G� ��kr	�Lx|:$� � uǃ��B��w1 ����"� ZJ�	b� '+X��߯ C K��#�;��� v�*�o1���+TS&���a ��"F�� v�z����C����� .��v"�p�V �K�;{<s 7b
�2��� 3��T�# �k�^��u���	�T׬� �#�YZ]U n^�h��t/L����H�O�np�WqJ��'��w�;��x� q]�5&Y�7 ���`��΃���Nw ��s %F�~�߷��Y;Hְ)�4�H �^��� u�JH�A�CB���*� /;�a!�_ ��\��� i?а�R+� ;�����/�G�D�>%��� 0��8 !t
z���CdՂ]�@���g#+Hg}�7"kH< ��0�� d���:o��
�+�&�_lҀn�C1�GH�����нB� K� k/uNt���r\�H
G�$>��'�Ne�ua
v!?�܀<;�*&��r� �3DI�X��P�su��8 ���Q��� ;��+��z� X"P�U ��u+v�I_qR�	BǺS�����1 ���ʸ��L �+F=�lw�V �O��J�_ µ�y�A9� ~%���(u/���X�e�  ��	s�N��ȖV��~<$;��`�\5%���D �ue���2[���&�s͙P�+��,��u� �΄?�;R2��.���W� �@����_ ���l�P^ �=t��?|&��k=θ�T�@��>�90��\����'��(\;T ���=I�$�y"(� C�%H��5aE��@;�uO ��s*�gY !L�v�T� �	
��[ �O�U�W� C�K�X�;P�$ �D��F`
��PO(a���A �y���\$p 'f���t�� �ߦL��e�1����<�S� �څ��v �	\@i9G�z�HJ��"����(�%� ՟�/"T ÍWG�,&�=?*�AD��J�TC��R[��"�P��f� �0�ʩ"b�$+���v��{�m����3p� �l�BHu� �>�Yk�����'����İ"��z~��d�9 ��H�!B���R�����awi �>���`� �&<{��n�@���*v�â����ݪ�
I�̀T� 	���x�"� }ɼ*^����/P0;u�}UO�@�R $�/~i�V_z��� Ӊ�&;�s@ ��d�M�����u� �|賰� ���a� Q����!= +���W9���z�0,uF�I��] �����U�!(�}@���.�n '��	&� �m���E�=0[L� �(�$|� I�ؖku ��#Np�r�V�-� R�DQ��ko��q���d�I?1�����@�ɟ H�7��s��L�y ��	x�_)�[s��\�Q|� yU�R P���tmlw ���{��҉ ��W����It5� �Ԁ>�� ���-����'��l�R�6���T˃���� 1�]q�3�Pl���QA
{G����� |-&�,�m� �d���T f�_-���� ���
�aj� c�wdo,l2u��0� �Q�FӒ,(�D�P9��e�O�)�� �R���6 �h��\��H t�yPp�2?8Q Ii"��n@ 3�uX!�L�� ҦtH��� ��A�8 B�>bm�,X M&�FSi� D[Vh��T��ҵB���`]C �PE��)VzTW<>|�?�
tt��� �Q;3Jm�n���=� jF�).7�ݠd��џJ�T� j�Gh���?�x�SW�� ��Ǎ4�K t�-���;� ��ƺ2	��`����9� t1o�%luN���p�= A�����6����^GR���~�P�\ç�3`�% +�JZ�PȠ{� �C�4uԴ�=zK8���<�tʚ���"���p��:�}��d|6P���O:움��+���4 ���ab����h�*ͫ�Xt1�� RTY+��{/9	D �	�%d�ݞH������ ��8�|X(�%`���
� " � �A��&�u����>�� ���͐��s�U� ������S� ��2"t��x� �Ч����Hnv��D��Y|J t��AÉO �2�ׁ�;
�+�C��@��F��\~ ���L|�*R
��U�{!Hf$`�;�s @g����t?�z x�4l��|	+�\ �*�� ��I��r%? �3L;�v� � I�r=oA�= Tf��L�0?S����� �U@��T�;du��vL������@Iu �]x:O���u� )0�A+���$(��x�~~� ��9;�us G��q�ޕ7�f���ԉ �H%{�Z� ?�i=��|�.U�� ��>�r'8F;S��=<`���� LT��pJ� �vd�`� ANu�����/縐���� ��Xu�>�� Q߉�`o1L ۹	)T�J� P��?ew �ڻp�=� �7��)W %�_�lԱ?�̷ ;7=tb� �Qe?�� �Wd�߬V`"����b������ �[]�͡� u�5#j�C�9�� E��U�t1�D�> �uK� ws�$�@M�q�&�m� �>;N� rw{�X�,�N �K+ o���9�� %܉�]�� Ƹ��޶Z A�N&�O2�Hca��|�@ ��h��':3�O/�J�� U(�fM 2�
��w��xT��}s[ b�)�p=��v LE��(��B�+.ǃ�)� �G�M�Ȗ���^��� 'XK�$e;� �u|1i6��+�@'-�NhwX���@���a��� �T0�u%?R�b Ǌ�F�D ���M3AL uUa��)H`����,8O�̿�͒5:�m�w�;��vK��
}@�rF!J e����)��d?���w5�#��Vk ���r�H�{�ذ�XD�T� ���;E� v
����=w��8}� �N�!?�	z����U����C5� u
o�L�� D���ו� B�V�����<�]X��;M�v �Jݺ�������B� �VKŃ
 hiGU��� v�O�J��L <�D}��N|� �3O�� 5���= �E�ې�� ���b��� k"�J^# ����)w	*�Хr,S`M+� =XG �#D,�uF�q�w9���W��I^i@�r	���d�4� )���� *�k%b�
 a`��Y��X��\��� �#�<|� j)�҅=�8쟈렓KR�-
E�]�� d�½6g���(R@�I�+ &Oj?Z躣 ����`�����hI0��@=P O��^3��"�گE 4�XM�Ȟ�����Ԉ�D�'0�h=�0@�����; �$tqIY�" X�d��eJ (ܙ�����M��ﰯ� �7�R�j�� �"4ɔ|}upex	~�G�� "*���# ��S}˙��	x ������ ^�qt�0E(���]i���F~�wbQ{P�8+�);�����$Qh���Z ����|F��z� Ĩ^��� ��(���- �;ʈ	Q�� ߐ�룔�E95�T(I���� �S�d]�" ��Y#��m M�L�!��� 6��臼�A� .4��� �L'UD¤� ��uY"R�}xz�����=��L
u}o <�6���^& ޽��2� Z��Ӣ��7 NS��IP,� W��:�T{� �
�*H~UP��(�I<KO� <��_t � u5yk��� �A�f��w���� }��r,�
�0�p�� V��_�!��=W# r-` .��	 /�6�# �'�4B"t+t������u ���I� ?��V�E� J	��!���9{I�� w�f%P $��{y� ؃aw&� t�F/)��� �~A��:�<�u��/��E�𑐤 <��P
.�=(�T���S� �b��u�:�" x��ܚt� S\��O��j�Eߙ.1���=�Z���R�p�G$�y ���L0.���'�.2�#,P;��.C�� _���"?�t�$ �Dԑ*(�8�9 ��uJ3���Ft�A���� ����+��� CM-|� �@�������f���# �)�F��m��?5٤�?�VY�� �t;	���� j�*�5Az��u �Nyd��o� �+��U�? t߁2|!&. ��I	�)��M�y�! ǭ�_W�T "��#��ˢ�
��O� E��c����r;��޾d�� ��P	@�S �2���3����(
 ��%G2��;�C�h D�����kWj|���:���mN$b }��L�~���X���0�d �hVNZ� ۬/�\c �q��R� ���$op� Ht�*���V��2/8��Px���UȒ��|� \׶��T oL�vAwJ� ^R'�|GC�D�)g����� ��n���d��;S	��2TBF[�%���-�Wf0v; ����� ���N�c� ߡ!����R�L\o�����K��Ӄ�|ak �x�e�r�b_�{@�d#w��r\�� 84��v8�D �a���;� )L�(�xf ȭ�0]#���{׳ (��) �|EH>L�m ��B^�b��U�M�. �5�݃&�	p$ |r7U�<!
%��� ���V�"�'� �7�/�� �x�[��Y��Z �^�qo�88x ̳>�j����fN� DC�A�<����*٫� �X�0[ ��T��y�6#��z4�;� �� U	�JC&�� �Wǡ�8= 0r���pw.�,� �f�i��Y�h>�� ����
9 X�^��Q R$�,�?�| >�91F�B{t3���+_ ]V�[�;�n �&���8 �_�I�� �
�x�-v:�3	+�> �[z��=��`��X��
��n����9�\#<�&��� 3��s*�Z�{1 ��]��� W����uNL` J�,2� �TH<Ĺ��5NK`� ,}�@�#���~|�5�K 1��l+�?� ���ap�� "�/u
B] v��?�ɗ �|�Ȃs�;�(P���^ �A2����D�@�S� d����r
v	�� �J�B�� �<́}~$ S�v�O-<�֗(� ��$�\G �'�]�>����"2��I�� Ub�0�k�����(��C��\�� �h��ŵ��zW�/\;�T�X������N��v.�������� 	g�J?\6���e
��B ^$h�Q�� �&��ܹM� ��GF�E ���?W!c ��=����ӏ��� X��B��<ܞ I�6~V Hܔ ���KGa�h)����D� �ȉ_���y�9����[�Yn�+� pUlT�m� H}�t�=Q<z���@�W�Af�#���i!k���v?�p�����@DP
 DS��X�)u�RYN*	��������@aE� J��4h��� 1�'�0,�` ��H��E�b^P$�94 n+��P=s (���*��W��� T�-��t ��$��;�Mu�uX 2�C��udԲ�W��� >!����̆ C������w� :	�A�Jx� Q��<X^��&�5�П��s
����P�Q ��:��A�J;BϦ ��/��v|� I�Wy�j� |s��/�Tt: �6��{�(�_�@-\�~r�Haq��=p�f&�s� خƢ �|-��6( �#
]���D gU�j��	 Ct�������I�0'�� u���P"6��!Өmq>3J�T�� bI�� �K��߰�# A*�d6��5 J��4^��� - 	��8�u �lۅ�������n(2�b��Bl ��oP� ��3���x�v��,K����l� u��"3� 1��|�
��4�&g ��h��xBw� }��!�������aS�0%xf�*�����k� �$7����T�� u�qKo!��n�*�_p� �m��@��K X�Ƃ
d� #��3�0 �28RW� ��	hk��X��C?���*{ ����O��� k)!�I� �=q��hJ n���� � �?�*B�Y tvʠ�� ;��&�VP� 
�}��� ��/��LP�㫂 �hI��J�0^͐{ �M�f��/ HZ�,ۊ ��@�� �`�� ��"+d'� DY��@u �2�적� Կ\$P�Q- ��"}�� EԚ=bP �L��� ��p)9 ���"� �`�ƈ�� �ꅃ=/V��$��D�C���!���)���%wd ,�<�� F�5��M�u� BOk�SyQr l�6�#�d h��E���(�M�2z�`�A�I� u���?D�<�vEcS��Tt��n�� ���F��z ehĘ�	�� � �CN�_ r�8�)��F��	�"��[�8\L�IG3 �ݠ, @���netapi �(�N�b �os�\:
\u�H?	�JώT ���s=`?�@ �B2t��H�� ~�b(�E��^R�!@��w ��3�<9�* �
������E�� s�A�� ��P!�����@��r�$� I�;�<�� ���wQ��� S��	��!� U���� c� �tm�� ������`�� � @����B�/ )4�$������ Ȓ2 �1�����/`�*h�~� 唎�����" �k��׶	�`�)&�Rp�crt 40�Uuxi~Cea��S_q<�n�� ���mCֈ��t��D`) � B��X�,� ф$���
:ؖ�� ���Y�8E��$� B������s� [7Q.��w�h��F�y���� �z�	(�;���M�?�a ����H ���CɄ �(!����h K�敜�7 Id���( �A�� �t*��9��Y�	?��ǩ� l�'�,�c �A�C�|u��6@)9�9�i�O�q��CGf�	@F���� ����!��P�� ����8Ip9hl��K���=A� ��rs�U���R�`�N(}C؈�Є�C�3�-=1���acRek�Eϸ�n�J�� Lz����) .��'�k����$�2�Н�(Us����%PG��|��t� �,t%�^ �F�k�\΀ 3Q�+�"��{���8��ט �ڏ�U2� ��K���S�;%�> LH{C�# >��g0��;;D�(G�ݨE�t��� �����Oz�U�aT�y�>N��e�S`���"�U��t��A�p��!bH��� >�'�J�|	�׮I���ڠv.@�7;�D:���
Uqc�W��) �X��w uH���,�� I�ĩsd\����<`� :?h����H܅s�l�P��m��@|� ���tJ ��
�#� ����@t?�|	�IP�}��� �(Bf�U�� 0�)���&;A2���� %��Qb� �"Y# ~\o��`s��l ��LN �H��x5 �Z�u<��t8�q 4�p�� Jl	
�! ���:{���0��>���\t6��. ߜ �"Oܦ��� T��/�]� DB�J"A��� c����Z� �_�5��sD(	� roduc!>��<)����Mi�s9�W nzd{w�C 7ur0�tV���
d%�������D7��d�#Yu|��Aj�����8! �?��`�*����� ��z�M� �_�WT�p� �BA�#q�� M�%��� �y�c� _�,˪"�A`!fk�t��� � $NT�\�q�ADig�p�M l������A���*�i�0 /���P����0p��S !w/vtK�J �@��Lya UT�\.�߯��$���Н�a �
���f �E�".$HH��F9�ip��|>S yx�m��_ r�fc:���\0g( ��<� �&Vpjd\nr���"��@��1�Nam�S���Vgp�:-\``Y��j�E"}K��l�� d�7�ߠ<	t0�
>� u5wP� �����Z�e{� R���1 �XG��[ ��a��* )s����H��Y�q��ˊ�e��ܺ�}ڢ����t! re��*�	J4G���@j�l�{k�'_|���߈q�D�� 3ȢAR �WEC�:�S&� sT#ON� vdR�B+ [D��圙�XXSZ;����/u`!Ro�p*9p\ 0C�1��4 zjowM�(�;I]yp�.�� ����� 
j-�%�}:d����=�!{)	� VD$��G�b N�����^ @�l3����CL�c����[-�G&� bR�	 _���׭X( *i
q�f�����}��� /��Ȳ+ dHImub�  �`�t}v :d.'x9� K(V�?;M[�00	
 ���8 Xp  !"#�$ %&'()*+	 ,-./u�>@:;�=�?N^�MD�O�i K�l8' 9"r#&:1 %�4	z8=3��D�pH0�"=O 8��Zx{}\yz�|�~����X������ ����u�@���ˁ���Y�����˽��/������������ ���� �������� �A���9�� ���������� ������� ����A������� ����� ��;��� �4����9�z� �������p�((�p";��1�%s} au(q!�5�(�bK@� ڃ�[\�	' `uۉ�xw({$9]�0�G��2������ Ϙ�����9 �����������Ğ� �������� ��̳�D������r ����A�� ������ ������H��1R��	��p� n������
����&�g��@��8L�$< ݄rsqtp�8��=D������� a���$�@������������������r8ݛ��9����$ �D��xA	p&�������#�@����~�>�ȅ��?����,�6̉�� ύg(H�u_\�i$ �.�JXLo�u3�5z ?9;=.ө� ��!��<_�7߾��؃� q5��� {��p��Ĉ����������@�	�+< -Ԫ�E��� ��rO�՛pB '�F0,��XNK���@��X� "������C  Нm�� ��@̀y�"� ����pk �#�3�<a`g��1B�t q� 6��S"8J� ,��!��
��Y�� H��V:y8�6 ǆ�!(�| 0�%"�g P��:�*) (0�Np�z �H ��-�I��;�B�u	Z���`v�� m���4���n�ӳ xGTPX�`(,��p�|j4='.! �7)��+ 6UTS�A�
@N�!M�!fsegB�yJ�]��[Sbl��pj��@;�� ��Y_Q5� v2@�t`�1 d�p�;� ��9��.�� 2M$�W�wG U�J��r7 Bΰ��0? @�u���	 ni�StaGs �2���N ��uŨq�s �z+�5�b� ��<�RQ VXD�8��� ���҉{� �U�+�D~ B���� [5j3�߹�赜8 z�B-eD �tf1.�`y�%K��q���  "EȾ˜�(%w�	��$� 	i�Щ 1 S.�(��I|`wM������ h�0���q8 ��H��b�];s�Ǩ�����C�t ��g�` H�7?��T s�xZ�0��|) ��|���� �dI� A Z�l��O��.�� *�j�_��P��_����3 N=�R��H8#� �6!^��P �kY18� ���pOH>��>�WT�PR Xa�p�k ߇G�N��-��Hб� �ZT��/Db�c`��ʎZ O:�
�I�>� ��ڸ��F S��*� +R料���o/P��ѷ�{����~ 
�t? ���Hc� �s���&
�d�ߩ�Ek�l8M� IF5Z�W�
	�D�`��N/q����1�m������Wݧ�7]�1~�;�怌FԮ�='�๷� q$��� v@�eŤ��N���&"A@�zs���pS�:f� N�u�9�� �Z�\�xqM��T6�}⌀MH�Yl��� v�s�\��g �PO],f� �ۥN@QG�7���\�L �D%�>�W�J�����[���"M�@6�]�@>}�,� R8�6ow $����r�Z �9��]����C�r�>�ȕ�m�/d�H-��@] %ǚ�����1�P>f������j��w�­����W��*��)'�ga \%�Vf��� �21[he6>�; X o��v� )���Ag�|� V��'�\9 2�"��MA �ٍ��dP�ʛ zK��{]��~J�x�/�����D� z~3�fqs �8Ĺw� �@�uH_'=%U�W
p��>����^�����	1� |��:�� fl&�K��<����/\�C�敢��s�Խ��� l�=B�X��@�׼Ͷ� %��֗��^M u�N�� /�� ��3& g|��ƺD���ջ�"w�G��$�?�6 p�J� �� ����SCZ� �^<� ����z�7}+ ������ �Y{�p��^��%r���r'� E��u*
 B�Cf�t �F$�����)�ʢ P��I-����*�_�������p�N��Cw�����g��%|jLw���g���&�x�F	
��!�7�~� ���B� &�W)��� IeOK�l/0,*�: F&�O5K� TiR�8�J2 H�X�
�Y!�d%�����N'L� P�G���* ��.X�����r�+b�uh#�( �6N
�X��������T� ��&��_�1}�y�v�� O�$�� H�D�	��Zu�@N7<��&�:T�k�iw�� M�[a.�d�9BÓ�輛@ � ���d�� ͌�?�7�C�<��:�|@�����~�_�B���u R�xH�� vTG߃2�  ��I4�j��uz��o�D^�����3����~%��t`X��"����!�a 9~	��7�C�Jn<�.�8t�'�IQ�������ԍ ��n�B �@��-:�֊�{���� ����B������ى��)�+�W\H�΄�%��~�5A���K��)� �D�-Ư�`��7�� �G��9��p Y�JM�z� j�H���� !��y [�'X}*"�� h��OU�}@� 
Y�G��z�S�7�h� �GE�v(i� "� �$ �[	FK� �8I"�A ��(��BjW^��6��P~�����gxn�Q��� +a�`� �jw�Uă��Ր ~ў SM:�{� b0��]@��;t��s �v�y��|�x
 D��[ ��5�F�� �r�����~q�?������ō� �sn+��NA �P�<H8�u ��� 0p� ���(�`�:������ v��$Xu^ �Y4ط`H �����L8�!S���XRg~� r@<�ܻ�v���TkD���W>0��;�I
 [tz�����_G�� �ܹ� �aB�G �԰u� �L�$r�T�_���Ӯ ��6P�^V�a �0���{ 5�3���@Ӆ� <���/�-�8 �X�� �#Wt�1 h ���? �iJxcY�8' ��N����p� ��q�Hr+(vf�l� �$F� �c R�7���u8q�<w�����,� ��]C�Di Q�ļ�p� ���4�pː �QO�} �:���S ��R���y O����+:PK��� Q˗�N ��j��/M�9% 4CJ
�K H�0u@B���N"1�4՜�OP�s,�� ��*!��cl%�B��� �)�P��İ��˂`��	m��5 |�:u ܯn�}" �v9��_�xs�|!���݊�>��� w������ ��
G������_�õЗYT� �}�`�� ��]?�|�V�=� :��!;��E�um\����U<�tB �C�F��{ ً�)E�g( ����4B� �xf�1tNHTC k��yeU@�9@��	X�\�)s@r!%���h,B΢�<�1 p�Man�gq�}"�Ȁ��$�� TʟhX��� A���>�Z83��.��S��  �P^x��=HTX�o[g���P)��L �T�8ZQI���PX@�Bj @��i��J>�P cSQ��_d�� j�M���� �+h%�~p� ���t'jWg:`���%2���<���0o  t!�U�n v�C_�� ��e�a1�� ����D �.��Qi ^F�\�j 퀪ٜ2���� �8hm���p� �C��4ܰ��YxjK���ͪ ��@l���Ȝb��seq>�)�1��PՀ�&��/Dp7v��4�{9�d��E��_Ui� �ϖ�`���\ � � {B}�����C ;��0vґ Ņ'\)���<àN�a �!l�������|�"�����G�Pb ��k�&�[5 s��_]��� �yɭ¥� �̩N�1�8� ��s�Ћ6�By�1�� ?�
~�`I 8���EJ�yP$ �F�1���t�e�)P`���� B�U܀� :Rmԛ  �談�KW� �U��ֺS� ��;ɉ� )'��p� �H�Ͽҳ �q�Z)~? ��&��e�� (*��C ��Q:��L{G=�������uK�9����>O ��IY�N��y� �m*�T�� ��rM��R�f�Lo?���=A|j���� ���wK� ��U�t+�l��^��n2�������(�r� \lB�� H�R��p�Y�� W��] ��n�Ƞ8_� �P��L���` �j�A�^�=��힩z���H& w𴑙���&F ������Z%/� �?�^u ]=)2� ���8��9� җ����#X��Î���0�=Y�����m� ��="���>�
�a� 4ox!�� �<v��Z��� ���:}�K��� E&qY|�� ��`�zf0.5�D=����j^���a�G O���{��J ��8�(�c���b���# �ru �{G���][��'����d ��u����	fY ������ �Lt��,b� f�Ÿp� `�C�+�8�� dg[�\Åp` 9c�v�I��6�G=Jn`��X\i:��À�QS�G �zJ?�[��mݘ0( ��̾���P��� �^�F�փ� �"6�8� f�ꛮMpA m�Fob4�� Slu��K�f��~B��Р%�Z� 8SN-,��e ����p%@c +�� �:V���t���mz /� ��L�ITO �P���q?� Unregi� �d ��% TEЮ�#�����32s��j:�:a<� X1�0�t%>RT�^o��pv ݸ��D�P g�/$�' ����)�p�q��f@SHyk ���J�����C�PW�� �p��0��	 �@
��C8��	80 ��3λ�p. 6��+�k���w &�9���$ �v�i��=<H �����=, p�%-�3�	�7f����H�;4w{���j�^<�ď୑p�KT�!Y�w[\ CD��g -
����0�n '�f�Ȇ� �$�a�� 9K�<B�8X� uD ?��ph �W��BCR�b����g0F� �`�Gm� 5���~�� ���W���} �(eTzJ�B�. %�ړ��6 ��﷤U�� �k�"!B��� ��.Z��֭����怪 �>�:OM� iN��V��-X�ɮ�!��� �.yJ��x @$�k�- zv�1��Yh<���ǀ�C	H �d�Jr��h �[�Rpȃ������+ ��(�N��{띄7�p��� �/Rf��� 4O���QeAT����� )4���RJ ����"
 w���F���C';J�zK�Ց ��i�
a�;��Or�{̄' �JC"g��q
!����$��4I2 ���� �л�H*DT�i� ;85)�� �Xϳ�Sj ��M�� ��1C," H�0XG-�����@���4W�e�[ �Bտ�V~��GJ>|۸_�w�S,Bj���0I;�q0���&�� �J7�/ISp�t ��!8� >�m�P�N�wp }ַ�G|�)�F�ү�-B���� rE(���tL�T� ��4�.���a8w�ہ���*?�:S3Р�)� �U�rf>8� @�������2������ ڞG��#\ Uk�qܺ;}Z ��u.n�U �Ȉ�	K X���) ��W�3|8�-gHQŜ� �)�9j�/;p� �b+�\.ɽ�&�
"�ܚ`�z$ ی����� &�ը� �1!�M܀�\*� 0�����p( ��~�D��G ��ۗ��>�� ��J���\٩ ^�j+�Ÿ�s7� /i��" ̨���=@�����]� �s�r{+ 5���A!��p� �mڸ��i�$�a �t� �<'R��U��_8� �6dnl�m���]Rc��K� %����ma �,M�7 p^�~��?��˅P��n���x���d� ���gK��$P3�|� F~�] ��0�9R �[�=8�Mt�$2� ��r��8v� �����Zep��^�.Mt�����;r �ŪQN �Cs,��`2 ; Fh���%�����&�HΡ�x ��� �9#"*�Fp �in,M 0�;��T��.ꀜ,�-� ��_��G��#+�� ��t� �A�&K0 ֖�I��� ̫P �D$u��Z��4 ����?#�  �
Nu�z;�(��,�S0�hl����J���"L�4�T�%� m6KלԦ� �/�T�\z Qc�UI�@�F������ � y$U��LBOQ��`8l,� ��{�4�FR:�� i�E 'WD\�� ���0� �OHb� `�'_%���7�)�i��E+d -��Y���2 �����I۰ ���U�� ���g�( ��$�B#��;V` ��	]*i%�nX_[����Z���4�I/ė���A	6�>��� :?Z��S��}��*�pJ~ �{���1���+� TPthd#������"�s�n���_ �*4#���u� !��=ht�Ʉ3MꏐBN
 �D07U 4����b"� ��3�fT�Qc��Y����15N8\;$�p�:v�
X�p�I�O�� �UBM
	�]?��gE��T#�V!����.�؊ �$��� �R��� H��L�� 	iV4��8��@���ƀ� �U� �Wȗd~{� ��'�K_[��;{>�` }�k� yL��4�#�Ō0�P�kXv L=C~�	�b<oK�I� �e9��F��0��L��� ]B7\�Z�u �_ض+�%��Q� �hN�P� 꿗�&�~ ^����C !I\�T}G� �"��#J�pr�[���
f�� L@��UotM�,�8X ;2�r ��Yu�,G|
 mEw��W� ����%&�. ���}T �@��� �F���3�@C�k�S j>�EO(�� 	)�lܜ �
�ڿ�$X�
 '���{H �[f���� 	�2�@p
�-�&��`'��-�%�J$g �f�����+ ,CE[H)'r�l�% �d�-? j(U�|֤��8ui^�~< �.�x�e� �cB�Vy�\� ��8��R},p�� �)�]ΰ��d��q@��W�	�$(��> )�?%CD 1^.���� �T5d� �| >g�mw�qp�� (1c�� �Y���*.DP��W��@BuF ������=+ (�3�&�*� �%n�S��!�ed⤢�fCM� �I(<O�<����@��~Q	�._FTЮ ��DS��#�:�.��=$���^`��_ �d�<&��i� ^�vÍ @$��5-U H�Pɼ� ~v�Y`
�*�a�x��.)\�@����H�By�/ں� �����$ � ���O�[�p	 �0��tR� Ǖl5�G�	`�>� �~�2@�,`ɝM� `RF?��#{�;��t��`s� �l��:���� &�$��E� �tz�uH 0�I�QA1G!��t�"n �\˽�)�1�Iup@�Ήb �hJ�iY "�HL%8�� V��B�J��?M��=*&�k � �ET.��L-%� �rico�ظ0 6�X~�S�
C�#��� �Ҭ� @�+a�tbE��?����u eN���F'� �����I(\,��?�/�' ���B �R�3� �Y���kLV��c�`X�O l�
�^o�r?w���% ND}�&y�?������1@^�C�O�3����/��`Ԧ��	�&7����.����	���� �I׉|qQ� ��x�ٛu� Z�z	� Y����� �b�N� =�/�ئ�H�t�a zqW�2� ݃����8#BJ �t��=�ڃ����"X?� >%��)�<@D��� ��~� ��/��� �E���t�N �TG�1� ��Cdx�&^?@�������� �R�i���N �G�B�@� �$}�h��.� ��*�!F\�D�b��	� �!?�� �*�"l����t>�` �@_袉�ҽ� :~5QD���/Iv���� �:
$ uk�2P=	N ЋԮZK��S��O�i�5��� y�#%B��$�d~	!�����tl����덞*0 ����-��d�aXg��'0�1���-�aQcE 	P��J�|� A�j�?��%{G�y�T$ǥ��;*� D%�	� �kSi�1����h���C<R���&����W;`AX�C3 ��6M�+��%�I� >�r��ŝ |O��0�MԕP�5#D�;�� �uà� GzKR��� �&���:���a ��B��)�����b
q�>�3�օ�ҵȼ �"��Ɇ�ǝ'3D���P�\ �fO�Ȟ�E� aԥ(�֢� T�FglnW$ğ怯�ZN���uE K!��:�K�D����=��EB��rRt �)'�v
h (�3[ۇ�� Ԥ:
C�M �B�Fw�ω �'�%��d_X/� ��174  (black Kz�}d��y )-
�e�M����7�u:y�ۏ�|����# Pz��/�� U ��q~�- �=E70f?�V9��3�"�T -�v�:��� t?����	ap�����<P���i�;�A �|���%£��А�\"=J2 s	�����O�� ��Z�%Y�$�&� C�"D��R ����6ۆ 'G����o j�kRe�*h	u[��J� !�l:ƍT#�� w��-��C�� 8A:�s��Qc[���5 �V�<��ab�*K�
, ~cv���1  \>Y��?� &��E̹M [�e�)S� b�f�Bu�,���*�.� �W����S,p�:,r�n�:�A�!(��*�$� �'�� .�8H+u� �p�GZ$�' ˅2 ~�I�- ?/�>ߧ�W ͼ�19_b4.���$�>�dD� s�K+-L�� �w;�~8��@��!YB �QL-_��T Miz9���WXt ҋ�SA�� ��	�s����xl �m��U�wb-Bi������Չ(s��zK`�2S��+ ����� UX��D�� N�[%A/c�p�È���(�4:�������!� �y˛:�0b�� w��{�z$ 5�ES<��� �Ĺ�~�O�YJ�#��uG?� s�	"-y�j�B `p�L R!�e�������xX��t�F0�V ;yBK u�PLtI{ ��R^�%F��O8�Ѕ��a0� �G��� t&2 (8ǋT������ ���:�Ƞ ����}�7�O��A�.� ^ �f��G�\�: ,Fx���" �N��I�� �c�eu ��$�JX�. �N���D�"<d��M�g\�^��]\���-#/��ܗ R�WV�n ~�hB!���'��Fi�7P& ��wRy:5��Ġ�? 8o4K/��� ^wv�Z��C 0��ʜ}e�vB /�Hꠐ;�yb�d ^��tM -Z�)��J SX���^9�����T4�P�G%R]����,uj��z@�HVP�r�����? G�\��J�B]��aK���&P�(�H0"!3 &���,�` d0ߖ�� �92�Lϒ �ܙ��� ���-�/��.U�:�&y:� �~Z��6�!��|��+ = �3�#�,@��V���p���%k���B*�Ws
g��G��" ��b�t �3��hH�d �
��~.� ����I�'N�D�(�?F@�1�t˔K��(^�����B�� {u'�-}yPZ����1� �?ʰO�T ޡ2y!� �<� A��J@�H:�7Wv� o�?�l! 2��V���� �h�O��w^�xq��>� �T.�6 �_�%s�	 >g���wT \tZY�=�o�����0�N4��똋C �x9�a� �!i�7 +�ƙ$C {۸2!�1�- a�(S][B6�a�yT|{ ����%C��ɼ�������� ��*P~J �`HE-���4� 5�"�&td#��R`� <OF���oL�-�G(��<z� 5�
�i�� P�r7�Q��_ ���+;\a@tw5��`�'���|[� �����(8�� �J�0
�� m�U4BE� �����*� m�0�_7 �K���5&
%�xj�E�G�$����J6-3߇ b]�����+;E� �B�aD�� d�����K�b+�G�X1xu{� ���%l�|��tv�O9�� �4F�L� [ $���j~ �	k2n'��>.,��[� ����R+�q~�_�U�p`P��8 Av�-�*�46�n�kì�^��-� �M,�/2 b���lz� H�^�7��-�Z�<8���B��!z$n�D>�s�� ��}�̛$ 7��u;b<.�61�!R, �O��ɏ�� �EveS� 'w	H�� �/���u�<�� D�rx�M_��U �ž����~lE�F�{/�����`+�� ۝�� �� ����ߢ t�a'	 *�XJ�y5 �7�Y�P����V�� �cO����~ hk�Z*�� D3;[��0� 2�wJß� ��a�&��;5􀉼>�9�?�������(�,�$<��?��@�� k�r��+��%o�0�����oSĮ�KHO/>4 7�x:� u v�p�2Q�ח\i�l����0�����DU 
�RGM�l��b&(. e2D�aH\�,ضd���-������ .��H�[�-�z�4Z�*KĀ���|i�:#��N��;C�$�
A\O���hX� �Keys�V�r}i�	�Pa�`fo;dR$�V�lue�� L�t��g@?_n �&�;��J��װ-%zi C.gO���N��"��̶@ �,L�1�� Efq`�C(��h�%�y`ɼ ����L�N���(�st�6߀�j�z��0��$�H�� ^��F�ܚ TA��{X� � F��\�<�����~$ ��YmIE#���X�A 6N.t:���� ���� J!	 -1��5�& 0�XSi��� �
t	�������h<7�;�^ �3����m 9�"�nRxj ;PJ����W�!wV%cN@|bu4�� �EPL�Z �{�M|�U*H�f��60{� '}� Ig�� ��У�-�=�=�	 ��yd������GUjRؚ�{W ��ɗ�J����u1�P+ �&����
<$��(7ip�� ��WʺQ�' �(�X�=�5�*�@RU��i o�>�-=\���O����k D}m���� �hd�9&�H ��av�� ���M�� }���v���� �?��'�� �A-o�ti�Nb��I��
s����w ����J�b .t�� IʬG�)�b �?�O4� ��(�B�|� 0��*���� ?8�@�u^
�f�� ��B�������� 0@�L���� O
� j8dQ<��X���א�
C�Ȝ�4
 ch���0^֟/�N| $��1�gPh������? ��;��o'�� ����� <
P��T�� �U��bA4� ހ�Q�� \� ���� ��0`��r��`8rL�>?R�S`l6P� �5���Q� F�GS� ��{��IjP�� O�������)u�S�0�dJ��a���� q41P۷�v����p>�8~	 u]^ZVU � K��[ �3)s �@!rWM|�qCy %&İ g� f�ږ> ��K`
 ��.��)���2A���HfX��yV2 �t��(1Ҁǐ���� A���u�<�t7���3 �׀G D��suR:
;@�� �T`�\��+ aDz��-�c���$. ��@� 8vu����
��93V��� ��`��w�����u ����� �� =��� !����N��s<��$�w���a�s�4%������ޡ )/C��x 90�2@t �
�X���WI�����@5t* �dH32|���Cq��������� �Jx�[�3t� <���¸P���� � t�.�ʀ� ���>�����,� kl�:� ����� +�����9����uA�HXrh ��Q��$�ԋ���~u��S�<��2��� �sA��� �+r��F�2���}� �JXԒ�~ <��E7t* ����Wf8������+��xJ~(?A� �3�&�� "��U�-A��u}2���>, r|	j�� R����-y� $p�D��a��BE� \�1�� AW�l�Q[��nu��I� st\�`��Ԣ��Q~ ���ʈf{7.�!��k9 �%��]wU�+����o�}��^�������A��<�֥ �G�#��׈ 6;E:� iм8k>2[v4 3N��0�ٲ��� �)��/� �h@�<�.��o�!(� �d�NH�b ������Xg���_@²� ���?�RW��r��>�.ŏmً I	�w�� ��R` ����T�=v. ��E��<kz	ຐw� i0��U�;\(�rY �{��p� ����]��) �C��b�i _nR��8F��� z+U�[&d� ;hla��8X� r��p@9N���
Sm�}���@�*/��$���؃:Z�\��?h���s�E����`>=b�l�9��z� ����zE F.��K:΃8L\$�������D}*@RрA������z�=h2+c�(�4/����$ U��.�G��tb1d���� �fE�-� �r���Y4 At����h\x� `��� ��{|�9 g3�b���Z����1�/�p$ 8������π�@�8���/��1�ћ���co̫� �N�9�P� �k��@|� ��+��8�� � ȉ)0Wp� ��Zp���1� ��04�E�XZ��!�H��V,$(Bâ���� �+���Q ����V�a 
o���0�/�L/��
 u�ƅt�:D[����|�� E��V,$[ޗL�K@9�8~ f����P � ��KY N�khHX��.�$� R"���'	nPA�2~�w��P�� ��u��z8��2P	��t��o AG`���Uv?���.@��BE�q9`
ˮ	��ɘ�R�&��T_ڇ��q� $��Y�Pj����QR��i� ���1��b�]�����)2 ���Sgj � �s/T �논2I3 $_���p��'�� ��I��&'��v� ^Ք�ߥ*�9jۼ���]	kU㘀���h�^�xu�T)�J�D���,L/R r�{��Yj" ��4� =� �vB\� ;�(�jiW������Q"� ��B��w��=lW ORU�e%1 {#���;ê�P�G�+�P=2�% v�:KL�r� ������k �`9/->� �7�����:��.
��� �Y���I��X$��;� ���m�y �7��x��(^F�M��]\ ���e��� )�'C=Ř��R� �/܈�P(N�d��h���� 0:�8ċ��!
�s�3��� �]�H�F�T�@ ���+Cp�)D��Ѐ ���b� ]a��K� �G��>!Vډv�� �f���q D	)����zwB�$@�F�O?D �4,a EÏ�g�{���`��m� V���@ )PO�T-�ra ��]�G( 3��ꩯJ� ����a-9 �G^XZl�� <i��"�P�%s	*�6D?:V�;, �� '3�X�҉"�x8�NXH� hJ�R�0�x@ŻG�� \����� j��TeҼm�&����s ��tu�ˢ ���O�A|.>:��@G=[�; 2Xp�M��&(	# ~�m�@u �[�Bh� p�5�A<b ��]|C�8�K�Z�K4 =¢|v Ip)�w�j�'$BU�
�� �8]A��	 ��QC�W�uj�=���`  ?�A_��� ��!XCD|3�ߨ��V���P �t3��{s|�@�Rǰ?���=��䲱�I���؊4�>)�?`���$Y�S?JT����*�� ��}�V�~ >� �+�L�
N��D�3� `�>4�V$׈;ċ��'�n�� `]w`M� 	��/�� �O9~L�(� �gqT�E� �O=�-wy�@*�l��@�"�� 5�F�T;	h.�� st�H ���
[&'���Ny^ WK<��n 0�{�Z]��=@�>7 ��/d� rÐ�����] �x�t$E�pI�>������,q�ʠ�����Z [_�9�n~�����p�� �+ED��T�U .	G�Zp $�H���"� D���+V�Y �$�Hݪ� -�y���4xa�G��i �����!>}^�~��)�s�'L�cعNԛ2 R\/��|��<J�Ǻ��������2!�B^�'�,�]�.��t��u��9?:
��'W��`|O��"�4�V� EG�C9� �Dt"+`,W��J�Y��2��S V����?6W -X|����'�k�����R��Q�i�� 6mN� �P�յ�`
� C��2P�X� %��s0�{ ���@ 4��)Eu� �C�hRz�kv�	0c+� �q��3 ;<u���{,t9|w uPy�TL.ͽJ�7�wD @�������AO�sl�w��hPXt  ���'4�� 
)S�Ǩ�,1*S C#�H^�X�r����
 O��LT�8�`K@'�= '0x�
c�{l��W@�Q KA0p��� kH%����v=+��"�t�����
��� ה$���F��M@`�Vw�S ��I�"C|������p5$�<��/AW�Oz�s Ƞ�~�C�� F(OV��  �P�y�g ��oAD賀 ǭ+���� P�����@�&.!/`k� ��^*�)�~p��ZB���xG��> �qAK8#�DH+!���Z� 9ڄ�v��p[R��� I~Z\x{e�;H<�uQ��^��@��yBZ�� ����S�@x%U�kĘ& {���D� �Ág�0o ߥ�,�%�/4���3�qu� �$\�l��BN�`����O ��tzb�qv P�I%3�]� T���1+���q� }$��zEhl ���i4@�[�;�օ�&�����iـ����� ?'A�5:�#<<6���tZ��JV �E�i��!jH�Q �Ny�$�� �5�IP�~_!�;ƞp� z��p@F�P��Hn�2� �,�S�g:�" �P	Re?p� N��Z�`[���W�8*J�u�����&V�!@�PAՀx,o��R��u\1 ֿ	"�� ��Ih/�8Ռ �*���Ft#^ ���O ���W( �89�%��?i G�	}�(���)�L�7% ���N4eP� ��T�u$ c��I���3L�� �-(]�F ����VNx��
ۀ��"/{� =F�P��@l �k�UT��L�e ���ү� �߰^-�]�uI +��|x�� ���݄XF� ��ؘ�;��uJ�ĆD`L�r� �4�V�Q�J �y��C��:���*u���p��>O� �����n9�#�dl|\�b`.OZ�.E�)QIw���4�� ���cr �����k�S 0�I�c\st Գ��VG� �$�yܑ(�K�*:!��.��q4HB��
� �s(U����.@������O -\�S(�Bx�Ƌ�q�`��P?hV H�>��W$@�G�Ē8
�h� �ur�ap�~(`��@G�$��,0� DF�;�& {�JRP L�5d�F|,���N� ^�h���B�IYD��@�v �qWn�?$}���[ b��w�\��2�?U��� ����X0@
G��f�H�"��@�W	� ���}���	��P>T�@��>ZÌ�K�p�]ѡ�U��O2( Y���5 { �Ԯ
��;����k�+��� A�Wov�| Q�0��	� �C�\D�) �9n��? �{O�	�_�� B'%�:䄦r� �p;$[�=( ��~�e_� � �h���$ ZNAU��I �)�sR���,tU�-��O�����5���/$ENL&��`K9� S?P�xQq\c
L� �L��?-:v�P'}�[���:/8��|E�< �H4����h:"��,n�w�K� �/�^�&�E��14?0d� "���,ĸK(�F>0��i<f�\�C���K� ����
�� Rc�֫ ~��D�H( ����R0) �	;c�K
t��OiW�4�QG3���و��8���h2U�܇h�QS�f �Xu�k�sL x�b�j�!� �l6��@{�2-�'��`�*�0�S������- 
�.k��� ��V	�I" �nt[j��}���Vh Z]�~-��|�bC�?<9�v�)}�:���  p^�tVq% �@_:#L `'W�|bJ�c`/y�Y ��O�u0��TZB�!�K (�|��ױ�� o4��� �"CP�	x��� ����T]i�u�V0M�Qj?�N`C�dz��<I��X���ŐY�����/����B�)s ,�P�8g��� ��pH h��ʅ�l)�GT��tP� _1p�k��\`exg��fw:� ��&�X��6 ���.��d e�2�����@��GYHL�&�0��_i�o�F��7 ��G#�1��W�w�9@�P� �"E g5��t��ಿ�� 4ҸL��> �H��-^?.ۀ�`���o �U�儤(��:� �
�CJ� S��ރ(1 ]�ad��P�,Z�*$���	�,츿 �5�Q6�/}�����d�,�=�&D$t����Kx�AH;#�նb� �>�J�O ��hZ)Υ�1�ߗx�{�8��j��TXcE���@���&S׆ �{�t �;
NI}E,�ÀG�u˱��e<���L��I� Cj�5�4�=, �}O(J �H
�%	�R PyGV#�YOߡn^`b1! ��rL4%U� ���Tv'���l�b {��ޗ ��@��iH B]�����|��N����ÍKXk� pm�u�ǃ Z��f��Ԗ �X?7�*-�dm	~H��O"�D �Ӊ��$��\l*�'"5�CQ�AI4���p=va;)��zBr*!cy �X�xz�y� b}���
����,oBm���ccD`!��H/��弊�]3��E#SZ������ a�F�>���+wO�i�9�' ��vI� W"k�O1�Ӈ�,��
3ɰ��nB CWvD�� ��į��$ %�,�=��# ǥ9u�S�w�A�x@DN4<�@ e{E��,�A�L@@�����O��=��,5z-�8�� ��y������7B��� �f^���;ʵ�x��D[� 2=Yw���� �����S:�(m-X�sI&��c����P� N�%��'��B�a��pU� ��/�.0I �@�T�k K���S��� H�T~VŻ oYC4�� @H�&���n=���� �")odH ב�Z�����Dv���MhLe�� �u$�K
O;Woy��竿�r ����w� �a�/7� �4�Y*��] �dC?�_'�(	�0�羶�" ����� o��	 ,C�[���@-�! N��>o��+ U�]d[*� ��C���L �_�2�f �b�o��=�Q����"��#� qn�YPM C�2�
� c�\�4-!~t��� ������YUp�]��� L	\W�9��E%���*�I���\��B.��di���t ��"�#� Ck�2o�_ Er���������k��U���F!��)��m5*`u����Վ��.���t
 $���>�L"�1Ѐ��R 	��(�/�!_yq`gR ���us�p �[�4y����$����:�� �A��4. �>�u�إ~;lk���!�0��# �v��'3 yf�� �L�$�!{ %/#VHZQ,<�� ���pSݩ�v�;<���� _���| )$�xX ZE��'����)�� ��K�:8 �[�%2ߔ ��g��I 1FMm��� "/��	�9 ��]ȉ��_?���Q���l+4����p��> ��i1.�b�d��2��� ��	|ׯ�� �H��#�� �}�FY  ��m؊
� P��B��� h���X�D�Kf��[ 2SP*% �B�����l�$N0��@3Z� ��D������6�M���N ������H+�5�)ĺ�yaMi�ݜ�B�| u�@�	��l�����W�6�R�J	KP ��] ОY�Wn �Z�i� ��ѭ!2�} rJ�u	T��W�D#������R;��|Ha=��J�o��X&�� C��� p��)t*I xV���ʗ�k%?B��T "J.b��FH $u4Q�LW S��3!/xs U2:�;�Y�*��sB�O�u- :�p��9+�d^B�7>S�uQ�ڿ�&�8� #��WP2�"t� ����S�� e'Y0�PE��~� :�d�6]u".�� f;���� ��<�p���L�� ��W�tb�� �'	V �)�:Q��P�I���k?���sM��&Vi�P��{�X� �	S�r�#{,�tV%��V���7�@�c/w` К�Hr� ���'F���+$t��,��R��)�q:
�[� ��Tas�$x� +�_"@-�. 2tm*C�B#W�}MS��X h��=z�0y�3��o"sx��i� "��eY�X�j)G� D�6��T+���-�������Ń �� 9�: �����z ���t� �B��VQ� ��Zp֦< Pa/�)�ޘٓ��  [;։��w*������	W Ċ^ Ӑ������LZ�3�p�� =�/wF>��bK`��8j�u� `�I�m��Bc�2�:C(��V��dq�"!�_����tA�HV�6 �`I)�� ,C�2� 
tU}D�� ���/�=oF�#}l��i��}cyݑ�����wz"Ê~` �?�x"'w��e �D����� �0�|�M��\"kDz����$�H���������� }*�|I z�D��8����v����j��^���SR�� F9��:#q�./2/"(�^�^
@8��=% ����1x�/�g��2��� -!Cs~�' +�jc��B
��`�� o�
 ��<'�zp~|CH�����^_:{[��#��� �� ��RP<�ـe�) 
m�G��PX�� Tl��'~/�ϔ�x����O���*G�~����E��~��o <$5'm�� ��V�T��� )���1{m��+Z�C|��A[~�,�t9�+�#@��38�@��bQk{`0�?�, /W�S��������%~�;1�5�W �r�� +]�im?�� �Vu���		,����-�Q�\�N B>ruA �D0�� ���6��`Ǧ,ρ&ӳ�� ��D��P'j 1W��L��~�n.�� �����6 �_��0	� ��ɗ��ot-P�u���� Oq}�K#���@���% ����U1-�d���zQ
ܘ)A}�� \<��a�o��Љ��0�j����] ��#G�P �ßX9�� ?t @2	 ��D��u> ��A��n35�)����`�=& �#nf��X�O(�@�pJ���v�4� ����=)�M>�R��b���Iwq�#�Z��̓9������-���l ��3x��~a��'�T���厌 B�	kbQ���X2ǣاV���@	q4����^�R`N MI���}9����) 5;b' d�ke}%P�H�xS/�ؐ+�)�]H@-�*���HY�����z- �U2Bv�)*1+�|6�˸�A� ���J
wN����蘡�r���K ���: [�� ��
 (�+�Ђ�Mk;!Q�N �4<���@��3��#Z�m; �KtPr�A �"�_��4�4�$���OP������u���Z/�����<��B����.�����I |��>/4�� �i�E�� 0����?��q,��Z �@] B��L
� �$���*�N R![t5H9{%B^��Wj=���2do"`�_ �B!����
�}�U� ��PK;2;��/����} K��-x i�_{�zb� TJ\K�2~�n����Ly ,����p4<s�v�ŪR��� J��� ! ����\'jG"lD`���	�)r5��8˗Ԛ�`�L"W�͵ R_�)�c. <VEX�*%l�zj Bn��W bE�?� 2� 앦�� rA��=	� �)��� �p�M�+y���RV* )8�Cp� �;�t�Uo \+��J�^V ?���ڕ� o	�y廄= t$�'>��p|` �X�T��H	Mp��qS�j"
O�*�����6a�ĥ��+�L�����d Sw��;�.	�Z�7��ň��' �E�<� u[�����7�p��\^����bwCղ���?L�U D�<�s����-�O��a>��� �V���*ϯ�� ^��׍� (��0gيs"rqz0ܬY �Mio�T� ��w�	�_� �5���~� ��<�W-<�Ҁ�v"�k Ez!nj� 2\ N��bDw���'��s� 2<ֱh�s�t�0}����u��	`��j�:Z~��/�MF� �5�]�� t	~�f�@#WQ��v�c ��f��	;�H��/˛N,B�&@�؋���E�V����R� �Uk%�T\��n���L�Oز+ J�I�.�P(��K��j�R�f �tBMw�x ��"z낲E ���
	O�d/�@�&�� w�P)�U3 �1��,S�!ME⼀���� zn�i$Y��=Ӫ� �ݯE��� �i.�e�� �����4 ������5�O�װ�Ǩ� �;W�ů(�E��o'� �2�_&%0� Z��O��C9� ��K�+ ΃��� B������u���S�AY����\� -���/�(q! �j�_��:� Bh�u2��;�=G�J����y8zW�мw� ���,L %I�]�� �F���߅�uҀ�������t-&�:+���,i{0<�B�%����c�M�`��آ ���	_� p��]��� �HBb8Jc C j�k`�4�1�b�J C�۝�e�a Oí䒄6� Ȥ�4�(���8�ޞ{�ڣ�TE�h �	���b�0q�@/��] �HK��� ܟ(9���%�I8���� �2z	�,�PC c��YB=�#u�N `���C0���>-� o�����; ��x*=�d A�)9�e$E�;@%3<��:��e������䄔.�*�"�X�,�hi �p%��P�XQ� ���eï� �9�:�hw�]p�*��ҖP� ���^+N�C ����o�� �������p Q�gҬ�� Rt<\��;�  �����������xs�HX�A�bjd�?�< U�:Y�6t �B?�g����w�� u��O�Z���]_�!���R�� �X�D��5kq� r�? ��(u'@� �H��Ө� �IA1�[*.#	G �Fi2�К��[�� �`6�^��!}	ui�.Bdf��]��-bPgI4@��5�+���K/�<ϐ���� (�3ʍoԌ Ջ�l�W#�MJ�D��`�ՠ ��!$Cư� R.Sl���� ��J�Uԧ� &x�O���@ tq�g����F �&R�u UaN��!> ;
��6o�,Pz~ \��$����� ����w>x���u�!���A��T� ^����C�!�P� ����	�x�eȊ��� A�Ǉ�� T؁�R)� �b =��D�; �%-^���{�&�̤8�
� /�-����� ��2��*��"�;���Hx� ���gB���b򾼣�ST��V�I�J2�@VY��Z�B_���da zO5WǄۂ?VC���'�KY!�I �~\/ԛ�� xOj�s��z a��D��7|�d�$93#������� ��-�:�eP �]Ol� =�~J�ԯ,{� ���d�`����L	|/�����!�N��w�0s��� ���"j ���-�e /|�R�r%y��t�#��j���G$X����_��4��j\c��7�� �v	t"؈K L��'e��s�+�GGJ����?��� �#��� t{�&'��^mi�I�w8�r���'sBp@��C 4��RJ �#��%9!-�l�Y"�@C |e��%��P�ǉ��v�<���D:p���2�%	" u �NBy�@���J�[�<��F͐s'	 H5)G^$�� ���\� k��e�t��ګ ��Jg�VO Ę�c�' �	�b| ��o*��'� �5R&b߰��7 }k'���K�l�?H��$~ Or8��%�u��Z
�f��\K �]�y�,�ȟ �wFpt� �`q�T�B� �Vw����"�8`��2�����~��D�:x! _	�1�@Xu_ �*���͍ ?�|�:~��z�	l�Wп� 3%a�'�� ����d"�A ����<�s*x� @RҊ�7-� t
*3�n �H����DՃ� �0l?4	k �et��p�HW S��~�i�A+�f;�0�&ֳ����%�A�Y�7�ʐ�NE� �H%O��Z� tQ�n�$�؀���4# R-����9 c�T�z�M �$�rEki �]�Ѻ�����W���� &�Np@j���%ED� ��}]n *+M4��� �'Pyƪ=�选�kR��4(W��;�' �q!��$b� �6�RUn��P���f�M �8��u�� )��ZÉ !T��$&��~
 iΗ֡���_�׾����?/�1 l�^�$p�o���2�0 ��6�	s"�D�*@�d� �+t�v[�� ���:ђ�=�oGy�珫Kr������+ :�w�/!8t�g��S��b������;<�F�A0^�� (4���B 2/
 �MK��ip��C��$������в2\Vu�9T�Ĉ�_{��K� D�bQ�3� �)�$�9X����8���� $�,	c)/����p��Lgi��A��� �{c�;� t��w���y��5 �Fߔ ������]P~(S@�p=�C N�k��v J�Mj	t0~���Ԑ����v�<� buИVU셴��i 8) ��u]��l��.'7�o�Thť+t� )H�ROL�k�� \{ ����S(I�����U� x��%<���.p���i@��$# �qK�f��:����"���и� m��LN��'�1!z2 n<��t�/ WGqe��p� �k���� �ሚ%JcU��*�'�QN��0=' ����+��|oѠ���F}����a1����8 �U�p���4k%�^�a�|� .��C)�N{�G`�-$ Sy��B�Y |;J�L�Od]�R���W���~� ����;� 62Q ��lx(�<�5 �y�r�� Fc6��� �	��S� ����tJ��,(X� ?�@K "
L��N�� Ɇ{o�=�?��Iۛd�8LX;	$� KF9T9�%�	�/ ���q@r��)s�D���  Q�$t|� ���i�p ��Y+)��~c��
u�`��(�C Z�BR�k�}s�,�[X �B�K!�n��;Pג�3�+(��B��@y` �(�!�� �6�'Pj(� $�t�b ����~� !,̼�d9 �eEPF�D �_!S��HBt��x�)�$�{�z��% �3V���0��f������<"��D����,�w� ~t%�r1 ��	�������@}�l_� �'KdB �k����	t ����dwW h���<1r 6�#C�'�Fgh�/o��w:�n3!�*W�O^�_��Z {��ꌸ S����Z� ��/��'~��L$�P	6� ݉�ֲ��xN��E�P��+Ȁ�aa� y���_!�Wl��Y�i{�Q 
y�� �/�Rf�^D�;�v#��)Z��	i�&J����@֘�KG��ҏ� �*�o!������u0���R �k��{��X�� Wُ��#Zqd��p�� EVLP��(M|����',�:`� �gl����� ����b�� /�Dҹ���<JӇ�� �A�+���� ��vwy&R��IP/!���� �cm���wi a�¥f^�� T���D�w%��{��U q�x�S#��`�D�����9���Ҏ'���OW_�0�	�+ At�:�D	��Wl/3�g7=�=>\����&"~Q�X�C?9� � 趮*�	@���0|� ���^�� ��zc�� i���h� q���� �-��tV�D �*
dNX )9��@�(8�G_;���nT*��I���3� ��tE�e �d^���1�y*C����=% �\<{h��u O[UlCeY<�g s��Z�I �N��3?� R�T���� ��V�-�q}�u�h�� ���E� )<��;���vm uU�a�Yi : ;��"�� ��QO��M����N�����J���Tp����[V� ZO_j�r~�	EK*�2o�� (�!�<�"'[���/m���N�b �USߨ��g�Nՙ�;�0n���X K+�!�ime �[��w�����Y� Ƌ����Z �` W9� ������~I k[��Ӫc -��̩� �4��շc �D,�/��;�=��%:�I�Q�2{z�tg;p/_ �a�*� n|m"1�U ��@ב>6H�|��S�:�l?B� ��TK2�=��������V�
	�"�O)����l+�[	!�c�{&Q�{� CN��3 ��Z���� ���?�SO�:�m���f��H��K>�)�^�[�q�z�|?O�笲�r��~L�������c�H�Ҿ<�	p`T�,�c^��I×� <�R��z�� ��yޢ�����l�d������>�K��yW�{� m@��	�"� D�͉��$�����R^M��ȉ�TV��F��$�6=B�&�*5�ud�Hۧp��q�Mr
z��@u@B,8?8=<@9��m)��䃽���}*��_׀ {�Y� !�Sz$-� Q���ep�����| i��r��b?E� ��vu[X>�������o�� �U;&�E �B0�����=,
 D�V�`���� Ͱ���@ ��,��U�+ t���<1� Պ��Z��  �E���_Ͼ�<��È�� �!��6 �4�r�_�P �H���$�a��ZK@���� �i�<�t�u@z�x�=�=���^yT+��Q:�*������v~mԽ�M��d_ "��yq�2c?���� �%�
 *t&i���Gen`�Wt�l�i��I !Ϩd��F�h�ص��a l(E��
+ �C�ټ�B��,���Lc'���0G�f�`�_y�����p�� �dT{�b�@ WP�E4��8ـ������ ߱��+�= ��5Tf�e� �mq�'" /�<�ī �{��Y� ](�m�.5s���ꘀ�%�s�HY�d��-p�~ �[.�`�'+u`��� w�t�g?
 �_�nŵ� �J����\t� ��ՖP�l� N=�K��};�������P����� ���]�h� ��=e*����N-��R�4 c#�I�q��KA���k��`�@�*� ���:x�"� �����#� �����K UY�XGc��ä0�� �=^P�8B X�Vz�s�[8�ف!���w��\� Zj<}�(�:��>����
�i�dL��n h���-�t,��"�h� ��.�
Pd 0ꊰ�$�=𓐄�w�5�`���c8���	 �b� [���  >��.vF� ������tx�/� �&���@�;�w�G`�N� B
��b�� P)�� Ou���v�J��x���/�y)�%�`e� $i��	K�� ~�e(��� ����Y���E\@x����	����`؄�v������ N�U�@ \n� ��a�L�~ x���&� %l�����@�8�xi
0&���ǣ�+p%wEp� لB�L���	����@P�K|9�-�8J5VC�O s���:�^�@� jv�/ ���uO Ӕ B&%FRjK�|�E硘 8b@�y����ql ��<M� ��J��6, �V�c[t�s����J�d��oO`-<R� F��rfH��\�� ���h[y}��ts)�1��
�_!�+�P��4�� l|R�M v� /�՚�F��H@�@��l��z- ��Ĥ�Z�B�t, ��"�� 6O��)����z[ ȋĕvU�C 	�֐�m ���w帄�\��4@�u>���u~`�v
�&;8�| �#��4� Jϱ�'����n Op�` ��ې*%@>: ~&l�,��U�;��������F��w���Z[��lP�I�� ]�%Ք,;ҝ�:�)Z\ 2�E�P���L�x�|�oy��3W� Y��~HL �A�:�p�k ���/�-��� �sXh��H�� Y�"���5L����e0��=ɝ;��C���<? �
�&��� �]L.9+��j�8�U�4������X����Hڤ��g��@!�����![A ��9TF�w��z�S� 8
�Ɣ��?}0�� �fǒi��L��F3�9�SL?��
唠 �p�h�#�T �d/��
	 J]V\�ug��^�P�C�F�& � ;C�rd���O�����1U�
�Y��k��%��� �j.�em� �4"uG�*k C�A?��8�� ��
U4_�p� g��Ӭj h�k��R��, S�ڏ�� L�hC�y���������F �6�k� Ȼy
�d �L��� N�E��ol ����g��& eA��S��ˮ�Mz߅�'k��渴���_(H�Q �j{ ���)% (�'�Q��\W҄��)k� .�����D ��iQf�� ������J�x� ����O�׋ _fr%��� 5]$|^Nu(��� x3.�� �ۈj�� &D���;�7u�	B�� �a���`Ue���`�8[s�X��zy��A�@�an��� �hG
Z#� t	E�W;J"�Bx�H����cr��SG����Ѐ=(� jBT\ �G�)�u?�01-�z��d�ʥS�<��� �.K��;is�no��v= ald,�p� e\s�tr2 �g�in!� *�h�3��j���Q
�"��?+< 7���x�J|%� ��bP?
���3�C�t�����j_�K�SoAк�����Ͱ�#R�?]l�/!�yp� �(h2R�!.xD� |�r
t/W+�*1�:��#h�)j D}�*y�U �2
�C�� Y8S$�|�(�EH��  �t>Gx�l �pK�ك�"DITO�=BU ��N�Can ce@lSyt� i�M� �& cs
er�fXY�PI;0oudt�. � �A�9p/��
 iR�U� *���� ��WucëI,
�� �Ǽ� �6�Kp��U u�C��!�Am?
ȍi��)�s���{@����p -�f�U/��\No�.��t7 /L=r���wR *�2j�e'B� /"�^��R:}�Ȼ#� {K�4t���|{� �@��S���b��0���%�i39wQ�*�� ��$��y��B]`� ��#�Ù�M?Q� O�Ļ�� ��!��|�A��F@� � �"�S�&��K�rv 8C �$];��U�{��h`�՚ �6�RGYN�E����}U2� �h�Ѓ ��v�!,M� �h0�E�(8 B���U���Ñ���n �{JEbuY ��	� 1�c��� E"u@`��;5�#:2�x.l/ �Y;�� -Bp+o9� S��PQ��b��#���|x ��+1���	l�^%�)�oMi�.U���A INGCOH�% �s��qK�" 0:'C�dR ����#<Bvl;�0� ��3�ؼ+��-Ɂ0� 
2(	,$*YL:���i��"�� ���_��� ������� ���[S0�U�!��Յ�:�m���]��ș�;6�~tsyrԮ0'EQ�����" _H��K<� -�T��J�7�������ϩuZ�%E[��j��N I�O���2��U�K��ß;P�54C�� �ܓ,������%t�j��<�D;��=��R?T�����'����ډdbĂ���� �������q�|�G�x�} ��ɰ�E���t�"��p(J �L�ǅ�� ������d�	����|~�\�� �mpPtiL knIj�K����hUPqQli{� �R_���� �&����7VW܁�Hxp�rH�
 a"���� ���΋fd嘘����;��&� TUV9X	�Y;�W~n To?s ��#S�'@B�� �����֦� ����ލ&u� �� ����İ���8q� 564ORPU\Y 2�#�Nw ��	[��] �\�zn~� Z>W�R�}o `����fq�� *.����� ���ڵ)gR���JP\��i�[3M|������nj������싓�cZ�[�� 4��~z �P<��� 8����7+���� w��\�� 0(3��?����ܩ��_퀺�ɔ�� $>�yw vqr�� �a[\��>����`�HI p�DR��T� ZU�SQ�/�����w >o�[�Dp�8�X ��24�� ���(�恤 ���*�RE ����d�?8����@���946F"AT��=	G�x�?\d` f^�v]��[�� ��S��F�@ _��h���� (��8���X� ���F���T�����}<8�_�`��֩bfgy ~}������SJ �R^c�s ��yY�X�	�]���0E_8�� s��T��34����d�� \�m�u�$eI7�&�Pr a����pn� R��S�� �� �x�:��� LG~��a�� \���N[�� ��cC;:J ����u�� V�[`��B��&��)�S� :H���� @��.u��d ���� <9;����*w�� IHz��b��w/=�c{�e��i��8L�\� dD��]�� �����>�ϓ�� ����t
,Pmg ����,�	�q��Ҟ�mhjȥ�g�l�v8Ȁ�z� e��X��T �I�ZD՗�ʐ��g ? �р��14 ��T���`�
�#�� 9�����/ �����(u� ��'����8�Vos2 �r�W, ���@� 3���<�e��>�������� c��"36�� �2���)fŏ�{�D���j
��'³���� ���G���} �������MQ ;��u��_� �`��d�� ?e�{q9� �s���a� -0T�� �Kr�H�)$�W��'Ljs�����\����z �a+��R����� ��%*�o ��v��w��x��y�Ç �t���� �f��	�$�� ��7i ��z��$Ա;�� ���y���� ���CHF ������H�� #<Z_K{}B0"9�pm@wtCus��$ EGM��V�� &9	<����� ����{�� �UQ������A�%�,{�u� &+)���5 32��ĳ��H� Bxy 4�v,zs- }�;���L��;QP�~|������W��i�E� �r������4I� ����`0�� �WU6;9 ac����tu�% '/2�� �y��p�� g��J�?�� �Hvw �`T���� �|8��?�j SN�_b ��f����.N@LK������a�`�c(`i�H];ol* %DG������h� ����g��� ��25�� �8��� �S�ݼ�|[)��`�*5� l�ȴ�9W�T��rUS R����ĕjqlL�� 10:B=hm û$��87�� ��m0���y��p�@��13�����`�6�0���l�� ����w՜�S@���ȴ���q�L�񀿽� yzxv�ͺ����1� �LƼ ��<?��ql ��9��zPet� �)
21�� �ś$~��Z<��?����*�s j܎8����Lqew�؀ۮ��GI\JP���  L��_�&� |W��C����}q���� ����+* ������I�s1 ]���[^�)y+@RN; ʢh���q( DEIA&@8B�������� ��dØj���[pX8&'�0� K�����"GEu �@��� �JR�-qY� c~�K��� >��R�Vl ���� �˰��5��l ����| ��S��Oc �R�slg\� 97q��~�-� l�i�m	��T�L>t��̣V��*6_N����w�0 �sX��Y9g���p� ��x��U� �W �n��88�����
��u$���4�����& �ƶ���r ��uoZb{��V�� �k�pf� ������L;Rs��"��٧��P���͸�� tO�S�_� $�r��iߴ s��D��Q����`Z�xp� �b��I�z'�tg 9��
�>kO���H�fe��� ���� �å��~�����܊����ŵ��� �c/�jHW{L�XR o�Ҧ# H�k��"?��Z*$���lp�u��Ƭ�i�b� q*�U�s� g0���}�|�ҵ�ߤ�k l��Y��Z��! M�U��T���E?R`wH!�,J� ��i���> ݸs��6>�s��5TZ�bI!�*t���M���,i��˕ VfIt��~,ܱW7]���r��^�ʟQ�u(�U� ���G������� �4�]��~k(�e�j<���mC��g�2��rg+:J�'��S�x a�n�s�
�r�i�f��\8 �P63�؃ U<tnY�`�V ,hΈod �P�sw2 %r):�FQ ���P
�.�rx�?HJAp�3��l|����C}$;�<o�'P�@2�=�֌6���Uc ��d'��� �I@�0�5 ��)�*я�?xn�p�6�2C	���0�]������>����u� )�1q(�`u ��A�; w?�ֹ�׸� ���d E�̺_X�uP�p��>���&a+ �}B�` �N�.P?V� �M�b`o�=� �!��P V$���;� au	�R^ �x�������#���P> ��8��NQ �Z�,��~ S��R�n�7 x0hr�dW �I_wYTD ܪ��v�VS�1 �-�f��E��M������� g�]�;u� ��.�[A�<<���U��� �H�'ؘ�h��w��/��J�_�W*� ��j�>���4E���� ����OJ�� '�����]�*�=�?@�Ŝ^ ��lLM�"9 � ���� Activa?�n z2�.w�T �������L ~:
�y-0�tWH/uw�{�c6��s� ��c�&P�  ��uS�7 �׍O) :ht�n�*� ��N(#0C�u h�鑈 F�s
�%ZX�2 �d@Inc or�e� >� ��!_M7 2dS�Ҵ��vQ$�����l�/@���� �	�@t�P E�rz�l�������J۸ �ӸX�#� ����ʄP� q�3�Q�͘S�H �(�LK^�} �]�~a�� 1��uV{ ���A��� ���/��� _�$4ryp ���<s�a |��f!;�d i��eߖ� s7ha��m �6��q=s� u�-�@ Ns���(�)�Xgh��1b^ pr㞔7ly��,��.��P�="��u�$�A7@�N�8��� p4�{��H� ��.1� T����\�)��J�3�쀨ʍD4U�����ҮrI�����{�YvW -P����	 I���'q�B�� F�Q�M� ���I߯� W�ղѫ�$�6䇕����?��Q�j*��`Q�\,k�Ե��M$:تu���%S��, �kG~�I���֓���4A ���W��,�� ���
�& �K�ץ�~' ՜��:��I+�f���ߐ��o �
�7b�� `~p펤1aj�֍�G)��
���A�F5���� ExK�|2��<����� �vZ�@| �7����U� �+����� 5Q��v ��&���� ��*�E( �~�,K)��k����  �5g��6�V Q�!`n�t� ��SN�� �E�iJ�A� �
�~� ��t+C��<�i �uW$
:�&��(L� �A�����%Zv@��� Ǻ��~O��?W�`�d��t�@�8���: ��.�ԍ� ��e�� �����I���� ��@�C�f����_ �);��A7n����l�������; ��a�� ΐhR]L�QwB�c�:��Hs= $�
��v�x �&�"X�T���w���� 
��' ���o��@�FKu[��D���tM�B�����)�l�TK�F kV��E+�4�`�$� 9 5U����OySR2 F8�C|}��E	�M� �NT�3.!%uJ�f��5 208`X@P %�#E)�� ��/��s��B@��'�˷ �j�_xn��M�������&� �)%�3��� �hj��'�;�� �}�4u]pZ�OD ���+ �`HV���?誩r��`�\8 l�򠍻T���Ӧ�zSp�k�`� _�8M'���j����; \uF���" ҙ�?�6H �hp���� S�����{ NH�uQB�o �ގ ��� ��kX��6$90� 	�#�*$��* [(�����Z�e���"� {�h�JS� X���4� �bG��� �qW���VZ �$Q��H�� UKD���� 5���S0�!1TH�3�`�m 
��z����X ���_�����⡣p/�� '׋Ht� ���u�P��o �%��TXl U6tg�WAe�@�`� �ͺ��+�a W�T%�uB �=pɦZ� �4���zxG��Ⱥ�[rD}/ X�]T�UP��*�~CW��' �(�<����.[3W����&:�s"<�>'@	)�`{U�t�8��� �,#�O ��zi_q \��d�B`k���,:1�y�1" +��A[�Ǫ@��=�p� �2��-�/�6|R(�H��������4 �IDH=� �w�VvC +G1K^��� <u(f�F��8��d
��:�=MڸAg��  R?ݖ;<�7�Zd3��2*>T}�O�%�zp=��$@��[ ��P��Q�d�w��5��� f�'#`�� ��
�,�����x��ܙ�A ��EZ��N ���W�X�T ype�i/)]`��}d��lJc� Sߥ\7� 5eO��%s �WINRT��SE�V��&���LA?NM��(�P媳L�9 10`�
H  ��� i?ߘ��� ;�E3K�	c"{D����އQ&Y��T^��z���=�H$@�(� ,�0�S�{8�4���)�cAN�&��. �t�,�l�dg����1�~�=�P�@���� ��g��� ·�r�uZL��I�@w/
�yi����� �Fl�� QO[26 (�@�X#p J�o3,�W�rk��J)���pv�}>.��� Ad����[  �u��Ho~m Edit��� �fesq -alX�D ��i����Y	Jw�����B�s�=�q u	r�2�y���}�;]9A�E�.����i�X��ul`DV �KqJ`��� $cja�k?Ui �;B|����9gI�@��S�e}~��C D��P*�\@rYTE Mo	[d&��rn h����)( �����~, �Z�c:Mw� �Be��G� �7.�[�jX�4 SPhL�� l��/Z��:���%���bC�;Az&áR��9 �u�~���O��K��=D ���ݒ�Z ,tWNQ��m�
"��򂧸0�� ;0>}8��J �R���D' B�+�W[@>><���;�}
: ���b�� V�Kvc��� �u����Z�n1���zp~s�� U���B�JY�Fܸ� ��0���l '���x�AO ���3�+� ���v�9 ����x��s� ]���#w6 g$��/0�� .�*�PI� �}�$c
t j�;�l ��!�C�>8��ӌ`����_ �j�U�Z��O0쪀�r�@{1�? 4��-� C_���3?D= ��&r� Y��F �P�����"��2|+�� ȁ��]�N I�ià_v� *��"�� mV���/ ��< 5����� ��^Cv] �1@Ж��L��H�@�N�K@W ,ru��]|�}���IX�����z[+ƙ3¼��2� �RYf,@! ����k+t� ��%u��ڠ ���Ĵ=]����ad�1�������b�+��@| ��o$Du0R ������ (X	�~� ��+Z�\q �)�@SU�P	 ��F����Y6PB���q _ Ak���� �jC� x�d,|� f��w�4 �o�{� �n���h}J���md��A�����wQ�$�(��K@� =P�YbHk�V�Kh`�+ �z��y�"H�D1�|<>�@Ju���$ �����C ,�t�J�	�%����	.? �N��%��c���76H����
	7 -PA��U ��{6��Q� �s��G�\��/!�x`��D�ty��9P����퐐|�� �ɡ�J�d�r�'f��	�
y��Ȝ�imQ4[�$��'>^�b-��H�w��;�*�<,�d@����ڗh�kbq
�d�(>_)pKt��R	V��>�����Am|80t�d	H.�\>� j�+�ev� <z�֙�� m���,Lٱ.] 6˻f% b`�
,�r �$+�3���] �<BL! l�;x"*��L)��$� ��h,qL/5 
�P��I �W-��T  486DXiu ���V�r0SL�2�.z�`|�}yvK�Wri���b��T E nh�W��J�4.`�P�] ppm��09�^�w�IxB�C ����Vn�� ���X�p0u�1t��@�v�$�&P(�� �%;�)�H�4ؿS�� �js�Ppޗ�XF��`��>�D���T	��������~�q��^V�'�,
&	B�Q���8i%�F��� O�\	��K� :!@�)��û2bx�糗<F|��B'�� ���Cy�1Lrx$�M�2a�GX`��S06���C���>�PZMH ��"� Ӭ�����	$�P���4�� �ȨOp@�x �P� *��	��� ���x@z�����){�4P��		�� [z�Kys�?d#�7HC���Y�j"{\E�Q�>�b�`�\8��u���d�`S0�B�
81@CL� D| <��"�AMz�\�m��(R)J ��pW*��y-KX�Ԣ0�ӝ �1?�2 �3�R�L|��0$j��� ��`d3.�U nk�ow� � q��l0� Chip��\��� �Q�L�} i�TrW�me t�>C=u�o�4�N@�T���E�X�\��` *1�v
/�]��p.�r #tu���x\M�|�E��̄@�?���PۨS QW2RVvs# ����5�h:(P�1�iKH] z��	�v}>���'U��M�}� �;�������zdn�����	 �pq��iIXA� h��$c��`O� �RX1uL<�r!\�3���ad�*H $)��� O�����c)�p�Ћʽ���ӌ��8x���;"� �]�O�(9�0�$��~��6 ��%>��s1����t ��CԍS]� ��9���!,��*O0"��g#��Q Y���T��P?�du�f_��"� �Q��;* Pu'�Yf0 �gH�m�� C��L~��*,�9� ڥ��p� j���!�
���]��؀T�)( ��[�Jf�Ez ]��@��)� d+r��:�>�� <�@�Ɓ���� ���E3L fH���{ ����G�t#��º�<!��V+|`�X@E��b�*�⊬s ZU��^��_YH[�t �U�0Q�{)��N�а� �Hʍ�t��{P ���6�� M�5B\!�X���������{H��^)T2Q�� �b��+`N� �E���8���W쀳��0 ���}��;Ë�ⵏ��%\��}F&β�.� �^6�4QEb �Y~J�V Z%��7�2N�\=x��s�nSH.TM' �8�+�E����J��`O� C卬5ɺ ${~���|OP������� ��J�>؜���&h 凌~8Kw�9d����=�A�� "���[��?�؀���j��J�� 	��G�c�3�s��"�d	H!�*�:D JZ�cl � v�g���Pm���d���[ �@FR*<�I��	���B9� �d)-�'�R	O2�$� ���� ker��Nl��D K�/CY�	 ��@G'zW<
!8d4,0!oв(B$ Y�*R��6q ���l�� ,{@P ����Q@T�3J ��؍@;�0�������z�%`�d֨ X��G:=3 �UMoĐ� 洗�*�V=O�3X�h� w�Z�n�� ��U~'0�?��Pͭ/�$k.!� :��dD��� K�'�U ۮ
V6�s=D���n��3� B����v% 0y��!�;� �^�e@�S�� IA� �R?h��ɴ~�b���� }%YZ�LV arFile"{>|� O�/�ԟq (��U�����A�t�`��Q?(f<7��ο��$⡀��#�z �p��WXP ��|�� ��ȧ$���p�� �2_��=�ڸ� �C�����q� {P�eh��1��Y,�a����W ��KZ�投 2,�)��u ��ҒA� C]���П^ .��g[P�m���e�O0?d�$��\��H ��	|rG<���Q��R�� 0�Com�,48sS@�+#p	@y}��,BH�*���Y�ma%�L�q��>����e2�� )�/+�#�G?	Lp O�,�TiVE�YȔ���$r�lK���\0�� �CLegPZ�p�[-p�0�(�v�w�cd���ksJ�!XqOr ���Ľ-�#��k؏Q /�`J�\� ���%�� <�$Dv Spec^J
B u�dlD<� 0M�kҁe�� �[�3�C j���_�#�"@/C$�gN @��_�'��)͜��3 �%d.�s ��qt�S4�2�x�І�\ �F���Lib !��y.�$h��3'D��+]Ԅ���U����?��N=��Uy ����3(�|���^`���8��>��QR����B�d X�.�˕w �8��s RN��?�6 �Hχ��q�����1�_^Z ��X�8�� �9V4t3�u v��D
GgL�"�MX�p<�Pw��l�uR�i����& 6�C+�E�:�� ���B�,�H����CȌ� K)*�� ��N;�G��M�~�B��zFՑާ�������a�;�0 �ˮUA|��� ��w�� �԰H)�di=��C�����$ 9�f	��
/�zԺ �r�� 끜j]Y�M�z� ��w� $���+�� y��v���0�E `������ .�P@���p�~,��Dûp}��m <�u�]To$~O�����S �2< �,� �'j�C*\�$ F?9� ��T�C��* M(<0�.� N�� yf�ب��b�4K��= z�|^D� �v��t;2 u�F[Ãjz Ic����= 9ps�ҋK:ª �Z�R�
]O���d \D��0���� �t�3��~ ?G2Ϩ�e��xO �.��Ήl| JG�^3#� 2'�.�� ޞ��W_�Y *kE�$,�xD|�C��ɂ�� ~#������ �p:��3֍ #��(�uMN>�@e2�1 �o�4G�ڮ����REH/l���w&$���
��!� �ͤ�Ԫ %��T��� ���-!=�ꈀ�^@ ��"�Z�9 `Ǎ�0��� h���	�0� �jD��/}�� �Z�qH�( )7"� ��B�U�`��m2 ܈�8��˵p�� e6hl\ �.��C��� 2�WT�S"�� (#I� � 0�M�`G�ؐSޣÑ6���"�{Cz�̏۠�xȓw����'����=F��_m@�<D�3��)��C���oQ���_zO��!��#L���D�1�����4?S�?oQ�,���GP�-E���������l hatp�kb q%eiuw�W \ ����K� r!"d�4��Ox� �l�nfh0`I����R_�%Ψ��/(�� <����\)W��@�J�l j�;	FO�&�"e ԕ}��-ߴ�@+>� �O���f#C ��p�AJ ��O�����r� ��l;=P(h�)��qe��ET@Y�8�]$ �!W��huu�k����6 � �Ő?�߻��# ~]'�/h� u�X�i_�� ��}.(�Gt� ��J���ȾO KӸE*+� '_GZ�m�O���n���ր��(x��\!p'P��G����% $o��������� r9�8� #�G�-�� iw�tP�$��o��������u� rЄ�v;_��>�O-]|X �.u��w \{�tL�? M����� �鍇S: �)
u�� �	\5��!N�˃�Օ��A� �L�,@��u ���i�#$r�n^�@d������?%hH�,�0u��u ��1�\�U �-�7q kF%�d�IWYL���s&��֦[�%�� ݂#��R~ +������&_j� ��.xQK�`�(�T	zh f�բ� �7}��*� �/��|߶���tr� �%祹�F �~��� �{�p��5�(�Z����)���� �ǍcuN� �_�YPUS G�,�ϋ 2`7[WV� mΐ>;���� �k.�N� �x��Tu��H@I�C�� 0����;שLF�$(&&G���: yP'�x4 �A�D��� �B~�&5'w �f�9� ��֊B�$ �7��j�U���������� �'#Ҥ�=<B�𜟀t����vi��`�1J <W	��!�#��`� ��TD�K,@�FX�c�p ����g� ��ְ"��E�4�W+�`���������yU���L x�'���N ����E�sG�q�H���P {��A\��0�ETr	u-�
 �C�Qc�_��� ��x�- t׸�]J %��8�|��B(��4�E� �,ɫ�	� �H(��eX�d �K!�j'	 f���?� e犎��(���s�7) 4K��W�T�>h> �R�P\B��1$�� �+f	�(* )�s~ $B�D��x 0�Lz<2u�*�m�&t �����>��_��8��i:Ә��u�V�Gf��{�PD@HELO@�Us >.Wi:th���u� L�$[B��wq������ 8�����x ×���9~3��I<}�CB �+� �)��.�P);�4���L�_T�/O� '<� >-|���B !IUYЉ/ '�M��x�X;8u �RL{���pI+�O|#o'�@L  FRO�:ڷ �ʼ���� +��RCPTx  O:���>�D �މ]y�=�������*�8)�Z,P���2��Kue�^�M���,ܫ��;l0����(p���i���@�g�h�� �%"zVP
m����eĨ �k#� �o�`�DAT ���"LF�	$m���g��~�	�S9ub���*�x,�� ���(-�[� 2?x</�l|�;c��g�$�=IS f8�5u9V1L)!��zC�@��W `�od�pg� 8XbV_�90 "}��,��C-���~�Iٴ����-}&��h@�;8%v ��4.X�i�>��Q8h�>�|̵ ��
����bp.� 8w�&��� ��.� ��2a
=,�d]Z/��s�P� ��/�d�T�ڰ8O+ k$�H<��>���o�p2y�T'xt4��.�#���pu bTm�t�qR���r\<@�s 	P�J�� �o�r�Hu� �����}� �A�ws��0 (�=��Vro,DiNZ���;_R� HhU����>.�P  & ��, r��QW��C�JP��R� �@x��I�>�f�&�Q�70�� 7_�^�~� ��9u<\����M��ܽh^zZW���w2Y �c�@��}d Ȉ��b�� ~��a� U�y��k&� T���hP� ��m��{%"A,�6I`�~d(l`�|" B���#��0t�� �ౘC2ihy�a���W� ��?Puj� !r]��� �3�O�K� DN�Ԍ� � �/a�ŵ h�2����</	��w �_���&� U��y �u,R]:ɺ�2a����	� E�'sh��g�+ (MUX� @)E�>�Hz>~�w �'dqfK� Q����) Յ���<?aL��3߰>h� ���`@��� �F/�,NC���g���	4 ����E�ݸ�`h씷  RH�I�j �e����B4��+�|�uǷ$���8 � On;"Q fqrm�`V gdl��XOS<�$��M�%�G���_�@�aH �4jx��N��9J��@X5i ���p��� E�vC�  �D���@� ȉ�́� ���$�2 ��H�d� 贯��� �!5ĭ[l�����j�@E��G��5 .^�(�Q�u�iHp%x�� �L	c�d�b#si��? M	�~� ��!q6i� D��8=��� T9@j2V�- Pf�O��0�3���� ?h�����9gH��� b�+7�����ݢ�h\�( y/.�3(u��6 ���� �EWh�:uH m�x^4�7� qIi��-1 B
�	$D< mq@k`�?3 ��\�,=�.���@"x�-���)9+ 8I�%�^�_���ؔ9)Z+���_ �H��F��젠��{0kXu� �Z'����� wLej i"A���*$7F n�"`!c%(�5hԸ^w���j�
�1�p�|k�q2�:(�S\�� l1��Q� �����7� ��	�=�W`<�h�F�7(P���ޝ�B !�ة'�f����L��Q�7 h�gt'�� �v���d)x2 ר|�C �#���ȴd�r���9��!$Đ�@�d�2�%�������+ ���,nI���g�@�9\Z(r�L�� 2�DG�7!{�@�&�X�9���4#����G��� �#Wdp qjl�b�o���H@cefA�uw?(. �N�9=[%�]�`�����x*<$-�_s��P> N \����� R�w�XV;GC^��xp�=O����S`�Q	� C�8&�%]N �d�0�S�AlX}�� љ8� ���%"D 2���x� 1*����� �A�|;+uVU.X�"Ш8� �a�&�� e ��#�\+� A��5Oh ��,�]B;QE*=Y.�����9,�� ��T��-x� $ul�%�!v :��;0A pDlic��� d�R:��,�� �<)��-�?X7?��T���A���8�) ��+O���:%uƳ��,R#
�=���_ d1�f+�P U� )$�t"��2�u қ���XS�k�dI$( J�E]�=�'��� D�� �<�8�C����0�:,5�* 6=(4�tr� rgpCbw� dfm(�he\c�
�P�@�H 	nj`e�� h&Ubxg{}��Ka �=*|RVL�5���+Ql%j@���I�� �p�n5193�� ��#j
� �%��>zx� �b�=ep �2�d!�D�����1QS��$9qw�s�v&ubi|)`��$.Lk�o��(�{�� *�V���$��5�"t����<jp�C QY%~�ĺ[Ve���Ք� dr.J��V ���P��=�a �/�52' k�Q& �\OC���a��M�;� Zi'w�R�����^����DO��0H�[���I��GJ uS�Y�
O �։B���D/����Q�� ����/-��*���b�h�S��'�|C����]�Y����H��	nh�%���O�� �u_cQ�� <-����MZ� H�Jץ��yW �'t�@~�ivB�2Џ� /�(����� � eE��[:��*���BN��?��q`+@�"� ��'� K���Pf@�
�-3/���� î�:�m\�	 P��2��� %�B<��t�?	���PS̈́�x �)nD�m*�>$��8!A�|hB�����3� �H�<-�f�8@��$� xL<6?�p �h�J�V#��>���b r��W�hZ� ��V�m B�1��GeŐ�/��u�J �
K�c��9xI|<N�w�-] '��W��Ų:�f�g#�G�M� <�w;�s�3�ѐ �:���H8 �<��L �[��&��u��>\�%B��M ,sTH�X�� �����; �G�u�C�n��ϨK�h�B'�	��S�� W�b� G��8���9�Fs�VC�^�����1�v Iz�����J��� ����f��� 	�5 ����u�1r�^ڰ� [���щ��n�G~^֐��L���� ��[�� 6��� T�?�� r \3S���/�Y`[?�x�R���H��{=	���C:
 .�BIu�$��+��JZ�e��� C��$ B�32f�_ �Gd"[ {YZ��y �u>�T��G�P������x�/ ����  �p7�;[4}� B�ODC Ư��1�2�:;�u��e v7s3Z9��G=�����/��H���P�� -C�k�� ��&�;;X��+�$_� �����Dx#yB�~>�� �{pP X�vE�4F���ܛ�2.����'Ҽ��	��ط��u�B��[w�DQj�ο P��=�`�Ð�p,� %���)ST
����s �W0�u� J�&_x�c 5$��ɸ�a:8?�  �=�/�UJB�t����PC��~} �Q�ETP D,�%���i ����0�F��]���f@�D� �$�U�|E
&+ƀ��˶ ���K�V	�7�Õ�D`v8�0{ �Ձl"��Es[�C�a��K�' �֬�� ���)� R�H�%�d� ��`�|� �,N�4X��� ��	���.�@�* �GPj
��;I� c'C����v�$)HP���A�,NA ���� v�Hܺ�<�� w6|0�ߴ �Fo"� � ��w���(�r;77���E �vF��}8�� ���'��Sw����_� ��J��P& E|p��ܙ [(��Wi��8^)P�<uh���B�U��^�Yu��@�
V��}�'Ѵ��� �a�t�/ v]�U�!} T8���� t��bԪ �6
��k0^�q�@;E� ��u�՟�% ��t,I� $�X�ݫB�@P+ �M;� r����>]=.� <�v9����]����y���M���J�� O"��4���9� �=�%u w�-��: ���,�= $���Q~�s	�*���_�)�"��3d�	�]C ��I�}�; �战O�8�9�+�b�� r�v%�^A�;9 (!�׀8 �u@�.tf�ǧ��@�u��`�����|� �S��C�u �	���b�T��?]�) -��f�$h� l'����� ��_m0�B25WVh����p�K ��D�ȍ�,t�]���بG��p0��hS$�$��r j�͜"d5��@_u�`T N콙�b9 K�+�>hJ� ��\MC����|�8����P` @���B~ ,RX�FlM�f#&"8�(ǩS��5��Wx�J�.СZ4:�����*��� ��u�h |���f@$��!p*
�� ٘I�4�<F�!� ��YN�GҘ :H�Ws %D�9� 
Lh�ItC�w?��B,��E)+�2H�z #�Y�:� ,��8�2W�Q���+�/�7��dU.N�^ ���M4�*bc� �;�}�."�K��OL@|uD�		�T� �A�V�PI�GeKt����d{ zqs� Rai��Exc���_��] ��ŤS(���81������� *�59�L.��(>NG ��� %�n�xL}	d=uO��!@K^�����a?�� �����iY �}�۹ ��=�~�<�Ǻ��C��bD"q`7� +8�%>5� ʃZ��ǲ ���D
F� UO/�,�� �_\��� I�U��� H�R�m ��'�0� PS�w��B($tv]�A#+��솥x�|� t	�,�b�8 �j^z�h �G�`�c,�
�FH�s%P���m8�61��B�<D���']� �����h  ��%�Kӻ� ���j�c�:���9���
�� �o��-|k(�8�؏ޞ)2 V��3� �>����/9t�
\��B� ����T�^��`�I]�3���z�cP�j%�JЋۀ/�r��><I�j��\�%Q ���
$RSWX�� J�↉]� >{<�|;x\���sa� _[ZHJ��h ��{����=���Q�"�� ��P�y�� ��hR-��� >�Ek�v&m �M5�G� z��F���O�������� �X�Q����@�r<��pThe�x�_d�k�2���ul��	[۽}�8 7~N��c�y^m��f.  k����}LOƆ���y�X`�d]p �g�um/�{�| �x�W0|�� �Љ���3;7���«�L^ Q�J0�M�g  �C,v ţ��}�� E�u^�W���H���������}��` �k�$��~��	ur�ȀP�ɖjK��k�p �%}���d�G"@�XL��CD@�5� �t"	6�:�7: 9&�]g |*�"S	 ?uR��M���d&Uٱ�ܦ�Ჺ� T$_� ��t�8BuC ��kJ�)b���K� 8 ��B��tWE:J�ʈ;�]:f	�S������ �pJ���q ����;�t ��UwXz$Q���	� (�Yu�I�	���0`8G�< ��w�\�� ��O��ߘT �~�����tn����<� �����Ʉ� ��FZP�" /i��4�k	 _w0����� �E2=N |@��,�RU��/�~�A���FH��g
+�L�D���<a. G�4@�` FD���Ʊ ��:^7u �b�PU� d�z6;B.�2�a8�$|Eܑu &�>41�u ��0��� О��`��P��BJ����6��_4�Ā��&] E
{��HP �:8|CV��� N�D�1x���'8��W�Ҁ9^ w����������JԸ)�������kw ��=�$ > *߼|z>ut��Wŀ/��G�\��B z�=�� ��L��Mh/�W8k�@�ڳ ��,�>R� ��h�W� �%2^���+ [��֕�&�s��;:��%�lĔZ������`��<
ˀ�&/V<!I_5`�Ye�(�ش� 9�ӨD����"�ăȡ��̸� H�;�N�� ��mTq�8Y ��Sޠ�L l<�ܻ��� ��u�� S��T���p� <��/��U '��� 1~��c�� @#�G���T���f������yz��ڷqp�Ї�<}6�5$ �Q.l|� ������pk\u �՜16���H �&t�a��G �b����9c06z��p$b -��^��8�� �9㠡��pP �1f
�{Z���}� ��t�y� ֨���nh?�
 ����q mW����3�p� ��NAH țj�`3�\. �+�t �{���Ya�1�u�r�e`Ϫ� �oAؔ�qH1�0_��P{�h�s���� ��D}���8�# �e�$�u� t��u�s9j�C }�Xk�� ��Ou��� ldC��D���1��x	�X_ �] ;��'wL���	� ]Y��KP�&�� �t7D ��Iْ�*o ��؉_�:W� �4`0�&�	9=,���߫�ט( ��%TR-� �G�9��tw P��u��B���}���p�� |��mw���ƀ��0;,u ��bCS �NU��~.�	��u��W \�AP��+� B�r&���'?e��,c�~N� I�v}���ܬu ����� H���K3�x�{%����D���3��~F ���i/� K"r�( ����:�u �a�������+���f�IK W%����� ��=��)u �:�Χ���
���1�#R��� )4a�:��98͜ �	�ݸ|�����
m� ��ܘ� 3@�P�9]p��������' ��x�X�� X�,�Ac��S���0b�]�a�J����d�$�bx�̠Az�-��^�9� ���B��� 5h��s�Op� W�Y�qV��hU��[|M�lA :�s2� �/!-��� E.����D >���	h �%a9(� �S�,���8� L���uٰB  ���p�6 B�@�����m ����_�S�u���ͩ �L���@����X��0��z�)�x *�F˽��1�� u!�f��= U�mnj� $h�ө���< cdVj�!�  ��q_ ���� �sۦ%�� `e��qu�`hL��)|� �^D�N���$L�
��r� �U���K[8u� �����
F�G�s�B61�.�V�@���t	WL) �_��N3�� ���P��<w�X� ���= �Ł�H��}�,�X!=�}� �s@r A�o/�P� J�=w�N)L�1`��V��?5� �(]Q+� l%_�D̟������� �<| ����Z�� ���.� 7���X[s M�_*��j �ؼ>�B XR��,��8[C������^����cTJ��4�}9Y�!@ q�hx.�d� �^=X�B 0y�\�_�	��� 
h7xT������U|�R �8d�F ��>t��9�0��~l�v = Q�{p �Њ���% ޯEI�\��`�)NwY-~��G� �]Z`
n;/c��@Ӏ�D.th��L����'��L� ��
3_ T��^RТ�>t"�%�}�����$��@�W/N� �Z#	��� �"�%z~Lk��|����H� ���8. hV����~ �� �vB�N�����p�% V#�(�if;*�]ۘ�ߤ |�_'������Pkd��ؓ�2�� +HhsO^� �����-4 � �{��i&�� �C%� ���c`SR  ��C���V (ݡ��� �u�#-M���P� s�� ?'�a(<�%�y�����Y;� 4��W�dX53��<e��l�N�( ��xB�a�h �!Cb���(�vEH8� ����`��� �b��@Ux�8Lc
�;K 41a� �_���֬RP���:�F ��&�� C-� �T�9�@~� 
u���b> �S]��Dc� �-L*���H�� 5[��!Zx �|� z� �)�u��i���7� Y\J��L_� ����!�8w^ #�XMB%u�n>�ȸ�.$  `��	C� |�
�6�� �TR��J�&� �dq�+�\�� ��yj��m ����ձ�� >�,͹P�O %u���FH�@���TĖO�+=�)���N�d�Z~�0V�tf ƊS�qTx07�PL�{� ����`O��v�hk�(懎��ڐ�rU�A��t���(���+��2�?�B A��,H�V !�@���� �N�~$[� n89�*Ut�_��c7� ;^�~�)K8��#@V|.ң` �dh�Cl_�%��y4�P��}y������k��'����&�^ �������6Uspd&r�J������pM��R�'_�|�V ��>cWx1�|�< ��K��pa'W���T��/e~ �\C1 +p� y���,�K=��4
��[�AI`�4�Ԓ.��<��ٜ�dL����<~�� Ä8: �u ?@%L�+��0�Xtw��{�|=�@�<�Y c�_O`a|���0��>�V>�0�� �w �C�W,��נ�d��ˆD�k�.�(YC� ��ag�ϐ� �����>Y� ����{���0�����y��z�
p�HB� ��s�5;X�]��ԟ���� ~+s�������8T ��W��yb Q�tkpC d�	�H���"�E��%�4� ���,�~��8��� �RF �<$�NW>{*!&����y ,$}���� U�_��
?t@'�,�����( ���� �����!'�*D�W��@�3x� ��ZH�=� ߗEe��� ��D[ 3^������:TЃ�u���2��I ]g���DC��W<��=�������� /����t!�@>��d�BL����i��q�￀�^ �)DB�+�����r�% �Q��B,�O�I�g�1���S �Ƴ�� �Wi-�MV� 8�Ȧ��Tt`ʊ�� XP�� *��1U�p����	&z�� �Qr� *�-R��X� �zH� \۴ )�2��?�$��H��,*8�p�DL� i�k�H� es˄Z-;~� �����<��W'����#���ʇ|Q�^�p��
�@��s��+������<���1 '! �BԎ�G��6���wԗ��'�H��T ��ߩE�/ (u��2X� �z��)U��� D(9H
R7� r�٨�W� x�8BQ�z ��#H*bW9�`ֺ��ӰO��xY�n(��� jW�R��Z0�.V/aѬH-[C`�i�N�ȃą 1SH�yU/H�JG�����;�V��I��! p#"��&��*���H��+c/�@������-JҀ;��>� ����T/���xY��� ٬vLk��mĩd���#3��^x��!���x� ����W����&�ү_�^�8pE��I�������!x� 	.�K6�(T�X�rc���Dn�r�g���J #�?)y ��Z��P �vDr����zy	��� C<(����H�'��� ���M�įg��L@�#��. >_�y�[���v� �MY=��J����!8�(9DH�ߓ�����.t ����Uwe�5k�g�yH�{�� 8�������:�K �ŤݦJ;]$ ״'�t�qt� ��szrS�$s�<�������o��u�g'��$�@S�7P�?f/w5u� �G[` T��<^�d�O'�H�)L� ���z�y<A'm&���-��W�����C?,��F 1���+)�Y
i�W��I�s�n୳-}�}L?ĥ�0��#?��_-l�>˻g�KuM ,%5�)�w��t�T�W+�^/��8�� 	h[���� 얄'��D�� �d./EP��� ��$�,:��?_B�=j`hs� ȺJ�y��Ho�u:�n ��c��%Z�\���o qeDb
Ò 	��W���C1���0�b D��
J��.�\Å���� ~
%u�D �JT�܅`� 1����'?r JdD��l��� ��(�<@ ���K*#V $���ͫ �'"LO��� 4$�38�� �@�ty�� O֢
$#C�uP���E �W"-�Q�� �A&t��3!����1���Z_����ܥ,}�]9�!^
��GɤQ�l�+ �կ� Ȳ��§ ;'��؉s Q�	\� ^��,����yr˻��L<��]P b�Y* se� "w@ ^�L�������
��r���s�`a6�08���~V �U�Ye� 5���Q� �t� <�'3�= ��0W~��B �̔�e-�� ۓf�~�X�@ 8��k� �:9EȔQ� �Js��\Fi���ީW��݈Ob� �CdK�� T^B@!z�0tx��|����P+�9( {���8�� ��C^�hY�x)��w���X6�& �Ұ�W�� pd���* �uj��T+"�W�K�!� x�
�"' ���o��ɨ P�������� �] ���G /�}8�EH�M\i=����,��X �5'Un���i�s��pM��� �;E㯼}��F�t�`�?� =� {��ߡ�ˉ"� ��Z�#~G?���z�x� �|���=�e,�o� �'�z %�*��5 ��M>7i �yeWG�T[4�f�x���B��*��2`JE ][c�� 7�Ǜ �$.D�?�� �*��@BH �D�kߝ �d���b�  �u�t�7�g*q��TB�R+��w�H�����G$P$�	�K �g��Z �V�J���r t� #�� /�ޓ"�$ <�%}���f*Wg�d�� Yi$)�_y�kG�/}�����W �+FP������@����}���� ��) W����ZxS	9��_�b��\� �!T�<)��st�,��8�ah���z({ "�T v_ �L^�?#R�@S�HK�9?{�?.9W _�- z�$Ҩp���I��Ly�F� ��*��\� ����ڪa	�)�����G��R���x�- 4n���L&�@ �rU��� �R�u�;8�����'��C �1V	~���߂�@f�%O$�H��I[�	d 4�s03 ���e׿�H �)tD��uoz�N� ���@U~��y����Ҹe���D"��B[%ou`=2�� f�nO�"��� �K�&�iJ>$j�����y)n^Aࢪ�t	 ��)�� ������ O+*��Q� SŒ��7">M�E�����S��'�� ��o�[`<� R��j��w<����P�6�K��U�cB�Y�#� 	N!ϔ�� ��k���tz���@�? .����d�� B��$W|�q�4 d�H"�1�@DO[�gs$���篻���� ���u�� G��QU�<�7 �K��vDS "j1k^�BHs��F���:��r.1�� *�#�
 �[VQ�=� ��2]1v�I�j%������� D���_�� 
�j}P��� ���z]��.�� >� ��n/��QW��^�D�2�U �c[r����	��|$� x,L�S� N�u%�]� o��v�	�����#%�_ ��G��@�u�-p��D�
	S�{�����W!  o�r�ah���A�`�� Xe�#jKظ��(� ��s�/ ŇcK!�� �J[qb�����尸*�PH7/W���`|o��YΩ\_W0�������� ݇�O� ��bw˴� ��sS8����We� =��t^�X 	<��#u� K�w5�i���R��4�L )�?6d3�7 ��ƕ<�
�YZ��$��9Oe �*C�DKg ���l� W�>�=8S�N��V)� �B+�w2��y1cG\X@�/��LW� �0��������� U�$�� u�(�Sq�� V-����i	Wf�R�J/���8�sI�V�܂#C��Y� j���[NWa SHy&�o<%�CA�4�k�:q���'1� <A�#-�:�r�F w�%W�P\�o��(e���V[ =$���9: �R*�h<� dU�_T�D ?΋
��Xcw�U��RC�p����� ��燆��G#@����J�� I���N��*�a Gf�: ���u|NH $t����L���@�7uHr/� ���� fk��_U~8`�����WS�K�� �`�����(0/3�^�+DM��]�S��v F���T��2` �3<�9q* 4
��P[_���$�\*�H ���nMq�40�G��m�>$����o�H�����������Vv�� �� �]�d��Փ� �Z� !%���dB	�H Ԉ�F"\Dh~�������$}���� ,�^���5G�n���Q�D�0���xJ�Z��8
@�r�/��)4^��x7��� r�"!�x� P<)u
&I>Y ��r���=H� 19e}OSf�_�E�ld	��������\�^�T�|P���9������_$�,?nЀ��^T���  
sǇg⍗�H��p*T~ �Ád��mJ��'%�� � 	D� U�VYMw�)�q�@�SX?I�9' �-	|}{ZX�� *�mw�	�O�UX� �JH����� %��Z�܄
w���� �D�W�� � L�E/�+��h��U�3�G�i@^Q������+�k�sC l��xJ=� m�;]3n v��UEtI0����� Ą��	�����k�&�rǴ�I���a� ��׍�f ���:9 �E���ɗ� D��e0T+���6��� �3i��<GT|���#z |��eBUj �T���D[����@1l4>t ꩫ�}�x��J�w�g�,��0";puа`=<MH8l��#Z1i� )��C�o |]4�
h����5@:=�<�7��0K����x��s�� �!$R�q�@�>��p� "� 6�Dt� ��ާ��-��}��i�o�����]���k����y?tZ� ,?���u��a
�
 (��@�	S�\���+�t�k����
_�~P� E`Z�%u��v�P���� z�:x韅e�E��r �' ��/� =�?t������Й�s �bo.�e��?>2�"�� Q�f�1-�E�`W�����=����T W� �����%5 �k׺.~�Z_�W P�#G$u<!�/��` A�m�G +խf���T �9�UVj �5 1��q �EN:��� I<�$��{����`��%��pD^-0_��e�	�'���(��:~vGl�B��@i�H�C< �1�	Ȭ �A$�q� �m;�PE� I��bÜ	s���6��M+�K��� "U_v�d} �Q�jArI�$/�&� O+ڰR;^%�{�J�Lu�� �"2�fw|�H�D�.�z^�i �J��[�� `K���U7�HF�	w˼� D_�f'yK ���T> �Rb-斟: �ef@����Ԁ�?$Oz�N� ��_ 50�t��G /�)�Y��1� (W �#'0RE����� ]��X��v" ���_|�D0���4 ���U�t$Q3eod�@��Hq�J/GI+�!�l �<'sSw�>g8K�]" ��%�� �*f�ݙ�(;�J �Ж�����,�|X��K� �$J��`���	8C��1�c- B)	P�^ �"dDu�� ��$�B�� �tJI|KM�
L�� x=F?j�w H�d>�,�S�� B�R�";�1Z�� 2�^� ������ ����LJ4d���(��\�] hHy��"�|D����$�����A"D-;�S�E�� �K}[����\l��;Um�Y ~BJ�7b �9CK�(�Xa���U;d��s����� �#��=C� ∗b��1�F�!����}� #�[BV=�?x������L�� b3�^�zw���eQCĒ��,'t����^���3� ��t� �ذg%
/� 6P�_龠 �l���=�y $�6jO� �����W��z�[���V��I�p�� ��m)�u E(� U. D<���R T��?���b'U���VP�ֵTSpx_��a�<z�����;/������0���2f���'�  ��� tT&���_��0��$�g�~T�!�^2�,$B(�߅~us���v��_��R�� \J�t!� ��m%q����_�� �].�N���*	RD@�իj&�L 4���C}H>�� $��W�� �-�8!�s ���t|� �R������'cn(`�=â� rY\��0�{��� <p���%P洌$������@� ��	���" �=�JW&$d��~�瘥@�T�� �ɼ��鸞 )�t�b�x��?'x�CH�wz� |!�s��f����Yį�2L���C?'��bK���ݔ�@ϕ��O��� 	�1�� ���;��	Hw7� ��\	�c@W�N�YZ w��_�l0 #&�v. `�ШD�AH<0W�l���v: o-�D��(P�~@��T/d@%��� t#�?
K�~	�&��OǮ �9�^C�T_�i6��w��- s��0�{B SPōC� jb�v1�Ө gl�����G 	�祝%N� $j��F!t O�sHbwEϠ�Z%>U�D,���h���p��@���`�8�T� 	J� �F�?�. 9,�(`	�W ��נB�� 1Ё��]�p �?�C��G ��>��� �� `�J �)w�%�c� �h�0ls��C� #�@Ph�>�F�=�3����6iLלV�8�\D:T�<a�=O������].�д� u��\ ơD)�V�J g�Id��܈a<K�0y�
'�_� S��C��b�`yGNu�������C]��lb���R A��1�� BT	��� L�S����iP�� a{�Y	� 2�v
0G��a��H���H�
?BP���!��C/��� ����E����D@HO����G 4������	=a����Il$� H�ڠ��y; t
�eb "�8����Z ��,�ȧ� ط�N�@S*���R��� ����3>G 5ܡd 04?8�h�����(˝ ��.1� �Can ewA�d�9*:��Xð�P�PT�B X!,��?�ۋ\�@W� 
u�Ѡk� �'֞Τ����ظ��Ѧ~����vj/� x��� ��{���
 y���=���� Hd%�NW�'~1)G��P& �=���Em� �aܺLA  ��}�${��ݏ����"R ˀg_�:g�4�pC$!(,�0D4��Ђ� ��s�R�fF�q�g=6(}\t懫����E�j��-Ln��P��>�@4,���0ݣ_y	8ࡤ���o� ��!bk}� d )H�uZt�2���0 8 �2�W��� �&�,� �?��vRW�F14���z��O0��l��p ����P��a��T�K�������! �{�� Z$��,�K��X�L�|O ���jk/p}� lhD��?L�c������8k, +���	;� t4�l� �p%�73 "K�5�I��0_�@+�,AO?�����w��>_tu$ �=!�}��� ��E�Z� �Y���� ��b,�&x�?N[�¯Y6P� oS� Z�dw� ����]� �U��oЗ�3�b�@�f� ")g�hi�H�0�P��4a�� u�6Sg%j֑����w��c} ���� ����(��	s~������U e'57u_A Ӏ�P�O� �ïV�����@x7*J�A�i �d�������T �"W�D�ԕ���b�J��G е>̲�� �K=|��3 O��;X s
h��)e�RF���p`�0+�A丛�zO.�U ���`/ 0쓜���� �+�؋ �@�O�N �%1#_� h!�u��0�Z�A2F%!"1p�0�	�`j�� �,�%\���^_O@sc��M�� a���gWx$0^p �ۀw5 ������	�_r��	R�� j�e�1] +zI�����hBC����T� J�R�!�O� ,b/r���gy��)4D:��@!�� WZ�C��r�XJ�{a@��� Q(C��8� ޟ%dR�� �{�$ū �>�f��7� P�h���/� �W�Xk	&9 �'7���4ɱ$�d���y��I�2T�"�$�<��D���j V�a��zJ' H߾!�B��;�:_ �8�0��J �E�z턾� �y$"��]�����������E���W�dcrMv��k���� B��/G��	���� ���pB �X^t%ue�3} ���GZ\��t��8��=/~ W@�E��Aw��F� ��j��*� &�_�J�x�0ʥ����� R
�D�l�  dji"wyt ��~%��
�p.�İh��Mvu ��J{�#�X ��G F� ����A�����H�~��%G,JW� D������V��������OR�W�h[� Dô'�X.���-� "g���wT ��)���(� ��E�,X� ��Ph�<D��W藻�4���1S90
����HV�q������ ��[�Hv ^�l��a���`�� Z���K}g��@�t��� ��B)Ы�~� �� ����e����Up�� xH%@|��y1��Y�@2x  ��3��|H�>���kD$l�)x���ǲ�G�u`��CPV#��%�M 떮"u�+�5 Ѐ�;�w2�  ���?u� ��s#y*� �c�<�ͼ	��Ai)�G8J8Y+����_F�(`����Qz�p��8��R�0*@�������T�0�� \ˇ	���B�$Fi�`鸪'��-��N� ���I�Q�CB���4'�n ���A��~� I	�W�0%U �,ҋ}��c Nu�T�Jj nA�;�w %?���V�@��:+�� �$^�fjP �� ri>Rz S�W�!L� ����u�bJ��,O�L2!��. ����} ���K�H1��+@�;�XZ �m"�D����~�����>�l"��� �k��t}a��p ��:2�-i <����? ,�㟏�*) w;<��X��0S
2�  /��(�R�:Ǻ����B�]�z��V��!��^R'���f�� vt
ʚu �M9:�� �+'Ȕr�� V"7��TL (S��O�9D z!t%��p7l&��תh�@'\�w�����L$ u ��xh� �JX�(-܏��]R���� BЂ�s@�S��蒀�	�F�TD@�O��/(�C���:���w�@���� ɂ�GX	�� ��UD�)F�� �"��p��ʃ/}�`��`� u\B?��0�8z ��ׯ��p $�\�Z�%` ��G��R� ƙ��$� H���I0� f�6�,Y}+����$���|�q}�Y�	_��� ��E���R ��t1q5�� Y�)~��% ��C����� �A�<�)�$��= &�;��h `N��ϖ�� y�8�P�G�u� �����[�a ������p�v� Iw��5Ԟrj�������Z�]	@X*�IbP4K�^�Ǹ�M��0xG��_&���� l��~  Jb��R&K D���;} s�	�P� �O�!cCX �$�028�� ��,����u ���X@����.�ڤI�| s#'U�>^� *��k ϡ�CZ{P�+T`M��7� ]j��H�� ���(IH��Ci j$��P<�����ø� ��1����͠�s���@&#��E�
I�T�8��N��+8�}�Z����=�,��`*� ��i�޸2N ׂO��<$�P���*�[G�"^�J�:�)�����ݶ� M�H�$�# ���P� �Z�[�z�ͶA���.�*W #��7� Ц�%���:�@�(}\� k�Bv�������ر� K@�Ń2O!"u~I@��F��� �
�	��Z�t� ���+m� �L	�MQ5�wU������b �
�;��d� ��"XP*�� �\��t3`	�۱��؍�����@�YL�P%'�	t���N&Ҥ� �7MSsC�I��ϸƿe���`�y�=?�<{�΄� ��]�n� p@�!Z�)'\GP��� ���*�"� ��`B�U�)>���s%� �ӕz�S�J �D�"�� *$�!� F�i�:BJt 3Ku>�q 7=[N]�� �Z%I�� ��m�o���0 2�����$ 題�)Ouo�gRi��=�(� �G�!��} �t �M��d�% .r)�PI �]��VtM'���Jw Puc�"��W ��Ζo ���p�k�Q u^��<�)�:�U�����LXy ���f�R�� b���j��=�꺐 �+���B� ���Lug
�3b�]�HJ 1iF^lX=L> ��(%��� �6�BL� V��dX|Z� �KP{�TF oM u'��>���������!�+����� 310�u}`��CQ�y Vb��S� �;�
�,�m u�}� .�xI%� h�Ћ���a �����DOp������K 2��� ���	uf�!H��(��9���=�v8 
�p<�Bh* ΃P~�uS �����Z�_ ^�|=	�� ���f� g`;E�t y����!��U�!��(�E ���3� C0�;:F5�t 
6�	9���J�fO`� �T�S��2
:�E� Ǯ�[�!��� Gy/�jeW Y���%�G�)��U@�� f�}�@rv ���̝�b)�
T��.]u� ��X��u �� j
�NLq�:Ä ����}�/�P�V�9�OW =��u�B�})m
�P� �>,U�Xﳍ�!�q����b���о���A��� $O���C��(�� Ǥ����4� M��J7��BI2@���K�� F>U3A0���H�
s�:�#W��pJR�� <��9�1� ǝ|sZ��C���,S H��ҁ�<8u '�Q��5KN��Fx;[E�{N�uRc:M� �t�5.D�Ă����Xu?�� ����� jECSh)��<ɉ�8�p�_�,��l ���È� C��g�=�\z�з�y�
��[	h��K��]�K�����@�X�)�S4�W�ă; �d��E �s�⓯�� �����S �� b�v{Y{������Cj��� Q'���xE� +z�����'{� �.(�� �2��_Y ��r���� ����d1,=��Y��0��Í� �2�X�'q �d)�7o� C�S$R����;�(�a ���S@����l����O��
��2)�' ��o/s+�3'j�� P������iT���&
��.d�P�=���[;u� ׀{���< 	?3�Dq:LA� u%V� mv���K j˂���u �
Q$~ �)�Ǟ��	� d+���ʧO��@��cCn h�B;�taw0 �'�_٩ �d@H��:J8G��~Ce�b��z� �f��<<�B����`�px�i%����p���b��� o\�[�� ��>�#N� 3&!\��M �������=��>���.�`��ص V�|'�Y$?�0�(��f5!,�iqny�'�%�gu�~� �e�ГT,�� 3=��g8�߳�����| *��x�K��~�Y�V���� ϴ��$�/ �4����y���r��� �c���� ����7.8� �?$WjhM��@<ƧU- /%��j�� ����a���M�[e����KT+��]|Y��/�H � ޞHx%M�QS��n�	��tL*� #�Uq����+/GӉ��G ̉07�Du� 8�V�Y�;]�>�T �����68}��Q� �z��@اB��� ��G��kޚ �{@��φ  ���N�8F��>(��� 퓎GŶ�< ��ΰfk=o �5�|�b G�%�U�'� �?�=�h + �sV �6=k� (�PM��=��(�� ����K� �d�6<"+�	��|hx&��-x`���k	 ��L ~뽝��ғ��$��� �e)(Rk�-Hp�C� ���2�T!� f�N+�x\ )Q8D�� �ŖC, I�l9�� �O�Q�@�� '$y���b�U� ��*�#���$� 2��  �v�p��`�|���^�~���Kܮ� (�����k��C��ų �: +�<�0!��Л�@��4�� ���y8!� oP�S�21. �!��� PW4�	�R (E����7 _b��:B�� lu�$��q ~	�,YN%t�Th����5$�"��� ��])�s_
���A�=+B�@�aY2,�L���_���P ��f[�S��}��-|�`�� ��O�:CKuz)���$��)G�{PC��3&_���A��;1!Jd$b CN��� ��sU��j� I��+���5u, ��	8�U�$�>;� rMs'��ޯ��f�~�i ��UBV��-؄���R��׊�����W��^L�5 ��Zg��#�pK=Ft���:I���2䰮� �m蓹8�<t����=�x> (w���P ���9;k��v��Q��J ��	��!�v�'��U ��Z ^[��d������E����a �#�{�
�}K�I"���؝ 7s�[�wُ 	�V@Ƙw�C�F��i �n]+@ ��>f%W`7�:��_U� p3Ҩ�� ����qR�=X��B��\<�Ɏ� �zGc!-V�d�� ���6�?��ߙ�_��^�� �PJt�8 (�7��
'���s@�U��(r� $F��D�i��E���I ��5��Lq L�}<	�� d�J�vm� #�����~��d�����@��t�����<���$ �ĐgP��L ܄)��� ��l�,!� ��j�_	�2R NXU�n��`Că*$�X�PR�&�� J��t�	� �ShR����~� *�4��{�:�`�<�a�,|�#N�ˇOd �{��� ���js�8	r ؚ��p�Bp� �g�4c\G�% �]i�jM�L��`R/�: ��Է��4�� ְ����4 q�D�3o���˻ =��`-E6|� c��%�#� �V�����/ C��KDk��ǖ�0ַ �b�q^
�z d����� I���/�t\�P]�p��� R_z�yBH* @��U��a�c�?%�" Å�uًb� �	U{�%�l ��W*u7� �:��X�,Ď�r ���
���$,0C�=��I����֣� Ff碑-( ���@+�;U
Gsz� ,=�*S׀�RdJ<jN�m8Ms��)0��2�"_ ��2�Āct�%ؔ� 54�H�I�?����Vrz�)���P�����
J �x5�,�!y&�	���̚�|M�g�3��]K�� ۔�H���{	�Jw�].0X@�HU"�V�BY�?��~,�;) �J��/n �L`���� D=0Tޘ_� ��%��a �<p��! ���̐��E�)�� *�� P��qU�I@t)��B`�*��  �w�JH+ ��LZ�> �b~R� ��w׺�� �d�8^5�r� ��˹?(U>�R�|x(P�� ��׃� �$��]҂ ��Z��w� n�J��l���8� ��TQR �q�|B?�%�g� Ei� �Ar����Z= ��R�8@� y�x
*K �<�G�����Ev��k?� `�p��� 3�*�.�E����-��< �{��&��� �C�=�' �9�n�z|� ��	 o� ����+ ����πr���� �i�8W��x� 4��� ^	�~o� ��e�Lfh,���%7 ��.�uUP��,B�` ��
�� 9$�l� ۻ���	"�(���p�2=���!�?S� pQV��*����ky�1�	��t9x7�<�a��p#Buz6� FI��� }Z�s�:U�u���� )؉��'r �����[^ Y>����'4W��Ғ�q�xFHQ�z��N� ���;6i ٛd��}�hp� �NJ/����"g���,��;��n��� ۱��C��J� ���H�p�9��<BE��Y�p[$�f6"�p�7���͑���� ��$��h� �*O�q�'� p
�Y�N�0�"e��6Q��#u ��O�iA�~��I�P�o�9` �)���� 6\_��7���� ��68vl� ��bu�0�0$Z�� ���\�P\�	�Z �р#5�g�� ��WR��|>�x P�4.�� (_�a
`c� >��Np^� 9?A�<�6� �V5q$lE���ς���� kC`!�?���2Y �"�r�\ �@=;��� �d����-�2�6��_� =��
挳[���7����� B��@�^ ��/U!3�S	P � �0��u�:t u[I�m 5���~;�~/� �ܻ��� v�jʫ`W�F�dK�.S�������j{�+��:] �G;�	�ϓ@`�9�|J>�� �HP��p Cm<M�Ñ ������� *�9�\��1E@���Շ�A��ܘs �-Xj��_� ǳQ��LD� '�qsv�t$>�AK�B �_ߓ{ �'$b���w���O� � ��6N ç֏T^� �\��yϤH ��BS���
V�>ةw� ������}�/�R!�+�Q��&� u�F �j��8c� =Gk�0g�~ fQ��_�聳���EyPF�� ���9 !����v�����;>�0 �t$�B !����Ib����]��}o�? �p.�#� �ZJ-1�7��}���u#�4�(�׶� �Lj)��89� �a'Eg< �S8TJp �L!�.����{��]\t���� ��Y�R�y��d�U�]L ����,��^.ʉ#�qb�W �΂Ԅ�`�����XM��K u����Q�p� L~�D}��� ڧ�+Q�� ��T�M� �k2���-\�(��3�{�/��H�ٴ��\R> mP{Չ�: �քuQ����=2�X�S��K�!�t5�㲰� ®��j�! s��P�� ��h�D �R���,��uS_��M9?&G g�W	�O �wY𫭅� pbKt&(�)�GD/��\-�fx*t ��I���(�`�u���� �g�WN�$��"a�
6	<� ���S%���v�o �pu���iR �tž�&25 1��Q�+ �T��*u ��ڠ��x �#� H����f,�'%�`�� � (J5�hwb $U�G)�<�R'V&@<��v M� ��\� ��E.�9ɀ$����Kٓd�p�b2<D�O��K�T�Ph,i�E�S��ˠxLT��8����1��^k#œ(BG�!�`E�� 㜓�x85; �P���7 60� �h� ��_��oT F�b���� "����dwt K��*Z1
~� �/�X -К&���( �?����Hd�@�'��: ���6�] ��@# (*�2+Bb",�eܙ@
�r�o'��bi�vy� �;H0u	�����(��4�jI�f��	�3\l�v)h �J��4�6��7U=/@�_W�8^���Q����&� Ǻ���i� ^��v89*� ����� O�Ar#�z H]��<�6�39� �dh0m�vN1��n�� ٩ 80���$4��3�! 
'����l�.��� ��^�q �������/��!�	Bx9+���-��Fj UWH
��@�wT�Y��+�� M��P�k��� )���p9�}��	����N@�;�%� �t'��kp9�xz�C@���J˃��dj �U hqK����8 �0'�j�D�V��a�1 �A)hX�BC #Lg(:��Z� +d�	�k�PI耝���]�Ӂ)����� O9�&DZ� ����PC	 *����,�� ��.)���= @�%��1O HX@ha�[P&����(V@8� �X�th  \�����?� K�+z�6o ێUt�� �&ݹ� �\���c?Q+���&� ��%���>)5��Լ�� �n��c/� ���$�4\L�� �8��J�K #^<u��IMqL3������^]ꀖ�crX�,� �t���)�� }�ʫ� S���2X�U`\��,�83m�<ˮ Ҏ^ ax{	���|�:� �������
Q�J5UÖ� q���h> �mO���8� ����C�0��^o�� �w-�"�WP@_�8�O� Ѩ)e? ���m���{� C~Xߓ8. f�gU�G����(��@���zP�����nɩ��.� �}����#����i�v�_xq�l���*0���:<��ut�yXj_�������-���� �4TN$ R�d?k9�@�	( �ɪ�����pI� �\�J�o����x�y�^��=>V mr�3�)�onÔU� ������ ��vmB�Ą� U<� p8� ��>i]�D ��������� Ea� ьl8z-��� K|wd5��y�� �x�$��Ɇ `%���r�&pX VC�F� ���DG5�L�1�)�^�N��d�#4HB�8Ϡ�0���_E��Ԧ� �e��dP��yȉ�c���١�BQ N�'�c�?�� 0|���q .��/�r(�)u�y��O`��?;�ev��N%� W���Ӝ oKwF�6�� �d�\
 p^D���:>��T�,�W��[!����J� 6��y��H�K:��p�/�+#���! Zjedʠ=����&�H�' ������p�� ���SF� Q%IE��Vx���M 	�  ~,����C�8�� ���O�}l k�,�63=4
�J��g�l��|�-7�"��
; 	0��>�=�`��yz��O�	�J��3���`�e �"������o {�ˋ�Um�(�5�ZNQxא��h�$H�{�8�&- c<I
?�n� �4�R	�b�@�{�;�U�!i`d��A� }�a� ��	!�\ ��"� ,�;����{ݩ�ߴs�R�%g �d8�а���X#�is蛖� u5���Y�3Ҁ��6��� �=�j#E x���t�����0CYd�Z+�m�;��h�����HlNY��\��[ �mD�|�� �dM��� T1��h��_�/u��v��2i�h6��nT& >`+�I �W=�7\#w �vX2QR5A�6��*�{� 0�O`���� PQ#�l�V� 8
�-CG�8=�� (08@P`p����,�9�� '�����q�N	�
�O���S�4�Q��V���W9J r5S����X� @�\D��n�N l������z����0/��;�s Ұ�xr�' +�R �� �%p��x� c��>^Y�3JD���������A���+ �,��f �� UV��W�E:�.�� ;�,����ì#��%  v��:8�\�(C�� @;ŉr �at$ (��Dh3>b���I�>v �*�j('>��4,�����H��� �8���x6 0~`}]< �'��^S@ �$l|M%�uyD�\��㘕�}��p% >+���Q��ӵl��9f��?���� ������� �OQJ?�@I��c�	�R�̘ ��FV�� *��2�[�&si K�#��v;�F� 6�Y�(" �N��
`�� h�H�;m7.�!G�8��A��r ����Q�$fW�� ��r0� Њ'A��� ����1���Uf2P�̠� ��o�1}sH��Ч'�;fL$+}� D(%��M\"Hd$�)N㋁��ߊ .x�;!F,s
� (Ғ ���0^��|d ��D�8�:�� <./Ty���
� [�q3��_��mC �D��-�� ~`�Yõ V6D��@�h$t� ���� �*�
� �y���	:r���OPP0h��� |����jv�\�v�@0Y� ��`k@N ��[��A�� )1'W�vB�k�� W~p�FTH��QDA����PT��X��` �\SA�ʪ��t_�'��b,�;�) �k�jz ���W��Q �6VSjX�4u Ɉ��� ��r�(��uxT���������P���l 1�	��hRvQç��� 4$F� `u?(j�Y ��0�~N�"8�� }R�L4#H��M_���e6��j(-�~W2 w8ơ�$�FH�q��B<�w �\�8�K R��(�$)W�P"��|3qQHF������d0f����+� u5`�)�$?��e�����n���@ANu��CT�%Jd ܐ^��h	D����]�� ��Q�7�W�� �e�5( �CRyN�h�t=�s 0ۈ��A �(#��� 5ЏO�YA-� ��L�� �&�.(�Z �@�!��� 3�PM�%N v�	����# �r2, �� �Z����=V�N�{�ο�@, ������g����mR�J�z���� ��aw+D�?���-���hX9v��l��K�{t ���rq����o�D Zf1�.�x�$k&,\�� :'J1������S�W� ���8sj�y=�+ �����F�͇C�$��Gn�R ���[����  ����F: ����Z� ��V%��P� � �s�� ��ж\0� X�ʔ��� Ȓ`����X���ݎBP%��A��8;\s���`��� P�~�${!��-0� ���P�0 ;n(�&�� �:,�8��r ���(RO�,:�BDǌh�G @s� r�(�����>��c-� eKL#�Dl+u!�8 ���4B���
C�����
���+2�߮ ��%X^8�(�	\[@�Z�0bte"D ��g��ap��n�!xF���	���Ŀ��l��� d��"� 0������I	(��z9tA���,O��sN �W�p�\ �"<XL�0Pz0]�  �^Dh�lbi�N�1�8 C�<�q"�qD�d>EB,�o |:�g>@�h��#�bvx�'�Dt.�D�h@$X��P�t^ �]g��fȩi>b" l�k6m1� �of� ��*Ԏ�@��ʱ�L3�� �0AB�)�h`�����"d��ߜ�@�0� p�h8"��`�@�z�������ѫ�!x��H��X"�������t��(�=pσ@����� �hz#�c���?�ؘ�`eڸL���$@V��U������4>3s
Q\,� �Dd̉��H�G�I�1�Z�Y3L��fQ
����,�$����|L"$�a�,b�@��4P�ͷ:1��@�,`�x�4�$�<P: b�꭬	�>��,�D�hHp�$@� �x�$�T� ���  �Y+1�M )&t�@�O�����2 ���@ �ƌ1 !�$2�pH Runtime  �r�o�ڃ~a �0;�@QE ��1234586789 YCDEFW  �U
�N�� ,]��\D`��'�E �N�<�
)z��Top C�c0�	�=ˤ�L \&%.*d� �.,���<�XDnsT\��oloto|������$�߬ߴּ�;����������� eD�$��O4�<\+� ��� rd9ej�+ �h���0 ib�8<j�G �#술k�X l1��m�CČFn�g���b8o�&?�T��GHJK��MN�ع STWXZV@ �AEIO� bcdf
ghjk� npqrst�w xzv aeio#P�"`�l�Dx�/�B �7q�� ����0�[�	V9� FY��?8��>^������[���1$��}Ut]�r���쀧 ܛ��7� ip�G�� Ɲ�̡$po ,�-��tJ���\ڈ�vR�Q>�m�1�Ȁ'� �Y��?��G ���Qc� g)@�
�'p8 !.�m,MPz��$s
$ ��jv.���r� �迢Kf �p�`£Ql����$��օ5�p�j��H��&l LwH'�8��
4��J�� NOʜ [�o.h� �tpc�x䠐�ǌ������lP�����xq>�h�d8A1�\$m��i�� ����� 󐄏 ��	?��I�? D8T�l�$�H$�"��@(��\$tH ���g! 	+A��� �� �!�]�6 ��N�� ޸b�	|��d
���CBrH����i��j��E}	Z� �Q֏ U���9[0�8��`�?p ��S��� 	xd� �DL���@��	T����Ʀ�?  |�E�-� ��V�K h�x�	 �"�D���� �$�H����<	!&2�PL��LX��C
ҒY�x�}|E�ڸ���4F��J`QK ��H��� 	�M�LP�@vR,T"�D+�� �?�|6� oW��%���w���	X$	
 $ �V ���(	�@�8 ]H�T�� 1��"� 'd� t�s� ,��� �HoV �9��x���4�r��A����/���M:�b��h��D�� �c'�b�|���$e3�)8��I��1���c<@����3� 8)�b� h$|9��F 6P��Yf���'e��a�8A���y�8ud ��Q��a�Z���iL)��v��� 9�� O&�A.f !E��1���bh��A�&�(� l���i3� $x!֡��� �t2,Q�&�1>(�Z6�!- �b��F�Hf��1Z�:|)d�ܓ 0<X9yl�1L�h�߼Z��� E�Ħ��! e�i�%�<�t�@�Ѥ��f&ġX R� �T��@��ډ�� f<Q�AT�� �!��͙��	m`1� �cl\�<e��3q!�2 �.t&�Em� ,�$����0>�D T�	�a4�8���(%Ы؜��p��fY�U�Х �($!Sz ��& V��>:'��z�>�
(&#�=�H$��)�`<-��#�裘�oP0��LH��\�q�I`j2L	d �H���"$�D����%��0�<~H~Zl$~ǐ����������� :&H(�4�PDbr�~%���������&x	� .O�AHe\�l2�$�c������ %�1 (&}" 4D>J�Vd*@���?�ҿ�� )�$ �>	J^ZIjH �"�D�����ڏ� *�,"HBXh�v�Z��������`c+���F�Z�p����$�H������y@,Љ0>�N-H`xhe��������F,-qR3�.0�Z��t�^Ǣ\q2~�H�J.d���6��\Dn����$���Ơ��@/	�(XO HT�h"pD�������Q�P.��GL" hdv	�H��z�P���$�֨ $�J�4`���n�l32ν�}G�tCu r=�n�Tha9dI�fD�F0 �Cri��ca �S��on zeDv+pm E~�J�I�x' $Rz5�V�r �u7"F�8QA��oc㫠�-L*Q��y��Wi d�h}aTo Mul�:ByQ 4]�.!0-�st�A�n0c p}y�{�z��i0��/�ExI���e 7��GS/ u�(p�fo}A �Pr>�d� Rsi6�Mo� �Han� A�0FiN�m ��Z�M��A�Er��ȓ��m�G�J5���� �,d}�� �j�C�2s �T�}���� IW�S�aUnhM��dF<p���3 �tS(&5Po� vE�\Of 7=R��w ������W�Rp�b��	p{C -S�zENy �mTi����$� C�z8�� )ԩI�ur 6��Kdyb�z��ML:�j��
ng���=;auBoxH���N�ltyv�pRi�&�&g \dV��� �)O4�n�� �!��#�0�
ht@Sjp��Ã���fY:o0�I�d�(4�^!�aeҚD�.���59'�-�k�T4��5΀]G6�d��|����/@i�>��b�U �%V&v� ��um��L �;�H�3�� 
�of��(�]b|� ��.kr^��\ ȫ5S�� �<vDT�o ��y>4�]P ���e�a; ��q&)y{ZEug�\���ƛ ��IsBPRo��S��G��b��Ø��ꠔL>�TLT:)4.W���w;s D�r����1 V�6�ɹ� ӡyAMC� sI�J=x# 4Ҏ��T�;pP5@h��NQ^ (��6����E��@��w��D��#	{�] Bk�� pac�$�� &A��֯+�IE��C�'K�B��xA<{R %�]�?�, ���DUV �Y-���� C�;ڤ�E?,'��9zv$Ce�02t�?l{�r[*�Bk� �!��i�, H�vlu�)����qA#�`;��0=�� ��,gJd-]�R��D IQB� �p� -��T@�ns��C���>p�=yY ���HT�, �S�P�': �AduXD lgIU	/�% ��ipq#$��R&j~�eA�57 -(X>iȟ��j} ��tB'�� �rR��_�psT�ڃIc��� ��s���j D����i��bW��R"�!6�Z4�ِ�ch ��9��G$�HB� Y �tk	�p��C0A �z�=�� D�V�gU�R��L � ��M8Y�}�t$�~Ғ?J3xӔ�FPZ �pLA���� oy]Q� fu ����e^�&,n�: �t����� �H0G��_d :J8�w� �k�*��4 $ep@WSA�^ ��lBj0J����$��f!��th�3?pH.\a� }m��v\`��R�$."� �Wn{;hu��s��Q2y��+�����p�Ln 0',G 8g<�@�D�H�L�PT�bj�rz�����������������ʟҟڟ�����1
���"�*�2�:�B�JR�Zb�jr�z����������������������2r tvx&z/|P~XN���4� ��5.'� G�a)6]�i ф�7f8 ���ʞ�ݟ��@��9 '%O��B~HV\d�v����������ßɟ�����:'G0g6�>�H�T_ڋ裢ʐ��" ;8ɇѧ�� ��<r�=�6�?�S�\c�r�yÛ����>ږ��a?� ,�5�z������%� ��ID � �(0rBt lvux�z�|�~������I�4?�����  1&N8�P �\dI{$ ���F 2
�<`�~������� 3
'G g)�z��Ǒ盓�����õӼ���m 4�ɳѿ�� �!5r't/v RxjI�8?����� �7�NΎ� ��8�C�:� �%;5�K�i ������ �o9=�:� >*N^��� ��?'O GXg���"�0� 
���� �C1;��� ϰ#3K�i�꧆�n�`��4[ 'nG�g���	����'J�G�g���5 R�8C/×Ӝ����ȧ����B��
@Y�"�'�I@W�_�d9�v:�;� ���97F9w;�@(���4� 
5gNv��� 7$�k��` :���u<�� ��=MN Ğ��Ϸ�Oޏ� �ʶ� Px$5�0Ƌ ����X1r� t�M�f:��3\4����6��̣ݳ���!�*�c��;�N� '�<gM�c<�&�}����������9�:�;�<�=�>�?� �����<
 ���(C��?�V�^�f�n�v�~ӆ��� U�&@=Z?�vDxRMXT��������������1�<> >/�;�H�Z�b�|#4v���N����G� ���� ?r
tv x"z*|2~:�B�J�R�Z�b�jMr�?�'�G�g�����ǲ���������������$��D`�0���� "�*�2�'i�c� s�&��c2o$|�@$��9��:�;�<�=�>�?�?�?�`93�B��<$=,>��~ND�LgT��Od�l�t�|τo����Ϥ��&���r�t�v�xܐFX�:�4�aGNg���<�D�L�T� L�:l?t=|0^�O���Ϥ�n���M$�H9~ 5N��$,_�:�K W&d��|��Oj�ɸ�@a~���0���Ӳ�����6�4>�<�@�D�H��P��;XJ��z|�f�Ӡ�f�۰�Q��L������70������~DNL��T��\�`�d�h�l�|�Ҥ'�����ҶĀ�c�t8 ������ �$�4�T�\�`�d�h�l�p�t�x�|����������dĲ~�~�~�$��cA���� �$�(',G@g`�h�$R�	&x('-��T��$���ȹ$Ч��O�����|:.'2�e (�,�n4�8�h�p�t�x�|Àӄ����������������������������; N$�(�,0I4A�<�@�T�z;2d��H:���Y��?�N؎���������	 <,�8�@�D�H�L�P�{l���$d�o�Ĕ�.<�����= �� @L� �P�Tɪ\9�`:d*h�T������������������, �>N��K���4X�t\v`xdzh|l~p~t~x~|~�~�J�-����������@'��p9?%�R �$�(�X0�4�Y�������pT�dP��ðfH2U�5 ^8�9����������:�
�������"�9;�\��=��(�2� �3���딤Րé�0œ�@�1{ 3b4�N�L5S �6�� τ 7u�l�����r���=���sk=�%�1���������8��S9 w:�&�\
� '�<;2� ~��I��) �A�qم� (=.IB'Tv ÁX>���Н 9��L�� ���N�E-�$��2� '�J�y�*3F��`찖� �4*�ƃ ����Ƞ 5�ɈѼ� ����6r((K�� �N��8� ���"9O�T�n������	:/�K��&�����B���.�$`� ^��i4Y( �<=�>�&�<�π�ԃ�F�
WH�� #t@vIR��9 � �&:�;� <�1����A�T�lǈ�r�t�v� ��2+�?��٩�It��� �a94s:�; �<�/5[N�����	�$x �t��2�A�K�0~V'[Gaef��s�yZ��Ϗ�����ş�ڇ���6�� 7t.�&�U�^�g����X�
98(:�-�0�Lɴ ��R=%��<7�E�`�i�������'�G�g�	��r6 N�Wk��$�ԝ܀��X�� N�VkIs �ȝ�^?~��<���=�>�$�Ƴ�@���0�r[T��O���\ � �(cb-4�fX�\�`�d�h.�6RQ���tX����� ��O���ϰ��������ȟ̟П؀���AZ�9�� ���1��< �� �$�,	�0hjH�-HpT�r�x��~rt xY�P?�$���r�t�Z�X�O�����D�~�J�%����� ����Ē�� �(�,��8�@�D�L-ٶ�h�p�t�̮ ��X�~�K�#��=V �bvx�.Z�x���A,�ɵ���� ��5r 7JS�9�:���p��9�,�� ���� O�����d <rtH%; XaI�&O��rctmvwx�z�|���V���ۗ �W����#=G�OO``lK�� ���?��� ����"� � aXw1�% `rG92n! 3�NՀ#4I 5�z7s ����� ��8_9;r �ik�4�a=�Y�$9> 3:�'!�x
�dԡ���*0�<+1qL��-93�:�@d4�C5 f�����vr�X�. 6-'�D9� �x����	���3�wO:�/��@,�;R<W=j>oЎğr�t��8:P'�G�e ���;"�d, $�*�� <.'sGxg� ������Z Qb�I>� �i����5���0/��� %'1u�����2>�M��H� �3w����U �N�i��� �,'^G�d? �`b�.8x��� K�'"����Ǔ(נ���> � ݎ�8D�X���q�Ȉ��'B� ����Jt ����?փ�%��8�<O|D�H�L�P�T%��9�l,��,4?�Ȝ!���	n0� @P*1rWt� v�JLs�	w��?�3p/ �AkP��$�����A:r,;�^@&���"�P�����XrF t��7����������txsf*��@�;G��Cu��&��� W�[c.���g�k�o�s�w�{���������������钣����������(�\:� �9/
z �ӤA�E�I�~.�`�N�걊 ��&��v X]\�>d'h �p�t��|�i��8�'� �"=&�*,j Xy$�N9	��h���%������KP8�� �b�a��h� ���6N �A��( �%$�T�0 ��8��GH�yhO� 2���t�AԔ	h���j�t����P�~��*�$ 5>-@�H���p�t��a�h�O�(Z� �����(�,�0�I�S@WDqH����:��,M x�?KZ .�eA�,N3JLH`j�n�~ 0P|!w7{����ہ8����� F~N�� �����C:������;,L.�����@ß������ �=�J ��O Z�m��N��� �/>E�M�o �{���7 �L������̇[ 0� 1�2J��� `%3M� ��Ϛ��4ưVo��k6 ������AR �;W4y �`�iV��J9�L�OF� ��.&��:�*;nI�P�x�N�	V� ���C;= sTj��>.N�@����c� �p���Ie ��y1Z2r^\t� �x�z�K���_�@Z�4E5 �'�G�g� ������
097��x z|�MO� �c9g�k�� x�z�>:B��C����Դ�9Ҿ IJ���m`�?9-̀рѼ �0�$I�� %T��`�
3� Sv_ ��肌4��D �����Q 6U'�G�g��8���<���Y�(��� rSt�J7���V���"��� B�����=��8��F��J%���6?r].��K W�4Zv%>��p �1�N�� ����O���2p,�>�.� �j���� �rJ*	��;,�ר���� �;0e8��>@��H�-Ps�X��%`A�hR�p��Jx ����ذ�f.�����l5��\�ب���A�`�N��P� [�5I{ �xz |@~rH>L[�*X�\�`-�
��x0���BZ ���˘� \���T9K���� �$��@ �3;4G��f� %aZ�+
XĦ~�(�0�T8�<��D���6ι 2�?c
��j<�( �.�T^]+B:u@��P�2$9��ޠz:����[� �=�A��ɩ/:���R�M ��B�!0����1� hȸ1y�H�>.	� 5{'�G�d�Җ�T��� b�����4t�v�x�z�|�2;O�w�(�	 )ထ�'/ �a�~�(z�|�O�#N0� B�ac�Ű(�������/�0�pħ ��1��X5~:&�� �����v��/�4���Ì�~t#HY  /OhGz g������� �
P0N�� ���_Xptx I�%�a��>� d��#X �;N<l=�xy�͏3�u�z���� Q=�t��I ����J(
y���"��T4�0`r|q[v^B1G��_�x��|�~�N܃�Q��0�3 Zk8��[��hD���A0�(&	:f'pAa;6,�J� �PrHY{\-���`X?Ɛ� ,��_��7{��� F�f�B 3[q�>Hu��7�\���D�F��§a��������* 2p U �]�TZ{�
 ���'��r�t�v�s� :F.	��'
����vG���<�+|�DA�\8V��L�92���P*�����?7�H����<>x�:��1sI��J����&쾆?	�X��Ϯ��J �R8A��x
�`:O*ȖH���ߒ�� �P �x�zɡ�@�) |�LR;�<��t >�\ �H zi!d�f� �N��6� �梴V�e�:�R�@�/m 6<"�=r�p�>}���px( ��@0��| x-X���E� ���2v���c ��,c \�+�T�n$x�tO#Z	̰ἔ��d�R�Lu:�l��Ԁ��X\J��D4�YI N&$@��9 =5%K�:�l>�	?AvX�̻O у��'t��s x�z�|�O�	����]�dp%@�*0�� 3
5��^k �w����B���΀fN2ot� �����4ߜ���q�0�D�� 6��	8�$.;>
��9���r����G�g�K� �+�=! 0'GHg�} �M�҄��d-����`��������������5 �	�a��7r>t����@�=�9��KŔ��(>T�m
��H�v�C���'�"���
0?%� �,1�p����&SˇP3A$c ���p:t�v �x�z�Z*���g��� ��ȸ%�;$�:;�' �a1y� G����8����9:,Mȓe�����;{ <�=�>�?�>)H�p v5[98�Q�U��~]'a�e��� �/=9>:!;%<)�-�1?5�9pr@ X��0T�a �j�� � X�J$	�,=E�v �]�^ �R!��)�r- 1�~9N=�4E�IS ;����y >ܑ�"< t2��V3� !�5���=l ��9���H r�%e�ֱ�U.�B>`�� �x��0�3 �4�7X&�	>α zHT- 1A�/�9&P�Z.������4> ��A6%ɹ$���9<Z:��J.AR� �ۃ�"x d�23#��  �)���g� �i6m�q�u /	�}�HK���a7D�b�:S� p�˲���/ �K?X�JN�(��"�>	9a�rяk��yY .`�-b��C�0VF��Z�WP� �ve� �L/�aR�� �D��n'>� p(�������93���%u�� ���A�4��+�?�a�������>E1�m�C ������� ��6>�Q:r�	��v�lh$/7e I�_ψ �K�Ph^o�������-�AD���N��:jN�#b�=�Gt .]��� �~'����> �:�"$ �CRq ��d��� ���֠�	9;& @�IOpi	��A� ?"��~��|� �t�<vx�N K��f�n�sÜӺ�P�L� �h�P8�Ґ`t	�� �i�q=V� ������@ ����j[�RGKS��r. `��6ِ��\�b�j�X{P�Y�ƀ�:I.rN<�+��ª��� j�A�;~	Jk�rx���� D��XO�� H�<��#9? /%6�(Z� ���$Ԟ] 1n+�� ����rt! ^9�s��Ow� �Dp�]�f.\�� 5-$���� 6N�A ���#{	8+���7�=$�US@x�p�������~�?�7K*'�`@O	Їϋx8v� �˛�ް��*T����Ȩ N���2�>%��d}: �Q ��/VJ<�x$M��{A|,�%4��`���hZ?�:��%�	��ZP=�� �F:1;E< Y=m'�A� 4Ю�����%�����f����$����0.zt�y`4N����xr�1-��U^�}�������|�\��a|Uټ@�� ���6&I Hl$=�<�� ��K���I ��*�|r?� %��$��� '��L�]�n.�Nϡ@���A� �<�&|h'� �ӈ�����0��2�va�/�:]@eA�t �y86,�v� ǂ��~��9��/�@�� ���!� 2���#>�( 3��OC�&S� Ne�b|��{�Jȃ��P� �P_��*� @O`�h ��^p��x�,��܈���b u�z^	f� ��71.*X�� ONx�� ��%;����9:2�b4$wZ��/�t�y< 9'�A\| �*n�JΦ� P���.8j:u��V�଄����ZO���� ��Y��'mA :}{#�������=�X� ���3='GDF�܋/�a��tj�;֎�������ȝ?�N��25��иbr YJn	(|��7?t^�`߶��ג��W���D;q <�-���9 *�X�cz��O�T�� %:J�a~� 6�K�,t}]�('��Dh�}/�x ����=r� 
>�hK�Rv�k #�0��O�h��qBM �l9=:K;Y &gj���R ��%�� �&�v���&�-O ;}5�T  �ˠ$���*@�E���� �8fXh,;�xPq�<��bK�Ĉ���.v:7 �Fʷ� ԼD*��N% �0^x"J���9?�;ҀR9�'U�`��-;!T�d���*�	H"���_j��KBX�\V��_���@�>^����`?qNw ��ˋ��|� Y�`-�X��| <�L�(H+CH� JZ�؂�V�Il��&���:����QE4�j����Xw ����/4� A$�+	|�Y np:5rEtO JZ�T}Ҝ� �a���� 7r�t�v� 8�=�HV �zs��9 ^{��բ�I�%( Of-q� �|�/�aا9��&����� �<
�$ �")B�^� ?�G�QOc ˃¦A��r��Ѯk¿H�k �����l@�"x�z O.>'�B�ȕ����~a$��S P�N�(K4��o��}�r��/ʄV� �%5�a� tb,�L��N��8*	� l���7%$S�Pr�:#�9/�����*� ��>�� (F�S��l�~�����=��=��?�l���\��d���K^ �p�|�2 �v.�;�G �T�f�l�1 ^�n"`��b	G�� 8p�& x�(�l<b?�\�8��ZX�$�� �O��q 'ȿDF�PҎ��e�ޱA=<5��,LN� ��7:�?��9��s��� ):O��0� c�AD64����� ���C^ Q?u����� ��X�% O���1�9{ �}��J��	t�I���<?�'��b�=�R	{���A����x��a�y� z<Z�Ȩl��$�`ݘ$-�� �2rK+ �`3��H;� dC�GV� ���">9��jlZp��0&�*�.Ф?6�:�2s�w���<"����W�rĽ���b 23�"t  *�.���6PĶ�ٹ�N����[������;�;��L<�^/�a�����'�?+�* �;p�[ C��Ki�S� �/Ȥ" ��1��` ����[��n�P�~���_ �4����l3�@� R5¿d� ��9)/1�b�� ���>P ~[r�x�Qz (�K��`�R\~�~ ��)u� �<�*���"L�!O��ĜU F?���7 ! �9�:��r�JC�f�6ɞ��$�pHa��xz <��p������G���B~���I��Hc%��w� 4V����tr�萀Q��G� ce9�V'( �J|*���;�I@�`>��w �|P�[���xt�� a�0��71K��3Q�t u����<8#� ]B�=[*Lh��T�������W�`K�^��p~ �-���@X �|Z[i�y�������� �l�% �p�H�2~M �'Ca<\j>	�u ������� ��<'ż �TU�a�w�=���~/���W ~���VX:,�j�I.%@��'0�F�a���h�t쎨�:�;� �'�AT�/ �N&�6| BE��z���J�� M���8 _�¾�Ў| �[�$��� !%0I�1rJ)��M��:]�0 %|ؾ~�K���VNܴ ���J��^� u��� ͓� ��x
Y'0/��^��� �4.*V;'j����:� �����5�"�Q6����q� w������� �Z��&u� QC�N��e	TP�������,F @��/0 ��A�W�: l�w�ޏpnJ� Ѳ�O�F�@�o���,ti,�; ���V�9%�!X�T ��\-� 
W�d/� {��A�� :�0�|�;��$�B�m�� ��T�(��� ˿r����?�'�a@=$����r�B�P(��	���� /ȾD+	8W A~fJo�� ���0��T�V ��D�Wb e~*y��� ���ҥ���,����ם <�'A@/�o8�=�ܭ� ��$��a 0+"  i_���������1>"�
%�a�	/$�}^������@�Y�X		2T�9/�dSI�l;��a`��<p�>�{ ^��T:u��-;� &8�%Ga�`R��j|� զ��������c��(�, ��4�8Ӫ@�D]�V�o�pO�x�|V�Xx�ɐ�6�A$�z ����q`^����O <���$@�	��v��� ��~� �H�L�XT� /\��]� ��+D	H�sX I�?�-�� �tvx_ۼ��K �|I ޠ�䨯 \�ɴ�"�� q TL8$.J�M4|R�}�H���D��1@0W�>dX�:"�z�p+�F|��V ��&%�y( ��*��^,Db�B.�0�z����4��$�W<  JT�%l y����� �,'30X�v 8[H��o+�?�^�ʔ�+�~[�� L�v���� ����R%�JY��̫ �m��8�<H�<=d��X�_��b�	\��d������̔!���� �ˤX�Z�� `�W���hJ���4:�'Gg���.%<�2D�^L�P���]` �?h'lY.r�$g����-�� �,V/�D��d ?�-�A��,np���+�N�A�:�Z�o&� y�\�?dݒ l[+JN�|r~� �%�Y�D���� ����'���q�>����^,��� C1 $",�0u���*�����`�@��D��ېZ.��oM�D)��+�q���0���/.��>;w�0�'P�� �1}�`�����f�S-C�6yy(B�!WD}N��IjVjh��F߫8mLhB&u�:E*�S�t7��Q��A��#v��6P�W��Q���
�@<!c A8Ч�9	��T:�W�3,.�o ���U*��tz
��� Y���1�q��>��j�G�@�<F	�h��/P8H�Ua0�V��	P���PQ��8��� -uL��@	�>P��7�ç׏����|����U��?3 ��tx��} ����CI ��)�� ���vL����`9Xb�H�6��� ��w<�^S�P�������}�uz=���E���d�)��UK��+�t uA���F� �g]#m:L �t��TN� sѬ}ʭf� ����tX�XP=� �,/� ���y�uy~��9-F�� �ٞ�a
K�� `��@q�S����آ� � &u2S�) nMJǴ;A��FGf�z j�W��~ Q��A�� ���Y�b�-�u\� C�SV� e��P���g[uo�%*�W��9�e��+41B��*9I6�7S܎ u$Z�J�⸖	c|?w�f� ޡ#_�ZQ!���K��L �7�2��-J� 
���� �$��DeP�=H[�`/au�"�K� +Ó�X �QP���Vv��B%H0�!� '0۔J�d<=�Ѓ �_jL0�<F&� ��G,��<Q[ t)��24`P��� Ķ*h�� _㙰5�6� ��b�aE� G\S��4h� ��;5�� �� A��L�=�� 	p���OrY ZbX�n59͛ �V���.!<�����{�,̨:�m��"�Ƞ`� AYZ�_����
���*�0� f^{�����&/� �s�(=�t��= $��):��� ���|V���;�S����
(p�q `�~�3}�>A' �[�i�0�p6� f�- @�<g�5" Cч�}�� Z��e�<����Ҩ�DхC�2�L��n����	΀=�1�- �B���G2j�l���}�e]Z��4�d�9�1�
>���� ��&��� lR�����M ꕰ<�՟�j���B>��?-����LY�>�́d���u�e �����H��>����x��! �ڈ:'�� ���kvD ��<^!�,� H�g�A+���UC���"���@b��O9�|������� lL*�͵X7$30z�i� Q:s�� B ���Xg� ���(��\�7@~�c�p� HRn��h  js��k�� �%����B�!F&��t�K �|#%�/XC(P� �]�asYg���8p��R���h?�� �kjO�A� ^�1�� ��􃧂8" ZB]M�hyu�vQ ���� �\���Z�> :����$z	VhQx�@�@�� =����|� ��=��sT�*x?��C�ǰL�b d�N��=_8����F2n��# {m}��� DMʢ�6� �/�%嬸 a3i�,$�%�KO�U��`�4;�}��Ϻ���u���s�PJ3W�$�%�?����tW+��_Ž렅�;>r��߅(�h ɇ�V��+���^�X��\:*�+��1Y=�}�6s��AB@���:w���b��3���t���� ��{]�&s�<�a��y�C���s_l��׷Vi�tua�A�occF�e�cP�o��c�Exi�^�8s�Eu�C�M)ag�{ÉA�w�printfLO�DER ���The�p>du���|Boy �S�%s�c�uld��еb8M�a�8��k�y��m�c.� kb~r�uh�Qo�d,��+uC^���l�	�ElG�L�A���f�#(Mo�~l�c?}FcA'Lo߮�S�紳f������0 1]� ���0a      ݢI~�}vG�+=Eݦl-�;ԛ�g��ft!�
3�S*��� �n����<b_Q1)�P@�����=���uf��Nv��@�ʅ����X嬎0��b�ld޳�og��=��C{����;�ʇB�F���_�Ih"/�gS䵨p�J�}J��] m��������b�͐d�w�
0��n��2끶���sY��B�-I�a�d^�ة��RX����d�!e�#vi��y���ٍ�������-Z���1S�g-r�� ��l��k�cˡ�~ꡱ��_Ă����#˴�'�oc�� �	�W&`�㍉y��ى}����"LA.gj�,e��aL��Vp"<lkS��ns��ܱ�x��X8��{�$�7}7�Od^7�����!�V���}"�O�1��9���99ķ�KF�x��g�򠩊�<�_�͏�U�֌�[�U (�yI�!�*�|�a��qu4�PjY<ٿ�=���n|0���zBC��pq�0(h,n��&�\5�.�c�Y������<}gzg�����g4�x���Xa(O٨W�� ��|xT���O_�~q�(�7�������6/_3���1������v�[!�Yke�P�Q��Ɠ׷A����Au��U*�߰�;���� .���.�2�È�:�1 8���f�M�<�T�z#����nlx�α�VZ�I��i�ϵm��>t���Ai�ҵU
�$�7���y1(i�|�R���X��$��^v2�:#��4��3^�~٧"���%vĄ�����խ�5�/�qM�Z{f.��{�b/M�Ò��^���T5���D���wb��a9x@e���#P��.�F�gO�M�De�[���ݮ����4�O^�I ���sf����	�m��7�;�ą�h?���w �%����54xc{;�c.W�++�m�b�A'�d9�������s}�$ ��+�}+Xǡ�TR�����.~lO��HuҭnMj����bK�R	�ķ�4�ֹ����u�j^��:��"�#��V�fԧ�[�Jβ��
�� ;��2"�H��6d垎;{D�j)8K,��:�� �XO:ί6��Es�W��� l?��q�ƌ���S"x{�8�`t����`V)���k��?�V�5�\���@(9�����3	Ll�' ���Z�>�"�j� ��Ϩ/���@��@��}�fK	�.fѩ�D�]��8/�>�^:�(��1���mbo/Ϻג�Ɵ�V�h���^�����p�bY���:�us�g =3�SJF�g��8����>Y�8�G�o�ˑ;k�y���!:v�V��Ϯ���vW{�N}�5z�hQ���'v���TY�7C[���M/ܷ 	U	��fe��/iHT�=��(h<��������M��f�MS�#��C�⑬�!m�6g�Z�
�!�7�+�:�0y�f7����T��n��\���6������7��t����9_�t��i �nr� t)��\�����]�{����A2r�ȗ�>7���#ʞ�(�tn���<�i�:Z����cO�s�F��y�ޥН���!Ӹz �F3�kDޜ�i��$�C����v8�d��:����_��[*��xn�*�����۲\��Q%������� & �X��|�ho\���yAN��Y�N)%`(3P�[�U�US>��~��m�ϑF�قj[�-�[W`e5�\:pk��Oʯ���Q_c��Oi��5]�����0�d|�߿;鑣>�،�#�6�9�a������pt��xJ7҅~�/��1��hXa5�n���Տ�0g� �������v��o��K�s;�]�4����ߥ@hraXq��A�D����#����P ����'7�AA���$�Ǫ�JK��������
�B�>@%�4��G�,�=nE3�vs�T%f�9�(�(	P���������ۄR���/<�c��ʹ^2�jw���x0
�N?�K�Ss��)�E�����N؊c�F��z��w.�[W?#w�Ղ ���4��	�th�4��T|�٥'Ju��c�V�B�?X5���<t7���V�=�8T^|5�_���9��q=�4��0�'c�c�dmY@O1Yo�F�!�bl4am�'a����TN����G.��)�/R�M}� XcĹTkX��φ@f��� �0V8�ӑ&L�pY��Xehg����IS�O��Ct��'�λ�~���,�Յ�7�8�['waj^'�8�^�,Ra����M߳��/���M� �e<�׍�}�����2���� �2��:70?x���;�Ĥ��*�~�:/�@�t�e�%�N|��䀏��}�3����ucM�S:Gi���L�n"����Zn�#a��6c��;+�r�?Km��fn�m��o�".$*���L���!D ���05�O��7M����"w���|�! ���� �)��A��C;��$�^�����Lߛ�&�w����#�nR`9����3�X�x!?�~�P�� '���Z���j��������F�o�7�L,�{	=���@���yf��BQkp4�Xl�L��p��V��0b�r�N*߮B=[�u��V^�D�a��Ӯ[��e��uƪ>��/��
X�ヘ��rE^�'�؝�>c%�z+j��'�~��Z�ip�� ����V[)��-r��-[�6m��8Y9%kq)`.���io[����G�%E�Ӂ b�G�����'�0���ތhz
���D�+�[���K1t����]x�'Y����.�Ԍ���S@-�g�/�U̩�}R�Q�_	z���u'H��b����fKeg�Ŧ���w4g<>{�?F`~�<����9i�>7d�p�"l�[z.�j�V52һ!��:~���q,D��n4�u�g@���#����{�ʟ�n�F��'��Z:�o�Ʀ��y����[]o!dM�$\$W��:���� ����k�6��?�,w6(ǚ|4,���"�U�Y�oU�a,C�Їs7������sR��4�#C�����h2]��v�?ҭ�9Ɠ�$�	�A���#5� ˖��-��q¸L_Dw;������:Re��꫷0��T�[�i��@N��Uӯ��Y?���x�Us��1v��}ޚN����_r�u8b:C^%yŲ_��_�I`Ln��M/�ژ�qt8(d�|/0����%�6_#dt���s(��X�J��O���,S~��CLIt���̉ ����v����(��Ca���.~��(nV|�hL�$E���%纆�(��c'q��m����2��Kx|�Lۀ���w�y�^ ��kz��V�.�X (Kh��Z���P!:�6�C�O�����y1&R'il�5�;��S-,��Z>��`-N;�E'��on���M;�Y
����׼�a��_g�^ʢJB��Nr�$���&=g���ꧮ�� � g�N��w0x��mUA�E%Y�]��9�
��u�REѰ������q:�������q#
�l �'���Etϸ�G�7�a��[�X<iC�Ö��rĤ%m�z��1#��_�^v g����6�^��U]HX5|F���5�~���4�iHy�A�	!T�m���������O��j��>]�B4@rxCq�b�%i=����x=����>V)����R���/� P�?@���gY���M8�� h�V����#��ܙ[���*��gw�jO�^����ޓ%����{�mkI��U�Y�PQK蝦�����2��s��UqA�$5{���^�QD۩W�i��ICB��y�lf
�c���=�|+HQ%�ײO|=��1�!F��������*[�^1z���X�`�~AҠ
��D�hU��8H�0���3�ً�f^+F�����"V��,7���Kj����W��E��ǚ��1Vb�F��	 �e�T��2r���T���>fŨ{�~/��=�6K�,��0�f��-(%{� ��i�"nĂɲU�!��z�ﱮ�����C���8�Dֿ�)1���а����>�E�O�ܶleE�8xe�j�gL�I�Ɛ�6�{��rSU��/;DA��Ɉ���L��-��^ģ����ДN��+?�ɸ�:v�'}||���j~�����S���EX�Zx7l����SP�S�p�T�3`��)�>7�L�:P�9?��M�`98��h�q���\�	%�=����NQ�V��'�K'�>a�	]��?9!�+#�S:�n���:s�I�E����I��+���	�8���
��K�?B?X�Ao�Ǡ�P��G| �e�NC!**��9zhD���q��Xd�@,ډn`���N\��|e��I�1��ZqS\g�4z�����>+#�]��U�A��������|�{a�R����ˡ٦p���� ��h�����5��aR#_Zy�E�i�E�7����s=E�֤ЖS�,��PM��� 1��Ws���<t�Qӯ.�)pjx;&��E��a��hd��O�����f�]w�s��T�0��!��t��W;�n	�`�Fz>I ��)��yN��-$50AX�B�c8�i��/d�b�a!���|�3%����Wnt��`���e1>d�������]��]� �j�4@^N�� ϋu��������"=��av��4E��B��k,Z>�}��KS��P�f�C�*y��*X8|�Ø�Ԋ�" ZE�ZE���8�K�`���	�/����p��UO v��l1Ⳑ���W�=�N�K�}��&bI����x��֦U�O^ Xl�=R��Zp]C�L�1�Zj:��RƳ�d3����&F��h�;�����O~����z�<fH�rU|�E� ��2�7d:��xh�]�� ��!�����t$J�{�����o�=K^���Ŕ�´�َ?���cK|�d�U�3�ЮU65�n�*��ܣ�r�����"eL+A|[�N���3	'�a�-pR��2�ek鉑	d�j�<�!bǣ:�2kg�8���������PJ�5���h�f��T6+�D�)=��;��F�%;��d��y@2��P��
�s���l(�
�_偖cʨ�>�%I���?���!�ͣ������?�<��-�����+(<�&3C�6?|���l���X����د��~�N'��xl)�4��d\���3��|;YR�FŊC�S�+ד��ƙ`�q���phM��/N�C�5�؆V�\̀�+�~[Q���1��m��$��I��A�9�vz!��^`Z7�VP�q�9���]�[�oM��&�u/<���哨��8�e�X&w��Aۆ����%\O!�W��Zt�˜{~���2÷����;a�>�կsʔ��\�f��׋�P��'}� �/�1)��'�)���7� a�@�K�� R�` ��|�ŝ���N.'6~��)�ځ��s�xa�7ZZy�����/�o	�����	�Z�W0��Ţ�[���}/����ْX}�p0���g#(��9�#v�[ݬ��?���p��TO	/�Q�z]��(��0-L}*0;6~je�W;��Lr$N�&��@N]�A!)*V����܎p��>�+k�l�r~nv|����=��S-y$�"�۸��ܓ�8:��~Њ���p��A�t9<"����5�cdf�9xk>��y���X��Չ���539�1��[��Q�'3�G�OV�&+��A�������r���q��&�[,�>����#�h�D��"MJԞ�S�/K����b��_ƽ�3�ic�[bbjP�l l��a*��Be��خ��ӽ|v��s�k�H+}T̋���٠�����S��(��S�z�΍���J��S(BM�>Mp=T3|���}����,D�Ŝq���w����̽�L.�#���a&�Y�z����=#N��'9|p�Lq'�q�	��ʳ ���}�{��G0!zNm�2P����_�q�����.0�"��ԟ9���@k[x�0�:E�=��>�ѝr ��D���ˇ��kD�8���\�eV{�C�<������@.cB4!0{��������$y�KȧJv3�8���a�WK��%U��G��ߝ;�i��e��w���{xn:�0���.
��fvC8��,�l6|����p1�V66����ݹ�>����+8�k�.�ѵ���K�;؛\w��_��<T�Xv_��}{>����Dԇ��?�1�k2~�g>
j��Z|�~�ۀ�	E`^J1��C�:#��lLe$6kA������.�}eS�A�N@5fl�c����7�-�֘-�*�{�v���H�[52��R�ܺ�g.������W�!Bx�)Ú���!_铻YR������� �nY��6P̳���yL�������%
���p/:��w�p{��<y�zP?7\���<q
��������ܚ��8�F��j3C� 9��QqR�@�?`��5ǖ�\�5��	s��H7+H�U�^�Q�"$��0��޷�5�~ڿ�-���Ŏ�4̝3#�"2��j�}淨�s�.VX������b�P�rǏ��8BIs�N��~��[��c�DZ���d��T���g�Ҽs���<#J� ��̎�nꔟ+��mK������zg��NruX_�)��/%,&z�i��f�	r{����et��:���j��5�m��F/#�� �G4�
DJ�tPSD�ri8,�ig�ǣXί�_3�jfK^ԛ>
	�����NY��u0���=�/-��3����P
떴gA�
���_w�8������l��t�$L��Dɋ@Du�6��+h�ܲ�ʍ`g�M05F�.!��a\��Zw�-�1���h!�Ų�z���4���/p6��w@υ�h��&�-�h�rPH4��������8���9]�B6�1��H��/�"-t�m�k��'�s��>ҕZ��IH"�7E�&�h3���D��z�KPB����_�nð륱�$������yi��bj��22�'�s�Jĥ�mQvUC�*��.L�v�i%�޸�>yu9X�E=��~��_i�>���c�#� /��4^?"�	��q˨��$����K����㙧�-��QR����9N����g
��`W1�Hw0,+k��۷�y}��\��X����i�K&i+Y(���#낾;�|Oթr~p�/��qXDC*:���p�H�R���ȇ�3�!obRQ�^��:�S���LL�4���\����6�q� Y�Vd�A$�?A�'�Jqć�w~�
��.�7w+@�T�hM�=v�9\>�Ζ�'a��~�|ek���b��S:���|�E���C�X�f䦛oci�GN޵Hd�U)-�O/]��C�	���k6��J&rS4�"���㹠�ǟ��*�M�}��)}�:!~�G������_�	�0���*�P�^Rj�c����5>P2�)i�jJz5F�Uz�����,Y�$�� ��d�-}@��5�7�Xz���I1��,��;�������OK�����9g�j�;a!D���b��n]_��n�u��h�@��P�M��l|��Wq&R���z��E���m�ė%�핱�W��c�$�6�H:��gq~@N���-[����t����?�Vx�tW���x:]I�1-����0��t��\c�GY��s��e�W~09x�0k�K2pQ�홁�w��j!�\&N\�U��<1_×��S�ZBj�#��/)�6��8`9�KV�׵f�q�����V~��ѽ%����s���fG<��vQ�P��c�|A��e�7i��}(��X��u �yݚ�}��(������]��&���[��Y:��.�Kx|�7�O���(���P'��Ģ��p*�|�y\N���?�JE���}`0�Ee�M��0�.��N��.��w�GC.VJ��`�>��X��e�h�D��ciYɇ�&6��ݑ�$�R` Tl?��8��B@&�g�z�������$x���ϧ�����u9�2�%҂�E��Pf��$�ͅ��p�]�{qGH�縟��7�P:�rYv&�1j��c��t�?wإT��C�۟!!�ih��y�կ,��6b�۱�{�d@~�rV)fJE���t����9��O���O���I��l���v[;7�A,�N���ĀȤ�%Tb�r���E�`���{>���lI�ЙͲ^�(<(��,��ն-�\�E~C�7�q��`WP�)j)�� �(�_�7q�Oy~=gń����[#��x��EǓo�Hc��9�D!�\�u�VOoP�uF{����J���{J]YԴ\9�8�]��v�1|��O:�q-�6hK�p��ce���V~X�i���7���r����(�e��-�W�*�H� :E���d�/绿I�Ue�[��C��):t���H=�u' �Ŀ��Z���H��U��C	��:5}|:�Q��m�"%y����`R���{�◄�˓��'9��ۆM$�u̲	��\$��[3�V�Nx�pI߭q��S�(���G�O�i,%D)��[��M'���#�n��y+�1�0MX6�d��c�-�JQk6@�'�����}V����bp�׼=���/$��%b�5i�{!�c�{��ϓ2f���Ek4�a�,��q�"l"���̟���M2���߅�s�{4�ծ��'�Ls>B�}���'
-�(����d*O�C�D��&�B��9�\A[.���L4C��v�!;�x� F/�"+���Y0> q�^@؀!�؎��r4?%@Z\-Q���.�������B3+ѹM7��Тp�Q��̱��.�zF!\���k*��ͩag�� �R��^��3MOb��`؄M�$��NRX��8a�L�k<Q&�d0$������;0`
�/��6~E�k�8Pq�.�wz?�T!/��8�yh�D�|�i�!�x�o�4E�$���~�T8��&?��V�)gt�xkeN\#�3NLY� �E�o�&�~g�tGv�*���#��O:�}��3�q���LkWV],8 � v�Ǉ�*����^�`����MzmkA�t.��/�;2�X>7�#�M�+�*����!�:��]A�"�����0�MvG�]�A˥�řgcv��*����L�=�21(g��B��y�%�2��[�fx�4�>�}�"�TO�;j�?�♎2>��5f]����8�a��p�Qx٫���qM�E �y�a��}��w��C�tiߥ�r�������Y��Q��p�e�u6`�:��Ј_�4~u��۠�=�w���Y��8��f�>����^J�}9�|H�JK���Rm#_��-���f�x�{7�V;g�Z��������պD�t����Lt��	��%Z4�
{����u�|�Lew�6_�M*��/����J9\�[���'(|����W��u��,o��I�ƾ��\k(b9���P4�"F��w���E�5Jhnh�(�l�L.����_e�T����FRe�
1&���f��f�)��-�xr��,Eu	��P�M~鯋sۻg���m�OM���<B_j�V�F=ʖ�UK#�`��\�_c�g�MA�cqQ��Qm ��Iu<�48w��wP6s��N�ܮ0�4��p=�y?����=��tos���!�\���.L.&�m��ml�0�v5�Z&�B��l�(B"T�oS�!�J6�a�X�]��}����������"�#�,�o\:��U�^f�� ŀ7�Z�Ag�����H)��c������C�w�c�䆧ɕ�sn/���+f�}��w���vV6�����I�Ao�ִW��V��x����x+�ތÿҍ����ze���}T@?��9WnaG�%�R`�c�-�<�mTH>��T�H����޲~MN���ULYr|Y��U���]fD�C�ٜ���G0{��߲��g4�r��*B�w])Z�®̹~u��A>����:eʿ�c�O��`l�Y��)�9k�~�g���(�<�� �N"v�A�Z����D�/yTEl�d�ԧ��=0hV%�y$�Xc�O�l��}�ґp�xf�z�Z��� )Ū�r峙P{S{.���u�	U�tQ���sI�g�%�P�ЖP�9�ժ5�CWl0�?NZ���R��\4�F�l�,�p�h�=TN*텨*&��WaV�AF�K��N���9	0� �?�B�:��	�,�	�+�F���9�a�N���~$}!���TgL����>z���� �{.M@Kh���L8�� �<����i�A+������Q��xs����%�	,�t����������瞇��5~�����]{.�f�y�����k��
9��f+c.HB��!'��m�ݰ�vr��4{� ��`�;Ap,Æ`�&3P����{c��ƣx��m����9k�W!��m﵀* c+�A,����[5���v�b����z�sF���4��C�Y0�^9��]d��z�h� k��Q��+�e�<Q�~`e�h�̘�,���_Q�����6�4(�g��1���t�,��)"T��R�������T�Z/�o�,��j�e�W�n��*%z"Z��3��>h���A��?�N�qhXM*��h`�s�K�ܽ1(�?��̖K	h�UK�K��ə϶�N��"W$�[r��SfEE��I�\.O�]Ǥrʗ`21	�6ƃ�6�J6�-O�'�XJN����d-��;��Aa���ݦ?��DH�X�S�ɣ��v!���3�wc�7�C�X�ɇJ����[ج��<W����jx��A�b��DIm�*j�L�g�͜{�Y=�:��u&�L<QB|�:����Hp��'��C���=��k��E�c,*�+��Xfg�@��W�k�J�c7|,�G�wPvpLĒ��p�9���l���D�}�-���c����H*/7g�O�$�ϧr�K��ު֑�q\��˗t
�:�e��|B�v���.�����[Ai͓2�h:N����� <%�$l(��9I[��	�{��?�-�� 12�Y��#Ku�p�g�J������Op���F! ��`�^��q��W�@ǟp3$�q/2�\���V�ia�E���%� �,.�U��P��G���2O#.�1 ���.q�s�!�;)R�YwR�>�_�n7�*9���pk$�����5:��񌃭������==�`��\	ހfZ�I,PFY����1![a���:oOfCq��#x������*�!je]�l�:��ۂI�"����]�)�-�E�a�L�Bc�T�8�uN���3Iw��w����|4<Q���R�*Z�6k��;íE����������c&����aSK|�l�O�?w��ny�N_�E��P1_)�>$�����t~9K��6i�a��k�4�p�a���<��6��s�OA��W���pA���0[ͻ<�SF�&��7��#.�`�*�Һ�f�3+��y����A:���>YsC|���lَ��%�F�'/3\�&y@���)��G��hԛ1������	��59��;j7�����D�[OT���N��3��j� sU� L�/ðYPX�b�&��S����#��b�������C"lhv��j֠߱�S/���͹�nb�:Gv3��7�={(�(��e����"�O��d�휲��Y�3��7
e)t����ڳ�k��O���C�X�&a|h﷦��`�����}4K�����q��'rQ&߈�����B>�aM6=T^������\5�G�Xtg�C�a���Đe��H��؊l�f�3R�����ڃz�V[���5^�kY�>T�	��%�������ـ����Y<)��X|�E8�@J>nƯ��V�����>�ϊ�D�Иj�귺�
󒥟h� w�+� �{�8�k�1e���御.s�/����ܧ֥�Ҝ��d�%����6�9��~�
51<�(iE���q�IĹ�oE�[��\���;�а��V�Xj�m������ݸe��L���Z6sa���� �!���֭�'�O�����į ִQ� �r�Y��6	��1R�N�I�t��d[�f�:�+�H�=�wso�5�<%��������	��jM��P��{����C���(;v��UwP��6�Q�������)yHs��Dv�#O/HE�-�/�}�T������V���1�j�i�ڽ+;���������獂��\��\�S�Ds�u ���*�D�BZ6�:�R�Y�eA��?#T{h�Tc~��Ѹ�� #�'�2���{�$�
�ye���C��NDv�����4Rs�N�Z9!��g$�e�N���_��'���:�7���
[oo엦��]�,�G�u�����94� ��/�WN\�o��Q���$[�Fej�z̏��?/�a�p�W���.:fp�*�����"ѣ�e�W�]�J"n�=ך��������z�O%1�Y����v*�5�֬@&��j�M�]�*@�$M�`�2k�;��zۿ�	�E�Ea�Zڴ��5:|O��~��"i��\8j��_�碇�}�"�&K� {��m�Y��Knփ��r�tN�	�� ����:u{���߼�=Ɩ�!r�bX�y=�峗�e7Ԥ�VQ����<�l��� f(/�o�O�%|)��ѯ���\H�P��dNY�E�}^�7�ؙGf�w=nO�ɟ�=AQ�s0+�	��0������0�K�ov�j�R\�{���=���-�Vy�	���l"��^���ն�����]RkZ��!A��d�=rG�����!SV{g�$׋��Y�^>}k��묬�T�2\cC��瓤�$��_���g�����-t���q[Mn�@�#ؽ��j���'a����	d���Fy]�̎�fo��s\l1�zױ�W�R7읅���Nh2V�`L�;-}�*y*|Q�WH��,����i�����;�*X��
�AϜ �Z3�w��{˵̯۩���b�?�m�jH>�[ڵ��MO�ڟ�����/���<$:���$�����6��c����ϲ�Sn��Fx5�P"E�e�m׏*��iG3�Y6�����a����'�C~+؏��})�c�K,�̸��A�I,��z�f���n�YbY`��;߁+�'5�������I_h;�4L4�Y8s���Ǿ���pt�DoX�S�j�&�Za���t��f��%����Ð���PD���\����}c����Lڰ7��($w�iڛ�ߠd��/,�L��R@�p<��t����bE"�Ď�9�?O~.^���!�CH�4Ľ��<���B�y�<��c�3 2�f��C�.�VYV����z��ܵ��;���3��eAXvB����� %��C+f	\��dΌ��O5Pix�X�h闼��#��i��܇ˣ
�F@f|���]��	��f���є�!Z$�#�N�'�"��+��*�Ӯ���+�w��H�#�79n�;�u��YD�RT���q�@�erH�8�.,���-���5���~��&]���3ㄱ���x��T^�6gDt�b�x�f|"ko�ŗ/��Ыۢ�ǏB;��U�(����k���hRt8(x3�3]� �Dʖq{�����L>�=�) ��z�,���
�aޒ��<w�t`�P�	w�Rk+m����L&яN�5�q{�B�ݠ�ڽIf��'���(u�X��e��0�𰃍��Ķ_��L�__C��A��/�(n�gg��*�~c�|���`��D[F� �j�Ή�>
q�r>�*t��R��L�Di#(+��5C�λ����U��ϛ��5g	�;�y[3j��)s+����'��,��W���Ț��G�yg&�Z�{W�%�wk5Я�D�<���@uX_�X�9�z�n�+��z_�#�w�$R����ƫ����*Or�	<O�B�]�w�gΡ�V6;o���tLm��Փ8=�񟀈���l8p�?}d��B�gদ:��^�u$��q�B6�G$�k�N&g�[��oԪ�T��ĩ?�����6pvl�\ea��2z�A�1��N�<�i� 3|�	M�b�������.ޛ|,}����o�vK����#1�3�sk�v:5$�Z�8ШeR:���{ۼ��Hr�O=,e�с݅07Nu5ދ7���c�r4�-�@�=c9K��j����3�!��T�v���Z���N~2^	���x�I�@ʐ=��Bt4t�w+gpy{3(��y_��2��_���b�v13����]$��i��.dI���Ő�w�+�4���k�P�������4������s��X�?F���:�\��m�.�2X�[���J 4D�(��OKr'J��$��H��~���X=/8��{���>Z�aEu�r^�:涭_�ү�>���soM�՘��^�v<�0�Űc{�昆�5��/�\.���NLoLo�����g�G �R�3�ǲ�ӡ�^����RI# 7������Փ�[T.���QuUF ���y�8]�P�	��F��Y�9��LH����Y�f�_}��b���ϐK�������A���_�R��q\�	H����:���F�D8��f�N37�&�>�䁔B�q��� R��c{޲��&"ʉ^���J����J��y��	�3����c�������Txߕw�E����"��Z���	���R��-��v%��'��U���7؞0A}�b�Z��M��oD1猞B����%K�߽j�݅�p��#�T,�`D�&�Œm�%��G0W�l$
����Ȱ�|���^�r(�G8����0,�N:�b$�D��2���k7R/�|+����@���R��
��!�?8����LlV7(q��		IZp�����Ȑ��4����*��`@��[��_�@�c	S{�"��j$�\�Uyk�nբ��E8���"/�)y�2��U���<x�?�vA_V�
B�g�30�Q7#�z{K79�+a�-�;�Ҝ;&DŲLA!���-Pֳ�Ϥ6���'8��|���8�����
�M��
��wZ��j#6��ۼ�= I��D'���)6���Y�~	��&�Ю��-�R����3�'��Cp�s�}��75jHu�N�!�ُWZ�8���}��;it�� �k����_]}���op��K�$Ao���H+\ڲ�G�����x�$dt1�b�����ދ�h�D���=:�f�k��P�{�����z���ol�ɞ�u�J�/��;`��%LC�i�|��=���~��ΰ���_����M~�q���*EO�ҫL~ʥ�>oH<t����,�r�a�W���@B6�%C���i�0���/i���P�Y�wJZY�ȩ*\��g5��ǅ���b��f}Ap�|�Y��{VAa�Lʯ�@ij��<�g�qk��:&�Q����)̀>zO��%
���6�,��� \��/|��>5�q��Cp�%��`5]�Pp�
���g�Ͳd7;OkYȸ栙 �"yXV�Y)�#�MU�y�r��+��A��H%i����%q�A����1��Y��T�##K-!�Y��u�3��q�Ԗ�С��y^"�ʕeG�G���{:n~X��8v�{ _�4b�#P�����z`=�a��.�9t���$B6f���V�a$�N!�$����R����UG�ۺ���W-`HؕE`�U:m�h�Ŏ\y�Eǰ_A�Wl��b�#��5c�ڌAx�m"���4g޷o�>^	˶<]m.sJp���+��CƵ����yCXp~5˅�[�1�Б��&h/���ln9����h��? �#Q״7�)/<��Y>�&i�h��"�D��&k{=��F/F�W��U�%u����ts��s��-R�5e+i7<�����2�cEw�\�ܫ[�`�հ��3���y�|�s��^z�<�y0l)d4��T)�R�T�ͽ9ϧ6�MW�H�Ȳ ���>�c�ܵh�c�x�T��XY�"��,�:��8[�4ۛ�=�W�Em�K���0����c9u1 ʻ�Q��8Xȗ��ɼk��n�B�E�k UZ�6�C��h
T;Dd�xy����[�ſ��Mb)�p���BZ-�w��p�g��fغ��m���Z��'J�}_s�� 5�@Ml[@���@����-�u��Z��ݤ�)[R�QS�蘐  ���U�&�r"���j,Ҥ�.��\A��~���=i��[˥����0�͐`Aq�3^�ׄ���&3��T`�������%ha79~/��/r��3�����v�R�ɫX��qr�=y^+��� )GRr��qu��h��xC����xd�-��0��q��_=���@W��cs�7��J6�T�LT��L�I�G ��Q�xv�(vZЫA��~��V����21�!pL����+T��Ǻ�N�nX�,�˷C��AL%Ǣ�.�o!�,�q%�֜��D� �GU��)`��1��^�a��T���ֶ-�(�Y\l�2��w��^/+���s'�;�b�M�`?Y�,`��*|�dq/M��MpF+81y�6�4�w):%iC�8�]j��û��J>f"�"�CG|��Թ�٥�G��UR�=��� a�\���D�hK�����~{�k��eޱ�\��Na�6�e�^~%>�x)�rz�j����� |/�����@�����NjT�-�1�\>�,��C{27g��� ��c{��>9�[J�s�u���\�5���i�!���u64??���/��?����;�Q<wz#�c@9�C�ڜ���d��[fE�{w���cD�-�V�e�籘�"Ȓ��R�{\í��f{���5M���ɜ!�B�]iO��9������R�����~u�3�Z� W������vH"xz�.�U���p�~�m��H�+��Q�3�%�V���,�|����� ���6'!�=o1�A4�nЛ�u.�U|I�3�����&�#H�/5@��t��a�gK�p���@|�~q2<d:~yB��c�9�R�;��|䍤ZѺ���ι��sb��!�: d��L�8I�ԧ����m��}Ba�$�}^�V`'.I���y�ĥ�x�<^3/�VK�1��2�z
���wL���9"���f�"_�K�Y����ː7��JK?V�6�X��x�� �
'5O`�y$��v�0mq��V��b����>�B[R��N��:��i�G`\\[vy����e?.�QD��'������A�7o�	��8�n�~O�լ�܈��W.*�a�������]ss��^"A���a�6}����:�N��1VW@��kWv,��G�b�e��X���K���Q<�'�_eZ�*y� y�瞿�}�ڈ��}�C����b�^2Ӆ���\� �X#��	$r�OB��e���1OQN���u�"J�Z�Qư��S��'9��6��ǂ����^d��>��S�v�7���l��PN"�B�P���1A3�^������q�8"n堏�wQ�CO��%ߔ���KG���ks�2��!fs�H��<s�<{kƯ�:-	�t0Bԋ�P���I����;��հA}ٛE/ܻzR`�+�t���9���#T�ٝIV-�#��Ru_�J4]玺�����U4�p�n7I�o/@ta�jdq^����uz2�Vo�63������K��H�M���J�Y�� �)��Nl{��<D����E���(�b��#� ���v��i�D�hW
.��0$�^�<�&�[##z�)��1S{��¢��O�rbpL��l�
��_H=�W
�=��'�H�3���%0&���	g|)���
NivGnM�)t�ٱv��N���wv�q���E�Փ�{i24���(��Ry�iûq��tRX��:y��F9G�ƀ�qS������ ��Va)l^���~��vU��Y��G[�i�/ϝ-/�Ga��	$��֞�z<��1 �,����h����n��k �Fk���s���;G��1
���H݇��0��6�"ܯ��.Ҭ�\]�ȼ���+(H��R��Zf�Պ7%6�! �N�6����ȹ�y��2�+]�/ᯊ(���؞�3|}���7�x]��o%�[6�8�u��ϙ�u̲1�QQ��Tۖ�xS�s{׉Eon�ȑ� -y)O.���)�qp�b.qTAS�ӌ��Ҥ}��"�����B�uU��c�&�g��U;%��i�w�kԇ�{�S1��oh�5ў�n6���B
.w�KX**�f}�$A�F�a�/�w̃Q4ZI�5���g���'�*H+�Ϯ�է"<����،�On�30�O��#XAe2��¨�ɮ4����9Ai�-hfb��dD�zl��
ZެXh4��Ø�3!�?<4+�^$R*�ޢo��0���>�%Q+���s���:�OC��IN^vS^��;��+��|u���ȵȌ|���Z�W�@g�K����=#�MVB�PxW
�	rx�W����3+~ګ�d�d!�Sc�7��ᷚ�1ү����T9�>�
-Igm��  JDeZL3�BĚ�|映y�3��o:,�H�ң�S����d���lV*{���L���8l��Gūhc��CO����%�/�t-hw��|/{$f�t�l��sX"_�~	E�Y$�>�5�Tguh�T� v�(p��mh��&�� �m�\Db 2�pęG�d�l:���>����^Ƽ"���|��|��&5wc���4�|�����#7/���'��{9�D�=��gR=�M�3��.���c1�0��bs��4 �$4 �I~>8��=������xPqg��*���z�yj�ʸ�����l���#
t�|�Ȱ�!�����ײ�_S/��2�4Uf����������Ͳ���&r刴%�^�#B�W��hb��1龓L,�X�vg9��ۣ!� Q:�Ø�1���?�,��P�����-{����y��Vjљ��)tg(� a��ۜ22�jN�A�TP!��zIB�i,̼2z�g�����I�Vc�)j ��1I�1o�DQ)J@�ʟ� ��k�"�2�͆d���*"��d<��h�U�&��t�ˊD\"/_���'��Ĳ�N���f�G�B7F�W�5�OŰL����e|�ČLje�jYe]��W��F'n�w��"�6 1Z�Ew��S�x
�0�C]~ꑔ�y�O#)�>-�,�aIKl�x�o�I��;Η<S7̢uA�wt��n�ݯ�MU[MK��t1����CF����~�n�|�݃������@I	������)Y<,T��{�.t�B8vP�P��)nrR��(v������.W��D
\�R����f����Y�klǞ=�`�2�@�4npC!�tL�,���o���Ͼ�F�O��<�V��[���ݾ���rĕ;�DxE�NXI�AX("��q���rW�����${���,�0�tj�1���W�]�����"'��@��u�]�"��QhфU�ͼu���7��%]8.�q���a��69~[�l�U��Ц\P�A����S�=��3�$ۃ�}�h�Dr _tlqqh�Gd�J��Y�ߥ]���]�P?�T�2���{]T�*�ؐ��p��7P���~g�!�H�
�f����X/X�����Rp!�����J/Ñ,�g�t�j��\1��j���d�%VC`v~��R���_[�ts��Z��k�@	lQ��8�k����#�˗wOk7"l=�#�e��a�9ن\r�K�$�:	e�/ )��#xE�ȯ�7�-W�����T_�W<�]y�����qz��V�y��p����ܦ�zF�R���$rچ��ʯ�[]��Ni�,�?�'���Il��+>$:�U�+�^���4]u�q�j��l遱�%�����m^�J����^��d���Z۸��c������5������n�9"�E���Z��N��t��ں+V�4���o=�bu��/���ؠ��H�dUh��F�*;�oj��^��|o�$D�r�,-�7z��>�X�:��N.�v� �2ѡ�V3<
�Ggdg����1�si�w�\���|M`��b�fQ�f��d�Z�q��4�Q�A������O.�:N^@f"�0�P����،���iLQ������'5B������sΌTJ>�)"N�^/HI*̽�-�g5�e����U K�Wo{C�i1��7� r���{NK/5��"b��¿���%\ř"�v��&B�"b^j�*��|M���ܺ�$����v�� 5u����dz1�3-M2�7�9xAH��@
V��r#Z2�~E��d���jzg���Y�)�r:�Ǐ�|]���1t�y���n��U��a�s x�$>2��䣖 Q�v�<�.��N�³z���D�L����,����>���m�B�%V��x' ��`=O�Y�C��/+�o������ ��l�����m9jn�h$w;_N}:����g�%��HH���vC΋IJ?�2�i�2/í�`<�㷉�׬�
��F�v]J>���wa#��#b�]�=g���2�5�ڙX.ZHmPK�P�s	�̢�{�Q��U#0�t����Ш�N�/ި
��9$�ICi��I�W|����[/�|��]�>��b�?��df+V/$�W8>z�k�)�;MY]�[�"\�%����NO�v��\e��x�q�G"��D�s�����
��t�ܖ�|�=i�03�:�̀�	�0�a�p�0b�9���uޑ��k��I�x�L�)��\�����$S�Π�F�����
r��C�;���f#a;�� ��Q��3��.�`�����	��n���?2�􂱧�#-*���@��p9�����K�в�P��� �y4<�Փց�z�*J��\zU(8_RW���a��ؒUJ.l���⛆*���:�2�ͅ�L֠eC���E�į�B���9H�J�m	#9��*dg�Z�i�;RE�V�t�e�Ɛ�	2����!���1��J�JSNz��e��Y��j���K���͛�e���9�n)�̕������AŘx�eŞ���鴯�H�dhBk�0�����������f�P����k3�dL��p!)��r�|�����G� W4�j�R1w϶���"����#�"k�������@;����ʃ�J��N{n�!/#\�� 龜]Ƙ+EM�P���[�:`S_��|J��FO\:���涺�� �~r`����D� ��7����`ڷ�.7���c�'�f�q�_cN�`���*q�_�W���vYv���H�����u���.�fq��e�t_�1@��p���C3�{E��#�Ow��W�+���+����hk��a��@w�{��X3I()M8�z�*�[�=�!f&��؎3�^��3���\��j����5y�.�+P����NJM�}�c�Eȁ@3&��ZMu��@c���k6NJ��t�?�M�ZZf�ؤnau|��̧/��5!Zh�6�~ ��j��}e���3)�ޒ@鐟qD�{�%�s���i4�	e����/*p%B갠�yұݘ�,,����a���TT�`w:{���P���
�$U�0���&���]\?�'�;�jJA��u�d�9֠�H����:0tY {�>]��9j�%U�u���	��FZ^��-'�8u4H�j)�(��7���w�F\/�C� �iTM�ʔF��5�p ���Q���4qظ_Q}�ԡ��C��nҥPr���[ՖV����l���$�.��ݹ�-��{PsG��z����-6Ъ w+:е� �g�$��+�)� �0w_Ȉ�G�h �άf�D=��7
}�F�秺Mf���Ɩ��sS-9����3����!��M��j��T���E_&k�~3qrln���KUz��pcc=Nߴ���i�n��#}4l�ma���2�x�3��+�oQ|��x�p�&��뷶��0�gn�@ZOp|�\�F���=2�J��$1��.D2d��85����dv�|CF�eԮ8�
�:K�2���"��L�����_:�	bp�c�s(���������>�{�� 4����%���˹3��u�� �1���-%XvQG�շ�e` ԅ�[Re>�|R:8��"^�����:�OK[,I3s�K�T���Y{���������{��VQ�V�{�gb(�� ݅�k�� R�F�хZ�9=���\_� �Ẑ�r�V��v��7|�<lI�Jiq����)�,@�$X>�Ǫx�ʽ_�{EJ�G0�h��n+�ǌ�ofVV��s�&o��_��B�z�L4j�s��TR#N�y���E��W*Jj���G��V��������O�s�ʨ�:x�~�_��'j/�cD{��Q��y�cY��#Ua�
������q���RzH5$� ����FJ�0�r^`]�U���Ѻ���'��l�BUV��֙w�h���D�>2���9QqwG�d����V"��F���8���T^	�p�k��q�3��bt3�ڵ�jo"��7�\�NB9��K6��9$u0t[Q��h*�p��'�g��X���Ti([#���ݼ����Iϻ]�n�Dv��2�����#�"#uO7Y}m���]`���|�ʲ�f��H�d�� 	��~/��7w���f�aiF��VSe��M���.�
5�C���=���w�
�d5�URU�w0�W��NEg�e�A���HX�Q��u���Y�W\� �I��)����|����q�+��� ���R�	!��J��h�a���=��l�D�Ρ���`���,�nئ��9x�����wr�ɐ~%�=p �%��0\�ȗ��gK*��on�|���y����ϛ[����B�o� Ɣn��O���>Ci`-K��͊q��>?�Ʀ��S���
��c�4�Ժ�n��,	�ӗ<�i�ۊpɢ�W|���f\��#S=V�j�9&��"m2!�:����ڝ���fɋ}��/I�K,&aV���|(�y�rdT�-�yf��pd@+:�%��_OA��Au<^�ں��:���'<jbO�GʘxmP^�A��j��}�����52�����޻�����o����.Jk�>�O�J2�V���3}���v���F|��?Xu^x�(4!`Cd���]G��\�w�X�^~
r��ϣ=��W�c���H�K�F�C3�.�q��KG�s)�˅�����Y�;c�j��.0fs4�Q�[�@]��,�P�x��~����XL�:U{��5��Uƺ��9>�訝�3@��|���r�+҇�/����*�,B5�|E�P_`>)k{�R��H[R͓�!޲�Y糳@�Ւ<C7�U��ҳ+-�h�S$�@�r�8���+�_*�GVFz���C����ވ8�L�����6r���Ljy'>��4��Ѓc�ųt�;�a���Γ�C6�Y��	���x��]���Q�7�6����Bƻ���J���O�T�N-��o`�'�\�"n}В�2u��6w#���d0���s�d�o��jQ(0>�/$	���h)F4���i��Vz(Nb��"U��ڡ.v���1%+��3���M�i���l������0 Fw��vz6�˯�����Z�#��}����a�a ��7��ka.
(F�T�2���5JM�������8ǨuE�U=��R�\���]��������Cf�g��S�M�A(�`HMG���Zϙ,X�o4.������Rwɵ:��D9t,}5��*-�>�56\��w�?k���FlY��% zJ7Q������.�ʢh��1��.��!=?�8�5��eD�;@�G��G3���q�.�g|�csa�R0����Q,���`O�0��=�L»��PK��ٲ��f��3��C렎&:���R{ IkAZ�&�9h+�t�7<jk�ϊ�ߗ�A�h~�������E��-��q�n�F���y��ڵo�RJT�[!�"t���~�^_��hI�D��=�Z��������M)�齳�YQ�"x�xBW���� ��q���;m��YO�X̙�����f�����̰\�����lG���N��vGz.�9p����b@���Y״�}A��I,�b�¹9�_@ڽ���ݤ��Ʃ��p��ݬ�5�2�{
�������M���r5�N�w��z������Dg.A�\�?a�~;�\@T��;Z�UY� 8&�	{]���=V�K��М�tQ�y��O��� )}���Q#<���ir�����r�Co��0�NX�?��("�H��,�&(oz�	 @����.�Ȯn3��܎T��[+E�nh
ï?�ű�}�=���lJ2X�Kݮ~�F��+�3͡�'ԸF8z(1$w�B�mt�_I��d�g�����y�~��.��	y�~����6�Q4�ag�|�2���r�:Ԉ���#7�i֔ YR�J$$r5�I�6Z�?l��)ڧ��ߊx�ut���m���f&��~6=�O����@���<���d�����9��}�e���Ml��s���)�k�i�j�U�$�r������⓱S�lM&��;yF��0DUs��sd<|��HlK�S���ƽ<E���6Ic�:�Y�n�e�@�"6I����Su��*��Q��:2��iL�C�l��7$��ac)2����ɟ��j���C���cV��Ƭ��^�[��W�а�.�Yi��M��p-�K���ڨy ĉ����:.��$H�m5���\~�q>�)͍X��~���D|����I��/طb�����ē��l�y�~\ʭ;��DԦ嶓�{0����˘�;'�2�A��
��
��ͅ�z�2I���J2�Jd!3���+2��а�P|4�G��&cQ�0���Qm!�%oE�J���fٲ�7�i�����R�]x�	�5�Ƥ]�`*�	��Ɔ^4v��
�Ѭ�M/��Y�j�*>h����m�XЅ��.�/ �4�SO?��sI����/�n)�$`������r�#D}���w-ذ5=�#��^���^;o��j�]�o>�l��9J&���Q��a�I���X���ہ���W$�4�,z6�!'������Gua�B�͝�0g�v�7�����s��$('A�Y�T�y���%����Ew��=�p��\�>��}E�B�w��EM�5<�:g~��j�7�L|���hg�on��8&�Q���&�i������W���?����yE%-Z��<@ܚ����ūy����n�6pV�E�ɂ���ӌ��3â?EL���r�cEv.荢�Pi�x5��c�tD��S��?�~�lS���a��\F�m�BL�
Q�a�a��c��5�I��	-�-[�Ho�j����5s�}�ď�F9��Olc4y��LЁ�YA�u|<"�np�S�7�7��ސ�Y��H���da���W�J�����«��yV�)	�ґװ���NI�h{�^�B�v�m
���V��f�{�jU�ew?x��|��դ��/j��|ax𘥼k��9T���{�'&��!�� ���麔2MXE\mMj��=f���Ґ�v�E�2�n���T��k"q��] �`��"��=^Cc�\��N"Y�0d�G�� r�֭s.���r����!�I�PL���L�:�SR�����	󵱙�E�cP�������Tex��V�!A6B�W�^'eZC( ���א�}��̫��g��E��B4c��Q���G��ifE&È����#�WԼV�²��a��v�8����.������a<w��zƾ9�cfa"�n���x?%m�X�����K��>� �:��O��l��M8;f�\Ps"��A�-�Sv��-����n�m�`?�B���#v�w���?w�AM���+m�����A�D0�z!�Q|}Kf���}���X�Ê�:���5���o����}q1U���Or/@���Mq��q�2�����|�]�����(�@3�{4Q.�	� >�6�E?$W�#��Ia��%�W���jà�]�]"��T84��^����&�v��Aaϝ��tS��*�9�k���SCc(�=�o��%]�u��v� ��Ҵ��^(*%VW[6�L������yu����C	����������1�+j8y�gN����-�ݠ��0�Tȁ5��<)G*�1���ԁ:u�+*B�h���gn2ۘ�6%dX������u����@$�c�V����`k	>������s'}�WRry��IO�����+1t�قiOo�dWF���:�R�q�i���Uǔ����
���K�Gҷ�)��'�6U
;HY�|6F�
{1���8�6�گ�-џ���sj�:28<�����ė_{�Y�\FG��f��EO�%��s4����/������G@�佼�v��9H1��сSH��KTi:3�����X�D>�q-��\-㝿���?���"��^`b�Z�edɴ�K����R
V��gKVQo�ܣh�`k�鞤�`b�Qq�GIB�}�k�#�ǤdU��ώ~���=����="2��S	�&^\����	���6$aK��-�W��F�譼	���qf�әS,� i:U�x���y��C��(79fV��dY�اS�� ��V���ز���V^�옧���3�L)!�Br
�SV`������9!��:1��zbSԗ:y��+5"I�X�B^1����IL��fB�EQ��|��I�w�U6�>e��\�1����[K	=��>+ߧ�֔t��آnV;wc����l1ց�W
 ����d9��i��E��#8~�z�$ԅ�w���d��۷�P_�_�
��u���z*��� W1�1�s�zkԒ=�B���jXe�B��-�.`�Û��r7�z#��l�?����Fg�(��)�P� �S7�}�X����Ş�*Q��>ޗc[��Ш!��8vs�b�e��X��	n��\���Wq�EC��Z4��IH�0��F��&G����&���X�A�tX_&xg�j�8s%Q�ǚB�\) ��)�TӜ*Dg�8P�ܚ���"��>8)N3�\�vk��j�Ń����Pu��7�2�q��S�c;{��ZqPο�Z"˞�D�o��q'n��-Op:b�����!e���0\��Pl�$��l
�,JO�����z���Onz��uKc�:���f�ZKU^�F�����������	�xs��6#=E5��!?ı�-��U�L���_�����`>ɫ$΋�u�k���k:Ps����n��Y�C�KA@I��ۮ�w��ơ �}��˦��~�׹;{��b)��
C(0�^�6'�1�a�b��ݖaL�j4^feXhsIv�|��7ߎ5(�)�����z(;u�Z[[}�IАw s��N9��3O�d�Y���{�b�Q�.�F��������q����b�T�����?Ӏ9�yxƺ�&D���R[�)����HS��ݺL#X��Zz;U�bf���9~ߏKk���6o�`3���裟�&�;�z�ic`4�& K�n�ȃy	��!�Ab���j��u�Yn�
� �����)��5a��� S1���L��2m��NyD#Ѽ�A$Vxʢ(��E�h�m,�TvCl��*���Bo�����yI�Y�9��r���573�뱔kc�T#�xR;vFk�~u�����v8jKn���'���5�A�& A/��|sA��V�x����X'� �1f�9�i��ʌ��*�y�~�G���)�܅VՉ��B�������j
4�N��v�#�|�2�H˿�P.��M��]ۙ�Z�~,b5��Po��Rc�[�[L؁
P�XHh^�K��3w�,�V�S�c�,�
t[�t�0����� O�K��$1�t_��ֶ�̖ �ND���ל���Ů���m+p�čd(�ꞧ� �u��k�S�Nc	�x��0nݮ a5]F�P�+c��SBU~԰��aEGr��,�T+�����aׅ��n�3����]WS�o��M�;Ɍ&����ŶXM���A���,�v�E ���sD���iQ�r���Q��<F}K�c~ƅS�Q�p TE.\S�I��J���s��h��hx����7�#�������1��ڀ�>��
��'���-��;���׍,Dfܰ±T�(�R�ؐY�d��ǰ@�ܲ����t���=�Iu~M7
�XC�����Wop�E�f���|�
��Oj"/��/w�-�&W�`v#�J%�?�vU��HV��5]�Q�����*�u>����L2Ȏ)j�,{�X5
6�e#����k���)5��Ph��X��[[U��[�/K'i�����`;�[��Z��L�M1�qa�I%��ǎ
�/�~5L�s~U��VQ>��k�ٛ��D~��
����џ(}�K��FKq5ɦ��0��h�ןW���gI�W�s�P���1e�zT��O�����\�	awu}��$'3(H�0jL^`m���s����|�<��~h4� :����M�W�B�q����3���WP{��P��)�$�*I�����Y1����6`��h�Dn��ze[�/~���ӛ<%�Y�?�����j����~�������):@<��K���̒Qyό�Z!��2���������6�F�b^�s�u�B���&��8q��Y&H�/!��̉����_�ᅜ�	v��ѹ�q�"٢�������8a�y��{A؋㨛���u^K���81�1u�H�F�GH0.e.IΤ��̜ɔ�
,CR�߳���9�v�I�$/s�������{��x�^�	9�Of���o-�,��e�[v�Wu|0<��o�]:��cb��k��<
��� @��u(�o�V�_��hĎN=.��q�T�~�t5���%�̊�<d�ֶ+-X���\#�?��"���t�ܿX`� �O"�Q؊��O��& �0��IX<HI�5�#[=AH@|��J�eo�&E3�Jp�-� ��YMv��J���0������LO	�h�\�����,qv���wX��������=pJC�;��0�Z�æ2=����>p�� ;%��ӓ8�<�hT��ױ&!3;�2�b�#��G�J�2V�\`�rַ�FGs�w�ݪ�7��?�j��N�<e��5W���fV)+g�4��Hj��`�F�(T��o�=�sb�#p��1C�Drl�8wz��]��~g$3�K���:�v��y���"ק��\���n6��q=���>��L��сנ���)I����$�Zp���R���<�M���:*\fǥ�t���>ۅJr?�^Sd=d&PiS��ǍV/WC�{\�u`�Wb�`�D��\���Z\i��ߡ�a���L��f�v�9�]2�����7D�	�b���YژN�:y�����-!�X���q�� VfTDeK�t.����8^���3
-9>Y��i��N��7�<ᵋ������%��S��'�>7~Ldx�P����qk����e�i�e$Ա���柭��,P����Z_n�Тċ��JU�����Nf&��~t�蟿{A'���P��K� ��lS.t��R EMh;�TpVH�M��xD}G�1q��`*Ϡ}�*�ePL.O��!t������h��`H��f��2MϬE�����ׇ'Gȥ�zx�v�^,H�"N�,	�&�qگz?Lw"��)Fr�`���/Y(~���t�a��#$��O��+CoG� G�7d��#:9вX�EQ�M*���H�H��8�SU�{m����Ó;GeiT[Ɗ�6��hF8��'rO[1R���&�����
�s�R1u)�,9h���,����v����utK��q�!�5���E�s.��G���Q</��C����j���I�6�H�w��j8����@�F�O��D�])�c�c��8�6�������y������|�S����Jgi�$�.NE���|��%oi�O���-���C\)�t�?��q��Q��u'�jWL��і�v��p5ߍ;�������|��)�V���/����DL��T�Uܗ{J~ϮAَ.{�A&�ȩ��<d��(�TC���!��8�F�cpг|w������Q7�nSr��
R�L�|Av�(�\/)��u�F4��Ӧ�Î�ԉꭐS�8�n[�6#�����G��s��Ή+�;ӑ����������C:��V'��x^��zi�Y�xJG�w�,������N��9�W���3	˷��^��]v� �WTT�+��O/q��Ž���Z��EE���JyN��s�� �m�0:1~�/���_�R�X'��r<���T��>$�.��&�ժ+ul��L����������|�y���Q�=da2"�\)�ĺ����l��/"���d�}}ւ0}{Z��U|�A��]��k�����y\R�u�*���9�2�,3�O$У��W\u�a7i�'3�jbڏ����q�q��7�!*���U��s�h����r�{��^�ι~_�j��_y����t)꒸HQV�y�T�,��c��-�yB�Oԕ^���bx�+�gUc��j=�
u`l���k] �#t5�2��xw˲�_��~qO���$'��� `�Hf���
�M�8���_����(V�����L�V?V��+����Y9��?���@xO�5�5d?SJ ޹���ź�,d�3F�e����W�\Q���}	f����9(E��AX\��,<�D���1�_��yi��]��p��B���K��++��i��ފ����U�\t���c��R?Sw�|����鉸� 1���]U�6�1E���[���[�?�1�H#C�%�.Gcy�5��KlRBS�	�Iv_����@	��6�s����4�A�Q�{��K�3��S��vx��F�q����2��}�rmϕ����T%�+�&#������o��I�Ӊ�S��iq��*x�3 od��0�mi:��%�C����������D=�z�khܷK�Y�Èa��¢z��@�+����LA��"#c�,bϣ�ߙo�Mr�n4@-�{����HN>~ڑ�*��.o�U��N�_9E�u�z+�؃eu�D�Fh������"�ϗ_�o�cVRk
6<��{$�g�q� ����g@]���c*�T;�ØQ���e`2��r�9����q�ŷ�}cćb[~Kyp���iݪ���B�U#��iք���*�Е��	kH	�&q��x���Bؚo�=d��_Ǻ
p�=Kd�W�Y�.��܏��佨�ݩ��n�p#.n��9R��?[�
c��2FK�tM��&�՛��K��7V�G W����+d��l�RX(òQRIޯ�0���)�R�>,�E�)�' �i_-��I� ���p��`��i֌�p���U�g�����,]��|d]6T���0�㰅��%v/yE{qv�T�񑫵l*q�F� ��|'��� >h�~[ӸP-���@��)��kc>?̚�!u�P��}`���䲔�``�& ���	�@��R�d���g9�<զ~�	��}���6/��N9�( �i)�;Vg�S!:�T(u�����z�c 4�S�D$L��{u��?ї14�^���x[��KɊ[�ȗX��%;+�wz��^.�(�2Or'�&�^u�{�]�D�H[���!���Y�Ȣ���F��('��<y�I��������.:5�)�1��[��s��n�v�OIB;MX	���=dG�hǍ=?O!.�b�\��q~�6N��HТv�ի.��gǑYnǢ;iW���,�p/4�Ts��^��m��]D�V-��p��^w�w��pr�{0��6q[�����9x�'��?	�-�Z�Ty_��t6
S�ʂ�E�0���-�B(C�sɆf�;�ͱ9߀�XO����!o�|���o��ɵ��,�D�¾��w�Ai�,k2DxX����~Օ��N���luc5
�l��6>�
���+q��+���Nx��)1��.���S���M�%��)V�1���}w㣜@��AOξ.Jf���r1J�3��O6���»��qFo�<�M���5[��Rن�0���4��t,
Ί��j'.�[��� S�A�p��|Х?���d�Ѐ��]��ɨI�8!��f�;���G|�sq���r���(BI���Vd4�d�,�V!�B��j��	�.�U�M��9��^_���8C@�Ұ�u�l�����L*©05E��d�}sO�ZU8[���תּ:-�Jԯ�9���.����S�ze�Z�|����<5���]�
�KǞ`�֒ymV�n��9�0��v3VmylLOM���Y@�y�:�5��ү��P4������tK��4�q��#�~�7�(w��}X�{�]'<��/;��̵�׬�?�,VAEG����&�PÖ7�X$�*=��E��m�0��v��N��9��^���J����s�ruMu�t��:�kl]C]�V�@=�����X�c�����VgLqg��-��O�v5]^�ۭ��4���{}�ھ��ʗ1zK`g)�N���7I�cd&<�|�y���,�pP����c�<���V����jb����g�͚CK,<e}NZ��0|��x�;�M$eD8�uCﴜ,N�]}��z�ÓL��*���	�Y�����x �GD8C2{k̯�{J�B��-9y�u&��.��XRR���c$�8���?]X;
�<Vyʃ��B�ݟS�7��!�'Dqf��HI���澕�_rBoY�o
�b�i͙ɣ���*��^����xv���	�X­`���;4��@P9u�ů�%��4�����֫��[Y�%�L
���[`�P:2
�ټw�?v�U�����)/�����Z��S������FwG3Sk�d�����<���>f���T��9$c��c�xn�O����ɒ����"]�o_�L��@7�;0��(��Y�ʑ��#?���lz���o��r@�6$}O��4����/Kh�H��h�[N xB� ��"�U@����SǢO������O�
z������7��F@��6Y�d�59�c���4�H��(D�q�(�-6���OK���������QZo�Ԗ�0_�Y�D�w�b�B'Jx�H找��lI��Cz��]�3����T���`4v��az�L���C��G%Sz�'8��k;[;^"hCu�c<]19׬ ؔ#1M_�G��-0�Ϣ��9�D�,o��j͌����i.ez���4$ahi�N	��P'��^��~n]h���Vq�Y#�����궆N��5��y'�Txg2pKs�q%d>a�ܮEa e69����B�;��" /�1�d��0M�'
�qߢ_��J���S�[H*�#y�=9�p$B��G�Wd�ZZw��ΈC&�����d�` Np���ñ綈j��=/���J̾�Sn��[F�D��*lO�����hܴɼ�n�/�N!��{��j���b�A9��A�#�)������F�e�帑1	��4����lZ����
�f�,F�j�^�7�b���?��)���0%,�<^���z�����u0uE��Ϻ=b�Q�- %�C٫G)������R�fnƙ��{�]��ɺ f�ˆ�q��Fwn�7�$��ef�\L�s[���"�-��#�ʕ�*���
��d`�! r)M�,�����۟�AۨU*h�ij��O?�0�)�b�H��]]DԭM:,r�%�ܾY���A�@aMn����g���+�S�"����2tbH�|T\�i�G8���Հ�3m�RP��/sqK:�e��X0�$:�=ApxF�Rk�'EQ%��2�]^�EZ��g�e�MH���~3�3�j��Ik�Ξ)���D��*ml�(N���W0��+[��!��H�<��E����Z	A_���)�3��_8���~f�7�|G�rg�sJ�*��&߽.�����x/wj����|�X6���e�)��j!�_r��6�vO��N��T�����g������6WòK/�ͻ��r����o��اXv1������ƿ<��7���H$pZ��C�5(����q(������X=u��()��@0�*�(�ή^����1���Xg�?��!���Ք2H�����uzIw>j�A5u���W�����3i9gP�yl�4��7;I�B��<�'M3��5�/���7�H~�R?�AP���R�3��|+PEJW��|/K��QGy�m@��v��^^n^z�1Z)���rXw��w�G�\.N&M��|���t��_�����[�K�p�D)e��X��(��>�����f�n�}g����kqc
*jc'����|J�΃O��x����T�o�{�mzV"��RY�u
V���c�S��9R���ޑC�Iӳ�^_5�\�Ѫ=����Ú,r�����hE�";)/�#`���h���G��oZf�,,n�[1 �87�v$|�`�'�h�(��96u����Ğ�H�;v���MD�Y�54�D��6�Ů�-�3x��R�n+����&����%_x�(��5�2���q�e�W˷�ҿ;(	�G�q�lSD������h���zrRZ� ���ç�P�����@wAIx�ȇȨl!J���<�L8�Jl���ULLR�ha������X�=�5
�wV9�s� ���7+�w�KoC�ڽ�%=յ ��C�*|�x�GmMo�~��c�<0��L_P�#r"���,h��;:�h�Rѣ��yyC]�F��%JoL�0��=��Ɵ깔��m�\�1&^Z��{+扽�o�A���Kx,���V B�MtZ��r���)����.��V4��p!�H�ו4V{i>������T����e]�[7�|��Q��$q��@R���g�X�8ɸ'�T�P�S�/��G�K��'o�����c�;:�	O�s� i^m3r�>.�Z��r����܌)b�Z�������Q�5��g�������!T��b���:t4���Iz>�=�%�n�V������q�ӶW�'�x�:�)bn.(>5-��Cؖ@U��I�.��<7R7��i瘣��{J��)rӽC>��E��w���і~׆ѵWl��*t�L}z�*m�b�ǅ�[oDrnx�2�$������\��Cǔ���N.��2-"��d�h���nx6���%�g���sӣ����o�<�e��a[���6�ہ�֡~�L��ٺ�u�\>
��9ڧ���?R�ɐV� -�݆N�����2F�����Z��V��mܽY����2&RF�hjQ�)Z��:ʩ��JЧ�)�ޤX��^�]d�� ��q���Ne�v����ca�U:Pp<1�&���4#�}u���F���.�p֒����!���i����DnoU��R�oDz�7#DES�
����{�e�j�v�۫��Uk�C�٤�=?ÅC�Ԉ����O,T�ιy����H�)�i+qV�`٢I���PW}SQ�0!�o����5~%)+C@q��5c$ԣe�?n1��m��TY++��FNJܾ5mS^�X�c^���f1j�;V3��4�� �ź7Η�%�W�:��a������^�N�ر���G�L��L��m�Y�	�=��4�=���0���lP�[$�W.����-{���Ȅ$H��^��+O�x��4���R@w���?�E����t]7)�vNp�@�����)�T8H��H+��T�K�l���}���N�Ep��n`o|�q��ݢ� I�SCA%͜+��m�%[���wH���*��^?�4�Uy��;��5z
�!g��%J��(l<�.�x:���(�7 E7�N���z���9�3@������mO��
zBsX�<$_�FKw%.��R� qu��e��{_�(�N���H��-��G�7~��y���9v����/�{RER���L?c¤��Y��G�ú�@Yp��9�����1.i�A�z�ؘo�ұ{�A�#�k��:�� �[qr� �R�U�踹�Ō�UC�aTemlܷ: �p���1h�L�ޅ=E�`�6�u}|&�*��0����i��u������2$�[t�6>ERc�C9UT�@����g<id��|�0��R�1#����;�m��Q�����Z�1�kcv����OWӌ�A������;#�i*�ւ>/�J�L��:�Ǿxd���0(b!EFW�^#�Wxqg�g��T����ɏ��|nP��ǚSh����Us�BF1���z4�`�<\4�hV�M.�NEa�ğ�)�d��k>����JkK��h)��b%�M9㻲=�B̑�����+x}!]�d���t!Ї�o�4�*�R���Ռ1~>-��Y(�����=�=��.�8���71F;�I�l)l��vY���(O���Y�>~�y(��,P).[x�5u&Ӂ�l$�d��WyO5!��,]�8ɦ�an�AqGk�.?]{�٬j���x�}54r�2B�˯_窖�kO��1��SG��q٠�e�HEs����L�Y <�GvF(`�~�p�9c���6��p!���+��;�2����GpVa��u����X��(�x4*�CWgSފ���T��ew�TyQ1 y͗w|�Ջ�INՊ�c��t���ůi�Fբ���#�N�����\�1�����D ��G�-4�Zn2Pt���R�nµ�J�KB�7JRP���(\-G)�EX�鍪�LJ�m��F��x'I�4��ä	�K���9��^H���10����Vq�JSW#iƹV�+S��4���s��n�d���	� �꘧ `�4�%�:�IB��E"�xq t��~��WI���Ro�S���X�\����:|��7za�����`apU� 	�p�Q[�1u���}ttoO�V�"D�=���~�����s�)Z'�[��D�ක�ީBF�>��^��ӑ6��}��H�j�������k��\��ݝ=���8Y�@f�x��T۞&$t�hçkd�r���rwCA�0��P}o�eaԳz<nȳ�Q�~@�=w��n"��c؄�l;{��7l�Ͳ����<��Clm�����MV��$���NM8���Q�Y����*��'��+�3װhG�
̒ѷ/NxV��e׸),2(h����TG>�W���R���uY�nн�<K�s�Y3��.�%A�����Ě�Z��1/�`�yH%�LlOs�ڨvp�#$fƄ���K��"�%�ǘ��5xo�&7�R���7�'��X!a�a�/���s�w8a.��O-��X7P�����x�ɕ$�2^,E����/0��q�Ď��n�_N3��ݲ����Š�V�>cl"�*�{�J�q�U������.I�a�Re�RTW�'Q�H�id��om��M@�i#A�ᨒ�g��^�31t+앯��C5g�)�����.ƪ���4���ݘWǆ1`��!�ы�FJ�3�f�y�'dҘ6=�L%+�e>H�k��*�B��%]�U��� ��%�j7�'��p��N��-�Y����fO�l��ϋ���)������T���S!."����T�I���T�����j�'t��ymuE{H�x` Ǌ^���e��V7{�!��#e��4��ͱ6�FV�g{%r��|��^'�x����ȹ��9��Q�Β:p{��*͆i�����e^�Age[�K� �9$	w�a��
t�~��*�˂���U?X��/�ƻ�la��y7��-�Xm���h��h����FHb�s�͞g�r_�&�~���$SUnY90}����ǲ���4:�d3�ݭ=O�Vj�����oʡ<�����X���rz"�6��^�xz� ��$5ç8,X��M��vau�I{���gWر�� ���fГ���B�t��-=j��Is�WN�>��]�n�C��Sќ�>�2���T����{<	Fa;7������0� ��]?�'"|���+�b�I����<+9]��r�e�L"^'�[�L�_a%g��:6�M�����Q�Ŋc���)~�Q�6ŚOr"��m��)g�hR7`<�l��2%�1��������S�Ц,�Ң��Y�he���e@�7y'�&A������>���_N+�{���XD����j�_l��֞xa�E�aD��>��m��=���B5u1�yt�;�}8>�[�n�[y�d��MB�.���e�ۅ7$����x�}���wD6�5�*���Q�2膮1j*�9LTMH�A�	�,fh\)%n�bXm)0^�r������lMB=ay�@MDh�&�Q]GQ�������eCު�&����d��*����@�����8AKN�J�[��3]&� �PH�c)v��Y�����)c�kQɠ]� r�?�&1����v���I�C�Isz��o�k/$q�#r��OIS*��,���a��^Gn,�/�W�t��9Z�|8������mmٮ��!�ӊ��X%��S��,��=�uv�k�]~_c�B���'���� ��V/��Q�g�ɖ}���¬h�R�c6a0Bʣ�z�9��? 7���ż�\�;#�j<1e`��۽��di=����k�|�}E�����<WW(1�^��0�_<���TH(cT�v�r��8�D�F�.���c�2?}��I��:���fG�p%�Ҝ����1H�`7��n��
��ٟ����}�B����y�3O΋M�_:�'b��;ƿM�#!�^�	��戔ᚣ:��K�<��;A��1�>h�0 �U�������b�P�fuմcUy���.�'�07�,�@ˑ��������\(dW�`��(�U{�.������>�ב(�1��o��v`�JK�V �S'6%7ntU�NuF*�r`"���Z���Z=w?mVg��6@�%œO4�d+�����ʒ'��6�x�Lw�V�πT#��B������� ��kD����@�g��&>�ҽCd욀A�f�qEZ�=R��1}k����C��8�$���S��G*stDtڇA�
/NQ0d�i*����yP4�?�L����ӸR���a\��71+��9Y0��u~�jd���O� �����Tb��F�4�p��{���ML�����9��(�p[���3
��F͔Z*��/���wf�5g�*�dJ���A�DKV�����#K�@�T�|���I�_��؎̦�N�E�d#K�/м8
K\:�1v�԰����:�!���d�}�Q��BH�,4�}���'"X!��mLF}y�O
 �NDK�c�;)��v���"m�P��`8FE#��N*L��j�u��}a3�i��0�)� ֍Њg3�, rO���KL�j����5�E�����4����/U�=j�酆�==��6{;3Ub��?e�vO�	�Sf��V9���0�or���{�#S;C ?�<H!��A��@�J���F�=g�~�8.�WD�C�_�)ď.H�:�qz� ��6\�OKy��>��'_�:� ��?.�>��]쌇���*W��9ܗ�J��L7�F|��� $�K�l���4�d����,�(*��#�+����Qv�����º��%�8��@��h���-�9z���B�5��X�&soa���5<2�PT��
��#x^��ۂ���R-�w�0?c�s���[lT�R�߻b�PH�M
jx��L���E~�Z.�+C�Ώ�b���@i���v��R�P("=��oZ�{��t�@.�\�ι�G$���\�>�(y��akWA���U�+Bwz�o�R'��GIU��MM͏�M'��ثm���w0͏Z6�~2�Ym�!���ZM������� ���������ƍ�v�F3�]��lX%���&A��
���MB�������X�WG�G��]����p�n��d�R�2W�H��[�����j�O��E�ML���aI;��WrM��x,H��G˚�1Ȝ|�"�+��|#�5�D�e�~-�5Q������2� ��0���nO������\�%n��k�C�{����������]�V��R��ȳOؘl!����h���c�Ǝ��Pz�����5�m����FV/�<w�@�LA����a��	���=�Xo/� D+�`S�Bp�h_	#*F�yP����<���ۻ~�s��k�+�c|hgO��	�-���,)H�{�X�l$" ��w
~Lw����ł�#�u�-���2�ʴ���(T)����nm �b��)�p�k�u�,<Y�DP�$EcBE��$r�u�s�Vgҍ(9
P���ŘuW׼C������d�6F�4�#a����)1E�t�Q�(���h�б�(G�>Z	���^���;�W��JR/Ղ�foh�5�wa�� ��Ei�� � ��*����u{�6�5������GLQ=Ո�a��bM㠮��M8�0	���%a�nF�R:��M<�#�a>�Y�F�f����L==�ɇ
���](���͒#�d
���O'�b����)9�s�Y�ݧ���-ad��g5%Qݫ��+'��@���]E���`,�^��O^6	���y�]GhY�F�f�0����/���
�,vV�����O����:�����z�#�!�d��ʚ�#[���[y�Ԥ��AK
��7��sV�]�{�Rb�񒝜�\��2�ہ� �l$�t��J�a�Ei� �	C�l(;D�اX��*����t�zS�!X0��%��]��4jw�pĊ%�Z2��d�̦�kʯZh֑��D�2q-�(�$:	li�[z�m��kLϥiM�swX$�zN!Ī8پ���Ȭ��}��ܭl�� ����ig�5 �x'[�qƈ��n��׎���x�KF��������,g�e[�(W�m}������Y���R���QR,G>>}.G<n�qW��`��Ve|�Ih��}o��5����͠6�6��5�� �����h����ɿPL��E�B8�]/����z�����q-*��\��8���5||��eʾ�~��T�
\?���DJˇ.��lMp�Ml���d;�snd��F.���0���E�X�аj2��&�4�ν����N�e�|(����2Z>�����v�0@���X.��!,3x�"�}:� ����JP���x���L�6"pO�?��wڋ&�^�������O�k�M�'�'���F?h�1o�p���v�L}L�ĺ�CE�4R#��`��s��q���'��<�|X���-I����]_2E�Ŏ�k�B�R~�&@��ӝrA󿪃	��v[yI��8<����{K-�/��*,�m2�w�ê{��.P@��	h�+
?�Dz��in�?)]F,%h��9�5�?������lf�ǒ���O�b��L�����B�%o��&F���qJ��||o���ɡo�8�(��d�!K��f�pΕ�Bg���5�\��}>�.�phaM�j[�?�p��f����n�FZ�G;.��<��_�:1�����*b9��En��*�F��q���
t��U~� "��eVj��~��j�,�@(��/E`V ��m�N~as��R�{Tҗ	5�R�QRu=�A����a�]>H�:B�%�/�I6��b�ԕz��*����thkS~q�z�O�%�~��7�բ��.8}(J����G`��ؽv�d��&�;J"PCB��vgj�ϵ�o_�	Ȩ�16�ܹ6�Q�I��%��/Xfԯ��ׄ��f���9��ఁ�G�eo3~1���·��:9}BA�����W���!��jb(ڷ�U������E�j�)J*��N����R��t��.0h�u[�k�3��j����Oz���}'y���~	Km�*�7�� �r�0��Ox=�FE�Kج95e�>W:j%P��5�c�("_��׸��g�1�s��v/�[�b�6�˅�Qx�-1�P�EǔZs�hb��S�О0Ȳ��?(�gɥ5h�O+�����.8�!��*����b����p���2$Zw�<Ķ_:Wz��
4`_t�h=�gcD�I���}��cr�n�n߼j]�g+	gL"�u����%6~1l�FO��_qv��K|�#kWJ�n�s�"��0>"l�l�O��_���[%ж�U,Y`�Q��C#,�\����r��5�Q}_P���1H7U�2^'+�C3����z�1GW��K���fk���=o�&�vfb	=����!7}C�С�r]p!R~ogn.&��#$|���YݥK;��PG�,�s�>R+}����D��=��UxF��@u9}�e���Ml��C����Q����e���nnim�����. �T!��bNɰ��$��@��l�$���]z��(%��ڙ)j����,���|�Kֳ���p'�}ɀ��������2F9STn�!���Z;�дG�Mh'�n�C�%A���gY��d;# J���F�
�"s ���8�Ry��j�].�4� q�$�*����ׁ���8JX�L��֫\�~�L h��iR���h�b����'������X�*8y��ߚ�T�Ι��#��~c�D�p&w�Z.�&)p�㿣���p�)�?B��Q�n��:�R��a�V��G���h���p�A��;6έ@۬2�#Ө{�w�K�FW.DhY+*����ѝ����1��*h��Fy���"�F噯�����J�(R��y�*Q���FE������v+��_6�������6�\������m%��n.ʳ�Q�H
��MP��b���_�<�� N�;���b^YN��Ɠr�ڵ��b_�T��m�wE4,Vȹ��x��!t��H���$�I��6���-l� w~�$�
ͮ����_v �Em�N*d�">
����8�8۪�M�_ ��������|΂��f�6����|
����ө	#[]������X��J)��#��ѧ��k���w�W�ܒO^������Բyt�����{�>��؈NwS�'���1r_'?| �5%�g���[�h�v�k�JTG���wa�:'"��p��Î�@^i�R&a�Q�\^
G�F��8�g�V�>	�Q�go&N��;�>Σj�1���A$�o��n�����'������:�퓗��:C��ǩ=.��D���,�%]C	�x��X�<B�tUL���Nx�<���^L&|r�Mn�[����B!��j�ձp�-*-(K�h�@���ಱP����+p�w�^dŢc1)��֤�e�e���C�($����j��"r��ko�h�6���?�[~k�HN��3݌��L����y��q2l���Avlm���������ERZ��R-���l��p'YfsO�	>������>���B����#*m�I�㴕*ԩ%�;����=9Q�5/�yi�sq����3�k-K+�s��
s��C��6m��&B�6�#�j���	�[�N�C��A][C�ѭ$�Z�+��d[u`{ +��؋)��{���� �\`��훶@�����̘ZF�� ��)�Y�5��Y`˰h��ó�R�<����&����H_7h��Q�;����r$-b�_�Xa�|l*�&�O���źgx�"jnQ��P�Y�Q��,kPjα�����$r�F����*�,x��AsxJb�'�'_�)m��a�er���P6B�m�bDm/HT�k�]��2/��\&��'�E�A�Y�d��Đ5�B���~���ж؅��u[�33�vRX���������%�n�m%���k�j$�����Dr�m�}Z⿓�r�5l��Nqx�,����_�����h�Jo�t1�e��Ο�R_�<x��,�Tф�����,	7���˶�%��>��H�_��F�u��gdg��p5�N�-3�W_�Tl�U�6v��*����T�=�M�,��DQ*��B5u~<;������Tx�~Y�4d�Ҵ��H�|?{5
 c5?��T�k�g�PcRM}�(+�IboГ��mX�l?���J>N����$&��1�Ծ�/K�{�u������v�Ns�7Q�w��F��sG�}Aʵ�	
�/;��և��|���IΒx�����3,�*'�M�c����c�~Fm�P%_1G� ���-I7�rU�#0��_���X���d�\>3�I��nY �7���/w<���Һ0es�e^����g��N �S��\�������~}	���j�a3b
[�g~Ì���[�e��i�!��_DBWW�k�����R�j���.񱊨`Xa�
� �7���i�����i���	�޽�Ĕ	!��/A��:�Sr$��UPI��nW��a��)y��Z�U�եrX3JGA�
E������LW�li�<S-�kG� U�.�@Al��As�Q�Kz�|8��0�e���P�Y�[{��H�^P,�D�V�h��OV[>V?��{0��=�X՜y�A��*��Zφ�@��~9f0�_zX���YA�S.���,Q�lO|�u�4_O���$�QNj��=��d��e�_n� �d�Sx#RM_a�>��KV�4{V oko{�t�L����ޡ��]A�7G��Z��S�,y�>��Q����O~���1bmP;�o�	"&|`A��S���v�z�����R G(�˶��� y�U�"�.h�^�P5����� l��]�BΛ"�����EX(�h�%��f��
h�y��ߓ65ז�+d�a�H��W�-��H���)�v]�}�}Mt4k��w�%v�G��^�.F]�>�͵������ewWp֏UvO��E��^MtB���`��]�Y�9_�(�T�N��s�_��aL�\3-?�6s�ɺL]8��Y(�u�G��_NS��C�G��!'��Vzm��[�˼3��O��a�[�I��E��\�RŅ�R�T��v����A�e΢#�B��#����YYn�_�[�,:�L���.27��'FUO��R=����V��1` I��KnNQJX��U�U���S�fҎ�y�3Oc3�U0��sh	=��XVqK0�F��{�1䟣��O��JH3�
M�P��R�.��npw���8��^Bk��7Z�D#�ڛ����t�c�1Ѡ|-��X��~�x�#͛x�}TS�����|Dyu���I��WFQ63��/7=������������P��O�~j�!uHzыiA��e�N*��x���z=K�oNWR�/pʆv�mQa��x�|av�����B�8� "����S�[	Տ����r=X׷wiˠ12'������(��4Т8N�K��
�A��z��(��FV��a�Ϟ����tZXd{����<�Z��}��Ơ�xS ��tC���t�u U��3{��c���6O�JK�DE���b1N=�����B5�d���g5�&Ү��Ku �� Ğ��mD��G��L�!ϺBҀ��ź��^���H��\�{%92�熢�~�D�8��fPgj?��m��n�Ǝ;@��|TAT��žA���K���C�26�mm��CRpCrzP�1���l��� ��!S
�=.9�����Tw���$�S@��Q��c����n�I)�:@�<�Q�s�m��W��5��3�U����0]�A�r�j��i�t�	���&�T��~2]Mqh�1:���=ع�cc�-�_Nܕk�v���$����~��03�}�J(PV����v �"M�o�m<���+�+Ҧ�-3V+���� an��k�K�;�A����x���I���6����U�:�ݩ�md�V=�^�#l0�H�~��OʼuB��Ir5�=}�*F�Gn���h�]�w�
 ����дE��>}�2��e�Q*D�!xM ��)�5�I��$ ]D�p�55��8�?�����-;L��:�Dg�!"+��bZ�@�z�SE�/z��?7�c�z����sՏ��,�B�Y!��#Yz��⿴T��'� v�oĝ��j���\l��p��4�Z��v�6:s��+܂�V%�KR�׸=-~�֒10g1��`�ia@�N����&s�pwzdkG���mƖ��}ʼ�[�Yz��>�ӆL���8�kꃁ��&q��G�r2�z΢��q��\�Z&�<�&0�/�Z��u�+�ʌ�b�L?�}x�݊9����M^p����'�1Mxn�k\7���:Ȓ��D�,������ǥ�4d��{�/��Ļ�r%�:��`�&J_g��\3��f�=������i⭸�[�d��E��~n�-i��q%��ݩ�#o��NV�`��<�Z�Z��g��Z,�hOb�a�~p����0��.;G�� ��)Uq��r�u^���g�Ӟ�Cϫ�8�;F��*��Z�&R���#��c�� V7�s��W��7�b�W�/l��0l��P�M(�������{���sR��o������'M�׾�f�:,*�!�yf�m��Nl7� Dip�{�]��>��н�n]����ۺ("أ~�j�ً�(%�L�����Q(�	݀�oBRa\{����A�:(>���P�5EQ�k�u��G�}�[&��D%6����&O�Z?U�\�mB���;��T9 �74����,���eP.t��ݱ�m����؛��v-�/i�����c���0H�|爳�������ɫHٶ@��J��O^��|�d�Qy%���$'����^�]��q��^?Z䡴�<�����
���f`ɋ�����]u5��C��;4�p��Vo�%��*]�F�rY}�"��ܜ�������������\���5q�ߧ� ��k�4<��D���|�=�l	��^_��P����>��a���o�rRD�}�ԭ+�� T?�x�-4�`���!~��Z��V��u]���_�
7z�l��	3���F��t�H��J*�Z �����)3pkXH�+a�R�BQmn��Yp[���Rk�]�ߵB����G]�<��)�G&�t��?�X�X��0�Orq�\�+Z��_���WEg^>�U�[�c[��?A�Q�h�B,��{ږ����1��L=|�n��1��hW�\��#D��s�2n��%g2�`�~Ś�=V�O&���ِ���:^��UWR�˳�/��㵚����bHf��E�L�ťʗ�+���S"����H�Ky���X�A����4�`>���$�Γ�B��4F}��u�w�c�i�����R���6����yc�h@�%�����Ǿ�6��\&�����OD~�Y�I�d�J	�]���	��z��������KB������O��a�vL����W� �7���r�]�ye�GX��[s*����c�uZ"l����ڜ��?
����pa�����
�R��ň��t w&�L]��?XbQ �����G!�nvm�X�;-��i0-ƝH>"Y�X,�?�X�y[�~��O²hF��ϥXKI���T�-l���p��P]]!Gl��w�NVT\U�Q���t�Z�a��Gp�ű��J���f���QĀ�I |j��E�]S�4u��1��;9��s��NE-%7Y�����{��ρ�a��fiA̢�yY��G(���UZ5X�#��t�@ط <��k���.<��2�h��|�h;��s���A%��m(���|���{+�9C�a�._���_�A
Ɍ��!�?}�c`�K_A>)���ĉ���}�S�,��2��(_A��dZJ�9�#[��"�m7Jj�c�}3�I[�?��Twt��}I��)��B0�}�jM�Z۩��i7�tZ��/ꁬ�g�$09w��w� ��� ��ipY�T.�pR����aMƛ8A\Z��6o���(u�k{��v:�Mw�5ߛaEWe2NX�E����2��7��F�>�ʒ���o�/ߧb�t� `UԂA�FՒm����H�֭ti�S�	�J"�ԑ �Y���b�톭啜|~�_Ϋ��(B߄{̲Q"g�{�A�9GU��ˣ@c 1	��so�2����h_Fd ��q�a��L��Vhp�W��x&ʊ�ɯ._I�H�Ⱥyv��W�ɭ3�V;���!G�ThB�]T������P�K7!����}9Ϳˮ�g��i�a0�ǹ�,�7Y� `�~�s�zʐP���W�H��,�]/p��ؕ��y5b�"�7��p��8X��j3S]e��I0��mA�"�^~���swW,�4�w�����8˯�2�&IM�`/�Z��}#����Sb��'n�b��]�d+ ��
Өn�������L�q���m��r����>�U�@o�'��VV�4��{`�b�XgW�ueA8E\��wҠ�8Qd����꣫Y�IKW*����d![H��X�نM�`�a^���Dߍ�	Vy(�Z�����D_�"%ps���KiMӌȂ�N�.���SOHy�`=t�24A�w��� Z* 0��ƛ�AT��W����:k�d�j��c8jI�~�D�%lI������rBGٍ2 ���i2AՂ<���PDqͬ��.�����콋k�#�7�̹pi���
_mØ�'	@K��+oO2ƘXLg6W?4���uޝ��t�)w`U9����_b��f�U�&w;�U��G�� ���I{��0����G%��]t_7�Das�B��|�:������Դ[:�/��J��)ft�L��ߤ��4�V�z��PaC|�6ޏ=���ޜv�R:nW�� ���rv(�Ş#^/�3��4������D1)�����_��8%kMƴ��[rC&��b	�A���uO�m�ރ\8��eK���E�,<_�1V�D)��z�T?BeWs�p�
���3�ʕ�����ӀY�6�-��S�?������ު~o �QIyl�^�m5w�'I�����D�R3ճ�Y
����{r�%WM�PP��G4�2!�P�_�p_�H���R��X�(l��?[��5������I[n8Y���fI�W�g/��qT"#.�0�XSa��\:�Ǒq�X��R�[�C4'Dbs�XW}n�8ӏ!���xO@��"��l�R�c���F�/� ��:0�^hlEd[��j�'�ݳ9���"B���"T/�H�?>M�P
�n&5&Ya�і�մ�h����ڔ����Hͷ<U�"t�#Z`�;2�I9;�n�F�I.F���m�/�ۂ*9Q(���x�!�(H�k,���y�"���3х����\\���RX�}	='WH �B�C�5�.%du����Z�U���������M>#�i�J8TzU���h����9.��_������5�A�LG�v��Ԛ��?fmLdFs���PV�:E�t���k��IPtybY����1��D���P:ɕ����<Y�2�W�4udE{,T������e1eeue�jD��Ũ��������i{�?7�>�	��u�.}ĩ�N��oK�O���ƪƪ2��1�5Ϯ�+̯�mߋ=��u�À��|�����/�E��y2ky�Hx5����1�Hε��L\c!��Q��5O=��K%k�zGB�j�ꏍ��]产S�;4� ����s뮃R��^_�ed��M_R��	��%L�x����&�z�b�4$�܇���7�`BB��t}E�z�Ȫ@�v���hB��`��y��Fs�V+Ӳ��������
�"��bdE<���ߤ��4����|]��ʆ�u��22k�0�ͩ@�.������@[8�x�FA��/��{�P��n����cZ�	Iv���#i�$`���������9�S�ڳc�|U�p`�t���� ��*rB֣0o�i
Q��� ��1�����_�%��S��녊���2�6ߩ�"�V��I� ����Ǖ���fDL�!��z���gɇ�*	��M�U���s�����8�p���3ϑ!ujK��i�������;�����J��i�r..Z"��~����l�`�J�������o���	�z ����{F�B頭Ԩ��i�m9An6�>^dTh�ӌf��<Ǭ~Q�ڋ�J��P� �F�t�5n+I"P��B��*wm�	z%��觝[4����}��ʮ��f�b�2g��$͠Y��
���
_a�H.��L��9�(4�946sې7��6ɽ�I�"�S��)g,<3*�;�T��X�i�y!#w#�U&��,P�Jb�~�3�S�g���KZ67��i�+��['���`k�b�v��A65�eј�X4l:�@\����r##!��U�S�9x5��%! �[k���ۑ�!��a�Q@��;�����,.u���1J��o��6܊Տ�$�l����}���:���K,�b�4NB}}h׳FX`�e����N�x����-ԋc>��$~`(���@t�Kn(]ȡ~?[���R��u5��KX�:�2A���eVޜ�"�0t�2<�]�N@۾���#���� �h��^N��=��w��_�7��`���`���V�~]��W7v���۴�Qjo�P�����y�]��PD��o�<�,t�(u7a3����<�I� ��Ur�ba����+�M=�B��&>3�� ��Dw����͞�́�`�~�uB��ϴ
��i ��(�M�|���m>�	����
��K�k.����{(H��:��eA�ɞ��bTJ�r]<��)��:/���bw��v�d�0ߔ����ΑIX/����(	ʅ�7�@�$��m��u�ƚ����*K������]�'ѽ#Y{Q�
E)	�����^���V��:}��duuݸ��t$X<QA�N��'���8w�C�>u&V�G"��߮ιo㌩��\	����[��B���8��"i�������<go���t��?�R�QK��{)�d[Ӗ�k@�J�Sݛ.�7�ةX��]l1�q3.dR5����C��<I5���L{�"���heX:ȸ�и�j�)L5�L���Ժr5�W����8&�v�R~��\�R�<#�=��>��H����>��{]^Y'�k��������	�>���\S(~.o��z���~eU6�N����Q�JI+���4KT�aw1L�:R�7��fn#��}(C���K��?��Q#÷RX��& g��΅f_>Wʐ�+�Bj�2�1.a.W7E'�+��[�1 -���5T���T�E�Q��J�2�`.�������0b%`h�Þ-�}"E��!����h�;�ϊ���ΐ\��U�$���ɞ�Q��?���$lE;r}SJ	#��#�l)�^��y#sC��zaSS.(��[ͼ�nX�=q�]�4�q�.fq<�MWQS?�+I:[��kB�����ߓh�������LT�,/�����h�14cc��m|�w�����z������#�\��q{�?��~8UP|Hk�_�K���!��e+T��n}��Bپ;���Ƭ���G�S
6�1.��X�y'
\� c����fhL�Q-s�����{��� 
����Qj�u�pQ}�`F&��1�)kg��xle?����2�Jx�.���R6�7 �u�8[ ��g,�:�Z�e�\��g���[΢k{^��D����X��� c���6�HMv���ҹt�_{/8C!+s��Z���t����2�� Ԕ�淮ʢ�ۂu3;��@r������;��vs�.��6�n� �.���7r�H�f���Px�z=2`���:����O.Bo'�@��	^N1�]`	�i��P���ED��W�~";�EA̽-�.�Qt�*v���i��n`}`yq>Nr��@������վ&'!�1R���%T��Js��+����O����y�MW���Z2�ON}g����).r��ܩ`FOh���A��X^v��N����n��uH_�����y�<x[���_{�b�J:&����ҽ�@�F5l��5͘E6L+���@�,�j����k͒�Xr�P�R��Doک��mX�Z��_w�첆N�I��zH�DG3��(PUo��D�,��W�u�����(v%^8���R�:v�w"�[$c��a2�6�l"Ld=тe����]���Z>�%�7*k �;4�D�
N�r��;]�*r&����G�1h�B�#���?�q���(G斓���j��B��@�9�4!��k�Ƥ���^s�L~;uz���V�Q|Se���!�긫��JB�$�P����F�j�K�	��
�hi՜u@ə���٧bE&�:�	����3���m�cm-]�B�`�!�8Vj�a�l���_N�}�T!z'��%*K��JU,����F��+�m�MEZ�P����2Y��"���s)}X���;�T�R�G \+n�~�G�(�溗�C����@�^W�eIs��?�S���b��ݶ�	#-V�ؐ~�����,]�&q��	C��=��WE�w⧪�@�C���^n�����'$X26�����ϯ�˚�N���	(��yo���=þ�{��L����'FR�������{St��>{�V���ΐУ�7/����(WC4B�O�.0��P��&7���&��2e���I��*�:j�p�dxc�[8����=M��V&1a�	��y�,-Y��]���;0XE��nCS���g����j���"/�~"����p'���Wȉ��+��l�I�W�|^t��WwF*�*�Ұ9:��Ļ#A��.WI�L��B=�F�8��
��=NǉM�W�H�\�#�[aA����7L�}��W��� 01c/�$��#O�gP�>�&�ۥ�?�6�ŗ�H_I�����=�t	���C��(ɗ�u#�wpSk�i1`�EaK����JJ�:�Ԯ��QD Q5��%��]�����f�mm����v^}֕�J�b��>$�����YH�a*�(�!pDW�1!bṅ.��\������|��9���e� -�:�p��T�~�����d#�4�Ce�Ֆ�@�7�s'���?ir�[��#]��t�i��������jX�� 
Muh��t�ѡ�>@��W� ��~]&���Ϲ��
�暄�J���#�)��W�_6�ϫ��Gi@�Im��+=b�3����Y��s�4s3[��������J��a�',~z��u�,�Az��z����	a'gs�4}&�	�0���Q����닛�� �8r�w��vc�GN��H/�z�Ra+Ϣp�L�Pk3auj��^��J�y%�ơ7i����{��`�Ss�?j��,N�Jx�h�n�F2����$�l��i�kWǈ�G͕��S���a���h���ޔ�2ka %�Xiot6k�w��3��}����n��;���%u��!���2E�g��(�dY�j~sV 4ØK
hu���s'������L{u/>�����$�F@�����;r��͈L���R��ñ�V߁�v�G�L���=�;G�[(.@��%ʳ��F��+��LM!X�Z�$�s�e��.7�W���wd��=��R ��؎�.�����dc�#�xOs���u��h#�|�ʸu�*z|9~_&b�p���]#��F�VW"j`��i�m���c ��y��dDA�S���tS�Z2ZRpӘ��V\���)!5]H���*���m�uo�Tj"AU���ty��V�4)Jݱ��W�Q�6K�D�C���I}m���Ht�O����Dy�v~����_�IEg=�Z)Y\g��D�#>,*��vt��c<�"q.~���c+����D�yٙ�P )�+���!ǩ'��wt�*�Ye������6����#y.��[~�����t�î�@��Fy�/�+�m�K��3:���*��R���_�dPz�;�㾒՘D,	e���P:m|���6��2�f!.�uh�m�&���/Fq���3׸
╅�/V�)Y�q�j	��{~��W\�61�h�S˂��%$ϧ����>�w��FZ.�櫞���ܿP��؍b��>yf$��#�p�7yD������\�(��v�-����[܁Zq��<�FI?\*5Տ��͙o͞�~Q���xgh�*�4��l���!�犈��<��sY�S��'ԋ[�0�\��	son��*'jj�������?�*(�����t�$����%p2g��c���Pm�'�����g��'+��P#�[Ac
������櫴����V�V�Tї{� Bt/�&�j�U��ï��T�4��u'P�MU.�6������$���x�	 �=��]�x�S~�^�T-U"�Ա�<�p@h��3��S�`�-dt�d9i҈��"ց	>�� �=b��?�F3�͟��oip���z�ڜ��8�F=��R�.JAI>S���I�s�A�Gh�eT��Ir�
��c�N�QmP��FE���r�G��8��XÊ���S��
�����'�=}�i*¾���_	�w3�΀(��ံ2���T����i��~�?�x���f��8�hՑ~5�L��'f�:�;�Iz�|��� �(�4�*)��f�	(��$\MuD�����	�s���RbN='Kv�V�$��yj���Ȼ����M�Z�T��!j��dN����b�H�f �d!�`$H���s��z�z6���L��N��������k ��w9HfN���H��V�$�,Y7�?�!��4UYc]6�U���/�H=.�M��� C�e��J���[q��d$^L/&�aW&�i�,<:�8�U�|�Πޠi�lX�����s���V�a>��|,��@�%*�3dЙ��l��'���*Xn6�)���ԕc*�e�-�����[�
9��µ�h��N����R*|1`e����9�|c�xD�T�U��z�!?��o-0y/=�b	���Wo�<A}� �q��@�	�PZ�F- 0(�W�j����IլnQ��(@N6���jj���:���$�!y������]�s����Ӈ5�{��d�[ͮMPᕢ�C��g��C̰���������24�-��vJ�)�m��=e��X������S��A��싲9���T�4	�`��x�Dc�*g"�9���P���o5�c	��L�����r �����p��3�b���[NӍ���N�Җ����4�R�ѧ�WS��z�L@b{v�e��1g иA+��q��Ӈ>�B��[� �S<�E䷇n>��̃[��OA� �a'iq*��H�"p�`ɇ��}xп4g?-B��ސ�����4%��iՙ�6�{�ݬ���_���|@�*�a��T�(C��8ӼMѺ3�%'�+/�xŵNl��q���]�"��J.#�ײ��tI�L~͓t�����d۬�Κ֯�!��I�Dn zx�g��E���.n����@(�:�M�F-Eȼ*�Bt�/{%�!�y���T��>H-�����7�D��~�v+s�}Ȁ U=��ҁ:�̜��W�D�}���B�����>�4�0w��׊��0��V���Q��gG�f��^@Ӗ()ٲ`�g��?�p�0+�&Κ�G��<C��Ǟ��d�Ms@��b����
Ш�i��1h*�%�BMe���y�Fj��u�Nxu�NĘ�'Ц�����w��N)���;`M8��q=?�)UG� �Unq��Au��ԷsF֍c����R"��R��)��4�WuI�6I��gA���D0P��v��(�
�0IS ��P��D����@��&n��iA�"�1us*9�ȡ��C�� ;�R԰W�yf�K$VH�����Q�Yr)���ʀJ�x�p����JRn�%ȡ�l���b�Ĭ��,���e�T��'|X�s���Ȳ�����璒9!lD���,�a�y��Gp�+t��R����4Xc>�W{��t1j��HP��n��3̎#���Ϙ��D���׏nIر{�U�fwgA�4�lӠ4�X�%�d�PP�}����<BHa���_\�'�O;!
;��� ڡ$�飵���	����i`=�ć���D=�0�Q
+�,0ڮ2q�T���z���;�`�;�>�]��ik��.�^WQU�/����_���������Ż��=P��!���(�!�@����T�)�t��	�t�1`�.}�.�E�U�<4�Fg�#m!N���t�F+T�l��J���H����E� q���kh �ӄe�h=2��=�3���+I��=�MW�d%a��гl�+˽`+��҃I��.n�5���}��wV�
�4��5��ɄW�?�/���U=�k��&�[�y�_Kµ9ֹ�N�z�*z9���Z��1�R,�Ĥi�3{�J���6Muø*�]�&(44����O^�i�%�I�w��y�}3�h��=E2�>���Q��z ���к����T�^@ x���𽡥�?\���Om�LX~�T23�0}�9�3�������rX��3#� %��9I�L���/����K�:�8D�S���,ӄ_�7M���FD�\��8R|�)�|��X���8XvP�3��Ö���GWPt�����b�RicG:Ԍ߳���I��~���U�1÷y̾�Fm�;q�z?W`��ڷ>	��Z:�1�[����&��}���N�?���M69k-���M<j&�8J1N��z>��M���4�JW�L���`��^ױ½vA�㢒V<�EPb�6�k�!��q��&Hyȴ#�p���f��W�ӂ��ؐƽ��d('"7�|A.�p��,]�F���|��l���C���|�e��Mm�|��<�t٩i���$xp��C�<o�j��,�T���;��_u��T,P��fP���O����������[k-�sztYy�%��Q�M��p	O5��IaW���n�l-�{��.��	i�f(<g�s��;$C,������N�&dc�}���N����vm�G�8N�C�IMe�6�6s���[I|TY��I���K)wk$J�=���+�3�i�q8ȵ��[�h$D4���|�Ů9*��`�3�a���svLn��<6@�N��c
E/�)K��� 3�E��
@,i"�(����N�/\�Pj���J�_ՙt���)���O��Z���/I&����X��SS�l�qx��f��ft������q�`����8��p �v���n��I,�Z��`�I�o�K�m�ĚL#
�@���2_dp�?H�[���@�U'@�+
c�0e�ya�Vh�!��g,����D9��R�(��(�Z�`�8��F������������p����� E�ߓ4�~����\~U+J��W�$ܵF���� �Mb=��l��4А�(�5����/�!{o�p9K32�3��R>��3�^���raJ���Y1
���IF�cW��ϵ���3��?�����%�V���z�d��>C���.�����1?aq��M#8�k�,���C݇ȐW-;��[4�$�R);�e��){�V��i¸��٤SSW�����9W�`̧��Q���ep�b4���_ $�������g���Љ�Bo�1�~�A4�R}�:��_v"#����?�v�G{��dZ3���2�ǰ���>/F�x (C|#w���+d�כ6=���uL�^"�fȄ��Y`�ӭ+PP���Qo�X���p�p��@���w(�����?ʁ"��n#��߳m��{���R��ޜW���	dz
^n����`Ź.{ FHW�0_�i�.)�U����\ʹ��of^O��+^LPqϛ���@����(5�]�\h��AU��{ou{��DOj�V�~�Υ ɘ��賞�/M1��(�pW >+_��!ŉ�w~����-��]_��	��*�uf����s��3�A�3�+mL�7I�#��sZy��FI�.�y�X�e�0FLމTQ���������7µ"G?�,�P��.��k�]��	\���ط�C��d�A��f0���6V����z�#��OyõXAZ�^
0�K�ݹ�c���� �������("�{�?ɸ2��� �;E�O�C�ь��p��L0�ۡ`|ig���{^Df��SbD�2�o����KN3L��,��:.p�	�� �M�7��1�ɽ��]�*�IV��IB&�>�@w���&��Fx�H��ڐ�ʦ��t�|Ah��t�@�蜇���y� ��o���In��Ʒ 2����y��Ɲ��EnN�p��a����?������2i�G�H��z��$!�K���)�Pݻ�j�v)?I��2�UR��6>&C�?�F�<؄'��N�������w�[��	��e��4��ޑF�}s8\���cJ��K��6�de��{���R�vיz W�$F���bM�?cHW9w�f�����>X��,7��8��W�6�?�K]�%'�^���M@<fB���U����ɑ�+�Lz)C����(iЉ�C�<-e/carÛB�j��籙_��CH5WP.)*����Q-��(�s����Cy����G=���J�,� �6�����+���s��Y�|0��P������\:>$�*
K��&�腆�pg�#O����\A5=����v���5Y����m襳
.��=�t��G����وۻ?�A=���
)�	�7��&��D&���f��6��u��H���a�28)�����Gy�LNb  ��#C4U6�`*�/�B�ue'�s�iO�N��5���L2B���uG)�RA}ǆo��˘(�I�_b%D}���ӄ<���������ۡG���jor�G�X�M}9�$�m�\��o�QeU��� �a��8��!F�I�ƙ�J!��Zqu��"˃d���=�n�L�<H|���) ������H(��Y��-�L��qJ �W��r�\X	���p����x�e��@2�6߶C���ES�# `P�_D5���w#W��^aH�ƞ��Rp�Oj�sBg�N�P��*�7U+ƒe�R�=�J|$C�Uh��w��/u}�@��7��,��A���GN���=�(e�*��I]-dD��I P{��y�t�xh?b�y��.��7��UqY?��=X7|����k�S�
�>Ȏ�J�nï!�MGw�.K9�z؟R�
�%YY����LF�������XW�v����&�1dog[ڠ['��gP�m֐�ʊ��m��}�� ^��S�v����:��l޼�9a?��*� ��:v֣�dg���zڗ<�
�9�.�Y��̛�]�&;�+����b%uK�E5������?�lnӨ�').�B�W��vRԴ�
mU��yF����*�`���;zJ��1�#F毉�#���g���{�hb��"�V�ICo���Q�(�p�����1$[��g���� ���D�@�X�^���}���Ў�wZk8��}B)X^��/H�b�L",\�R�廓/�иr�P�~��*�(p��t����ͷoF�Q�0k���mG^#+�� տ�)4qt�`����=�Dg�q�3�qZH3�w#���
1��}̴�&N'�|pj�R_4���Ǒ��P�`T\�\yQ�ɫ�:�Ɍ�J��v�j>y,�:u�Wg�;�%�۴�sDS,�x�$Ԍ���T�i������g@��k�
�E�+ ~�v���R�B��WW�=ܶ��D��Վv,�#��>��f�x/r�`>:�WI��$я�=��]�����̶]�?��9<�@
�({��Zm	!�����H���Tu���
96	Lj+h�4W�m;
nS������O�̡yN؝��Oh�ɴ�\���e�	/7���� g�=T׶e�֚��i��J�+��ױ�9��\���$��J7ok�!��]b<�8�$�b��Ã᧑��E�xhܹqx��7Ѐ%���8�S�P��ٙ�@Ʊ�%�|q�����γlf$A(�R�X!;WZ��
�Ʊ-~6,k{��u᤽l�[����"5�m씮?��PD	�tk���\ 2��*iֳc��ӗ�+��L�|�k"��L�<�0�j��~j$�%�V5AY���]�j�;cB���2����C$ݞoM���+<�Y3�+��U�N�Nlgx�@��wt��vh�+�$au%Uϕss�dn�O	�R'P��bKž�jY��_��U���d�5������`e( 8�WN'�)d�2+��/y�R��J͊��$�nL�cm%tڱ�p
 ��'�0��n���X���&H�M��p���) �"s�>�A���YI��� �?���͍\^Th�=��*�W�Y�z�~\K�wkꍓ�Q�Rk�h<&���q<�O�{����Ed�j���*�Zq��a�ڃ�5P�Yd�6�R�w�0z*���@,����s����d�RF�L�]$tJ��'3�\+�>�j�����V$e�UTS�S������`�~������V��0��B����������H��*�]w7_�S���-�B�b������B�BumN-6G���y�O�i����WV�(���d�CLPB@DfFn� �"��uK_:����X����2N�_h�&*�1���NQ�<��']$?�5�ri�Ju�ӈ&��l�4/��gôa ��N����N1��y�Oo'�x�/Jc[:�aA�e���y���:���pj�3���xGW����(�ͻ�������a���QcB{���|Յ١_k'`�8��vH�Q�I����29F˕�ol�a� q6F�d#}�QX�wuc�٧F�o ���x�é�@���狣r;�x��2���J�㓡��%���F�B鸆^�{k+��>f�p�8iOE���}}h�*Jj�j��άP�����ƺ�9� BʚW0ap�Sa��|��_5ؼ;au�G��}�rW!����MbVSn9��f�����Gb
lV��(�d��\�+k�,YE��� �Jh�2|��ڗa"�l�b��'��i��TeN$��.�ДWY��?�-��nc��,�iF0I�f@�C@u���Ȝ!�J�N���1_���֞9,�Rװ��~��ė��� `�f�!�l��SRY�v�h�a,�c*ר�G�iQ���&e��K�R�o2�Rl9C,��Cc*�Z߽�����I���L ��m&착��)�}�Z�X໻mEW����#�x$7n���)&/Ww 馨r�!��>z0�*
nF�+���NpO��z�,����i8�{~�o��*Et����	�Х!_�H��R`z� ��Q��}��9 ��p��r��=����) [H��ҝ��3\`�h�Tk����Z�Y�fZ}/���E28	�0�ou�܉�`^N(l_Tч��4�_D#�
?F/����q��� 
jw����I�}.��?�S>���J1\���u�5R,�������Y۽��X�qNǓ��>$�^�p�z�x	a�!�3�l��I��3�*�*�b�J�ɫ�%-�l��K���<Ma/��ȱ��!i<�P�%RB��TgR
�r�� ֜�l�U���7��������ioz7��Ka4���mB���,q��eDpt�g�e5"��yD�* iM+�H)������
�����i�[T+�}�"5[
4�����<�,����J�Ĳ�p��fvj�2V{��#����>]�	�L8E���ר��J$^�w]���������Ј��5]�<d����P��A�NeʗҜ�� ���%6˩w��韒�N���]ף�x���w	�l��rb�FF�l�9nӳգO��0�D�ް	b�M����\<�f��CuC��X։���(i8��6H��=Ks�n��gl��R\�@sh�QZ��u� d���V����rW�e>��!i�,h��������S���:������y��Q�6��b(z6!�������7�7S��n�U;7�D/����������;��j����VN����-�;�C��촉���,$�y��?�f��p��2$:��MB(��c��O�+�ŋ%�r7��0��r�&�g��O��Ϻ�����q���������i�!X4&�m^z����5��\P�֨�?~v��:��� Tq C�7C�A�f�Xt���C���Xۡ�']���,�\	���\����jNX��&��|�j��=��T�y)H�c�������Bp��^f�\�LN����3�x�7)$�cqhv�p�h�XpĶ���{�Y�����[�˘��kaX��4q+fK%��	*Bҁ?��>j.���p�n ��U��И�06�3�u��0 �I�P�]���cW�)�����G�,
]E�A)rJܕ*.=����}	���9|�%���#ă��C�Hx}��5��]�:/g�+��ƃ�������[�.��cv5��% R[1�)��PI2��Ӱ#�<���z����c%��Wqc�W�Hp�T�ʲ��8j��pNoj���Qr�6��q��wx�Hx���~�k�_IB��0uµ7�~ob�o�I����#B�Κ��ߣ �x꼖|����-�	�]��hW��JAZW�nC�����{�'޷\,�T42&��M�Hȸ=qhWh���d�AO*�����h%�fW��!F��	����a�� Krv�pP�[���-�����7(K�R���U�0�"�h���o��@���p]"9���6���B�$J��v�*���$e�c�C�z�ƌ	_�)����恑/?�32.W�uX	p_Y ��o��L��:�w��H(d��{&JU2Nc��X�@\�yaU\�j�F,�~�4P7fϏ��D(7�%d� �D$�����̪�!�$�qfE�x�$A��K<A���I�Aײ��ED�o��:X�s���;���2�~+�~Lǂ��<�e��Aʉƞ{$X-3��[���h��ui�N�I���}���u|�[s& c��G���������!�U�G�MӇ `��|}��_0��|�I�fC�FD{3F����c��t����D]Ut�U%p��8aAC�����{eS��aML��>��$:O�iL�s��_*iKg�L���7�N��cݖƊ�YS0>i@�+�hG��\��lL�?;�y�����Aޥ�"V�.Z�s�n�*����>��y(�Rsd*^�]A��&���:ed��Op� Ǧ}�l��~�J�{w�#����.�����"(�������K��Ԑ�EgϽ�к2�� y~�RW�K=#k[Tͷ�M�.�D���8�s�p	n'G�E���x�G�9�˧c��2�ّ�Y�!w	�H�1%L�`i�T��:����� �+��=bN�b�(k�ލ"[DC�b���窮l��Yoͼ��$3�%\�����Y�����<�@��V�PY��0����wp�m�@�:��S��r�,L@��3��Qj��1�uJW�������
�k�r�ƵH�]��v��Z��0�b��5GN��f����χ�A%����\Xs�bܭ�T��V/�di�W-�YÁ�w�3e끒�&Q#��P�(�0(/CpҌ(���TxN~�x�4�;��I�X��'X�"�366�	}YȒR�N8�Ju�B-���hX�	ƻ6�k� � �l��M��V�������	ߌb���zU��L=��r��,xa������j-��Z3s�6:iCQ�ULb�`z���w�[������W��u#з�$5���)jl��\�|Ńk8��3%g��ئ�"����h~�L�eWT�0-��X%t0��e���!�ףٵ)��m��ސ���03�o�Q�gz��W�%řM���������ǀ�b�
> oP}bU����MJ�T�_�NZxf�{���*�*�1g>qu}��a���1.�,���5:��I%��Z�V|��ŕ���X�N�(�b�3d�qɊ#0���$�W	�anEf�8*�����5�*��1дH�J��*V\0KDGOD}�K�#f����h���~ճ�����<��?�eV�v���M,�}u�4���m ��v�������W)cP��M��$�q%��x�:j|�DcK��z׵s�ߋ�����D�c�3�=��Rv}��U��U�I�%0#�)o��I'z����S0ض��\��N��9���A9��_v�%�����MDq�/��u8`L���Buļ�ʂ�����Aym��	�:Sf,,��#\*h�dijU�P@ �sJ����k]�H$��0�=�c��y���6?���[�п�iS�ꋇ&H�{M�J�����a$�ã~�/c���Vy�案!r�Nr��d�0ּ��?��ƍ��V�q>���L��%'������w))	�C%�sHX��5i8n�׆9�7ʨi�!D�� e5ˍ^aS$���_����ڀ�i�#�:�AR�Wp���ɑ���o��oa	�v���	̷= X��z�y�˘.��I\�kk_õ�X�����.ڰ���Xf����z� �P}�2'���xo�L)�3�3�q��;���d@B��e���׽ 3�S�ؽ����9�槗�+I:�1t<��ұ�����z��K�ђ��{nϵ3mp����E_���_��Ηf\��S��8�k����1<�=��P�-� 0���6�*��u\�8/]w�٘���pɡ�Z9ª��U�4�I7�i֖��t[k)k��w$4ăA�*Y�g[���$��|>���k����E+�8o�cn���*Ur���]��)[��0���$�c��ɐ�J=�[a0ت
mM�r������b�FH���L�t������9��ll�(USm���щݽiʄ9��K�x̬������xMS��O3l~ ��4n�4{2�\O���G��Zݯ���J�ņ�3�D�D������O�w]{������~��{��*ou	�*�m����m��0v^,S��l�\4����}Wlf��
&u����qA�7����d��L�,(��|I��7��e�$����ؚ�?�¸��#k����L*mWIx�u�l5��f}V��K{Q紗K����V����ӂۅh v�����39�)-�VP/i����Y-#{9;����e^n���{�_���ę�'��⹦s�}��.����.��9?�S�Yēex�xG��d��3�w�X���3���^P/�e����+�����r�֤�����:��hHXм쎂q?pw�/�3A.��`R3W���G�y3�lO�41��#`����8ZQ���R�������ri$n�\���g'���	l�B�c݅�M�Q,_���9�+�B�ux.Ͱ/�!BeUo�肝Z�\&�<8���J�C ��pY�Br<A�����c�����5�'=��>��
E��&������l/�e��=<ߡ|���L��w����gO�׵�]d:��W���aY_���ސ�y�e_��_`rmd��S�o���NP�Т)=�'$��Թ�,ۛX����~���]�5�E��0^�=���i�5+�|	��ZS��M/���� �|u�Ez&W��G��w��l{*��^ᒮ̧K�9i�����S�&~¸���C֩ڨw�>���!�Q���+�}n,�=��Rj�P�W�?	��򘥮I�Z~�w8����z����	�X?�nr��'�N���m�25��Y��U��3d�>�<ֺڈ��C�opmf4�O��H�+cR�;}z���=_��L��\�y���򢘪��g���*	��ͨ���n�H��
��-�i�^��G>H�NE��N��D,��m놞�ܮt"jH���x̵5F�����!MFF�ao0������x���}����~�i�!@�1
��/�`n/���&bFo��KD��9��˦�..�Y�R���ee�o+����	��E�f��EȦ�;�8�E����=H��N����h�3�K{���*��T����Ŕi'ȸ
O��.�WbM��I!��Jx3�����j�@��|ǽ~Ux��U�C �B�5�%T���y�<�]ܡv��!ѥ�_�y|`ʽ�K�~��d�8�T{���G��[z��'vx��#���^�+�5��%�f?�ziJ��	�+x��
�%T��� ��F����#��O�W(r����&
a��l	.��h�ƣ������h���w�P8�d���~.~�T�Ǹ���K�fŨ�ج���}\Ĺ���~�Q���3R�
	=ި�LIk�F�r&O���FH�@�$��34ʤG$[�"�9�שׁ��F��ſDh�ŋՍ*(YN_�bH��޵���o��2����>Zݝ�4�sC�Cm���\�'J���&�Z��l����?R�y�mh�'��:G�&`,�4h��1��o�f�M�fr�XKF��*_.;�P��D/���t|nz�Qu�q�Q:�g��E���J؝z$݊��j9�RD�.���_���r���pe"]I_=�L��r�4;|sk��иǖ�xNcA@�|��G���؈X�
{8�z�ϟ}�B��~ڹ�략rK�_��Ҽ����K��q��a~q(���ׇ
�Nl�b*��R� _�F���Z�g'fqI�jf�S%$:���P����L��)/jq�۳W~�cO��D��]�2�kr �	�q�»?ن���9��pz�������|U��ϷX?�v�Å:� �b�d����������Jk�i{E��6�F��n�D5@_8��Q$�A�1= ;����}��Ӝ�)��_6/;�r5�d��B���k���?�ʙ��׷�,j�cId!�J��?�E�5�tO�}���b�5��� ��V�{���P��H�����6Kfհ+��᧴��L�ϺS�-%�J;Hv�E���޻�Ke?�=�/�ņ���<����T��6�"�A|kld�����Nr�ǧv�|�aI�K�/�D�
Z�06��i��$��f�^�3��U����w&�i�*���<��~��i��Y���n�9ViC|�˘� l�B��Gc�\I&&8\�=����2�P���$z�TU�X������J�sɀvuA�rB`��B&F��p�a�jQn��ђ�p�<��D@N��_à�+|��������Ugj�9�ky؛�;�=�.�^s�ŗ��-�)uԟ�z�1Y0�x7u��&H��DyY7[^�y�#�������qX[��B��M��[�i�s���!����K��oNpu��P7��<�x�H��w�-���_�pr��q��؜%�5���|��o)1�Zf,�}���v���B{c�];�-&@d�|��AUwN!Q<�<���;~rA�^
@�/R���šy�	�a��x�Wll���+�-�:A*\�x�$8�@����K�K?������
pl;w��v��-z��G� auPDL-������-�q(}����g��2L�]���_�@?�Z�XF��n�r����}����'ޥXv�q�h+6�%����ۘ�`8��x��"��5}�`ls��j�¨�	[��R�Tr7�H�0��|#�H���ظVw_�O�X��<d����8��d/�3� ��������o%r)C��$���<$�]&�r��{���d��/̼u��E[<�#�Y��HS��Ȗ0/�ԗ��rhX"s���1ō&1��Jcޤ#M�DF��'�K��d���jA3�P�vOǻ�����Հ��A�kx����^��߻7H�}J�Ρ����l,���$v0�Z���s���^iLL�J-��L�7�� ���{���N@/�y��'�q5h�v%�J���)�(�8�U����p�VBD���? �=�ˎpt�����E�
�r��F�Z�:JFm^��^=��W^�哇}B��k]��2�Xħ�=#�(Y�����dd�Ws�b�fb_�@DE����ؿ��D�ƞ��$֜��gQ���,�+ a
uBV�7��C �h]VW=�"b'�Y]�i z�
_��L���^R,��2?��t�U�@޵�@+�w>Ght��}���kU|C¦\M�Kb�odL���Z��B�1�Ak1� +��xd`�S��G�fM�;*�\W��i=��
jep}ށ�zDRE5Q�Űt���9�ܙ�2�o�������h���}��[��tOy��Aޙ��z���wb�?�J��?�\գ�X���;+��uR���a��X�0T3��Y$E?V��`��[8��G�f��ZX�x�k��&g)̈́�Q���:}�(����ikhh��}/#�FT��/�npS2�F�ڞF���c'j�	�%Pn����ưfM�i������ZeWh����@����r����� �vЖɉa/�B#���h
rq��kf/R���M��D��f"��sEAW��k����/ٞ��{.�#$)Bv썞l�$kq�=(��*�b���"Tb�.w/~K�HmS"a(z�J��*��*��u=i5�3K�}��=B#���=���Hrb�m�@�6��s@^���\�&2��g���5Z֊�XR�HD�� �B`Y��.�')�&�n��:i�_��ާ����������Q~�/ܕ(��~�%d���Ɵ�1
5�ź�_r/[�R�K���SZ���V���%�\k�����T��'c�7n�u0�ҫl,��E�~��0�ݰ�Q�h��5t���z6�W-	�s⢜�>,б�>��d��sz$[Ƹ�V�47�.by���W�%f!��+�Y
@Їʠ�G1[{x����]��j�;�.@Z�t�+�4�ظM*;aͱ�I�����9�\ξ9�ӑa�M�6�V608J�"�JW'�%��+ë�yώ�А#]YI9��Y@bj\q���%e�$��E��<�{_�J���t�w�#�:��Ʃ��$M�a��lL��?r����d��L�I�t'CXxƘN���*@��"]���+|�?QV�\��of�-�\��G����ޏ$g��'q�a�8�>l�47�W?(h+��b1��TW�8!�eG(vM3�-8 z����bqYr��D2ʖ���3�jj��GN�<D�Ԧz�/�J@�!��<�ܵyX\�Eg�#pN�)�;�ݡ��,�m��9���홗���8	FRj�~!�ng�iV���������K�j�3��I�'��o�.����CY'��G
��e���9g�K�@��,���*��n�����OB9�|V�ƃ�o���W�j�r��}��$��.>̺)j25L>�����XPj�rc
���T��U���(+m|o�����/&������#Y��'U#�YW��"���֐�K2J�_�����t���=v8\!�)5��.�d�=�QS�/a��[~WL�r{�P?��KkV
b��Pk9��I�!vws���Sx[C�7�-[4�W�L��wI�nUq@�ғ$����a�⇮���
���7Y���D1�	��p���߅��+G����*])4���/�x�M��;��r��w�n�{���K�u^�{q ���p%��8�	�����P[�
gU��U�L���n��uY��//�>	m�$-w�8�]ħt��bZ.m�|�˕!3�u~�4ʽn��kЂe��]��!(9;~cv��$=m>!3���<�&+��S=�?�Y	L�j�	�T�Ђ	%DQ�4���&����z�`��<�k����%�R�V��+�ݎ�@��յ��Ω�����T�mϘ�/���Ҧ��*`�5R ��-
|�d�n�����c��f������`7Ӓâd�3=�E�ġ+��qf��	�~
#4�Y�*/a�aj�7,�- $k�s���|�?_�r��1�@�C�=%{l��{<x����L��*D�S�}_GW�. Avh�HG�ߢ���&M�JJq:,�d��\i�� :��9�)�V�k�1J#�Tф���#kV��pDg�P9.]�r��d�F�l��ޒ�D;������� "�K�(6q�_�lt���y��xت�~���`����б��kHV�	���#��jB�C�g��<��i���z�AzV�of��׶�<��Ș#��KJ��P���y<Z�؞��
y�<��S���Z��3�0i�^S�$��Ra�&�ݏ-Ɇs��j���f�皝$X#%Jj���G�/��!S���J*ڕt]�*�6�A�
����Hfa�=�k��v%��?�߽�"�b��T��L���>��4����.�y�fHt���-I����2b�:������-��E&�!m͐ݙ��g��v�
K�i��)��������v%��^��d�<@ϥ�`�0S8�6g��I�+��]t\ث����� �N����V�l�b�Ɔl�*\X�M����Yji�/�_ZA?����P���X\��M'����Wm���)�i�%�m~�H0ҩ��t�?���&�H?kC
��Ӗ ����\̨��8z�8�^�ƂGM���n���C�l�2Ĉ�,��+�w/,�Z��qnQ�a�cI���X�Sm{���
��y������/��<}��5Is
G�#9Ư���T�~,2M{V�x��B�x��v����I12Q��i�q�N�CM�k2����b����jV2���Q9��|)}fy����/d�}#rl�Dꯈ	B�pZ�}��i�?�S_���Fә�S��8S} �����Q�oަ���:j:�?�;�B8T�Z͔/���Q�x�ՀL��v�e@�%����s�V���x��А�n��G���}H�3�Z��o%���1j2MA��P	�����c��F�8y��T=����{唘��kU)��� ����QV��˗pU����	m��>�����G�#�.���T��J����+5�φ�����΂zH�O<�Q��S�0��.�	�H/zo�T��}��Q�.��}���PE��L6vm���?Q��3D4���i����1l�а��^����AOFM.3���2�`+��c*���G��[nq��v���J7���jW�����n�. �BRn���]��� 9��Ӫm��x�L<l�/!�ԤYb�2�2Q�'�;QiY����z��;�D8�ͼ�R
�>'��``.��ߐT�����jF�*���-d��J�5�%�1�o3/�?�m�a���=~��mG�5C@�%�9j�+¸�g��v�%Z���'�&�%:���"w�[욻	aO���>��ŤD
�^_�w 37��	z�M�5��QG���75�L(zT��o,��&LSL�`,Qh�1'�>(Wda��f�L��0�X
TO� t��"9��/q���R�ú�|%�v�ӓ�-���iG�s w����Jt�鲍φ��w~��f���}3����)i�v��h��\"劢ف����kw ] ����=���R���̯_D�����IP�R�~؞����_�� ��}�4��ޅsHSQGb�82?lp-����%�Q��d�P��:�^T�C��+��X�1ʒ���e!n	IT�+�[p���c}
��e�DJ�y��&�?@�M\t����7���&N�M�u�H��:�q��'~��5|��+�";.
N۟�;"}G���r��1�Ph���sH�1�[�A3M�;�����o���ܙ���Y%�cZ��U3߱2�s�w��s.Cߔc��.'	n�ȹ�_ǧ�%���W�ˑ� A� ��CѠ��՛�5��1n���i:�%eܿ~=�ȞO�ae���?kgɃ�m@��9��3G�YɍmvMX=Bޘ(�D�h5a	UC4���8�����p�7Z�r3���ͻ;��&ק�苿/f�}��G4��[��}��o�к�-0�J'(k�)MBO5-���̈	XE-�u,�������
/eO(�,�ik�qL �˹��Ju�O�K��?����o$��i�-�D�k�~�=�q\�}C����B���Y��A^�� M@�|�8���Lxk��Ҳ���Q������U�&Co4�|˭0|����@��*�5@�x�Bv��GD�0&�`"�bǸ��R����\������2D�!�>�G8F,����^A� �\�ǜn_(��,EM��v�g��.P�/�5����#�Lt*:^|���G$���5_��e� ʇ�JK��ԛQ)��AT *��m_��m�ċ�2��Ts2)wFMQ���+������*���D�B��he�X=E�g���%8k�@Zg3�1�g����nK0�w�]� ��҄��"Y��<���2������Zj��gּ޵��1t,9mܜ�K�2i�������"����*��u6I�LY*h�A��j6۞4A�gq$�D]v	R��Gر��0�8z��]բd��++�f��T�ʤf�7Z��abq����k5�nѶ�/�iD]S�ަ�~�{	�r?s�4s��E����.o]K��b`��f>5%����S~� �����y���z-�$���*��{��h����H���>�琛�1�"��p����C5�4_KE��$�p��#��^sB�V��]x6ۚOXi���v%r��JZ`'�9�J�	�6I��k�aC���S>��3`��8u��.�� �!E�q.y��_	�MD�$N`%� �R�
��ПA �8�ȓGS�Z��y���C��\&"`wCT<�2�;7pr�������kTA3ېUC��F`�C;E�����A5:�{7�z� D��$�&��u���gz��O��(HIY����'����<6��_�r\��^��?f�f�'��ŧ���}���u/��;P`^���+Ʋ��d�2	lzX��kX=%�����J�<��u�~+6J��.����.��V,]��b��T#�u��o�Z���c����-}�͎@�D:sv+���*;J��x�5 �P3�UJ��2�����@�o�R��@�H�b�B����Rd����h��)��,V|/@t���^ng��m�b�0C�dA�ߪ6��:oͬ
��ukO8j��FE,��,!�e��u�(_�轇��`��X9���* ����˝"JE6�sq7;|�|�CN�x("N�� ?,;�?�D+OHҞ��O�b����"x.W�T8[4��(J�~͎��?4x��~��s����94۶?����&�R���|����k΢�cY�� @"PHz�q�J�30���↗��A{8p���6��C�k ���lr8��j��r�s�&.�egȑJ ��*m?|�� ��i���K��u�;�lz�FnC=e����:g^c���wZ��J ���^� ^�n�A	pӞW6e�\�2�˻U�O$_�Dmߑ�w5-����B�4�5!8�]ӦPG�K��͆+ϔ�S��� >	r��;&�#c9A�N/���T�U��&�n,�a�D��3%�T�!u�Ɇ�L�["
2Iۺ��6��g�L�Q����M�DqP3������JU1���-)���O��1�J�8�Y��!������"���ڨ׽?C=ia@g���& ��1���i���Xx�C%m�c?����8��T�
��O�ɋL�I�nE��T�?��ɴ��--V��
=L�@r�e5mq������C�)z�0k!��g��V���z��ʴ2�T�-��p5%!On�Ht�	}y�zĖ�=u����rSp6��p��3A���7cw�Ud0��s:D@'�n�%�M�*ՈIV��M���浝fXK��MЋm����I��X[��GrI���Y�J��+j� ��{Pq���m_�e���K����5銋r(A�.y��v_S����7��J�D��T�b�0�]��g-������qDow�u;����Z$-2��i�d�1�e48���{)R!�o����H|���0Ԃ���^��n�+}j ���p���6�Q��4�/�gPn�rV�X�3��,H<i;����(�;��Grb%�$p`?8j�����	=Ǆ�+�����TQ�.�5��'d�i��8�_��w��������>�W+��QVh
�D'�,���9C�J�c�k<ov����,�v�,q���D�e��k�ܞ��z��ܑ�L���$���.�"�7`W}�|q����(�ص�!i1uU�*�D'�jɁ�X���l�:�/!�#�>���	]N���p�^�����*KH�|�J�#~q�{�N��Zv��R�g$z������g����?��Mj�Aq��<u3��	����vV��I�W��/�ZrĤ\6��7mè�ٹ����"c����W^��]�s֍�ٻf(_eT���I��ʞ�Dt
�c�yU@Q&U͕nz��&wg��_Gג������@O{&����`�K����.��N����*���Vn =1- ��Cx'�F��{�y�� ��~�qg����C��3ϿG�A|�믧'zǈ��,�����-7J��Ύ婨]�$��h��V�{�zܙ45���
ie1p��K��j�n�़\.�˪��'=?x�d����6����u��C$��2���{(�f`fO�zqF	@�KN�\^F+`�i��ܢ6�A�����K�_�^��m��
�� C�ެ�%38���wSu=��a��zm�X�m�K<����FJ�����`}s2��o��=@���>��9W]G��tĠ�%^DKͩ��4�Ӓ�9�3C��������Z��u��,۠�8=�o�q��B���TP�`����KaV�hU�h�M3��v8QKgr9�t�7h{F��ș�H}|�*�)��%Q�,��8fW��n�/P�|����~���ϳ?��$�q���hWN��#�8�A�n�9�+ML���Y�Q������Sߞi�� #���rڀ� ���� i���1h�&�����޶�"G�,A׆�Y�P\ٯhՉ9�T:,�~O�Ǵ���Sl8u!c�� r�SR!���I�E�d4�w&���/�������'N	��[)
�:�.�P�ׇľ����u]�ԅM�ek��EpHAGO\IXo@����eQ���z�w�/�=�p���W��eqMe��҅{Jֆ�͟�a��$��Ͱ f��w�/��,��Gg�]�{|�R�7F�MU��S�:P�01��2�ZM��*?â�]��y���˦B4�Z��>���9���I���aV���V'�~i���[uD�-$�ߘ��@)҈��
X\r/@I@����0�D��y���Ƙ=�a¡�L=`�`��J��yN����u�OH5��S6R�v�qHn�y+	`>�U)SK�p�FL�������!�!�1��0;Ȫq�e��C}�����W$���}��UMp���m��X4x�"�B�B�Q����Ybud�֕d��o���L�ܸ��3|�*�P*WR�����%O�l���z�8�u����!��T��9{]��]��-�����=��H�%C`��tV:�-��:���N�0jɺC���l��E�I|�UJ-��iqs����P��7���%�ueH��DH^Nx������p4���y�b�0[f���y����^ ��Ex�o��|�ylC%�b�sP�*��?����D� �H��o�Ѡmhz�=҃	�`�P�����\j�E���G*���F��6Fh�DL�IdZdz�%��Gf���.�:��ʶ�[Z���3�S���YP^>!_���Gײ&s�]^�� �����-�q9I;����!x����(G���φ��m0��K�:��e����4g���*jn�l1#��M2#:��e`yH�-�/r�T���҄#�m��㇒�.�ʽ.��x�u��V��c}�_�?;�?�Hf8X���~�>v�+�6����t"�lCa����QsT�{F$�E	��X]O�����X�#cc�ϱW����R��5�͜��{�F�[,S"F:��*�5 �@fw{!�0O��|shF�^[!����|�o�Pv� 	x
��`_~-����V��]D��b�4�t�)��t���C�fq�m�x��^���j�Q�w��U'��h���-�󝏩Pf���f'�5DN��H�8��U1�e��ؒ���F�z`a���:�� Lm-%����߇�S�D@Pڀ74���<�ү�Mpr�JR���҈�X��?�0u��Mv�ӄPK���md���XW�O�.���b��f�!��2��`�.C)�_��r@�ѳl�p)�H��WE����{�%�Ft�r@.
K�s.к,'ϳGz���T�3�?�6E/����ևÊ!����~s�[�<ҕQ��k� %ƛZ������+Tr?+�I�et�*�x��W}�p"\w+?��͐��ݺHaɏ/vp��8�'���a�����ɹ��IV�f[>��:���<K����YC�GĿ�(���j���n01��Ɇ|�X+�rL�I%���@��㮒 �eL�����"�A@��VYe����G�N��K�$�Aſ�9��:g�(e��V�=]�.�ߋ���W�.|*[� �Rjeг�Nט��mf�C���:P�!y��v�����[����L�~y�*W?sYhb���6A"�0"R�Ԟ���yh���&���ry�� =T�'�& ���d3~��[�^s=.���T��v�4E�u�	T��,��LD�'XsRT�y�>��6}��#�XB"(���g��Ro���$C̞
'����$J��l�fs(F���ߦ�Z�S��K��{��I�7�q��d��y</�dc�E��|x�h)��%@J���6v��z�%�ɧ�^���/��c��2���a1� ��J�������O�E��� (K�%��e��|��3�8.��Y��w�Eh�(N{b"�L����D�����hyB&�|�K���i��r(�BwF.�����-��{�Y�*�+�n�˶>��頼�8js�h ȩ�^�:EW��]��Q��@of��fp���l^a_S �>W?T&��r�UO3{�G,h�N��I��6kɨ.��?���]
q�:��w>�Qq���"Ho�^�P�S��Ǎ��ﭩ�F簵�,j��������Ɵ���]j�?�P����W{H�p(,FY���Ù�H~/�6F^~���ӕ��S��
X���∭b�C��� =}�ã*H�N�O���\���PL��n4��l�N��B't��7 �i4�iS��>c���v\�5�$4S2a��V�Upt�N���cw�j{bķ�! �Jnz�Ɖ����ʣ�s��c�]2�&P��7�)?�Z�RFܯ���1�%0\h�� �@���Q'��m��Ա��m��� IN���)��7 �Ś�1�r흟��~�O��	6D�����(C۶y#Ek�䘡Fz�'�::�
�ýp��t��t{��!���}����c����� �+�w����	�)'ޭ�B�ͰBM���1�}��27�E��V��ȗ,(��l�JQ�8t<������h�������,�Z�kY  ��RFfx�|Dq�=}l9υ�3Y���Y,?R�ܯӑ-2�� 0}-!J�����Rʤ�?�͋�1�y�|�Yr>�,&�1�!d.e(v�����q-��W�M����e0��+�Q����ڂE�AR�}�U����9�'7~'��^�����؉�U��e;�x�U�e �u��D07��Lj� �.�vn8�>��_I}��o�tM�EM��<�*w���~�1�6��%.�I0M%z�!(7f�^�?�^�y��I8{[J�*IU���;E?<��"㞜�N��"E��u��ޱ�w� �Y�C��O�b�;W�>��8s2��#g�o�Z��4]�4xv��{���#H���n�m˫4.4*6�j'��V}FٛF�Gm=�j��t�yNד�	B�¼�sA5��N�a�ـ�N��{��3����֠���D+bVy�Qٶ�f*�j�&�U��̍�V}�(ύ=��_� �0ꦶ7��_uX�~�+ӧ�l��-:.�GPgZy��SǿZ1]��r�?��N@�.���p������|)��<����Nٽ-�۵�,��\�k��5��:�z刚 j�r�����`X�;;��D�c�G�p�
#7�[�K�;��:L���.�Q�n������6��'j�"y|vپ���\I���݉��Q�0V§�W�1�R��^�1?��4�Ths]"�i�q#tk�°F�-X��0��ն*42�\�Os��J��%��� k�� Ci�d�IļG o�_/��	
��s��������ׄ�U����2�!+���su=����D�
&|���X�K�2�n6���~���>Ͽ8��ٸu ����c�%ä� 4p�֦jno�h�YJB�[��nG=ܸ
�O���:tқ���g,�R/N�CW,�
A�X>k_(p��?�)�O �YJA9̱�UtT@� �r�\�����sz]�+|CE�b�L=}�-�G�� i�Y���q�=P,�X t����y�S*hXU�	X/��"�C�{��m܍��`�,�Y��L�q|��3��K �yؼm�G�vܭo
$q4�;� �aT�)�T)�sI���3�2L���'Q���;��G��!���x�����J�6�',ų��R؉��MhmG�UWt-�JWJ�1�K$o���Xԡ�76 f�֜"�zJ��}�?��M�dڔ�3%8��n|a��6H$�7����5y*0��M@��![�}i��F��l������dĠA]��75�P?wY$�&3�FG���C�[k��Dw�Joʩ.P�;�x> ��g{�c�,���0����,`�Xu���W��sM馮����x����6���ϊ�wο�M�H!�}	����~���C�˞&����}u���m��B�2��ݡ1� DD;����9��?��W�`>.�2�H��%.�^��˗�#}͆,�s.}��Lu`�&���PLm�_bO�+�)\f�%)����<z��"��ף��.����@���E9hq�I��D�g�l�p�pU�Jl�2���k�(5�>�ཆ�m�2g�e����m����2�KD�����d�U����	�V����T��������C �!H$7F�x��1B����x�{�?E����[X]2�Í������z��ڊ�d̰�!���c�	���g�����f^�"�M:�tO60q&S`�zRz �D� R)�9��5�XP +0.�X�[��ڃn�T�'a�9e���A��_P4����dH���`���|�������Q�����@�3
�k�a1S��-��� K����(�A"�8A�S�NSjO7( ��,)�p�?֟��5�����7�Jb�e���Tױ6�pV��r�;'.�5/*��(>D8�iA�.FI�~���������
m�F�"״��~�0�+5�i��a7��Z[�#�%m�iW�0����\@=R�[x9_7��ݸY����A�]s��
�nw�X]!�����61�zý�͡pj�Y��4%��N$���B^����,�#��9�l"E����l!�x��=�\�@�*rֈDZ�+X���6Z�������N2@��~8,Bah2�9���Z1`�e=�x�+q��F�/k���+���2=8��0B���Ɛ�: P*�T���%,��ܚ��&����3b8O�+��Q�dP�q��E��2ȴ7���ҫȳ�s<[�>����M�];CF!�骚�PGљ����+z��x�FPX��	B����dOz��9�b��m+yl���K!�x�a�bl�Hא1lD	fM�x�[#GW'��|0��� �r����5�h�<�9���t_��*��	i��#��pL/|�貀�����3.�:s����R��[ʲ���L�)^s5���%ߥ�=�~�j�E�ߕ�b҇y<�H���w ���d`�$]B,j�9��ȓ�(֌v>����ycr)xo��=���wv�$�4\rw?Kы:d�$��Ay�fĆ������R\��Ui��w$�;�hk�+�LDӿ���*U��zS�x� DE[�T����I[�9��c���s2D��NLj-k�R����+b>w,H���nKJ�71w�>�/褶� b��� ��NQ�w�����[��h��nO�O#��nJ{
��1T�Q���z�)wv�=]�CC��@�'Y¸֝����>�j�[�%h�����`�����h��|����KG���?y�G�����t�Ni�N1�*��4,�;��kr�Ow)��v�E���Hr�%/ܖ`p��	U`����fI� ,� ��7��x�]ʠJ��w�Sn*�(L�+<ǘD
I�z��=�x'�N��|}4qd���՜���7g������{���!��&Bc�*&�W�`��,���&�7�E�00f���$awD�L0^���c<^�;t�V�r<�m��ܑI���
���:�m�Ku�LO��i��U�?��]�8�i�x�p������c��yA��34��`��j����ͫ�󁙹 ~���u4(�J��ja�d0m�����f=����K��U�4%����b�
��*=�[.z��b���D�a(h�$��r�j�Y,IC2�I����;�R�����o����8�]��ѐ��6�r^ΩOv�H�=b18�_B��buYsǳ6�{�v���Xۀ=��3?>�v�����&^�A�P�V`�!LQBE�D��%����a,�m��7�/Ia}Eؔ��gN'��t�|���8GX�{�����3$v7�v��M����g��E4�5P"ظD��L[��`XR��e��@�c]g��I��+b[ /�*���xL����
��4���)��\�W��L�TX��������@�x;!�Ʒ���fm�D��D�"����&\^����v!�-�E�ZJs0q�Ș�֐�٢emj�c`6�'��p|D�����jʵ_m��=e|j���	��R�X��Qes*k���s��gQ�s��҆+E��9Jn�4c��/�-R�� S�B��\�C`��UE�y�᛬c����m �a�����R��d��s�#�=��̸hn2:�!���A���<�n���k)�^MEHa�ǐgM����R����nW�
������4.i�4�F}�R��l������|�D��
Sѝ=����@��d&  ٳW2�=h�U����-Q��K��	���/I�g�$�3i�LZHa�a��C�>���Д!�ڐ��)-����v"J����n%0+��Rc�f^�f��U�G�{���hϐ��?;�,g�?�l�� �_v�'3�V��@f�b��褲~uC~Ȱ�Ω8�h%6_W�J��,o:؅K����`�����*��E�XJ����mZ��6'y��8�X:�f�4�Pn�n��<�w�qM]�����xSW�Q�����Jz3�x{?1����g� �����ڳ�sx�U�(eM)źw�h����:\ʤ%ie�~�s9 ���n��?zu�߇:7s�Zw��	Zuf��Ac�ȴXH��u�/���5 �r����mr�&�mQ��ݲ��4ˑh=?�ѱ�n�����
,���g?��lza^~$��#�zK1���x��9�D��<�	H9xyIg�m0	�h�ܙ3#XQ��7H+�e�_�.\�bL�������r^A��p��O�kk����a� u5&nʮ�_�k�d
��4�������J�!��b�k^���"O�E�Wtx����
���OGW�a�}����1?��-VՑ��+F�聧�T�j��0�=�Z���
����2a>o�Fx0��8�e�U0%��H$�:�hq����������
��]a�)������wG�.U��:X��ᾔjm��Z���<N@T�~rM���@���:&�j�d/��B߷i�����s�02��!͚����@N��(ɒ�]̌
i�sw�3���2�
��~Pom_0Ł�7D��`�[W�D�.A�Q�e;��6��Z�=�Wp������e���N)-�4��Q~��c�'hfS$�XJ"�;��l��(�%����$��k_��G3-����-��8���%X;]o��[o2�/��^ �{�Fph=���+4�$�.��Z?H�F��F&ȧ�^��sS�/�Ǌ_��JM��Pm�w�`$ֶ��H����_6{�%zd�v>3�EA�-bH�;��#H���`����yIoU�.����֧T�1GQ�"Ͻ4�� f��I;=��fT(�g���3��(=�R�F�q�\S���"8�f7���Kqi�`S�{9<��|w���c7{:NmZ%Ff�Bxl���յ?�C�k��x��C����r�S�;Ų���)��뙢+� ����do�oiشb��F��@y�v�6����urȧx|)�(����!���d��/�2��p�1�,�9���|򾇳�Ꚙ<jѮjg �����{��p�����?�	��ο	K�"�&f�f�����JѪ; ?0r�D8XK�;��%e\�FE�F�w����@��-ջPmA
H�Z ��-r\\���m.�xt���۔��?8�V}��`5$y���t�u�7t�Fe j>���nͭZ����F#�f�p���$��cQ��>;��Ũ�B犙¨o�:G�{mc ���2��Ҳ~{��72n�>>���n�y�'@Cc�(�!"��)��'��a����i��e�K�5��T��A/�d瞶jh΄��� �-+[(���q$�A��4g�֣ΐW�qk#3tͻ͚�ÆQ�`�t�P�^��L̸�м����?*:�[��On�k�+8Z���v��f����d�i����Wgx� �O�?�M��3ha(��T��||H�p�b5�ы�b���c�c���X<Ϋ%8����QA���B�d�yt� 3�5��/
�X�r�pY?�u��J1H�TP>3�.:�n9��M�BĒ�ޛk�+���Aj곘!��j�)L)�oA�qA2ߕcAIE���&��JBr6ԕv��5�JzN�,(�S�0jN�de��.ԙ7ݱ��i��ae{��E�]�c=���y��c'+MD:��^�턮&k@�&��Ӧ˅��H�Г���9X: ů]y��	J+����~ę���^4W��A�C5|�F��U��t�;\�o��	eأ@ε�0(ա�5�HX�޼Sßس��yu:r�����^�IS,R@��~��7�Yl�fx_].S����x�V)=���xF�T���A���G?�NJmj�F�o��Ar�${L��p|@+_*#:��gR7���� �s#�4���֞f�����n��+������R�HY
hhh!��]j��演�7�����im˹��'������"g�#X��ՓW��p�Cv�i����6C��cu��ң���/K.�?�$�b�p��� b	j�/���Ț 0i�R��y�r�_G�j;��b�r�:�����J_2Q��`��{� }7��<[��z�Ԛ�A��_a�ܭ�E}�w�-��\�����B�EP[��K\Y�[\�8!��0����b��K�g�/��[>xL�dl�R���?�#nNJ6n�uF�Me8�����~�ʉ�j�̨�W�e��kQp�n�c�f�:�0p���:f4y�HBt�S#W�w�`�oM����k��pN�&Ǉ�"���-���Er�j)lL�C*���&o��u�t�����~�#`���T�;Mh��u�,��E��/.�p���6J��X�x5A̠bw�O�];�����@��X�{�!�X��.gh+����X{��@r��?=�5�e��y}�-�V7��3��W�L���ܝ��=^fY`)5}�f7r��gI}@;�;^u��-`O�k[��@���gN&�&z��L����<3�Y����DѤӯE�S��w�J���7&���;y������9]"�tG��s���^�j1�_����׽( QW����{�6���r�ܞ}Q��+����`�� s�8#��6' �Y;0��s�S���,��c�8+�9�Ms����`��s����r��׹֫�{���.�E���=o[2}F��Q� ������	�zo�,�8��S�#������U��%�;chC=�9�{H���H�O`�w�1Uu�����'$���`c��{E�}�~nd��vD#~ð���]H���u<�ĩ�;'��_��dHΪ�?�f���b�bHh;�yfe�{c߂�I�=��,����Q)k��3�gD�0��q�G3e�|���s�K��K�:Ӆ�>��z��0��<��w�X"��*�rn�Z�&��EP4�m$|?��~��TH�\*���D+n+�>@���lc/��&���&4\@mq>8���i!t���V�hϚg��#�Q��&78��渕��|��ͣY�:�d���_���L�=M�1T�w������U@����ģ�̅
���,�6�_��9&˰�b/�{���ʥ�@�0�EONş`�᮱l����� ��s�L����wM~��j(�?�ˮ<
:ݣ���zO���a�g*p��G�۱=u�H	���&.`O^O=%pĎ�
�(���Zi4��>D����m��3�°��OϲVi�Xt���H;-��>A�<%0F>�i���iۭ�t'A�/���ֈ�P)Ij�ݣ3���&�4��i��H�q�7P�}�	�[BVt�(��������G7���y�5�����yh�;#���rX�ԟ*����%�w@�Je������[�%���0ۓw3à����Z��|*��x�@Q�s�Q�fz�ٰn�iA 
,sb�]�}���x�1u���';׭�a`A����O�}� n�4ו2��D$T8�U/`޻��2s@���}�l�iHZ�!�F����%� �[��L):ؘ�wñ�Ȝz�n	��_!Ez�o��u��Hc�L{_0�]�A~�e��c�a=ĹL8�����VeuՁJ�p�(��x��B[�{1�p$U�s�����C�m���	�2�s�q�_�l/� D������ʗU@d���$�����H"�N�`����<U\^p��0�����N�<
�m#~�(��Ror�$���ywW��	,�2��%�/�'����)���ԑ��#Lc�����J5�Y�R�h����`*O�T�	��ټ�Z�dSN儳��j"���N�]L�z���T��{�j�2����F�WVK��It��&Ҧ��+�te�)����L��:������������X��`�Q{!������C�P��MX7f,�Lt�*h�}��b�/�u�)��4�!�����v&	{��ip5횩�0#{�(.x>��U��%^��@Z2��E�n���܌�A�
p$�B�<ŗ��N�M[����)d�����Z�
.k�Qt`�|������؞�#d��%���x���jh
�2�Ӣ�*��TkI,�A�-�	e!��6NB#Ō��az����1H�ԘN�"���QS>%fw�4�x
�O4�s��]o���oG�$"|��8}��yt���F��I��Z�t���76�-SZ���.L��ϑW�J�jc�W~� �cS����l��%�۷E�-����0T�����o�^���H)�0�F�F��ĳ��S�*l��� ��e�(�:��B��ø�m�ǭ(�?���I���+���Z�<⯺����Z��
,�B� ,����,�Y��{=�v'���s/"�}�j}Rc*J�͹2J�Q��_�D���ƌ�!� �?x�&H��}R��:j�٬�#d�_/��h��*=9�ѥԛ@�р�n�"|A������&�ݿ�u�)��L�� ��D��{����!dҔn5R��\u�5���w�k�}�<*�	V���?=~��d$�w�	��#��q�;"�2�'VP�P��>��@�^p�����usu�E)���'p%r�b BJKq������=�{*S��Kꕿ��16�P}s�=-O�J�z���yg1�S�4���
��d�Q� h)+6^�ģT&~]ҷ\Ȯ.e�9��Ũ&��P^�����%k�ZV�q`폞�&��H���O�+�l����F�eR*�ݫ�<@�h�����Cn�k�'�w��"�1P7n^C"A�9Z�O���'K�b,�q�cN,�sʀ�s<Z�A�����"�c��! �Aޡ-X�}o�%1K��tQ_�d��eu�yv@�F�IX�����eMB��n��
aƸSA!/��PVX1�Q_Nf���J7#6Ҿk
�W���2
{{l2�k>1�Sh��a�DȰ��l&6�*��Í�Q���%<�A_j|L��mj����_ry���UZ�0�������O֕D"o����tA�G����`����V�m��.�.�a��#_@<�
��e	�ŕ�6�gZ� ْ����4����R��4��y^�̧1��\S喇!��b���i+%xb�v��ID�=˾�\7��\`p��AE����w���U�%[T{	�d��&H���29��-�n}�d�h+��!�\���؁>�AQ5�!�_ucQV3�]`��B��u��P`-���,�5T�үCr.���^l�Pᜲ�bVeȁJ��(�	�u�[[dk� �r#t�[��X�P��װh�kx���D�[GV��� ��V2��55D0�C��h��q���K��E�&��Rbן}`n�v��+H)��i�g�d%��m5H)�53���.��*�Iጫ��|�gy�]pQrߓ�j3H�n}��g��TvR/�'&��ޜ3lr`���,����_F�C�D"���Z�fdp~���������g���i%_ĝM2�wL�s�k��nT��R�PH���x���!Qj��}4ߐ�b!�9Ð�X?��T���j(�YQ�u�r�Q~p�p�� ����Y��#d��v��k��]��p���Y���L��Y��
�z2f�&�!��I/
��F�5��ÿEj�t��b�4گ��|���u"����~�o��Ƹ�.�8rs�=�p�[8I�*�A|���h�A����w���m���mQh�}Zt��4��t�0��&ZEq�z��5�Q9yѧ��V����$G��t���t��٫��ji�<��9l�lc>"��6(��S����󂲌�޿����WE]�@��C�$gt�f�4*u���"�:���)9GM��NZ*Q5����ft[��	�Z=��}��]=�-�6O��Π���J�JxEA>-�;�?����~��Ԯ�\�(�y%x4	W�~��4�;�I����PZK����1:sl��b`������Ǐ!��j����R{�b���9�?
�z�:���/TK|�h1�A�'}��3��.��rsZ?�B ��i�:\�+:�%S�}�5���b\e��V�Lt��6���eއE4Ix{����8���t O
�@�͂���*x�jv����WR�.��Ĭ��x|{�[�Ϟ�Fl�xx������͉�`55�_Qs��Ա�FoԿ�V*��G���<)ߨ�B7�+��2��ٽ�!E������I^Re������ש�uJL�J��ӪA���`Yyxt�����Wv�i�Xׁ��T�~�G^����#��D��b��SC[�=q��5@��\��m1�*UU�e#(�8�m:�Q�@�/$�goO
���o�@2T\&K'�9o�ѨcfQP?�����s#�������B~{(ج�k%�g�`�cw[�C�
���hжcu�-�I�j3nO�[XEw��*���ǟ��
2�Q�z�z�SN�E��z��ӹ���;'��Z��@i���;��<��M(�D)��8)|)Dc �G����F9��x.'�H�p�N�pLq�����qv�f�*��߸������[Z�LT�s���T�i�a� zQ]JxS���9c^+3J*ljul�D�� 崂��f��2��+|�����H,O_��ۘ��֦�
Ay&�B�v��{��,��ZJ_4�V��C�wr־��?�TPZ��H��쎕cq�Q�a�˙��;����&�+��Z�
���	��U�:	� @��;��eR9_���7��z�E<qj��K΢崙ʥ�4����[@�/\�~�o�����Z���6�DP�i����"��EDd��׳��S�E�}�ʺ��+����*��c�,�'��ջ;y ��/��z�֏p{Ő5�E*S�=v|D�z�X�HK�hf3R/�TDE�/됲۪u�*z4�W5,�	�
�z����X�	�o��ڇ�n�8���6�C\h��Ɵ�B���(�8u��+�۳-� ��?� �<��~�P�ec(}��nN�l����p�m�,ʋ�;L�3�����P �k��ן��/��I�����������,�(����&��B>#bwF�:~J�+>Ζhc�l��.�9�O�Á`���~`�iy`��=H�S}��:�x.g7~\�fr�k��OZ��?�.��mL��w��0F�N�iE�@�b�,c<�%r@��Sn�~N��)�Ov(��'�Z�ʥ�s;�t��[=�/Xq��;X���dc��Y��|�����Ǵ���Xu���#�h*g�1U��S8%����ܹ�Ð�./;u1��(���s���]����͸>v�vx��b"��H�	���$��LRJC�Zt��V�M"z.��Y`g-�2�2��P��x=���# %4̦c]>�i ֍r+�B|1K�Y�uؖ��#�a��eRر�E*Sb��ɡ���7��q[]��H�)%xHY��{��F*�	���o�\"���:ګ�C�>T���;�tD*`�}1�p}䃿a�~�E8p�����g�>�.�kb��	�%G������%dZ.ƏN~��"�D�-�-�Ps���F�#�}�c��1|�`t��>���9��Q�a�љ��?�4��� ���՟�M�饌� ��j�����C�c�O��3v���/��(Eo�إ��j�e[X��y����l'<lGh��]�Vc�j'Ɍ�l#��ty��T\��OB9�5�R��~���G��AZ���R�9��5W��\[���M�z��3�"�'^1��>k�Uɀ�z�
n���h�2��%�5�W>1@[��\1HХ
�c�p&�rc�j���)�cp�#��Ұ�m/;�h��:Wµ��Ig��Ӵ���}�^��\����*CgPD4�-}�E{��TEf7o-�7��s���J)AKO q�pӒ���L�jvX���'{/6����C>$����\j۔� ���=�ŕą���ǺsM6F�&[j6}�G�nA P�6���.òF���2��r�������W��A����rS��87h�!Q,c�r�@��g��A!�î��Ps�(�v�x�nb��S����Z�r�ʒ�rx�	���b�Wy"���8I=3�H�D; �Ʌ*�y��4���A��ԣ�Е�}�h�����t_�x@?M�$7� R<�!k�=�=+@��o&B�)T)�3��2%1X_ *�
u�>�"yA���D�ʦ����}��8�Y��@����~���ؠ���D\����4�a���ʜ�c�e��3Y3���"'w~ ��`�P����vF0�a|c�eF�-�%��0 �k�ۏlBAN(w��X/T��n��Nh�y�AC���Q�f��6)�?[|�1��7݌�J��Y��;���Z�4�2�=�j����
�z�R�&������<n �~�-�!��O�>���k:�^:�n��x{
�6��H��<A���o?��b�8jKJ�O��|��nF��=��=���kvd�5�g���ҏ�v ^�Ў��Ar��n��Z��&���&���,!WkR�l��q�m1�@��g�&�E~"����<�˖����®�s�&.���?Q�]p6��4)�k�1>�ZlO���w<3I.���zv)��g�8��z)R�zi:��ͦ�m�*��#2T|s�Y�Hv<E���`|�^��9�Pg��Nz�ly8K����.��W+���y٪�$�Bq�؇j�숫�f�5C8I<��a�K���`,������k|S�2��u%(��1su�M>4~PG�p&�cK�����w��4?.f��#�U�zXH<�s���#�Oӓ1l��2�[B�Y��A�c$�I��~`����ӐaY����H���i�^X�YB>o=� �ٿ5Á�K	�lN�:���R�p�'�*���F%	�0�����{��|�MO����Bs��[�uƟo}���CH�up��L7�߾��>�PQ9XA�E��W-(�jo��[�w!��1�1��@�oV���I�;��L0��OW��T�C!־&º� �y㎍��-���4d��� ��ŋ�	!x��(��j�"��d���q�L6sc���ī����Y��(��?��'�����|�2+s��G���Diz'\"�m�W����������:r��1�Z�)�9����;'�Åue1Q)]I�"��@�A�imZ��j�u��g���bE��m�8LT����Ʒ@�r{��y0(��NCT�ap���*����������\����ֹ�I�����~r�K�o�}��5����K��>`o�q1��80�ޭ�Z�t�!C3��"m��Ɛj6`�IkE�������p�54*�Gt���yp��h����z��vE?�
l�$�sk�TU���4l�jV�G���oՓ�"@c��'�9��N	޾Ɍ���p�a��_�sXe���Hi�/���$
~��V��1Pn���ky	k������~ɩE������"P���!���wGī�$$X��@���Bo�W�-���D1���@TJTٖ2m���10���hr���B�T��P��&(��l%o��P6�;��X�<t�z-��;u�0�+����Ȯ�ro�*(��h��=R�R�y�ց<�*���#�	qW�sz֒���M�rl��#V5��r B���Eu�]�=���^
��qG���5�K���m�	��>a�H�H�i�V�l:��R���lJ:�k�7�LD�[ w@��񟬱6#��F�|)M�\M��Oo�Z^u>B���� �E�.BJ��*���K�Z'���}@�_�Z�7E��f��_�"���@	��>�$n�&�x:�ib5�˹]��c?�3��u�;G��r2�A�c���o�[-^�]�c+�E]{�g����jMo��e�hX
��兦p���[��h�����է��j��E6/P�ܹ9�(��,��6Y��	�><R�@��x�f��A����5��
�H�F�Br�b����«�P����ۻ�@i�� NH>��I�'�g�u�5Icat��~��k��D��������M�p*{	��ըvexB ݟ8��q�p���D�����!����x��qǦ�}�V�Z(�����:�w�;<0K-`!l闍��1�k?&м��y�,G�׈�P/����o�_�K,h�Wj�UlF ���PD�0���D��wa�-6cp���-Lh��Q,��H6vy������<!��uҐ]��GܢqO�#w#OV�{�.����$W��qr����������Oߗ9�)�h&���@���J�'g'��5g+ZW�׽� '��4���5�s��j(��tǥ`��)��x���0��+�3�4߹�)����MY��\�F*�A�QL��[(�Z�<L9=Sκ[��蛎m�F.BN�|c<����Re��H�;�8��^�X�)�v�<7�AX;z��3���s��3��h�b?߀�&;��b*���2��x9�����@֊���^d��wZhUџu*E����&�W�����CGҬRo��L
��Td'�0J�R~ɑ�t��a��3h��K�c��~�&}A6���T��6K~4O����@�0��E���yZ��<����[gxǑ��.��`\B�<;�x���w�hȪ����בs��ZY|���4�2�����s+]��#gl��k�N	�7�%iC�GGT����%��9�Ѯ��H<NO����U�~܆�ob�6����ef��E�a���G�~ݴ�c�����U�9��=�Y�ڽ�;tE�v��٬����H����ʗ<�7`�(I���pp��6B�_�Tj~�f����Q��`Uљ�c�0W�0~H�2R/48S�����'[#'a��y��]�?g��'�:�Pk8��XZS%�4��p������W��H���f�z���mBEjbRlȮ�(E��D�;��}�a.8��o��j��/@)�#����$�b���1��������ԯOU�?��ݸO���D��<a�Ϣ�~�G6�G�rk��=��gL!���,ǽ�)K��~R]���Rnݴ:)
"Q%��[���&�*ʛ�Yu�P�:�9��k�����Mn>�e.Z��˨��uYsJa|{��/I\b4�k
s:4R���+s�G�}�LM݄�՟�g��<E
�5ż�Cq�nbu��̽�>��y{F;�Y;�pA�Fe��)Ư����W՜��@��\:e`�UwC�!�[��3������3�y	���ǅx)r��Zⱌ�/�X�BsC=���9�YxY"Oi���M��,tV�ѨO��6�L��q��(����U�
���ؿ�nR��(��*2am'�ya��#Ɲ��xɝ�ee>�^l�e�}��()����'���اg��{���|
S Vy7%A���nLS�����us�Hٻ�*�j�@p�]i���n�	v��|��xf�0^4��+6O$HŪ�#�w%>��]���AC�\�e���GJ4G6A���lq�y��(��]�Jlb�[���Pgg�:׻lk����u<k��	G.� ��<Ζ����#���OT�g 
��@���+�p���8��n��l��9=�a2c}f6ia:X�>*2�Ȯ�{�ɽ�{��~4�7 2�t��Y���i����� �F�f�Z��� �H��c�����#����/]O,��֢1Y�����.w�!���e�5vڪ0a,�!�����$������	�9F0��!1�38{L�3f�%}��̀�7PwK��9cy�����*�-J,xL�pU�Զ11Rfc����ܩ%�T; y����-�@郾ay���\��2�R�C�!�1a.�q�&p*�e?�K#r��XD�*�-˹ܼ�~@o����^���B���u6?"0��TE�is�.$�'�%��VF����r��@���@��O/����P�ý�4>!�j$;��O�	��>���x/�VTz"�I=��q�:'���p<�0%����L�FYRe�2Aˣ,s�<�.��iy�a�Y�'�:#�2��Ħ�!�c}^B��?��ס?����_�;	h����ӮJ䣢�4����a��+�j>�݆�(����g�
�|��[?s�b��9�J�#;��ۙP%�"y��&�@��;��Jp�|Y6���e�i9�ɾY(���}|0{��[ן�[W���W�5�fa���gGa�2����?pC�7+1}��HS�(�O�>�}yiwT05#��p�!�}���BZ��Ɓ<���O�i�!��TX�4h2Pj]:�=|�kr�O�+�����7�;��X�$]��اI/��H�n���G3��>)72���akz%G��T��I�:N��dA=s��˪`�U:{H�]��B�E��߫ogB�m��ku�K�1I��	�mR�V�[���R�������(���VG⮥'�/��L}�:�y�B�` �;8)���qΉ�)��K�XDpN�p�0�p�'s�B+]6���R��8��K��l�F~LYo��C�ۛ��Jn1k�A���.�t�� �6>-�b����Ðm������[�v�m�������q:��	I+:��C��D7e��2��˻��\�JJnM��������ْ0�)Y���@ʆ����,Ȓ���"o�m�ܰ>��#�Jr, ��aq�y��j���?�,�z��0��6�6�l��h��빮�\�YU|	�Vǰ���X�C�RF��|U�47*�tۉ/YȂ��YDL���&RRg����V�PǇ3}���
�k��Ua!Xj�}�:#�? 7̵�����{��"��2���ɥ���ѷ�/T�W`{�T� Gڂ���z�/��`�zWI�5WG���~�Ez�I&f� آ\���sA Z��A��<b�*�~�xE�H�=�5Дpdn�i�d��<��?>p�~�H}g�:�\���tq�0qj��"i�h�p��
-4W:�1�"�;Q������Z��5
4�SaJ*�&Z&A��z�Gԅ.�^uÑ�~������k��'Zh�Ĩ#ى.���5E��'����#r ���d���Ρ����4ku��՜�WT�R�&S0����y	 ��rx����$��K����r���r�m>�
k���ʩ�)��Q�P�����.��Jz��12ՇaR�1O�x�J�b���H6*@��;$;�ԉu����%��U�`�+Tz<!�+����?�+���{�C̈́����Z<���vg��+�)��i�<!4��{$�Č s�
&���O��t|__�Z
"9s����|K��L8�RKC)v@�׃�@�>���\Fު�@Y��� s2��D���O�6~��M�8�l��<�Ly����-d��ڈD�琚�8F%�	�r�Cq���/ �jGX�9��d&�Ť����D��n~qä��6��;ך�0^rj�7�`��޶����-����ĭ)�I��fS.�: ��жG5�+���0ik^�x5�޿x�d7��֐��nA��ϟ�(�|�A������lp+{T��v'٩L��俞�ٹ����N�O��<)};(3k�F$�W���P���**6P$:������˘����:!QmlQ��H�g�5p��
���;�!0���_�TMH��4ђ�ѳ�+E��T����g�C�oQ����g��tV����7 ]�P�x*c��P3�w�χ�ӂ��6��GZ_=XF�b�̖����$x�:c7�O퍴���<j���[\�����MH�KЗ�z�2�sp�S�B{�KL�v���4�=��Q׳hXQ����;s =E���:X���)2�5���K�S������)�w����/Za�r�9�w9�"S����+�)��F}eG�r������(g
W�P�g��Y�k�?A|Q&��+=�c_v�^��Uc�m�&}1�u��d��ֺk������Hջ\�9?#K^�lx��3�r��$:��5�p�<M��/$g�i�H_�%���)l��2;zX-q���I(�|[�C{�dK�$��+��{�2�
.6�LS�ۈ'=�N��;����kK�����n*mt��1�e�bs٩��p��c���w� p����J�;8)�˗��8ڿ�C��X+D���Gtg�&2���'�B�<�A���ƨ+%��i\O3�?�]^ˌ����pg�]5;㤲�G	!Z��@�`Q׫�t�6�~�����~�̙�vq�Ir���^���j�ȕ��'��-�	��No°
��=o]�2jF�/2 �o��gs���;Pw�Y����kr.�+HQ����p_y[�<�$���q�n�(��r� p����C���M�o~X��C��	�ʔP�������|J�����L����Y�ȱ���6���IW��ն9��|�J:��Չr4Ѿ���B��έ�:�&^�V1j�8�S"c(ak����K��ȆD9�+�~l"�f"����L���#B����]计')��� �@N� [=fC�\]��p�*y�/|wE	hM �3��OK�r�p�����+ڜ	A�ϡ�4Y��g�Y��B�j/���n��\�����t����U^Pi��#đ)}�J.wȱ�X0�`�	3_�S)�QK9܈N�F�S��R�Тw��7�	�����i=u���k��8��N��5��J���Ab�����y�U��"�*>�P�|W���i������N�a~�,���J8:��K��3`��"U��Uę	cU6�M���g��ի-9�E��=W�&;O�K�,�!�}�U~zX�G�B�D����kơ1w��0=,r��P��c��b��DE;8�>)�dc�Z�u,�����ޘp�Π�̛�Q�Q�K�i0�mʏ����(���pȘ�f��=�!����|�X_��@1��/bR�,�uTVM�-�8 W@�U����ҍpK����������%91�~�w��3)�P~=���;�k�_�I����hUX�4���o&��������V�m����!�)���`Ƒa:Ś�����=z����,�wIĩ78�?#l�!���K�3{�n��-m��ύ�f���b8���k.j�LA�[
gr鋫�_�d�G� ���b�]����қG���D���ZA�<�q�b>1l.=�6xo��x���61�ȣ-_-�e����'�?��A��1�<S�1�����e��.j҈�m������r��(W��"@g�#�z�H3!�&#Żʟ\���K ^ ��P�An�j��`��\ts�z%,7dC���e��C�\B���Kg�N�}}[���8���"}Ӆtн�iQz� 35�C�<�Oԉ�}���i�1���M�ڙ(�1��?|�Jy����UU\ ����n���V��;sy�����({{����ɰM�
C�J�ZF�ϊ���k����%��'
Πbf|2�p�[�3�0��v8I$����SV+��r~ч]���yg΂*'�*H����N��z�=����'=�(PJi�Q�i	 "+4�;��?q�/+7*6U�n����L�$K�*-�Tyb�Ƿi����>�{���S�f���~CcB���]���[��A�G&'�er��<'C�5��כv�IW%�n��/P	ȔL*��J{�(S��q�J�$� :f�)��Y�z�$�1�Z٢�M뜫��<f���4�����p���h��삐Vp~G�M#�<z�JYA�
~�4��r:9��c�[��	ԽMㆽy�6���>I�Տ�D8=��ĵ���&��7�{˓�
�����9s�t���fC	�
�/+Z)[�r�a5��_�v.T֯]b@�F�ۭ%�h�QV���)��_óYE��c�=�H�a
էx��slI�W^#�H������r�������"?��2L�F�ޭJ��M:���md�Z���5֒�QT!�+�b`$��i��?^q�p�{�jY�	N�?(f�D�>���/̠��ta��Iu�uҳ�� ���[�=�*�z����LH�b�QN'��GI��E�w&�+֜r���#Z�Eդ�����}�ѡ�kz�l	��$cW+w�f��u=��/
?�L��(��3�V����2�������k�
ej0��XQzŝfT,Oġ6�B��������:�RBJ��)�����<bM�IHކH-(;�v� �ӶZn��Э~/
�w��o�e~]x$X@�;X����ll�t!��?{TWBJb��#C��>/��#�oB혇��$����;��A���4T��4����Z�3��"��S��[G4��,��y՝��X�S4�n���,�p$���@Y�fNK�5l���6o�h�hdw(HH��*�X���L�m���O�_\xO��,5 �����=2~i��-F'�LP��kA�=H���ʖ�^K�Y����7<���9F�[c�&aާ�:H*Ξ�|ĝ����ZvN�������	�.&f���Ƕ-�Z��*�d���HAto�'�	�Y�vM&��EA�%dE���Nʦ�!
b�� tegk@���Ѭu�l�ף�W�o�\"<�d����A�������M��c��Ѱ����Dԃ}�Id�a���(o�+}�Gm�O�f���8���r���,b0k{v��\�{#���7v��G�@=�y��#N<&�����NnB�Xpoa��u���2��}�=��|1g�b�uL��"@���~[�����:0sC+�8�ga���VN�9+��φ�������8��:��"�G����q�v���o�8fg�u2�P�+��^�H�Y���O
2\�����W6<�Q'_��3u���GpQ�Z@�bS2L	GB�A�RR����щ�_����n��j���o���%��z/}R������`Z���E��^ڣ?�h�\)��>n�s �D�����(#��0M���?>A![R�ҏA3�n�)�3Hṟ�$�x_��@ѱ4ҹ40}�e��%�CI��i��q�I|3�J����/[�ib_]�@��?���n�_��M��4q�-C'����׎����r�'cFfK���E_
+�4T@�+s#M���Z4�k��r%�yh��I��Ӗ"�s#I��z�Gm]?��	B��j��<,�{��o��~�"��jw*�3��Q��=�K?wQ��S3���r�5�^�ѱ9�4��0#`�(���\f�o��P�q�Qi�*PG-�H��C��_��:��7&�e:�b�Ǻ޾~1��|{�ER�r"	�s���C��T�{R,g���	py������[:�v���֭
��C��V�D.UCC��ڿ��>ӑ�z8�  D�Ft*�1KZֳo:�v/Y\��u4����7�M����k:��^�Օd�(���i��,]�j� ����S2Y��%q��)}t�JSW��r��	��,Ț�,8�.�|�\Ť�`�&j|r@�T�t���=n�1d�"N��@���=z6��W�T5?�����z�d�b�bt� ��:>�n������}��Ov��0	�x��RAM#����q���b��#�z�U�ݺa��@���'��_��8�Yo�YQ��|=��S� �d=]�}0�T��.�p'>�8lծ�V�I�DX�1js<r�7�]Jb���Ɂ4���ƍ����������d&+��{��s��F=�h���sV�F��p�ڶ"�e3Nc����ni�x~�d���v!G{S�ㆠ��yP@��do��n=6�Au���g�i#�q`F���L��^\��t�{o� �Ǫ����9�������yf�iy�SBg�a����� �&��sM	2iY����nJ��V~5��m���©�oջ�G�"tRK����l�QͿ� ݎJ�����D8g!�Kphp'�� 1PF��R@���R�Uη�\�N�i'��uMHv�!h�@��{ �<S�Ne����Ҕ"+�ca޷"�Gh�N���ɏ	��@,�2B���emkL@^�@ѥ�@���\`��l4?F��C�3;ϥ��)=�z�?���]�1D��c)����+{����&PB���Ԑ�#���k�4g��zj��6֚[���|E?�Y���$�w�M���#��Y��|oIaBW��P�Ԑ��E~�sN�w&��FB��pN����vk� ��IQt��0�r�eO�G?8�}A!}�"�-.>����=��a��O��c�C��S/���������P{��ݴ�����Τ-)��C5h���3قZФ��HI��TU���YiBaF����@zz�Axs���@y:-H_d�����2Q\j�� b��u�L��2~A�
�Jȵ�Y���Ѱ�$u�c�; ��*�{<�#�R�e��鹁���Qe�U���`E�_r����rq�y~��`(>r�M������6������^�+_GQ-����"4An�$?���u�����a�sލ�:��z���3ӿ��N+�O6��5���/V��ˋ�B
7쭙�c�PU��%������9����2onF(H5���X"V(�2�wML)Y�@Nx��	|$W�M�&�����x;t$@�|6�8�9��%���a鎔�4�]�#Mx��'3�u�=W�eR3]�%�xV-u�i��)�%�ŭ}����5���{�%U6�:���4��~�d���������BM�M�kBX4/��o&��"!A
�=	�hNm��k�<����vrx��-v�'\��ࡦ~R���&�B�ԁo�-�R}f>�s�����n�y ��q
_��˃��K+a����/D4�˄f��.V�S�t�'Z��#X��^�i1�r��u�yI�� ƴ�r��X�f�@�=k����>�|>,�1������/	�௓�hހ�I����P|#�"�C=xb:,P����1�tM�稕>��\��>�6�ئ�����-��<�n$��xmm�½*�x ��}�6Ȳ32U�.����ey�Lw3��#W�,��|e�*p4�lTe��(<�[d�a��`����fB����� �M4�&��}}S���5���B��0��_�0�����>�	[Л�;������on�=��b�QNڌX���H���
�ƪ{F�C��n�.��f�1'r �����w+�bէ�m�:^�b�D��
�?(�z؁`�T�N����X�:ڲ�qЮ�;����ܷF
�Nh.	�o���}�	����$?�}��{�]Vdb-�F�O�Hl%驆!��`m���|��;P,6l�qQ2�g��lI`wօx�Z�T����z�ݮi�	Jɉ��*�}�۞G:�:{���|�ϴ�'�r����Y>�J�v��vCX� �8��M��'�����&ǰ���0ͣ�M��#��?�X����K�^���kp� ��-=kq4�!W��<��}��Գ)�'D��ꋒ �$Ԏ`�E'��@��%L�4*�X���\`a���R%�N��y��/��a��i۽`�U}�(�M�^>�">���4'~.JʜT�����=ԝ�m�ܩQ�	õJ����yN�F.��������k~��;��H��\Щ�q�w��i��J)(��MA�n���H�A��I���\5�ht`�����OmV_9*O �u���0��O���R�+x`hQw%��T��/]�<�����xB?g�������CwBS�цxn[V
�||�v3[冑�ȏ�n\b6,6x��*i<n�YѯF/�%/.^Z�~5��_�a5�5�"sK�����V *�h�9ڼv7�N9=6A�C�������R8�ٶ�@�hw X�+���ͩ�����ndjDC��hC��^A�UzG2��_
�z�i'N@<e�qS�����1�7T����{�ӦW���`$O���Ǟ������,Ɣ�ض&x�l3�ް�I�����%���G`�b�0�-����we^�<a �Z6x��qk�ț�!��b�X
�]Y5�a�F���'��<�ΠË�A�9�K���U)Rm���hɛO����)�:��Oe�S;��Y�J�ƒ�ωѪ�cjS�te`� �1~^�U����BDC8��9�ϕZ ��id��ʹ"��23veT�� �Og9U*Qwk��F@/L�@�/#qp>
���� ��q ��*zY8�sq�!h���q�caef��"����5|�QDL���$M�~�i���|����L�0�<���}�v�n(���I�I����ͼ��bWU���� �[4_�i���Ǯom�~OBT�Zm
 �v����ve�p`
QL������Tӌ�뿓h8������"@z �!Qnl��p0�>E�F��Ʋ��.��X]Gk��1c_ĿE�N�{�s�n�Sۖ�yU�|� 
n����:O@��V�H�<��e����Ʊ�G~�fZ.�.\vp�F�XWU���q˺Ѳ�R��͉�f�d��@�!qP����"�[Ԋ���i�f��+�'a��I�H��̨y�/�v&u���f��8�|=�8��P&�	J��8(k�a��QgB$�3S���q���f���n�����Y�9�?5�����k�)�(%���kU�ҟ�����7��IM]��-V���ة��j��a#|=Nt��q��w'Q˱��⠡FS�4��U:�z�b�SC��#`�v@Sϴ
c��-����o�i����_[�IH�!�M�M�#�4�zל�|6]Ȱh5d��kj �mo�>���`^��r�8s܁��C_���Sj��Q
��5�u9�l&����ag��%,|�Һ*�ka���B��z�{ǭ�Ҙ�h�	'5��k��K[;6�[��?4W�8�MFFD2K\���-��������Q,�Fc������~�>����)�޽����+m��ŀ=�Q��y�F(b)\�ФR6j�O�Gc�Ԁf���n�?7[��R*��.D�?²�o��\:�����z<4>W2�{��5?;ټ�7�AoΪi��3}��q6j�(�^�&@���V'qa6����"7٫9�tw�J���g��S���.�[�	��J���U<��ۆ��.��C�g�hݍ4<�(%�z6����՟��w
�!na����ޙ�V��.���K�C�yds�����ڡWm��;y�Z�C3��?�#�E��W��;p9�wƧ��r�\�}q1�c��~�ב	�	+ǅ��/���^�hߓ���N\@�����,/~Ek���4s~T�D��>��ɶ�����wMs�ҏ�����Ӎ~љX+�y���� ��i��2#yIC�]�����>���yR�	��Dx�Z��Ht0����k�$^�S;�nv�Yĭ�w����헃,�5e��Z�N�ʵ����}�t�*�³�@T�����������M�\��5� ֲB��h�7�b ���x�yU"(2h
�"ύ$<��Ԉ�B�sz`#��'I���TΫ��lɍ��о��
���=�"�'OȮ=b��fDR�ұ�Ե�y���27��
ܶ6�y��ڙ�k�D�/�ו�N���^0�㐀�����������k�&�h�	Z�/MB�	!T9��Y���U&"���m=�����a���D���%+;?���E��	^�=,
��%Y[���
90Q+@�,	[�[k=,ҭ)'�@N�=,{ڨ��t���	4ruF����=���!��i�9�.�(M��G*1�y]@l�eX+2��k��O#���
V��&��'���x�n��c�n��'��e|٦�:4(.��>��Si��� r1'_p�f���~K�V%܉)󤱼a�����$���!�2Br�	;w9v�&9��#I���{`�<f<�� Tѐ@r��X;�J& 30'"~�σ�
^�,�w���H��
���Nd��ݽ�n@b�J]?n��kչ�30t
��t�{A�+�e�x�=�c�ci�S��*��X��c�䎂�	q�;��
�5iL���8ߏ����5���섫-�)�ΛM���0��\7���[$�]6��zN7�7M��:�F=�EN.��	�V4��P�,	��ʽO��,s	s�7��"��$�ow��mwe��`5����^�ۻ�v[�jX�ł�E�j�B��W�1�T_�px�Ʉ�WY���=���9��/X����u|�|Y=��l/����M�͸��N��6����@��5�ȍ��By����[�y,?R��s�ݖ�/���M��S�˫9���a��B��.+��W/��yʾ��bx�t�y�J��y���f��,k�Ƴ���F�T��c6�$�$� XĂ�wN�����:u�8��������B3٦���/��O&㱤g�_�^�x�#c��+Y[vB>�?�5/ (���ή�s��z�|�&�i��O#�����>w�G�U���g��̖�Iۛ�f��Tgz(�W�+�3�Z��I�v�[�k5���q�29�Tu� ���y�j�֨�:34%��E�-3 �y��hPBm%�ᝨ�b�cj�}>�)N�WuΔ����s/n�Ib�kf'ݵ��79"�i��C�:��4��w����� ���@=C�x�VX��;C���o�I�ʧs�GSPO�pk8�W��m���6�����
l��<>��sG7�V��0���b�	v�K�h��̣9�Gh,bL����c�rxl��e
�EzF�E����.d�_\
��V8�V�L�D�.����k���v�*l�{��߿,�_$��Y�.���s#�&��	��X�+��l��Q1�\I��M@^E0��o�)U��=G��%����2$���/\�������gT�A�A˕t4��V��&׋6�I��@P~?�6�����m0@�-x��O�ey��lP'������W��e��;V�?M��;�\
j#�5��v�0�·����2~[ZM�����.�l����Sҙ�=sRP�8+���(�v�	���`�,���J'�)w�"��"9��j7�s��vg�'����p��3Z�/��"kVS��<Hv�΋�xHE)�K{��2&���&'�K����yw7����A�{�#�����֛H�T��fy1LJ�
a��~���,�fAS*��#x��v��T	κ$���NL�6�}ۧu����`J�	�fA@�ǀ��Oʡ�mwl��uկj0l�B��.DОZ{ظ�:�x��vJ�L˨t��C)O�g]�����Wz��/��,��D�Q�����,��Y���<7�\��?��+�$�.ms܋c�'!���(T-gS�L�?a����T�a�]]@�\=��@(ۃ�=�y��m#A����}D'K:��?5��@�9X��T��U����֕�Z�y(N��۰M��?i1i�a'���J&���ॲ$�[��y͂y�~�U҄]�w^^����V�o�O��0���6����Q��S�5�N{�[�����Ɉ����M)�N��F��?��0�� ߸X��2�G�)��E ѭ���^�R���������)�-��&-vP�O~��?�x�;ڣ����t�a5?%�½��/f�(Q�ͮ�#��Z�UØȠӡ>y�(�@�x���"u�.�(Zܘ��������!�E�A�Iq�E�Q �ME�-"�a��D�%�%���v�Z,���XK	������/;���i�}.�!��2k�b~����&�@c�F�7�`ƕyk��Q���:������u��&F]�%�� ������BrPM�x7u����RS:�\�I~�`O������`��&���T��+�5K��ѭ�g��B�^���r_���F�GΌ2;���VH���{R0v>G�Ad�g����i�0�f�>D����'2�ip�"�l��S�x��~�@ �A&���=�?d���?z�k�k�x�:�;�J��U��֝5y?���OK�|���HXhD(Ǝ�?��8���W��Wq?��K5�_t�q,q̑�����>2)A3���u��ڐ�N' 
0с�$�B�*!������^'-F-�t�ET��N�#=̘_�F�tvU��Me���!��gX_���suT�o���s1�L�<2B�~��SM�K"a3��6�.k�V�X>2޲u�/�p�)���5����%e u� ��m��j[1D��D���G�� �bf��,t��&���C�A1��
?�D�0���X��:���%ԓ�aB��֖�tY�`+Z"I�D�oQ���Y\ICH���T���j�8Ο���0]a#�?5�������;=4��r��"�
uM�r�Ja����i�=����q��N��<z�g8���.ޠ@�hY��S�.M���[t�2�u$�'!�n�ͣ)�?�H�nW�M�I�]���ʆ���&�S[@)������gPj!=��i�񆖳��0�y�Ȅ��zc�����q�G�%(dF+j;4�C��~�#N���MB�ji*]�6�R!l�]{��
�i��B�j.R	;ϿD�3�Ts�\pm�<�5nF���^��P��WuKpIs�~  ����f4`n�|7?�9�/�V�M������3���'��#���8��Ғ�ޅ	;G�A'3��C5U���	��]�Į&Y`~�A����n.��4.���v�I}E>W�&^+I�u70�!��`�6Y�>540�r��o��������S�g��̝M5�X�z�����f��2x��+� ��▅���Vŋ���Fx�Cs1�m���L�I�K�dF�ƥ��Q�n�,�%����,�S�8�Y�?'�7������ �5>�.��>����>��d�$ǭn8W�I Ip�Bg�D�Rٺ���j5�˓sSC>/���/G^��2ӽ��wɥ����匧;N!��QZz��z���Ȅ6S\���73��Z�9B֦�a��d�S�@�m���9��G����OO��ggxl�c�8|������w<�6��"�s׀|�&�L�{K]�^΋�8"�6WY�3±�5���p ������):�JG	���̉?��+���;�K���6O�,�F�� f��Q��O��m>ɯx/K
�7�'�`=F��Q�U�ך�y���9��]��7M�cRݭ�Hv��d�32����2`wYq ~]����DL��/�\���/dn?�&_mx֥�X�;�T��e���e޲��]"#ȓ��Z� �9������C1|c��h���Y��,i+��4�
�3��_R�����xR�c�l^7������g~t��\U�|��VM�	Z�,O)����h�f�Gӝ{���a��Y��wxe�*���-ZR8)g/Nv��Y�p0t�d�RR�#� ��m���1
(,�6͗��f�6��:���i�`��&h��Xa�	� �	���/Ω���,�!P�`�9�7Xj�x�|�'�!��҈H
��	�H���[�if4��c�>���w����i���|bL�@A��I�?���:e(�R{�}�eo�SXH�W�޲�̳w䌵�0���U�h��>��Ԫ�N@�~���^A��ѵ�Ł3Ǯ(���*���( ���6�Z�&�Wz\�6��Y�uZ���ĸ�Sa��1r�#�c|<����_���&�Q�_e�������J ���=�|�(�i��q��;���X~�7e��j��FA�IGɎ�ư^�q�E�o�	�������,rZ��f�$�!��.�!�+ڝ��òO��M]�|w�m�W`�6�R���g�˗Zw�+�rc�C)��ˑX]���Y��~�����6��웱9��$�'jۂs�VòfC�"�MD�)r���s���y��{�ƶ��xM�J$	2YT�Dǔu�7��B�
a�|gSN�Q�nU�+x�́N��PЦK�E鷫�Y��t��p}/j��[r��G����;S���0Dy��[�^T��>b���Eo��D�NM�gF�l��P�~Y���EHF}`�k�=�F����R��V��{��i�aΊA��:ۤӣ�L�>�cȻ���cо&F;m��'��`v΃*��Y�N�q�|��^��I�걡�V�AiԌ(��h�3���}>z�ɽ�g�#HJ!�� |�e���~�\��(���!�R��G/l7Q��N��~H.A�ᩬ�$]���Q�ӄt�����wOG�g]��|�nѺfJ=+~�U��&��Š~ @����=G|T���+V��x1��]�ၵ/���a��_�?B�[�!���5��m�% ���h���*9���S���G�.��B�Mb5�0["i��G=n�Ѽ�����;P�'D���c���l[G��U��W�\���X=��{�p�')����AE��3�����2iŪ���C�������эsf��\u�V���Vwhi nM\Q����$�25k~/؈�8z��7l�"K�^mY�-k�T�_:客a��ؼT�����^���՚����$���M�f�X�%"ҰW���O��e���n%�W��|hy�
�7F0�I���>��T*��v�G��hz��´�(w.�)[�:t�Л͋�hQ"A�ϥ�U��4����RKѰ�Ӳ>����s4�dŵ�/j&y���򲪓8�t��"���`[)�7��*,9��B��_�� ��˰�Y��i� �K�+laJ� �F֎��Fb��}^z�p�Wc,"�2пf*�w9t�&Y}��k�p��r�&G�T�=m���%���o0X9�߻��;W�ܷ���D��\�F�.ɟ�ذ(*���s(�k�7F.p��w��Q`�U2������Ɗ��v�������Y/>¨��r�'�Zс�%��R��tXw~3��>(m&��3����*����5p��c�m� ��W��VZ�׉<�͵�frle��<���pQhk��X�!~E�[�0fX�=ԋ< �� �"!`]Ѡ�|�/qXGU�]M�rpy�G���A��t�o�*�3)]1�9I�V�c7\'``u�S_?�M�ܔ,�B����^�fIw�t&��4@�23Q��P*ҨE����ȼޭ���y�x�!��v���6Ƙ7�u�"����~-�B%�E��yҤ�qR5��ŋR�x¤2ݽ3s�+W���"���0�4���<o�8\+ٽ'?v8�m/n|�./�� m� W*�oqC��s� ����Ԏb�҅�RC-49{`�PP�c���8�B�_$��}�s�;��Em
�͓�O��訪��}lD���%���4
�&�R�g��a#�Zc�LM�.���{��l����JH����р�uA60��L#[xҍ�L���	���=-�sA��N��L������ȵ�<��ܝC�fJ�9{��e0X��Uc(g�-�y�*C�Vq�gWɇ����w�D |k�y��gA�� J��6,�Ҳ�S�%��5~��B�I�"ôuaD��T]Kt�����%��eI��!Jb9EvbOͯG��WþY^�S �jZ�hǃN��w����)��(7����m肣�{�M����U�<eUK�-e�"q+F$ q�52�p���
&m��$AN�<��&�4q�E3�G#�Ul&nۇ�~��( Az|�o�����oF0�E����i��x���J�ȢW�8�<(�D��Ou��L.��
OR�`l*R�5�K9���M�\��\pʀ\��A��l�v%!��Y���4�f�Zc���>L6��=�і �+�y�-���$�����gS0f��%A4]I�d���v�Ɏ�����Qޑ"��4�lG��>- �$�`X1>�_�#�:�V:c�	�3&�o�U��߮��Z��M�(b���n�T�ռ E����%G!��W���R"?��_�r���v����A�mB�������
-/}9��)�5ƾ�3]6�9y��ǋ;^�$���g�1��t�|$H����@���B�MC�g�)w}��q�S >�km�@C�n�o�Ö>�.svV�`�n9���Gb�U(�WS��~!���i��)�\�8�(F�	k� �+�h-wz��y"/�+C����!�Ɲ�)w�HF����I�=�._nt���/0�����8O��z)��1Zv��(�Q>,�������1$�Ę��Z~b�ɗ�ѝ���9�DD
8<�`���� �a崝�)�y伲l�U���;Y���	 3mƧpu%/9k�P���U�.�)�1�O���GW��{_��|^��0X _�V�����8�P&�n�0�����?.�9n�����>1��P�mJ*ګ��h�_��4�=��A��竽�j�?0i�[2���b?˧7r&D�>���&Z�+�i�P��Y�K xz�N�� 3��S$BPoc�S��zhW����/����.!:?����}x�K�Blo�·$=��eU�I�-�DA�y�.�?�c�)Z,N_N"^)7EKX�-�uo~'�B��C�W�Q+s�$�J��-����d��N�g����e�#Qv�G�ԩ\��Ӎ=e����� ֘	���s���XN�"UQ�Id'~�����<�bUa�1��rH����p;�Ǐ�/�@<�M��˓g���a�y����s-U��`ֵ��/8@%��#�.�|�<�B����-et�;��涎L��3�Y~�Q��i�3	@}jV*��jBWL�N��^��S�o	x>) }"`�GK�Ԭ�C+����L�j�� ��.Wx� j*%���Г���b����äghح�	�<(�xO��oqTM��	O��e1M���ü��ۣ$��2�г���2Ζ�Α8��z��X!r�3�4��W_Vd�E��@��s�'n"�l���� �l�Jb�>F�����t��b�ɥ9=����%����*Y�B��m�8W3�
���^pK�i	�s�`���˭��,9HN�:Q��YqP�7s�oY7M�+7��{�~�¿�['�l%hA�@�z:�Xʗ�9��3t#����2�=Z&���v����Y����#�kK+�r$w�>�-��Ԅ�:ʷ�N�`A�ٚk� u�J�r�~W*���uBr�^`�(��9��y����po1����&~��t���V�D{��?����I::�N���<�F���Y�,x��_P�]U �^�6�	@��RH�rT89>�'��|��v�?.����yă�H�t���0���l�%E�,3�%�HAm���߳,���X�)U�-:�A���g��1�]T�ͺ�'��7�D�c�̷+�FX'$�2��#JiQ� ��(�t �	�P+]�f�m[N�0��Y�����$2���׬���_�}- ��[�j>U*� �(�¦�'U�z-�ǂ�alL�LA3�aea�����c���<���cB)BS��+��u̿�r�e�R��8�=����h�wۑ�<����|/�sDmԛ�ե���xEd��n�b*m��F�Vf�)=�ˢ����f�<�!���S�O|�䝔l1��ʒ��$v}Jr�N�L�+�FR��}��!"�Y��g���$)����P��Ē��M�&u�%c����a-RQ����(�@�!���S#�XS��b�9�с����Y���[�����Rh��>Kx�m1Z�Ia�"%~ʙ���2_^d�7�-E�W�!�u~�&��O���2(G��m�J��,V�}X� ]��=X�}"[C�Ek�i�����cj�ꢌ��b����4����M����YOc>��xd5@+�	�{M�>V5�ۏ���Cq��`�sle��N����u�ӑ�̜�gob��PV�|9�l�oP|��s�ަ����=$��B�㎙��ΰV�v�[ÿ{�Ν�h���F4n�gL�O��_ �q�s}�{v���s[x�eA��k;���#�~�YQ,5��~33�m��h��׈(�U
���b*�ewG�!� �9�������st�3�A_�w+0 |��.Q왌�����P1���~P2L� ��U]G�B�S.�6p<2J��>b�7L�����Ł��wj���j����j}�Q�e���#!�=�5Z�4��Iş�'��ͱٍ��tl�fo��r��z������Z�4�G�Ss�-&�e��N�)����w�q���`-9���܃i�G:��������ᗓ��JK(���/}��~���6	�8��<��z܋���K)�r�JywIr
5d�6��A:d�����6��W�����xy�y����R0{�Vt{�ed��)9�[�v{�Ѫ?Wl���� �,�9A7f��G�@����hVd�^��U.aZw��|�h�:+����`��<d��
0g��b��u���A���J�ϟeL�8TQօ�� �/��.�O.`�l� [�W�������
�U� ���,#{��V���t1����;d���w7��(P��Qv�6��ui����lr"� 6�l�f;�ix�a��x���ۗV���:�IU����_'A���v-f���ͱ�ixK� ������]]�j]�wV9��j��v�NCǎ��S/��gQ��3�"Hzb�s��E���{�I;^0����'8m�u3L�zw,��s�����rSr��FRm��*��Y<4�N7E�1��ïB?b�־M�C��7Ґ�7�����uòU����U��m�ҼDD�-��5i�2�$Sy��%mˡ����"W���yp��gcI$eWU�q��D���6�+h8��[ݷ|�·����WdA��;E�����bG �Y.�ZL=��:�|���R֠h���
:�~���,���7�7�4�WUCz���������i��"V�1���h ��2���MO�����ljQ�R@9� �.�lou�Z��WNPR���wD�cR;Pe��O�3h���1������@��-�צ~&4�u��CW�Y�g)S���*�r-�i���ű@ه��7X��=�ƙ�vq��<ĵ_�\��7 g	�:j*`1����Ǿ�W�d��d��R�]�Qh5Hڲ��u�$���'�D	��7ѧB��_�j ���m�>[���Ѝ�j]����j��;�����k6K������qO�V�Ԛ~�����>�J[5��z_��5<�	$N�`Ճ���H���d����Q�}jqk�� �^����/�c����������-&��0}R�E�=W��)���rn1v�u�B�>R0��GX����O�J�2b���2ʼyK�hj�kl{៨�v8m���/������ʧ���8�^���C������c�:�I7��!�~>�  �~�iҹ�̣�7�X�\8cr�I���&-_�����\�~vV��%c�K�QJw��*{��4����|���}n�T����?�"�3��_�$�L`�`Cj�}�#��'*&��>+2���:�I�U���3�y�7���$��q@� N�m���}�$[�,���^w��C{��z�H�>�2؊�(�O߰\�Rq	eg��� �/�2(�
����pw�"	��l*�l������y�E��I�	D]�V5���ߍ��/#��A<����9���v<�fBn�Z�0k��}���o��Ƙ��5���I����^f��A�����k�c-��+K��:�
W�687sn\���2��P�d����sv%�,93ݢ	`��臠��\���6�m^B�rH_����z�%Y�4l�A�ո0qn	"�_�,�ki
p�A���#n�s� {�e�=����7�*Ö́�|ζ�O�����r� 8��pk��y9<��5�t�呹���F:ӈ�^~�r�%�U�gW�m�T�G��oG�r�b/�����Ic���oW�f��W<K��N�L47���#�r���ڽ��F�5X#���
����R� o]h5'�ב�^-��x�1�=V�b��8.��8:�=n�[>��qCkk���D���@��^E4�H���gFx���i�^��JO� o�Ŕ��s!^k�1�@u\�S,`VC�H����h�05j�/�j��%k�$Վ	.<Su
�f�Ț�Gg������CKƳ�Ii�W�ȸ��v@�1xn�;7�V���uMN7d�y�&��riS���XI�q;�֟O-��T�J��{�#���0��l}}Z,<-O�]=����8/-+K{����ׯZ��N�M��b����/��f�!#��~_��'O�t��!≞A���V��\�A��),�H�?�]M��NnO���Y�꽉\k&K��H��yR������6Ĝ�e�Z�^u%P��QIC!X��wGK���VJ��M�7x;b�]	�Q��Vt�|M�@��8@�]{��	3�V���s?��<��>k�c��g'�I�\޼%�[��wp�Jە����<�C��iX��m�^.�>��Y�:;��L41���C3$ ��oO���h�_�Z��y�-��S	O��ir���K4�H�m�N���k�Ӹ��T��M'S JeS�ۛYG����vA�/N���T������Ʌ�G�����[�ᙰi�!l
��f�o\e���o�w8�@��TP�r��Z��������4���!1�藺O ���`D�\�o�� �_=6E�{ZSU:�n�nXE��F�2�� i¥a���.C��K�w��aY����B����Mf�OF��ʁ�jy̆p�:���J�z��ҙ��c�RI���^.p����-�Z��&b�;x*�/�i�r��G�+��;=��:_B�gw
ue���ʢެ��\�J�<,�_���ʝ<�M�"�z����7DA,$�OJy�mΈ�B��PM�����)��G�-vc �����UzƗ�= �0���w��cT1�eYk���{���u?1�r���:�%��_A���0���(qR���F)#Po0�f��Ovf��n�XtF*a�4D3E��e
uMl&���a���e���tK8gY�b�9�)S��Y���s����g��R�*��l���ta5�vP���pĝg"L�>����ڣ}���wjGT�G��_4��f�����"�`�6U��{|���	%4��T�x�_��z6�[�2r�#�(c�,�Z�_x�b����C� j���v��kxH��qJ��b�SQOKx���έ(z�)�/{5DK|nF�c�.���n��d� R����[��б
z|^ *�Ț��U}��!���GwefࣀX&\IM�W����H����U]-e��iS^H,��p ��z�:�wk�I1�{(�V@�����gG�Z�i���K
�q����>�E�l�S����+���7�bA��i�� �Љ*C����|h<+O6�J�ʬ:W7�䧗���x��^�����F��J/�]b���+ud�p��������9�d�<��w�Q!�tv�"� ��7��7_��I�֢E�s��0���_�i=8�p�R)�)�Hѐ�e:�!���(��i��P{o���wk������T�^:=�ED()��Z�0�������[�Y���EO�g���p�TM{ ֘.B��aaB��{����VK����o�׋�l�;�ʬx:�<�n��⁙��.Y���$�d��}�,q%�w��l������2���x.�]�������wy�[V�v���A��.���q�^9��Y�׳��PE� v�� nU�[��0��i�T�E$BT�@���Y�p0]��A�ӗ�s:�]H�~����?>:aP��n��gc5�$�ڑԏ6��m��2����RA���)�MIC0RU��_XLl���\Ȩ�#�[�&(��دiW4��L�~�%�%�2|�rH)�(;{�|��<i���h��α��)|�H��a�ܝ����V��E<	9p:��ͣ�����D:��;n}� mS|������ٱ�}駞����-tl�H�;���r����U�2P����V$A1�])�qg�y��Q��F�0��]%�ԁ�1-kv��x2�#��ͤ2��kEvUL�s�n�.�~W��cY\����uO�O�@�H�Z�f�I�G���?�K��&@b�;�~g�^nNp�d�JU����>��_�e�����2�?Q��#�Hl+>��rG�9�yj��]y��/�y��7断�d~�S��>�ȣ��hc��ȱ5,����p��g�\	��Y]q�/)o1tC��t�	�L��p��ps�D07s	����d�^n���T��jnk�h�ŏ���S4��/Ӣ�]{Q���k�D���;�������Z4�.���k_CZ^��eJ���Q��#�%W�8��oo�c�o�Z��cZ��"Ag_	��Mj��/�`�ؓ����pQ.ߦ��.��dJ��h�DG↛K�����	q�ʇ��X�V�i�6-6?5/�V��m5v�tㄔ��v��q��R�e�^�i��W�\,����R��|���%p��Ւ�Iv��+�����!~������H;���6(���+U�K��r��)���>MK�"b��t��_��
�nU�W�՘��|��>ܩ,�������mg����>ť���~������Ϭ�/��*�7�ýc�V�(��Cb/3���%��n�2�Q����#z#�%_���	 ೌsP�B��ִZj��4@�sP������Vm�|�M^�������@���ȭW��O�^����@�#"�A*��H��U~��d����?�t�b���@�;�}�(7��T�.�Y�{��{���w�o�҄���~�8�5ـ��#A��s9!Q�AMX���m-
h���a��z�ODQ`N%�͌`xv��8�\��Z�9�D�f�f�8���4������,=�:���Z��m���@օ+S��Y�����?��e-r
�ֶڹg=����J��6�� 8�����`)z{�EW����&C��Z�`� �(�\����x�ֹ(3�0����q Ӕb���K1p�$�+��BBt)��M�`{�ȱ��}��uXsT���$]�ea�����I��g�h#���T��jI�����	*JoM����"��u�Iܔ�c�{Q�2���lL�5���NK�׸T���z�ԃ��GH
,R �Q�0��ө��e<$��ށ�/`\vm��|&:Wb ��W�zi9,�'��)�᳏⇖D�5A���$M�������V7��R��A���)]��lt�|'r��G�}�{�rc�����:-�Í��
h��l�|[U�7�������I��XI�����Y5�vM��;[���mi�{FSD!��?��M������J���3N�s\�A2�Tb�E���#Ɇ1/�~�i�*t@�p8|�4mQ��bAw�ݕs��([PqS�.��V������=�`g�>E���0�/
�T��t�ur2��e����&q��щ�Z�z(ɪ�RK�PZ��SM���%c:�T���:xD/y���Ǆ��ہ��+aˏ�	�����r(KAx�Q�=\�����Ӿ��+�)]��V��G�iȼx����A��
t���UĔ�\iB;�yE��1���Q6�Q����K�Ƕ���7CF/��VSMñ����a��!�p�S#����y������xY7�3�㸬~;�J��i=��i�b�-���!}�U7Icj�G�Y�:H�(��8y�Ne�K��ܖvHi�q�»X�C�X4c�YJJz �wh0#�?}Q5���0��q;�#A8s�~e?�-]D�h�f�Y�K�;,�]4B�Z�G��Q���L�jr�{5�f�jM���ֱ�އM���y#���RY�@�n%�6�2s����s��"%%h���2�\oQ��B�he��V�xy��/R�D�����x/��tV|qjb��p�n�� | ������(:��8��t��0C4�l��]�E��R�/|��̛ĥp�Pj)D���Q5}��=Ƥcq�@$@����B"P(d�H|V(�q�����E�+���=�i�Ƥ0�b�h�r�g�	uW)��ߵ`�+8�.]Q��v/���&������Z�@�@(OD� ~\��)��C�!�0)O6���l7c��X�7GEhY�������{B��0���0a�O���ȿ�D�>�4H]�,=-�P���Mu��;�`mΌ��ʰ�6v��8��߰Y��%�����Nr��U� �ST��z��Ɔ'eb���-���T,�1�xG�_�:<i��Z<I���M��:]N��$h"0{�f�z���7�{�;x�� 
vD���KZ��]9�чhP��_�a��)�J��&A��E���M}�ږ�#-m�!�˛���gw�Z�;���]�G%�&��g^��:L7��ko6�]q�����KD:�d��zɁ������#���J^R�
��Z;�,�ӈ<p�NJ�|�Bl�m��k�fh+͉����jM(�����Q Ge�&U�$�����蓈�X�vc��=�.O���#�&{�nOg�{�����B�~�sg�$!=z��9uW5*n+�̚�F�t4-PZF3 �	I�ÁX����Ge�X�ZtwM ��Hڐ�C�3E��B�n90�H�4;f�hd3��"�i���~ZR�H�$�^i3�'� (���q2�p��猪�e�Ň�=�:�Z�h��w��&�C����w���#�`oy�k,�I���7�����{�P�J�j�^�C
L��]�+�|K���S���#�1���r(rI"of=�*ny'4�|��U���a�>L�����{<-�_UEv1�R&��Y�	&'������uR�r�w�X,�F=�����Ҙ��Q�����uyY�{s�J��g\̹�l]�%�ꪜC�t��h}8ْI�����R�)�^eFd.П�&-�������lrk?"W�g��p��M�>�?%��K�nL�iWam]_E �/�&����	�:ơ� T�+���	#�$Tܶ7�sk�NjK~ݾ�P��X��L
��#x�Qλ�&��P�cꥱ�m���@�[hb�,L�{<�������gN<�p�JMKeᚹ�<H���O���AQ2:���Z�����g*Y����C�܀�����h���v"��4�ݴ���̽���;�G�i��=F���Qu6���\�Ή���~�-��:2�����r�F��Rj�4򈰋��!/������ ��$��Μ��&�M��}'�$`���!c�6��B4~���Ŕ��.�~�����u��u^׋8J�	r��G���Ժ��l!"��$�ʋ^Mf�����}[��h�XU�M�)�mw}ׄsDٞ.t��a�$�ؘ�X'9�W�TpI�.m3oj�F���&�������'���^4�m#W.����dT��&���y|Sު����h��K�Jd��_�"��⧟:�:Ѓ|�b��`���{(m�O	��~M����:��n�en�̞w�ݭ��	[4!�Ԟ��ih��Gɢ2v��%Ht+IeÉ��>��pb?^�_gl]lD;�S4���jbI�7���=!兣�]#�7ʅՊv	��穳���"��s0���-T��q�!S?�T<(ֹ@�/AV��Vʾ�FH-�P��R����]�';W��g{6Yo* �L����M�m��3K�V�?-Z�.{h�aWz/p�l�Cн����*rJ>%1�I��I8ɡ��Zw���ID�-
�DC�!�~y?c��}��<����vcŷ�)欹�����������2�?�>��Ӳ��7>�b'�r���A4�Tdq#vG�-W2
<��a�KD~,X+�.�~M�3�ǭ���kը��Ė����Ejű��2�h+�����*��W����C�E��;��2Z�~P%7�o�b��eP��j��r�c$���Y��n��� p��^�_O �yw3�>��"���{��ն�c9��ݗv�<ή\�V0����s5�,�-#�r�Ig�f�+PU�Φ򦸩_GW���5��y�
?:�^x�4�"��ϴ��6]u��%�ܕ��e�����<�]�8��d���3.8�73��{�8Lj鹅=Ii�@�#����;����Ę��=��}�4q��o0>Z���Ъ؞��S�v?��)0�@��)���36�l�Y`Q��	�S��`2v�?�L��&����	H}�,Ȅ~d�������m-���ˌ��&� �2˄ x�X�lU^��L-i���#N���5��w)�:��s�z%�F���8k��U��kff���h��u%Ap˛#�ԣlj�:�0�C{�WW`㼇�4�>�5��+\W��c�
6��W�X�;���&`���7�]*f�P��A邐�u��h۶�_����{��`�u���hʎ󇍪3uC�������_�����z�E��o�<{�5�kع���|/���N}s�6����ue`�wԵ1]��e�a"��^���f*p�jlh���X2�_��%�x6���+��@_Rz������ �R}�5�-��Ḛ��"�M�
�@�.��m|仛�o)�:Y����W
˔�"eɜ+��I������1I �� �[� ]���¦fk` ��/�z����C�<cg�lD�����H^��SO����[�����X����3B�/Ѳ�����U�H��'����̠ȭ�59�S7��_�xHn#~��VrJ�h6�¨p�+RG�����7 �=�C�5b*Gkd��y��ic��ވ��m�f�f~
4��ޔ;U��q��x#�����n�xyX*�$�B	������Nz8�Ab3�SL�HI1b\��!r���,ͥ�F���a:2����\�ha��>��i�V�,��/�<��z/
)��Bz�Q���4ʄz�7Ҝ(�vX��ԃ_+�p������
.�2X�S6�t" M�?_	�-*k�O��b�t;,��oJ�FP/��+�KG¦�[���+��MR3�q��W;��_P��e�E����c,�Yi\2ը������o�h���
u~J�_<�]��X���0��4�>��;��p��S����\����-)�T}�7n{Zs�U�мqԚ��K�y��|zi:�Io9��՛@ժ�v���9�	y�]�DV�Pe�($��L��)�5=B��\�'�Ի��x��5�&��Th�	�f��I��<.��8p>x�X-��j���A�����o�X��P��9�\���k�Y֢�7)���ۈ�X1�Ä������X1����ܩ�-��]$[~��"r%L�k�nf�x"3�����spN�b��G�2�������`�LYLu���?|ʮ͌�����Pafʭ��O�N:c��[�Λ�?ŌV���x�$?�cm)� �v𶠓,��v~�	7A���-&� �-���	�?*Ȱ'�]���yf~�5շŋw瘅{_d`�c���;s�����͇��E7(�����d�{���s�ܠ5���,y�+`Y��Kq����,�ڏ��!���k�0�#J&��랐3DX�"N	��Y$�W�
��䣪u�zh�4�P`�/ ��O��9CZ�i�=���V#m��1_�o�ڙ��h��t���F��Z���<�&��I��4��l．���ׂ���� Q�K/` �<9�F¨�wK��(H���o�����&��z��f*��f��bЃO��]�`Y1dN�|��`�Y���6��$�X��yX�F�$���uK-S!0�]Ò�F?�
����n��p����7Y����9Tft6'y�\�����[?�����tf���Fd�Zs_Ҿ��D(�Z��q^��n�U�7|p ��q�˙��
M}tl�;C�ĝ�����D��-t�D�3ZC[A]5��!,��51�Z23wEؼ#��
x_7l�oSHg�yBw�8@ϗu^}YG�����F�k(�l:����M�^;�6��r[ �ΐ���r��]d�%�UK��ǧ������E�����R�/Δ!%h��ٖ�����TPe�ԡH� �J��`݃�-_P����\������B��;
@m��@��x9���{�x:0�9���8R�$���`�ވ���1���x�����[��>x��O�HE2����:����|X�Œ���Ԍ�����ڟB=����*n7��$�lW��ݞ���|{р�ϩ�:�?߭|��&*�)nL/�A� �-��iR�`cϊ(�Z��y�{j�!qؘ��(����G����ঙ��̆KH^:���������R��a�AF9kW��=�!P�e�|@6���?�/H�?a���v�"M��K�/u5VjAY��j�ڤ5#MKyUԔ�b>�)�lK�ε1L�W��g�j�g�p�'���c����x�����=�� ;L��m@yKe�?Cj.j+j�iM'���sL�����QalSĦ��rm��g�>'�n�L�@X3�D��b�G�!Ϻ=2b(�v��5GXv��o�/����i��y�,Ǚ	tr�d`��̨t��q�c7��W�>��\�������K�q<��'��<��@�0E��\?l�]����.w�Vz��:"��i�k/z�ɚ��K�D+i�ۉoiL~tz-�z��Z�Az�����8�˙K��z��9�����L����N��}(�8����@e�?B��6̔[v�mu��z����뷌I��2���[g�D�Ĕ��j+9�f�P��k�su�Xҟ�޼���&
���'���fY�k*t��4�B#dgVy8��u;{ype�'����L�^l=�	,�:VL�i}��S�[07�l������e�j,ldJA�e
1���� ��p��*1�ǻgZN�v��s����*{1��ፈ�@"��:��7�<g��C�Z���*��1�쩇�5�����7��i���[�-U� "/�1J[�Bb�8_��-P6�b����f!�d�AމͺR�C�Vt8�ۺP\�h�2k��5��R%B�I�&|�����a�e�݂1�#���(�|,!�h]��1^X}�qRݎK��)�3��O��LƿK�/u�#��>��;Z'^|��r!i �?29��('�D�K�0	���1�[�7٘��3�vP���n��	����˿��R~_�ͻ�X��I������VM~�~ <�"�@ WѶޘ�v��;P�i3Ԍ�i�ڊV�z�G�O�M�ESD�^F�|�m�%O�K�vN�I�eE�[�+�5_��?�����L���WO���s����s�)��^�|�3?A0�[s3"~xޔ��+���k'��.���J�\�_ڇ�9>D^5#�^ 
�^���6bVP��§� ����T���͋^	���T㣯:�VF��	����Tж�y�Qy?�y� ~kO3rc�2A��P�G�R�)�⥭��NR�l����F�+"�f��5	�d�1:ds���3#��}+.�ݻ`@3&U٦�oo�o~	mNλR��
-9W�B�ō�r�A�p~������e�b�<�����@����g��;��O?���U��7}�_�;���m[�2ҌP�rN"}*���_70t�:�:d�i��+��wQ������t/�.w�$�TJ�H|���'B��_r5�N�R�]�;$�S�#���$��}�l�p.o��0���O��a̾�X3I3lA+q�˩��+��.�S^fu�y�k �Yjv�Y�5�>f:���yi:��/G�zu���F�p&�Y*Y5��ު7���]^�s��}t��rīOD#$o͵ݴ-����������~�Eʄ������<�-KQ��� ց��y�^z�\��j�Df��Ԣ�p�\6�f�)��#Ec���0(��M�jl�pG!��)�f߀N�~�hgp�����K�u����Pb�~?�Gz~���|2��3X*�m?��
�qN�2ŧ�fۧ膚I��K.�O����I���Yl�n:�v����&������[+�ã���@��0+�c��g':�F���ER䓎*�Yd>p�)��������NL�:�����jĤ��	 10���9��5�9x�Q�E�QjC�Y������#���c�hq5��oi��tHA�E%�����h�L�T[5Z{�nh?xg�M4;��k�jf�<�C����*m��ߠ���?E�X�P��
ȼ�L�_Zۄ]R�2���v���4��h�ȡV~�P|ykvV�<#��k�]��4� �܈"ɓ���c���-�9c��8v��*�����MnY�[�@��|����x����}+�����?���53�%Ǽ5=�vCx�ۆ��CJĿ�6E�$&�2����m�rb�֪K���W�~��_5�<]8� 2C������`��M�j�q�g�|Z'�%|��q�����i٪����k�y�*���s�������"�7�x"���Ï�Y��[���ٽ���Z�V�/�����Y*�r`ܧ\_���1h9f�1+��rl$�
�W񩦴��fe�-sW��S�un���7�\Nz�T@����=��*���i^.�h��ݏ:=��6d>�ɞ�Cm���bM44Mћy9�R@ܻ���Y�,l��"��Βs��C&���5���o7��ޡ��D�X�i�]�7�7��щ��C|����:	%e�l$�Ʉ'҆�~��0��Z+fƑ�!�\����g�v��m�?�K$�*jDo�L�QdWR鋎�@�)q���B �f�GА�����6�R�2Ua����~�?c_�H�����̷3�aƂ:r��U��^,�/�'���z�� ��8,қ)1*�H$S ��-�� �PR)au��x��h���j'E��P����&joS\�xyo"����c��)�pТ�H��my$�.$>��o����	��y}[��\��b	\�t$m�A|�<L�� �1�1Xz�`�{Iܵ�;�YW��v�5s|������:�9���Vb�������:%����b�<���		��Z�����\��K�"ώd��{�sL=�dV�����[�ᖺ�Z�c}Q�}��ySk{=ly@��֭��`�&=/�{��Fe~���ŏ�s�I)jʡ�D������|�����r�km A'�Ē?P��r�Iq~z�ھ�4��.�_堊DKK5�B�y���c�}�.v1c��§K?6hC/���>�`{���U�Bt~L'Z8t8�0ԱC��y��D^K�3ۘ��HR�g[5�,�'����+�Mp�����۱�
5&�3;��%�}[��bh��'�M�������N$�����X?Ȉh���"t�r�Kg��67�`��{��ϔBP�`��n��P잽z�G*���H)�S��1�IK�sMyШ��_��j���q�arNq�*T]v�����8��=�9�&r�V�Z5i�<}<��2���<��dI�+sYX��#��.Q�{[�rH�{H̔]� ��էEW�ӴN�-���o^헶)������ﰺ�[LUeҞ��g~���g��ԃ�'C�.��֒��J�iR��%2�a@�	i���1w�ŋ�4�k�εX?�E��A�)�탃 �k�e���qE��é)w��͕��ϊo�ھ�����޺V�
AO*���+Ԋ���ƭ�a�)��Aj5Ώ�A,u�i0�|9~������W9�1�X��A+@mD0�������6�A�gjn��H����c����;4T��F�9i���ejL�� 6���2�0�	�e���tD=~6E��jFX}�Q�vH{�x�	HU��!H��}:j�<�2��q������9Z���7T�e�D~�Y�M��:��52Bd"�fዀK�^�sH�I���Sn��*d,p��lv��}�x�g�a��[��.[Y��>���� F4��ȋ���l�f�A���Xt/�f�����!�Τ���I����ث��@��+���"	����返.������5�Ҋ�괠B�����#�ۛ-���N�1�����C��O�R�i�D�r��"gf��J,���W��0�J�I�w��o�66��f�����_뷻��K���PG�O'T>�g3�A������Cy���\��|��c��	�4sL��o3���+�=)m\�$5��$�c�-f�MZ)Lq��ng˔o�3>��'��/���f��p�6g0P��9�O쏨$o���ya��A��zń�1dS�*ˏ�����u�v������/O�߼pʓ�/���(w9��UXb98�?���%��W�|��xu����1�T1=��ck���VYqg'�49���u�z�q0���N�c�k^��~|>(��/F7h���1Y7�t6���W�mg�8�_L����Tj�w(Kb&\D��sʴ�����N��轀�#U�	RB�φ���b1�5�H��IM�
�NՈ�K�Jr���{��1�p��ٗ����<4鉌��6��Bꂰ��/hqbic>E Z�2��r��@�tai�dh�>+���� �c�b8'*}T$��oUrZ��hغ3j��2v�rg˭�d���,2�Y�u����ZÖ����W�5m��W�E`���E�����K��
�Y�q[�MC�c$���/��+k�j��r1����VK�����2��H,NM"f�[�e� ��c��krf��c��Se��G �5�.��)!	��nF`/����x{�ą�e%�`?�*���X�6���f+��j1"Oՠ�Z�\]	=Y�r7��}n�=�E�ӗ�*z�V�:4�=!���:�H�M#�c���̭ݔ*;n��H_"���f�m�T�����@�`ͽC�o|�j~)��[WH5Bh��>k���W;�o�8Pu	�$���Ƃ	ͮ�x�؋lǦ-�ʚلa�ZE~�j���#���P05VU�/�2�6ja�n	α��ۛRF�.�~o�@?�%i ��fp�Z�Cz]I~�u�5"��?`�PQ���>\��D�J���u�8��v����SZ�f��@����(A���!] �_���-�}��fl�8�LY,҉���� ������[E\P c�.��
���p��WDې�0�#�`c#S��}����L4��ۮs�{��Ѵg���(�H���a�-��(��%\M!G��&#�:��S�)F���_Z �/n�>X�'��N�N�F��4���*��;�>a�8���iX�Σ'�����Лߴ2���Q�O�;�6��Z2k�w����4ۖ�}G�/�+�!�K�����237.d�C�U�,Cz�Ū�W��Rc4����ݺǆ���\��H���>��D�����\R���E'^��ИX�D�K��; �d<������;jT�e�66c��u��Ļ���2^�p>��Yx��� �9�0�hX���^;�@�)q\a*�|=I���%vB{���ІQ��O��(�P+3��`�P���+x�:�U�/	-q�_9��Aެ��%�1��h-�/��]�H6M�A��SE��ۈ�E�M���������p��:�F���u��SRd��M5����e��پgfD��y�sp
?��ʿv�ڠ�̼�Cd�~��9)&��cW�'�O�/
_A����3����nxA1�1����f�.|�D&Z�E�ӗp8Crx�b���8^��
�2IJ �	��FtL�$J�è�a ����X�L�ҏ�������f ���w*�R��y.	v�{�`����2LCw�u�JdqE,4q�طC�Ǧ�}#U�p<'�h�}�p�4��3b3Ot��`��'t 5����LE'&D��'�!�O������<�u_[���#A/ca�M.�j��}������0�q�ڪ+�
h��f��v�ߛ,w�8�x��@�9���]�Va0|@���r@���Slq.41]q�3�^�x%�e\��}��%�36����,O��O@�C�s#�����(��p���TI���=E��{�*�QG[̺RfX�.`-���pbט�|�l���x����oP~�sPz�����O�q�����r�����u:�`����M�U3Y��Z�W���щ�b��e��mi��ކ�t���e@��a~N���m璛��_t=<{��>�!U��}�Yk��ܭ���z����3������=47m����A��������O>��Bzԣ��Il�=_�Y���P�{vNam)��!ʉ�kY��$@��鄂z|�E��OA�7��ǈ@��)̷�<�)-S/�| #� H�F��(��<�6�3�W6���� E|�.d�ܜ0�<8�5��)�;�H֌���)�N�[<���-�K��a�u�u���F𸩔a���YH�*P,�U�b�e�ջ9;N�c#�.��LՁ������/���Fy�����Q��\��`{?�՞k#�%����
�����1�(��L�Ag���7�f{�(�/ss���Nku���k���.�߹�����/�?hjG��B5�i`���d�3�m>qe��)��]���6,v��AP��lL��L�hNI�;��:\�߭�ѫđ���P�2�V��	��m������q	y��e��,}C���v�1H����Wˍ�Q\�D�
1��x��.*ش;z>*�l���  =WhD���P�f �qn�ݗ�_�%U(�ϪТ@Ӂ{�٪tV�Ϩ��t�K(����Ѐ�ɐf,��X0&G��B���<ЕGE4_�<5����������n�Ja�γ��!�I��*h�jS8�k��->h�x�P��qLx�Ir.S�j�^�|��� ��hC�z$8~��D+]�*��<��/S�CC������˪����O̩��2ϙ	���:1�'����xj	R��3^�3U��*�z2]�?��܃av'"�-m]�K*"<e!���g�����p��s���<�cy��hP�w��r���[�#@���<?G�˙���t��o��G�-Ϳ��aId�v�A��KQAH�X���a��YA��ȥh�.����t'�t�����EA��o`���"�l�\�_�����V�ۺ�������V�ފ:����7br�	���G�n�m������>��/[3`�����ز���ݰ5�C�rX
��?Y�-:	�ACH_�w��rƱً����"�5��s����AR����G:i��RG,��
U���cg��,��*������Oy�2�Lx6�]~4ˇ�0/<��pG<�.�o 8� �Fk=ۜ5��l�ߚ�B�N��U�HA�bJKb��݅�^StU����.Zi��	�pYQ�O�i�9m����,UTWE�!2��S+XYA��͓RHڑ�㿵�c5�C������$���YW��7���=��<�{RaD�!�z�w�<��)6���O��*��TB�Bd%�M��g�c`�2	v3O�;����3$��WM#��UBp��d���E�̄KT�T���69Z���£\0��Q��	���L�>��LMk����5�^�P���r��8t6�V��Y��j���7� @5%��_�}!�\�Kn�H�g-؟mR�����T��s�4�K����H���x'����d�k��#a��06�u�D��$�?�y�9(Y_�L7;_��h������v�W#���1I�:�W�`
�j�{C������V����O/�/�������g�u��'D�!��9��5נV3�`
�}�p�����"DJvN���
^���-�@"ϿD�#?�&�Ͳ幩3|��d!�����띰����zk�����?7;�9e��x�T\XD���mV�J��A��a����}K�jXf�L{�"°G��z��g��]i�"Y��f�E"�ܦF�rA`����F'd��3K�2��
n҅�G% C���؍�&t�]�V��#ևf4���v`'Z��\o���=�#�r�}�ا���͏��ٗ.C�aP�����r���A
}�9	�������|�s̬Y�i��rN�爥���������h�WA�kl�-M��2J�/�r�,�Y��6���F��7����x�Xs�*	��yC�'5?��U��Dp�O �g�r6X�ّיO�Iw���^ZCC�e�!�jG��	�L�q�쩻hӗ\��N��@�e�'���3��驊=_�q�S����7�S2�k����v��f�����>���֤\� @{(M��H����|�Z�ܙ�ӝ`� �]H�\���tw����ҧ�����m9 (���-�͠��j�}�՘}�;�Ҿ�UL%���YC�O�7�L��MƲ�xY���d6KF����	�y�&΢���lS�&C�b�,��I�� �!L诣��o	��ԙY/@��̯����� ���}�8���E��Q$�_�匢-wc��<�x=de�%�[մ
���<dq�n�#�ơX��@d��ǺHL��y�Wߧ�����hhF��5�0�.�=W�Fz5W�Ʈ�&�����f�R�Ơ�X\��|�;���۸�@ؒ��a@�Jr��ݍ�>5�X�t�n���Z+���:"`0�K��
����#o��:�i�W�!����u#A.:�q-���G���U�J��J�& H#K��#R�>ؒ˩��1�pD�:֫qsپ�M�����z��H�u�+8�J���D�c�@����k�q*ۛ�n�s:���OY���],M`��ʳ������t�hiY�|��
���m�i\�#t�s=-���E�s@0���BK�a�B#��t�9�}Q�ե9�3�׀�K�x7V�8�21(*����q���sB2���A4�,�p*�S,����qԯqߦIS�W�@Q�X���3h�ڊ��C�:�ds�!�>-A�|]�ÜӐ�{�B �m/!��XG����}<�ki��p��g1(@��oD���Q58)@�s��O3���-�$���b����T�*�9�+R��/��fDy~؁B��tM��w1]_Yzޗ�R�^׷���/����)��aV�ֽ��7ƴ��o�Z������1Vml���O��*�Z�a〭v�׿��N2�avq�Ѣ0^_�{G	�Y�k(}��b�b!g�]";.���y��'�M�u��>�ob�7<o��d{�	����H����*ʳg���	�;V��l
��@�\d'yd^��j>�R��J��U��)�+F�-J{}K"��J�o�Hq����a�g1\<�
5gG��Ӹ)D�h���y4�e!�<+Ӣ������ê'�� uu�'�bQ���\�5zDJ�߲�f��7�d�I&�Rϡ1���C�f���@�~�����$��E��3�*��>6����fT�|�D�Fe��F�- ��\�w���q��X�a
L���?
�PmZG�x��2�9�i7� /��hh�M��<DO<ȹ�kb&�	�������ibi�w.�,��^�I�'��H�jL�
��۬r��C^�	�._��N��E&^��{+��')����³C�3��ԕ�q�}M� s!�R�K�.�������\B88
���9�π(��J�k|)J�[��h���M�ΌE���c/�l-��l���$SY���L0_�/'�@�n�/D���ܢ)QC�-�2�h��&v}p��NfBU�˚z��o�p��j�p����~�Ϫ�+%�Ӫqw��c�u������//b�.рԋt����B�C٧-�M�r�L��6F��,_������_ ��e�C��A���qL����2Z�3���7�I(�E`�X����&�D��ޗ"��߻�o�ϸ�c������0�8�<pi��-E3�?_	8�:��`ǯUk�	���R�uOL{:<w�l����GM�֗�Gd�����DL�T�p������@�Y����.�
����7��S�9$X��+���2�S�`��#i�^!ݚ�0���^Ya�����1�^M4�ϱ�Pv�4	Z�2>�0�P@��T�R
��J��63���+N�yO��0q��X�,�!xVg�5���
���������)�O����K0�'�"�j����'����m��V}��Z� ��O�]�ʇ��B�1��t��ߐ%��N���*N���$��U�N�U�/���e$Lp�����>�"�7��Q����!ټ�qptm���.Do!���s}%T�㝣y���sP5+��D��e�A��d��ڃ��i/�8$բ�M��0���gz�L�Z�Qdv�H�m '���y+��5mw�bx��!��+��"Ӯ�U;�+�Yp���u�����X�P�@�  c�A��J�����Y��-�")����.[x;�]����J��L��;�w����/I'��H�~P�C�q������M�z�3e�_�0�?JG0Ρ�����=^�~���qvD�>n���*߾�Ȋ��};� �> yB�G'K���{g���j+��2�cה[���r����|����ar�L<� ђd������ĕ�,�^��:�-��A��$��G)x{FyW B�E'�2�©���=��)h%N~�D��R�cw��}W����J0���UZ >�}������i���p]e�� l�i�W��8` �".51�aTc/�.�p]�\���;�X��Gy�#�g��$����G�Cf����.4i�����$KT(�:�v���hڠ|4x<=�Q'����h|mk4n���#�4�
lTf�eq�e�&���E�[�Z���e���a��s�S�]t(���\$R*�)J��f��(��PM�����@���.���������U.��Ɠ�ܐ�i��+�r6��N��ͽb�x��d����;E��r��p�)?����A�CeN�8Pи�4t��L�� Q!w�Q2�U�;���2M�����wM1��З5���7�����>7����Q���Ŝ|�r�]�X�R�F� �?fO���9wl��D�&���m{��y#���ظ�k��uK�	s�"�o��[���؞�3fZ�JYtLf�����`�SpTZ\�����̑�^��h�Y5\�ȫ�D�
��5��t^����4C�\ǟ0�C J�Z1��᤼8}�徂����Tz�F���M��M�1�>St.A�Z�6h��r�)�B�V~ �j��W�\Uߊ���P�:�L����Hv�Z��"��>��(.�6Ĳ�H������ʪ��]<��h�u��(���g+��:�l��'�-�ۓ*{�R�d߈���ULW�#�:��P����i�`��w'Z^��";�rn���c�\v��o�����Cv���z��-@ #@��r�X�e7���=��44��Į<�wԱT�%mqY��Y�Z��S�"5� +@�A�h_��:�]$E��z�Y3,��B���[�c�v�is��"(^b4���vb"y��[FN�~�à����m�e��0�ϥV8Kn����!���)���ƆU���ɧ ��[p�R�B�k!U�넀�g����܆.19*(�m��S�̈́�̪�!2����nbdK�}�����J��u<�4 XKԀ�-����Z���x��v�����FS6!�sh|i�$=b#1:ţ���سNZ��FQcD��y�Ժ!���SK�Y_�
�/.���7AW���	�"���-�A���O8��\�uB����Xӕ���/�mgEd@+�T��*f�O�C:�HY��]�v�(A	|��b����U{{܄�ܭ�O��*�� 8��j�76�A�s���;WGw`E����F`S�=�Ēٶ������'��2\$�X��w�Fk���ݩ���#*2ۮ�C�c�u�������|��� ��?|@�"nKG�W��^�3h\��Mnz�/�@���%��dҘK�j$�mf�^�#�Ȋ�������W}J�V�Y��Z�#bX�@���y��-ob���)�O�$�vP����v��6�nJ��u�)��)��{�S���܉H=N�194�UN�Wܚ�ᰑ7�`�K(?ca�KV?�u�>|�AE�F�jAi�t��WQ��<X�ֽ��FBi���;�e�Ts��k���,��s�R<�������C0}Ǘ��W����	^��s2�W�q�ө�~�0;k��(T��Dɤ�"�D�;�C`$�O�h��+��)f�.���b�u��P?�KG#A���A4;��ԁZ ]��!���M�NҐ���3�A[_���C�I#��Pdg��o�+��?[��t�F;�]��5���5  %bpҀz�t��l�U߰�o�b>`uZ�/���	�T.�q2?sV#̸�.pKa>ḧx��-�c�x}�f��
c��a�)V��@O�P���lz���^�?G������3�6(�<W�w)
�wɵ%�Az��Pa�u�~�#G��nR��ME�d^�=}�=��.���c��ԧG�:l#�jG�ja�y7uqϬ���
�"�i��1 6�����7��Wq��9(��BI��!N*���Aw����#(�j�7<����$8vUL�%1Ϩ�殅J�h��<�S���$�ǌ�-'���L��Ϻ5������9сX�)\����<1t>
�˘	J��?��Q"�7�$,��g�p!�[j�ɗ��p�A��y|4�8��g��@�[�L��2���6��PX	����l��o��O���m�򹸉3�t6����l7�-hN5�D Ula	��?����p'B��}!.d���o�)�ix�U���/�v��,i���=��y�;�m���X8q�^t��q�W�1]���Y��у}�
Ɋ�g'�J�\n��J�8`��-?́6����u�x�F��l[bdJZ��q�J��'��:!���ҏ�����H�#hI�W�:�-\&m��L��<�s�x!q���x��И�ݼt\�%�M���*��9�Ў�?d��b`�p"g�Y��\s�t�"_ʭ�SϞ覐:%����l�GM. 
eKJ�!��Q����%�ӂA`/��d� [���J��JUI�ö,�Oܒ�)��$�FxU��M+$�B�/��W#���%>�Ќ����Q��aF$*��vR㲣1�����*�d��"v�f��]!@��-�+z��k�0Ru�`����;�1��c��x#`��^��4�?�fX��cv3��*�BRE�h������ k��n @iuC*��>�����
K�L���~�r�Z����P�0D�oG,p�?;�:|�kO��.�J?p;��l�7i3Z�R��	莡��/X����i��N�1�h�����#�%�+�;ߓ�q�l�l�䧨S��Ѵ���ɧ��hJ;�4/�v�>���l�D��&� �����LX�I�*��O�P�Y#�V�{b����.���ĩ��^��5�=y@����Л��^"���G���_K�\3Y�ٰ��f��c�0y�fz��`�&X�0=��	J��$}+vێ`�@k范�:���O�@��ٔ.>�W�8b�<����!����P
W����� @��w/������BHgɥ��L�'�~��J;�XM�>����qK�ݮLjө�3�?^
>t���c�>y�C�D�e���:�7��;�X]��QE�(��YzΥ2(Yi���a^����NTq�%Y6|�N����&��ݏ�|T��YtL�8�H>&7,��i�����ͩ�=m����]�������+KE��G�升9�@`L/�K���r7����CG6`v$JPY�mP���NN�YF �]��,m�HH�����k�nx��,�+�f4�Q�\�HSк�O�u�*%d ��"��
T�f���}w�/���`�?'j���q�C�]]C*��ʠ�� 1�bԄ��6j�:V8��B@����`�N?B��&m��	�f/?���Kw�t ���	��6��%�G���E�|�v`�X�+��0J���&^�����B���3%"'���j��\�ء	q�[8k��v^�%��E�]ې=�Fį�*)й�}5�@� �Xq����ן~֛73_�-@�"嘍Qz�B�������� ����67k^�������B�.�8��.����jХ���9	s���{+��y<D)���o��b�a��
�i��m#�n�������!�Gh��q���L�Fҭ1;�q՝��ҧ8��GX��Ƨ���+Tp�MvWC�����T���.��e��}�7�Ӕ��g/�S�.��J��xTv�q9UfL!�ަXT�01]g_iwX�hE,�-�د�|�_A�"�k�eB�k9��+�]N+vE0�N��}M=�+S��>pK�G`�C�<���7q͍�}a�ą�P4�i���������3J���B��i������voD�'f�����E0�m�KI0�����l�?贈�DKn�x�r�K��c1�/��2*�7>��=��:�}hF�A׿L�{��PQE�
�n�k(|�[��'��qTR�!a�����TK<����H�^�׺CG��-d�o9Bic�fO�M(�2�k2�଺@U8R�5}Tғ���Ko:�a~�b��j>�.�ǧcY)#6o��z���R�m3�`4ix���֡��Ȱ���W��������:T:֙ы2O�o��+(����S�Ε�1�Б �%��<=ʧ"��M~�\����"r{r�������4���W
Y����б�;���
��*<�(�ޙtR��q��|��?+��L(�k�5�ؐ��CJO#���lͳ|z����RFu���&�f��|Е(TS��Ge�s�6�#��{�9l���1{����  ����Ԅ���#$��W��i���jz�C���j�*ts�|V���-�O��о<���V?O  �������56O�`�n<�t�A�^>aGs#�蝍��|��?y��ՠ�(fyp�?\ǖ��"m�]�OZ+Z��K���CY�3���5�4�+]�t�h��ӄ�L��KE�����^��*��j����_�������`GSK�(���b�w����Y�a��$_'�ͫ�#�~������FA&�&$ �..������.�P�j������g۝���91��m|��-,F��<��V��p?�5�7��".���w��/X�oߩS�5�`��/�j0o��_�?�^v��M$��`��A�S�\ ���p[m���G#��L^2%�
E����eD��fl�Yw���sš��:Y�E���=f�c��K�y�x�i�d�b��_�o
�c-���v}��,�Z$���b-���ORnV�2r�#f�%(�	 V��G�K���UCeE�J���������w�L�tC�_���AZ���.i��s��D������S�ga)Lf5�h��N������[y@���%�c�+^����~�%���e9��&���,-�>�f���Sa'2j��ƿ�8��c@�x-�Ny���M�g#,C�_^�k|�c�N�q/a��RCqǼ�������X+:2r��J�\�h�2�Nj��pDѝ{%�%z!�z�,�G
�#׼�{�:V���Y����
�M�ﴤ	�v]._�Q"�K��d�X��%���2���<�-9�~=�CO|F ���G\0���5��G)b_M��M��W��f��"��Y����I��$�f"�ܠ���Aq��ZL��7eϞ��>�%�4$U�kRW*T�����	�m��g��k�3+��_7�I	�Z�8�u@� �����3�yڗ��_n+ۧ�s����Ϗ���ۺb��f4�T.I�����?�]�WE����\c��=�I�#qh��e}`ɔdS}��2�F��t	:���2x��Ѷ��X�F|�Y���^��Xq]��j�pM �������n��,���������F�&�Ļ+�*�d��t+��Z�~dI��!�v�`��(i�5���������Hۥx,;��S%���c�n ���+:�trh��@[gR�*$��8뇎Kf��o[1�[�V��A֊w�	,�@�!n��Qc������:��=/^�����Ve��/ �}��&7_P�a��)%8��|��kBct���;T��6��b0mW�uv�2���
t�d�ϵꪦI�u#��:hM[F�L���q�A�h=헆?»��$��GC؍�������|�@�P>`z�>}�y=��&�'�P+�w3
�r��V����+a��U�%�/)J�A���d�ڢ�D���ȴbJ�]g�m݃�_�uˎ֡�����T^�� �H�L~7���,��b^%�ͦC#*o�j�����o���ӯ��m���Q��u�*�26�V@��ǾPBs��4��c\�w��z�U�"��99?s�F?y�޲i��!׾23���ZIzgc��_Ê��P$$�޳5J�G�\d���-�"����xT-xCq���(�y���3��e�E\����Ր��#n㾕S��^HV��9�\,��I�N�"��^��-Qc<:Y��CQ}-l�<p����J3{����'<8��^Ά|�>����+�^`!Z
p�F��IӚCDp��!��K�ʂ��݆I����{)���#D��[�'�N�������X4W�\�R��^��UXh�E����-���}t�X�8iT�q�A.y�җMwS�X��7��4^����ѝ.�h���<����	"9�E���q#�#���11���5�:�	R�E�}Q��?�]�G�du����T���T�h���G��F��\D�d�o�I��ދ��p�U����6� �yØ�O1�MR,�<���h%"ͩp�������g���Nx�Ӵ^�u�AN���KC��Uރ�׹�@6q��ԩjk����	��`1�2�q�+��idJ���ItC��X��~[�\���V�����߹�l��'e�?GKno���袞��ޑ� �����+E�d)�gZ�y͸߉��!�u����l��k�:�j�s��S%ų4r;�b�Zs%�xͲ��G*���7x6�C�*!净�yH�c�BU�9���Q9��>AȸõW"VaTb[�rb �[�v�H7�2�{v^K��p~��_j�g���46���Zyt�!O/�nb:E
�G�%�O@��P�Խ�����9H���Ny���������Ȃ.}� A�J���V������	�3������4��?)5x�x����޾>��א?s���&������T�>���gQ_ǔ	�j�'���{[V2��-)��`�%�[�
v���d�������e^�o���cC?�K����	��gϭK���)�v���9_�I핚.|�t^�0�P#�:
}�����1�Vi��$0Ҽ~Ҷ��
�r�B��۳rr�o����ߊ�>�q<�`%�F�uELr���J�Z˷�~�WvVS�u��W���_+�ݙ4��� ��X�mp}Vܼ7�V!��o�EL�A����H�l�p��,�ɲҙߏ�AApΪ�`�N� f�8/�ӯ55��H�9HǾy|��I���(��a�0��ju'F�!r���Ry�dd��G\h���������Ip��d+�ds��W��Z�Bo�:e�z4|Z��)�����հ���_�4�Iî�HT�l�m�ˁ}&��oN�+�\$h!���ڈ����.7�b�}I:��7��D5-�Yc[%�w�k���vV�n��q+8�V�}W;�=�Eǃ' &���_��]R�ԇ6�ق&��c�4bU9: ߺ����Ϭ�O^!��K�����}�%81��X3Ö辪���}��,9�G_ ��
\���4���1R��g��T;��%'�?�L���~��$��t/|Z������Ԣ��؋	|M����7gVO�w^�i��JҤl���y�)g��7�h��L���|e��B�o������uS���Pq�O*�_�N}��s��P'r+tRael�*�sW=�V��;�Uac�!Md�� �iI��[ � �&T�H�2���S���D٢h����j%`�F����a�z�B55�<�0����+�l�&�Q<��Ѡ�²H�P`��&��;��9�� �Q���"psc�~�$�yo��A!۾�/�DX�V��f�5*�౬Ok��9�i�=���T��~�I�X�����"�[C؅ы��6�4�A�Q����K؈9��gT҃>h�����L���XW�)T�p�rS1�ۡ��:6"�$�^�^�l�Â���B׾)������a`N����F�ȋ��Z&�Mș��ɐ�}u���F��+\0�E]vԺk.��:�)�S�<�El�d^X%���G�y��5�/���ȣ%.e�w,}1v��8h}k�	�JaN���s���\��Jr�E#1�5�H�����Z �>�Ȱ��:����Ɍi��s仫��<��Θ��>�>���]I)}W*���b�p>������*�v�A-ꤔ���k���7��'N>�t�)������Y8D;(����v�،�DZq^�r"��5�'�hC��Ψ⢤q���3y�oA�A��u�9/���VaP�ċ�"<��2N({���km�����9�.�h�H���(�MOվ��߰��������[A��1c��Ma��RFߊ+�EWP�1�G�2�#
̶t�3}9A<؇:��(�<Nh��dg�(d���8J�Ҫ<G����$��a��U��@7����EH�h+-חT0�<bUH_-s���
��ڞd�T�;�g�� ˦:o�% �J�L��ۆ�vpu�y=J�,0���7,��{Ж�A���K0���m���;��pD�^���ٛv��;�f��ܴ����F|FY�"A��׸R� n&��aK�����>Ǟ&��7�k��r#�3�@���Ǟ��K49�I�������<[˒�AM���yρw��7)v�b����������O�4�~�9��3%WE�j8X8�#�	�K�8p.���b�9ؚVp�?���c�ŭ�-0��.����9WK��_���M~!�&��p��GO��
=(��P��(����}GP-ڳt��+DFH<.�Z���B�~��+W�*�y�w�EJ����0��5�8.�U`��RQ��$
��
�1\mm�<�O�ouu���xٻ�$�~%��م��^w����n-!�O;�t��zEVt�"Ү�V7�k��Z���_�~�zc��q'��2!#���^�1)93��l�������Xy�����So���V�����9���!�S%N����(��41��2Wi>�Ö-JJ�|����.��;�+ؽ�E6�� &��X�ZRT��x2��n�x5�U{���Q_����TH4�4H�e}�%�C,;qW���nm�/t2�j0��R����`�T
�6�a�/����5 z��ℝw��&�Q����g6npH|�+���F���-��ʨD���H:�^Zc~',}ᔊ���+$�"��|q]WPB6�v�� ��&���-�Y�,�?r"�R��f��J��q�j��_�".'|F�n���~�x��}-G�J�ؾSj�k1�q�X&��œ�C6��&mR'?xL�B�R���Ko\z/R~	���%�x�:y���ea�z��2G�9����<������'�en��ص���6��v�ڸ���ѱ[�����<�F�U���Bd������,�U<����7� ����=��Q`�K�R;mu����re���O���݉^��ĕ��M���q���S`���A &7�Wb�z� ���� H��`-�� h-,1Z�d��tƬ ����
N(�����|���ڲ��H��ګv��l�΅�iU�B�P�}���(���QP�������*$�
^���/S�Gƅ�yc�|�8E�[��\'=��a�"�P�ĺ�J �������+*�ށ�,��~�.~5��2\`""~ˍ�.m0ί85\Kf��I4�5����"��a��
U�ÿH���u2�$`��}�?��ӣ_A?����߭ꈆ�&��	m��
G����g��d2���i�k��#����;�پҶm?3~<�mvoT|����_V|<���?L<��Ӂ��ӈ}$=����Ә5���@/�����0�$������.wc0�}�	���>RC�d�,�?�bL|l6�ӄ'��A�)E�����6�O<��K�@��I
���3��QK�����f-�JS<$��ݡ솕xE?z�ًn�eU��&��B��k�$���⣬AUH�����K�̀��7����sҷ�K��%���~��ȈVB�F5�,ȸ��_fEo���Y^�,I�~zQ� C���^�d9�m��?�B4
��9ފ{Zݷ�R�U�U�E�)�R�����׍�}��iF�õ
q`�y�9�W��OyI7'�m�2��$���1ND��I�{\չ��6l3Qwǡ�'�����,��&FS��kn]8��b�U���g��r;�d���m�3�7]0Cp����C��h:�����\EGp��K
�Xx��W�%R@gb�����m��C��qQa�	E�	���5/MC��mQ@�lT�����OO�u� sY16ve�/fd��1�&�>�v-iB�ka���	��i�dX��<�]��@>)s� S����7�Ӎʎapه�#=c�O9�Te<�^��)���%�HYL�+�Hd��^ܻMfd�9�"z��V������l��߲Ča�L�K�L��8��=<�0�-.^�YeMm����P4N_�,p"�G��Y�C#*%��5��&a�-[�~ �@9��������Jq%��([��Am�Rك�qL�J,��fؙ�#)�|�-����h��s�>�Q�9���A�eY���҅i��(9[�"Sv���l:��Y�j�hx".��(��3����wL�-��xx�F���,��'7�XX�������RL���I{��YE�e����!
,j�++vuY,�����O��"o�l;,|�,��92u\�V߳�d6�bS�g�.�� �9�g�	�af40 ��X���0`f�~
X�iV��R=a��C���*p'��*�i�>i1�o��i�haOv-t��_�!���Zr͆l��m}T��/+�hHe:���=�C�l�/�إB�͌��P��n�Tt��F%�Et�Mk _.�\ '�:lP�g��5@���j���%�8��$ډ�~�^l���}Ai;u/	�U}�X�^л�c�����(1܏�^�JYx3���[�&�Ύ��VNRH�C�8�$ ��MSf�pL�*�t�U�\�')x�B� ��Vj��qjD��nŏ������*٭v:KH�[:�&�nX�xu�VR�ʀ��}I8<sd@\vj\�M
<9���}�lo/*w:�������>�Dn�'��C�$��6{Toc��="z��v!gd�'Y`@3xmvxG$��]�`n�����"%�3��倢�_�R"8K.Ps�Pu�j���%_9�ul��ٟ����,k��*��I6!� s�cpyyf�.�^p���e�!��k�6o��:�ԯ��f3"�'W���am�l)IK��z�%�������f�f�j�@��ۆC�he�iM��dt���2@���˶U���>�w�F��%�JC���B�'T@y����,�OՊ��F���n��6Q8r�&����9u��F��ݙ�VO�j��䱻M��E�^�X��!��Ϟ�I��z7Ա�á֐�y>��qُz�xꏆ�~)��V���zt4G�/j�r��ݨ�+&����ZS*�K������Ԯ��Ve��j����m�\x��\�ȃ%�⪣5�V1_2�c\�aS0nP�IU�)*���A(c�/��E'ҧ�3e��_e��w!�����R푈|*���eˈB{y�
�:S��gN&�r�jJ깑L��o-'� V��@:K7l���	7ң.�u����)���!p$�\<<��4hה�79�"�_ �RP�f�Ҫ�y�իq5�HU@Fw�g�Hs��!Gp��=��{��	)6�v���p�HbϦe	�CΈ�I�`[�[L!X'G���ܫ�ެ��J�}#��e8�����S+��x`�rm ��@�a�{�����[K��m��셔i�-���!8M��S���]�����7�u�����P�Ey!�Î����]I�ϳ;�$X'?���^�"�O��_Xq����)\��{���)ۓX��;pƴ:�����HVn�},G����m���&�m&���GSc� ^��	�l~�gc ��8u��ƥ�B��CH�Z-z�o�C�bg��;�W�jj��mRɅ �<�!�1���h�=54�O˚R��WK�T��vPOZ\&��(U�f�i/����G� ��hf"{������P����]�p@���>T;���s1+h@Bp^�A8c�<��݀�'�yjeU�Y]h'`�k�Q�>�|1MW
�N�,�Y�"��$��|1�j�F���P6��S�!��)��er�bRbB������0�n,��!i�vⷨI+��&/48�N?����c�F��������:-�ڟ¥��E�w���p���)gG*o� ��5٠���k��0?��x'�����xPi�{��$?�N/gG2�́�7i�B��	���!/��	��TLn��`�c�k���OYȵ ��K�0  ����ώ��W��D}�0X����}�0���mR��SN,�Ơ���C�̦��7��);������3J��:d��#��y�
"K|yd�kh�aDj�>v�aC��O����6�����[Fh�7�/9���8-=_�X��0c�1J-��wkrD���v��6m��H?�&�e-aBژ� �7�hޅ��i_�E$#�\0���x���$>�ٙ(@�n֮=w�Q)㋭�L���$��x|��ø�U�Ѡ�,��7�K��Q�u��E)��K������G'��и�9 O�����+����P�����v�;L����h�� :�)nUol���� ;�-|�A��v��⦅�q$ ��Ҕ�!��������1��\���Ո��<�>%	.	(�F���HTS��e�{
Ȉ�V��,Ӭ(l\���F�l>��������>�M��ڴ��+���x��L�w˃�Fjp��lQ��1�>��bb�	3M�_��L�Ra�� Lޥ>�q]S�Q�6x���@?x�c��|/�>ȃQ�)8�� e�:�e�EV�� _o���Ac��y�	���:J-O-FDݨĄj��z �
%���ږ���%_E�&�z~�0'(n椖3t<�"3��Ag ��
R���V�n$a�+)�Eߴ�4���N�H�C��<l7������E\%��-��s#84����2�Z��A�R�D����J���4tmL!��U�)�M-��?�ċ5e�z���Jq���+�1D=$g����8O��<9Z3��p������S�����������Ĕ31�M������ի�V.��Vs�3'\����I�'�5�ګ�G$o���le��Ӟc���l�gԦb�*[�xnl�( ��ƞ[N��$#��1>�ЃA��.n�!y����A��pԙ+���{ �?��r��P���&@���f��L<�Ј+����n�1��������Y��S�`r�	<�F��O�]����dRͮ�D��� ���� �6�j��q�&��-d��G���6S��A��ĆRb}�<O����JΪ!��+�R��2��
�H9}��9�pM�
�Xa�U�<>7����n6���wQ�H�y=�FL7��	�J�s�f���g��;>ժ8��%jD��G���L�iͶ< �����o��Qg.�K�8�
=Vz��w�Q�3�r���݈ѽn��W_��C� di�D�?�δ�Z����@?���:��a��n$*�e[r�A,6�`>�;_�J�G���x�r�s�z�p�Õ�Z�D���pQ"�פ�a��#.�8���H�P�?��B�%Z��jP@��D�v"ܤ�՘*� u"��nZ��y���з��߶�$�bR)�U���j�W6`B �ybvf�s���V5q}���k6.���o�蓕��E�=��Y�Y�W�l�nZ�E�oMSBO �_P͌�r�m2�b_������"}�����(����US���0FK��	�~�Ko�&���z�>��ޟ�gԏ�W��b+\F't����:���~U�
o�=Ɠ��b���#�9�8���eY�ȳ^�Ũ��=S�fg+2̗Y	��Oq� ��`":�1)V�Y-��/7���n��*Z8���ؿ5'�a��q}T�KlT%�d�
�A/X��TW�Kط��Z h�uS���)�uLrY�z�/2�N"(i|
3�]��l�~�OP���o�W�i�<��>׶@Z@�~�����Qcؓ����ܯ���4nv#L�D�8�Q����j�@τг
�x�D�m��)�c}jX��嚥�PϏ�����{����
��Ƌ��=R�N����ľ4x^%��֚��G?#�K�ik�}�Q�N��r�<�#N�
�\啥>;N''�E ��!'��:�����1S��-"��^4A��M�R8z�[����J�{�.x��P>� -��G��[;{Z�"T<��{�f|M�(��5p�ɲ���Q��V\������q���&�yA���W�/d�Y+О�����/�^�1l���]������D�n	�NCzɢO8]"&�w<&8�s�-�6=�J���7/HK�cKw��H�sT��0Ѧ�������J�Җ=��Pd=n�.���ψ5��[U���3�*q�?�L�P9B��g����j7d�� {�l@1
���0zG4�z=|�� ��JH�	Rw�?����*=P�eC�;z�B�Ͱ�_{I3?�ͯ���7M����~1�dɆ-7l�v��S+�ϗ!��V��	�)M��b���ׄJ#O�R[ ��ϯ����C�G��MK.��T���bH�3���k����o�*/���v6�k�6H9�ڠ�+��%5�,�8�$�X�qN�D����i���GwEW�M�n]�Q8�-�H�NH�7�\���4Ҙ���<����@�B�Yw�5N������q��;����~R7�Jin�{՞U��	�#~Ƈ;e��LȐ�~�"�H�ʞ4�rh�{�WYЌ�#g1"� ���̩.bVh%<ȶ�\�	$+��0��U?����p?5IN3��0��<y���a���6JC�GE��k��k}=G9j��ט��ߑԜR��`��	EL���!��"V��6�Х2�ekΠ�̸6��{2s���@[n��Y��|�y�D�݀���B����G�_����n!�S.O��I��ܼ������5y^9��5��T=8�{0Հ��9�w�� ��(ٚh&��qٝ���P췫	a�H���K����?p�c�O����Q�}��ŨO��o�p��m�D��Y���HK��M�e��G�G;x�? �HKz6H<�ԐM�����~6zȉA��ţ"�(K��4�����ˉ��[9���m � v��	���z�B��N5JJ=2������$���v�l,���LV`*�{b$ƻ {E:l��Y��f���]�3n��cg��Oe*�V-|�P��cN�2�g�u'"+���`�:�/-s���1�ɾQ���NT`���� P��8����)&��m�"��~	.ԗB����D��׮�Y&+���d�g$ds���obj�lV���S���ώz����p�q$�������v���-?yY<@8Z����2�Z;�;k&d�Dݻ�sz��ޘH�ST���5ȵ�N�t�P����yHbt�4��6�/�� 
�aoJֶ�hWm�N�w3Td�3$eP�`��i���MI��2ē^$�m��B�"{m'�7m_f��I����N�#��7ڪ/.�o`�����5��AD��;/�$7݁�^��#d�I���fأ���_� ۗ�_��g�Yjv-�����O�#1Ck���<?��=�ʲ��� ��.�m�V:�֜|��H����g��$��Đ��;"Hj�N�!�8 �	�K?X�JF_X%9�#S�\�k�CX>��s,��h�Gp11�Q%04����?�P8
Y�s3H��ShJ|���?Pfh�Yۈ�_oRް����9����kr_�o\�\�~�&�`�47�6~�_�G��(�<]�Ņ7�;�=_����Q<a�l��{��v��K��K�<z��ݦ��(P,mcy�+�S�<\2��Ѳ��%1���m
s��l��[S�|V�Շ����Y�d�V�Lӭ�Kp#�/_#��dc	:v5m����k%"��!�<��Z����]9z��G�Jt�N�@0�0�t^fk5���x5��;~��P�	�hӠ�Er!k�� k_�ٶ)	�\��=��៏a�=����q%��CN�:�*lm��L�<Ơ׻|&''�v
��30���1B؆N�����~�(%q)����1c12;Jvu���],՝�|Y�P[~� �}M�b<�p@k�	i��B�f�&� v���JC�h�[ `���|P~�A��j �y�@��Y�0nV++}"+�(܄�|~�Vě������6�oB���ћ�KJh�Msmtt�X�(����͒���DWW�$�c����zqnw���#���ίP@�8th��w���c��q�\ޏW%^��Q�t8��p�ֱ�?�z�&á��A�RV&~x�p�wʀ�9�J�<�=���i���w�|?����P�d���ݰ�-�W?��d��'���j)�Ӑ��u�xhz	���_�! .L�����c�;��e�ī��Yz�qfuS�$S�%�<�$�
g����7ր�4��[�wN�G�P�^;���`?`2$�۠��|��Zp������kמ#��Rrے`���l(���9ǧ��`טy���Q���yь��3y�ϬȮ%�w�	�J��t�z�+E'wm�]%=4�(�ݷQ���^1�Y{�Ac6R��61�&,
��i��I�ʸ3�ԉ��o�H�/ +�_�r>;�;�u�"�S[�DǱn��f�:��uP���՞����I!6��CAKݿ����+�g�r�U�m�ii:�^�B�M���<�1��;�\�w��������
ƺF2f5	JI����=��ज़���Tm�t"��T3����~�}��kR��u��_!,8��y�h%�}�M����}	!���� ٻé���~,��jmÒfV/��vcj�<Z��ނM�hO��ӳn�ho-2�F`�!2�ק?�Z��|n��&Z�jZ�B����S���q�,�(q`cD�hd��ܒG91�miD<�F��W�{�tlI��>]�8�£�c8+�_)/��פ�b1gh ��\�Қ5�v¿���-�\r�Ȫ,�o��d�uŊ�6�Ax�G��
d�Z��mT�@vC� FB�|�O�D���
@y��5�9���	�>yGʆw�ƕ�Z�pT|d`��	��zv�Yn�Q[)#ՆZ*�/X��J@1�_���z1�O�8V�
�XS��{9;���.m��s7j��FΓ1>l�Z:L�˜�2�ygDJ����l�� �@R����C��d7�?͋�^��
Oc�����í��.tCn̽���4F@ш�[����{b�5Z����(}@S����la��^3*L4<���8��k"�DRl��E9.�+c�]؎����~
�>,-�V�_{^�`��$q,4��g��.y���o�k�4�ҙ��F�����J�IC��#a��ΗCQ@��.�X���p����6�8$!ܘ����1>����ƯfYMR'��PA���o��q������O�y��h��q`
'��Yv�-�/�\8���,�G�O���cD�%�%���Ϣ��x�r���X�vg@J��~�ȥրB�0��YI�Q���������-���\!/��d���)�&�i�f�pX���P�:�!��3��e���¡hrj�lH�F_�cȃ�:U�d{�h��Nu�~�D�]���< ���4ʦ�2���BV\h�Œ�y��a�[=4_ϛ�<$���� �a�_/Z�m��	L��3�"Ej3�[#	�Ӱ�'#��+ä�d�In�X�����MސՓS&7����������2Q�3���g���bd�%=���g���'އ�FsZ@������nc)b̼�{a� ���b�
��TV���Q̆r�ݚ��Q.	ԥ��k7[g�����9��!�y*71���Qt���I!T���1 ����>(81�+�,���q0�ke:���~K0�vs�F��C��3���(lM"�K�<i ^L������l�����{�I�V9���Q@�j"@`��t�H�����ʡt��A$FF��2�Ѱ�n�%ŀ��9/�ewf�%��r�lͺO���i)�Q d��*=���0���C����0�5Y�s�W,Y�_ 	+D�vE�ĝ�P����}0�`9Pl�GZs�{C-r�HZb��I@�%L�f��t�u���3�ͤWD	�T�
I$j'9�B�B6��`[k�k1 3,e�C�<cb�X�e��{��Ӕ��G8�C`b�A�V��\m4t�Ȍ�M�;��>����z�pH���R���$�����*�����߆�ʡ"�հx.��V�R2�@<�M�ÄT�P��j�K��&6~_�K�|����:���4ۛm%�	�o���6G��I�b[��ۋ�~���K���|�x�.4��>6���:��Ss�_�J��8p���w���.�Y:����,/ǿ�� �\Q���"h���z�vkPF�<$����4�'��>���H^�9�����}Yx-v:�J:�r�������d�R�-;"�
vԿ��9K�hj�q0HX�{j�9�\���?�y�y��L���OFT�l)b���%�s
x���t�r^��-�X*!��}~�Vle���Y�BI�~�\�"��R _m:�I��M+�P�e.q���9_A��`V}Z���hg�������'t�-�{�V����=$F���=d�i�.�x�=�*9�[�E�)}D��MIʔkm�on��0��*b@��S�5"���� 3=��r4�{E��$�Rt�}'ey�%)tE���Q�U��ϐ�:1~?�*�*�~�ۍ�7��9/��w3���S�]|_�%BU�g�Z���oOe�~c��H8zJ�^�_N�1�c>�G��uj1��ۀ�>�(�3 '�Q�Bv��c6H�K��۬�<��.�X<H*@Af�܄<tq5�@q�=�y������xo�1�q�$S^�l[� ^x��RY��9dv,��±ա��4]tB�{�V����{�QEԔ�p�ŭ�P��ZH��Ϗ(9�����3 ��
�G�+�P����j�!#D�MF+�8	�O�}oл�O8C�{bӂ����s}G�r���x=���P��z��Z}/��J�u��P�3:c�3�!`���9e��<pB��<*k���~;1�i$��l>�3czU�BX�,���p��3�Ŀ����Fp���o����cJ����VS)}={�����d�#��>W
������CY��$ɻN}�lZI��q܃����W�>tv�A?Z�M,�$��xR���?�%��F��3�?�ֿ�N5i���S�.���7��x�0N A�v:�C�gET�ճ�5].�E����������� B�y��v�L�Ӿ2��a�mHi��^�N1����'��;Tv�c��޸l���"���d�~��B�Xs@�*�g��R��Z-�'��9�p�%n��}8��Y=����c[�a�CV�\��(��gD���CGy��eQ��(�����W�rA�d�L���XSv0�C�ZF�Wa�Fq���ȮEM�F�n��| o�Ȫ�&h�����0���fK�|���j�u���q(�D�C��hX"�P���w��ɇ$���T�mO��u�d��r�����y�<�����Ǜ[�AF�
����D�y��d@F�r�J�͎U�W �ja�&#(Lj��E���8W]О�����8#�dE�_-K�8��{��J	���D'*�v�/#�,��>��(z�"g����v����|%\��K��a�?�R!cT3���;\$�ź7����u�k�,u-�	y����JǙ�����0�R����O��C9/�`�9�*"�@K�*���U�5N��#L���r��� |���	i���6�Be��9��l���W�J��}D�I�Λ'V!��y·x�" 
�7�XPs@�?����Eǟ��B��1DvE���mV�R79���P5���Ϭ/b5@���w��E���;��x��<�V��Z2��iѲ�mH���:��E��Q%]����J\�	S��eJ'�nU�I�5�)��p�������|Ol��O
�"9����{�l#��{=n�R��*��D'D�2�+�A�P�a�毵�Ɣ}��ԮΡ�˕KԐ��Y��o�	E�J˫ ��~ͬ_��?~r���pF���	}��F"�4��_<N�����Td� WFJ�!vK���R�nq�/�z�t�e�1�/J�PT�%�P�R( ���u��7�)Q-���)�Rh�&�e[œ�TF$���X�����[͡���pr���B�Ο�ۜF�ձ ����횫h�0�=�?b�/o��K��?��
�_~2L�@t%:2�F���Xd5�����=�|�-`+���%N+b3��A��E�*V*2�-m:Ix0�W�I��c���qJv:� 2m�c^ro�V_���3�������B��BKpiA>�M����݅�ح02���Wdeq�(3ow��,z%A�T�B�!#Es�����͔g6c �1c�t�&g�Ę)�� :�WE_>��-�;�d�)H����0��*OVl���7D��G���9F�	��&iIȯ��D&\������gؑ]��ᏨGYY�|Q/�ȣH�_W���Okzo'�
�!��	�./�ZEf7��8��8(������wmlfB���阒�1e�kлR�cօF�jc����;&ZTƛ��Pf�c�ވf؍఑<���c���6_��"z����[Y�x�'�u��U��)Z�nI�y�A�z9a�(���S���SSQ�E���!�>�{%�rL�l�������"�RϏ�w��eZ'FZ@ߴ��[��#�Z�S�#H\�M�n#ScP�y�J ���p�Y����y�-1!�9������L�2�AqR������=s
j�;%��9_0���:�F��)j��I��t*=+42/���#a3j�(@Lu^g��Y���|��/�Ad�=��Ѹ5��	m�S��/BôEU����d��^B�y��������l�^F  ��,\~p=���cs���р;$�DW`h��r=
L���o��������������)�iF��h�vZ���1l=���\�l��6��o����6|��N���{;}�:6����K&j�ȩ����o4�.�3㴄�gl��]���1��wA��~8����~���� �� Qڏ���/}z��;��S��E<�K��2��%>�m��yq4�[�g3�JV�=*�{��׺��J�hWd�!��yHʒ�"��V`���I�5�`8�;4�a�޹K|=u�9k���SK[�p�K���g��D>�x�~s��G? ��C8+˴���ˢ��(nyvJ����iF)A���^N��s'ْ��q�N���ϐ)Kť��o{��
4Dn[%����$��?%H�N�8䕆]H3�b�&@ o��@_Y���`��bl(�<a*m
�!�%m���=����#��f�^Wn��"��N��PSoYR�u~�5�����H%��a�&S~R�BG���C�6�d�J"������G�.�g|	�D�Y�����T��P[�}$)�a	{���}G����m�Ru(�8腾N��g����e̼<
`B��~����_��)��g�ۜc���c�Z��jZ���N�� þF�i�]���$9*l���t��[1�����:�c)-�0�T��j���r���׀�IO�8�wP�V�������`��&-Ů.'�4�jc1���ӫTVuD�D�q�5��q���\X�*&��d�5vU��0Nd�f�R%Y��.j�jg@�E���)�9_��kt��k���	z���#n�)Z���������P/t�e���m�U,��HH��1Ŀ%��׸�[�� ��-�/C�Ŏ�>0��sz�ۮ�����u|":Ur����܁��m�(K�!�T�]������0�ohz�`�0K*A9ё��?G�?��kK�0r/ށb����y��+�I(E�M/h�tŌ5q*�N�=���d3�Z��Sj]��)�b�a8�	(֨�]�]4̂ul�SӴ?���B�W��(���T�w�b��ok+NnO S����U�і�݊�z�/{���6�1�}kP����āw&Q�T�}�ړ���Ń���SŹ�
�|e%GY�������Z��f�wZ8���x�Ǐ����Ë�]Ǒ���C��+��_�k���U?��^�$r�G^l��.*9�
��G��	�J���i<S�yo�"��|�x�A��R�a}��#�_����z?K�eVy��Y]�ج)D/�@���?�؞FUM�,�<:��l���#�!'
Y*7ߏ��AP^���<�c���?����r�Z5%݆�7\��"���<ɚ��j���"r�3K���&��톀"�o-]�E/��M�V�$�����px�/GV޳v$g��;�O�������շ����(�ےbۋ����:5��N��?	��&��B�O�,<؏�:ɄT2�I�����1LVne%����F����������qcM=��?1	��x��S��d8͔���-�#8h=xTI�q���<��G��7V�i��t8O��<nv�5������\6��UIqE@��O��ɬ�����.b(�8��f�E���,J
�b�{V,o$�ё���]����rاӉ(����ؼC+	��꿚�)��0u�B���R60$��uF%$�,��Fj� +�U���Rt����>%����m�D,�6�v�L9>�>�p�XD�Ϡ��`�ł����,����B_y��L|I!nG])=G�`~t7ؼG�c���&v}�LNB�˷�w��kl=��� gd �`�г~��Ҩ�0�0�I��mD}���M��2����zY[����C!��\+��M�AX���$-���~���t�W�g����蝁�zby?�>wd�c@9��h�@a�:s�fƤ�j8^>�f��%gdV�Nt��}A�O�s���[)�]#�;�r_eF{�D)���uda����+"_��$ P�=��u����'�ͼC<���9�]�*�&�>�c̤�1s�-KBi�^EE�
��>��0v Q�|�)#��&��Tl�H
�^�L��`�i���陴�fC��VBV-�/^�M�m�v�~a��Nn�[/7獘�!4�R�bj���P����0V��hEm�BB�\<�\^�����e�*o���e��a�xVv�Løe=+�4��v��m�ni���WyR�]t0M���6�$���aC�[�X[�y�.
�넡+�(	�Aq�g�X崻2�aKz�IC"�*��gQ�p�]m*"�)��g�d���	N{�\����au�(�j�: ��MbQu*���O���X�[����N�;rg�5x��v���}�_%+�Q���u�slC�idM�`iJB�>�H>O��a�dU,��k��J�ɇW͛C�"���K���ħ���:՚��M}�^�f�z-΂hW�\O��
,ce-?����b����}�ay��\L�C{;����y%K�ha0�1U��n*�aR'K�����)CZ:�u�M5ͫ�;�
����Gգ�ϐFC��w��q��	�.��g�f�C�%6�ZX��l#�Z�]���A~��vY#(�॥��*���I��Z{_�T�0z�("D�2��˟�U�&'�)�u�K�d;�@2?���]9�.��HZ]-��L���^ ��;�o>:�4I�)�Ho�w�胢�g����:&Ay{��m�h���7��b�)+*HpT�.Z+m���F��C�&�p���$�Y/<�ԁ�O��� �偲�1M�$P���B�{e�O������M��$�m��ų^M�af��y��!p¸fMNĠ��Њ�N+�
X�e�j�S֌a�W]G�L�VYv%�oA~�.?�9$O���?.ː&q�Ʉ�[�&�hR�2fה�G��w	��Wә��x_x�r	��U�LإK�ٯg��>z�0���M�^Y���X�5���/��)n��?2I)e/����c�[$�e�������Es3�狉&�O��.x���C:�䰷��o&�ĝފKn'n�XR���I��h/"%ˋ{���}�BU��`�Z��:< tIy}`����ƥ=R�G�';��z-������N����E�ֆ]�� �@����oMF�N���%е(�Q�O�p
�?s�E�@�.q1��a�d��F
;�GOYGr
 maa�*r��~0�Oٿ���;cjC���ӱ%�B��kl�|���������t��>�_3���0,�t����+��Y�GL����9��u8����b�\��R��ڽ����i����5�smk �D����	5����۷���YE�ƵV۲-��L�M?n��<�_��r�h.�k��5�������d�κv��[U��m���fĨ����&>E�	�ζA��'��P��y_�2q��t���8�y��T�K��4���vHC �� 1'V6�t�72�G����/��I�u��I���W^H:����l��`U.S���&�~!sܦ:}��l���xO2��([� ���ͮ�_n~�����s!�u�k{/������wJ;i��(SQ��#$��z�4l�ѷ�˲��^�<џf{N�h����u��ma)��]v^��Q�Ǫ�x"[S|(�[��6��.:vs��Y��Yk��DH��_�ǃ��ဂ��ڷ��=ͩ�_��8�մ���q�@0��qx�Ii|=O��3������o�$������j%��u��+�,�1�ߖ�75����>�ux��7:��!���F�OBS�]"��1%�;�Pt��28�ԅna�����d���+�#Q�#��M�ګL����$yQ�����l��v�4X�rp#�jo$����~�3���Ҭ��Dg��A�>��R�Z7��e��x�܎z�?�����H5�����2L�-���G ���2�3��l���?mR򙀌���/���u`D�V�!���{>ɇl�JyP+NO�rZ�"`D�?D�8�.�p���􇫅�a�QbL�EW����u{h�h
����>��t����hW��Uؘ�h�TХ;������`U ݿ�n�d� ����jA	:M�,�;��&��zA��������̱ ���Z-�in'{���Y���5��h��T�i��b��dN����tf	;Т���y]���S�N{n��r���wTS۫wu�s���#�'2�M���j��$���ߩ^��'G����"�pk����(|@f~�:֊�FrZ��V1;�$�p$M�u���Y�c���1!�������x���³A��$�cZ��a?�:N�
�m?){ B��k-Z�y�i�]��VU���>�=�K=|�M�4��ԟ/Q�J��*�5C�tX��Z�;����<A�� 8�)Tt��\)���7!	]/<��-��S���1��M�u2)Ƙ$�c��v��<�o��vy�XNn~.�\x5�0+2��l�:^i�)�.�����\	�E�c�=���iA@R�9[ ���w ��5@�^i�^7�p�p:ԥ#��3R��6��H�κ2����Q�ѽ?l[�؁Q�q�>u�ټ��n���w���6��yrd��*!�5G�q&gX��1�������&ěT��C�|�Ug�'ֆ4X�\#� ��`��*�������-�����C��S�t,#��&Eɯ@W�_W<�\��S�E�t�\��w"�:�0B��fQ�W�z� ��&J���Я|�<.I��t��]K�y<�^T�s��t��ۧ�"v�U%�2���
 ;�W�����M�Jlo�tgJ��b�?�Ō�I�Oa\�[�р术���XP��$��!	<2���>�[Q�A2Y̗j:�B�$�6#�<c��4�J`��H���D���ڋ���RA;n��C�[�y�6A y �wGe����-d�uSn�î'���JkgD��s_e9��{���I��^"�?����@|p#E�~�J�ǡ]<j��v�>�_Ӿ�m_>4c7!}|�>$f�бTJ�(��X}/����4��J���E"��q��-\����sć\TC5i�������'�9�9�چ��
����<ݰC��}��љ�Ӗ��]FnFbf��" �t9��L0p���]45�)}�$k1�]�$��rQ��'�Zâ/G�awA�c� �+���@�\}b���~Іǒ�\��K}���:dχf;$_��F�a�>S�О}�G�0�Cr:8̾۶y�L�8f���;�H+­˟����Ɠ��������?ٗV<�凔>_Z��w���xԊUa��]3�x'7P�#�ŗ!�m=�����N�$�]n{�˺ꇷ ��{�޵g�6�US(������GH�Yj*oo��|`�:N�w�P��q��-a`v�1���+[�ƀ�.�8�hX�G{���������J#�Fa�>�M>�9Or+��� ����q���`�Qpn4>��"v��H �0���m��D<�7�~���ޗ�7����s�·�)߳�yѤ�b�_N�E���uo@1��UE�.BO3�],	�NGڭ�
̎K�|.Ha��vЕ%șd��Gj�~�,D�`���5t9�슢ڼ,�2q�����`vK�*�.X���C�C$���AO��ܮ7޾W�+��ǳ�*~d��P���-��ThO��6�v5�M7d�qx ��V���h[���{.�\���=���f<�X�� ��Ĕi����aX���N	�f3z������]\;�@.��`�����d���b��!�	����ҵ�y.��x��8o�mR�����5�UT7ut_�P�xK�2~����w3�ZG�"A��F��ퟴ��ɢ�л0�����@�7���}���]�15q�WTa.t簧��	ӷ�u��1}�J�!@�=��P3��m� KY�p�f��)�9
9Ad�����!�/�uЍ�j�R;�ݒ��
�,��UQzo���/̖!Ʉ�h�k���`��/2���I�ۜ�Ҧ�N�d?gF$(be m�Ȑ#�W	���u��s>:2�^	8�?02��c(q�К�����:x�L\�ǆ��*�ZeI m-X�>�*UV Wi��Q����3o'�Yi�touu��ϗ���A�z\
>��� 0G��x������3�[���敼g�k��狭NglJ��s6�=�t���rU=�aaC~t���"o?��B��bٽ{^Q`2M�`�Szw��A�0m5��Fn�c�%<����z�A��j�W�$!S�ڋH�0��4��i_A�?\l�+��x�LWӴ���,�몄����;��zP�e  ��4�9<���Λ�ޥ��]�+o虼/�P\�,i6:��"����Rq���f�Ō�W B�R4�g�!����&� ^�>�8�(��b��0�|��~3���k�e����}�5:�CW��סChi0�L�آs=�O~�b/��\<��M�/��v�-9~��3��B���W�`[�t�f�vb�`I�>�$�uD����Z'%gM=,�v��jc"�u�T�����-�����D�9��������,=?7�K89VR��i��R�t��0u�A*y�XW�ISil^�cz<!�f�;�>[�}�7d������jjv�uX<r�A|W�eCl�����'�_��Qq�`�b�ar�8ۚ:?y8}Q.9l��FE�LP�3Y)����Y$gU?��d���Q>�,�.DF]ڳ�9�Nu��`A�9���O�O��<�z��{�ȳ�x�qro��M9-�C$Y!-��^��_��s�N���6AĬ��3&ި�Ar9����ÿ">� @���P�F� �C��oDN�4ОۍPZ��?�i����8>�\" �&���^��Y��!a��_5|��)��T� ���证��� ��Hy����:�-�� \���9���,u>�bP�Gh[������rc�P+����&�E�A[�OW���k������<6�战�S@�B�(]o�̷D�#���nRG�r�m�'T��?��:oU����[��*����@�͌����k��T]{�8�7���'�mD W���t������)l�8!�9Tq[Lo�G���i�6l]x���vΟ{9�U~U���.�!��{�Ur"�_�T;]�0m��
Y�&6j򠵶�o��:fƔx(I�LZ����"��%�
y��-��tՖ�v�6׉��p#�:Sl����b���'���2�~���\�f�Z���5�)�d��~jO��\l� \
�.�5+B�ڴh}�s���e#��:���S��O��#�$~^�H��"Xz)��9风�q #K�e.��N�]"���ay���3>O���ΐ/�.�R�Nm��W��JY�	��>/A��H'����4�UZ�����r������F�[:Lg�CG�'��l�ni+h�bc�`z��ϋrVS���4Yz����� ׷sG���۲�j�&d��H;�&X��H��y��c6�/�lu��)�4��5/t��.�Fl�61�}�����H>:TpE)��Qd:�$���#ะ_��M.�����2��u3�!-�>��^�W⮨+3~�����|��E�-�ش~��M��dk8��ZG����O��T�2�,��^��1�]tA���O��UexG�b*s�=_���" 4s��Z��Ez%w�̆����:A�/Y>�J�T���������r���'�ឧ���9+���됤��X�S(��q������	Ņ83�c,]L<
V����2iC�ѽ���|V�4z�u����ɘ+�w���N;�1�߂%Z>��r���n���Pml��Kڰa�����Z��k="��OԤ���P��/N�������t�X4�H{DXg@���b'/�j#}h�@Sm�]?嶃[ �r�}=��|�ux�,�xi$���C\�c/�[��7-�慳v'�W���/F�I�)��ѣ{��x�a��d�0�y
2�҄�����XyU3�E�����T��]Jl�Б=l����^i���Z��-��k��S�|h&����A���0�ᑖ�K�h<}��L�/c\��;W+4������CN!R���������O�/�g��e� \dj&L\x���p�U�ݎ��*���14؃�w�3볍�v�h�h�y��:F�	��4�z���60��(v1���L'�O7����PX����2�-�1>�w�0�&�4���_R�W����������x�ħ[ីE���z�Bn��ą�bSc��d�F$�u�4��'�1l�T�4e���Y��@�tV/5��1b@�.$o1���)^v�W��I�_����8���,E�ꭝ|�xI�����]�������7 >'Q�n"~�&ė҂�@Ib�!����\Y��S�V�h}m�����Z��Y���(�������|YRrR��!�)�⧸3�g�̜���W�b�?߁���BO�e��	+��ݪ;v�6�C�>�Wȿ��V����@�ɭ��iI4�U��fM�Mډ��f��h(��O�UVɶ������B^����j�k�ѕ��m
�rЖ�@���U��Uh�d����z�hi7*��� N��%�|g4��`����Yg���Fs�!�#H�M紐���Q@~P�WY���B���`j�C��R��ߦf�Q�D7���#����2��=<�a���t�\C����pN��.nJx���mr����dm�ܴ��B�I����dbԘ&��s�_y_��0�E�Wal:)j̀����N���d����\O:(���&$����=b��i�`�'1��4�M��*Ļ���ŠN�.�e:�o[��=褄�� �8�x���.��ͤ?���R����w|��ɢ����+6��2�櫘�yO+[v��OS�-�\4dz�mV�=`H�A!��u���!�ࣁe��[��{���WV�M���P�&����Wz�C�k�y�V+�y|SѢJ��E|8U�v��^j���ޣc>v^dgj�G������2y�cg�άI:nd�O�����:�Le��e���d��0"�E2f|��%�c->�4����7�!�P+�T"�ɝ�r�ꦤ�}�<S���� n��N��\��Q/�?�a�-�Q�E�+��w�/U=�޽>&���|
�����)3i�Z������	������F5���Z�gbx�,1�����(��!~k��'������p}`>�4`ѐ9��a&�2�FL=q��h#���kn]�u�� 6�Ħ$�=�iQcZ$�ll���C�O���Ӓ�oÄ�l-I�V��`Lގ�t�P�;���:��_w���}"����R+n��b;���,y����_N4��ʞ�H/�r�a?�˽a@{J������H}c"�41آc�4�k��o��9��T�	yBq"�� �x���6��%��$_���K&2��X�@�~���9�l���)[bY��T|�d��lbD]��x�R�oz���>���`�:מ�]Ne�-B��FZY�LC_���Vx���8��ʐ��*V�R�ݭE�Zw���Ŝ��b��S�c�i8з�B�o7�A�}����"�9�ɼ�1���6ǯ�8�v�1����©;U��vY�T������
*���{�5�q*z��ϐ�
���$����FM��E 
��_��Ac�Wf�g�2��{8}{���x5�=��}��mAtv�	�C�����`k��G�[:Y���7f�w��^|J�(ӕ��e]�]������3�Vo;�W�!�l��ِ�	�N�ˣ��HRe��I_�D(�Fs�+�����_s���$�����ч�V��Ý���v6�m�˦��*wp��ߵ��6��v9��au��A����s���|'^d� �^��m���}i���<pv�yL����I!Ea*��7��>ʥ'V��VDӟ#��۷�͗�h&f0J�yR���8/d'�C+�$ D���q�x�Q9��B!���c��M���I��kV�:��c@ՙ� ��G�U���a��&Ȧ��t��a��J�#�r��m��N�7b2pM������iE}V��1^�
uK�0z�����y�?�j-���35O�^���/�,,�@�w>��٫Q����]� �П�/~�;�u�����7��d͹ZݏO���*��l��X��%�9����w+�g�W����Ə>�����=mD����r赢��ecz�\���O���.#�(��դ��۵�Q*^B4���|:��!��wf���xΤ�P�{�4'����9���S^��<����uFP�I�6>A�$��p��8t%���a&'�7�T �U�$��+�foz�".b!�Dщ�dp��[<�Q.�d�
XǍ}a&��8�
8��^(�����%��Tǈ9Đ�F�f�~����5��8���e�PaF��3�*��!����o�
����s��m����")���r�'��3�y�>"{��ұ�͡��N�m��0�l�/,t�pK�(����LR���F�W�JO��~Â�Yܛ� � �E��zn�$	�W�D�s�,p�;��O�.�j����I�9�i�e�0E�qO[��E�S~�_%j��zh*l?#zV$�ë�"H+ �x���~�����t�RA*asxy%u�� �ć��@'�J�Lg�%m3w{0�����L�$�E�XM��Х�T(E{����%
���	�^�{���,�D��ɪ��.K��KeVبmWk��9�جxS�f���^��M��o�k��?� �����d�fjQs 5�>y6�A�����nݎ�nps���[
�ޘ:���G�a՗G�-��A�P��X������Q��t>���
�hΚ��N�&]O�!:gT��<߂3Ԟ.$���y|��s$^{3���v��dR���3-�p�u�)��R�`��c{�	�Q�����z��(�n�d�&��6��~�N�X�39�7�YgS�SN-��p�XeAL��u�3 G�J����m��ic��� 9ӧ��v�V�n�]����@Ґ��.�&���a?h�����)�H��N^�B$�vF�.�+XC.�+$w����&�k���y_L<%QF�O�G�[yY�ٔ|���kzvkZHȦ��*�}��8��Y4��