MZP      ��  �       @                                     � �	�!�L�!��This program must be run under Win32
$7                                                                                                                                        PE  L ^B*        � �� p        �o    �                         �    �        @                       � �   � 
           r    ��                            hq                                                    UPX0                             �  �UPX1     p     b                 @  �.rsrc       �     f              @  �                                                                                                                                                                                                                                                                                                                                                                           1.25 UPX!	hF^��b�?@ �_   �  & ط�� 
String�%ᐋ��2Ȍ���2� |xt2� �plh� �d`� �2\�X�2�TPLH2� D@<2� �840� �,($ �2 ��2Ȭ�2� ����톿S�ļ�
QT���D$,t2����\$��D[�c� ��<y2 ������s��mV�l�<�> u:hDj ��Bmȅ�u3�^d� 8������3ҋ���D�[��B��du�߿����+�� �@�W���J���>؅�H��P�V���m��0X	B�PP�����
�Q���G��WUQ��_�]�$i¿}�-�G�;�CO�S;uG�����m4�F�'�%�v&;�u��;�u����֋���4Z]_���@ s^�����2O��^�;�r�J8�kk�w^o���u��~)T�{��`?Dd�
�r΋�ߵ�n;��)s�&A�$+�d���|$J+Љ���4�l�m���S;�u�Y��/��ڋ��� }���n�)����	���sjh ��� V�|{�;��t#�Ӹ��G@c$����P&��cU�ٳ�o����C`jOhUR�ɑux$�`oN�; vۍ��k�L����7�� e�T$���h�m���N�Q�s���_��wF��v;w;;t4�=�m��v���`tV��
�E�}�Q߁�Xu����v�/u�|7���8׵FJyH+��Yl{������m#���� ����e6���9D;خ&C+�E�5ζ���c^~��v��;{��۹��vW����+�WS�|��	6���=���s�g�8+���%C��4��O�$�u�+A�8[���$s�;�s����@�&A�ݍ�t�7D��P�%w����?�� �y��3;δT`7�TR��@��vt�FHFt�!�>5	�u��gש�.P!�̹L���r�<$-�P,��1a�6[s�	����>�a�S;Tu�W���4�f�ߍ٨+�����sU�3���ȅ2u���X�l��k�n�M�Fa��4�f�J�k����
�H�R� ��6�8S(@N�IxQI6���"����;č��5��p�
;�s[��s+�D{�x��P��\M�ɾ��t�ó8����s���s��;�y���]�ր�Uq�d�2d�"[�
� {��= 1>
�n�d�`	�P���I|h�ˏ��Ix�=A/����K�3ɿ��@=������<`��0��m�l��ZYY���}��ʆ������-]�.���S%˄�iѳ 6y	��g+��� ���tr��G�Ƈ<�1���ĥH,��t�`��1�8]u��& 	�㤉��A�[�S;�lu	����Ul�H���8��Ml9y���[�b�̈��$�n�bx��.�����@�G�K���|�J��r6�p���u�+�xqh�ƍËʃ��ߢ��؋|�&����͋�,O| ����-�����Ѓ�����T���
u\j���;6|��*��}�
�I
 ���sG��3|t)�S0�߾c+V�3���������� E�r;s�7"�;p{	�$���Tc�3-��K�� f%YhW����g�c�1N�#�;c.���!
��r�@FL>�{ۭ��7+����+1ƨj���}jH
t��e���(��,�����ޑ�+�YpT�8ŷ}C��s
�]��7����楗բă/�IF6��8ƃ�4pM�7k�t�~��K��Lq9�q����\�[u�u���:�C�Z0�t�,><|8`�g{��2l�-�X�`�p ~@os�6���+;0Ǝ�p���t��tiҮ�pw����jf����N�l��4�|�#�C:R�;�s
�5
��)G9���+,��>��\<.t4y#�X���#l�o���[!\~��&�3�ԍ�2�dG75��t �$bp���RȮYQ��0��P(�_�����]��9�$�T�����u]�X��c𿁽�zZ��dvq�'u�Ǒk~{
��p+��-t��cC;�`f�@�*�YN���c�v[Lu#�)�}w}�8�ZbE �5z֐F'��	����Y�5�L�=�z��ԯ�;�֒�
�L�����X΋<� !LaM]�TJ� �������8
������e�A%�1!ۭ��%E���ިû,����%D�|ty^��j�æBO�uE`�)� |2 �Ձ��˞=�Vx9D�
�M�-7��`�R�Y`0��<�H�c�;pJ)S�{)�����T�2���������*�*]����Q�|���9���Ɇ�8�-*�J)������~v�}B	;��ȸ�����))`���E��9�h�f���>
���!��;"���V�[�0�@;�tu,��'DpUp��b��
~�o��$�}ۋ��t����7��)�>2�?�x�\
��܄#��1��k:�$������1]��f�؁�����������c}��^Z��B��;������{8�p�8�`�؍ft||�
P��)�펋���P�'�+�:�N����@3���}-���͆@�4;�=j���g-ovj7;|S�g	Y�fz'{�5O��c�޷%��Ư��+tm ɔ߰핡�Mw�~�-��;�}�r7��{�q��^����?��]�R��:��(�N�.U!�	���W��a�t	vRX:���!�s��!O�A�!����HƂ8�]��6d��k7�W�Cj;a=}���ˑ$�z;Ӊ}�ěr@7?
��vS�		ÃL�f���u�^b���t2{P�� XK�; Y9�#-ݰ/9�Q1���j1�����}��VZ��H�yy�Ϻ4�7����������cM��������������� ��WP+�߾�"S��Ɖׅ9�w����t/�x*������!X�-�t��G�m`p[)�����g��E�X  �E�k�<fE�K���1�f�U��i�����/��,��Q����نZv[-�$�
/o�DYXZ��ǈ������f�ј	�Ѫ_;i�p�F�B�
��17{;RW��֙1�)й*G���1ۉ��:0�C2���u��M�-C�G�(��.�� �)�~�c��}O�� h�D��GKu���5��Jc���-eP�s1�b�� �����F�� t�� -ti+tf$k,/?xtaXt\0�'�R?�OJ�����[�]4�;	w,9�w(�[�����)u���i|����Y1��2�F���~�x�[)�����'���뼿N1t�Har�e{�P SvwЀ�
���^�Y\��ËO����3�)���~uj$��Ў|t�u�L�ЈI����[���� ��	�P4Bhr��V�|hN���Ԟr�U0 l��X�/�P3��sm� �@2� �-\������f�pf%��V�f��?f�f�����[�OFTWARE\Borla����nd\Delphi\RTL FPUMaskValue� ��p��� ����_��Q���%v�a�>ޞ����8'aHw{PPRj���f{X��XO��vOPS��Sɿ���`A�9�t�u���AA�mKvC}�g3f��QI QY�#!g�ZX'R�g���L�:����dX��@���;a��8�!�o��Mtn%��3�}�e����'��	tb�s�k�}��9���t7,�o7v)��8&w (P���,�;`�� X���zd�g��
:v�5�q1�P<���to�HSt%[gxd�S�(�P-��@�R*H<(���[� l��o�_�G�Ku'�HS��U��N F�&��� ��A���/m5�/t�J�j�MB�j���T@��8����W70�@'Wf���LSnB�`�wZ߻=t�u�[-�[)�Y��R�g	̋H9Z�d$,��?�]�h��ù��+�H�����w��26��R�O#=�}����,�=�tW--/K����=HtN�`qj?r6�=��t0�R=�)t=-�."���$U-�/'=t&��߃���*��d���"���p���������������
��ܰ���Z���R���x�]���&�d�B�#t�ẗc����A\�;�S�Ctƅ�������ߑ�5w�!|�y��0� 6�ٙQp
C<l_��`X�
Zv�T�h��B��gsw1
"9�ud (6�op	�|t9u��oG�K��G	]�\��_cpsw��~��~K�D�#����m��5������v�4\=�]sfw_��8K�0�O��x]�;�~����C$�_;��c����$��t���CL��
��?S� ��8�u�ib��K7�#|��(d�(��Z_+D3�������P*��u�n�Mx�9��-Z�����w �7���}��֥��rA�@�w�{:��7�A�$�6ޢ{Q�?Lzݭ�bк|��u�����1(G�$�]��0��(����Fw3L2���������H��K9w��Ik�
�L5 ybt���Wv�Cp%�LB_@���;PtΘ,R=��u�SJ�t~Xj��fx�V����^�P[���ons Copyrigh�(��-�c) 1983�9 8 �aR�� �U�Ï�6>"��Ⱦ�h��� |J�I|����w�B�v�XK�É�$wK�)�{_`�(�Nu�k'�Q�$!A�7�D�� ��XH��ok�
�-;6�{���KC
~)��Q�~^����߾	�Z�P���f����$�t��3�W����n7j�Et	���OF�k3��;o�� ����@ًꜛ	�B�^�"�g�]-��},�_�/�U���{�n[~!ǋ�n����#3%��k�!�E�'87[�R����.b+1�!R:
t:5���J�t9�F�K&��B �Z)��.����#/-Rf;0 ݆�,�3���m9:;��ųO�
BI�W�7��nP�A��X��cvX_��@s��e?7|����u�y��V��bv��-w�$��NzVh�^�▻n���CaA�;�;�5�֧v�4:n"0W1/�Ӊ�PJ�F`ǳcO�b�؋K��bSإ�XH]O�E�"��p���P��?RP�AkR���[��A�J�Yƣ;���(�'��͵�bST鍪UI���JZX�$����ðm��9�Ə�j��ۮh�k���W��w�R�����&��9�uXJt�v�;�K�Ɔ������G
Z)~Y���"+8A8�u:oS���ځ�Z�[u8'q�#`���n�jZ0-����ԃ��<5��i�#Ya,aI��S���R+M��x�{X�[��D��V�-�X�4&J|9�})�@Z�v|�J���d) ���i��G[�B�7@y1/�O�W*w4h�Jx�F��h��ݕjw��cA�Z1 mɴ�����kݏd�i1�LH�VZܺ#�xu�J�	��_���X��p�0�
U��(�;��X1h��9�|��(�+%vt��{��o)ʞ��?�2oY��[K2�M�t�[<�� �I���k�'0��"�<$��+�u1����9�'۟L �\�X0t�S�`r�r��b�Uu>8���	���P�OaM�;�%��ddk�[(�a}H &h�+��[r � ��i �8���Cc�0� Z�׬X�d��e�=bJ��%� �G��&��S��K����|
��BM�-A'�UO z�mp��������7s�V��
�tF�R��tXtb�{��2:�lf��HX��6#	OX
��]'�!Z�c섳xNj%��Cma� ���n�R|U���.
\.�۱[�.�&��]�4��f����1�|B-F�
oy((�4�3no�I�+��n����u(������r#��XGukz�U��fV8��1���D@����'�h+3
�h�(I��3��G��և�ZX��u"ז^]�0��jKR
�cV(�|$uB]�+�3!'�	�B�~p��O��\�+f��F�j�C-hAgĠ��o*(*�W`��o�8S��}��,hፅ���:P��U�O��}/��*�8mܡ��8x\�%c�~�(�;Nt`��C�a�LZ�]*���+u��F{�`�\gc�8��&�0]��BX6����@�6{֧2�4@��w�6`G�s��gS��;ˈ�����@=a���MHƄ52\ U-=��@�6@�߶�`�ƅ_���C8b�kernel32.dllo�F�GetL�gPa�Nam��eA������� |�jH��E� Ķ#Hh?o ,h%Cv�t$�و�r+و��*���nc��JWx���$XD#f���+�&,�Tj��o�E���3��� ��g� 8�}��
� ,;,�=������Kt.�����;�u�	tmC<س���StjF��k��uFh��%� r� #��C��	�Software�����cales� lR�" �)C7�����e��9�,���&�S!8��
�~��Y	_8u���(Za�$p.r�f(.r-U@��l�,D-;8��}�" D�����;U�:Z�j��!i��l��w�A����P��&�G`	Q���s#\���h'���Pz(,�R�PR�p�@_���]���mt���ZsQ*f~�5S��HQ�k2h#>k0GY3�����쟫��HuÉ�4S�F*�j+�-�!GH#����.�/I���D�'�=�F8p�'@ۑ|_�(��$�x�4� ��~H��/m]�i�QRCFHP7Ŷ|�����~�+����y��m�߭'�6#(@!�-�9{r�s�PXc�E��[�W`��>몖)R @ZHP�|��6�L����(-Z@��+�I%
gE	P)h���"Ŝ�����.b�o��0t;�:��^�6W�u��B;[�3��'{8�i6���ލ������fx[��˶uN�	 $iH/�����@t�z�	���H�(���J�uRPY<�v�����g=B&��$ �S�b�k�)�4w�n�S��S$���h+sU8t�>G�����x$u�;S���sP� �����o�U0�Z<��J�7h��3;Ҋ��M�2B+���f�h���1y��1�@e�=�t���P�XKr����o�@2:X�RB>��f�Z�
�R	%
b��7����{�H��Z��&`+�SI|��h��B�<4�N�ˀ7�vJ+Y+��X�u,��6��`�������h�̝�t���}<bw��.u�
��Kn�@�b��ڋVzey��
)���_�Ɖ^�V�h��f���du�n뾺����c���F.����xx�+D�?�[�����^3YX������=KX���u�P��X|H��E:t� v�7/���F�`3@~!����@W�@%V�u�>-����,ՠ@kv3�`��꽣'�+�~��4�љZ��[}�^�]��S���7��H}	�g�ƈ�A�'Z��a�����ɁB���Ɠ��T+vQ�y�kZ�Z��K�,����ߢ�����IZ+іa)�C��6�h�X��jo�m��$2�6d$��`���� D;�"U�3����2���1�~[�\Xy
���5�v������ۃ��\����� 9���o���������;�rw;�r+��@��[�k���|E>D�;q�����[,A�#ɃRu�6��C�Lun���WH�^�i�#�_3d���/+�uX��C �z�Ȕ4]YB�/�u��@H7����~�#�4�3/v8 �ʏ��� |@|">��nF�����������V"�����#�4v;��7����b�^o�6fbE��u7`W�
7�3	�I�l���	�B�܃6mM<9`�]g7X�-�D'����i �_tr(,�2����34f�k���� ����حC��'�	Fpƚ��آ�G}�����,�캺�d�/n��}O���	H.9`�-d�7_ {�� ��A�������{�ʺ�_ACv�a
��^B�먿hj@M����7t�S�0����<��s�:��ӸӼ����z�,���(4���4��d�L���� �J-W��2-�=��h�NT�+�č*Hq���
�S��Z����,�A�1��<�
7l�w)��R}�`�B�*8� c8 �1��3��8��a@�p8��m/R��[l�����d�A���� O��XT �2PLH�2�D@<82� 40,2� �($ � � �2�2�plh2� d`�2� ����� ���� �2����2Ȱ���2� ���2� ����� �����b2|x.M�4�]c��4 $S�q9�����B��K;���;v��L�C�M�5:�U��UG��ʭe;t�	�+�@���t�^&�_	(;E�r�`B|� W0+�س��O��R�v t�!���ao)y�)���#��E��}���m��������2���U�.ar
2�}�z{�m� ���ۿ=� �":E��E�	�Yog�l�.9��o!��E��� ~Z�vY����H�;!] ��@#H+4@5�����E���U���-��RM|;���J|U�T'�M�u׃�X��*�,�����sA����"���=ԃL�= ��G�$ZP�hVz�F�6{ք^��Q p>0y?.����!͘c���!�!��v�i3�!��\�OXn��<j��j��8v�Ye�q�gl�ݺ$P�)d<�\#\�~�ܹ;���3� �<�t��� ���%� ��2�3����r� ���2����̃l�\�@@$���
 ?58��NQ���@� ��WinINetз���nOpen��;Inter
C�~f"UrlA#2���nadFile	�lK9RGoseH�-s��%['C�ݒlooki��3ȑOGni c���ize�S�5^ml�E��BlU,�;���0$͍��������A�l���W��2��%��}(�L���z��b�`8�
�;O���+��9>%�%mnb=(� �m�T��%�i��`��߯���tyh ���toh)���j�[)�L�/�{w��v-�Ƅ#*�x�t��!���n�0i�b��~c�>u�Wȋ��E�A�TV�p#�� @N��1.0��B3%d�B�@�7=��@��D�u��@�|�@�@���@�����@��� r@C�9�)9C$�U)9��\�9����9�)9���)9��̐9����ȔD�D5��K� <�� 4Y�?��IVXLCDMTC�6�+�0��b{�O������@�_x�$LO�@j�� _2�
����� ӡea2���eO&�D�!��GD8 /���R����~dZ��Y�9�9��Q~��R�;T���/�: v�^n��4"u����&���C�=K�EN0;%��a��[��h w�\�G䜐#`��F��T��u(���V�9+�j�&|N ��F�P8d{��
�`�E��Qt�n|�:t�;u�
�Q_h6�U��3+M��'$}�K@|B�8�����|�"V���ȃ��P�0�F���+���(@����m�Fm�����a����� 8�tڄ��������:\ |�!����Z��BX��sB��0h �Z�f�C8����PȔ%;�ޡ��t?:�v6jE�LN/����|�*U�4��]N9��jaMTO�m6���@C]2zo�B	�᪫aHT�^lY���_���U�a���Dh���~�UHHY�/�u)7aϟ�>��h���?<6��� j�
`#F�ʶ%&UF����q�G-$�@F`�zD�T!���K	�� )��Y3g$�����T���!	K��"��ړݙ}`E�FC9h���o�L	�% �?g�T��_yH���@���u-�dd���.��e�m��X�3�S���sԧ];��JHm�k���@���g,�ܿf�8'�3\�x%���6@8"f�DB��O��;B�	)�� �L�<
<��a���x��Tn@0�y^�~ ������DP����@���0�`tH[}D�{�!�i+m�9�O@N�+�"��h�5���z��E���gyi���63R
i�`���F���Eݶvo�9��`���L��[����/���ˤL+��LkG�6�n=D�E"N�H�����	�LraU�b3�愸�8994723#�l�088193913;Þl-#0H�)s"# ,dݻk4�����M�uT�l��=x] �|%T�4���'M�i�А������'���0#��N\h��߰�F��t�/P�r	����N�N�Y� =�dٍ�p�$E���6#:47&{��Nc�%�.	-��R��_3\�� �gram Fi�7��'aded Pro#\Do��wnl�N��с����2`O7OC7�/�>Nr,�Iu�Q�R����kZNV�I A�DM`�̈�\npR�R��������6J!��\�?���&�rSS�4|.{X��t8�S 2��4H���s�xq�STl�d9�|���|��8�K.���q�d9��@����yF.�����K&���v ����T �8�s���Td9�(qؔ���T4LԌ\2���\L �tМ�<#�̄���̠�tYF��OxF�=�ed�4�+YF��"��I`d�kFv���R����� )}K���#i���ܜ+SApRA��I#umEn���K�lA+sEna��nnec�+&{m�a,CC��R޵�[y�pert�P��c4fa�`'DialPa�_%���(7S-2���2A+B���kngUpJ��7�xHa��Statu�5��l�k�]��]���Devic�ؒ�'Ae��x@y��VHH�>d'��,Y'�t��o��OA��e۫ˢSb�'2:�&���;�k8�8m+��9�r0�
�����Ur$�V�*�	9Y���&�����:~�5����]@���|jt{[;Eu;M��8[R7 ��>�Ȳ,�%�M�������ȰVKHw [�����j�Z��b�i��y�u�3`��A�A����Y��l��АA��x����n�f����-� B�VR� ��<a� :cr���:X�=A.P���j��\�}]S�$չ�#8R�q�+� ߉�ɢ�X�8�x�X�U�+�=���	�;��e�e��8�T�V<T�撚�![6,4�1�-�Ĵ�l�����@��Y���Ud�Y`$�Xȼ� �5,y�����A�Y��KH����d�A���)�K��C^;X���
�6�g�%����,�[� ����Fܠ����OՀ�֮8Ctp:///`@.�ht�|*��u�C3s4����'Z�|�H!ZgZD³��
Pd�F��������B'p�츀)��G8�`fS��rI�
����uCM��bAKRH�l\�H�Z2!�3J^����G�%Td�I�NCKWFAW�o�sep�tout�ٌ��s�owb�~Curre�VsnY\Ru�k�A�M<s�%,U\fd��cՑ�[��[9%D��[�\Hp��\�4��l�'$D��R�It����R�G<�`��{I���J��T�^1Q�H���hU��ÆÜQ��䀥[ۈ> γ��X���(�d�32`\�SuO��]Q�h����	�� d�=��Y担x��t.�dd`l`\֐KFp\�������.|���T�`�����jC]X3���|�&����OS=+.׭������M�SJ�&'�U�^��c+v�r�P���o�J_nx���� !� ���X,�ʚ;�Yl9�U	���>��_8�`�g�6��_l���󵏐�x��|�<۬��/���y�d�_�>�.\m/_������\X_��XN�0��Vx���R`rʭ[@,�;�-�` �!#\�ʃt#F��^�к	�`�ekModem��$<LAN�S�N���`[�,�T�k.h�Rn+.2�� th.phps���?�e=1.8o��&R=D7S�&9MP
Tipo����ln=	Univoco('_����(=7IEA��S�$SiC��[�=�ɿ�
�\T�s�'��amp�W�apd���C��*�$$�8ub�^�a0<�����a$�hUO�,�`����Kh�	H�]x�E��8}��ٝ<T&Z��M�]+*�qh e�0a}`0`��,�ﲗ|t�AT �M�MD/U��E'߈�,
r
,r���B'���0���A��W�I�ݰ�0��'�$��d�Jg���*�2=<1�G/u�V�ࡸ/�D���R��D�>�3� ϳ��xaT؈ݠ׬I������[�uøR+1d��څ<��*8��ټh2��yy�<�A&����A&�����A&�����A&�����A&�����A&�����H������F�`+�4B@9���I��.Ћ/-d���M�uJ.�H��;}�g�0$u��l��7~҆��AR��
9, I �d'��IJȤ�d�"��G
���Fla\�0z^$'G�e��e�ɮ��f�,u>�fs�R�)��f,<@���P?�H�G\�@�uz��V�pzD�2Xw���8#��g:�U��$�x�D���n�	y8�Hw e�9��%Ǉ��Jj ۇ�9��h
\^�5�x$tp��Y�h�h�h��2��$�(� ��8���FV��,��5���ٽ�h0i8i1��i$�D�y��:80<�h!4�<��+2Xhx��MI4k8h"��<�2n;��e<��<�e�y�;�����c@ihX)`%3�G2Snapsholp6z��3�Tooqe�Ԙ��C������'irssscFjE�u�!���2Next`���4C�
E�6n$���^�#�I��䓓PSAPM�7`mt_���A;ul*��d�^��;����xSe(ܲ�EKxZ�7�J�9r�������y�f����k;��8�	0�(��*�婅�P�Wu2(s	Cq�2osMp�sUHN�,�wG�c�+
�D��(���kԣ�dۍ]h TD��gQ�䒑	���#;B.�0b��0-�p��kB|铊���� j���^����ly���ۃ7^��9�8CWс���,HO*Af��*�� e�2d�0�F�,5�3�x�x:�+O���-�;G���@WfK�Ϩ��-�����W��B�/�FJ1�[���[~=��l�b=a��;g��l�@Ht�i��gclkH ?$C{�newd>�Po pay~ �MtIE43�B�C�1.e��^[_iޗ�eme/2=�7���&�89n�����|�!���	�����lhO��Dv92��0������u��na��ˈ�K�+X��c�]���� �I�o�A�rE�X4��?\�1 �Aݠ�9�1���܂��C[�&��h�3R�\#�#�%{8�q��{�9�M�D�1�_=��a�ˈ$Ez9�lbF��5�,c�7��e�Y��o�К���S�[�h������h�pj^��)p0pP�|g�+&����p�`	��p���P��n^���KhY6�����0��p"s�3!uQ�Ua-!��o\Y'�3�XRq��@�T�|Y���3_�w����̏qd,��:�v>Kպs� -׸�J���-��mitX�h`�[��xv��Á�qE�P�])�q_�E�SFr��$#��<�@M��w�6�������E��$��U�j�B�w�	��w0h�<فV���<.�r�PdP�|p�v�W��7]���VT��}���bc�B0��Id�Ć��4���ˤ7�������O�@��P����CI8,����/s�[��	�O�Y�;�I�e��,- Ɓ,ȸ���ȼ���r ��Ý�a��f+	6�m�ۃ���8@�
�8�������#Y�
��跱z�d8�]�r ����Lr ��p Ȝ����F�7�|��Y���a���IB���9���A� |f�-�� ��GH�ȁ ��.�aS �-�@.�٢�"��@����@�!���/5�쀀G�����
*%��q�f�7���|�2١f�tle�[Ht���X����5�L�6��!1�#w=��逶�@�H��#F�-�d3�7G�QNw�J�(� u?U�0�l��Ē��x��_� �&k����00d@�123@d@45d@d678�K91w1�11��111�111�22��222�222�22��333�333�33��334�444�44��444�455�55��555�555��t��|�jtO���:�pËxwG>S0xjh^fg<�P8��3c.�,i{{��5�u�｣@"pj0O�m�\w� accede��w�ll'Ca risvata!�R&⬧AyF��|n�+ݠ�t	���I�ѻs\z��l���J �r�W7�	@��V pH5�����|�|���s<��P4f���� �QI|uLe& WS��#K�K�?"����or.e)G�ItKpl��M� D`��G�"�H�"|���9�|j�0P�����	\�.L��0�=�`PР�)zd�hd��y,)p��~߉�oXdh^|A�h�0�!N6���9�Wc!l)rY�W�=�+�b��
Ĝq*8�)hq��9@ �|/)8�HXo�MIp3���H�9�t!tqm�f��#c��~��%S .���P�P���h��`_,�]�
={����1.�H��d_�	���"u���(0�a<0�	��HizY��CNE��XF�. �IK� quCl�c�3�V
�� |�t�	�}�!��h/0⠊�K8�"@�)�Tm�)C��ܱg��+
�+.ދ�h��|�����hȀ\H�]���%��<�c�DG6��H���$#_̓Ǘ��lN�TJ.�܃��F]v`��'��H.��$�4�=[H�(5@L��.%5�16, �666Xh�"��r �6t�<�¨*݄�&؁�9@��y䤴�<�d�D� ����g�\H���9���L�l>�؅��$3�@�P`<���0<L5��� lВA�gXhx�<3� 8��d��l����ˆ$�Ƞl�d���$I��<{���lS�R� ��N�è�drcA�B&�tGeɗ�Z�OSle��=rcp�lst�r@at���DE��Y[1dX�U˷h���H3�]v�M��AS!թ%S��&�S�Mov��U#�lSC��%'shyAS
��7ec+!Ѭ߷r�'kpu�sageBo�U���,�|Tr�-�#4#�DC�۔�W��YbT�w��@�e3��I�>��jPY����Μ!@c8_���Q�ɓj 	�_��Z1�d\W)�i;$�
����t�4�U|'���mOtE�A<�#�ܰ�!��J���py��ě� {%�mzY��'�	�>G�F��҇f�ܺN��h�YSTEMF|����t_l\
���nla�\{4D36E96D-E ����5-11CE-BFC1-08002BE10318}\X��,DVvD.&)�!c�UhHK��InitBak��LM��������䱫�dB����I�ֈ���v8��PL��&yX��"�p��dx�h�2n���<�
B�o܅T�����oT4\�I��#��y�E���"�vFz��Q�����|�,t{��� u]M��;4@t$ Ga�ĭ�ğUua�0���)#qBץ�`�4���se$�l6r���x��{H����T���v��f����f.d9y��ք�Ȅ�<�LǶ�c��B(ch��T�2S=f�քY���L�rՀ]��>4�j������W;0�C�.,o�V�[�&�͸/$���,�ui�ODN��C&�SDNO��RrH����F"CSfd�Z�AC���8�ٍ'��ުPeIʜ�*���;E�vaM�I����v��'�EV�G��l���s0���X�8�S����� tQ!܃���vF��L8��0�5��Rԭ����$��r,b[?I�#��0Q��l�m��	k��z���xP�|gIr*P���T6��7#��dS� ��e��u� �d�s�
,�ڳJ,^(0C��4�ɔl���xx$Ms2���x �rC�<����jkU�g������v�eU������u΃=�-;�s�>�{�xy���3��ŭ��IBo�́0#����\��ј��z0G�L2ȣ8^� ��$'�d�8^dd��9],��]�b�0�F(!�.y.�(�Z�����Ɛ=���{�s %�T=�ɂ!��L�����[��*Ȑ����-W8�x�ɑ�'���5��n�	���)�-'��-E��V��(�ж��W��6!p�����뺅��\�#��d��t��V9l�����vp9	���6����5y!������N��������v��9F�g�\�!0���#����sQɑ��mp�p����B��Te�M��)&�=D���%�0 �#^'p8�32lG/��V��#�G̦���r�p�pi��I���p�Dl!B�Nϓe�~��l�샷�>ݮTe�Dl%k0g�حW<Έ��h�A�,�%��u��a�s�&� \����\%�g��R�p�*�xK�����d��;� f�|":b�0�� K&c���ѓLr�����+������`Ų�	XS,`��\<$&�8�H)�w�l
��^�}]�euf ����|/gF� �gE��cj�-�nR�<�
��$̎��}pd󐯖D�Tw6.�����b;f�ƄlZCl<�`-FMClt6\#�>���ũ`I,8wB�m�iF�4W�$���
$#�M���[�cHC��Rp�\XtM�,꩏X<�5Ay���\�g�A��`�Ը���d�}�P5W� �}A΢m	&�,߷�$0�<�H b@�Hg�mҽ�.��پVwM��`΂�S��x,(�0d�9�����9�U�Q�J���B�������˕L.(1.1)(3�e/) (Y���0)�w�\2E-�ktoH�Z%	�Dț��Ȋ�ɘh�h��D�h�h'�ɘh�h�h�HN$�h�h�BN��h�h
�!�h@��0(!���	�	�c�M��KL�!�j{��kA)�[ �]/��ϝ����-9��ȓ0����c <���p�ݐ����K�2����`c�����Xb(e��Q$g�!�b䇘��4��B|��a �@��!_l���	�7�A6φ��T�|bA��8P�@�2(�q�*G0�` \ }dvK���O���jf�.traff[]��gtob�n��`w!?D=;/Ac �_NySQL.IVRMw��
C=���Bw/R�cW�	ecugF��a �� F6�gold��0�cj2 �M�9$c#�x�rHv�f�@]�ȭs�Sj��N���(�.G0�Ф �0{CHNн��h�z����9@P �%��%�l� �\���"�Ul<]{�fv5��b��� 07�D����������� p/� ��W�n���-�蹆�ؑ�(�f�P��h	4#r���l�����էd����]'�uŐTz\tG�`F����`to`��K��t
�k�˶p�$����d5����5�Ao�a�� �7��e|`�M��J�P"����\��f�r	Kh߁��a	n���?��䬬V�r�tY���ٰ
�X ��� l�ʆ����P����������Ҥ��� 5���d��`���{u�(h$�2�	����=9��t8��pQ|!���%rĪ�����D���Q���\� yf���;a<�@F�H���B:u���P-�3�O� �!bKN�r�t!������=��3[�t\:ӄ"Z˥L�f��S�����"2��耉��&,vɲ��L�ʐ q��DL"���� xo CE��? m con�gur���� � sistema.���S!%s�o m��a.`�i~_��(Z��>��l709dia��p�fBUW��|#� �rm+�in�,���j3�t�?�0��oCs;��jw ai�1nu�IN�˥�`������P�2ֈ�H��cM@^�Ѧd��@�osVt�}T�6�;�T@K�� �#�P��wz�,BU�n��i{���AvQ|g�\�b���X��I����<am��7��6��͈��`OT ��=�HTR`lvك�T~:Ժ��6y��P_�������4(d;ّ�/n
1�1L$G.��L\�mxp�
1��`��%3 DS%4��p֌�JfUx9d{�����H��^�����lG$`u� D�I{��@��9�Sq&�y3<A6�C����dѱ<�D�R��cP�;{%Z{^���#8�8̖�uSMa�uU��^�'0LI�f�����!00�
9B,,�H�d44� ݒ] 
j���P��V Y޺�����$ i�����?s\c\� ���\sy�32\d.9�py/vnͷ�
�mX�sn.9V�/m+.��?#[	o.searc ��~+�a7SI�r�ONVET�sB�#N���]�JX�)��~�<AÍ劒���_@�y�10G�R���m�,~&�,�e��Jc	قY"A"� ��t;��d 9K'��#�T%�����2���[=, �U
J�a!��ߊ��hH"j_	��e��S���A����9��.�(c�u',���T�.σ}�L	T]���F4YM�xK^�Y�" �`�p�u�r�� �,��~<�zg�D�\�vnXغ�_9��@9TCM�V6�AԺ���\�sRH���k0$&P�p�	AŬdY���^��`�uH��w�@;;4� h5P(޹����9X���.�Oo�#���=2]�~0�P|C+7PPDAT-���);��a�Ex\QF��uk Launch��Ɛ�Y���O^EB���찓#'����HPd�H�����P7��ړ�S�A8�1���>S�8{b�َD��h�c4�t^9t�h�/��"��-!߳QI�s������IyЖ9�k�����A�Q�Ar���ɔ����Ar��������yf�<U�G&)�S���RN.�,���BAK&�(ˁ`����.� �x� �A8L���f��X�v�[���8,%�d�������f!H�x�-���U���Jt� "+5yXl A���f=����X�b�J�)������
&�M��Z�.���U�&�'y������9@��K�C���X)9����ɨ���-	��7����O�� �<����2�`g����� �����,sR��A��j�/��T�[�����һ;�v[��Grp v(ap
�@2�oups+���C��\.lnka�@w��>ll FcU@*p;C5fnCG�J��r=M�?��ݾFavDit)�D	�K��Q�-U ��>,� Di�ns��T	�a�O����g -AӘD$\��±�� f�\lR�6�p�� A�|(,���� ����f�c,.��Q?-@��X ِ� }��wA�$�l���4M������,��������
�E>�B[��;�wK�06<ƚ�iBHNT_"22�Ee�h22GCNF)����r���]�}	j�$�rX@"���0��/p�<gD<�����b@��Og��g��<�����%|�l�y(h~
����HU����
�ʜ���d��쌂�Q͇�Tt&���/��ɻ$�0��*{	�Ԗ,@��X�g�;��<`H��<#�����rAɑ2̐F�̉¢���G��H-���\�$�S�e-�n`gs��٩�� %g���@�K�g觜V�r A�U��֮&\P�Pla�� �form��΍�\@Og/�9{`�r �"�0�{s��y@7 �	KVW�5vH��0��C fģK R�,e��z T��_ ����u�� -!�����2 6	�sI0aD����&�ITo�SS���Z#d8�˭�4�6p; :�\.��=$<�BA�i��H�P�Msi����CР�uM�4h`0(�\�n�[DC�@Lt�u��M�WNcN��k�gO�/xwK�]�u������������ �4ߓ'<푼\rl����[`w��&�����+�I*�0�Nj�ݧD�=�¹9B������}����R��}%���1TǖUp:`����v$��=VEJ�⣍xZ0
�P��H��˲������
G}���w�BFm� ��R�;LOH�G�����]�l
RQ�n�ni,�P"��
 �ũ2�r�d�##�����2�t�Va#� ���m��z � 0  E����0123456789ABCDEF  ��ܡ
�  ؄M�	�� D�G  Mw�L���CH�������4��M�����@J7<���} ���`�tF�l���4M�\m  0@y%M�P`px$�i��0<HT`��i�lx����i��i������4����y M�4M,8DP\h4M�4t�����4MӰ����i.M��z��i�(4@LXdi��ip|����i��������B����_
���GHIJKLMNO��[�]UVWXYZabcdefghijk�oT�lmnopqyuvwxyz�i�g/+/E���|�i����T��ו0c�VD�4]l4���i6C�Px�"��,t�	� B�2 �v�(��Z�Լ��e� �AQ D V C L A��� PKGj�-�I N>O۞ۨ�MC!�¢N��WE!#x]#���C��i��@&���%PgT6BUp�_�fb KO3CommDlg�Sf;��7	�GDK8&D+���ΰ
(ShlObj@sAv;�K?veXDrl
���*�API
�RegS����?FPe�U#r��Mon�RichEddsDM���_7_sv9kAUYoX4_Vm9w�ߚ�H8d�Uhls_XuR7fdu6����#J6_BYh6tS2Qq3 A5�_pSw7gSS^��7��_xVTMsE57#2_WnBygqT���CB1_DxDO588F�5QX�_BkuYQ'���U�(�l�9���\P�	cmpi
N*�{at	TeP�$�<Lr�B�Library=4gDir�a[go���`�Ex>T=S�JAsf	���WAddr[��1�ul�AX��4x�W ��C_,�vLa\�Ef���nv�ymT��=�iabH�W��۾nFre�����To�o�UĲ�}���*fe��[7ipWeK��^l�P�z��Tl�Ţ �G��KnA)=7T���gPQTh�dIdDe��Zk'����@uWS�e�W�vEQ=��i$�P~�VirtuO�������6X$Q�{?dZ[(lTh.eM�R֒�%�t.
v��py
A	�H�v��{*���up�foAeT�2�E�h}���F�OA*4ĘxxX�{�IeWesUnh��[d ps��s�j="PoD����E)Of7Rtl:w_���
aikH�f��d�f!��&S�d�$� yp��Ns����e�!��P5�aFKeyj�3" l�,fq1�{��0����ى�yg�&�6�`�ȱ�l��L`j���_Z�R��q32��ck&z6l6��So _7dBru'�5ޣ�]#�ҋAQGdb�f[(������m�e�Og�b�YSL6�fk�a�Dqg��:^iv'x�S�=g�lzm��&�l�ux��T���{�˫�	(���i�YsoR�8�{ܥGDC
f�LU��elX��V|NRW�Box��sL�4�Kb��I˶ba�gn|В1K��! -�csXl�f���:�~B�U��^spy%o����\oy!6�X�f
4���cHHj��#x��p
���^b�rdB�����N^
 ��,	!h�HwOFv�_��DA4��O<

����
!����@O �3			"Y�l	E	����93**		<�/�* $2$Z�\�k<1Qrh�(����:Z#!�4�E?Q����:44 C-	2	5(N(�T"1�ۻ��+K4k�J���"
�����[������KC�K@	q�)�;O�g��2�v�
 
�wk������vmOH1����#	k+ A��v�?+�' %m����?M&*X�2!�.J��� Tv+���8$h)���v{��!�Pp/oom ��$� �7n��S4)]*XI�g��1�e#B:�	KFČF��� A^*�Hw���-7%�E0�·��0�B3(4�.,�l�&3�|���YJ�(URK[��!8c3�#�@9��Q$�m��
E�8>#B=\6]95c,#�2Y&=,,��ȶ5J:f3���� R��>�e��߽G8-=a^���-�� �L����;�"m�. /57s�W���&�D���	[�_$d)&d���l�	$ғ%�!s���WYKH�g7QBW>y4��-H:5qNX3�����a'KA7�Gb)���}��p�� nk���O�� $
��ۻ" .�3'��[�8`�N;+B ��
��0H.�J���5(%�~7������ݶ8 �I+%�e�o�� @e����f%�C#$("~�!`)$z�;��n�{7i<�+\�q/!QO����oc'�(&�-m ���D��'̹Y:�-5���a_0�! �超yv?8	��y��-�L |�Md�`<�� P�L� �_��^B*�w���={�\,$����Q�	�=l�<@��w�4@3	h��e �7j0(Ю,� L�+,���6�
CODEо����}�z4/��� ��#{���'��BSSv������.<s�5*�� �����O.tlsN�le�Or�+i�'@P�	Xe�K '�{�4�sr&������'��  >r�74> 	   �          `�  ��  ��W�����������F�G�u�����r�   �u�������s�u	�����s�1Ƀ�r���F���tt���u�������u������u A�u�������s�u	�����s���� ������/���v�B�GIu��c������������w���L���^����  �G,�<w��?u��_f������)�����������ٍ� 0 �	�t<�_��0z �P�����z ��G�t܉�WH�U���z 	�t��������z ���^�1��G	�t"<�wË����������$��f�����a�[��   �q �q ��                                                                                                                                                 �K�6          (  �
   h  �   �  �    �K�6          @  �    �K�6         X   T� �              �K�6        ��  �& ��  �    �K�6           �   �9                �K�6           �   : 8              �K�6       > ��  �    �K�6            �             D V C L A L  P A C K A G E I N F O  M A I N I C O N P1 (       @                             ��� ��� ��� ��� ��� ��� �� �� �� �� �� �� �� �� �� ��v �� ��w ��i �� ��h �ۊ �Օ �Ϊ �֔ ��~ �ڀ ��_ ��x �ҁ ��i �̅ �ʏ ��[ ��X ��v ��s ��x ��e ��k ��u �� ��Z �Â ��Q ��M ��P ��i ��b ��T ��L ��M ��H ̳� ��` ָ} ��W ܷ{ շ} �d ��S ��M ��` ڶu ��@ ��R ޷h �^ ֱt ϰx ��A Ǫ� �P     ��@ �_ ��: հm ߱f ��> ��: ��: ��> ٨u �R ݳZ ��: �E �W ��H ��� ��8 �< ��9 ��H ��9 �= �> ��A ��s ��A ��3 �M �4 �3 ѥ` šk ��B ��9 �/ ��5 ��= �3 ��C �K �1 ��g ��; ��q �. ƙi �F �D ܨB գM �6 �/ ��> �2 �5 �3 ̣L Ɯ[ �9 �7 ��' ��& ߠG ��s ��= �, �< ��` �4 ߨ4 ��$ �+ �1 �/ �7 �: Ǔ^ �8 �+ �9 �* �3 �3 �0 ʚG ڟ7 �, �4 ߘA �$ �< ܛ: �/ �5 ߝ2 �2 �( ��? �* �( �- ޞ( �4 �* �2 �5 ͏J �- �( �/ �+ �- ǑA �1 �/ �6 �- �& �* �0 �' ݖ' ��& ��3 Ћ8 ے& ה# ܐ( ސ# ��T Ӌ. ��- Ή0 ܇. Ĉ3 ��= ǃ8 ֈ( ׆* ԉ% ψ( ��3 Ԃ1 Ċ& �~A ц# �8 �{? �{? �}3 �,     �z% �t4 �x% �r4 �p5 �i= �q �o! �j" �g �h" �f& �c �_+ �\4 �\3 jTD xX6 nT: xR/ oQ4 iP2 eN4 bL6 iK2 uP" `I3 aE+ X@0 IIII�����IIIIIIIIIIIIIIIIIIIIIIIIII���ǵ���IIIIIIIIIIIIIIIIIIIIIII���IIIISx�IIIIIIIIIIIIIIIIIIIIII��IIIIII����������IIIIIIIIIIIII���IIII���Ӭ�yfXKN���IIIIIIIIIII���II���ƥ�dYA0$D��IIIIIIIII���I�۴�������oY8't�IIIIIIII����ݖu����������oY0	:�IIIIIII�e��u�������������b8	E�IIIIIIr[��}������������ª�oA��IIIIIIe[n}��������III��ª�oA�IIIIIIaVl��������IIIII�м��u8j�IIIIINR]�������IIIIIII������i��IIIIII`Vs������IIIIIIIIIIIIIIIIIIIIIIIBR_~����������������������IIIIIIIWJg����������������ƾ�zC�IIIIIIII=Jg������������������^6�IIIII7II>3Fg~����������������kT�IIIIIB(II<.Fg���������϶�����k��IIIII (III1,@p�IIIIIII޹�����k�IIIIII%II11,O��IIIII�Ĳ�����k�IIIIIII(II1*-���III�׷�����u��IIIIIII#II1*3�����ɫ�����}d�IIIIIIIII  II&&.\����������o��IIIIIIIIII  I"4Qmw�����l��IIIIIIIIIIII  
"4Lhmws__��III|IIIIIIIIII  -@PPR`��IIII|5IIIIIIIIIII   
!22=�c�IIIII|GIIIIIIIIIIIIII     +H/��IIIIII|vIIIIIIIIIIIIIIIIIIIII?;)��III�|ZIIIIIIIIIIIIIIIIIIIIIIIMUU���{�IIIIIIIIIIIIIIIIIIIIIIIIIII??9?IIII������Ǐ������ ��  ��  �  ?�  �  ����������  �  �  �  �  ������� �� �  ?�  w�  �����������������@;           �               � ��             � Ċ             � ̊             � Ԋ             "� ܊             /� �             ;� �                     F� T� d�     r�     ��     ��     ��     ��     ��     KERNEL32.DLL advapi32.dll gdi32.dll OLE32.dll oleaut32.dll Shell32.dll user32.dll   LoadLibraryA  GetProcAddress  ExitProcess   RegCloseKey   SelectObject  CoInitialize  VariantClear  DragFinish  GetDC    `    �?   p    h1l1p1                                          0�	*�H�����0��10*�H�� 0g
+�7�Y0W03
+�70% � �� < < < O b s o l e t e > > >0 0*�H�� ����׾8�?�l�k�ZU��
X0�'0���0	*�H�� 0��10	UZA10UWestern Cape10U	Cape Town10U
Thawte Consulting cc1(0&UCertification Services Division1!0UThawte Premium Server CA1(0&	*�H��	premium-server@thawte.com0960801000000Z201231235959Z0��10	UZA10UWestern Cape10U	Cape Town10U
Thawte Consulting cc1(0&UCertification Services Division1!0UThawte Premium Server CA1(0&	*�H��	premium-server@thawte.com0��0	*�H�� �� 0���� �66j���[�ځAb�8�IU����G�H5:R�+j�;/�V㯆�����euM��	�!Q؛�gк�sԓ˗* �\N��R��Dn�Jn�/-���:�s�FSXȉ���s?���BM�@�7 �00U�0�0	*�H�� �� &H,�X��t��_T?���x`^^n7c"w6~��4�����8�M��BC�ZF����J�(F���B}���YnշQ�㤅k�L��餮?��Ie����>%�����2q��^�P'��#��˦B0�N0���
0	*�H�� 0��10	UZA10UWestern Cape10U	Cape Town10U
Thawte Consulting cc1(0&UCertification Services Division1!0UThawte Premium Server CA1(0&	*�H��	premium-server@thawte.com0030806000000Z130805235959Z0U10	UZA1%0#U
Thawte Consulting (Pty) Ltd.10UThawte Code Signing CA0��0	*�H�� �� 0���� Ƹ�'`��ie�~�������m�,�pw�&�W��?0��!�h����.K�5� ��J����ڈ� �!�	G��	�y��L��nT�i��L�:A�}�d{cE�``1�����n&$�����Դ��P`�Y ���0��0U�0� 0@U90705�3�1�/http://crl.thawte.com/ThawtePremiumServerCA.crl0U%0++0U�0)U"0 �010UPrivateLabel2-1440	*�H�� �� v�����-4��Es4܎k.\�L}���h�י.ȵ��͊�I:[� �mR�v���e�"g�SS7F���/�{��El@!�]uvf0�߂�/���۟��r7M�wH�J?	�U,��$��0��0�@�;����,.m�F�[_�$0	*�H�� 0U10	UZA1%0#U
Thawte Consulting (Pty) Ltd.10UThawte Code Signing CA0060113000000Z080113235959Z0��10	UPL10U	Warszavie10U	Warszavie10U
FAST TRACK Sp. zo. o.1'0%USecure Application Development10UFAST TRACK Sp. zo. o.0�"0	*�H�� � 0�
� �pjLfe�枭�"�b'C���N	v����:���j��C,�ֽ]m�>/	� �j$���==�BE�	�K�z���d.NE����q�PŶ�ȑAd��L��7�v��Q�\�����=�m]t�GTWܣ�:�)�o��Mu��r(Ҧ��+��ӫ]����ݶ,�V6��4�WMK)&��6}n�v M�]՗���5�!	�Eb,k���p�c?-�^�{CArJ��޷�R�?q�-ZH�QVS�C��oS'��EV� ���0��0U�0 0>U70503�1�/�-http://crl.thawte.com/ThawteCodeSigningCA.crl0U%0+
+�70U000
+�7� 02+&0$0"+0�http://ocsp.thawte.com0	`�H��B0	*�H�� �� ��uk��F�(�#�r�"��,��JԆd,�����(Tqj8��®��>:�{)���(��8���Nh�8�9��4���y������wMI���鄆yK�26B�G���;����+��{���"�[1�0�0i0U10	UZA1%0#U
Thawte Consulting (Pty) Ltd.10UThawte Code Signing CA;����,.m�F�[_�$0*�H�� ���0	*�H��	1
+�70
+�710
+�70	*�H��	1[vᲖ��Ӊl`�0&
+�710�� F A S T T R A C K0	*�H�� � ��K;�G�"�٘��lr�=��(fA�x�̍�LeW�L��� ���;̶0P�`N��7�%�;�V�,�o��β����Ġb�rKps~�A��(k���rvbm��4�{�"}p(�⎻�nj�����/ؐ҆�*����.e�P�T��E����]���rW`I������m�k<i� ��vJQҡ2&-�c}xbڴ͖�}N]4Dl�;#�R���A�d�S��mn΍�K2�T�ೡMU     