MZKERNEL32.DLL  LoadLibraryA    GetProcAddress  	56�kByDwing@   PE  L             �  % Z   �     q^     p    @                      �               @                       �` (    � �                                                  �`                                                    .Upack   p                        �  �.rsrc    `  � �                 �  ��`C    ��B     ����                @ @`C �`C �`C �`C x`C |  �  �@ �_C �_C �^C �uB   �`C �oB �_C                           ` �0  �   p  �
   �  �     �    �F4       h �H  �    �F4           `   ��   �             �F4          �  �    �F4         �   �� �              �F4       r ��  �� ��  �    �F4           �   �l                �F4             �l �               �F4       � �8 �    �F4         P  ��             D L L  D L L 1  D V C L A L  P A C K A G E I N F O  M A I N I C O N          �   (       @         �                        �  �   �� �   � � ��  ��� ���   �  �   �� �   � � ��  ��� ����������������������        �������wwwwwwww���������������p��������������p��������������p�����wwwwwwwwxp��������������p��������������p�����wwwwwwwwxp��������������p��        ����p�ffffffff`wwwxp���������`����p�������������p�����������wwxp�����������`���p����������`���p�����������wxp��������������p������������`��p�����������`wxp�����    ���p��������������p������     ��`�p������������`�p�������������p��������������p�����������`����� � � � ������� � � �������������������                                                                                                                                ��nd��׎�A&��vN����p���T/�Q�΀�S�
�S<����#���$6F[�/�Y�ؾnA��xeŀ�<Ԥ�����<��&g/�=�I�V�PJ8=��Ч2���4���{JH�[�7Z���7��D9#&h��n��nŰv�1F}�g$L�(^Z��|�py���J�W�z�-�aK�A�"��J���u������}[���	����26�C��_ۀ�M��2���S�0�~�y/ ���A�}��+"�<Uu�"�A��;�-9�5�UV@�b[q�N[l�^����|Pt}�s����I������V.N���"8�/c!�k��!@u�����p	�n6�Q��� �CZ7��^�n �9��n�
O���q#�%���8f����&�qP��	Os@+V��y]����ɛh�p�R��]�V�,_�~>3�!h �c��z����2zۤ���齬*u3{o@��g��e�ٸ�៖[c!�nΥ�
g�h���sJ}���Q��Bk���9���s١��y�Y�LկUU�"DR[�����o�(��K����ϻ\�����4Qg��~��E���6���x>���2�r(b�`�u�!��V����'�a7m*���}"p�5��5��Fit8���z�o�+��פ�1�%������QH3+���>y��o��'_�H�w��'��R稺
�!��S7Ci�|]��3d3���ǰ,׎�h?�������3[��e�I���g��PW"���	^}WU'��6�ݜ�GO�wJ��x@)�̄|t3���(��K먾�������|�?�� eFzH�c��b��6�CvZ�l�^tZ+���v'\�\CI�|�G�:�gݔ(�H��Lv/��i�M*�,��Cy�&K�Y:�B'f`�麂��{D�WDvh;�ʽ�c�/�?`�sݤ��x��aY����vC�"Ƿ_�W�*ۖl�})��z�æ�����)�]%��F7��T�tſ�7���A<hD��-�U"���pF���\���TL�)d� �3���n(e��j���ޞ�t1�׀�p�i����������!� �	PM�_:�7���-S>��&3�7c�K��& ��쎖�c;�� u�ռ���� ��X��8���?�䷴�����J?�IK$����Gy���g{�����]-E�ߗ�ϐ��H���?����d_��4NfS��1��JRkQ�P����[/�%�>���k�H��)�k���0r4����A�gpobZ�F5����qn�/�(Ed��?��e"',����\F�F�@K1���n_i.���Gu��b��+[Ŕ@��* �ANoA����Pժ=%�I�F.��Z_�.+5�҉\�k9��0�a�K�c�H��Q���ߕ�j�q�q	9���'- ��)�E��;&�Q�Pr����]Z�r��+��+��ۭ2�OC�M����Bn�23�>�z�і������m��zǸ٪�~w������U;�l��S�%�o%j2���T'�T~������O�x������O�S�ń�wp��n��T�b�+��9Hh����a��D.n�=��s���/D3���c�i�9���`�	�Q�����q�һx��&SM��:�K;�C�gz��&�#���GP�
��B\����Y*�+>� ����	6��}���-�95�	E�na)ۛ��LnMc�X��X^�*�746�SHN���Jop�!�%yN� W2�u��dF�>ɛP]�a"����xe�b��
��윌z�up�|`&	��"��X?FRJpzQ�*�X�4�y?`���n8���c5�����$�۩�j:n%��,>��7$����I�Y�(�[1�Կ"P�]s�>r�I�u;K�A�P��G�^vCm��X�<Ϋ�ݍU�t��KJ�#�U]o�c�G
���-�(���|u3�h�_P�&�xlU!�oH>'�m����>��]3r_T�E���PI�͇B��� ��=�<X�_!�gqb;>\�$&�}���1t!����/���/V��ꉭ���ݹpYm����D۳7�=��&	��*�vͲ�L�{��qV���n5���1��ŭ���ac��%Ӕ�v����f�"4��[]��g�LെE�ٝc��_EC��D�.�'����ֱ���Y
q�P�&�<"Ѥ9h��7�g�a;�KOm{I۱@c�����|�g�1,�."]X�p�s��1A���z��
�_�]a�h�(WP��I�n���!�s�lRЯ�/ظ��$��.L޵�6P�©����(%ߦj��֝`|H�L�?��]}��o5�'��i O;,y�B���k�)��̴P�%��Ât*Yv�i�-����ײ�>�ي;ܔ�A�w�M��	H�p�R*��Zc{!�����9+V�q"BicP)C]��j��K첞�Ը�E�d�4�li��F�#*=�>��.�e%��|�X�N|_G���}�?`j�MU�|>�j3V/�%I�eWh o�W���]����9�p4}��R�*G��Dړ�!�z�f�)�hd�z�iU�`Q�@e���Y�%3�Ol$���Uv�0�ř"�Ɛ,�`�>#�^.eG��~�Y�8�s�_򺙲��&xR�Q�Z��UR-���-�;j��^=Tl��.b��ŧ=W�H�r�@ԧ�7�O�|��y� Q�uh5q��8���;�ƌ�e����L����'0������h>��H��k\�n�"WKz&_���p��p��8�`��3�fw�_�K�d�9�23q�U����!��,!� �T�g��絧�?��`�M�������5�|�Y�CF<$��p[R<d�c>�A����Y\�"�������/.�����eA���b}#�S�L��d�V�m�LȨ�J��4��N/2��
��*g=��-�$h.��љ�t�����A,l%?eo�*�B��Xz���:L\��ƾ;��$1���>�F5'���	PV'kħ�#�G�q֢�wa�iGg6n^E�j�i0u>�p��GCΤ����6rGR�޼t;IF�o?�`�0K�
���e�w��m�#��T��e���uOU� 4X5/��yGF����
>Z��P��N�A	���~鏌x)���V�����C�vg]${Ӌ����i�#D7u~�O��tm��L�(�ͮ�Y�w.�����^v��������^�>���֧b���͞+�7��}N�z��V���<p�E��QHY�I�{��ş��!��ް�Uۍx� ��{0s'�ľO��c���~�Y�����I�}�Ŏj���v�@dP��4�h�$��լ�"���L"��0�H�롸�)�Xt��U-���N�����+�+Z�m"�z(��3%� �g騾ܯKa��bL�B.���ј�s�/��������3�\����jt�c�ۿ\pچhR���N|�A����ڳ��!{�R9��)�'^Yk`���ڬ��<lЉBd����z=Ţ?$�:���/��V��"6:Uf��λ:"���@'�������M���3�F�Qc���*�vx�J�KD9��4�gS2ы�ϐ���T�J��j����/_f�;�F;��O�L������0�Y�r�䥎ڢ��"�R��y5Y���i�pxvj�c����I�������(��)U\��@t��	�F�X8��]��֙�ԣ�9%u"��f{��m��6<�c���?�f iv3�`�Q�H��ֱ��`�����)	�KX��Io��;y�?�J��͘�Ւ�eN�#�<N~DyWN��me2c�2�u�~Z"�R��+]��)׵f4 z�2�f06LE�6�&ݿĔ���H,b��¼Y����B�q���p�
#b)�eW��q�MA����{���Ӱs�Q��?K�Æ�0����Wl�-��~�B8�$gc���Qo���m��T��ka[ʞ��Ȱ���4E'�b�'��m��?�.�}�6^YI�s�G�[[Q��O��|S�:����������h�Z�L�:�۱}|��SPTz��o�c�*9d���֥�:g��j��̸ ���D���c��A7ݕ(����jM���BHQ �37<T��i0�x���/�%��գІ�B5�H����	�t������+��߶��F�2m?w&�g?뭙~O<��:B�������Ht7�/_�����]�"� ��^+������#�L�w��̡���O�]�F� �h�AN	�_.4x0~^�������۳-��noN�ͽ�ۻq�K�}��Ss�`"�Y�O��H}1j�"��_/�wbB�B�ލ{�����V���#���&r}m�+�z��� ������c�4Y�����|}I�~X0d�&�����4���D�����7�7H��a����X�f?֥x��k�V�eTn &0�ˢPfE���@�W�c�7C$�v9��0gW9(��J��_}��^��
�OT��S�n\9�#����m�"���*ӣ#�ţ�Dc����`V����I}-�?n�}ƶ�cm)ُE��I� '����0��x$�x%M�qd�n�F_mC��&�0��Zm�$Ҩ���q_�=Zy%\��v����n��4��RW��K�JS@�N�-����csX���]3͉�:�NX��-� K5�J(ϐ���څ/e���Č6��gX��N�G����)甔d$pC`(K7������){�=�^�렧"��y��ٓ����آP�co �\�x<c����ʾ�^�����9�����ޒȪ���o�%���L�cJP~�C����������a~�k����Im��lb؀OZ���Z/h�lnz}HH��ʍD$�|26�i+�HA����Q�����;2�;2&���!��j$*��Go����m�D�Ȩ"��Fo6�l�� ��͎�%���ܗ�aP�z��G���9H\`�n�E��O�Wx��%�ꮺ�Q���Κ:N\3vs}߯�l�7#h�>|� 񬏫���	W��yrk���O�aC�Ù�
��Y1��G�j �!�nuz�I��=�����"��LtL��"NCe��G��˻pȣ���pnr��,jhӐ�t�MTwd���p��_C,�l�Dr�� ��#���>Nӭ�@27ؙ`�qoly��lb��K�%X��&Ef�����4��xP�F8E�9�3�0�|�2�T���N�%UU���T��.���1�n�HBZ{Y�i�W��wi���fo��ޛ?m���p�l٣��^F�"r�C�sL��� N����E:���_��|�$q�^o��?��A��{ךcE��V�Ȓ�i����hC���]ӏ��T�:,N�e�3Zi	%q;ӄ<*���}U�p�Oj�!
��]	=�&�<���D�擐=�X�w�f��ʗ��iɯGiu⹐���Em-͌^�h%�l�}b�N��Ͼ��}�M3r$(����5��F�O!7����J_���}����1�b?AwR�W*a�L�-���V(�pf��j��L�\8����G��C���=O_����'����Ͻ���]y)�&&��4��X�rY$�T���o���[�Fk�F0r�����@�a'M�@��Ȗ
`�����e/S�̒���K~b�}Ln�l�*�����ig��q�� ������)ȇ]����(x��r�a��?,Bw,dD���Ey�6�p���]���L��8>֢Q���ޤ��AX_s�=ߒ!Z{X�_g1�&z�5���k�IaIfN��sɘL�!���
 �N/��)k,��I�&+�+��n��X�7�zJ�5��Zt��DZ�m��KCk�)�n�i�v��k4{�S�$���1�ɀU����n�-X^�C7�RF�֎�ӻ��i�S���7ƌe������%�`�=::�o
4�������I�}&��C�e�g���������`����M����d�,�S
��%��ף9�Tu#��9�͘�i��k �(c�M���J���;	��X���vL�Ʋ�U����9H���tP��O�CM���ۜ4f�5�`�:��_9�胆7�2��p���9i�3����#���$p�q�'jB`��-"�����]���ء���NX�i����:���u}y����OHX�Z����xo���*b#HJ$ٳE��1�C<��m���e���{�I姇��V����Je0�@�A���n}�,�������w�J��e��yoJ#8�ҕ���l��]vC�qv 5�����4LpOAu^��MD����
�W�tΰc��D,?�5���?�hJʈ5�5�$;�pWo9�F@@�Xa�4���������M�T��_ ��?��T"M�98#��3�Y���@+�_�3���!	�ߡ�/Rk~�)b��Bb�Ѫ�0'��A���W������P�ebr����X�6������*���W�Ʉڵ/2���6sM������I���_�vO���X�&ۓ���̃��t��RqW���'N����Xv�m�|휆�5����^8���Ƈ��E��A��pg�0����p*�@��7���u� s34>�$T��ۦ�@��A�H��6?�Wy5�Ĝ�:U~�d�e�Ɉ���>m35�g���7��8�B��1��Ev>��ig�4)?����T�ɉml*����*����~����ݮ���_���}���WaK
���A�G��d�����]x("�%�\<�Ϧ�R΄\7�F�1��8	�����nv]�F/.b��L3���;M[O�ճJ�OCo��_ݺ
K��GA*��� R�mS���1z?���gc��b#���,P.Y���a-�Z����xX�P�a@�.��C �k'��h��h� 7p6�25��㗙�ɠ|���Z���6�2��MR*<J�I.�Ĭ�W�D�~�0�$]��?��/4�ǪW�8��ےodLeY\��x��:�꘾�xمV�t���y@���q���+�sٻtt,a�+�֥ �k@#�}����N��I>���R ��fX����#�k���O�$q�-џ,�O�V򋍝�M,kB��@r�数�4eIa++/�T�y�*����?Dv�?�#�@~d1_kP��a�3�X S����Vr��ٿ��Y�@�1�q��5*������3)V!a�W�Ԉe�!	���'�U��7n�ȇ��1��Z���(��:�	�.�q��:�*?v$�'D��;[
���K�h'��o=�%�_N���#'$�%f3��b�/��#���u�2,5f�����z8�^͈pr��)��N>K�������"���@�$�Aq"`�_&x��قk�
����z�]�5�Y|����$�=�Ho�$t���EsJ]vo?=#n��V}�3��ǫ��b`�����<d^�V�1����MU-7���2�\5�h׊>[��!D7�cNnR��Gu��<�o�?i�P��K²R�8�)d���N=erz�$2$���Q, 0y���&�S�%�Zvfя�p�Ȉ��nxNc܈��6�ݓ���ՙ6,��f��Škۭ�68�J���DN�����0y�-�mCW^X�UPv#�	p �v�[G�b��v�>�SY��MT�1��!~�l�q������(��7&U;i��=�\�	���(C	����ow�n�`yy�<�0y7���u�D\�����!=AұS;��i[����ͦ/�<|�Va~!��c���`�V��J(K �N�CǦ:$a��ӏ��QiGO��r-��@�����V����C��xZ���h����2�'�_�yD8̞m���)��&=R[N]�b��ڴ��]���lP�t@t��p�OL��j}�y�zcZ���"�Pti75
�(�����TpP�~��U ��������f�Ӹ���g~�7#R*��k����ߧ2�A���@�q4̽̋n;���|�r�R���m���<����.[T؞D���Y�-�v��5͞2�Ċ�η��3�1�}��y K��Y���b��(j��˒���H:�?cC�E�D���iv�$遳�ǎ#�������*uM\�axy�h��8ݹ�!�+U�L�Z��}��M�o7,��}"=�ikH�h�8%�7L�9���х�(�#�`�^�/yƧĒmTڶ/�&aX��H.A�n!9X\�{��Q��Cy�=jm	�e?�gqTKn�ٰ�$��"���-S��'-<XS	�W9�����,E`����)�M-����	�$#tk�
�e��Q��bT�,��?�he�"�:iz7�Q�w��oY{�����:H�0(%P�P��AIj�� 7^����i�`Yc� n�j艙{�`��aN�cl+w���d�\����t��o���W�I������W�}��[����J�,���4�!S<y��8B[��N,i�*�N~���'��h"vW|��W�2�.���1qN�黅{�Ȳ���I�\�ľ���v)P�k�#�6/��B= q�c`���`k�XV��F/�"w��N�ω"�f%��7�v� �:#�6���>��5�1�U����%9	���lB���q��  ɩyڱ4C�|�8�>E��W��$C<�[
������R�^��$��:�ƶ�d�Cٕ�!gʱ�D�s�m����`o�Gow�B܃��Q�!ß�b�����;�D�
��^;�vd�y�Y)�4�v�wH/���1C�!D����	�$ڬ�7$mjM��v�|��\֏.��p����{0n�B�e5���K���	��J�x�v�5��a��x�G��N�m�qA���<��m7yS��r[��$C�	C�f�,���+a`ټ9hT���<@���*H�"����v�Q�� ��v�*{���5+���*O*3��iA��w{ iʤi��D���,��?�-�P|E4Pq�� �z2~�;�ꑊ�O�	���:Qܷ��-V�$'5g�&���[N�J+��Vae���Qꇰ��
�&{�%���W9Aa7.ƞt"K�+�n��������%��>���h@Gﯲ4��3�*��0�6z#���J]p���5��~�]���vJ�Ry��Aۄ���K��
��\�i�H���M����L]���S�J��J��I�� �o��⥐;�:^)�)Br����M�5MD�Ö�B�9B�`��ͩ��e�bk�Zw�^�20��*��4dP�^��J��׀&u��f3��;Q4�d�o��oK]YSP�z@9�^�,����y��=���E#W���4��=�����4���3ːۻu�/`KI�&���!�w�F�X��p���%����y�/���mB�|z[��F���b�&4~�@RD9 �ƪߢf�ʹ����d��PMD����v��yN�Ma$�㧛�ɒ4�Q�{���q�,���������1LC-�ɡR~~�|�B�`�;�[�ݬ�lr74�3����OX!��m��2	ͼ��۲�Sc�M)�ET��*�7�s����r;<��"�p������C�����Z�\�C�M�j!5�3��ފV5Q��q��}U���h.�@��m���p��PY_�y�T��0
�X+a���b������Eλf��J~�x�c��E�
��A_{��E������Vdp��ѣ�m�}5ۚ��bU��U)�Z��?Pv ��E��]�S{��<:�b��P�R&<������R��A��\�#��9�������[p(:�Ci��K=K/�Qh�������8c$�e7q��]/3�A����i�J�:e�|R�����=��!�h$̮�1�8
�#��Z��sD��.nA� �:{�<W%�9g�N��Lʻa�C�a��dO^��!7�ęTf2[���LMH��`���!��׀��M��7~Z�����(7�R�q'|wo}E�qq9���$�2ga�1i=j���	x j�q�Nh~��
��"�q�CWm\�>k��_Yc�m����_83�
Tz��)�&�/�����W'�q��P�(B;/��`�ŁD����E��˰�����>������Wx�.�h㽇x��FE�$A�)y���|�O��t�;�ķ�:�?W[���S�KC<�>a�9Ýc}	pQg���Ao�$8~�ŉ�` ��8M21 �*~Q��6� 5�5R�ނgd����jલ��ҳe�d\Ҽ���\���H��3��1����ϓ<��=	t ���vߞPm�`�>� wj�z��+5jq�:�VDK���/E��ԭ�Uv�N&A`���#���� ,!��X�=��e.F��R�]�}��>XK�L�"5��zan)+^ a!��N����wf�QJe3%P15m���W��w�J��z� �
	��n���YEMz6�G����&"��o�2L�ь��[����"A���r/'~�g5�&~���m��\�����I��M6���w�Ḣ����-P)�����ә�< �ph��r���@zr�mA	Bs�B���vO�q�̀iBS4퉷�9��4�f��Zz�q4�u~�v����&ˁt�6�������L#Q{����͟�	hX��Kj�t�ϸ̍��?LF�ڨk���mo�[�{Q������C�6͡,0E_(�����	B_�jІ�=�v=��dwlF�Z ԑ��~u&l�ɘ�/:��P��v�̆����Z�c�2$Ha�-�_[��k`�
�b�e���ʠ2���$�z�)�䱣�%�w^�@L�Z�z�$��<B� �Oy���Oޏ�j0`�O�e���F(��OK0�fᛝj�7������cB9sK����.P�cf�/�~h��n�#����n��IS���]�P�(_�9ӽ�Q6~8d&[�e�<�*�%J��0c[�?�<����~y�zY���%�9J��Bj1�=T�z@v/�p��r'th�Qf ��uj6�˧��jKr��4Wo�X� �_������c���IF��˭ލ���=�"�;�!IJY`�Dŏ=(�'x.�e\��̏Jt��T�E�)�pI�c*Ky[�DV!%�q�ޟwc�T��y��,;@��1�h�煂n+��)|���/Ol� ��^@Fr=(�JGEBvA��a�ɔC�X��W+.��J�'/	h�I'R����b�(x���n���S.(�|<��&�H7$����i�T��<��L�ʨ����}���evQQ�f�<2���������E3xP���2�%mCِ���)�(��N��S�����hZ��;$Bff���f"(�ۼ�{�lRd`!Oȱ�n��\l5�B���d2S��'��H���(���w��\���B�}���1f��ڜݼ�o��q�D-Í�]�p��ș��r�*��Bn��:��y���#6�����d�����i#�9�{!���v�����qe� I��D���������_^ �-P��P@^C�@|N��P��W��Ӻ��x^
8g?�N}�J1�{�	ӇiyD�y�A�����rfG0e���p��g�&���q��l�SOJ*ըſ�Rq��F����B��UzfU�])�>�1n$�N�2S	O��N���Ԏ�����@@�_|���w�U]��`-�wWe"w_{	��5��c?��8m�ָ���L� �j�j�vC��DmU�..b������B;1p�X6���)5��7�yX� G�5E&-zO���`:[�5�fM£�^��4�0J'0樉Y=��Qꐁ��<#/���^\��v�L1�u"�v]֒k4��	��zԹ�i�y��2�W1{�����,�@ƴ�?h�6�I���㎐5?gۖ�@MO$�ꈡk(���dcضaw������K~�� �_#D����ד�լ�I<oQ�m�c�tGY��^~,��I�W����}�m���}@��;e���6���<o�2H9�xe3b��,�ڣFŎH���퐭Ls�Hs֘ZF)N�����s��\�Q������>s>u���q5Ѭik��m���a�p����zo$|"s�ޑ��?�Y�+�@zb��wy˅U�����R-��#�t�DsB�Q�OZ��{�P�(iL�}��mpO���2�W�J¤��u&@*���up<�-�1>
9�H�l��E�g��ڜ�Y�ƶ�W�qn5�i(�:����=`@�P��"���GL��xU$J?�W�ya�@�O�!�bz�bt�˜��.������
R�f$Z��ߌ0knx,��w\ ����0�m�v�.d�,CZ'��QY|��?�E��IRvm��E���%"O؇0��5�L�-���aײַp�-e��u�~���@V31j+��!D�H�E�������]$�t�_�E��(|@��,�hk��f2�ġ1�ԕ9���:S'.%��g� �����:�_sj����8�f�e�X09�gu|�:���HC>�`O	imwN����V��ڽ4�"���bm<�Ue
0-�����B�ךX�^��
����oi��$�-}�[�,���eۙ�>�ӓҲ�/歹橓���@x*"~3�Ҳ��9�I0=���X��f��&���H,�ڋ_]gY�����j��,�H>����NƅO���I����d�+ќ\j���(;��(��n�R-d_R�e^m9xZ֑���.�M�R�Z��p�V���+�=58�/����7�Q(�g�x4���Jm�p%=.��=��y��a9�!t����)������z�ݛ�:��h2.j�jH�'��r�>Qt���u'qx��6l�4>b�g�',6~&8r�v � ��Fĕ��{��a�:�����6�+-@h%n@�E�ClN����!�F���,�!� ��C��3C'"{Ԡ���x�^Ά0kT�+�=e�7&BtO����a��'�*�Zŀ����x�?��5.x�O���>}�����"�[���`-vI|��:IM���c|�c�f�������N~��>�n��a����+H��֮-;�F�=�c���T���ǣ���Q_��c7w���(�ަ��@�R@��'�R���ކV�HxZ�?+G?�ڳ`r�c�4�ùcV(7��oXe�9Ձe+��Xt꒘���OB^�ՓH;�����Ŀ�])�,���o�8�|	����	_d��rk[Z|u� nU�B~.!��>�'������ˉk��LY�6�q/�����DXd]���$��XM�tf2��̈́÷a��T]poA���q}M����q�
ֈ�x�͸sI��3X�V�V`��^w���*���<E:ט���7�U)>�)?�Ϲ �̱X}u�_����%z3ﯠ��9p��?��E�w��E�@�4�S�� ;w��g�H��fʪӺ�LM��V��2�@���K��8�M�Y�ذ�m�������*M�����{ Bz�sBd(�כ��A�
����ܫo�L������̓m%��$b$&�!�]�{6
�a���g�kZ
B{o�k�\q����0}��s�cd{$�:��,\�e8| �z���h�a'Sͩ&gLlk��Ď�薮�D��&B+��Z����zMp-8-?��"'��]�	�Н��R1S�����`P�4��t4nz.C�]�=�0ek���M"�o�f��B�K�B���O�\�|ޱC$�hF����q���i�z(%��z��+&�=��x�?���F�	�?V�0}q
�$��:�d/��}�������a[���S0�+B�C���	Q�,#:9�)M���I�
r�ψ���K�(����O�`����_�����U�NHap��� 縃ą�����NЍg���B8�U_
��ܻ���z�����D��o�������FYX����0́�r�P~(��,ا�����;�vY*E�ZlG��]t��osI���/tfEmd�12��aV����z��5��!�ǤQ ���������QI$�n�a4K�0�c@e�4=�}�L�U����-\���IR�2��>���4ĺרή2��u��>Ȕގǧ����oO�2	6�ZrJokr@�EUb�$� ك�����n�ɟ��*�=��-n�j2g�7�{���]�\���?�%���ۍ<y��U�N_�����Ӹ�yuZ�R?�t5=��7/�숄J����ߨ�m?O�ɦt��"���Yvv�â�Gˡ�?_���sI'�]���
�"���g���`��o�L��6FX~�����*cp`�]�Dy�6���'�E�?u��$��I&�c# MK����Kt�CPJ~�B����?�Q�ʔ�ټ��u�����q:�Q=�	��{���a�K��4ո�,�����
Ҿ�\9oc��	-����Z�zȝ��S�E��:NRZ28X��R�����2
��z��mH�"[�N��)�u�oګ(��'}3�|/w��}q�hj�
���5�Ww�L�:�G-��Q$?��H�zp���k����!��%��ސa(�5�ؾB���C��p��vX(�*�S� �@�Ŧ���w�5���RϝźWD��e�_ڊ��0	�Jd�C4�ս���ѕ�(&�H���ہ���*Y@�ڇ�]�]|&��`�������ω�SA�_'>�g��hu�1���>�J"�z]��w��om"<rg��-�����i,o�2-Ͱ-��<sޔs�Z��;J:o]�>\i�6�]p�����nF!`Y֙��EDZY����ğu͞����R���QtYyv�ht��Ù�_cZJu"�W�=�w��z��_р���`vO�����vJL%fX˨�J��:��t�j�-:�����Y�E�i@H��u�c�3ŸM�Y[)YZY���&.���S����M�C��	w�=m�
fy�;���y����ڊ��f��8�W�;��ib.������R�A�\�_�4E�o� �.��7���b���<:���,/��K�.��lI�GqL�2��i?�/�܀"R�ݵ��T6/��(�y�&Xa��/%�v�<�]��/���M���@#+V�<]�>I9��ǵ`���u毳b3@}#[m�{׶�;�m���i���*gG<��nsE?�N]�n� ���������:6-m������f�ͲGk�B��M��,� ���P�Z����$Ŀ��G�VK13�X���m�o*��m�Q{P���k�-�!�8mUU��>:�'�+������r9�����Gcm�(+w��Y������\:��f��Ϲbv��X-�E �P�v�3k=��;�B��n�z�;YͤC�&����W/Y�0�HL@��h"7���v��N-g��a7+S.P%�$�ϩ��S���O�n��� ���DjnK�P`�|a��,�Hu�U�d��XÅ%�D�[��ƅ-AǮ Ӥ�Z?$���U6WsЯ7�Ygath�h�6�\�q4e(��}W�$|��\͑���Y�%�,y^bZ^��&�40�7���r;<��xy�?�%��Z�=_� "�ӱe�S�������~���,�Ur)�{���YI�Fn��Z�$�{	6�4��\s�6=-�,*�3�C�J�a�q�@�%ʎ_�c�?t�B�p�[+���;;I��?�!zQ����Ź��^�Xq�Rq���h�(h����7��00\m,n6H���#`��A!(R`ig���2H���e�����T@�n�6�iH�ځ
��\Ť(>�����>��?�	L��O�&��֯�+k	�E3��Nb��rB����J�eD	��q0_��x���/��MAG�.HB؊��|�V��K�-]� ]��e��KLZZ�LPr2�q���Ӆڀ\P5��m��6�wh����sc3`PO�Ze,d'�IՃ�'\�͏r�/ׯ����\�?��<�@!�FW���$d�]GzM!���WRw.z+c��� F^-���h3LaL�@K�9�L�}g{  ���:�Z:ƪ�w�|1�րOv��c �ޛR@�/�[�������+��o:��.�~p?Uؠ� ?5�M�<헫�z
�^EU`�����~����R�/t�p�r͉P�0���dP/v�:w���3Y֎�I<�v�}���N�ز«����%�mtHvjs��x�3��^�� ́o��aLH�h��^�׹���4a9u�0l�t����(�4�a���;�<��X�`"�������nP��ǜ�ڑ�8���u~�}P��#�W�Z���+�##�)�]V���Z��@����)��B��$�W�$#yd�x��%/<��{g|�_�t(pz�v�LC/F)=��1��°�=#����c���N�!Y͍�G�fa�R8�Oh
�~Y`Jf�Nv��.(J��۔���6}���˩��z$���7󇪬f�IOZ23�����

 ~<}�� Q�eA���m��-�����`�/�o���ޙ^�w����j�TY2�X�K��H/���FlԻN�%�M���\-��
;��Ѯ1��t�+_S��j�L:�5���ś݅E��m�C��tg��Z��Z
���a�=UK��/5�l��F~1��E�߫�É:C�T�6��.�v��<��<$v]%6�A��f@r|��fJ��*0�?n��8�pHݨJŤ�?O)~��bb�C��_��ٹ���i��X�M��]�m�@�;1]i�2Z�U��A�/�E	�A��H!��M]eA�1"M:�˯��c�Cr�;xO�O:J��J�a�N4�K'��g�k@ծ/��(SМd����b�}�h����Kf���O�0�)�v�W��D���T��Z�;Hn�
ix�ݯ�f¿W������o�g��q^(Y�����M����m��
�N��'�n���)1�n3rȊp������a(�?�A(f�|��d�*�\�*��j�9Wk�1�<���1j��/Ga��#�\�,ΎՄ������J~�)����ԀY` LD"h6;Q�f҈c��H<��E(�_]���]�h�<iLm��n��-�˵~��U�Fs������)��$mh�X�}�w�1x��t
|�h恲&�N�l(�{�@s�D�j�"��7b��bC::���_ًYT�2Uzq�$�~��?� ll*݇{"&c3Q����� f�G�ȐΛ�������~�_l�߂.T�N��^�
*̜���ǡ�{��ݸ6*3��W���Z5�C���ƞd⭿)ɦ��ZH]vJ�'����fH�T�L!T��(!5��"ε(Ү�W��j��nu	W>KZ����[Z�N߄����!�oB�~���r�8���{��R�hL%7�P^��3�^.w�	��y��vsئ�	<�����M�ɉ�^_-h9�QC0�\�3��[O�6���Хt�N�^Û�&�1�!UL��� IRڧ����W�_�����ja��Y�j�+;U�<Dk��)jh+�J��W��<^�J���_j��#Z�L�M<��S�91�|��d�.��������pH��[�9��?�^�I'�1�Z��U�@� r�Bpt
���w]�;)�_�ea%�i9$2*������!_f}c:�H�6��Y`b8B��Ϧ�h�y��~�F���уG�>��س�����m��p��*w��Û;�����P�B��� ��ޫ��"� c�
)q�N��Ĺ_�O�52�H�uW�	�1�v�T-�:ohB��=�"�lE�ʡ� ����V�����Wr�Ĥ��r����\j%�7Êk.&�WnK{0��hDU�/o!�^Ώw��>��֨`�)�:�����6D�Q~Q��}��\d̨r�PHZ\N"tS�k/r����5���?!M��R��-�$��AOgSw*�-M�����p�r\�8��B|i���mw8������ڿ�T���0x[ym�$��v�L"������([z��M�H���ve��
�_�"�vV"�,����0�<�;J����n�/)$a�2�,�L	�l%\�#d	�v��$N�Ӥ�I���q��\�e��4R��.�����n϶z�$
��l6���{��@���ނ��G܁�7�p��t��0e�>V�P�^W�o�ݏ툨�Ii�	:\��I���Vyۥ�4���u�X�C���fĥ��� �4���m�`�w1hZ�ڤ��
���ϳ?�I�"�ۖ
�B��y	��,���������|/�ϐ;�#[j�Z��Oy lJ�����\@��3�cNA\���}C���L�=^�*���<��+�!�� ��+��nB�l;�rl��yp[,j ��L�;{W����D�y���`��+�Y�yK�g�u����o����f�2ũ���|d��X1(؋��0������QeO�O%�� �o��2#
��1[�ۧwː5�>d���%N��L�ts1��B���S 1氦Ň��
����#{�F��e!��P�����p��.�!��P�î\�X��p��o<�5���P��_�A;�7
�M�*�� ɂ�i�%B+��6}3x�}80i簤�KY��[poΔ�!��c7��*7 �ARb������ri��9�޷�PV���tc����Ɍ�[.�,Pm�"n��'v����~��4�1ή����`���x�-���H�%3�H��c:e�9a�Ti�}��厥���h�P`�����[��Ոó���c���q��z�]�+�
;�R��Q�+���_)XaU}�N�*�wN!]d��19��'�˵H���Jt�qUo���dm������qM$�����LW�;0t�%���4�
�a�4E���y>��5�%:�F?���<y�M�G��-��L4�^@O(	ҙ����������BG���X���i����$�O��Jy
B8�'y���PЧ�U�����,a'&\;�����V�p��"�[��[�:���#4��x+X��<xҏ�cĠb���b|ׇy�Xɴ%�\
c�v�mb��&���o��=;��P�X�0���A��a�h�D&i҃Mӂ#z��ё)@�W�`�u�ս(l�b��rR��:���s���]WW�B�����7#t�GJ�F�(�L$f�V� �T�㮼���mj�Uߧ��:KUrբ%�J��(�喺��B�=� Xٶ>J��s3���ם!�6	�2�d�f:��rx�mg�Q���
�s�����|�ڌYr���Vx��ұiG%~`a�1w,Q4��8�� �my��W�;�%5Qu���#LS�ȡ�e�>� �@�`��,>� ���|����;ofv�*�?:�+_bU�(f���=���u�UcHvx�	w���]V�tH�a��_�K�8�ޢn��w=�rӰ�g��Z툇=>옩���Op���5:�֤jP�k�*Ƃ0�'�Ia���%��#N]��a��s�m�h�~�g�9��0p��,Wkk�!��m7_5�G��EÞ��ॽYh1��Z��	�d�@����|�fh�I�pm1�k��� �y��{/�"���G� �u����.�DBy��[㒩vD
V{�I�'$`����ӭQ���&-�{|���p�B�8+��*c��@��}K(0!�z��c�����j�K����l���D�6¡�Y}bJ1cx!.��6K��eE�i߃�Fu#2�U����_�QVF<���P�%�aݸ��dz��9�Q4�iz�Z�tFZv1�i/����h���x�0'M�U�i��D�,L��e}�����V����-��k�Q��#'�����sa� ���`0(D2�֍�R;T�����T}w�(��4���a̱U�o���lɈ�c���!��y%�.KPs���?���T�,�����A�޲���	�}L0���X���%�z�H��|f0�'½	65mi�Cc��*LJ��=�Mʴ�a���;C�I9(�I����?b��)�r�EBG1ɼ5QS�� MD,��P��MCEs��w��������k����5����$��!�|{�]��\F��Gڦ!�k:T]O�S]y���"��~�R
����|���ڰ.#��	��zk�~F��r֟���0�F��Ă�lǼ1َ	#W��A���u�L�07���>//���I��#;���a��m>aG8T�gd����L��8L:�Z����xr�;�WK%j�L�a�F����(� Q0�]\������n3�a#���w��&�ʯX�|��l{��\g❬��1��o���u��=���NB�7.�D��1b]tʳ��J�l�d-��yy�2,R�w��ɎSO�e�kcM��n ���Z$"���Y�����;���ֹ$6ArZ�������础A��c:]�ѣ��g	�W����Z�u��)�Fa�C@e)A�i�J=�b4���0(��#!7Ұ�ɯ��)O�����'��N@A=ξ]��kr�3{y�~YI���Ԯ��d��J?�yGS2;<��jAThL�����2��@���͑�F|� 5�wbm�2G��h��c���6������q�b6*y�Lb�{��1
J��֣�^5���c�'^��|�0�1�ZV���N*���K4����ȵ��St�_[ˆ��%�:,�;1Y����d38-���ʌ�����wl(���F�}��"�L]٢��V�y�g�$��Z�,&�l����%�CRZ�>W?o��m�B͑=@I���.��_?�^��K�8��}�"cL#��R�U!i.��;Ս����Q"^�������RypE�:�v �~���LF�%a�>a��H�ņ�+��Gb4j�9tԹ�iD�(�ʀ��6�� �M t�w���^E=~:9����;����F���gX��`;A�9�b�X�� ��U��M�5�]�1y��f 3�dW�&hO�a(�{D~>�ۣo�:)Dms�-;NXy�sԏT"��z� ��Q�ZW�+�ʖN���٠w��砻i�>ȿRx�c���c4����<W��uO��@H�ڳ�Κ`$ �X簜��v�zK�K����� $;uD�!I�6M ��&;��<P_����Z�Z�i�Y�9��j�+X���x�z���oH�/����|VP��>�d��1���>oГq�ES�4����Lqd!냳[FS�O0bT�N�P|tQ���fE�Y\��}�L��KMg���k\:�φ�E�̗ h7QlU�H�\�1J@�����~\�8��p�ˋ@ ��ũ��}A��/W'�9V�Pp�&�y�?�������s��T�^���qҏP6�za�G���_��	@��]W �9D�}K�:�;�8�f+��U_̢���Yę59��Y{ҡ�)�����H�3+���}�>����L$N�HU��&��XN:���^�u�lp�h��&ȱɭC|gZ*��,�+PUS��	
w��p���}�KM�O����P_��J�J�{�DO����:�m�}��|���5lmM�l�;ҽ������P��n]����l踹oF�G�YB�]�wfU)��7/��k�9��s�z\�
ځ�ˑ�D�����b��͖=N�u���)��lY����T~��E���!.tT ��b�!1@|�^y�Z��
F���et�"u�|6�L5нm n��B��3=A��>�L���H��W�ye�N��������V�s"�:��d�y�%�D&����o���ҡ����~�5�s�E��E+�_��&���ۂ�뭲Ƒ�<�v�u-��WN3X�k3�h?s_3�z���x-[>��C ���(o�0V���T�c8��U�R֑�v��K@��$93H�N��@!��*9<mݠu�c��|�#)��P�1��C���,����M���?>�)�F����n�g��z��o�h��L�pL�\�"���E�K��C |Fw���r*@ �/��p&�c9��$F��~��/n'�78D��Ê��oO}p�܉=Yb�)tg������7���7��
p�SŮ����W�q7��R�nQ�i|yq����ݿv��E�.<D�(�f<82�E�Q�X��o�\�zt���x�G숂/�^0@��xUf�2�����8O��e8S;�熃��<�P��K�7�s30}�����7:�,�-����6�dy��-�~Q�#�ȴZO�X&��o�rZ�v�r�ˊ��X�@��Bm=;2�E5�� ����䫴ۢ���ǵ!��o�(
>�+'�_�7������7�[(OC;!:�'t=��|V�f�h	�V�+�{��^Bܷ.���Օ��OBf���hl�Q��j=�R�9�L���ԁ�n�y\�
IBb�Mwx��{H'se�(�y5u!s�}_�&l������� ��y1��=�=«K��kˀ)5��*
��<�c؏�I�AoI��N�N�?粕�}�-E5;��xۧ)���Q���������r��u��sD�x����~�d��>��A�NW)p����>�'۟~b�2-���c&��������-�(�/wՆJ;����8i�����Lq��󘌙�����Dz�[�J�����V�������05�Q*��N
�
i�~=�f�l�b���c� 1}�Aodn^tWϡ;�o�:�RK��Ϣ�z��y^�E1�Z�gI-�r������	ޥ%xy\���y6eP\̤��R��dF �(]ɏ�Iy����w�Ǒ��b�2���14�D����`բع�5�i:;�rxl�^AEw&�1�ٳc��l�S��ZE�'�{:����z�*t��PE�W k�uI|����"��A���4L�-~�͠��x���~]���$qR��ಖ0Zc+K�_i�i(�7䛈5��Z��`��d�ݡY����Q_�����8����0������j>'"/o�!�ƔEi���K��S'ܼ��5����Y��=_�X>����-?�1�w�}\8�M�uF���R��S��g���P������Y�~V����dY{��*�.!}�?>)�>-��y�ULst�#~�/:��z�U̳�ږ<6Gξ4<o"��k�t������.D��U�!e �zbm;�Ry�e�u&g�m�� �ժ���n|C�M�խ����?��!܇��b�n��q�E�,I*�!�r��k�)	�7�n*�^k��)>k��C���&�y�v��_��whU*�lȆ�m)(���Ma��%ˈ��k�n}'�a�a�|'ȍ9�>��Ĉ��2ڤ@�+���dѻ2h��D�L��g\�}����A�hy(þF����Ud��!�	[Dv��80�^I�Ή�9[�3�͠�;P�ePB��00L~H��AD����:��7ɪ:L?�V�00�/��33æƬ]�ִ������ɠ��v�7��8	K"�u	�b�+<x��k���fB�*�͹��b1� 5�ɞD����u�ZG�|_��䅌hE�3����O.	�􋕭
Xkoß�}�[g�`l/W~�4�-<�,�ӂr&����mFRH��t�rB�z��І/x�v����֏%O�E��d�$���潐^���|���xV'7�<MrB)ڼ���
�l�B":S��n�zB�B
�^&����ntыq����m�0˖�Dx8Yz
D��J�Q��t�N敨AA�1W��M��a�e9�Slf��&�
�"����f��y��B��(ԝ-�/����ds}�y/��,`tכ�h��h���Qq 0���x�|H�M�O(��#ۀ�o�O����3����īRZ��y�p�f���œi݈aUĸ{��ә_-�|�\�d���2��+��*����`iDZ3(N�v�bz�pcrʊ�8��tG #��#�� ��堳J �$��Xt[��w�A���CGV`������xN��m��Be˃Q�Dܓy�j�&�����M�'��(��i[��OL�%+e6���Nt�7Y��\7���;JRZ�,�*:Ի-��T�P�vc�#����tHY��w�w�C$��{o���Q�\��8��'�Ml�c��`h4vf����]}�نe�߉����i�Ogj��`K�"Tߡ��*���f��p�e�Q��ئȧ!��-�:ٴI��gC��!%�.�JY��m�A\Z����,\�w���!V١����%��[�K;x##��i6����O� o�{��@���f��p8�j�]���#���,��;l��Vl�'�L�v%];�#ap�":7uи4��~���L.�u����W����I�����(:�wl�h��>}s���	.�l�'�'�,a���I�F�����y(�m�K�:������V�������z��i�pX�1p;}Ķc�|��:>�.��3L�B,I��wU���b��M����%����c��43�u���o�㗅;�	W/�̑Nsj��C���*g�1ig!��!c�q�غԌ*��;�P�]�#Md;��)_^u\�ۨ��Z���o�*������g���}�eoP�����:~S�;#o�ɸ�8f Ӵ����-�nf�r��,�� y��|Ґ[���#�C����*�A�b8�T�]x��楮(ە/lm���k\�,FJӅ�-��k��,���J#��H��z�&&*���J*[/-�@q���im�=D�)K�5\L�L�Ԛ�f7T:g����"���tI���Lܩ0�PT�od�-wf@�

�e������*��Z��M���%��Ԓ����c���v�����:���5��U0l�\2w�zh�,�Z�4W�۟��-7�呭��co^+C�['̫���(�ی�{���,�?�+Fj��cf�SI@�t�>����uYQa�ɕd�>8H-�Q�-z�i�g+�E�d�0�kWL�W ��������%�Kj��:�TP�5UM��6Fb��V�`��cb
؍JG��zy�����c?Jݍt�@�L:����U��A�0�����7��=�S8�B�D��ܹ��h�7ʐ�� �u��6�ݒf���ޖL��(a��	�!�E������ V�Jw7�p��,&Κ&��r7ɝfR8���2UY��q�28&�L���͒��%&~M��z�E躨����b�o)\ľ��)m�=yH7��e1���X%�֔
�|5wFo��FwT�C��@Ξ�H�Q�	��%���cx���`�B5����T��2b^���a����n'�����+�s�2j`��f�FW��� -�X��{�$�L@��O���{��'Sc�nU�7͈�@�Y�V�4xH̤���E�doQ��bh�r��'J0<rs�Y��Q�4���׌څ/��Y���O�H�$#�o��H�T�H�ת����`k\���ݪ��:B��jV$��M'�^�ܯ����%A�*ߪ�����n��G#�����q��'A ��@ ��A��Ms.�k� A��OIȭG�+���՗W��ނ�|.��sď�< A�0�8�<��p��!�+��q\e��R���!�4gkf�Y���FTarm"	G��f�8v�"�9�K�����k����W�7 Z��qo�����U�cd�\E�;dv��MSB
�WA�%>Ű��&	�gn�� .В<�+��H%I�r�JV�x{0��'71�x��N�A���Z�	�xɿd��Z��c�2�F�z��R���	�����ap�z]����$q�R͖j
�.��J ���� RQ�Ĵ{��h�!`%>���D�� �f�z
&�����PŸS�$�Z�I�I:��3�wpv���"��Ux|-w�e�
z�Đ��&�r�s'�[�do����hkC��470@����n���\�5SD��E=m�Y��kXw2�˃�cH��E���P�.�X��
�gۯ��������h)g7l�wM�P|����ѭ���IN�1뵭�f����6j����>���[�
T+72.�� ;�t�W��ݑ	g�=�q$� L��kc�Δk��J!mF�[��uC.ɿ�[�ߩ=~I�YI������r,��H�p��/�(�<F�����5�G܁L�V��V#�v�v�C�Xk`�Nc�)�WC�m��d5���$+�S�(=�ί@��Ի��E���Iu�zd����7$�.��K� 㩲��J�4(������Dj�@��x?Q���DK�F!%/	���Swp]�+�.bEAK=�(�W�������dJY#�����|h�r��E8ր���Z/�u��M�gFt��kk�{����PvM�$����;<�U"��L?Q>C�p��[�N����Þdl>|�#/C���n�>qyy����(��1�;}W+�̅)J|�v�Ԥ��&����6�'��w�]8�t��S=�_M\�(\f��/I^}f	�zҎ#R5a9XI��Ax�{[�ݺ�i��W8J6��6�8<2����̊��ꍧ��
��Zr'����3�I�����}}�b")SE
Ф.u�)Wf�Q��(f_l�`Gd[¬C��~�����*�Jr�PX^�?N�T�eod	&�׉��R���k6�Y�@�.�,Q)7��U�K���#���!�:�io�]uc�'|q_�z+�H}���Mב�{�gltr�<>��r��2숨�x�Y���Lǻ��"ɜ궬b�FѨ�t�+�Kb��.]B[�p�q�VD���#�/ś�ԂC�|�H�ʼ��L��"t��i�K�3������m@V^ί�� �\�2&�ۋ)��?A�%d�S�E�@�Q�����7#v�s^t�&�=%�Crt;�0�Q͒Ȱ(]�hH�E��6G9���׍�Y.�X�IihE��� ݞ+R��)p�iK�oGY�����Ss2��-	��JK4��+�s�J�8'7�����@
���ev%2p�?_E	�w���p�9
�rS����پ�����}k/-a&ppd�cZ�o�^j�HU�g坝R�������)�J�ejZ��%t�0R �!*���A���0KJ�l�*����Q>���������*����Υe�qU��<�W<i�UΣC�5����b�K���zB����-.!^���5�#L����@U�#0�6�t��&��o����EJor�^�"�)o4�GR�~c��SG�b4S���P�K~�Z�zN_ϭ��=��n�[����L�`O��X��ę�֜{�(-sQO*+
�.��Y*��F�2�R#���avz_C ���U�ǁ��ֹ�Ǧ��|�;p�bln�`h�A�5�S{Z�=:��Kh�k�"����`â�BO�����N�F��Wx�y�]VK�6@�DL�AF�pewi�m �"��L��f]��Lx�^b��#��k�4��i��]��#����{�7Q��gf̂7�;������l;���#�8&��>ˌt�uL�w5�m8�C��]Mc�+�=Ёܰ�N�!}�%��T���u�t�W���9����;ZK= �[9���٥�Ť�rL* 9Z���~_#�C*�ꋒr�r ��"�B_$�K�_�X�7�g���支�)���u�z0�e��GϬʪ�s��s�}������+K����gQ���������404� *O� �l�!uono��!��k4yk��$Q�Һ1�`���u��, �m1MazV�"�X�
��q�D딳ׁ��Yo��@�{d������y�ߨH���F�-3QND�-��+r���TJ��ƕ]uK�/a��L�u�[��x<E��bC}����Xm�ߨ	?,s��M���A��f���V��e̓'Щm�MF�y�?������͠���
 w�n��8S�tm9������j�����g�N�H�~�]SʕU2_&G�h4߰��j��ph��a����8���m�ˀ���~'b����n9��R�1�Uֽ���LQ�H��^nA_�;��i�B�m�����l>���>7�
x�����1d��v7��� ^W�;3���g������� �eu��J�<���u���wI"�8� �_�>�hO'N9ؚ^vJ8���6�9�B��zC�x�Ԕ{�Z���)/�6��;K����B��)���ZS�b�pKo8�]���4��>1ќ#�];�*��2�Nf��=��8JF��F�毡|�z��E/h�~�
�Ʉ�k�m_�cy؊g,��"���ُm�f����ҟ�����a3��6���	��/�#3s,����{�$	���X���Q���k��r�$�K�����F
])�W`Ko+�Gu��ϛ%=A��́��1h+I�f�},�~�b�\�Z�y����.L�&�3C-v�����QpK�"�n��D�\�/f���!+=���U4��IH���(8���+e)��+6]6�U9�D��&�0�M�wf��e��;���L���G�w!FA�#C��|�gς3s�je��)u�ƂkKV( �'�-�_�7{�])c��c�ч���9y�@U��7���(;g� r��TE�����/�B�s����:��[Bm/��
ex%���j�w3�h��%�+i�9��%"�^�=�Qpj^E.�D�k"��ex6��Ey�~��u��9��������Pʒ~�yn�aN(c�t�����xS��s���$���j:r���A��PZo9Z�=P;8	�{X�.B�	N�'Y�8E��/3�f�wq�Ef͈K��<$:�/6�7�����_�Ѣ��Ӑ�xt�,�9x��f"0(}��Y�4c����q��È:�&�&�A�0�:E��r��}T�Kg*��T1�w'���#S��4#��Ҿ�͐,u�b@8�?���^j�/��ġ���Y^c`�>�{�d��,1�0`��}W�۷����l����y��>k�[���eIܧ�}h��n؇|ˏSY�a%&��q���|\n�� ��C��J���.O����"M�?݁�Н&6`Ha�
~x&���O)��,-"7l3�)���|Ұ��:�O��p�D��w5rM,�aKQl=���%j[=io+wl��5�_E.�L�5�c3�G�'�a�sW�հ@!��w����WB�F\pس��hR�V��p���$�WY$Xb�*��hP|:�'��>KV}�����Q+~���,�&�4NK�����%8@����.�(�4{�Cm�B���zJ��-{'���슃$W}���sE���@�����E�w��m>I}�s�T��.2mi�W.0Denw; V���!���o�+@���14g3�J�;d���lp�N��%y�Y	H�OŅʡ�3�d�|:Ӭ�_.����)]4�ŀY�aa���H��x����B?�Ya���Γ>���Y���0ƺ+����o%n'&�a�;���ͤ�6�e�S�g�Z�ƴС��=�Ͳ��($H�� -rz��n�Ҕ�AP��& ;�f�����Z�:�Z)��Q��XQ-0T�|�H������䌆k�QF|����$b�\��M��v�r����[A��{�]Yn��u����Nl���u�#�]`{�l�2�S��)pr�3!�}+*��G����Η�^1/X����2�����ӕ�!;6��}�V��f�#�1��P�A�vėÝ�milw1=8���y���f/At��x8=�b��j5lo�s��, W� �ʂ^�����ƑƣÌuTT�n��z�%h4x�9��3y��+%��E�����t�Ѹ�/����ӿ�S�ҍQ�Td֌������?-S��O�~2��P�t��qL������R�*����M#��2$��{��C�Y���|���hH��nB���H��B��-9��=�:��5�c*6vK{!�%�Kl�~�Zט��*{�A�{�,�$�J蛞���4�Z��{�8�W��/������uђV�ԣ�&��1��N���d�v�O!�H�],}� ���������D,��-a> Q�#�JH���\knD�γsu��E����ԓ�gR��Ń͋�N��d2w�d�QA��$��	�h�<u�����`E��&�� 0X�
}��L�����%��	<B/4�?�3�C��_��j��n���|}Z"'�ԧ�����U���ӱB��,��C���� �cv��P�˘�D�n�&lS)0W)3�E	��p	���s�K����a*���R��H7�!�jj�C�T����6{E��8w�W�@Z�pI�m���}ܼ�jtuŢU1`��M��?3�0�m�TB��9�U��Idr/9z��c�B��'h�(���b_d��� ��#�nk"~*���F�|b!�K����M�~��峲��͖,!GL#��EZ����`��W6���9��a��"��O] Z�&n��wm�P���E&x�
ɨNѹ�p&��<�� cP�A���]������C�z���<r{��&�	j(��Lm�����%�6X��m�5�����M�
g��bh�?(���� EV&�A���"DA���&��ju�9Ħ;0��D�ஒ�#�]�rs�7 ��乛���:�g�s�#봚M�p�ȡ,F�4ׅ~}����ꑱC�ջ�³�*U����+m̍�f����'�����f+���rE���!<,;=�b��v����YvI�����0u0˗ٯ�S����!�������� ��k�2N��Ƴ�7V�p;9"[��0^��|y
������ZL([{����^:�b�/^��
��R�������xZ�oF�8��'d�0���Tr
��N�T$/*iy&�|�gQ�%�d��]�/H��J��w�I��ǲD���O.F�[it�1&jx�_��'��-�;㖎'�0�kQ��CM���i��9�S����>�\���<�\J�Πh���2�3��".��{.��w�?���W����]O4-Ni:_2�i�1^A�9�E/�(v%<��?jb���HLH9����͇p��%������q/���Y@��||L!�v	�&}�J�5��_���	@kS-Q�B�L:r�����C�����Z�Ц����-���c0Ȝu_��@v!�#'�d���2O��2X�d+n�W��l��yDϷ���h��
,�V��f>�|����`�p�D�᰹�'{oϮ��n��P�<�}��j钛x0�Duj�����אj�h��ځ����C@eI�|�'ĵn���q�a���q3�J'{�1�j0AYY6E����� �7�����XC���Ȱ���J�#��N�j�έt�|�)%7�h�i� �,8f���t*�y�[V5(t�!��:e�o�����lg�ٕ`�[�&\+\&	��:��TI�.���O��O�{���-䗜�`;�_U��Z�Amٸ����vV��Z��Q0E1lw77�%5��T	n<hWS@������ܖG�֒A�^��˧w3�^��u����۵��ߑjZ��I��0O�����`��=>�C��i�3НB�W���T������F\��������ϡ.6���I��!$��Q�J#a��:����u�=�,D8ѓ�&
�_vҢ��qN����5��V0�c;&	Ϊr,2�T�i
Z�φ�=��P��`-i�<?�����O[�VB�؉���V��|G��l2��"����t� ��G��5�I�z��|GA��79C�@' 9#~Y�7�簡)�P\�b�u#�<�@�܎}��.��44���xa ������oߪ�69Ż�R�(8T���Lv�rmС�J{74�;�v�>�|�"�AU������+i��,DE��gM�	x�d�y�B؟���g+�{�0��˂��eR�;Y�S��ގ�U��	���Lx�'�O��jۡ�hxӈ�d���B�O��?��+V�zP��A꜃����q��K7�=��X�V����Ҙ�0���\��W/�9�m6<�?4��n{Mt��X���e�}&4�lҲ%��TJ���a[��MՊ�����CC�ĬFUI�N�υ�eu@�}ڼt��>�݁:���`q�ֽ�Y��;��n0�\-� S�C���.	��"Wf+{o��LL�|d-C��&�|�)3�%ue������{�'o�[�n/��U�;ZlY_~i�,}L��bU=���}s�~�\��1-�<�ML?I_�d��O��_X9�A����[� >�2�x	��q1|k\�8X��tSԕ~��'�S�ʇ}�ĥ��Be�|F���C!�qfG1���|�;0l��eB������H�<0S�A��,��OMP�	݌�����&Qx�)�	��>+��p+ݸ��PV`}J�|��=�'z��j�0Yn���<�A�^
��X��*�I�1vy����6%�8�,�q!S)�Dr�2.���h�(�R�hٱ[{ؾe���UDA�����>�N�KR����?�0���7هu."�A���SC|J�r�ͫ,6��.X���.�p?ן�zC�R����@9�dJ��,g���f.�:sm�[�B����S�8���\�h*�>yf��{����oUݍ��J_����A�z�G���=gd`/}�
�DM���T|���n��i�1�kn1��-���- ��u^A�
�.>��s���_�����z�[:nlk���'�
ڪF�X���~�޲��BE����#s5jg=>g���-\� V�OhkS��X7P��y(�d�J�R
�����C[t^th�]���ƻ�R�ӯ9f�lOt1)��@0
��ޢ+N��v�c���%�{H d����I�!��k}��=�,uxʘ١K�>eܩ���)U2dZ��I�[3C�!���g�26-���$�*�`�o�����I���8�YS��b����"���nϢ^*Uy}f�[X)�̪��qL����2/	����5�6�d�٪�(����?��[ǧZ샻H6(��@��6�a��&��V�,�<�B����g��_M��{kz�k�l�
��5����f���OH�u�_VG33����7�R��'�����S4�zu� ���&K<yz�{歭��CVS�0u*��r`�S,���rm�
�Se��?���nw��e��Тa۩��m�~�֘$�s�ƈ,���r�<zc} �°?��kWIҫ�k�����3�x��g)�����f,��3�f�����x^7`�\��P�MD��ˑr��2wM���B��5�n��'TL&�&�5D�'O�f��T֑�s�Nc�\X}:��j�6�.ޠޢj��z��}}����+ד�c����.�!Q	��}	�L�� w���(�mG�2��ʖASg��N����HTfg�u�QŴ�Ev1���ݩ�!+T�/蔳�Q��O��r9�X�]z�Th�D�>c�9�Ѓe�4ĭW�TT��f_P %��/ (ʐ�$�_�Y#�*+3�Ii6�,����Z�CdpUR�`�~z��������АH��L=d�1ݹ��L>�ܩiF�,��uv_&�{[2���G�7P�%l�=�`��<���G����;�I4�Zo��5�u�)����t�R301G���db'��Y��� �}���D0�-#7�_�[w>�����������ҋ>㫑>�ԶZ7{�8G �<-0�&z��Qc` d�0z]���OQ3e�64��JRƘ7S<��5����M8�~d߲�B���Gh�=Z��J���4�%u��|-ؙ#K��*��O��=�ܾ�(`�/����F�J�%i8�t��`-SBo��ϹH@��#�va}����8��!�����������F(����1L�O��gBU�xa���[�̫W�-k���*��:��Ud�*� �Y�ܴ���Q��q�; ��%ty��7�!�b��i�Gc"�h�F��0��=bl��?;�,��N��f���Q����"��p�h������f��
A d7ᵦ*� ̽�6к �a�z�[F���e�;S�^���I�W�,G׉՚������'�]������HF��ݥ���gC�I	W4��-?�����મ��X	����(|NV��B�qf��uc�|�,e�B~[�^��+;c���x�gL."/�3l���U���eEu%h |�σ����������GUˑ�S���e�ޑ��`�Z���z5Ŀ�mcD�S0bi���}��7r ���߽��7]��.'v��;S�˛h,�<p ��<$ki�Ӿ�v8�P���A	�����L-dP$Z��������<C��
]���$����_�D��g�Q�5��z(<�邫X�H�w�s���L/ �|v���­�G`)"i�8����Z���������ЙQkv5v2k34�E�SF}=Dэ���Q���Q5_��?��I�n����#��x��'����e��T7u��۽OE��m[n�
��X������0G����'��):��m_�4i?��������.f�z�^�	罄M�N�a� �V��[QK-^���-�>��˔��@GXxxR�E9���M4/��8�6[�g\���>���i�k�i�N�X��n��|�A���*����>7��o�� �up��d��g������-��%��"�4.�@�>65$��z��/��	d!T]s[�/����z7(a�T���N�	�w��@!�y�.��}w�SC����f܊�,���u��\pׇ曆�_kh�Y��}�h���<��N�~^�ro�_��Yy{�l;����)A��o����s��A���:0��=N3Q�V��+FD��ѻ!^�w���W�2�t]��u|q=��_�[U�0>^wD�����;z_9�C�O��{��\�T���S�`GG/�K��7��������)�8Z�5p��8OY�`��j~Ԛ�����U�ǣ��1-�#K��!���M��&�d�(ԕ<3�fCEUW����?�#�ܼ0MH;H9��T�Sc��G$~�����ܗ8�����_��0M�x��?2�W_"�~����Rr&��{�H��PE���C�9��ex\+U���-��Z5g�"�if��v39C�"m��i�&�'��3y�6Q!6�'�ʎ��:ҧ�6pz&��Lr�j9栉��O�{���^�C�i��à0 �f�ҵI1	@?�-�lW��W9r+T����ש&G�V.8h�pU�:�C��$ڽ7u��v���a6l�^�t�"a�s�R���و�~�Xݒ�(�,q��jl��М��* =�qtJ� ��a�lB�7�\7;VvZi0d����8@�{^]��_��^��eyD��ކ����_�cm�=8^�4�ڄ��=�	NS���˃�U:�!��ת����s!�A���H�aE��[�Ru� ��Ј�v"-
��
^'�>��wN�nb�
���؍܌��[¨m������P����a��*����?B�;��+���,,���6��,G��b�2���:�o���s�Γ_��ζ�cg6}��=�Y�Dc���֏�/[�^�gIUm����r���nm�,�zG�!�cd��`�R�i����Ji�V��	�}�+��=^��(��W�d�D�~F|�����Q��ќ���#�M��X�t�8����t��\9���8�)���H+�T���A��a��c�����fH��=*��i3�' ˊ�C��d3�l�uX��R*�W�+#�րJN	�7�#':Q�19�l'q����� ��,�X�0�uӰ�F����#y4�V�n��i��*�Y�b3�~���Ϥ(���"~��o�!r0�@�GS�eo��5��F��L,�7���"�Q����{�[���p&"�2��9}�g�l� ��5��x.��+s��_���A����1��K}1���c2+JgJ����N}};!2GRcFFbu��
���ֿ��T��	 T��{.f�k'�^�g��
�n)tL�taNDKO"�%�.�_�s ����Y(�'�(��`ߝa*���p&��s�2!""|W���r�^��d�
�1���S����ve1/�n X��j�֮����o�,.��z��S�����F�Y�R��,O
A�5��'1���U'�z4Tb6�$�P�w�t_�#8�@ܭ��8m��x��(�l���Kq�!�Og��]�� �k7�MM�\?�J�<�1�F�p�?���+4=�Òm?��`(O-�������,pE`G�;Y쭴Ҭ��Ayb�-~�(��K�A`�'���;C�d33A/�F�?3t1�塠��&ׯ�:X3l�MϞ�ς�䆶|���"b�6���%M0/F���dT�ay��?���y���t=+��G"��]ڠӢ(�(vQ��y"�a�{��^/�H<�#p�`�2�\�/��P�������%Ͼ_������MZ��r?<���)�vԳ4J�d�7}��x�Ϋ..�+���{�H�a��PP��J�	��x�V�W#��)�7J� +
�o*��E%S�����-��Ş���-pH�QW�_�:���#���>FK�߂�_Y���RI9�����";�lfP�՜ӿ�܈k�D)M��Wm�n�Z�rk|Ƽ:�챤{�u�7�]��'@��
qB�����J�0C~|N���H�K�u�ޝ��U2����>���o���F{���.#����yu����+5��d��>0�b�wX��-�����h�v(K�-�V�l��G):�{tBH��D�ʨ�<F�<�z�P+J�|P�e9Xi�9�*��Y����P���tT.���P�-���N�BӴ�՗g�LO~Ģ��Po
�$M���J*�~��˜�K�8�qt�%���=\d\ޠV��-J�s+*D�����2�;�\��sF���(N7�� �\ 1<�)I"I�bP��
����u�;�]d��{���4�Q1`���H���,	�m�2FO\爟V����qj�С^^}!"w�b,m�Q��෕q���J#�H��7��Q+G>^qU�&��D�CS�f���!�pHpٷP+[9��~��@�>�GȄ7wW��D�S����j<��<.�ƕ���i�ѕ�}�+�H���B���6b���L�n�b�������`�/���=���r���0�&����ܥ2���ST�r�f2瑇�)�L��/�Gܐ���(��iV�}�X�,���,"D��9�M���w���pS�ʅS����L^{�N�����R��� ��t�ɮGu���~jJp��#f��7G�>@��Xc�3w�pm�Lim�jz�jm��y�G�\��<�7��fܚ7r���ʅo=�������Z���ȶS���&�F�� �%1�k+�솴/��������Oq���@K0�Z�m�[} � �s�Xt�;Z-+�K'���� �=����da�\�����,�S0�a#�1�;C"+�zq��R�O� �6
A�.DyD	B2��tw��:
9����<��L@�؈4���ݳ�4p��y|��\'��%��p{g[���ό���h�y��r����4�b02�)�`]���`@�Vy ����a5���e��ax�(�B4��=��ێm�S.<�
6�ƥÈ��сy���P$-S�o��rM���c�]�D�D�`-h/�Bv�dQ�-8��￯��S2��[0z���֨��I������<��	����J�a�u�>B�J:������I�˄ nO0��lU���v^�4_�k(ƲM��٤�L������'�j�z�u5-3>HN5��=^/���Y��N�Sk"傇 �6'�H^�Ͽ��0������ɂ���8r���+��NO�Qޅe,'o��WdCt���s!����:�ޮ�o��/�3-ǝb+�~0No'���3�qy�:�z:�t�J���(��;�M��VN��.o|ۖ�e�.�fF���i���ިj�`�i؆ָ��M�j��$,*OG\\N΀l�|ߢ����p#X2�@�a�;*���]I�O
�i�K�9Myk�6�G��I)�F������Zu�����垧�`��%?��כY�}^�B1oA��I�����!����#�ل��+cUm�U��//�l��z�ϣ�(C�����Ru��?�����ߣ�챰��&3��<F6��V4��V���q*LQ�U�炝u�{A~�عJ�t#��d�<g_��[�M�����PY^���L�Ff�Ty*��O �s�B��X���q�S2TT���9���v2���Ja�W��Z�Qk���8�R��ulh��<*��<6�~r񫧽.?,0�����{�f	�D[��G�8{�D�t�{�ߒ�� ����-7��~���LK�)��`��v���WG���i7'o�ͳ�h�����bz����~��S--`1l��SBq1�7&�Q�M���ॻ�@�
1Y��G�w��r��|$"-��Nm(�N<c��;�q�ϫ�q�F�ǒ��N���S~�߄<@��V�6[ݽo}�xr�#�g4�n�.>s����'B�Nt��ف]_�
��>T��2�n�x��G׌�޲r�����y]���v��nN#�e��/�fb��N��.��L`�n0�݃��G��GLw�c��Ѥ����P�!�̮�p>�҄�����B��?^qTc�{��L�^7���lM���݆�R�'~��7���ӹ��Ԩ��K��O���a�!���:!W�����q���-�c�?�}��l<�y�%��LX12J�BY� Գ�/� [}Q�>����"��f6�P�4��D6������֑1M��"�C ��1��"��D8rE�a ln/�G�Yם/�<��P�����2��t���5eX6�\��H/ �f3�;�i�3F�	����,=h�(�!��+zyc'��߽��H�+Hc�x0�s�Hweê��%�
#)!;1�*�"��b�Z��B����9�D	z�7��M�#��n�c���A��nU+�ɿ����sW����b͠a�F_c/ rPA&����2�~��y6BKy��)~L�"W�_��\��</_�.O�A9�Fݬ.�s�e�9ᄊ}Y­V?�W�ތ38G��<�"��@w�]^���h�V�Ғ?�u�$:��4��e�_~]_��(�2J࠹����E�&/�W�2^x��$�g8#z9}p�dn��C^�9��XF��f�8)l�U{�1
�w�����RU�r� ��F���fGo�U�*gi����ۅ�7��"���U\�҄�9~��"襘ŝuUM���L#����s��\�<�ݐg��l�vmR���I�ҩ�%[۠�=��w�	�10mu����R��>��yUkq����q��:��0��8�����Ȱ��&�,�p����e��~�"O�%	f!�y���M�PR��ݐ�����n嚅!¦��9��׎C��ϐ$g����'�^�o�.D��8R�[�kE���Htu$�9@@���r~QM��L�FV"�
�,���`�A���'��z�[�uޚi�ѱ����a��.��;>g���`�"�;��>�m\<t ���L�����9Zt}���:�V�l��:��M����s��Aݺm}�0�굚��C�:T^����>�j���y>�\s��D>����sR�?ߣ~��A�(~�:��VԈ�*h/��r�$Ω�܍���7�g/+Z�l�9�[�+����r-�6�n0Q�^�׻'AM����L�G4����O���	|��Y[��=D�Bu�yo�]��C	�*n�:�k|ȬK[����d�G��d(�����Wǥy�b���V鮒w�Mb? 'C�Ta�n�ش^/W7gI�S$G��lM���.e(Y)u(�-F��b�^�t1)��#���r��{��ll���R���'K��P��F�����dGT�OR�;8�ly/�|�6��s�Ϳ�i ��͹,e{�z�:�6���f���NQa�t!�����4�wʐ�xsK�[֥�f�"�~�G�vD������)�#��X�Ͳ���[���+���6�D��?�>̄U&G1�yA�D�W'xo���X����<����4ߏ7=���B"QM���s�#�!1��.1��Y��m6,��􍤽U���Zyu&n���ё��&�3�M��SA�n���qp]�;ﲙ�Bp�{��!�4c�U�'�w*�@Y�G�P(��'�<l�d1�!�x0��RǛ}dn�4�F�[4#j6Z����QS�Csz�׽ӄH��'m�nn���u�{M�U��ӈ[T��F�P�IH�C�yz*����x
�yL�E+�F��b���*sn
�vX7V��j7��"j\��Z���!�˴�h`_�a&��9H���5Rg.�N)93�񔲿�+3�\8ߴ�ߩ���X}|�i,��.m᪤�&�1~N��e_��T��2t��/���W��rHÅ$P݉~��x���$��M���5��4p�v�D��b�!�;�+��v�.�����ǂ�Ӹ��NƯ�c�ߥ�3F�Z}��?��=6�B4C���ܶ��+�Il&&?���:���W���T=a����O�3rB�Uz!�����Ŕ�ދ�[�e8-�3�sA��?��1I%��"�EOC��+�L7VX��qT�[�hȋ�g?����ӃW��c����}}S�r	�6�ZY�_�@��g�@-o��r��,�Y��xh����q��z���'�!>8�i���g��dY+�K�"�HI3��n�1Kz�1ҰkU<>|<z��A����(�_�f@�#tYl��zR�y�\�)�]Q��f�ze�Is���d���u�)*���H	C�z�;�q0�?2O��n�!��
��G,�r�ܿ4�s��6W�>������}�#����gŔz�А�@t���-n��a2]q�L�s�Iɕ�I�������H7B���C4s`���%U�+"�Zf�En&�%ܔ�!�p����K Y&�Z6h�k����6R&����2�Cm�>�� �M�~;��ъc(�2Kx��6B[~�����R��n��@61�$#�^VdF^y��.Ա�,�����YT}k�y���i�W�m�h�<<0�;�cY3�0xu�-���0�+�BQ�eY����;��I�{�:>�gD��'?�s���� �O��x��f�-���ط��q��E�sD��`�����鰟xo(��Y^�_0�:~@B��3v9��)T4d�0֞�$�>�{*�����O�gS̈c\X��sۀZ���3"ȱL�j���m�������r}ģ@r
��ZZ�Lm���K��C����ݘ �.�z��)�n^��R���#��>ޮ��t*z��v�=#K�"� ��������l��ҷ��ɀ�uO�b��mMل��5N���[�j�S�͊e�ӧ��$^���X��KT�~�|:99����ٻ��T� I���_��و�GhL�U����A7RJ�Īj���m�����Tǂ�-*�$��ny$�Q��_Py((�����[��GB�P�֊���sE�an��W!d�I�t-犂���ָݓH�9%7����KQt{a����.�VN��,��º�"G=�с�����[���zmf�M���b�'@�1�B��I���z�/L�D��ޓ����4Q)��_�����pv�H�*|X�6��g?��>��5��tY�/��*�͡���D�1��"CN��.˱d`6J�A]����.�e��0��:������}L��h.�P��xu��$Up��8�ީ����Ok�#�	}e�n�(E��l��ߙ�s�ϺF2��t���ݘ�o�<�G,�8��(� p�{5J�Ob[�-�:��t>��ę�/����c��ro^�jS�A�~|Ȕ�#�3�Yg�V_��5���~l��&r�6!j��7ry�;{pP�{���
vn�~V��y(��rnh�ϡ�P�hn��^�77�W�"�e h8���D�����1�*�C��S]�z1�<����~ҟ=m�㰷W�>?����)�K=q���pCY���$�%=�F�!m�����]mUm"���>m�4NJ��e�_���h��$uA��m~�+"J�������T����tuw���̛ɘ�y�*�\gEhe.1b�����℻L%��$(ip ��?��x����@��F,%���G0�����bݞ�+).��̈h$f؅����`��P�w�E}O�X5��0R]5�ď��e�+�p{n��"���Q�su�ldfg�hK�
�w�{�s��۱3�����E��Ix݈�h`�5��u	9Q�Tzw~��kμj~`�5��
��ˈ�]��� �)t�����ӹ+,:���U�S����L�K�E�����c9^dڻ��9���DT���T�/(��*1���~l<��55d�m�(�ӽ�~71��c�朗�����F�HˡR�	Kd}��-�3}�y��##%$���}nt�z4�y���%�M'����X���V��&���T��g�/���/%bK�1�)��-D�\L�́*$a�m^f
$Z����0��Ҩ&X�OV~���e̔�T`lF��eU��.���.B�Jq�%c��ҹu��8+kJe������}C�& �:��s��+z�Scz�,�w��Ш���U�BE�,|#�� ���t]��*����Ӈ��1׺����wD��g�qF�	�X �b���G�MX��o������[#��`�-�u�{�������weˡ[�d��'����ZY���q@�5��U�Ѭ��K^�s�Z�`�
!{�*��D��j�w������Q��V��f�����țqP�� ��,��UB����ތh�A�\I���Ѯ�x�!�櫁$��D��;�-W�_r��h�4K���# ��pU����N����.ΡH��hBGR����CQ�"x�:�8��]X��_U�C�P�"����>��Xф�	���򮔊����I�����2�� ~����U�F.C�Hq�m��{���#j\Y���!�	)ƑoS#?6�P�`��`-���c�u ҍ�e���@QR��w��)�8���"\1vL%'+6�&b��4l�*�E����=Vb��|�����Gr<U����2��-��0P���ZQz���z#���Q����Uq��} R,��B�Q��`�vL�m��q ��G���ف��B���wԯ�թr#~Ⴏ���"��?瘬?$ViMed������t��>�3�z��>[����]�qo��^\�3L�%�Fׇj5ԁ�ڨ;�]MƯ��E 	��1ʀG�$�w�z]�0i`x���My��m�=��7�Lw��xVCL���J3�R�����6��@�w,��)��WP�^�}��g���V�|�Gb�@;�|r����I,>_)+��B����n��E�ڽ�#O�QF#��M\�W�Ha���8�y��,��ZOM~��B�{��.2��?^��r%Ձ�"wM�A�g�Fn6<��2��g98rν�8B�ت���|l8����Ò�(L�����&��!;,�h��S�J,�p��ˣ��lU���hC��� *�k��$
o���ygw��]mz�v�6����p
����w����B'j�*�"���w=?�=���Ա`��$O�Q�.^�	��(�~��ٽH��f����Udav�vo���t�(*g���Vn��xv�i�:Xdoҟ�4�v�}o#��%K���4z���~$��$H�3 u�p���zF�0�ᥴqTR�1n5�p��#��ެ�4��x����yo%�6��v�ƽ����̒��F����+�c-�h�\ʱ�Kp-i�J�=[���	��J��+zy��U~�����sz�oLñ5�J��ER����N܃)�r��4�`F+��/�kf>�A�%�d�|.KVN��XA�>��=���?�M_7az_���r���u�������F
����u�B���of�g	p�Y9�?�����m�ql%OIܺ�m���*jMw�Ne��׃'��+GW���l�zc��]��4/��S�%QR�	��8[���x&)H��_�p�.#�9��l9<���(�w�������<LE�V��|��O	J6[�<y���*C���; P|�N1��({<�τ�
��t�m�*Y�$|��ע�&���J*��sD����+��Sr�G�?�����L�7:�=������t_N9��p��cjh.)I#A=�����FKP�k�Ւ���L�.�Q���G�n�Y�မd�����PFJ7��ē�%���$�-���R��v���Hn����c����3���Cpe7�N`P@���Y��E��<���a �"�|�}(>Տ=]��!�k��%��j�	¨�ɒ �/�N����3I�~]��Wm��&��(����C�rc5MHk�s�qd��Twg����oq޴�y޾g]"�F���=���˫�$h%;��ݕ
���-k��tw@r���w������2�#�9[/Hɀ$�>, �ڔ���WB��h��(��%��/�̛οO�D����W
O>��;��]z$�N��Q���I��(`_�
g����_+`�����ǔV.?�)�RUM��1V&o�g��2��[_����Eۼ.�i\GN��&K[��H��.�u�8��X��ٯw�K4�^�gq�TPNŖ,d��U��o�/�)�V��ܡk��dJ����r�ڪ/���.'���5�u��kQSaƶ1�b]��nJsn5�{�ˉ�`�R"3;�F%�PO>�ݑ%�fPd���i�
W����n@8?5XGgթS�,}��XG:������Z�Ԧ	I�t*��E��
}D-��A����nS�X�[�
^��c�Ѿ%����ˢp޸��S�\Q������QO ��"|g�⪀�_T��#%��i>��<e�;�;�����ZϓB~}qnB����`pb�ׂ+�����*)��f�S�w�c���z�Κ]h�*3��I.�z��O~�1�EA��w��f*��9*�'��T�*��on��[�Od�~{2/�t��������Y�}�������J#���=\��s_� �E� ����[�ҏ���-@�
.�����;%������6��[8�E]���!�X-���6�LLs)�^(�#7Cǥd��R�������B�INV-,��Ө�P[8I�vu�Z��ծRe%�k�4B#��tn�%�� �q9 N��ߖcTBR�]G�>�~��@�V���=h��1"D�/	�K�u��5=VN`gܬ��\��/��f��&��
����W"C��N	�����w)~��l�>N���jڧ��㲈���{�b�ר�n;��0p��C�U7��9��Z�̋��x��i�&4�%��=���R_g�����u��0���P�{EM�вv2�T��U���or/Jx�u��jv��O[���|��{��H�QUN����� ��.�,ɳ�.; �g��W��]@��׆�J�
mS(�0�G��|�_V-���l�Tg"�'b����/6����$R�Wrm��Ӛ�y�wf��\�=�����S9�b�������m��,P�o���e��m\�|�!�����RU!��x��l�ƈ��
k�b!Se�#Ձ���`a�@H�Ğ�v[	y���|_����4kw���B��Ak@��<���7n6�A��c>6b��#�w�?i������sQjB���th���6C��ʬ��\��y�<|m	²��fܪ�Jh)��,c�Xb���S�$���+�s���6ܭX���葝Sތ.7u�Uؾ�ͼT�����	'�y+v;,|>Д�rU �|\����Ԡ��Q�9�� L�-�z8��E��U�x���o�Á�4�|�^�+�G�`y쌤���g���� L��o��\�D�#�e�jɢ"�ܓ\4���;��i�Z{�t�0W-����\t=x�G���GGR�M�@�jl��I�nVEBh��y�]��p��_�;edM��*��r��-��(CAq��l6�G�3�
<��F���ȝ�bD���um=P$wJ�����]���f\�ԍ���k@W���I��-���o�~���v��Z�3O�vl����S�A#��� ����wcv]�y��[C��)zd���g}�^٦�E^	5�����������n�4�y�Xw$ҏ��!���:�Ԏ�A�T�_˟����r����%�-bI�����6C}�q�1]�=hQ磉��m�o�������qP�>��U�,��Cw�*��B����"�u3]i���ϣ%8�L���[��R1�S���	�χkM�q�� �"�p��rR���j�)�>}P���@Y9I�؄q��m&���H�����a@s7����vuS����K�ʖ�vVg>�C���>#F����_�t���"#��d��J$o��<fp����*8LJ����r;�, i��0�עEre�P���c�&P�"k����ȶCu��3I8���`���sز�C�j����I��k��V�Rc�Bn���D'�����;�˻2��l*�n%&r5�^�)�l��\��Et�O�7{�ϵ���|ok2���j��Y1ȹUk�P�b.���:������p�o�ڙ���3C&��9��G42�����	Z��z���<n�&|��
�$�j�vQ��-y_�嬈0��h���Q�0�J��}�vy0�齄�t}"�HJ�ze�cOH	�Rl_L��$�-���%��^~r�Gt
Eߝ��� e�
�+r�#D��?U�*�Dxn�d-�֬�4�ř�0k
��7o>��kh�dzu���Ɖq9���:3rغ��j��/nz�F١Y�Ô������un.۟)�c�4o�7Іx�.��/S\�'<�q�/���v,�έF�:"�I/��Z�j��$��uC����Z2�bҴIAzC�i���tA<W�r:��ٱbx}*�yzg@&��3f�����i���=�8��=X�)l��P�&\�@��4�nc�D�ўΥ�a���E��@�r�e�����6R����7�Ϧ�n�B�����e^2s���3�R�! *Y��M�����YЏ�_{��ޙ�8f���� ^RFnڿL�7���f*�!!-9�ǖ��@T���5}���4H��2+�ٟR�/�r{M�6�m�q0��~�p�SنE�fN���1����
�BfX�81ʕ�}Zq#��}lF�� .���V�4��H�0�/�-�ōC,9'Ri��4��D=�!�������E.m�����|>�;D����5��
x���G����#)P��u��ݐ#K%��:�������q��YTH�m�DzQ���
Q���|��˽�n3��1�TрS����q0�T��h7���$&C���� �_8Y|��ɲe��B�O5����k�n�*��W���C�* ��O9�W����������m��B���f��N��a�bP̎�x|x��yF�7���"VAnu�}�����F�8�F���w��z�h̹ӱ����*U��04��Z���V����<	��ڨ �V܆R���r�z޶�*/�e����=$�*Y��ɲ�
N�Q�-Vwc��N��Y۔7�&X�H�d׊oє
��7�Y�p�LqJv�����ǿM!�"�<	�M�g
��[B�ER)�^YΝm�O��?�W4��j��yR/�ˢ}���vX�<@�t�6!x��{u�k��`:;�EV�l�yJN~��(���_�㍹>L���K��rŊ�~ԩx�� (���
������*:iE&��YW�+����U�0��6$�@͎�	�˶�8��	�෾��d���"�����%�; x��7�+M�m��:\]`���p-1mK�	�
%׀(׺9Y�^�x�~�����n}�xcGnѴrԎV6�PĖ*a��p{9R�]m�X3����5ш #˜���n�I�҉��n%����)U-c�6�}h�>�lAGq���h�^"���3���y��f��H'2�w��
"�E�V~?�.$�o%;�'	(LG��U��������Y�ؑ��
T@<��]؈��L��w�'�|rT(�\'�%�e]u������-sq	c}u�z���wh��jx��Mګ�ML�����p#�t4d ��nP����/��&�Fﶰ��oȮ�-Ĕ��p��'����T��;�*�i�ȫ��<�.)���a�
���r����u���,8����R)7��sȼ�����C���hw~<`1_PS���ow�@P�K���8�9�i�)*!k0�5��؎�'���#EI$s(�d�<p�|��]T��C��}���ƃyA�5F���S��}��5�j��T�s5v#1JE�=�؂�ښAc_���W㺶�p�Ҷ�9:Ӵ��i9��T��d��(ԓؼ�����LkW��.��r{Ȭ���_��b���D��#�?#q��F@������S��[��B�]/u���u�V�'Zi������7��ǒF�b�^��Шc|���l
c�3���Oz�A�=����BMM�Zz@$��P>�C|ErZ�:������h�=���8����S��{�f�;Y�8��J�gC��#�]$a��o�Q�g���3����}�ѣ�09���-k�F�y��YU���/?�hay�5��3����L��E��/�~��T2Y=���r꘷\��_uz���sbb~�J��W�~&��}���ڹ����hGP��J����g�����hQ��X��8=8�'�Z]s���="�`��>��k}o�TK*FO�#^!�z�}�����G�G�!�/Ŗ�p����ύ����5A^0��Sm�0	  ��I��vruw�YP���*#s�ɇ�e�����>���LġG��	C�G�*���1y���9���n�W��cց���]ErR��]$��}Aճm���*�}��϶���!�&s'��S�0TweJ�A���vd+ʫw啻p1rp�h)A=��H�7	0��������1=k��V���r����B�F����ؤH�*6�M���9��~
�Ӹq�|E�����N��M�n��Q��kv��lƾ>=���G��D��V��Ɨ��+`��ur���[͐K���e�ό̘e-*p�tcm��L�䩤�e����1�h��	��L4Ԧ�9������\��֡�y?R������7����w�}�"Ȭ����*M�M�����^LX�U,+ڈiO�yI-�(b0���J��bZOeQ�w���}7LwB��L84���i94Qj,�9c����FFM��O\8s����f����)�,n����,����!ڝ��
0m���ah�9�T�J�b��v�ιAZ/�O��.D$��׬!.4�v4���#QQ�:uhm
�4��G��P
j�a�Y�9m~����������'#?����	�m9���P6�D��-�rk,>b��o��m�$�Fȅ�+��g����`��d���B���5��N[�h~�����볓Y��X����>�"��K�˄�N8��
����JN�D�@�������}_�	>�����q0�X����_���`/Vm,i�'|�E;dák5bb'1A]y1+��jrr�s5��Pn7�.P��3N�3�"���nM��*E�a3�~ȫ��.���"�)�	C�-P7�[�R������*_��Z�d_:01P�����)���ǯ_����n��o����v?�	�c�˒���BQ	{9��A����^���>q�,�������Վ��EAQ������yO��{�/�(52ؽL9L��!f���U��M�-#>l}��c��m'	,Y(\���rM��5�	(��xu�EI<����G��,.ɠu
�_Y���v�4��c��x9�C�~y�����u�-JHY*O(��:P8�sѴ�J$��kzb=j�7���T�v���g���s�d�wy���!�[J62��1�C���%Ʋ���u4~�dٸ)�a�K_�ێ<��X&+|�^�R����SС��j�x���jk^�^��Ǎ��ę6g�a����qG�
y���; �٦��s('�ǣV�V7����SY��b���SA����;���,��Q�>U&?�1%o0�IR��V�r\��T�]{�$ ��u��2E�dL�=q�B^æ�C�&)5�n�-�����u��ƶ2Qv��\�**����Q��}Y2j\��5^.�=��Tz
���R��*���Y�k�����Wt��g�1Ԫ�k����5�a~[�������f�[x?|�Co��Ы��l���mW槢�d�dNbu�4Iv�Ұ=�O]����H_�R����-ӥ�3�#v.���O�·|�����X1�GsR��4)�l��۶ωɻ��\L+���^`�Ե�F?"�Ͷ����0���ϘǸ�Bp��"�{2� �n#D�"����a�.���"F5*#%��oщ����}���4�q,Ԫ��%N�*��b�,\���y��?^���96���:��X0#7�t�X՗���6o��9;&�Z-�R�>;5��ז����59���;����UTV­Fi��Ɔ�>+@�������J��=_3�U"�@�g3u����e��q�ꇜ ���b�X�RC������6fG��C{&>#�o��0�`�B�hƉ��	�̹9-[k�z�X�[�x������l�
��fW��3��^�����?��+�s��u	<�]�SE�:��4oJa^��3�i������<���w,
hG����������֭���0HibD�-R ���̤�%�)����6��`Q�c��.��}��W~'J�5���q�!��n�Z�#[*�@n�:�_��>���(��z����D��C�H���k&�)�h���p���*I9ǋ��h�Vr�\1N$]������ć)ǫF�ڼ��X�ҩ�U�� '܉#KO{�ks�5�;w�_�o�j�{6�M�3�8�!�ED�Y^V y��j�_�q���F��t%���t�n&�,6!�7��*�~�(;�:�1�p����A��yѱ6�����j�o�xݧ�t��)"�W`^�6m����헰K
O��>[<�=9�S�@E�O+��ackn���UVm>�b*k�=;��C�cu�1����s��[}i�7���Өd�H#P �"H��=���Ffi,`ƭ��@�<Z�����:��Q��;眂�3&kt�"�.��ȱ���h�:����RʈX�U9Y<OU9䊆���ѕ���z6|Uc^�p�Xg�(~��Vl��z%��s�
��K�d��_��,���-�,��%��LMN��u[���}���9��u��Ucޙ������I�����)]-tޖ(��r/eH�4�q7��F�*9��r��$8K�J����졣�3��ژ���Q�$�(�Fi
"�s�1��(L]a�n���\r��d #��.80'}�JIM��_���@{����\���.u3���c٤ D+I�`XR��Yl$��D*L2G�%J�E�%�I���l�N���+�s�#���7�؅�������0�P#B}�^��<�o]q��،g���΢�iJh�����		Y��+P-���q���+�F+����8�{��cX�Sf)�{pS	?_^L�����X��l.d��~d��|aT�D�'V��q�;���J�Y7b5��S��n��o���]�uw
|��l\�#���o=\\�w88hPP�O��Ue��c�_�����l�� ����waO�XB�E�E�!\V�������Q�vw[�AP[�6�&a��~�������}�#�#�)�.T&�"��[[Ϡ!��g�O}v@{�_�6up��~}n��-�֌H�n>DR p��2��û�z�gv4��p;�y�n�����Y:C֣�^�\m�|���E}�烼q�YY������w�Y@2���|3�J翗�(ʼ�OQ �k��\W�5%�x�{6��u&j���{�>���ɫ�Y�������L���u�jQ)��'��o��㚘�`Y��@��������a���"�B�s����Z.����,mRa�G����m% ���(m�K	���mU��/�U>ivȚG���qt��@%������r�6����#,�)[=�_�3�|�%i���w��
M|x5g����k��/���U���Ʃ3�((rM���F���<�q|P�bAЭ:`��a�q�6m)����C�W��EH�|&�u��$�YT���hꂮ�^h�|���Aa|iOX��q�\�1�/\���j4冐�;���8���}�D��3	@���q�����ͫ��e�P���+�'�"Mf�q2��:�Fa�uD̑�#�FK/���8���.f��/;K�a{�y�⸕�P�4��g�62
��(�����[Zc�u��š�@�
Z�[���,1�ǹ8�) 9��݌�B|�XR�[|��gA�%BӞ��Y�S�@Dɾ��~�,�hr��XT��7U���E*<�z����)����6�[�_#��jo�a�M���v����"���vX�'~:�w����Ԟ�12	��V�$�������t0;���eO�wPn�&ap���P4ν({�����nK�D������IJ��T؊΀��?꿡3b��]F�-*]�~i�AA��LO�^�]����$�ĵ�Ud��*=�)M�|%�R�v{5g�O`(�Q��N�7.?ȓ��	Dh0�:u7/���ؠ�3�̀"JAj[�(�Q#�� �(�4��[]J��eT�0��gM������8�鵷�����{4ݫ	��w�H�]֧�t�=D����<]x *��
V���;���K�q�Y��0�)p�L��s?9��5^(��� ���ݰ<�~�s��6�=b�ŵ���I�����굢 w�DG(��Z��$:�?j��CmD�s�=�_&Y̇M��� ��k��@,GQUB������mp���K���	J,��'�ϱ���8��A�GvS6�Dtퟲ�zդ0����p���0��jEr��X\r���������lu�m����fe�8	��+j�':��%�x.�,`)f���!9s_Qr��-�=��)��r���=F��.��?yFz���$�|59ѧ�r���(㡋QZ�5��C,9w��⦳�F,�a&�[��Os;O�γ&:�	��+m��-�a���g����?AS��*��D�N�5���y�;}�Z�tQ����̛ 	��~�F�u����ռF�K�)�l(�	��|��|��s�2J.����)z@��޵�1�"�ċ~ң�񢕹�*�-b,6�)_���待4���|��^_s��kt���|�H_0?�c�״^�_M�lğ<�V�#�!�i���;��~���{SPǕ+0\�����ت�a�3�t��Tњ3e&� 8s�H�l�y�@��{�4Ơ�F_=P|�O@k�d蠟W�ί�6���[�jk݉G=��o����s���ν�`���d���WI$�~1E�'=y���v����Y�&�|�#cJj�
,l��Fx���l�X�f���"��f�B�i���f��:,;1���8��byu䡺�o{(�7��%�[G?^?nHi,���9iL�,�82�ׄL��+����d�Ba�="���d'�� 2���ZI�窜�A�P�+HG�.ʹ"�~�d4`G�� �����(��A��GTl�����}�} rτ|R��Я;�D�8  �J�'���/@7�`�
����)WO�����ki�0�&��T�k�AYl��������,�!�]T���܍����y"ǙY���"��f��]�����B���&-ω����	���)���^��S�8��.�:��}|]B�I����KD�֒.��3�a��x ��l5�R�n֎Z� C �͉��R��c�4� ��Gq�(���V^Q@�G�*"�Aճ���s��c��wju6Bj��:~<��=�c�{�5O��@~@&ACCP��ܘ�ۅ]�v]BD�YjY�&���G��T#B�F�2����r�s[r�B�\4����X��U2�N��֨���4���x^I��R��|ŬJ	Y�����A
�kg��o��m$�Y	]8#�%��wZ�x�R�Ź����b�S3���J=�� U���_����<@��5d�Ow@�m�v�jʯ>̾�,�6�P� ��>q�D�&���e��Ck�eEAi���-ʇʱvW��w�
������.:*���� '�q׺$��/�?/HY��0�����f��`�kxqo�i+
�`\pH	9��S9��д̅(ϜʂJ�������t`:�;�DZ���6�T�\����4?
q|�* H�J�Q!���ds2��^��|���f5��������{o��A�*����OϢ�ğs�k�A��x���V�RJ���}����Tj.��[�B�!4Xٶ-FL�����[�v�������I�Jص
�R�LO�_{�/[�A�/bz�I3-�2��J�&څ�M��C%��s8.��4���%H2��\�#���:A��N��1��d�����}�N�0��A��p�O�aF�_��]K�P���s���8J�z%�ٕ/��\*����|fc���-'3	:�f�l��y����{�$N� �\�=*B_���.�2��̼��mu�?.ۺq�S��F��o&��6�]��$g�fR�.�*v�جU�r\<@t�ﾷLL������Zq��'��ɤd�>U�`((k�	2��y�n�(u�`��̍+�Z�� ��0��<�F��1&[�x?��+&2H�x~���U�`9/KT�������ak⯱���2PT-ݹ�ح��6�d5�](~0 ���0>E��t�coK�tES�w�`���!.��X�v&bвGCT➅���L���z]�t���]��\����E���g��EK��.��[�����=�g�Oqy�m��ubh�0�x7��N2��k.�<ޯ3Þl'Ș�����P<[�> ��@ ������󥭵�P�QX�T�\�rW,s� <r,P�_���� �[���  ��)��+U�*3҄���R�ƊЍ��Z����t��t� 3ɵ�V3��f$�0�]��sK��r��r)<�	r�P��+E� �f ��`��]s���]s�]<�r�PS��V�V[��f<�r�
P�]�]�]��V�VjYPH;�r�����@���|  �V<��r_3����HC�C������|  v.��3��U �m��+U�;Ur�U@U�V����؍U3�S@Q���ڑ�V3�Y�����[�CY�]V��+��^���;~,s�f(X�N0_��G<s��< u� �F+ǫ��^4�v8F�������V��S�����u�8t��yF3�f�PU����P�ER���"�U ��+U;�Zv�E3��+���E)E���)�X��} u�E �e�e��3�@����;�r�+�ñ��R�s��	s���P���V[�� �@ �@ �p@ �@                              �`                     